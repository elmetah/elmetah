MPQ    ��    h�  h                                                                                 �A=�	��Ez�+a	���?�'%�d���\�G�����gV[:��ب�l�ݰ��#T���&��YԔGu|R1Ҫ@����E�lύ`��l��+qԐ�Z9-�V��h��W9�8=��Jɚ����]�TæW>0�3&[C��ȓ@���
<�ic�ђ�i(Ox��$�c��]M�i8�Rs��T#e���Y����(a���k���n0٢7#w��"1"Ƀ]Zg&��'r�<�g����vc��8��6���ށ�´��D2����xV��i.!R�+��?R���W}���b?�]��.? 4�f�����'�p�n:`q���FNC��LQ瀣��Q�pj�2�Ի,+H��u�Qq8^�� �B�@��o�4��e��T�D��aA	��B%�Y��z�>�jכ�eQٖ���z��>�\*�J��R��A Y�3��u�C�� �~�ej�6��>ԋke���(?��K	�i�,;惮ZYzᗍ���c㌗�4�"�Z�_����ת�I�"Lw@�E�٬�����C��M������jv��Du��V:C�9Z�7��n򆐬�+��ǆ��1���C՚�d�ºb�Ŝz��o���{JZ���ڦgטNp3eIr[��%�����D(��N�]�3�:�jb
��+w��F]������4�3^����_魌z<�Ԁ:�%R�,�k�T�c喲�Xpe��H��J{���˝5�hz�B��&1����cC��)�y0O�6�y�\m_.���46.*Ci�x}���#�z��*a�)l@��_5��;�[�����H�!� E�X"������q�$�{�C���F���YX�t�h�'�Ī�Ja�4C6~�NX��A�:]�5��Z���Q�4��Dn�y73���b� ���k��Ғi��pIl܆X�rG��u�n���0h�s�U!��&oy��\�!��d�?��2�5��ğ'r�1�@�����26���:��K�r_E�v�+�
B�L�7!�8 0a�D-"F/�"�a{J8p׶dn�X �;�<��+�IR$�h���T����&��<��AI��F�!�!���ܧ��ܪJL�]�ޔ���'V-���vfS���k%SG�N=�~��)����1_��ɧM��%mtA��r	Z]���B�'<��W�=.H��2�N���炒IA5ʄ?�-A'�o�^$�T�ȸ�%T+L䭇�aV��x��S��*~n�2���8�ߗBL��zJ�Wbϵ��u���Vsa �V-�ȃ�X}V�Z�ц6�����6�mz�K{���Y�_��^.)�"l�ĚڥF���y=�	Ce$��"��:�rK|�w3o"zwK��]���XJGl0:�/2:}��g-������x� $1��J�hYD��mخ7F	��:�D�@��[�:�oQ�iNm;��o�O�I����T)��G;7#�!r�b0�c��77
�㗽�_iY7{�h�� ��~Q��@;�r��	��]�ކ&L��Zt$\��l��)�"5Eu����;��d���@B,�\Z��p�Jc��fq����)���%F1�-k@b���CM�V`O%�ŋ��W罍I�AN`���L�]��X��Z�9��l�a��0����@�j������@g~""X0��Ÿ�a��qA&m�x�	��)�mD���[.w���c��}��0/�J��/6�$�U��L����-� 
���Rb�P[6�<�r�9ϵ"D������6����(�}{��hVE��ሒ�k�n�%��/���^;��U޷fϱ��U�8��ۅ~H���?���R��\sYZxgr(�˴�`�����਄ҷ���K0bhb��ji��~!Y�^tt���F/�r޼���wN�Go-/7>�|�}�ԗ��VL&�������3�4�2���JS�͌v#/��[<$E����h��.@O�GB�� �ۑ<�K��[��y���x����G�H}%ET��s���.X�UaE��}p��V
���"�id�Wx�j3����m��@���D�b��-͋�i"��x6|����I�"ܹP.o�ߚ%���_a�,�8N���Ol��9�C�Ux�E�I���S��<�//�+���ZTҼy���@14�4���A��P�{�b
efa�@(HhЛ4z������Ji�=>�\�_3އ�ku-�E����g6��]m8��"ټ� O2C9�B��Eʸ� }�#
�E(���.%�>�$� je�s���ܰ6�=��܊(�4��������	��d�}��H��	P�N���ݏx߂�_��GI
:PW�ˠR�e�`U�U\
W�y/ I�~���nؓ��K���Ev8=ʹ�����
��D�������!�lhg�j ��[�ċ{ҷ�������8�L��Alxg�.z��-���	���	�BV��)�MM��Ţ�#c0�'N;9�>���fP'�_Z�oɨD- �Bo�Z�8a�A�\�kd�?�x�a�P���R�Q���."���L.��uƬ1l��l��{�W�*&FaRd�5(��Ci>Gjq�M�b���m׵�2_�}t���g�
�C��V�N�P��*(���*����tf"y-Xf��f��l�D`A�@�T&/���XM�<�t��C�+-Iե�e��������F��
ʧ!L�L�?V�;܃jel�(��� ֓�P�v�7#QK�{`|��ޡ��v���8����h ,�$�s�����l/:���+t!���==ƛ̫��ʾ��<i�$�<��׶����B�ی ����
F+��� �)qC�8]�!����N�>s��T�f��S���р��$Dh
��*�jq������Ȣ>�R�����h)��o_jˊp���@ا�۰GZ���N�e�6K�4�FѴ����&x�'�6Η[��f���1���Fċ}���M��Ix�A�V�|}��z���:���F�{�ƣ>�������M��hG��%�=��G��B<�6��f�h������3�3������^���p��L�v�l� }��RD[TrרRVqMj��5�,Zn���{����	���&`�<b��6�����/�\>���֍TϘ�3=�zg�e�6/._t����B��NV���Y���,oft*�ߊBX7!���wR��S�ۢO!`ݽ�8.�}:���}�ÉX+�0�r��Y�$��pt�?��?C��r*�LM$F��E&ʦ_Y��)u��Qt/p����T3\�O��+���z���8�E��_m����p��a��p9��� \s��5H�������}$��|�-�E�E1���M�K~܀�,�5�O��4eY'�[^*�R�~)x��E�ꦯ��k� 9�}-HJF��,��^jzf ps��[�r��XǾ���Te�l���	�T%�;��ς��mf�@�n���|ä�9V4*<&��Z���\@®��unTEZ� c���`��6����vk n �JU%�j��V��,��UKH��&�k����֒��Xw��Ŝ�!0��E=j�	��5�����рL��FVMy'��9p��z\v�vuУ^ЋɬC����rn�C��i�O�ņ�:���X�U�cd�w�b]�z�C��7e����	ۙ�E��֐�pNYr�Z�%��3�-��Ь!�N�,掸�%v7�C�w"�ZF8̛������3�^�YY��Y�G�<K�:%W�Rq�ÔU﯇��c�cֲp�p &H�C.J�ip���R��	���F�&,�ؾU�,��CD�šO����8�\����X�T6)?_i7-�A��9����*<Sql{f_�>�;�;v���"Hr� `��"��ɘ�q!�р���p��$�SXq�H˃!7'u�%!F4~��zLՃUA^�]C3�u�z�́a�D�b�7������bfc� �{��N��M����I���XWk�ہn��0#��p�+�� �Ψ�\~�d���房���5M'ĺ��¬�3��r��{�� ��9�:�bR�-l(БKp҅i�'�5!5+�0���?��F�;6�bw{e�8�1�H�3�H�A8�<#���D����۟_w��lƚ�����J�碖c���|ZdЗUy�6bު�T$]b���������Q�������SbA^�ɐ~Ʋ��/������|����x��t\!r��J��b��be꿣�8����=�	Ѓ��*8�3�5��r�hu��I+Q^@ ���B�h�+g��i�zVa{��%�Q�|Q�n�,�I�����L��RJ|[/b�$U��es��$�s\�P±�Q��sX�=�Z]�7�0 �r�����6��1Φ
��:�t{]_.�jl#dK�5B�F�4�y����H$j"|Y�:��|�o�L�K���XZX�#0U2�2�(y�BHs��sӐ�&"�����h`�ۈk�7���� *D)���`��+�Q�Fm�e��-D���S�4�Tdu_G�*##��r�Y0����
p���{ZYr�h�i��E?~�Tb@��&��]�y5��a�7E�t�E��g��)N��E0�f��z)ғ��겲m,ʴ��V)��XKJ���!D���!x�|
�� c�10�@���> �V�a,�D2���O�8FD���L�~L����SF4��rs̬|�?��������89�i��;��"}���{s��L��@mk�'	��~n'���.�~��� c��տ ʁ����j,$i��G���#�����X�P��?ܚ���ܭ���P���Fi�C w�\�䐘���d�jEޭ��Ì��.�n~��C���m�;,0X��XUf�{夐��I�,~C=7������h\��jZ�,Fr%F�+q�����۳��8��^h} vj仯YA|����ȗ�RF*�-�I��@io��>}�H|����2uVG�f���g��4#��2#EpJ.C���T���[7�����h�H�@j��Bl�����ڑw'/�0�ް��F&�xך���G��TX��T�ǀ�# �.S��a���}�z���h
[ "a�d?�W��3�s����@r��_|X����f<�i]�xр���FH�}s�P�s��t�p7 �:.�,2���!�g�g9/;U3��d���V����<բJ/dt��Z��O4a��[�7򓸭���9AKvkPzH��]2f�Ȭ(���O��_�?�%7!x��\Eނ�`ƸM-�����_�����Յs=�����z��2��'��F��`���38S}�G�A]o(+@�)�>�u %*�s�wa�W����^��Ҽ4&�����;�d��#��Ə~�24ڪ)[�E7�����7�
�?�����m�=���uU7/�>9� �i�~�Q�R��N K4��WْvӴ[�7Ď����.�ݠ�l�o�j��|ֆ��Q۷���z'd�Π��x���z�-�"��D��ؤ�V���а��g#~�1_UeN
��y��OaYf7��� ��*[DH��B�)Z״��|���s�kb��߉x�~OP��yRC�(���R0ݰmCh.�\��N������PWo�J&!3�d�Bs�p�>B�Nqq����15IR��2:Gdt:�fgp*C���LPu�X(� �*�g�O�9yh{b�>�����n�`����ou�/�F��3 �<Mґ��u��NI0n�eVW���J��S
�%L ��?�N�6P�j�_�(g5 ��˳��6�Q�l`��ޜ��vݰG8Fx���{����NiF�>�l�p��5�!���=�:��Ƣ�9�C���$Ζ�zy�����B�O� a�)�%=�ښ����I�)��K8�ƥ��Q�NT�,�TB���a��#��q�`�@ �D��%nG��;
��H���H���&������
Br˅�����b,Űb��r
�e�a�ں��׎��D&�����[Aܷ��[��o���iDAŞ��ќΞ�S�o|�xMzA7��y�ԁG�ǣ@Σ9x��4�!�l:܈�ᝊR��=�!��:��4}f�z��Y)��S �3���6��^�\_�T���F�v�Å�{I��sT�&�Rѣ�j�wi�g�D*{��b�k ��~��`�B^b:M�n�~�M�U�ʠ�>�e��v����AX Wgv..6
�t�r���),NQ+�bDb���,�v�*i��B3���U�Gw�?S�`Q���b`�A<8I��:*CR�X�o���\��������TEp/�i��p?��{M�L���6�&ŕ&YQW�u�d�� �	�K���\K�2O�p[+���z�8�j���"<]�K��a�
p��1�����ZH�I2���P�X��Q$.+|��x�@�1H�Mk�ܛ\�ڰ�g�pk�4I��'W7"YE`R@�M�̖�
ê�!�|�F��97�^H���'��^�� +ĩ�vR��eĘ��Y���B�T ���ģ�	G%p%E�k��"ϲ`$=�
O��,��4�'*�!� u�w\O�)��uI��Q� ���[�6t=$���%k;���šW�E�0ԑ��,qC�P]r�M��&=���X�����L8�\�������V���O�����9)PMTY*���l���v�B+K��F\CC-��n� ��O��d|�䭂�\s��Sd�L�bؖ+z��ؼr�k�����u�\B���9/pi�PrQ�%g��hA��Gw�N�����������w��'F�
����j�V^�-��s�i�؝<�=:���RL4���1��9c�R��jwp�o�H���JqI���?�޸3�xݏ&'8������C�1{O����\�;���6$t�i����VT?Bp�*��l�+^_k��;�;�BÑH-�S {	"���դ�,q\����YW�z;̖�X,@�˞N�'�EF� �4���������A�\�]�>����G�/�]D�H�7Tn��[�b�� ��R���?d��A�I��X���֭�nV�C0޸5�������΃�o�z�d'c惶A�M5���չ��'�r��� ��E����:Hd9���Ь� �8��#!p=�0;�B�:'+F5h���{�v�׬i�����|U@<�^��?��3��Y�"v�v����	�Wr��=�8��H��C�R#I�Q秪@}]=.�� �B��?���Y�'S}���D�~����j�+g��5��]ޙ�3��tw|Kr��D���̝�M�>�؛3��m���>���p���<Y5��Uѣ����^�0�
�|�#��+�&d���V<_Ȕ`�]��Vn�F���)�U��LԴ�J��rb������G֋sW�����>��X�D�Z؆t�jکI��E��6�����u�����mP_�BU.ߜ�l^�����F��Iy�T�n�$9G�"��:�r|An$oX?�K�Mf��X��?0p�j20�C�����	��QE3y� ��hϛ�ۣ�7<���\Ddc���)*�QJ �m�,����`����ŻT�!�Gq^G#�O*rbOY0J�5*�
��x�Y�ɉh�楷2~�@�r����a�,��<��r"tZO��b��)���E�S���ɵ�D�,�K�ː��`�J���6��ln�����۟=1k��@���9�!V����������S�h]L+�D�N�XwJ-|���
��&	� ��s'���p�6k"�H��u���W��g�fmF�	1���"���.-2���#�c�U�{� ����̥?$M]�B���~�h�v=y����FDΚ�&���o���9��o��)6�	����`����E��������ny/�Lx�Ȇ-P;G�*�K�~f�eB�����Tk~>�O��M��/\�1$Zn4r޹�f���$׊�����m�]����h���j_�|4������2.�F%���r����xl���o#�>X��|���͂;VB�%�t���"�4>X�2�MJ	�(�쥽elG[2,�D��hs��@�fB磠��)����Ơ�|����\�x��&��7�GT�3�<T//b��n�.N�a�D�}�]� �
���"<�dzOW�G�3�`�#|�@-��z��w�!�A~+i�i�xl�������*}P�1��o��t��P,m)݄���bs�9��/U�$�Ì�߮�v�<6�/� �D�Z
�B�&�v�#����ZA��P���X�f�(��2�j�a�� �� %��pf\��n�}��!.-`��,8�]�6ҹnN��X0)�u^F2�5��g�{�ʮ��}o��|m(ƴ��$�5>^w/ ��s��n�ҏD��� ��4��嶡�w*ڒp���g��~��:�S
߸m"��Gg
�N5Ȋ�h��C��V` Ut��y Q�~�,C�%��	��K,qǧҹ�v��(�VF��jU��p|�f���[#�l���j7��Wq��HX�!Q6�u����ϠdYOx��tz�-�h�����?�V�O����;��#��[��N����� ���:f>�P��HDc�.Be��Z�P���⏒r�k�����xF��P�}�R��p���R����.����b���u����dW�>�&�$�dpҼ�Z>=.q�jƍw�0���p�2�ztuQgjHC��L���P0��(ߵW*~��*֠y����ٛ���l��p?`�5�ӊ�b/ʸ��<� #�4����lI�V�eKw��E�<"�
�ÄL;ߖ?��G1�8js:("�  �Fͺ��~�Q�`��ޗB?v8�a8���"P��)]���le����_�!RbW=��:���yʴV=��"$	�;d����B:� ��@T�������M)�-�8������N��S�S����Ii��L�p�{�D��� �:� &o]K�����4�S�m���?��DRˀ��a�����}ꪲ��e���a |��Ǭ&.��E�[1Z�y���we�����U�|r��9���e|�&�z��L��Լ�>��4/����'�.��z<��~E=fa��J��l�f��N���h���3Ηҏ��^�S���t,�'`�v���5R���T��wRL��j{����ɟߑ�{�����J�9�`�(b��IJH���H�e�D>�H`�C���x��sE�g�[6���t%f��x�SNL�=���ʝ�,���*�&]B]<���Aw�LS��â$`S�08d�:����3����#�f+i�C��[p�7��?9l�(��L�,l��,&��)Y�E3uT��������|�\��!O9w.+���zL�i8u�*�������&�a@VpoL�����y�Hd���Ng�LH�r�6$i`�|2ǃ�;Yv1��M&��ܶ��+�+�K�4��S'�~�T��R�������%`j�0�!-9r��H��G�"��^ �Q �4������OV��T��9T��ֿt	�G% � �˕#������Y�Z	���	�/n7*�<
�І�����¤��u$֣н ����V?�6σN�o��kV���@֖ �|��n�,�*�K��ᨁ����ƌ�������������{���QN��
�U��H��+�M/�p�54}���v���B��C#����+n�t��y����@Ź�eB��?�dB3bS/%zds���-�L
���v,ڷ_��L6p��0r��%BDt�������VN�4��D)�������wF�	�PQ���^{!!��Y���\<:��:*uR'�T��Wg�%Z'c��	�&	'p�ّH	fJ��m�\9�������&"­�`��=&�Խ�O��Ka�\������6�i��Y��֏o�o�/�*�0l��_8�;�[0��� H��� �x�"7�"�q��݀LQu�u&���NX�Ջ˹��'6F�� �4�ǻ� o���A�;]�7��79�����J_DO�7�;����b�� B�z�*u�C�󭪗AI�kX������'n��a0��������t�^��Җ�d��`�~��C�B5�q���¢��ڟ��U�^�����:�� ������1�{��0!�o?0�m�5��F��^S�{�Eb�'����䷒�<YC�:ZX�y�8�E�=�͚�s��>8���������2c�]�l�9����]�R�@l�'�̆�M�w[��v�S�A�����~|���S�"��ɸ�0���Bt���rz�J�m����E����.�W��4��>��R�f'5[/���=��^���ew���+�w+�_��Vc���q>��Fnʀ������&1L��:Jr�"b`b��&Z����sR�&�g����X�k�ZS�=��ĩ�|T���6�}u�\�_��`���_�R.���l��h�kq�F�J�yN�ٕ:�$TD�"rzS:["�||o�QSK~���,0X{Y�0���2������+�2���I�[d_�[@�h���۾�7�Le�D�$��,�zQ�{ml������ym�^v(T��G��#�r��0Y�P�&
�z�S�Y�Fh����I�~b�@lo:��e]oD����st�x+�]C)�qE�۟�5Y�҉+�h��,@o-`��툓Jt���I����rE!���1���@3���4�MVq�@V`׋ t��.���F��k�L�=��I�Yk�b褸��J���L��{:i�5
�U�%�1��"3�4�0�\��/�⌙m!2�	l����5��qy.���Gb�c-����\������B$���=����ȭ�1^�7���h�����#��φ��}����Rո�]	��qo�ZW�E�K��9�w�<Ynt�����A�;b���ƭ4f`o��'�AB~9�P�\̓��\��Z��r�n˴�񲧿.��)���l�|�$h�:�j�<Ჹ&���F �7���h�C���*qo���>3�&|4P��h�PV=i��ϙ¥��4Yې2�5J�.�'z �[-�ɪ���h.Vl@�u1Bb���������f7�~����xM����HG~�Q�pTj��Y�H.I4�aV�y}?���D�
Q��"�#d��WI!�3�m�~(w@����������yi��x�2����3�P_���0��f�d��'�,���R`�]�9��dU�j���␇�Q�<K��/�`��ZZe��������e��y�A��0P�30�SU�frY(y3*���E�U?���2�9�\SѰ�x�D|��-�y�G����r�Ҕ'���%��p-2T��s�Ȗ���)��}J�	��>(a{���>�P� �ms���M�m�Ρ�;��4\ȱ��d�|��"��}ْ(钪�g*���S
��w�
K~��E�����7U����� Y�~�'~�}��,�KG�a�M��v�ϴ�Q:mݾ��6��p�Tjl�ߙj��_�2,��<^I��.J�p)��I`Q�x�$z� -���ɺ����d�Vϫ<�^��#���U�dN���0�䅨Tf�dc�p����=D~��B��?Z�u��I��-�nk��7�P"x�P�q�R9X�KhˡȔ/��6.��wƽ樈0j?�(�We0&�6dU�E���7>8��q'�2ZK��H~�2��t�jog��1C�!b�_\�P듀(�j�*�u��>Xy�!W�tf �ඞ$N�`r��ӥ��/}m���%Z<Î(���t|��I�^,e�^��A��
[��LvX�?'p�,��jv�U(� � '�R�����Q�i`M�nޒ��v�M<8��?�*,
��F�q9=^l >`�ǩ�!���=n�`��V�/&���EB$D��o���IB��i �V&�[�+ڐ�����)"Ӷ8.@v����N
} ʉ�����Α�'���`PD9і����{0c���΢��V��H����u�@g
�{rN�����İ�☲h�.ef�P'���&�tl�g�t[L�߷��ӆR{7�<��z��w�R��ɒ�|���z7:?���`������熣/[��Ԡ��E��3#�H[=A�Cم����,f��L������3�;��,��^�j���fx��v�},�1B�Ń��T�$�R�h�jV� ���z6){�(G�!O����`*�b0�w$�A�þo� �L>�Kj֞�3;+��gglT6��t`y���RNG�,�?��EE�,��*_z�B���ȯw#�}S�r2�`�e`��8$: `��mx�	2}�|Χ��5�p���:��?�U��L�`��l�s&��hYTXu�Y�~���@\���OԝY+{{�z���80����6���aW��p
�L��Jr���H	0��5��M ,$��5|��&�6�x1�kM�[����Uڦ���&�J4�%'���O��R�MmZ���@��q����r9�_�H^N�ͣ^{�W ��ʓ����[����o��Q�T6S�ֺe<	�%�%�Z��(��V���u'�ۏ�M]`�**c*Mx��-���8���&u�F�J; 4���Q�E6*�8�*��kqI�ǻ�������B,� ��F��������s�U���?�Ҷ����� '�
�����"��/N�M
��p��T�v�ί���м��C>"N�#�	n^: ��1� ����ùxՆ��d(W�b���z?;���NC��4����������p���rG�%�<�޽��}�N�}�柑�Vq���w�j�F�Ř��*;ܠ��^v5��)�j�x��<Um�:�ÒR�%�<Q���Mc����ǖpQc�H$'`Jg���7���Twר�j�&l��fI*��!���ifO�*<5i\Y��)�6>�iH
��rv�M%f�X*�P�l,,_��;����!�H�^ ��Y"���Z�Gqҥ1��hK�p1B�5��X������'�F�� @4/�͌���ƥ�Aog�]tx��Ət�=4���DZum7�)��}bwD� �~t�E�>��l���RIX�X(���e�ny0TF���f�u �9 �!dS���y����5~S�������zv����{,�����:�Ƨ�^R*�����������!���0qZ�0�$F� ���{�4�ע� ���#���&<�G?�5���A���T�X�͚�
�]���"��s��Ws�A������Q��6.w]��1�{�h��i��{.�H8���S���:K'~W�����6�gK��2��G��<t���r��\�Hl)��пt̹�)~��#L�:|��4]�~�!56�,�Ҹ��^�E���1��L�+��:��"�V�X����M��n����Z<
���HL
MKJ�>b;1L�aL�}��sM����~.���X��Zλ��>���1��{rI6�mηxi�k;ű._��.��bl�DE�9(F��y�����n$oa"�:l:6�-|��eo���Ky9ߚiq�X6J�0��F2&���X0�m�2��lj�A����hEs����72�Y@sD�_��zu7Q �m'���g���9GET�gG�%8#��3r��0��9k��
��^�.�Y#��hU����-~��'@'������{���0��t��1�X��)_�0Ea�B�P�w�� �C�P,{|��(���!J��@R|��7`S��9��y01��6@γ��/�5V�X+����/���-����La�C�D�6Ƒ���D�ͪǪ�F�VW�c������,KH"��6�떗��ĺ];�m���	��AO0a���.��g���cH�ͿqV��p-����$:��8���4�����Rʂ<���q���^(��!=��x��T�T���q��}���/Eo��t;2�ײ^no��A���R;}�h�A�vf;�,�AlI�N�~4�T��l��>%�\�ՏZd=r�Cִ�a�Z���̔%�#7��7��h��jU�{�`ƹJ���hӢF��(ɞ�������o]->	�|o���]V8j��*�Y��"�4t~q2��*J�dČb�����[(����!�h��@�%B�&?�l��(��**���W)Vx ���	
G�lB�uT�]���k.D�na�g}����
�v�"�d�W��3��h���`@�;	�	km�E��a�i��x�N9���쎎��P�Y�K�i�O���T�,�<��/
X��9@�Ud���R�P:�,��<��/5V��?�Z�GIe��𬱳�������A��APK�\�N��f���(4�����1�Н]ƶ`�)#L\��
�s���B�-����b�k�Sr�o �$�i�v�k.2����.�6ȱ�Gʤ��}%s����(�ai�M>JC V8&s�K�������E�v��4����3�u�hP�s�%Ӓ�s���A*��$����E����
�͓� .���G��L�U�],��9� ��{~�Buc�W���KbKħ��Dv�<Ŵ�|�p �����`�Ѥol�GIj������w���W,V�k��0S���Bx�e�z���-sT�����u��V�'{�z��}�#�<(��&N�<�*}�� |�f����3��[��D���B[#=Zh��-����;k�묺�s/x���P���R���&�ư>��.��p�c���q��C�&W���&�hvd�*ͼA֬>3J�q������f��ë�2�}8t���gAI�C��3��.�P��z(@*t�����_y�O�Q)�ݞK�`-g���U@/�0B��Xm<���j w��IA�e��k�:���2�
6_(L��?�0A'l^j��(�߹ B,0<`���ppQ7�u`�ލ`�v���8w�)�E�=y��ߤt�|l��T��i!�`=)Yj���ʪu�$R$eK���
-B�l� ����v�;��1�n�B)]��8ɬ¶��Ne|ɴ��V/�?T�� ��0�DԨ��oV��Z������{�*'��#fd�T�j�۩��v� �ؓ�ڰ��n����eA���(����iq&����"=q[g�m�oZ"�-�R�w�2+��r9�ѭp8턩=|���z��]���U�2܆�tk7�*��E�������R��W=Y����/袠f�`��jͬ��&�3 ���#�^`�ڜy��]�v�
���n��>c�T��fRB��j1�d�v��{怣�|����!�`E��b����Ck�������>�n0���x���/�g�G6�M't���̮�*NB{��s컝 �0,�f)*���B���w��S�+����'`Ɍ�8��:�|���ԉD{k����+G���fp`|��U�?/_>�M�L9�b���&�"�Yb�=u����3hz[�_$>\�[|Oo��+v�pzMh8������D���a���p����/j�/��H���
=-��(:1$�*�|h�a�1�1Y��M�����ҳ�!ܷ���4��'(n�JV�RQ(]ދ�[�A�����,.9���H�P-�a^�Ͻ \v��J���ƕ�{�3���2TѰ�ֵvq	XVu%vD����
ʬ[� }���%��%�*����F�����m[�u���F� �ǘ�Lm;6�p���,�k���6G���6��B��,B���AS�^��Ws(����v"�_���y�ױ���	=I�U��s��==e����M�-髮���v��P<��w��CYl����n9w�� 
������~�m�,�A�dC��bI�|z#O�#2���(���/�m����op�Ũr�(;%�Iu���8�N��@����.��w��F����#B�;��^qiY���[�3��<pc�:}�R�x��A@�[Q�c�-�ܥ�p%H?J⻛�A虏��Ia�&6��R���V��
6xO�vt\��v��N�6Өi�>��-6��c�DM*�:0lg;�_<��;��Z�S��H^W ̜~"
���5,qֹ�����k\���C�X]a��'w���`�4j4�UE����A�]/ٷ���긯"{ �D���7%7��>b�$� �j��`z�937�`��I�2>XÍ����ng�}0����gt�����a�H/Dd�q�t[��l59U��&�U��Ub=�Xc{��� 
:Y(/�ߝ����qG���>�!!4n0��+��FF����{�C���+����-m�<�l �0���/�QKB��s�u��α�8�%��^�	��"�#cЃLQ��6�����]Εa��r�]�ކ��B-V����S��H��X~2�@�p�8�r��F�n'��d8�t�Mrp�z�#Z�NJ��Λ$b��~����J��O��H5A �T��Y�^<*���T��+�y��U��V��ؔ�{��+0n�T����n���DL%��Jh��b Ԥ��ї��sH1��cx�orXZIt\�ɩ����a6�})����&6~�_��Q.pkl%Vġ UF��ry�����$��S"hQ:�|��o)�sKt���ֆX�Z�0��2�-�󤁨�:�*q& �A_h �����7��XVD��bCFp[�Q[�hm�@z��e��o�8TP��GB�#��rs��0{�v���
⎽	+@Y^�<h���5~�)@��޳�e�!��HA#�t+,��S]/)��EK��k���Px���,���c�W��8LJ*^��M�R
B�h ��lr1�@i��*�V'�U����6~�$h(��u�8��L�r��?~�!O�^V5��*Ū�3��1 �$�����y�'�"顸ঊV�'9b��	#m�MY	�+z갤��y�.>��?�cc@ƿ�o��Kv�V�$կ�3V�ُ%x���s�mX؂�m�L�Iܙ��ϼ���s.�����Hg���ŒP��EJi\᯵��rt�nj��]��ȷ,�;��ӗ��Df㹤|���z�~/}A�,F���\��AZ߂ro8���=Ń�d�~!͐���h���j�=�� *��<a��mFB�ރ�4��ZJպjo�8�>�S�|�|�ԞkcV3�J���p�Sn�4�AZ2,J�ZꌝY�6�o[#�Y�U�nh���@ֱ@BX���G���cXŠ�mU�̌���`x�a���Gt)�`IT�$���.?[a)�}�m�,-�
G~�"͠�d+f�W4�3��H�4�J@^�0�x��=*��GiI�x=�����[��P����f�\�y�,����ES�b9�O�Ufp��2b�82���<���/а���9Z�\ }���W��ͥe�[A7��P极�I'?f(j^(�Z����%�K�Ƒ�]d,�\�}�n�2�-�}�j���Q�J��_�a)�p�f+|2
����mD�̄��} �-_(�h'�'�>oc� }�s(�CN��sܱ�`4������}������2�T�|��;:�Z�߉�;��7�
=sȻ�d���/���U���*z� P��~�}(��r�:�>K}��C�v����"��"��w��݌�l���jvy���NĲꇷ�IZ�f���� ՠ��x�ؚzw�o-N�8�0gO�V!V�����ȰlU#��KN����e���o0f���&z���uD�-B֏�ZC䒜hi�c.ak�~��&xw1�P�mR/���H�>yR�٩�.����s�ш����^��W[�E&���d˷h��
�>.uq�`써�o��H>��2�z�t&{Hg��,C�'��!�Pa�(05*ݻm�yTH���[
�|ߞ�h	`�/���5�/s�����<9ˏ���r��I��ZeB��U��MN
]RL�?]�"`j,ml(S�� ]�5��k�~�Qrl6`��ވ�vIj182_ث`N��=�ֺ���ol6��L!c^�=�MX�2G�%%��#R$�?�?���_�BKa� M63ؑY�چ7ٍI1�)�}r8d9���N��T��a��nߺ�<��9��,!rDo���Z~�1��n�I��P��e���ѳ�v�q�[r���N�T��2-�^8MeM���M�����&?������[����|��Ĳ�H�c��m���<�?�|� z-�������m��� �%� �X���Ɋ>tc=�����~�=�<f�B\����?sv3��"�M^;��@����l�vѷé���:�T���R���j�جSLj��߈{����� �j��``kxb&����ı9/Z�6�>����T@C���$�Ԙgb��6v��t����IT�N=���ιD���,��*U�B���Ae�wY�S���i`��'8��S:�L�Ĩ����7}�����!]p{�pw�?������Lt)줢��&���Y���u�4�����t:(I\7��O
K�+qϸz]Ʒ8�=:L�z�ŷăa�~�p@aH��4ކ�+�H�H>�%d��`��F$��|5�,iR1��tMW����ڜ1��ܾ�45FR'�pE�iR�"��#��v�Y�����99#�lHQc��y�^1�� G|��2��Q��V���[�Tl.�ְ��	���%1�X��Q�L>ʇas;>Y��V� *O��������Iu��Z�¢ j��G4m6�N����k�{�Ǳ���A�}��,�}�<�ṕ�p��9{���[�:��H[v�L����b��;�E�X�?�%�M�`���'��! v����(��2�Ctָ���n��;�V���й���������d^�bĸ�z�*l�^5k�ꦋ�P{��wʘ}�p�Ar=l�%���T��гQN�o��U�Ĩ̸�Iۂw�g�Fag�=���6�^l���s��r<�y�:�VRR��ה|dA���Bc侙�7��p��HZ	�J]�����ʵ˨�w'& ��|ހn�'�%"�O�-���\��Ǵ_��6�1i��7��!��(\��*�D�l��J_םo;�{Z�� �H�� �^K"��0��"qH&v���f������XWo�
C/'���l��4�y�����rA%�]�YS�����3K�VD�! 7�d��b-%� sv��{�����;Y#IΣ�X^&��n¯{0�Sk��ժ������x��d�u��o�rT)�5�v��A^���g�0n�������B�:����ԋ��`�����n�=!\��0��Q�&�F�Y�9!{�rט�¦zo�h
^<*�Y�+�	������Ś�+���CS��ľ�}�C&C�>�1��;��,_ ]�M���%��+��73����E��S鱇�0u~a��V.�R���XV������t�(Vr���g}̉������fd��2֨�9&�j�'�t��5���яZ:�P�j^K�v�� 9+�*2�ЫnV�.)�L����(n����ϳ�A�$L@e�J㸺b�.L�׸K��ܗsC���xg*�X��Z�p�7��5�m���6����m�ݐ�P�u�_xXS.Kp�lJ%��<(:F���y_V�kE$��X"�:��|-��o�I�Ko�Ț\�X���0�Z�2b�剮��㢶�p���l�h�ʃ�+�7(����DP(����*k��Q���m�����d��~�H�T��G�l	#�+.rΨ�06nw���
|���AY��uh��摿�~s@�%�,���J�ި�B^P"tƵ��N�)m�E�2�Ԇ����|���8,��������J��O�A��m����m�G��1W_U@S�%_:V�����M�Q3����c���s5"L�=��:��|,�߉�˪�׍��_ _�&5�"�"D���a���B��S�ym��	�F�Q ��-�.�?T�x�Uc~��g���&�.̑o�$p�\�.�m����b$����.�2���'����&��W
G�nx�
������e%E%(���O��V�neæ����rld;�Ǘ7��f�LW�����P�W~*]ʱa�ʹ�C\��ZZ�rJM|�R����H���^��+��RLhjK���ݹ���Ȟ�F����+�t;��o41>ľ<|�B^�9�`V.����Z��
4�$K2�e9Jup���*(ю[�K���h_�n@��B�)��"m(��4-�7Ѹţ\�v+x~��4\eG����T1�*�.:��ag
�}pz�G��
¥ "��OdfX�Wn�3�T����4@K\� c��ͭ��i��ux�w��g�DH�P���Á�|ת��,Y�l�#/8N��9���U���9�A����<�/k+��sZvB��<b��1����@b<ArͿP����D��f�"K(�)���!�ƺX�lU�U�\$c�ism���-L>����I�]�%R��^��aZ2e���G��ʚ��}��ZhY�(2�=�!y>ʜ� ��Ds3$�Ͼ�q�_����,4-綍nD�+I�Ƒ��M�^���ªpUZ�?��$�ɻ���
\�r�vV���P�B��U~�7�e�' �/~�ؗO�����K��᧾{vZ���B3k>���H��hb�G��l
x`j�$���X��`շ��V�a��Z1נPGx	lbz�)-)�1�k�`ث�bV�L�o��'�j#��\/N]����u��V��f홼���$���Dϖ�BQZ ڜ�������k�o��av�x2�VP&oR�~��\�yҰt��.����λ�a�7�y	W�#&h,ide�w__>)��q8H9�crY��l�f�2���ta3gw�>C��
�p3KPM;(KJ�*j?Bݖ5_y�=�E������5��`�&��5�/�|�z�<t��!_m�I�72e�Yp�p�`�(��
�zL'�?��t�j� h(�� x�c2sT�Y�Q�P�`o�ރ��v�(L8��J�{}"֕l��6l�aF�G�!�G�=�b*�M�[ʠT]�^BB$�9��`���gB�uG ֿج�����$�w)ӂn8��#�Q*Nۮ?��;V�5������g1QD
���eb���I$��2��� (�م���P��C�l���*$�	03��Ӳٓ�e�f: ����&&�U2蘴�[�P��e���|9����K���h��c'j��6�|Rz���\�OԨ4�Ǫ�@� KR�����c!�.����=�А�6�����f�Dn� 0q���3:���6^oݜ{����v̄I�B'OŴ2+T�vR8��j��\���r�K�{ܐ0�2�'�%�`{E�b�����N�t��ю�>��֯N�d�ߙ]g��6Q�ts���.bN8�!�)�-�v��,��*�4Bz(��|�w�[�S��f�q�+`?�,8Е�:��)�v>��m��-w���Fe�pֹ����?%Ҝ�L��)�=͛&� �Y?Hu@EG�pd=L$\rz'O���+l)]z�_�8a]-�7�Y�Œ�Fa)p�R���YΆ���HP�˻@�u6���l$Uuw|�y��'Y)1�)M�Q�"h������4p�'^��@��R=���.�:�R�����9^aBH�s��o^�:� �7k��:��̽��1�"�2�T̼֫��	�%��7�Ʋǔ$�b��v�����*^�W�����r�~u�Y���� �_�B�6;�x�[0k�D��, ɖ��Ը�,x\��7������͌�T/Q�� ��S�]G������)����s[���ugM�2+�!���%ւv~Fg�o���RC�`j����n�PE�vy��ֆ��(�#oշv�dyVpb?�z�Rټ�X}��t���.��#�8e:p�e�r��g%��6����N�N��氊q���d&�w�FZߦ�<v�q��^g1�:g��q�<���:P�R������G���c��A���fp���Hu*J�$���������&*��w��) ��@.�O|Q�QY\
7��q�6]6iYׅ����v���*^npl���_r��;���	��H�L� A�" B��Xq��f��o�av�F�rX�lC�%�'�7?�G@4���������A��~]��R�X��16�D�'7[��� b�E� .�z��A	�/ ��/�I	5aX��lֽi�n�0�
ӣd	��	-��B��G�d$���ji���5����\׾n#���A��Lx���d:K���X1�3Ė�g��I��!�xm0B��!ȽF�%�?�O{��&�U���<�K�&z'������[��轚v���1��~��D�,��?��Hc��V��`Q��'�]�%��,���'Q������2� �S®��%~~��'���n����b�$����Dt�#�rfOۊٕ����E�@��K�4֡�kHf���i��K5����N	��0^���ѓ�ʹ�+	��K�PV��I���	��yn��.�k�ؽ���L[!�J^�b�]��ù�N.�s>��Ӌ��'X:HXZ?��l�p��LH[6}�M��H�����_�-.&�l�E��O�F��:y��n�&@$�x&"^<:�!�|h?o_��Kj���z^Xgܧ0���2���d�ށ٦��ghѦ��8hv���*~�7�f{�C�D�i����&f3Q�:mX��,�I�e��y�T�^�Gx@F#�rr)Ϙ0�_<��
�Zӽ��Y�=�h&���Y~�\�@X��G�\[��ރ64��Dta_�I�:)p�nE�:Cԡ���u�����,,d�����huJ���Ԃ����^;��"��1��2@��r� �VV�okBS�l��9�>e/����L2(��5���)�ԇB��x�����E���c�����w"��<��`�]o����m��R	X>� t���.����3��c�L/���h���,$��)t�EC�n���:͂�:������v��&�i���e8����:b��FU�E ��%
�W@n`��^��-��;�ZB��ׄf����[)��3�~%]ﱼ
��o��\0<�Z�m�r%���r��+̈́����4V��h��h/Ujƾt{�����9;�FN��9i��/<(�o�O�>�I$| )7�ԦVV)-��;���e4�'D2�RJP��5l��[�Y��uh�@n�BN�w��MH��0I��TT��h�hL�x9���O5�Gj�zXbTV7���S.5|Ha�-}+��b�_
=��"��d�j�W���3}�}��@���F�B�͈�Ti���xs<��{v���PK?�Ü1R�?�\�,��R��^�I��9Q4�U������|i����<7��/�Y驉Z��������X�u��E�A�-P���?y�f���(e1��W&�Ay��G��ڞ�\�ө�d�]���-�&��V��ؕ� K��Vn_:�\��2��F�_A���n�S�}������(�ի�;�>%�� �f�sN@��9mK�:��'p�4�Γ��S���F���h��ӕ�K���z$V߿���w�
�{��1�k����+�UY��Z� ���~�S�t)hذ�K����9�#v5���}�#��Վ���-ns�W�l%@�jl�Y��W��(���(�J�\���aY�Dx$2zm��-��ɦ��FǼV�[���,��q$# ��A�uN8���!����f�@���fz��e�D�pB���Z�;��f���K�k��4��'�x��PA��R%vb�C����E���.��C�)���I���u�WQK�&C��dA2ܼԜ>$�q�O��eg�94��2\Խt��g�C|���eP��(fu*���qWy��1���T��x���`^! �V�/i;��U�G<��ǔ;��hj�IR��e��􋭻�
�
ǸVLb}�?�2l��j�(�� ����,i�4�cQ�T�`��C�~�Lv�'8��������&��p H%��llXC�(!Q�=Z���h����s�9�"$0T��K�i�B�� ÕP�ǧ��|L̍��*)�~8��8�z��Nv:)�4ʃ#��߰����C��adD��*����)�S�MC���XJ�����(B�1\�g��(���Đu�b�Te�s<������~L{&�5�S�[��H��MV���(1�4��c}�Ѿ2s��|:m�z#�7U��r�E������V�dH�IX��4�=��J�qu��s,�f�f��{����l�3UR���^�ǜ�o1�.��v�qK�����oJ\T/��R�r�j�"��&���I{�Haʍlo���`�?�b�7�����l�>����
嘘2/�~�gX�16,�FtL��)�N3����v�1hD,,w�*KBUk*����w���S�Ƣ��m`���8�P�:�zdK����m�v�w஡�)p���㦣B?�;�o�:L�q���&�ϾYs�mu��1���R���\�9;O@xw+g�]z�8�cH$Y��m��aC� pvd$�ݞ:�@��H]�[���,湧�$�J`|9���"i�1j��M͆��=i�ڒ<�(�4��U'���;��Rbw�F��Q��3��h�A9�LlH����	��^�0 �H��c\�G�߾��=(�T���֦i�	i��%��g�R�C�BD�=��� s��?��Z+*��{�wz�q��@ukJ���� �"�="�6��c��Uk�-�ǧĖg�*��	,[x�2i��o����i�o�������ׂ�q����<���j������Mv$��\������vy��M׬Шl�C�
ğ�<n���Ry�ކ���~��rT�d���b�	�z����ԛ�S,��,��~�q���5p�)r3S�%�¿��6���{N��g�s��B����w��F5}v�w���^b� ��z�d�<�8:�i�Rn�I���,�c�\&�� �p=�@H�k�JS������@t�&	T��.����[ZO������\E�F��3W6R�i��v�^5A��LR�s*9�(lk�_׻;��-�d_�H��# C�"{R��ƪ�q�&��S��\�����-X��[�@��'w�;�"��4�_�&��=�A���]`���20s�)�b��DFN�7���Abㅪ ����]��Fw��$5ID��X���ָU�nxfX0@�ޣ-���z�Υ���d�ܞ�e �
6M5j��wp3�	++����|N��&���&�:j�JEQ�NH������$�k!�J�0ݭ)��FWF��{"1�׎x��0�)�ޤ�<`�Ծ!���@��|����B^��F���~�����߃R��"����д����˪"�]_��g��.�N��s�>>�໱�S�&Ys~Æü�
�	����*k�����Nt?r�������ȿ�Ν��Nꏙ�&wJ���ӂj�5���c�����^�A�,����s�+$�I�ƴ~V^V:�����"n������ݽ�=�Lv��J�W�b���M���ns9�9�.�V����XUEZ��`�eJ��F���$<6xmJ�#vҐW�1��_n#[.��l����r�,F�19yk4���$��"�|�:�q|�Q�o���Ke�"���YX"M0K�2Yc�?���Y/�P#V�8��"�eh1���E�7=���`D���3};a�$Qlēmu�G W�����ʙT�LG4�#��r�0�q�� �
r�罚��Y�dh�_��v~)�p@?�b*a֙}�^��4[t�(��D��)˅.EMb�Լ�����'�Oa,g�4'x��0tJ;T�>�S����وQ���W1�oD@:r��e/V8bV�T�������r����[}L�2c�08C2G�P_�9k.�~��o�\��\ =�/�"�?��%��x:k�I5Lmh�	����������.O���{[c���]|���l��w$�2��$3�٠�H���S��۳�(����=�J��ύW^�dl ���y���U�Ӓ�d�E��`��Cy&n[MnR���K�;��E�-2�f��¤-A����^~ }��*��*�1\K�HZP�r ���b����x����ҏ�}�#^�h:|ajA�
V�5�6���ԝ�F]ޔ�7��\�&.o��>z�{|[/��otDV$�L��{����4�JE2�RxJ+���N-��p[��f��h�'�@'|�Bɬ���N�M�m�'�����Bx�F��j.�G��U�T�:�`�r.0^Ia-J}��}yJ
�T#"^E�dܜJWPAs3x�҂Ef	@�ڿ��Y��c��i��_x!D�v�Q���P��÷�/ͅ$�7H�,��l�Y�FD%�9��/UP�!�!�@������Js<rIV/����{Z,��QY�2��� ե�GNA�iP����:R`f9�( ���2��W��"X�	\Zdd�_�jC�-�;�μX�?��ۣt˂�5��W�2,��[�ʐ�}����7�(h<r�uC>�o� B�si|Jϴ,��̛�b��4c����XF��q�<ѫ�������&��쵹��Z����Gd
K���X��*Њ�8�^U4����p !_u~���#C�kI!K����v<���i0t�w��������ݽ'nl@(j�ۦ�y���c�̷�b7�W���[�Ɵ[x?�	z���-߫���J@��.V�W��%����X�#;u��?�N@Ռ��
f�z�7��G׈DɈBG�+Zԗ؜>e�4
�k�s��Mx�ǖP\�R��f�J�￭���J.�G-Ƅ���М���W̭�&p�d|���hr>*9q�v3��w��{����271�t�g���Cw�Ғ&�P�h(���*`��L%�y�z�{;��V��4`J>�,��/�~f�0d<��֬~c��I�haes��������
�1L���?.sU��j=�?(�� ��7(��ԿQ#y�`T���yvZ�8c\|����Kr�K��`�@lo���!tz�=�z̃w�ʖ����$k���d���B\�� ~u���~�������)I�85��u1#Nѹ�����>��+�Ȯn���ݱ�D@G\��^�BD���h��y��%��@���G�L�b�������زϪee��w����y-�&P6����[�6��[4Ն��`�c��ͮ�^)�^�pD�|U�lz��
����*�y�D����3�d�ފ��.=���٬�d���f�������p�3pP
���K^̼���B�ə�v�~ɩ�_��*��TJЦR.�
j����Ŀ��M�{� .��C׈�lI`�Y�b�;Vk����@��>>�:��e�#���?g�)'6m�t����D�N.s������@,Gg`*���B0���?�w*GS�O!�'K0`�[�8,i:�X�Ur�0����{���K pLw���i�?ūJq	L%F��sd$&��*Y�{Su��L8�f���J\�#O�>[+b=�zn��8��Nc�fx��H��a~�%p����#��ؽHƗ�v�k�d�a�$�?]|Ԓ?���1���M��c�Xۼ����m�Z4��%'�̷6��R�ѝ���ǮR�~3"�C�=9�W�H"[�k�^B% Hyu�3����4&�����x>�T=g�֡�	�W�%bs5�m�Ȳ��o�3��A��T�{���*�?�2O��4�!IuF[B2� ;��8Ik6���ѳak�6m�"9�BfW�.��,�yî-[�����C&����&�u����|������
S��p�s���lR[�������xMQ6i�#��[�Pvt6��^��c�TC��ş��wn��N�쪭'b���Rùٳ�-RPd��?b5b�z��������2��J��ٯU��V�p&�zr��D%dո���ЄNN���f{K���4��w��F;ք�H'ܧ�J^]y��_��L<�{�:���RI\��-�p�ǿWc��F�H_p��|H��UJ���~��{q��{v&�Ͼ-����i.�v��Or����T\�Kt�086g�iP�u�!���*"�lS�_�#F;ѻ��>HJ�o 8e�"��hա�Tq����C�WHE���(XI���[
�'�x���x4VK�����A62a]�~�M(7�ݥ��D��7���Ղb>�� �Y����%�O��:I��X/�Pֳa�n��60�׎�H�>�y΀�84��dZ@��`�e��5%�Ē)���Q��5^������/:���RU�i�9�]%����!==0x�ɮ��F�����{=���	�ЦU����<�>���7�7��߼��l���B���z�0��%:T�c�oCk���I]:5A���^��#��A-���v�S:B����T~�Iϼ)B������o��H=�P��t4zsr\ll��Q4�:/8�{�2n��|���Ҁ��e����5}���@���!�^�7����@M�+?���A��V9�����T$n�|�!ýr�L���JT�b�U��7r��1�s4�K4��[qQXp��Z5pr����<��!�6s���~}�a�L�X_�8a.�^ml����9F���yp%:���u$��"T��:}��|޼�o�a�K`���0��X���0-��2����؁����`=�)s�}�h���`�Q7�3y���DL���%h\��Q���m�$�b���[��;'T<W�G�Gh#�`hr�{Y0g��i�
�SH�u�'YJLh\�H�U�~�_�@��س}~�Qqt�9���et�[�?7)&B�E�����G�k���,��?�{��J�;��YH���T�ŕ��Y1(�@�1���V�t���)��5��ζ�Ԅ�$�Lh]�+�l���J9�Tk̪����+������x-"U�����{��%)�ă�mC�	��$V󣖲	�.��g�z�c��8��K��ْ�B�w$A���W��^��aфٜ₣㿚���܅�F�(.�_����4�ِp�S�<�@E�$(��#�޺�nV¥�f�ȣ�;iї���f�J��hF#�!m�~��ri����\f �Z�؈r�K޴s!�a�$������
����hU�5j��l1�ٹq��o F����sN����A[?o��!>U�C|�UE�
b*VO���;ϥ?ݭ4��N2���Jr#��^�8L[pʪ�z�h�~6@B�@BD����o��O����3��4�Yx�(�GG`[k0лT́����.+`�axnG}�`,�}�
3��"9��d��W�ڐ3s[�����@J��7u,��4�>ˢi5V�x�%C�q�1�U��P�$����H���O,
c���b?�9��Uݏ�<�p�r�s¨<��:/<[g��IZ��k�j�3���kԯ��jA#�cPR���5Kf�(�)͛'nG�7V,��%�P��\�7�Z_��S�-}�U��B���K�ҶK_K�Q��R�2v���Ք$�8���\�}l��א(Ð��2>�� ��!s��0�/C��ܝ�F4��U�~}��<6�� D��H��
�c��n��U��7�
m:2ȧ3�E�����U�1��c �&�~թN*>^�&��K�j�/]�v�F��4�-�z���ص�xhl[0Pjb�߂T-Ğ�v�^ �R/��k"ޠ�,xZ��zc<�-��|�,�|��V�sY�C°X_�#VS�7�N�H�Q���'~�f��2���e�iD ��B�Z���T5���gk�%\�r��xc�Pw��R��mq��*�	�E'.�Ē�߰%��xU�ʓ�WG0&�ANd�,��H�>r]qI��������*o�2�\tlgH��Cr�P��*LPM&[(�I�*�(��'M7y@����4��F`Ԓ��G��/_��7_<%�ϔq�^��I1�e.u���#��GX
}��L�χ?��Vp(j�z(?y ���������Q^�B`�q�t[�v�#8F;��y���&���8�l��E�t!���=�`�̞�
�����^�$��R����B�r& 9u~��u��r��)�R�8Ы*�p�	N,Y~p*ÃY��ߦϤ�I�#�"'D۾E��Ew��5zΤ��s��u�j�R�{� ����]��ު��:�&�:S7�Jf�e�8��l{�Ύt.&�Vy���[�٭��:`�t�LĞj��Y�Q�t�e�+�|pi6zC����o�Y���{���f��!�D��*v�*&�=c�.���)~f�
��1���+�83��*�ix^��j�,�F�d�Wv��éS,����TeR���jxJ�?���i{���C;_�VO�`̓b� F��%������>����	�I0�\gN��6�D�t�̵~
N)ԁ:/)��9F,bw�*A�BQg�-�w��S��x���r`p�T8!'+:�	�0��k��������(�W�vp����Ot?�n�%J�L`:��&���Y)J�uq�g	5��_�w�\#�Ov%�+]�rz��8�~|����#�/a��p����ӈ�����H�G���@��u)�o;=$Un|oOs��V1 	MC�"�smcڈ�Z�H�4!*'/�?1�5RL��z!��+���Sj�܉9��H��1��P�^��] ʐ�N�=�X�°Q��tT�dz֜�@	(+%O���;V�8X����'�����b�2�*o|����O�m�#�u!��m3� ֩.�3��6L�y���1k`;ǝ���BT�i1f,I�f�(m��%z������.��+y����4$s׸����M:�i�'Z�������M,h �Ґ$����voޛR�rC�o��^n���'#�����*�4�X��o`d�uSb��Kza��J������܈C�4���i�XpAF�r)��%?"�@3Z���N������x����Ǵwu�DF�Ƅ���By�^XMR�Kq��M�<�w:x��R$�|�h5��b��c�z�����p�=}H�M_JI���Y���PA&��aȀZ>N��O�D^��\�����6��-ij$����q,x�H)J*��l��x_C�h;̻q�>�H�� S�"q=~�|�q4�p���j�RG�W�cXnX�v7;'mI����4�&!�\R��IA��b]֜��h@�����v�D���7,[���b�f� _�%������3��p�I��lX���֮�In.��0���c������[��o�}d��s�[�e���5�=ĭ���ڜ�9�<���ۊ: ����~=Є�'��l���Z!HO�0A��FKppX�{Xo3ׄ}���6��T��<���"*��mC�O���V�����x��/4������H��oD�*\�)��A�]m��2&d�ц~/��x��1C�SU��� "~y,K�Bg:?����|p�5!U�k�tO��r�*Ǌj���ux<�������E�Ũ�4���! �`�5X4�{��cq^�'��R��F$+Z/���=�V���8l���L}n����|t��-'�L�8J�v�b]���á���%s/j������X���Z�Z���!��>�6n��ٴG����g~�_dn.�Cfl6f�Ĩ��F{jy���Ww$�?"�]�:Xq�|Ho0T�K[�욋�qX��10H��2�����}��;0����:>���?h����{7�7J
b�8D<�Ԝi�Wg�Q"[&m����}<���w�[�dTwxGI{M#��r:Z0"�#��
h ��PjY��h�|	�}��~�V@�ؑ����h����J�dt22�:N�)��E�i��Rp��\�eS�,�k�j�0�� FJ�B��La��<��σ敳�1C @pi��V��s0���G6�b��ϼ��_)L���&Tr��BŬo�R���-�x�K*��KB��"���M-ϸ�0�?�NmC		�A�`��=�.M��d��c����S�*���i�}�+$�)ަ�V=��N��}Y����E����l��$֫Z���v����.���f;���!E�c3�����y[nQWH$���^��; �#G�f]4n��k���9�~��ȿ͠�\�ZF��r��	�>����������E�ސ��:hpv�j7� ι�$��
�F��p�J)Š`��\�8o�aJ>0�{|ћzԥoV��Lg���A4�_2v��J��į�=�?[
�,���hK�k@]�$B��=���ȑ��ՠ��w�?��y��xj*C렀}G۷$��T�A��c�.&�_a��$}\���X
���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4iy^�����i��]|$-�'��������f�j~tɛ��T��h�6]�X�_3;B�s����ݦf~��fcÌ>��K֯c���y��b����PW����ܦ"������T���
t��hRDj�Ŕ��V�2X�u�w�0��jH��w���vF��P� CO�2����E�DTr�B� ����8-�����-��
z"1Y��+(h��D�}1��2[+R��e�{_�r���UOʖQ��˪Nؙ֬߂�`�����.0��0�C���T���'ߏ���(�1�`YpN���6;z6k��I#��Ʉ~M0�]c�F
��5�����}�o��P1
18ѓ�dΔ"S�F�.9+Z]WX�.	w�⤠�bAM�ӹ�����D��aYmu�[�$۠�k�k��2@�k��CR�y�pۛ+�m0f2A9!?Ç>�TUG�ֶ�&|1�+��f���3CtRD��q��0���{��'a�P������bC����P�=�Ŷ�T�c���^JUP�$u�Ҭ�LAɱ,�,�����Oa�5Ɖ�M���q���E�x,`����1m�e�j��[(j-oհ%2����]{��l�I-%��<�m������т֩�9���Lu�OV^v������牫�#���"�w���U�^$lC�M�pw*e��M��x-`Yr9n���`0�u��޼vE���Ɯ�`�NS��(HJ����@���$�����Jp/]W�C�V�g_�0�Z0;в�w�i[$�ʎ�J��lފs��C�_y,�d�߱T����9f"��̀l(��9�v�����?F��e�'/}y9-��~�<`#�-��cw��<FH�ׄ|��|ؤ={���X ��G��RHx~�}�9e��8$"�힘`._	| ^�(E%�6�)`��91zØ.[
��Gw��X���2����]�H�?zz;��߭ڜ��V�+�?Խ���Z����|5�.t�d RXM�3Qbb�Դ���zy���f��oEkO�.ce��!��Ӊ�9��s�z򆩝{� )|�qQ.��d�@B�_��7R)ϛ{�'A �u^͗S����U$ ���Ɉ�*%����#|�y��
⶘;�u�UG�5�>'4��&`�/?�p�/����G��d��Ó�#�<��]��/��4%��'*��}CR	q�p�td�<'jL��Ω�٭I��� ��!*	יN����5Z�Og�9h'�X�����{d��O�YǪ�	�>���N��
�hhj�u5x���N��Q��3�+��n�n����y��wJ�=+F���$�:����6����w��nG��=Jb���έ\��-�Q�\�̋��Cb,��!䜋�`�Z>(vq[2���QI�k6˞��L;��{_x�q�C��N�C��<�)KKCq�L��\��?'�Ԏ͏�/�]'X�>��crK�5sЈRҝ���\8ޱ%��fF�EX,$}�z��e�TI��i��0{����%r�J�^��R\��h�QDV�t+'�8ב2��Jc4*���-`�5�~�b�Q�u��.
��;v隙� �d_��^D�\Z�}Vz�fa��p�B٢��KT��ѣ*�Փ����5��fBK�+|x��Ǘo�6��h�a8�X�]w�8��Z�$� �7�T/��vy�����vER�������1	��6�d�/�!R$-K_
�v^���g����x�I
�o�m,���ˆP�t�����וg�L|l�<������΀A��pԀ�tm��^���G��\^l/ن A�<�#Y�𣡒X�K��L9���ٸ�t��!�yR�(����|#</
��em%v�,9���6��(;WM��2�h�T�j�侃cW��\z���"v�1� �У��$D�P�%���P��wʙ��?�3I7ܪ������!���^em!�7�`��\����j~n:�d����"n��@M#T�6�����4���A���
{��,�$*>���لґ6<C��H�&:g������e11�-�p����`����V]O3��y���?�s"����<D����"]��"I��/�{.U�R76�����"�O���U���{D*�(eUD7��<��J���p��94��Ҙ�D��f�W=ְ���1@���ln��]DS��V�{f��ba���cm��9"��锃��*�"�A������ۙU�X�!��pb��=X$��-%�t�����	4sLҊ+�����R�B�3�����d�����|�I����� ��RkF���podK�#�����1�矄W�����n�0� �ya�:#����[�Q-�>�����G.g���yp�*�K����L�S��T/�a3n�떑���%79Y`�fRꖧSC��ذ�{�'�d�f+-
]nn2[B`�8��Ȩ��4�Q9æ��PU�X�-�c+�-1��G}\���a�vw���n�V5o1=N̰	�k0�y�5~,�^3="��Y��!�S��^�,�����P���)~��6�n�0��ڢ��MuD&|˳$u���
+���꬐�qM�^W�N=�Җ&NG�sl9��q�޳�k���^QXsw�8tHoU&p�.x8Տ�W�^��ha�![�hs�ͱ����ń�&���uM/����ƀ�>˥Yl+�_q����Ȥ�y(FMʮ6�U�g_M�'~�%l��g�?rÝ�X�9/4�<�UO.�'So,��`y|�=�qj�L��FF�48���A�����WG��9��[���)�FV���z��R;:��৴�� R�ӓ�sHkh���;�l%1�?�+�~��)�N`h;-�Ϋ�;}���J��m�EK��z#Xi��0
BOv&#���w��zql������k{���t��B'��e�T�K��{�Ԝ5k=��.�\������k �P_ia�*q\��a�A���.ʯ:v}�rR�W��>iX+J�h�;چL��6SC�-�D�A�����ۈ� �'g�)P�f:�S��C땭�V�X���4Td�F*��^P�APu��u"�����A�A|��ڋ*=7�YJ�;��7����0�Ax2�����B󣕼�H[.3�5�K%�����w��HjI�y��NS���҉�z���+�u��^�8��|���-��8��|Q"D���թ�[��^ꔲC9��p��u����>IVY��'�M0������h�����rƢ)����ݮ�xJ�Y�����"5�Jv6�W�+Vls�_2Z�`J��8w[2$&�;�P�/l����J^_�Sd�ث�����9�,��l�x����������ƙ�H'�|b9s��~�5��4�p�,�=�BR�Ɲ�Y����{��eS fA���f��k��x�eR��$n���T�.eN� $��E�3p�o�<̑Lz��[�[���� �̿�$�P�ǣL�H�=Xzu��3r��+�XԃWA��t��4�4�*EXӾ+�y�yb��Ե�&ys��f>�Eq�.��C�]ʡ((6�?��s��*Y�S��> θm�,��c��<�"Ok��l�+�Q [x��0ԜnO��x���G�k��a�A��݇^|�W�E�}&�Q��x����ar
��i$�����Y�iƟE�
�
�=����ҩ)J��/��<�7�mJ�|O^��,��6M�;v1�$=��q=�#�Q�
���9�-},�DN�]8�sj��Q����]��r{�I@>����o�0J�@�����P�����;k���������B9�+�iӴ�XR�N%�u��	��;`%����*�=���r&(��Z�:�Re��6@Er��YL`~�߇P�N�:(1��2��L�?Z��
I�?��O&f�CM#�S�r,a�"�����`�9�ݛ&5��@Q
�{�*O��aޏ�n�3��˲�g�;��8<'\R�'X��(�� �%J�HĐp�/�;FC�	���Q�L|VAL�VF1�H*�cmvS�ڟ�f9ѹ�cʃ�`$��ک0��@l�����{Bp�S���F!�sB��WS%�������<=��,�AT�H�B	���W3�i�����6���f�9m���V���t�L�$F�g�>�x"���E�m� V;�I;�4|h,�ȇ�\�K4�Q�[�G��(?��ƴ��}��e�hu*������)0B������
G��
_�}��iB��O��N��WM}��v'
O�Ao3Ps�|���d8}�(�,WR�\��E����b+�1���C�dۙ6	K2���l�X�B�E}�1:%v�[�N�tF@E�$J���ģ�=�)������C͢�����ʐ�N]�P��B����&�0%y��=�Ȫ⭐	�>r�8zS˨��N9*�.�i�_�g��Lۿ�
@I��r�YG���*��	N#i���������{M���Y�+�aP�x����Z��t�r�9q�!q^�[=��A&N�J�������޵��k̓���Ѱs94�tJ�&�����8���W�}���
!��rs� ���p��ƴĄ"�M�ˎ�E����۰(��q��]����uM�]������'@���'���5��?�����_%�;/G4�<U�6s'�,��y�R������H(4z�H��Vƚ�ޥY/�ɬ��ݢ�uFX��Ӽ�DR�Vۢ������)�sʨ}�t���nˋ�_ۉ��O��p`j�-�H�ϵ�ڈ�o����i���z������KB�O�#����9��zsm�>B��u^X�aS:v�BQ"\�|��Tm��}�1�w7D�M�ӏdo��DT��	� dzi#	�*s����O�A(��.�6x�s����W6%�iC��j�;���	O C|V�D����V��
�r�؊'i�[Pɘ���C�`��X�W��dT�Қ�U�^Rp>P��7u��.�`�A�F�4G����wWW��=��U���y,}����x4}�ܚ�uS�r�T[0�gwW7%:�*�������I5k�D��������ٌ������JCu}"^DH��"Y��������X�"�J:���Y�]_�^,�2C�d�p"���F�G�Yz���ޚ�0�S����ڼ~䮅��aƤI��V�q�0��J�Ɏ���H\n�,BB����Jx8nW�m�V���_���b}9ؠ�w�!$�Z
�R��l�<��6�_��d���A���9n:���Rl0��AB3���a����c�'7<�95:?~��+����N��D+ ��
1���Jجei��� �`���i�ј�3�e���$��E�HڂkK�j�A�c\�zC�C9�E윔��g�ן�����1�p[ι!fz~�2�f屑G��~���]��`FR�K�}ĹK�p���z�ᴛ
y%����b�j��F�vL+���XC�w�z�ގ�A��_�V1�,��
 ��z�m��;�M�àeųp�2�����2����[���mx h2��d?D�>ٙ�G<��ȧ�k��+_����%S�˶-T|��u��G1��L]���bl����!Җ����$T.����"���E�\y��{&�!�f(m��8 r���'��������2p������^iv�`�+��gV�jM#�FZ�B��Nt��)- �T�����ub�>�CDrl��1&����rfD�-	G�U�0�U�b��'�DSt9����r��ݨ�%�̯�SLm&��@Lv�fJ��e��a �N�l-���97nw>{=�&Z���[��a�!�c�VWd��J����2��(��~G��p}�_�Xc�J��X���t.un=8A~"Ńp��'��N�Tla��l��۫�\=�\.RJ�l�[zo ��4k$��H�/��~��'{@�7$��E�X�4�a���iYkO�쪲�.޲=c�$Bdɴ�䶩G�F��~T�����
��6="��?�B�l^ˡ&̽WO~��ec���kл�C���� �yr��ڡ�P7:0}��܆k(���4����V�H!jĚɷǑ2��U�ťA�j(�Mw���v&2�0�{ #��2��%��D4��"R_������EA��^b��Vt�
uYڐ�	��$��1�" ;���|���"�G��FY��M���+?���� �38�4d���d˃���XP��/�@�QA�F�s3<���N���M�DO�ys��N��	@�Fle{��c1.9�/D2{'��~Ғ�{�H����+@�a�h����Ǜ{��q��ϛKu���Y��{�����S��^�9`�x}6T�g,��B���U�-h��<�ce3�KN���'��61Z����}u���+Ҝz�N�nH3ԨN`�������3�I�Q�� ���a{��j]u��ඩu�����1>�:�*�X��V�%�.u��9:m�hGpFIF���O+���jl܈�pI��d���֗<0�h]T�/N!4h{C��y���	�r��7*�<J��N[ΌG���j�]�����	k#�N�����0Ze��.��N�1�f{g2���;�m�+�au��7��1h��]5�5����;�|�������EX�`Y�o�K��'6J�F�+I{��[}��)!�.��fZ�s�3�صJi����!\C�$� 7��H����"�����·u����(!|�q�&������I>�U���Z&I�������{�Y]Ժ"ݲ/�4�.�F7Jh�s�&�,O���iHK�**D>�Ee�6 7/�2<N|��7�ȓ��H��,~�D�%��s���J������5��w�g�lVLJ�2��b��}�ܙ�\2��[���Ұ6���rc�������5��p���= 7����ň0�U9�}��}w�?`-�<OR��3|���`���j��芖��]��;� "�R��l�~d_N �-�s�ŭ����Z������R0d�!y%�3:�R��� �Q��(>QDH�w�gF��y,�پ��K��ʡ�S"�T���Gq��*����7�3�`���~��SW�r�D�ȥ;ĭd �-I6n��`�y,�\��H��Q�[麲����R-�#������[�9�A��� �@���j�8ŞG�ĝk�*����58�r�v�<EY�������rC_��P�[}��8!��{�2�Sn�W��n��a�&�:�!��2�-���\����n�j�S;%s�󝟗'���@�i������@x�>A��ޕ#���xu�Ȭ���Hn�Z�]�s�H"&_<͠Е�1Z\�gCѬfμo�,����"�hv���;4��}�F~�|\mT��u�o��dt,���g� U�I0p
Rz|��!� �	8��m����7 �Ix���՜����J�*#��]$�.%��������i҂0N)���Q#���1�~u�F 4w����S>���0��U�C�«�N!����	��k���X��fҚϚE��Z͙�X��劑����9V�ߘ�;9����3���t]��i')ʱ�hu���]�Tr���������mv�%�U_��>��˟OL����/��E�G��b����L>>�V3#���P�-o|�F�E��9ۀ9�[���/�-|�O֖e~�G�-�H��ϒ�q,�*�P����\����e�9<*�̻7b��6P�?1x#�;ۚ�̹!WnPQ��A����LK��m��4?�u�Di���y���T�2��@�JLuN��!zV޻�뽝Pަ��~�9X��^�r��O��j����[Qq��٣�t�J�������ז�a �v�/{?�<XZx޼�E	�4����0� K"p%��l����s�Z ��;����s͒�Nt��NĞ3�ç��(�=Zx���§l�9fnE��j�գ�-�7��/ӷ��_x8$���B����|�YlF=�%L����op_h��ğƊ��S?lmҏȐ[� �\Sv�ط��� �1?!A�h��t	�X[���\��T��lP��5���v��`h
��Z�a��^Ym���Sȣ���5��Y�%��A#,�_&Ȑh���#'0��OX�s�6a�2^= �,AJ�f�a�|�v'r�<��%*=���zî.W�j�v�d���`����.�m廞GY:��Þ1��Y��v���[w+�$�`�z����q(��OvSHK��m��x�ם�x�ބ��9Wk�v��b�0h�C�*��=�E���t�b�hvoX�	n�,�w��0�&�V*�]�9<U���b_D��q��}w�FJ|{����W6WQs'�r���A�)O�[�J���p��R� ?��?Q�g�>@#n(��
I+�@,�]Y���ɺ��)��:�8����>q+��İ��N};��<tyt~F�J8�y�]~��x)�fK�
^�s?|bG{��*A��ߌ��@��ߖ�`U�2�}��o}٤�Q�C�_/�hv�i�(ߣ$h�"e1� �p����+Xz�f�2�Q����~a��]�OFu���u<�����Ë��
�XΓ��o���jF�v�+�ZX�uw`"����A��"ږx{j���� �m�)ή�����!>����2Tb�@�������/�mD[r2� �?�a@>%q�G�������O�_H�g�l!���TH�5u5F�G��nL�`7�.���g��!����Dz�T�9��G֧��h�eN��YA�rɧ!�n�ft�R�\zmra��������n�Hߍ��%���'U�8�ϩ ��Za�O����y*�ⴗ��3�fU��os>a'23O&�m�/�O�E����AG��n�� �<2�]UФ/Rj4c�%e�;޳	��ʲ��<%�������'���O언fL����	�g@NJ�E���ZQ���~�[G��E^{"T������E�<pё����-h���5����V����q-���R�,	=�
U���ʤJI+ɥ��`����Ώ	8o��̗�#�F�J`���l��\^ӆ��פʫ�����S9i�����X g(�߼q�/2���J5Id�6IT}ֱ���*_6�tq�9���bC ����K�ĖL͹w��j���Kr�/�MX����!,�Kz'f��s#��X\�F�%�K�f�(�X*��}x ���I�Xo��0�D�K%����L��P���0���qH��_��k���ē�scrv_�j$-'����*�sQ�����ٹ�M��D�VD�h�Ǟ��}��f_���.�d� �"?Sq�~�a*���:�f�s�Gf�cKs��x8_ݗ������a��ӳ�x8UtX�ľ�ύ�c��;k����4ϸR-ܘ�=6*/$G��4��\�RbO�_b4^zw6g����UGC2-	s,9U����Zt����_�g��l�^�O��l�AG��_�tk���"ܤE��p�Z�H/��kA��
�a�S�g��:�$�L�d���lA��fg��e����(�P�:En�cb�S6�m#'T���݌��l�S%Zetʡm��6H��w#߭�f`L+F��7�&��a��C��쿘���ߺ8����1�v�p^!��gs�zA=��\m��J~x� ]��F��c��m湮�����ʋ��
�S����˔��SFy��+�f X�a�w�j���8A�^�9cco'��;��Ѕpm fW��L�?��6E2k��74��d����jm�>�2Lw�?.�3>\AG�8��SS�\H�_��
G�&���{T�l�ul]�G��L�!~�|�э!5���TQ-Q�~4o���\�0�)k�!dG*f�k�ԣr�?���X���E���+�5��C���!DE��é�J�Ji�����M��IWZեf{C���/-�l
�d'�]�XbXLCG���H���f(d��[����� �0�[gb8R~�G�@t��%�mX��E<ݨ`ͯ�줴��:ɾ]@Ol��r�J����sGa�A.Nk��-;����[wA�቉�Eν��[��ڤ��c{�d�E00vd�5��(Q�$G܄7p�F��w�c����[W�4i�t1d=�5~��p���V��a���ʻP����=&߸� �me7u�R���w�Tʃ�/ W��a]?{ޠ$�ĒEU�����Qi��J����� X0$0�f�79��!��E�~����R���6 *��b�YB!q˄�� ��~3 �c��ސ�u�͎��>y�s˽isPz�� ��܉L� S����wc�˵�j�����P2�$*Xw�s��j� w�Dbv�� � f��2?N��(sD�����7�݈�q\������џ|V �Y=���ǒG��1<F:4I�G���;mG�Y$�鞲�+bVz��:3��o4�;x�'�ˆy������@�v��ɳ3����!�{LDR����cNzX�@��e����.1q���5�{M91e��UhS�k���M���D+�h��ƚj�����ج<i�K8e��|2������5�N9�7�x�$��xz�����F;��}��Z�evr�N~���*4���0�ՠ����'j��#����zN�,3��`���6�V��I�e��/L ���F⬊/�uG��l����ʹ�:���W���$��(�u^��:0�5G��FbJ�O漐В�� �g�]KR=}����\�a�}���Ocf�TЏk�6���p��)�W�uC\Ƣ��X���������;m)@ng�:���Xz6��A��Do�������,�� s�%M}ű�}}2�X�u�fU��3j����X�|�>)5QuI��E>��|j���K�����ӢzMF�*#֮�\���8�{>jm9�Al_|�-J���K�f�ʷ\�P��@d	*��H�y�5@sRʣ��-��i�v�Vrz�5#�h�gRK�������i�c ���r��k
��l:0������0$�<O�RxU��G�k�8�S�H�-f!|K �E�/���hx�v��]�L
m�itE?�<�����E	-
5�2�n�r�y�{��Ҍg�7*���̡��ϯ�,��BMC,��+v$�4q�Yz��_;�z}�T5,�ѭxs�ô���!5�|��[���2�>��|˿d�J�A�CRԠ����k�khC+���Y�j�
��X1�{�d��*X�ق%I4��ӑ�����㠯�z4�� �rvb8Ѫ��:@a�*���"�r_к��~?,��jڬ��P:x�����L2r���<�ZO����6�� 5��q��`�A���a`m�"Ovz�L��9���&�����{�˝�O,�&aϰ(��'73�E�;ؠ;��<w ��w�j�xҷ �Gx5�H�����;�.�`���L̾e���V��sHzm�c����9Q5a��^�
't�5��<��2�)���q�p,:�ӄ�K|o�,%Sd�@�)�&L�	���k�	1�A�x��at��֊�Z��)����J���em�(�V�lJ��h��t��d���r��򾤽��V���;�,�h|��o[��
�Q����� (� ��81�4'�}4i�������"vBل��g�e
����Z�W}�Y�B��O�7JNX	W�Z��*�
���o�8�Mo!�V-�di�@�x(iW���\���W��c`1K C�f�d+�C	���W��ռ끾����O1��]v�7�X8��@���tί�գ��o�yv4�9��2��R�	%!�-#>];��kT���&K���Ϳ=�㱪2��	�b�r���S!�垻R�~����B��mx��4\@�-�r�W|�+���ܻ#�0��n)��_���|�F{�PC�����Z�9����q�d^iL�=��&&��҇Ed-�d�C�kʸ�0�Gs�Nt�|l&�'J�8�s�W4�S����!-.�s�j��;%���ބU*3MA�n�M`J����+a����q� ڭcn�K6CM�v��/ִ_-A���'٤b�����
��e��dkd+-ua5�w���V�'Ys��D��G�Q�}��Y����wO����n^��\��U�&AR����q2^��_�9�cn�FS�t	��6��7�:�f�li"����D����t��"s���N�*���Rq�A��.-4�9����{W7K9i;)����K;}������Ce�D�ek�ɑ�(n�O�'� �P*\��V>CN���b����T�ڹ^�^�|?P�Zu%���/��A��&�$΋��x�&�~\��o��=���#�x��1��țv=��{[q9S؍�%����8�*�Z�}I���E��1Pd�N��:���}x���8u�T�^�%�����F�.e�L1-"G/I�f>E�h�^��C���p����Ȳ����Y�i(� a0x�}��b��������{鸷oDݱ��JI`��=�)��-a����J�eW>��Vo�_��h�#����wި�$	�Ó �lGY(��;_"9�dq�B��.`���9�[.�X*l��r����_z��ŚoƼ9'8�d9V�%~ ���~�s$" �<Z����ܦ��ͨ���� 	���Y�!�F��eu"�$�E����.�g ��tE�	�������z�ׯ[*���C�c⸿5U��S�{��H�~Tz$�߶���+&=�&����+=�{��k�M�XV�\ �bӈz�X�yv��f�7�E4 �.�,$��(���"悚rs;���{I��|[�^.�em�@k�_9-ꈠ�)���{2�� ��ỳ�r� �BUM:k���ڈFsb�9�̂�y�����H�~�nUpEz~P�'���&�.�/�)��û���_G��N�C�(��<v�] ,9/E'�4�lǁ1{��'W	�>ʽnb<�����K�R���%r������2	1U�NUX��Z�rZ�9���@�!�c�w� {m�	�xg
��*��H��g㳩rh3=�5�	���ŽB?�|�'�5�C�е�56�K�nJ+O~��M���t핎lpɗ9��O��JK	����\	����"D�5����z�~���T]��C.�('�9qGVI2||�7v7I/�6t�a�.����_��!q�W����jCꆆ8�K�qJLX��z���:���u/0�XZ�����K��]�Q!��q�\A��%�Ef���X��}C|��+�IRaJ�ֱl��I%��~��Z%JT�G{4�����
ñf�O�?�@���Q&����� �[>K�#��tP���ouB�<g9�W���eZ ��Qf�Ye�e�6I��lx��z��{0�*Ofŉ���&����ߞe�S�*k0i7,dU6�w?{�E�����Wx�!�H�%9]L��m�c3?�N�D�-��ͤ�Y�E���&�L?wB�+���h��'=�Z�p��j^r���I�j�@��~��F��>02��p�C^I� �� w� �9�9�/�xh}uE�P��?��Z	��< �%�H�����oZ��(;P�8�}�U.'�cӞ=ଧ,(�0	ZB�Z����l���ڴ4�խ�<��d��Q��J�<8mH�R5,B�<��FDNY *F���%����Z�oz́��y�R�S	�ҙ�J[*\��l�[1��,U !��?��ThN�	��L[����Yƭ�WlZ5�5�Bv,@�hԼ�d���Qg�Y�%n�	���25湷��S��W���N����w�]�'�1ԙ)s:|��)�=*���x��saNN�����Ϣʪ�Y'�>��;��xҤ����v��)�ҏm�FK.'���h��:波��V����vu$@['=�n;���}�ЕX�q2��ÙE�H�U��6�Ԃ�N����E��,���b���ͽ*���ɲ���bz@lo"v�n�w�7��h!*��y��<�8��� 6��dХZ�w�|��6��J�aw�Q���Jل�^()Y�,�����ђ�(�?��0Qm���#8oȢ�*L+2��,Z��޸*e����+�$�68M"����p+�Z��3Y}^A<���|Faq8�)]D��)�^��MsIe����ʴ��שQ��J[1���2`ߣ�����y��$C��2eDsh����1�h1�D/p�����zT*S���㑝�Y~�Y]�,�F�⪧Ӝ�a�.�����w�]
����봦�@��Flg+�8AXY~.w�t�t�A댖�l��, ��ˤ#��mӅ�#�J�����	,�2������W�n�9�Nm�aJ2_��?�"3>/KGR׌�}0�Oe__RlD�����T�u?�[GGI�L3�������q/�!�C����T�N�Q����4���\�#��|l�!s�f�2e�&��rk�~�&+��E���o̓��R���p�4I��|�o��}�9�@FiM�4X����X�>V 2��-v%.������!NbK��C�����b�y�����~��3u�0�x�b+uǚ�tO���}�a6�{_����)���A@���%WwJ��j��&�avcN���-��-� �w��̉<��Ѕ�[Ff�w�c��Sd]�#����R('ZG��p��d�^c�Bf���&�'$�t�}�=NT�~�:`p!��R��fa�7�ʮN��j�+=�%�>��$�H���d�
R��v
@/S�9��6{^�$!G�E(��J����i�bͨB����c��;�$���
������zu~�����_����6p��՘�B�7˷��̓��~&*�c����q�v�؊_Byȭ���ݗP��A���7o��Y,�
�؀���jڌ
ɍ��2������&N�j�o�w'�|v|/�FE �J222!��{��DJZ���w��P�ĭD�`󣠄f�ђ�#S�Y�	Yޤ����1RQ�Y���u��G�yY��Ԟől+��Ī���31�4:�3����ٓD�n5����@r��᜿�3R*��Ѫ�n+�D�m��HJN���@P�=e[F��#8�1���W�{[�����h)���|�� ��w��hW��]�P��e����KK�������S�E��C<9�ߊxӨ\�}�ǂv��A������R�e	KrNqґ�}}��L���|�D�=�˛9�P�N}Z	3*-`���@���~�I�B�#�� �)V�9��ݾ�u��U�7���͇�:ݤt��y�7�{D;uK�:C
�Gy�F5nO[��%����g3�G�2�\��1}�6mO��?Tc�(�)�	���){�3��N�\9��h��5�ͧ���={VV�)2��nz���#�z	��t��|H�Ў�����ș�l�8�w��C��-�eW}�� Uu�����݃b]�?�5$Hh�s7A��j���K�ݮ_6������*��Rr�*В8d2�j��ϔ�|��&@r�~���9�⷏l����	RgH$jǑ�ԊR���Ġ!�i��/V�0�5���v������u9�|�`cs7�E�k=�il͏�� Ipa0יUO#�~x��)��pkx����\� ��|�3�E��/���1x^M��0V�
�B�ik��/����E���
H���1��:��X��w���7}/��E���ɳ,n,Mq�p�$ �q��)��{��� |�g�,x�Fр���|1�4�ֆ��V��L�>�¹�2G�J�7�vf��3����O k��"���=�}�c�o���N)�7ʫX5n%<[��&�2�>�[��F������r��q�=�:3˳}�5�9�rr�e.�~�B���q1߯:k<ן�&�L�'b�����=��bT��WX�&�[�S��5�a&v"bEC��h�9�ݼ&��#�k�оOE�a�l���Y�3b�̲��; c�<
$`�j���� ��H��H����R�u;��^��5�Ǩ�L��D�/V��'H�Pm��J�"ff9�������]��'v���L��������Wp������������Sw?��T�E��`����A�����!-�Є���{��vlۡYXA��2m���V�1��q�'��$觛k�GC�9a��P��V~�;L3�h/Ä�������Qǲ�ʂ�("96�ô�Щ}����[�\L���4�B�(���
�5V�C%}�0�B�O[��N+GxW�RWؽ	J
���o�'� I�i=�d���K�XW�)�\��2�JQ���1������d��i	n�������O����� N�1=�8v�B�I����� �v����<ˁ�,Y��,S"�B���<)����s].��`����&^I<��=���e�	��Or� Sn?)�Q�|���	�"$��|��?�@,~rͺl�~q����P#̒�̋�������T6��Q�n��P������*Z����5TXq�7[^�\�=��	&�|��k0��Ui�k�k����[Ts��t-vz&���N�vU<yA���M-`��NHQ@ko�eֹd���1?O{�`]�{Vf/?�G�#5��לޛ���RE9h�Lj��U��r¬J��K�'�
�L]���} ��9A��x�����D��o��\���i��-�peD� N�x�w�����N�_*��J�����#2N�3%��`'�yP���hI\����� ՞��ԟ��n�u)pa�:җ�����h:��.�%�u`��v��ul%V:�/G!V?F��O��s�`����Ygy�`�D���R\b�}H:Oq¥T�mV��G���)�ҡ�}��\TQ�������c�w�Q2�)��[n5���>/�z��O� )�k�i��l���/������ ��@���CX�U���=�����+Z��5�?l��Y�|j{j7�KD��	<7�H�����4�G�b8��$j�j�Ϗ�|���ę�B�z��jH_�Ĳ@	�1H=9�C7R�L ĻVUi7��V��5��HS�>�H���3�7��c�9>��?{k^�l~�/����02"�O�<3x��p58�k���!�Z��{|�gTE���o��xyC۝�<
{+�iBo��}C���E�Y
l���)?�J͠M�~�y�7x����N�����,��kM�f�ԯ�$[�q���� U��"V,����� F��fНoS����Qz��;l>���M�3Jm�&�Q���n�!�b��k��.��Ϸ8�&���Ё�Y��
aXp�z%����!�˭�W���(br��j�xC4:�ؒxO�����r-�Z7�y~��!�xD)l0Z:�˟в:L@3W�o������e񇭘I�au���00�an\�"G֔ڡ�90:&���^M��Y�Ozg{a�����3}�����;���<E����&���� ����FH�����޷;�/��.���b�3LN#�7cVd��HOm�(��R9��A�s�X��X����_���ai���bp�Gɢa���ʹQS2����$��)���w��^dA2`���:��+�Պ�����'y��v���w+m�DV����ɂ)�߶�����������4VB�;G�Sh�Q��=Wְ)ewQBgl���$(]���]*;��J}����@v�w�i�p4�B��ǡ5�:
%Gl먈�}��B�Ov�|N���W��x��ޞ
-5�o�7e[Xһ$8�d�bЅ��W�n�\��:���T� �j1Y��a_d���	�v��ezCՊ�(� 3�`1��v�,����Bl���k�7<Ї������!�&�2o�����]ɴR["����&pW��==���@ �	�ܱrx��SiF?嬊S�L=��=+�Z����)@g�mrh�K�yC����#�Ϛ̦���b0�ٛ^�t*	?P�����
�Z�ƪ�P/qm�	^wN=���&,Q�����w�ӽgk��%�~HOs�~th��&������8��xW.���!{�s����	E�ŤᄣuxMOP]����2�y�l
9�q�.$�;+����M�Yw7�Zu���'�Z��E���?��J�5#f�Y^�4�O�Uo��'sʔ,�u&y�W����8��f��4X���aA���A�w�鎧���{�5nFv4-Ӛ�R[�L� C������v]sh���%a�����_lH�?U^�ItT`�Z�-���[���������e�&�zC3��pBo�h#:$���"4z�Ұ�K���0���� B/jH�NT�����U>���e]�|�5�G��O� Pi�>)*�kY��T�A�K�.��d�x���QW��ix�\��"�;��>����CڈSD��Ƙ�ۨ� 
�'�"�P���s+�C*L��=�2������ePE��)���}����3���G������E��-!��`C?��M�j"h܈�݁���n��M�6재�U�H�!{��Y<w{��$�Ȁ8�#��v!�6`�j�H	D�g��&����1իփ���(��Մx���]d]s4ƞ����d����"��������+>ˋ`�]�K"�i�/�ʹ.�_�7Z�&������O����ym��kDN;�e��7?��<)k���ȣҧXMx�<U�D�s ��N��T������d���Z�w%RV\1��B�;b�!���/�l!5�#���異Fς����d����E�p�o=00���Řl��\S�-f���/�O���K6R���3���+*���b��ᅖ����۸� 21,R��ݷ|��do�U���=������j줿r��{0tmy5f�:ǉ���9Q���>&�T���gV�Ly<Y����K�ʱR*S&�JT��W�z�:J���v7݊�`��uSg�@�TTN�K�d&�5-.�n�0F`��7�lw(�X��Q��$��L���A&-����jQ�k�D�Q-X��3�P��zj�!��ԂkԱu�5"�L����R�7�	��|xo�N��AV�Kg�����Jow\�~;}J��O�VT k�����z)���x\�o���O�d÷�9V�SzY)�;�n�4� �|z�d�����Ҷ-�[����6���u��n�9�5s�N��{�U�]�Iv� ���=5�|�#7���;j��K	2��K�,�ʐ¯z�ڮ6���Ga�8!��jaBtϑ��|'�X}���[���{���iʼF�	z��H!� ����R���}�Xi9nmV�[�5s��ݭ��q�$��ֹ(�cPfy��kZ�rl����spOw0tX'O`;�x��e7�'k3=O�@/�}{�|��EF�0��^Tx;����z
�ԓi�@�Ҍ�	�:EY�
�.��%�+������+����7z����#�,K��M�����$ݜ%q�^����b����#,U����O �v��u�`���SZ����>,�a��fJo��ӓ,���|�$+k����!����5�L&Ɂ�L��T]�X�dO%�)�#1���{9�3Tq��Q�*�r����`�:��Gz�D���
r��b�o�~�Cg���%��:�$K���L��q�1���M������Q���Dٰ��2z4a��"�ߔ���92��&Ձ;��!��)O|�laz*�r3?�{���e;=��<�;���+��P ?a�]XHd4:���;�N����ڍ$��L>��'~V�KH��m��?��9��q�+��Z�S�j��I ���O��c ��S�p|��#���޴W5xS����yqa����8(��Y� A�=����u�m�	���S��=�Am>��VG��(��ġ4a7���I�Z�V�n��OV�cl;I<�h��އ�92��OQD�J���(�Kc���f}V}��Ű9���r��B)�G����
�$몦�}!�BBT��O8e�N���W���z�6
�<Ao�7a�XN��@�d�{M��OW��\@+���T��_1�9,��ɻd{}`	�h���?�w���~��1�2Sv#��u����0�ĩ�^Y@�9�C��O��i���_�(jfY&_�}N<]�D�]���;�&� ���=?K����F	>ޗr:�iSk����4M��/��O8�\$��.֒@���r*���{��R�#	$��h�G�d�I���Ė9�˒DP��L�8��Z.}"���qo9I^��6=K~&�h����_���U�fkm�ꀉvs��t�7�&R�T���87-�W��րJ߁!}%�s:L���0x�fhD��IGM������h~��{��Lޤq4|���(\����M,�I�2|7����T'�!��ǺH�Պ�?�B��w�c���P4� GUqn/'��H,]�Wy^����WF� ��G4f�c��:���Z͎i�N�}J3U�F����\��R]~��BpS܀�Ɏ��/sj�'�$�{��!��A�ۋ��`
��-����]��V�M���'�(YOz�� ٚ	�B1c�#<&��d'z]��%^�������AB�ը��T; �q}����zA��O�����a]� �Zi�Č*�-��sA�B.,�����T�EW֌�i����
�g;�Z(����C��D�"����۪�.b��'	58Pi��u�CM,���#�m�KT�z4��^��PW�uD���.̸Aq&H��#�LҎ�����N��P��D/����x����|_;9��&[�u��%�Z��7-A�91_I�~��-�Ѱ풭��yp�������u�<^��a��J�я��$���ܣ"fB��e�����^�C[,�p޼�svθ ksY,�~&:0WSw���'�L��1���D���O��4?JH�멷r������Ik����J��W}ѲV�Ղ_�����1xԔw}�'$�����l�@D�6��_!�dP�K�����4)u9v����lТ%�Y��^��ݤ��{��'�#.9�~-��Ŋ�Q���J���{K��L��M�k H��.5� R6�%��e4~�$'�Fd<.J� &E͟޲ѿxn�zk��[�,��;�����tG_�r
��UH��z����U!�mr+���eK��+�z,����Z�X�o�۔b2��ԗ��y�Z�f���E�.��f��G��?j�፪szp��.T�{H '|:f.��'�@�}m_����(�)��8{1Ox d�z�?����iU��o�9�s��p�9޻���y�-�^r��}U��K��'�R�&ǂ�/����Z⾈�G�����(����<�[�]?/X/D��4ͳ���S��%�p	[��<�'��~��Q|���ڪ�b_����p	�2�N���ۙZ;�`��WT� ��6H	{�*��SF�R����1��q㲽�hю5�/�%����b�����t�T��4���*��J�_3+���ɂg`����-���U�8��.��J
�u�V�$\�Ɖ��k8�t�뜦�}���3>T�+�(�_]q�~�2w�פv��INf)6sV@��}G�_ ��qE����ԫC)��·��K�P�L7���9���|-�us/}FIX^<H�%XK�=��0O���[X\��%'g�f�yX�=�}bU�(+I1���ꛓ.�!%W��a���������������xQ����"Ľ�=c܊o�7-� �&6l
X�Q���H"��A�A#{��R�c��}�f	����J�)��`�(�F*�P��d�O0w��)���(P?6�.c�Ȭ��_�!�q��t�n�C�Ԡ�/=1Kc	/L����_V����77/�	�X�n����aK��Ш��
�\X"7%���ffd,XLh�}��i��iI����&��%�{N��J�r̥�7/��q<Q��'��=�����5�DcT6Z'w-�gd������QU�N�m�[�����5��U�|��}v��f��rǐx���!�c����*����R�U�f%�eK�x�0d�� `��X:aX͍�}�r87<�z�� �	�t�����ר��R�0�ZHEo=4��<@p^�n�$4����g��|��9�/�o<
�tͮD�׮� 6^,I1K�
=`|�L�!�H/����1�%֪^��⏸ȿ�b�2\���# ���?�3�U���o0��6"K�Pʃ��O#[Z%�����q&��^P�{=�)o&E�*��탙v-�LJ�kD���7�Esp��taϻ&�2a��8N�BW{#�!��!4:�s����O�ŽU����aM�Ct���??ӥ2�3�0jq�!&�T}��҄�MC����X]8.~'w�>�e�,FN?�h쎨Ҏ�4_�U(��'LT�,�:�y������]K��.�4�e���日p�
��i3���lL�F�6v�3;Rv���^����y���s��͠+�Q� ���F҉��#�"Y�`�ڢ-	Q��Fĵm?#�����A0��0z����B�!V#s�"���z
��7ǆ�$���z�2�BH�d�S��T$[�+3��n���M�U�*�
�~�� ;�'i���*
{��hSxA{.���@���x�W�i�÷���;�!��`(<C�Z�D����D��=y ' aP@�W�,OUC�*�o�x��YOT�f��d�^�UP.�>u�,����A�Ȫ+C����-��+]������:X�)�5xK}��ӝ�L�ܼ)�9[������%�~�Ρl��8�I,u��*���^��nFP�?�Sa/�$��uˍ^U��R�Ѧ$�ãb�"���w+�tԢ^#�(C�{<p6��joJ���nY�>G��Z0����	�U⠅HS��;�ͷ�݇�J�̩.��?���'d��~J��WT��VEv�_+e
�yg_��ww��i$��l��vl]"��l_�Jd��[����k�W9%H ���1l�V�������L��Z�Ҟ�'�9�.~vI�����IG!�V [�3��LЫ�D��c��Dw q-����������:e�X$^Y��]��.�s� �j	E�#/�h���ۆz�~8[��P혩���9�K���)U�ǜ wH�cz:+ߌ����+|̙�<����&��uR�Mt�c$�X,�ȡ�P�b)̡�n�yL3�f7äE���.�菶��">����sQu����{ߖ�|��o.�<�C95@��_�\i��k)j�{Ȍ� ۂ͖c��k9U�=�0�\C��Tb��y����O�TLSUN��k�'��&~w5/~���&��V�G�u6��V˓~�<��]��j/���4D9d�&���\aX	0�:�v�<����pb��Uh�h�薹���ήc	��N�U��p1Z�3J�x�f�wDJ��J�{C��HE�Id���^"��I�h��5�������D��o��K���g��ˇp�U�J0�+%�ƽ�Ă^�=�����B}M��K��"EJa����\�/����ϤK�ŢQ�Μ���.�Y��(�ȡq��2nGۤM�oI�]6
��/��L�_WD=q\F��n2C sF�n��K���L��u��R�$����/t�iX5�|���$K;O�Ч�n��.\�b%>l�f�PKX���}����vI��Ȳ�$��e�%1���XF��7��v������ʇ����t7��1�c�@�{��-����<��1,Q��x�\�����8��e^Q�	�u����}uw�f`���Ou��a����ܫ��:*[����_�T<df>K�[�xy���X=���a�����j�86dY���߇؍���gI��z�����R�Z����0WV��)��S�R�.�_�-�^�g�<?��1/H�@N-V,z���%��t�]�K�g׬@lǤN�d�����A�2�s�t�e/~���j�^7�[Y�/��,A׏���~o"�������k�H��c���=�� �a(t9Y��Ĉn�̠4"`m$�*,H��Xq6Z�G(��rMp����R@��fYc6������>Jǰ8X�/#��c�OP��M��8�V�A��2D3�X@�)�!�G~]�`�8�}�H!��+`~�!��:(j�7��b`�ben��MB�6�Sŗ�)x��Ҩ�T��{N����v��>m ��q6;'�kH��g���;��1�,e��56�H��_�d���j]b��� ΐi������"�3%�[�A��G���N]��T"��/H�E.��z7u�������O�0��qa�hD���e�#�7Z3<��������Y[��7�<DK����Q��W�P���������\VW>��/cb��>����3��'��Մ���EE�}�c�r̴���V�`%Yp�.v=%�ؚ��3&�����h]���j�#�!�R��h3�΄��J��T��O���n���[�F�Vڵ�?x�c�Y�Һ>�[P<�\>##a�y �:t?�kqhOu	�[��G�K��T�l��B5��pv4�h�,ۍ�$9���#YX"���Yd�5�f���G� �Ɛ���S����[�'�4��Z�0s��{==KQ����Q�!aϸ�!��鐱0��@O��b��^���Y�UeGvB6
�s[Y�A�.���iƎ:h��)�`�D�zv�p [���/����vЖ�qS���.�H6g�[t��#�w��~H��`������b<D`�.��*B̈j����U,b[k�o#�bn�u8w [��*j ��<`<E�͜b��\��7R wEV|�u�B[��Q~��+믄���)z�o���&�ޝ)�?<��Q�x���I#9IN��D�+s,�Δ�9Z�x!���v �(�8Nm ��s6+j0��6}�A�<�F�DFB1k8���].B��U�=)uMi�U"is�ɕR~zʕ��ת~��k(�!\>`@=�e\��F)��/C����3���2�.��s�1&��pR4�����z5�����Ñ��;~��x]�g	Fi��t4��":��|ۗ�xqY
�t��,9�����F�4+���X;�w�r��u��A�����Kc	��!\f�Ĵ�m�st�C����*�z2߹��+�g��57��M&mO�2@�?���>P~G�na�ޝ���ж_�G��lx����TMu`N�G��L���y8A��!��w⯶xT������~]��\)ќ�. V�1-�Xv��b3���g_�~"��z��g��,Á�O�� �׹���,�����]6�P��厾�&N�,�=�0۪Um	q�jr͠�S^{�Az	��1�6�������@��r�D�n9߄���#���{��� ������M.^-�P������Z�r��%F�q�g�^���=~��&�����������*k��J��zs��`tR�&����8���W7��]Q�!�ٲs�9���c��������M�E�P���{S.���D�qg��ڐOû��5M�l4�J���	'����]6�h�-?�~���u����4��)U�ke'�_>,��y���e�O���4-
��֬��n�,	�����p���F��E�o?�R�>�b�ܳi�H��s]�B�g�g�����4�}��
?�^�K`=A�-E�m�PL��������:>��bFzX����;jB�ۇ#/���,N-z�pχ񯃆��o���5I��B�1ۧ�9T`�7�Ї��*�M�`
��͗��܉���� ��ti��*�����5A;��.�bK�����W��Giqo���U;�ں��C�E�D�`���۝/:�IF'�T�P|���C �+Ԏ� �/TyT��	^���Pjn�u�����^A�j��g�r�?��JN�t#�-X��ex���M���e"w[�C�*��%M|��
}n�l{6Ih̈�����`��������`	�u�	P^Ck'��0���@S����N"�頫8K��0&^_lCNUypr%j�&�$�3ӏY����Q�0�&%�+���	�����M��	���Cb�Jы���{{���4�ׇ�J���W���VƠ_g���5���kwp��$�&{å�Ul��捩a�_�!d�);�K�f�'^�9aI�j��l�Tа�1����&���'ʛx9(��~2n��Z�����^�(��i�n�؟��� #w [�1��1o�܀�Xؔe�	�$-� �.��r �E@_첤m>���z��[�m}�ԚV�uR"���2����O	Hԧ;zv��H�W��t+8���x.��uZ��M ��	�����X�6I�.:Fb��Ԫ��yc�fs��EF�.J���r��݇����s����{:W|m�F.6�M���@=i�_Ke���4�)&0{�b �����⇌��Uj��
h��ߔ��/)�KyǓ4��2���KUB'��l�'�$�&:��/��ɰ��Q,G����˓:�<Ȑm]�(/TT4 4ׁbڃ��t	l����nC<���,m�$e֭$����
��Dl	M NgJ"۬�1Z�G��c��37s�ɔ{����J�� ��ؑ2���thE�
5NI,�zG+�]j��\���e��sZ�o�]@�JUrd+���͉�λ�Ʒ�����K�a	�J���I��\�l�������
�^f�PIR�fГ��(�J�q��2*(+����I��(6Fs���_¹q�{��K�C<�4�*�GK�.Ljc`��G��o��Ȓ�/0�{Xq���~�Kw>6�cj��9݉\�X;%z�|f�%X�PH}��J��KjId�)�(O3�!��%m,���� ��2�����؀O���X:�r�[�W�c����-{�{���&=��Q9���ţ�6����O�>p��op�׎D}1>Lf�*����ٝ�\��;6d*�`�7;Q���f@X�KP�Ox����5�XX�aS����A�8�م�>ě�d�O���#���A�ՄR*���Gli���%�*�R�_��g^׊�g�e���u
��,�
���5�tV	��4g��l�W�Ln��IAĻs/��t(.�:P��}_�_�Η�</t/�A�2�~�}�J��st5!)�'��#f(���-����Ը�(��[ɗ�������ȋm`�,ԍ���n�6� (��_M�3S������a�c���W��Y����������ϟf�P|���%�ޔ�'h3����e��:Ϝ��9�#!��Y`:�����jـ�u��nJ~�M�V6��L_���'�{����?*��z�k���6w�a�MH�o�gO@+�wpi1Lܟ����_ך՛黔|�]JGc�x�Ԑ����Z��"W����B��˂��]��]"��/��,.p�57�����E��*t.O�V��PNf���D�9ep�w7�,�<`���#Ț{/Y���D��2�r�|�+0ֵ
��q)��
`NԌV���C�b|���C)D죮ў:�2��������9O���\-�pO�뜴6p=�=Gs�����o�pKt���t�gj����J��fR�h3��t�h<�^�������d]I�20K i��R�w�s��dF�y�׬�P��L�W��H|�����&�|0k�y�Z:~���^=�Q7F�>}3o�w�*�gM�*yr����K�h_�(P�S}{�T
H:n���1+˷*7���`V^���S��؋�ޥbJdk�-��n���`T���b�yQ��ٸכ�0�-����������ȿE$�ӈ� X�����u̫7�k�4YQ5�܄��K��Y�$������Y��x����T�kt�>(Z�yn幋�uS�H9�&h����Ҟ2E �&/���pSn�SBㅀ�q�^���m�i	 ^�O�M@J������6�

��?���S'���nlZ)o���(D"Mf�Ԍ��m�QZ#�}g��f�eo�?����"�凔�4�:��_�|g��U��o"��ts��=ܵ \8�Ij�
�	:|]��!�vp���PA��A71|I��-��d�h"���CL#@�$'��$e4��f��ue���0�!b�}��#Q䱨x��u�`�4~R��Ȩ>b5�0�X<U,ο��!���0]k$��ʏ%�-���AҒ���b�V�Xy}��X���R���q; t �B�����&��Y_q)�pch|cG�D�	r�~Q�ͬ�$�>vf�U��b>����
�����|�u�w��κd��:Ҍ��!>���#�U�Ps2EoCUa��#b9b����A����T��V�eeЛ��9�����@'*l�ՉW(��YW���Je�:�*��27	fV6���?������i���Wugo||"�b��L��m�?	�D����:�� �!����L�=�S��"︽�L��ʷ�~���^�����.j:���ҹ��������PѸ�x��]if T�	���I�P�x%�GE0-��Aͺ�L�U� ��%5g-�5t��M�$ZGߔ;%9��>���v��@o���+�I��(aO�Z��Կ�ccl���5D˴�	�*pP��쉬vݿ����8�-�B�^��#��Y���F��]%��3k�ow.;�~t��QaSS汅����6m��F���I��]z�7�!1�)�)��!�s6�!�������v�ַ����}`��C�1���f�U��D�C<����z��7�����Yg�1�x�p�kT���z����~�
��~�|�].�F5ͧ��w��f��ȡ�D�
<�W���-����F�<�+�0�X�sdw�h�A�WAX�Q�y����������Nm`���P!֠���vov2��
�w�������&�im��2�Q>?n��>��G_E%�*N�����_?;5�ɢ���qT�΁u��GTtpL�[w�E�(�^��!u-h��8vT��h��{���Ŝ���p�fiuH!���f++���Yr�i�!˩�C��܋��ud�����a��X�܈b��߀��M�M�����8�����y�-�	�����"�b���C���Ո�����ɧ������5�@Q�09�obx�Ǉ Qt�77���.(���X�_��֟9	�3@��!���.J���ȕ�a�_N�N-{��.0w�N>�ɕ3����[R:��h�c��d
��p�v�ucN(���G�up���ac����t+@tqn�=�b�~%�p�����1��a4fN��R�W$=fq�1������Q���D������j/@�ܡ/�{C�!$�&7E�a$W�=�Ui<a֨/]�_)��@�G$pqi�w���̱U�ɿ�~7ߏ�	#��^�C6@Ļâr�Ba����-h�@Cv~s"jc�ͦ��F�F���W��y5�|��DP���`6���֡�@ֲ�7��M� �`j�f�:Y�2Ϧ.�����j+[w��]v限S�y ��2.�h}�D�P��%@��k���+2 ������~�@/�Y}=yJ����1|��^�R���%��}�G�DYdj��H+���M��3>�'4�u.��(��C6������@?��	��3_�:�H����D��3YN��@��e�A��0��1��z�8�{H�3q��ҕB	߫��ލe���h�_��� u��|;�Kx����>�L�(	�Y�&9�x����
��EIt��(��g>�_��e��xN��l�j>
�ق};&�ĳ���'�����6N�.93eW`Y.
��Ũ��UINA�0�� G���T�ʹ�u[A���l�\N,��v�:�{C���(Ʀ�h�5u��:pQ�Gӥ�F�4LO&���0�F��g	h����:V�\�CM}:�O���TJ��v�O�ջ)���O�\�@��Q��CP�T�ζ)wC�_)��n�����4�zv����A����Q���$�&3��el�^��hQrߩ��*�U§ist�)y��!�5��������j�K�Lm�;cB��'��jE2�&��7��8v�jQ�\ρ��|�md��K��~�����6{~	jH�
�uR>R
��m6\i)a�V��5c9*2���0�֩�"c@�:��kJ�lz���**y0d�dOP�lx�հ   �  z  �  %  �*  �6  NB  �M  �Y  �d  _o  ww  ��  ٍ  3�  ��  �  )�  l�  ��  �  ^�  ��  ��  e�  ��  9�  ��  ��  �  ��  V   � �  �* �5 D �N �V ] Vc �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����O��=���Y�+�F���eIq���JK\�<1!( )�%p@�ř'#�ܙ�TW�'w|��I�E�J�����{�)"�/�F��B�IX��-Iӯ�7�ة5�Jba�u�	�'XJXw�
P��-��I[� �l��
��� ��{�*\">d 0� o9f�:�"O8����e����!(�"R �R"O
=�kZ�t�:f�C(kA@B2"O���1aT�l��yj'&�8l��u��"O�"3�	K�,@A�˽\u���%�'�剁IQ,h�A� 
��T@* �L���'!`5MV�+�z�i�ݕ.G�P"��HO���Q��cD������z-�"O�܂���u�0"
]�8�Z���	��0<��	XX���0��r;�}k�c�F�<	E/�����b��B���t��E�<��NʭZ� �被�������j�<�R�)����ɀr����F�e�<IcY�n��,��%�T$IUF�M�<QCK�@�������Ip��EB�<�e'��%�!A�*Q�)�THX�@�<Y�!]2yΈ��� �I/�P����p�<٤H�<��y��фk���Bn�<�1�D|L��a��=�m0�yB�E�`+X����I��A��y���':�kQ��h����y�+�F,|��Z�0�i���Z��yRE�!���h2ԋ+
����y"��;(?�h��c�!T��	i���yB�N4�M(���M��9�����M��'7��b)Ÿ4w\��!��=L`����'@9{�`4Lb�,`�թQ���'���(6�Ӿ�x�J!��:����'*=�� �g�H0�- <PMz�'y�0�q��.)(�� ,׃
��"�'n�؋��O�7G��\�*T����'>ys����?ڔp��o֜��C�)��<Y퉟:��|�go�)r)l����b�<!cn�/@���bd��u�*E`B��x�<!2悑D�\)��D�2�svMIu���p�{�cY>/QB��e��0"U𥣗�y򥟏=Ҧ` ��Ns�X���=��'+ўb>i��C��0���2���?� 	 �M7D����ǔ` <2A��c�� �V����xB�Zv�L$��,Ωw��TI2KK��y���c�:|�!K�>̨)�d0-M�=�'9P�	Ǆؑ0��H�Pm�;R��

ד��'��a)�A	>#�����9!�>D�
�'�����I�O��� 䌑�q ��'p��˲d̩��,�@f�Յ�;�yRK��|��� ��wI���V���y2���q�h���F�.#Z|XƬȻ�y���L�\�c.M�%�������yRdհg_�Tٗ"�>�IEfނ�y2��^r�9�%�/�0�0e`Å�ybOڪQ�n��T��"��Q�տ�y�gS�+�T�sdo�3_04Aլ��y� �?/l��nK� Jǝ2�ў"~Γ�j��q��	���[�
�)|R��ȓEA�y�h5T����Mȇd������?9g/�r_8��֎ط1�@PgDx�<�U�ъl��fS4+�8 d�r�<!�B>p� K�V� �z`��$F{���Ŕ<M\�0�	��j�d%��7�6C�	����b�)u-&�:��]5C��/}����LϪm'��9�Fߟ6 D����<Q��-se��#�_>v���z�<�N�	s��L8'U��hS��t�'#�?�hd/� d,��7\�xiSp�7D�� >}6�ͫP�D��#�շc�`��e=O��Dz��IG	�������������D�Q�!�$�]�X�k$">n�R(@'.�&F�Ї牑I�I�@̙ �`쏨V�C䉪&D$![a�!��E�	��B�	�N�@�0s�E�$$K�	��(�pB��Z�Vi*R���N���F��C�I�q[�0�*��Y�0�I=��B�ɷ)�b}�r*K��
�ę3�ZB��8Z���B���Y�&�Q2,6�_8��?a�@ăD�X�@'�!&^�vc�}؞� �Z��j�41��p���-VH=��<���ȓTZBmqB��*J�����i�&�m�/1�	[�Ok�̸��&Ze�πri�	�'~l���G�E]y`D�B'T�
�'R�}Q��8k1�X#��)3���	�'3ġaǦR��jY�ťܱ|���	�'2\q�Y�&S�$T�BvRt1	ϓ�O���#f;�6���F	{eܩ9�"O��x��Ž��,Jc�ךw}�!㗟|"�i�2��>}ȱ�U?Eɴ���Δ��@�1�Cz�<�gC� 8�`�_'/��I��u��u�p�$�>��O�X��̙ƌ�(1�q��2F�zC�^�C��R�z���!@ǐdJ˓�y��S�\T�d�����C�G�q�:C䉸:��br�ʄ0�l��G��dC�əZ�*!h����`�H7cǚd��B�	�>x֤b����R6� Aj��(��B�	!g��F�P�(��q�M�(��B�<6e��b�D<h�p,�y�B�	e�̉����<>�Xt���J�CƲB�I�Y�X�;��ݡc� �;e<]�B�ɈZ<��4�T�����$�B�	�Qiڹ�R�D6U8���_�K�ZC�ɐ_�Ȭ�JK�QT��wR -�"C�ɷ8e��X��F��Ԫ��"6C�Ie9he��Ԍ��ȉ���3lg2C�I�6��$��CT�P���:�%�7^`�B�ɶId�h� z��L�< ��B�I
T-� 
���d(fp(@��F��C�����
�/"�bV!.��C�	�	i����S���t��&��nz�C�	)��4��J� `��f��6B��.�����A*b���ʒ�n4�C�lR9
$�I�T�شk��B�	�+� � �BO25h�!�5N��Fk�B�I�jhy����8 �!�*Ћ�C�9S4�@��4&��p@�*W��B�ɑ�H�CA�u���+�d9�6B�ɹ!hآ�R�tȐ`��=s_>C�	�~���'*�=;*�P�`*T�-QJB䉠6]D�jt�9:,�T�k�?t�(B�	8Y=��Q�N}�,��lN_#�C��"�*Hs@�C�l#����L�4/�C�� X�@Y�cƇH��<�Gi-�C�I�<�Mp4!��F/�dA�f?\e!��� s.�IeD$-,��GŚ�@/!�ă�C�5@3l�})r�⣍:i'!��%	�4Xg@\*&$X�c\��!�DΛcT	�m��.���!@\�!��]e���ZP���J}rS���0z!��P��[���;w��P�Cτ:f`!��6�$)B��.�:�P��<w!�d7%6���bސ����v�Mb!�� BQ2Vk��48u#��5[����"O����(ð��4���Gߴ @"O�X��/ݷ���ÖHڤ6����"OAQ͆�a)��PDʜ�_Q.eS"O�Ժ�坎z	��;��k ���'r�'���'�b�'��'a2�' ,x��u \aZ��S�+GT8h��'q��'C2�'B�'b"�'���'�T��!�	�ȼRm	%xmF����'��'�r�'���'�2�'g�'�&�Z���=7Й��)�
	���/�?���?���?����?	��?a���?��E�)���Eo͕v.�����?	��?���?��?����?Y���?aAO�+P`�|8�LN�n��p�KR:�?I��?	���?a��?!���?���?y�$�3X��[��[dd�Q)`D�/�?A��?)���?���?Q���?���?�� ȣn�$s�[�S�t0��Y3�?���?	��?Y��?���?a��?��׏������[Z�*��D�L$�?����?���?9���?���?����?���C.8b��"t���b�S��?���?����?��?q��?���?Y�f�L�� ���)O�z��TL�3�?9���?)��?i��?���?���?I�e�N����ݰ\��	��%L)�?���?���?����?����?���?ač��d�4�j��@�^��,r!�E��?���?1���?����?������'�B�Q;`@ah� ��0�%�m��B�˓�?�.O1��	(�M��5m-��*�.I�$-gAOuL�X�'��7M<�i>��4�5�$8`)�?Վ�[3+Jßd�ɑ��m�T~R1���u���b�~,ZeA�� b:(1̒���'rY��D��
3g��va
0j�m���7���1OT�?A����K�,�`H�+����.���%��?���y�Z�b>�ґ��æ��a�|m�4Hīpv�A��<�
���yr��O�ɋ�4�����!���2!�""W����B�kj��<aK>�2�iQ,���y�R�b����	D���ف�߮)��OL�'"��'��$�>+*Q�
 ���sNl���q~��'�(��@�C���O�*��	�)BǞJA>�h�O�Y���5��(@��y"�����d�#l�Pj�z��4G�S���DϦ��b�"?��i&�O�	F���Yf�J'�4Ec������O(���O�5�a.b����t��Lʳ�P��r=�𻴯4������4����$:I:��L��|B��C�;��m�'�7�,?�1OH�?� J@_#B*���x�·̛����O���t��$>��������MNV�F��Ӄ�!y�l���bk�@���
�m}2�ƾ/"����'�l��O�,O�M�W}�΁rVm�77F��P �O���<��W�mj��`����ݬ9���tK�8Ռ��Z~�D֦��?��<����?��6����"�X |g��v$F*,d����M��'ߌ�HU�'l�i�Sq���lc#���Ui�C	Pz�K�Iؐ>k��K�;O>���<A.O?]�F�E�hYЙ�A��ļ)��0���M��i�a~r�jӬ�O^�Y MŨz�)�hGXH���QMg���'{��'~��J�N��1OB�d�Or��ա��F��)��ڔN@j�)�&���?a��;��|�.Op�$�g\��/ڥfĮ=��5a��%�d[�e;�j#�	}�TmL�L��!K�B��h��
��ċ\}��'��:O����dN�.��8�B�_�p<�EA�Y\��Ҙ L���������$1@�+IN�	4��ɪ�+�4(X��Ā"��������˟L�)��Ey�bnӼ��1��mi,�h%�ʎg��H� �U$Q¸���O<@lZT��/;��3�MSu�N7\@|i ���Z�d���ЦM`���'N�x2�i�D�O`Q�?lJ`�S���P��7��q1df� �H��Vfe�l�'���'�B�'e��'��>!h�1�i�9T�|��jD	w3T�2�4.�h(���?i����'�?!S��y����L�"a�M!4BPs��¶	<v6M�����	�"I|6�p���bGL��)YB�]��@8�Eb�����ߜ$���)OD�]y�O���R���-"�9B�.�Ȱ��D�'��'��ɳ�M$&O��?��?97��:>��b@e��6�hpׇQ��'���z9��hj���IU}��#i�H�cnP�cs�Aڿ�y2�'�%'�?4�]s�O��	�wZb֝��?�vD�$�.�5����>�c�J�2�?����?y���?y/��p��?E�Id���+3l��J�r�REk]� �e��5�M�"c
.�?!��&�4�L+�%V:B��I�v�I��R���4O"�oZ��M��'���1�4�y��'DR��U�WJ��R��Yr�l�����K�f��&D�'��i>��I����֟�iq�̍<3p��kS	|�*$ӡ�<�B�i�v�iu�'�b�'~�O�r�S3!�Q(#(V�lPư���Ó>�l���Mm�8�Im��?�	`�^\��o�~2D��`S&��0������8L��!��u�o*��<9áٽ2�t�{�)Y�K$��Eƌ:�?���?q��?�'���¦��o]ٟ��[��!��t�ݙ��
*Ulv��I��M����4�����nZ�|�(EuN�0�P�:z�+�gЊ
�Lm��<q��Fl��GR�>�����?U��@�l�8� �y23��i���A��'B�X9Q7O(�d�Of�D�O���O��?��anC�z���i��CMߟ�I�d�ٴM[@�ͧ�?AW�i^�'�YZ?j����b��S��KF0O��Sۛƌi�x��X�87�y��sB/�g��q�_�k��Usu�H�N����F8���u≃��4���O���|[Z�XCb�A�<�:��Z�����O��c5��
-��'��^>!�AG�r����Ǘ�")��e
=?��S����4T���8Op���I�`h!� K�36���,O��4Q�b C56�D�`��\��k|�Э;S��'��Uu�+z�����]�^&L!��'e��'�B���O�剡�M��Ψ9#��2��b:1a���	�҉����?iD�i��O�=�'��7mG,T;3m�:S1������j�x�m�˟Tr5Ȉ���Γ�?�Pm޵�lU��O~�A����"dDw�-�A����y"]����ҟ��I��8�Iҟ��O�^���g�7�lB�Z8<��+u�v�<���O����O4��������>hXVXQD�%������m��4{��&9O"��|Z�'�?�RkϚ�M��'�D��FėzP���d� /�}�'cD,��D֩��|�V��S�h�"�B�H��P�S�ƾ@ƾ���(U���֟�	hy�Nq�v|CS��OL���Ox�JB�+��A7�F8k��4�  ����d�O,6f���'��-�&̏�3����cםadP�'�B��O��B�E���$埐=��#j�}�������t'�'�}#S�ٵ������?q���?)��h�8���JVZ�����B�,��k���D�=���ş��I��M��wo0F�,���/T2�Ub�hJ�y��`�]n�p���צ���?��. *XR��S�k�"hƄБ��]���'�U*c�f�!J>�/O�	�O����O$���O^I��U�5
|�5j�_�$D�0f�<YA�i����'�B�'��`�E[	E_p:�iG�FB|��N�J}s�6$nZ�<I���5%U��4G�J/�@[b*�)}'�mAU (^��I4S:L����'��-$��'y�k力���0�E	�	4H���'���'�����_��۴<��������1�M�
o��	��J���<����U��D�vy��'����'J��Um� mz��b.R��d0���Mw�V�����LS.���I��۶�M�i`�	����*�u0adI�<����?����?����?���d�5hz�S%���tL8#��#l���'¥g�2�B�ʹ<�r�iZ�'D��S���k��9ɐۏv^�D�44O��\ڛ��i��Ɇ�$�@6�1?ab��
Ls��*�� ���S�M�#ԁ�%�O� �I>�-O���O����O�%
�c�`ɡ6N�,}1��J��O��d�<��i�<����'���'��S�4�H��ϯ<[���d��0)y2�R���M+��i��*�Ӯ>wl����f���x�(��Xv��s�� ��c��/?�'R��$��>u�yK�$�	L�!
�`J'�j�S���?)���?Q�S�'��D�ۦ�3���#r�Z0�R[8U��	ږ�e�I�$xܴ��'HH�]4�����tI�lȕt|��2W�
M��6��O�@���b����柠:	Q?"]�t�<?	 aB�'d9�T�[�#�<�����<q*O��d�O��D�O��D�<�'Rx,�
�l��)`�.8\جP4�i�z1{��'��'���y�n��n E�45sQ�D����#�)�1
�n���M�'��)��QT�lZ�<!�T�[n��/2g[(���O�<	��ޱ�,��ƹ����4����ٸ�er���4���ƣ�$f�<��O
���O��w��V)�_B�'�҆øR��PA��!�p`��Hn�O���'`�6m���ϓ���� �� q,:&��f �I
&�
�8r"­3(c>Q0�'���		��<hc��x����P/:��IП|�	ğ,�	Z�O$��<@%��;N�Ƙ�@��E�r�n�$!X�	�O��$�ɦ��?ͻ��u�k�P�7Fִ	e����'�z7�զ��ɳ9�n�nR~�B�	F���S�nv0��@kMx�21�R�/��Pv�|B]�����������IɟlZ#/_ މ	gL����;f$Wry�D�䨋�`�O��$�O��?��f/�:0Bq#QhH<1��=0"������ɦ� �4�yR�Ӓd�	 	�m�	�ʦC�����i� �
�I��\��O �K>	,OH����:G��`��䋯h�Ĕ���O����O&���O�I�<�Q�i�`Tjt�'2����A3|>8ۢ�6\��U�3�'�H6'�	����O�7��Ox$����se�Q�ӑ�Nx���/ ��7>?y�A^�J0��8���5f	0WV��t-�/AR\شJG��yb�'�"�'���'���� �ZY�E�P In�HC�O>%�����O��K�U@��y>���1�M�J>��K�U6Ѣd�
�C|��d!���ybU��m���MC�$mBݴ�y��'��Qb�
�+0mD����@x�h����H���"L.�'��i>��Iğ8��=�ȳ�?s7 3 �-��Y���l�'x�6�
�kB���O��$�|*�i��x�!��#szV�pQ�OW~G�<����M��'a�O���h�%Ĩ��i�t=�Ya��#��1P�IޫU�V���Of�镽�?!��'�$�2.���(���QDP資+�j�f�d�O��d�O���<y�ixZe!�N�'�:�B"�~l�d��Ú���'iD7M�O`�OP$�'�66�����
�b'H�fXpr�ШE|~�l��8HE^æI��?�����8�4���Q~
� ������"wZ�`d��6��b6O���?��?���?�����F�",�qg-
?i��Y!�ںe`6�o�!eܮM�	��p���?]�O�	x��4?�pePF鄐����-�K-zQo��M�'E�i>��Ɵh���p���;OV���ɚ^\T!��G�2�4�`�1O�Y��%��?irm3��<�'�y��B�R�` ���=������?q���?�������z�ʍUyR�'|t�+�(ݫ'Fl����:��ӗ���I}��}��nZ�<!�Or��/[(��  REA�G������� �J�_���ys�;��_�B��< P���m?6�yg+or�	��П���ϟ��I̟pE���'���se�O�`ps#T�`�a���'p@7�Moh�$�O��mZ^�ӼcT��^�@I�-�D�6����<�C�i�7��O,�dӤ�C׶��0��|��I��]�\K�)P�|q��Ţ����4���$�O��d�O4��	SJi�!2M�4�h�j�:� �Tћ��	5V��'���IW�3Dh��b��N�(���8!{���'à7���� O<�'�b��-�>������h�a�ӊg��,rFFq�t,�*O�q��]��?!�"���<	�厪>��xj���i@3P�V�?���?���?ͧ��D�ܦ������g�?r?Ę1v�A
;�n�r4@T��z�4��'����?Q�4�?5̓�~R���'�J�E��4"ՠ	q�P)۴��Dӈ4� �����O���آe��8׍`W��H���Q� ��㟘�Iޟ��	�x�	_��tR�	��!f��M�0�)8�QP���?���&��
��I#�M�I>񒎊�Fr0u��(ԍQ�2�s�fЬ�yW����4n��Oi� �i����t��p[�G�	�d�#T��0�	���>Ux�N{��y�O�"�'��AͰuut��5!4^���˄�ĈX�'S剡�M�-�:�?����?y-��M@E]�#<$��Ř{z~Th��|�O�Yl��Mc�'!����`آ?�I�e �<zt6��_@��ta�M��i>E��'�&%�4r�M�d�7E�=J-��vb�ӟx��ƟT��ßb>͖'#�6- �^ޒ`ps�%>����u�M.^���"�m�OR���হ�?��Z����4�|���d�@�!��O�����i��6�V�N$�6mj���	�&[Q(r�O��y�'h�A�'�_$��(c�"�����'���ݟ��Iןh������a��1h�LUi��{��!�&ؚgV6�$L��$�O��d%�I�OX�ozޡs�(��rt���QL�T7����MS#�i�ɧ���O�RR!^Ǜ�7O^L����r~��U��t���� =O.����?�V(��<ͧ�?@�.5ٺ<Z��-!@���o�1�?����?��������R�Ey"�'Sڀ��ի
�X�a���!L��(J�d^\}�Du�|�lZ�<��OpXC��5!�4�*]U����;O,�DN-�tx��Q�~)���?1ж�'�R���?4��xB(�#6n�!�s敘kn��	Οl��̟��	q��yG�V�j�dq�7*ûY��� F6e�*uӶ��&K�O��^禡�?ͻp�P|j���4<|?},i�f�u���ܴ 9���'m�({��i
�$�O|��u	E4��)�!�͂U�ݩR'"=0�b^M�x�&�,�����'���'n��'|�T	s��]s�!�ԩvM�M�eT�t�ܴ *�{*O�D/���O����ؑ/d��Xt�)-訠�a�E}��e�>�n��<�H|Z���?��nɠ_	b$�e�W�%���	J�;�P�� W~�i'A���I.��'E�I3n���PP���7�8Y���#A�U�	՟���ş��i>��'8�6��k����>�~� ��D:2�(��Ꮫ2�h�D�Ǧ��?�ES��qܴj�&�'H�IRWDF"�0ئ�ܩ=���kԆF�B��1O�������'��	�?19_c�@|�1�q!q*�_�@cnO$�y"�'��'���'�r�)T�"+��gnN��*�8#��"2�'�"�'��7m�:LE���M{L>ѷ�^�~ւ��i��dQ!OB�yR]���I��瓀_�H�oZf~"o����8A�LAq6Y�����%Fj�S�r�$� ����4�����O�����I��M�ץL��F����3����OF�Gԛ�*�f�r�'+RZ>�T��B���CN��V�d@c��>?��U��)ش+��&�|ʟ�
�J�+(Px����O+hi��n�(M�`�4��3��i>2��'Q��&�8�
Ar̈́qa���"�>��������ß���˟b>��'�L7�)iBe�%*�G���� �z��Ųv@�<q �i��O���'d7m	�=�� r�ߣ~ޤ� ���V}o���`�*��'�D 2č��?���n���Ԅ$�����2`�5ON˓�?Y��?���?i���i1 ��Y�Ƅ/2�!�V�A)qF�}oZ+5O������ ��~�s�4q����e	V�y�1 �1Ա��ڎz��6Kb���L}��D)�)S���:O��VC>[��aɢC�V��ՈW2OD��KZ�?yd*=�d�<�'�?1�b�u�K�:O�^�*��P��l���������yb)�Os��'���'���SJ�Q9Ʊ�A��z����$Uj}�j�2�o��<Y�O�l�t��%)tMs��Q���u��Ț�C>>v9�I �S�9�K�ڟ�"UAJ�,B��!C����m���t������	ğ`F��wz�;S���mHT��k��)�r98�'27���|���O�Xn�N�Ӽ+�Ȅ�@�,���D?g��
U	��<	Һi�>6� ٦�KaUߦ]��?�A��,A��	�`�? ��SD�2:5R	��lϿ�Ē�g0�D�<��?����?����?�U�ۑ	��`�W$-�pp���L��צ�	ǣSş���ǟ�'?��I;?|�Mb5�ԧC0Y�wDS~a���*O�DӬ��U�O���u@�3E�(R��F�ęT�� ��Oމ31�ο�?)#�(�Į<�a�jV}�壔�h�HQK�l��?���?���?ͧ��d��d����O䬒�kT b�A����{�g�Oܩn�p��W��	ٟoݟ��1��=�b�IAY<F�(}w
¾B\�mi~rEܙ�lP�Ss�'P7k�ݫG�b��e��]��	iFǩA��O���O��d�O��:�ӝ?d����
,:I^�	t�@�����������Mk���|���x_��|�i�_�v� ��CH��XYR�C�D���>Q��i�66m�O�� ��u�
�I�\�ʗ�Z *��gx��F,ܔ�%�'3�u$�����$�'�R�'�1�c��+����������'k�\��#�4 [��B��?�����0G�б�mG�Bp�"�<iX����$���J�4�y��IK�445��,�8@��<��kD
i���K��Zǜ������=&7(MS�Q��=�RR��\�P�$?tD��۟��Iٟ��)��Qy�w�r�P"N���-���Zu�Zr0�M�0��O����ئ��?�T����4ca"3� ɇ!�J��4M1{�"����i�r��}5OL���tK��
���!Y9Z%�.��P�(c�l�+�	RyR�'���'��'�^>�9Qꚷ_�����%'�-�A�?A�h�ϟL����%?I����Mϻ^���ӡF��\�g&f^A��'�f1O��S�Ss>�oZ�<9U�]>(ǌIc��T�#�-cEc��<�r��4w@�Բ����4����٠,Ր�AtB��SŮ�Y�ş{�4�$�O����OT˓u����(b����"Q�A��,�U��o�N[���]�A`�I�M[C�io�D�>q7Ì|6��BB��"UHl�;���p~�/EW��P�l���Ou���I+���Im[�](ũ�?}*!��C�� ���'���'m�����3�I��1zW%LH6q�g�Eɟ�`�42����)O�\m�I�Ӽ���Q�\�P�q���a^�ucg�G�<i�i��6��O�,�Cw�`�f^dp{Vc�X���gڰnL��%���	��Δ�䓑�4�.�D�O��$�O��FnZA1���<$�AJ��Fc��4S�6eR�B�'�R���'�:ʥIÅq(:`ˉ�HL����Ȧ>�v�iv�6mi��D�$�>YVh"�&C"v_pШ ���d�t�����D99,�����A�ԒO�ʓ<��#r`�3r/�ij�K|��Yb��?)��?���|�(O,�nZ�$�.��I6D=Ѕ�I��X��x�(�����Mc�2@�>�b�i�7M�Ox�1��9`��U���97I��i��f��6-o���	�?��8���O�����ѷƆI�c Z�f�Ye�3&U*�0Q6O����O��D�O���O��?��C��f�I�M:C�d���������Iޟ<�ܴ)	�X!/Oho�q�@ ܩ���=;����iV��D̓��d�Ħ5���|Zc��'�M��O<��A<,�Ђ$WR}�,J��˗x�X���<Hp�OZ��|���?9��6_>A�����d�p�cn \���1��?),O,�n�$�"t�������l��n\�0��adµC��x������� N}��h�Z�o��<щ�D��� �y���+n�acF�$�J9P@���S X0J�O��@��?y��>�d��(hP��x9��A�k:����O��d�O���I�<)��iYtQ�+��y�ą�lI�Ni8���E�%���'��6-,�ɰ��$ʦɡAK��KO(h(��6^dHr���M+��G��ܴ���ѥGr�����ӓ��t�tO�fBN9��cA�b�'���ßT�Iٟ ���l��Z���c��)�_�De����OG0'W�7� $��$�O��d/�	�OtElz��bo�C09"AL+i~5 �ˉ)�McA�i��>�|B�ɂ"�M۞'���̌�}�>�Y�i߹X�4xK�'��xҗ�۟�%�|�[���jw
��ZX�d�Be7^F��D����	ޟ4��Ry�u�@<�"��O��d�Ol���ʓ�N�I��,��,;���O��OR��'��6�@ئ-������~)pB����YEX�{�����O�I�C�ƘHuN�q�����1��ş`s�`,�%'2.��%���2�$�O��$�O��$?ڧ�?ɑ숒.�4�+�$Ώ��Yt@̫�?��i���!Q��ߴ���yw���YCmi'h^�2P�J�Ǝ��y2�pӄ�oZ͟�Y���Ŧ��'=P�A��N�?U�e�
bj�I��O�sV��*s���W�'W�i>�����`��ȟd�I���.�n��V$?7��ԣ�P� �۴>��)���?1��"*����q�E�rk��m����8�.��'K�6���%���'���#��@J�rBx��I=,;���4���8���'Pv"�K�쟈�W�|�[�dV睊1v �E	�֠`I�'�՟��۟���ߟ�Yy�b�L�ÃO�O������-Πت%$5I��ّ�O�@mW�{�I��Mk0�iW��X54P0%O .�ʸ2�꜕X��	e�i3��Oԝ�+G���a������5�iY[<U`��s��Ǌ��y��'�B�'���'�	˯#x���+.-�I
Wn�����?���i�FU`�O��pӦ�O����!�0!X�\;��C���rcj� �'������ �F��p!#� ���'M�Eո	�Ն���X-�A���?AU�;��<�'�?)��?1��_�h� p��L�{�apOƻ�?	���?��l�A8���?1��?������3Bw
I�	XP��!FgQ���@y"�'��f��OM�$O�
�*L4��2��#ե	f��ݸ� BK�j��O��i���?�j&��(���qG�d���J�ǚ�n�l���OD���O6��i�<A��i3�4j4g�tH�g!"��ڵ�I"Fp�'4�6m3�I���d�Ӧm�gσ2g.�����y` c�nʦ�Mk��~��Xݴ�����i�����'�������!�߄J�\Իd�I/_�|+��6�=H�LF�A�D��bͺ8�F����ڎ^�4{�N!C>��kS�W�M�Ҁb�	
ج�b zR�� -L��p��#Rر��T�a�b "��?�p!3��ccx��6.E�:ڨ��@ �Ɣ(����&a/6�;���E<���͋�%���r7��)���5B����;S��(}f0{�߰k�pX�E�E�La�p&��3�R��Ս��T�dd(�g"k�p�QB�ӦG� ����@�XI��ҧ��/��T�����"��:{9$�iG�|�eC�/r�6-�O:���Ob�IQ�i>�[�f	 ��[��?-l�����MK��~�[�\$?�Iӟl¡��-4����B�* �rMbT�L�M��?Q��9�Iu�x�O3��O�����1r����	�"�8�K!S���'Fբ�y��'?��'�"�����q�nX�V)�"m�t(zccӘ�D�)7��'���П��	my���*�P�7'/0A�����B��7��O&e1���Ob���O�˓8��I�����y pF8LN�m�1��0J�'�r�'c"S�t��ݟDS�AVu�]Ju��yz���=�Hc����L��ey��dr��DG�`a�c��M�h�@��?H��?����䓟�_+K)�	1�޴!��}F�24F�C���?����?�.O��z�H��7�
p;��}K��*	�Tb�
ٴ�?�����O8���?f1�<�pGH�nT �cK�$t���������'VX ��*�)�O���ƶ���JZH�@���w��X�xBS����9�'��t��>��삃�&V�8��w�A�M�/O ���i���eq��p������'2tl�w�ϩ
TR��Dϫw��0@�4�?1��\�~Qp-O��Ov��x�J$|:�)ȃ+A��k4D�Mۀ^�g&�&�'���'��t�$�4�v� �^�{���ja�ZZ]���N���-��:?),O蓟��OL5@��ɗ�=AnN�?2�U2������������ N<�'�?�'�`��i�$+R03Q��}P8­O&˓w�Zu�<9���?1�8��,��\�t�$�&��kU�C��i~����D;BO�	�Or��<��EH -
��F�J;V�>�9��F�M����'�H��y�'�b�'��>MJ1����gF��*��ԝ4� $�	���?���?�+O��d�OVa��B!=ݡ�.3"�I�eB�}@1Ov���O��ı<��/�}���N�W�Xi�!�=c���'�W>k���͟�	|��My�N�����8\���C���w��	B�X�8��՟<��ßx�'�(1Ҍ.�i��'����'T�2��%�FD�[�ܴlZß���sy��'�����O'��@6�"H�X�d�B$[����ٴ�?������ƫo�-'>M���?ט�-�<�UΠ1�n���/�i�Ot�q�E��ޟ���G
;rzm)Sㆵ`$��cU�i=剻RϬ�9�4|��ݟ8�S ���X@�iS��{�д�7�^�=1�vP��vg5?�O���M�0C����ӂ�2Z"yzt�LŦM�V�V��M���?)�����x�O3���� �b�4�����=+q}�Ӳ$ d����'���yb�'��'�4U�!)��S�|	
%�`�,���O�$Ȋ"�@��|z��?��'�.Њ���P�-qd�� �~�X�=�I���h�J|*���?a�'Qb�Q殞�֩�#�s6�:ٴ�?qӦ�����O����O�㞴�S����!�4�Q�
�m�GD�>�QFX%vs|p�'ZB�'��Iџtqb5-ZX8[4���3I�c���=0kd�'���'�R���O��qYk�|�8�%G�x1�a�d�ȟoO�A p~"�'�"R���I-�x�'f�KV��O�t��lѸE�jm�ß���֟l�?��;TH�R�kF��1���ߌU�<�Ђ�#D�n���>!���?A.O��d��aX�'�?���ݗXkN��$ ֻN�`��)
�
��'��O���B���`x��x2� �&���?oJ�:�����M����
�F���M������	�?q	P��"!��Q6i���ȗ9��'�R ي�vy��y���e wI��`T�1BY�����#^����m����՟��Iʟ���NyZw��+5K(NÒ�Q��A&^�:�O@˓r|�AGxJ|Rw�F�~L�f�ӝwYĴ����)r"m�����Zy"�O�i>y��4$y����Β�s\�4 䞤)�eJ�4�L�aTb�S�O���fD(����©�t�+F-A1�5�4�?���?!�	ұ��4�����OZ�ɂaa��� ��8� �b��W4	�0��yb�
0x������O��ɳWp�!��ôIx8��P'{��6m�O ��%)�<����?�����'�6�0��8K9�I�c��.�J5��OJ�3b�E�l3�	D�	Ay��'} )�G�J�]��8��#�m˸����}u�I̟8��ϟ��?���Vi�|i��$L)�x�tdV�CO(��V�	9వ�'�"�'B��\��Eu� ��)%� o0i�HP1)�2�Y$�i�R�'#"�D�O�	��N�^��v"״	aj��u�J�F'�� �lI-����O&�d�<���aP!)�x�d��0���G��`���a�^�R���mZ��H�?���/��5h�_≀\�� ��S ^$��T�Z�P 6�O���?���	���I�O�����	1�
}p�LAd
��ƪ��Yp��>��B�A���c�S���7�����6o��+į���O�����OT���O
���,�Ӻ;�	��P�𡘸Ae� �S�~}"�'@����#����O�-�EF��$j �S�Ѯ�l�ڴA
l��?�-O��)�<ͧ�?1��	�{��H)��ݮc����w":��F-�9z�@ �y��i�OF��`ۄ�E(�A� U�=�#Ǔ䦅�����I�:�<�����'���O4�a�5X��A�
1m��	rv�LE�Z��a������'�2�O<���b	�y,DUwf]�O�p��i2��=*���ٟL��蟈�=�d�i�P��pӤ\�DU��u}�o��ig���Oj�d�OF��?Y�/�/\ϐ,SD ճhX�vK����J-O����O��$7��ߟ�{��F���$�ЉQҍ�*pZ}��;?a��?�,OV�DF6D����54䜸�qnXh��(�1|�\7��O���O8�8�	.Sj����y�ڜPi�+EiX���h$'���:Y���	��x�'��M_���㟴�� A1�$�a'�T1Fg2}��� �Mc���'B��Y:�`2K<�cf�3dؘ�K(F�n>�|����ئ-��Gy��'x��8#R>�'0�4�٧"���# &2��a �N�*o�b���	"2��HY�`?�~���.�t,�6![�6V�[���[}��'�\� ��'�b�'<r�O	�i��A���E�J�N�m���1��>��t5*!��q�S짓]��u�a\��C�'9���..���'Z��'(�d\���ş$�fd�1}%vxyև�?� xQ$ۈ�M�tƐP0��<E���'����%j�7kҤ�4_;f'ıA� |���d�O���B��2��|���?I�'&|���"C�u~R�yR�H$1���-(�I�>\�d�N|B���?y�'yrt��Ξ�uL�c��]�>X<%�޴�?����/O����O��$=�	�hQB�c�C�-�(�U(¹C���HgvX���W~��'�R�'��I�W?:U�¡��\�����6K�����S���?1����?9���ذ���� �~X�@MͤY�h��ӄF�?��?���?���?��J����i�t��ڼ5��ͨ�c�,C��R��%���O��O����O�y�i�O�@���A���2U�ݝ^Kly!u�Ǧu�	����I埸�'����W��~*�n{�hX��@>J����_ 8�XA�i�2R�4��ʟ��	$R���I��CT�K�*+6�R�FiCS��%m��X�	JyR�F3B��'�?����ҵ.V	K����Ď�u¢E�/�=8��矨�������o�\�'�B�ן�5caI%� �q'�F�����7�i-�ɣO�p[ߴ�?)���?��'��iݩBP�I�W��Ԁ�4��XG"}����OTr�1OJ�İ<q���-�KԺ��TM�*Q��@P�폁�M��7'��V�'r�'��d�>�(O�]*C�ZjJP	$>�>,qF/X��ͣ��n�,��GyB�	�O����
�BMJ�X�(W3v`�Fϑ����I�d�ɀR���	�4�?���?��?��m�0XI� �~e��b�KM�4�io�ǟ�'��R�����OB�$�O2X����#Y���I�C;d���Q��0� ��ܴ�?����?�R��I?�����Z�H�E����	�'\^}2���y�\�$�I�����sy��:Z��~*�hГ	͕����%ΨZX����d�O���?���?��	I�T�<S%KY6K  ���j	�!͓�?�����<���?-O��Zᬇ�|����{�4�`E�d�Vt������'J�S�����,��;j���	3�-x6/]�M����8%ر\��])W��':�6f`���d�D��ڐ=cT�ε�2�GE�],�ElZꟐ�'+��'�����y��'��$��`�!�(�DEiI@�q����'U���I�9��)�O��D��<<��Ӑ���I�b�<��95�_}��'b��'���c�'��'��ēH���(��I=?�D���ŕ�4o�Y�|��n]��MC��?!���*�U��ݔ5h�8��T�P�����I	z6M�O���2��@O�D
®+�q�����熛^PL�g�[47:���i_�y�ajӬ���O�����A�'n剁?�
�0Ɔ������B�K$��޴,r(5��䓙�O�ǘ$.&#2B��eܤ0@��/2�BR�'(B�'�N�+SO�>)O��ļ����l��x����K�R082AaӜ�ġ<�"S�<�O�r�'J�l��$b��Î~ct,�Q�CBb<7m�O
,��oSN}�V���	by���5��M	t���Yԭ�2�~<��Y��D�+7��d�OX���On�D�O�˓>�2X!���@R����(yӪ�2B�>��~yr�'o����������uB��JQ�Jߨp&��,t*N�	�IΟ��ğ��'Xfe��e}>a��X�<���; @ѕ^e��F(eӬ˓�?�+O��d�O����g���0��36ed���U�GԆ6-�O��$�OR���<Y`��F��S��`��/�s�U�BJ��I�T�@�M[���d�OX�D�Od�2O����O�eX���*�Za�j�_JP�j�#�0J`�D�O�˓����6^?��I�L���� ��K7�a�,3�G�>�B�]����ٟ<��#~���d�?��å֒AP�@V�؂z����{ӺʓW���s��iGb�'Q��O���Ӻ�DL�*l� w�-^."�AƬ�m��͟�ka�g��⭟�d:��G�ܥ���NiC2���� 	~7��$1�j�m�Ɵ��	ǟ��S��$�<9�N@�P���"4D́}f�m�2���Y�&�]��OD�?)��%Z+�gX�^ V���*_
�]��4�?����?���У7��Iuy�'|�$�'o�l������w��ph��X/`���'���,?��)R���?��o��4�W��R����7H��z��Ƿi�Rk_/| O����O&�Ok,��h��B�^ @�4�ؗ {�ɲ*�,��	ey��'����f��.Mn�(��k�h�bg
�JD��R�6�d�OJ��4�D�OH��[4T�(dXD��"��&(xl�]i3�"���O����O,˓4�4��@5����Q�M
!�
< �)W�d�S��I���';b�'�+P7����l���٦��e���ⷩV�3����P�I����'����#"9�	�2f:T�M�fA����v^x�l���%���I��,.:K�d,}��?.B�����:X�@UigK�M��?I/O �����W�՟ ��;.��d�#��D��·ac.�2H<9��?� g��?9I>�O�>i�K�.G���P�)�\e��4��I�yxN�nڡ����O���n~� ��x՘p��'+�DP��!�M���?�ׂ���?yH>���d�z��p
.k������M{�h�,�&�'1��'�J �$�O����Ζtx���B��.�ʠ�oP��e�tCm� %���2�[��E��2AȔm�0���-F0�(D�i�2�'�$�<}�c���	[?Q�
A_�Z@�� ��;T�rEN�9$�P���$��'�?9��?I��b"�v`�:%�H&�E�x����'���X'�/�	蟌&��X5)kf��.ُ��T�d#E�&x���̓���O��Ohʓk�Bu�"���qa�-^!\Pp�B!(��'���'A������۟�R��4^H̘H���UX�@�%^/�Ly2�'��Tf��Y~瓍	�<\ۧ�[�w�bT��	Y����?i����$�O<���Ora�6��O�y�3�!J��R�i�za���Ts}B�'�B�'��I�v2-�I|�b�Ṭ̌GE�B���a5��2w��'��'��'���sA�'��i�u�G��1 r,��o��`�1���~ӈ���O�˓��������'9�D�U`^�p0!5s�ViRS�X�7=�O����O8%��O,�O��	6�έ���4R:����)��7ͳ<��$��Û�j�~��������[����c�Pȓ�t�6�#�FiӒ�$�O���OВO��>��f�T�20�ɐeZ�	IjӮ��J���֟T���?�RM<��7�͠Į	v�,r�$�	]��yҳi�H�p���2�Sџo�=:�����Q�2�b�R�����'r�'(i#3�7�D�O��D��4藢�4L��8Q&�B����/w�^�O~�$�_n�ԟ4�	���h��ՒRR�����2����)�MS��=r� d�x�O:Q�<�F�N�6)��Q����9O�B��>�4��?Q+O��$�O��d�<�d,�xRf�< ��$	�0��@�x��'SўH�Y5��RЫњf�`���4�"To���	؟0��͟4��p�T�K�y��J�KI8H��E[�y���uf����6�'z"�'��'{2�'Ba{��*�MscIW�/���Y6�P�/�"�(w�T}B�'��'6�ɐ�D��H|/�-/�V�d�P��H��DÏu���'���ā�^|������¸&������s�h{��i���'bb�'��lʣ[>��I��8�*�|��LJ q=Ljq-��~�1PL<����?Q���~h��<�O��my��F�-c2�#���w8r!��VyB,��*�7M�|r����������	AiH�ᑉ�T�	;�cn�"��O2��)��&x=a7L�8����6o�;;#�6�F�Dn����	ȟ��?���?��:q�<�S���[6.���i�T������+���l�Vp��Z'�@2�
���M#���?��L��%@�x��'�"�O��۰*(T"�0�N&=iRe{��d]�a�1O��d�O��D�*0:��9c��_ڌ(;F��huv�m����xn���ē�?�����ct���� [��J�H�b�\]}iA���'���'tT����M00�R��1+l�d�J��\��L<���?�M>����?�#K�������ܯBR� է+[�J��<��?����6!����'}� �z� ]�gU�x�J\Qa:(�'�r�'��'�b�'e�\9�O��c�O��mA���4k�ZTz�^���Οė'���P'����O�����rA��EH�]�H������]�IW�	Kyb/��J-��I<Y�H�ƺ�ҔeQ�$��!�K��A�I�(�'h6�K$�#���O��I�b�.\�e��P�2(��A�}�� '�`�'��)��D�?i�7�X�:v1ӑF �8�l\���i��ʓ/���AR�i��꧍?9�'X6�ɺ���$��,}o�A����D�7-�<����D���O��d�H"�w�K>G��3�4@&hc4�i�'���Ot`O��v�? �B��		��0�5�D�F`� a'�ir&]����蟈Hw�Ź'��i���V�b���L���MC���?q��9Fs�x��'��O���roN�D"��`J��@��#U����1O����O��$˽	�Z��1��"!�4�Ůޒq+�n�럴�� �����?i�����Ü�_ö鱣��
�lyJ�B}�h���'���'r[�xB�ˮr��%���Z�4<��j�jT�"�1O<i���?�J>aM�d�/�54\48��� �t�41���>�I��	�t�'�� ���?��	�<�z�:$��k���	�^������'��'D�ʫO�y���ӛN�Ȅ�ר�	Th��[�L�	��	}yR�
�����"ؑ ��<� C�����{�O�릅�	U��t8� `7�� �x!V����t�tӺ�D�OHʓHX���W����'��4���<���[PL��'}Z1Љ֩�fO���dH"=����Ƭ�X�^�rA�� 2��W�J0����M��Q?a���?�!�O�Q�V�מ(&��,�2�i�iܡ� �ꊰ��Qt�3C��k̛րB�6��7�O����O*��@~����QW���r# ܓQ���A���#��C7�?���U���8G+�x���EX{}�����?9��?q7����'���'��[�Z��q�Uo�!bT�te��"�a{��'���'�J�&M]�K��Q5-��J�aW�cӢ�d����˓7���H'�LSWH�|� �K���}��AK#������ w�qO����%N^9z�JH���(4hI��Tn������yr�ƯW�H-�r瀭�6x+aN����O��j��/p���´���GJ��\�\�C�͖��ȡ���g�a3J�3�4�Z�B� �F ��;�썂bȝ�/_h�C�
�;8�ٰM�-"Q��rc�7C�P�s�d��(W朊�FI!-�[eIǾ{[�Xa��̬"@Ρ{��� l� b4�x68�a�:qh�	����
X�px큢 r�'?��-���g	4�ص�e�
 !V��'\�標uH�^Nf�`�Ա}��DDy�G�h�:(�NΞl/�l����D�p�	f�R��-"�[�X�"�s��6j���Gy�H�<�?�����Ollr@�S�D@�/2���s���<���mـ�	0�H�vBd�p�kI8@����I��ēH��`��6�\��]������<Y����4�Iџh�O�L`���'r�'��0σ�$�h�
'H�)A�5��D:��J�M��T�F,[I�O��m�矸���HwZe�͞�ZH�9P� ��p^05򗡑�r�|�F"��?E��6�����J(%s�M93��b�Iݡ�?������Ԝ|��4��&���`W���E���y�@�pZ����� 0��dr�@�=�O�FzʟX��� W[�,�2DJ�*��$�O��Ѵ}r~���OH���O0��J��?Q�jH�V���{�' N�W@K 2����"s�L�z��J�Akv�g�'���%�/q�C%�[�`JDd��m�O�L��!�!D�p%c��	�����þq��h�" }t��ǆ�Fe���a'��'ў�'�҉�Љ�=n�V� +��3I�b
�'�����ضk@���䆚{2��!� �S��U�������M�@�D��u��{h|9�q���?��?9��J��I	���?ќO8���7���k�M��Krl���]�판���Wn!b0P��'�R@�1"Z�YG"a!ct�kFd����B���$s�u@5�'�������?с�X�$m ���L�D��5������hO�?�˟�v�BЛ��
T"�[A`�^�<��EZb��З�aL-3b�X�<�aV�h�'&�x0�>i����	Ţ=���J'nG��jQ!�N�O�T	�Ol���O��)�〻w�L	KF��>�h�@�t��$�u�J�Г�6l�P��a��#�(OH��t��e��4��I/]��)�����߱0�r�!�+
p��y�r�I�/� �D��U����"+;���4,_�R� ��fӫ�y��'��}2@-S�욶%˷P��d ��0>�B�x�,�9��!k�g	��x��@���y"E�Qr�6�O0��|֬V�?����?�0�5Y���$w�86�� ��2v��8h����O�@��l���A r��1k.�3�.d��M�x^��4+ޯ&�䧈�.�2�N��r艜h�H옐� �L�F�(��'ٜ6�[ɦ-�Iy��?��Oʧj�y��j<d�-`CO�<	���>���?V� Df��%�^�˷�g�'�#=i��'�?�0�ѓ��uy�)�-O弩� ����?���^�$Qs��:�?����?i�K��埠����8pW��3���<0@Ѝ��#�<a�#�&S,�t�@�1P��EB���d��y �=+n�Jw*�/ U�I0WZ��B�ذt�*��hO(��a�	4 긼%�,t��:��O�D��On�n��M�gyb�'p�I&l��YC���
�KFm� !�u"O�yZ����"�l��A�A2j����AX�'�<U���Ė�ay�}�{�? ���DW�>����S�;��X���O���O�$ױ� �$�O���$��$�O��6刊j2��Y�m���X���'*���)OhQ���:d-�5C� [��ۤ�'h����?�	�<zM ĳR튱���A7�E��䓏?Q�������ܷp%��ǌ�t�F�C�e��(&!򄒋*�r�0N%�Zx�eo��~}�Q�HR����d�O�ʧKM�c��3��	S-ٶ �80�O��?Y���?��]6C"��'��M c
���ɀ)B�i H�T�(�ÌQ��Q��¬��u�BqA.�Tv6���?-#�JD	f岵��8sb�V�&ʓc�nL�I��M����W��~�˒O����4(\�i6���OL���*^gN�ɲ.�(AvU8tG�V9a|BD=�\ <%�g�I1%��遦%W+N�dOU1���'�b\>uS6K���d�	� �d���4ږC\'���B��	&.�4H���IV��P�F3�?�O�1��E2�V$5��>6y�����Z�]p�Y�l�9c�8T �ϨzbF���O�HfI=u��I�q΃F�V�rbPUa:��BԦab(O�Oh�DS���t�Fb� ң����L��!"D�dK�V \�l49d���Y�>y� $?�	X�����a��?d����#uJ�{�6���I�D�B�Ěc� Q�I�p�IП�s�� ��UGe"��i�	-�$��26���O{D����I�,�T�)�۾N����6e�Z�I�8�8q��^��Z�%�,��@�@��-����']�(Y��?	�S�'+S��
���q�P]�Pa0�E}s!򤒓>�D��F�A&1�R��GM�X[��Fzʟ��d%\tz�4J�4��:1b�1�N�DԌ����?���?9@���?)����DKC��?��t��8�*Z�_��Ȋ�.�L̅�ɉpʓ=���E�I=tni��ގj�E��Ɂx;��D�O�+�%��2�`��� 1����"O��j����~�Xv����R"OFX1��%i�I�-C�dd���?O��>��̝�i���'YrV>uQ��)q�Z`1Vg�
ܺ�Bt\%N���ԟ(�	�g(eP"��0B���@Ea]2�p c��ȤycTYV��2��[�����I�Y� � ���<�1�ڃ9>y�O� ����Vr��"%/��sV$��E3n�r�ӞGh�A;@ׅ�6���i��\��C�	�2.��iu�-g�*�8ŉ�L� ���V≚f��`[��H�V*�q�[<8�Xc���C
�j��Fr� (��W
K�2C�I9x3Qp�ϛ�{z����]��B�	�9X��!R��x:f��fЮB�	\ b����&_��ѦEU�S�B䉁l@�x���ڿ'��c#〣\oRC�I2l��یt�p<�r�P")Y"�����w��#��'�!Ot䄆�!ی%:�m &CT���q�$���0�⤘s��3^�@E��I�<&B����j�uNU�g36�h���z�J�3�"O�"��]C4C�)כd�Hp�T"O0ph��P;z>|���C�F�|	`�"O��p�F4Y,��e�c讐��"O�us�H�:u�����=�ԙI3"O�	�!��W�ʝ@g%�}���"O&T8�R,hg��r�+%�2���"Ox�d��"Ԛd+�b�~���"OD8���$��Y�D��^
�h�1"O�D�����#d��%�2��"Oh�9p]�"�d{Q��06��A"OLaх��)VH�dA���"�}�`"O����ǂC��Ȼ�*���"O0̋��Q�کS6�Ο#���"O�ۆ�Â"�X �9�z�:�"O���2�th�񬑏�P`�E"O�P����>��La'� �Xӄ"O���t��2I��K���\0I�"O��Zү9g� �"d�p	ZE{"O�`��X"m*Q�D�d���P4"O� �����<	h�!R�#_��xe"Od�9� �Hwʔ���N_��SV"O�HAƒ�M4�T&ܑ=�@�f"O�$�&�"j�<+�V$o�d]hd"OLu#$���y6%��&N�@Q"O��㲃�� ��I�1@�@���'����F�'�إ�F��K�~@�!R'At̓�'m|�zD*U�C�Z1ȡ*��:R���Ot�`�KE�t����=�'!��M�C�P�!��"CT��ȓtDB=�T�ٴ�l����j�FHC,���V�R���P�XJ=��'�ʀ��b�ἳ2Ƕ3G�\X����FP�Hc<�6� {v��t�Y�	�x��G��5�D�@2g�k'e���ϟ�?7E;D�f�p�I���D��NQ0,IҪ[
hmvɺ��5OBq�iX�UBAi�C�<IC ٰf�.�{�"��9���"�`@�*��<R��!�t��I�Q�<�e�Q#}�y�2	ԓf_�z.-�m�cM�-)O�踶��h5��$�"^���o�)m���R��$ɠT�24������@���x�CàA:���g	L�HM�'���_�|��"7	�^�2 W�N�h��w	i�bQ�1�>�`�(��A��=y�'�k�΄�V����#B2z�br	1���h���*�P0!"�'p�eƕ����P>�*L�q�F�ǆv3
�is%��Le�0���"�6��U�^�k�4d(��A5fP�����R�8d�p��Sh��+ϩ_nz0i3�ZoW�`:��Nx���w�Z�L��ţ���1;Ԁ[��-?�C��]�v���T|�]�������<��j�(�p�J��҅kq�}��ˉ�~8��?��]��'s>d�5L� �t���+(-C�u�6�S�3�%
D)�ҁ�0�W�L��e�3T�@@��#m��tɚwM1��Ł�9(��ڤ#D7X{�չ
�'�0��M�}�� %CV2	m�p1t�C(C��Lх.�rr�%�Ҧ'#���1�E�$=(�"!KFI��'�l��F̇E���ï;\��k	�j�>-�DM>>�� �&�M+%�pYA�&N>S�=��fW�#��A�U)�? �r�p���1���9����<!'L7v���E\��Di�c~r��z��a�$���BF0zj���'�<!+Tg���y5,Bu�DXA��N�j�s
�'R:���"�!�|�0S�P8�{��C?=� �Ė.gt(UH�'���'A�ďC�P�(�9�w@蛰iи^� ���)��_�6��O�aPCRDX� {�g�k�Zd��ǒ7!�A�g/Ę �,�IT}�i��T�i�`��RQ����E��%2.���6�^�	C�:P ��Yf�9���ax�n��B���p�	?/D�Z�'��eg�(�bfR�hl�X�C�Y#(�v�Q�0i�6T�B��~��4�F�'��)�fn"�i>��DE�1flu���Y=�=S �"?� �^=;j)9� %?��zB)Ѯ	*�����D%6٢-xF%r�t�� ��q�4�$ۀc| p�>E��Y^���*��5d��>A�� と_.�(O��"��u��w�lɣ�R'��X����q�zQ�Of���/PmX��!��4��I9тʟ~@�`�b��;<�@��搧]�;�GکV���V�OY�e���y������\%��%٨uH�%� OZ�q��ڷ$#� ���?@�|�� �Әe��8�U�F��`*ϥt�<�[r�#�@�c �& ��º!/�c��P�z,[�/�6y�PA��M�a,f#>1bO�%����"�
�ȁ4���<	���m4�Y�=��2��T��?�ƣ��!��O?{S�� 9��[��W�`�P��x� ���k~$�HY!}�yW�i�"|�G�S�>��ǘ�8>B8a!y�<٣�ֽ?�ȸc�^�Q��$�B	Lw~r�֝L#B�K�'��aaA�1�����$�89;�d,889��6V�MV%٘j �]�NȉQ/V��
�'�@�0q�T�"�\-��f��Ezji���D4( d�:T"&ʧCf�`@�_�Zl�ل�;T���EG����̿MH��ӁŽ�oZ60�^���i�)��9ҥͅ6 ��x�pA��R����4D�����E�Q��W�E�B�Ra�>��h�B�R�	דha��1��� q�
Aa�.�~���ɶܨ�%|���ȑE��]~`��p�]4vB�pd"O���Bl�B� ��R%��%j��鉖/�Dh#��ӹ:`(C�V��lhd���^��C�"����b�ڰk~�jAO��A���$��m��">r�ߡ���'�`E��&*���B�_*I�pZ�"O�%k�$���C�L��#bS���'�D1���m��.=
V�O��G)�$��)3�Q0&)��X�x��6��5ّ�˒ �h-����[4�kgKs}Bc	LL$�ڦ�,��dʯl�<�s����Rf�k&H��x�L��ōgܓC��� �$A!�CHXYtd	�n�nh8Pa]2t�b�3��'B�(�g�s��ɪ�� �m�@,*�'��H2�xR�Q(Q%���*::�s�bZ3�H��U+MFɚu���_d<Ȩ��������'"��䐚X�H ô�(�iܴ}��P7�i5B$��eNp
�x4��Gbv@S�+U`����Hq�%�?s(ܭ�u��p�T1aB�'*�1#�'�\t�j[	*�f���K\�Z�Y)��D5~����a�9M6�D��ぷ���5	3�I�!�xB)ТR�)C�dԁH���"��A.��O(XP�-}r�T2G9|7m@� �|�ḱOv���d��1�I��V�l��<xpd�+mD6H(��'��sM@<t�lp��,�%��Ҙ'W�AӒ>���t���Lɲ�IXZ��%� ?0t����N��3q蛶q�����mH<�����)"4�T�7�8 0���9[�*��MsU�̧c�+1�0#CL�s$��
����5棗�5��p��
W��B NR�0?#!�?YwKȡ�x�h������ ]q�8�Kɣ�h�*f��464,���Q��W3���I<�h�Q=��VcU	��8���c�'�̸%�>9�̛����Ǥ) XhK�);p�.���e[;/H�lڂ����ҐC�郈?Q���
˓_�����+�Vo0P⎔��@�̓k>�bI����c��M4�ԙ��c%�:T;n�ö��p���"��<������S.L����l�CV�C�򌭱�]�t�t�o�-9H�tJ�4g� 0 7Y�H��X�
��1��*�\cL�!6'Z�o	��F�'��"�S�X�ad��0���B�,!�+@9�gʍ�t7�se7����	�{���	�3�����/k��'�=���[���0�۟~]8Q���M�G0"�A�g�5�?�ק*�vW�{���gK'd, 0Æ�;��T��Щs�T��&� ;|���H�>���Jon��Q�Y <<�	�
������Ɯ\՜��C1j>��[g~���X4,5�$���%�ubH<2��E�`@3�ND��OR	��cH6�6�j��� ���i�z˚'%2P���T]҄R��ƒh��L��*�u�L 
U��5�+O��i)'ɒ ���l��Ѱ>qY���#,����^����Dl�t�1��D4��|��M�M)ZE��BV'b\�,����T6,!�'�r%���5��v�ݵ3r�t�����!9���j��
y����9y��$P�b�0�c�ҠC��#�aY,2kFR<b�0-z�L�2f�a�E�'��!�d,�&F�6L�/)2
��Frah&h��!C�����y� �	�b�V�Z�L�--:9�OJ6J��sBZ�s�X���@ʌ�l���%$�'���TJx
�@��s�>mLpӤ���R)! I��ԅ)I�(z�N)�0���:�P|��k�C�RV�G���w����GG��=�|�=Q��I�b��;(�x"N��+2.�[�b\�N���5�Ӭcj�����Q�������_�(�z&F��k�.�Y��x�(�
I���c�44�膦��O��b��Ak��i���P'X�h�y�U�xㄩ��(eZ����1#�1�편m��Ҧ�l�=sb��d�����yT(R)��\5H�؃�0߸ʕO�"aRx�Q���}H:`�U�(��B�,\�V	�kTĈ��)���Z��U.�L��&���M�B.\�a�N�qi lOޑ�2)�;ET$�A�oǳ0T��ZH��6Q� �7�X\"PY#p�͔M���	�9��4��5v ��+` ِ��&�m:u��0>�C`É/� �z��7R��� �9Yrx��Ɗu���"qe]�L8J�ѡ���iR��<iEF�<&��&I�s�X|���y��("7BO,;Tqs��x�����m{D �f������
d�P��4x�x�fΒ�CfH������p���)�<١I�*�"|��O�hֲ��$�QG�k�t��Q�΁Pr�Ԣ����H�RD�?[M�=J��]>�j�;D��<�U�Oz�C�K�vH�yk&�.a��D�U�ƣE�x�"1O2mv��Rv�L�\M|��*��="�YiT�"��&0Y�$'��a�|ᑑ�i����hX���D� ��.f���kA
��w�<���d�2��T����|��벮��h'��bDӚ-G1����9E=+	��P.�}��n۳����NP-Izpx	�J�Wy��O��+)L��mܴcba3��81��%�	�dB|��������~�r	iC�3fI�ܴX�6��;��m9v�M"3�\��𩇶g��'�ܨ2�JåҎ-��$uS�}(�}R�B/0_0�Z��]�x��'.��We,� �S�%hP-�с�=b)y]�ybP�dT�aO���N��P�p���ۦ>lD����[�eTDmAGLA%ǪM�CFΰ=��N܇=��H�#	�ʝ�6	LIo�|��;O�p�ѫݛhХ�pN݅H5�+'Y=ڼ��5f�Ȳ:沥afʛ�6���6+��0>"�P���3ElI=;<�-�u�\n�@�[����C#� [��%�2žqV�Dd�������@�Y��/EL8��+΢=��9��-�p�l �瀖�(&��Dx�Y�&|q��K
fa��B&��?��#�����O519ܙ��\��x� K/L}�P�kп��0�E�ڍ# �ԂTGu�c�Xa�O�3������ n�� f�5Qf��:G���)�j-��֎�?�����7�8	�(sG�Hm���@oK���x�ќ}%8�w���1��/�-���ɟk'�1:��Y�<�n ��`ޞR����A4c�L�@U�rؚ��do�2JQ!��A�{
1���Q>rp!�O��T��ڵ� �K�`�	7b|d�K��4�Wn�ɒߊ�1����5&2��F���/�������e����ɍ�~3̕2��!>�6�j�O
ܙ�3�L9ac*�7dC���<� �uq�L�l�Zm)�̙-s.�`S��a���h���'6̸b�i\%:ݜ<T�؆�2�b(����k�A�A�<Yvh�Q*������'yޮ|�`ŗF�<AWŜ$fr틃ee�B�Xx�<�v
C�=+cZH��:�j��5<!�D�=��Q�"-'C"Q����o!�X(U
*!V�b1�܉��T0 !�ګU,��
+e*�m�Wh�Y�!���c�@�2>3�T`�"t!�$��F�@�Ƥ1�b�*� 2$!��']`!��&��<� �9�Ք !�$'3�y{$��2�Y��!�!4�͙0�I���AD΃�!�DϺT��eDIR�S���9�1�!�D�4/\	�5�?^�����FF�!����e8u*ut^�p!�Y�!�D�"#�v���K��zg0=h��U9l3!��C��:�W�;H��R�%ݽT!�$��_4d�i�B5�8�C	F�!򄒬F^@`��7Mf%�6�R�(�!��Y��� `��B1�P�
�?�!�DL(U�����6_���kG���x�!�$�E��JAm��*~���7b�Y&!�Ĝ�
3��e
%Fq�&��+
!���4���0�ÓTp�rg �?O�!�ĝ/\B����㎈�D�80��}�!�ę�0�P`Z�A�l��4�!�䂉J�M�Q7�9�a�F�!���_��dW-�9��үQ-Zy!� I��D�
�Э��n�Cj!�Zdt�z�J�� ��Q`Vo_� W!��*�Qd��=[�v�z'�*`3!�S�c|�2���b�p��.;Q!���"�b��q@ʅr	�%�X�bA!��z���O�\�<�'�&;!���"T��K�0
4��`�3X:!�Dm�x�$�ZM�m)a� 8�z��6� �#� O�S���:s_0��}}�@-��q�5ʆ.yt�	C/D� �S%��${
� ���6�l\i4d?D���.,4�:%,\5<��9�1g<D���(�1*����h��d�b��:D�hp��	#t�����͖�
ڼ	�#D:D���1�˝G���AAhU1�Jŋ�b6D��1fƁ�Z�vtr�g��X�v���0D���B�J��(!�ڋj�F����"D��Z�X�p�����x�ᄋ"D��b�l�>���e�֥X�&}��. D�\B���F�BqkXٶ81 �"D���W �v�|pd���w��`2!>D�k�Gߺ���Rv�&I��yzf� D�$���֋���B�+�4��ݐ$G D�\Pun��p�@Q�J�4F�~�:��+D��Ps�ĕq� �"�W��H���'D�� �	��n@�E�Եtd`�hqI D�Dȅ��=+�LU����vta�"D�8E\�Y��8�C�?P؀}#w,3D�����7^TH�#M�	/�zm�5�2D�L+6N�:MA��$�� ���["a5D�p��-kC������7*s��j��6D�@��i��8��@�P�Rc/D�P��B̾0j�4w��~�j��E#D�x7jU�.�,enO�|���$	,D�dy�@���@�2"6Iڥ�d�?D�� b���C�'��i'��hi;�"OL\V���~A�u�� ��xEy�"O�a"�g���q��V#jر�4"O�s�	ŸFizB���-����"O��0N�	Bx՛%IS�X�"O|� Qnʉs��]x���D�|U��"O�a�ӎ�.'L�af�g:�kV"O��p¯E�+�Px'@�pG��C"OTh"�����)���-=� "O,ȡ���8�~ ��b�m���"OT�R��	
=Ty��,��Q(L9�"O�)"M_�����K',p��"O��Á�oJ���@NI?>"�"OD���H[Bl(%���|��j�"O��XD�#<��A�����R�|��"O�8��gѾX�	M�z����"OF:�(��9��PSv�;�P`��"O��j�.8��c��0b��!�"O�tYqA�%SR�B��1-B���"Ojt(Gb���'EK?W/�̩�"O��XQ��3״e�JX�t��d@p"O�5iD�
�
^��v�O%-�*��E"O��#rʗ|����N1Y��!8�"O��k�DBx�u���)����A"O(��F�Լ��r�웣���"R"O�
��).N����jA�YT�yIR"O����LP�*��š�$�0�>|��"O4���KU�d1�1ٗb���C"O��%m��#x "f�V8 ���"O~��T)j���r��,4�$9���F�����k�"�D��ũ�`��u)G��y"GG0�Ƹk�e&l��X��Å��y���j�`ibt�ǈOpD0�q�=��>���y�lL<@��D��D)����ʒ�y�'؊T��r3�Q/;.����!�ē�hO��>Ir5Ō�g��`��/�z�Z�"OT ���@-����O�;�2���i!P#=E��4�&!��!�p胠䃱>rv��ȓ$NB�k�IT\��<�ϙ�
\ȇȓ;�trg]�!����"��C��ȓj���o>�!��yHf@��B�x�Y�A_�l}��X���a��ȓ)u�A�!�D�	�����HJ/he�ȇ�ʈ�� �ǎS
2�?.����G(<)ɂ{���	�2n<� 9D����`A�)��h�§�b����D+D�0�'.���ꂥ*��K��)D�d#���Y�ހ��I|��1�5D��02��0��
fN�F�9i2D�yc�ʺ=^��f��I����L2D��I���5���[���*;�޼���/D�ԨF镟��]�� 
���``3D�ܣ圣fJVac7c�4q_tt{6(3D���4d����Q�XZ" e��0D�<�a8z�@�Z�1::���!��On�=E��� ���Љہ-�xZ �"E!�D	u�*��C�
3{�:��
�X�!��OR6!;Mcg4�� �G�L��|�x��P~��4�R��W��qpb���y"�C-w�Z����%��� I�y���#A��R�k+}��]��	��y��U�f'j��RaP=s��CŃ+�y"�N�D�E��M$g�hI5�q�<q!�t�8H�1$s`�
7Uo�<� �yC�B�BP��z��	;�,(:�"O��� �Ȣ��퉕�F�Ga<��"O� �jD�l� HR��v{�i"O� ���-5�y"�*�B� ex"OjT��[� �h��SI+�.���"O2��� �R����G�a�Hi�"O�	��Q
��зD�(m|XQs�"O6l��l��=�1�&$*p�$3"O��z�f��zG��d��13k�h"�"O$mSU]�+�pxC��ͥo9X�iR"ONP��!�5Y������jz����'����?���h�Y�<��!�
�~�!��h�ȢGV"l~<-����%xT!�dR!3�܄҄��u¡�A�\OS!��MU�yۢ'�|�S
^�UB!�d�&V�:��# [��j GʼR?!�$�1<$��G�_�g�:�+uHէ!�d��+,�=��P�os �A';d!��F�T���[��_�`j,�5����!��<SBH�:�ɼs��GQ�kw!�$�L�uhW�@��-�t��Mr!�D bF&mB���\��#T.Ær!�Ě*_z�l�m2*�Hx�d
�KM!�D̄h@ Q��"\8J� ��(�sI!���$"�J��z�8��Y0!�d�281& J��32 �ĆF�$i!��X�``h��bD۶Y#�i!�DѺ;�!�D*PR1,D�5�uH��(�!�d����q�͓��0(�l'>�'nў�?وbB�#q� ���a�D�>���#D���%��T	�(�b�_J<4!�L D��ȁ*�p�Q T)$��Źp�#D��s��N��i�֪Jbʝ
G�#D��8"a��o6JQ�h��4h�T��"D�$��,ʂ-�
���L�H�L��!D�)$$�v�B���U+s� �I .>D��#0�	G1�<����*|J��.D�H��MX���0s<�&�PWD,ړ�0|Rg��s��#'M�����3�T�<)���_�&@��-s�<�K��[�<��H_�1��0��ߦ7�h��!��b�<��!W/#O�ԣ%���-������^�<�pќ2Іt�V���0���P�<!�	؄?�  T*G�n9�M���FM�<W$�
ϴ�Z`�7=�TH��K�<I��]%��<�&睴�P����[�<!�d��n�C#lOW�*����E_�<٠� C���Z���:x��p�<)���q�
#TI̬@����k�<I���dD���j�)A(�R��e�<�5b*T��Uc �Q$B&9���W�<�ń��'`���H�(!P��$��j�<	�� -1�8M0	ی/�Aa���k�<�4�[�p9n|�6�݄��|��Lh�<!�߭H��Ԍ�9������h�<�a�;*��0cS�J��5��|�<1�OR*we6|#FL�w$�&O�<q !�8)Ś�`�i��&��'DI�<�O
O��!��`�*��+���F�<�t�+L�ah#���d�B�+a�F�<�5�X�Tu�|�a,��d���
�I~��'��x�E�� Ԙ8J�!ʈ&e.4��'��� "�+�Na�oQ!�>�9�'��)UbV�YE)�Ԁ��)��� t�D�M���̃��Y�;�q�R"OR���j_.VC0Y���Α8��yp"O |���܍iM�d�P͎��`]�"O��Aib��"v��6z$�Ȧ"O��!�;�F���A�==a���"O�͚�)ս`j�%���Q+!.� a"O�0�Iޖф広(T� ,�B"Oܵ�H��P��!�AhP�*��"O2��$)/��ib�!�e�f�p"O�ڔ��2��%��K��p��0"OF\�!�
�`��CoR;��b�"Od@�ã\������
9�mҀ"O��p*@�|Gb�Xa��)�C"OP�q֨��^�, :��\>?"� c�"O��1uB�u�F��r �"PS"O�;vG�`��:ǏU4 A�"OzMc�h�oTY�@U'1e��"O�=@���,7��c�ʞ4	zD�"O�����E9#9��{�
ژF�f�{F"Ob�;eU"Ru�I�(�wՒ�"O�0C��'�F92��\(8u^%zd"O(�#�A"Y?f�
�����d�&"OB�*a����Ze�À�]��$�ȓ(�Z$
t�	�T0[�;6M��X��a� wh~}뢩 �CLdT��!�fH� ��?ֺ�2�h�0��p��϶��R ��Z|1j2dlP�%�ȓ/�\�	VOmunA��?yΔ�ȓ ppK ��Q�lh:���f�����1����dܓKД��INzчȓPd,��m\�%J:%�5�-�Fɇȓ�T�JpX�i�ᙵ��	_��ȓf�*���H�y;�A�f�i�<݄���M9�)�0VC>�@ϖ �RY�ȓ1�DʖߝQ�Vd��0e�,��ȓ4$�93HW�)�x����/~�����Z6��V�F��Q���,:�
��llDڄLޅr�H0Bu�L4.>���ȓ"p�Xa��9`��9u���E��X�ȓk��)��Ò�m�>G�{�o.D�л4fT1J�2u�"J�4�J.D��J� /Q �;aJ�N�N�s�H2D��q�W7;|�#�F���F�z�m-D���we�7 ��H��(�W���`ԋ*D�t�S)I�\w``�V3|��["+'D�X��-��l����9����P�#D�p��(2��Yp�ͮM�j,aC�#D�d��鎛"��3͕"j[��$D�D��,@�Kw���%@�Y$���/.D�p�0/�3u�D�"��F3�}a�..D��[���S$:M�'��9`�.��7�(D�D��E]�+N&,!�L�NJ��$3D���T�|n�C®��yh�2D�l��晴
U��ҡ-��D�F *D��K!aھ87�H@�Ѧfsz�k5�)D��Y&oW�i����$Lѹ[�:����%D��ѴH�d�NP+̔�B����-D��jb�ԓ),Blۂ/�{�Y;�*D�h�t�^6f!v��5�P�I��r1*D�h�Ѕ��n8�pr�`�}�5���'D��a�Z+F~:E����NP�5ѷ1D���OI�Y��X��>��]�wF0D���CiZ�t� g�Laʙ�A�)D�49��Sj}�4��n��eS�$D�� H�GL�NB�bT�6]�"O�XB쁘U�H� �OK�4�� �"Ob��N�`aS��=��#"O�H���0.wn��5@���@b"O�M��#�_��LK��z (P�"O�H���Z�.4
���mO�<��"O�=(�c��7W���5NZ~<���"Oh=i�ٱ�|݁C��WN��@"O*�8�l��&� �pn;, �5�"O�=:�D�r1�d��ˀ����"O��C�˓�86��f۫"ዟ��y2
;Z�t` %*ۓ���*�1�y�A��&��-��ƔR (�����y" +gN��) � }@jD�yBF��j������K�t�F�)"���y�/Ѳ]� ���M/i_����I��y2)17R8��C%hl��������y����>1�g�]�*mrJ��yR᝔>�pb�Ф }�Уq���yb �8���� 4s��@ �yA�2f�lDI3.�$�V���$��y���+eF.�
f��3Bu��#��y2�2ln�� N�)\`�� �y�":��w�/�ȹprD��y�A�r<2�Z�ɏ6����aD�y��RQ�`��$�_�T0��NA1�y�C�5#�~��#�
S'>�u���yB���`u4��¨��Cgq{b$�8�y��&oB��6���h���y��7odI�l��9jyqA�^7�y�θ=�ȕӧ�д`X:�A,P��yR
�6g4�X'�R�d�r!�ׁ�y��OF�Z�����{�E���� �yr)^Ly��q7x��Qb��,�y�b�L v�B�o*RPHp�H��y�l�2=d�Y�w���a6��L��y��E�s�A�wAYK�p��6KĴ�yRo�&ww�E'�E�K	R)Q�ï�y�P�h���#7��^!�E�؄�y",�
?/��2/Ynt����F��y»�T����`��t@��Q�^���ȓ
>�$bsCܬN�*�+�I�7_���ȓy��P �n���¢%�����>�x�y�%[�G��!OA�P�1�ȓT�*�#*O�3
8sՇD�UJ����%�����dA�;������_����E���т/E;j��zEJ�1!�ȓP9�= QA����8�b>���ȓԄA�ϭ�LXI�˕X���=��]ZVHht���W��K�T��uiL�a��6?D��8�*	]����s%�qր�dڢH�`�-�
L�ȓ�*1i�iP6\,m�उ�L��I��su���W ؔ�����ʂ�-��=��F`�"� ˞�T�!�#L�E� ԆȓwN�QYE�I�C���'���sDJ��i�
��	sW�:V �ȓ	3δ��F�240�b��V3N>L���eT �3�G���$h�G�X��m*��IC��-\x�㠀�N�<X��9����"#6nƌe��.o�@�ȓ(sj�p�˖��u�r�B�	kx�����ʖ �DU*t��-өe��ȓ�p١��ރ6�xB��L
=-&���S�? &��5N��?�6��Q)x�	�"O�e*'����
�T�6%^�qS"OP|C$����牛}��3�"O4��)I�W ��#lJb�iU"O���d��,	rQRˑ bh�"O�vB��o��,#���3���"O����/�Y�l��ӯƪ9����"ON��@-��y���Ң�]'B�t\�B"O҄��
�G�ţrA�!�rȒ"OP�@6$L����S��y4~�Y�"Or: -wv6D�� :�tp"O��,ΜzcF�z����uc�"O��ʕ,�iHe�8Z�$<qC"O��3"��*l�ֹ9�F�?x��<)"OVI��$�������K�3�����"O���B�yUj��#o�Nx�0"O&|��k�B"���h[�x}��"OtI V��-j*�s���si�P;�"O��ZQ���'�~ t�W3BTAx�"OBh��`�V xM��f���"O�˕�_�~V���VEJ"L�@DQ4"O45���U�s��i T�V�|���Rr"O ̙�lŉ-e���Ö�7w�)�"O@��BQ�O��
e�ҡHY��q"O�A��¾e6p�3��[� ���"O4�� kX:D��M��.M���"O��G����4,��$C�x�"O��z�d
�]��@t�A�<@E�&"O�M�5�ٛk��C<��ы"O�}C�F�&a�f���2��["O"ݳu�V�A�z��"E�.E�"O���F����i�3o�#�U"O�x�­��g�ܒ%�I�u[nH�q"Oлvg��1�Ο�/�Z`�"O�|@Ręg'�t���)���×"O��0���6�Ft�%-Ox��D1 "OZ��("	m&pB�J
%_�D�Z�"O�ѓ�ޅ"��\�k��~��`"O��j����.�+j.)���je"O������O�R���Ʌ-{���%"O\��˗�&�{��+9`T�!"O�0)�OHPz�I�_�ru�U"O��a�A� �|��sʔ t���	�"O��`��[<`k
�
�B�`�کq�"OP��e�1{�\H�Kҋ��9J""OB=;���.W<=i�	��n�\��"OH�ok�F�`$閻qXLs�"O�`A�j�^�	�B�D�
l "O>�i�蘤6��U1���+<P��a"O���"�ޛI�����ΡS)\q�"O��Łֱ7����r�q���٠"ODź�莧lL�i '��h�	�"OF��'aP�}b�$`Q���Q�3"O��P�bY6�D�����Ny�s"O�C�֓d�A�fFY7�x��"O�=*a��L:j2w�
T���v"O��SA�g�@93�,�V��� "Oz�P�#գ{�N|y��%n��U��"O����,�6< ��1���f$8G"OL��B��Y�*-	��X�Ua���3"O �#��K�N�r"nU�[SJM g"O�AJ�LX*(��Q�oG�^^.	 V"O��c�KH�� i�tn˶r]�@�"O�@�����LHh�Y͆d,\��"O� �����Ln����	 �6"O�<c�^�T�r����T�0�Y�"O��%K�z,$�'+\�KvT"Ol�2҅����Y��HI9���"O�%���8~fD��F�&H�ԓ�"O�ʑ���!�uO�i˚��"O�p���+�0�sO�8�,��"OȈ8'B�	h�����R�Kq"OQR5.X4�����\	Zt��:"O���!�?B䚀��h*���"O������*�b�;'@G�g\�b"O�|�7B"�(���.V�����"ObQ92�E����oN>Mi�"O �`�	�\V4�V.�,VjI��"OF�Ca���	�´{'H�Fj��"O����%�0 �G�[8A"O(�W���h�BD�Œ��̨�"O&dA4E#�@U0���n���&"Ohdy7�I""�$�D[�3�BQx�"OD<b���7b�z�K�d�.{�\ "O���/�(�L�)	�u��9�%"OR	J�HWJ�ӴRx���'ؖl2��S��l4��n�r���'X�9�EC��V1�G��1���'�$�aC�X���VNή]��k�'w�t*6a���f�@�̂���i��'1fa��I_�5�uz�gߤ~�p4�
�'��4���ک_�lx�Ŏ��i�%�'��|�!��.y�D�4N�6D�
�'|�yA'+���F|a�*��;�5�
�'�<�c@��)�B�H��I2K��h�'�Zp"��=IҠ ["$[2Hڥ��'2�"�,]�mJR��14�~���'��ĸW�uQ�p�"J@�Sf|��'o^I�Q��
L,xB���!=��r�'tt��ͩE�B�q�Q�
/����'m^-�2˅�{,X0��m���'� i@��X>E��䙜'��=*�'Bt3 �_	"hzB�!A�����'{�D[������[w�_4&_� �
�'5*8{��'S2�p��`]��j���'���A���1A��b&�΋W�q�'�Dd8��o�^M�	��{����'���U�=��|T�8
��@"�'RB��&@��|� qc��~��	�'���QG&ڄd���b�o,!	�'����7e�~P b�[�j�pPI�'�H�iQO�?+^�+DM'Cn��
�'�L!��K�l�����W����'E�Q��ȅs?H�K�H.|���'p(����s���dU�VQ��'��q�$�3�����+	�8�J�'� 1�d��Xle��.r�j�A
�'ĜJ�6pD��L��S6Z���'n��Y�ȋsKVU����)#�4W@�<qS��F��� ���.?�HP1@��z�<a�h_�5<���!'�qT��u�<�a*�.%�����mn��$�m�<��i��C��+�&��gN u�FC�I�M�Jd�A�+���so��`B�	�ks|	�G�'��Xr���|�BB�Q�R��T�Ǯn�axr�M�m�2B�	�j��%�ƩK�γp�jB���h[�&-����:-LB�)� �UX!E�gg�a��ꆧ>Z�	h�"O�l��G�7J�p�皢jBjػ�"O����C����R7,,��"O�%{S�͎:����(/N�k�"O2#�>c8�u0�e 8�,��"O��#J�*%b�B�K�Q|�z5"O�����H�ի� ���L�;4"Ov	������c�V�)��"O��s�T����[�R޺|��Z��G{��)Ql��)0��#h��H@X���'���#� M�:4Pa�傒�\Z���'�U��j�#��p��NW�u��'��HT���)Jeb���I�L�	
�'���dX �<I���;�l�
�'݉�)�+LH��� ��7S,�J�'���{Ui�*]�h�x�
9db�#O>��0�ɢL�M6,ÚKC�yD��?  �C�I  ���4�֛b�8��a��]��C䉎�x�S�ƨ=�,jՍ�7<�C�	�<�^���G��l�!L�C�I��N���n6	�y&i.!�lC䉭?�Dq���7&ڐhsR�ְr�|�pF{J?���.�(������7da3V��<���?����?y��	���d�P@
F�|�� z�I�o�!�X)��D�$��i��hߊw9!�$E&����inh;�MТ#7!�	.jvL�)e��m/L0����l�!�ۇbx0%�r�ܠI�xi* L�^}!��Ixe�hJfg�B���Hl�	�!�׬6�:a"v��NH$�M��:�!�Q> ��L8Δ��w���{!��)@�a("ƀ�Ch0$����!�2-Bl�T ��T�J%S�d^ �!��J�|B�9�؁�w�C�P!�O�l$QV�W�-Xc��@/>!��	wup����	�t����-&!�D��+W|u�"E�<�b5�B�_!�D�3�(�L� �R��x�!��H�H���EIM����ck�L�!�d\�Х��X���G'T!�4(�'<B���.\ ���1�
�^�T��'�2��b�60_Rer&
�X�'�&�C�g�1��q��]"x$�C
�'��Sŭ�y�Ij��9m�A��D:�'[�Q-#ER�%C��H���Tl8�RC.�Ä�c%�̐C��9��۸X����,e����p���Z/r�W�V�l`",z�j%�ȓV5��fS�1Oq��.�	m�C�.Ҿ E��&�U��f�q�B�		%XVi���')撚2��;,0��=��hOV�#�
0ֆ��Į�$�.���.D��[�"Ǝ�T�zg�C\8�ŰrH'D���	?T�Ќ!0�AֶMʕ($D��q�D#Fn\P�I_�@���C0,-D��Z��F"vp=��X:=|z�f� D�0�u$��o������V'X?xq#"�>D������	$�U�0E]�V����O֢=E���6R��ڦ,	0_��pTc7W1!��2p �1���$��J25!��0����"��к�z7�̥,.!��,^w��p%a�>[&���W=v�!�Dˎ�<��UGS��ى�n`!�$��l-;�JOj�a�P�C6!�� �$i�
I(M��D���2C��Hp���O@�}�T��=@2�T+WR����J�-h�l�ȓ'On��h��Q�H}����5����;Et�rōSr�eIE&�'4�N��ȓzkf\Z���0?wb���dޢP�@5��xv�Q�Ą�|���!C�\���j�Y�WO�o�(A�u�ŸagNͅ�J�&�x�� =fka!X�<�X5���c�'�| ��ڴ`r�B"@T0J	�'s�tX�I�^���"��g��)	�',�!d�����d�P�D/�X��'" a� 
7SF@�Z��
%kjp:
�'�
\��I�i@�3�]�"�%��'���b�I	�)`�a�,����'r`iw�ֶ���{S�	���h	�'��$J�O�?���r��9�؅��'� �Pǫ%T�0��W5��@��'�`9j��M)b����%[���'S| 𡙆AS�eaQ���"��
�'A�Y8�*�5�<�5@�gz�
�'�:�1<<���K��}��'�0�!N�I�Nh�mF�e��Ѣ���(�8�ډH4�ɂk�^Ȑď�1`�ЅȓR�AFn�N�c�Ĳe�*�ȓ�Nd&�B%�f�C�W	�v��ȓ#�@9�UN)���۵��F��ȓT�,��%��L��s���pZ�\��<Mbe¢��4�ࢶ��Z~��ȓ��qCpg]������>�V���y��;`e�7�I �ŕ@�u��W_��3�%�N=n��J��ȓk朐O"!��IPɄ�s&*4�ȓlInx"��R;��q���.W�P���6�
3��
|�b|Z��X�a�"���4�0��ō)-3�ɻC��$/��H�ȓ������q D�QȚ'q����ȓF�18�͎v�Q�� ��iX,4��{�8@`�"8�:�����ty�A��CIvE��\�Nn�jp�_�i�1��4�Z�Ql�z|��
G
y�����#��0P�#dJ4��~�0���zv(�:4@^�<�J@i�)�"+��ȓm��QIGAʊ)(�pI,�<)�pX�� ��d��$"�8Gm�6=x�E�ȓW�ȶ$��H|@���R
M}���ȓ=�t)�O��]�� H�{"O��H4������H�� �FT��"O�E�&��?o�J�+%IX>���a�"O�ts�f�5Y�n�c �N�b��U"O��@\�f. |0��s�H��"O�EY�@�V~�ECBOI���q�"O���F�;gxAWÈ�^h�܊A"O��  �-�D
#��r\���2"OJ��
�rނ��IR$<?y��"Of]Q协&��t�B�k>� 3"Ob�����m����ߞO��D�"Ox�9$ZF��%C`��%,�|�"O�8�i��l]�ف!&>Qp�p��"O� k&�˩L�JX !�Q&̄���"OZ!) ��y� )2�$O�zt"Opm:��(�D�!J�TQ�Z#"OzM3��R3C*a�oD�I$"O��+�LL��`�w��t;�"O��������,��ЏC?u�0�1"O� ��2%�Y,tjE�&l�����"Ol{(�(B��x�q��)�.��"O��'��-F8�IY儇��@0�Q"O��l�2jW���Ea
�Y�6Q�!"OހqrKºi3�b`Y9��Y��"OZ� �m$�T�"/C�c�(x��"O�,I�P�L4  ����P�#�"Od�A�#�����¥Z�g"O�5+ZH��&b�'	S.��4"O�;��/0��A�n6.`�c"O*�;�*��5E�Pps X"Ȇ!�"O��� �% �>M�p�ɴ ����"O�`9��W�&H�(���$J�`đ"Ov%WON2ԴУ�F�X�$�U"O���a�ވ��- ��/,E"���"O\�(��D����2��W�5���At"Oؤ�rNO�hw\�����h0�Lҧ"Of=��N0B���s@ѷ=,���"OP�RDXCV�� F.8]+3"O�����"�:�nؑ9���G"O���� K"2���;��۲w6)"O�h0�E9UF�	���04l��""O'	Q3+k���l��.�""O���e�UB=��E�	�,E��"O�ATE�Hx|�1K�?b�,�r"O�1���|uԈ�rI֩C�l;�"O|ms�Ä�e�F)Q&���Z�~���"O���l�7p��� B'�<>��)��"OH�s�gÌr$���D3e'��²"O�0 �O�y����d�m&�	 0"O���/D��L�5d<^) �"O�q3pK�n���0��Op�p�"O�\P��F� ���جbL��v"O�<����3!��	��H�'|��P"O�E���/?m��8��E	h��4ڢ�'!!�d��0 �kP�OB��2�)#%!���V�zk�
#$P���q!�D\�xnA��Cw&`#+	9_!�_)K�.��F�~b0��j�;^!�A�J�z�:U��1Y��jc�U/�!�C�*|��)=I�D.TA!�DW+�~i	�%�a&0EY�o�^1!�䘮<*� x���<0�Ը�����!�$H .#9� N��z,<���h�!�� e~5�#�M(ܨZW$PHL!�dJ'0����E3J��)`��<=!�$H�2U2ʔ�_ �X���ތ5"!򤟧/�ҵ���HC��@&�!�D̤J�����q��D!�(��!F!�DQ�<X��O�;�ꍨ&!���Py�6��!�7��V[<o*M�ȓtY�`�V.�@�0���EjpT��+�����b�'K���TO�:�R$��=&�5Kl��T(�ՍQ^T�ȓ��4�S�ɘ~��g
1. P��d2έ�Չ�9^�i����p\$��aIv��ȥ|�����j�?mE&1��)�Ԑ�r�ի}��i��)M=W�RQ�ȓ44\�2"ϱ�������8$�����o��wm��*|��g�6pW�T�ȓqz�i��҉Y�`	��\�ȓҺ� ��܏���6� #Yn��I͟�$��D��'4n�Wo�:Z(�9�"��5��|��'��Z7+�-L�DxY�lV< �V�`��� �d��L�sM�1pWB�	B�Ѐ"OĬ�4`�i���TAR�3a<��3"O��YF�D�nt�A!��/Z�
�"O�4�W.�x�p4c���<�ek�"O*�Y���zNx@q��48H01�Y��'Eў�Oָ 
Q��$8B��v�6h�X[�'�-�1�ۍ�*�����X�T��'j4�"�'��B�h�"��U90�@�'4����I�Bxx���T�J�B�'��ۓ&�V��0S��$��	��'��=�d�_ C	(8҂&�x@4ܺ
�'5��@!k�.qe�}�B�@��3
�'M�H��a]�47ܡ!�E�e�H+Od�=)����i� ���L2��h���D4�`ً��'D��d.H�}�r]#4i�H��[ud3D�P����X �lɂU��񣨟f�<��I�Y\��"'��>z
u���c�<��M��6�:M��B�gc8�괌�[�<��C�j�A���/F�zQ�M�R�<��%í{ju�W��H����u)DM�'�?E�uO]�
d���J�%���n%D�`K�h̄�∛����(�(a�� D��j`��$I��B�F�R��K�<�T���[D��+c)Q��h��MLf�<Iw�O�3TP��*�<��TL�_�<���Ʉ;HN,�AB�q>٣�XZ�<���T6^�Pl��ϓ�긔[c��\�<�6�����w�'8:$+WkY�<A�.>=��Ps�%	|��\�<񗊍�M����L^69H@�b�T�<�g�U ƪ�7�t��tRk!�B䉼+z���.Q�)Ǯ��%����B�Ɍ�-���/[������JQ�<FB�S�h�`)��a�y�`�`2o�l�JC�	�"�4�ԃ��_ j,�� ̜J*0C�I�>D�	IY�$���՝��B��b`��1������P�F����B�	#*9N�s0([<w��hZ7F��)�B�	�e]�hR0^�"��83яqKtB�ɱDw��:D�W.qN���I��ozC�; |Q�`!�0*��TA��T6�B䉀'!\U�����8��i-8F�B�I6ak>�qr�۠r^�P�eK��LB�	98�4�0�E�R�2�Y��>xB�>X��ȓ)�%�4�b��ӷI8B�	5g�J��2W�Q(�	 h�7��C�I�7s��6���A+�1Q1J�)�C�)"c(�q MM�)�ꡰ��D0����Op��yb��C�^U�J��x�xM�t ���y�ɼR�,�z��!hX��l��y���3LüPI�DV��~a��C��y"��
6IX�0u�[�s!�2��%�y2Ɓ���F✜����^��y�%N�h�\����)�]�r��"�yB�R�>N<b�,*>��"ȓ���<��$�f���;r(�D�] �E;!�$�PbAP�l�6E� "E�!��iya�c� $�3 @�	P�!�K'V.���)ʳ7��q/� +�!�S�1TBɐǍ�71NT�v�0N���Kp�I3�J'���	2���?I��)	f�(���A�f�<�8F㍮p!��/2V%�v @�Z��i��8?d!�$ܤ��مL�7'���z�NcY!�� ��h�CY�Nf�Q�`H�*8��UQP"O�����H�=|�H��E��,��"OZ=p� ���d$�9|x
��"Ol]h�`�-T%^�c��YuXxF"OeI��+h  g N�Ar����"O�	1��*.��+r��>)�H���"Oph+�`�(��vo5,��E�"O��P +O$c���0�>e��y0�"O�Tr�*�>}��`�s�S�_��t��"OB���Hȉs{�Y�j�[�nt#�"O��F�S�4r>��+�	L�D��w"Oı�g����`L�6�C"O΅{d�IĹH�JT�x��S�"O=�aC�p�s�hK�~�D A"O�)����
��سs��)f"��"Of�x/}
\}�2&�#���P`"OP��e]
������8��\z3"OX���w�N�
��Ibo��a"O,�!�Ɏ�|��!��d\:��"O����V��7��"B���"O�H�jV%��	1��:=��k�"Oh�
&n�0|���dd�.zt��F"OP�(RȉE%~Q:�Ϝ�ʰ��"O���Ĩ\�8V�=��A�
n�8�ɗ"O�E�p ]�S��Uڕ��y
�Q�`"OT��C��-�>u)$�W"�^P�"On�2
6=}xe۶C�� <>�0#"O�Ħ��s�b��R僝[� ��"O�!����I����P�щ{񶥱"OFܣ�Mܙ�	+��&�:� 6"O��s�����K��Z�?R�*�"O�U��P�Z���
��+d0�A��"OZ�
G2>�'
o?&l�"O���'V�Re��a�PK�X� D"O�� � 
���p`H:o����"O�L;G�0\�H)��͉��� !"OH�Cb�E�Y�������E�"O�aڲa��*Hf�E�*x:��"O,i1B��#7FH�R��ax\(�"O��HՏH�J��������2�!"O��hwmC�4:I��1+�
8�Q"Od�i�k��H��a�#	k�`�0"O�(�QȈ�Z�8��U�X'LS�0q$"O^�9���Eڈ� ��7f[9B"Oޠ�a(�u	4�Qu�ǰ>ޔP�"O6a�4KȪd�\����ӅD6�!p"ODT��M:6�<1i���F]��p[�@F{��	�/?4x[u�R�?j�]�jݱnT!�df5%H���R��p�S�F>!�ӒKTa�Ś��>�s6���@�!�$O?�D��刅>,�����4.�!��͊1T��Ba[�p��<�f�Y�Py�I���a���e�"��QA��y��c���"2lU㕨G'�yR#�V#� �co�8.9�ԣ��Ӽ�y�M L^�Xw�WdF�!5f�)�y��Ͳ\�L] ň�]���j����y�'�p�T�b$�fdr0p^��y"'M�"I���oV9b|�̠�,��y2�Iq< ��A%D�V�����y"�gU�3�j��LR"�!E�T�>��<y�����<yK~W)���Ɖ>��4�Mѣ�y�Ȥu�ĵäۧai�i�ɥ�yBk�fN0��`
Șf��h�U�?�y
� FU��!�&:���:�b��2�<�0"O���5*���@߸4�@��"O���V��J�&�`o|�,a��'wў"~*@J�{��Ӵ �0��K����0>%��?'�����mV����K��GT�<9�-@�gNB]S.�4؊d��H�{�<i3,J��E���F
�)K��Yc�<��,��a}�<
�b�	>e���K�[�<���a�#Gk��4�D���M�<9�ƽo{l��	X�B��@t%J�<��!|WZ�v����T8T�ş�	П�&�"~"4!��.�D����T0��Q.��y&@5B4NԉV,$~�5������yMڵH���b@��q��̉�@��yr��A��P����m�n<�I��y¨��Ejtz`��]ajis����y��٥Jm������\l��)�a�'�yr��%�|\��m�\R|�QE�8�hOP��	�	�*�wnK/g��q�iN� 	!���7�FA���[�l����W�!�$YI������DD Xh0�	]��!��J
��u
�Z}sE��-p!�$� >��=x�+@� ���=;l!�d����8RGT(��[A�ɾF\�'��)�$/זhS�'��8<=�Q����O����A�b�FPz��$���b�K�I8!�݉Hh��l�*UR@)Z�D�Z�!�d;n��kPl�E?���1�E*-�!�T�f\����(��!�,��Ζ�F�!�V�~C��B�`T���K�y�!��*YL�Y�VϽeSX�t �wa!��̹0w\�Si݈/�>u��ȯ�!�ͯBH�[�.�(��ѠEnь�!��k�G�+wP�I�m�	\�!�$�/}r�Mᣢ�8"�i�e�T�!�$Vb� $a��ٛ_ФH����0�!��ǟ�"e��*M�fÞ���T|H!��	��	@�Q:?�PĻ cB�`7!�d�1�]�'�_>�8�J��0U�ў���C���jqf������C
�~�FB�	�p̦�P��Z;wj�d���S�B�@B�I�3d�څ�PdM|`S',P7L�.B��	�<��ʆw�j��EPB�ɧRH蹳� �.苁.��
�.C�I�rI6X
����FK@��$��+4ZB�I/Rd��B-Z.H(�r/��`��O\˓�0|"�&�4��㇂&�,x2�No�<�e��s�<����S+v̹qL[h�<Yt�F�(l#�ʞ$N
I+��Gf�<yrA��CY���1�N����}�<�uN$9�գ#D}�0)F�7T�ؕJ	���(���6a��@c�%D��a�l�;����D�kZ�M��"���O���<�M�q�kD��d���H1)E�<��I���$Z�ϙ���K�C�C�<A�ܲe��I��іr�f�s'�Gu�<�	�,v1��%%	 ��m���x�<�&�f#4��$LP�~��<�yB+6u�D�aǊ#: 9�&�ĉ��xB�b����V��\���T�
�BT�p��R���ӓg}9k0�%h�y�$.j�C䉑7�V z�FB=�Tx��f�\UHC�ɮum`�����H�V'�$(KfB�Ƀp�aZ1FZ#	?��x�G�BB�)� &���dD)!0��r��|6n�Z&"O6H@�"��y�t �cP&��!"O j��r�����X<'�,�֚|�_����'�2 �`�@:���G�C��/Qi�������I�s*̩,��B��*�`���/�'	ʺ���T.{�B䉪"�����Ϻ.�����<�B�ɖ7q�肷LT����@dS�B�3;���䮏�X�H�RL���B�	5Qyb�AWM��d���JE#GU�B�ɏ����2 0�r\��O�ڔB䉠e��k� E�U@؋�� �x�B�	�>�Ĕ2H�R�����%�nB��`����A�	�y���@+��B�I<5��U�`
�3K�ؐ�/�]^B�	�] �y�MH�Fp�`����e�:B�	Bfܴև��{���a���c��g����m)�d<��I9�h�R�K5D�$Rqh�4	�N�B'���f��7�%D���tc�}����ӖV�@��aD?D���&���"��ؤ��+�4U˰�*D��ql�_n\P�ŏP�U�a�v'D�p�/FK�!�IΆe�����&D�\�����N=B6�ם;� rs-��0<�%��|�S�f-r|QbL�a�<��!&����Ɠ�hhCЩ�v�<YEMF�[�v)��>�H�'�t�<�j� $�tpaN�%=���C���V�<D��A�
=rt��;b���֎O�<	�U>#�@1��b��'	�+�ƍM�<���B";ߠ�Rw�d!0�#�ȘH�<B�Ŗ	��Z�l��'�L=���{�<����2��i�U�,(��jw�<��.��E] �k�"3��H�l�v�<9�!C?wth(iEJ�����y�<��o�!-�
퓀ϔ�^��Đs�U�<��o�a��(�r�R Fn��
F|�<���_�X��B�}�,����a�<�ͬ)�>����J~��f�f�<ٗ�X�A����/Y�sP�;�hLf�<a������q��L�>�αKqJB|�<���m `$�L��w�d �B��q�<Y�cFCOf��/U8:���k�<ɡV6�hh�F��Mh�L���Ig�<I�K��/vԨ��,���b�<�k�B� U(�$ؠ
žh��v�<a���<'d���aCuDV�*Q�o�<1Ӣ�4�J5��'?��9sjUa�<�P�kI�u�".D -FQh�cPi�<��#�l�je%��ŒB��h�<��(�(D��Y�C
�Y�<Y%�c,~����Y��UK��FW�<T�3�tP�	�C[e���N�<�'I�3(�Y�D�4-�4c2a�L�<�牘�Q�8ش��&~�T�rj@t�<)'���l]XIߥkm,q3EIY�<!�D�q]�9[pc�}$Dcr�XX�<9`��6WdU(u͙	:I��Ru�VW�<�B�s�D���TYjF�R�<!��4][C�U ��"f|4m��|kr�(�D>���7O M�̆ȓ8��|h�F�7��Y��WL��W�|��6�J\)8AKԁ::hB�	�da�Ցe��/M-��)*B�)� �LA��I1-��{A��C�j�p�"O,�ʕC�+V1B�P�U��Y"Oh`CBM�erĝ���y�%��"O9� ��,;Q���AR+�j �"OS�S1-}�ո���d��Tx4"O��P�B���ݪ��A��^Ez%"O��xT��&@0��@�;�@@�P"Oִ�ĕM&,��),Ik`�c�"Or�	��{��y���U�Zt\	4"O���#�� �$	�M[M�	��"O����*wCRI	��̒I`HiZt"O&$�����:}Be��kR�O`4D:�"O�X�s�Ŭlc��yD��"O.��fHS}i�0�j�2*�I�V"OzH#��W> 5��
�u��2�"O�iX�"T�	.}j�Iװ.|���"O
̃��\7 ��2rb�9bu"@�"O���!t�6��pB֢u�PR"O��Y,<hZ�H#�9?{d�Q"O�jN�=G;����"E}=~Xѷ"O���EI��A)䨃�b�f8xi�"Oڴ!s*�9Lm}��� 1�ٓr"OBT3�l@4NY�dbF�����""O�!�B5
��@�E�#��)�"OP��5'W�3���u�B33���"O&�8s恆!y���h� �"O.Ak�.�����Omx%`�"OA;#hG�\<��PS�U*�"%"O.�b�1J��d0�!]K��H"O�@#DD�G��q���4���	c"OD4As�;$-D�iG�)�r%�"O�+4�A�"��P"Y+G��x��"OjY��AC�\�F����ɠTJ���"OH-��.�L�|\�A�E�L0nXu"O��p��7_԰�%�Y�4��"O��j��O5Q���ǎ�5{&�Uʤ"O@��C��8}�زD� J���"O� �k�3A��=ѥ��6�*�)r"OT��/�L��M���p�s3"O����ō�$�jm[�
�ނ��"O���)Ͷ���Ql y�<4�V"O��3c��<�@��%��X�`i"�"Oha0,֬bB��C͍X���3"O�H
��^#�4)Àc� dK(��"O*�s`�C��K��0{��`[Q"O|`ZQ,n�yWᔡ�P�k'"O� ��G=E��eSp�ۑR�>�"O� �bg��k�4���H�<N�y��"O2�"s��~�#��9@�"Oz�D���=:��X�GǴnJ:hu"O&��!�Br�.u�/�"
C�;4!�J��f�x��L*ބ�R���|!��P�~RHu�0�xۦ������
�'�^���3G�$�AɄ>duB�'�� `��0�p|J� ?���k
�'���j�(�H�zwi��f��	�'���;5�F�t�hr�8Zֆ��	�'u:|X��6*񨅙ql�{Ś8�	�'�-�RC'�R�j�'е#��	�'���a�	V"/m����)�fi	�'��+���.uO�k��: �\p��'��ɢYLm��n]%C�m��'�(m�#��
�(A[A΍�*cЅI�'BP�J�|�I��ǌqF������ 6d��,�$��p��G�ip
�0s"O��ycB�y6X�l	�sZ�$"O�%C�
[�O�v�9�MM1I�@p�"OZErr�Z�%�Ɂu�%q9�Q�"O����${	X%�'��4��5"O^u;fi�
�PêƷR�A�"O���b$V70��d��	F�*.FA��"O��6%S��	��Ĥ/F��c"O<³�ll 1rf%�Ġ�"Ol�4�ߒ
oj
�G]|j	�"OlřSD��6��	p��� "O��Z�L��MJ�aI��!S"O"\w��l� � G>)z�y�"OM	bC	&U��S��۽	���1R"O�8�"/W|���|�ڱ�@"O��Y�+�F���1�9b�r(8"O�E�(A�J�,�����7W��#"O�  ����*
6���D	4���%"O��4�S�l^I����7/�B�0�"O���1�V4P �p��V1f����"O���7М	�|� �Ϣ-�0�'"O:`�De�}�,��L�'��y�"O2`g�H) �P,z���=¨��V"O�iJ�OH eJ��3�C�q�V<�5"O�}�U�L��l��*��,��)�"O��QU�(�д�&@(W3hD2"Oba��:V�!S�r��"O��0�%~�T`� e���֠?!�D��<6i#1�ek@X:C�C�	�Q�0܂BƻU �d�l�0bb�B�I�
	�4pu+Ҁ^����v�#B�B�I$CBԊ�F3:�~Ȼ�
��d�:��q�!�S�d.z�Z���n-!�d�bo�U��b��2�e�W�GX!�ӣz֚���[v����S;
	!� �D���q\�;!|qyKU�!�$҅tR����W
H+8�8�m�!򤚧vs� ��*�T5���!�ȇK�XJWA�>�@W+��N�!򤆐Z��H[b�ؑC�T�@*۶6�!����ȲЄ�!�$�
D�j�!�$�	D#X�D�$��L�'�� �!��x�b����9CyQ��f�3]�!�܃c��T#1� *q��'��J�!�Ʀ#F�S!ڝEf�I���Z%^�!�d�IM"T+��H&d���3�
�4�!�$��<��C�W��8��)ݯ\�!�*{V�d�P�T�+�����H�M�!��I.j�0B޵���VE^��!�L'���ړdӇӞ� ��}�!�$ַd݊�l2R��Z���/!��4-�d�r�� ;��#!�d֕�N�1�(ġX	r��,)!�X�e3��&逼Z����Ԫ�=!�d݃#�v�#��D}��H�a$�=�!�$LNDP����X�C�(髠 N�+6!�$_�s�DC&���e��9HT���?!�D����B��N�h*!��:ʡ����A����8s�i̈́��y�nʲސ�K)-L<�8e ���yr�M��~]��l��[`еx�P�y�.R�{���i�QW6<��O�yRŖx �B䊮TX�H��'Q��y�G��@�p��� �
e���y
� �+�h�Q�nh�ւ\y�p�[�"O�1چÆ�gN���<�����"O��+N.�5b��Ğ���"O<(����g�t8��X6^���E"O�����LU�D��Q.D	"O6����Õ*�2���,YȆ"O~�;ύ�y	���Blǿ�D�"O�,1r��$`�օjU�w���"O���c�;�T�@%	��W!�U"O��� �BD�$n_-L�ji᥁ܨ�y�R Y��(�ҧ^�B����F���yR@��V��j�AN�$>�m�4+��y��]�G�~Xk�&�!%k$�Q��)�y���+����!����	h����yr��,z���b&"O�BX�uQ���y"cC�jY{�,�,��Dk��N3�yr�##�h�2��P#�4�xc��y���!�L�(�kD�) F�J��2�y�^������<(@^���4�yf x����,���B��V��yl{q���򋎡+"��;�Ö�yB�� ��@�@��)K�a��-
�yR 9#t @:Q�? I�(Y0���yB���zBf�Y� �ư8z�' ��y"��
�X��#�<��0� �y�$��ْ�װ��Ѩ�-+�y˔%r<�W�*]<@4��KS2�y���AO�|S���F�N�c��@��y"ɀL����Q�Y�.G
�
��ـ�y��pS>a��Ę�!z4��WG�$��=)�{I�&Cd"���e��0��Wk�0�y�$ѿ�$�MN�g�ɦ@[�y@��|U��#�a[��2��ǡ�yR@�cX4HA��Y�_� �(J�'y�"�S�T@]	3��s��	VfP������y�B;~=���̀�HC��s����y�	��W/�JB�69K�i[��<�yl�W��BG?3�F��p/þ�yĚ�4S�)���)�6��!,H0�HO��=	1O��(��e�X �R
�;�"O"F�9v���I��	R1"O�\cӌ�x�Hq�p�� �
5J�"Oq�F�:p�P'�s*Ļ`"O4q�Զ
����GA:U��XsO��vKZ�"6�, �W5�(��7
j�<1�.����ᅮP�%��Иa`6T�p,M�l��K�5A��$�'L��Lk!�d׌P��Pc�������X�xNv��?��S�����+�,��D��a設���+F9��
O����"b4H9�1�!C�R�7�'����d�v~�	��$%"�l]<X�t%H�!�0>1N>��m���p�/dY4��S��O̓�?!�4:7�?�z�E-b��qq�oH�\]$�U� ,OX1��b�C��RE�O,h�0.��?y���V��;t'�z��4�g�B=VÊ�<�d�g��mZ�<��O�OcA�'@�WJ��+#&�5`d`�C(O���D{�v98w�F�A�nP2�G�U���γ<Y�'�.��)=�s���b��:���8|�is5�[�^�hd���L~���-ei2`'ڼhw��1�Ղ���7�OX�!P�P 7, �!&I؃( �c��'">d��+f�HP�g��.a��ͩ�o��B䉷g_��Ȁ�E0j5���	ޫ�C�I?�%�L�bj$%C����.�4{�?O���Bi��J�'��O��䰅$A�hț��'��� t���BݸeѦHȟK7����"OBD���t3�]?�ĭ�&�'��O�`��ՙrr��+Ɠ�Z#V���O��.]�DU�JF+�Ax��L�!�֒#:��଑�?��@iVJ	c�!�$ή<�*� �	y��;�瘭Y!�ע{ x�  $͌_��"GQ�g!�$	`�L��Y�l�� �P.ED�!����~��5���g��/n�qs���OB�I�Ot�-��IS�H1lq[g�fi����'���%��_�0�b�D!��'�<ܚ�.�>Pcp���V=��'*�cFAJ�H A�B,�N<q�=N�l� "μc���I7�˥X�T���JHfMh�&T�P0����6��-�ȓ�&���D����p2���:�$��l�G���O˘0�fc<$}�t���3&/�qP	�'����T J1n$��ҋ� �
�'9������"f	>�h�Y'1�9S�O�<)E-�O��	TyB+��[�O �C��}��D �m���,M3>��)aw/�/(�!�ߞdQ̊ba � ����<�!��+N� �A�h�Zh�4M�<G!���
��ĨO+�2�a5
(e<!�$ݽ.�4d�U��+�\�;���<M!��H���=c�d?S}0���^U!�$��^m��e]�e���M�!�dA 5r�isĝ�\�T�mN�^�!�$8P�Fl(�naNV��W�(�!��B	*��%i�	\�LT����C��'v�|�"R�^���cT�'�R]�ca\��y��� ��܊�L�a�'�y�9VY��0�%w��I�����<�S�O�P� ���V&��7$��}�P�C�'�	G��Y���v]��KF�jI0�ь7lON��:7K�b�r�� �.Cr
8C�3D��h��  
��1b��R��a��/?)J�L�	c�S��AB G��ޢڦ�M�y2��'ɪ���l�M����F���y�́�#�,S�.R9@_XIg�yriK����w��&
�48 �� ��'3�z�l�z��J� ����H���yrF�S_��kSn��ȡ�a��y�
@oD��Î�/~��ئ����yb��RIL5)E�Ǥ	w6���'�'�y��H�9�ބ)��U�J�|�')=�y�nN���5r׎ѲB�t�yl�$�HO��=�O?l�I�B;>i��!�d��kn~�B�'h6$�7��5� 5�s�� dU���'�yKW�OP�p�1�Sm^eH듆�I&��i`�ʒQ���+�G�re�C䉕B�za�9ip
�Q ��
[����:�I�-Ԑ�#eF�K^��v+��	BC�	�J�|��5#B.KP�PN1ғ�Ov�'n��H)��N�e��5b@fР%�͓��?���(�i��������Y�<��V'^�̴�'��L�¬1�UV�<9pʢ^��P�AXZ��M�V����xR,��ĒЮ߀1~XD���Խ�y��S�r�OZ3*�xhbȜ��y��	l �҂��5a�ы�@�!�HO�� ��4|�႐�b�*-�6L��]��LA�"O8�[��N�8+F�!&�ݵ#�D�7"O��� �ͩd��g �!;��jt"O� vP�щ�hP{ ��BU�����4�S��\���Da��9A�����
	��B��<`l�`�	�~�������Jb�Ț'��O?���s� �(P$*a\l	 e[,X�O��'��O��;��y�JL�Cl���
:�C�@��<�5mƨ�*�"����֓O"=��O����@z�/M�g���IG�8����$���A�*��R��%+��x����A��lE��k�Kx�q�ьW�Xبu����y2��"��h�E�!L �5J0/����>�1?%?�	i�LŜl���(+۞��<AN�hE�4�9t}ru��h�*>I:�H�K��������~��'����ۺ{v	�2X;;8��	���'j�0�R�߹)D!B.N2\����'*Dp	����uC�zª�'08t���4��"<��O��V�]�VH��K��Ķ/�b%�Gܳ�y2m��\B�<��ʅ
W>�)Ô�ő�y2�E9&���AȷD�4��u�$�p<������RQ�fއq��hr	�#!*�	���|��Oo2<�pJJN,�5����HO�ҡ�4dTc��kR�R�n��Y��"O$��U`8-��8��2@�4��C^�$�S�qOp#<����X!����#ߛx��;���t<A�GԚe{^`tO@.6*��ݳb (�ȓ> �̊��>J�@�Fׯ"�x�ȓd��m2Wj��Ȃ4�ݩ�4���6��ѓP�=W��ab2(2|�ȓ�P�jO
<�r��O�����ȓ[�f�鴁R�K��%�����u𸍅ȓS%�,0�G�Dn��7�� G��e��~�p��G��(p8X�g�Ru�@�ȓo��K�!D�́�h"�ꉄ�Rx��WTm���w���"]��ȓi�VXi��I�c�B�kMTƮ܅ȓ	��D���\�h�c׍Z� ��?��<q�Ûu��XD ��.�6u�ȓ
T�Ɓ�F�F�J4�~��K�_�<YRiŮd �ҳ! )O*J�;�K^�<!1�]���	����Mю��rE�\�<��E)G�8�"Pt�HuC�(�O�<aիR0�X9���4}�=�B f�<!Æ��Rޤ�!�a`�d	��b�<A'�0J��C'}�����.\�<Yap�c?n)�ɂwJE�dLj�J�'eH�V/��2k���W�vk&ȹp
�'1Z�+�F+6и����#YR\B
�'��@Q��33֐��b��Bn>5��'&I�0MBn>Бv�]%9#�`h�'�f����!u�T����.�2���'L<a2Qd&P�d+�?(�����'B@=��E	.L?�@%+ب���y�'{��h�+�-��	
�Ʈy\���'&\����]I|��W�Ƹ4��'��@آ�Go�"�J7EȂX�\$y�'��q#a��k�N�BgLGT� ��'8�(��h%n +���,I�0:�'.fLX���x PXcG�6BJ�i
�'g�H� -B4_�`$#C&�-X
Z��	�'�^MhvK�A�j9�ш��JD6��'�j��M��C�BX��	jʔ��'�z����]]8������'ov�w
K/�6*Î��XhA�'4����hP�=I�e����'�)�  #W��� !�y;����w���%��	7��d 
�&�!�� Du� �� \�Q�5�¢V�����"O��#/W2x�rM�!�Z#!���� "Of��3ǁUkfĘu��<�"Ol�0��)7R�j��#c�� "O���4!�pN���ӄ܈y`Z��"OL��Q,WGpX����\��2�"Oօ�e��=o��@�H$8J 8�"O��0pC�V�vuȦnV)�����"O&�FM��'�ɧg�$<$Zi�"O +��Z�4u�;(��"�"O
�ا��	"�U�#�J<R"=�e"O����NؿC�|�v$�X`�u"Oj���\�Lh}�p��1@��r�"O���0<J�X$a�p�rɒ�"O��{�$�'q�e�R��**�x`�"O��('��#�� $o�Z��q�t"O04��5W2ZDu%�,��f"O4��PƊ.dV6չ��1��ʒ"O`�YdD�VG�h�.�\���"O�	�tkL�B����G�"�>q�V�'C����gG`�ɺ(�lM	���}�ls��^%tC�		l2�hfj�f��LA&%�5P�F�'̈́%��,��j�p��ᓜQ~6��V��l^L@2L� hC�I�o��X"�� �PB�K�1)�DA��I�<Y�΀%���"���Y��v��[ǫOu|��F�$<�>��RIyx���r)�9D�x�� ��{�2B㌡EFĩ�w �5�l���Q)"5�Q�*�%~�Fx���?[�"����*���0�ө�HOL}۠o߬o��Y��j���^��Y?u�U.�14�A�w�W�H\�ܒө^�z�1c\5z~��	7R ��,R��4��K�q�ye� k7�����\�@[��6S�ɞ�S��,����7s��y[c��eH��V}�L�r��P����'�V��Qg̃u�|����.}�����Np�4xG*��,Aբ�m�l�X��ag�<�"�X̻�N���$��C�b5�v)�:�*#5o�w�|x	ب}��]�d��Y��uP�k_~��� ԬJ�_�r�eN�4��q�g�'̮�ѥ/�#_��Y ���qO���ǝ+�zT����D�։i�ቺ0h<��ώ�R,��ƢƂ^�`��F�\��,�!�3�jX����	6�C�b��Z� i��WA�����'<@d��L��p�t�c�ς{�x �c*�Ec��>�6�ǌ�9Fl��,P6q�z��<��"��{�,�������#\&�yB�#a~r4�y ��3�I�5nj"�'�"0�2Hا�I:3��UÇ���MST��,	��R:m�7��E� a��o�1O�*��Gd3�!A�-PFX�\��o�(m�A+2�Z)y<��f��&��1C��-총
�'C�}cRr�O�0d(�B+s((���L�&��a&?�FL�>^P��ˤ�כ7�r)ӑ��I�';�L
1�x�� �IL�3g,�r��	$ӘI�7/�M56�P#$X�ņQ�|��R�4J�)r�Yh��_�,IT'�Un��O��Q����#\�k��]�(�#U	�zrae��"�R���)�S��M��G!U�;rL[�<�c%��)�0�  ?,�Z�!B"/X�䢍�R	������&`�P�qO�(3�[a�h������B2�Y����Y�uH�	�-�;䣑0��c 囇b�`ز`���F5�q�h�3 ]������FxI�֯_
v�kD�[.:|E[��t�'(0�Eo�l��4А�ׯv̭2��ǬPdJH��@E�,q܁"�G��Tz}� �Ͳ[x�R`(Erx���@�$�/���zBl�A5,�ڲ���~%Dz�kAZ[l)	f��Ji�B�LI����W�/|!�w'XVG0��1A"�H�b��z{��Ud@0*��,s�"
5+j���Y�SM,�BK�C&�D�R��w��I��ŗi3��z7��	�� s'o��V`�VCX-v��7�ߓb����cX*�t4�5�_��1���;[3��I�a��5����k�֥��c[�p�p1f���)�i���X5��#G�)�9����&�ߞ(R��*�N
q�DlZQ�ѳ�ŋ�X������xX�1��;_���@�ߺ���QhV��GI�K���-��Ԣ�O�-y�N@I1��+�Q�d�Q��,.� ��'�E\�u�$�fe"����R��]���_MtjA
�f�r��1�4+�"��Pi�I��PJſipZ���ׅz�h�2�\(Ť�7I�/;�-���D�;'���@��ɻU�Q�'��]z�p8�"(^=v�V��Mí\�,�1��O����kճ.�6��%� h}��ȟ�u�F%���,X�8�Q"F�K���[��ɣv	�=�&4!I������M��(R`m��mCDˊMl��9O���9mE�hI�	M�[�bN̎$������4
.��H@6p��� Ҭߍ4V`�p!�+=�D[���!����PC�6�u�*���������
�ܔl�"�q��:k�B����F����8/lD2G-܉q(4�C�(�;+�0Y��"�&t�ؕ�b�?>�$�ɶg�>F��\9gc�';:\$��C�hs��SthN�r5Nh��c:�4��u'�Ӟ �9AL���քՠ�xre�7yR����M�lJH%�Ѯɦ�M�Ə�2��!�-I*B=�)��LJ�`�`S��2<d`qpF	{4���"^ z������c��/O�K��U�2��f�S;"���Xdv����-�7̊��.^�Dtu"Ƨ�(ׄl[��Ⱦ��YrT ��cw��Ჭ	5��ԃaΟ'@f]z�*��%�D�I�:Z�I.� {&ᩒ��N|�����'劘�Ӻ��S%�KS�8H�	w�����l0� ��� ���k���-Y�� a���*��@�o�v���mL@�,�R�Z���+�g�[��9A$�Ҧ	5�<An)�G"�>Y�����{���Ɛ�~.���Uo٠�K��>Ed��"�>X��-��`�1QV��e/�P�� �a��T�Ri�F(\�2aj5����uhT�g������&��dT!PIH�9��v�Ⴇ�^�1�꼪񊞟t!���V/x��PS������iw��9zѢ�!�0����1ʟs*�3@�|��:�g��Wd�Z��*�  ��+upD9%�ƫ���V��4�"��̺Ù'`8�bU��Q���$����"&�|I�@�À�5i��:
��J���
�$<X�A��#���@+ܢ%�du����˥fŁN��÷��*I�tYT���d�Q�}8����OX�
C��&��	/Z=	V�֙x�����LZѨ�IGbM��s�(Z�L��D���G�ƕfC�����^�B���{�rh�d��S�h�n�_%Tx{c�ٌs��� ��ʠ*���$E�2���(�k[q���Z.NL۴�zasNC@W����,�~5Y5(�\J�z0�kQJ-��/P���Ť *{H)���U/�n��2C��������s�$�5�Pw�4,+�O
�/R�Y��S"[��a�,C�B��؋�O�r�$�UJPu�><4��aln�����a��N�f4DAfƗ+>Ơy	˓�`�2�KQMp��ֱ|�n����^%O�T��u�h�'Ȇ�yt�a��4a��(���Q-�y¯>O�22�wM�3�E�?��tH�-H9	�h��!�,�C"!Vh�`J�I {�L�aAo���Nؙb옦&���lԚ����@j��/}rr`ɡy�B�Y1o޽
�Z��L��0���,�Ҽ"�iA�M���Z D;�@�!��
(�b7i@)N����d��	`�40���0��遬#��y�� �Rt���O�"�+%�Dx�%�t\L`��N�zBz�#DX�,	nڋ���)��q��I�k�'D#���p�Xp���x�VBa��_Y�axDCÿT~K2��"E�X�e؆F66��Q"{4�y�G�V/���d�C"���Y~]~�ɢk\�M�4�@�R>Y����-�����~��>q��#$�ʼIV����۰>Y�"��Բ��.
&�|ڰO�$;@iY�y���ڰbI%�nT�!.2����j����O(�qt�A�T�:| �NC�	l�0q!8OPZ�샇��E�Hdu��԰V��0�C�0AD �F�:X��{��tӠ-��L�.�I���6͜�o�!PӓlD��	ӄ�?22�jrA��<���m�4d�t�g��%YE2�2'T1Ԓ,	���'|trtҥ�B�(zR%a��Ȑ4 �Pi+��B'T�':i
�!2|O@bR �'"(��fRy[)��DA�k\�!qA U	a6��w�P�A��楞�@����{^9���oV�)�@T�k$�ؑj�\��c��	��5[�&��K�>"<�S��!���c�ƙJ��� =�2]p�)E
`�x�#�Z�����=�R� �	0,���i�),������U�A t�0P��_����MO|~�*F��,��	&H�z�����`�>�R���0+� }�$�W�<��E��&�N��B���D�^%E�>i�v1r2�H$n9};���3S6�f"$t�d�c�0�|4��I�_ku��U�+����ԣ�v�ɜ@�.d1h��)0���6�6�1�J�a�x\iA�сD����ĜP'�QxWFG���y[�@�N�)U�=,O"Q��hV�##N��ê1#�ȉT�]  y �"i՗J@*�S��J����#�\m�Ē7*�����""�2�4-��@�s��CF$��V)Lg���
R�{�,��?�Do_$<��|B��Ӛ�x2�O�(�!T$�9Cކ}��JԐE!�@���kF�9��~�T5)�"]�F�q��B݀q��*D"�H��_?�I�Z�&�:rn�88����G�"zx������cӨ��x���A�Ȟ�(�h��p�H�0����'��4��呚w�xMr@&H2�$Ģ�˔.��� ��'f�`SC�|��|���ˌ#�џ����4)�b��BI	�D�}o�Aj�.,s�.UbH`�Iы�$�ɱ�\uq6�zg �(�)	!o�1q��£u�@(0�E�a����F�
������*	�V�+�X�7��d� ��Q"k������W)@��&�)��܍/�h�QB�',	F=0�-ШG�.���\i�"��=�anI�M��A�� #k�H)�6���P�T��u'L0X�4�a� �}��h`�㗹m�@��Od��M�w>��9O05���T��Թ�	ؔJ��Z��2i�m�N��]�TM�+`6 )���ZTⓂS�|�]�n���j��� ~��dRK��P�ɣw�
�C�'�\��؈��I>Bi�l������ �dl��?�:�{�O7,�:`c�`�E�X�R��å��b��K��P.P�%�����M6W�޸����:��lc'KYџ�c��NhV�TJ�Mݭcydh�pF�y��H$I��U�F4R�/L/p ˷���A�4�reM�O���P�G1~�� �i�<�O 6�`V@
|60�ؔEm�v�`N<I��˹+�2Ÿa,�$�Dѱo�����rmS��J`j�̎ ������D�A�V��s�ˆh��(�	n�H((k���?�$$�Em�8R��]E*�,,��l�cɃ�Zݖ�UI�S� 芲�ͧ9�48�u-�|� ���0���MV�B"��?��u�`Z�$��	�5�` ,O|8!��_3W�q��KX,s ��[Ri� e"�)sE��5o���7"�>'�$��ޱR�E�6K9�	Ɔ���gV2T$ �z%���dY�ɼLZ�H	~�ZL��� ��;D�r���؅,U]� @�P�F��p��_�P��DZ�62DY�cE�A
vg(ƓxRK@��|p�,F�	ej����ʩY���|H�l�5od@�!&	*��pզ͗oA�[��0D�X��n\�\}ss��0G��Y�7i	�	��}AE��6��Kt��y��h�P�$^��?o�m�wL��UD��,0�$M�5TXx�	�'=*Y��	c��z���;� ��Œ1�$�0&��+B�4A� IMfN q���f��:���:��icHܘ;%�	p7Ă�u�yB(ܙ8"�)0��C�v|ȩ#��6e$��Q#�|�P uN^�0u�"��>�5� ΅�p=a��];;����Aظ}A8�f�|�|B0�3�=5�ֹ��ю�����d���C��];.TTT1�NQ���=�FW�F�T8��S�? ����i��8hC�H.�ա'����`㡬� 6&��*�\�|ߢ�ѐ	�w�4��8��
�V��ɉ�V�`���@ғO�p�ɞ���O*B1�W��
+���~hy���Q"�|A
Q耱1�6M�n��0j��X�K&	�ـV���ѣ�tQ*aH�9Z�^]p�.Ȝ�c�S$�p�����u�>Ip`�ͫ;�0�Qb�W8X7�ܨ0���y�n�Q�L�$%�xT�"Î���\��MF�W�\@B�'3���O6��b.O�)��<!�u��	C�lE�tE`B�ɿ�$��`�.ɔ8귯��F�@�H�,	��Кq���4��OQa ��h��t��<Q��Ó:�&4U��B�x!c�-M��~��I�H�d�@SkA�y029  ��s\L��l�
7�̠�#ҁ�ʈ��G�L�t�x3끍�u���11�d�)�wd�DH@*G0t����Dhլ,[��v機�����'F�vE�r'�q��{b�	>���6�I)�8,��)	:"�ܘ�chg��2@iB"H���s��_6����F�+�68��	�8&� ���Yi��y�#����= �Id��<RRO]3:�]Fy��$�h%Ha��(b�oܔ6��m�E���U�m�D��f� !��XX���aەE�HZVJ�`��e�e��T�}i̤e� $�'1��fJ�42�~����-7O�u�'fB��
]c����F]0^�X����8�:��UF�8hi�1���8Jf�S/Z�3�||��Ğ�`X��Ä�?`���RS�ƥlI�Q F�i��~2.�a8�[G$V#�t�b���\�ĸS�A�;vLv�a�	�/�����:g,�cD�#	�`��>�y�AyO��âg��G�T�b��( �X����/r։[�䋆(Z��:�g�'�@��@��b�rѲ Y����c��l�3������U7 �akǾ%�=� !̐[����#@\1�`V��T82G��2X�����!�f}Fz��h-�ccix�! ��B+Gh�B��:���U������1��A�.�
Y�s!�:X��*�wGh�b/�9��ÕM����9�OKG~�!�Bk��#&����
B��V�`CT��o�0h���;AX|�P�~�,p���HE��	�5"����lF��*�!&���-I#0Hj)��ې5�q0�i����fߣy�Be
�(�<z����ϙl��1�g��'���c G������!z�Ji�O~���aoމ�oB^�,AJ@+ţ�*L��˹ � ���'�H��C6u��]�'t�[�Lȡ+�N�����@KǃG>6ʎ�"j�-?,p@����w9p�C�,!*�J̮��`�L����W�Z��QZ�^ʈ�UipQ��.=�Xg,���`xӎ�@զW�0�J&Mé?,�	�tJkn�9ꡬ�/e�2�ғ߁O��u���ߡ�"��-�*9.��*����I�D����� Q+��D�:џ��Fk�E�z0P����H�c,KZj���J��`�,�d܎M�X9��EF���1@� 	<D���T�C����?ef�;�(�
U4��hP�҆&���l�����O�E��ጌ�H��8(�]�	\�tC�v������j����VaK�D�~�Z�n����QE2��"Z䌫vi�&=܈�V�ܽ��=���H0i3��cP٣�:��Dd�>s�2\�㍜7i��ܻ��C��x�F�4 cF�Q�P/1R"�å���O���͋k̜r1�Ha�siZ��`�����j1 r�&D���j"Xi���%� �J,�x���@�p�R-��ؼ[�
ҧ�����"2 EP�É1,O^�Z-W��ybGϕj$�J�ċ9$|��������].����Ar�h�V��`�^(Qr�^�R�J��ȓ�Ѐ�0�݉N��ȘƦ�52	\���aUrPJ��d[f!rP��0|
���F�X<�U�
;��|�S/�/7s�Єȓ���sw��U�.��%�Y�d�X��W2	�F��`,����:v Ņȓ����4�D#[������0`�:5��C
N`�1��W�4۰��3~�0��I��!�CN,ˮ���@�3X:�ȓ&R�P" �J74����^����ȓj�&x���C�Q��\��H�8.�|��	��$��
$� �hæD;�8��%�<l�p�N���
U�L���� �^P�%�ͱ1h�
%AA3��,�ȓ|_��s�ҙ+I6�B���7X���)F>MB�зnX��z'���.��B�ɿy��g�,,l�)RjĦp�C�	�*��)��˜3H������C�	%VH���ɈOH��E�	��C�3�D{&�)w��pv�E�BC�	.�Q��G�~�a9�F�B�Im �gN�.D����G�x�C�	G��2ꀷ �����e�	u2B�	��lu{4+á#�\$H�@# �C�	g$��T�=U�(<�P��B��5g�X�1��Z�?B�cq/�� �LB�:GE�\q�c�0�k�L�&�.B�)� ��$h2P]$���LD]6<��"On��6���*���<2Z�h�"O����!D�,���&@�6#@�"O�i� D�L
�n����"O�}��(
+4��ݱVmÖ�l�"OnI�WHAB=ZԣF�@(C���$"O���vc�o�vH�GN�`�n� @"O~m��E��
W:�᜾ �b HC"OpH�gJ�$B ��4B �FAPy�"O�"�M�:�LXqZ8JM�Y�"O>��Q�A�Jt��"�~@��)�"O$�S0+�j�z�z�Ϥ8-'"O� ���
`�E�e�x�D�@�"O^�"��5�|mJ�r��ؐ�.D���0���u`�+� D9z�����,D���f�5�*$�@Q��D�Sm$D�@E�����́�R�n��!�(�[1��	G���
��]�!�$�*�؅��
l���D�Ѹ�!��Û2Bi
p�U13��]c��CGx!���]��"R"�$�(�>_�!�݊pH�T0D>T��%юSw!�$רk��ׯ�*p���Z�T�R!���Q�"�ЫA�<�D��L�N^�y��=�F�'� �G(�=خ� ��S�� 
�'G,��VJ��!(t�HB莓N��+O�����&�MF�OJ��c���dr,-S��Z!C��0i�'���l�-/��1�9?�=�VɎ`��čb+D�ۣ��k���g}�g�!e��N0Zf�v��$h\��� �-Z��}�`�[�2�5ޠ-�d1JIpm(��ȇP��ʐb�P��Е'wD}�GH�
0\D�FxB�>��j�i��//����֞�HO���$�AWwJ)�4�ڕ~h}x"[?śT���CǲI�P�E��H��)8�!=wt(��ɘ2⭑�Z�e�Ļ"�Лc�,�!�GޛKڮ�!&�.��yFnҙ3~�)� a�܃RmPa�*�![c� QGH���|��N��;'Fщ�'\�W��xӄ��V&�%��	���ԓz�ġW��inZ9+��JR�g� �<��&2!��9�w�F4��CJ�`�ƨ�G`��&l�a��,!���!^)�q�Lwl{Sm� T����"�NF�8`� A67���dܰ}.<��Ĥ�rpSc-/�ɼ'�s&Oq;�=�rԌ 5�"<�! Ɯ}ZyV8�h����)nБ7�&u��r��8?�drV)�(o¹I2�+�8�c�ͧe�`����:IovIckK&K�֐y+�:I~���f�C��P��Lq�����:HmpE{$ˋ'Ϙ'oN��ɍYt�I[f��.}�B���"O��e,A.?~J�烥[��9f\�^�����3Hx*p�U��b�����iy�XV��M�	p������Kޒh ,��T��	;�T(��M::���R�p=��'	0��h
�-N�IZ*�(��z���S�&0��E�;���H��4��t2���8K_ �'�D�b�g\)
)�ܚv��8�������<�u �WBL���t<ѣ!��Q��+�bT�g�� gNX7[�� )��f RFI@�w�m��H@�c��ʓ?؁;��6�TZ�x:Ui� ˢt�jU�g�Nd���g��S�
I�4OwX����|.}9U 
�p�~}��gA�La���7EK�ϬE�@�ҽd'�0��GU��b�캟 +��6�$&?�<B���B�IQ�t}��0#��"�(��ě3>�I�4k~�9�@1�T��>��8q1��F���싅*���A��<T-�@Q�K�Ůx�����џ��3�Ѯ-�p��!�;D��P4)� �e"��Y9^Cf�c�K� F�\LY NإF���e�V;E��	x����qr$X�ZDj�[���Lo�dZ橄�^� ��"�gC��<B'5c89�dïeJ|A���$+�XC�E ۧ���<�f�q"	����,��`�3~��X�)W �����I�{5��.ϔ>�`�Yr��� �� � zhZ�+P`�r�+N��U{�L@=5���q V�"����i-���=8�b�T�W�81�Ƃ�yoTݲ�#	yy�j�1���3�.M3�`��U�ېa:~J����N�|Q����-tT-
�_���1�`y�"\����C�����_�gN k���Y�4*��ѼI�ם������!�8l�:��HU�H��I2�,٢q�z��f/9T�^Y����$a͜R��V9o��}�F)K��l8!M �}�ȉٓ�&l���qq	��<�g��=��u�&�����Lhq �[��6M�,�
��K�p4xU��\v0h���1;`^%���� �|��ԍ9�M�U�+D��ĚbiH#f�(-��	�m�<hsծ6=��4
�3����6�C�T�Ld�󉉡e�,)�	i�(De�E49��Z����\d�8��R��ͺ�l��(�<�ŦK0|p�j�-Jɛ5O�l	�`@�L�U	�� Y �9D듟|(ZȪeC%Z�&���j�,.X6��Gb��]�&x򕩒N���"ER�y!N���L'^�,��TJ^.�~"��x-&�+�F�
l����ȕ*��Br�̈G��U�j�B%�/�Jp�ר��{&�h%i�-Q�e�bO�rE����3���P�.[C|<x��Q�,r(���O p���eD�vM�i�u�ӆ�%7�;
� ����O�j���
A*I�h��P������G�;��nڂ*�1��CϷ���7G��T� xB[�3����D�'j�\h��o�c���g�Nhl���Fy��`p~�qi۶��a4�����f���Úm,	���^:�x;��]�.3�}�q�L�Y���x��@�Μ�Ԧ�@�Ɂ�����Z!��A�1-�'���k�(EC��(�nW����Z���b��$�p�t���<(WD�/_����ܻ^�Zl����Ol�$�7 X�]apa
¯x	ڤɄ��| ��{��х�>ĊG`Kd� �����TyXQ��|̐�T�iJ���	Y������҂92�L��'ʤ(�֧EC�ԩ��ʕ&�]�lˀ�ۖF���1��'�i"���$����� I,�AtgݏB�z�!��[��qo��D{��`Di��#�剽D�1'c���b�R�+�&�ё�W �0�(��		/�"��R-C�n!A`�ËF'���"J	*�,��1���&�hTBȊ)�<���
)<��	�Vs�����lE��"Ì`��	#ۂ 3����u�I�W��8�&��i���p�B_�� H�k	�n�*��6h�7)���AJQ����LS�j���s".��N�^�@���LJªd�#g�f�O)��8��
f��~���N�1t�U�C!V�.L�U���KnղwԜ�� ��^YH���4�/|�R�-rXI¯M- �FIZ@�V=b����VG@��M+t���Bk(t��FU�j$�at,�Z��ͪS�L����6�����̇K^и"E��;M��IqHN�XD�	+/Jpm��`�*:\���r��f�0����H��s�ț.^J�I�+#ғ}Rh �s-��e��p�5�ؕ�n��%�9���;��K%[e�QQA�|Q`4��\�f��l�EF���d��W�G ]�$�p�a�!$ݱ�#�eM�퀕3�m`�'�U�!iG0w��$A�eN�*�qa���xc�I5_�����i/�)����a���2^�2�yxӢ˼��p3�#5����'d��wK�!cΨ��Z(O��� �K���Ӷ��H)M���&`��L������2����d�� k��t��<e�!#��Kn�A�ƆXZj�n�U`��Fy�ȭIk�]�F�YRz,�en�Qh���TF�&��5�a�����&�Ǔ~N ��gȀ:vJfi`�'�~0ɷ���x��s��	�+�0$k`�� �*�ye!���6-��f�t���ڧ>�8̰��!]�I`�
�I�Ê�?%�"n��^<�R ��O��� fM�F9*��K'T���$E�02�e"���uI�E�B��qF�[����Gs�<c�4*8~y��W>�	,\�nڸ��խ�� ��nN}1�q�v`ںW^�p�D�-�O��ɶ�K�aS��Y�$ܷ'(�k�m�L7�!G��RA�Ic��:p� ���CoQ�bk(!�Q���V�Q!(;�L��A,7ڐ���u���CN�Nq�IV�5(���>�"�C�0kd�)�.ZBT�������t��$(S�=rTg��HM(l�5]����'R|!Q�,+`Dh�-��x�4%�����C����=�S�*���(K�\>@쨰��<)n)�2(J�%��Q��BKru��N�4j�4�T�_U��L�6΃!J��A��䒏���nx ��G��|֖��]���BQ2db����yل��E��*���F3^sഩ�-H(^v*���v�2��ݧ[X����%L�"�Ex�)��5�yB��[�M�����J�Y8C�ФR���j&��	n� �C3j0L�6ԑ3.^-b�F��ƫS�2����C�8���:�ʄk�4�C�б��$AkLN��dDU�S[��FL�VX����MND���A�y�AAhK^�ɫ)r�H�&L) LKBM2��})Ug��5 �}2ae����0#)�Ps�I�`ۥP��AÓ#�r1�nC;I儌���		a�X�v�qZ��M':CH S�x�`�!]&wJ�h���6Z:4����� �E�@��@�����MĢ �J@X��>)ltj`$�.����F���c� �*p�B@���]�\h@�It�>6�"W��[��!�u�՜C���C�����M�@�Q:@�ڔr���!g��k�g�*�D}�`H�w��u�FȌ(E�@Z�j2��t�FnXzt���e���v(�*��7G�h���%HG��0���?aD�H�~��iꤤYw)�s����fǪ=�9`���<z��B}mf��� 3��xQ���&�*��F��<�=p��Έ�4j��bޝ�#;]T��8P�K�d��=:KW韸��ىY�� ��! �r�F-�0�J���� �tʆ�`Ҕ��HT==e&\��@˥hO����1�@�ۛ'�H�v�g܈�J3��#���A&�A0g�l�ye�Q#�p$!r�'ϴ�Js�!C�� �$Y�n(q�𯍎3U����h����Q��� s�O�1���X?j'I�0�0T1��S���F$��j�?ތz��� lN)9����U�u"�� ��Ԓ{���=�̥(��R2�Q
G�A�iP�ȳm��v��	q�c�$r���)��<9&W� :��,&߮�;�&agzSQ�gp��B�-�9'UXzV�W1�OF�8�w�Vl(��֪*� Ҕmċ\��{�'�PE�u鑤h+N�j�@][�'䪥(��D���4i�.Ǥ4����U�`I��L���2�
�;E��U,�G����4[��]!�Z�d%s�n�����Bf��q�m��%D`Y:���CI����X5>��%��2�����ӏS���b$׾PO@t��(zg*�p�Q:/G�D��3���'&�V��~Zq��ւ�+�E�2~�|�g��F��"`�h�r��"ݛ��ڰw`��a�f)��Q����<{B����b7@ �����2r�b��,/R}d`�+H}ӧ���DSh�!߸:�c�N�e���ަ4�P�YrM ;E"p��(;�uBӈ�� ���o�����wo\�{`�D%%��U;smU�\Zf\xL���V�Z*b�ay��WK��a*�I��CU("�h*�<�Vq�t�ٿ5V��NH$TC��c��UL�qO>��WHL�B+j���� L1#��'�P�*m��82�F�&T�	��NϽ_�����K�4g܁�1"ɱ)����]�а'���f�z�m�K0�5�խ��[�\�A.����<������2�%���'��	�Ӌ�(|,ޭs�C0�����-Z�Ip�t0Z%� �"O���!�P� � t��v� ��I9AK�*�@T�(w�A�Q
���Qc����](X̻V6�Y�ۍ �������j:|��Mr#�J�Q#�5;d���|cƥ�3�@`�"�1qE���a�6bVj��T)��{
� p�cs�5���@��=�Z��6�'���0��9�J��vd��6�����.�b�<�j�@$*ŤHP�
�*�A��/
H�
דO! ��L7$�Z@h�Lج?��X&�Dx�̘�<��D�D�B�
��|cLr����*ͤM#"����;*��ɠ�*����Bw��T�<��hR�5+�H`f�]�����AG�i�,!r�b�f�Б)�/np��R"4)�ӽ\02���w�v��C�N-p���g��=J`h)qJ>�w�E=Kaj�?����8r�q��!3l�r�dZ .���3G�f��:۴[l�@�et�)�l_Ae�4�/����s��7K�$�"��7
��XQ���b)�p��.)�(�d��aa�!
���7H�tIv^U�|]z���t�n��0�f���xh�$5�J�i׫̟dqX?�aw¬<ͧ(OЅ�J���S�BV*z���'(|�ֈĮQ$��gE	;��Yq�bWa�^�b���{WҪ��X{>$���ªV������p�|���C�m�"�Ru�X Nz�)�X7��T �%$�ꤲ� 
�:5�;���:LlLb�KN(O �Ġ�#Q�E?����$&���)9��h4�qޙ*A��,Ȧ]�焹^�Ĩ�%�L��~�R�; �Պ�F�.jc�3�	)�F��S.\)t�U�����5��;Gʞ9��ũRG%U����vݰ���/�u��@P4>��C�J>��%�	T�rPz����>�~��S� �Ju;��7rTt��d�68�j��M��\��0Ç�/�@��tH�/]�VĂ`挈9n�2*�K��К5�E�dƜ��")�D��4�O,X�ZКp֟���3�R�1�2]��G�X������l��)�<�
l��ΐsH|��f%M���;�K@7P�� ��ďD��� �MX���Ŭ�R&��H$�LZ����(MU��m9EE�>�I-Z}�H�)�!p����P(3����u�@�G�<R���\؁Bs�[�\r�$ɀ�q��� ��7���B=���Z�.	R�l��D�\8��Y��U 񪓣3���� �Q�L0���Jo��cD*ܫ/��:���\=P�E��b��"7

k�37c Q:�y��P�t��d�0w:R9P��at�)�@��Qx�lx�	i�j�3򇙰}�@Dz2e�)?C&�r�E�M���S< ���*kĺ';�s�e��`�Da���V�+C	3RQ�L
�a#���
��Ļ$:�,%%	$b���$P���y�	*x3f�c�ҋW��'�b����$�0d�4�Z�8G,��OǮzI�t2Q��M����E J?ho�Њ�E*8���"&��_���&�M.T���h��#au�e *��`?9G�ɜv�s�l��*�*�*@�q��aAA>˦��R�C) 4�Px��Ȟq�k�<�(�2 C�ļ�ȕ�D�c�%��BֶQ��TJ�Z%R�@�: T|�J���'hyZ��;ֈO!�'�H�fU��N�"V�Z�Hy�+�O�(�pAp'�(pV���GѼPE�8���Wź[��k4�	�oՓB"6�Z��	e���$͐!1� �c��C�7Z�"?�F�L'h�7-�G.2��W
��ES�Ѡ�B�8�Q��c:�J�@��.>	9�#\�~9օ��*EAX��ȑ"�>�Y�/��R	g���eę�P<1q2�I7I'�y���f�Fm���	4B��t��k���!�:m��9#��H�(�!HȚ&c����P�2cȩF��O�t0c1�Hp�RaM�k �>�i��/Ø�dT��f�i���S#Jj�h��ʊ;�X���D#D�87�-k8t񇖁(Z��H��Rg�'"��H��S�x�����$��|��R�XJ���WmQ�F$��P!&ĄS��ҖlU�����Ő;aFDp	�'Wf�h�l�t����DJqb���d��|��ؐ���5*�b��~ʰR�=�����͌�p��h�g^�<Y�i'�t�Sk:�n�05+��5���)@B��8���O?�$	@�dӄ+ԒwWT�
fCco!��/�Y2P�@yH��
�ħCV�	1�)y�'��qr!FU�P8��I�R�X�
�'\���&]^��q�;dذ|��';X��vH�;�� �_!W��0P	�'ͺLxdG��u��0�U&��	P�'��%qp�Cy���(�.ì$��'��X�A��N��I�)^Gx��'��]�V�F��&t���ZW�P�8�'u���		2N&긠".ӞN(����'|f��%u%�Ń��4<B�p�'������\&o��Xmg�)f8t��'bh���h���>@����da�<Q7 �I���I2�9���ʲO�W�<��� �xM����]Ÿ�
�J�P�<Q2�:�l�	�m}$(���j�<a�dS tj �"���_�x<J�*OO�<d��DH�Xb���Z���!���G�<�Gn�A#��!��2�����v�<���7	^J"B���;�No�<�B@�>?�uR�;N'���ƁQl�<�E+ڀGfp��I�7H���Wh�<�  �Q��σ�:V��!a!�S�<�ǎЖ�{d�W�y���qf�SN�<�b�C�G�TTғ�\���CG�g�<� �ɂT	��[��sA͌ [ҭZ�"O���ӬG$=�@��3O�/}OJ j"O���E�՚Fx�y���1����"O	7�ޓ? ��H��9)6��"O�-��E����:�B�81 x��"O�	K��2?����蜪mU��w"O��Bd�;Z�P�t-�`��1B�1OT�kQe�&H��y�ܠc��:��	�v�}X6.���8#R#�T"�p1qǜe� l�<%>uV���Fd���B��`�B��� ��Ax�� t��	�M�G��0k#(6�0|����c�8�
$�a�>�1�R-!4�����N� ��T���0�Q�5�F/���Z���ɋ�!VJ8O��|1��e�		���r�� C�V���=^7a����8���F��:��,��@�<-N�{ kN�o�xe�é��9v�{	ç!g���&�0! tI0��j[�Abƌ.n�k "�i���YD>)�.�"`�(�G�wz�X�u�2Q�pl(�rax`r�G˵X������s��j�%جG4 �"�B�i�Z�0�M�)vX��rT���H�ç9����QIb2��L��Z\ݑ�{�@�.��"~Γp��(;�NL�&��\g���2��x"	��`
�	8p}��r�#�'��#�#kb� �"/g�� 
N�	�AL?�bFJZ�T>�[̟���` ސT(�8"A?@��0h&�'�	�#����NfRa��O
oqS��i�>a�4����I�jҼ���S�<I���~�C��y��3U�ı}��h4�B��u�!Oµz���Fb(�G�D�Nٺ[g��>'�@��҆@+4��8�ҩ�u�n��'X�)��N|���i]64r���BxI���G��Q�Io��C�Կ,l���IĦ�ٖ�*tNL���\�ʣ�m(��J��i��Ʌ!�*�?E�DOS�\Vd�l^0M�To�6�uE���Q	���OT%�çv�aB4��<ݔ��#?��p�q�\�DBZx���'��5���Nw>�+�#-z|s1g�"3
Y�R/:b;�d���r�)� �е)�P��)�~�𝀡�Q;�|u�٤7����4�Ms�:(�Fs&�MG�O�=Ғ�_��E{�,@�v��Pi�"x��b1�4W� 0cG.MF(Q?9ڂ��i��_qYp(��m��'2.��,Oaɱ�7	+�̰�s�0�t"R&�$�y���kTr�;D�T�¥�'4�`ic!ӣ��0���4D�T(U �;ҪX���>Ā�#��4D��Z2��z�ԉR�o����{tL1D���℆z0i�!���*��tq�	;D�HC�H��
ѲxI�.�f�LxS>D�Dx��Q.��-[����C?D���p�W� ��'�Aey�����=D�P{2��k{>|�`Ք�X��=D�@{OG~d�d�2�� ���:D��Qd���^�@z��6X���p�-D���Gω8�Mc�T�Nj�Pd�7D��X���%3����nT�d���t�1D��x��� �}�@��O}�L�F�4D���G�k�0�hrJ��C�N�;��$D���'�\#�6Z0��'"D�|��!ˎz(F@֍A,t��k�!�y2�O�R��Vy�����M�8�y�m\���|bǂЏhRR��/��yb��	7gh���H[]��
�J2�y�`���P-�TX%㗆�y���5���R����xL�H�3�ׅ�y2+L�}��Q����j�p�������y���.&	�IX�
\h}N�R�,�yrF	�j��u`4C���y�`��䮴9B���C>!Y2C�:�y�C�]���Y�.G��98�e�0�y��8M���HWP�t}{�
��y"d\�s���2����]�� 1eA��y�Ȉ�*����P�T��e�  �y���z���HJ�y��Ņ�y��[X��O
	) y�E#�y�Ǖ� *��Ug�Y����B��y¢3����P��Q��H��y
� ��P��N�R<��P��Y�ltm�R"OB���A+=�e[G�T=n´�"O ثaJE		�L����@b��q�"O^��p�ٛ�H�[B��#k�7�$D����T$'Ѽ�p��Y7L���-D�����T&X�ҥV'/���!�*D�l ��*	�Ȅ����\F�!;tc)D���� ,P�a��� G�b��(D� �h��,��l�Vjԁ{�dg,D�\GNɗ)A��@�F�<�ҹh3�)D�TP�@��@��ŕ�b����3D�`�bLH�|&vx`�f�P�R�CE0D�HK�Ý�GĽ�1�ؚdB��AL.D�
���!a�
�k��sJ��B�ɭG�����@�+䰭��`ʄ|i(B�I	V0ب[0�[6��xr	�n��C䉓,�0"0�]H���H��	��C䉍B���ݮH�d���y��B��V�8Li�N�$_q�%B� D�J�B�	'H���#���h��1y�]\"�B�I�jp��R�����"�ڭ5g�B�	8q&;��^�������Q�$B�ɄJ
<�H��L��$3���C�I�\:��/�18�<�r�Ĳ!l C�I-?�ndx�(Q,-ltX��BB�,B��D�vp�#f�4Ԋ,p��C��KT�0�� 7ۆ�sR�-mg�C�	/Ft�Rg��4��jPf0@l�C��)_����!��|aI� �#2��B�I�)
��C���`��c�6�B�I#>|@�p��_c��#F �4\�B���JG�ӵbv���bP�z��x�
�'?Nl�G�نh� �J4�#���	�'O����8���SO G>*���'��s�h�yJ��sS�1;i�}"�'H>d��C��?�p�
�} ��'�	Sr��\�6���*e>��	�'�������Q��ʤ&��m��'`D`:a�M�Z�,CA�C P=J���'3b�KF�M8A(�Q���0I�fu��'�Ԅ
��4#�D
Ǝάl_:��'��$B���=o�T��+ aR�i�'jR�1AI�#�\���X�Y�'��uC�!�[d�-���@�V�Z���'�t80eBW<�@��S�M��M#�'�m	��?,���6C֥Bs�x��'u:4sңA�/t���M�>�j���'N�sAK+1�ix5$�(��$�
�'���i�J:*����E[���݁�'�٫#���d�@�b�4m0,��'��9���	�0���1A㕑vt`��'�ty6��]a��2gDߟj�A
�'~��*�Յ\�[���aw�!��&��Sc�8?%ܰ��m�PV���r��h��M师uʜ�X� a��st` À雼"�t*��/T&���Z�fd�#kB)}v��)�g �DZ�q��lRv r e�|���Q���ȓ�^����+1}���"cN6CwzŇ�&&@8��c�j�P��.g�I��|�<��n�Dp��T�����ȓ}�p�2�S�Y+bqP��$�ȓvj�E���_�Q���"��1�ȓ~d,	��T�12=�C���#p`���S�? ��	T�ե �vh��� P��r"O�l�t�/��Qbjٔ�(xU"O��s@.� 0�H�1�(��g��J"O��3"�7�]X6ϱB�F�3F"O@l�jY"5˲1#�Asy��"Otۡ.4T�s�J}���"O�����(���k�6��"O,P�Ձ8@_�� �\�f���D"O�m�� �&�� �3Q8#e���"ODh���&�hՁC 1����"O��J����[!V-�� \#��+B"O��k��L�M@�Y`.�&E�Pe"O���RmS��Г���,�c"O]���%|V�<��b�N�8�"O~0��/L)�t�pp�ŗu�d`�"O��S퉧{����f�^<-��+�"O0�B�J�x=���JV�B����"O���JhP����5v��1�"O� �5BF�2=��H��k���"O~Iڡ�s����-�3tߦ��"OF�;G���.�l��w�_";����"Oi�14z`f݁�DU�D���:�"OH�BG�T�/\��W�F���w"O,�CZ�j9 �8�˃�l,H�"O��@}���� ޴P�(�7"O�}���4Q�8v��o��U	C"O���&@�#]x rh@��8�H"O�1�D�m,�@1� ���]@V"Oj$PEB�1��p���<{�eS`"OP@���b��!pÈK8x��5;�'y� ��0�+�τJ.��'��t�R�ɼCb�(I���;<�v���'�t0R�)"ul�Z����4� �R�'�4��c���.�`�^9�j`�	�'��[!o������6!#�'�Z@R�M,5���beHˇT��R�'�T�0g%IE��Бt���V؎��	�'Ԋ�S�ƀ{lV�@t�G;N�*�'z�)��fڋl���@朚7	����'K�Tz��_�T�$)	�X>6�TH��'�����o�*T9�	j&����5��'q���Cͦ<+Α!}���b�'�ja�Tϗ�Y�bԆB v �qK�'�Τ pc
����R�w�b�9�'�:%�֮�Rs$(�a�qP晇�_��TK�E��|�@B�]|�$�ȓb�ЩhR! =e��b��5bC�8@��,�ЮO?2�$=�v��5(��C�;h�8�f��<I��,%)�>_�C��9Waxlz��R�HΕ�v��"O�=	v� �i�r���-��'�p��"O�1R����X�6�R(�"O U�e�0E��QJ���'���"O����嗎t��LᑊȖ7�8�)"O�]� ʛ��c�鉍tsN<�E"O��A��zO�S�ǃAX���f"O���p*�"q�j��B��6AF��"O��*�E��m���EO1*5:�!"Ot56m���Q�.  x�yt"O������ `V\[@,�"O@�����UR�hc��@jա�"O����e�0B�v����E�5���5"O�PH#-M�)�<��*���B,��"O����Ye��a�&��Lq:s"O� ���h��z� ��"��9wR�i["O��:�J¶������!t7hp��"O���	�<�v bd�Ȃk���"O^�˃��yt䈦d̓O���0�"O���Sk�0m�4�n�U�4�� "O��Yѡ޸@{.��g��1(�@a�"O
�����>W`����Y���0"O^��q��Yh�����8�ŀO�<��b�4ʰH�j�*O�����]P�<	D!J�2"��aMϤj�����`JI�<1F�ܮ�D��fQ#d�����}�<! �)QiV��dZ�`�@(��gP}�<٤�O���I���!���@0�_�<�&o˚X�b��rYC�ƨ `�<�#l��n��O5??hp�BY�<��L,gļ`��N1`��U���L�<Q�;6��<��ٸ�6��n[E�<�	F�x�z2ٛ:���`E�<!�Kұ���a��1;���ȜG�<qr��Y?�U�����i��\@�<qE���uPG�ǥ&�)��dTF�<� = o� 3#QI^J<�ȓ1�nyx��v�B��N�:^`��L����v ��g�Ή�3�F�,�%��W�P�3'g���J�D��>MjȆȓW%.[�l��`9<��u�M耆ȓn�A��aŞ�9���y#r�ȓK^�	��˶u�����JJ�ZE���ȓM˪��&��.�������lzn�ȓst�0{�	T�c��a�I!��%�ȓjm�Ĳ2`��k�x���Z�[j,8�ȓL��H�d�ߚ6������ۙL�nȇ�Iy�FK�1Szh�q%�2ڬ�ȓQ"i@�J�
�2�x��ʖJ����ȓ����s��..��2#�_�{Ld���/Y���	C�PЪ�m�"�4 ��8�\�� @�?+��d�dBG�"9H�z�;D��1��P�c��U�E=%<�1�9D�����E�+��X&��L:D�pX�n����a���9���q�*D�,��A�0����Ԯm���#)D�y���
6���H�w�`4��O%D��* �N���Ҥ-|�6��ҥ!D�h�1��?��H1��
�N�$�8u3D�T��̒NzƸQ_�$�T4W��C�I=[�x-5�։j"�=z���p"O�8R�ͼ
J��L7(��"Op�*�F	T��u��悖$:��"�"O�;�E�N4ά��/�O�F�G"O�!�#�V�&9vL����&m�hb�"O`��@&E=*Q҂c�b���Z&"O� \%�c��*"�%�a4>�@e+�"O�I���p����p�jL�g"O�0��._�;���礐�$.�y�"O��7˘J�m�D��J6��""O�L�h΁���7�7?|�"�"O�b&�wP����� 8�DY�"OV<Ɇ�\5`����P���r1"O��THݵj����Ј3�N��"O^-;�G�&�<��û&��!��"Oac�oG�J���&�
|�:�k�"O�mÁNY)Q �H�\ 3�2e�"OP%ipg
q���2$ڕW��=A"O�@A���8Ed	VC�f�}J�"O�AQp���#�СT%qH<S�"OrS�T��6����TZb	;�"O����֙_���y��1I����"O�|��5�6�h&	�,3�a)P"O�(r�@As��`��Q)�Y��"OJ��BdZ�7Z�L��o��>��0�"O�l�%�:t��9���ƀ`�f�#"O���ƣԍB�0��Եa�:��v"Ot,@w�O�L�$I	��
$�dL�@"O�zԫK�[f�����B�_�~��"O����i9L��0z&��,���Kq"OP}�+	�` ]`�O�&H�t��"O4)ɱ�֓*^�	����j+>�au"O�x�ՎTBT�s4�޺o8`q"O���Β�d�����#48"�z"OT#b]1L�^�����/d2@���"O�!�!� ���k��QRn�B�"Or�
�Nʖ>���o�&�Q�"O�%B�!S@��A��a)+�a �"O�� ��9��l���T�OR-��"O�%!�!��T�*幕���oZ��SS"O�Pᦩ�|"Hi�A�.�`D�W"O��q3�V����U���r�=�5"O��RN�m������'mEP�S�"O��`�W�S�A���R,�吳"O$���G0.�n� 1f�4v���"O�i�wE�>��b;<����V"O��;��ˊt��W�#~b�:w"O�2�(T�s�P s�E�5z:Ĺ6"O�� ®�L|�,WG��Փ�"O���G   ��     �  B  �  m*  �5  yA  	M  �X  ~d  7n  �w  ��  ͋  g�  ��  �  o�  ��  ��  b�  ��  '�  ��  ��  '�  k�  ��   �  B�  ��    �
 � � �" �* z1 (: B J OP �V oZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��	��M�#�?q������¦Fr��,/`,4��'�6m0�i>�	��p�v��.E����w��`Ǐ�����-��5$���';��đ>�R�ӂdY��N��Tf̓�?�*Oj�}�0�^.8�����֘{78�R7m̋H��$�'��'�Hnz�5�Т_v�x�ĉe�n����Bӟ��I�<A�O1�����<1.� ��Y���ؑ���<��'^��D��hO���O֡� Aհ_���xZ9��2uʑ�<Y-OX�O.aoZ�,2b�4A�DZָ�b�뜂&S^Bo S��Z �Iݟ����<�O�4c@o��d�lS�_�W�d\ ��	�6�>��P�>�'Tl������dTC���i��
����]
�,i!Z���'��9O��Ђ/�?X�ań�.�Xh�:O��m?Ϛ�3|�V�4�8B�` �j���H aDc��R�9O���Ol���2�6�Ot���J� Ҹ;��I�&˔n!Z�(�B��}�"�OX�S�g̓W�� S�
*��r]
,n(�'h�7͟Z(��D�O��D*�Sxê�q`l�8#�jyxG&�	 �H��ODm���MC0�x��d.Ёx
z�h˕��\�f!P�:�p�B)A�7�剄@��R�u��|BR�T�e�O�m��}K�/D�
jK	�*Da|�a�}V$�O�t���^�l}v�k���9|�Tu�p��O��lZN�u���pnZ�M�It�4���Wt�L](��H9XZ�K>��R�1��^�S�ߙxr�	g�V�"P`#	�0��Oe�����3g^���W�=F��peC�TRj(��ϟp�	�M��AM�dBg�t�O4����՛@2DmJ�+�
'
�:�!#�$�O��4���3�''���4=b�G	�Y�����k�iM�A�"�P#|��IO��Py��d�/Rʦ�:�A��pd	%�� N��,�ܴ9	X,���?�����	T l�
l(#�
$1n����l�62������d�O��� ��?p͚���-Z�͊'+vi[����YP*�ş�����D�i?QI>!g�S\:�\��FU�C"�L�1�?I���?����?�|J.O�5mZ�[��DC.0A�IGA��@$ND_܆�$�Oڍn�F�/��I�M�N9M�ea@AE�S�d�	O�i�Ȅ��%3��œ@X^\0�'w���B�N�2�c��H-HјV��	ܼ����D�Ol���O��$�O��D�|�D(��r#.���̕c���u�ˎT��V�G P�I�t&?5�	�Mϻt3�E�ǋ�^x���Y�1��H"�i��6-�g�)�}���'������ wP ��ֆK���ٙ'L�A��&C?�N>q+O��C���Щl�6�i �O@�̄�I1�MK�d�?����?!Sb�"7��+�蘔)�.��@?��'� ��?)���J<�s��[�x�0�ȇm��)�'6������1C�t�E?���v��ْd�E1=�����������?���?���h�����|��ֆ�+��`�'eŦ]���d��e��۟��	��Mc���4���Y�Zφ�j��� AV��g��q�d�5�4A�����?X�Iퟴ���\�P	��B>9�,�W#T�x���ȓl�)a��O����O��xcaE�7�|K�-�JiP��0&i�n�r�'""�I[�p�P�����l	�@Ґ�'%�6�Ц��I<�|b��<ک:� 1wڄEJ�>,������/{��@��'&�'A�	<��T���*7.����N�f��ݟ��	ϟ�i>��' V7���F2v���C�pc�$F�&h��
E�g2��d_���?A�]���	�0sشp��U�7$��]����Ŋ�Q����d�,��Q0��w�����>��=� 4�y��^�d��Rd�T�{�2�+`4O���ć�K���+�gT 9@C+-�t��O,�DU��)�a�3B��i��'3�Ы��wP`���ܨB�Jt�(�d���� ��|�G�)��Ax�s�l�2T�:��,�z���O:I��ӟ�����O����O�dКk7���T�`i���w�W�\��O˓)��AC"C��'��V>uQ4HC<uhe��bݪ(3 �-?Q7^�����CO>��?M+��Ohf��wb	,k�v�x�eL�b�̓0���"��*��O�.6�D"Zz2��@�},��SC�Z�P���O����O��I�<q0�iC�pbQ�x�U�e	O,-�m�5vR�'.r6�$�I'���b�P���l��=޲C �0o�� F+�ڦ��ݴC��1�(OP��ޚk����	�0{�b7�=����r��O���	hy2�'92�'���'n�U>�Q���%f�8)�N�)*f�œd�ې�?�� ӟ��I���%?�����M�;rߌ�bgd�fL��צBTD#��'u��1���tꖎ{��I�1&��F�΃q����աbgt�� j�� �'X'���'�r�'��l�!�T�4⣣K��Mˆ��O����O�$�<���i ���'���'4.��k�=+h�{���;S�D ��F}��'�"�|r�\/D�*%�qZ�
��DT"0
8��f?�4�H<��'��NײO�a��L	�V�����l�"�'���'t��S�����'�0s 6@�&�6/|Xزg	�ޟ���4hb�����?��i��O�� ]Yܙ���Y<I�2�@ڄW����O�7-�A��ÝF�@���O���խ�.T>��q�)YO��!�Z͟��'C�i>�Iȟ���ϟ8�I23�(B��8~�bM`����Q�ba�'��7m�'z�"���O���<���OD��d��YЄ�tO���D�*Bx}��'B�g2��!j�����e�Z6���n���(�1�J]���	4-[��3��u��|P�P���="���'\�0lni� Hɟ��ɟ �	���pyBKo������O,��W�#Nm�'mD	O
����O~<o�A�F��������ğL��g�&"�ht�S�ը��̚$�*>O��'�bo�<k&��`���� ��/ N9���-%�9��;>����O��d�O*���O
��,��@�R�	�p؄Z aH�#q ��	џ���&�M��C�|*��!z�֙|"A�_������^�&��1
g2@O�o/�M[�����,O �����$��ԭYA��x�v*üZi:��5E�+�?�h'�$�<����?!���?��I͸�	���J'�@����)�?����d����#v@\Ο��ßt�S�?�V��QI��H ��<@��1?�#]�<b�4cܛ64�4���ɒW�v@��	(4��Z2#@�,���V�L�M#���ch�<Y�'"�.����O��C�ǝ@r��[�l�&a�(�ON���O���O1�(�*]���U�l��Pa����v5B�B�:0��f�'��E�X⟤ۭO��oږ�B� 6+_%��U`�gE?:��ts�48ƛV��\$��柌0F��$��dfEoy�Nٜy�Y�s!�nQ��x���&�y�]�@��şp�	���ӟ�OO4T��+�&a��}�f� fy��1'`�,U86L�On���O����D�Ц�*2��(!O.g�j��$C�K\b�)۴{$���9�4���i�����d�<A6f�'BK���� �I� \�0�	�%"l����']$'���'�b�'Զ����Y�]`�T5i�~4V�@�'#B�'�rQ�|��4C����?�����)��/�4*&�I�4����H>y��Z��I�M�i�FO����F�N%�ƨ�8����8O�Q��4Aa���O˓���<�I�q9��rC�¸i��(p�@�,[��\�����ʟP�It��y�&�=Oն�1�ɓ8�,��d��`�h���O�$즥'��s����]�o8��w�J
oT�*vOf����43����{ӆ�y@4���7N�0��'T�}�c��FG�q�"�M5<�TRd�9�d�<q���?y��?����?D�Mo��(�I�t�}�Q	J���$�঱�'ŃLyr�'���^>q��H��IR��K����+"����OXn#�M[��x�O���O��a�g��1�&�[���1;SNöm�RU�<"��L����#���<YAZ�{��piEzH�!)��=�?����?	��?ͧ���ԦA�C����s��I��P��Ô|J`Ѝ��H�޴�?�J>	3Y�H�	֟���15({P���0�����:I��D� y��'�$�[�l�E�+O��I�Ԣ�%P$,��qH��+�(p�78O��$�O��d�O��d�O�?tm]�R��J-+���������ٟ(j�4ydyϧ�?���i��'����S�m܄��h��ƞ|��'���'���X�^�0�'40��b�O&[�n,Hf�&h%�Ɋ'"�-�~�|�\����������� ����?�;Q�/N��ek�����	~yreu���!p%�O����O��'+M�=�c�
��ل{�(9�'����?������|���_���A&�f�@����q\1���4���O���M��D$��S񆁠s?���b�Σy�Ib�A��D�Iԟ��I��b>��'�b6-հyT|H�4��[
�/A�>����SE�<�զ�?a�[���I"0�4��B�6$�
0۾e��t��ȟB��ny�П������?͖�� �J+��R�M�싽;vL�x17O���?A���?Q��?����	A�ߒT�$,�a���JgfW)?^h�nZ'�U�I՟��I@�՟  ����3�"Z5�|�B�(�CJ�?������|���?��&��
�(C��b�Ꭺ&��$y�b&.�d�*��z�'��'x�����I(��h��DU�|c2=0Q���T\ @�Iݟ0�	ȟt�'IN7��D�D�O��$H���0���!��<��� 
�xH�O���O��O���&^�e���[ÇQ�~$�-PĞ��鷃O;�tZ �>ͧw:�����Č�~�JDy��gyt-��?v����O �d�O ��.�'�?�'��:�t��-g�8��2�G0�?Y�i�� h��'_�dhӒ���q�:@P�a��LH��L+�~�	��`��ş�p��D�I�t����O�:�`-���N�[�h�`�ny�O�R�'���'�RJ��y�~�a�Ԧ<0�T��.l�剆�M#����?���?QI~�� @�T �Ϟ
g�"���[�5�tq�P�������%��Sޟ��	��nXP�J/BN��We�3�ZM�PJ�
��Yg��
��O�7��<1�ΕT?��q1��/|@����ׄ�?����?���?ͧ��$�֦��qLȟ �iP�5�Pё�Q�����Sҟ�P�4��'��ꓦ?1���?)DJ��h��p���2.��CG?+%�M�(O���Y�"�z�'���?�]"L(,	�ًkV�b�䍈#H�ҟ$�I���柰�IO�')ҩ�"���`�RЈ�U]X����?�����& ޜ��I��$��:F�<^ ���S�p�xb��h�I՟��I���Lny��'�����ӳp׆(�U/Y�F�(@��kʄ7n2)�	�[��'l�i>��	��\�ɰy9,}�oX<}�8�4%	U��l�	�T�'b7mP�3�N��O��d�|rs��<Y�T�g*��!�4�H�a�O~��>I��?��xʟ�(��A�0R�2�8�.[9x����"1�dP�����i>m����u��|�M�~l|�!�Y^�����U�1��'��',��Z��۴j�X��s/�7@��:p��-5*�+SHΊ�?)��_�����i}R�'��9H@Z�����A��^N�"7�'?�7��%g���?Y -C�|}T��,}r�ӱo��y�s���L�
�P�yb[�H��ȟ��	���	ȟ �O�te�V�:�^E�!��?I3I�/tӲ�"Q��<�����?T��y�%w���ibm�
0T�ك�G�R���'ޒO�I�O���ʀQM��2�>��U�)t�l5��ĕG�ϓ^�����o�OV�yL>�/O��O6E�F�Xp˶�$I�Z{�1�J�O��D�O��Ŀ<A��i. q���'��'��㳧ߙ3w�2�Z.�����ĆC}��'�b�:��σ7�hal�2tp�gx���Ox(�'D>�p�O���Ӎ9Zw2�AK~��Ʈذ,���ä,�7I���'���'�"�S����a�T rjP�E�(|c^)��OʟԪ�4Z����?��i��O��;/���ȇ�
h9P*�z\�o��l�1�M[恏����O�R��:�����E�`��[dIsQ(���UK>Q,O��Op���O��d�O",����x��X6��_� ;q(�<�g�i,�4�'8"�'��@�"b�}�Q�C.˜.!�{e�\D}��'�2�|�Ou��'���ÈؗEے��%jRj1�A���V8*��U�Of�d�-�?�;�䓶�d5a��6�W�o�t�(Ѝِh>D���O(�d�O��4��ʓO0�v&ƣ�R
A�3�B�h%HƵg)~��b��� l���
)O|�Dt�^)lڒ[B6Nq�}8�Č� ��J�m�S�I� ��}) �O$q���.�i'���ᣏ�:MP �bV�r����O`���O���O��)��?qT�7��D����ԏ՟y��e��ԟ�	2�M��*�|���<ț�|��&)8�a����%����l̢Y��O��o��Mϧ"��!M>�u��0��S�nZ����Պ�#h\Q2���O�%�J>*O�⟨��\4c,E#q �lgF�x5`>����U
r�"�'�2S>	`�EO2��惀 5b$ 5�=?1$X� ����('��'��A�"E�����6,j*�낺�dq�����4�FԂ�' �'5XL��S�D� ���c`�q:�'*�'����O��I��Mۗ�Q�;�.yU��-�*u:�n	�U ���?��i�ɧ�4�>Y��*Tf
`�z��1�
 @F� Y���y2��
��Ӻ3��ٹ���\���D��~���(�֫@v ��os�T�'���'Ub�'��'�������N�i�$�*O�b4R��Wf60������o�S�8"������Ir��Q��,�h`��@��?�����|���?1������$��\`=K�l�0C ]�"��:L0�dֳC�b�'e�'��	ٟ���r�x؁"��q0<l��� `���ԟ�����Ȕ'n�6-\��d�O����<i��[��$�U��j�5|LN�`��O����O�O^�� ��A�Pr�M�
���P����L]�.�����y�1.����O���B�#�6�J�Ĕ�LF$�p��Ob�d�O��D�O,�}���0���Td�ȡc���J�h��[ʛ$�;��Ŷi��O��X�B$�'(���yRA��$5��$�O��D�O��!H�<I�k���H$��v�� ��@��T9�^E�Ď� GD���.�$�<ͧ�?����?����?�"�Z/|�y�4E��tp��k����$Ҧ�B�@џ��I��l&?���9'�̨�*�.�\��V�I�y<T��O����O�O���O��䙐4���)E��D+�"�xd����/�O��P>���K���$�ԕ'�(���C8������4���ar�'Z"�'Br���tW���۴m�p4��`:�{ Ϛ<eVX`"GcO�~�+��ܚݴ��'���?��e8��\57�ءx��ՍR���`b�����|Rb�
�A�SK�'��{#h�f~�P���I#?ӄ�i�j��<i���?a��?���?����ٝ)���J�֣�e�r�ݎ/�"�'��#~�>d���<Y�i?�'�b�Hq�[�"��`E���`����|B�'R�'D�*�^�8�'&)|]�pΐ�J�lsԣП,D0RR��%�~ґ|[�p�I�D�I埀��Rx�<�`@A\?�9�M��t�	my"x�v�d)�On��O��''�N �Gџ@���`�� �J�`�'2�듊?q�����|��\��A��R�6�`҄T3~|P���Ñ.��L�����������'M�'c(I��)����� Oh *!z��'��'B�O$�ɗ�M�(KDȔ�ՎM�l�dY�M	�Q1܅����?AW�i�ɧ�D��>�ir��R�P�?�VTi��O:"�|�)��p�zn	Sح�'�2�І?�TD�'��̕���[`NC:O���⃋/[L�D�<q��?���?A��?q(���1��(<fb9j��]�0 U��\ަ���l���I�H'?���M�; A$5w��¯�I*�����?	K>�|
��E���ĉ�nMj`LP�U�D u��>7.�֤5�@�j�'G�'��i>��I�O��S+]�;�1p1`^4]x��	���ʟ̗'��7m
�@�\��?V��"g욐hՠ�`�+���.���?	�T��hߴ&��� ��*:���`'��(9N(8��D�W�IQ�r�*�噠j�0�%?�2r��u��'e�R\tZ 5(���)���y��'�"�'���'I�>��I�~x�qJ�#�2qoD`��&��y�I(�M�)ƈ�?I�3���4���S'�/'O�US��Ҕ��<J�5O����OpEm>K<0�'$�)JX^1��:���b�#֭?�r���	�O�D+�|�W��ǟ��Iן(���x�I	d��82�߁7n
̓W�cy"�oӞ<�G��O���O���d������ƾ �� q�'T9Mi ��'�7�JЦ�"O<�'�*�'"(8dSte�[�I��Ǩ�W,D��?�/OphؖC��~b�|�^�8!�ǘ#"G4X2�Ӫ���w�ڟ��	ş<�I���jy2�b����N�O��Fgӻ8�*�pf(?bƴ3=OB�n�D�I��I��MŲi� 6�ߕQ��!@vC�		���qƈ� u%�P�*�<1�Lp� g�?�'����wj�Hq�P�l�{DJߩZ�}�'��'���'2�'���䁤��1~F���-Nd̑p���O8�D�Oʽn������'�\7�<�$
��(�d���2���a��P�T'��mZ)�M��'(1���*O���
�jϨlY3��$j�����Y����/���~R�|�T����ܟ��Iڟ`C�$��-�� �0gÌd�����Dy��hӤ�҆C�O,�D�O�' �q���� nQrܫ���(_G�y�'o ��?	�4�ɧ���|0p���mS��ɞ�&�FQ�8u���[���p�>�Č<	gDe��\k_Ft31�
�+����O����O���i�<ђ�i��a򉞤tǾ�c�͒&���i� ��&�B�'�R6M>�����Ħ��s/=*����E�
�TARRk�2�M�W�iw���0�|"���4ڬd�'���@4Pak�.��7.������t��<����?)���?����?a(�.� �K��	�F9� b/W�����lE˦	�Q��iy��'�O�R�w��n�Rtɸ���dn�P�Q��xͦdn���M+`�x����*I��	�x�F pG�G[�)�����I��ps��O��O���?��AB<��⏬c�ԁ��_x�a���?1��?�.O��l�E0�@�':�-ϝ*(�xFEM�I^����"��'�$�>Qc�i�6�K�pФ�EF�
 I6�(�ȑ7 b.�@mh�J
8>@�\2I~��j�O���O���F׾R�9���J�a���8��O2���O��D�OҢ}λ}���+^Z�9��5,Ҙ`Jwa������4�������?���i�ɧ��w�Z���iKL��K�m��X�5�'x�6M���eܴ"f�HK>�&�U#ʈ�i&A��a��`�����4J���^�YN>�,O���Ol��OL��O���V$S�q�X�X��<� �i�l�OB���"��T� ��s����̙q^�U�#l}��'���|�O1��' �	k�Ô� ��,��`	�.bv�U�6Q�'avm5&w?9M>1+O���H�P~biK�Ŗ�!.t��PJ�O�d�O$��O�ɤ<qջi�M"%�'|�i���&C8H��)�#%����t�'�,7&�4��\�'���'Bn�$�r���<��eQ�x�X�0�|�eј딹����'r�"��0E�:
.���q$�8e�е�I	�O|���k�<��[A�찙�G�0�	!�'�6q���K�/̸:��!#0�Af��@d������-�l���rzf�r��S�<aX��C�ί82Z=�G�5?��ǘ�]w�HsG�=[��ژAN�eٱf�3}p� X�D�O��]�%�]�_����f�4�ߒUf��3c�%р ��Su�@�,��A{W�-.Ş��B
=["4h���a��B�o�57`� ��G�0͠����':��	�� ��oO�TkvcH�Cd��C�9����i���'aB�>T�����O��Ɉ*,2H)7��z�D�p��LNxc��1ӦS�	���	�ȰN�|x���HW�<VP�!���M���%5 슥W�<�'�"�|ZcDX��'����O]$	4���O^�8%��O�˓�?���?y/O��!�ǎU�u��o��r�@E8D \3���'�	�P'���I��@v��:/���F�@��5q�-�(�$�����x�IKy��4KF�S�>Q��ҵ-�W;6���A8)&6��<�����?���?���'!��W��E�&�!Т̙�@�"�O�d�O����<��Č�E�� �G-�5�P�@GDˎ|��dP���Ms�����?y�
� 5Љ{B� %�>�S �ڙC�<1�W��M���?1+O1q�]R�$�'���O �Hl�l2l�!��ͼkq�qq�&-���O��H�
�㟨��3p���%=A.L��خ}>�nZAyr��p7-�O���ON���n}Zc
�}
Q�]��V���]S�LE��4�?��y��(������:;��T/M&}ؖ}�E��//țf�\�7-�Ov���O���R}}�[��%I�u�Q�e!�?u�rH�j�M��K'��'T��������bdW
h�&�L&c�>�l���I͟��$���D�<1��~�c��y�	k�g

v�T!�0	Y���'�D�Xd�|��'�b�'��u��hԹPT4�h%d[�z?v��(l����U�a�'��I���&��؇#6��PAK9���ZPh�=Ȭ�A�yq����d�Ox�d�OʓA]����1F �
� B%
$�1�&gJ/U�	ay��'��'��'ި��F�r#�Q  �F0L�x��J�sh�' �'9"R�@�ˉ����C�!�
��'�
u|�z!���M�/OR��4�D�OP�Ē�8��0�޸s�BN��ҡH�����ꓖ?����?�-On=B"��z�S�7�����SX�س��0G��ٴ�?�I>*O��S��O��O6rl�F�'F�
�IRM�}���4�?���dó+8�@'>����?�؆p}����b2|Ollq�^CRH6��<q���?�qk	��?	H~����aπ	��!@WMD�=G��{@�����'��i0r�}���O��O���gޤ�ɱʣm-��H��E1Pp�l�Ty�͋�&Rb'�i<��iy�Ȃjԕo��$_�V3�5I�4S���2ǽi�B�'I��O�O��G�9�0�6��91/��	c���t���nZ>3v���ٟ���ߟ��S��R>Ya���N�� �#�����hۛ�M#��?y�Lبis+O�Sv��ma(�e�̆:
j0�C��H��m�<)Em�7C�Ow"�'\�-�a@��V&F���E�� 8��7��OH-��(N@�i>���ܟ��'�)���%�v�`f$єpm:-���t�<�$_�k����<ͧ�?�*O���8�d�b��=�Di��.��b�o�<���?Ɉ�'b�i��(��ˌ	`uѕ$�=D ؠ��P��d�O����OTʓh�,%B�6��Ly׏\n�}��@'PRF0PtS���	�����by��'��! �" ��s޼,�U�N�$x%eH0IN���?9�����O�s҉�|���h^L*u-�&Q6��C��bU�БB�i��O����O�rB��9��'m.��EC�A�>��B�
-X���4�?�����D��&>����?��	xqv�# N�0ia�-v��#X7�<��?I�E���?IN~���C6[��^Muf�o%�hJ��Qަe�'�B�"(sӒ��O���Oh4�A9��gB��`A�S&@':7UoZ��I�t@T��ɫ��'�(����>v��1���X�m�>4cT 
9�M!�9?����'�r�'��d�2�4�k��YP�!1�ω�e�|12G�H�DK��'k�'��X������N�2�A�����RQ4��yo��8���@���Ҍ���|����?�vLU����4��Ri��!B��Wś��'�B�'I�	3��~�'��'�*J I�pk��	)^�"��A�i�F�$N�S��5%��̟���{yJ��,����$�F]�W��%t6��O��9]��|��'��\�XX�(�	`�\�{#"��Ԁ�?~� �I<���?Q������O~��QBv�� ���I������ӡR�E�G'�ONʓ�?����?1)O
�!v��|�e�]�K�FX��+��s�9Y�fBD}r�'(�'�ɟ����9 "��ie\H��G�l����B0Z�؜��*�>i��?Q.Op��:ns��'�?�ҐM�i�D�E$1-I"fJ������O~�@6"�:I�xR�[8�NP�p������C�M����?�+O���-�D�S�� �s�	[a╕zzݰ,C�N���17�!�$�<�C%	�?�J~��O����B
I�0�ֱ0)^0��O2�DO����D�O����O��)�<�;l�
<3�ʑwRtJ��lRTIo��D���N�D�u�5�)��|G�d�A�F� �̠x�I)U�7��%\<��l�h�����S����|*��+�s"�	aa����,D)r̛&O[*{`��'��IN�4\�x����tC��8�b0k��K Q0"��ݴ�?I���?IT
n���xy��'�����eJ�h�A�5(�rU�wn�&Uۛ&�'��'׆���)�O���O�)��cת��2��N�%|q��o����	w�<r�O�˓�?�,O����� DQÊ����p{#f^�-���a�i����y2�'!2�'F��'R� x�.����>Af��A�ԅl��E���°���<������O,�$�O]i6i�)���aj����lP*6���OB���O0�D�O�ʓ^��[�:�v�b��&+k���ab
Ѻ �iU�֟��'Tr�'[�'��yb��1�Y(e�8.�����W�V��7��O�D�Ot�d�<�6�Cc������<�:�I��1X��%5����7��O���?����?IwF@�<!���~⁘����!ȒO���r�A��MC��?Q*O��2T̑D��'y2�Ov"� �aš@˪���4�v��!"�>Q���?��v����Om�IH�QjK�V�J�mǉag� S�i̦i�'j�P2�oy�(�D�OT�D� קu��P&a�ƠCf�ӚW�,y���M����?�F���<	���-�ӟbr�� HW�V�y�rE�5QX6��<J�n���p�	ԟ��S7���<ɒI��8��ńL��i����֏C�y��'l��O���?��Гr����a�Ǚ}ۨ�CFbR�9 ���'8��'��#�h�>�)OB���4pg�Np�,�����yd�2�`����<���<�O��'�r��9j>��s�]�B4֭jc�v��7��O~��D�z}�[�x��wy���5��E
1�~�����gc�K��,����T,���@�Iٟ��	|y�k�hdr���O�0Y
�I��E���F�>�.O ��<����?	��S�!�����Q���ly�H�<)��?A��?i���$˪pF�1�'F�œ6g���ة��B�6v���lZ{y��'��	��(�	��@CM{���WÁ?RӨTã��211�Q'X��M���?���?!+Oz�hrjDX���'�H}٤�C��Ai��N�^���O`��d�<a���?Q��&S�@̓��i���j��B%��t:���+x�^�r�4�?A���L�в8�O���'���ɁD�R�RuGS� ����4�~��?����?�����<�K>Q�O�	HU.ř9��G*��o)0ݴ��č�y�HqoƟ,��ٟ�������Z@B�k�v��l0&_6v�z��i���'l�@ �'��'q�X�k��)����g$)�v�j��i3����Os���D�O��d��I�OX���O��"WMV!��;���>�h$��n�˦�A����p��͟ s�������^�]�^IӐ �8-~Ъ�4T�n�����ϟ�pT�
 ��$�<1���~����ov�y��. �@i����Ms���dɢ:�?	��؟���o�D�������3�D'CzX�"�4�?���A��ky�'��֘)f}�)�5��I��iЁ~���F�����?����?!��?�,OԼ{!���֤��R���	���b��>�,O����<���?���2��"`%ܰRn�)����QX�dꄦ��<!-O4���O`��������|���ʛ�j��?
	�౱�Aئ}�'>bV�x��ٟ��I�`~��I�76�-j5�<�p�g�4��0[�4�?I���?�����W
���O�Zc���$�
�3�~uv���@���hٴ�?9)ON�D�O��d�b����Op�Ċ������.��r�pcw���dZ*�n���|�ICyBl�K�h꧂?���"r�J(�H�ʰ�
T!�iـ$	*6�	Ɵ���Ɵ(���z�@�'��֟\�cUR)�@2�NW3zARb3�i��Ʌ[�=ڴ�?)���?���[A�i�A{�A9O�$rp&\�>)(��Gu����O�0OΠ��yB�	�t���	���%���
�j�����%2��6��OR���Ob�i^}R�@S��L�1S��C��E鹄�	��M�ah�@~�W���R��vc ����#�� b#O�C�^����i���'M�ҭ�������Op�I�	�����H ��6��S�$�6��O˓w��S���'ur�'�� 0W��4H�r��7�a4jx����(\~��'���۟��'�Zc��a(�'�
N�x�k��?ɲ��ON5:O��d�OB���Ox��<��	ǐZ @dE�Z��@��Vo�iBQ���'��U�����4���6O��@�1`�j�nQb�:�
`�c��I����	���	qy��2NR����p"�Fr��)Ë&?�7M�<Q����d�O��d�O�ыR7Obi��V�F�\��B �d(\Ij7����	ԟ�������'�S�n�~2��+��m��L�1U��p�7a��9�	QyB�'��'AD�'G�s���P�'����@ ��&z[�9�@�i#r�'	��d7n�����O��IC�p�K7#�;�����F.syR��' ��'cr�������#�0�y4��+A�$Z&7��(nZFy2h67�O"���O��)f}Zw�B,�K��vü!X��Y6=S��i�4�?���S���ϓ�䓅�O��0���p`�g�N�4���۴&|��Xưi���'���O3b�� �!(T���Ͻz��}+�'��MKD�<�O>)����'ц�Eē�\}�1�f�	�Iz\x��m~����On�DM:�H��>Y���~B-_�[X6��֛7��cI8�M�J>q���?�*O��d�O����TmZ��D�D,Lh�C.:h��io�I	5xO���OH�Okl�?��e�'+�-���2��?��I�4�i�	ay��'���'���r��HZ�m�/�luva� <��Z&�����?����䓟?��=6Fd���)/1����q�*�2�䓊?����?�*O���@��|
���%(��`��5ne��L�h}b�'�|r�'��h��$� ZuX��ՍO��Z��%i�x�qY�d��ҟ4�INyr�S���t���ЁF����a�}�Bm�Wn�ߦ��	t��	�����i�$A<���2�ݷI�x4���qu�f�'"Y�������'�?)�'�d[� �	,�����Px+���f�xR�'���߮�y�|�ݟ�,K��7"P�B��M%j2��i(�8�v�0ٴXJ�П8�����ÑzdJ}���B�@����&�G,(7�F�'��%��yb�|�iV�J��pI�CR9i� �F�(8��( �.jp6�O���O��I�N�I���B�n�z$�[%"�d�XŴi.\<��'��'�Z�$E�֮5��oW:-����E�8m����	�����-��'�R�Ov�ꖤG\�  & 9eX��ӳi��'���b5�'�i�O��D�O��'&U�8Ј����G�F#"�Ǧ��	#q�:���}��'�ɧ5F�Z�J�q��/{��,٦�Ǯ��$�2+��ĩ<����?�����$� P��J�>Am:�a�50���1��j�I����Iy�	�����<ruC�%���w�99���r�v�@�'�"�'�Y�0�1�$��$��5U��"/\����C�����?�O>����?�ъٯ�?���B$9<IC�л_��Pr%�+�I�\�Iß\�'`�,sw% �i��F��P��$̠|��@�bJ�?A�doD�'�g)m�B�'N�$ْLЙ��F�e�*՚��$13���'�\��fHI��ħ�?���ö���`rDE�k�5�\0bǧE쓗?)C�ߔ�?����T?�%y����h:�>e!G��>���rA���ʟ��I�?���u�]�Bm]�MIq)G-� �4�?��Lݸ�Q��l�S�q$�M�LմN����B��M|�o������4�?���?���OӉ'��m
�j"���/�#���6Ɂij�7��������	�9�v�ݍ{�04q�f�ZP� RG�i�b�'JR'��DnO����O��;��M�fg�	�i�^]0c�ЊFJ0����ܟ�ۆa�A�T�I$*Z�v�&]��P��M���X�D�,O��O��|�iP�N�T�!�NYe-X��.q2�:q���v/�z~��'#��'��I�V���*�ڶYF*Lywd�$J��m�4+�����O>�d�O��D;�ɹ
�6dy���VT������@�D5@���S����T�	؟��I蟈` F�C��O+y�F�q)�e��}��'Wݦ��'��|"�'��E`
6�=\ Z��f
ܞ]L���&��$n����|�I�� �'����3�~��\ ؐ0r`�3N�x���9*k0u�s�i'RW�T��ܟ��I3D��Iן��I�� ��!z1�i�`N��]X��M#���?�(Od)���H��'{��OB�A�*iT���OA�a�	�%�>A��?���V����9O��ӵ9{,9߻D��}�%W�6M�<��-W����'r�'��d�>�;jP&xC�L�}�d�!�"^}��o�ğ���u���	|�Il�'G�������E�,�AR�2g��n|Az#�4�?���?���g��dyR��!I�P��$fʜрӫC�xl7m�%���9��3�SП�Bd�v����_�a��iB���MK��?��i池�_���'�r�O��	Q���
�����HA�Sp�"&�i'�'ϸ��S�T�'�2�' 
%�B��]i!�/t:H�b�
b���D��g��i�'���ڟ�'�Zc������w�H���47ڒ�!�O��h>O���?����� �e	$��+u7���iT%!� !��<��Ify�'j�	��	П�ap��-f:���ڗHrƜ���
e5��	Yy��'��'e��'϶�1�ҟ�y�wi��*�&�X���7-���E�i�r�'���|b�'���\��ݴ���3�i�P�z���&H{8��'�R�'U�Y���/0����O����	�Tt"1�Ye$��`��@��?����'��x�&�$]�d_�����Dku8L�t���Ax�F�'�r�'�"��l���'��'�����(Ⱥ��W����@
���(��Ob���OҬ
�(a1O��;�Є���LaK:tH��	�Q�6-�<ɤ�*XO�f�'���'����>��u�f̩PhÑ(p���皍m�To�̟h�I�nט�ԟ�����0�}
���� �ڜ w��>r��8AU�y�`��/�M���?I��:rR�X�'7�������@z ���
%eh|�tӢ�<Ov���<y����'�4f녺K�H�G���r�2���&u���d�O��_v.��'K�I���;��Qi��XA�ă���rc�4n����'�x�����)�O����O�Q��#Ρ?WVx*�
4r�Lh�&JEަ���a򐠚�OD��?�-OF��Ƅ	�n]�Mu>�B���5hXpek4V���oy�\�	���	ß���uy����^��d33(��Z�~p15A
>��%g�>�.O��$�<���?��"8L��[2.j���Պa_��٥�L�<�OB�8 F�
I̠��ooj	;����BlV�:��x�	�;�U���+9|(��O�-���"]͂��U���������K
K��q��n��@4��l��k7T��l0�.���H�_�(J�+ؓH��:��י��	�D��j��m)NQ�5ŔMx3M�?7|�e-׍t�<���ڃ9�<�Q����4��� � 8�4�
#"�].���SJ�X2�P"�j��1N2i@��� �PY&�E:��{�N;dM'�"��A�E��p���m�X`R�'N��q��
����W �j�r�X�.�� `ts�L�-%Z3�� �z}Y��>����n�I˱D^^�D����T	*�CC�~2��ƚE�P��Q�Ӷ.��p�t�D��m}R�'4�>��>	|k�$�J:�"�F��=��C�	�]t��Af�	�����R�r�h��$p�'�V@��`:�6�X;�*��ei�>���?I�BS�>��pQ��?����?ͻ �����H�} e��ѿ�@z��:X�F����&P�g��83� ��Aj�7HC<Ds$̀v�1��.����:���|�� �~�%fX3=�BH��Z8}�����O�	=ړR���vbZ�<��	tEW:7?���ȓ*K�Ĳ2��4Rc�NQ�;����'��#=�On�ɶ�*�zs�۬2�Q.SZ�Y!w�*Q���Iڟ ��џ�z_w���' ��b��C[�[��Q'�]"{6|�8��K%JQxe�׏݄A,��ā>p�D���C�-��
�cD� XJ�g�{��t� K�24W���{}֍Is�]6�V�8�]�=`(���'�r�	}���Y��bT?d�5�WN	'�8�ȓ�� ��=)�b��ë��h���<)4T�Ԕ'd�x�HhӮ���O�<��t_����AN��Da�`%�O��d�����O��B0�m�_�"6	BW�n�4�;��B����$T�'�lc������8Y:��1��9�E?O 0�4�'�rT��" ��oDP�`��,�k��~���	ş��?E��a�[�*I� \1�qrwJE�xR�~Ӣ,h��_6�@x�$��*%�AJQ9O��?T��Q�|�IO�4gŷJA�(қo�@�DH�V0��I��I���'P$ȖEV�D��٦� [���T>��OH�@!���",U���T[R�r��H�b�í��}s��F��/�Myt#Q A�"h{%�����ɛA�P��O��}���X��p��ؕ��]�%�O�S��d�ȓ@
T��"F�����oֺ8� 0����HO�<S��&0��� �<8�@�Ӧ��I�|��.~�yR�
����	ğl�i��C�LX�
B�K'` �]dFc`7>�\c2�	 Mk���I(����|&��1"g�=D"���Q@�.V�de�O		>I��� l��Z�[?{�X�>�O�)H�� �`��oǬ?�"�#�?�	�=�*���|��ī9�,`�Z�q&��`�`���y"���e��	@%�,�9�V�������8�t��cM�Y�JVW��\�^7Af��$�O��D�O��dB޺S���?Q�O�������=2�:i��j'	@9���O}�|��Щ:[˸�3�}Ѵ���I��m�L���X�*���qB�X����p�M	�$E�q�A�@A�p�'%��6�"ؘ���-%�����m�e���$!�O�!�X+y�6DhCJ������"OF�Z�ĵd���(ЭQ������R�*�PÓ�i���'���e^2~^����.�#0d�����'NbڑM���'<�	*O�j7M<��V|"<��'�1a��}p"j �_i�x���Y��O�A�W�Ǎ^��a����F���"u�'6x�����?���?iwkʱUD�p@�,��I["�W����Ob�"|z��T9T�q���A�p��B�n<�`�i:p���F�a����Д
�-c�'��+kP�ش�?�����[ �`�$�#D��+��F4� @�O�&ky����ONX:��O�b��g~�r!���c �j(f�������	�C��"<�*tnW��@* ���dF(��'�S��@.c������~ԉxu��b��T���ɯB!�$.l�~8C�^�b #̘6.axd?ғ��%��ףiʐy
0ş�j�YгiX2�'1bA"-x�H��'��'�w�J���âS��a#�
c�-��
U��yV�en`��%"&X��ǝ���'Tr��ϓ8?�`��(S65[������5��yr$���?�}&���1B�w�LE@v�#	�hX�0�<D��&U?,V	Ѓ�@�^�[#�4?���i>}$�T���@�r�P���o8$s��/.k0� �@����I柼���u��'�?�6��B��8D�����՜y �xk㄁TN4���'�O���r�*s�p��'.ؕ����QcL$�'�pA̡�A'QTX��hF)б�B��&?]8'��u�
��,�O�iSPOB��15��	�����'w�'B4�BO��n����l��]~���yB�p���OꄹaJFA���'��P��DO+>���I�,Ȏe<��3P�'_2��D��'��)�3�r�K��ĆMYNz��`�p� � ��m�(�	AD4N�jP��'p�7�Y�&�x��Rk%kV�� ��������wB����#$�'C����?�)O^���C�;�� ����m�|[6��O����68ƅ;l�*)��qr��+H��G{�O�7�D�#��Уu�ݵv#V(2��"0N��<�f�Ʈ}@�&�'	�]>u�1�ʟxX��=5�"caD��ȩk��ğX���w����z�S��Oڐy�%])*OpAi���[~�)3�>��ȍN���O�� R/[���eNoo�٫N� �j�ON��O��� �ӓ��1���&�h���p�c�X��ex�hK�Ď�Y�,Hu,�}����<O�1Ez"Iӧ]���Fcý+rp�w��^�66��O��D�O.�K�4�����O$���O�N�y����˹e9�L�*�2$��@����v�h��4
�uSF"�F�g�I�0 ���B���f��s-9`?�: �=D-���i9p�l�h�g�I4n'���E,��Oǘ��UhV�i���<�hV̟�>�OȜ�Ѩ�+q�bU@�d�<|��t"Olp� ��dG$�K'Cˌ�F�w���Y����~?^� �l\ �N,�f�+sH��A��Ň 8�a������ݟ�^wS�'���]�!"LQ�Cn1:��l�r.���aO�퉐��M��� Y�)��(���!�d�M�N��B���jS�,+ᡎa��y�'���-��C�Y��suB�y�o0E�����ѡ8p :V�[���'ǎc���!�O0�Ms��?--4*\[R&�:;&�)�a�A"�����,��\����|b���+{����b�ȹ6sb�HѤW��#G�Xr���"���9 l��d�"T-+�4q	h���F��<.��hi*9��@�-ڕ=u�m@�%5OF���'@�'*IC��	@�bSń*tq���'>,+тL61�kbLǰ�|��'��7�+|<�,�cݤ-�aj�"��u�1OV4�t��ʦQ�I˟h�OQTp T�'L8�S��l3�Q�w�ݪ�����'�2"�.MCb�T>�9iX���̏�2����"oF 7zrȥO8Q��)���Q(�)�N�=E����#�_#.t�'�����Θ��O�.��cZ	��Ҷ,͡q$�'�Ƶ��nI?1R�%�Q�@|��A
�
����KUA�k��X���٘/ΈtK���?�MS��?��e�q˖B��?����?��Ӽb�Y�S��[f匤y2 @Ǐ)��'>� ϓi� �ӶT�܉`�	�Tm�=��	^x������+�f���d�p��m:S �G�s��}�)�3����c=�(��/�(�  �ߥZ!�$8k��DA+ׇ)�D�ؒnY&2
���HO>qj��À;�� ƃ��a���^.Y|x��Ο|�	Ο4��q�$�'X��C�/\R@�e��!1��Ų�A�:u�x�Ɇ�)�O�&h�#!��3Sh[\:�T;7��i�<��r�ݡ�l���'�^}!��!��=bh��3� ��	1�?�2�id7��Oʓ�?ы� ,�0���QU<�a�Z��Oʣ=�O۾�P�F]�e���_�T8�����|�i،T�7��<���	�A���O��7i����0+T��͘w�R��z�D�Or@��	�O6���O���C�K�C��O���0䘘t)f88)�K~\h"s�'&9���V,sal98������'ǊPv9P�C6j�d��Q8�D�� �O���W˦Q�I.aE�l���Y�F6��En��_�<��'����SJ�����Y8?T�x��]�-�T����O$�n�:" d�Z�L�4��`A��G�j8ڴ��d'@,8n������b�D�R�[�t�k�oD
0�l3iͳZ(��'�� 9R�'�1O�3?FթZBR�g雁E�Z}�CmZg�d��2���?59�� �
�h4��:w��I3n/}�Ĺ�?a���?�����OT�qi�OV�Nt:)H���.(,�ˈy2�';�y�h��\1�^΢�E�՛�J��ቆ�HO��I<%[��ht�+�����Z�e����@���I�h�)� �՟�����8�����r5L�a��F!� ,L���k���)D�0�)�l�g�	�Y��M�톫"��5(�*yV=!N>�B̒Cv��>�O����lԍS���j_���'7�����,O<��=��F�N�uŶ�ʴ-�-aTC�W+jq�Kϲ^V�����������?I�'���c���>( J��$�[$K6dr�@�G����'��'�x�	�I��<���D�� �奇;T.�Hk�b��1��XQɓ�e~���ũ@A�3 m�/'� ���S�]���1�C�7캵SF��f��X��h��p��"u�N�HH�a�D#<a3�7� �����W�t�ʳ���z�D��Dg�O��DW릱��iy��'�����Q<�Y�'J4 @ׇ��8�)
��H�h��h+�'w��#]�,�&��_��H�y��;�,X0ņb�P�dTL}"[>�2��)�M����?)$+��.�n1���Lui��c��H��?i�P851���?i�.춵aS�i��'⢱�ק���ڤK#*Еm]J�zǓO��4B�� �P-|���O��X&
�%� \X���jʌ-'�'�Z������f)pӚ�DL�!zh�U���s$3��!>�ʓ�?����4�'+��ED�P�j�Ȳ�Yޮ��	�'Ԯ68i48�E B9���qs*�	520�o�[y"�]�{eNБ!�'ARS>!(&HF� z��� 6�
�F;�\����^㟰�	%I�)�,ؤO8����0t|૭���'I!f%�$|1���KJ���O��rRL�3B�A�2o
5v���B�(��Md��gdK6V�����<V�'����l#���'w����'>�z1�u��if�H�eت��'���'p��'&� @��ҽ�Vg=R��a�=O��FzR��%UН��&�3o�@���C�p�z6��OR���O�=��I�SJ��d�O�D�O��;|Ϟea�Z�1e�P	�� �l%�s�yrB�_�ʏ�D��<
J\R��	6&��g��.!�Zc���J�& �q��'*�Xj��ÎG�*�
�!�ͅ�:G��'��aZ�:�)�<1��7�;�)�,-@bJS��b
�'�U��.��}��Y ��2��p�O$�GzB�AZ?�*O�4ш�D6��"��Ҽ��J�ݢ9F��O����Od�$�պ����?)���̒B#(Ť%��B5)'*pC�'���<��+p�1PÌ�N
�0��R�~��A�4S�8{���g��uR/�E���b�=(�l�cڂ5ڊ,�Lɭj�,�$�O�	lџ0�'���D���|�tjW�L�n	ī'd��*�ODyХ/�z5���������6,4��^��j�l�Ky"�M�1�םퟬ�ɶ;V�2���>lg8��*T�n�����	������|�b&����z�*]^�Ԥ�4J�d����Rr �C�#*h�	��6\�����؁o�b$�F�����Q�I)	,4�P���]p�4���:O ���'���'��ҳj�Ё�A`DR�&�8��T5L��ß �?E���O�LM#s�_�G���-�xR/p������()��1�᪖�Fk�s<O,�R�Ցb�i��'��S:/W���	�@��� W8E��!_R�
T�I؟��wgިB:v=��)ML~*�@ʧ3tހ����PYb&k��(�bQ�O~����*V>�ŢA���r�"}�U��� �|LXC�$]���2g�Jl�Ĉ;H�"�'��'o�Dly�bI���Tԡ��o������O&��8B�$CG�U�}�h�j`ߦ�ax��&ғiq�Qp��Un(�%"3�F�-@�\�'V�}R,]	g�2,�WF]�/�ثMN�y�m�dL�f�� 8Ā	ǎ_�yBKBJ��%�3���[���3�C0�yb��}&��zO��|�d��R��y��Ғ^�(��"��� ����y �)>�I�5-Cy�qF�=�y2���]��uB�oW�Nf~������y�d�b��ҝK�r8��k�<�e��(A�ਇ�!� i2F^u�<IT��L��u�R'w���cǞu�<�@�N�ꕁ��H:���P�Yi�<��  B���9tA��J�~�<i��ڪg|�ӆ�����a�x�<�SA=w ���s�߁~��s k�<�udJ�Gt��1SA��P�$��r�M�<1!]�&����`J_	"`�-
��F�<iP�ӟh6��.���x���@�<�c��	��M����%0�(QI�o�F�<qKοyDUi�-آ-8�@���w�<��պA�H`�r!�a<]����r�<Y"��4V�} �L��8�*ݠF�X�<�"G 0{+�P�$%B�Z�������N�<)D=Q�\�Go�
{N  K��u�<�"�\�q$J�䔂^՜�Z�L�<Qp��=�^��d�N����W��M�<iGN�9=���(T�0L���I�<� N��E!A�6T��/Ir�y�"O�lÇ�D&�xi�Q�ǙX�T	�"O"}�����r�D$�J�'�x� 7-�j:9�'>�����O�Ϙ'*�@4�U�3<~��e�M�/L=Q��g�T��@ҊH�.�rբ�7��"��1'g$����zxs�&[ʠq.�6/m�t86�Ś#��G~R��0a�xk��Ñy����ן~ ��؆�H��L�h��
�"O�8�B瓔M�r ��cI�(1N�!1�O�m���_��E�q��Y�]G��%P%��f��ՎlI�*1�yb���"�`���G�x�<�kT��".�Hh�8`��S��u�-�媘�&�p�э���Lyp�:�㝑2 ƀ��v�azr�Ɍ� #��Q���dȥ��4���� ��u`�K1�V:�L�5}�RiKU�'�2]H&�_i"�	5n ��x���y�n��hỗ/҇`j�*Z�caɴ��?q�$�K%<؉P]�R�d�I�H�)�y2�6�� s�F�.�S2/V	2{ � í2�h2�.B e{r�b7�-vT�O�r�`�w��Lan�k����F�.�
�'�20�I[=l��hjw
��'D �X#!;��r��r/�{D��U�"�7IZ?h��b�����M�����ewV�#��0LO�UI@��?��税� hP�� � "Ϣt�փۖH�.��s�0j��!�$Z�*��l�דT����&hA��"F�ǡ|^���<aƆƣxV��i������`������عBԸ��u�Й��=JF/T)��ywA�U�<g�>�ژaӠl�H,�5xF`����+R���0��"zAo�~��O�����wFp���Ev�M����O�DY0
�'b��B�έn�`Xاj�6+�U�J�>h����� ��"Fh�D-D%/j�ϯj�px�=�qB�{D��ՂȈl��9z!kAO���*�dE4`���5���w��M�@O�k�\([R0�43Kє!�t�pǕ�eՀP��'��l��j� ^�f��42 (H�y��0:�I�x#��
䩙�ֺ�J'�����;�x4���{����Φ=�C�I��l��vy��eOB�D��S$�A?���R0 ��M�f9�#2�Z�8	����'b*����n����(�%ޜ�s���t���+9܌��AK�?���|皕h�q8���!��1;�`<���X�R4�Qc�8b���38o��*A15����'��{���3M�8��@�[nP1�%�G ��'�4�H�@b��7�F�~�Ad�Z	���D�>zm����F[���k���-D��2O���q ���:!�I�������ɩӮ���MоYW�tsm�~M
����K�(�͛u�]'qW�i�Ӭ��_S����E��9�qOz�i��E�#�:��`�X�B\J`�Ǧ��F�^;ƦӉ�p>arfԽl!��p�� w5ԈpOf�F���*��L��,2QO%�3������m�Nĳ{����ҡ 3>��2|Os`#�<�:M�FT�&o�X� ���J
�"�H�1�ax�Κ$ ŜUP�� �R��� "A�w�r���?$�h�k�m�&�$�G��� ��Q	(�6�b�D�d�P(J$�P.U����]��@�g�H�Oq:hiv�<)m�b->�뤭�= j5�1OD�'��qħ^6�xH��U\|���]Ct�E��')X����^�<���s��NE��yH�y2�D�NUPa��Ό0N�& �wJsN��P6Om�	��	;&���! `��kd:)������aF?F���®��MS6j�ߺ�O*C����Zc}ܰ��eB�w��,#t�9&p>�;�'��c ƵG
XA�AY�T�T���b���~b֕�X@�II�|��.q�|��ʒ�r�����H2uMVAS�y��h{e,��f+�(	�#� xAcЅO����!;Q�8� tY���"�  4lD\�@��x@aԍ_���'(�P�@D)I��PX��3��y��sB���R(E�D��	���'����,��:Q���v�ɐ^(ljSg��~M�9�M�/'�{"oK%,?�I��ݗQ�r��FOY<9r�U��+�@�|��9��'#`䔧��c�� DY�!�#��c���C(<�T���sR��p�aK�&��EЅ˚*2�#<QA^����-A3_"��a���0PuF�t� �ƍ�4�U���%�)��.$���t�Z,(h�-C3EQF� x�e*$ @�H��zt\ݲ��!}���}u蹸a��#���@��$��'dTX�]�h��u�*[�1F#�O���v%E�"�b�0B`��J+8���'_Bdi򘟼*Ճ��(8�Hr��W��D٘#BӋ�X���7�|���V�my@�f��/#Dq�"��-aj�ے��!F�Y�6�'���0��OqP�Z挍++TQښ�y��GeB��@V�ytt�ڷ�V�*�!��7�l=wl�j��pY�O�7Chh(5�Ǳ5O6X�Rf�Qt4�9����V��t�'m�q[�G�w�hi*�O�B$�O�u��1�C�T�U����I������P?'�h�d�'IH �ELh��E
穑���g[R�T��N柨QЭ�Ey�1�M<�=�Rd����v�ԻJv�]�6��U~"��3���DeZ	k܊�0��
��M#���=5��Z�n�eS�������G�ŚO����6�M!�zx�D��==�a|�J�e���#ŗ�
���r�.-�(R2�^�|�|��ϓ�y� U��Q 0�
�H1"����HQOT��Z�9a�4hcZl�Z��v��H��2�'�5jkJ5,Z��r��`!�Rb^8^#2��[��Г��2U(f�Er�ؘ
�n��H_:bJT��1�����c$ұ7|z��邟h�(rT��	}���X��E��M��jN�]�#���Dy2m3<�p!fiB�����õ�����tr���t��4�2�� ���}���K�i�J�&�VX�$3oo���i�&*$m���:<8���r�@��b	�shJ�G��`�SFq�O�����>H����D�z⚯o�8�����������t�.}���V�yv=�=��F�^�v<�0OlPK���7K����8�% �E3���Pk��WZҠ�%��U�'D���NS�=�^hK��x��$=6��e���;"~Ͳ��W�]˲�a'�Mv?�`��?���|�<�Q���h��)�Dٳ\ff�tn�L���'9�d�l�3}��3�vU+�K�no��	F�D�D�Z�@�dG�?$����M~���]�BVz�f< \���R��69��7�:���<��H��v�� ���Tw?�ӥ`�u@ᢕ,1[hё���M2�$3��,Od���H��ܸ'�ȅ��!z98�C�MP<�ez�)H�H�����tX��g)���?ex�w�2%!'g�X���s�P;4x�J�O�L��������T�ߩJ��&䇡Hr���у|?ϐa�E����u��Q��Z�;yx�ܪ1n׉��@��a;�ɩWF�A���|2f�|�rcY�[�t����Cj��ap��f���DǏ�x�;�N=lO�N˰gf����e
�����$솃��yJ>� 䖣B'�d�I;hۦ�)u"�Ο�'o4����(X'E�����E��R J3�	697�^h7�� �(���o��%rV��흋P�.��gU�yz�Y&oE,\޸
�ү>�V��S��y�h�5~��Qcs�>+
���j ^vXᓄ6�n�㷪�;)(F ���e�D3y�,0b�ݳcMp���#
�?����"c�<9���<��ם�SMў�9���&��01���<)��y�@�q�{�虼�?i6f3���Ӽ#BG�.qK�u�ӎ˿)��$㊜b�D��,J��hO���gZy��� c=��Ѹ� �C��,�ݖN�����'F1x��ڲ�l�O�1`��#��*H*6�n	d"V��J�cE�U2�؀У	Rh�r ؁ҧB� �b+4�D^dc��J~��}$pB��_\��0��"��$�+IB&]s�r��"�T?	��� l�UZ 9O�չ"L�IB��5l��`�H�kB�p�  DzhQ��f�"r�O�-�ED��Q;�b\�r�8�(Ѓ��e��?Y��jL�28�*ԋ�B����s& hT���e� Dvr<�5��	=o��T�I���yc��!Q��Z�`P<�B�)E�?8��(���e�"=��8�Ȅ�W�.?��nѰU{�M�UDޝ~�̍pbϓ�2�'����ۦ�9�iʂ!+����$'h��kנ�*c*��#)�	�j�*��+��1jMp��Y�6ZA궦#?A�i\�DT0ūҀ���4F�k~�V�qODUrA�âF����0N�4�z���V�!r��Q#*���iX����ja�G�4��c�8{���?˟����C[}�< qd�R�#O&�p��|b�B�c�&�r�+����Dӣ�2��'�Ƥ�!
D��Fx��֗/x��� e\
��'��>�I�՘Ł��E� d� ۥb���xT�I<Z\u
D���qO�Ӑq�2qϻ���$+w쉷M
�F�h�����O���{��}��6b>(4��E�YfH�ӌ��y�1OH�ׄ��9�a!�R��t8����\oA,}��jӕ2�^(��΅�Q��y�bõrS^)��ƕ�u���,G� ��EpjU�gLؽ#/�$U�rU��O$'!V�{�b��IP���?���`	�x�D�$,h4Li'Kݡ^<��螧T�I��FӴ62����$ˍEQ �p��F�7��t�al�+���Z�DWAj��>�Ą���&�u�'bJĊG�N9-�\����0xj�#�T�8���&�U)/�.��=�O��� P?��YK���-6�䋃M��O�^�"a���d���`w�L�xXy���Rf���O��PS�k�*\_Ȳ� G#(����/�I-c�����u8f���M�+�rc�<�E��l@&�pB���q�z4 b`ΓQ��l�<ӣW#`����9#P�;��F�`��(��Oߒĭ�9���+R�n�
�A�"*z�,K 薼S~�xR#��>dV�Y�GQ�}��(���0d(���5����/�)�'(rpd 'jV*�=i��Ζ&�:e�㉊��e��zۚ��	�O�8�(�Ν���Y/;�ڙ;qI^����e�̉]����{*�j�1s�b�����]4��p�@��F�\pȷ�!}�=x���gQ#�޹E��F6�l�ÅD�*=�މB��zi1OވF��:��aa��V�t��w�ĜN� J3,C�Pɦ��	F�y���� ��tC�$�'���A(��dJ"ɔx,�h��bX��E([
R*���gy&�B.��z�Z���(U�"��ys��'��` o:_�1�I�)���GS2Bx��a���1S�@�Ƃ��4$!����y2AK�v�V�9$��+E]X3W i�铗�' F�{���+�X1S
6�y�ρ�`IV�+C�����97)�UV�$e��6��H�'g��]*i$,�ƅ��1*�kW:g�d�DàjT�A���F:v�qRGF�?-�&��'j�$�3u"���tt "��|$���#����%EW'��	'�?� ���J��� 䲀O�H]�͸v!�p*QOp$L��Mʬ+��I��A��� O�T�S+r2"���	G,	���sF�ޝ!���I�=pŐ� X'$�S�?Kd�)žith�R7�+!q�9Qt�8)F}"G�5CN�/�3E��郗j���Ϙ'αؑJC�;J�1U�ì' ưX�O�Aa$�Ƨ�@�c5��;3BI�=Y���]qΡC��l]&%�,�v���Z���@��mBH"qF}R��yg%�B$���kX�6���&)	ֲ�"4AC;��c�l�T���!��-�'D�$�-{b���dS��|�y����#>�aG�Au�m�j#�S�u�������Ov�p ��ϔ�'��H"��(+�f����|�uH�~]�"R��<���<���5>�"d{��3}��I�<>c��c��)YH�k#ɉ\��ϡvn�{����	Ь����-��鉠!�4��g�L��IS��<)��
r����b�#۬e*B"�b�������Ğ�,��٢�	�4{��CvW!�D<M����p �+x��T��F!�$I8|ڄ�[=&�|`:�%R9K=!�d^�%M@lkW�A&L�y@1CL�E�!�č�3�֕�K[�0�+�G� %%!�H�F-hD���y�8bU�B5);!�dI/lX��X��ıyjt xI �!�D͊њ�ҧ%�sc���! �!��
 �Iz�MN����i���MY!�0sY �ф� �z�@�b�ƞd7!��d��X�(�!U%���R�Bg�!���0����� �.\""�ԁr��C䉠>���3%�W�F���e�?VFC��(_ƹҧ���v�t�#Q�˧��B�ɯH�zY�'�ץFVJ�b֝��B�I2jݦ5!pJ	%&I�H��һ��B�@�NVR�@ L0㣞$��=��'u��M�;P�'fG;�H�'r�k���|�1	�Z�2�yr����$y4L��afe���>�y�ϚWS��7#& �:��1�yo�$:�R|�Z-!� ����yN?i�<��(\�D�nH�f(X�y�'�2��i{`"�9�� �T��yB�͜e�,Y#Ç�$�pq�b��yb(�Q4�Ԉ^��Xly1���y2)�(K�fG���D��s-�y��
�]y\e��!��h��T=�y�`�*j7����l�j��e��y ���Ȩ����^�dA���y���0P4uC#�� VIЃ�D5�yB^�N�F���@�p���iC��y�$��O�L��E�Μc�y�s	�yүD�dļ!�dj��X���S��L�y��=�����|��$�B 	��y�dN/f摸e��:{�q�򭑭�y2DT�,�R蛺)'��� L��y��YR�*�H�"�v8���4�yr��	�F���K�o� Us�̖�y���U�h��O��|�\��R@���y��	�&v����\�r4����Z=�y2I��o(杀��"m�ƙH�چ�y��
�`��q��bܘQ8��	�y�Q��1"O��H�%�����y2(L�X|��JBC9N�����mė�yR"���V���_[��$̎�ybO�eޔ�5j�&(sR���S��y2�Y�R��:BM� �d�Kt���yba�V� �"p�ˬGҰ�j��J��y"�M2B� ��@��iA�H����/�y��Ɉ0����3���54`Q��P#�y�%*��t��Y$��)��͈�y
� D���B�Kz����p�T;r"O�Z&�0-���P鞗o�,��"O }���}��� ��Q����W"O�\�q��(D�����w��E"Oʠ�䯗�� �#7!DV���"O�Y�s�W�Nfh�����>*&"O%����q{��S���$D8h�6"O�ա�����e ʕ8#B`R�"O`���#2)�}k�,v��cA"O$q��*li2�K'lh�\����y�n�2f����%@m�9@�П�y"��d�����$�pTcB ���y�@V�.$xh�Y�s�J����yRH�;��e0!�;3�}C����y�J�'
	Н�!G�@r���D��y��o�ڳ��"1��1��(���y��=qL�c0�_%�>��@$��yr�Ɣ�^�hdȜ#����e�&�y"�/+X,io�p�t��H@��yҫF�9�q�Ҿ~u���	�!�yR�H�g$�C��R�w���dg��y#�?�|L�V���&!9
����yR��	i�tS���6zB���Ǖ��yB` /ZS��)%�ě1�1���4�y��9KIҥ�'��<$5ڽ�����y�� �Ʊ���Ѿs��bDE��yBe֯*0�%Y��\(�u!���y	�*[�֡�D��#N6��9b� �~b�)ڧtZ�`�E�"�Iҵ)��~�P��=9������A�NDf��3M�3�+!%����R�t�8}i���|.=��Ɩ-!�d��� ӃǍSQZ��A�@8!�QPd��P`��S�PKR#n!�D�;B,�LǪG� ���U�!��=��Ȁ�[(������q�!��-�ASbə4������;�!�D�~����u)(�ڤ��a��!�DR�d�̌ "��x��#�b��!��.�N�RH�R�����L��!�$v�i��MH�;�@ȑ�O�	m�!��3d
.��߽|��H�CC�B�!�D�8a����׬�Ш:em�,F�!�D�C#���e ˶c�p 6�[�Z�!�$+f�����3|�G�8
��*�S�OZ|�1��t>��n�D#Fy�
�'�m�T�9S�<��敕D��̳
�'�N h����{-2E���8*c
�'*�`cM��G�zd�G��2&��S
�'݀�c��)D	�	@�2ŀ���$+�r��(�x�9��E�(,(AQ""O:I�3��0�F\��₈{��F"O�˰���c�4��p�v�
 "O�����L|
��1�8X�P�"O�����2A����M;���Ж�M����ú>]�0�U'@�lN���$D���'GR�݂���R�t����'�d3�Sܧl���M�P�,�bΕ�|�XL�ȓah8{�H
k���S"L�����ȓt����p�ƥ��I�D솴e����<�* {�팈��x1�@������X��0iT+�R�:Ԯ�0( .q��	�I֨#<I���]��I6�űM��В5��_�<)�bص#@x�HS/YIx���	UyB<w���Ӟ|��)�Xo|�9�BR5F��Icҩ.I�!�� �� S�[%:͊�2�iĢ1�
�zF�d�z���C�G� Q�N�����D��UG�+D��)�(��ؽ��Y�mz� G�.D�P87��&��M��-�0m�k"c.D��HU�N+b�D�	�Ɨi ढ1m0D�,A�с;~�j6�%4w��f*OZ�i��R鄘sc�0/���t"O�)z���Q#�t�&��&�q��"OTLɆ'7B`~	砗(WiAu"O�yI炙ȩ5b�w$iAG"O��x�h��C�K��A�$*�"OR�R���-&��ka!�!�R���"O�m;j_9�܄����-?�<ĒB"O��g�$
�f���F�-x� ���"OV�c�jD�y���s"����@&"O�DC�l^�/R,!�%"۱8��Qr�"OL���~�T�aR��1,�����'#!��%J�ҹ)U,Y &�hi��	�!��	�AT��l�3	�n����v�!�D��0H(�S�G?,��ۑ��Nz!�77h��ǬR�N�~:�B(�!���$&��+��yY�a�Y�s!��^%X� ��S5x�`p����V!��*A�R���Rp$�x�C8)F!���1#
���`y���(��ךW�dB�I/Q�~���fՈ�¸ʶK�(�NB��0w��$ N��h���ϐ|����hO�>)0Sd_8e>2a
ɺw��Xe@.�O����5�M;y?��h�A�7m��ȓ=��9�?|�2���ȓ|�p)R�f�(\����M���JX�hC:�����ǁQe���x���hp�����k�M�1��Ia̓=9P@��6|�t`ۡL�)z܆�V3R�fж�*@���ӄ	�����ܛ�S�a� �z�J�Mn̔�ȓgV��	�-!��vAۊ���Ol�=�������`�B�5(v#�]�<Y&P�v���	aę=1�Vū��]�<�%$ɫ�də�K���rY{#���<�*���L]�u�ڿTtNȋuIU@�'��?��yz}3G��OފU[�>D��"SD�h'~e)�.^*4�hU��C���F{���_=s��QCu�U:"8��S�[�lN!�$���֐p
H�k��xc�Ӑ$!�$N��=
��@$p1ˤ��z��	h��H����-
��y��n7�!�v"O��rPi�xr,I�l( $�"O�X#2��<����	.0�#"OHM�fՠD� +�B �=�L��"O�6�N�&��;��Y>Ӑ�"O܅i %	{~�C5l�JWPC"OPʗ/Ɯ3'*����M�sT�Љ�"On!c�`��pHx����ZS(�b`"O�#%���d/��m4LJ�H!�"O�MҡI^?���0F���N8�&"O��{4C�h�8��=��"O@,��-��N-�DIH�X���S�"O��b �Ԋ  �T�a�ƹb���N�<I��_,��x���R24���b��K�<1�}hB�#���9/R�Җ�_P�<@��>���@��;I����kQ�<����#�����X�3� �O�<��ʛ�Z�����Ψ��Pw�d�<� m��j�:a>&	ۓ�c!ƍ�"Odth�/3�P��A+܁3
�ػS"O�̒2̅�Jr�Ջ�»2�B��"O&H�A�9%�B��
	w -��"O�HFȏ	 ��8&�Z��A`�	F���i��1� DҲ�!�����	 ]�!�dǋn�Ҁc���8A�~b4a��"O`���+@6�u�cD�ߒ�K��y����^��S@E(!*���'���yb�]�"�d�'+��r�y�Wo��yb�GP��DcQ�4���b�-�y��\e�ᙦ'ŗ~=0�I"���y�΂�z[��Ҁ�$qU �k!E���yB���.�Y��탻j�:]Y���y2č ����rW	�<�A���y�F�\��<xw�ðG!���B��y�R�إS&��Ȑ�A���yr'= :���I[;|�b��yB W0R� Kb.M�)��!�GH�y�JIDz14A��~T�ȃ�y�H�6��}
g)Y)�s�F���yb�Nb�|b@v8`���ylFL��H�V�6��`'�,�y�W��*d(s  [��AW(�y���&���"j���zqB��̞�yr"�
SG`��#��f�8TLI`�<1�oqP��`��ˁR�f�iv	�M�<�``��3}@��f��@��R��M_�<aB�ya7�s`�i"CH�AJ���2��t��;|�[�mޅ>ȓ_��<�3$�5$�p�YL��~��T�ȓ�4d8��T��Ixģӽ��m��\���J��''�r ���:@�hD��JB�$̭ k�4�(ŵzhZ �ȓD��x��b��[�
dC��ȓc���H�p/ZQ�ABY ά�ȓf�,`[�@�6WU& �6͹-|�!�ȓJ���q硆"&δu:&d��V�Đ��F a�Cc�,A�6�`�Δ�$5<�ȓ?�V���n�1�$	�	����C��A9���h�VY���S�+�̤�ȓ'��m(�Nަc�&���A�[�L�����ـ6D*hsj�27�DTK�AZb�<I����6a5�[2��]�,�v�<�U-Ørb�����Y�8 !	�^�<����M!������+S�U�%Z�<i�e3$��ts�A[)��4�HZX�<q�a��J�*p�c��%��:eόi�<Y�ˇ:p�aB�L�!Є���M�j�<��hX��n�*�E�a�ޜ*lD|�<� %�f$jj��__��{��\�<�!�.~ap�k��Vp��j�Y�<1$fU�^I�e���Y�p�v��'DM�<م�O�z��ǀ7n�����E�<P���(ǆi�&��4��1�� �C�<qԥ|����̖!fw���$Rv�<�A��2�x��h�c�����X�<�`��(���P�E1XB�)��c�X�<�i�7�<��a‸{HдeWT�<�E�1�}2��_����V�O�<a�lGt�X�ŕ	+�XT�@/�G�<IaǲT�ȸ���C:ӂ
���E�<��I�OO����%AzX��P~�<��C�ۂ�(�%��#��mIT�{�<� .� �+���he��WKS�X+'"Ox1��KIn ���!*�',B�!qS"O��*�+��g�X��G6++�-b�"O0��⊌$�=�d���iA"Ol[��?VXb���&�$66��2"O�A�mQ�]�)M�m��B �>�!�d=>Z�qN�2~��py�Z?}\!�D�#�`��Rl��B�����C+\P!�d�.qZ0��HE�[�@pj�V�?6!��J�?����&��%�Xy$�L�.*!�$W�∹3A(+��9��ܦ !�$Q
A|��p��&!���c�Ǆ!��֚Q;E.�B����!Y#!�D��K�Ɗ@���@,Y!���0d��ؐ��R�4��xH��U"�!�Ӕߢ�ƅ�Rt�r@E�.-w!�䆹W�@4��e�zM
Up*�`l!�$�~9�������b/\i�j[$yh!��ѹW��X�D. @#�i2iQ#K!�d�@*M�&�P>-��Q�NW 
1!�$��V�X�k�o�<b����ؙ'!�Dϭ����k�$�t�v�	!�d��6�Ѐ I�f��<�iV�%*!�Ċ�S�4YҡŀM�Duا(��R�!��[�8Y�ɖC��i��@0g薵&M!���VONA��8t��P�u爡qC!�$Z1,���@kmb���+5!�Dܗ[�|Uh��#O���/xO!��F�Q�rD�ud˵e� ��ƦFD!��]y")Q�-
�%|h(H�ʈ�3=!�\�Y��h�턮;g>U�Dǐ�!򤚼0x����j]#+�\!�ǙMe!�V�bz�uˀ�¬}8���Gғf5!�DV�\�@lS���"��E$��"�!�D[m��p��ίJ��IjD,R#4�!�D�J{r��LYP��}Q���!��T>)���:����X5!�d��VNQ��K�' $	"j��z�!��K5F`0!m'f�8�wBM'!��A�t`Y��;b`jq�۶�!�D�j��!�'�N�(����!�8Gh̙�l]�p�ʙ1��œ1�!��>AS�8`�:h�blxu�9	�!�$���H��]>'�С҅��!�bݎ��&��(c��E�n!��/^�Y��!��;$+h�!��L���� �	�88	����,�!�D��/H�,�-8zp��JD�o�!�䈕��0�$�B�%��X�S<u�!�ǞIQ�M�����'aD�Pn,|�!��X���f�ݟ+X�چ�џM�!��1�)����BK J�F�c�"OD}+�4$BHCq!�8�h��1"Ol�9f@ϲ��ԩ�@ r��A"O
��'�8|�H����J�h�"OȄ/��80�E�Zv��o0�!��	�(��9"�ӭ$0*�$��O�!�Q�Lxt��fG�s�|"CMY a�!��|{�s�@E�a�vI����p�!򤋞
Ș� Ö(2��t�7�^	�!�[�j�h���	o,V�� ��,:!�dD-� ��J�	 q���r�!���:+TTK�O�Y�`ɰ�M�S�!���|5LHdO�#�&$Y���!�� ����q�ظV	Z�N����t"O��*�&�	7V�T�EW�i "O�=X��� '��E�ӊ�O�Șt"Oօ�U��lf�)5�X9z�d�u"O�h�*��'v��[L�L��Ȁ�"O���c�M� `^@�sDɉm j	iV"O~\)�(M�<a�r�b�`���"OXc�w:�$�c����y�"O,d��`V?1!�	�BP�[T2	%"O�h�dY�dhʡ�� ǹ=���	�'I�%q'E�,���� @A�',h�Q�l�h�"u!�yx�"�'�d�¥ꉴE2iP��`��
�'���bC��$ h:`%���	�'��h�@t�-���V�h��'� �� �_�h!uŖ:#����'i$�P&:����Q9�<��
�'�T����.�PC�!a���
�'g�|����|Xp\�C�Y�J(֠�'A{Ã/mj�Q6�<�� �'ڗ��q��� 8%,R
�'�]`e�]";E\��B9-�"�	�'�$Ԑ!�W���h�--j�,��'x���w�I�XfȁY�+��T�r�'ٺ]�2�]�[f��a �7V �"�'��SȖ�G��t!�POA "�'�da�B��(��Qg�"D���
�'rbx�q�	`ܦ���<���
�'������#�)��)�.1��'
�4��	F1�p8sFG&�K�'��TH��Ư7���s
U<�Z��'�ν!��tt���mY .�L���'54`mX+�����6r�> ��'\��Q��,30L��%ߊl� q�'��!�D�F�Ja�H��W�/5Li��'�l��Y86$<3�D�-/^��	�'�2YK���|���f�s�&H��'#l�$%Ό,�8`FLÇ6ZE��'�>����W�Q������,yJ� ����Op��0§�
�ۣDZ:<|��
Г6�T�'�2�'P���O|�J%�u����"j������.28HC䉺E�R�͗]7�(�GeD�BC�I==Bpiu��	���Q/�	,�(C�	�9&�z�@ӊ͌ �F-��}"C�ɜ=ٺ=bq�Nt��OǴ)��B䉮a��h9R-��R����'��l��?A��iO�B`�c�b]<���"I$E�S�h&��gܓe�F�PT,�P��X���	9�ȓd�m��
�GƠ���5�Ň�8��%�g��#ae� F.�&kyR0�ȓE�>��JU$8���M�O�xT�ȓ�=�fÓ >̱2��rWb��ȓV���8E��G���Y��jJ���T�����؞�i�@\<"EL��?�ӓ^^��5��5�
-q��ȓ\� Ȑq@� x	p���>���ȓ`:���Ț '�\� BJ/M,��bu�pv�Q�3�h��4G�)��(�ȓ���RE�Y�8<3�l�4����>�l���H7�DQ+c-��PӤ��FL���"�Ё�Z���<�'����Э�0@�0h)���)`�C�ɮZ\"�[���7�b�1��[x TC�	�	!	��d�>�)Q�k�tC�)� dX���ȹV$A�q�ʶ�̲�"O�|���YT= ������ʵ"O�`��G�_��)�C�/����f"O2}��j�uN��d��={�4�C"OT�[���`
�[�Ⰼ�Q�^J�<�!�]mAP���WrNS�TE�<��oՕ;
v}(�/�e4�]����|�<�w�.{��L�%��<H���s�d�p�<Y�e�\��9�d��?lV|k���m�<�A��k�z�CF����n,#e �O���,��@>y��%F4?J�=�"��Y�h�"E1D��*穕/L���k1�[13���P5D��P[���0,�4[U�HQa�0z�,C��/n�@X�\�{̼��C�.O�B�I&���(��t]�M!�,5�B䉃|R,�pn��!�Y����ra�C��	9�����O� #�œŮڙ'^⟬�	D>e�`�z��D�Dم=m�\ۀ.1D�4³�R���E�w�ظ�ĲRD$D��I�J��(򖨪��*2D PQl!D�$�u�� eU�2\���
���y"�2v^�Ԡ$��O~5+�J��yR���%v��X�H?2��HEj�2�y�GG�6��qCNY��q�gDP���hOq�lI�!D� U|� ��e���C�"O�dpQ
@p:�X���G+P�-"3"O$"�+�\
DF�0���X�"O�UB��X�R��ɂ�D��]��<��"Ol) �l�)f����������X�"Of�c�J�1'¬�T�Z	
�~� c"OR�����бo�Ќ��Y�xD{��N�R����Bo�L���9��]�!��>Q����Մ��fy섂�KڂZ!��S���:ce�qL�A�j��!�$� V��ѐ�Ί#$:"�7��7!�$�1d��VC��<�����U�Q!� k��``N���
y��־�!�D�g�.Ӏ+�)"�`��A�P+�2�)�'E]0����@�j�,�#�%Q����'2��⥝�'��ccOW+6!X���'U�K7�0=B�$C9����'�TMec�X��9� �95�v�!�'TV ��e�0b���۳d�+.�����'�r,a�"Jb@H�83	Y�z���'|��.@�T��D�c8n��'���+s���W����U�9#&�
�'�z�IQ�Y�r���3���7�zi�'/��W!U�v�PLE꜁k�� A�'`L�HA���>d���#{F�l��'�	2e�g�5�H4��GaU��y̋&/���hH�Bj�Y�����yr��6N�F I��Ǩ?�I�G��?���'J��i�^}�� 5Z���t!\k�<A�D< O�-#Rjͫue^��7D�c�<9�����n�*�o�L���&g�G�<Y3��2[�8�	�5P}NdZ�A�<��B�q��tG(c{"xB  {�<���A���	�,�����%�x�<Q�  �-�$������r�(��q�<����bl�xp���9��4��E�n�<3�Ͽ�J�2��-C�����j�<qe����!׭5jK�bK	f�<�"��;4j���¸iJ��V��V�<�䪙x�Hu��1��ݺ�.T\�<� ��" FP�9�Ty�5l��w�b@ Q"O&��$�� �YzKF�(��)y�"O�|��Oլ��Lq������Q"O�$22�ݭn����� г/D��J"O@಄�>�<pzr��?"��t"!"O.��P�̅#
����ŋ:�R�a�"On�k1c�0hOh�rg�<(��(1"O�� ��V`��&�\��"O���dl0%ۗNu6�iY!"O��h�0o�,+��ӏ ���"O��"�L�#h"��K̠X��YV"O�5c�PE��H{j^/Y�Hc�"O�pxl[u�dhPF�Q�*Ժ�"O|,R���o�4���G�����"O�u�D��-�@-	UB;8h��A"O�`Z�aEK
��D���3�
r���O���2���"!o��5v�1���ص�N���%��i88����N\��m��P��Ș��53\
�����X��!��y�t�D�֛	�B�R��*)q�-��:j8��ƀ�<d�d
�.'zj�l��'���Q�K�2M����j3r��JP�!��h��D�93�oO�d��0�?�-O#~��XK����	t������H�<Ib��Eh�Q����B$4���j�<�צ�y©��͇�l�jۤ�EQ�<�ȃ1B���u*�1��ݪqL�X�<9� \$Ei0�y8�z���V�<�T'W�>
ʵ���B/lI9QGJ~�<�C�U
����A�M�z��$�TO���?���ň�b��cO	�T�A�'KE;�&��"O�i�D��
.������[�]��Ma�"O�$ѵ�̥d����H�A����"O�-���Ȁs�J�s2�89j�"O�!ff��.���EC
Eiy��"OΌ�U#I�_���C�֒C3teA�"OV�J�"�"%��<[Ċз	-�`f"OR8T�6Ÿ�Z ��2�P� "O�Ak��K�|A�D���R�D@!�"Oܜ���܉���Cd�$�g"O�H����(u�\�s�E�vn	��"O��ë]����b��N��Ʌ"O�%-R)%=H%���@Y���;�"O�9�qN)q�9Pˋ'0l�aA"O� �%�2�-Ѕ�];�N�U�|R�'�az"'�,ph�V�����p����yҤ�$/VP�Q��&�|+����y�-�I�d[�E({�YY'�;�yR�J�{������ku6]oJ��y�g�JN���s!ɏ]n��S�	ŵ�y���25V�1�B� \NZeb�-�y�AX�4tZ\p%��#D�ROF�䓥0>	D�7���Qև�c�x|�uJ{�<W!�{j�)v��	o`���'Xs�<��'?i�!�4+�-	P�@ K
{�<Q'�v	��(S�|w�(H�u�<�se��D��p� [������J�<i���:̜D�A@Rlơ��A�<Q C�kG��P�gV=Byv��`�	~�<�4IהX���Ygė6k�B=c��{�<iH��	&����C�6F)�y���t�<���I�X��h��m�R�ҐH!+ Z�<qA�+K��X�Nź��a((�q�<a�Yƒ�w�
�bڌ��Uw�<� ���	\y���z��g�2%��"O0"�d�n	���GMkJ��v"O0Aڂ(f�ɲ��>DёR"OF�DE�6u&hS��R�Ftb)yw"O��c�/Q� ���k,L-
�q�c"O�H���!���Q�/�����"O��X��
�>�*M1ʃ)��S�"O��8 �0/T�J��E7t�Hp7P�,��ɴ]�J�Ƈ4�l�сF!��C�ɉYU��{����pe	c��C�I�O���XbH"AX�W�.6^zC���,��� ڼu9�����̄.��B�I�6��qq`��#d�9`l�,_��B�ɂd���c���OT�����"Y)����g�(*�����ćU�%�h��8D�,ʄm�-�:���KR�2�` ��5D������2S#2l)u+R/]���hp�&D�\���{<q�&!\�?3����$D���hG<얥&�@Y��$D���  �w(��#,V��(6 !D����M��e�`�q@�, ���
?D����?k�l�!6I�-�ހ�/D����)<(Ķ ;�KH�}�l���.D�X&�ٔP����c�)
�����-D�<;a�2բ|�oF�R|xz��*D���U���	yn�H (EBh��b@,D����Q�U$���- �A=�}Jm4D�<Ah�4i�~,��X�Z-���&�O��d�i�B�L��@����R&�	�ȓA��0��N_8]X0�;�C�,��ԄȓNDzz��C58q$�;p�~U��+�Z(є�?$��(��7hm*U�ȓit䉻v���Qx�����X5���ȓ
�]��,B�+��3E��2cؐ�ȓ:RƸ�4o�l�Y��g�� �����I����I�<�6���p��(hf��We�B��I�<��L�$����g���W��l"�E]�<1U�ڔ~c�݁�n�&R��Ѣ.�\�<)�a�V�&0�Ԉ�1o)�I9��m�<�EgK2p/�����2A��!��u�<!�CWd��L��'�08����&�q�<��Z���pht�N$j�b�B	�Ex���'��Pő�:X����gO.Z�^ #�'{Z���ǉ��(������W<$��'X�y�tCD��\Rd�I�b��'���蟶9��T)�([�x���'Le�e�RD�PX�cC�Ԩ�'2�����t�U�GJ��R���'4D I�A�a*�X�%�$E�Ɲ��L�H���KP��z��W!d��݇ȓ�xq�s��ee�ݐW HqX$��:�X�2�#�~$�V���{b�Є��.� �,���S �	�t@��U����h�Ly�mS�h�`�ȓb�EJ�&�U<��=��ȓ	C�=
��I�v�*'�@�����ȓ�Tإ��u�TM�@�d& |�����c��	k����W��z���$��,a�R�n�"m�v��H����Z&�;'W�d��ʔN&M�JЕ'�a~�Iϛw����O?`ϖi�c昚�y�g�3e,à\�OjL��3d�?�yr�Y��lk�A:���q�@��y�-\'A& ��b��2�b\y��E	��d�Oj⟢|� Ɓ��d/y�@�RԤ�-�,*�"ONR@��,4�3��CY{�	�""O��cT!>�arD��Ef��"O� �� ��%���`,�o�����"O����@1NڒD�kg�`�X"O�x���+)V��L.`�\�R�"O���S��2))�	�> � x��D>ړ��D�3xX��ڄt���yA F�Y4!�>桠�
�W��p��ˎf!�d�^n�k�&�?U�j�Т� �.���'�a~��J)C��أ&�� E<�+V؁�yBc�%f�ډ���K�S?40q��ݷ�y�չ&�
<`T���PӞ1걉��yb(@�1���`)]�EL �с�A��hO*��I��~�5	��	������!�d�
8�K0�D�cLa�v���!��8d��L`r��.�^9�p&��!�D��L��֪M�v�.T�4��+]~!�M�!���RQ�Eln���eC�/�!��D��8"�i̝Wax�@�ݸ
n!��[�_�	i��K�riq�8 �Ox�=���
5���v�d�mX�@�VxA "O���2�������b'.�ȷ"O`U{��OB�E�F\��R"Od��¢�8�U�-Q���ʇ"O�-�Հ�%
��d���VF���"OYZw�Ƚ&��#�f�*T��I�"OD�����L�qY���_�D�#"O�s��Q�<��l�7P3`Ⱝ��"Od�q�O1.2-�W�-OB>��G"O�}�g �)����_%z�c�"O愻$i*aP�¡N�!rb��"O"���F��>Jb�rB>8S�la�"Ox�ke���U��p�a��w�8�"O�q�<#VV*�O���y�"ObX�G�E�2x���Ņ-�`a�a"O�V����������o�` �"O�XfNԸa�X5 ��.��Ы�"O���+~,����n�1a����"O�IQ��>K~d�Rc�L��Tz"OX �@�0 H���ޜU�r�C�"O"�xw�C�-˶���6�4%��"O�(S��AD2Re�ٽd��0�"O��A"]�h�� 9��)FBE�"O�!�nS�9	��B���8�my�"O���+�zh�#�oTA H)k&"O�S3���=��������C
2��"Oƭr2�٬'/h�p%�#e�� ��"Op4�@/�-[���A��%Ҝ�
�"O�S�R���a��D�1"OгũW� ��|:��σD��h��"O��Yd�����w��0�.��"Ot�;�Ǉ�1�
̀���?Y����B"O���FA)栰PL�Ny��&"O숑d�!w$��q`X�5[$���"O���U(۹l7�0&m�}<�Ix�"O��rf��,�OKֱ�r"O��p���Lq�3���f5�tXV"O��rc�l۲	r �C�Y2lQ8�"O*�[�o�s YKi�0"2mJ"O\�ȴ�
��@��f��>�#7"O�Z���+e&"I���
����v"O$���n�<1Q�1Q��Xjt"O�*�g��t�f	;�#�<w@@�d"O� Q��g�V�� ��A_�qY�"OF,��Aڲx����g�*+"�x�"O��9惞:��P1��@��^��"O>03f+�*m`B}��Ř��D7� D����W/����H�"?l�I�m"D�4cU��8H5�C�XÚk-D���2녫b.���@N�;W���ɴ�*D�P��E��y;D.�9rFIե(D�����ptj��]��%ʜ�#!�dԺk~ )�@�·dFN�HQAQ=}�!�I����A��92J0ء@I�-�!�d�o���W�ǿo� ʗJ��!�$D2J�*)F����R��!�K�4�f����W�=�f�r�	�!�D	�F)���	�w���8�LD/n�!򄜶�n-�W�G�G��D`r�˱�!��Ly@.���JX'Wm�(�Q�[l!��"�R�dؠQ\��;b�]�!��@j��@�L^!ONH��5�Y�[{!�(	���%4���� {�!�M�F�xQBCމu�n1��x]!�ĔJ��h�#:���#�V'Z1!�dM�kҌ��.L3_��-`�&�#!��?�P��D�c���Q�E &!�1��+Zo�n�бNR�!��>�:1P��Ύ&R��Q�l�-�!�D�(���4��'.�m�Pl��X�!��s�p�D��L)80�Ʀ�!򤛲U*.�"�.u��x���=MX�C�I1.$�أt�@	aw�5cBØ�_��C�Ii|�=j��Ԍ<�!�'"�?�C�I�E����u�x���߲V��C�I�u �yQa&�|�F�����1U�B䉫!_���.qL��Ǉ�dxrB䉊H�
t�E��<e:حkV@�>�lB䉌O�.�
��XS~ĽK���oJ�C�	5rȍx7 P��^]sc�˷Nr�C�-c2J��I�B�2�Y� �&^�tC�I�='b������N�X�Z����q�RC䉙\���&	N�$J]ʑ� &2fC�I}*B1�#�D��x��BU�JjB��
zT��%��[�P��"O�RN�2?��$�%�7mD���"O��s�jֆt�Y�'�E�j��b"O� +�
���`��@
�&hXM:�"Ob�0aL�-���ToT�R*t��"O�A�Ҋy$�`QTI�~b\�w"O2i#���B���(�G�>B�]R�"OJ��_�2�p 4FK�uX���"O�!�P�ZR�=q��R��y�g"O�9��	�t�����!z�l�؆"O�|�s�]�|V�G:N�
��"O�p`�IY�}R鐧�A���$"O��0J�:o��a�GVi���2"O� ��jS�+Č������`��As"O@�Ґ$B7b)�5�0���'���*2�'�'�B��>!a�X�<(�0�Y�1~<2E
�x�<�SF��j��Q��2���#�u�<��	&yx@��(Գ+O����V�<yf
��|�,�EN�/�@!�mSO�<��!K:v��erC���[�x��E��D�<��J�y��R�٩-�\���
@�<�J*wr=P!J�;�v)��~�<Qs�Xf�}�Ɂ;U+<񨇅�y�<� ��+Tc
������m �=���s"O\�8t��9=�ᰱ&�,<&P�k�"O�qq�ZB���AS�=�$"O�5B�,�S�~teɌ*.؄��"O|�����:S�5�v�K���2"Oh4롊@�Lj%H�r��3"Ot9H$�ˤ$δ`
Pi�/L��څ"O�8�'����D�"�K'�( �Q"O����!]7�QÇI�R�"O�)2�Ĝ�^��5���&K
�ٓ"O�бc�����F�_`����"O&��BÏ�g��u�Ȑ�A6%��"O���5��1���皱w����"O^�sCoY�Yz��YUg��HFY�"Oj��f��a�f�a��Q,�!�"OX��"ْ|�� ���*G;ؐ1�"O.9�ǖ�p�ū0��0���"Or)	5-G�tMq�%��G"O.�;5̞J�"���ܠ)i�"OԽSĭ�=<�����X (�6"OT%��d�CV�S�쌸j�= �"O&���Ϙ[1���j��y����"O�|Ҁ�h��*�X���
%"O��Ti���T����[�A t"O>���_T� G,�&��II%"O|�ja䁐j ���ʇ�D�j	y�"O��2F�ֆg�Ȥx2G�0�(�Q"O��AF���_f�ak�*4EJ�!�"O(,�*:&�D��P:
�@X$"Or�+����#M"�8vcAI�zEr"O̴8�O$P������1]��Rw"OtU2i��ZR�D���A}�zD�"O��ҋH�[��:��T�Hqc�"O�qPP��=>ߘ@A��)�N	��"O�t"F'O#w��[E��y��D�3"O���DҤSB�i&.�dv���"O,q�
�*-j񀃂CYj�q��"O���T� `b6�[�yp��ۓ"Ov�"V)��.p�5Z�Ŗa!zb"O`ui#\{&�k㪈�bRR��"O���cDJ�^��#�g�3@E���"O֔[w�=ԁ*cF��WAưK�"O�ЛhW-�e�d>6�D�'"OХYPV"\y��r霅"��B�"O��TeF@�\H���Ão?���""O����@�"9&DrV�3
���&"O�Y�Ӌ�^�P�����&в5rR"Oެ��+�,5V`C4�)�d� �"O4!�M (�j��/P<�8���"O�A	uF	�y�x�2,�"n����q"OR����@�X�	S� ��\��"Ob�zV�I_V��������7"O6�� �$eEV����J�^� "O
��C
�Fp�`�Mӓv�p|y@"O��ѐ@�Y'�Չ��Q�KEr!��"OʙӲcZ49|�T��K6_�%R�"O�țB��*R���pNI[Z|1�"O$J2m=X�4I��qR�T�p"OD��4�ɹ��E�m�6:H�� "Oȩ�6�B��|i���J�2��0"O���"N�ܔ�eB�)HՒ��V"O�9�%N�J���c��9�f}i�"O�$3ǅU�c���p��	/�.g"O�a�G����9HT�#j���&"O� F0�m�i.�h��_T�@aI�"O�tP�C�ď�A�Y�e"O��b�.J�=��+a䛡5qP""O,,R�J��-����0K1��b&"O0� ���Gr=���m��PX�"O� Cs���;pd���Y|@D�#"O.�c�%{�xaS5�� �U��"O�Ē�,�Mv���!$A��"O|D��,i+ !��w�ڨE"O5��$[�+䦑*ԏ$d?���"O���@B$+��Mx��@�A��� "O���H&?�05� �(8+F��"On��D�ǥB'@����:z�H�"OHZ�E�m�HX�H��Q�	��"O�fG9	��9�F�=.���"O�Eu�G,Az
�d�@/��0�"O�E��lQ 4�N"� �`��"O�I�G4B�<��!մ���"Ot�Д/U-$��]Ɂ!�:~$"Ov%: 	M�|�x�!���**�J!p"O�𠲨�q�����7�8 �p"O0HǮN =��b��պ
�v�"OZ%{T,՛5(��rƄ�@k�T��"O� ׏�!z��c%�A>���"O��B�a�(l[t=�ă-(2�Tau"O���� ~ִ;�Y�!�zR"OV�X0%��ab�-9�]8;/����"Oδ�T�5 �jG��HoJͣw"O.0��#u^�dn�"md|�q�"O���u�_�BUR����	|X�0"O�%�n! �u�q�%hV0Ա6"O49S`Ç�	�&��_C4X�"O疴�B��IװZY�a�"O^�S��2-�Xq0��H�=�%"O� �g�X!Ct���65�Zt"O�1g�-�4�� ��.(�"O�x�ĦC���
Jt��%"Ob-�$I�3TJX(p�I���C�"O�D#�# �*Q�G$��t�"O ���	;v@-Pn�����"O���edǣW���Ҍ�E��B�"O�!��ںH�ܳU�'"�m�"O��!"M�p�pykSǮD-�U"O
0�4�{�Bo�L�"O�Q8 ��	0���j�m_�A�b�H"O��X�W� '���$7M(�"O�i�0g�&@#e�ˢV�+"O~Y�0�W��)�U���|��=�A�|"�'g���1�%'��	�ΕMff1�	�':���qȕ&F:����:V�$�k	�'KP�7䆪Ob�4���0R��]��'��SSL��rN0'��K�.�R
�'s�ى5��(s�<��Aqx$�	�'���� �*.p�]rT.�7C�5 �'r���r���@Ϻ�#�/�?���K>�
�c��ܣ�K֎��FEY�[ ��3>��U�ݽ����̀) ���ȓ`��I��1m�j�"B�?u�J��ȓe=�-�$�?*�Mqf�>>��!��p��Y��#<U4���ȱ� ��W���b�<]Ԅi���)U,���Ed���d�Z��yi��ܧ�d �ȓ���Z�@�q?:$�DdԊm��(�ȓ\�" v��c���@�炬r2���S�? "�P�'Y������#Ϛ=��Ī�"O�	��ْ���RF�K�/C��t"O:UZfm��n08�� �v6���s"O�B0�K6�٠�^4"�3�"O�pG�W�Q���+Q���I5��"O�����;"����KׅxX$2�"OȽ�#@әH�N�P��]k�Yk "O�3h�(0hY ���<<�qzV"OB��&n�'�rdQ4aW�h��d"O8�@�-a`�Ж��5-"@|ك"O�ap�H�7���vN� �U+�"OJ�3v�?42�ӊ�\�4��"O��P����a�ԧ	vø�r'"O�}Sw�F�x*�@� T�"w"O������:��1aۀ[R�e�"O��b���8�� ��^)6���"O�(�5��Z]2e�uo[z�@"�"O���u,A+.\������Ig`u1�'���q0�-�.ē�7 ƌ���	3D�(���9?��&�ۜ �e�1�1D��C��F4?�%$�s�1S���	�y�&M�.>�@XA�K�RD�rv�1�y2Ak �u��'\�N��@�B�Ɖ�y��I'B��kH�AT�ٳ!"�y���+@��X�k�&=�h�Cϐ��x¡]7Rp7�N:d
�Ea��&�!�&N�TPVa�� �)ai*`�!�DH7T�݋��X?�48�h��{\!�$D�f��)0P!�?m�<��)9A2!�NBw�#e�׏Bp�xҳ�SF&!��t�J��%kX�4Z֕!)��!�� �{�<�g��::jh���x���1Oj�P��O2v���I�o�0��"Ol�A�&�8{bp(�(,B�)(�"O"t끅��(���bK%K� ��R"O�|#��S![��@Xfg�@�N��"O���D
4(��`�����k��3"Ox�l� �qf#ة	�Ԥ��"OF,b���⎽��"��u
"O��JE��2�@�	ʦhQt"O0�����k9А�ԏK1.���"O>���Ρ�	��OE��m�"OKF�>���3�E�d
��K �L6�yR�Ɋ^^^�K�e�]��%
��y�a��xS�nR�b�3�cK��y�؉�TCw�}�2������y��V8bNw����_ �y­��l,�g�oi *!�L#�y��O�R�����jG�Pjp��ʁ�y�D�t��H6GR6��A�W'�y2�˕~��"���'��ţѥ9�yb
ڼg���X�
�	B�۠Dߎ�y䖌?*p4���ܜ_z��`�!�y�W�9����u'�+4V�� �@�y�%�0� �0ŏ�niq��U�y�4	���)q��H��,rɕ�y2�� ]���aJX�m=�q�v�C��y�՚Kb�|q��/\A�( ����H�<9��`����Ջ]D.�ȓreva��� �h�2���)Ȝ��6����Z6j��f�w`X��ȓ����`#.���Ĝt�8���iVʕ3D�ԖX+1� E��d�ȓn��U@��K� �G�G�����S�? �);s�ىR�FU��h��	%�Qȁ"O���iJ(ZX�$+�ߧf�!R�"OF�Q��z)N�[�k^�s�VQ��"O�Y�#�̋@_��j��
>a��b"OF��@��W�,Cb
Ee�����"OșdF.��<BlS1^�N�t"OܠPs%W:xh�%!�l� ��c�"OR�` �Z
	�H�s�I��r�,�I�"ORՒ ��k#��ZT#�^pbذ�"O �`]���yyС�:j ���"O�1��@	+l�@g��b����"OYW�O�R��yG�� �D�*C"O��� W�JB�����ԕQ���3v"O�p���)X�%J� P .�X��"O
L`�K&J�
ШP/Q'��j "Ox�U��1pT�MX�/W�&�F��"O�-���ݼ4P,�D��mwT8B�"O��ǫ�E� Ô ��[P�X"OH!�vj�36�b ��(ƩkCBI��"Ot�%̘�9s��²g�+jasA"O����^,sZ��� ���d"O���P._�fgi����H��"Otʂ��f��p��S:/e�&"O�-;��[�n�|�C��l��1��"O�8�"#\�m�ހ�oE�v�t���"O`����F�p�C��C����"O�1�j��������\N��)f"O�Y�cK!,=�e���\��}I%"O�`@�_h0`+w��Y����Q"O��ض�؇Q�D�чF�s� ܪu"Ol);&�� /��5)�̞���"O�m�%fL}��Gk�- R��"O��H���i(6	 ��O�<��1w"O�±�\1o��ɸ������`Q"O
F���w ���f�4���s "O2q��#Ǝh��I�4c�Fd�Ҕ"O������nX��9EKW�xӲHJ�"OX�U�Ӹs�b)`
�Ϩ�0P"O昂�e#6e��3cT*_�م"O��3�IF�F�T���Ѝi<|d�%"O��� ���U��4��"Q"
#P"O��F�c�����f�B�X�"O�-9��Q-aFH��l�J�:$ g"O�l����HHBv�օK֌�05"OE�����h���Sv��j�\̨�"O�Z���4�fu��/��\c�"OTU P�'������ Z�6x�t"O�9��9+���ňBKL}*�"OⰂ��+�1�3:�3�'���EF����,�P�(>�<��'�u:W�ȏmc�Р)X�;^4�[�'�F�SA��S�)s�!�=5��ɚ	�'xj�A�^�h�u�;+�4��	�'&�����+�$�H&e�>L���"�'ʄ�d�Դm�Xha�LB�Iun�x�'����K�~=�Y���A+^)�	�'�R�!Pj��5�ޘ*���:.�J���'+��o�Q�[�|TKa��U��'/���!�E�!�ry�'�Dd���'"��a�L�Vic�/� ,�|�
�'�.�T�UnUr����9�	�'�̫� R�r}��uGHuC	�'����d^�F̩��I/g'�ث�'���B�+82��X�)��Y�@�8��� �|�+JT}����٠m�င"OH�X�F�9�vMk��Ro�x�`"ON0	Ł�� ^��#DB|�|��"O֡����@���C+�:�Ӥ"O���c̥E�Z�׆Y'."O�`!��h]���2�\#"���V"O�ـ&/,I�M���,X*��a"O8�f�ɖ5�r9ZE	J+ބ��"O����0��gƟ<;����B"O>��. �ri"0����h��"O�9 ,��'���"c��8؈��D"O<�C���% �D��s���,�$�`�"O��KA��c���QE"�=	P��"O�Yr�oE��s!�J�
Yiu"Oy���X)oj� �7!�mި�Q"O��y�J�E��F"�o;�98f"OjX��f��U��k�斋 ��	�"O�����
c��J�.p8�"O�@CE�Q���@5�Q'89#$"O�9�u�V�+6�Xۥe�?i�!)"O����l��T����ì7�����"O�H�$I���y;&�����s"O���ă5�֘"@���v�r"Oށ�d.]�x=�D���!7��z�"O�l�ԗ.�2ԑV+��>�X@�@"O��X�*N-;3�k kB���:b"O����a?F�����D\Q�"O0���3uO,���.�Eh�"OT�5"�4&�dL�6G�w�Y��"OI�+\�ѷ ݣ0�
�i"O��3iD��IpT�N`n� jt"O�x%��[����Tm�.Y�"�"O�y�$�J3�T��NwT�i�"O4ɠ����LL�	V�*fj8I9�"O����xӨ�YCG>��� �	1D���g�Q�as�U2C�!_���"��<D���"�G�/y"�9ϕ=�t��ą5D�iF�6yjĳC�)Z�r�j4D��B�A��J�!I"K��E�α�4D�@��`A0I���`��Fm��%�d<D� � J߮*�ȸc�����i��9D��:�nC�~m��w��71oؑ�b7D��A�4��1F�Bs�U:sG3D�P�4mٻcì$�2'U�d��jq4D�4ɡ��)}�B�f�my��xw�0D�@���? ��\��E�'*p@ Hg�4D����BB��^�a1*A�B�>�2â%D�
G�ݫs�N��_9�8�K�o1D�8�p��zY�T�^)��Đ��-D��#��ӷ3�4���!��p�s�+D�D;�ʷ7͌My�΃-?h�,/D�hxv��<}P�ܩ�L9� �kD�,D�Љ�b��I�Ƙ�PF����U�D D����oU�)�T[�DI�E��UR��(D�`�¡H_�Xz�b�2p�\�J��<D�@Q2b�'��q)AJ��~  ��j;D�$���'.��1�u"��F �1%/8D�8[�
\f��ؔ B''��ca�5D��!�ʍ')�6\��!�N�Jp��I/D�TI��a��iP�D��>�:��(D�x�ꈿJ̀J�<Sg�X'�$D���an�)#��fG8.=*�s�"#D�Ђ�\q��蕦32�&��6D���	M�j#BmЦ��}_^���(D�� ��Y�A#n������GP8�a"O�)bQ�E01���j�CN~��Q"O%ꇋQ68�^̉�a^5i�� �"O���W�he�B�P	o��ܹB"O�5Sq��9R���H%����<D� +��L��t��ѧp�P��<D��s4sV]��O]0*�����&7D�`�1��1BN\�G\)&����J*D��8eFM<-ab-+�NZ�2�d!�)D��ūW�^�eGbR�l\,�;1�&D���c�	f (Q�5"�_j��� D���b ��&���r��0|Fc�"D�l{� %A���R3��#�J��>D�$
�hO�`��2�@��s������/D� ��85�PT҄拣L�ȉ8g&)D�����H�z>�)�/�4bU�A�'D�|Sb�:2�%��2P(4H!D����G��\f�L���0���4�,D�$�`�N `n�(T)F�*��̢��<D��y�%Q�(�9�G�sa.�q�<D��9�!դl�=x2Ƈ< ��k:D�$8�GB�\�ȼB�*
a޴�4D�i��Y��6N�o��@@�%D��C0J��=� �c��cN�QN!D�$I�$͇6>��3$R�/<R��#!D��Zplө�6�$�ĭ%�hQ�w+!D��c0$�>ɔ19vLC�3j���t!D�|@W��n�RM���b�(0 �=D�$��i�l�h43K#�q��<D��4�n(�UY)R� dx��>D�p�4(	��lx���Z���ҡ�;D�d!�-�d�L�����B�P!�7D��R1� �����?da�qs׀;LOH�@�7��34�XQ��A��sF���v�;D�L�A��)�  ���@�"��m�!'�IF���ON��XV�N.\�*��W�P!��'ŢMX����zd� ;��N�z��M�
�'��]��/p|d�A6���\_�,��'	T���Y�IdA&Є[�(�c�y��)�ӑF:���CZ�F=TX��M�-q C�I�k?$`�	K�LP�8��)9��C�	�IE�9�qL�|:lY��lC�ɸR�࣢G��e���{"�Y9�pC�ɭ�pYqU)�.�m���2Zd��'(1O?�	?gr�2�H���9����Y�JC�	�m�j��T�'S��UT$Ԙ�<�Ip��໔ϋ TTB5�
�;]��� 1D�T1�o	�t��؃��g���e:ʓi�xˎ�=���9��� K������y��]*v"�M�|�Y�с�
E��i�|FlA��&�1e�֙Hg�"��	I���,�ɯm�-�Ӄ�@����󄁹b��B�	 /�Q:�c��բ$��W|���u؟�i�����=�1�����)5�'D�(V�j�Hw��,Yt\�P`(D���U�^3��}PA/U	v�ڰ$&ʓ�hO�&Z�����X�X� (#��RB�	/\\�Aj�
Z$D6�Cb�ϭS�����.�DJ�L�
 D�92� ���u�!�R�ԤI�+"]:��4:�B"�}�'����+�!�&��'a��%�x�� �)D��(���~B4ق$��zl��E�&D�abΝ �|l���J�QMh�&�/D�8� �_.���֕7�F<yv,-D�� ���2դ��!��t�"%i�"O�!C
�[�.�z4*B��
<$"O�[�aԾ'�d)׈*qX^�8��'�(�<Ad���sp�P��	?|��8�HF�<	�8z���@��$(����JM~'?�S�O[6�	�A�^�r�ƋD�1��H��)��<��Ʊ�΁�C�K:sn^ ��RB�<q�ᔚ�^�Q�+W�I�A��ʔ�<�
��,$8�Z@.���bcم�FX�$�O�3R�K�)}�5�%E§Z��@��'��'�i�v����`�`cW)F� q���'�S���C9K��Yy�E��|7�Уa�X��OF���k�-�d��fj�@�|�q�DyX� �O��9U΁�0^j����p����7"O�%��ގ+��	��NNF�4%I�O&Ͱ$/� Fn�8���70�yy��#}"�'������,D��݈��++�X���O������}�j'�� / �CP�D?C�a~U����ꏩ\+^:�H F�Z��v�>�
��P(&$��7��dB�"
���g	�p����'l$��'���
H���ӮeH&��[�PE �[4w;0�ȓTAf("V���/j8`���f���'�a~��>mP������qT��а=9�{r��_�i#��ݰ,[���D�	��y�b��+@p���0k�y�G�D���'���FyJ~UC�0`c���R�����`9&�UV�' �O��'źl��"G���@���WB1Dy��Q�ܪ��%���`Bǀ2Yݔ���g���?i���CRU���
Ul�i7�X8,�V
Oޅ���?#�V-#Ü	Щ�|2�)�Ss �LIe�j( ��z���'&n����|m��:�,J�}, hs�y"�'�,ѺצT�t��E	{��k
�'��X��1�v4��ũ:N��	�'�>��6�L'h�~PZ�C��5�ޡ��'0��@"Q|�4{Ҡ֟*8%��'������YX�P���ة�	�'A�Q�#�.<[�0��w;d`	�'�`�
љdxȅx���Eb�{�o�'<�'�� ��N�"8�
�K)"��
�'�D�(�#�#y�(�_�Hٖ�u"O���e9>���ҧ3*\IJc���'�ў��,!A�<F�
ё%���T�RX8"O<1���x�&@s�Q<Q�T=3"O�ݪ��-3[jX��F!z�޹C3"O4p�2��7 *a��F0e(���"O�h�q�S�0%KkL6y���"Ox�)�b�1V���P�I�;θk��$8|ODZ�(ג(cؙ�È.Hn���"OM�5�οc�\a:#h��+�yqP�'�	D
4��a-��%�Ш��iN�*����q���qJ�5��{��]�g�ȻM>�������|����0$� � (ɳ"O�i�'��*3�`1C�X,m�*�PA�6�SⓥS"�d�a��Q(��Q#k u�jB䉰 �>�u�SM��yc�n<�C�}"�i5>�C@��V��9J�M[tM�o)����f?i�� |��<��ů?���Q��M[�z�Z�RK�4Di�Ӹx���_�O�h[�j�p?��j�d����,�١FN�e����!D���'͈�-pʥ�QbȦ���C�=,O����Is�
W���Hءe̼8�p5�M<�O�Ϙ'�����%X���kg%��7��MQ���1�g�? ���`��:d�� pQ�R�a��٩�:O����� �慪e�>����&+�44y���$>�ĝ2$�+ٽ-�2��K�[D�~P�d�fعl|X�s���'�L=���*}��'�6�S3V� � ��]۩OVc��D�T���lU�U����8�#�eΞ�yR�T�s[>��eC�-��)���'�ў�	�䂔��y�B۠_��"G"ON}�!�Ʊ?����4��*^0���	g8��A��\��$�!ԩ�Ah�c3D��ذ'
�p1�y:��71��9�2�(�	a�'�N���'֒�܀s�Q6=��,P�'�EyZw(�'~��P3��!�S��km3G�!����`�v��I�r��w.E�l��I.�yR�/ғV�Pa���(ƈD��-WO\$�ȓ$4&��#��$r�V��)W#�6}�O�=�bE��(�Gb�C�АbJ^H�<��:`�Xh3���		���)�o�Fܓ���hO�%;F��2����L/x�O��Z�b9�X��.�E�"����6`�!�D�51I�SFD̢m��LPw����'��'��?I�Dd�"�bAJC��)&�aT�.D����d��b��AwANh �G�O�7�<�S�'��^!+d�2�C[�xp�uΕ r�!���`��0U�?�jq�U5=��o-�|�DؖtoH<�a��)#�y� hӶ�0?�,O��1@�Z���X�.A�W6!��"O���-�;+����gKD2(��+�"O�� �'l�}k��N.
�f0" "O8���LUdy��̐t�"O���&C6��5��J��b�I��"O�s��T�y�9s ��e(���"O��sASB>4�!��S1C� ��s"OT(gl��\� `¥�7�Q��"O`L)2�/aH��Eg�&���"Od!�W�s�Q��E�	w,}�t"O�e��Q7)����پ���!�Ó\uԩ�fɑ�)+�Y �ժ!9!�$���p�I�`O������˿3!��=��@R�J��߀{�,��<!�K
{6V���-�*�}SҊ��&!�$�CJ�k�	I�P�0�)���q!�ѹ+&�	ԠE&D�
�:D�`!��ϫ	�����#5.ʒ���<U!�$���֌�@�E)t�.�ʆ*k!��;y��H�R����ZL;׎4cb!�-p�qu� �<�ܥqQ(�7jI!�d
`�L�����$�28�pD(:!�DZ9:�8p�!��{��t��E!�dA�Ww��J3C�1O�Xc1�	�p�!���;8�����;]d^����D�0�!�dŪM�p� �&��uKv���
�9.�!��N	P����/eI|��)ġR:!��@v�LBf��n�\�q��<_�!�dP�`Dp��Ð_� Չũ��!�D�7ij��)��A�PD�v��?�!��'>�[�D��S�� �Vh�>W�!�d�9=�M�#H��w�T4҄M�2�!��	1Rk�5���	PE�����H�!��9��)���i;�t+u�	1D�!�d��Cdlu�B��>u�V�7�!�$Wp�dʥN#�
�Q��%J/!�H�Ʋ�����l�FY(�g��9�!��R;êm*͎� �Zh�F��i�!�� 4���&:rVѹ�LT�!jp��"O0�`�䕃l&��+˄�s�N��P蒌AF@��J9%�R�A�'�&�PnU��"�5a�.�@��'�*��4[����eQ�����'Ȁ�#�
ϫ�N-�U H�}U��[�'h�Q��ނ\��6���jy����'���"��5C������:g��9��'�1�V��&��!�^�g�T��'&�������9qV=i�ԜZC�I#��"��^|!@�̀��C�	;3S���F�A�%��1m�� q�C�xo�$�GW�:�=s2/� 0�^C�ɞSY��s-J�NΑ����7�C��0����BtI�hh�NI�*C�ɒN�0eqehAL�Lp��:*C�	}�ܐ���˨:�oʔz�C�I�s�b1됎��8�$�¡L��C䉿Mf��� ).p�؅�BڈB䉯(\P�,I�d���P��(	�B�Ɏ����Ǚ�0:��J7�X�	/�B�I���Ī&D��c��ʦ�ܮY^RB�I0���2C�=Cf��#�e�(.��C�	2�x�g�ʚJ��'F�8��C�8��Ei��ܤcq�2�K�	ntB�I�d>B)y�j�h� ��d�/�C��&8v��1eT01�Ԡ��'��Ms B�IZ�a�&� �`��NB�I�p�j�1GM6og�l��`� !�$߼pݐű$�֢5|�i���fe!��'Rc�)(��3|
����Z�W!���7<�� 5+	P9K���!�DM�i�x���W�,�|���ϋ6/��~���5��q�!dF�OS8�9C�.s�T=Xe��u�<IA��4PTL$+n�=�E�S��Z�'jV�rmԕ���~��L��p���m.N���Ya	�W�<1�������+kRl��b�#.Lȑ*\_z����Y?E���[��@�,#[@U�ҌD�i�Ʉȓn�HA���H�q�dh���.Ԕ��:��8���'I:���� ͉��O��(�-��O|0*`�C�S=�H��'��1�
��N���u�hY�Cʌ	B�M��oXI�'+�Ȩ@`V.t �lK�"�#��I�r��"�Z��с��X�H���\�Ӑ8$�u�S���M��a*��B�I[~X\:#		K�t����葵G�7�����J�&U���+�g?1��x(��s+�':�p��L�<��%�$Bm I+#k�
\"���B XZ�D:��R�6�����a+,,��;��O�|#�o2k�*�!A!\76c��'24 ��dg�ę��޼�rE.ƥK��]+e� =?���Q�ȠV��~��PxfHa@l�u���C��4��'��1�p��J Z�����r����>�8�Æ�E*'�NKA�Z�G��B��?=��ZqT2�A�5�� _U���à)\iQ�N��\4��UE,�'�~�o	�	BN��㜠G-T�Z�n���=���X���]�ȁ�7�G�{���U�	:������(~�v4�W^���c/�̺+���ã�؉q����]�eA��D5sKqO��s7ڸ'�]�qq'�ŷvG"bA)��4V<QK��8?���q�)� 9x3E�5�p?�򈇇}��xz3`��uӃm�#*�v`���<���7d���Q^,"���Q�n��hs�8�Ī�"Ϫ0���Y@��0p���SG"O��{do[=Q�����b���ŝ?F���u��<I0E`f�
)]��K�/�?T���˟�D�4u:����$ljݐJ�~;azrb�3�vx�r�?i`�u�jd0��K�̬{������A) Z�t�`��Ե5�ϨO��Rb�
�HEZ6��-ߜ�{���E.Մ�d����	�_�-q�h�5YF�z�n�S��1;S)i�9+�G�U쀉��	�$��DBR��1�
d�5ə#xX�)&��F1��"�$JM �����?a4��B�4J��}����<Y�
=��cRk�<�wf�6x��,�vн`,���n̸yb@�׉�o��� �Rk?�@�>OHh�'���S�? �)"�d��3CoK�f�d�I��'񈍑�Ř2B�Ҡ���2�a5�6�� JZ!s����'�`��3��h����	0�<��ФI�z(vu���['���\¢ʒ]�,��z�+X�0�>�@�'���vg�;V	�e���9D��R��Jnʰb0fU�%��A�IW,dJ���=ф�<�`LS�[��Ijâ�3X��8�5D��H�)�)w0� �Dʂ;=>�9��'�K��W}B�P;��9C��CO�<9e��1�d���:f����@��H�<)6�,lhP^ؔS��/`c�!��b���+sC�UY��XKA$;#FA��p9��%�B9�Ó@�'@N��ȓ@�|m;uH��|���#7��2������R�`q��j�x��	��,2Uy�#%�
ap `�!�YÊ{"���c�� uX` �ޟH!wI�;IQ��P�ᖩR�D��)D��C���:�>i3w�,�us�q�ܼ�G�&o��7��9a� [��5:��S�S9i�ȵ��_�-��A#������DK�o�T���C#�ybOK�����G�� ��{�+[��|;���~�ʓA``�|�'���6bʠS^*!B�χ
�yX�{�gC�(�"T�Ht�O�p8r ̞v0�a��a�e��NǢd��١ǀ��t��d�O�iP(ׇ0���ٕ�"���O��09��O�lj��V�mf��T�i'lz��F�4H���F�����y�'���:#��*�@��-�VSB�-p:z��� ]��R�T3#���:��<%?5��l�6Z&q`��¸	�t����=\O%����(���q�'" 1�$�6wW�ٛ����{Z�y�B��D�IC7��<�r$9�gy�_��8�T��33�Jt�'�����''2��@�Mt���D�DJþ,� 1���+~,p�1d�\;�6�� Γp����"7lOtac'���t��U��n��'f�	s�׷u���[�߅z��d���'{�^,R2&�3`v����S�T�	`$
e�T�� � X!�Đ�B>}1j�67�ZŢ�nC�"�F��&-&L�æF*Z��a�t�!V�8�O�i�O_����j�#-R$)��Ϥc���3�2��D*I�pX���EE��IبD���4+���9F_0vV�B��!X�ԲS�_�h�qFBC�^�=�3�/��4��7�����%�܇y��LI�@!$ވC�	�Ѵݠ�I�)8�$��T�+�z���y�\��ӫ���)�'m�.%���a� �r�A��6��dJ�'g���	�
����ï�&�tC-O,�{3�μp�h˓0�~�C�k��Nd	����'ꖡ��ɭL`��	%킑j��V�?�H�&�	d�ʉ��NX3����SO��sꛭ �*�r�A'(���*Q�x򂃋LU�ţE��9kZU��X$��O�ԍ$���0����,[����	�'s�|�fo�"}��=R�B�c��TgK�i�1�'H\�� ,�.�¸O�'k���(͖[7�W�.E�.�3B�,�<�sc��rr�-F���o�8O��A��ߟ(O���@d��<�����8���HB�p_69�R�ZAA��"qh�c|����	h5y�� Kd���K\�LOڤ�S�@���(
QE:�C֛��Q�����z�D�@T �b���H�D�!�4��ɧ}� h�Ֆj�>�ڢ�S�?VP0��dm��ɔ�o�RH�gA3D�t6�C�	`�/�FL�wC�(-y���>���WV�d!�k�.
dqO�n
�)ڬQ�n�;�j��c ��S����n�v!����A����O9jN��*B.��תE	���q�jҶ(D�D�M�Ffh��I�w�����6�p<��M�9$��!��.?9r�Ƞf�Dh���Nv�D����R~B��>��x��4\��dc:���H�e	�8NO�œ�ċr�O�ӆ#�mZ#3���C�T]©"C�1	LxB䉕	�r�ڂ�	���8g��#L�JP��{b��&d'��vј�a0+��l���@19���ȓ�J4�6�ޟB�����N����'�F�����yWl�b6����@9����'q�����<To*��UďE@jP	�'��Z�՚$;�p��dC�9V��y�y��)�J�%��Dߠca�haJ�	�C�	JZ�(Q����L���Uƅ|#<�ϓ��]��F�$7�T �h\Z����S�? B�Pvnڽe��˔ �k���@b	$4����=>�2D�u�U�iz!F!$LO���r�� ����'�QS��� D�����Q\n=S£B.^����T$4D��K�Á=g$&����D��DO5D�LPT��u�Yp5j�'Y\(�b�>D�D▩^ w���6��0�p�B9D���u� j�ʇ�͇o��Y"*=D�p�L�M���wI	48���S&8�O�	���~��Ɇσ�f�@1'£X ��'�EhS9e�j� �#3>�iN>�#�~¬@�@��9�D�|��J�4dA‒=�d0:W��/�$��	a��u���>S� ���9�$=*����!�"�LKpt�s�c���� �<D���5f�=��c2�"ԣ�+K��O��`C����O�@أ���lx)@"ȧ`ͤU��O�����ŒJɖY� ��yq��!�@>�4��m�!�SvNi�A�H�n��0�t_���êqA�'�e E��F��'Ѥ~�.���J��E�6��HMw�H5:e�P�&��QQ��C�,��LY��4}��i��|���K��^'��\2��Q2�V�\�R,�'�3J�����cPꙠ�OŒ\|:5���4+ĳL�T|h���8���%
���Q�P� HB�@���Od�e'#l�P	��	�'�^�c��L�s��#��K���,ľn��Q?���X�x*֌!@��xH��Bg/"������E�
ܱD:8qb�>1b�����(vv���$�';�L� �+ĸ1��,�e��.5F"a��8OF�#Ӊ
]<��BC��'<�R�P��y�ԟ��j&��||�Q��>$�����,d�i���F�7l�D��"1��
�n�R"���A�$�N�=Zq9�/�)zB��F�ŀ�@ӧ��Dx`�Z�J�I���Mh8@�∥�\r�>`4�tj�1O8�1��§p�(�k���l\):��m𕌂���ɵe���W3	~Vp"��חа<%E]�� �p�Ax�y�� �<!����`�A�$xɦ�J!�o´I��u�
;v��z�ɇJ԰BI
�VoB]���>�OFM�b�_�2�m���8IP�-x���;?�Xh�-��~B-�gr����i�m��A�9HQɧ��ʟ2��y��E66\���AF���O�!�Y�_^�ih�O��H���F6%y��V���JU�"TDy`�'��xu�Ii�S�O��	�X�;�1�t,�%5G&X0�O����/�a�.�O�>��s⒂'����OϘi�l��)1D��y����)�y$JT�V�G�.��U�R�˓
g:��`��~8��C�E[
B>��ȓF=� ņ�F�>�[e*L�Z��ȓ~xA,D�!%D��!�6�T��ȓH������N����T� �T��чȓSY���a0W���P"��%��+X8��l�S~d#B�нB+�!�ȓPvN��O�&��ђ��	?-FH��	���+4��->�d�:p��9Xh�ȓA���ȉ��cP,F�_�,���x�#ef�^��'Ɯ.r�0��*}d��;?}�գ�@�f��h��I��+��S}�J�;�H�`�(�ȓh�Di��F��=�a�
|I�ЅȓqW� ���	���UxD�B&(��ȓ:��p�W'Yc������%���A�U(��M�1�`Q!��& B剪;n�$!���2=Jؙ�,��l>D�؃����{���"��Dq-�1;�?D�X�d��Z��d{d"!z=i�H)D�$"��ǚ<�X����U�52����;D�������4xG�9�J�@�ȗs�<���#oߌ��*�ilpyPcBD�<cn�)c�����[)o�>�3�+�H�<�5La�ͫ�Q!
jl�I K�<�c��26qpb+W����Б�FG�<!�g֜N��f�ܙd�	P4	OA�<)����\�Ru!O�1�8�+P�@G�<�o�t|3'�Z}Z�I�u�F�<�%s���ʑ�(Wx$�2��z�<Qï�
�����JH&�����
r�<� �p��2��p�f�:K��M�"O,�1@��P��s��K��ҡ��"Ol��N�o��t�s�!|��b"O��R�AX)f�ؕq!
%��"O
yK�Z*L!F%27;_�2�"O�m�2́)h�hbi�	�j��A"O\�����,�@�]1Ko(�(�"Od��.�Y�֌ �eD�uAd���"O����+��Pw$�&OW�0)`"O�-��G?%y�L�`c�:A4��"O��%O�}=@�C�!0�a(�"OX�S$H�25�`��"�)(ȡ�"O����%� ��U���k��"O���6�aO�h#�[�M&��!"O�T���_-)DxD�Ԭ�!%n�*�"O�ju�W�mKE� #څ����yR��.0oyR%W,'�:��ꃤ�yb >(/�JF,/Xnij6O���y���}6� ����w��&���y�%�)� l�b��)�ċ��ɢ�y�1]��C.A�O�t�%��8�yr�ʫI����k���Q�@[�yB" jDޱ��tݲ�U� ?�y"'Д8Q�2F��n��DY�%��y��E�&4�aJG ^�)"�H�^8�yR�ٿS�&5!c�%�8��2�y"ɖ�~\��@i��x�+�)�y���5�V���۝| @���O�yBɏ+&�ԋ2O��v�,l�K�yR�ԑ޴�x���r0佚�d)�y2掼nR"����]x��2�A�7�yb)�L� l��̋9�D���C�yRgɀ=��<1	"Q���yb�/n�h��%%�l `��y�π�y�r�7'D�y,�ා�2�y���4鰁%Jެsxʝ $�y��E��,B�B�4Y���:LI�y2�Sbd(aR3M/]��i2�o��y���	Y�2�3�à �fpI��9�y���=w-Ra�i�Bm�!-�"�yJ��F[p���ԅc��U�`g��y".��)M2� �ҟc¹�0-P��y�[4����C�g����铏�y�k\�;�|�@�
�
���ؤH� �y���*��10��U�t��8˳e�y�D��:Qbad���z?
!C����ybK�$h���VM֏h���X���y��	K�@9�i�4l���#t!��yo �CFT�2�$E"�����y��(tnpM�ѷ"���R���
�y�,G��ٛ@Z%V���J���yҪ�� �\�V�Y�<99��Q��y-��D:��CN�9�0���yH�l��LN��$=Y$C�2�yr�W�;UѰ��t�H��s�@��=�N��;|�W���N�n4D3�͖��X��	��c��!9>���L�2�6��=iDHtZ@؍���B����M�1x�ȃ�	]!���9wK6�H#I�x:�
t��XyP�K�����	��"|�'2��)�$ׂ5NL� TY ̌0�'�0ژu��� ���$�0}U�� %�����@x8�TY�kU<�:���	O3���&�6LO�L�$'����Y��'�)RЬ ���D�0j0�P��'�4%e�b��<��g����y¤�
b�ꅳ���p�π �I���'+�z�Ç���:��"O"��*��S� %h&��6K�(�0��O�\\+M�X26!?�g~��˰��M��ʠs��;�fʉ�y"j�!*18�f���,}��J:L��ePrᓁ7mα��IN�p�R��}��2� �%|x���D�	<KT�c�B���~2���q�0�S��Ҏd�H=`��С�ya�0W����C��P&��A������'Nְ�m�	��?�:��:��)
E��E�޸��j/D�X��,��I���
E�C��(3_�X�="�>�#Wa!�A%���yI:D�gM
a�<���9��E��K�s~8m3�]i�<I�ر\�z�*��7`t��Zg@�k�<���_m�N}p�A�&�@�;���I�<a�D��2��u�۸X�:��^�<F��<2��)������P�Z��B��z��)1 �Ц���x!��
%�B�	�w�h0���M�#�����%�;`�~���*��+�)+�Odq+�DXTB%��C�?b��Yc���s3H��=�O|���Ⱦ`��MC�o�O��y��"Fc����Z1ex�4�b"O��Fj���jL����Y
��c�i�L]��bV�Hs��(փC��D�#�ڨJ��)�	�$*��2c�lH�I���z�`[�z�H�˲-��<A�HЉrOؙ��K� #�r�ˤA�1@��xW����	�Q>�n���Zfj�0d�("�.C2��H�=q���rt�P�t4�'��l�"�@����-��زp�'y,���$Ș�a{�3?a D��.�8O��i�,�V�X ��� %��ɠf��-2�AW'��G�Z9�4Em��X��۶tg�|hm�{60��ȓ�~}j$��
����0 pm��h�I�C>@�� �L��}P�L��`}�S���~�1R��������ҧl��H�'��(�4��-9	�R��4���Y�$,�"��="D�aU.�4��Y��0��<A�#Į*w� h�l��?��0���W�@j�T�ժ
�%r#~��oF!<�H}Bre�1Z�%p�L�h�b �3o�'P����'w2��d�!5D��H��-��U��C�MO\�qĜ�~��D�P�h�b�aa�'��}aB+�!B�E5�[0�&�8�'���q�@�b�x���+K+%m�!C�4��-0I>�d��%U7ǔ�)dMc�	��T�+
��$i��_�FD3����{k�{�(�4b:��F��(���B�C�F]���%N+&��b@mH<9rm�o ����0rj@�+w��_�'}�D���`(5�~Z�
W�pw�U)�\$�����X�<)t�ô-��X��C�\�2-�R���D��k�.�⥚>E�4-�0_��i���-7�����%ϐ�!�J��e��苄?��]����7��$��
u")�V'���<	B�F�x@�$B���R�]x��h`O$C���"���6<4�x�H!mY[��X�f���їȁUn!�dQ�t����s�ҍ|.K4 ��y�'��L2��@%8�<Z�ޖwt�A���d��=%p�A�CEV���ʦ���y2� p�)а�fA�6a���U��p�1��"F#.h;��+ܸO�' <8�va��'v��`�U�g ���'�q��<T_H$��3u�8�Rr��9hz���Ĳ :�({�����<� 
��[�.5��#V(і�j��{8����
�^� Xs֪��c�:��3f �|��y�2��	�ň�?�!�Ė
Hf��t-.y漈��\�	Y����#�>���қ���!�E�f8(�����!�;
_*�`C���=�rq�e �>��Е>��J L��>�O��b�'!���S�ٖoIb�;�
O�U���^�G[&l��Q�R�6�J�샵k���(4��'�0?*����k��1�
��D��v8�L:�o��e��:𓟔��L�R 8U{P-��{N�p�*O�����AO���R$�/ �Ǖx"�H�4Z
(F�|��d�ߗq���0lK#$�(pN-�yŔ�L&��B����v������$�DL�g�D��z|DM��KM�:֍îY�!��:F��t��,�Y����P�>�!�
*1I�5C��?.b��m�!��̄s|�UG�3z�f� ��0�!�� zM�r�
�����Ƙe2Lk'"O��S&l4;�б���	*�5��"O`��[�Q��́1CT8s���"O.8 tD�	�vH2�HlbD�"O�t��VEӺ�SF�'dN8�"O.�)�h��M��P�#kM�$]zD��"OA�cC+-9b5J�*�* ���"O|H*�E�<
p"_�]u`)Ic"O��L�r�FE���dPl�U"OP5IbCV"r¬�P�C@pP��"O��R1��5�t�u��v�j�I�"O��b�Z�����S^����R"Ot�k5,;v��rF��o�Ԕb$�'����*��x/��2g�yI����O���{�	��j�WN���ٗ2�
\E}2.�!)��a��i�9,��)�9�Cr��TX!�D2k+Z����Lp�"�T�2H�	<�l`k�7��)��3J0)��Q�Hؤ<���  �2�U��!
%!�PΔ��(S
{E��A��V�ɦ�4#f�!�2��Aj�3?�i&���>cG� ��,Q= ��{��-L\�?�#�E�:�[���l�Z���(6c	+7j��U�!HR� �E��c6��J�`��\�S�O1ƹA��]�w����@@�b����]��U�/���pk�D�i�*klv�>�r�N;Y�|���ڱ �Xy'n�<�%��1o�f��"�=,O����Y`.�e�1S6�يT4O4���f�X�Z�۬ID�'�F�jF6Z���[��K�v 䨀*�h�"5sfm0�P z�1�\ *@�� ��(�%�%/E#�G�H"�:RHk� y�"Q�6d��`�, ����^����?��*J�<t�+䨘�n�\x���<�{��|��'�3A���i�_ (�gj2N1h�s `�0�4�{��B�0�=�4�ƺ.jC����)�'	H��5�L�rb���闩KB��'d�y���D?K�F%̓ ��J�fX:�T�>����(L�����ٯC&ȕ��Ƣ<�S�Ra��*/,OBi�S�_��EK�G�}:Z��!0O�����5�n��g� �il��Hw�F�38��P^���Y����[�|���F#"ܽC�&НP�����	Ň��l2�ǟ0X�����h ���}8��m�����BI�G�i>�X�ŤM���q��C�4V�`*��!�5ZZT℩ܟ{>�DT�Ѣb
%(G�!�F�F8<�Z����S���Ij�l�����S[B��"Pa@t����-�2�
2����]���S�O	�0 E�b���"AE�yf��1�'v�ECv��J[�A���r]���N>�šs_���dB7`�������{�蚃A~!�$�(2�D�R���^�,��uA1k�!�D'7=pTKr�����A
�W�!�$�{�tZ� %aɂ@B�V�!�	�"%�wOZ/�0�o��!��6cSB�QA�_6f��Q4��6�!�dE8H{t9��T>a����햤�!��7O�6p���	qgDh�K9:�!����(��&WR�����Y:G�!��a=,�� ص6w��#�#�yM!�DL%�����C�xt��2$��'#!�ė<g�l7� �G3��XP㗘o)!����(�P�H��8���b(�0d!��O0(FA����2:���S�A��!��P�8�B@'�u̔��Ꮛ;�!��?y�Ȭ�$kĉ ���RV �e�!���<{F@�buC�� ���`!'�!�d�L2ޑ;��[�4��� ��S�hq!�51j�P7劔H(����@�
l!�d��P}�E��
�qR��C�N��!�D��2�2��4�Q�	$I��nH3/�!�ϖ}���h���#4�������N�!������bo^S,0Tr[\�!�DE �p��J.>A1w��!�!�$��K,�$qw�y�i���+i�!��Fg>�Y�ׇ.L��LS!�!�� ��dsK�9��F�%h�$�"�"O�󀝶K�L����,���C"Oj���)F�;�Ta�O��v�P1"O�1B�g![��U9Pm�{��л�"O�q�6`"*�X<J��L�h�:<�"O4���.���˧צ\�)�"O��i��Ƌa�@0��HI��.���"O �p��"w�.@�Ԫ$��"O@�1�kL�Je�A��A$�"mc0"OV�b��w\mi�#��
'"�9$D��lA<<����a)Z$Q"p�;Pb�0{��O�SU����2(U�Ah2����4L$ Y՚>�Ƀ�!i�L�|M~�iLeRr��ӏ�-M�.��� RB��_�[��YH��A$�0|b���T |����&Ul�j��|?	�C��6�:p�6}��� �5	Z�iA)��,���J��+<�S��U�@���>E�t�J��S+��Q�d҄ș%1F��j�$>� <�M����.6Mp5�ᓬL-dD����=�����#!9����b$M�-�JK�8�C�~z��)ϵ�n� �J����Q��%8�X���R�V�q��]�>+bDP�S?�F��ɜ[����R*
 IZt�	�I@��?��

�,����e@��)�GҜ-{�L�\%x�	���X�Xp4�2�}�E��p���"�f�[6�K4xB"l���Ǩx�A�>e��@�7�V?1V���L�$��@�"�lT�MNR���P�@��� ԭb�D����t@�~�	&�I�|��)FT|���umn)�1_�4���/txY�۴R�a@�J?֝ݟT�l�a��}��JV/s��!@�J~Ӕ�)!��`j� e��]I�O��Sm��T��	��լx@>�O<AJ�+Y��xn�:�PG��)h�*Tk@�@6>�"@�� l0�	� ���i��Ȏ���d��B��4,�j�N�gBҊ��	�nԛ<�?O��AH�<t��wl_�)o�Z\�|��h~�a��F�"D�E'��t�>ɍ����D�<+�(z��%O���k�����0>��fķGpe9��A�0�,�`i0.kDx�a��+� ��C��S���`E��j=:E%2�ɚA�LU��S�w��eZc��;���bP
F(�O��'� ��Hv˧V�$��o&b$V�V #����F��8;Jr�'�l:���l�����>﨟輨�.۾4�J��b��6i>B7�'��CÍ�*,�ʤa�Ɠ�t"a���ֵ
��t٣�M�h��y�Ҋ����h��}�
�Jf�qP��ˁB�xS6͇�D1xu��?N~Lb��؊lZ����)�d���ujJ(�A2)lZ}�ۍo2Ɇ�����r�˖���P�AS�6u��Lj�
�dV�Wy����
?�D��ȓ^��)c����LW�T8+��C�fD��`q�I��O$�P���	;>/&���OD�@�-�8��d�7�2%��]z����&`M��PîB�Tơ���e+��H �0�kG�!��Ćȓ]��'�7l��Ҷ��gt���>�\�':SeL�F��?^z��ȓUa����Ί�p�H�fE
��@`�ȓ�H�SSi�zP� �P::���C�^�CtH�M�����A]2.8.Y�ȓ���'�ӭz'&X�cҵQ�J9�ȓ \�}��Gεw�ACA�\�p�ȓu#jm!#�1v��DCƇFK(�ȓ	���{Q�Z�3�`4�p��o�,��ȓ]���Al %ˁ#J�%.���p���cI):�n���"R3�d�ȓ���0�ˋ�t�Υ�t%��-��b��]8q��XDpS$�]	�͆�L� '��p�������Xc"��ȓc��,�"�ޞ+�<I1$��,ex��ȓ�e�a�FH}����fV�]jņȓ"�H'�J�Jf���uL�:F����X���)��#(�!�"GW< �&̈́ȓ3��\*�k.���� xp��S�? (�#`:6���ِHƌ.�ͪ"O��vE��A��QBBH@0��i�b"O`�[��PP��eSe�*���d"ON{���a~,H�W�+jd�i�"O�av�)=��V��-�BIx�"Ov5����a��*��w�����"O��a� �`=(���	�.[3�y���r����c	H4�l����y¢�'`��
�ʝt˨1ᓉ��y��@�������aI�U�r�T>�yd��L��H��� B��8Â�̖�y�'[��D��ʒIU�8C��yr�סp^��d�A�@�$��a����y�j��7BPh1��7h�ݛ!l_��yR�҇!�8�0��_�,a�9@鏁�y"^!8�tX�G)���,(�Pn�0�y���IHbY�T�D&z�vؐu�M��yb91�\[�b��ZD�o
�y��>`
Ⱥ����"�L�Ys�ʊ�y��</�Չ�E	.n<pg���y�&r�� A'ȸ_�$�	U�H��y�3s�1��	͔,Y�<����3�y�tb��!�������/]��y2� ��l��	��n�n�94� �yr�}�B�1���f\Ą�I��yrǤdL���K�O8�))`����y��P�鰤��HB'L�h	ڒ.@��y�g��g9X�pK�:���/W�y"*Z" s@X;@�RW-E"�y�OL�p��{��Iw���y��	G�&N�z��|���_+�y2B�h�r�3��=��2&���y�'M�>�2I`�O�3;��P�Iȭ�y�޹Jf
�x�䈧%@���Vg�,�yrj���s�J}�)�����y҄��7��1�!�;�@� Dᘰ�y2�M�D���0M�70�E@���yR���Rd(J�+إ�u.�$�y��K��<� P(T�o+�Up5Ȃ��y�"�k�F9Jq�C�c?j$)ƦO��y��!�viI�⁻*�2�զ���yB���`�|xҠ+hH	E%���yb��{>��H�ۺo3�m��*�yB�o9Ry�cM�9j�H�C!���yB�@_u�U���aݮ��B��y�6x��`�LU�x\	abD�*�yRhӆf2���eӺ6g����dҥ�y�X;����BC#,�(!���\.�y�8m�������e�֬܈�y��:��A���t4����y��O"�R
� �-`�N5�A����y"M�*R�8�x ��
D�Q�1)E!�y�Cբrj��6�Rx��(��y�`%2]�����(�$�I�K�'�y�mN��������Z�qa'J,�yb�6�|s�DX�0��s�̏�y��ܮKN�	@�1�6U:�bP�y�J�^��'�8?�jXB���yҏXK6��(�hC=n�x�Æ�7�y�L%M+�;�/�Z� H �́��yr�It�.� �ũW2���*й�y��\����MKU :�������y��څEl<C&�E#}J��'̔��y�	�R��%��'S8xܔy��	��y
� $b���X��k��[9�ִ1�"O>�iP\A�5k�C-\n�a��"O�R�e��h��䡕���t\��1"O��;P�؎zMĝ�6(K�H �d� "O]�3l��&�zI��ң"O�kS���+|��s���4)��"O��rf'�'LBtɂcfR��U�&"O��(� U�C�Tu�S	��
�"O�qSV�����W��~����"O�����8�P,�6�	��9�"O������%���g���*�I5"O`�4�G���٠�bD�w���5"O�}�5�ٶ[L��y2�)�y�"O��"ca��2l9vaӼ)V)�W"O~���M&R?.����T�z�"OfH)W)N�S��d D������"OU�2%C vm̅����%�^��"OɛN�5H4��3�]�TAn�w"O +r��PJ؅�b�ݭ1�42s"O�q
�扝w;K嫐��Z�"O�`�V�Ӏ7�d�4���*�dL"O�u!��Xh��aM�G��`"Od�B�">
Za�j��b;V���"O�E���  Dz�oL+N4�u�"O*����.'�:���Ͼ3���""Op=��� �9"�m�JR�$C"O���`��b[�,�
K'h�Q6"O:h�U
��W��$�P�̴ 9\�@"O�<����¥�T��RP��S�"O�U�E�Z/T�M�Pb@�5����"O8�"�n��`bZ�q�BX�`9��"O4=�0▐V)2$c���p�8�s"O�d:�BƸw^
���]6[Vvݐc"O�\� ��S ,��E�+p���"O�[�c߄)}Ȩ��c��X0�"O\U��[��	�bB[�8�=X"OP���bOزE�G}ܝӣ"O�����������%΀�}oVB�"Oh<�Eo�$�@��*�3r_(\�5"O$��r C>����@	 
�x�P"O�4`�Jͤd�ء���6�@G"O��``��)A��B7��k5�(�"O��x�ǅ��2ex�L��w����"O^���Z�T�ܤaQ�V�uV��c�"OD��bH�}�r�P1��j=T��P"O�A�ի�1�riQgFC�uG:�"�"O�Ir�lF 1��d�
C+!��i�"O���+ X1������b"O��l����ɶ)U)%�
i�5"OR!g��0:H@�
Ȭo��D�Q"Obe��섳�����]�wκe:u"OT���#�*Yv�����N��x�"Od��gݨ�l}HA��<q��Cq"O�Dz�E!fY���fd��k��y�$"O`�җD��<�\0��ɽd���b�"OHɉ'f
3���t�̡in�� �"O|����׽9��[�ɓ.[�Xp%"O6��F#V<I�j\ң'�/@Wt���"O
�+CK�F%�PF�]�8YS"O���� ��q�"yq(7~Q+�"O����P���F/$�yV"OZ�r��J)&����&��7��D+E"O������|e�4y��pwAk�"O�#�_T�q���˯FEu�Q"O� ��k���qh)����04QXd"Ot5
W	M�(��q�[,#��H1"O�9��є&�vh�&�pe�t�"OTxf�:��	�� 9J��Q"Ox�)A͏�y�赩����"7��W"O� A��Y��
ҋ_	��R�"OV9@,B~���sT�N.��	�"O�ų���:F�1�D!��!��"O �A��̈A
������Q"O�|8��J�i�p�!��O=	�N!Z�"O�RpEPvA`���(*l�܉�"O�=���k�P��凗)>�-�"OrqRf��+: 4����08�iD"O��,M�i��+U
&��6C���y���$j��	��Ӆ*D\1'��y��ռ
EP�R�'l���5��(�y�7f�H�2큼m60��,��yb�^8VVb�b)�0d |�	�b
��y���̚%��Ƹ���O� �y�(�eL�	���Ѩ�3�Q�yB�M�L	�)RL�< h�"��y"�x\��0%�!a>e�!!G��y�̎+�n��c��щ��yRP���H��bW�I��ba�-�yb��ZZ�C0+*FKJ �E�:�yb��6hW��C�DJG1���c#��yr,�:�h�c�B-P$!���8�yb	�*2D�7 ��At �����y���";gT�X#�_�c2��� g�2�y")F:Uľ(P!(�_��R���yҩN�7x<�bo��Q{��( g��yR�N��x�A X+�d�I�,S�y�m�Pز�k��`���X��y�Ό�1&�`j�g��+	��RW�M$�yrD��zNR��!�FaA��yҮ����ӥ��򩂀O�.�y"�C�>���
�$�����,�ybo� ������R���Rb埂�yR�?�Թ2�E�8S���f
G��y�HG    ��   �  i  �    �*  �6  UB  �H  �Q  X  J^  �d  �j  q  Zw  �}  ��  _�  א  1�  s�  ��  ��  <�  �  ��  ?�  ��  ��  �  ��  �  L�  ��  ��  ��   ^   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n%�^L���ܮ*����EK�0�RP�"�%?���i��O�9O����-t<���C$m����EL�d�O�$r�r����$��$�O_�h���4j���RɀF�b0�yB�'��V�O������^�q$V]*B=h_�1A�l�f�s#��4�Ӟ�M�;U�"M����-V0���L* ��P��?љ'-�)��8'y ilZ�<��!�=�e�APht��d��<��'�$A��hO�)�O��Ѣ�АsaZ���v-���0O˓��ji�&�2Ę'������fڶ����"${<�����e}��'��=O,�)9�<���Єum�u�Q��Ar�$�'���,p��,���#��(5�'�F��7gş ��=��L؍cT���]�<�'U��9O�Til�*�~����Y;��q�:O@�l�!x�x�=_��4�F|	�"R.r�����X��-A7O���O��D�>Y~6�(?��O�B�	��|<� ���f���``�[�3}\qI>i(O���O����O��D�O��G� ���[r艎K�~��pį<�0�iG��;�[����S�ߟ�qGJX����Aȓ�c�4�jQ��DLΦ0�4g=�����O��t���<siZ�CZM�d��=8&И�iB����ZX���1BL?�I���R�a1��icr�k�b�=a�d����؟�����@�	՟�SOy"}��	g%�O�a��d5���A��9v>]Y�$�O�yoW�{��	�M�R�i�47��J>�!OE�v���� _
�)C'`�6物9U���̋#���B�<�+H�����VQ8l8!/�6g��1A!�U����Ɵ���֟��Iџ��	s��%�j]#��Z3X��P�Lު6	��y*Oz�����4m>��	��M�M>Y6iAD>*�k�Tx�.�d��'J�6���i��(} �l��<��f�A9��K�5�*�A�^�-����臬rO��D������O���O���6�:����$�A��		�~���OF˓r���PA2���ЖO��� ��P�XsF܀�oD3o޾���O���'~�6�Ҧ� L<�'�Z!'�*?���y��[�1�H�`C�?r��Z%Fݓ�M�R���S�1��D,��ol�J�G}&�Y��1>mV���O��$�O����<�&�i����ƀI04 ��
�U�~(�R�.�&m�'D7m%����$�ަիF(��M~mGte����	��M��i�u���i���O�`b���R�o/?C��4T"���ڻ��-	��|�@�'���'bb�'��'Q哚o�� `�`RV!�9����4���4|9�H:��?�����<����y�R�^d~Y
�Oڔ%�F�:�ʐ8�(7����N<ͧ�r�'%�f b�4�yB.Dh�u������gj�Γ{�����On��K>�,O��d�O��qSa�y��P�����򄬩���O���O��D�<1T�i@�B �'X�'��t1�QN�|1�Ϸu���s��$�^}2�q� �n����]B�)R9�Q�����J�Γ�?IC�
o��Sp�4���
�a��R�F��$m�"x�)֙c3�����N�d�O4��O���2����*�V	XTJ��P�L�*I�vL��?�7�iو���Y�d8�4���y-�K�)�5KJ3Wߪq�ACP/�y��q��LmZ#�M���M��'s����-��'j��<�u�ʁ0M�p�M�-��L>�+O8�$�O��d�O\���O�0	�EȚ'�S�i�I%�h����<���iw~9#A�'T��'���y�C׭���'����yFJ�.n`��?Y�4S8ɧB���br�D<	�c��sօXKE�NP C1AК��A�Q�xQQ��Fk��O|˓˜L��`��U���"fCY�}.��j���?Q��?���|�,O`ql�Y�z=�I4)�x]�w@eY�����4lK�;O|�og�M��	��do�4�Mۢ�s(=f��0��5��y�|L��4�y�B��V�������?mz�8O����he�=� ���^��Ea�M ��8Ѡ:O��d�O����OL�d�O��?��-[+l&�+g�
�\�H���-�Jy��'3&7M A����M�����^�n��$Q���!dW�;�h�~y�'��o$�M���*cI��4�yZw���G��e�H�B�@9l2Y�g!�!Y�x���'�&�|�.O^���O����O���!˦j�n-	�=I�]�Aj�O��d�<�ջi�dh���'��'��>U�|��� Q�i���I���n7��S�ꇱY��P[WCB�u�2X��+�z�~P��H�
em�&ȵ<ͧJ�\��y�ɢk��y��� �Iy�N*�t�	��h��ݟ��)�Qy��Ӭ0��&~�HI�cnG�

�I8CË�a������DF|}�ak�l!@��P�>�J�C����3�A�֦9�ش4k�iߴ�y��'�,�f�Us�,OT	��f � ������5��?Oʓ�?I���?	���?����) ���}�7��շ���m�Y��ij�&�'�2�'��y��l��&4XdрS�8�˄�X'3�mn+�MӴ�x�O���O̬*�it�Č�6�2HXW�T�.����D>>󤃄85ڴy�o�ؒO�ʓ�?	��S���r�.�'E@wc�����?9��?q.OvhnڛFv@�I� �I�	C�5�5��&�%��h��w��I�?�T^���ݴ}���"�>��������'�<�I�"���O(�V(��h��Qͽ<Y�'7���H��?)%,K+Q�$ec�6p`��e�E��?	���?y��?1��i�O&����0o#ȸ�׋M=&�2u\0�$���q���Zyr�d����,=l+A�r�P�1�m�,T=b��ɦ�1ߴ#'����b��=On��Ή�T���O��u؆���]r4�9E��;I\�qs�|rR���	��X��Ο������wg�3��3�T;`�N
$dUyr)i�J��p��O����O��?�R��	�P�Ԑ��%�/?�@�V%���T����4cՉ����O���Z�):>�P���)z0@�&O�(:��Z��E�=xbO�y�Sy��W�.����6f�_�X1�,\�&F��'F��'��O����Mˠ���?��!����Ʃݩ"�����?Ɂ�i��O:��'�¾i�26�$(�ҭI4V�5�l�#�ݣg-��Qw�x�4�	ٟ{d�JZ�dh�~yB�O��
�0�,`��K�\6l`A3E�%�y2�'�2�'L��'���iJ�Y�m Sa��B�N��V@s&����O��䦩�t��Ty�"d��O"];Q�צ�c*R�+�|�XbRu�I<�M�ǳi�����s|��<O���ҵ^��4�6I	�|`�h"*��q"����?�&��<����?y���?Af�^B��A�DW$N:vD�����?�����dXЦuh��쟼�I�`��?���	�=�u"� �I
�!�a"'?��X���ٴ`q�F�%�4��I�;U�A��c��s�n(0��88��G%=
�HCǪ�<��''���+��L:T�2@N��F�F���u��T��?���?��Ş��DĦe0�R�Jo�lV�.+���V�I�,��'��6m7��-��$��is�"��Nh!��)�5h��r�թ�MK�iV�x�e�i��D�O�|D������<1��D�e��3��O�s�꼓4��<y.O����O��d�O��D�O@˧.�TS�*!_���%l�1tHdx��i:p )��'���'W��yr�o���]��CW�S�+F���#{N|m��M�t�x�Ou���O��}�Ѽid�Ĉ=�1�nC"bTڸ`W�~,�d3�(��t%�O
ʓ�?I�WE2�����t���"W�QފI@��?����?),O��oZ$kBܗ'��!��u��u$�$y�u�6J^��O�'��i{�O�apR�˦UHe��@Ct�S=O�$Q�bT99�'�:�@˓����O��Z��%�A�>��L���1u�� '�������㟀�Iş�G�T�'�<��n#
m�ݛ���,!�I��'��6�DS��˓` ���4�P����ݰo� �d�Tk@���8O�o��Ms4�i��ƹi6��O@�`Ҍ���Ŗ2	�m�$N�)�Ht�"�)@���O@��?���?����?a���X�a���^.��	�OibT�)O��m��i�u��͟���A�s�x�1ߧN݈HTO�E0�Ǘ����̦AIݴ	������O;��#[L����+A6(-��٣�Z|F���Y:�� *j�e�'p��&���'`yP��Z�X����@�U��`S��'V�'������W�`r�4a��,Q��s@0�j�.�'2�b,�j������'��'��k����~��	mZR��0���9!�v4��厏]�b�sG)�Φ�͓�?�+�!���釅���䟸��N�R
,J���H�}�7���e'��O����O�i\��'��hy���zv$ȕ�^�.���"�O��d�OB�n��6@��'�6�4�Ď0*^V��u&�Ȳ��$��'��شZ�6�O1Vp*�iO��O�3䥁=�v�hՍP�nn�%�(J,ܣ�'��'�	�t����	<�֝���&m��T��b��p�I����'d\6m�&�E�'���'1�S�?.0ɘ��>n�f �� A�mX�o��I��M�ѷi0�O�	���y�@''�:Ǉ�\��A�5�3٢@i�- t����C��O�UhL>�0j��i^��i��_(Ҧ@������?9��?y��?�|�+O�$nZ)}T�):�/��lahZ�/��9Úcyboe�h�H�Or�nZp��@�ah��c��P�[�����4E6�&O&�v;O��Ē*s�8�Oq�)� ����%�4ֈ%�0��?��\��;OJ˓�?q���?����?)���?iMI�|�:�Vj6��2խ��Fl�E/9a���.O�ܦc>�`�4�?a1.^'Mv�C�@��i28`�"[6⛦c�<$���?M�S`�d-l�<�d�<o���B�.̽	}�����<�V
�/J����H
�����Ov���/��E2�K��Vyps!�.$���D�O��$�O��H��&HҨl���'����o�Ayw�BiE( Շ�^[�O���'S7�Ŧ�H<i���0��e�H�%JЋ6K��<���W���0pa'u��M;(OR�ӄ�?�7��O�I�3��/�Ҹ��b� #�Ƅ"�N�O����O����O��}
��w^p���P f����E�5o`��!ۛ���	W���2�M[��w��0Ư�>�9#ժP%Xp �'\�7M��:�4v�I��4��$�!������jp���/��Րg��
+��"��/�$�<���?���?��?�b�\�lp�pB��,9��Ӗ��$Iæ1��BIџ�I�L�SG��'����?x�F�*� ��0yk���>�%�i+�7��f�i>����?ɪ�A^<����5���Ť{�R���LayR�ߪ�����2��'���$F����D��Q���Ba퇗1z��	ٟ�����i>=�'�6-�#�"�$ݓm�
E1���̚����e�?AfX���	���cڴD�&�#&�˥5i�h���X�v�1�۠�M�'6t4+U�%d�8�'L܆K%�O�4ט� F��tO�VPI���r�f�	ϟ��IɟD�I�����s����AQmR s��� ��C��)���?Q�Z4�v��e3剰�M�M>�".L�l���+5�qk� "M��)��'b�6����ӭM��oZD~REܾ
������V�s
��[>�I�����!P�|�^��	⟰�	�x�U�H�fji�0cK�u�"x;!�Zڟ��Izy¨a�ҡ�b��O����O�˧4�Ҽ�2�-<.��#�X� `��'l����{Ӵ%����?��HI"F��ru`�$	a�Y룪ѭq���U�=W�e�'�������&�|R�
�J^����%*�Բf�@+M�'���'����_��۴m�5�R� ��aL6��q��?1��k���d�F}��hӬ�1��7�	��e	�&�<X�L���޴D���ش�yb�'뺽*����?	�EU�4kv��4~��X���YV��``|�@�'��'���'B�'哈U��KRcX�x���	2ǈ� A��Yش}����?����䧽?Ѵ��yg�K�q�n�C'�G�:G0=�Q��,;�6mKͦ�I<ͧ����)&A�۴�y��G;=vȘÅD�71Ѽ4Y���-�y�̛\j<P��� �'k�Iȟ�	�W�)�b*��y�� �Z"�%��՟�IןĔ'R6���zV����O �d��XA�p@�Zj�"ǀj�lوr�<����Ms��x!�a�Z���m � �!P�@� �y��'�H
۩Mi��*�<����F�	ğ4)���B� �H�aĩx��D�&ߟT�Iğx�	���E���'��PRW�Ʋ�А0� ;2�	+��'�<6�\�_b˓hh�v�4��x�h�g�������"����O�7�E˦I�ߴ�^M��4�y��'��i����?�
d�9BZ4Q�#H�|@H����΄G=�'B�	ϟP��ßP�	۟���1vQ�i�aD	+t#�`5��-��ԗ'��7�4f���O��d5���O|�����a��".�q �$ �G�\}�n�b�l����|*����EL�S��l��+��P�
� ݂,{��wO������0
�����6���O�ʓ^���a�� 
w�E �.��7޵)��?!��?���|�+O\o�U����ɾ�^�ᑍu��e�7e֫D����	�M{��>�g�i7m�ɦ�@��]y��re�`w"� G+Է�,�l�<y��:�z���h����/O������=y��A?W'^(8�c��&���Jt>O���O���O����O>�?��G �'`��	Ck����A�bJ�Οx��ß��4~���)OL�ml��� ��V&�Aī��c��P(I>Q�4ś�OXYt�ih���O �0T�˥,�3r�ؑqK<�0U�ņi�L���$��O���?����?���xt<���x'`�Dʳh�4	���?).O�mZ7Lfl���<��B��8��p5��7f�@٥�����{}��~���l�5���|"��H����s��,	�8�*҄ũ}cE��	!�l�bjR������F���N���O��4�؏}EΩ*L��9����e��O���O���O1��˓,��&�I��r-X����St�s�d��_�%���'҅pӎ��q�O�AoZ<��Y��"��Z��P���W�&�,�A�4_��V�M��'1")V(xab���1^��I�=N��Ӻ%`���3�6�IHy��'r�'7��'�RU>��+s5R�h�%M"Mb����M#��¢�?Y��?�K~Γ[&��w�N��f��]�궧 
=	�@Ӄ�d��1l�����|2�'�ZD䕗�M��'��%A��֚5�,9�j<Q��ؚ'Kl�Z��S?�H>�(O2�d�O���)A�}����G*֕d���'��O"�d�OR�ľ<r�i�t�*��'���'�N�C�"%_~�;d�כZ�*ͫ��D�g}�HzӼ!n%�ēQh�H!�ȅO��0��'�;e���͓�?��_��fa
Ԉ��������iD�D�4@Z�ЀJY�
qx'�֜n����O����O^�d*ڧ�?�Ō;l������N��I��o��?IT�i��I�Y�d��4���y�CG�d���ӧG.H�X5H����yB��Ox6��립��k�ܦy͓�?Y��R�:]��	�M�? ��B�5%�.�@A��P	�y�F�9���<i���?1��?Q���?a�ē(X=���~�:@��X���D�Ħq��$Jhy��'K��e�W��C��]��%�536PT���tyb�'֛��:��O��$�OkҰB��[FH`���V�= ̳Mþq(gU�H�V������*��)-�uГ�IX�P�;��O�=��O\�9m��8$�H�s��ܢ�1D�lx�� $0]Ft�##گ�D����;�	�y��l�	�Lj�����G0W'T�8�j�1��`��K
�nk����e
C 8�di�	���H�'Z�E�RW�٧��3�P�5�U�;1v�A���w�&�ѳ� Ԃ-�@̇-,*H���'�\�a����T�"b�!%]���\�.���c���L��1�Q<�Rxl��Z��r��^��ڱ �!خ�Y�O����O��O����OUʴ��ON9	Bk�2F�m��Eьc5�A�q}��'��'.�*+���I|�CΆ^��̨�CL1|/������iכ��'��'���'����'�� �*9���W��hg@H�m�x�IAy2�OC}���d�
9��HJ��EҲ@́[�&E��Xt��؟H��>�`A�	`�Ip���ǌ�� b���v�l)D�զ��'�T�J�!i�\��?��'sJ�i�%�v��?h���c@N�k�Ҹ#A�r�,���OlI���O��$�O��?��T���:Q���&JМ��DL�~�D6-�&F�nZڟ�	�Ӗ����<I�'��N@*���? :�=����>R
�f(N0xW�'}��'��Oq"�'��F�\33���p��	
E%�=JRE ���	П4�ɸ ��ۯO�ʓ�?I�'�
]p�R>'¤��A�En�3�4�?����?�cBX�~��������۟H��I��	��F64���JR*�dK"o��*%�Ҧ�ē�?�����{�EEX������0Cv�@0�Uo}��Ѓo�[���	��t%?�0��A6�ZE���f�Y-�(Qj���}"�'0�'x2�'*f��%Ҁ=4��j�F��c�]JB]���I���Iuy��˽:>��U�~��ӎљ
Ш���LOK����?�����?���k��K��W?��Hbf��ԃ�㎎ah�u�gR���������~y��Bzx��?Ab&�'e�`�F� 0b��p�S�,���'�	ş`�'�f"�P>]�I�ϸ��s L>,P, � D�'����4�?a���?	���t��W?�	؟\��;>�$`R�jL�C����GI_/t.�9�O���<�@-���	�Ol���?!0F�V�WnR٨1@�CTx@�сs�J���OX�`��Ϧ��'lr�Ox��k$Ǳp�<��"ͭk\-x�#U���Iß`Q5K��I˟t�	Z�cr�C���e*L!i�-\+:�)�4s��Z��i`B�'f�OÖO�)�A��)"�ֺ~�V)�����mڥ)gzh��������h�m��W>���Nj�pił�%{J����ż�M��?�3�ཐ/O��I���# b��``�� =4���#��L�O�������./jQ�J�&I<���+�M�l�H���Gy��~��B�?���Xŀ��aQ�@5w�7��On@����ܟ��'v�C�P~D�!^�C��e� 6F��m�W�D�	����?)��?1��[(Z�$��G��l҄�V)g�4�ۈ�')��h����s"�_6S<�䒧�ϡ�6�������ڟ��?Y��?A���]}򊕘h�>��PbY�>@@%{�Oŧ�ē�?�/O��ŧ4��ʧ�?y�U��p	V�״ k�x���"2��F���O���ւ*� �O� s'��K|��*q,qi�#��I㟀�'` �bc(���O���Ƽ�#Lx�8ę��N�k�=`��x"Y�� #�ӟl'?=�'d�LJ�J�&`भ�7�$ �bL�'#"�U/y�R�'y��'��Z���07�n�S��N;�(x��P�<�`7��O���G�\��b?ɐw�1,�!0�=)8�ȉ'IxӚq3�P���IΟX�I�?��N<�'J݂���_�W't�SCڭN\4����i8H�'P��'R�O��s������+d�̴��h�
_����rΟ�&z0��'�ʼ�2y`0���b� _�ݙ��Fv"
���3W�lx)D������6e5'I�uJ��T�@����vo��2��9K���ŉ���м��g�)�OO/'L�+�䝱?)�l�숎,A��Q2C��Te��[�a���hS�_3<h�皿+� ��.�7������,�5y�#�y0�	�"�0��	ޟD�	ڟ`���ɟ��I�|��dЍ?Sp$���� p��#��\�d�ް��ݟ��%�Q�\�Bp��DV�N�X�f�JQm�����PXt1c��~\��bG@8n����Ǔ<�u�	��M�G�4<�M�0��<V���DbҼby���dZ^��yB�(���n�y_��"�y�b٪@"t2fa�<6��f��y��>9+O6HC�d���M�Iߟ��O�
p�CD�:e�MkƇܥps��▊B�2��'2��_�� �[C�24`�kT�K�$��O�jY��܁t�vi��� �lo�4Î�D�]���Yb
=�6c��;iT�'!NB���)X6ɂš�	@�HGy�a���?���䧡?9b�rV8�y��KL���r����?����9O0��6k@$^АYsV-<(S$`�'�O~]�)�|T��*�?q4�#�<ON�[�Mզ	�I��<�O�X5�'���'��d�Ȇ�d>�٥,�"����H�=�l H��{�^�ԧ��'��O� ����ԭ$ܜ�3�L3E>܃&K[)���:�/�&#��J�O?�H�$R *�q�x��5�	����i"��OZb�"~�	*hu�l�g��}<��,&C�5J��H�����1.}����v�2"<�$�)*G!OV=�+*�����K�<ivG�Q�|DK�G"J�����`�<1�HXc�ԑr2큞8����Y_�<��fW���������kB*��\�<���ڂ4�!�D�iB����D�W�<qfd9qH��R�P��=�F!�L�<��:�P�Gg��S���`��G�<a�G�J� XA@�^�^A����G�<�V$�8iF8u���GCT�`#$�]h�<�GOO?��< �J
�\V +��a�<1��ۀX� @:�.۴e������`�<�6�ҟLt�k#�
e��X`�r�<)DLK0[Q�=�qB�{�RdrQ��j�<�^XS �D-fuz����>u�h�ȓa���z�Ʈ+���	��&\lΡ��u^�d�S�ͧ>6� �Ӌ��~p��0_��*�Eǲe��p��]�5����%��F�3F,^�]¹�ȓ(��cE��,)����1�B':��ȓ'�
)Y�%ٯnL��PB�~$�ȓ�U`�.��<����8�"O�q�F/�X��)P�T�����"O,��Ӄ��F��I�&Ne��9��"O��â˘,<��waA�i����"O���"ۍ	��̉A'�XJ��h�"O �,E���i`�"5y(�i���y�aJ& �� ��`�3% �Cdc��y��W��ճ�>~��E��y�"ݏj2J��0ꋦfFN%�b���yr�'Z3ZQ�gƣfK�@rE �yr��3{�(�JT
�Z�����y��ɑ{�H�{��E�Q�=��ԙ�yg�0H��Òk6D�$��3a���yR�)H�HsS�^�5����w�ؓ�yBf��v<��V#L�`�lI��O�yRN�AK8�����Q=bܺ7mT��yBgR
$p�XQ�fF�P&��ö����y�eŖ�R��s`X-=�0Yj&�R�yi�J��4�P$Ω+'��K! �yb�&���(Z���Ӂ����y����mx�t�%�PC���F]��yH�8�84�-��ҽ��c��y�
�zx+�.�-?F��#f�y"jK8�x���	�2�y�֎�y���w\p�E-ājy
�Z�L� �y@^�6x���"�4��������y��ԑp���Q��%e�@�J�y2�W����-�T�\�3�kD:�yR�A�\}B��3M-�ݙ���y�e��	�g�I�H"���Pl���y��0V��)Qh��>ּ �"��yr���$N=A5ِ0Z:��r�K!�yB"�75P�ȴ��!�@4�2`�7�ybW�W3�u��n�R��R/��'F(SR�2S8ҽD��-�Lx�z���3*�����y�n�)��"� ������k5yl����B��	�]T�"|�'���"o�?�rq��A�  Te��'Ѹ���� �)�ȟ�����Q���uP�1�{��0�>�!���B�AYvIP��p=񷌀�Ж\P.F؟D����Ĉz%.�9-�����.(D�� \�0���<����@�F2
b�S���VD�b�Q��E)i.�}��l���(!$&����d��	XC�<�3��0h�F�"dI�Ϯi��g��~s��rc��򄞾%
>�snm"e�ܙYv�͛�`�Ʈ,�ȓ,Df����ވG��)@'� ���Bl�<L;�z��"��='I '2a�DÞ[I��FG�gX��9օ�`�)+>�� �C���&l�A�N&�y"�]00��ގf��<+�ֺ�HO�\ ����h�V�SR��C���3��B6ȣ�"O����y�~��K]�q��ȁP�iS"��%'�o�S��M����Tas"X�i^�qS��h�<�c&�!WlQ���ܼFx�D��Pv��}���i��Q���V`OR]QC�
��z��R� lOh\C�hI��J'�АRi���/С	A�(�B�Ԧ[%�Y)I��S
�.�$d+j��_�f�hDO)�~T�>QEB�_պ]���P�5�~�����'�j��	:S�t�� ���M�x��	�'�L���t�vT�0�x�\%Kp��$X<BsfW�N���	bӼ`@��Y�)I����^>�$���"�;&R�{Q��[؟8y�CO�P���+e�G�"`��Ytd���1�4P���	R ��Q�k� qf0 S�F�@��!ӷ�8��է'{�Y�S͹��0���QmQ�|x�o��y5Н�����A��ю�O^؈���{��8`��Kݺ�`앭��'�.��)7�J���<i��P�vi""N
j�0�NSW?i��X3Q�9RT#�95��Rs�H?��̙�:�L��ҩ��S���K��!�� �n��>}�Pڒ�&4���&,G:)..�!��b�~�#�DE�(Br����z?A��jZE�/�$wWP���A��s�:���"P�ADj���o_�_�����'=�m cL
(M",H�(�<V8�D:A-�8#L�@q� ʒD��b�gE�3TB�1�$G�"-J� ���E8M>����=h/�R�e�u�S�_v�'�݁���e�*IRb`@7|��d��0�Z�� �X9P^$���M�%�$7�E8kR
� �Iʋ=�XQϓ"���+D��.8���G�2��'�z��q�ɷ�Z�+��H�/��|�O>��צT�'
}f���wdT�1�N�)Uʠ�C�:�JB�ɎN�<L3b� ݢ�{��"q���`��cV�	��%�[?�1b_�&��t�)����g͌f�����:#`drc�x�<Q�I�D��E��;�޹��dE�!K�lٲH����72�I��D��[�)��p�Ç�	���1QF�_v쑆�	t�ʩ��Þ���f�Y�8��_2;w���*A�;6����+)4��S�ăC� U�X�p�O� )�	�{�Rizq�4�']��
���_�f!j�l���q�Z�!P M�j��2 ��l�MlZ+{�
�+R��s�h5*��֒g̾|�e�n#6�I`"O���)Ki�=���&����^�H�T�ɸ05�{B�P�"IV�R�z���K��G�>��(��v\��$F�D?PcW��@�CF@֚a9!�Jr=�=;�]}0)�Ta^:*ב�P�R-�^K�>�t@
9D<�ȅ�T�[�9�);D���sI*P�2�ҤӦi�j�r`�e�.hA�E��������چaD��suo�*-\x-��cV;�y�kM9^L���hrI��Ί���d�x�D��-+B!��F]�V�`	1���Y��u��I9G2n���'$n���@�2�0�aX/.'Θ�'
A�2dA�=y\��#-��r���2��䅩L y��	$?EjH(3�3I��PN�rg!� n2ܱ`�N��ꐓ_���]�{�LX�=E�ܴh�&�ց׌#s|`�%N՝*?�����كN�x_|���ޱ*��(�'<�|���'����׫wO�m�1D�c�����'L2ء��o�l���)��S�'Y�!ÑdP<�$����wm��y��Ip�%;�Q█b`��!�yҮ7�D���J9L� q;��,�y�\LLEZ���K*�pL�/�y�ĈA��rԩ��N@���f)�y�˶Jtd ��M;I��10#0�yR�H&B�&�)��>�^�4�y�]<�
��a��f9`���޳�y
� �(yta�Ml���L#l�m��"O@�ѲaB7AR��BCI]�¡�"O���7Μ7����+խ�t�2V"O�y�.�A3` ۖL���݋s"O,�����	(q�ņ�Ȍ9"OH}z�A����h+�� |�8��"O��`ή1���Y�d�Z� tP�"O�\۳��e̼P��@ج��A��"O��g!��9�RAW��� ��1�"O�����"bBh	�-�
u��a��"Of����� �/a�Nm�"O@d�ꚝm�H0ӥ䋸%z\h��"OVH	T��.'w���D �JF6�Q"ORܢQU�H� �H8���"Oh@��ү~�*%&�-!R���"O��W̋�,o6�Y�,��	d"Ol(�/��Z�tIժL�H�=��"O�ݓ�䔡O+\�D�� �$��y� �����[�6>.8(�KG�yR03��$*����'��[�	ޡ�y⢜�s�`*-���n�0Č,�y���xEK���J̘Ӧ���y"'��w�T���)�$����<�yr��*K�\�H�2i)"o�:�y�ʭN�*���<R)�L]&�y���m�R���>�P��h��y����_> �Y�V
�(чل�y��CKl$I4!�~���4�y<a�y�&�&8�9����y���'���QK(`����U��y"�޵��m����/h^�tٶh[��y�-�|�6�KW늓*�p��P&���yb���Q� ��-��R���'�y䆹-B�yӐ�M .r�(d԰�yG_+6����G��~9 
$�C��y���:c��NH>he���y�f��#�Ip�m�,����y�B��VMīW�C�f�aÀ���yR�$ֈ� K��;ʞD�RB�9�y�n	�ʬr���!=*�#�(_��y"�L�\�`�A�$�fU�D���y��
7(���BQ+{�zQ��:�y�H��[]����]��Xk�=�y�ǀ� ���P'[?$��� q�Q�y�C@+	�5��K-kMZ5�͟%�y2!����)��K�K~������y�&�JV���B]���q����yZP� �D��t!"T)���"C�Ɂb9��xS	G��ݣ�v�$C��64����Λm����s�f��C�I�R�rm{pN�W&��ifi�	<"C�	� �P@�g�D+1`ŋ4�{UC䉦P��С���DYn�?V;�C�	�x��I	6�� TI�u�P�~èC�	#Z��a�M�H7��� ǟ:z��C�f�E:�+�L�!I�_QC�C�	�r �L�`�X<�,(�C��7:82���@�.�F����6zC�I=X�hF@�*h��6�V�j{2C䉍`d怣PjJ�)����G�7^C�I�t�� b©F#�i%F�O��C�I���c��.����DY+ǂC䉋]
�bD�Ǧ[�~Io�3Sw���ȓdl]��&�<&�yg��6f�H��S�? �C�mH�B��{��q"OI��`T�2��Lp�"O�a�'�� �r�ل@�T�V�S$"O�����B��
E^� �"O��ឥ_A`a���P��<��"O�Q"_�M�!����:�&��"Oҩ	g��J�05�P/��h�"O�TU�ا$H�:���l�ĵ��"O�����о3��ſw�\D�"O8Ա�hK5�
�&��L����"O>:w�J�sXr�EɧcX-�"O���eoL�:Pes��Te�C�"O~X����!l�촩f��;F��g"Ot�+�N
�HRm ����Y80Xҗ"O�!�"�O*���sr�R,Na��"OݓTK�BT����˜ �A3�"O>��QKP;<4,��ᒖ�X�"Oh���ÒH/ ��P ��v<ͺ�"O΅X�A�s/.��#NJ�2H���"O�����a<r�,W�5��c"OH��䎣|�(�;�I��0Jh�"O2�j�,_<A�z00�G	cW��p"OH��e�9]ʄ��V��[4R ;�"O�(Ś�eV4�(�Ћ#�Ft��"O�t���*0VY��蕤ɘ �b"O(����҇nl>����X�b�T��"O��(û)|.\	�,��	�j0��"O��A�腰L{�D)UkQ�`�c�"Ol��*�3
��`�	E�T`��"O��SGB�ma��S�G%�U%"O`�X���KP@�����/0x��G"O���p�J�@��FB�]v�"O����dޥ7��ᅌW�ez
�@"OR�el��d`�X�ą(uU�t"O�逕杵t�Nl�"�6qY�s�"Ov��p��r�vpd.ƄlV�] �"Of5�O���}��.�9��"O�{���~�Tl�����q�"O��Wj�/4u8�B��b�K7"O����Ȫ��y�S�g����'"OI��U�n6&� �=u����s"O�)1�ω'A��I���^�0ؓ�"O��Y�d��]{��rn�	�`i�"OVt*�ˋ*�P�mW�Q
�� �"O�s񣃒b/�Ål��Sb�q�"O�����n���Q�LlAn�V"O E�udԞ~2ȀG�w"$D`�"O�����<q�xcDmXsx(�"O�01���6���d��lb�Cw"O�(�#�"e T�`oY7EX��r�"O^����ҖBRHre�I.�0h��"OL���8����E��tk^iKu"O&��Ƈp�m҃�
����"OЁ�p<]l�ԓG��f��9�"O�J� ԟ4��[A�"~ŔXA�"OV�Ar��=;�U��1W
�͋U"O�x�����r̆!���;Ljd��"O��e�	<���AAŸP��E��"O��ۺG���q���6�B�8d"O�$r@�ѻ^��`��Fz�
#"O$�"ed�-~��bD���d~��"OΈC��\ jnh�C'ׁ;��u��"O��V��(i:-��ƀ�|%���`"O��c��O/c��r��;j��Bw"O� *�j�E)��xDS**�ٓ"O�\k��30+�Z��W��h��"Ob ����
ir��Y�6���"O�P��g�*^<�D�=P�p� R"ON�і�߱LAZ�ȕ:\s��y�"O8}EK�U�M(Gk��"O>��6㝸'.�V��HS�H�"Oꀀ�kUM�ipb�rƝC""OX4��r���i�b�(NS�� 	�'�p�� �ʦJ�$Ո���:W[Ą)�'���[�ˎ���1�B�NU�Ir�'p,����_�hse�M�K��@*�'������Q\ ���сm�����'V�i�#�w/��0�L%̴���'bd�aĝ�c�R����Ŏ �U�
�'_�4Yf�o ޥ����.%�e��'���nT�*f`( �� sJ��;�'�aᦩ�� fm���d�✈�'Vt����);�j�H�%����'M�U��a�'.���&iS��4)��'E�H�GHh�q��J���6Eh�'�@s5�ҿ%� ��&N�uZ����'���$�	BJ5Q�h�'�l��'�1c��;�i�V��Cn�ӓ��'��(7C�0:�jٸe�6\!Y
�'�.9�F�,Np���&���P�'�h$�a$CFl�l�7J]�u��(��'���	���$>�B$��,>����	�'������`���N_�NXy�	�'w쐰S�BBԀ��o�.����O�왕��`�$_'uFn���"O��qR́1=.�84dY�\��z�"O��K%5Dv<�EH���� R"O �B���?<ÄHH���v3�=�4"O����$ޮ
�	���Iq24�#�"O�T���S;?��E[ŀM/w0�l�d"O��h�� ������4J�J�"O����<F��ER���]f��"O��u)�%!vq)��F����!"OJ 4HܕC��@(4/H/I�@%��"O8h�6�׉0�(�0�N��y���� "O���΄�N�{f$��B�XX�b"Oި` �u3<pCp�F
�0�a#"O.X�U��(͈�`?
h2���>A
�CPbE��f���e�F��A�r݆ȓ07r�A�)�]���Y�*�	�"\�ȓ'�����	p�)�MJW�V|�ȓ=��uaU��t�#��9��1��;k��GE��H�\���x^Ty��b��Rf��(��u�k`~���7@�,Sd[7������?t��(��P;!a �ǚU�.yDÔ�BF�� ������)���ĉ�t��WRv@gŃ��d{BeQ�'�-�ȓb�KE@���֪q_���y�@�NΈ�!���S�`h���Í�y��ʠ<�
�p�J�A�4����y�F�:/�^\h�ئ©@K/�y��Z�{����@j�|l���yb' N�E��{Ҕ����:�PyR�	&S���R�dn�pƧ\A�<I����!0��?g���XƊt�<�P�L01E��xR��V�����Hr�<i���+��r�KQ�{Zn�"�h�m�<� Zu��� m|�5�ԃ$3��\(�"O��G�� ��]���4^��=��"OM��*K<
x��aU�S�Tq�s"O��C�.(�V�Q�+�����"O���E�z��x!`Ȉ1�t��"OH`
��us��3��tm�� 5"Oqj%Jڛt�l�)�*R�{:�䣧"O�]yw'�":!�\d��/.Yb}�"O�2�->dz�i�4b�l�"OHY7 }�Rm`i�"�����"O�0RG\�Y Z͐�CBJ�m��"O��؅V�yr �r�8;+ᚒ"O<��`]M��` ݫ%^� "O��s6AS ���r��	:�1"O1�E(ѐ�2��$d4��s�"O*��3(ڒ^�B�x��q��_��y¥���L����i|�P�͉�y2
 f�%� ��X�$s�� �yD��(�
pxą
:�X��Y��yR	��*��p
�c[�	�<���yR�)8��1T���+�0%Z�,E�y�(S.ϤdP�'O<veH����]�yb���B ��8�ɀ+qh�� ����yR&U�a�p,˷�͸Ln\/�y�.֎K��b�h1Nؠ#tmԳ�y�."�u��'T�!E�a��5�y�B �QE0��Ą1!��@�;�yBkL<"Җy��F�rT��G���y��Z']���2)����#���y���)���󀀿�D�(�n֝�y�E�J��i�������Y�y� б��(�uC�$�Duy��	��yr���D-a��єLz�ݲ�#(�y�JɎH^,\X!��<��<+����y�EN�3��/Q�-:������4�y��1����dF�3$�}1�<�y�(�]�0�j͡`Z�H35�I �y��)K��U��,Yb�b���y���b�˴��O"�ġ���1�y�	�3C����Ą�J�%�R�Ȱ�y�+�A�<�����::��)ǀ�
�y��̝i�̜�&U�H�����\��y���B��QR���o�؉X E���ybŉ'�
���� 'dĺP����yr��6¼�뇁עW�V(H�a��y"C7By���q��6Y��uK��Ņ�y�S�7�V`Y��A�LISw@I?�y���@1��ȁ�69�	P�HT2�y����Ґ{�eL�vE�?�y"K�_��Y�CK���rqp ����y��S;�~�Pte��w���2�-�
�y��YO���k��R�D� ��&O��yr��{߈  �nR2;?��)����y�Vj��Y�k�3����mĤ�yr`]�a�4��< t 2��y��E�$$�w`�&���I�yҥ	.\�����z�tT���yi�@�S!L��'uܝ��F��yREس�p:JV����I���y2B�m����'�4���$���yr��0/ �{O�j-�8#��9�y" �!n�Q�I�*hT��!��R�y��|����,�M��DjX��y��f
�۳�O�O|�وt� >�y
� ���3'���i�&Zt�$ v"O�m;E`�0g���P�=:��("�"O4�*��d�^���ăRS
�E"OD<�.��8��a�Lt0��T�<AЎD(~.Ź�3@ ��
�Q�<qdnթ�!z0H
/W!������V�<qR�;P����l�g�<A4(G6n�|c�Gӓ�j�u��l�<q%hș��-��ܦ��EQ�Qs�<a�K�Eh��Z�&��k"����W�<����Q�a��D
Q�1d��J�<��c7ms:�K$�("�,1B�JE�<1�"J9*q��j�#(&B�H�l�G�<���6D�48�vjRIܒ���#NF�<a�N��Lsd�H���:h`pQ+��<iE�b���a�lN��K�b�f�<��n��D~Z�(��ŵR�"��A�a�<��-q7&a�DW�d����g�w�<���U�j��B�6�4��F�h�<aT,�W���q�E��5����y�<y��Vn|JE@$iȹj�V����x�<a�-Q?=��k�B�?�,)�d�w�<����(؆���*X<1%N\��l�<I��FTn�XzdJ�8�l�p�@@�<I��Z�JlXI^�b�p�}�<���K/B
�yF�M�,^�u�uÝO�<A�ɛ�LXūQAlJv}�7JXJ�<Y�#j��RPpC��A��G�<ARaD�lQV�!aT�M&�t"�`HE�<�b蓘o\D�+��T��"�&�C�<��[=gˈ�儒35>�f�x�<Y���>*�q�c�':�{�ii�<�tǖ�{(�h;���A���ӭ b�<�6 
 T��@������@m�a�<�4�ɱX����2DԐzf/a�<�.���i���ܞ:d��PG�[�<�᥈>�V�Dg�0���7/�\�<Ia��=;�����\T	��0�(�|�<��֥^)�R��$�؀��Oy�<y#�^*z���d��D88PT��u�<Yuf�8 "l i����$0x��G�<9���n��A�J�8`���^�<�r���=<6�@�B�6d�	�mFW�<Y��-7����˻`�ʉ��]O�<!�� 0Q�U��M�8;f��b��L�<)&$�=�z�ۇ�*u2^4c`#LF�<i�B�q����-K��D äh�D�<i����7g�x�%,׉_����G@�<���۶/Ct��B́�ZQ�Q�7�GW�<	�L*k��m�F/�e��)P�T�<��ӎ�v�aq���Ƭq �v�<!��N�=�����79Φl�.J�<Y�)1����[�y��!QWH�<Q�LG�pM�q�(D�N�_�<��C��J�L�9cNˢ)<����r�<RMF�w������Z�Z��W��r�<�pkE����Lː�BDڥ�Z�<Y6� �<_�����=J�u ��YT�<A�,�� ��P��@Z!"�����eR{�<�!!�`�D��S!�r�<l�d��y�<�ҍ�_r�6��z�ިAF�a�<��l�u�ș�-ōM�E��O�h�<��쐾o=�4� H���S	�M�<�d�6*��H1셅�,�̈́`�<� 0L���ЗZ5��C@C8$�h��"Ou��D��T� ����4��Æ�^�<၌�J�nq`UG�>����_�<A���Ŵ�b �Đ<�*(e�W�<���	z�Yr�-�5h1��h�V�<q再/0P5�G�	X�4q�3��g�<���AϤ����Y��т�f�c�<�q-@�J9{Po��7�����k�<�4/�<CJ�A�a[�n�X���&�g�<����w�nI�CO�IL�*W,	L�<�$KB,H@�D�]4'U��Ba�<Ƀ��97jʰ`%ШTl�B,_H�<�����d��x��$��1��Yy�<)wh)0z�4����	B!ڴ	�)�o�<!r�[c�mR�K�;�ai�"�S�<�2(S%L�KӮ2��w��V�<V�ͫq �)@�N�d�����CH�<ye$Rx�Uk��
8 Z�Hd*Y�<A
oa�/��q����T�A�$q���{ȴ�I�$ˎ���KV�X�n�.M��iֵ𐄐�GJ��7��5U���ȓS;M���I�lTL;��� �:���-�T�PR!;n?����l,K<�,�ȓ\��=IR�^$sF��Wj��LVL�� ��(R戠��q"Š5�q��J\�ej2-�:d��OɁ	�ԇȓjr�(r�%�=�Z򇋇{�H�ȓD��l	�B�0>�ة��L���NL����u�Ѕ�G�, <�������q�R'4� 1	ƫU+0t�-��"�8 ��)9 �u�!��Eb�'>�@��F�S�H��Q@I^|���
�'���Jʝ~�
 a��?hFp`�'P�E�1%�7.F�[�œ9�E�'D6��ec�?\
����K�)�����'!.!j��]'M��Mۧ5
Vp�
�'�(��ѫ� 3�> a4��=6``a
�'��;���}(���ˌDy�ٸ	�'fn�	�&�y"8�JQ+�>�ʘ�	�'3��"��4d\H����ȓP%�-JBER�E���rGE@����]�R�b�"K"�\س�ļM�,܆ȓ"q���Ð(8�u�V��!1�e�ȓ{��u�����T����H氅�}�����żrt��B7>������d�Έ�j�i��]'Fn�ȓd����KN�����iZ�]sH��+��B�,b�@���8���ȓL�@��#!�b0���7h<���\y���A4�����2g@HI��#]��#ϗ.�8��A�(bx���}�����!�9;�%��F��m�H	�ȓ/�ZlRT�ѲZz���C�?���ȓSV`�q�%B�aԈ��EJN�%j��Fh��O���'�P,<��]�ȓ�ؔK��4�D�ӕ�̦|Z�Ԅ��j)�a���	��i�"���h|M���Ԓ!W~A�1��Z�@`�ȓ�(�Yb����T��ȷ_�t`�����cG*G])�C޻E�@8�ȓR(pP]y��(cQT�2ئ$��"O �Ic�I�e�Mh�!�!M�ʹ�f"Oذ�6W�����֋3{�d��\�<A�KJ�3�hi@(�]���J���B�<� n�#e�J#:�^ �i�w��5q�"O��I�`.���w����䐓"O1�m\�cޢ�1'_1d��dQ%"O�Lk�'�59:45jwK@m�"O2����r$���f�� f�h`�"O�9)rN�c�(�:p� {ʥ��"O�a�!�4��šp%�"+`���"Ob��C��Xa���s�7�b���'�(��!�5�Xa`0%T+�J���'��e���#�x�K�Qh���'��+�`�i��2ք��'�|��ubZvA�tX��A!��\��'�`["��xt��D	�ܚ��'f,�ch�7@m�V�(�bT��+��= ��G'H�mA4�	�ȓz�����-ѷ9\2���&����|��@a��>-Tj��w(���i���CX1�Z@��o��@���ȓB="M�s�'&$��`&$�%����ȓI{�@���$�]PC��ä���%��"lڽ1���Ɔ�P^Շȓ,�1!g"̺[�&h� �"O��ȓ>R��W��$r�BA���%#�4H��!�8Ê:v�@��Ս^Ϯ�ȓ2É�Z^��Wg5��a��v,�!!�u��v&�>:��ȓ@����P�ȕ:�~�2��G:p#̵��*�Z`{���W�$��+�4z�"��r���Ru`Fk[xDBh9=�Їȓ3�R4�FBǺ�E��gӴc��̇� 1������7R�5lU%F0���l��̰��@$�"��$`�����oQ�q�d����!uE������D�d����l�j��3 �3e�LՅȓ�2P�u`�	t�|9�)̭iKȘ�ȓ �<�d�^������,(>���e�s�+�1S�Xq�C�)�Ć�QX�Qr�7S��0�B��B����ȓfR �f�W-3ޘ 1�T�=��ԄȓpŊ�0���Z� ��<l��̄ȓh��<XB�5�]2�H�Y9��ȓ,r*i�ghly��] 1�,d���� X�>pH���ǿT������{�,$"!ZR��;/�r=�ȓ��0�K�^�NL3�(ǾM�p��ȓ+_�����i�t��a\?|�m�����B��P�pd:� ��v��نȓ"_�u#��Q�F��\�;�R��	v�������.���� �L]d4�-�;D�}��<D�p�H�eR]B��K';	8�q��/D�P����'ZR�����\7I0����+D�4R���xpnEX�+V�m�9��)$D�D�򢔀4t�
�\� Ai4-/D�lc��LE.��fO^�3�����,D�`�V$'pd+��9,E��Q�?D��D,P�
�ɫ6B*
t� C#c?D���獢1�mф�@,^����<D� �4C�/6��� C߽#�:���9D����LØ2��g&_FP��+D�d�0%��O"�Q�°$�N��D*D����U+&�@�+�ø+D�z�h2D��@!#E	\��9h����D��i�O@�=E���&&K�0�B)��\4�e�R�,n!���[��z#� �y�Æ!;P!�� ��Y�~�<uǚ4pY^��"OtX�V��
7ܞ�a�����"OE(҆�-��Q���ļF}JT�e"O��#�R�3�n�"6|��
�"O�H8�����Xx�MHSqfi[��d�O���Oj�;w��J���HE
^�*��)��'�f���o��'R�;Uo��z���'���vNȝM�f`�A�ϝw>l�B�'��ҍ�~@����}'���'��ybEAV�0���*�v�r��'l�lR���<E<��۠=F�8�'�l1���I���H�� ȄʓB���`u��u�fZ2)�A��ȓ� )�S_ N?2(��н]�bH�ȓ.��-��
Y�*�hѓ"U�I��`��w)��
'.ƕDڬ	�#��}�X\��e��c��ͣ~�$|pփ�)C�����!��!�Q�ld8�b�*H��'����ԔȠ�ϔr< ��"�4؉�EK�"�I��T�Q�Xi��:��o��8�ұ$%�@���v��%�@�L�~�J�z�W5�F���G�Z8�ǩ��_r�
҅	'o�9�ȓy�ع��,q��)�ACT�Н��FN^��$����Kw'�G�ńȓzLnMI���-+���E�T�9�*��ȓ+/ u+A�L�_�̱�MƎ%,B��(�����#ƫLR�1�JF
6�0y�ȓh�ɒCU�3��pѠcɜt|d�ȓ-���!��T�P:|�6��(��`�ȓ����݊a�RZ�KYT�d��ȓ5�d*D�H^d��ɲ�#F�rp��/��Mң���X,yA�X�F�h��!���Gɋ&r@��x!"\08a*Y��af������<Ft�H�c�*nN��ȓR���E�4%Cf ���>K�4���3&hy���	�c���ӀO�;gH���ȓo�X�9S�БOs���զ�7s�4�ȓ�*PbG���OCL ��O�/O�>��[8���5�b ���.t�61�ȓ?N8=�P�S4(�ڔ)���&)� ��-�09�`/R�Zd��OH�Rt�Ȅȓ3�P�Q�`��n[�$r4GҊw��l��V͖�9���%(�pm�.R@���ȓ�(���۳_fB�i�CX�ZR���i�����טPÎU��<�Ե��/֩�Vb��6e԰i2jF�%���,��+0'�'wV&��t��P �8�� >%9��ɿ/�0��M��5�ȓT8��r��';��p���cq�]���r\�`�_1I@H��I܁p��ȓCӰ��rLI;F*�s�&A?yVv=�ȓ�⭃�K%P�Fh3H��(�ȓC�|��$��!h�-��dQoR�!�?9���0|
֠R	3����G.!�H!���d�<����K� x�4Ę�r�DXaHa�<��	1o�4	1�b��*�[�<I�쎀e8�m�T"D�F^bh�L�<1A@�1)����#u���(7�P�<y�*�^������S�
�8��[W�<i����>�|��X�u������m�<��%\�J!�Th�"��� ����g�<��ģ,�, ��l�	2@ +w�]e�<�Ύ�kT�(F�ֶW����BCEd�<� ���ĕ!%@�h��J�q"O pAPf�o�J��P�!s��0��"O�ݻQ	�e����m�x�c"O2P�[6~-6��cϜ-O�� x��$�O���IB�+�
� ƕ�v� �X�aȋqў���I�+(6Qi�E	�:ؙ�l­w]B�IX�D�KEN̋} ��P�E�1"2C�	�K\1�rO��hXN���l�<47C�ɪEEr8�ǃҋq�,* �R�B�ɷ^k���$K*d���J_����$h�P��f�.1 4��$D�)�t��'&)D�(�f=R�|��%��g�(�4n(D���t�:WF,�aw.^�
$�(�E!"D���r�TyG��`�%юyK~@h�B>D��	h����Q5R��K D��2�J/��aJ�P.t�t��g�0D��!�I7s��PǪ1Kz��/.4�x��Z3(�$��9	�����ψ|y��'��83�.i��a�FĔD�FHH>I�
tC�O�z�V�ZP�òY��X�ȓjɖ��p�O�D�4-Rd̗�~ނD���"�z���vp!:A�"Fв$��AIEK��kr�ꏢG�Ω�ȓO�f����?����MJ�!-�=�ȓB���)Q�+B�Eт�	�hh��7<�h��C�>���!$��bٕ'�a~b J(�4�^�����%�K��yb�E�'����,�X��� �!Ƅ�y��FD\q�߃}z�A�'�5�y��Υ���G�6f�\]b#�'�y2�~n��;)U2�� R��5��x�V?z�� �#Z$�("F�V w!򤚧zh`a[�j�-%V�E��MS!�$O"S���e�*h��%`TJZ?!򄞂<6{���8}N��FI>X%!�E�m��L+�  �(�V����A�!�d�-!`T��V�=/ڬ�1��
�!�dD�l2�����X-�\J��n�!�Ę<Z��}����;��S@����!�H�xX��)'�_^*�k�B]>�'a|�!�2�	�B���ta���C�y��firAk�,Y4��`V�3A�����2U���ȈDp��#��2<(�%�ȓV �@e|o2e�b�+NZ����}K����:b0�;���*"݆�Bs��2�2�b���lI?��5E{2�'}Hq���"ŜQB�&ɶ&錐i
�'�r�Y��u9�	Bo�H@��	�'h@�5��7\��A2��F_��I�'�6������^)80�7C�<KHb)a�'�L�G�Cz���V�š7���P�'$b��ˋ*k�"!3����0�ȓ�(���̔�_���Pk@�6!�M���g~"�E0��]����8G2\������y�#��^dɁ�P�A��qS�;�y2���J5(i�H�#���y��č�y2ⓞ)V��3��Уl}̵{D���y���g�\��]�9�S�^�y2�L90���YS��]�b�s�I�!�y� P�f��$IfU�0�7�y��2n$f��*	�����ꘕ�y��N�4U^����*����V�y�e
)W��!*2+$�L
w��5�y2�K$Fh��R�#'�𐖠��y
� <�i�f	�����S��}�"O�ʅ�^\Y ��BjR��ܸ��"Of�1GO��V3*�0G��-t+����"O����l١�(H��Z��"O<āGA�$Қd��C�h��"O�=0�G�x��A�U�Ț��Q�"O�l9��'E��P��n�L��졤"O6�I��);�O�	ƌ��"Oz�ە@O薌I mηP���E"O&H	�
<u� =�a��$4�؁y�"OL��u��>�n
����HC�'��Q��Y�lA&C#�T�C�'����	�+�<h� �ن�p�J�'8�"V��',|���k��?�Y��'�p�iVn��3#�U��c�;}@�r�'�$���ʠDSB,3��i{	�'jN�̏-;9��0�mK((qx$q(O��OZ�}��0�����,h�V	�0�
� �vm��~R>�C�֘[�n��%�E�5��i�ȓ��WH 5���x��4 7 L�ȓb�p�kaF�W~�`A�%6�ؠ�ȓ^�zYi�P�.��$��F9W߈X�ȓ�r�t��Q}¬�U���ȓ@�D��'�S&4�TMIV�ͅy�����|����z��# �|�@IAL�
�<�3�8D�0C�;>�:���� 3LLu"��!D��R��%CW�y�aO�"g��)�&%D���F 9ig����М�,u"��?D�\���ڷF��PY�G�%n�b99+?D�dK��!`�S�MO�3�P�<��Vy��58fFE�2�ҒUݲ���(	�˓���h��d����%�ʎvevP���K3�!�&!�T�� ���Qba괧�&�!���K�>�[�ށ�l�b��R�!򄖉}vޠU�3>�p 
�e�2k�!��R����d-N�5δ��E_:Kp!�$�q'.��E��� �T<c%�H~4�O����|
�O7�H�gl����Okux1�	�'*H|� Ɛ�j(�%�>s��A"
�'8�q�������T���d����	�'qt��e�\�N��Q���Z	�'�������z�3�o P���'�
D+���Xn�a�PH�y��er�'14��G�^;\N��w�FgD��[��'����|:P���<AހI��>'#�0�t�YV�<���4f��kd˼Q��¡)�{�<����96pMb'�ܶ�J��db�a�<��c�gb��(1-b���֍a�<���
�%� �It�S�|{�$Z���E�<���I�Lø�1��V!:�)��\�<a��^+Y��W�&XZ�Ы���X����$2�
S4�'	�*IwA�A)�v����L�H9���ߍ~Tb��v�4I����족�˙',�e��/Hz�u�ȓiU*y����P�b��,��v;Q$/r�A+�.5Qsv��v�`-�2L��1xz��f��<{j	�ȓPa�� @�	<؂�
f/5Hp6��wwr��-� �N�ʑ�J Dx��	{~r/��FF��.֬z�b,�Eg���y��� *)R�["Z�m�}�u��yb�޻#�L5���ߢ<�"���Ԅ�y�h�)��X9 �K	0�@ѣ�T��y�@�L���K+��<��^��y
� T���D]D=�� �r��D"O�r���:R
�q�N�O�8EQ'�P���pO״�8��ݫZVP(U�"D���#@�=5"��P�`	t�*��Ӌ%D���3�I�yn���#�9v�u�1D��x��ޑO� |�F�\�Wn$��e�;D�Xx���'_[�y�CN�q��AIt�.D�,y��L+XB=#�M־�� pv�,D�p�ć&-������T��`�!+D�|�W�S�(��,�rL�+�\\AF*6D��`�D.\��4��H��I���a�9D�\I@e	�B��z5��n��D`F�7D�<R�n]4䜌���D �Ԍ��+D��R����d2Pܨ���#�b��7 &D�䨆�E_E���~R��ĥ$D�XQ�
Y�V�l���I����O�OC��<^�:PR4k�*�@�
\abLʓ�?��_�l�i��J�6�bF�J6s�����;-Dp �kL<6H@�鰦P3v[��ȓ`�|%�E/\���m-X��9�ȓ~��ɢ��Fa�LA ��"\�Ru��%5�łBJ�V<�F(	H�.5�Ɠ|6L��*��n$BD��z9�X�-O���΄k̥��&,�)��r���d��@��g�P��m�4�PCY��j>D��0j��m��p�Z�~�t��i<D��ئM�q�H��$��`)ҥ��.D�� Eǫb�\�.�!�E��c&D�)3Ï7�tA9��x���P�P����
|�i�E� ��`Ѝ��/�B��ȓlt��ࡗ0Wit$z���>K����?����hY ��>ju���|�x��ȓD�t� �N����(c���P��Մȓ%�x��$Vy�4¤h[�e~ƀ��ON��s��ܿ4���)ѦC���d��9\*E� b͌Z�,�	�G�*3$���;2Hy���Ѻ>�lX8�m�K��<�ȓb��h�F�!M�`��fL;I$^��ȓ�T8��M�NV�����P�x,Ԑ�ȓ���b��8��t#S�l\|(��nވ�G*��.���#!S�i��V�qr
ز�L�@�&�n��ȓw��!��C�":瘈�g�U	��ȓ&6����� Z���t��+���2A̽����%�p���<s��J0,`#  W.:� ���$ȦspD��tY��"<�&����8t4��)Z�L�����35���k*l�&u��8bPia(߂?1�ET�/���ȓ)�]Y��CQ��bǂ�@�f��ȓ-ty���¶ckZeK�(6X�l��B-�A�R�Ń} ��f�浆�b�����V�zAƠ��(��9����P�c!�( �<�p�®E����!����J��~R�*E��O5��ȓ?��bQ�ԌZ�푫l}�	��=D�d�"יTg���O<n㸑�Ԇ<D�Tz�G���1:��M#<�X� D�� �J�U�݊0e^�{�6���@3D����НK����U^4,�;D��zTĐ�?�y��[M]���p�<D����fG,F�i���x���:D����@_ �4�����<���,D�T���̃ ��R2*S�z�����'D�� \5b�gZ,��H�!��W��X&"O��jq��kײx	Ȍ<�Eb"O��aW�؈��\
'���`E!�"O���`�kE�Ih�+��f�ni�"O0��&H���B8�d��H�@T�%"O�Y*gؗA_N�[��#q�(��"O��b� �1��3��;����"Oʽkw���4R�J� �F&�"O�M�f��bӾ���	=$#f�:�"O"�A�38�С��)��0����"O =�W@!~)�acwȌ0Q��
�"O  �e�.|�LqP�G�n}ހ�"OĜ�p�[�&���K�M��ڜe"O�`Q�i���R޶	up"Ol��7�H>4��D��ܦP��qxV*O,h����n�ؓBX�[����'K�0P�� �% 2J�K�^)0�3
�'�!���:��@�$O�L���A�'�\EH����x@ C���{��a�'�=�7ˇ5�V�*7�ԅ!E��'��h�ӧ�1A�����o��ɒ8�
�'��0��K8��pHV��&Җ��'�fi��8pB��u�N���9��'Uz����+&�����c<�����'��l+���g`�(Ί�}�`�
�'�� 1K�洂�'� z�j��''�<�vn� l���e
V�>��9#�',�Q5鏕KA�c�[�3��l{�'�r�YG��N���k�ȇ0��
�'�M�$c��7]�(��7��i;
�'ؚ�P�ٌ
z���Bҿ�0y��'b.U`���@���N&u�K�'�r��a�Q�n!�E�į@$���"O�� ��Hq��d AP�F��""O�@�ZR`��8��Im�� r"O�p���E�f�z���N9vɠqx6"O��؃E�Dj"u�U�����"O���GcX��u��&؀|�����"O��0���!�Ba�䐫+|x�!�"O�����Py����7�E�x�FY�W"OV����x)�!�!{��[�"O���W���-� ��0����@I0"O�,��*ޭ*�)�Yp���"Or�Av�?�8��l�-�j��"O���/F�e����V',���.�!��	��hc��.h �� �ϑ?2�!���FC��"�Nꄝ�A��~!�D��tE�,ƥ�;u��aVMV0,i!�d!ݴ�ㄨ~�$�� ��vq!�$a�l%�foR$a���c#$�>5!�Ę�@�\�� �S�>��DIO��!�$B�pU0���g�rYR�']4B�!��-
�x���k���AL�4�!�$2X7����ÓXʰ]��do�!�DF�tT�"��\R��p䋋!�$Q's3�!�hY�RV"�#��Ppg!�C� _�yjflN��񁓠S�-Z!�$~�"H6K�8I'V�!v���A!���0t�z��-�>'�U�r�Z�9'!��DQ��e�G!2�~$8���!�ė�5;A�#�a����!t�!�d^��R��J�NҀ�U��'�!�7k�
1���N�Y�amG�r�!�	��&�9�L�m+������!�� ����APT�,b"D�ar��S"O\�
w��=+ؼ�@@Ǥ8�Y��"O
T�d*�3L��9Ơ�[o�	�'"OP]�q�Yw�l�UF�u˄b�"O&��3 �<�ly+�D�_��P%"O�)��,� C����PW�Yl*ȑF"Ob���")4G��;��zb�"Ol��r	[^u�À]|�: a�"O�ڠ� �{v���Z�{���"O�p�q���������C�"OL��Z3�RܪԢS�Hֈh�"O"����2����'�b*P�� "O�*Q�.w�DY��f�.I�=�"O�{�䁚0A�2�f4<кm "O��be\�4��kA��:�N��$"O�E�C\Khp��@��z�n�g"OI�'�\"��q�" �p�r��"O�<"����5H���-���H%"OPdud��
$�Qɀ�˵>�j4I�"O �3�HЬO1t�a��1m`NT��"O8`ꡈZ,0G
(e�$S.�(�"O�𑬁J�t!oD�"CP��A"O�qREʴc/0�nV���.!�dг<U�eB���F�b�͌�Ar!��4�L��É&�R�X2J	�4t!�dP������#�l�&�"?n!��Û:�:� Њ��z���ɶG�!�ʶ#������9�Nݪ��W�J�!�d+�J, �dG�?�����9�!�dڍ]������#5�I�|ќC�I"�����ŉg�Z�A�41ΞC�ɽ"H���i�-PFDxD,��yP�C�<T���c!�̀<�D Z��̨u8JB�I;x?�Y�K�;m���g�~} B�I%d�x��_9Y�������,B�ɯ�ua��	y��qXE䋳R��C�	U��M���LI]�1�E�՚5�C䉪wU�x�&�M�	%�� �m�(#M�B�	8�t�5(F��X-]P�B�L��K��	.Ek�y
���9d��B�F4�	F�42|��1�jB��,th���z����^�KDB�I\��T�h {��ȆB�I�lݪ�+�-�(b�.�B�C�>��C�	+-�ʩ�Ն�d��8�PkT|��C�ɚ4!����P������L�<B�#E�Q�%]�NR�q"a�1o�B�	�^�HC3������Y�W�p�
�'"���[b��h�こ�L�RU�
�'�6b�![�?��`c�o�(}`
�'�ؐ�tgY�`R��˂�:gI��'��R$�=,���Ɨ4:����'�H���Δ_����"Õ%g}1
�'.l�3BƆ�.�v���l�P�*P3	�'b%�aR�y��i@>'�1��'y���sD4)aLa��QQ0pZ
�'U��R��6c������)�'����4�_�.F�asA��-@{�y�'�����RA]�0��j�6�P�J�'<����X?m���uHU�𲈘�'s<��_�$�z�c�
(��'6j�X���	��d��|�~��'��I�C$[�j I4�;?��k	�'��mȤK]?D|8�� &������� $�F�&� ����p7���c"Ox���|C�\�#�Z p��e"O���1NO�,L��Џ!���"O6D"�ƿw"�A�t`��-�!�s"O�ڰ��IPB�ޤR�`hw���yB�<����i�}��|��K�y zIr��D�ܼy�A+�䓶�y2��bY�!������F,�y�'�<.R��ˑa�,
�R%*����y����d��P��4�����G܁�y"j,1���6��*2�2����ԅ�yR(@6�^��d΋�3:�ٻ��O2�y�H�sP($jsl�#�2���e�yr��/{ )����!v�8�a&X��y�K��N�LMP�΂��	8dJ��y���0:�u�P�E,	o@�ϙ�y���6��2��(w]`Px�R�yR�&����Իpx	��!�y����1�Jv����1���y���y�v�9P/	��\<2�*�3�y�c��x�0�D�ا'��p������y  n��p�SZ#:�$��	R��y�D�&<��qɇ`
�P�V��)�y2.5�ś�G���h�㛵�y���,&"X���ҹK�-ڤ��yb+M�e�j��emw�ޥT�� �y2��rȤq" D4m��v�R6�yƃ�?��8���7���p$�y@�sV ɷ�"6���qť��y��]�v� �!����3���;�F�2�y����m� O����ˤ���yr��i����)
#*�&�Db_6�y�
J53�̸�b�&4����ȅ�y�Mߖ2�L���Z'O��9��]>�y"fX!¡��Τ��Ȣ��yrK��IZIzw�:��l�bJ��yn�@�I`��{�l	�c��y"kC�	a����\VU�vJR��yb�%AY���3N�조ࠋ��y)$���I�<�������yb�D )Լ���������#�yb�u�ƅ�'pq��E�y®�6�tzt�+��� ���y�$A��Y��I�|t�u��bX#�y�d�2 �R�FP�pN��xv%�1�yb�V�o�h�&�e��� K�y¨J��ġ�N?aI�]pS��yR�;A45�J�.��H��E��yB#�u�xpG��[` {�n�"�y�3a�:AY�C��y&�)�	�y��ߖ5����&a�����SsϚ�Py�
�T�#���J?@Z�ώV�<A�Cӊ_Ȩ���<�l�f S�<Aw*�'��C�B
_�i�T�GZ�<��	+,���xRe�2[�j帆��n�<1�Dk�V���o�+���`&Âi�<����*������'t%�� ���N�<�P�^z 4j�l��>?"ٳ�L�L�<y$��H33�Ě
K��1G�@�<�s�ɻBa�3հ!G���%�Js�<1C` 3>&@Bb�ߑg�ج��Gt�<9dKI2)�B	���P������m�<��ǌ=ҡ���D���ف�h�<aD$���B��Q;y�L9�&Qe�<� L�3��֢R���%Η�
IDE؅"O�m8p�N�<8��l��@��Q�"O��2U"Ѥ	|�ja&�T�~��c"O�򓇙�Im|b��w� "O��V��˄�0t*_2|�*��"O9��m��ZEkħF��"O�8�6�ƷJc$���L�D�N�	�"O���E�^jr��&�L��,+!"O��sՎ�q�܄(c �[�N�0�"OZQ��iT�����l�
�zW"O�-Y��9
�&IU��'Q��8�u"O� �Ů�d�[���2ܼ*�"OR��d+ݐ-R�ݲ�o��e�r%��"O��	e�׆\�Pq�`E�-�j�:D"O����e��d�t�p��Ђd2P=�2"O�ZW�P[�j�H�)S�Z.1H#"O���2혇�XE9Ї������"O ����F.���>T�N�yt"Or 9BOS�7�H �D�gODm��"OB4!�F�ґ��B8`>ʹ�s"O�X1�Ŏ�$� �JD��|�`B"O�1�U����f	�:R�`�G"O$�[pkȕFLFHq� 9��5"O���e-�M�,�zfCH�K�8�"O�]a��D/j���DN�+�dՉp"O.���
c��#�⚣2|nثS"Oh��pG,<���7Bd؆7�&D���G�V
��Z�LX���ŉ&D�h�ǧ�P��rT��G�\5�N#D�pQ¢�J�� � ���i�$"D��)�$�2,��9A��M\Ҵj!D��uj�*��؃�ɑ�jH�V�)D��&��>64�HD�.;ht	f�,D��ą6Kn킓�ěl��H7�)D���L��Ҡ��3-X^���!D�@ e߇��Baf�
I���0( D��Q��A�<�+�j�9�q��+D���.R�}ɲ�Q�
H��|�6"$D����9��׀�8W����*"D��ba��+�M���8D�|b'�-D�ԑGc�H�h�X4�7V�q��-D���sR9v��ԁ�`Q*kV�ԈS`*D��P���	X�5�'P4
z��J0&+D���#!Wy؞H�!�_j���'D�8	Aa� E����HL� �P��&�&D���gBf=�P+�.��%������0D�@�w/�>O�a��D#tb�9���0D����P6�T��g�]*j'�d�G�-D�@���\�*��K�k,X�!�i-D�Tf���|��e�4]�py�%D��n��m놵�P̙�GN�b&A#D��@���:UM���T$�2R�� D� X�c#iB��Yf#O;�
���I>D�\�#fS�/�b��F�8򶀙�'>D��H�@ע;�H�qFE�j��ؒJ?D��@V��]A��[1���r��(8�d>D��(���N4��(����,���׮?D���&b��Ea0,�㥚 +��q`�=D�عdMۛV6�� T�>r���EN=D�@[*ǜg� �I�K�fR*m��.:D��B0�V3��h�$�MO�`�,8D�� �#�6
P8x�j��|���0�6D��h7c��5�F�H���L�F���B4D�|3S,�"|`� �D����$7D�� �l s�3�)����za|�XP"O�� �AJ.#>��cd\C��0�"OZ�&�Љ�IZ1��.s9�=�e"O4�8a'V�v�Z��ŭѠ`%
I�0"O^$�%�Q5n��騶��:F,6M�p"O�Y����.5e�5�������"O�m�f���
��j4bf"O�0��H��d��$��l��T#�"O|�z�B��W<a
�dߔNE2�"O� ��'�#?�0�I��=���{�"Of��"S&㎙ѓGA���[4"O�p���F�lL0�Z$�T�gB��SD*O�1�J�6B��h�\��TmC	�'����o>en���M���M�	�'�՚���P/D�ITc�
�����'��LA㤉 �v]Q����xI�	�'v����H`�c�E49��S	�'r�p�b�A
pyF��� �H�!	�'��@%I��q�E��	ML��'\�	����1��t���3l��'��aP�ڹu�u�4�ъ}%��:�'t�-p�ɔ�<�|�n�M�r���'J�8���iz�$���\9���'��tXF�=�А�6k��5;�<�	�'��D qH� D�pt�f$My^� 	�'D��A��-@�}a�c�.E��,��'�|�(��OHL8TK*�\�B�'���8/Aqzļ!�g�-/j��	�'�l�����-V���4>�`�y	�'�H;��:4�H*�P�:hq�'c.@P���]¨������`�,t�
�'t��*��F>?�!gnQ��j�
�'�F��&
�)ف�@]Y�@h
�'֘񐎓7jԠ�-I�]O�]��'/p��`���krmTaj�A�'�H܁ө 6pA��a�I�2���'tx��S
7Z�Y�pk!� i�'ڤbv#ݨSܨ�B�����lQ�'\xQ륉��/�$1�RDΕ|40���'`���2�O�+x�IKrdO�c7�%��'Gt�J�'mrf q��V��<�']\��#���9�a㐿�\���'�h)k��X2,��0ao�v��A��'�P��D�U���KA j��=a�'�:l�T���Y��03�Փi�Qs�'D�9�r�ݘdB�P�NZ�/��(I�'�,PA ��!^�Z�Q�L#.�l��'=�H�,S Q"n�HRA%-���
�'���¤ �;�H��dȮ(��@�
�'�-���L�h�x���A%$0L��'�D��&��'�%�O/�x{�'�D��ĕ�9s��[�iH��RU�
�'}� (��G��aJ����9
�'_PX���U_:Mr�ɔ��i	�'���N�$�q��	*G� �'ւꕏ�=jA|�b��F�#�X�'�(p�Ë�'�XcP˅�+��I�'�N��C#N�.��;n�'��9c
�'*V-�D �vY�A�Ҫ-Y�5�	�'�F\35�� ڢs� ���%��'h���4,%�(�H33�`��'~6lke��+$��pt��W��Q�
�'f%� K2aG�ir��D��
�'�1�L�E�D�) [�Er	��� $D9R���^����cd��H�K�"Ob����V�b|�P��l�^L+�"Op�q�*t�~�p��[�X�����"O ���d�(< ��@�Ə7��"O*@ b��f
�5k�e�:"�C�"Oм	�E�h�X�d��r���@"Os���"[֡j�?Pь0�U"O\�����$ie�F�W3H�F���"Oޜ���=���Xя�2u��`�"O�hQ�B��m���`�K�v�pu"O4&l��y��T9�8~c���"OF�Я�%���K�lL�]_�"O�]�&K7Y�%���&Qhj��A"O����p肶�J^��5"�"O�XZ5lW:sT�ö���	���r�"O�@ NB����C��4�=z"O���ȇ%S8��j3&�75|�(�"O�!F���#s�	��'�3��V"OKB/l����Ť��A�N|���C	�y"�K#�Z,H���=Z�t;vLS
�y"�E��vȩw��0�,��#�y��4;#���!&è�j!ZBOC��y2'M�|��D�A��pp�NP��y��N'̙��W�4����,F.�y҂גt2�K-t��o,�y�$O.��I��GW u-��ꂨ���y�+Ғ2�p��R�یv�J$XŠD��yRHqQfE�RAP��9�CNH��y2�߉T���CK��J��FS��y��P�u�� ƌS>��QT	�7�y"�+D�@�JV�H�j�@�B̈́�yr �@9�F�O�dX�y�	ͽ�y��QA�4���Y�[�\m�wO��y�d"��K&��/T��12����yb�N.l��ty���9�@�i� ��y��>Z�y�N#Y$=��Z��y�Gpa�J�A	�Q3���0�����'��dEGP�(�s�ٶ%�ȉ�'R�܋��.G�&e�EVlk��K	�'1�d[6h�zb@X�A�*f��<��'������(2us'M�9[lʄ�
�'%�<���4aꈙá��`���	�'X�H�!��1_	&XB�j�_c2�R	�'�z\�-��։ipN&Q2�uI�'i���$�n����<J��<�'@밉P�}�d��sĒ B�v ��'f�Ʌ�K%	k�!S`E5f�Qb�'��E"�A���6���](bEZ4X�'�� �)
5d&��{�LP=h+ ��
�' ���&�[�ΘkQ�20\q��'�*@�ۡ;��uh�C?�����'��(㠜��|�"�δ]a X��'�\�qj�< �"lY�ט��'�z5�A�0��*�W�x��
�'$��!��A�/��d���.�x���'F���qd�$W�,�֏N}kt��
�'�X���e\�1T����'�����'�
lva�Gv�@�@3�:�	�'�,d��*[6���!0x�n1�ʓRH���uØ1���$b9?�Ĉ��H	�u�%�:n딴ZfB۹S�Bx�ȓj6���b,N�|�£oV�T����DVN�x�bH@C���n��H��D�ȓn�Tz��D�m� !��=����S�? @ pBa��IB �ajM���52�"Oj�J��!�R���h�5̢M�"Of�P��q��S��N�@��15"O�$@I c���3���>Ԫ�"Oʙb��O,W�	�*]m���"O���a�"C]�H`wV���qa"O}"v�� 1���sa�E��@��P"O�)s�O�e�:i[�
 !q��"O�w˝$Lo��롄G�un���4"O �Zp�2�`�գ��S1V]���Q@�<��M�2eZ�z���[���U
%]��	O�)�?��b��X����j:�PAc�<!D�L�m���a��LFʌ,a�F�C�<�)^�B^x���WP�\8eC�|�<��bҭ&�n��F"����c�y�<y�+�:�ly��/�\��� &��\�<��@��g���
1?�| �e�Y�<�Eg�>��w�V�Y�`�U�<�����D\����� W�����H�<A- ko�4�G�� m$���	P�<���
v��-�P�K�K)-���f�<�E_(X{D)��8�`8�w��m�<!pN�;�ʗ�#�~�A#`m��X�>�f��>~�(��� 5�����)�D�<i���A�T䛧�H<_\	�'�Z~�'�?u�q ��;\���>](���(D��8#R	n��|��4#�:�>���"�0� Ƅ8P����^#V���ȓs0p���%'�J�#/Ou44D��:�jՈD����d�c/X,��4E{b�'�� ���v����!C?']$+
�'X<@2�j�#�n<At�0 �E��'�F�G٤�p�:��#%z�=R�'�.����G�4�TM[��đr�u�
�'Q��B2G�0lZey���&J���'�
0h��ٓf�����aT\"u�H�,��IC�xT����}q(]e�@L,�C�	9R� b��D�G�1 v�D/CC�I�}<: �aΊ�p4u:��ś0H8c����ɐ(|�4�q�Q11gh���	7�C䉬[��]�aN�6c�Zٙ$G(��C�ɻJD]`w��~8�ڴep�d"Oؙ��F�0��
�J��*iY�<����=��,(x�0�K��7�(t��^�<�Ph_�Q{6؁v �	a� ����V�<�r�\�ju��e"�_����-�x�<��o�N�Ը�b�?u��Y��	t�'�?%���)I��M��o�2H��R��7D�P����=@ 岴	��1���2�A1D�@@�K�TVH�����{B`$D�(XS��`8�������E(�=D����H����qS�L�M��ݰU�-�O,�I,Ph�P����6(%��2�bWv�v#=�'��>IBt�=C���酦�n�`�)�O��'ޞ#!E��-�L�(bPc��J
�'�(���C \�A�
K�0l�*O�"=a��5g5~!q�L>��r��@�0C!�D�-3�����cŊ��1Ԥ7<Lў�P��K�M
"�tQ���W:^�b�"OJ���A�ܨ� Z>:�a
P��z�OY�R�X	p1W�.l�(h�'�6��1�E�$�����kK�a��%�'�@�a@�2��A��gָ�^x��'�@�Z�Bž�8Y���0?����� �I��%[q��*�ʇ�H٨��"O���ːf=����G&8J��"O���1��/�"�+�ɜ�>y6,��"O��c�P�Hy"Ƞ�*��8a:�"O��zҢ��u��5�
�R��!�:O@�=E�dI��WJ*�s�l	�d�0m
@��yb�ԴP-ܝ���NmY�A)���y2kT��D{g�?b����p��5�y��ܧ8���pg�Y���P`Eگ�y�⛈�2�౪؍PR�pp( �yr͐��d;D�.CR渒P`'�yr��1p�T�Ö��2@� m˗FD"�y����Yi<a��%3}C��:�y�'�M�1R�KĐ��L�R�yb$��������x2�wLG�yrnI���J�E��aNQ�&E��y�%�\ҔQQDS�^DI�a�Q��y�7l�U���T�aF���pM���y""��(���3��5H����@4�yrfA W�F�2���X�N܁�@��y��_�	���tFK�ebl�p!!F��y�ELhml0B�nͧF��؛PR�y�B�m.IZ�+��=�D�6(U�y���*�Z���+��4+��%i�4�yR.v�� l�&3@4���F��y�H6X4�i� *��Յ�y5L�b1��0�xk��Ǚ�yRD��~$b"$DC�l|�:��\��y��/	�܍�S,U&]��������y"OǜC�\8������P����yR ���K� �>3H �� �y"���2:6����C�#9��r&^�y�BV� j�E*@�[�6kvF���'5.t*��Y�$�-`F�+\��y��'��͑S���g���'`�L���(�'�H:��(GZ�1;���<�<��'�؈�h�� � 
$�A/EU���'E~�����1��`�*����'e�9Q�Α4z޸�VLO�$ê�'~p���ς
��ӕ�$n��	�'�dkAZ�8`�M)��V.�,�Z�'�L�qa-�t�j�r(S)��<��'���Ѥi_�$��`2�<I���#�'l��{�X
7#�-p���?�l2	�'Nlآbu�h9�Ƙ<���y�'r�}�2�L�æ��,�+,Wn���'{�y@e*�G'���ƥ[0$D���'#JM��,ޘR�,�8�dYs�8C�'�>Uq�0@��F�s�((8Q�m!�'W�ŉ�ڨ�@��Lϓ5z(P	�'�А���:!hF�Y�.��,��'@\ݨ���<t�B'� $�<X�'$�<�5&	�#j� ���s�<Qh�'O����]�x�8���N� �`���'G ��aG߃t�i��V� ˒���'�<�#��A�	}�Z��ي��tq�'H>\�UDN'%�(�v�]5xj����'��بp�J�s��`���\t��p[�'���O^H>,	a�Èw��	�'��#�X+�$)��-�0�X�	�'���ˢ��798`kL�%;�Q(�'���òˋ5E��!Z#�� 2����'h�����5Z�U�+���`��'IvA�cM�9~p �`)ڜ6|L���� �!:��@�7H �4��	h��"OdXB@��N�X`�0��J��݉!"O��J�-$n�¨S�៮h��@�"O�ݘpk�P����E���"O���c@�w���P'�S:f"��"O��8�+JF#���5�/h��z�"O�E���E[t�8B� ۱*��� �"O�0�Y�y��]	dbƧz��D�"Ot���%O�JDH��c,� "O<� ��T�h'Z���f�<U����"O,<x�c�# ��5pƜ�|FPd"O���$ 0�С���'xY��"O�a�eJ0L�`(Qe�ޢB`�V"ODЂ�A�y�F�©���l°"O�q�r	�'�05Cc�F�!��I�W"O��Z����� �h��JN��y"A�'z����U�f��}�����yB�+YbY���ϕe���Y��� �y2j_@�hf��g�Q�î�;�y���}�nK T�S�V���,��yҪ�������F@�P�`�!�y�Sl?������g|������'�yb`J����J����O�\���L� �yb(ˎ@�9�#@�B�b��E���yR(��9?ꈡ'��3;������y�Yd�%� Ђ;a�l��m7�yB˘�A��7KP,7I�T�����y���+9v�����+��0B0��y�&F�tb��	Th�VU(�B�O���y"L���I��o˳L;pࡃ��y�:]�q�CX>y�H�z b��y�kޚ��I7`K�x���h��A��yB��#��p�ړ�-�ge;i���`�M��0?ɵ��w��h���N�5@ihqC�r�<a��	o�t���-=B����j�[�<a�-�	�(Y����6����DKl�<�F��Q�B pT꟠��y�m�<�REW�P�@,�G �!#�N�0G&Md�<1D M.��R�[�o� ���c�<) ��S�U����0`�|�R��Z�<�E� F����\2��U�#�Q�<���){`��G/ݯ-�Z�Hu�<1��)G�8��uj��W��Mbd'�o�<a1C&oh�0�`��nE\�Z�fCe�<�eAB2+m"�����'Z��a�z�<A�n��,AȪ�'B�i;Z�֥U]�< ���/߀��g�E_
#%mLg�<i��	�L�f�A%��m��=��ȚH�<�Vd �1ؐ%Z	L�X"��D�<y�I�J�T!!J\�:�@]�GA�<�՗��\��8R��j��K�<�ը�Nutt�"�8� �q0� ^�<�@J�$�xe+��YoܠYe�c�<��f2s�x� �� �c���1�KZ�<y�eN#n>�C�Hv�\�Q�I]�<�R/Q-D>b���WQ�6|�f'w�<�3��#>���`T+~� ݀a$^s�<!D ۙ(&P�"�\.:��aYD��g�<�K�3Eǐ��dl�Z��Ѐ�j{�<iCP*dM�e	�ɝU"�}BC�j�<�g�Y��\*E��2��"�%T�D���ƲM�fT��`�LZ�YQ�2D�����Q�{Ĉ�Ivx��7�.D�<����eْ�����|�\"�f/D�� �t{���4lxw�(�,� Q"O~2�O�@N8��O3T{�D��"O�aY&cݮς�;���)hQ(�"O
HU`�kî�� -ú,D2H�C"O��BW�@�qR �1���9@�5є"O���B/�6�
�)�yF<��"Op0�5�F3E�R�K�ОB��ɰP"Ov`
S�S���Iʗ'�?ky��"O� rc��"�6,�����f���"O�4+��B�Sy&�"F ��]�����"O�`!�aû*B 9�O;k���2�"O��ńG�*7�{R�N�n�(�B"O�\�F��8!ƍ�A�� (`���"O�$���J`��i$B9J"O eG�<w:d��O��`���"O��R�K���eX��J?��ܒ�"O:Lũ^�M�=�F����"OP�����Xul���ڛ@�x�5"O$511��\�tU�2E�O
 A�"Ob1�!7D�Ȱ"���)#"O��8��X�X<"��D��-�F�W"O�!�3�F]E!���1v��5*2"O�9"!�O)���A`��uҜ��"O8A�-M�k�1���k96�"O�j�1S�x�NG�/p��"O��I��H5���с���)��'��P�G�a�S�O�P̛�O��vo���1dK�`Z~��a"OX�b lA �����cV-2�Ĳ��O���>�ny�	�*�f	�d0%h���㇃&�l�E}�IJT�	=|>d�I(�`YcT	"�~Q�w�N�6`��ЁL "E1!�TD<`!��)"]����dR��� �Ԃ��:�X[҂VA62�4ZR1������Ǜ2AK��G\��́]I!���m�(�"��x����~+�,���ۀQ.��ߴy���? �BO�z����O�@�&94�v��&坴2���"��$�O���EV�_#�� ȏ�F�dp�dF�
dÎ��1'!a��y��FMa� ���vz��'�D�@k� �`�5f��Z�l<��P�E����w`��M�!���z9�QH^4U� !��Y:=�����'�DŐ��\`��C�ɵo����`�-	��S �7H��jk��d`�)��CE�K�u�Af�+K�(�`Y|��<�
�p��K16�@�Ѭ͉ �3�"O�|K�K.r�dm� �҉, �T���50��j�W&�2��2"�%X��4�K�p�jM���S( ��x�A 9?�=�V�M0�^���I�F�ੑ��\	5��m#�B��������>zF��p�](©��J$`��c���uY��	�lj$����:A��!�b�;f7�c���.Y~���Q��)�]��
Z����ˁ��`�QC*�o�(�v	��A�"݋f�֟4����I�D�W��.d�4"�aP�~�d|�0dN{;@�B��A�@��M��E�l�'կe������+��� �n��"E��^Dt	(qDGw�'��@铨��l���,����"����P�v�۟,�|�3���C
`ם�"��Fg�-�T��Z�h��&<s����w`�Eu�l"UEa�����yqO���ɡ�U�T:�ɐ�K�oX�Ѷ(,b�~a�����q���Зf��i�4�z������ɱe����g��*C	4��AD���T�D�QlC�&ds�^���7m�
=�uP$��mΆ��@ҖW�I�Pf΅��(��耩k,a��G Za{�Kp��(�"ѤyXǏL�2���Q�6�t�x�{����FO9\�X�Ѧ��@�A������;`�F�H2���:C��)g��Z��F|2\
C�D�TK� �uC�eO P`���	M��" �sU�<B��ʟ��\w��{�ܔ8�X�y��>q �ݘx0!�F��2�đ���<�W��#l���;��h ��6%� 4
7F�=qeL�C@':VEpf Ԓ��6�L�|��g�+
�
�J��'>F�;[Ԗ�ȅn�5w���խI�D
i�$����:4P�K���<��B��eKB�xe"��$`�`�`�nJ�TB$#��_H<�p�X*J�a;�l�8m�qʒ��b�_�$��S��p�gLU	$��.eͻ|��:Bn�!n^�˦.	�%�l���%N��G��Y�`A�� ONj�n�	^��t��k�.n�h�'�6�� C�b�e�&9���h,H����R&�ȸ��I	Y�L�C䗛R�6er&
�%�μ�ߔ=�61���g�!��U
|m�%�p���DkSD��Ola
�H�)$� Њ2�3� � �%�*X���#�! ��͓�"O���d�D�]���#���35��X��Z?J�B����I9��d9�g?ٗ� G<�z�{��('O�U�<q�]�N�Liq�F�K��	u/���?����AdX���[R�*�p��j"&h�㤝#�� 7�Z�&:a|b@�8(Ҹ!�Q�M��q��+�~���ʇ�	'.b���q�ѧM���Lek��ضC�Y�����H��(O��9�,go����ޑ٘O�j�!⟝j?��q�dI�X,�2	�'9��s�B@>=�Ҩ���n��0z��( ��KM�xӧ���aG�b�F$b���E��q�A	"D� !⊂!����)G�"D��"}2����A�鉉h�� �uh��h&����B�|�C�$����O�<,��AJ0G7�C�I�L:`0�!עd�����2c��C䉔W#����a��@�c�Q�C�ɸF�>)��̴X��\KqA�8]�C�ɞ4�������M��Xx�IP�2��B�I t�<�9#���P9���4%�9u�C�ɦpo�D�V(�&�����I1:�B�I0v9�i�V�?7��4���	�mO�B�	\u�%�%��>Mv����>L�C�	������h10L���ǂc�C�	�p��؈��	�ӃEPۤC�	T,�]�Q&$W��%���Q��C䉱Rm�Qb`�
1���2��+.�C�	�*4c�Y6�����!�>*�B�I��\��݊1��̘'��_޲B�Io+|1�a��b�̬P�c� -ԂB�	%��Ш&OBF{�D:�a�I�PC�	�jP�#V�X��$�ӏXwKtB䉅.����n�#��qP��*�B�I/i�u8!�]Tȸ@�cۮ0V�C�	 v��`s��<"+�]�sFU-w�C�ɴ���S��4�pm�Ӭ	dC�	 ��ʀ�׸G�^�b3.N�OA�C�I9ĆT��#�R����}n�C�	�n�(��Uj5�\Ej��W�g� B䉀<7�zU&W�GO���K�Q["B�	�<!>��#��84�eP�d�4B�I0�dE,�!l�t�i��7��B䉳)S&��D�G ~��0*�>)�B�I?g�:������5Bqx�g_�ٲB�I�#�rhkq/&n��JBn�'m�\C�ɑ�B�a�X8M����ca��"�(C�	i��	82c�K����F�+�C䉜��u�Q�	�b ���䇓��C�	�|OZ[!%�=�$�ۦL��}��C��6��	��.�;*�w�0>N�C�	!VY�����GG>���M7(��B䉊<>6�@��O���m�� �:2�$B�,j�j�R��F�D�hj䌷?\��D�.6j� (�OB�N4� dE�aW!�d�G��颖&ģ��[��]�!�]/DS��ȖLL��Fс`ˡHw!�D�5,7�QVL����@����!�֐y�PH`C�H�`�\�A��k�!�e+�<*�p��L*5��@�!���8`-��/F��쵙�#1!�$Y�m/�h�W�'�n� �Q��!��� CU�d0vQ�)��A7M�j�!򤑻h��5� �;+?V	��@;y�!�Ԏ.�@�ŋD�f�J��
j!�d״l8!��*���"q�Nz!�$��tB�y'@� �Y�~!�� �x�@4it$\Z���C��P��"O�uce�T;iN�9s�eյ ��'"O��82#�	K�~t���P�)�"Ot���ŭ���c���L�
�"O���aB�W�	aw5�]*2"O�u1���I�d��4 �7�ڌZ"O�l�fOG� Y�1��A�
?Ѳ��p"O�d��j�;n�)s)�(q��K�"O@�#�W�Q����^>�b=;`"O���tę'ir�es�:0�>-��"O
��ѫ�&s��8�G�[�´S"O.��̛$c(u�"E+3�`5`�"Oް�%��E��J��P.�7"Oܤ"7@.2�"9 ��/C��7"O�L�wΜ:�ٹ�d@.g0���5"O�D ��S�[g���wC�%A)l�; "O�T�&MX��Q7�J�EL��"O����$�1m�+*$&1�\QG�~�<�bK�+��P�5eU=?�1��t�<1$"U��zs���J`��PC�k�<Q�'�	3zB� "��1'B][��3D�� �O��������J=�G0D���7h�$j����(�O�<5���/D�X��`3./�	��&I�/�)�r@ D����U�me����X�frrx+a�>D�4�g�ڿptdI1Mݩ"n���+?D�t[U�&w88�P�[�R�r��/D���wB�+W=*��H̽7Ur��9D�L��ގt�ŉ�
�&�`���1D�@��K�j�@����?ht���("D��9��F�1�p��&�=�|��n.D��X��`b>dI����b=����(D���&�8IF��g	�t��ru +D�8��"��b�"���-���1�)D�@1e�h�����M�8��F�3D�l�&�U~�b-k����dճ��.D�lC�IE��xT��![bO�)SA�(D�<�!)� =|DH!�d�!O�ƅ�bb=D�D�S��&Hb�9jқ{�B$[��:D�jW͞�H�T��`�R�d���t%2D��𒁒#W16����kT��E�4D��$`��e�#ច3�$�À$D�����m��A�I�m�� �"D��[5�� =/��c��ض[/���I%D� SM�C���PQD�6'�p�r-D��K$I�j[��.1�&�(C��
4C!����d ��e��~j��
�Iܫ)C!�ٻNO�ԩUoځE�X��t)!���9­�V#�(��9�m��7!���>O (��ц]�Bz�C��׏=`!�
,���p���bǄ���I&@r!���w�P�o�q�2�1�@�#_!���6\��+�3I��@���&J!�$�f�X�P�`���S�hJ!�đ2,`J����BM�ZXB�g�!T!��
��H-Q"��bؔ�БE�*4.!�J�`��$��l�3�N�)���Y!򄁽o�&�+�H�H���@��#c�!򄒳4S�$����q�*l�UfR$ j!��fu:E�D*`���f#��E�!���Y�%L�\�D;�b��_�!��1a�F�R� Q���J�O�A�!�A�lr���4`TBw�*�gM`!�DM(�4��ūN	h�3\!�� ����G)?B5�F���+��#"O �cgV��м�p��j��\��"O��@G�@�@A�o]M��r"Oƴ��Ũ]�"Xh���<-'�yav"O�qA�W	F�0:%��	Q&ò"O�� �Ŗ1h��iku/������"Ox�� �_� p����� E���F"O"Q��i1��<��J(c�&d0�"O�E�W��8��/+�8ˆ"Op��S�E��:'�pJq
F"O��`�aA"F�����jZ Y}D��"O��0Ğ}�� b0�FO����"O%��L�6X�ʩx�ㄇ2��,	C"O��:'�?�h��њq���`�"ORq�QF������Sȃ�N�"�w"O��1�mΑP��)P�� >h���"O��s� �`�����E��"O8L���;%�b�Y�%ހ���"O�������$I��E��}�2��"O�, p'
]��R��	1�ڭ�"O��*�,C��$#m�025"Ot�vf�����,�)�$-�`"O�|���+i<��jły�"@G"Oh��#��<�%[B(�1:��}��"O���v)ȓ )lQ �gB4,xz!6"O�@�`@ΑD%�6Ǘ+�x��"OR�[���h�p)�E�90�0�{D"O��$&�o3&@  � =L��"Ov�I���W��E)�OKN��9P"Op�����:2B��"�]�;���u"OlZu�^�P�}��X/*I�"O4pA3���(Ы��d�=�U"O����D��r�n$H��A ���i"O�����Q�`��S��t��"O��c%S�p@�3�	Z�vy��"O�m�-�m��Qg��;	q@"OT�P��7��U�2��k�̐�$"O�v�ۑ]d���gԸ\4��U"O��!�أ!�T0�E��]����"OP�䙈uP��# �� ;=�U�w"O�5Q荙�^��Ղ^9Z;��Ң"O~�4 �,,�L�I��2"Oxiu��=~3|�cΞ0;� �"O��)��^
������ >"e.��"OL piУ��<` �O
"B����"O��+7+�F�<���͒�pNBE��"O����x��,��J�1)��0�"O&�Aa�)�����J̻L�h1"O�M�w��:X`��d��<6|��"O�s҄�:5 �B�.4�䱘�"O"M���#��yc��O�f( "O�$s��@>T�0Z�c4[���Bw"O��Y�`�,-8�`b�-h�^}�"O8��8=��ᢌ�_[rMB%"O�P��`��*'�%� �ǉOM&��"O���&����EۚV:Q��"O��##F�U����aM�;�rq@�"Ot(���sL���<��-��"O�}r�����`���&��%YU"ON�[��cD$#Vb��Da0h��"O���5�ʁ$�)��B��C�����"O���RI�hXN1!A�ҫ	�
3"O E��E�S������g'�,�P"O��(6���7�ʔ���R� `���"O� ���Bس1݆���Օt�,���"Or��E��5��%��Ż�"O������(A�gjI�O�P��"O>�"����cƊ2$4��"O �J�V�wU�H�.� �Ț�"OZ4���R&��f��O�#�"O(�� ��A*B��� p8t�r"ON�ё�0T�,�R�Y�d����"O"Aᢍ��U�V1 wI�n��G"Oz�����H4��!�h��Vi~!�"O�0�@WK���S��(ED7"O~���4rw�-âM��H@j�b"O�@8�	��H��͘�/��Ka"O�i��E� �e�wPD x�"Oрb��/����J&j`SA"O��'��(Y��X �G�T\���V"O.�0�Q7��h�	�15���"O��b�.�L@8�C#>&���"OfԠ�*��IJ,� fE&0b�yg"O<tk3��>4��"#	h԰ې"O�P�$���-�@jf-�}>�s"O�4�+��R����A-^;���"O�41��s���ɀ���_&8P�F"O41��wG�p�c
`����"O,��Ƥ�Ada9ǣ�) 
th�S"O���c�Ae \("!ĺ\��"O�q�ă�4�ԢU���b�,%2�"O4���h`�MK�l�:��A.�yr���i8�o�[��A����y��3rq�S�	��M�`!T�_��y�iT�{�x���i��K4.C��y�,�2w��87TX��r��ȶ�y��qx�cVp�"c
��y�gS/wі�Hi�Kc֙3vG�yB�RD<t(��ډi���⩌7�yB�:5<�<ѷΌ�{r|ݢ/ϱ�y�,�v!�p�AE�ioP���$�y�����߉\���s�+�jfh��`����J��f   �?ɸy�ȓ{�~���l���Z��剓!���ȓ~Z���F�)DԶq{�_	[��ȓ-�Ό��ҴEt5�'@W�Y�ȓk*�8a&B�3�����D�{V4��jz��giַͶ�p�An�A�ȓW?^�:֦T)w�����6B{N\�ȓ2�t�@�Ț6|؂2��j%zL�ȓC�H)��k[/��K)8�)�� W��@�G�z��J�
� mȅ��*���tb
$[���
�.e�a�ȓEH��k4� �\:uO֍H��i�ȓl�d�Rj )zp�2h2[�Q�ȓ�.���l� xN$Uy��� �V0�ȓ?�A fb�	8���b�@_F̇ȓ�J���	lB��3c^�}r	��
�H����Rt���FG5(A�����E����%VR�s�E1���ȓ��q�S�II�ʁ��i�)=����{�hs��P&V`�˃�B�PX�U�ȓ���Tk�:b���Q�A�x��ȓ P���"���F�1۶��`F����IR�|Y�����r㩁�x�bІȓ \�(���Ӡ�~"u(�%l��m�ȓ+IT\J�#Ȧ|�9�aS�<V���ȓ3����j�8&���!bm��cm�P��S�? D�&h�&���� �Y/T�w"O�0���D�@1�4`�#7*i��"O䀲jG���@bo�2��s"OL��Ba�,{:ܡ5Ė�~>�I�s"O�L񦣛�^���9�39>��W"O����3(D,$ Kӧ%z��v"O���Y�VP5�ʬY��Z`"O�]�rn�Iۀ�����$
��f"O���1�ݢ"S���,N(t+d͊�"O�ų ��)��T�����`*x�4"O�CIM��V4��#*Dv9��"O��Ibo�)X�tZ#�·a>���"ODP��LH�h� L#�ɋ�S�Z��"O tإ
�
m����Ǉ2u$;�"O脐��=LԹ�ɢ'���B�"O������,Ȧ��
�*g���K�"O��	'i&mVu�D	���5ӆ"ODXJ�+����;�fЦG�4 �"Ohp����Ӡ��e��o�\��"O�u�3�\�*أ���z]��
&"OqQ �,. u���I�P)
"O���Ԩ�6}>9�sϑM��-�"O��(��Ru~��CD�<�I�"O���R��l?��+#�/9�jܘ!"O�� b� v�,�©��eٌ�@g"OfE��'%���au��� Ƙx:�"O4����p�
&]�q@ ��"O��S4oZ*=�|U�f�-RƌK�"OHd�g�]DN�
B<7\Q�"Ob$!6c��^�@4��Z� `���"O��R4B��Q&��֤	�}�t"O$p`#hE�R����mH��6+ "Of��P�&| �O�62x�Z�"O ��^_���`��<Z�L��"O,�ڥ�W<�2���%U��3"O���s���>��#lZ�i�"O���ӤL	��+P��-V����"O�sP-ԊG	։q����O�<P(�"O0�+�N�lF�(���1v�b-)�"O qr��/?����Eй�b`�"O���20gK����R&mn�I1�/��<F�''
8��D�2H1��@BDY<��3�'X�8�@�U��ē!H%,����'��-� m7Ux�+!	� <D��'p0�*
�c�*Q��=�jI>��ν��<�}��m\>@}�rG���]�~hqr��Gyb�]�v�t)�y��)]�d���B+�:���μf��ɷ>l����.�)�,vZ�"֋ .R��AeN�X2��r�Ũb�
�*��T��)��� ��)p�m�qv#C�lRl��q�Ȕ8���6Q�<���v*���Z�"�0���IE������#<ب�"b+���`YdoX<[�<ʓ�Oc~�������mV2R��m�&�Ǹa�R$���Ͻm�d!+����0|b�I
�k�Me�N�uv��:ZR|��4%5����q��;{H-"����~�K|�uJY�P��Ͳn4}�X�֎˕Z���U,����S��M�;j6�Pt	^�1َ�I��٩t=�$i�F3�	�0|2�K�MlY�׎]{f�J�B�Q��P�X�J|j%N��l3�Da�м��D�P��	2ê��?�~��f�,1�U(���:^�2H��TV�<9��=A7��hS����H�{P�BR�<��,ܭl���3%�}�!�Wn�r�<�.ՓO|���&B[n<HU��n�<�r`��	u�0+ �Z�~�v��C��l�<��Q/b��
3鄷#z��3���e�'~ay�*�Hx<��MՋeB������y�F7&,� ��'����FL5�y
� ����$�T=k�iV�y��Mb�"O��1C��7( ���0(���"O	��"�9:��]��m�6$�	�@"ON�)�'6���(�i�'n��0�v"Öq��^z�l�	H�<@����d"ONm���ߓ{��q,J�|d�Q�"O�� �,�#`FH��̗vY�b�"O���S�ƞDj~��ɍ-s<���"O���c���	������y0�Ub"O�TI��U)1XP��9x�@1"Oȸz�Y(�2��)��5Be"O�]b.mjn0ڳmL�0K�H�"ON�
ce�@z2�C��,T/ܬ2�"O� P�'G�8�4"xJ,{"O2y��s/��Jo��&���'"O �q��N>P��MC�" ����"O�Pk��%���P��e��H7"OL�0�(]��9R����E��"O �҉ZU�����
�%
�}��"O
��AEߤ>����
-M�|"OD@��gӼp�¬��J4z��bF"O,��6 ��t|�أ���Hx9K""OB�@��}�^Q8j4��B"O�Lk2���\�s0g],+`P�{�"OV8�քS� ��P��8PL�(�"O�UYUb��U~Ri��'���Q�"O�)P�Z
7�P�M:l͞�8�"ON%q@�"/��J5�>�A)�"O����hM�C��XX����_Fl
�"O�1C�]�S	b�c��B#��K$"O<܉6�B cr@A CdB%�
m�e"O��؂Kώ�6l�K���|5"O�q����_p�(�2a_����36"O:0�5䉻i;>�ɤ"')���q�"OpK���8�D����GQ��yТ"OȐJU B��I`#��|T�"OtL�� ߏt9Z9I�O�D}A�"OL�ySG�&8���q��|�䲄"O�<X$N��]�t�igʀ�{�L���"O�$Y �ØR#`I ʙ�;~x])�"O�5���-�� !B�%>�I��"O��� >:���Q�m�|�uzF"O"�x3,c�P3ƥT��;f"O([�DU�@NA��g��\����"OP�C���<ʄ���L>@m�Ts!"O�qY"�ߕ#"V��ܼP\��`"O����+ S�TpWʝ9.바��"OhE �+ѦZW��(P|�*h�R"O��eRP�=��7�hI!�"O cC��%#�B���eڼ5�����"O,�(�=G��� ���L�(@H�"O�$�2d�h�4dw�r{̅:�"O�x��O�t]�
��* ��y��_=�89QʔS�ڐ� ��yB�K<F ��ʧ*�2OKZ��rͲ�y�m2Yih#)� I��9b`ݶ�y�J<��0�:qb��a�@��y	��k�0��a��,`���Ja���y2F~�F�p���S��AY`�վ�yr�L��� d��a1��q�ӽ�yˢ&u�����C/`�P$� $E��yR�Tbj�!��T0ڄ��,�$�yҭ�P�Y��c�%QP���s�O��y���=8��;��	�8BY0�}�<� <���׊q������JFp4�c"O�,���ŷs�ވ�����3.�5ap*O���e�9Ea�
��\`�'"�����&M���ˌE�@�C�'� ��!Q<r�� Hg��9.m+
�'�p�����7�^�&�?*ݖ`Y�'��=����-ub�	�#�z�����'m�Y��A�k���E��xO-��'8�$qJ���t�vl�4_bΩY�'�J�0�Ł��aBG�W��m`�'dp��FK��Q���H�>�E�'  4����>��Y��(:,\���'�z)1�cȧ��*UJޡ!/Li��'�E�'�§j���HD�^�J2Ʃ��'�fٹS	��,�æ�xa��{�'I�m�u��6����E�o�p+�'\X�7ɇ�ow�9*���`��AS�'�h�K��4���F�A_�d���'rh��.��x���LC%V}8��'�8� �Kګ��!P��G�M����'�REHq �/4P��gX�L��L
�'rn�`oV�ܳ@��H��
�'���b7�ٹ#U�g L�9�|��	�'6���KBt|}p��2��	�
�'�8m�sKB(���4�69N�z�'����1�E�MRp���3�(9�'��d�V��M���E;�}�	�'�N}��
�l^�Y�GL+ Q�t��'�.y��G61u���	�1u��1�'�`P!�R�l�L� �o��k����'i�h��ɍ,�~3�/ݖa�@��'�ny�E�H5*�@fk�l�����'�B�y���5b�K6�ːz���;	�'K��q�jNx����]G��q��'O>!B�l
�M����"��<��`2�'W|���/����5�ʑ4	�(�
�'h<|q&¥@�� Vk�#�f��'�J4��Ǉ*_��3���*`��'tlQ U��-��Lha�1�N�2�'ld�I `ԫ\��S�iY�_�����'� m#d�݊�b��g�5H�p���'W�|��$Ō`]n���I���'S���ǧ ��cM:q� :�'ʦ�qn�3Tea@��
0��)"�'�n=+uL�;#/��bJ�$ݺ��
�'����qe
Or�0���L���ȓS�<��`D�/t�1t��C�Z��ȓK����&\ ���Q�@e�x��X\I:+��s���AQC�=����K�>���C^~x�ۂ蜝}Kꠇ�[C*Sh�� ��X� �K��x�ȓ9O�IRp�2qV�%{�A� 40��L(Jxg��j~lx;eNb;�y��y�0�t�%�P�kE�F�|���ȓm;D���>8�r5�1�O15Be�ȓ��<��bD�o�^�SP�4~.�Y��eH����X �Qs3�-� ��M�r�-�I���� �*�z��$���a�郯9����XBT�A��5�n�EE�'*XD�@'�3������f0I��2/"Y��/Gmp���'G�<Hb�͘^^3#��1I$ʕ�����2�X��X��$��1E��I�ȓS�ư+2a�� ��oC���S�? u�A�ħ+� KO�_j�Z"O�IYB�ߢl<��Dt��tY�"O8�	3�¹h��z�.�.9��]b3"Oz �6A�H]�b�,�ɒ�"O�ظ�n��,ش��Eg��V^�"O����`�3�p�2�(�Vيc"O2H�S`�a��f�LP��e"O�	���e
�� �+�%b��d(!�$��&�Dd���~�:��T�U�R%!�.Ex���֎�'�,���2!�
.u (�#�>R��`P��I2ko!�ބW��\�AѠ��}0��֎!��D�~	,4�������r����P�!�ߓ�n����$u�3��ي?�!�w��Mp����>�* ��� (�!�D�	\w��@f'�=�X�� �!���,�t�B�'�ܽv
�h�!��E:�ج[V�g�M�T�R4�!��T!8��m�r��m��U�7�E�g�!�׉�DI�]�}��(6��Q�!�$�Ixy���t�Z�j�1F�!�%\�f�a�Q�y׊z��L5t�!�DU�0�t�QT��7<]����A$�!�D�H����Лf2̲Sל"�!�d��^�4�6EIv0�7ki*!�$1I"�A�F8F�Ī"-��8!�d��&tv��WgM/E��Ȧ�Py�ءa?�)�M��'&y*d�ڮ�yrf�
���DF�l8�֒�y�B[9viM����H�r��:�y���r�ة8B��6QE�k�E�y������Іޡ2� ��� �yR(�)o�UH���h��@���y�i�-@�(
�*	�j���3C�y�����҃��2��pi ��,�y��K6y�(!t1>�'	���y"V�8|	�S�� �@�뀍�y�<8;�q�Dqm;&��d�!�ߜR�~ٲ���%M�*�'@'�!��5G3^E�G�%�n  �hB�	�!�$֘�ȡ��d��B��mI�Y�!�dJ�!.4��+�?��(;u��SX!���Q��
0��+�����;F!�D�yw�E��̊�yl��H��!�P3slZ��«V -s�e�JJ;S�!�$�:��CS�N�ȤٳC��>�!��:wݎ�*����_HU���sx!򄄯{�����^'BR��%��Qj!�<L�
�+�n)G�(�k��p�!�d�*0GB�{��O�cj�P���6QO!�\�=�6d�C�r�"Q��aV8R�!���X�. �e���X�r�A�&�5!�$�O;^�s�m 5S���9���!�D��2HB��A�_M��; n32!��˰EK�T��ϫ.� �I�ķ	!򄊵I�D�C,�	��b!����!�DL�6���W#��*`��F�U�!�^&V��*�
��]�U` �.L�!�ҏf�fDcK�lYfx�n F!�DA#��%�V@��x��V!��X)
�jIJ'g��?0d�F+��!�䎙�]�CkW�	&h������!�J�+��h��_v��*��E�XV!�DB� ���^)2
_(��"O� �Q�N�r�% C>��`@�"O�t�Ώ{'R]�ph�FHXe��"O�t�$���u���Y���}�"O���A��	g~a�Qχ�"��@
�"O�}`��g�mIԤ�.b�e9�"O�qC#�5�]�2ꆾ�M��8D�|2�
   ��   J    �  Q  �*  �6  'B  yM  W  &a  *j  �t  
�  ߉  <�  ��  ��  A�  ��  ů  �  `�  ��  ��  '�  n�  ��  �  H�  ��  h�  C�  � c � 0 �# !, �3 �9 1@ �E  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h%���븧�O@��1�AE�8�QP��Z�	$��
�'q��&װ-��J�gI�H�'|�仳n޽�j�R���*[�����Z6����C�k\���T�[H~�B��D]HV��
	����2�W;���'�^���d,�'HW�ePU�K�D��!&I�� <��6���$�8x
�Q{�/gY���=��^�б3�)�+("�F/W�4}����ys���Lס8����R�%:������?��.ߥR������'/�F����j�l�L<�@��=l�{�nM%VZ�����i?���S�^
p�Ė='�:���l� C�I�HX���4������ݽ}z�C�I5n(]r�'oϋ%P:ӣ���?��Ob�"~���/Xr(+��ˀ*tv�	s�E��y��]Te(���aE1#ǒH��f)A���F��4�$�͌]a2u�0��@���q��"|OHc������Ţ�\�?� ��>�	�v��yh�5��dY�eݽf&:P*�Aޚ�Px���3:� \I
�<I�y6C.9�֑���>�4�*lO�0�±�
������ڨ����c~�>q-OT�	�F��pa��G�z�qf"O|	�t@1����v�K%H�J���"O�كh��<������47u�HY��',h�O�i���B$;��hu�Qzj�(�p"OheБ������ �_rW�	��HO��/od���
b~t�`��~�B������*� 5�d�h�!�(ǶB�3L���a5���Q��?�RC�IM�R��&l�����G�g�I���?	r䐃]Lx q"̖�G�flpc�C�<���+��XuF�/�}����}�<��){ji��eH�T�H��R��zX������ ���J��ZVvE�$���m���Q"Oظ�AQ�W�4!Z��۶7^*8��x��)��!WI�8�Ȏ< �����)J;JW�C�I9~@ h�)N�̖��臰T$����q��G�y��N H)�ݨ��ב5�b���+\܍8�X�`�J��0l`2�D|2�S/����gN^+z1jE��>�C�	'Gp)��@������;W7nB��+O��Qp�L�*�m�)�~�BB�Iz7�l�E��BMx�{����<6m�����'��\�Aބx�8����ؕ2��H����$�<!aA`}j@�'"m� 2�U�<�4�C>y� �R��ČF�ȅ�ULT�u���O�����@�V�:a���?�X�
�'�` �,�.��ujw��0s�Ԛ�'�V���*�^��s��Ŧ,N-+	�'g.%�$S6*i���Ԥ��]<h�'-�$��WC���R*7Όq��O©B�ɖ�U3�C)G"t!��"O���Tc��t�:���Pέ�s�"Ox�r��f���&���\��8k���u���'C�ؔA��V���RBoشo=�Dn�R������OS9� A ��C.����1�8�<	���O޵C�
n沉ar-8�Ȅ)@"O�iS��#df���Fꂑ$��{��'��	-26pQ5%Jl&��%��ZD�<lO��<��h'��J��[8<�����9D�<���J>{y�R��5�μ�p6D��c∝e�tLڇFK�F��@�.D��S��xj���`"	�{�̹7G9D�d��G�6]��uL�. Xr����5D��s�c�d
D r��z�(P��.D��ؗi�7$��m�� ��0��|3S'2D�TyϘ47���8��B�&����*��j���'U��(!l0&]X4�2c����5�}�%��$W�ژ#��7K����)����`h�3�6M3��<aj����8D�C' ��f�t���C�sQj��/�ON�[
�1�5��
Հ��to-QML=��>De��)4@��"%ȫ|Zͅ�b�:��r�HvD0k��1� �=����D�8&$���i�e꬐���>�y�
�=����`��I����W�R�y��І���Z#FB+X������6�y�n�	h����P�:T�r�/y�����A8�x$Kk �1��P#Ԇ4�����$@-Jy!�#�G&�z����<$�0�T�sYx��C�Y���'�ў�|����#v�ᙑ'j�C�k؞��y��Ω�,�BT2t�my���y��Pb! ���#�<U�!P���'�ў�O�x`��Ku�˦�ϟ�ex�'Q�i�@�M�E6��Q�A�	�4�'V��QDJ;���94L�#9Oʰ��ј']j�3BNߨj�x�G�#��`�'���jP+�-gN��jP�X����cӮ�}bn̊#2�m�ǅT ����Zr�<�a/O(1�ޡR�'�Xy��	V
ָ��D{TO?��ݙ3y��$MN�!�d�C[?S�!�$G�y��qFb��0P��0�F�*����>��M�6
�P�ꒁ�.j���W�Nr�<1����03��ǡVQ.  ��q�<��B�Heb}2����2����To�<Y��+Q����`6XF��F@�n�'��y
� ��!ыe�he�1GC+9m�t�`O��j��0Q���F C�
Q���ج��T8����I�'9�p��e� ����+4�Ot�"�'��l�`�[����s��s�|j��HO$��-�3N\��2���P%"OޘR�CKe�lm��FW����c5O|�=E�t���\#6����/�n�`�N���y�M�fs���7j�:zl�������џȅF�:�(��4gE6��3ED�	���$�<ѧ��1$FH�xd$VNΠ5��a�p�<��A�O�H�2	 �(=��2�kQ�<�1ˁ�r��y�vʽYR6!p5a�M�<����C�\��J�9 L�8sd@��D{��ɗR%�I�e�=V\��O]� r�C䉲#J�Q��G�x�Ԋ��.B����	�7;����~��hOj���L�?}�4���`��K*���'�2 ߳
4b�얏�lՋ!�Y26HoP������� )|!@E�Z��v���
 �0=u�?�(N�Q�Q.�o��ݪ��E�V�,��p?q�F!���{G۸��ؖ�]cX�,�O���E�M�a@j�a�	#\���R"O� ӿ�Z�00��H0ֵԐ|��'��O^b�(#�l܁2P�*s�R�\��ǩ4D�4Y��y���h�Ι&a��0D�|Sf�94�,%��`��w,.D���K�o;�0����> ��b �'�I\kQ��Os`����4$��M_'>&N�P	�'Wf�# S	���8����*�NE�v�:��h��_�#�����n_�AF��0SE;*!����7� =� D�"	�H1R���A�'�a�iZ�UBج��S�Q�� 8���y"��zh��Fo�J�d��@�y���Ql�X�P�4��͂��Y��y�ܩ"Pɩ"�J�5Cd�#��+�y�
�����2��=Wk����:�y�@o��:pH�H���$ �<�yl�aEX�9�o�2H�\\rtB��yrGOWG$�(CfR�sܐ�6�ϋ�y�gJ7.����F�q�Q ��ߘ�yƔ�P��<�1�A=�`MYe)F��yBV0D��t��(�:/�e�"P>�yr�C�[
|�p���#$�4Qd\��y"bϵ>,�]�aW����#0���y��K%Y_l���,O� GNL�B�M��y�8c5:5��	�#�!(g�R��y�^�6�Y &�ӱw*1&		6�y�j��o=�����i���y�F
H7^D���*E�PѱaO�yr��*8�(S`���^8*qL��y�CE�UI����Р�p$�y��D��Cr��4n/�`�Q��y�I�1A~�"��s�p-3`�6�yB**t�yIB8o�q�'nâ�y�9�fȢr@�oa @ʖ�yB��8^Jd�1L�,�rk��ybF�l�8�)+ ��Aqf���yr�?p���1��p1�J��yRĈ%�!�i��"�.
DM)�y⣋��e2 ��	&R��b�A5�y��I5hb@l��ٗ#*�[��R��y�FD"?���-�<���H��y©�Li���-����/��y����e�E�S�U�)Kp�QBY��ybG��N<�PN�n�t���(X��y
� L�����S��z�ŠdrR���"OJ��4���C��5�i�j�5�$"OD��P%�pD�P�b-�蘥 /D�pQA�OY���JN�77�����@?D����Cͯev���R~ְ���O���O��D�O����O��$�O(�$�O��(d�Q��5���� � i�O��O����OP��O����Ox���O��Ѱ�΂�R�@m��,D�RM�O����O����O.�D�O^�D�O����O��@�؛���"7�������O����O����O����O��$�OT�d�O���W�M�Q�ҝ���1X8�tᑻ�M#��?y���?y���?A��?���?����^���P�(��|�"�����?9��?����?���?����?���?�VȄ�|Qth��
�w���ڂ��?���?����?���?����?q��?�5&R'q5�|36lL�)���;�?����?���?!���?a���?	��?qD�>03J}�hL�B�xтB@��?i��?A��?����?	���?����?�DO���[P�\��*e)o΄�?���?����?	��?����?)���?I���JQ�HТM�q�t1����?Q��?����?I���?����?Q��?!�{Iʅ�/���ӱ�P	$x�	˟��	����I����	꟤��۟P���n_\Tq�J�);8��;�G� -p\���ʟl�I���럼�	Ɵ1ݴ�?A�tm�(0�/Z�Z�,�XQ�Q�&� @��V���	Iy���O�mZ
/����ށ�Ր���?9�E���<?Is�i�O�9O��DQ'6�΄C1M_ {0�����n֔�D�O��!Q!g�����$!��4�O���`���'N�8� �J��S�5@�y��'R��O�OZ���_%_�e�Dۢ��x@��i�����d+�� �MϻC��@���_8(��eMR�P��D:��?Q�'��)�S4:d�nZ�<adk�5 ���&��Dr�L
b�E�<a�'�����$�hO��O�1PL�`^�1!�Q(`2v7Of��� �v�M���'�����h䴄���X�܌a2��l}��'��>Ob�V�RMeˏ�~�����K֎>b���'�b���^�H���d����L���'[ܸy�,�
��A��ǡ+��Y�U�X�'���9O��ZC��`�]�F�D�r(�Rv1O$�ozK�j�Bӛ6�4���2`�	e�8
 Եs`&@�E?O6�D�Oj��	�E�P7�(?ɝ�៸H�� �e��L�t��Sk��(��P9������d�$�D�;bk�t&�jS䅭?����M��!�����O��?A����P�V�ç�!�!�����$�ئ��4%����Ox��s�N�J�j������M�6K�T����VZ�����Z�Z�'{�Iky�O%5��p,� �ۄ��-/rх�*�M��_��?i2��J�,�ȥ+T=dy>�Z'���<	��i��O:i�'x2�iN6��N��$8���9��e�Ă�����){�Z�h��%*6�?�'?e��	p�҅����5�T�hQʖ�!���	x����PC�0�Ҭ��4�.Ո#��NyR�'�6�]�p��4�M�H>)�$1Dʴ��N
|%���?���?��|��S��Mc�O���cNf�X�-ˏI7$�Ҏ�3vRfk�$��h'� �'��Oΰp��1lk`)3�E�0|ɖ Xe��M�Š�&��d�O�ʧ:��5Z����#�J�s��U.wЂ��'*��?����S��aͮ[��\�A��Z{* ���I/�T����$Q�o�<ͧ_���^�8P��,��T�G��Rϒ�~����؟��	Ɵ,�)�SLy2r�D���C(~\��������ae�%rY�I��M���* ��̟���&SU���"Fp!�*##x���ݟ��u�����̓�?i��ܙJ����y�]�����g-�24Q�� �'@��y[�@�	ٟ��I���	ҟ@�O�B�0��@��x�+� 8h��Q*r�F�`h�Or�d�O:��v��L���	�l�J3 !=�9C��G�9�^�Iԟ0�K<ͧ�?�'>��Qٴ�y2LلIfd@�K
	���yRFV$/|���� o�'*�)�0�"w�;���B��tK�_E��9ڴy��,O(�d�
��`A� ȁF&U��8Y���O>�$�O �O`2�לLNLQש�)Z&��2���B�Ӌ#��mڕ��F����(* 3�>�c��O2F9�2�.]Ɵ��	�l�	��E�T�'~ء���>w�h�S*�s���v�'�6͚�p����MÈ�wcȉ�SI�$x�A����?jT�i�'��'fb��Uԛ6���1��Z�Uc�i�}޶��*�2x�(�b���m#��O �S�g�<��8{C N�Hst#SF����'	�6�C5l@��?�����*H�\)�@Z�Z�(�IA�F�!�P�
ћ֨b���$�b>	���Ѥ&b���ND�k���*d	pv�lZ����U�I~���'$�'=�	�?��C���V0�#f#�C�x�	������$�i>Q�'��7�@�CN��\<�X1�hSZn�P����^�����Ȧy�?A`U���Iٟ���4�V���kL8P�̚�ّU"�R�!ב�M+�OP� ���0�2������ X<�D��t�͹�J�P8��;O����@pz�P`�3F�:���b m�x��?9�i�N�͟f�nK�	�r||��@� ;�|@q��9��!O<���i��6=�*i)��f�~�6��e$^�Z�"M�c
\�1j<_E���������O����OJ����6��I��\�K3N�`S'W�)2��O��Da��jP���	���OM��"B� ?���H�) iz�O���'���i*0�O�D�O{p�c�fӖa�1['o��:`0��,&���Bu�Y�����|m��f��O"�X�G)�"(�%�T3#.�ebj�O(�d�O"��O1�~���a�5�b�U��r���l���$*��'�RboӀ��q(O6MX�"��(
�i
,4���� [((�m��Mk����M{�'��\t:"��r-�'1x�F'�7cFX8��%�T��'q��n��p �f*[�D�H����MK�M�ciވ���O4�?u*����� �uwЩ��Θ1"�P�3���?Q����S�'Zt�Q�4�y2��M�D��I�3]��`�5�yR��I�5��������O���4�V����C
7�x��n\	(���O��D�Oj�R��-D��y�'���P�Vu����M	(A'���O�H�'��'�'����i,_�.1�G�D/^x�<Q�O]R���Z��7�%�S�&����O��ѤvB Cv��
���b�O��D�O���O8�}j��+%zu� �%0����Ģ�L�nh��'9�n܁5���'�6�)�i����"�z���	[(m�2�����Φ��ش��ش��䍄�y���
��5{E)ПrުiTaJ�&aX:[�?!,O���|���?A��?���"^�<��Лu�|�)��'¾ѣ(O��oZ�-!�4�	ğ@�	z�ğ���	^d�P�jn��XF,�pr���?��fۉ��OGBI�W��5G3&�4�F�2̒�y%��?�JHS�O�%s����?��L&�Ġ<��JQ	>���j/:z��P�\��?���?i���?�'��Ҧ5���ϟ�0S�̧��p��-ב�ʨ���o� �۴��'�
��?Q�d���W�#z\I��l�/#o�����#5�"u�Ҿi:�	�#����E�O�q���.�'&юI�嬅�5�Bt����3w���O`�$�O4�$�O��� ��f�����gǇd".�6�;C�@�'�}�8��s�?��4��1m�1��M2s�&ur0]*(�h�1K>q��?��)��H۴�y�'`��b�Ǔ(�x�XTH�|��!��'i>M�ɊE��'k�i>1�	@��:=DE[�Ή#4����"��+C�������H�'�l7M �����O���|�V��OXm�w(�Mb0�I�`�M~�J�>I���?�4�xʟ�	�]�^�H9�&�V�fC~qҵ���x@�虖��n6�i>��c�'�l�&�ppC�TNf�(���
���"�
I��H��̟d���b>є'-�6M
oh� D�n�(��V�n&��P��<�i��Ox��'>�&�('��h��}�x\p���.��6��٦�����Ц)�'��(��DB�?I��Z�#�d�,/]K�(�>[��k�HH�$%0���#Ҳj�ʽ�!O�@�����&J�*�0G0�6��Zađ5�4&��Y�.��j�����Zo�V���k���j	���ɀ'�@;9Ɋ}�-Z�q��l���O(���d���C���hW&hIB�%�xx���> t+���bb D�S�m�ԥ{�BL^�x��@� 
�@�  ��/&����iEaܼ�����_$/�daPE��`���%:���RRjBI�A!�1.��̪E���
v�����Y�"� 0qS	I�M����?a��
U[���'�����/�8|dv�؀�
�V.ؠ�h�D�G�,�	�'�?!M�/v�,��� ��j�:r�M�r7���'�Z�M�S�蒮Oh��?q�'fNX)Rʹz<��('��
�N�ٴ��4Dh�a��T�'~��'W��K႘�W��=Ic�	�,y�,e�^��V�2h��'���͟h'��X�;1N����
�,ѓ�˞�l�-\e`H>	��?����$Q�pdx�d��b
̈�dJ��-��LZV&YG}2V����z����I�~d���I��5�<HQ���$M4�vO8�	Ɵ���ٟ�'���qP�z>����  @��q�"!�9�rȲCKc��ʓ�?�N>���?9��L��~B� ��䑢�M�Y<-�Wa_�����O��$�O0�&V�	P?q�I���(7�^# ��kpL�J�\�ܴ�?qM>���?9D E��'�f�`��+g3f�3���<�Xa�4�?�����B�X2�Y�O���'(�ġB1`)��W㎙i�$p�
L.-��OP��ON}�Vj%�I{��.��S��mP�ѶUFD��צ�'���Nj����O����NDէ5F�A�H�	��=|wF���xyo����,����?���D�\'*U2�`v'\�d�(l��+��M�`��Fϛ��'��'-�T��>�(OXQ97Ȕ� N�����1W������EΦ����v����O�H�p�q� F�%f8���%.U�7��O����O����Sq}2V����o?yC�d�����-�] `Y�D��a$�d:`!���ħ�?1���?Ʉ��l�!�3kT.8<�C�L����'O���>�,O��d(���ڥ�JY/���ಬ
f8��s�W�Hy3��W�	㟠��ß4�'0���h1�o�袕+��H�x�`T�l�'�B�|B�'�r`�Y�$��kJ�2m��f�(5��@ e�|"�'���'��	X����� �Hx��/K�@� #��02:�x7U�h��ן���{y��'_�"�/�""L%��8
e]�Yl,����;D��?9��?!(O.� �PE��1�����F�9��`s I�[�`���4�?Y����d�Ob�D8V���,��,ׯWb�q�ժ~���z%톊�M���?Q-O�x���
k��s�����X���!�m(3�ӌ(��7-�<Q��?�k�&�?�(������k��eʚ(9��Z�tnH�〈�s���\�l*'\��MC�Z?���?A�O�)HVo'M���2DF24�<�#�i���'|�t�'N��)�|n��h��=�G�V"H� J��^)P\6M��j�����OD��O$�I�<�O�������p�)��E��!{�iӖ!C�π�ZE1O>����̭uL��H
b�z���B�T�ݴ�?���?����*i����T�'��-ԏ�L"AoW�\W�����bl$7��O����O�qFJ�d�T_>���^?9�K��pJvG���֍��+�ݦ!�ɼk��̔'��'��'Y)sb�X�1�@T����
.��Χ>�k�9y.��'��'O�P��q�V�"�h�RŒ6d�h��	EbE3J<����?������O(�ʜP� �qІŤ����B� �C��1p��Oʓ�?���$�O���v�?ݓ�K�Y�\T����,���n�L���O��I⟔�!�] E7���|�n��7!_�*C�X8 ��;�	��d��џ �'�p���(�I�8ϒ|�ӯ���Ƽ��O�oq`�l���Xy�'	�"�UO�~"�F0B��Y�f�fF���¦]�	�d�'�FE��M8���O�������q���)�M��MCm֔r��i6�ܟl��;`E�m�	^��?ט,��=I!�'D��-�����6��<���Cg���~����2����R��
�tŰ����(���£}�����OF��O.�'>�	i��4��jAL��]L(`ZҁE5c�lo�x�Q�۴�?i���?a�'>r���\cn�� �VP�6����:iΎ�3�4>��B���?Q��?��'����5�=۠`[�3����p�H9�M���?��)��i0�x�O��'�<�6�57�� 5�֌Q(l�a�}�����O$�Ĝ�a@t������O��Dȍ,�p!�P%�;]"�����v~�4l��5�K���|���?�+Or!9����<dtD�fU�.��t�u�R���	�T���IWyr�'�B�'\�I�|2Z��c�N;��l0���4a�,m
w�Ń���?����?*O��d�O�yv�H��[g�Ϥ>#&�bEOZ8�$���<���?1.O��D]>{���Sr��M��m�$m�y9�
N�7��O��7�I���I�^+Ě�lcӆ���.��qachL6g<]S�X�t�	ԟl��jy�B��.�
�d|x��K��q���`\���Ŧa�I}�	wy�AF�2QR�~�DjƵ���ɣ��j;�17����u�	ByB�'Tj%+%S>}������s�ie�\�9�6�DG�L4Iz �'��O��$��2a0��T?�Pf�^:�p�*
y0���d��ʓn�T@��i�J꧃?i�' ��	m��ѹ٧C&,Բ�[�9466�<qGM�?����TR>���z�j����Cd ��r��.i�Rmnڙ0�ܭX�4�?���?y��i�Imy� W:���ɍ|[�M�!J7�EY��D�O0���O�?��ɆNp�(PV��X,29еΖ*.�Z��4�?����?�0����Ty��'/���R��x�a6�`4sF�_b���'�"�'�r`���)�O����OhHI 
�O]D|RDҲ!s�d�J�ʦE��$Hd��A�Odʓ�?�+Of���XhY�����m�0b� e�R�b�V���1�y� ��ӟD��ڟ�Iry2Ȏ�Ib�\�)�;IԳ����������>*OZ�$�<��?a�f̆�R�
�NV��& �������<����?!���?����3<>M�'p7r�������#��'1)��mZLy��'��	̟���Ο��`�l���5�0��01�F6t@����hֿ�M���?����?�/O���D#�z�T�'3��p�c�v�j�(�;UU���j}Ӵ���<���?���a��h�O��Ą�1��dYDˊ�X*M�3�v���'�[�`ޢ��	�O�������;%��U�4��W���2��}
a�[x}��'��'h�ʟ����$땕YF,����!�i�g����M�*O��������	ן��I�?��O�]�9ǲ="7�͞v�P�1�^+k�&�'�bM��y"e�~���O��a+�-�x��R�b�]�@�۴���!%�i�r�'d�O\�듿�\!:%�Y�#g�8+ u�S��C���m��:&�����'�����j3ph{�)�D��� 8�p�iM��'�Rg�����O��IW��" �jX�ԓq��r*꓁�@�Ba�i>��	ԟ���p;�P�W�,D�hd��'Y����Jl�*���`5�Q�'��I؟ȗ'�ZcNx���*�vM�EIZN����O��38O����O��D�O4��<q/�(.ܠ�v(Q0MvF����RE!<\A�R�H�'��[�L�I՟��IO4�8��!G-"��P���6�(�c��k���Iʟ������ly��Ǧ
^��V�ht�sj[ 4�T)x��H�a��7ͺ<)������OL���O�E39O�����]ZD�s�̀"�<T*�L���=�	柄����̖'�@d��~�����3nz�a㫉�F|��ـ�B��U�	Gy�'B�'�\��'b�2JT9��	��H��T�Vؑo�џL�	UyR`ݐ%��'�?)����P� ZL���)p)�QR�%�Y^�p5^��������0i��g~�ڟ�)����K� ۄ��]����!�iub�'rN�J#aw�D���O<�D����i�O��g�R�q^]�gK'� A�jX}��'��(@�'�R�'-�Q�i�pvV�4�ڦ9�i����wp�� #8(�7��O"���Op�	�p}�Y�d�#m�$I��CD�1Ҳ8dmN��M3  I�<����"����H��Ͽ[��a�l�	'2���Â�M����?��<!te��P��'�On��u�>q�V�Ai�+�ru8�i�^��P �b��?����?�u��)W ���q7�$����!��'�J���>Y*OL�$�<Q�����.�=�VE��x5�*�s}Bj��y�[���I���'?���g�F,��4���	#��?J��a�Oh��?+Oj��O>��WmT����
$��1!u�M��u��0O����O����O��Ī<�T�W3󩝶
n��t�Co����Q¿Dg��Q����Iy��'���'��,��'V�	��	��1G	4�s2e��M+���?����?�+O,��t�Ec���'$`��'���9����lݺ7����Q�u�&��<���?��e�̓�������ː�qi�ɋ�4���oZʟ��Ixy�k�y���?I��Rs`�(���b�f��Aj�+��K��I��4�	˟p�x���yBٟ\�`Ů_�����s��C�Դ��i��$\p��P�4�?)��?�'b��i�)�V�aƬ�BW#ѣ6�&�p�{�H���Ol��D����'6q��i�#(��3dxTk�G\�=l�Q�i&�8���l�2��O����H��'{��A` ��$�2=8���'_o|�)ش(����?�,O��?]�I�O�t��B �@St	��+^��4c�4�?����?�0���O�	|y��'&�d�[�bM�e��6Q�0���ZF��'��	PU��)���?���[��0� RW���%�D�^�v��ӳiBK<WG�����O�ʓ�?��S�B[�̃�$Z����Ɔ! ��'A^@I�'5��'���'�BS��I6jG
B���	@�]��h�?M�tD;�O���?.O����O>�$ӱgh�B�B3NP��
/�Rt��6O����O��D�O��$�<�q"��`����2z_|���� �oK^��c��ڛ�_���IZy��'���'lΨI�'��(�l����u���^����uӔ���O|��Opʓv
���Y?��i��k��8��ya �+J|'tӠ���<Q���?��iy�����dߴO0�=[U�	 ��U�%�>��f�'�T�T��Mڝ��)�Ot�������8i��hEL�Gp����,\y}��'3�'N.�ӝ'�'���A�i����7�6��� R�0�&]��Ѳ�%�M�"^?��I�?�)�OD���n�^5T�(&�V��n�B�i����lR�<aL>!���-:�X���0����Ҫ�M�
Ee���'���'��$# �D�O`�qڡ��R�k�����f��z�aI���'�"|���J���*c�?��Z�`�� �p��iG��'����&O���O&���@V��S�E�:��ԫ姅<	{T7�*�D��3j��&>���ʟ���c�J)��g�&������<I7��3�4�?ё�Ra;�'���'�ɧ5ƍ�_E�AIЈ\���T��cI����[X�'r�'{BU�|X�F���-��<�ٵ#��%ndQH<���?AJ>	��?)�L�n��%�!e�;h���� >9V��������O��D�O`�(Z�ᡤ3��˅`ܤNR��b�$E�%�TpБx��'Z�'���'κЫ��'�t����T�k]�����>y���?����$Ԧ��%>Ma%��� �4�Q9ॊ�7Oś&�'��'�2�''p�y�'w�Urx��h�5��Rt�l��nٟ0��xyr��9���p���X�Cы�j&r��.��)�"�"-�d�	�@�ɶ����O�	@R��#c�L��,J�gJ�HU'঱�'��P�(b�F �ODr�Oq$�0��\1D�C�/|��1��SU�̱m�ןt���i5��Ix��T�'���� �	
¹�3�C�b���nzq��Pɦ)��ǟh���?�1�}�\�z�NaX$,6���CD�P�2"47m�i����9��;�Sɟ�;��D%()X�+��]�D���.��M#���?��[J�Y����O4��p��i�"��Z��씷M�6�?�dӸ! �?��I럀�	�c��#��P�RN�j��C.o�HB�4�?)�I�)&n�'�B�']ɧ5V�M�yPx�cm/�J�7/F������Rm�<q��?q����$������ǈT~���-F7[����cJ�p��?�H>����?���%	މ˷οPd�\Y�m� bڱ�������O����O�˓a:�`�0�p�y���%H�AY�eݒX!���Z�,��Z�'k�*_�8"�HQ#m6�"�&A0D���T�U�1x87��O����O�$�<��Q":I�On6�E8KZ�2�F�D�`�q�{�4�=��1H�Q���?1�'������
�s�BӐ}����4�?�+O��d
>A�����O���O��ܮE��=�+T�I
�x�cӼ��$�(���s$�݄b��'L=>�J`%Q�<zm�g"=���l�Gy������7�N���'��D�>?W��1�M����/1�˦�	���3-�S�g�B (W�ʇa}L��D��&[)^@l�;��a�ش�?y���?��'0�'.�!� �����eRQ8��'f�a;S�i�􉃈��۟ Gb�7u�P���μa�`�F��	�M����?��'U�P���?	,������ܸ4�=p���0p�U��u�K2��';�8���1�i�O���O��w+J�+9�+�'���P  �O��D=��u�'���h��p��E_N�� ��',p�JW"7d�	�)�<`%��	����	�����:e\9:��M`ti� @�Bn�����矸��Gy��'��'!��O����ݕ,X�ZE��
oy,�JѴi�`H@�O����O���<q`'�`N�	Ă01�d�uj�AH�8B�&�}2��V����~y��'�2�'CVIҙ'`b����	O)�T��#m�����Cpӄ���O���O~�Z^�ej�S?��ɐ��"�@ƲvB\�0��Z�U:۴�?�.O����O��D��WZ�D�|nZ9_��(�/�8��d��&-�6m�Op�D�<!Eد�������	�?=�(ӶD�jU���Y~�0���E4����O8���O����?O��O����
^}�5�Z�Y����$�z6m�<�p�J7C*��'"�'���'�>��i	F�Xԏ=g@�c#LRp�h�o��t�	& h�	L��h�'w^4�#ϙjjڅc��(1��oڼ9U��"�4�?����?��%g��ey"�τ&���b �tR�)�> ��7mݞ�~B�|2�i�ON]��m��w�H���+�O@�+B�撚�����I��@�OH��?��'1JD���U-�`�@��6(4���4���Xx�S��',"ޟ��0��EdN1��br�Ɖ�M;�k 5x�P���'[�[���i���&mہ؎�ҁJ�Y�^@�f#�>�h��<,O��d�O��D�On�D��W�\@���N�:C<��0J�?Op
��"��O��D�O ���OX�O"���O��ǋF��XX�tGC�x�Z��T!�k��ɣ֖�X�	�`�IKyR�E
Q6�1f�=1�IS�����Z�K�6��O:���O��$=�I�f�ޅ��t����ő
gt�p�Ú/{�PU�'%r�'���'D�Dڸ3��k?#��B��T�d �T��F�^٦U��Y�	��P�I*)Դ��V�/��4r�
GK�g#�����C$oW���'��\�0r�$D�����O6��������8�4E�&���`�@ʂ�w}��'���'LޙY�'�b�'�Rן�6�
<�"�^�}-��z �}� ʓ-������i���'���O��Ӻ3�f�?((u����y4�CE���I�`�֬n�l@����8�S{R�13gV��T 6DW1c�`7M��%gDaoZ�,�	��������d�<�B�e��4�Ì<5[���l˩H�&-S�y��'q�	r�'�?�7N�$�j�	�h���B
��3��'��'�V}y���>i,O�����2���?O�qR��)T)q��{�~���<1��U�<�O���'S��1+�6=坈p���*	�U�7M�O�بN
w}"^���IPy2��5F�I�  �X��6l
D�uC�#���Q���*?�!��,ۢ�r�g�`Fās�BD�1R����k�H��DAR���PR�N64z  Ĭ		dLҩ�E�Pџ��!�Q>�Mrb���:u ,�>�2��>�Q2���qĜ���=�0�1�Ǿ4Q�9�޲G���a1N�.���Y�>��]XA�ۤZ\����5dF�H@�Қ+�F��b�MB�	�#G��N�!Ȱ̉�ц͒� �4@��Ac�M���P�������T�sݬQ#RIŐO�
isC�̮t�$�
�2��cdB�\*�I3���[غ)!^8�?I��?9�H��(w> bF-fKX�pC��#g�f�Ӝ+��)�/��
�z �PN� *�$�<!�Ό�P(�-� :����Sn���(�b	�7M�Ayu�� �Б妗� ��<1@)������x��C���9��9,?���'��TI���?���,Y0H��ve�:@3���U��+N<�0��W�22����6���tL��<y�
��r��	��O����'��'P����Ǽ0Y84)�i�0>)��D
 ��t
rCO�j�֧�	+��O�%� �K8
����(>m��P#[�8�n8�#�M��4�O?������	�$�ʸ.B���u��*� !��O��D??%?9'�ܫ %�[����+B�\7��(��<D��Ƭ��^��u��`D#5Ւ|!`�'�P����z�%94�:~Rԙ��P(@�N���?�ӏ��ℂ��?9���?������}�l�� �<|�J	�0m����0�)ߟ��$�Y;<� ��h�E���%L �e���y��3|sR���ri�M��I��.����?�=a�&\���&ϔ��.�r֍�H?��  ������'��ɵ|I�	�d�2$ �:aeU�M�0B�	�2yx���1��s1D��`�:�����?A�'H��P�e�"�j��R�|�d�Aŉ5+�9 A�O��d�O��dF�,���O��S%��xo�ş���I^-0B�Js�I�V��036b5�OܝЪ�>�dN]_F��p%T�jt��W]e8������Ob����(�t�"Tj� �����H��O��d�O���'\Z�E l������`�@�B����o���"đ:w(�E�� 4B��Q��	`yb��#�x��?+�p�0"���"��S�e���� �Մ_����O���H�w��̀Fg�,NyCW���' ���i&�ۃ��
E�׻Gtp�Gyb�Z�5�<|h��>�nk��� �@�G+E���Ɋ��ӑ���F剐k�^�$���������P��с�QF44Ic�Ӌ�yb�'�}���:�:��-�Y�!B3�T��0>�s�xҁ�U�X�x��N"���	3/A2�yr��[��7��O��D�|�%���?����?�#�W(em� s��?6����\7բ5sՆ��"3�MJ �5+MIq+��b>�D��_�z����P2�Vt�ĺ��3A^<h���T� ����'lD�`Q?�d�bXL��Qp�X8�@�-R���E�OFc�"~�I���YR/P�
���q��D�B�?	X�j����J���^��"<	6�)���Ӳ&�T1��N:(���#���?���;��"���?����?9����O�.؜|�r��VT��4qyj�ɫ[���@ԄQ�K���cT!8�y�	b$#{a�m8,ǀH��$蕽z����F�+���1��KF{Ri@r�
	h�_���́�l��~"�@;�?Q�0J�r'��ބ�Ԍ�R�q�ȓ ��s�V�����@�)q;\��)�'_t�X9�isZL���F:U��O�K�����'Rr�'�������'7�)Q�zCb7M�O�ՁR�".��(ӠE�>�4����'V8�C�]��T���-T��V��5��1�9�OЋ��'�2�|o`�rg J# =��#�ri��'�˟�?�O�䘱4�?Li�f�<�����'ۘ���ɉ��h@�`δ(��;�'qb������̦e���`�O�&�0 �%7�졥�\����0�j=��'2��e���T>��d��>*=<1@�U�h�T�k-3�E��	F�t"��'��+���OG�e�]��Ey����?�����s�ȸ��D�>v���6h[�[Z!�$��O_)ö]���2��RRa|�`*�$ߝ9FU���5�M�f��W��fYm���Ir�T�J;�r�'��F�rwtUQUF'	�� xSB
�
y�H4�'d1O�3�C�+�!_D��V�^k���gN�!bzJ�Gx���'�d�� �НmHVqү��=�\5������O�)�J��S�=hc䏴m����"O^���耜27V�ۆm�7�֤�5�	%�HO���OR�f'ͧrZBE�d n�`��O��d�<h^j�F��OF�$�O���R����Ӽ���>����,pϬi��lVd?q���d��`Rۓb���ӡď����ƾj��ke,aӴ(���'y!|�6g������(g�N��5�w��{��<`���ݯY|R�'�f�SEEͽv�L4 �`ʤ$�\�'�BJ�7S>)�.�x���p�߯k[�#=�'���b%5�i����t㟑x�yaK�1^�YB��'t��'��A�d���'(�)اq,	@��C5d�l�"o�4h/��8��P�!7���G*�(�󄚉XF��	"57��9c� I�ұ�tɋOYh�EH���$KNr�'�B��%EG�Qت�H��6w�b�'X�OF�}Γ4�����O �M[��W=Ck(Ȅ�	~�'�@���"�\ȹ&+k��PA�'�t7-�O˓s[\�%�i���'��Ӟg3B��fv�32�� 6),m�Q,ܟ�I�L
���ϟ��<�O��3Gn=G?�Q���#a(����Q���?��ChN�cv��ȗ#�t�"�H,ʓb���I某��؟0�O�U�ǭB�������-F ���'��O?�I!^�T�q� &�����1�6����k�I�bDPI�4ȑ�/ z=�0&��3Y�<dq��4�?�����IϷk�
��J��'��p�C��oϐ� ���
^U�d�3��oT�y�ʅ�f��A�� Ȧ�'��?�cl�(^�m���K�Rܲ�H¤8�������V������ȰO��LF���V�$�+Ѝ|~����,R��^�Y�N�?�y���'�x`�cnEp\����F�IA
�'
*Ʌ� �	ެL�g擇@Z,���Tz���I�$W���j'ƃ'7�|�sI b'����O�,��'�7AW���OL�$�O�x�;�?�;u�j�rV�ͮT2	#
֕s��5�y�5��I�<���䅇c�ݨ���1,Ȩ�	�C���Dί!�I)e��?r��B�DSf��J(���'0f��a$B�`Xƹ��)��uٰ
�'���O�d�U1�パ�f� ӯ7�S�O�1�@`x�$�)��	�[,��R��T(Oa��Bd�O�$�On�d۟ZD0�d�O�瓹x~��F�N�2B���n��5�7XH�tbc3<�D��˓?�H`�UX��a4F��VWL<�s�4_� �N�t�}Z��'�T�a��?� �K�ܕ���	p��(y^�|h�"O%[fi���-z$���@1NQ9�"O�Xc4��5]��̈�P�ϸ$ٷ5O���>�5��+b��F�'��V>��`D�e��*H��nBa�ɢK�$ ��� �	�7�F��IP�S�DG�m����S'Œ*����a��(Oxu���G�M��.�.V�	c��ڢ�<q�-
۟G�\�D2u��W�,�䔿[����ȓ�z"�T15Z`�;���9 �N��	���x� ��IU=?Zx�cA�I7�xy�N�Tó�i'��'��m�������@�	�"����3+�'zs¥3#��A�&��,��|�<��On5�[idD0 ډ(���Մ[J"@Ӌ���O�� ���!�`rTbϔݬ��Ԧ]pd��#�)�矘8e
S!G�4)�b�;,��]��H&D��C�L����Ip�_�7ǀq�� Qꑞ�'mNq�7�U[
���Q�����?Y�n�'��Pz���?����?1+���~5�QFB����#DG��yr�_�(����
	#.��2,�h[*\B��#Db�	*���Gcέ�<�{��*�^��$�S��D=peX�!@������?�����I}�F�w��Y� ��ny��K)d>���pcA�8��AC���0<ى�D�gX�t*��D	� |����6p�jl�$�M+I>���?A�'KD���Lg��Q �3h���bՎ���SSLß@�	蟬�ɝa<T�S� ���5�XA0�DU��䪔#W�� �8#��`?�9���3�O
ya���^��eH�aډ	������<��bhO�<slU�S/PX� Zץ�O���_4H��dc�6ON���J�+_�To����'��?!��b�5y�H,��OǛ-�6e�.(D�`��`
�>��*�'�$y&.)BV矌b�4$�^���GG��Mc���?�.���)ŮB�g�84��-	� ����!�)�2�$�OR�d��1x(�#�|����E��YthH�鞭౭F�'�h����i�93:q���P!;�>!�A�=$Q���C�O����O<�D�|�f�͠]�0��z_$�zg��?y���9O�XP�N�?"�'��t��8��'Ol���l"�$�K�4T`=�A=OV���¦���ǟ��O� m�u�'>b�'�9R�)�6��0�e*CVEZ �b뚹�J�zQ�!�T>i�|�I�5�n9c��3i���C�[kܕ�A/(��*M>E���1g���� ,|�n\x�/���Sf)�?����?������rO�,��a�p/6��{Ƙ�I�����ɥ u��8aホ����5 �0/��#<��)�� X{妈:�+Y�}ʤiq�`E,�?��� �0�2"e��?���?�����Or��/,; ����:y�N��d
�w��l�qͷjϊ}��
��J�ʑ�;�Ē��ޥF���jR"��k��u��� t�8�k�(P�"P�a;VL���0�Afڟ­��U��'^h���6:�Zm�S ��Oz"�(��'�Zm���'a��r��Y������lZ�P&�� 5II%9j����-
L��%E>?�ߓ{��ٕc�$E#L	[��!&�����V��ᖥ�&�M{�S�P>Q$� �M3q披)&��@��O}��'jI�?9���?y�2d��$��� p۴�?I@�^?Mt�l�t�-}��1d�U8���E���E8�Pa�	N�Sn��b�B.dO�hui�&$��
V���dҦ�;a"�%=���#��GT�Y�"nΨ�M�����d�Oz��'�<M���Ş=\]+���4w������?iv�G�Q{&L�C�k�:�K@��<)"��$:=�&Z��#��\��u��'��R>�C /W�h���aw��UE|���ۣur��۟���$r�~�kD�x� =�o�E����z��ulo�*��tI�	?��ͫ&�	�P�}����N���'���T�O(Ԙ2�H
���S��=_&����$|S��k��$�O�ʧ)���rr� C6,]0�f��B
�+��?����?��|ʊ��\�8|��nV�5<y@GϨH�a|&<�^�Z���[��Z&@�yQ&����.(�4�n��T�	w�D����'�� C�F��TR �X٘L��kڈ\�h�,˵w1O�@��/S�e�q�K�:_4 �R���!����a֝*�<h�y���'��D��K�.X0��U�K��]	��j�"�'�2�'�?��A��q@��C8��M��Y�Ly�$�Oz��D� 1��㋧�j�D�عD^������۹�~Ҳ����b�2]��	���O!���'4mS�ή��'�B�'����Ɵ��� ;��8
#,�"}���g�)À�ɣ�N����\F��(�B-�d%9�%c	vC�lK@���^�Y�d�+nT�P d�-0� �3ړy���2aʵ:�y��KNH����\����?�u���,O��d�<� 6	H�'@��@Q���&T=Ԡ��1|O��RC��4�<���Ҧ�� +V��I@ߴ��+Ą��dyB%��eM��]��r�RPk�z���8禈��$M�������ȟ(��B�ǟ����|�e@w��1�*^�!��2"ƕ045���W�śv5�1��$Ӷ��<a�aH�LP�j�$Y�֠:E�ʪR�l�1���p$�FO�1��<!Â˟���ӂ�:g`2t���� "v
��I�'����?��W��@ʸ<�-4 ��ʢ/9D�h;g�7��c��!�Lp��Ba�,��Oʓe��C�i�r�'A��i{��Q+���v��2e�@qR"���,��Ɵ`���;��xjR��K~*�T�s�AZ�X5����5(�tm���	[ �,r𥗔X�PlⓥV��Y0B�ۨ,�*훁�")8Ң<��#��������	c��� I���ڐKBk�"B��K*�2��s�T�q��4w����7� �굨(�OB�'�<
,�����	�!ӛ���U�i��X���Ms���?�-����I�OT���O6�z��?�2x�W��d�$9j�d<g���nF�S���d�b{�5@��;vt��7���*�@�:��1�)��ةSB	dm��H� C�=�Z׉�:$��i�������_��?qD��hiÒ�G���s��<�����>ɳK*G�xѕoU<n��[�`�i�'��#=�+�"`b�G�b�)󇋪!��p`��O"�dЬ.F���%��O����O&�D��{��?!�1yOHIzԅ�2u�Qa��a?A���zx�`��A�3�r)cVf�+0h8I͡��@W�5�Oz����4�h��Cﮱ���O�`���'��{bF�(0�
}0!���M]�#7�F��y2�ٴ;��I��@(A"��r�nUk�`"=E��E�La�7�K�{%�!y�U�Hx ��l�3c��d�O���O���4��O��w>�a"��O���4����ô@����F�5b�|2�հ��� 7�q��F4p��G���)M�|����?��H(��{m٫K�\��D�L�P),,�ȓ~����!KW���Tc���,AlX�ȓ'�K�h�2K��$;��,7<*��u�OșѢhݦ]�I��0�OúȘci�G���V'[�Sv%��޲9�b�'b�Z) ��������|"�+�(� �5�X�M�v<*�+�J�'���,�4GD�D�����^<,a���T��$���(O��[��'{r�'�BY>a;AO˵�
%��j�6��3/�<�?E��')���w�G75�U� 5sp�p*���'�H��hM�
 1r"'�4�P�q�'`@ � p�����Ov�'r�8���?!��|�c%��0d= <�͒�i���I��ũ�?I�y*���#�E�RT���	ŊE
�<jP�?[���Fx���'D�Y*J&�<��0�$9��BD�"(��'���N#|�I!{4��Ǫ����ؒ�<���Ї�I�A��H3r,�%�������DXn"<)`�)�R'D$N�u[��ŝ_�6M�2��?)�jF�mQTd̔�?q��?!�]��n�O����0,�IR��W�!D��a4nE/��$�	j����D��A0%Q� �5s74�#&U��D��3)x���ڸ+��HI3"E;R|�)B
Y�[��$ʚ�b�'��'��'��9;n��d���!��"�̒<��C�	T/�9c�%�9��UZ�<.�����4���ħ<��#�#��fn��1��p2�I�9iX��3� 	����'���'H� yq�'�b8�d�v�����R�f��(x���_�1�$J�#_
���JN_X�@{ᮙ�q�ʀ��Ì�*�"hbo	7ق���\��
��<14(����� �$!��VX��r�M��������h��dJ~�K�*f�6�Z�K�h&ܙ�	�'L�h�U)^jn��e׉�0�[�'j<��hO1�`�1q��0 �V�uDT%���y"Or�#�+��q�E�QYc��42�"O�j���ZyZ��Y�kx*��u"O�u�؇T�ER!!�~G��9�"OFi�N�&�����'U�У�"O>���شI�	��̥v����"OBİq��13��Z��Y���y�)�2Ǫ ���
72� �k�P.�y򡛈v��pi���*�P�$����yR�@3��L*c)X�P�P)���y
� �]`U-�Z�8a_�nօ`�"O8��7 Wei0L�ω�urj�S"O.LpC��X�%�/}��E��"O�h��u��ِD˙�7�qc�"O\�ꖮ�>;t@F	�q��"O�8�C�ݰ��C�n���"O��Q�Hۨ^�
b��+>�8�`"Ox�ޕl���g/��
�B�R�"OЕq��1 ����hUC�"O�av�Ǥ5���i����Lzcf"O������9'����</<���"O��G*�u�,M�՞6@
b"O�q##�59p60���v��|�$"O  �G� L���䠑L��9"�"O�I!d�ԝH��A��eI8�"O�5C�ȲC���ua�w+�x�&"O��$��7�6H9a�R�U�d"O.0cteȸ���Ǝ
@�U�p"Ov�Dע,S�#䌌h��	Si�p�t,�6͑��������j�Έ�p�.�kD�L0�#\�z�bع��n�a��O�aV�M�Vn����ñ���MK� 	�<).O��(e� ;�X\[x�۰�>y3�����$��+͂<h���&�v�pҥ��nH	{�>�K��G�E�xѤO*��ҥ�]"�p��/	�$'�px6��*h�Z �!����!Hv���p<�s��Q]�Dd]�dA�%�6	ۡ{G
 �H���tIlI*Q�̓F���D��e[:�{U)�|��Pk A8�L���)(�����٥7������Mc�E�=��t���0�)�����t����U�~ �3�ȦG� �:��Ї0cNP���'G��n�)
]~�B oƦt"���j�C@f�C�C6,߾M
�O�8B�+�:�A�reC"z��Q1d�d;� ���<����"�:�Y�HI�#�2	�6NY����G.ƶ

@u�oe���lZ�5����A@�[fT���fi��q鞥u����N8x���r�P�XXc�^a�'�����,`9�b��8���*㈘�
�`�X�
�3n������n�1S��YH�2BőQ}�O��\���Y�5P��6a�<9��'��%[~��DMqP ѡ���#f����/��� Y�L�{�.X�<�(�S�S�808m��;1B�����;lq������)W*T)�k����J�.2j��S� �n��!�NZz/b�b�P��0���3Z��9���A5��+s�E,s�̰9�-�9�Dʊq� P\A�̐���'b�R)��Dڪ1n�!RXv�͒���"JB-k�e�:s���c6
ڝoR4�3͕� �:yS#�"+����)U3zS\X	��p���G} �<h��`F<B3�P��W>�yb�)v�`�!0��>|䡂�l� �G���@��@��X3�PEp��M`�
�C'#��`��3G%�O2E@\u�lp�E[> �D��cM��PC`�SԤ�ATB�m9�	 '�6�'pSb��w̌L)��9R�`U�+�_��Y��z�EablZ!u���ZA
ʠS7�z�I� ��Y����O�L�B�R�!�
�B�"m��_zD�`$�	���R�>sV�г��86�VM1�\$]fQ���7o�+}��a�c�4��d��S�:{���G��M�b ���)I°0;�"�~|���p$�\|�� �c���F~�gZ�5z���Vh�,=���� �������vȫr�V�@0�=����9`�Pk�b�ܦ�
��'��4Z���U?\�bы78�iK K��i�N�S��'d�$E��0t/�MC��'�>�q�Y��,,s*�vy"����0ͫ$��ٰB	ï�M#��l695(H�C~.E�0��O<�)��'�5 3��7S�u;ōY�V>`y�$I	`7mK��?�P��%g0]��) �k���a��AC W m��N�/�jT�A]������қ��O�]�ѫ��Ib�E� Ǩ�Za/�7LP4��
�;/c�C�
��i���?1S(ݰs���jE�7���9�hR��#%0l�!�F� W��p6(X^��	,m�j$��n��IB�ā2K�6��F�G�k�F9T���u��7��t`�c�^��g��(�J�xG�\'�v,�`Y1v�x2�8��D)䙉�E��*��c�<բ���D�7*�8������O�8��Z19&6�p��4}P染��>�5Q�����16�$¤�G�9z� �"��d����DG����6M
?>If�E�>C����!ѱE��R��-�%rİ3� ��I�B��V�x�� i�D��g-�L�2% �!�7���yjS�/V�� �(u~��@�!M���Ir'��ɥ�_g�(<�M�r��>Ʀq8V�B��Ĺ^��h�S��J0᤟uAi�S�䚦�)��<�ǳi( ��j�S�� 6m��'x�x"B�F(�I��S�$YѪ��CE=iЀ;�G��U-���RDKLJ~�G�> ��!�I�VK��IhR����*["!�d+~�����߄La��i���7����>9�M����f����剬&K@�z8�dP)�+h�e�� b7f����ɮo�eT!E�Ɍ}�Z!�$�*� ؑiF��F�Bu����1:��y��I?i��<� �RM ��Oۜ]8B��Qy2$K<3��AhWe�3_��	�D��8ò�17'�6��9�'�e�ajFh-*�r�#N�?��O�:���y܀Q�N��i#��`�����8� �pI�vrџ�Xw(Y>޼���O&C���#Х�GU ��ś9m~d3&�OX�9��9O��P�.�9i�l�`�B>�x ��/Eo��$��J�L��T�����U�q�� *�C�a=�E8fJ�<E�R|�ԧQ�s &b��k��I�f1rQ曀AĬ���D�L� �;��_�^��O����G�/��JJS�2� ��Q�� lH0�v<�3G[5|" �b�~�ʸ�Bo�S�>uʹ�Fg߳x�T�#
�F?*��'xt	��J���&8��́4Nb"��O��+diITa�#kXI� * ��(��F��dU�9��'���~ޙY���7Ap29ʱ/B0P\Sb��O~\Q�/��Xs2B��a��x�A*)l$BA�E �:@�V���]��q��O00���r���~Zw�R�J���@�U�6�U=+�,I����;ԡx&@�'�,�Xƣ��T"Z��E�'p���k	�f�R�jaN�Q ���ǉ�uhlx� �d��)�Yܘ�1�ߴW�Rx ����U�DԈ�P��������@F# Ձ���/(tx犗&b��1�ө�4͸'u���Pb��|F |C�˓<4yS�ѯ*m6H�e ʧ=����Kp@��$U�T�N�pcF���)16_FB����+g�vE����V�pA��,E���,�Ԓ1���v���l�5b=B�`�gPYS�Y��hG�ZI�\ �'�v>�Ց7���o���|�Fl�'"w��3&[�8�p��S%(D&y voC�$��o�8~8t��ɤ81d�c+��U��V.0o8L�G-6��IXg�V>I��dB|��y�����$kN"/��;@�ՃLK(݇���xq{��&"0�{��-�vd�ƀ�O i ˪wk|�� kO&͸'>�m��/�F���	FņsJ0qH��
C�`!� 5Fax򈙫 
�T��(0��n�	EP��LQ�6��b�	?L"� �!"�	Q�Ł). 
���g�6���'V�M��
�B�zԹV��n^����O���w��=O<y Aϒ�I1�@�ET�p��-kj�ű1��FZ�35^�+l��2��[��d�������1n�z��$ӸZ�dF!�az13�M�u貌8�)V��2�p\���0收xنP�k�a�;��$ᰬٟJ^���I�e|x�gA?�O���B��o�$Ԃ$�@	"����[x6!PJ�'���J�'��;A˒!a��܊�C7i�d P�HQ�EcVZ�'�f�;��'bp�KW.�zk�P�CoN�݈�C5t�N$y%�	,#�Lce����',������**h��J�B�3b�F��J��P#`D9v.\V#�n��M�a�*u�Fe�g�'�� 颅Ϥ��˓K��b���� M�s�MR�n�b�,܊�i(O�Е�5O�ulvQ(��ҍ(�x�$T�Z]|Ӗ*HP�<i�n��,D���4�=)�j��RDȤqe�R)p�r���dט2.f��̘��=���Yv6���� n�� Rg��
��\Is��uܓz�$Tj��Z�+������<���ZgO�" �ι �+��Op����)�?Y�Ǝ��^�qT��k�-R��H�0%DgƖ	;C�o�%BΑrţ 4H��'!ҴP�%�x"!i��'g@ip+A V([J�R��{v�'7bdh��!t�D�c����ߵd��}���y��	�!��\I�gʗ~Q�9�CHA�'� ��;)�N�9_���qw �EqΜS�~�N��'9�)��9z|��@U-H(R#:�P��h&�E{b�?{�PT	�ĨN�TA)B,��?7���&�Q	������P��&~�z"#!�4��s���*JR�J&�Ū���q� NC��I����<���8G���3�ሴ���I"��O�"<Y�/�x����e��^��d�,J+ɸ'��@���=�`���k�x�8K>�Enۜw��D#@�[�GP�qH�G��d��{�C^,�U�?�F�ԗj����>YrO�}���r�'��;��� �%��ew�=��BG��	���_-�hO@p#8�9{���_8 �z��ϯ.���+$�|"�ߏn���) ��S�DƝ[Uj��?-�����8��b��9I RUx��$�%1�0�єL��!#P�J�����$�����J^:zb�问%mi0�
���8++�
R�@��O䤡(��>iQ�.O�Tq��Z�s&N\rԍ�/(���P>O�t:c��]��
Y�Me�Us�K�7.�O�� g�6/��Hc�ʇ4�c���x�H�O,�s�. ;���mӲW�LY���xr�6)RIK��-h  ,N�+��m�*��P� �q���'.J�O��(�K�{MR�)�JI.J��\�&lبB�5��,��b,��p���(O�$4��PrM9!������o�U���x�n����b	@����Πg�y��G����D�XS�xRH�y�S����� �-�J1��[p�O��*��<����8�.����:x^.��p��az��1�F��S���v��]`��>�	5��(w���	�!����M�iԺ1VkG������L��c���=)�o
�.L���UfQ
l��<Q&�A?��Ȁf����məo�=ڰ�,��j�	�L_���?ُ�IE/H����(�P��"ԈI=҈�`�@؊���[�B���KU>︧�AZI\T8FdFUK��:Fa��V�
�O��8Bi#LO�|�a*p|��ϸS-��j3/�_&��{*��	G! �1'Zɋ�ޟ���!�3��0ҮX��@!�7F��b!:g��/cm��(��O����@$g��?�KR�Q�Onv�s������D!u�t��n��q�ډ+��[��R�I���O�1`��z��8�"eR�!�j�i?yC��7iȑ���	3N�Ʌk]��<� l�:�oJ�d�kwG�}���֎Cz��$��6GqOZ%��O�b"����s�A��]�`�ӳ���d����P?g��y���}�:�H"��)��g�S����_��㢎o���C�٬�Q��8T��y�ᦆ,/-���&���G�/�5r�!ǕXX8��rgB�]��n�S�4gJ�r]���S�n��$\�f�rx3U"!���K�恘YVµ(�$��2 ��H�t���a-L�&Er�T>�'�n�z�%I�&8*d��������P�'ݒ�k��R�KZ�+T�[,%An�x��d��@��D�E�:M��!���2�f�I4ӄ���H?a*((�4irˆn�����4���LB�Z�X� ��PFD����R��1Or�ADR9�yw�8T�V��Q!`MzL:��5w�Aeg=^�` Ҭׄ
�Pa�Ϙ��	�.Zl|0���lA�����	
$`�<��
��|1���:,�c>�wO'1Z�ej�̙�O�
	�'Mª0��u��T>���@���G��<�X4/퉴�K$�`�T*�*0�Tw���K�E���_?�~��D��p �։�>(��3T�@��0�sdH��~e��*�ڄb��c��@g���	C�$�)g�p�)ׄ�H����y\�W�6��H��&AI�Z��%�	'p�iW��D�s��A�7A��zX�)Q�d�Ţ��)}��� ��I4]p�Q�D�E  ��;S�XQ*�-ΐu)��""�����2a��Z�[�J�b�h���|F|���c���H"��)¦�`5�?;�剄g�d(�v��6~���!��H>���D��)�XL��ן8=�U=x
I2��ٞ�h�AG��#n�X�A�������[���:�~�����'D���j��SO�98Cj���#��e����`�az,��Q���~b���;\�8 ���rw�Mb�fm�<	fʓ�L�flÁE1�'��R�mS�q�~��,�[���r �AU&��0L�i�a�� )��,Pm2�s�0#�/�&
Bݰ�k�\�@��cb{2h�d�>��� H����A�bO�|q@�Z>���W-��8V�7G���!��Z�;U�ȉ'HP�!e���+
0��T�U�0h+��?���+�HdY��I�	���%=���[��X"f#�){�\����	m�Dj���� "��!���څ�~��P��,�4(_����äI��0=�'\���'�fm�SaH�N(��� d�S�{b�L��(	2�S�d~Fۖ�F�s�}�c͜�G0\��b��C�S�7)tY �N
<x�5�R�ۈ0sNC��70b,���"�rD �X#Z*|C䉡o^����MǬM�d�����/��B�	��̩c�.�b�hYSŜ�%4�C䉙g,:DY�e�>"��sS"ז'?�C��\?��Bl��!p1��)2pzC��(�]A�(ʭm�E�$�Z.�C䉌8�L]�p�_	:���8en�>B䉕<a̰dMG,3	ReSG�PyXC�	:u�F�A�(�&
*&5�d�Gt� C䉈O�:�"%���� =�W+E�21:B�I"b����F�+ځR(�/P B�	2-�	�U�<@&^� q�Ȑ�C䉨�"l����3l4�{Q�ċS��B��*/8Px�ƍ�� b���cD�K�B�I�<4�	���!(���A����>C�IvU h@G�WU��0E/W/ErB�I7_�}S�@'1����T%�B�	2mwH�P�ث"�t�	\z�C�ɵ&n�]8rl��"3~�S�+ʦ4�C�I2g})U�ȪE芠3�'H�in�C䉝Đ�b	�h�ɂK�Ks�C�I�E��������{e&�A�\���B�I�.�%k���y��Жf?ŖB�	\P�<Ya��y�4��G���tB�I��9�7��G�h!łH�i�B�'@.։0��
������ ��B�	't\�� �@N&pܼ��O�rB�IK;$��
�z��L�U���1�B�!�~	Y�֬$���s�%=BH�B�I�3
6��]�dp� åi���B�I#a�H8��M$$F]�� ��hY�B�	�P�,9��A["�Ih4➣=��B��@��X
�����: ��ێ�hB�ɃN�nc��^�(�█d�C�	!.b��y��J�D�f�w%$Gh�B�)� �)�4J��(�q�U��#w �"O(�;wIDBH�H�.[�)ZV"O�#V�X�=SDt�T�O��D��s"O,t�Uȁ0d3§F�3����3"O ����F�u.F���G�j��eR "O���Єe�Z8�w�G�\�:u��"OH� �ݒV����(��R�)2A"O�ё�΄:j�{0�ۂ���;S"O�����	�A���Ig4�e"O��0���[�|�"�$ܘUTB�"O���6C]\�,��Ϝ�A�v"O^ȑ6O�>�.D�v@	cpM"OD�`/�5P1�1Yf�(YR��9�"O�����7"�`��Q�F� �"Oօ��/�\9��	�: ��� "O %��둡@�1W�3"����"Od��ƇA-fJ�&A�7;���"OR*NF�P�� O�}�؈3�"Oƅ1W�^�7[*�ɰ�>1�\he"OJ��r��9��I��E&8���a�"O舨����>�Hs�LG�#�5��"OP�s�G�r ސ)���;s��0"Oj��a�A�w���;�Ф5n4L0�"O��:Ԇ�,QD����
�mN��K�"OX�2�l�	I>�8�G2mHB9av"O��J��	C�#��E��`�[�<q�D�)%ٖ�0�	�H��I�`��c�<�c#9g����o�
����p!�$(`?��+�&� V%�(î�\�!��!]4�x�@��2!�Y�mH!�:VijQ��H�v����5��>;*�}���`���c�6H��j,�f��k-D�a��5��tB!T�J�	!�*D���N�>�T����:qq��z�n'D���,vN�ubd�9d�"ͫd�%D�����x�<S0
�� *�495%(D���D��$+u�ٻ��W�B�ɘv�2D�X���[
��@Ȅ�ԑJ
>#��5$�X�6a��{�����Qiޥ����y"�ا&偄aP%v��p�A.�yR�1=|�v�Xh�m�����y"��u�T�Y�E&Y$������y2��I:}x�i��J�o_��y2��sp��V�j7��%�T�p=�}rCS�V� ��ȤhE�U2��ɒ�y�D�?� I��	��o����%��y"�)�~\0�c���D|��9�*4qB��ȓ	iH�û)$��M�@C̦8�<��ȓrb�Smɇ;���p�R" 5t(�'(`�Fy��)�$ǈ@&̷��0k�M�"7!���	�|`�e��^��|��A 0!�$�!&�^ rV%�Ib6�k$��M!!�dğ8�Jl�ck�5YHj���f�11!�w��5#ϋS�4�)���Q�x�"?ʓ	��@�`��M(n�%��)V���;�8��Ba^)�X}���̥.<Z ��^r���3���\:�@�S�لȓ���B��Ur�����_hQ��}�ذ1煐��4�F@T��9�ȓM����
 "̽H���#I7B���H�zB��`JD-�]F_7�`������䆒�u����J�8��e�ȓl�|%��f>p2���׀O�g�X�ȓ&>��ҭ��>`;'�ԴT���S�? �����v8��Q�L�MɌ�H$O:�Rʚ�q��`@�</n�U�v�"D�9��\6J���r�
Hx1�t�?D���ܟ�jI	� ՜K�B�Xwg=D�$C��G9n��H�:Mb���(!D��1a��;L7��2D
	I���Q�"��ሟ�����Liȭ*4�7!Z����"O.��E��31�y	 A��h<���s�'[�ɤ2Y�y�1	
[�4@��E�/��B�	�X�a���ߗU���3�C+rm�C�I�YͮxB2�֘|[
�cł�8��C��]�e���XK(T��'�	��C�	;CR,����[336�m����E��C�Ig�<r �+ǒ͛�E����	>'�ɇ�I�	
h�"EIT���ˑM+p����!��m�w�H�cK�Iu ��CIH��q�p=���C��Eif%I�$�|�S��$j��"=y��O~���w�ҵ/� ��!O�D�rI�
�'�H�檜1B:�@pB'7D� Z
�'p)�E.�y"���.U���	�')l x�#G�?A\k��%���X	�'����GOM�S˾�`�>�.�
�'���!&@ŗ ?�e�&�$`�r���'�:�0t%�Q.H���KQ�ZDVL�'�T���cN�9��=K@A�=�]c
�'��e	l�1������
+Hn�j�'����/v�b�&�
- ���b�'g�d;g*ǎ;wʬ�$�D."�89�'}���q�{P���C��k�t�q�'ب�g"�F�B0ӓ�9c�4�y�'�>�#Q�
�l�l0�#��-u
�p
�'�n̰��S�i����
@�q"��'�Ƅrp*��=����5DX.O,�=E� I�-N
�yc#����z O��y�f�<���""�L�xR���"�y���8~�
��wL�{q�m�V#��y���~oF�*vid���e���y�FR�d% �X�Z�ӄO�2�y�@<1Z��
���-A`�dX�k-�y�h�8w]|��b���oN�<YfAJ�yb�>J>�p���eU�[�N�y�%��V蹥�V�)T̫��y���\�	a�C�)5���!+ٓ��=Y�{�/P'n����U+E'2z�C����y2�[)R}V`�)*B�;PMZ�(OX���E#��T�����}�b�Pjp!���*ˇJ���጑$9~��ȓ������� �b��T,�`Ą�Y��JV>56ݪ��B�m��I�ȓj�j�RBN'/p�(3��}�z�%����I�g"D%� ̛^ �Q��B�9�v%��#����̲&�1\��B�I9(��uF�4d��Q:���`�����-�Ě)
��1P�͋�'��0X,�!�d�C��A#�-&�VR�l9c�!�$ŢJ�P�B�ݚY�L��w΀�!��Y"0�U�D�Q&A��dˤ� �7�!��$P�Z�I�m��`�)B�7�͇ē ��B��Z���I��,�|]��	a�:m�]�mN)Es �aGАfȓX2�)!EO�
v� 1��&XT���ȓ.��C��ު�� �'� 1pD���IaܓF͂��Ⴈa�N��� �P=�ȓ'�r� �k��r�Ti3㌪"k�=��S�? ���A�EU��0�`�
;����"O�eba�/+.vEiA��,y�1"OJ=0P�K|q�o8Q"O�	�LK�&�$aA��ҡ�z��"O�{p�X�8�x�R�M?YC����"Oԁ;4���N�^8jD��@)����"O�l���VS2��T�C��b�"O�LkU���G �:G�<N<튵"O�� �]%s�"���M�;g�
� "O����4�X�%#�8r*���q"O<[�KП&�	b�h�r)�}
�"OhР�B��;H�{�g۲+<9v"O4�!�W_>rmAE@�t1��"O
�XB
�|K�XH�Ձ_�,�0"O&�hGgF6��X@��۴D�4���"OX	R��S)�y��S�xPFb�"O�����	9Y���&	�3r�p�"O.)����12&`�_%O��]�"O��a.	8|^8K@��I�J�H�"O�3�M_bb��fD���Y��"ODݢVneOJ�2í��eǮ�'
O�7$\��I2k],��(�K	O!�P�$�T)����.�:9�6̉"3!�d*3?&�I�j�*Srp!�Aċ!�Y ?�N@z�m1j���D�B0�!��_\��zU�
>[c�l���*�!� �L<�c�FR�WH�m2��ϤCX!�dH-o�Jh놅�oC�a9eȅ 2U!�D�|��2P�z94�1�P�$!��M-P�I�ϟL���"�U�/!�Z�#6FE��fͶS��Y��䕃i!�ā�����F�](�4Q���&!��A�#���3���sNԲ���}!�$��~\���ӫX���2��O�!�C/�f�NbvY�D�x�!�D�1p�V�rb��z�.����C��!�d	�Zl�R!��$��X+��A|!�^42�I:��[_ε%͟�=�!�dRW��)AI��W�|��,�av!򄁽L�zA[4H̺jN���L� 6m!�d�%R�0Rcϥ$9�-�-.�!�Ā�xf��#��19��P#�G�H!�Ѷ	���9�K��V�<M��
N)'?!�P.IO,-q0%Y�vhxI�H��z!���-�`"��Ϡz���H�&��9�!�䜕ys ���M�F��4�!��^�$�@�1ϓ&n�e�	�y�!�d�?;�zd�X.����f�-/�!��"�� ��Q�N� #�8]�!���F�D�媛�7�f@��R8_n!��V_�IҴI�$!���"�$��f!��@�o^5aR��"�X��b"7S!�d�95�li���	��P�A�A�IO!�d�(|v͋AG�?�Dt�� ء.,!���F�����h��K���iY�\�!�$ʕ&m�@����a���g�,	Y!���*-���aG�	W}����DW!�d���e�VCT���Mū~G!��)n�0�%3�Q�S-E��!�H:(��`Z������a`�(T�!�d�������L��n��)��AS7}�!�$�y7����^>���%�+�!�DW����EY#D��P�(	�G�!�H�MH:�{��2��a���e�!�� P���o�mlX@�FsvL��"O�����d�[d�Y c�}A�"O�JQ���P��E�\��I�"OX�ֆ�� 6LK�˚,@h�1"OX)� q�Z�$ǬO%Z�"O��zU� �g^Z�8�l��r䐱�"O
���#G(<N�t�+��5��u"O�@Z �Ǹ����'+��i����"O � C��-�p�5x3U@�"O�1�B)6nR-Ξ�b"�ZU"O2�r�*v�<���+�=\�Y�"O��ꢆJ�� ���$�#3��%) "O��xa�¯%k���a�r/Bm"O�-�dȚ-��� ��%-G�e[U"O�l�g�__v�@a��R\���"O��M��'�|1�B%��}��"O2$Ygj�~����E�[�̌��G"O�E{UZJ��V��nƲ�2�"OnhKBD��Q1����O�?��$*�"O�����/2�=��� ��1�"O�(�m	TP�cI e�����"O���b�Z�d V<�"	�)=�J��T"O4|R��"#����C��n� ���"O�L�Q�ٯ}���ٺ,{�Q�"O ��dg
O�d@���co*y0�"Op��r��f�AP�̄�PlA�f"O�(LX�"U��R����Q]HҐ"Ox{������ #l�40���a�"O��p7L͜z���"�\06��\p�'tx`�䇗/�4�u�̧M�:�Q�'(El'T��A`�@��q�
�'����BA���AE��:B�h	�'����H:?{�b$l��5�P8�'8p�eA�hptyCDF˛1��,`�'M4�0���8+��P�/�+Zt�K�'�������0}��U��-z��Ȩ�'�&�Q M;vsS�A�w�(��'�n��n�:r´��eG�%D1��''��HV��F��P7�Y�$��u��'�dP��N2?��=SV$�"����	�'1R|*��<q
���[ !ڜ11	�'ϼmrR��?6h|{Dʺg�'�f�HUN�5����4%R��@�'nR�k��'mt�C��O�n���'�(A
�CUu�2�IU�t����'S�mZ�,H�x(���JC# ќ%�'�
���l͹�p��ƤV��Dy{
�'0J�!���B̍p�"ʰ��'��it ̈~��<�%��/J���'S|�p0X>':٠�� �n�X	�'����F�;c�Xh����i�ޥ	�'�*lc�B���8�`�g�>/���'w [ N5�`�sH����y��'{J �A"o����%��4�#�'��t����|���B�W�2|��Y�'�0�QL�Wl��.��,��'^Э�ek��y���ff�9���'����8�fq�Q���L:�'_�"`�F0j�$���S�|���	�'����_E���R��ݛaS0��"$D�LP�I	d~p�����=�:�ɂ@ D�t�c�C�;PWw3L����{�<y���.0�-t道@�P��ץP}�<�C��G�ĸ[3�N�4��l��{�<� ���g ��T����,�0~Ԗ`��"O�S��,g�C"n���X@4"O��Q�d�.�a�M6U�f���"O\�(Rf��!y�$� F(pu�""OP%� ܕd�ƨ�`^�+��yD"O6$�$�y:ش�S/��w�́�"O�['����pt����8XN��"Op	&�7M��:�ź"Q"M�4"OZ�c��p)��ea�4��$"O��1 f���P�.��]ڠ"Oe�"�k)F�3�!�4��iu"O4���I0�%j��7<�\�)�"Ol��1g���$���C]��"O8��b��e�2�I�;_hÐ"O�u��ξ<��c��]�wU^���"O�\�� 3�	���l�lp�f"Ord�ыϨC�"�P%`���""OL���.G�lT����ѰF���K�"O8c�=���! MS��l�"O�AЈ+
��Y�5�����5"O��:R(0�c�Wc Z�"O�)��"D�b���B�8kL����"O2���Z.�^Q�� Y|@
�ȑ"O�d���K�ޜ+�098�"O� ���~�  :�N=a�B}A""OZ�{Ï��3�NJ�sḘ�3"O��b�|T����<�x��"O�0�Rj
�M��Z�,`I3�"OP8I��i2��7YYl���Wr�<A��F�p3"��N 2�(��6�z�<A�c�V�A��	kj1��f_�<y�mρ`���$K*W�t�r�J[_�<�v��!u�X���%3�R�N�[�<I��-=�9!��B4���f��[�<1 ��7��l�s%���`y����Y�<iSn��d�r ��P<3��H�BYm�<��H 7�����f ����E^�<��m"Ttq�!� ����Y�<1��Ȫb�:��	���}xuO�X�<9��z�b�16���PH'HWS�<�*:��	QDI��$��@�W�<��d�SW�"7. S��ZƣN�<�B�D$sP� �Æ?�T��(�J�<�f�[�|��M!�o^`��&h^\�<���@�	X���%l�\�0e�Z�<1e���(���A��/ =>�9r�,D���0Ɩ�xIҡX�J�����@�6D��K��ïm�R��d���Yg�%y�m6D�t��8�����A�.F�̐��7D��)��Z=1�@����;KJ̀��6D����cL�k`��aD���<�Á/D���rO�X]~���Ň	L�`E�6�'D�����υ>�إ-�O���##D�d҂b�-:s� �E+��J�̃�%>D�p¥(��c���P2�+�H6D��	�V.�x\��"L�4�.v�&D�h[��q�ڐ��F�yJ�Y
��%D���D!�,5Ta�T&�4>��	j��"D�x��d�3�$i���@�~�Q�2m?D��p�G�l>|�Z�ǟ82��A��;D��y$�%q�<�A��ܹYf���o-D�j@�T8���C��8� �|�<u�&Y����&׹2|��p���d�<�D�r�yJǊص	�틅VX�<� ���	K���!�n,݊\�s"O�x�
�g~�(:&��;%�d�IE"O��x��4�:�c��K	<��5�F"O�-W
O��n��U�b�^�+B"O�K@�΂,���EB*t�튧"O
��u�L�6�ɢ^?�*���jJq�<�É��"�@s$�I��q) m�<���A��ف��<u Zlrm�k�<��	r��I:v̐�VI0RPG�g�<�0G�BO���D ���`@$�]�<	�+�'96ыB�F�f��� \�<�Ӳ�A��*A�|0Y5 ���C�I�v�f����6|"�hK�#�+/qZC�I�pފQ�%

:˒(:�a�i�2C�1k=���,CFzT��E��~:\C�	N���B �D�>��5�6m�xB��<R��0��%}�<���N�S�C�	�0?Fxy`FN/�:LX�;K��B�ɮ��|p4��l5(�3�ȼ~B�I1U�r�q�� e�%'��FelB�	5��y�@��]�vQS:puB�Ɏv5�}�&�˫&+�YB��E�L�C�	�~�@9෇��d�s��f}�C䉯��1�!�&" 6��"X8��C�	�� �rA�2��t��U�\C��9=7.����?Bs5PFg�  VpB�ɩ~H���S36��`��\��B�ɘ2�H�Ti��:��r<C�	:g�fm�Bț$��9�B��F9�C�	�d�qD�'6�0"��E��C�Q�P!cp$d<�|�*��?T�B䉧5L���E���c��9a��C��9z��P �JP�$��t����/�~C�I1�4�YQ��,��ࠠ"ǀ@�ZC��fق��B7�İ�PA�u�hC�I:�}�6��tä�AW&R,{E�B�I0av�Y�2@�47@��Z���2ӴB䉅$.uX� ؂�vEs��N�f'�C�P�½S �0�����aɷ/-�C�I!����"Q�b\����z�vB��),�t�����s�1@��R�4C�	�K�����E�M��D��#�t��B�Ɏ(��[1�P�5�������nT�B䉉:l�� j��w�dXy_�Ш��"Ov��s	�:0�D#�Aæ�zM��"O��dUQ���Q��dcnm2p"O�x+���L�T�:�H�efջ"O<��N�6@�P ���p��"O��X��>q��U�i��N*�8"O��dfK$����'=n��#"O�t�ٜ"�^�;�FՄf�h�A�"O�)�T�YHm��+��ye�@�w"O����C<M"p���	D��!�DX&U^�������0�k���5+!�d��pG,�x�b�8|��e���!���;�8�ɷɁ.E��&�@?!�U���$��o��<(��$D�u-!�]R*Eh���j�읢��O
M!��:�@��$	���pd�! H!�D�^e��B1<r`�!�e�%3!�Ϣj,�b���s��ɢ%-!��5S �aroH ь�YE�A�{!�$@BڎDQd8?�ެ�Gݪ.�!�J�Z V��oN�E����%E@�M�!�� n@s�5���Ak\)/@����"OF����"u�Jed��8%�8&"O��2��S
G�b�[cK1c��7"O���@�<@'z����'(�"OF�`OȌN&ʩ�D�_�( ���c"O�HKuMW [�� �cՠE
T�8�"O�0�#OJ�.�����֡x�xc�"O�m�D�+/��t��ƚ�g��p�P"O4�B�J��,�$ �����"OXh�h�4��(�f%�+��H�v"O��$�֏.;���f�$s� ��"O((�#*Т!¸mX�E��6۰"O����N�(�lA�'&�	�!�"O0rS-��[o��Ř�>3�I�"Ob�z G��z��҆��b�
2"O��S,����p�^��t#"OR�ڀ �*q�T8�S��I��8	�"O`���>��Q��/z�\|�"OB�XP�����3%�]i�|��U"Oƹ�"<`{�1!&F�3{ �B"O���C�� �d�:���b�̌�s"OT�)�e�6!�Z��1c9&ĺW"OFe���$���!te�t4d���"O^آ���>���̈́�U(�Q B"Ov���ָ5��d-ȌO+��ٵ"O49+E�3J�MJ;�$p"O���	b����T�^�,d�'"Oa��""��eH��F�!�`"O�@� ��G�n�{�a�4^R$܀�"O��kCAW�Q�����6�H�X"O.0��(sc�0�'](M ,��"O\��K�g>܌���۫5 �(�V"O�xZ�KĢ$wv�+�)О1Ơx�"O�\(�.قj���1�	��{`���"O�P��N*x*p�Q��<)��9"O��Y��]��ӦX�W��"O&��Bϔ)mr�-U��m���	��y�D�i�I*2@B#}30���)�y�
U6��i�m�%ۤ������yRW��y�D�)v����J	��y�/��p0u�b�"W M�͋��y�,=;*DqRI�6t@B� �yRGK�,)~��B�Փ~�<�`�"¦�y�iE����5Y�����ă�2C䉮LP���?*��QQ�%�)R�B�I0f(�B&,h��Z�-[#n{�B䉭z���:Ia�5"����L�pB�ɒ8�̌���G� c���5f%*$B��Q~l������* �F��C��+X�@2��]!�Q��ݷE��C䉬O�#�I�V)^= P噣EܸC䉘5��G,R�|��+�*����C��j���Sw�Х�DK���C��l�T�A�C4q�M(���6U�C�#5� �愬$�89@�EB!#��C�	�CP�8s��3uO�����ޙA�jB�I�8B�HT�T mJ�@�X�.B�Ɍ�
ɳ�m�/S� I����|`(B��s�E
��(<+�[&e�24�PB�I־����+m�L�0�ڐX�C�	.J�Q�F��.�A��8Mr"B�I�mN(�ઐ�ne(��4K�	�B�ɫC��:���7%=άx�oQ8�TB�	�Z�΅I&LMm���9C�$V�C�)� �X�qhY�'��Y�R�jS���"O�-I�Kوu���d
�FC�Y�U"OF�����
�:Q���΃ �Y{�"O.�j�^�1
T�Ȏk��e"O�� �m��5�rȓGD [.@HS�"O�Ѳǎ�3G�N�*V��a`��b"O�L����"�F�2�����H��"O��QqCȸH�N���ŉb��@"O���c�� DϰXB��Л�"O���4%4���s���,��S�"Oz\�"�T�CJ:��L��L�F���"Olʡ��}��5ɱ��o�d`��"O��xb�Ԁ,��V��0_��ţb"O�DZ"��,�֍�����6"O��� h@�l��QS
Y��D1�"O��r�	�6��C�S2H�l�"O0@O�~���sb�o�ҡ"�"O
�%�k�4MH��U��[1"O�i�R�P�O�ʝ�婝+�IH�"O�]{PA���Q��-aR"O���GiG(g��j�fL�.���#�"Of���\�=�k� U-X���H�"O�1)DMø��K[u��`1"O�F�&h��hXe��%nN`	��|"�)�S�M� ����$8�ā'�K,/�(C�	0�j 
�
a���g�V}�BC�	&\؆�{�S�>�ʬk�J��K��B�	��$�#KT�=�j�yTȋ�B�B�ɑrf2+R�V+m����	�C��H�m�D
��J��G.�*D�C�ɲ]񘴫�`��V��`qu�C=�У=�Óo6�Q�CƐ-�6�%DR�[��,��(ʐ��c�-
��%"�Bۄ�F��ȓ�;�+T�6�x bU��^��܆ȓD�,�zA�:$��	�ᐚ5�~Q��o7F�bLIt��+��X?ӅLt�<1b�
9
X)�ع=W�,a1I�o�<� �<r�G@ܶ'`�� �Tp�<Q0蕋1_��F�	��"�o�o�<��I�85��I[G%͒y��
r�g�<�3BL�V%�$yF�b���eb�<����h�����J��F�欛�	c�<��eß9<�,Kpb��*X��B�e�<�T��\�N̺#bZue4��]��B�ɁE��=��@J)�8�S��*	ܰ�ȇ��16�d���J1�(�r�۬XK�C�	6}��Y�2�A�r����'����B��s�¥��/�Z��p�k׼49�B�I�j�BppACEK�ؽIWG�Q-�B�	S�u���� ����J=x[�C�I�\S,	�MV5^�ԫAJO�&_*C�1&/��3!���P0�D��M�5M�Ox���O������逑
_S%���4��*v!�5� 	�Ŏ��P�G#r!�dŜ��u��`��a�zع5���dS!�D�6>�*a��B��k��4!bk�!�QM2j�!��1���6d_�4c!�ů=,�P�"�ͻ )n8�҂�g�!򤛁~$���	H:`
eRp�O�����.j�]A&�.�\e*q(���!�ϡYR�Z�M�Kx>�꤇�T�!��S�hWZD���|L(H٣� �I�!�C�_|�7��F���Ŏ �!����"�^�:# �4��B�;�!�� ��a�Kػc!xɄÑ�=,�c"O����ѹ�z���V�2@�"O��h%�+MlI�@W�G��<Ҵ"O�T�!�Z�m��q�oQ�$����"O0l���N^x��S_�	��"O=�U'��'" XC��Ñ&�h���"O*�	F62�m#q�$ ��	y "O��5�\0a����Jش�&%Bf"O���$�a�� ��1s�����"OJq�S�6+>��u.�S����"OD�K��	�Ș*�㇭u�F�h�"O��BA��5��}�-R�0s�h07"O���KW9�18�!��C�e0�"O� s�FO�N)	r@�?s���*"O�p+����
�8*w�R3�L�
"O�Xp'IG����C(@���"O��u�#�b���Қ�f�=D����K60'��Y��te���:D�P�kX�D�H�f�ͭH�Bd:��2D���3��
pNF�����6� ��Ҫ>D��{h�<R��;qd�|s��Z� D�̱tc�+PT�%� �6�@�j>D��S��Cǆ��`hK�Y����9D��3��^"�u��I�-�蹑 �6D����m�}��E�E͹�ޙ��3D��*���<<��|����bV��#L7D���d* �yp��6䎐��K&h D���à�$ώѱ2��CbQ˳�2D�4���Ɇu���G�Xْ�M5D�� LK�Pp�dB��1tC.�t�3D�Ĉ7�3N~^-�I��#W�2��0D�1�K�3������<�,{��+D��:ōŖ=�~������F���e*D����kԟa�6Q℩�3@�����'D� ر��/��́�Ѥt�jy)�B%D��d/�5bX��Ui[�3	t�Ҍ.D��*C)�6P��(�)>���,D�<����paƉ�e�� u���P�8D�X���ŎD��8�F�2H��A���5D�@�0�޾[v��2/GN�����4D��S��Ѐ��� �2V]�Dʁ7D����Q9xb��u���t@j`4D��b�Ȟ^��aa����+s:Țf�1D�L��B
�ZB���hF�tܺb�%D������/�8uĕ<F�:�hw�%D� ;�I�3_g��j�����q �#D�@yGF��6P@rɘ禱"r� D��J%F(*�E1��m��U��<D�D!�G=Y��\) ɚ�*͚��s�;D�H�u*	#b����R��(�����E:D�4������TH�99�t��"8D�� ǃ�j,:�p#ˁ=�����8D���(�h����p'ER>NuJO6D�@{�ԅ����'�+��8�s�6D��w�W7L���K�++��,���/D���ď�8@���2��$5���1D�p�'�ʰs��py�)	kڝJ�l<D��cb�!<T��"S�rxn\���9D� �RmV�!�� z�f�/1�,��#l9D����߯g�,�A�-K$L�,<0$8D���-H�l��X�?�����M5D�\2�Œ�E��i�(�����0D��J�OMj���:�I� 1��E�` 1D����͉<S�Tp����E�)�e)-D�� �)#U��!5GÔ:�(�Q"O�L1�J�O���@ڐg����"O�0��2LLX��̈́tz:�a"O������a�l����hF8��"O΍�Wg��-҅q���z�ɓ�"O�Hō99�B��Ă�WP�}��"O�#�.�04 ȉp@M�1.=�!"O�8���O�`�:��l�++5r4	�"O����[-xBp$c��B�	"��w"O�0@I��=�~A&�/C�j6"O��Yv(A�H(�i����J�3D"Of��a��B���U��)x�T���"O��x�'����%�#: �'"O�0�fiI3>�^U�W؊6�T�"Oh�s��L,~�DI�D�/sؒ ��"O�Ѥ�
�6�օxS�,�b�;�"Op����@=0���#��t�:"O�mXǆRK8���C�R�8蚑"OU��b�7~���9���� a�"O�9'�T?j^�����;{J䊧"O�H�7J��%����ل)1v0+q"O�C7N��}�@���K�0�!
�"Oؘ�'i�2�٤��1+@���"O�hD) k��p�$B��ɂs"O
P��EޮňA� C�"�y��"O�9aTCH�wg��p��_�y�r��"Oj�����49�
�'��6�B��"O���0Ḷi�>9��Ǧ1�֌Je"ORir�J;P��x��I�>�-ӑ"O��AIW8PH����X�_6� �"O��C1��\�H(+d$S�E��I��"O�1�6�̝~�$Ȱ��B��Q��"O��ꦁL����$ɚ?��0)"O����C��z��PK)ߢds88"O��KSDV')(b���g����lz�'w���"��D�C�
Hvn�	�'��X
TM��.�su�B
R�! 
�'� ��s�Lt���e���&���'�"�!��8�)���-bmи+�'���$��p��z��֎D|��'m�My��EUKH��;h8X��'�f	 n��n���
���3#�1�'4JP�dIA�$�r�AN/$���0�'�~!�Va��G��<�p@ )F�q��'*9�P��ph|��qΈA��U9�'�܉PD!�	r`�"�Iв8bR���'��C���R�<��G��5ز9y�'��aW�[ 际��2\ �M3�':`q�P� ��ړFއX\	
�'�x`%J���ȃb2�I	�'���D���4� -�2�6x숍[�'c��22l̫$Lt,;q��i��
	�'�`=0��P�j����Q�a��i��'^�QY��^T�6���� ��'!^�
j�K���&�:�'�`��0ǒ�*I�k���{α��B#��`��\<ìi[B���j׌�ȓ^�$�>p*������P��c����*�w�����_�{V�p�ȓ]m,��C��P<�����Z�Ra�ȓp��+�$L,IUi��  ]b��ȓ*���[��R%S ���F�p��>x\P���>��IQa(XB��ȓ$�X�E(8�P�G �$h
)��S�? N�{cA��vľl�!�+`��j�"O���C�Ӏ-ɴ��S#��bx��'"O 5��(�,�J����V#�xʀ"O@�h����r�T5P�@#�0,m4D�p�.�r�^�QjN/��(A�N*D�8��H�� K�h�u
��r��(D�;rfҋD�t�#�
�v�>ݰ0&D���SF?<U�4�Qh*c�6E���'D�Ș�E�0WF������d�6���� D�4Q6G��W�@[G��F�AE�?D����ͫz@v���H7k��^�!�$K+�$�@�B^	G�Xr��W�!�$���p�A��ˁ�$8:�-k�!��AX���*��\*JD�ȳ�#��!���6'H 
D�;�� �ԧ�-!���;_z�0p`�@)j�]�bG��:�!�Ă%l��QbU$,˦��%�!��&
n`@����gK2MSR+�P|!���#t�G,B�r� ��,fZ!�d��]ɠ�K��s�p�� C��!W!�C�ը�K�L
P)�02cn!��J������;5�hW��wg!�݄ ���įG�%���o��MJ!��V;b錠��*҄C�����2{�!�$�5�4R�L��9~2��rM��0�!�$Y&]�b���LiG���%�׏#V!��Q���(ƅK�*��rTk�/_$!������K]�'�A��� �Z!��N�����4�ǈ}��dxe��)�!�DH.Y�~(�G	өa�f�)pȭW�!�d7?�x��(��C���V@?�!�$C��6��$�>�\ab`�mb!��8<.Viz��_m�\K��P��!�d^�F��ҧM�r���жJ�!�$ſW�Pt���X�6� '�\'|�!�ē+p�0|����V��:� ڟC!��63�}p�R�(� ;��Ɨoh!��Nm����G5E���)��FK!�D�=0e���H� Ϯ	[��~_!�dY� Yn��V���6Μ�P���|E!�I0�x����� @P�B�m!�$��E=z��M�LӘPA��g�!��L:
TR�Ȅk��M�1��|�!�	�P�|`Q��?���P�)�%�!��]gN�a���.y^�y1fӲ)�!���m�@�����Қt���ٚ�!���6$��$�R"7pV		�P*.I!��6L��M��?	��� �8}W!�Đ�K7�#��B�'���SԌ�%�!���[켈ʔ���>�z]�G�� �!���S�� ㇉\ڬ\J���0�!�	DX6��4��8g�~0��I��t�!�d��������B�6�h'/VUt!�D�D��%��U���#�C87!�F�G�6@��Iy��d�� L�:!��+"h�kCB�z
Eq&�̋BW!��gb��9L<n"M�# .w!���0U <�:��%d����]!�г!��9��W9ul���C�ټc�!򄇨��@�%J Px�so��8!���K*Z4zF!A�S%B���# �!�}�L��Z:n�@��N�Jo!�)-��s�-�a6�k��ҥe!�F�f�ZH��].W�� �o�9�!�� &}��J�/g�l-C��P$⠁�"O2��� ���X�� ?X¨��2"Ov��m�6:�a�FͳS�r"OFG��("/���4�^����&"O4)rC��30���G#K�6��`"O ,����RBċ�\�z�4ɉ5"O�DS�/�.4>�`XP._��`�b"O8U��a�&��$(r/��8��`#�"O�(rQ9?��A��>wk^ٚq"O,@E�4�����G'aZ)��"OD���L'��3�HL�a �"O�Բ�f��[r��Sd�`2��{�"O�%R�@@^x<�DH1u ��٠"O��#����xƐ�6~Q��"O�hw��}&����TS����"O"h�w"X2�m� 
r�d��"Ob1�G,�4� ��<��M��"O��@G�U;B��m���o�l�XP"OЭ�Tj��?�`C��N�l�Pj"O�(��F��)`*F'��-)"O�������� +�N��-���s�"O��qfT�4{�� ̒�&��e0�"O����(L�-CS�U�9{D�#�"O*�R�#�;/X��IN�mrY�"O��Xe�^�=v��1��+h<�!C"O2ܠ�$�/]��Z���6Zn���"O�|�GÑ �nyS4A��eet}�"Oк��8%�p ��ə�G� I�"O| �Ȃ�+�ҔٔJ#'v��"O6p���̱>�VU*�
1N�*��`"O�� �̃_�"�y�Iƻ�&M��"OT����6 ��dR�A�k���Q"O�`�*�&|�Qx���a��x u"O(�c&�J
�!����/*�R�"Ob�H��G�+�l<[$��x���U"Oܼ�s�βb�֙r�lY�ajɻ�"Or5���0 ��l���6ZY+�PT�<A��̹0$����bdiQ��L�<y� 	 -`�qG�K<���nG�<���0<����eHV�A�t��"�C�<�S%��,��+���6��҇/�S�<Q���y"�)��U�1 Ii�/g�<I���8���K4k��ީ[TJ�_�<)F=�d,�c$U9����^�<aCL�Lg��!�	�zĠ�ƭP�<������ �Fl�!~i�<���J�<�3d��'��Y�pD�Ds^����l�<7&�/,.eO �7������~�<9`��2�^�b��T g�I�U(�u�<��	'qy����]N�7i�q�<�ֆ=XOR1��%�5�L�r!� v�<���`(<@%�.\D�9�%M�u�<Y��>T�h�PV�	T� J�Xs�<	�	�#�8�N�$��Z�<	�� `���^+Sd$�Qt�	�<�v��ٌ<�ɂ���E��S�'b@q�S�M?.*��Y"e�l�-��'vH���Ռ2�� #5
C�ZJ�<��'�B]�¸P���SB	}��)	�'���k�C�������!�{6 ѹ�'���)��۴Τ!Rc˴b���8�'�B�C/f� c�-Π�[	�'����D�Z�,i2���+n����'����s/B�\>�!���(�*�H�r�)�� �@AÉ\#=>���p����d �"OR<Qs��6�te0
5L�(;s"O�QXňM�v2����T7@��bf"Op2�L������
F/T���k""O0,�2��To4T���U�{�H� �"O��q@*�?cS|��j?$�H6�#D��r�h׭J.ڠoԐ*�ƭ�p� ��^����^�Rň��z�Z��tM�
��C�	�1�*��@l@�fe�G���.B�I4wB�5F��ip�@<+�B�	�����/I�P���	^�@�
B�I�,�,�Ɗ_�k j5Y�kW�l�C�I�hf�Y@�Ȗ�F}"��:�C�	2~�܉�J�Z�&qRG��2PB�B䉗��� !�7y��(��A�B�	�T��x���S��R�VB�<� @�i�=�J�Ơ��$B�ɍJ�~L�b�˺�8 �~B�ɣW>~����4]�>dKӡ�p:�C�	p`H�a��&��K��6v�B�I\��`���
-��K�A9tr~B��3�B�k���EC��(����c�"B䉫7Ⴂ�X�@�<�r�iX�7�DC�ɤb ��qr�[4dstd����~F�B�	 b>V�SДv�K����@ZB�	�=1���>K�!��3}�B�I��-{���&E���-�(�HB�I!x{ iy�+u��D�S�Ů�:B�ɶy�8�!�K�����M!�B�Ɉ�us��N����CȲ��C�	�j�J��29Q|M�Z��C�I�[��"�@�+�h�����p�B�	?�� P2�K�踗)���RC��5�B�!�Jѥ���p7�I٬Ɇ�>�3v�H�Zw�Н?N�&���	{���	Ⴧ�F�����e��(�@1D��q�e��'���@��W��m0v�0D����2?�t�ѤP&�N5��4D��j�O�A����є\�R#�?D�$R�N4 Zy���p�BXDn?D��c1'Y3'�l�z���8~�&�"?D��CCJ�l۔X�w��X��i+�C�O,�=E����+n�3J�N�-�V.F��!�d� 1�E*D�&�(���T�!�Dʗw|y�'�Yi4�e��!w!��w�ڱ�L�	�@A��' :!��R8v����	�<��-;Q& "!���,��b+��c�&@���'�!�D�yA����^Zh����M;ў���I av�ɑ��H!�$�G�pC�	�����d)V� �$�R��ɕ��C�	4��鲪��Iqz��:�zC�?Q���穒�V��dO͓�jC�I6_�:xj�&P=��$�a�)ҔC�		&��ZsT
c��eĒ#,�8C�	+��P���ĭY�r=g�K�I�B䉶G"�����z�2H%�^2i�B䉉W�����B�hԝ�qj��a��C�ɮ^k��9���US�q!uǅ�C�I"��HV�-W�]���ĵE�|C�
=�<=�T�9rrPB�¾8lJC�ɏ.�rMh��H$%��3�怱3$@C�3�,��VH��M�l$�EJ* �4C�ɺo0��`�Q=~wZ4��΋'��B�)� ��-��^�k�]!0���"OJЋ��Z�h�r��P)�� ލ@"O�	Ǌ�G�d:b������"OJ P��w���ؒ�
�xȖ�X!"O�x#���;2I��"fD)v"O*蹢��p��L����|��S!"Ox�(&!Η�̤�th�=ٲ���"OL����5i�*�D�(o�	�0"O�K�		#�dY�� �_���B"On,���_�|��+�AG6	^�\�t"O�ͪ�F�n��DH����@��;�"O�` ���GҒ��A��1�$�Z�"O�`;d')_4$q�Z�C��(�"O�ұL��x�B(�o 7i�$�"O�,��"�:Q��A��n�f�ȇ"O�]�ŋ#I��E�V7OȌـ"Oh��A'�(�T`D!6 Z�P2"Ob�f��/[�6}���_
Ja��"O��9�a�
B�f�j'��u��T3"OR-���Y qTHr��ς�L	sR"Ol`!����~�
"I�\]>��@"OLHq ��KL�6��zL�4Â"O�1І�:I� ��"苊D1� �A"O���%�����Ef�7+,���"O��zTkۍ*"D�JvEB�
���"OtԊ�AȬI�:e�QBV�y�6,rr"OL��Տ��!��CU��68�p���"O�a��:E	\%h-�)ky�Y�"O
�������Y����?f�5 �"Ox;�C�F2h��OIR`	1"O�d��L��8X�Mbw��X:���%"O�	xu�Q�	D��2�ܺR�$��v"Oh�9 ��,CHlC���oϨ���"O�\AUk�!@�d=s�b�@� tʷ"O��{k�A �[thɵ$����E"O`���
�A���&9�n��"O"��%��
ń�(,
A��"O�xj�%\�{�����@F�|�t�"O��q�b��9�М�� ��%d��3r"O:�2rk��s2p����-R���b"O�H��k��xZ4q �o��3U� ��"OԘ�G�WH	,9�c�2��ju"Oj���@��5��� #�<m����"O�I�w�Nqy��	�n>ha��"Or\�,/�B���,D#(/f�[w"O�����X��U�Sj̇V<H��"O�p�G��z�؅�ai��Y���@"Ob8;ׂ�);^��e��#����"O�!�o��
j"� ���H��9�'"O�����2rw���B�
���@B"OB4h�e�|'��k$S�Xѐ��"O�8Za �3?�X�qa'̢c��xxD"O��� ��`�Di�&��PU2�yR"OJ2d@ߧ=��`(�_��Ux@"O�h��D� ��:T�H���=�' 1y���}�zM����B�\�'�2A�MȳI��	9�n�e�$U�'�z�X����ZIs5/� `|v���'��H���S�9�_�^M���'�@�G��D)h@.X�UW�J�'���6��+sG+H����'QB��Ï6z��A�H���P��'���ّ�s����2E��Z�'.�`!%̨uҮ����8GZmC��� |�!w��/f ��Sp͂ d ZF"OR�Ɇŗ�,��գ`Ꟁ7�f��"OX�AG��q�<���"2��DA�"O�)�C/I����aM$r��c�"ONTI&B&<��17/E�&��x&"O�d���8��UsDm^�a�"O0��@�6�f�JgJ<5���Bc"Ofd�n1'��\��	���X	*�"O��	A�Vԡ�4(d���"Oz�rT�_�'P�( �H�Kb�@r�"O*1(���t5D��gV+���"O2ȨT坸M�С8�*w���"�"O���Э;?$������y���D"O����69�"P�V} �G"O4{�U2{ΐoJQ�q�"O����<a�~��ût�U�7"O("C�Z�z� Q� Җ��у"Oʐȷ��4��`��n� �v1�"Ol�F�V�\Ch����\��F"O��u!�'S�5��ѵ3�*Ј$"O.�Pu���H�Y����/V���3"OJ��E�]����j
�v�X"O� ��/���S&ǹ&@�ʣ"O,9Ҁ�7?�`S��ҾK
��3�"OJ�x6Z5 ���閜	n���"O�$zd�@�� F��F�`�a�"O
P��I��8���X"�4g"O�t)�Ι�6�>р�F�/�R%i"O2}��5�~ث3CC�x�\�"O��s֍^+J�NI�F��9�|d�1"O.ui����ij��q���<�r�I""O2%I��$? ��X�F�b��tX�"O���Y9u2�K9���s�"OlE��/�9h�m �(O/�<@�D"O��[�
��@�tiV�z�E+V"OM14`�$/�(x�gS�&��I@4"O��"�ă,a9�)�%�9֡c""O>��	?|g��Jr��|�D#�"Oftz���T2�a�6��7�6!�"O�I1��3t$�RϱG�X@��"OR	�c&ɵ67b̡%��>�����"O�}��Ô�k����� Dyf"OD�����"*|�����!�.�"OX8��N�M�&�e��U&N���"O�PBh
m�D  Ww���"O���,�B'��hS .S=��"O����6>�EI׎�;d�f��"O^�"bЦ.��hF�ӅA���e"OH�"&��L�W��:>0����y��%E-��3�C+P�j0Ǜ�y���~��a�Հ%���	�Շ�y���Q���'��jdm�2�F��ya_h��a�Dβ�,���(��y��9n�`�$$[�w*����=�y���@�RRT�
�����@���y�o¶C���4P�F��P
H�zU"O��%�ޡ~�����V���a"O�j�F��+�T���Q
H`*R�"Opy�iF�E������_
$��`"O�Њǥ���F�)D�(g�`�[7"O�"��ԡ{��<��L'k�6��"O���ׯZ-z"�x��G���.�3"O¸�k� p� W	u�T�9#��c�<	�"
p���hؠ{�^ܒ"��]�<� �Qt �	�̤��G�6`ΐT�"OFi㣥՜v����-���"Ovi��
��b�T�8m�,1�"O�,��4S��*��8���i"O���2F��p-�BU�|�juQ"Oh�b�&�0+π(i'lĹ:R"�1"O��j��f+A��v�p�"O�Ljשا�R��iѵC��`+"O,h�1��-n\d�c��?q"Bl[�"Of���A 7?`�zb̀28��c�"O�9�d4dUMڱ =(��E"O�{'��C�$8`e
2�l�4"O�-�p���D����E:!�,�A"O2��F��U�
Ͻ9�zYIV"O~��JPK��I�"�����{�"O�Q ��QE(z��Ԯ:q~��"O�!K򤌀9�4@�rb�5.X�{�"O�eA�R&1]I�FaC�P��s1"O2��6CQ�(^*a�3�ً&2��"O,�[�)\�J�v��1�����H�"OV0��.�/!�AZ
���z�hE"Oj���+[�E���fɏ��8G"OQ9��,8�ha([$pP! "O<�+��X�6����Ԧ����d"O� �$��3��	A�@7W���f"OL�8�N�
-�l�Hu�S-	�tM�b"O`�"K�s| �s�F[�i�v��"O��8c�X6vZ�A�W��x~T��"O�D@��˶X9��@v��0Ts�ц"O�m��'��
��t�JKiΛ �#D� �e%F6�l��W�.gp��T#"D�H��*Ѥo��EB�. ��rA?D�t۴��a�ɫ��C�Ss�u<D�|���ܟj{�t�Lr��!��;D�$AS ՠa5���/��l��Pk0#:D�̊Vh�>95���E	��[����A8D�@�s��=�PأF��{gN�)�o7D��0UJ���)B���-CG�9D�8ڣ�ļ`�68�['R\�I���8D�\ìر=�Х9��7.6�qS��:D��'K4�Ҽ�Q��W����*OZ-��jP�_��@s!�:���v"O�I��Ο2�!��?-���"Od�����G���rweϳ=z�#"O�-��)���VY�D��w�ޡ��"O�Qs���~d%�����.�cV"OPI�#F�5"��=	 ĕ<j�i�*O���զ�2�paqA X�\���'�Q����9t4A���Q~&���'
���.U$9��q"�t֩y�Oz��䙙 ����A%�Ur#M�H5a~b]�\�B R( 0�hB흪s�5Y�a&D�4�$�ٵ>�b�K��LxA��	$D�`�7�Һ�Y� !_0Du*aO#D�t 6��(�|��I�� >�p#"�O�˓���r��1^�f-X��36C>L��"�.L{S���#ή,0bI�5Uդ(�ȓLu�L�tF��^��h�I��r�ȓq^.1����P��3�(H�ȓO�'�X�ص��/Y�h ����I\}B�D�>zA���R�K�;�����<�!�Ė�X���'A[�w�\�Õ����h����
$�_"��$��R;?�>""On�y���3VC�A���h}�5¡���﨟� �Y�pc� $�$�ؒ'�0�{�"O������?���7����i�F�O~Ez���K�k�������f?.8č��&r�y���c��1B�2w�x��#hY47Y$�=	�2��0�6���#hjy��(��I=��O��=�G �]�ŢT�{:�z�OP�<�3���	9py� eOXj1FF�G�<q��P*,�^���O;lc� x��C(<�ڴK�   ag��N�|9C���5����;�<��dD;Mp#�g�"Q��ȓ4���⬝;&5�y9Pk�3i,��=Qۓ;v�@qt�+z���(CIΘm&ȕ�OZ�<����F�[p	{��N�Y�P�P�ôV�!��	�lj,�qV�J�h1�Q��>e�!�D�X�B\a� K:\�ı��R�W�!�$�r�P���4�jY���
� �!��X�f���iX�l����.Ϭx!���6d� �t�=��( �͟^^!���42X�"F�����+��ۚS!����T/,WfС#i	M4LS�'����$GJ@ƑX�%޸*�4���Eӯ& a|"�?�D�N溜�e��STʙ����8)yax��5'�tB���$~�\s��H2'��B�	��
T
u&U?Ve,�8��F�G,���hO>��d��'~�I���ƚ ,�Rr$9D���� H�{3VM9R(�Q��6�	`�����A�!5+́X�$Q/y-��3�I�G�x"F��.��)1��i�e�l]��LB�I�~���l\7@i�u/��3�D�ƓBzN�!���?A���AP(	�x��<�>�ד"��ci��+-j5��M��CH~��ȓ3D3�aݢ��A�	(���h��0}���iu�a��?g ��#��/U�N��<����T?m�ҕ�S��K�r��3�
E��O���	ϓO��)��R�)d��d/��KJ�%���'�qOV;%JJ3�����A^4��"O�Q{�&�`���䯋%n�`4�&"O�-+ʝ*tW��A/�q�(t{t"OB�����+��H��@Cg�����|�)�;"�`�wjuf$�b�]�bM�C�I4��� q�Ϡc��ЈUC 4�O���$�G�,��G�>��xH����_��~��W�<iSiúd��Ȓ)ӼV�y��GN]�<Iԋ��$X��[�e�m�# ���'��$^	�(O��!H�צ!�Q�P�<N�T{�	��0=A��I6վ��E��b@@�P@��X���=�S�O���q���'�ȫ���&h�lx���'\�����#<l�r%݋>�<���'0,H��"I+�^�����*�Њ�/�S����G��`�ab�xl�%�˔<�y��>|z&����!}�4����>�y�I��� $��zA>d�q���yR��#<|V��3�O���E�P�N�y��-i���ʦ�%r����Z��y+�/D�L���ow��r�Ƌ�y���.0��:3�Νu�ĺBǞ�hO8�<٬�̈ ��M(B�ma�m�>8�6\0c"O�+a�V-0��� �Mΐ��9��'Pў"~2a��DЄx'�e/� K3HA���?I�'�kP��S뎱�@+H�.ݖ���'
0��M�|�Ѝ�GƵ~]p�'2��D�֐�{g ���r�'jZBu���G��b�rɂU�5D���!O�<�&`'JpgA�s/D�� �,"�)@�^'��!y՛��	z���Iųy�|P��)�/,.���f^�#l!���=x ��Ch�#@"҄Pk|!��7x�nUQ4c��1'rH���/c��Syb�|ʟ��	�,x�J\1	�<y���6rTC�I� 42-�0%�.)��C�%�RɄƓh���bv&�c#��)�h� �p���N?Q -�A�h����#q� ��B�[�<�W(�;뼥�P�ۡT�  �]�'ʛv��p�O��p3֥�f!�=C��(x$I��'����G&���4��+���*Ot��4ESd�d����}�'jQA���P�Гn����'��m���;(���#���<ȋ򤀒�0<�-��In�<AW�~�^��i�A�<�� ��zP�5c�!�BQ�P�KC}bP�$�V���'��Nƶ4����<��`peE0s�~��ȓ����CIܒL��S���4T���)O��Fz��i� T������V��n���̒8I!�d�1���"P��0[�,��U1O�������s�E�AP�{��T�qO���(��y��.0PC��kqF�����o�����"��4a�V�xa���X�US3'�Mk�'A:`;D��p��ŀĖ�TF�mk��~��^�V�ZIP7��(d����H�ybeJQҕ�l���	kv)�(��O��~��$�@��w�fG.y"VǇT�<��O�$�&F�!��
׺\����>�������Gi��bf�aZ��с�S��~��I1V�1O���Ih��������#!0|qtQ��&��㉛jr�$����Zd�2J��O�D�ʸ��O�R�X��6_Ϊ�Y��.�h=Q�'Ma2�W�UӰh(�L�0�J� G�A5�p>	L<�5BK&V�����ٖ�TmŚk�<قeP�A��,��mX�D� 3+�i�'�ўʧ��:5b�e���Z{
1Γ��?�a�Ӊ}��lzG��`מY`"����hO?����1���X)t>$`)b��-x�����2}rj�J� Dz�b��~~��`�S1,�B≞X�(���	���x���u���m�㞸���*i�i���L�U���"��<	r��b��IfE�J���)m�H�er����z�#Ƃ�8p��`��˴UG���"O�IA5b����;q �(��x3�Ixx��X�J�-.�d�C��=F6��Um(D�l�'�Z�5�Fi���/E�(�X�(D��a���$�r�K�y#�A#o;D��p§�/ :60
�/�6
z��c&D�`�v�kdfaNQ+~H���"1D� � ��'���W N7�H��F<D�Hj��W$`����˘
^�L�:«:D�x�%L�u	�C (�HR�/-D�$B�逫?h��T��->t�{À,D�x��B~�.��7�ѓ�(,�V�(D�l8��,����Ρ^�d����9D������7mZ!�AJ�Zlh�J+D���I1D�8D9���?`���%6D�d����&%����ů�	���P�H6D��c��Y:�����-p��#��2D�`�A$��zT��A��"o,�,9��0D�x3�O�4:4�I�A@C����+4D�x��jZF�I������!�?D���a˖�l3JE�3��V�<	�tb=D���5@�@��A.T�K5F!`Ƥ;D��#�I�? �BDK�ȯ)/EH�h'D�� �-{�2x���I�[dD�Z'"O.t��Mϖ ��SFC�Cn�<��*Of�pG$� //͸p)�-����':�4!#�6f<Z��D�'J���'�A���f�nX�����y�	�'��-�
��Tt�)���(O�Ȱ�	�'nX���  ��C`IػoՌ���'�z	�f��_��t��H��V���'��YҨtl���ǀ[d��Q
�'��Pɡ�]�j>$�
T/�#I�r��	�'�B�K��`Et���rP2
�'��9��Nǻ)cdz���	9�	@
�'�T�0�c߼C�@��r��	����'r��aw��;=��<�Q�/ԸH�
�'ﲨ@RK��Dez�:��A�~h,j
�'��yя̀lp�Bp�S#q�v�	�'�L�BlшoȞp)��=����' H|R�'���c�b�%B�\�����
(O���O^s�D�	S��,~�d�x�X�X&�I<��!���!�D́�I��"#�V����r\!��ˬbTpP@F\9��H����> �!�dɔ?��� W �>>�R�X��2G!�d��pS<A�Ī�s��� ��݊:>!�NI���d�υC���P%�Ū6�!�$��&,�7aX}h����)9�!�dxf���2�;�F��5�šA�!�d��3u2������pn���`�!��S�H�|t�C�W>��u�E2�!��vie�s��+��J�F7N!�dS�OEXy�$�>���1)�%w!��ڨ@P��̋$q�����IU� �!�D�I�!�F��R��N(Nl$��')V���K6�]�3�v��`�'<9��C�*0�Հ!Ϳl��q�	�'�"���%��#"�B�j�dh&i��'�*��/�V(�!pOHf�BhQ�'6Z���>&jP��+f���3�'~t	*R@W�+&``�V�[����'/~ ;��BR��kSᆣP���	�'�LP����RLD(H�v�	�'������'U�EQ��W6X�
�'Jޔ����=�� ��"I�A2��
�':�xQ���n��#<0 ��r�'��4�q�N>w��7�EyH*�x�'�j�ٖC�3il�����yM
H��'��Y1ć�t~�,�Q��s�\0��'J�1��mC�QR+<��a�'6Rx�t �
L�E�PeL�%��
�'JQZ��ĶdST̠vPV���
�'���H5�Ën�lA�7N�A
�' z<����,"�i���)�Z
�'
nY�MǠ8�4�F�� B�d�
�'͆��.��t��F�C�lCԼ�	�'���7M�<H��I�]�[<�+�'��њElM�N�J�(Å�2^�t5��'.��Ul�7���z�O�H�
 ��6�܅���5m��ibk&�θ��H�� 7�J�2���;�Y���l�ȓN4����#n�Es�*�Q��ȓ�v9�����s���"@k��l�8���p)FGU�d�hA���j���5J& �@�&i�0!I�E�ĺ�ȓ����Y/a�h��,O�����F6���*��2 �3D��)����S�? (8`J�
0�1�m��
�HV"O�0�#"�<��8aB�$h(�\b6"O\�� O�j���:�Z�L@�;�"O�hK7��CkN��F�n�`k��xrkH�W����I��1���Ǘ	���ܿ2+D���L
S���&��=��f앤o��-��kB'�B�	�]L�Q�����F`�B��-�">��+I�2�I��q�����C�J��!@�*i&�ĺ"O��b��K�l�heo҂ Рx`:O�}�䈗�S�*=HH�"~�e" @���a��Ґt�0�)w�Rf�<� �D�7��/�(!^laFǂ]~���6\Z���,E8�#��KV�T슳0�@<`Sc/�O��g�2~o�m9�L�
?^d
f��-@N���Px�jT5�!#���k�
��&���O^��"gip�#��'pD��a�02��U�7��	-P�	�ȓXĉ���`��3�,B<'N͓)I|iYfM3 �&ҧ���5���-XD�q���n�ZkT"O��C�C�q�й�%�A�|�����#���v� r�'?�i��~�~m	�Q�P���I�p�tx��_[T(���T�:���˗?��݅�{���f�6fav {0	�4D~��62ڲ5��\}&(x�����l"�틡�X���ʈ|\�|ە"O
�:�	D�<���kw�		�"�S�'@Pbbh�O"f�E��/�� hE�a�'��"H:�yb!ѽN!�`sNW;��q�C����TB 4�r����O�1D��O13���3�P��c��P�.��""O�H��X�us���r* Q���A�u���� A���9�BPeX�Dp�R�n����_7�h�'\O81ӗ����L��qa�J� !�deĔY����7�Fa���C.���ʇ�_�`4'��|��V;0� ��d��z���r���^�z���Z�lќ;y~�;���~N��>�C��9�N�@����ul{�ě6?/  �WjX|�3��-6����G.w|�m�fg����ZC/�v��J��ؗktָr��=�'W/��i߷Z��vG<}V���U đޢ)�%�^�a&�~B �<%-D ˖�Kw�ti����(J�V�{��2hS�8)Gi�$K(f��dmż%-ZӖ��v�nA��b��P�+KrP!�iP�[G����cKYx�T9��к_N���!�S�/#�"����&٤�(�ÜjZ�Y�oR�@��`R�[��>ع.O�>Bt�
^Ĕh��N�!	�Ԩ�J$����#���ʅ#C��̀���C��b>�cŎ��E U�!i�RM��R��:���%b"R	���ɟ��3�	,1��0keO���Q�%�.���Bc�0Q��D�1`Y�_����9��"Z�N��hp��愛�,=�d�p 3<:Ȉp �kI���	"��P�']�sBe����C3�x:Ҫ�$r�uQǀU�4!iD�#��T�;tW� 5�@y��^>�y�F�$Xla��W�|" 0��I%\fy�����z.�E���0�D \��<ų�#�r�Z���ӐOƱʑ/��8?,1�[��}�Ư�8{�Lt*T�g�(�a!YJ�If�"� ��k����*��AX8a�΂O�4G��X�1�,�HG<M�1LΣR�%��l���؝E���'
��6Z%2�A��W0zY6��@k)�}j�.��H�|�祃��`0F�#�|�C��W�(Ȁ����h���CA9�!�$�4+��aCX���l��A7.^]�J9>�J�L[� A��*���Gz�{~ �FV�37B��U�ø�p=�%l�R;~	�@n��M�U�v�NuK��D8R��Y��"Z�h��|7$�/��>iV��J����dȅ��Q�� y�N�ؤp& 2�E+)}�
 I�a^�yh^ �O┨����w����㒛"�R�[�'3��2�(�k'���ٝsM44�C�(��<�FBIN}��Y'Ă�l6�"|b�=����@˽7���$(݉�N��"O��bd@�T�B��`���������.C�Z�KD8	uT��-ߊ��i�h�'�.�:�IY�S���s�c�S
T�����^�R~�(���aD9�o�1w��<)ek��&D��X&��TX�|H5i�89>B�m�~��t�5ʓ@�TepE��;< j�H�}����]I�
[:�V��F�Js�Pd"O���HT�[�:eC%[{�a�uO �
�T�腪ҷC�2\��G_\��m�jm�,��`g�"5��GގP�"\�/#�yҌ����i�ҏ�~�ԣ��_��!�0އ+���A��C:�i�����w�zp��' �����\�3�h�l�:?W���� ��t�毒�6�|�����Hu��$F
��!?"�qOJ�@��3?� p�H���t�����T)\-�V�I"hrd�(��Q3v�>A`B�L,^�nQ���	`XJ�a
�%_�����'���:��Q2 �����ǽ����!ϝ�0S��^����|Vo��8��'�j�36�C�G��U��+���%	�'V
ș2���	v�3��20l���'��X���^�䌹1k4�I?	u��'%Z��!�&@�-�������#N�M��	�4B�X��˻8�4zЎ��a�u℩W�.Ţa��-!�ɴ-�Q>˓2.��reA
���S(W�lF{���k�XF���1]
 yP��������y�i�GJ!7X'cY ���*M�y"��*K�Om4��W"���yB�C9��皮F���k)�<�y�*շy��(�G��G������Y/�y���@�!X57���&/�yr��lI"]�r�^�֜blF��yҤD	s�pY"S�8(��WOE�y�$׉�H9���%'�������yB���~�|�D�!WW��ƙ1�yRO�tV�j@�AI�L_1�y�g�9�,`*�OX8\@+�%M��y��2?�5"Q��;$�x&���yB��;�0��D]�Z��8�Gݮ�y��(T0hl� dr��#4�Xr�!򄚀-3$�sFז'�̽JS�L���$�)���W�=���� �\��y��@R�i2�K=k�t��@)V������k�����b4�h�ǩD���S���5��O�\��5�jX�J�I
Ekq
��02��Pū��$�칔�tX����l�Ty��ӳn�%?�L�C@�,L�<(�=�?���S�<�@�S'�O�ku� <i\T)�$bLf�"� �W�qOT�Q��Y� �KV�*@i�/i~Z�a�N`�v�qJ���?�`O�4��)  ,7}���OE���+W$\"fx���C����x��ݼsDQ�4Z6�(M:�I�ZF��AG�fjbeA��ʶ^-��5�t c�O��R���E��HĒ����?)�r�g�B��p�9}ݤ��$(�8�� �>Q@%-���'S^I:����NQ�	��LGh��F���B���Ti�D� OMp���Ho"���P�oG\�Oq��x��$2�8qSAU�R�L��Q$�L�����#ͣM@瓧l�6�* K>�村 ��`���(C��1����W��(i`L��������O<�B%��[��6�)8x��CˍY�t�)�OHՉ`c�^b2�R�ΘZ��>����V�x�yP�Rz�d�s�2=�rdQ�֙&��\��x�Z.z}�EK"�7IVXb!%�Q�������<���'^��(U�ۭ}}�}+�ͶN��dN\HGB�
)֠��a��Q.���6��]�F���y@F�i�G�#
ru���{lL �M4D~�8(��W%t�� �g�&}���f=&@����´��A�+�'c����g�1�"��H����`FM,p\�'Z�&���I.#�lx� ��/eL����R��	�2ZƄ��OF�rMC�  @1u�@o	ڙzc�-�$<K!�O�pk�.�#!��?�Zd3�lA�LcD�I�G��_�<�������a4�O �J�*�`�Vp�$�΅9�`��M�T��49�EK���l�D�J�4O0P
F�B����@5(�Z����]�O+���nƗ�a{�)�2a�����OL�b��O9{A~@�ӁZ���x�"O$M�eA�Щ�̹C�L������1�A����W��ڴ;e��E�n#P�Q';�!��ͦ~l�@��*~���Eky�!��:B���u��s>��A��͐D�!�D�;��]+u��+J/�-�����~�!�D�����
���
�!�G�
�!���M�`x7�J��蜉O��!����t�D��!��]�Tқp�!��Ї�x�w-� �J�(���2el!�d�P8��`�������W�!�d�)�fL�6w��"r�H�P�!��m���X�a(S�"0���!�$�60��c�+�+>ԡ��Zb�!��f�<�B��O;�u�sjQ�L�!��L=�&PJ�ĝ!6ۀ�R�ŏJ�!�� F���A85�����'��"OHE���,=�<�9�Y+YJ2�"O����X=�"�S��F/�5"O4њT�*o�,	w�_7�Ċ"O��p떬u���H��F'�����"O�Ł�_�m�B��׬I��x7"OZ]��tq����߲�� *�"O�ۖ	�;��t�����=��J""O`|�P#B;j�X�9£\)�����"O��brNP�NPH�SG�ܖ׶�"O���ܨZ�r�8r��[$�"Ov�0�O�#\�25���%��� "O��B!�1h��#�O$-~��"O��5�$e����%�9$�`�"OEZd-�/c�2��^�;�V�H�"O�X�v" �A|�Tr�&[���@"O�h�`��4���`�B͛p���q"O���Ǉ8U���� ޫ1� �g"O�L�ĉ[�5x�*��E�DM\��"O�p��eя�U��:}( G"O�Bq��P�����D�qQ�H��"O�|���W
�e96#I�]���"OJ��aK�3vBx�Í�#C�l�"O
I�f(�5��хȜ�F����"O��д�� k��0ˁ��}����v"O$Hc�$�.k��@��Vp$��A"OD��S%[)i��-����v���h&"O<Y�q�[�*Yj�NN�x���"O:(�U��@LR��P삳YWj�T"O���6�7�����K�6�h��"Ol�*7� /��zVꁆO�VQ��"O\ԡ�m�}�6 ��'
�~t��"O"��6��-g���k	�'t|\�"O5!��P��H��ʘ�|2h�0"O0�g	�--�����6
hڽ)�"O���ˌ�'���#��H���Y�"OJM� ��Ȕ_�A�v4f�x�<�P��o�2��Ek�N/�)Pӡ�t�<��e���z�:���6NUڢam�<��ګs��H��$��g/����D�W�<1�B��fyj�eΝ�+)*�����y�<����n`[p�"clJ�� IRx�<q��`����X�KvLفVj�\�<���mw��t̓w�*}�q�S]�<Q��ƆF�uI�@.g�� E�g�<6�;(���p'(G��m���GU�<Q7eV�X=�VnW* ��!a�H�W�<a�BG�A�\(��G�+	�\=YE�JN�<�T���df�U��d�&u��%K�O�<�1-ϐ�Uq�j����b�B�<�T��r�蘛d�T�x��	��IB�<	�؞|N��D�]�`�r��A�~�<�"�h@ԉs��7n߂�sҭB~�<�4�O!,��%��f�%�Y�.]�ȓw�D��ej��B��x�@nƗ'�6���d�`��s��5X܃� P�<A��aƬ )�|x� h��N�S{��ȓ3��Ћ��[���d��D	�=t��ȓ2���k�>�%B��H#5����ȓ$��4��F��nyX�� �E�U�R!�ȓ&�
݀7'�.X����)	���ȓg�f��N*I ��	&cצo�8P�ȓ"�64�2"D�L��M� ����ȓ[��-�e���9m��Is���z����S�? d�ڰ�X%&o��86%��#�h��"OZ�败$A�):�$T9;��"O��EJ�*q�D��B�o-����"Ot��5����ܵ�BU�d��ip"OneA�+V�}u�@�P�&$t0P0�"O�����7�� ���[o|4��"OZ��F)�"�b���JE	PGh��"O����k�ȹ&��HK�e���xbI������	�Ux�\kf(ՒںB�#�??����ϱi\���8$=�@Y̑�3&�8BY梈��'��y���ʈH����r-O���9����m�M!q�����OxY1"f�
[����&*�|��'�f4��-��B���!�z���'� ��iE�ȤO?ED�&
k�؈5�I�-��9�5�1D�a�Y.	?��`��br�ڢ#)?ɑ���%,�̀�'OT���\�tKqm�ZJD-��'���b��8��@���^8
��(A�.��R��A)�T(<��
K�0�ĐDl��Ѐls�mHA�'[P}9҆���e�}��/\7��ҳ%Z'v�ĭq3�MK�<��·�#�����5#��,��L�<)R����7 ��ҧ��^H"dJt���1u�N#k�Ny��"O����(6���x�9�Z�1&���!�ۮ'uV��s�'V:	�7�ZJ� DKȈ��0�M�t�ޮ$�1�P*��=0>�H2I�b��B
�'H� @�-cMD`�)W�L@��$�t�lc��t��h>8��#��i�t\��`���yb�T����&��0�$TP���y�T2BA�,�`	�&hH�3�HD��yҁ�I�젳�%ش��Ι�ybG�,uV��6�G���2��ybD]il��&L��r#'�yR��(-��Ȃ�ӻ?䬑��&�yR��d��i.���bF�F�j(�'�10���ɧ(��8��0�*d��GLMz.l��IM��캀�)]�4B� `WH8DcH|�h���'�Ђő�$���OppR�΅Y~��x�&Ж~0�ȑP���l�4���$���b�`�cS�u��QZ/�!�#aʘ%�����LK�os����x��\��'X.�hi#M�A��1�O^\����=�&k/X��h����ė,oN��?�A��n�h����)\kt�Ҩ(�O�$B+�xf��1m_!;���Kѥ�>&|j����Y����C��Q��[��<E�N	&h����MU"^��ĉ2��O�Y"�J�Z1��酜]�ޙP�=9@�cq�^z�Z�?��`�:}K����'����T�4�z��L���|%A�'Ԫ(�b��U�O1�x1y���,M6��bÙ0�D����� ��f�B*3����Y#���C�b١(�n����Ӟ#��BT��2�eZ%>B�5{��}BF{�X.���O��]Y!�I%a�%��I��� ��~*�$
�%B�.q��ߕ`��ECpo��T���ԫ^��E1&h���|�B-O�>�������lrw"�7c(0a�*��2p��L�u%q#�"3�q��a6��R�u�:|JP�ƙ��I9�a�� Č��g�s�D�ȵ+�b�,�Y�d|Ե�'�8 S5�̫1�0���y�Ol�Ae"ѕr�8 ���K�k˚!*�%$R�U9�OT�:�#,�D)F��A(r�����@(�5��Z�� R����g�l��Ab/\G�2WJ &�C�IM־�+�fF ��B�=k��U��ʿbv�!�'�ԩi�ئe�
�,I��82r*UAx�$&`�"��$RZ�Ȃ�.f�����݋���k?D����4~*��1��>�@��<�䘄=�|zV*\/�ȟ�,a@��/+��e) �17ax��"O����Ky\\��&f��br�-Cʉ
��	�ׅ�h`�m)�35��3ʓ{�Z,C���b|�d� �HS���I%/��r5��d�����H����)�%q��}�d.��4����	8�OF�3���na���$I6�r��	,�J�� �o u��k˴'L2��O?�i�T�C:,��xu�T'�`z	�''$�����$�"��E�'�DE�u����aJ��B,C�ZTRb�T%\&?�� 0x��%w�X6M��a84�$"OR��4�
,L ��FM/�@�Ak��Nb���t 	m�0l8�"L����)$�V�bei���p��X/������D~x����I��%sij�F�Q���A���Q�'�B���ğ�r���ۀ ��E�N����Ԯ:�Z��w$ߌ����!A%4*C�X�D�6eJb�*�"O�u��M�,�qe�<�d���'���R���R��S��?�B�>9�|8�4�J�6�S���}�<�DD� ]@\��R�5d��<{�z?	�
�q��9���9LOdа੓u^��❲ ���9��' T��#Ɲ<5�bJ�ze�!����<b y�g-;D��Ȱ$�tLL�3���cM}+Ъ/�>(6$�!=�'`*!�SN�V���7�D#0�ެ����Z� =o�  ��a̲O`@}�"O�y�g�Ѡ}j���.RX���"O���� 	�X ����z'��I�"O.E�P��>���a�j�d��"O@�ECօV�"$�B����"O�0c�N�"*KԱ��!�h�x��"O*�c���`�y)��F�"Oh�h��� �r�a�!X&/?j���"O�M����!9����*�5H�jlQ�"O y r�SR¨��	� d�x�"O�����,� x�Q�� 
TiS"O,����&}
H�[3b�:d�	C�"O���Q��q� 1��/�+��I�!"O�<���b�h�H5h���y��"O�1���P�B̼���(�w�����"O���`k�s}
E��:i���	4"O��C��#7(ЙR`�.�g�� >6���#��Y�,��^<N��私0Vz�3�!D��A�ʧN��l�w�&8��SՆ&�h�D�L��>9�C��v9�ɘ5"R4h˦��C��T�4ڐ*�qC��O����嚪w/�*7"��*U�۩,]qOZ����Y����=�ָ1���K�T��n �	I�|�Rn�1\Q?aà�Q;�	�b�B8 }^$YI@6�q����px�H �
���[6�Bm�8�	ăd��  �>���1#�D�F���=��K7p��'"���X"��,����&3�	�%Xa�4FB�~�	U�c��iw��
��*�h�-�ZYi6AN�s`�鹰��'�"���5}���NK)q ](f(q��-H��ۡ¸'��a�� u_N��:-N�S5����
�Ӗ%����Ǉ'.��JQ&O'ΐ\9銨���I���O(��#��q��땍Q��C�?8:�1OZ���I�5"&����d����8b Ğ3��%# w�$��q��!V�A3ؿR0a}� �u(N��P�M���M� ��6]�0W��		����'b0]9�@
v"V���ˍ���e�pF�>I�$�C&���,9ZLE���h��0����Tݺ�I:O�(ʕ�,k�X�dJX"(��0�(��_�d��fK>@��=��
�1h��0�Oq��I�J�-K�����7�@�3���[�J*�)����y��<ϲ}�T��A��T�"�FoN>电h̂�i>L�8�>a������6^�����)�+��Q�j\#%��H�勝�{�V�IW�5�D[o�'$���r��`s��ϐ@���+��Z�HJ�|1��O�}���	w'�%0�� [����ؼ$��hhw� *���	�>6û�扬O�Hp��4�'F�fQ�i��f1=,]*i&lOؤ ��äI� ���ZN�@kQeځG�8���|�	�'Q�X�#���Y���>Y�v�;�2K^�}E�@E���c�H��`ۭ+���H�B��y��P�2��P&Z��E,�;�y�-_�i����s�,H��X��S��y��D1��Uk��{*0	u�D�y�/4�q���E�F0�����y�z���"+�qF�����;�yrf��O��Z!RanU�7/H��y�(7|��1rS��b�-���&�y��`E��'Ev�jq�'��?P~B�oP�`a�-M�a�M$C�)� (4����( ����u^�S"O���`�iLHQ�Eg����"ON�%�
ڒ�{SGO-b�Ց6"OΙ)P�8�Z䉔6h�����"OV�WjZ?'��!�2� "�ŏ��y�ŕ�\'��9�MЇ +��:"��#�yb��:ݠH����<���b]��y���4o�)2��<r5ƥc�J�$�yr�N%cqfi��H�=j���������y��<2Q4I;��8c�y�&ҹ�y�Ґ?jtB���;3���1��ؕ�y����7�#5��)Y� �ےɂ�y��F=E�0	U�8i5/Ӝ�y��Ֆ@���"�FѪLM�A#cC	�y���	!@�ąC��m���ߋ�yBE�'H���T!Y#��!R%j
��y"�� }x��{1)ǎV��b(�yR�A�7�W��Lia���yb�}Z�T@V���Y��(�&��yB�Q o��Ћ2B��J�J�2*�y�&�!b"�k�bńtk��#�W��y�c�O0���O\�a��-��f,�yBO��rJ8�q��"4�Q��,�y2c��K���PC,%k�M�5e���y��PV�ajRa�
d�ꥠ��yRj)R���6�l�=��	�"�OTq[�JV$�ڙRsmף@4$� �lU7U��q����-!�$ ���oPplR5[�laA�e]�|��Cs�S�O�D�Z5�ە;��X�O��gP���U2�Y�3��n���)O?��7+���m��ʙ	A�!3�E~�`�a��'���䧘O��E��T8�r�X�L-�)��b�!+��#l�ӟ���ق�~ҥ���0|b�N	�"tx��֬|)��AC������
"�dm���S�N��FK&!z^�cdCA�
&*A��!���@NP���:v%���x\<���MM�O�p��)��̅ᓨk��C�a�8��E�g��"�6Od̈�*ޱAQ���|��|�e鱄׼%��}2�#��?�7nJ�OQ?��r�F�4�� ⃃�(��͊`�E�.6h⟼�ᓌd�DacO�/(�29`�����c���3K1���f�-�{�I��ֽ�숞`�'&�s�E��=�4�D�t���`����M�,gB�k�e�:���W�m�B`1�{���ÄwϬe�L�$8%�+e��
>�����5,����=E�$2���.X�q��j���HO���ᓍ� Ц��"=�L�	&iEOmd� ���)���'qR�AR��3s�a��$�.;��'g�"=�~zAJ��|�湒�!HHz�G&�|؟`��)'��Rp!Y� ��Q�ⅆAs(��>q�����!;,/5HW�I�]��lУ��?��bt�OQ?����/jB9t��b����o��<�B��>�'i��0VJ�%�8=�CΈ?r��=��}򯜿a�����O,r2aX$e�́��xx�cy��'� 9�/�dd?��Y
������Y�)��'�P�p�����.����O|0�	E-G�
=a�����|�At�T%7�(sVd���?YPD�J��3"����?��N}ЕH�i7ؘ+rk	%'�̅�S"O�Pf
��Q����'�1I�h{t"Od�x�S6:P*�CP
ю
<��`$"O�*�� %3�%jӨ�~W��W"O��3����v����G؞BH��v"OP#攥?�洘#Aة?�Z�"O*i22Ń�mL�8�Q@ZC,�"Or4��'�?Κe`��Y��L0P"OP\�V��s��H��c
	Ӏ�jE"O����.V�p�!Z1Pż|��"O<�*E+J >w�u���͏n�v���"Oܰar��,^E����2��UAf"Or�w��23�؂��0p���4"O� ����B�Z����ϑ ��:"O&� P)��{����W�%�Z�"Ob�C"�³!������:}(�I�"O���[*j�q1`��Iv
v"O�ɶ-��Ɲ1��&�H�ѧ"OVA!��(����dm �;���a"O~0藫I��8,)W#X9Z����"O�t�w@�7OW�	#)��S����a"OzD�q͙�E���L+,j�9�"O��(g��� �a�U(%\�4[d"O ���LK�p>Ri�ň<#gt���"O�ڴդx��h�G�4>���"O�M�0��.>�����i:��!"O��Ab�1zy�`C�4PS�{F"O�m�٠roh�q1n�|;2л�"O(!�c��2sTdPP�,0(h�"OX�p �U- �~|�cI�@�u��"OX����^?{����H�^��"O��E��	|�
D%["~d�l��"Obar�$d�΀9ai6;d�a�s"OVEQ���
)���J�>[���"Of�C��C��~�B'������7"O�Ph�͋�1├J�O�]�޼˴"O�lp��Y�e���-C'A� �2�"O�dAw��B��gߠ~�0���"OH�S���L��}�$��uܐ-!��Gz�\0���GF�i�&_E!��=���F�# 2�H
V��y_!��6TL�:�"�u���"��m�!�D�?R�6ᣣ�!'�DbA*�.0�!�$�VHB�SF w�LtC��X�a�!�)n��L`T�$	��l����U_!���#
�h�I���+TM!�U�;Y�m�u��{���I���{8!��[)vS����^}C�[/7!�d�\���H�Nm$1'`I�mz!��օ �lI���<�� ���:mf!��8/�"�)@���#��r�";Y!�W����΋:�aѢ�Č7^!�$L8_JEQ�� �څ�����!�]}�D8Ï�	~����,��!�)$z�����
}�a�1���D�!��]<u�`[�K[���� CΑz�!�D��S��=�צ˶~�J�Z��<V�!��T��bG�p&9�FNޡ69!�d�S����T�D�F�d��<,!�@�\�T�࣎ �Z�C^�!��QDXQ�C�������J�`!��ꂠZ��R��ki�!��,(�V�D%�rE��Q�<�!�d�Aҁ�J9.����% �a!�DX�EM��3��r��!���_`!�ď3t< �91�JDtp�.���Py�lީ'Z���2$� L���'Ĵ�y�#�r�젡e±j�����Έ�y�Kd6��+s�C����8���>�yB�^�9���ku"P�fG�a�S/�y�DKAލ�ŀ�e\}#�
!�y򉛥L܄<(�(����i�@��;�y"��CqҔ
e��y�0�/�y�

�R�ka�0sT�X��!�y*�>_2����Ҿ4	�?�y�ߟ#V�3p�"��l����y���b�`��X8{X(Juf��y
� TM�Ca�XH�AMG�U��@:�"O�d��,{���];�`X�"ON@y�
���Ӵ�S,1ц�+&"O$@�P��@h��˒���Y�B"O(!���ĵz���8'��p�ܐ��"O�ɃT�V*�fK݅��ِU"O�Ď\1jh��%��~�*��s"Oje))X�1�r��VH��{VDQ�"O(0�)&���r��/Z�H��"OFyf�p/.��Ÿ[n�r"O.�+�aG�2^st���P[��b"O���"I2c��F�B�vE�"O��I�ɳL���!"Ƀ-ZqH�*t"O�ykB敾3�Z�ʕ���z��Y "O��r��4u��q��V�\t���"O��(3A�+kܼiL[|���"OdE�T.R�8��)A>5�A"O����`�0S1��:$Q����"O���i�.'R��d�΃fI����"O��S
1[�L\V�GJ&
IC�"O�e;phԆyx	y@͉�-j�"O``���J�cJ�-J�˚$Z�PH� "OH�Ѐʏ!EE3�6m4�h!"O,��V]�i��M�EΈ�_ҹ2w"OZ\�ƍ�7ֱQ#Unn�9#"O��@���gA�x�V��'YW,-;f"O0I�V���cPt���F-�\[�"O�	aT�ׂP���P��߯;2�i� "O�i�'���C��Ȳ�S:w#�aC"O쩀�"�Z?�P�4�4�QjP"O0��po��>�։�3&I/>��"O"53"�A>gi��_�|���"OZ��Q�U+}��rw��Y@���P"O��JBB�"��!���;RJ� "O�P�fe�+}�]���Z7	>��C�"O��jq�9w�"D(��ڰ	
J�$"O求a� {z����<ZZډR"O��{�HKJuA$��TIP-�F�<9`�$j��*��)`�
�q���<��Հ�t�X��F�
'�xyb(�w�<���ٙZ�� xRB]�$
��M�J�<1gͅ�)B�4آ�W%;e��B"@{�<QeF�������$o�q�-��<1Pb�;j�!U@-�<bl�U�<ytAN�a�T �i�K�<l�0��I�<�7�t�);�đ(�����C�<�Q*0v˾�PF�CS�FY�w�\B�<a��N.k�hА���\N�� ��T�<����#54�5D�:B�BN�<!����G��a3�
]�B ��!L�<�v+�9KȮ�+�e�+3�H)��C�<Yt	 �|��՛��@ H"<�c��|�<�׎9��}���xi��!EAQ�<��l�s �D�w��E��*Ef�<ه��]��r�Y�[+|�shJ�<�Aݠ}�����Y
7c<1˴��A�<�w��NR��C�~=��^V�<i�KH�8��$ʃ�6�`�12�z�<  U�`Ǻ-�A���a�5{�E�s�<)��'���3d]1&��`2��Ax�<A���h�f�ڤ,.y>�x�4B�h�<A�( fU+%o��>?"][�N�k�<��GS�>4����W���zpQ|�<�C�#<9h����al>��Fm�<� $زC��n�Hu��˫n���"OL�bW��4_`*uـD9wjB@"Ot��,�B�D��Ǡ�|��d�"O��ScႏwhJ�&�1AxtIR"O��Q�\9��8��$��fYzEؖ"O�p�f.U���A� w��#"O���A��7d�����U�U�4�
F"Ox8*ք��xa�ڠ�Ո}�����"O��01��$B��D��F��%h"���"O��B��D:J�^�����;f\���"O6e0��E�Mը�M­�""O���Bf�tn�|�D(N_� ���"OJ���[�I����A�-<����a"O�Qٰ���O�&�U�B>cZsQ"O�lPc��O���j��^�c�iP�"O$�	�D�K�P�#��(�Ƭ�"O���S��y���SbMO
s��� ""O�]���DF\[�k�*+��1�"O�Cd�N�=x� �/;�h�3@"Oƕ�a5d���^�*DT�g"O���H���-W�����S"O,���G-vQb� 1�y֢<�q"O�Uv�Vb�S��=4����B"OJ)D��(wVt����.1��<(%"O��͍�"��p㶏�w��u!"O���Rk�;,̀�4��),�j%��"O�U�P��KqZ=ʃK�$~�~���"Oҝ�K�4Xh�6��
8/��{"O�I �)T/ ��Ё�b?�|��"O8:�X�i�|���
$By�"O������u�2H��S�"Ox�'�I/8},01��	Nx{p"O���%f��#�b���B��Wv���6"Of`�7j%S����b�V=Z=x#"OP�	cbȭ��D�E�%d5�p�0"O`��A,ѸO\��wc�,
2t���"Ov\����.z��p�![�w9Rȡ%"O��C%.ܠF�l�afAL 9XӦ"O�U�U&\9] Ɛ�杕5A�"O8���Gk6���<P���w�Jl�<Q#G�����=�I��`�<�Ѐ�J�`�ͅW� Y�a�b�<��Ev���jJz�2��\�<��W�]T��@(�S�=b��U�<�I�Q�$ĹrÅ�STj��NN�<�@�3z�$�ih�t�cFA�<)��H	%���G3Ӟ��ЉM~�<a��>�R�QdE��Όx٦�I|�<�D��#i���B X��,my�l�L�<�5!?W+��C���9`���WE�<�D (�~X�&M�G)�}�&FG�<	#�ھ*w|� B|����b��y�/��4����.�dNӎ�y�4VO��x��,:$� Y��]��yBfN f �Җ����D17�ϗ�y"��6> P  ��   E  7  �  �  �+  7  �B  cM  �V  p`  �j  vw  Q  ��  �  k�  ��  �  6�  z�  ��  �  D�  ��  ��  B�  ��  ��  �  ��  ��  ��  @ �	 � � ;  s' �- �3 �8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r��EQ�( �gVlɦ�M,H"�O��@Pg�9^��@9dr<8�q�"O�Q3c茟u4P�뒤���%��"O��$f�2����� �IY8�(��"�;�g�6��I؀)?D���嘈p�l����J)�4rŭ|���=E��4a^dX�(�7#!���O�iV��p���%����'HN�+���?�|��v��6��lp��~��˙}ּݙ7�I�<.��2���?�`;\O��'�LG$�4[����G '\�Lы�������I~���4��;���5M]��A��D�>���O��u�T�Ѓuk�a�V�ѸC�00�L<�N��E�����̲d��b9���3hY��~r�)ڧI��q�ȗR��z�	Usv�,�b$�j�����d�7JC:�H��B�{�L�I�&J8u!��L$���W�۠T������,!��/��H%,����P��/32d�xR�)ʓF<�<
���J �*��Z�(�5�ȓ,o�x#&�En�҃���h���
A�t 9j��b�F+� ���?��nma��[ a\�0d�N}��X���O��8�AAd�",⑊��~h)�'��	�2�"�J�l2R�z$��}�F$u��'��� P3Ġ��g�D '4��'�@��.��e�5�V� 5�h���)�S��e�l�$� 0�!f1 �b��'�y
� R�Sa-`liV���{a�P���Z�'~�>�I7Bf��S�I
�#{ -�6%�C䉇O`�7��)��(1���~��C�	� Ǿ�ƭX8����ƌuJ.B��>0�հ0�S�{�t��J]�HϰC䉍q3���`	]-��A"�֓B��C�	 �&9�u��UJ�#�4A(C�	�Hl0�n@
R���v�7��B�I.f��U�P����@{0F��,T�#>э�~�F�1i/d���=��ѡF �p8��$� 1��U �T9G��(فB+D�hP�I����rgR3��|*4+D��`e�h�Ŋd'�FS`��Q)�a���OW�`���(��d�$�`����yr&�8��Uh��G�Z���bB��y��U6BT~-��Ѣ`�d@	���*��x"L:yTn�����/5�p!4�P�A�LB�	�faNe"�B�[�<�+�.�$���>�/O��#U�7d���4j��*�2�"O��P�E�碙�5*�6:��#p�|R���F���J�N�t�ل�ơ!�6���;�y҃ύe�8�� $�#������2�?i�)�e��|)�@K<6��XaK<$�,�(
�'xr���N"l�U�/��f��0;I>!	�[�Y[bB�0��e\����!D��9D��%`���U.��\4�@�3D�L ��f��Q-�}H�ՂC�l�3�O �>�k��)C���=�tyZ��V��<�>���/K`8
��Y<m���ऩ�T�<�`�掭	�˜�I$1��EP�<�s+	�el&�(��N�d���`�O�V�<��C�x(0J��
��- �G�S�<��1 d,�H�J�Q���APS��(Odͦ�����gNy��xc I������"O(�9�k�:et���BHJ�Z�8�c�2�]%�"}*�w�$� � �>	����栤0C�\(<��Q,����FJ�90�哑A��O����'���D�ɶM=�}9�n��R��0X"^�%XJ���-�$�t�j�j���1m/Xm���E��j��G{���/@Dg�At�̲�6	˥H���O	mZ[�O����`ΰO������Y�80QK��"R�p�z��DF��(傐ef���	ΛFV�GP�����3tR��#�M��O����X�rܠ][���-_x� Y%�u0�ɤO��'�Ѐ� �'qW�0��n�:r�x�`(-6�$��Iw�=D�y���+3�DyT׏ ȀG~2�����H!!�fpc�@P!M�㞼E{J?Ij& Ӿf<�z! Z��J$�H]��yB�Dr��i��ҜHGvhs�Ѱ<��,1��D���s��V�,4�;���( �B䉐!�<�0d`�ZȜ�&E�{�O8�=�~�f�O��zዱ�͗/bZT"!�MЦe�1�\�&�W�2�H����yOP���	A~B)�o&Z$�&%H�X
\�����y��*Hm��Y�$�W����T���HO:�=�O��(V�>�"	��$B09�D�p�'_���i��5��qpQ�8R��4�hO?7҃c��@IM��w�N����%X!�����cé\�}֋�X}����Ez�reA�9��9P�,�]�!��\�B�x���7,B���'�a�Շ��BTӅ��Ikj�[@�x
�L�ȓI(`�FĔ�R���O	(�>Ɋ����@�3`�02ԡ��e(ô�އ�y
� ]aՍ�13�J��#倻`������F�|�u�ӵP-"����G(����b�<D��"��А�B���9�ĥz��n�^6�9�O����H{�j)�£��4���'�*�zO�|"��74@�fѴsG8\pԡ)D��@_���	���,�aU'�O�qȄ�3k�f�B����Y����ȓ5@y�7��*L� �&���PD|�J7�-��D�[�<l�C
�}`L؇�D�!��CR�y
8r�m��[�,̓h��������X��u",t(�
4F�.܇ȓk�:�BŨ�k?�����{�
4�'�ɼL�PH�?�O�9���/:���&Α'q�0!	���94�Ea/@�F գ�f��5!��)t ��Ȣ�Dg���ƃX�!�$�"K ��`�^��d�U�ĸU�!��	Ғ(	b��SKҸs�$
�,��;����Ob(�W�G':*0#G#2?HQ(d"O^����<A�t剗D�"hD6�3�^�	��'�r٨0�-F3ʠ1B���n��Ó���\�K����"1iI�<T)���JZC�X��k6����O+�ܨ�MÿR�2�G{R�.����N�u��qT"�,���#R4�ybC�O�� �+��j���ML���'p�{�پU~$�(��]��*�ó���x��'#X}���U�s͸�ǟ�3xP���'e�8�_��D@%�
s�|�!�CAX��Gy�o�2sK�A���v�@�$��y��f�r��ǣ����A����y�����FF��zʤ��C#U��y��	h=+u���%n�\�B�y"�Y�0��d�3,zr=�G7�y"�ُ¤���Յ���zu` �yB�%r	JÄ.��=#��p��y��r5ӕƍ2��ҷIϒ�yb�kHX�1S��>� P	����yB�Ef�~l�f쑗	=<53 ��y�(�\j�2d�Q�
�v}pC%��y��4���r�	-@�0�l]��yb�ä*}|Ő�C�t<����R�yBL������DH�d8 �JK<�y�!V�o�Hr��Ô"��3c�?�y2����xӀT�2��1`�9�y�ʘ46�fh^���g�HL�<���Y���m�v��D��a��ΚK�<1�Hr�D*��?gZ�­E�<AchES���5��JM�2a�H�<���R�XHz��,�3d0sQ�E�<	�c
Z-N-����	N��Y�EVC�<	��^�G��eSc�5H�����h�~�<)D��s��� ��4�����Gx�<�"�/r�QY�]�4x�@��w�<�VE�(I���uEl�N�
�a�r�<�V��#*\��p�D�j��B0/�p�<a�'��|D���hU�B��Q�<�A�X�����2<�@�ʗ�R�<i��ā@@И��B� �1��TP�<�g	�/ܕ��Yw��Y3�Tc�<�1��Q	�]����:��l�]�<�C#ޣ[�
Ix$d��*pRHy�\�<�ce��&� ����	R���JS_�<�1-�2T�p0��#�~� ��X�<�a)L�1$gr�}�B�n�<�qc�> 4`�㘎�1��f�<� �8r���s�(��3C��;��(�"O,r�hS0W|.Y�Oҽ)Cb�Hu"O��C���dh�F�@ـQ2�"O��ąC�"J�#��1�\��"On5�@k��f-�g��J��D��'�r�'.2�'���'��'���'	`��mS"�hͩ�'ń�4�a��'H��'e�'�2�'�B�'.r�'n�MH n�?f�0�S�*ƿ7��l2s�'�R�'���'t��'���'���'�h��� P8YG��cd�m���E�'���'\�'\��'�B�'uR�'��|rU뎏C���䧃z{H�b��'�B�'p��'Q2�'�b�'LR�'�ұp�%�RrM�$�C�\�X���'�r�'�'<��'�b�'���'� ����O#
�L�U�Y�!�(2�'s��'d��'L��'E��';R�'a���3&H�\�Q�$��4�p��'P��'I��'Kb�'�R�'4��'/�5S#̨fi�%����k#�'#�'��'�r�'�R�'�B�'��Ӑ�R�YU� ac�.&���c�'b�'*��'���'T��'R�'��ث�n�&��h�Q��N������'���'��'���'F��'S��'�d�J�d�s��:C�fŰ�	��f7��O��$�O��d�O��D�O��d�O��$�K*vPb��
3�� �X*�h�D�O@���O��d�O�d�Otm����	\�<��ތz�:�q��\�1�-O���<�|�'��7�F�>m�E�L�J$� 
#��1��x7���ش�����'2/�>��-U2l�r��ҩ��Uǎ�����?�A�M��Oz�;�bI?=F�@#i��Lc��xs�Eg�?�I�@�'��>q8R��8�N@�'�îj����D�݋�Mۖ��I̓��OY6=�����OWƄ�&�_�.�r�O���n��ԧ�OL�sV�i?�.^�ȭxS;@� � U+5W�}��� P�=�'�?q�*O�1��|��nH�9�
 ����<+O�O��n� x hb����(B��\L�`k@�0���ZS�_� ��IȟL�	�<��O��piݡ1��	cAO9!�8Ð������l��}��$�l�����t�fM�5f�B�v�Τ@�& sU� Gyr\��)��<a���P�����[1��0�S�Q�<���i����OV�l�d��|�o��sV�1�E��V-*t�����<9���?���n,ı�ܴ���v>=��'Q�.��	�7��ms��T1P�n5�b�"��|J*ON����֮ہ⵷f��<6(�a~�'j�F����$)��I�<i�P�kHZ+gX,U"�@�O����OH�B�����I. �j���E2���ru���ku^��֯��Op��~]��
�6�?�9}�gyBB�!�.���JxZŧG�@��X��'��'16�e��P��i� ��H�.ݰ���@X�E����?��<���?���d�+2K�6
�����́����%D��M;�'@�9@�'����`�'<�������$5dD
.9���c�V�-���X&:O����<.O?�F��.o��JW��$4)@E�'扦�M�Q�O~�En�6�OzA�.�~��l��i.� �u���'���'�E�~x�v2O��$�O~ �҂�(kT��N(Oe,8`��G��?ٰf%��|�+O|�$����c߅k.�k��v��$-��զ��3�7�Q��o��+��q��8�M
�!A!���i}��'��3OJ�����*|D�8�v��G�`]��Ds��D(:�p4��8�	�P9�hLl�ɅH!\:0�;��Y����=Y�D�	��Iԟ��)�SAyBbu�P`���j5vP��D�n�YC��:3|j�D�O�9nl��	3�MC��>)�򐄁#ذ;3�+0���$`�ؠKdq��	ʟX	�� $
���]Ky�G1/ߔ���G\�I�E���y�]�L�I����	柨��� �O�8uQ�e�'�<��i�/�(����t�J��<i����?��yw��;S�� [&Yj�g)U9.�6mH��%�N<�'���İ �ٴ�y"���T��X �K	� �v<x6���y�ψ�0��h���g�'��IƟ��ɚ�f\��@�?��Eb&�X�44.��	��������'�6mM�a���D�Oh���̀�@�O#
���F�W�&�$(�d�J}NfӺ1n�ēF�tM��̚�
������ ̓�?���M+5���2�������j�0������z��9K�"M��I�Vo,�����O����O�?�'�?9#ĝ�(5������!j\��3C�:�?Q�i@��2�'({����]�=W�x���>e�B����u�牯�Mӆ�ibF6-ҍ��6�1?13"�9o.��I
!*��:�g��E:hAzqڵ �ZH>a)O�?9 �S&KLlL�3#��x���
f�@g~�$a�,١��O�d�O��?��G䘿�|��N�,�b�zd�����$�O�6��c�)�	L:#��H�撁&���h́n� ���Q F��˓7*��4N�O�L>�,O��ţȢ9��S�F˰e�h%���'i�7�K�J����D _<���Sj_.��t��L������?�2V�P��4,l�FBp�©�g�	 HEi�H�5M�L��%L�7DCX7�9?q+�0a���)��'�� �L ��ޞp'fxS��^�����:O���O4���O���O��?������{�"I���A�Z	���������T��4+�d�'�?���i�'����d(Dl�x3CK"҄Quk!�dĦ	X��|��)�%�M�Ob) a�يa0��"��rc6-AV�|1��P��-�r�O���?���?���u�X���ެb]�,@e�%�v,���?�,O>�o�$@.a�I�4�IJ�D�˚&D��S I�HH�ⓧ����D�t}��t�Htm���S��aA�r4��o�'���R�%KET+����%�Z��-?���x�	?}kh:�4��H`�B�Gɰ����8�I̟��)��Zy�x�rxt
� d�fsD�9d� +�n�D�D�O�n�B���I��M!B�4�Ucr'��(10� ��p �~��� m���I蟴����;G��sy���/k�i+���� ��9�y�V��I՟���˟\�IП�O��L�ALK�|Ä�맩ӊ#�\�Aw�k�(���/�O6���O`�?����ӗ�F��H#�K@��E.]؛6v��$���?y��mh��m��<�p�K+*�@��S�ʁ(Z�����<�b�I7����������O��dS1D0pi�t��y ��g�NwĄ���O����OZ�g���!D�G���()A^6'21!]��읱��S�@�I��Mt�izO�d�4�	&c����4��G��)27O��ݭy�,�z0�_ �fʓ�Z+�O�p���O?N8"D�H"���["i�6*p���?	���?Y���h�0��3Y���%���x ��*ԳC����Ʀ�8�$Ο���+�M���w�$9��[�F���!�L�GF���'��7�Ц�	�4�F�4���Dy���?-���Ćb��@�U���
ߠ�³��-ec�'��X�'d8���O�Uо�I���%��L��Oƕo��B��0�	��L��u�'~\,bG/�>nu�����a8�tڐY���	¦�I>%?� ���q�ji@2�L��Ԉb�)L�t=gI�Tyb��=�6���$-�'��	;NWHAt��*]��x�k�D�T��	ԟ���d�i>�'9p6�Q�[���\�?UF�Z�C��k�r|�Do��aD��$�Φ��?qZ�d�شU,�6y�h��_
���ȣ�P�b����-��y��� ��(+4������UG����) WG[� �l���d�d��M�!	e�`��͟����x�	cy����8y�$�#�$�	=V�C�I��?]��'Fgӂݱ�7�R����%�h�D�°V�4�ꄤ�>O"�E��D&���?���|"��H��M��O<m�Q!�:"n�F+м0�$�y��W0�P���c���O�ʓ�?���?������L�q�[Q�F1C?
����?�-Ojl��J2FE�	쟈��c�J�3겘Jg�7l��%`�� ���r}�~�B�mZ����|���:`�8w�дy�8�X��ƫ=
v�*��I�bQ�r-Ӳ��D���N�T�O��rk�
�6qҷ�Z�h�pD�aO�}n�&�డː����y7�rN�	�(ڟ�I%�Mk�"�>Y2�i6��'(�>xJ��΅Y0p��Ɇ�M��i�2�b�i����(i> RB�O0P�'�rP�R8ĸM #��~T�h�''��X�����9(�kE'�(�����͂��M��aϻ�?���?����hq��.o���S�׾s낑p�gR�H!��n7�M���x����I�	{��<O� �W!�j�d�!�J�|e�y0O�P����?�WF%���<Y��?)1���w�I��ϋ�|l����?���?�����ʦ�b�`ԟ��I�<Q��ݚz�h��� �
m"pYy���b��X���*�Mcw�i(�O0)�u��.Xo��EO/�4D�u���3��˭q�m���t�S+q��I柠�آbuqS
�L�h�h!D��+��*�J��0�
3h��YJ��@��4
D�Xy��?��i��O�NC�-ͮ�(T�2A��]@��� T��˦�S�4v������&���� J� UH�D�&!F�|��Î "�$����=���1cPI�Q!�߫!��,1C�-' aTFE��M���) �lb�`��u��y�f�;M���mZ�wN"�*��6���B�!F�ޙ�v'E�P�je�B�ޥqO|H7��F�|8�ܱ T�	��Vq���t��jx�M��֛n	Fe�7�5W�6� G�ٻ(mIW�Qm�2ICG��V;�)���,6E������+Jp�Y�ve��KX��%X>-��ą�zc>IE�&"m�5���%VHx�A�o�b�&��QX�x�t�XS%�/�t����5Ml&1��i=��'�"�Oƺ�_�<���H7�p�Rl�-&�<�l�ǟ�I�]R���I؟d�IП��}
�+[5��z�!ט#���" ����C�IX˟��	ן���?��'X�ӣ.�@9˥F�!�Uk���O��y��4C�������H�S�O��.��>ɢ� ��J)a̲��EO�	?S�7��O��$y�|��'�O>���|����~-�L�ab�FR�d�-)�D>
.,c��������'�?i���?y��+a	��Fq�x���eɚyH�<Ok�'~r�~���a	���Խ u�]#���:*E4=l�>�U�I�= P�'V��'.R�'��[��t��煦�1JҬȖrl��u^�H�'dr�|��'e�NI�s�耖I�g�$H�@�?V�:t�S�����O�D�O0���O��H���?x0���M �e1`�G�m� ������d�O.�$9�D�O,�d\�#�F ��iR�}FXQ9P��0`i�1�O�$�O����O��$ƍg�����O��d�..�0"9{�ļZ�� =kT�ao�Ɵ�'� ��Ɵ��t�S'(4�O� ��y�+
[`uє�J,j�֑���i�r�'�剨g�Μ�O|�����B���ˤE�!eh���g�R0a��'���'@v����T?e9aХ�x��c���<�qJ��qӮ�_m �aҼiE2�'�b�O�����S� F���kX�G�D	���ۦq��ȟ�%��؟ '� �}��A�E��у&׭�t�x���)��M���M���?���2D_��'�`3�얳bh�KSF#f�@ �Cr���� �Is���?tk�+3�Y�Эh�J8��iކCۛ��'��'�����>-OR�����b��#6f���ĝ5O���"�n:��&ֽ'�������I�k��$!��N�w��M�F�6)UzX2�4�?I�GZ����dy��'8ɧ5��Lcn���`�hOZ�����(���ԎX��O����Ol���<�eET2q9�\Ru�
�lX6Y��ˁ�K(�!S�S�p�'��|��'AN�k��q�OC�7稘X��܊�)�|�'���'��I�k�p�0�O4d�(���g�`1�!ݑ7F5�4��$�O�ʓ�?���?�D8���o��m�GB��� M��d�Oz�D�O@ʓqN��wX?��I������@?Z�t��@��B�`�;�4�?�N>���?����'�hy��d���Єp�.	VN���4�?����N+R��y�Od��'��ӳ$�&]���v�Թ���0]wVO$���O
���$6�	]��$E 4E���;�
�3-����'@�X7~�6���O
�����ק5f���C�$��B,�*�����C�M{���?	����'q��[���bH�����w����i���(5`i�6�d�O��d�!�'��<W��A�X�|���V����I��Md斡��'�����BX��Z�% c�4(�2�HO�nZܟ���Ɵ��ĉ2���<����~��T�O�*��PO5�N����?��'��l��yb�'��'�>I�&�^֜��"�r��(�E������p#�	'���ɟ�Iyy2�7%e@AH�cS�ʫ��D�<en���4�?��J���?,O����O��$�<�dM�%o�R9Ã�� �HYQ����]�ўx��'hB�'y��˟���6-'��@�3�P�3j�:}JX��������'���'"^�l`ԡE����ѡ �~��$)M�B��"�C����O����O�ʓ�?	�7z���UA6\�%'X�e��xr���>B��aj_� ��韰�	Ky�c�O��n��©N�]4��Ua�Bl��ӌ�����	��(�'�R�'�,�R�'�'��,��̭!���B!��3!w�\o�ʟ,�'���wy��ݟ`�	�?�ؽD� ����d�R�qT���Mj�O����<iЃ�w��uǎO%Dbf4����LJ6	�GB�����Oԭ;�)�OF���O:�D�`�Ӻ��O�<m�z��gDAe��x�s�����	ϟ8¢Q�p��c�b?5(����x8��7�<��4�0�{��<��O&���O�D���S���*&��$��bB -��)�)�Ly�7�x����W��S-/I���'f�^�"L��J*V��ڴ�?	���?)tB����?�Ox3�c��3�.	��.#�1l�O�@v2�Ɠ�T�'���'�rX9 G��q�XB�b�|����Mg���$؃`I��$������xyG�|�@�0V�E^"藣]O7M�Ou���OX˓�?Y���?i-O Xa��҆m4=��`ϊ-X��
B��]	�`$���	�����byB�'b�ސM��}C�N�[!�X㫖*j7
�`D�'��I�����'L����͠?%[�9Usҡt���Q�� _���I����@y��'��A�/
�%
�X�f�P���U���V\���?y���?�*O 5JQ⓼-��%a��ݺzfD�0�� d�l)޴�?AO>�*O ����OZ�O)��ۆ�N<�4h����n���4�?������;?�&`'>q�I�?�؂I�P���~=P����D*#*7��<���?!v�E"�?*�����kLZ8Q��h�d�$ �EzR����	�����	���	�	�?��u��]9��)����Q���7@"�M#���?)q�����<�~�Aȟ/��85�ψm]���&��=�� �M���?����"v�x�O���Ң��*�q���@:�����s�n�p���O��d�<�J~Γ�?qP������3ӀU�}��h��웈V���'g��'�v!Q�#�4�X���O�<�Ã�O�"��w]�\��ك�ަ%�	��j�T9��L^��'��'_R�A#?�����xd
h[��/��7��O�yY��A�i>��cy�ڟtHa��4K�@�P�O�[��1*�Z��X�̟p�'!��'h�Y�L֍W�3;d�p��&hm���I�Y�z5#K<����?qN>�*Oҭ�H']D�)�	G�9�Ҁ�FaӫJ����<����?Q���$�B�Χ�Aq"dO�lM �V�F�=��Xnpy�''�I���	��XC��u��R �Z�L<���+A<l䰤��2�M��?���?Q.On�xP�H`�$��5֯۰IEb�FB[�9Gv�s�R�M���d�O �d�O` S"?O�˧�f�)�B�>4�Ik�E^$�:��i��'��!DgܴR������O<��J�s��5����?�Z$y����~�p�'���'��g���y��|ן�q����1��$��d��^�(`Z��iZ�	����4�?���?����i��ɰ
ËV��x��EK�~Լ9��u�T�D�O ��4O����y��� (I�
L� �k$�
�����i��@�i`�J��O���� �'�I&T�a�F\�C��I2����o9����4S,9ϓ�?A-O��?U�I &�lX!�Ȍ	�����?SJ��Voc�R��O��d��`�'3��x�b��l����,~���B�L���l�؟0�	՟�B�'y��'�?����?Q�i�>6�
���oK�j�ĉ�",I���'�= ע�>�,O��ħ<�����jJ�t�b4h�@�_�P�[d �G}2_�y��'2��'R��'��Ɋ8x��'9Y"f�BhW%y�ʸs`)�	����<y�����O(���O,�v���(����r��ei�aC�d�Ol�d�O����O$���]�26��B'��a@����
GܼYv�iX�I�t�'Y"�'�¢V�y�Χl���G!Z٢Q��C.
s�ꓔ?A���?�+O�0�V+�T���'���,پ{%�<�C���L��oh�R�Ħ<����?A�HS�0�>!�Գ}�%����}���au�Ԧ��	�ĕ'�D@Ä�~���?��'ZϪ I�&e�<�Ӡ	�TX�b�T�,�	؟��I�9n�'���?m�\�������T"3�4�5Lf�B˓<պmXԵi���'��Os��Ӻ[F��4 �!Ç18�M�ܘ�M���?�B��<����$,�S!��}`�ɕ�h�<�QT$
s�6M��%-��nZ�4�	����-����<'��,aqĞ<l�6����J|��E��y��'\�I@���?�a��o��36��'e|<Ũ��#kśV�'���'���j�¸>1.O�����,)A��>T�T�#��g���ad�w�(�Ī<El��<�Oh��'Aߥo-��R'n��p�A�ǫ�;/l7��O�`�Ia}BR�l��VyR�5v(\���؄L�O�X��$���M���o"���?���?��?9-OZ�ف�>2r��t�f�����Ǡ7�Э�'d�	ן�'e�']�$�2t��c����6: �S�g�@���'��ퟨ��ϟ8�'�j p�gd>5�E'�H�昪��_��RQ*v��>	���?�O>��?y#n�<���8l�$[�OB:�R�!��#74�i�l�ן���[y�������1�-��w �xb��l��+�ߦ���G�ן��	�g���Q��}�|P%ዛ�p|Iӫ�iw��'��S��⦪��ħ�?��'u��H)�`�xRĒ獃9B�p��ǔx2�'��i]+�yB�|ߟ:��"=�XI6#�6V��� �i��	/L��9��42��ߟ���=���VB	H�[3��"�a�)�V�'j2h��E"��|B�)��R�bI��.Ӕ_�^�s��H-Qv���IU�7��O^�d�O����{�P���"mՀcI�]��_4����0�ip�,#b�'{�'%�0��@4q�X�
�!�>_�Pa�"Enl��oZݟ��I��U�M���'��O�	�c��%j)�ŮT�E�u"t�ir�'�*e�e�<��O��D�O��GOC@���LJ:{O�e�qh���	�_���RO<����?�M>�����v������㍊1���'�lh��'R�ٟP��ɟL�'���C�],Ck�ݣd���D�^}�H�4f�c����]�	����	�N��$�ʗ�g�nٸ�5UČ��S"�\�'���'��Ol޴;&(n>�I�	,'�T���܆s�sE* �D�O,�O^�d�O��iB��O�8�U�ƃH�jI�&K�9Anԁ�F,�T}"�'���'��I�S�f	 O|�� �T�y� @T(l�� lބnP���'��'���'��E���'�p���&��e��'_d���l����py2%I�p0b���d����:�G�}u&��#�G$Ț�؂ia�Iϟ0���ޤ�IE�NJфӓ�Xh�툃V��<2 ��7��<�<?�qӄ0�OJ�O8�.���V	��X/@��!DB�5�'	Ҏ�@��|�����,���nQ�Cv���3��Mk���W�F�';�'E�d�#�4�d酤	�W�`!�� �6���S�ey�#�ɟ���fy����OP�wd�2JW:$i ��p�"A1��䦉�Iş��I"^ٛ�O:��?)�'�>���WA��0�B�$"~�!
�O��l&\��T;��'�jI�W@Wj �ae�H��Xu���k��!
���'��Iޟ4�'�Zc.y	�N��
س��Z�v�"�O:�8#0O�ʓ�?����?Y��?1jkj��(D0r�HDv�da��i"�'���'<�����O��1�fV�vp P���7x]��[O��O���O��$�Oʓ0�@�7�h�1Ǒ5����"Y9vZl�R�in�I؟��'or�'`򍚉�y�&N�Qܤ A�Q�}=~i(D	�	 5�7�O����O|���<a�A��j���ϟ֘�p8�g�-��<�#o��kF7��O�ʓ�?9���?����<����?	��B��:�Oб>�|@��!q����'��W�����������O����$�j���a1`��2c��wUХ�#c}�'���'(��'��\����9<���8'd�}�tJת_�` n�gyb�Q,SP7m�O(���O|�I�j}Zw�DyR���8(PH(�`D9]_\P�۴�?�~,4�ϓ�?����?I���n*R�t1C	��&��²�Ĉ�M#��?�����Ov�'��	(Rnfm ��9��]�Ab�s�6�rݴ'�ؠY�(�H�S�O�����S�4rg6<��ۓ �	>�7�O��D�OB��1�p}r\>��I��D�S�H�Q���q���������a����'t��)p�|"�'PB�'8F� �P��ƞ~,6��SQ>���i��d��I&����O��O,)�O�X��E���B/��l�2��u}B�[��[�O|���ON���<����!]��d2��1g��/v�nDI�␐�ē�?����?9)O�$�O�d���C�B侼�cg��7Ҽ�[�.D;#1O����O����O����F��C�M�AA{jFU��
4v�P�ݴ�?q��?N>y���?��&�5O�n�3Ȑ�S�L{���� �hU�꓾?9���?�*O�$�s�c�4�'Đ�{�&�v�Y�j�s\@ ��j�����OT�t���l�y'��A��!��������m�ßL�	�D�ɨ|Nt�Iן�z�O�*{�ֽs1dT�]{l�k�.Qmn�'���'�*ܑ������i�d���!M�b����6,ϝPh�&�' ��C*v�2�''���D�OkC\;XQ��WP|�[��9O\�����7���;�h����i��FS��r�
c��9$�[q���!�7-�OZ���Ob�)�u}bR>ŚbJT�| ����LW�-i,�#�0�M�"d�z�'����|��'���7d\�\�<��Gʇ%9�(@��,l�"�D�OB�I ^���O�˧�?a�'��	Z'�'(\�H
o�����'�	�6��DKJ~�W������Q�V�L���\P	(��͓X\�B�\�G�Dp�ׂ��w��X�1z|��dƦ(t��ȦL� /�%{��Z%�z�'Hj͔��$���� $�)x��	���h�I�CBt�M"f���o��� ��?-0���&�#l�Zv��D��)r�D"J���/� X����J�B��G"��8���%v��}@��4w0H�9a-�
L=�
�㋜1���D$Z ��Ey�Ǜ<H�Hx�ł�|D�3���?�	��iA��?��O����#��C}��G�	O�������s�ϐ��A�u)�?V�"?qU�ѡ)�p�w��|�~@����>���ZN�W�(t��┊=�|$:cI�e���0;��O���<��aI�q,"%j����Ni���F̓��=)���i��%�"�,\��g�J<�6�ig0؀b���W�\��GG4���˛'O�I�l/�೪O��d�|���B��?A�N�\�.���	����W�L�?���e��<���P8NÈ��A%�>�O����\M��H~)��;%D� B�>�����A$ȴaB&I�.�Q?��!�N	!<� �� &��	� }cA��?���h���d��d�:��g̾t���$�
2�!�$Lc�Lu)��2�����ˁ�ax�E4�"X�(�	Y`��h�I��H��!Z�H����ph��
�L�|T���	ß杌v�����e\-mB����2S��pY�m'_0=��d7r�J���L�g�	}@����G�zm����n�6l�fT�_��I��Pc6��ej'�3�����m����
�qр.U>+4��9?ْ]��S~�'�dQS�QH1�B��C�k��8��'�)rՃܲ8�]�`�$j��9�O��Ezʟ��l ��Ą�2i�Z�Q�ɇnI�<{f�c��(����?	���?�Դ��D�O��S� �h��̎L��5���0d^���i��e��[+4oZ*�'�e��� SFb�yF�R�p nq�R�[���D����k�ȈsX��3$ꙩnH�1���ZŁ�@Eo0.�d�OҒO(��5�s�<�F��.xCH<�M����uHv�$D������T0�b!���B�^ �tc����4�?*O��z���Ԧ��ȟ��T�D.E�D��*Ke��d9̊ן���(4\���	՟��	�e���: #�V��0���M��b�\=J`��]�U�l['�z8����g�;E����oC��h,m�$2�8ٔ�W:�>���N����$�_y���:���OP�"���fr�e;uoġH����Չ�<1����'L`A��& �E�&Z��s�i�)CJAZ����|E��!�'>47�Xw%�|1�.׫T
8�B���0�'�@e��'�0t�gӚ���O�˧W?�a�HV�b�^�C�8��P�D�n�z����:o�%B�"�)�d?~X4���#]�i�4]�O��S'%�"�0D.ӆg�����M H��'���������ٟ)��G�ģ���J�����XΖ��B	&��w����5�)�� �&��3OX�yC~t�s&�&g�C䉹4���`{vfhP� ����$@W�'ն���4^un�а*� �Ȥs�M{�j�$�O���^<n�m���O��d�O��4�8��A�Ћ0k�x:afŭ-[T��Ҡ�f�5qp�c���q�I=L:b>�O�1AQA �D��˰.���"��Q�$y�P�gn�#8��T�� Q�q��'o��hvm�X^��6KH(a�y��H)a��L>� ���N� S���-,��6�_�<�c�3h�Z��so�		���D�^~!�S�O����f��,Z���HK�>5�n8�.^|�R�'���'��֝�<���|��՚K�,��U%`�Dp�!�O%Z=��h��J5��8�R 9���dP�p�'Sq<qu�'
(y���s�.�;��ŝ?ua�	X����*���)z��\5fF�)S-D�� ��&�;v��6́�y�����$^E�	�0L�G�i�B�'�Ԙ��ȈE�Qfe�5\�A`E�'�r��#e]b�'��i �sC|r��b��x�u�ҮY����r蝦�p<��\�[�Z%@4v���Z(szy��I=����<���R(i����BVmI�k�!��=/g��B�	Px�$�Sm��q�!�$�¦�s���m��A�5�/R�@�rWb�|�"u��z۴�?i���	�i����S�H��C5�lks�E`�*�$�O}x��OXb��g~�
�)&z�шOS�)l���ҥ���I7-?"<�r�G�.$���`�V4,��V@�Y�d�/�R��i]6��	���Y�z� �gN)T!�$ÝU}x��Wd��Z��!� ؜9ax2l:ғ1L�,���E�U�����%��^CN9XӼix��'����*C�iZ��'�b�'�wJp�b��&K*IŃ��\i�$3�;�dS�j����|R�ձ{Td�h��N�z:M1�k�g�Ѻ�a�w3$tm�6�M���|r�ɳMt��I���laŇL�
�1O�|a�������A��0Ӕ����̣��I��;�"���F�_��#�C�:��?!�i>$� �vdM�EI�Q+e@H�{��xb��[�oN�R�\����I�t�I$�u��'wR<�0�Y�j��P$��t���#�(�bD�m��YJ��do��p��!<OH�+R@�E1Z���^2!2j�q�N�iaD�Q�eI09b*�Z�E*<OJ�Q%����vi�8		���&6o���'0v�*"]�n��ڇ̌�*������DD<�S�$@^�l"A*�-5���l�ڴ��H�����ia��'|�C�S)C2X��Y�bY�u�'�#S�A���'G�	�2uU�|2�@�g�\prh�8KD����p<I�F�x�|�4�h�a���#��=2W���㉡+{��D)���OL�a5��K�\��Qx�!�d˶s�"��0g;�h�&�+FX!��ɦQ�׌�J @��m�J��[�f(�긅S޴�?Y���)��JC2�dU�)�(�q� _�i�LE�w2L�D�O�M�	��]���Q�EX�����t��R>Ep���"�rYq#���4�m�$}��#3E��b�z ��5�0ʧmn@a�D�-;����LU ���Ot`;��'���t��T��2$���� �n�Bx[#�J$˘'���'������K��b�bB|`�Ó[ۑ��b�ɏ�6�fe��*�*�*HR`���MK���?���V�t��P����?����?��ҿ�3�{!��e&F�S�Oɉ3j=	�O��yaE |1��'����"��Y�@�x���'J�Qo�������Iզ!:'3�q��'(��r�Y%q�8 �F?�p�e�{�~0o�ܟ�AЏa�n:�<)�g-�qk�.˹_n�E���*q7h�2�'��hY�V
��Pc)V�D����O:�Dzb�F?9,O6!7�ʪ[�|1pT��*`���(���*�pBN�O|�d�Ol��j�4�'��i>X�)����_Q�y����g�j�b��N�a~n�?iJ�r%�Hlվ�ba���A�~A@ ���0?i@�Z!PE����U�h �"���ޟ4�	ş �'i�ґ@K�ArL*;4����g�"O�iE+��U`2�{0��e憘 �d�d}Y�HC� �=�MC��?a�ܤW�4����P�5��=� AJ��?��xN�� ���?i�O�������Xf���F�p5���3E��ɢ,	���&��,MhX��?+�����&O$�!�'��'ܠ��ďQ7d��� �)V,-ܢ\��'��z3��z2�(/;�m�S��A<a �i�H���1�n��2ș?It2�ʊy�!DHr0듕?y/�h@b���Ob8�@ճp�v�8%�T�h|،�@��O��dEb0����E@�}���WgT*�M�Om��-ǺE��i9(H2-S%b�L�.�'V�#e�ɐa�:y��&U*\�ƣ|�.�w��g�K����.�E�$\�n$��'�>���!��s��߾z��Yʄ�ڮbK
���=��,*�ۉ]��L�8�$I�቞�HOd�3ģ�<]���AdïI�(��E���1��ޟ�I�?������`��ޟ$�iޡ�Y�w�DL��E'{�rU�u�a�X��ٲ^$ң?���6 ��y�F�U�NhS"�O�̘'���J��O�g�	�d���N�fZz�{O�23�y�	�0��8�D��)�<i�=�L����0q�>�(�K۾h��dp�'���h��ց��� �A �Jsl9�ONTFzb\>��� ޴��ܧ&$��� |��r�X-6���yfb�O����O��D�纻��?��c� "����`��d+s����\;�|Z��A.0I%k�g[џ���|nZH�n\�}����'e
(��aG�	c���pDN�G+�(1CLQ� �\	���:��
�<�B@#`ID,h$�0��u���
�
�D�<�����'� ��*E�BI�@��0z~pej���.ړ��3�4�C��QX���K�����Oz��G���1�4��)�(D`o�؟��IN<���dy��z�J�1V��E����p�"��(�I̟���BU9M�@{��+c�ZQ��e�sn���ǡM9���Q��8 ���H�I-7>H��Z�@��	�ʊ;4Xa�gt�CG��q�6� �����O�����'�F6�\ʦ��	�i����C���'�����^%t�a�'V�H�'�4���ʄ,5�� ʥrJ�-�
On7m��a�̙�'A�
?!���3CL<c�F�o䟈`�4�v�0_���	Ο$�S |>�����Q��,`p*�L���E =/6���ڟ`�c��$7���@�c�$P���)�|1�OV���z0�`��]��*�B�^)��q���Y!D�EP�\B�O��Pk�� !�d;�	M�8i
H��v �O0�d0�'�?��%S-Z�(@����`�
VAb��	�'�5#�Oǅ����� �쀳�ő��I�e
Z9$E�$@��d��m�������O$�$�7~ 5��O����O"�4�S7��W��C"�������(e��!1f˔�C���̳m�c>�ON� �,�<+]�� !� ;��X�	I0��T�%7wRD�p��C�q��',",��d�"2��P��Yd��2��'��ɬ'���4���$&�I�-��tzEY #���f��<C>tC�Iv��$ʉ\��ō6G��lF���'��DY2z}�`�*-����E��2X�\�@S:v����O����Oty���?����?�,+��e��h��IJV����ƟG,����,'�OP�+ҫ^cD���U�W`�4PѢ5� �XT✱a��G��_X�D±�ɐH9��H�H�Ԑ�egͽQH��ě��� ش�?	+O��D!�I83(�1�)� UV�Qf\τ�I[����|���&�I醑��@�JO��ᗃ'�DV��uR�4��,QW@�o矰��':�lJ��Ŗ �h"j�������C]�X��Ɵx�'u���*�Ď|�I�-���pf��)�h�C�Y?d��񤑦&��Y�|��_�e&V��]�-ĭ�EÃ��p<Qe���P�4{���':t���F�b�U0��Y�93eS���	M�S�OB���aΦBN\�C���{�'�86�S�$,2�R �-::�����3zC�<�Tj�4����ДOl�12�',�aK�d��`�+�!���'������ڭ�/L��8`�^�r���	��;�8�r���mj�H��D]�K*��0����M�Q���ʗ!�gZ�����+�!'��I(�"�-!���+��?ZB"��O�}B��<|D���@�,>;Ҡh�J��a%@���'�]#��ЧpD��!�J�r�:��'��"=�(�* �~�Y�nź3T������2���'i��'pz\����UM��'��y�擹�Bh��ip�Xx��?Y>*�O½y����I�Ԓ�1OBLJ�BAY���ʠE"p�DD���8Z���tC�M�9�q��')����5r�e��B�\+h�.q�6Qn�ܟȩ�.�ڟ�>˓�?q�k_���	G�>� tr� ��xB����d~B�'
�4�}��Xm�@�ɤKS$$q��V(F܍�Tcӯm�B�ԟ�z�O|˓�?��'�?Q.OrA�`J�IO6p �-�;��p�P"OP�1)ѱDz��ϗ�5�A�"OdMUv\+�%
c��Ya�!��y2���\�J ����)�Һ�yr��3������N�iۗ���y���4&����� ��xB������1�y�.AD�%s��\�r誑B �	��y��τ7p�`����d�"(#�L��y�FE�K���U�	/_,�{�e�:�yN� V8 
���	N�֭�2����ybƑ�m��$�W���)@rG��y�ʌ�o�I��]�m�q�F�ɮ�yB�ٛO�$C/}F��Y��y�fÑ'�������B�K�o��y�������挚�2��Z��h�ȓJ:չ�A��ל��%�8lb���|� �p��'����ܶkP��9�)i@�\/F;�8g���^E�X��S�? *q��Ñ6@�"7Mѐ�X�b�"O�8��(w��5a,��Bya"O�m���NC�$B�؈=����"O��`�A
�fm3Ђ-[�N�*�"O�L��H/6ƶ������Q"O��cw�[Kb��"t �q���k�"O����'�Ҝ�yF�Ŏj�֑��"OfHʤO��0m��q�Z7vkC"O�L
���eh`}qU(Dz�Y8�"O��b5S6α8v���q%"OdD�!kO-w���S��|�d�'2��pC��,A�T���0z������!jV@��?!@�(�0<iD�tll����4Z���r��f}bkå7\�Є�	v�H��Sa^se�	*�
�sb��[�;|��z�8em<�	�V�h��A5��̐�@���O��Ā� ��~�	�M� hٴp�X] �����a��"�MEz2`Z�6,.F�4��2Dج�D]�y����D�X5t�(�E�O��ё�|�n�|
じ�*h�R�服�U(�L��}b�N�e��Ɍ�3
����!���5f��qw ^>a�4�s�8V�:�'��7ޭ`X��d�	�=����7��'˘��!D���0W�UY�θѭO�%ϕ�:,2�(I�b?-a�o�u�Vu�2d�?��qI�`��T�J�Sc`EoÖ����$�ў8�d!���y7��:T ��$��)�!P$�8���R!A�(X�1��$3�E&��ASg�0,�xb�0/ݫ���>����k0@8V�h= ��IW�A���/M.4���8[qSu-�O���*Ps�	���iD4&j�m�;�z����D�h��%x&��6x�T!oZ�0�Z��%E�DOd���
$��"?�ňO�Gq�=��@�<.g��hT��K��y��5ՠ;W7�� ��G���yR�_/� b�ƾ5����B����P��1|Od<3�'?��£ɫ$J�E)�bZ�[|tѩ��	|z��H��O�b���D{R�?�*�R���3Ï��,��x��憛V�:�>!��^^�O�@��GL�w���������7�I�y Z	�'.�8���A��f��1����j޽B�҈`׎��B�Ҽ�s���N�6��ӧuO����͸A��A
@��>X�m��
S ��ڱ�nӈ�A���-�V`��З��Ѓ��:�>%V.L"I0�t{���i[��'�ɔm���s�!��2��gyX)V�c�C) rR �R	��\���fm/|O0�K�w("�PAȏ"_dY:�%]/g��3�*�/U��"�M��ܑ�8���������R=�
1��E2' -at)g��;Q�9�Ʌ`�>h1ݎ}����G1eV�t���D�+<`f��O>a�I�)]��M2��-5�ݲb}�t�'I,�d�p�S��fI�~�:��f ��f�^�I�� �<Rى���:>@$�^��ų�_f≿�1��)����I�>��[u#�����׃7���O>���'��㋞���અe�NܓB�K�K�E3���r#��b�8��'f	w�G[�Hp�'B�O�E���zC�Y灅y��!���Ķn,l��3��5�Xɓ�"�ax�C]�%|�lpI���Cl^Vmp�Y-f�$�)O�x'����O�qOĠA�M�V���b��[?;=��
Wc0Oꕂ�Ni�	:�ܙ��J_�Wc�%Ba#��c������<i��'Ҏ�ʧ\��x��\�z"�[���70�ЪO,��Uq-��%A���?�s�n�
�S�~��Ӻ���B�@&�3`��g�@T�C�h򉤧?�K�k.,�*l��6�[�'n6�ڔ
Nz]�b�n�p�bK�O�#t��%i��?�zFB� ����Ѡm�`��Γ��Aٵ 	�^�z�Ғ �_���ƃi?Y�e� m�V��˂,7�j�D	�5���%m�������Oܓ���tj5���[�K�WhH���-iC
�������0!p�,|Rt�e"!xZA��+`���츧�ia�Z@��3�%�]�pR�`�1~�
|r`��"�f��+��'���<Y4�� �>8��'h�L���DjC����N��w�x�f�O�:G�D�i�2���X���'&Z��!탕):J�!�%3��H�'R>Y��˱�,�%MT"S����'}J�l�.m��hٴ#zՀ �.b����E�y_��;�O@-X�����Ě6M��|���w�\)�a j�	Ņ 	{:�b�Fѵ"�!c�H��)�0��5���Oڅ����b�K�w���( 	aJ�Q�(�$�Ɏ��uY$��U0���MS��m�P+���>z��TunH=�v�v��18�H�R��!-o�Q)�����s�F��rh_�1z�)b�զc;�:�gTm�d��&�Pl8�k^����T?�Ro��_����%̄<0�����o��2�������C?b2���5ݟ����}��N��M�U@Z#BbaKps��w�L��ʟ4	��%1?�s�O�ZQ�f�<QL0'�7~��%�դ�_�f���1�|�d^(�y'��1	1j���Fd���zq-B���7Xѐ��ՕHi^��'ɀ ��'3JT`�HbLM�%&�D/$"*9Ҁ1�@֨dF��yB�6Ǧ��c͔!�"`��-ti��"[>��bB�0Mv��ͦ?�C��Ҽ)�J(k��!P�8L���(,̙v���np ��3扐f`8@�Ҧ�N��Ð@n`x�iV
Z��JS�WB:�OZ��BC��:���7f�C���s������-p ���8n�1O8�U�:j��a��o�>�+d��6�t�G��S�.;E���l�FG19�؁9��T>]2r�C����.�UтJU��P�\��^)����L���D�,O��#���`0�5�� #��re�5� c���pa���ڨ
"	�.�b��X��92��{U�*f�����ߋ160�cC+޲S���"��)�$Β}�� �Ù�a���gS�Ka�\Z�.߿��ͣ��\^2T��݅uj��iE@�:�b��)�@�>wܴ!`%B���3c��00��x�3��,a�#"��:s9�-c�+Rs�jW�I�W�qO�à�i\:h��1�}���5�]HQfA����F�8��l��⑴i]*ȉb�ZU��AD�ަ]�H�ҭ��h�qO�(d5�y�;5 ��'�%p-�P�&�I�E���Q� 4�|BU�
�<d� j���Y�p�p�ҭ��@Xd���/�V�Nb����'�RN�)7n]�
�M6�4\0s�B%�ĉ8�l?Ebɐ��!`4��M��W�&�O4��E��@&�Q ��,i��%�Q�\'�y��ɟ
,}�Q_���s�ɋH~����
!�l6 ��Fȅu(����w���&#n�ƍY��e8��Oƌ[��%��sC�\�1���ě��)���؅ *j=�s�E� 1O����L�<h,�yb� B>�!� we�98�)O� ���rN�:R�rasS��S��	��T>5������5�Z�X���&@E�ԌI���%y�>��7�,Y'T͓�yG�,Oj��N��DL!��xY��֊(�	�8٨�҂{�uX�F�4RP�b� p�O^�G��H�-HYC�����#�t5:��I���зd(��Y�P�ҳlݼ 3&C��E���SƯI��6�+a;4��	Z�&�%|���Ug��2�Vb����c���Ɛ����!d��c�EH��Te2@��#Y���ۑ�"���#��ٕ��fل��EECdqO���� \>��#����+f���;�R�j�B�?ER�c��S�LB���*Ыd�"��Q�F�E�V���/Ԛ
-�HB$_UqO哭F2�̻Ǝaq"B��e�!}���KPG� P�%[4+VF�	z�#|�'�v@�^k�$�D���{����@�A̓;�����H��]�X�_2	�����?牢w�x,:����{�I���^�~�x�5��r(���O�:��O�x��g��oy���'6Ѻ�2�y����B��W��c�[�jc�Q�#���*�������Is3�4m�!m�l�Z��w���$@>2P�9���(_G�	
���'� 㗆�A�m�3I��)�x���}h��O��)�E^�"�T�'��?'����@"���#*Y�8��q�}��xDCs�nޡ:�'C4|j\��@J��b��Uk9�ɋX�t�X����L�"M��݄I�xvg�+Z�|�9���J�I�4��� ��EG��3A���v���2u��k���
Hh3ˋ�y� Q�	�v_���s0����0}B	M��deZ��d�@-s`���#S�!ZT��*f��6V�Z�"4Y&M�$�Z�-�d������-�<����W#	�`��Z�l`ҁ�=m2<��'��5z��Yg�g�I�F�@��h�(h�S'��#�$*�9poP˓2�AΦ���4̫J�3��D�W|���hA�%O�ei4D�A�=����xA˓(@>�]=�z%�d!�9>���5%�0`8���M�+��Ӳ�+\E[j�S��O�0w�~�R�̟s`�x��'�p2t+��^��U��ד$ј��A-�$,���F�*oN��hÑ\T�M��B��`��6�������S�ڻ��8�� ��3w(:�ʧ��V�t��'n@U�GR!k$b�x���X x<a�U'�~�Cg������W䵫$b�jMt0ˀ�щN�YuMn�آ�L�Lh�&?�xX$�M�I-��3�h�$Z?>������՚ЪcFH�u㒟eҀyZ :O�I�[�-�'&E�$��%O�4�rw�2nҐ�!iB�b�]� ESK��Hؔ)R!A,���4FE�̊e,�'24RDb�Ik�ڌFBs�(S��)�	�9��A���ۀUˢ�F5<�|��f�����K4q���c���E|�!J�C��f	{�`��X(HQ3F�ւ$��r��>�b�@����!O�I��o��,�tn�;BN�5�Ƭγz�3�)��H�#},=3�eô%άxC�Y�FR��{R��u'̽RhڜAg/ޖ[�v	���T2��)�����l�ag��1	�QII|�>9�@�KDM1��œ?Jh%q�煸)ĺ�I�4c^=���G7�N�9�0��Wwr�$�����p�G�)1��q�/ٍP���e�Y
K'z��'_<��"Hߴ���1e��+$x�1���k
�l	�H9��0E��C_,�����<�򏎗cj%�͊�2x�D
� �p=�ı.�	�vy��,S�>>v�²@��
�m�O��d(��ƬWP�!
�G#{����~�v��N~�s冿b:�	�f���T�@Ԍ�\�V"R *�C/��;V$TnMh���Z�F��`��hh�ؠQd�/�ʬ��eժN��Z�v�`���X�g�3ʠI���w �}��
�[���r�X�	5j78{a�R9tiq���2���O�����36|��VPM��BP�[E@!I�E����ŔV���W��S�U��͛��Z' �g��$����
�v����
���Y��Ks�����X���TkZ/$@Np�1O6���MO�Sz v*���e �� �I9PJ�0�<B�#L;bd�Z����C%��B���`�ҕc�@Ǭ!z�h{��'��=@�+<���1C[��Zt�O�^���²n@bp�	�B=~x	�m͠dD�Y:b`[Nb��S�nt<U����-k+�h#S������ǲ<�"�M:th��N~�=�@��qq�:f ��x��[�cG�I$N����#� �&��Oq�(� ׮`X��	΢�b��Ma�m��JW�j<�	��b3�)�O$@�5f^�Mx@�"iڸ$�(���� �剄)c�e��R�� %�Sa'ZX�iز&X�E8Ք'��Q�D�ѥV���i���(��g�'.���m_�\^�B��Cs(L�$ͅ	=�$CA�C3`28�@�W�}R\�҇@�P�.��&�1�j��/OP����+G�h���ؿA#e��ύ'��	�?F	�͏;G��\b� ���O�)$|R�[��\���%��xO�a�wW��������%?�����*��cV�m��cnRL�c��|�`�O�@[��&�̄X�8�e�Y2P}�UM\����ƍS�^�Ð�E��pc$ȂS��5qA�*PE���%-��i���Q*@;�J��xj�����Č5�\@n�fOB�В���h�g�Q2ذ�IR-n���:�D?O@��Ȗ�jp���ǉez`5ӷ5)���*�O��
�rUZf�A���P��GM�B{H�ܴNü�p�?�)�I�|�����<�pP8ve�?��{�Z�t�ڴ?��(��'@q�T��O�>7Ё��a_��A��G�����<��=Y�Q>�f�nAh��ԫzH��c�2�N<�ȓy�l8h�$����eÓ	^}�Dn����{
�}���J@G�lN��ek_�b��ȓ:5"�a��p�Y�}�BŅ�R�h�'�5 ���S�x�.��-�(<��eS,�`�P�� mA���.��2�ɋeN4���<{6D���w�`����A�E9n����ȓ9����D�\�N��V�]Y���ȓu�t���D�m��b��;��ȓ	*��q��!2�8�e*dp4��ȓc�n�kq�B�2�!�&W.��1��i
�qd���%�B�k!�dr8�ȓ� ّ���YŚl�F��]h���Z_�]I����0 ꏱ��`�ȓצ�04��#H�DԪ�+7������������1KB8C4!z®��ȓ�da���Ҙ
�<���,��\o��ȓ>z$����Q��h��n��ȓ^TH�K����5���X�J^�x�2���}��}�dM�
+��HS�9�C�I:���	w!��A�a�	�@~tB�I	a v��u#G�R��� �1P�xB�J�V���-�th��k0�LB�	P�Ѡvn3l�K��-�LB�/hr2�{�m(h.s�Ɛ�tC�i��`����!�@�A���5"O" �@�EWp�l�bOҢ>a ""O�-BB���_:Ȕr�AZ�j�yu"O@���
v�^$�@�Ĥ$�̝"�"OEYbl8'$f=��o<'�E!�"O�Ey'�ȍa-D ۄ.�|]��"O��pO�hW���w�,_�v�"O����͟?Z`�u�A�}ْ�"#"Ox=�"#�JU���`a�%>���"O�My0�)`E���Q ��n
&�8"OL��S#�`��H2���"Ox[6��m���qvI��,�܉#"O6!FA��k�l����XD�"O%��e/w�jWiЕ|`ۣ"O��1#^����YW�I�|G��"O���3�J���r#�,M�P�B"O*廃�#!�Uz2�3D/���yҋ@�7��4@���R��� �aͪ�y2J�7�0;�%ױF&!8�kP��y�o�%[�dxq���pj�:É��y2"߭;&6��N�1��RCD ��y
�  ��b�}������C��|�ȓ�� �bF�$�=�ҠF�+,V���f��(�䎙�7ڞ��ŧ�5n���K�P9F�.��X*dfϳ7�����<��7X�����nA�"�Jl�ȓ-��u���R�Hհ1�%-P�kT�i��$�0b�����`����P�5�4��-���%闥\�Iq���`��!��-=Ȕ0�)�'A��W��A�ȓ#?$I �`_3zk*�p���C2А��,�p���#�7R&-�PPFju��Y`���`ǈY|$�r��җ
2�ȓj:e3@О4|���9�:%��4�*U��C�7�)�f�+۾�ȓ�BU�Gf@��%�zg:i��C:D��a��P�A9�!p� �QI`8@��"D���Ę�7�!�Nr���Cԍ;D��	%WxE��ŋ*:ޒ��i;D��@��W�8�8I0�i׌\5jiYn9D��� %` �bd$@2Bs4;�g7D��K�ֶc\"�P ݳ4��U�)2D�4����1T��Y��AY�M�V��`)<D�D!�eH;~���"eוl�(h�5D?D���e�"`4�|�U��B ZMJ��;D���C˗�h[J��t�CW��thӠC�	j��Pؤ���B�FT�U���8��C�ɀU�(=r�i
�	M&�@�J�'��B�iI�V���zZ����
=7��}�7"O��{�n��u$�7��}��{�"Od�a�KTF)� ÿ1�h���"OnpH�h=5�<-��8Bu0�"O��cO�w��H�c (<� ��'W�I��H8g���4@sE���J �B��+7�NU C��,aG��B�I�d�Bͫd�4x�h�'Y+A��B�	�	��chO�vV�e�QaU�gN`C��t���K�\i^Ĺ�N�i�rC�I$2���C�ʁJ�y�Q�ܿM�V#<��y<�z �E*h)�a0#B3wu����A5b�b!a�4�h �V�
�4ȆȓT�H��������C<%�ȓ83f4�P�ʰc�H�Ij�
�Рm�L�����V�Ld�Jĺ�JP�$�� *B)�y�n�6��eX~�H��H��yrl��F�)�g��*a82�d�yүX)ao�U�VI!~k�ly�O��y�G׀q�,E)�`�fa
�nơ�y��s�&M��i�2R~
(�1�צ�yB�ڂv��aj���0��#����'xў�O��};�#A6-,�(�E�,0��'Ff�
��Ҥj� �%��,����'�Ȃ���.��T�R��v݂h	�'&�@6'�P�bU��`�R��K�<q1O�16응��h$����F�<�T
��n���!�2t�(��u�RA�<	��u��5샰��I��f�<���38&��sB�.,���i��a�<��F̨*��C�.or�KC��C�<��),�,Թ�"�' w�9��A�<f��7g�=v$��J��0��{�<ѱ�̋7�R`��K�70y&(��q�<)�.K� \, ѓ�-*Qn����S�<�Tl��y!�h��ӧ[U�� ER�<	0��E���"�M�'\-P�	�P�<� �D�!k�4
�Lp���+� "OP(�g.��3�D0Yի��wE��P"O8	r��?}�lͨaj
'�!I"O��G&�2]�!j�"��d���P�"O∉ba��rf<
��K$@�H۴"OxUQ�NN�2 r��E�Y���`�>�
���*V��j�sQ�E'���ȓ �L���":l��و��'��هȓl�ı��l�1��ѫ%����ȓCY���u��)�&e��
��=��1�� ]��F��)i@�`��8�ji�ȓBZex�KE70�lg)�i� Շ�j��;�$C�"�F0sMO�pO����%��U�t�>{�  㰧���<=�ȓXJ���I�8P^�u��j-H�ȓPĤD�3�J!3��XA��'��ȓ&�Y�s��r6�y��$mNbą�-�$[���(:"^��'��� $T,��a�"���B:a�ҍ�v(ɹx&\�ExB�)�n��i�<PW*Rq� �i҅^�<q���Z��u��
H	��9��
P�<���D�g��-��i��c'e�I�<����9\@8���Т6�69�tD�<�2�Fg�	9gM��t�[��ID�<Y��Ф:��oB�q�C�k�<铩�Qv�9Z�oM�vaJDQ�\s�<�C*��I����T�WM*�:U$�E�<�!'	��!c#vP�JJ I�<9G���$��@QG�F)]��R��K�<�Gn��o��qҌ׀w�~u��j�Q�<)7�
5�*@R<.�
�-���x�C�F�����Ғt��0�^����hOq������sJ.���T�]i��s!"O��Y���@i0��GnŢ+Pn���"O0���Ꮇw��t8t���?�.�;�"O���F囙D�j�{�~��"O��i� ¢�6X��,3q
���"O�L3Tb�.ۼlJ�K[]W���2��؄�	4OBʀʢk�@�����B2<C�ɻb��c"!^�zQMk#�J-$C�	�)�ՠ��(����cSb�bC�I�N��Dcw�C����z�OD~VC�I5~!K�)�~+�첇E=L/��D=�S�O�T�+F֡FBpBw�"|����"O|5��Ù4g���%I_33
Q
"Ol�)�@�BFp|�f�dZl%3�"O |ñ'�:H��pk��8�p���"Ohr�I$7�2��eً+I�Ū�"Op����PH�7.A�̚�"OT���u��#�m� {�"O��(�@�eR�qmѲ!U���A"O�9���7�f���A��S��uJD"Or �U��1!r�����
4�Iy�0O���N�z�jt�W ��1���Q�!�E8�Q�kP�DB%3.�=�!��K�1PP<k��9.?���6L$��pD����{��iD䄔*[Z N���yON�5d̑5�
ROV�i&����y"�ЙPɤ�z���?4dTLQ���;�y"@:dr��3�@��w9"d됫@��y���u�l2R�L)���+�y��#��g-]�;.��K����3�O^�5��%$Z��:�e?�p"Oj���W4?�%!�kW��(��'Iў"~	� Hq���+KN ��(0���	"O@Ę�����|��I	�}֢�*V"OH�x�W:|��e�
��^�)�"O�آ«�e��9�'�֋����"Or��@�,h�~D���n/
��B"OX̣��"u̮=�U��S4^	R�"Oj� � rR�.��GT���"O­ �!M;d�|kE�޸Aء���	c�OG�qi�*�c~�B�G	����'.�X��`Op��=s��T3�.<c�'k�՘�kƇg�F�Hr�J�I��Lh�'\�mJq&[/��@1e�xp֘��'H蔈�'1W^:0/�<�� ��'	�T���
IP�Bo��7��a�'�����Q�lX"G��4�SL<Y�����3�1Y�Ǉ�i%�=�NY��rG�N؟(�EK�8T�}���n`�!���3\OD� &H5�K,W���:�,@�n`c�j�xv!��g_�و#���Cw(|;�H�2�qOLIʏ������j�ťҳ��]:�e��y�T5P<���йu�������ybkܫYH-aQ�]�p�>l� �-�yR끇a�B- b��pf��W,J��y�Q�KE*�Cd+è|~$ J�[��y��3R����3�ݞx�h��E)�y�*T�ƥ�Ն��l�&\ف&��yd��Z[�y� �P�7E�I�����y��P�U#@ダ����=q����yb⚎}s��E��#�(��=�y�����s��>�n)����y2F� ޢ];CU5�prP
(�y�f�``✁��J�����ဏ�y"$E�6�9�DD!�p!A�
&�yR��
�<��,\  &~q�����yR'֞q)����#�p�pLBH��y�D��]���a�ǌ�s�hs1�S/�yB�A%P�8]c�*�1́9�ʝ�y�C�,�)�`K�~�\�2AIA��y"�
8�hQ����*�����y�M�X���vlY��(9����y⬛�8�K j�Zk��96,S��y⭉���(B�bR�N cB�Ü�y��wN`�1B�:yB��y��E'r��RSL�7���ϛ��y����P�G	�-���*�!��yrD1B���l�4-¾��6L@��y���G-�a�"�? ."��F�Ã�y�G��d�2EI�I)2�X�u����y2���� 12��5z$n���*�y��<9D�U�F��D��l�$����y�e%2�XL��FA*>x�}S�e�.�y�
�=�J��7�R�J����`I��yb��c9�[d/�=B�+en��y���4��|JT`�7;������Z��y"��+�т�/4ĸiYd-W��yAT�}����4���)@��J��y"�nP���LZ�8{��@�<�y",��tl����.�#���E���y�CO�C�I�¿H�.�u#�?�y��W_�qH��Q<*El<U���yr�ZjF�*"�N�1�|�%�K�y�M��IԊ�����!x^liJ,�y��T.i�XU8p��$l$(At���y�ˀ�g��-���^�d�
�j�,̈�y
� (���/V5^v��� .ڄ �����"O�i����f���X�M�3��+U"Ov�3��&
��P�d-"B�p9�G"O���1(��F�-�+_� �Tz"O ��E��_�����)��H�Z�"r"O0�ᗉ>���1"͚u�b�7"O�$��ك2p`@z!A��8%��"O�T����K��H��T�T��"OT�����~:T��Nբ/[	r"O��6�B�IB�N�lR�X�#"Ofѱ������� ��,mD"�Rt"Ols��F,L�(;����3���w"O���Td�4�`	o�!M��y�"O���u!]�`:��� �3�~ 
C"OD�� �ש4w��aWm�7��k"OH���ͳ#�4%�gLc�X��"O�LW!E	�YE�=�~�@�"O|���j#
���is���\�8�ps"OV�K�$�&#���0Ȗ�Eh,�c"O�a��o�al4�C��Sb<��"O�������L�i�Q�͌;w����"Ov(�BN���r4��3^��� "OȀ"T�ɨq]�e�A%�y>
��Q"O���s�Χ ��5�Uc�!:����"O�h��ALV�4�KB���g���+�"OBTSg��bCdA��_�"eɧ"O�l$f�$�6i�F7#�F��T"Oȫ�ҢKL@|�A5V�|`:e"O�	�� �'J�9�l�)B�%��"OJ�ٔ�J�(�6승V�<��"O�(P O4{x�0�*3S#>�rT"O�AB0�07��L��I5*-��s"O⸩���Y|��P�C8T��R"OeB�>8M��j'���(����"O|-z�I�pP��8���?����"O������J�(���AOF��$"O4C�( �fQD��4��{��T�%"O�1���T@��@�3�f�zc"O��is�҆)�(I�]�Qqe�"OZ���hѹ,�>A�"��2U�9��"O�IѰ�E� �X��%o")��"O<{FÁ�o[��G��]�Q��"O��Z��U��=� �*#��9�"Ot��W��,d���Ex��(�"O�u���'�:��f#J�bt��"OF�� �S�R�84җ�H}R�y�"O(�
;=�r�b�`=�p���"O�])F�(`8>m#��Ϋ4�⡻C"O��� �I8��\��0�� "OZ�`W�	�Is�h�jć!1@�{�"O��bl��-�BT�B/%&��0"O�q�J���h���-橢�"O�����?2z���J�zE�*q"OP�hE9
=6P�t�)��ŋ�"Oh%*��l߲,g��	@v��H�"O�Pۣ��am��.d0��"O�����HN�fш�g��,��D["O$ԒRJЌ
�&�9%h�*���r"O�8�sK�|���gFI;=�"O�� L�+�H%S���S`lyІ"Ovܒ��G�S2�lXU��I1�{"O$t��eȐ"�`��*[h.l	z"Ox��fEb�x�+㊑$�$%�a"O~���J�~njA��>u���0R"O� ��͋�3�x�" ����r"O��B�>�Lk� L�6���C"O�]j�@�q$��#��=~��(A�"OpX#��\�clz��FiΊ5F��R"Olᱢ�X�E^�X`��96��R"O�(��-�)YI.�8��S/. �"O �����N=ΐ�«��`�����"O��
1̃v�$� �,��Ub""O�HU�@�^r虱�G�,�Dӡ"OTI�@�
~H�y�A��&ţ�"O̔���Y+
�� ��;��tzD"O�e�f�;I(��o�"x��i�"Oh�A����J��&"�4�zF"Op4hh�*vK���G� �h����"ONH"qhD�[
lxQ���m�f@��"Oj�i���w�����c���"Ox�Hf�Q�`0� Iw�,�V"O�ԈT�J�[��T�Hԥw^*ݘ"Ot�k�\:4�U'�[>Q�d"O���F&0B5
f&)m��"Ot��7L?!���ԅ
�8��"O���b�=� =�F��y��I��"Of��Y3�i���4	�����"O�"@S�q5R���\k��"O@h�r�*)�$����y��"O,�aE�	�}�T�� Ԅt�x���"O��R��V93l��W*X>3$zȈD"OFQ�c��hvHX�Zr̒�"O�mZϋ�tB�a%f�(>h$��R"O\ؚW��@.Hj%vs`ԑ�"O�����m�$�� ^�`� "O�3�AX��1�J]�o�&m��"O>��qkA�V�����U;l�L�"Oh�Я�?�,�!&	JLX�!�"O�*!�4f�,!�@��X0��#�"O���!D4d��e��W0 Q!"O�����(3P|�caTP"����"Or)�GP�^�5r���
����"O�=N�J� Qӓ�ڒ�R��t"OLӑ�:c��Ċͼ���"O��R�$*�Ku��Y>�s�"O5Z��'&N��&�x%4	@"O�Ђ��&4T��䗞��B�"O�zg60֦<q��phS"O�9S��>4�X�VTUJ0"O���0�=sF�CQ,)$^��@D"ODxI%��?ޠA��
U�Hx�*"O�p ���_��Ps���%Wvx�Q"O��xuC��+�|��B_;DgP|C�"O�Z��«[��%�%⊲U�X��c"O�%��I���E0(�L�6�� "O89s$�Xk�Tr�� g��I#�"O�uK� ��('y�\2of�E�W"O�S6���Xުݘ�#��J]8���"OT��)O5xJ���DZ�T
�+�"Ovy���kwr}#�!��02�p��"Ob���-2z;�M�5`�+Uy"O�J��*�`�sR�ٶeBșa"O�$ID-U�ll�Xàj��N9E�""O6M*ƯC�*�PA��I�.�p"Ol�0uH�y���J��X�O�ʌ��"OmF�Ѯxx��U*U��� �"O�K���$4�XZ�
�R�X��"O��`�E�-H���U
]&P�d"O� $(b-��?e�=�'�W�Z"�r!"O�=P�BLC��A$��S���Q"O��Yb��O�͈s�_0Ʊ�7"O�|R��ڔ� ����9w�`��"Ot�p��@��<˵a�~�0�Ȓ"O�2��O���rៀ	{^䠕"O`����\G�@�B���|�l���"OX��5g�d��o�8dv�u�v"O8����+�m�d�@��y�"O����FY�H������H�ܩ�"O<U���K��4���bK+|h�}�'"O����G/=��q���i)�(b�"OD5���ăF�A;��
�6%>}��"O�
�GE�k�Yh�lƍ"(�v"O�a��M�ec���Q<<V0l��"O�hVn�0�B���J/5:| �"Oh% ���S�¹Q,K��y҆ 9>�0k�z��1����yRE�@�.�9��Ҏ._X�Z7K�"�y2I��F���8��4%�*H�6H��yB��yҚ�Rw�^�!"�(� .��yBዌ*�Yy�nwa���y7�QC�'�\����<�(����A�� C�'96���F��Z�6�ig��S�4�	�'��J��#4���f�@�y@���
�'��8�惡'*䀺�F}H$$�	�'`�MP��D��iz�)S u��-i
�''a0��G�mꄰ��i҈i���	�'<D�pT �2HnP�Zc%*a�����'ԉ�F'�$��	ѮghМ	�'�KB,]��y�.�C&�s"��C�<��χf� %�dJJd&���~�<���Ι:���*R	s��)���|�<�A�ݹ~Pfب��^����i|�<�Ќ�=A�z�;d�=%���"'�m�<�!!�
@���
S-A�1�éA�<�a�RB5|����|H\��E��<�kE�	=�t9�A@2�t��Q�]{�<A^��ع���-b�p�	� z�<١���?��� .��e-(����t�<A#�V�IҀ��W�D�j�]�!Bp�<�M.s@jb��v0f��Ddk�<)�+	D�d��ԡѮe���z�	�`�<)�'U=#��Â?M�%I"�\�<!��f��j��C!{}#�AV�<����X+Hò�Ӗ\��	;�e�w�<qƋ�A��Id!�B�xQrm�u�<Q�_K�HeQ։�:z��T��(�p�<A@A+W�9!����c��A)Mx�<a B�Qټ����"�`�hEs�<��l�o1:|K�%��?{����S�<�v�͆r��a����!L�X�MR�<� �6m3n,c��&" ��� h�<a��|�P ���	2�ӀhQc�<�G	�Wr$����.��iK��w�<�U�[  ��X�Á�{P�-�c��t�<�Ua��.����`�*|��U�u�<)R͏&Y�֕8�)�8��X��.r�<���Y=DҾ�B2��PJB��G�<a��Nm�
��JΆ	��t�ԍ�i�<1Ĉ��B�Hm���P`��� u"�g�<�q��:qa�c�.ψ&��+�*}�<�w�J�& X�f�bݨ����Px�<�S,ԿI*6�3G�'e6}s���K�<� �9� ��̅ &�Q�k�N=ɤ"O����#��X�"|�箓j�t���"OB d�V��8�$�ss���"O��UDW��1�b��ccr�"O<}"Ċ�`�C��P:Px�+�"O���ׇO�,�@��J՘<Y�"OlQ��H�kI���âWV���k�"O�	3��A�x�4��&�M�����"O���%�(]n��뗛��))R"O�y{q�p_$���j,^uXڃ"O
��B��)kT��sd
3^Ϻ��V"OJ��m	����t��KZ`�"O���F���Ov�`I�G#8;�Y� "O�e�EG�1�9Q��b0bx�C"O "����
MZ���&^ �"O���B���A��]�D*�U T"O�A��a
,1@�Z` �%!ڌT"O"X�B*^��A��{-b!y�"O���D�\�n��<X���e4,�"O��ȵ"�>A���S�	��r�>��g"O�d�D.*!�jx[�.-8�4��"O�͠�A�Je����Q1v���9�"OL@9�Jѕ6��bv�^�%D���"O
�xT(R��i��F?\��9�"O���"4��<B��)jԽʔ"OrX`�lرBMH�s�o^�5_���"O:�i�#��>��I!�X�J?�٨"O�D�Fe�%$H�GLT�9 r�r�"O��	�aXh��P$b�?�X��"O��၄�0yp��d�K � ��"OشyF���_�B$���<�X�"Oj��c����-Y%�C�uטL�F"O�1b�DΑm�9s��=Ɔ��"OJ�sL�QJ���gᙴ�~�h�"O�׌Ηcm�`�b�Qn�L���"Ox\�I���T���^)S΀0�"O�����)g���P���9H�D���"O�ȂL�8@��T�ݴ�b�K�"O�X�f�l]ԭ��E�pԜCs"O� �b&�Z'��ψU��B4"O��RcC1c�@Jg螡2>'"O�,T*>ta���Q�sA,]��"O0���M/�|P�	E�46`��"O�) �ʑXN0)��)>	1f4ӗ"O����W>w�@���G�3-��H"O�]c�N��)!�AB�g��2&��f"O�hC'ȅ�fW �I�F%�9�u"O5�u�-�V�{G�KB��	�"O�u����]\<����ӏ�4[�"O���A��v��K^֊Q�"O��+Џ�C�Vq�՗73"�XC"O�mY���ic�A	;LN�p"O�-���v�j��#*�"O�pӯ�g,
8���?A�m�"Ob8Q��B@�\X��?)�lA��"O��avhZ�d/pE�G�Ӊ)}�x�v"O��� ��z�@��Ɍ|FDj@"On}��z�%ƞw�	� �;�!�$ɇ(����ܮIj�7M�;n�!���5%�]#ISx ,t�c�X�>^!�d�T
�#Re�`�lQ4JŪBJ!�$;���0�$�/��a��
!�D�p�y�d�5T� �ԏc5!򄗚�hp�6l !"�1ȠcE!�� $�;�A�#M- �G�)�H�PC"O4��R���!t�i�s��5�0�"O�u�Fj��e�^��6��[g,J�"O����D97(��V��zgĐ�"O�\"�ǚ+C{�=a3cC T�<���"Oи��,�+����rçS�:8��"O�M���ۈI{ի'j�$3f40�5"O�%�3d�<�����"J�)�"O6�"�E�R���d̮+@v]�7"O�	2�%������U蚋9�\"Oʹ(c��1���sa��#�t�6"O�dA  �5G��I� ��J�"O�Y���䨐V�Ç=�2"O��u�5E������B����"O&��$��m�ZHb�a ^�v�"O��O�1�B�6���SS>�T"OnA0�E˾��x���#"O,T���Q����۠.Q1/<~�2"O���u�L/?���� �*D%9"O4�B��:lv��'�؈\��!"O�8p��	��:F��%�Ĵ8#"O�Ӈ��/�0�1s��D�ʌ�"O0�M�"�����M����9w"O@
� !!s�p"�g����e�"O��R��Z�I.�yR�֥ ���"O�8-��L�(<9⃍��Es"OtTr��:|v \p�C���mHT"O ��e��)*�P���� �"��"OB�kq�M�y0�%%�Bi�,�"O�TR!��$~�n�X4d�xO|BP"Otݛ�.B�Iy�u)�B�D[
a�7"O䝱���%ikVY!���kE�-�"O�2e�Y��4�R���B*U��"O�	��`��@�Qqj��՛�"O(p�4N�x 5�!fF7i�n���"O����?8��E(~{&e!�"O����ET:=v%�u�^ �6x"G"Oډ 1�K�D���  oѐq��"O��7�̪:� �QG�����c�"On�R	,����u/�7G�@�"O�F�-{�PP��{�^���"OR��p#ɘp\�`
�d���6I`"O�Ƀ��гRDH�/�vLZA"Oh,���?X�\�#� �����"O����Ú�+`Qy�ڰ�"�x"O��Q3�A�9�^,Bp��>���؇"OJ�	�j�9(��(���V�\ �lá"O"�`���:9�x���k�9
"O�P�a��"u�%!�L_�k�Έ)�"O�R��I#S�T�����D"O��!��FҸ��
s���v"O, ��NS5tɈ�Ceo	�����"O�	�! :Z� �薟p�3"O�`j��!v+41���#˺�Xf"O�m��J'Ae��� D%��CQ"O�8�
�y��a"u*K3D}l�36"Oj���H_�0Fb<"��9$`|�ض"Ox4p`"݄o�5;��×Y%��P�"Oj��!ܮo�i{D�%K���C"O���Yi������ێ6ܣ�"OJᅒbς���Y��&`@�"Ox1B�B\�Q��c�h<A�T��"O����Ύ�6%�G�ŧ_ �LYq"O�Ȑh?T�0]�"B�j!J��"O� 5�q��i `i1��Z�&"T	T"Ohl)�� ET訁�I�"5"O�p��w=��1��xb�Hp"O�L7MR0*TX� �i�?S�V��"O�!�aL�]+�Y����m�j�S"OB���Sz��+�.�R-#7"O��)7�W�d��{v�Q-6"@�"O��j(�]��)�M�R|!y�"O��	QE:`��}"'��\t s"O��&�T?<�~mKC�\�"�y"O���� `��Ԋ���t|0a"O��s��ڵmMp��EFq�5;�"ON%ҖC�;J���3B��1\mv��"O����kI�&��0c'֦gN��""O �{��O�]��P �&ݟ~?�i�"O4�@�Z4���&U�((x�7"O������5q$X�A�̡:"�}0"O�օ�F�h��J3C�ri+�"Op!��I������Q0"O�ݹ��?ڦ�p�D��Q�
8	�"O$�p6�Uْ���R�z,��L%�y2+�nt�#%��Gaj��ƌ �ybKJ�WH�{ѧ�6F]�Az�d��y����	��:����lZ%�y�DU?"8R1!Qc�`{�G%�yrBQ+fbN���'��T�n��_&�y��
#m�6/V6���a4�yrĆM2�I
̱K�Т�!��y&�Pq��ht.
�pT#�B�*�y�0c�z8��%H<?����aϭ�y2�64Hk5�ɩ=2x�n��y��a�`2�O�9^�xJ�D�	�yr�Ϸnp=Z!c�/Z4�0{����ybj�K�F�ä�DZ�&��RiO&�y�(��Y�y�sJ��Kx�e�H��y�ƒJ�z�JE8E�~����?�y�.GW�1 G枱n�([G���y�D�t�*�`b��g���d^)�yB�@�P'ШT)ֲd9\������yl�[�f�͝�	iP��!���y�T�.��i�d˝�r���0έ�y�V�@7�u��)Z&d��T�p_�y��O7�v�GiC	I厡+�c�yb�#>`,�FGٮ<BN������y�AĸX)��]�K<e�S�C&�y�!��H�YJu�(��uX4�]��yb�J4-��!����;*��Q{Ӎ��yB*E�$8,
7OR������"�y�)��A۳w��z����y��Yan��͕�t�j�@��y�����(��� ���P�@���y���Z&@�b�f��ր��,V�y���/�N��Ѣ@��zȺa��y�ցc �jQ(|J���p�3�y��N�C���描?�"���f�y�H�h��&G�9�$B��W�y�c�<-��Q�$�L&_?,�P@(U��y�C@-*�1�BR�� �����y�(Z/�T`V�L= �^��ƍ��y2lȚJ���r��1' �x`��\��y"��!"�fH+qH\�n�|yaQ�	��yҊKWuBQ���	m�a0΃�yb�T#ʺ �� ��_�L)(�@I��y�+U�`l���K ��!�G�S�y
� ��"7@�>/�!!�B�I��Pa"O��*��
D�����Wl�!"Od(��D٠P�ޔ�o.?-0��!"OMȣ̃	/��yD�E�{(��("O ���j�1t��g�P�^$̕��"O���3�@LÀ�k�g��j��v"O���V�e$�Y"�-��z%i�"O:p�!Զz������3��e�u"ORsD�QR�	�d���`i�"O�G��3p�]���͚�XA"Of��H�5#��m��]�����'�Ԝ �](�l��.ƈQ:^�1�'��j��B%
���0��^�ԍ�
�'���1���?��q۰ȅ GlN��	�'��tB��LY�fȳu{�x��'������L<���i�M=k�����'?H髕��(rf*`e���:�v\��'IP�o��g-J�Y�795"���'����RL��y�-й6�Vh��'i�8�P87�!�fnȮ=z���'��}qR
�<Z-Z&Β:e" �h�'a������\~��"l�f�x���'R^�@�X�x�B�5I�6�1�'B(��!ʬC�2,�I/#��M��'�jț�U�	��h0���m�Qa�'�D��.J5IDT�� J%d���'ƬuB/�	N�P	�w�\.�|z�'t]�� ��N�F��6��}�<�x�'|�Ěf� K.��w�>C�X��
�'R�� �O[St��G/8?k�
�'�9��*J�\�|䱆ۿfƮ���'L0�ӳ7 d|�E/���Y	�'d���F� 1@A��T-i�'���(��E�~����&�fm1�'Y�r�k��Y�$T�R���J��'��TRMS�V,�+㏨=R!`�'/^�Z�l��u�*��u���7�eq�'D5W+֘�������-��q�'��I��
���f
�""p|h�'Yp9p%�/l�2�����XD`Y�'g��j���4{�@����Ml�	�'�������{2f��a�
��$��'�j��!�+F�0��(ǡe�I�'��(��P(ĪEq�KKo� ��'m�P[�����7�Z�:b0�'O�d l�OT&Qq�N#1����'#��1�(�=iLI`J̌+:���'E�ᰶ�Κ\p^x��T��D1�'F���%H�!h�!�RF �`�'�V�:�O@�5H}���I�� ��'��%��%��c6�;Qu�<�'t8�����s��0S( '��\z�'�D�v/�.��8z�O�MHx�'I���IY��ل� Rv����'K��3T�gUؠ⣌P�J�
�i�'w,y֦0 q�p���H�|I�	�'*
��w�|'|!+ѥ�6C/�4�	�'��<81(ǆ0������
=0�AB	�'J�$�ь��<8����O0�i�'Pd�׌�?}U �1r�9<),m�ȓ?¾t:�\�\�:q����)C]4e�ȓC`��Q�Γ1&��s��&X����ȓ:m����g�:�(������	�ȓS��9��ϓ[�<u�ѪMgx�<��S�? �u[�O؟FTF��F��>z^R�S�"O��QL�7�"[O��J\��"O�����b?��2�(��S�"O���vEǸb��x;��Tk��i�"O��!�A</"����%�h�2"O� x�%��&��H��ė~ҹ+�"OJa�Hێ�z5�A	u*�Ӕ"O����{�L��m�����"O5	��^�O{H�B)���J��4"O|)�C����(YU���Ll,K�"O4���㏌.�"HSE*QL�P�3"Ot�Q�J�P�P$)�.[�ڰ�b3"O���@ 'C"�8��řf��A��"O^��5n߯d&& ²CS ���r"O(�@1Hʭ�	��B E�@ӵ"O��Ѝε|�Bu�AY�obH��'�֔	��E��j�n\#՞t��'>�����L8y��)�+	�T�ʓ3_H��Vl����׌�^�8��x:P%�͗d�j๗h��H��l��%��	�l��%W��ѡ/�*1����WL��P�V�R4��K��
l�ȓ$��x"W ,f^ zW�Il̮<��D�NQ�5.�35�e��z�Lцȓİ��1�d$�Âߏ	�p��ȓO%l8Qa�#n�hɻg�ލ�^u��O:���U-�NL�<����)@����tɂ�CW)�OQ�Ӕ��ȓ�\�u��(cH:��W$Y�?�M�ȓ$h�I��e����e]�t�rx�ȓz��Y
�(��Honqɖo��$�ȓz����$K�;7�`a���& :5�ȓ��4����(<�\)���${V}�ȓcń��LAU��-��)�E��؅ȓp���aƭ��F�L���&O�,��ȓo�Vq�����N"@����4�ȓM�.0+`	��w����K�����ȓL<��G/f�c�H�R��ȓVVl���)U�`���#Y��ȓh��c�Z:nO 8���6� ��ȓM�b᱒�5�l� ��r���ȓ�d�JB�N�U��,B�	zd��t��PX��p	�L� ���d�L���L�`���e�h����rfƱM�����c��Ұ� )D1�[��`��ȓ]&@)t(Ʊ2�*�e��Ȅȓkl��Z�iR�?��<;P�|�n��ȓ/,���	O\��"'eL=@��ȓ5�P}btbJ�,P�b�K�Z���ȓH�lȑb�K�b\��#	V@���sf�4'��^~B��Gڽ. �%��-Az(@j+�j�G��gUb���L�ڽ�&&��|��9I	E��N�������K��V^$e�L#@X��t�Q��IX�l�: ��p}z��;�	(��\���!�G3�a�ȓ]Jș�M,,�Mr���Қ<��76�`��]�!�,
K�T��ȓh�\��$����i�^�<_V��	d��$I��c��9F`ӱ]�y��eHQ2�M�����c�̙�4�>���!s���et��X#j�%��̇�]�݊��Ǚz���p�c�:}���R��,�萈�s+�5��S�? Ұi�G5F[�� L(�ɱt"Ol�p���^b�h茮#ء0"O�e�r�ې4s�T�@e�j-<0W"O"�4嗢B��y"B��$hUB"O2M�m��a~�4����4A#�c�"O�虧@M�hEз�H"�"Oub�D�A�8�I�fF�Nh}8T"OzP�6g�
�t���;K�~9�"O�uk�J$`�e�C$)& �"O��s%]	\|m�!�ԷS��(	�"OF-���\�d�!#���qS#"O*!{Q�G�����C��6a��dy�"O�5慄#$έXR�N������"O a"�އz�r+��{��]�u"Ox�Dǈ�O��ڇ�R�QR�*6"Opm��3S�"�1 �
�D��"O�qk�@��"�E�B�� �dP��"O,�[��9ox�� �\H�~�)'"O���AY�eGTĳ�G@ �"O�);�)˲Z��谔/P,2����0LOZ�#ӍE6t�y`�͇T!а0E"O�Qb�'0Z�Q��O�&��aq"O��yC.�rH�q�C�8��@�a"OfD�"�K�u�y�Ս #A��$�"O.��t�|l���wB�.��e�"O��x3��F���
�AY�c��y!'"O�t	Ө�?U�r,��/�N֌�z��':ў"~j�H_/e^A���~!�Z���<�y���:n�xݱT΀*T6�����yb�+,�A"���)��0!bcC��y�J�v��
��8E��*O��yr�D�Zz���DA
��<�����-�y"�Y�a�ͫ2�L�xU��S�(�y��%%O�1"'�uۚ���e^5�yb��=s�fm�A�	@�Hp�����yB�K��&�;#�#P>U�4�B|��np4gǜ>M�\�H���?آ���h_�`t�4h�$|h� U�ń�A36��V��^���@�M�i�I��D�4SeG§8����m�pFꉅȓ-��`�t�#4l��î��}39�ȓC�Lժ҅I�k�z-���5<zP ��Aݾ�q�C���q�v��1�6��ȓ{xZ�@vl�=�))h
|����ȓ�B�Q�
��yZ�-\c�E��]�Bd��l@7��¦�טN!%��N(nl�T�2]����X�BMLl�ȓ�`��O�sy`���jн`�vŅ��
8�AGج�X��A�L���	�ȓ7c(�2���Չ@�؈�v�]f�<a�a[�Y�T�"kQ�mL�m���GK�<Ԏ8X m�7۠R��eiG.�K�<�i6p|������*�N��L�F�<��ꉄT�^|
� U� %�t���L�<�3�.�eIBX�_��� U���<�oH''��@�@E;���1��G�<���" ��yCiJr��׫�|yb�)ʧL�h��ǠU"���iQ�N� �p�ȓobԤ%���Ev���ځM�D�ȓtJ�Hs�G�Uf�M� 8x��ȓ�^LR���u���A7���ȓ*��L���c:�t�Ei	)p�.Y�ȓ/2�a���e�$��f�)j� ��^ƜL�6�֧���!�@?O��)�'�ў�|� �s�%�!r���'�Z�/�*I#�"O��Cb)޷n���3��$s�څC�"O������
}dx`�5��?�hR"O�l��A�6<��)94&�Q��5�G"O��K2�
q�&#�O�L��a��"O~�b�LA�v��!j-����a"O��!l���0�T�Pp�g�'}ў"~bE
Q��`���3T���&��hOh��O�q.ܑ)k�z*^����!��/g�F���!@9�Kһg��8Z�'�Nd1q�Ӆ�D���*d�0�Y�'ru�튂y��I�ͦW�q��'�����5Q�H� !N�Sz)��',4����S�Έ� ��Lx��:�'�l9�6.�|�@��ુ^�-��'� Y�4�_ ��pP��8H�f� �'����F� NhT���Br���'z�,�w���/����������]�L4�U��#ʘ�P	%�~͆�5&�if�M*�t���:X �ȓ|��M��Q��EζМ�%��D{���ȪM<6�P�쏛V; ��6�?!���'0��k��N�2��hz�o��֠��'cH�!�K�Z𨋴(M<����	�'j�k��N#/�^l8t�E?xk쀀	�'���,L��<�4oE�r4�L(	�'�܌ptlUSv�֎݈S�B͢�'r��	���<C3f�ж�O�bшH>y���iF�n[����6X�x ��)Y�Pg!��K�b�Q��F؃�)�DL�K!�D��-��)jC��$L�F-Ҡ@��2a!�ZLn�`B ��D+�� ��<=!�$èq�8�Zp��v%M�A*!򤓋dG�a#ҀpHq��-S!�D�-6xt풜/���0(R���x��(����p�ːS�R�sh�T���j�"O�H����^U���U�Ҩ]o��9�"O���'Ȏ� �0l�0+tUpH"O����p�d*ݜldd���"O�9� ���2X|���<G��H�"O���v`� {p�����g��}+�"O��r.�����K��s梑�p�'�ў"~:'�x�q)r%
��K⚇�hO@���7i�()�[�J+n� H�6�!��5yT��`יJ@y��"�!򄚩l��٠��ިD:���CY!� )(�ڹ0j@`R\��L�_�!�$���I�6���($�GL (:!򄎖"FZ�"���	|d*���-9Q!�dJ�zX|��L�)��q�U D*1!�$> JJ��Re�.���� ļ
�!�d�*T� ��,,[�5k&Oώ-�!�dD>��M����[�4�yc�Ւ5�!�$�(s4�{Aa7��$a�!��Z�!�$�`�-����v��H2��ۚ6T!�䐯�����] }���mE�:!���0���6�M* ���P�Q\�!�7Gt�Q���c�D\Yn� �!�2"Z�t�S]&�vS��\�!�DY�`fb��e�>��j�	V2+!�$Ғ7�1�D:0����Y�e�!�$\kܨ��'�5l��e-Х=�!�d�!y*�-��>�^��F�)w!���XU.�Cnʅ�Й�����!�� �uPaJ�8\f�!;�͒r���q&"O���ꊧT�������<ի�"Oz4sfH�K��r�����Xi�"O0��B���[��L�f^�@��aS"O��pEY�aȌX��kz����"O���4��cD�D�q���"O�貔OL�@���ã��k�&�	"OX��ƫ_(`��\a��C�qۣ"O�@�qCI7��ua�̞�q�mz'"O�Ig���@z ��K 0	���U"O��S3G5%�|��
PT�}SQ"O����`J�T� 0C�g��|����"O���)��Lߘ�*c�V�)�"O:�1��a���[ ؍U)��6"O�V��4Qʅ�?M�|��Č�B�<�#�9r?J�N:6��r�lVd�<ap��.r<:c$��A?�p�A�Xv�<�%fV6v:J)WB��&%���Y�<�#����p%�K<G�U�]"�B�	�rB,A��,[9M��5��d8�B�[�(fȂ$O��i��x�p"OȰ��� p��3�V�(��!Q�"O��%A�B�yb��?��D�V"O�@�whD��P��Vi�����"O�,�6B��"�P���IK�}�@x��"O�QBWU*�� ��@j���C"O줪q'�4Y(M�4��8dy䝊�"O��{�d�s���+�$H==z�#3"O!��
H&R00=�A�$"n���"O.̲���!o�%�12Z±Ѐ"O���`�wT�a�3+S=?�<�h�"O�����\Բ�H�
jzb�G"O�I�S�_�h��Q� �ōM�����"O�ؘC�9Q��2����#��8Zt"OV�sF�]N)�x�G�<5�^!�"Ov���JSJuf�J���?�@��"O"P���:z!^)�T��,�}�f"O��5��
=��lQAŀ��@\�@"O�<�a�	�dӪH8.�I:�l)�"O�{��@ ��䁀�C�#3 Q��"O� Y%k�_�hDܛ1h�ʠ"O��{u T��x%	�![��ɒ "O�@H��r���M�$\�i`"O�-(���b!ڤAVχ�c�y@"ONH)3j�i�h	��K��K�����"Op���NƦ�(� ժ۴!���"Oؠ��CY4-l8���S=����1"O�`���ۜpl��j3��8��|k�"O�UQ�EH�%@��j6����"O���ܔ-H��f���J����"O`x�#m�	b̬�%�\�F5�"Ov���Lؼ�)��d�Q5"O쑑���ND�՚�F�:X`�x�7"O���e+�;~��EXV�;S_�X�b"OB��f�8���.AVJ1� �y�n܊l�̬�U/��z%�e[�B�2�y�ݢ�
J�'G�x��0��k>�y�;4����k�q"�RF(���y2
ɔY�H"�C�m@�t��ܕ�yR酖J�b���a�
a��b���y"�*Ax�ǥA�()k⪀��y2��8i,�r$Y�p�x����?�y�& ,�Y7,��Q���2�yr!�0i���㩚��jh��ꐘ�y
� �!�!b�/_��S��5!�6|�"O�P�c߽K���t��'�(<��"O�![��Y�M�"u(�L�4K�TM��"O܌���I;L0�13�E�&�z�"On��̕*GpU��ݢh�VШ"O\�5��0^,�|!���[��P�"O�x��T04��l�s�֥yd�f*O�@qq�-8H�+sBM1��UI�'�4�2���#��zGl�!!��mS�'�>�i��9wy�xW ��-����'�(#a�+3oF��Qc��
i�m��r�ӇN�#��ؖ��1X,݇�_.�Բ�l՜�ȁ����t��@��HaɅ;~� � �M8W��A��b�HA�f�ռ�����[
�8��g�u��ب+A��Ԧ0���ʓu�)c�'f�rf�B3W B�ɖ|�PͩC���A<*�gΈ�2B�	)hEDA�s�U93�����M%n��C�ɉ\��BU�ۃ���rB�	�XK�C�	�~}�҈�3* ���4�lC�;H�����;i�ҥnн��C�7l���i���<3�1�A���C�	�v�eY�KI�B1
8�� шu�LC䉵:d�8	u"��)��a�R�8�(C���\1�� B�21�#��nC�/Ma�hC*_e�28!��v��B�ɘ��Ȁĝ�v�ͫ�Q8B��B��" $̤9㣊�*��  �#�jB��!/�J�Y�+?.N�X{���3�TB�I�,2Lr`��<{Ԋ ��Hгu�B��5O��1.]�rQ<uP��Y�C�I��|�`��[ 2=x� ��G[pC��[��Ͳ�"ǀ:_�)#Y�:C�I:GF�ٹdj*ogF��Qj��\B�	�y��S��`6���=R_�B�I%@�ͩҧ�1y"�#r*�fA�C䉮�HY���G��&�P�*ǃE��B�I�w�h���ĳo>M��@	�z}�B�ɝ{hڍ\70E��cH�h`�B�$+�5s��|6I�4IF=�B�I?�"\@%�W�^0]haP�3,B�	�RD ��
7ms$q!3j��h�C�<s` ���Y�Oz�����#n5�C䉴U����6�ҋf�Q��`Q�i��C�	��|��c��m��9��w�C��#UCfq�q�:@��aql�)8�~C�ɑd
c0Ve��tS�1p.bC�I�mg�I���!&\A�J7s�B䉍f:�`Z�ܣa䑷�>h��B�	�l�,q1�!��Y%O�.aЦB�I2=����d�;Ġ�/'`�h	�'��K� dy�s$�l�h2�'�RsuB�#kf��#��N�	�'W2P#����z��1���L�y_�c�'4��1�	4hx*!����w�ڵ��'Mj��ׯN�,����㊃ p�i��'P�c��ڶ$C�jB8`�>)�'���J�_}�t�yq�Gh��X�'�ZX#�P�.����Ց)/f�!�'V8� g;H���î�Ԝ��'* �Y�)�O,������ȉ�'ub:�	O�I,2\���!
m����',�(ID)=p�"���jf��
��� f��cf 5u�~`pt�[�<]�@@�"O��R���$]�X�ˉ}[r��r"O��CA3�0�ѳ˜w>�tcE"O|������k�xD���:LP#"Ot��7i�1e"ްaE#Y�&^�+�"O��p(M�2�҆��<5��"OB1:�ց�\�S�A
0$T��D"OHT�Eu �9#���1L�P|�"Of(����KvVu�##�)�l�p�"O���U�jIp��Ă��[@-�"O΀Q�08��y�bU&�i��"O*d���,�B!lOf�4C�"O�x��%M�Uľ�Rb���\�*�5"Or@��!Q�\��HT�z� �!"O�؋�-��Y-b�bU�O&���"O����@�=蔨�ƙ�4ݒ�W"O���4c�0$���E�ͽ7ɴ��"O �JJ��|��ʨ$���r�"O�IK�+�"�t�X7Ҏ%��"O<����<�+� �M�<-a "OzTr����P�Q%� ivz�"O\,;B/H�=N�H�Q�O�S�"O�+P	W!<�-e J
~�"OxM��"F�@�e�f$ѼQ�^@�"O ��`�>r�,��Ae:z{Vt�a"O`��e��DE�dpO	&�ja�w"Oj���n�:?:͈���	IX��T"O��cW"CQ�T50�cƥO.Q� "O�a�kX�U(����Û��j`�"O��@�i?"��q�| S�ŅI�!�d��.��#�G�Kb��q�V�`"!�D�;[�,pi��E�]��5��dڨt�!��3�lJ�G��Uw�8����-h�!�	¦�� �V��0��(�6y�!�X8Nr5P`�ǃN���#5ǔ#QK!��?�ޡc�$�,����A��y�!򄆑t��-�0�¥Rpp�0pDÌ.�!�d���X9�B䊻nb��	C*�V0!��63���F�LI�{��1 !�D�*����Gjә0;ީ#g�[*!�d����@R"!�W>����Q�I�!�䟇i>6�Q�+ɂo�8�
@�O2F�!����h,��KJ�l�<Q#5�w]!��@��l�R-P
rOt�ۖ��'�!��)���Aēx`�IucI!�!�D
s3�kb�[�X�<�⡍V�!�ʭ#!<�s�ٲ�Ay&j�<!��ϓ[�5q���Bu:r���X1!�D�{t��@�Ek��@�b,h�!�d�[\��"rm^	=@�c�ڇP�!��2A���P���'.`�AGJ�L�axr�=���̓G�è&nI��5��u�ȓD8t�P�W;-�`u���G�nLΓ�?����i��v)n�@�� v�
` ��A�n�!�T�r��GĂ���)�5���K>�
�C�B]���>I2���C�Ij3�B�I����Ğq0��d�-K�`C��z2�K���
A���ᲃ��N�JC�	�T��B�)�0h���$��=�B�ɺQ��@�s�D3 �^� 2&����=!�'^�>��$�t8�WWp�傴��JY�B�I =m�,�"��*��UQe��h�rC䉛p�R���=E8l""�Nh��C�Y��Q�,	0wQR4x���԰B�)� H�����ci�������Jx�0�"O�q�`I��-e  A�ƀ���a�"O�a�'��t��Fn��v`91"O"�xA`��Y=vѹf*Tz� Aj�"Oz�u��\h��jcn�9�"OV��$����"5H4��S����"O��sg� cl$1��-�rS>Y���i��dD�=��� �Ņ�c�<cm!��'�qO�9��ʧ���R�ߦ}Z�<�F�'A!�� 	zN�4Yq�_;0�i;f���D)a{����(`��@-�,^c�y"LLS��XD�$ď2'9�@���'�q��ø'�N"=%?%�Ӭ|-4`P�OI�ZMa��ac�G{���Y�=�h �0dCG�it��C�>�'P���'�����&��6ӄE�7��9����.��{/t���m�w��d#�	@26@�d��4g=�J�6����_�[BE{�Mߨ�L��@Z�o"�|as��/��x`"O�����C&�q $�%2=l	�R<OТ=E�4���4�"��$���8���y�E�A�Q �+��"uZ�2�.�>�HO$��$�?0���r�/\�'>dA$�r !���V�8-�4��u$��s���!�D�xv0���Mت:<�x�)$�<�<	Ǔ5��mz����(��\%'�Նȓc��|JpC�%2$$���ɸy>v���NUJ�b'��3b8����0�Q��x̓w�PF��O������mf�E0Fj�QvD��NQE�'�џ�jc�P�
Sz���L��6�Q���'�jc��i�[�OJN�PR�{��	�����y��خAʵ�e�ҹm�6Yn�9��'�1O:�|R�&�*�J)��	5L$P����}�<A���+�T�Cd^�%���� E�~�b8�P��Q9,�����d�+�O��O|}��ɲ=Kg�ТN��['�x�'1R�A�u�` �'� Q��A��';Hm��S�_ .���d#`s0��'Y�	�gL+��PeGB�n�Յȓc�z�{u"^�PXQ�M+:�I��Ug���	^8��ä��(dX���_��q���8+Z� ��
���I}�'JfX�v���|M�f�C_2uʈ{r�'��)1c���H���P�+H<�����ԸiM��ʒ�@� �,�q��8u��j�'�� Pd`�V_D���(g�����'D���T�˫}�x!e�Ez����'�zT�p���Ov��a���8���+��D*�'ED�!A�S/�8�a��ob�����r`h�F}@��� �K�x��=Qۓ]}n!7��1}8=���[<0�<���M�v��)��<��O�F��q�Lp~�'�0)*uiX�2v�q�"��72�E�
�����<������08���N-䀱���F�<Q�]7U3�q&�Z�B}��3�A�P���O5��g��b�4Y2��5k��1�'�h�c,A���� I,/:���'����.R�c:d���U�-�Z��'����ޮ* =��mG+5<2��	�'8]�+�"b�-!MT�� #�QD{������ťD�`ڡbW��
.� ��-#lO(�H>!v�˳��q��k��{��AL�<���ɑe��Ń�N�8{���AAH�<r'?P����gNQ�S0�9CB�E�<��@�,�v5�OJ%]y��Re��x�<� �Q���˸br��)�!`���@c"O��[/���|�Xe��A
Tm:�'��O���c%��v|XьD�����t"O��PU�>Xn��cӊ��y+��Z���O|��Z��� rU��lB�>nt��'~�����\&��c�U�(�¥c�'�T3a��(9��E�0�W�%DI(�Oң=E�TA��������64\�02ER�y�c� �ȭSD#Λ-�\�tBV5��4�S�O�&D�RfRE�������҄�/�O:�'2Xq��l�,i4�ajB	�5+۴�PxB���Q� �刻D���J�B�"�(O��=�O�YSL��T��6L��v�����>a/O2��$Q;q*�,����X�(;���7=�aR�OX�a�1>C�M�}q�`��"O(��c�>9�ڬA���Z���i�a|B���pƥP:D�:AS �#H�%�d'D����/.����[�MEȁ�U�(��A;�(O��x1S�kT�^κ)q�mH���"O�����UEP)R-ўnS�u��i���d�=�~���O���u����`�!�Di��	��Z�4$F!�FB��UH!�D��wn�Bċ�P-.�8���6u	!��F��(�5(�( 0��x�i�'g�!�$D�{���FS�K �=�ˑ�^n��*W�Q�"|�Gd�IN d�V���$��IW�<��g�}"�a�JJ���f�x�<A'���:}�\(��X�۠�H����i�)�=��'���s�g�$T�`Xp ��/Y��uz�'3�a��O�_�IY���V)"��'B�:P�'�Q+��7>b�����G��Q 	��?y�O��PG�2L�2H ��>x荣��94�TC��B�3:�*4j�	uz~���"LO���q��������֡e:DHi��c�hO?��@�	�l�Ib+R�2�z��៪�Q���剙jUN���]>ڌ�`�COy��C�I& ��9�M:��}2$,�;1y�C�ɭ|W ���<��q�1���B��,n&�KY�!��ؒ�#��B�I)=�ʽ��-ū0�����ݟc��B�Ɍ#�2\P��͕v@@�K����B�	$@;�oR>�,� �I_\�:C�	[�^13d">M{��
�(�<VC�	 J��Y�f	��E�0O͞j�B�I5��0��h ��(v����B�Is�9 a�-]h�T$ƇwTB�ɺM؍�S�[����B rB�
:���S�	�lߜ���ᔟ:�pB�	�;���̹,(��w뜴>�HB�	�$��$�6Þ�g,�yA��ABB�3ʨc�j^(,)�a�g��B�	�w1�ܓG�9�(MP�+F%f@PB�	�qq"�bV�=T���3q��B��<d�����ױ�4	�ɚ=-\B�I�oZ � �gʆK���  �1C�I�U$��B���$
�r��b�C�ɱlW�t�E���
�7/��P�2C�	%��q�W:T�2���
E�BB�I�o02��P.�o��e�( 0�B�!L6��2��
:2�hR����C�ɞPT,*֎�-��`!D�O�zC�Ɋ/���%��-m �0��W�B{^C�/" ��x"�-0�M� �LC�	�p�d��C�l�칡!�Q-`�TB�)� �	'"�����(�nPG���Y"O9��-�5�H��� �!�T��"O�(�׍K6h��Pd�^O��Ke"Oŀ1́�j���`�����W"OH���J]=�@ؚӡ2�x�"O�,b�˝qB�U`k�,iP"O�I1�g�+E���v@�3�H<q�"O��B��U8NO�A(���:2���"O��35H"}����ۛ-�r0��"O�г�N�8�Lə���%M�V�	�"ODTî۷]�^U����(�@1b"Ot �M�B����U�2d�@�"O��C�9�}F��}c ts�"O�q���(4�V�9p���nI45�u"O6��N��3.ؐr�Z�V� T�"O��w�od�e`˷0�:$"OL�WL��b�� 3���-rSR\�"Ot����;~LnTk�҂�x:"O\82�����KAb^;S�N�J#"O�ʤ���৬C�*�R]��"ONA�ƭ�������i];��"O4��&�G�pzU 3"�2+��#�"OVu�&fJ�|�A�#�ɴV�� ��"O�q���H�R���@!U*��"O6���d�S�n١×��j��"O�+��10�l���{ֶ"O (Qv	�.E���3�
� g�X�CR"O��i�%�!b�~��	�����"O�� @m_!ba�U�O=�PȒ"O��{�D =��6�]Tb�Y�"O��x0�B�cJ�8?OE@�y2"Ol�i�ͻ9~�dٕ�3)��e"O� H0`�N!r0��ܒ�`jE"O�4
RkA�*��U��;>��"Oά;��
��}s"M&�z9 "O��BEB�H놸��ރ�b �"Ox,�0N�<���D)���DR"O"���Țg�X�רŒ��`:�"O���W'�iܝY�fì��h�"OJs*	�b�R��ۀ0��=� "O��0O�:M�܉@#�w��}��"O�a�ƚ0&2�jcC�}�̽�W"OZt�M�#����b�ƾ�	�"O��*��	�i爁���>[(���"O�\*��:f
֥IЂH*@ı4"O ��E�w.Z�2��
*���f"O�P�󍈲bxTLs@b�R�ɇ"O$\�C�V�`����T�P($*1�"On��!�*Vl��s��6�8��U"O��!P�>�5ׯ�R�`���"Oa�A�k�zq�rm�.xvF݋�"OP�#A%I�?=F���[�g,�"O�-�l�
A��2��ۈKs`l�"Om�� � �`�����8ΠI�"O$8��	��6p�Zbl\�&Y쑰s"O��a��=-x��1kȌV2�� �"O,n ��x�cdϿ4���"O
�2��ӎ"�hA������R�"OD��刔�6/��a"m23�%�"O���VH���b4��G��Ƙ}cu"O����
fق HD���7���p"Of����$AOx	∎�x�"��r"O@uL�=rFB8��$.��3"O`�ˤ�05�Ԛ�f�>�,�g"O� �<��W5�"��M�9mV��"O:ܡ�̓"�!�E��͹�"Od�:��õ%)���p@��"O������)�: #	�*?�+b"O\�b��jB��
�S^!�@"O��k���3Ԛ��$���Sp�I�"O�;��KS��ŀ��W�L�&"O��c��B?g>V)�t�3t�>D��"O�()׿�����
^T�4�"O�}o�J��	+0M��xr�I�%D�����%E^x[���
��A�/D�ĺW��$xK�)�T��Ţ$8�!�D&.#L��H�Z���Y�@�(}�!���&��KGD�95�ȡ�ϊ�@!�I�k�zx�@%%���h�-�='!�$�k)Z��p-�r�tٳŭ��T�'�pѣ���[�SܧM�<:���F�MZ���?,~��x�ĨR� ���q�I}Dy�W@-���xNm�~&��ٱdU��i����KF�p��'d�-�Tmr�SⓎ$�P)C�
��!f�<��Ԁv����'�U�G��\r�'����Q��!{���J7i�cZ��S	o�I�b^���O��Ӥ�ָM�J�'���2RD��4n�XK����,%���
�'NZ��H�"I"�D�wk ?7z�EL��Z�J1�t����#cg�T�^Q�O��;ӣ��~�ᴎ��,��'�J����R8nx�P�'�$�Ӗ��s�2�I���9=ʮIK���:l���q}�m�V��|"��7m��)��ŌsMd�1�H����	���r��P�{Q?��
)�p�S��)� �Ӷ,>W��"�f�1ʁtX�H�4
H��Ç)��m��U�e�H���'�&���+�vbp��9y���)����H�	����H��æN ǡ�����h� ��X5�@Rc_�v�b���l
�P \��U#��g7�-
'���YϢ�S��*1���*!Yc�u�s�ܷ\|`-��ɪ>�t��vaO<p�p˓g�@	"ɞ�9�^��K H�A������O�L)�$g�g�ɳ%��� '�N$�lۓ�	!|��'�L����ɒA��	j���t�,Y���c'DTI����6P�ig����<V�'�؝�����q:���<k@]:@�ܛ"δ��j�yc�SC�4��5J�h4��gi}"��C]�[�*�9S���P����?�΋A���#��y��kEܠ,4�ӆZ<.�h�(�VR��B�ӿo���'�1�Ȕ;��ͣQi��8�+�G�
eYP�	�6�N�q2�U,3s���|���	@�Z�"��;7b�3֥�{MR�L>9�%Vm���$��,WJq���ޡ%�ڹ	�MT!W�I=�9����k���@ʁ�*��>m���5O��95+ڑ���#��6�T�T�?�O����ሖF�0�[�?!Cd��@�Z�M�|IM��$���#BD�~���'��	��3��CMR�k�%��|��h�S$	�r@��hd��AW���鍯���y��ȋC?]($�J���=���|pn}5fי"$��E�]�';��g病Thn�I��A8X~������j�i�j�^m�FjI=����"O��Kf`V�z��B����(��O� ��K7P�ӕ�	�5`�1 �)ҧ@"��S;H	j&BQ�:��ȓ/�d���e�}Y\�Y�I�(�r)��ˌd�aat*^@r������|R��\ͬ%k�@ݗ&� P�oQ/�p?Q��	(A@f�����:��$	�dؑ4Ԉ\X�)оn���#jLJ�	q3m����<٦��d�'�H�g�P�J�a_*,`Q��qR�� ������q��B�#�0���O3f6r�q��F`�B�~H<�΃9EI��C1F�M(��7�V?A�D\�2�8�i޽|���R�A\#!EԽ8�� �&A1ּy�̍ά� w$�7��x2�Xr�:M"�C�/�H�q���%j��iqg,%a~>��b�T�Jx�֊�s�>E2ַ����xb�2X���s���vp�s�,հ<�Ǌ�V��$��Y��j�pf�����`��͹~ViJ�@S���@AȊe�ҌYr:9;`-,Ov���Q3r� z"�Q����>��̖��1�GMqò8Jn�BH�hQAJ��x�� wlK�n�"|I�B�g|Z��*md��Ɠp& ����U����l̚"���X�`�3Z��IE��?l�ĠA�(�q"$����i���y��H�^��C�h�h,��"`ɂ�Pxr0	�ls��.�`H��' �,�s`	5��ʰ�i���B�=��k"�Fy���06�4�"�#̌����q��
�p<��k��6<r�2R����y2�-� ����Tb��R�A�l->x�G�*o�L�0�/�O@qH`�� f�� ��H�r�-`D�>I��`�8D;`hF)����R��0#O?�[6��C�,��ڇU����$D�бB��)hB!�gVh�"HXDg�.�&��)O�u��!��ܸ����c����o�����5�
��S~�aɁ�\�pΎtජ��2����e�o�)2�Lȇ�>i�f��'\�!4`ζsZ1�`E�hX���Ȁo�r�Q�T�r��N�&L�5ꛏg_FH�ō�<��W�n<�㞢|ڄ
 �+��1��AԲ4Ơq��@�k�5Ĥy�� �k>UYĆ��p y0$ʦ �v�	rD0�DȔOT��3�(O�u�s�
�N�ֈӤw*��c��'��q��A ^`e�P�� �8$��,߹Q���5@f<`��[A��vdC #ώE����x�'� ��$;jA>�|�1e*nK	|JQ��B�G�C䉥^�l�H�k�5;T��d#�I�<�ɒ]�䝹a�����S�O�XC'A4k�`��3Å E�6h�'�l囦��_]��B���en(qW�<���M�H���	�d=��"�7+�lۣ�E�-MT�U W�p?�ŧ�xд`!�nI�m�x +w�җg�X2ѡ�W�����y�byL�<<�Z�4F
K��EG}r���"�\��3鄞Ja�O�1����t9��$-0�	�'!B�Jv�H�^���#r@ܧ̈́�r�'�����8$�U��>E�t�^*܂�㞑�d�Z�BB
�y��K�H�y�qKG�]��鐏U�R�����Z?F��2ML�z�����(Of\h%�Ҋd���&��	DP;��5b�`T�=y`Bڳ@9:��u'\�5J!��ӰdS��0�dP��;�O6�륣S1s��4�#������ 3%�:]=0�̍���$�t�lLR��$Ι����ڛN���*��*[J�a�K�i��{�$��u����>OV� t�W�2,�\�$U�e����`�'�p7mN̂����Wv}r���7'�@��t�8n�#�f�/>�]�bj� &�O��b��+��-O�A��
!��� ^����t,f��sӤS8^�N�lp�OL�H�th	��pzP%0Ix؛ro#8g�$B��V# ^6�,O�!R�ݘO��1BA*Y�x$��#B�o��(ю�Bh����ƣx;!�DA�	B a�g��|"V�
���?_�0� ��4s�5�W�>�ߴ�M�ւ�9d�Hʓ�5v�ȉ(���I��\�K��)�v��;G����U�@߸�#�д�?Q���7/�f�b��X�[���K�<�"�+E+���*?}��T�\b?�k!7��A�g��b�
�A2�I[�@����.N��>��E-O�2�8�h%�H��bmcU`>}�
ԑ	- ����'�<m0��,�(����n�l)s$*�$��R�>A��>��.�(g�pHˤ)��&%(S��V�<�0��<U�-:Aʖ?�pDҶAVğ��eZ"�j���	Q�D��MU3���1�铻RE�C�	�@�t� �%�ArR`�/lˀC�	�}ň��V��>��t.�1_��B�I�.ZZ����ң^G�l"�+F�jB�I��(�Al�>������R��"B䉑'J.�A�l4�Z�����B�	���%*6�3����C�@�C��:�ڝ�E� ���y���>>z�C�	n 6H2c���kӋV�h��C�1C������I�<9hbђ�|C�I�\����B*:I��K�DO>OG"C�	�m�ؽ)���,8��82��
��B�Ir�6Q �dѐS�%y��^�Q��B�	��.Q �M�0��E��V&�TC䉙C1���
�(�b�B(KwBC��713�#',�
gr�2$ҨH5RC�.@����H˝\�\0sa)?/�B�ɩc�.�ð��$X�Vt�5jS4w
�B�	�-b�$��Nݒ��%�!�Y�C�b�4"�U�`p�}!N³r��C�I)����h�e����A�d��C䉕^�����IR4�� sDϔm�C�ɔ�vBk�����%�Փ	afC�)� ��1B���z��g��8�,�"O���9�T@qB�(�%�0"O��It�X+;�<�s!�\W��!7"OF I���$}r&�{��Dl~$�q"Op����t%�����KST&Dx"O�IA2�D�%!�#�V�1[�Yɐ"O��+�4�ָ�N��E6l`qR"ȎJ��Z-�����0H��HQ"OV@�ǓJ�0qcP�H">��B"O���O +�48��q�,��"O��j����(�fQ٧�ڽ?�|���"OJ�I�D��^�5���B�ǶX�!�D<��Y�E�'b6f�r�͂D�!�&_��`���J=�A��%�n�!�پRG�("��W�8�ndS�D�!�$X+3���P�ǃ/oKTb��Sq!�dP;�2E�8� ('�Y�B�!�Dս.��sK3L�Q!��/~!�Ēu]N��ǅRS(���<�!��76K��&���:��}h����-d!�D
9[�.p�ba
"%����g%�&j�!�䝐HdP����S�S�p)q�))<!�䑂.1��E/^'dǨD��ð/!򄌃9��p��*��1�B�qB��!�DH>=e"�jA�y\D���[(R�!�$_��� ��;{)XK�'8�!�D
�0mJYa!�?��T�34�!�$�a.����4E�`�,��+�!�N	4u��`5m�.E蚄�R�=7�!���X�L�S�)	�BAӕaR
�!�DT�>/xPZ4��.�h���F2O�!�Ċ$��E��:^�J�K�&
(�!�dЩSmXE`�����(�7�+~~!��O����"�����W`!���B�Ψ���̗M�&u�nĢ�!��l�2���J-U#��l� YrC��SNV�©�!+����KC$C�ɰ:��C��F�<
.����kB�C�	�X�qAr��*w9�<j�����C䉹#C���&/�?Z#j� �	\�q<C䉫`��a OM9W>^����ݿ��B�	�8%���'^�"�b.*G�B�Ɂg�6���'�!�08`��^[�NB�Ɋ�82�
��z�H��Kں��B�I#w�$}�g�R�v@����#bvB�	%P��p���E5�M��/W��C�	�e�T�3�V��0��]W�C�	�}�p��U� �m��F��qI�B�	/\��������{W���A�7u�B�	�h7x��`k�{t{�F��q�lB��_��Q	E��%0��AXQ���B�I!\?$%�tA�.n�`%�.��B�	1qm��^4���!$)-\�B䉝s� H���,U�IC"�0 �B�	�e���Y@h��dۦ!q`cD=v� B����e�I�6xy+b� NN�C�	:�|ݚ�N�9]�G^<��C䉖`�Ȱ��'Y�c�>I�e
��w��䆥5�T%�v�D.^��ey�˃�[�!�	���]���"G�L�F�K/$�!�$؜a�ʄ /�:gu���TEF!�D�W��8qC>���o�,H!�DB+�� %2Q����d/�"`K!��; x�����ۂg�@{Ԁ0!�� ^d�A�[��h���ñ)�z�$"OJȚ��_'U�E)�F;>܎��D"O����NEo�	h��2&��d`�"O�]�dI9��p*
H�.M��"Oj�����:l�x	��O��I�4"O�yz���=&�2��w��z�I�"O��j��
/��A5-�B�A!D��!��Ŋ�"�6�-���5D�D� 	̬$�桹 K@{�����5D�<�p莜��
��by�ѡ7D�A�DV)�F�K�&�m�.�z��4D�(�Pɜ&p��*w���iZ9�a4D�pȧ(�vq�l(�i�m��P�f0D��#!���i� 0	Ч�if
АQ!/D�$3����V�٣D���iSf�*D��X�'�	 �ش��� ;#�I�#�&D����H�+]D�����.3�݋��*D��:�N�4�X�X�MJ/Ð���n&D��2�M�NRph���3M,��t�8D�t�#/\����tl�0,Z���"�DF0-^���{��ԧUS�$m��&[��L�GD�?�y��_"K����$�,�j�+ׄM�+=�q%��;�$*���ēJ$B�8t��e^�УT�]?{Y%�Գt��>zqO�O%F䈣B\%98�0v��u�9�W�;-�I��#A�������>yz)�R��{sF��1'�>[�'rB��a��?��KЕ_�tĳ3��XCU��- �
 Ju�ܑk�ꥻ>�����Q�$I:��1d�e��� ��
T�r�d��B�q� ˜<Nt�`�>�B���
:���: ���Xg�U8��"c��=^�:������N�@�@�����7&�d�J\����'*Px�(�V�g�I�e�tCt	ƤR��i��d�l�'�4 ��$�"�@�D��l�v�(��U���P�A����<��@0gS�XvU�'�6T�B�kv���&P4��53 �$��� 6o��П�1�� �~d�I#�>Q2ǜq������5"V^��� [y(<�3���1�~Ԑ��'8h����w���{cjƏz��p��!�/R��w+[������� 逘���+�ܡ�KHb��xB�6�`�:ή��$&���)���V��"��*�\�1"��Z~Rj��W0vc?OL�w�ؔu�5����K�0�k�>a`(��}R�d����J��A��v�h�G.���Y���(O,�͇��>1�@A,o�@�shU�V
���v!Z9v�����7-B���I�@�~� �ܵ���@�!K��[��+&�P	`�n�š�$�*`�"�ʊ�=�C�m	��x9�b�/4���ɣ� �Fݘ��q(��)� 2BB3�V$h�ZMC��+x&��D�k�Bq#�l�*��d�c�8IA��!l�yf�?|5��3��
:>�u�<RS�E�¬
�~ɀU�&lP�|Δe��,ޑw�?%���0QȽ���?���[��G�AIޤ3�<�O
0B�$éE�u��B�^Ny��! H:��O2�E9�3}�m��)�>���"M-}ƈU�4����x"��F*�-���7�t���Ӳr���X�b�j�ʼ���.̨��m�d����M6���d��V
|`��<A�n�	G�.)H�ϐ"7s|`�K�a�<ɠ�a���Z���j�����C�j��T�ÁI5���� P0^�:5R#��`�1��"OZL�$!ٹ��ۤ$0���!�"O H�&�^�C�D� `�ڧ���B�"O�)�TH<c6�x`dƏ�_�����"O����Ĝ,(o�)FD:D��"O$��QC(G��:��34 քQ "O���BϹPVLyS���1"Ѐ��"O��y�&�!Y�<�`��K�8+,б�O��`�EЅ\�H���R[*4f�G] U��4�O��D��z�P`qIűf*��Y��'��pB�a�PT�'����e:K����lsơ�	�'!H���ɔw����eAuR	N��Q��
9�BlDI�Of�e�"�|1�ň���L�:��
��� 괈�̐;M�L�b��wW�����ω\���'��E�Gg�P�g�I&T�J1�jS�D�}���$u~B�*O�p@����8�ι{nО[8ne	�C�L��؃M{X�P�ub�%�<�q���]i�
$Ol�P�
i`��'�>Ⴥ\k���Cg��9�"�kA��\�<��!��}z�Ⱥ"�7Uu�E��^���l����B�>:"�0%�b<���@!҄e��\CF�T�<�w�ة)��C��[-�x�`�{}����[��x��z>q��'ق�䃔rS%����c�����'���TO�l���ۈ-u&�RF� "�䵺�-��\v���$ۓ	�`��Bҝp7,�kW+��8:ayD�%9�dL���Dy�L�$bf8�ϛ�%R	b%O@����?n�<@�{���CF��y"�K"_*y�ǩ�/��'^.q���D.�a��fяP�6���/
 $C�lI7�X7�ē J����1�p<%��3Kj	k�
Q�x�|}s‛w��<�T�MȪi�4�=j�4p��>���i�'M�!�ğ�#�l�bRǂ���X����5Q��2�*#<@�7��Ha*H��O�8:�҉)�^�Zo!�D��t���C��2h���E�ݽ>!��֟	�ؤ!��/��)ڧBYv�v�łd2��*���<0��=�ȓ/��j��6�ł���eH:��"Y�H�fK��PԂ=�@�~�?����/H@~xQ�N���H����O��ȋ��F)Y� �y��B�B~ⱘ�])`�
�H�C�$���	�3�e[%J�1&t�����@�>)cNѴS�\�qâ���'dԈ��c,&ɂ�iV)��F����QJ�A)�OV�".�9���V;���R�n�x"�N$��=C�S�"~J0)>�Y�`�m\rHr���w�<I�fHN���
�a�� Gvo�$V�
���0`��73,�g�'r4���Ǜ&x��8�n��`+�(��	�b-� ��B:~���h����P��$'d�n��G���a�܁f��L[��Z;R�C�Eӥ�ybM�5tΪ��'�j�kL��m�IK� j�Өo|���e�[��Q�`��ĝ�v��ɱ�p��iY�!k6d�R��| �����ݳcO��Yl� ���S�O���"��+�0ș�N�R܊5��T6!�Ve:�f�5�h��y���^j0*�M��bȬI��Y�����4G��Va�g��p	�Lئ�B󁞕:�� z"�	���$�Jl�d���7�Ҭ�gbA'u��-r�!
)%�F���7����h�#�x��6CWPmy���#
ڔ�Ud��M���)(E��"4�>)׭6C[@]BŔ!	 �OsZaS!)߫F��aP䃤K�& k�n�@���e���D�_d���r�B�0��e���'^�A��B�|�ئO?	�b,Fv���h�Z�Ψ(�m(�I>0 \Y#��#��>�z�NA�J���]�	x�c�(}��	�*F�'�}����)M.͙��Q7����/��F�Z�>��>���[?rU�tS��_6~.����]�<�qF�%�2Z�.�-��'�!��3$�4B�NVm�,����T�t���+ҭSVf̑��*D��2᪗���d�@N��@�x �6L&D��(���Q�0 � 3zj�I�'"D�BRˋaN���q D�&4H���)>D��	��Ϊ2�(	�J��.2(��:D�$�b�5GSYST��*y8�9 F�8D�<kE�˶E���D�ܺ2��i��6D��+eJ	&+������A.�Cp�3D�4��M��S~�����֤Z���O4D�ԛDI�B
d��$L���pb5D�0�tF�;qA %r�.�&*���� �$D��if#��"��RJ�`�h�X��7D�T�4΃������k��  2D��r&5ck*��ኁhZh��*3D��@�dZ�N"fYT ��u��(1,1D�X��ٽG����e]�x��$Z!�:D��kb�_2~��c/	�Lk�L'D��" �b��S���N�"$� �'D��cW�\�O�����	��.CJ\���$D�� ��k$�U��ᐣ)V�^Н3"O��qR�ފ�H`gIGd(H�"OH4�Kf�DD�
�b�Bt"O��C#IJ�0�s�ˆג��"O[Al�C��q���R>T��٠�"O�-��
�^��q��#l�4"O�:�Dϲz�j�������y��"O����أ�.�C�e�p�H�"OЅZ'�ɥnA��pѤGɌ}y�"O董e#r�9��AE�m�P���"O���ɐ�@V�q �+6����(�y���h��qIQ%	���y�ޘ�y�I�	�f)���%9��`�7�y��!BZ	��t�X遇�K?�yB-=$i4�)wc�a� pyb
��y2%W�(i��b��\(�|�Q�Γ�y�ɛ~�Q��쌙T�� ��b���y�NΣc5>��V$�In�4
BAվ�yBφ�J��@�&ĠO��X)�����$A��<Śr�D�6RO��dd���m����
&����F�Obl+��NNW2̀M��}r�O %�8h�gh��bT�"co�^�c��b>��J�#�ԠB����7�@Y�[~�I��HO>� ތX���I32s��ʥAk�Ȁ���ӷ��})fkH|]֘���0�\6m�x?��E�i~"R��?�AL#���!��^�K$>5��g�"�a� �����b�"~nZ`���f�U$��Y���N7u����Lyr]���v�O_R� ��5*͚�O�(8٦���)��%���vŬx �kUB^�p��"O�x�`�9kf��O�7s�2�:"O��Q).DU��i�[5o��@e"O��։�,b7�HS��!I�(��"O
h��e��V�D aa`ՙ@%�!�"O���p#�4X.�Y���j*��9�"Ol��7�#�L�reՁn����wQ�E{��)ьK>�Q�va�/Z�bP��B�7$�f��47$ɸ��=}"�1����!�sM6`�i�
���Ɇ-n��ӦU��0|b�EG8}��e��+�/:��ȱ��]}r-\ ~���f�M��S_�0AhQ��.FT�k��Q!:Ӿ6�[�,h���?�E���^���M�Fnδ���58�Xdn�5#��'������"�T�&%k����G��-�})rnEn~B�\ �?�'jS�%��H\l�S)(@����`00a6*�5�Ȑ�Ā�-�t#Ð�?���,�,j�l�9b��h҂�Q�{Up0���R τ�+v�柠�G%G]La��᎘e�Vm�d�v�Mh$�QVM5�O�ŋ1%�8i�@�qnɛ*cx���"OV8@��X!tuj�Z%y��YV"O���p��[p���h�"OHc��'`�\����@	#wda��"O��i�"�u�4DjUϑ�Xqt��7"O��Y���J��z�")q��D"O8m�G�ȟ[��R҉ڃ7r�1
�"Ot�Jv,U�d� 1k�)Nir���"O�铕H6w�уH�1fT嘥"O��0� ��H�����&Y�/]z$�c"O�@[�H�{; �q��>5EN�@"O�Y��k�?D$p���nW>��I��"O�1Z�+c���F#O�X��0"OVH�
�>�,`�j Z�f�w"Od�����e��'Ы@԰�hF"O�24A�(.� �+�Ʉr�(��"O��R�Y�
5H�N;%��ҥ"Oށ��K*U�N,;���F���z2"O��*�)'��yD����JtK5"O"H1"����P�«���"O|=bԥut�*G�Z&]H�Q8�"O� �h��MVX%Ɓj��Q�N@n�C"O$��A��l|��9Cl7H/P��b"OԄ�))F������,<��4�"O��Pi����y��K�(���"O�]x��La�2@���,k ��"O<ySa@����RmC/F⸱@"O�`��U�"���k��#p��c�"Ox�G��0W>��*����XW,A�E"O�̃�D_�,["�;-/w��!�"O�u��N�%Ʃ�&7Z��T"OX02u�]>h�tYŋ��]y%"O,����J*��U��
ʮ.� ��4"O؃�ܵo�����#Ũ-"Z�z�"O"���c�; 1�`#.Z3��"O�I�a �%/B��XG"��)7  Y�"O:��S�_=a�l3��:8P]��*OR0��ƙ�)M(�j�$��Xڬ���'�.����	�+V�E8P_�J�H��'�b��WG	/�PQ�B��>k<���'�}p7:����Y�p*�j
�'��#�Q-T̺l��E�tf�i
�'�u��
�6,�~I�@��
q:t��ȓ73�2ŬY�a��E�FA�tȄq��x[��N��r�D���J�K���ȓ#⦍�B�\ks<�1�h�:��͇ȓt.���p#H=�D!���ȓ��i��% w��p`�U"y�p���>�e�v���`.^0� ��)!.��ȓp�x�穇?
��d�X;�d����1�I�6�wʕ�yA����!FJ����4}�*|P�(J3 )��N���@oM'=�� H��E/G�l�ȓ&��r@J��SE*�ȸ��m���(ք�< �����J�L�1���X%��J�!g��ћs@�Z��L��V����': � �����3��p��v��eg �*��E{gg�M�$��ȓ@�., ̅F�Q*���)��5�ȓCP -S�I,FX�x�c��!�� ��L�T�x���D*&�R�͊}� ��6��S���h���m��J,|�ȓ&�Z\qR*�<������!coX�ȓU(�-�S����xuġ`bh�ȓX턐`���"|���㊙r�H5�ȓ2.�h�BK�9BD��b=1 蹆�8��<JV"��5�J�P��Э`	$��ȓ2Јj�!�� Fa�ȓ3��1��	��,a��	0�p���"�PQ#S�Y��R��aB[s�a�ȓ[5�+e㞮*�����*��.�B��ȓ����J/)7f5�'�øW��ȓ��C0����0���1]��p�ȓE*Hpș8R|�(7�H�o����ȓ&Uޙ1W���%�Ա�&Y�Q�
�ȓx��XC�'M<MJ-z���4V�=��V���@o���q+�I�/H.l��LØ��W��p���hʖX�ȓ<�̀�A�A�
����w��>!�ņȓ@�j�A��w�����a��;�.I�ȓ*{R�S��ȕ}8b�i�4n���ȓQ�:� ��nܾ �-4^D���cb��Q��JP�s3�ڸm(��ȓt&.y�ł�_��5�� �*E���p�J����
�CH�#��F$!��l��S�? ��4ht_<�Rn�~,���"OLqp7�J?^�ڝ�K߶,�j);""OV��Sgӓkך���B.�pU 5"OD�"b�(�V�1e�L��b�³"OHҦ�T�>� U�'�Ȩ{�n``"O(����X �,x�t/ēr��8�f"O��{�<>��m^ t���"Ov�pg�b��S1���Ѝ��"OĘ���/
6���L�K"��1F"OlA�Ç��6A�ҧ,
2���"O"��2䊄N��$����9��aK"O����$��a��!�cK�m|��8�"O����$mp�	�C�[|աC"Ot����Qn\e�fb��2�H��&"OL`�Q�<s���� F�@�"A"O�B&�"�f����v���"On�*�f�%N�t�Y�	P(����7"O<�E�D$k�\���ۨ[����"O��5�^�',~$r��.�J�xD"O|K�k3ZV���T�y�pE�4"O��u _�HA%#?9p�y8T"O\�`d�Їv�H@���/	B%��"O�D���6Z�Rʷ�˝GQp���"O<���ⅻZ�hB�L8���"O��0|8�9��C�#�8 "OH�ɗN��M��AX���d�S�"Ođ U�E:p=�}�7b��d�d��"O��I�l��W֬a�D��:PI`�"O����A�o~*,s@��4�m��"O@Xy��
�
������G"Or��q�E&C�� ������)#�"O���si�>(���/�P�Z���"O���2*��΀���3]����"O`�Ʃ�h� (��h�_e���B"O�����$l����(U�ZZr�zP"O"�۶dKg0�h�F�Uj���"ObE�!-	�'��X�aƀL7��I�"Odp�fI�{Vp=��䌮1D$�"O�K�/]8^ib�P�S
sX`"Ob�p���Gѐiv��\�h3"O�dy�)Q�D�b��DI'q��ѐt"Oa#S��uW,c�/̷���w"O�=�'^au��.�c�(�"O���"#�=�����B�d�Y2�"OX#"�S�l�t��v�]��a�"O�<��B��s�`X4��3X�]i&"O���q.�6�+%@ԜK�{"O�L"� ��#�V	�p��%W�Ő$"O�Dp�F�3ٖ(0�N�� )Ԑ��"O ����MQ\��cl$����"O�D��E��"}�M���<n-H��"O��H�c�4���� A�3p!3�"O�O��b�&0h0���Ɛٲ"O�	xtjLw�v�P5�ۃv�*p��"O�Ě��UR�-��NXK�pU��"O�D��+X���RM.�qp"O 92L��|s®�1OȠȑ"Oh(x �_%H��Ҏ�)�"OE#�/�*��u��#�6�@�"O��["�(
�sSHm��3"O�}�%�^r���g A���p5"O���ҧs��w��R�4��5"O:q��49�@uh�l:K"F�)�"O¬JV�V-�щ������R"O� �uyU�בJ�РWKZ&#><��"O���B+O�L@�  ��Su"O �B �#UJD����=x��Y�"O�yGڭ!2LPӥ� 44^���"O� �s/G�yO��"7 C""0@#"O��k6�
���|�­��->���"Oy��l�=n�氻�,a�U9�"O:�X��@����`�ĉ�"O��YA�8����y��"OְJ�(��5��p�@?N����p"O�zS�G,w�fR��F0p�D��"OtM�Ah��TԘ��Kq@�R�"O>�0��N���3���o��P��"O,,)�bJ<a.�� ��G�6�H"OhL�!�p{J���΄�o��!"O2A�roV9�\:��0b"O�l���Y@ܩ����Q�]�W"Ob@(W"+/�1U

�o��[�"Ovm�dA�f5���X&Y�"Oܢ�#H.8�6!q��δ��!�0"O�T�u
����v� �y��"O&d�3 �?�y91Cҳ��!J`"O����d�l� �BM4wɤ|��"ObQ
��D�0��u(U�@M��"O��� GLЎ��DX�Gʲ�9d"O6)�bd X=Ti����#~-AB"O��a�c17��h	�R�5
�D#U"O���7+	�&��Ğ�9�4$1"O0x􀑃$LX '���.��\)�"OV [RfZ(n�*��!^�$�$,1e"OND����`	���ŶP-����"O��s��w\�`�V���`#��A�"Ol8�T��1<R���Չ=,Xa"O��k�ʐ{L��&�H�G^DI�"O�%�V�D�1���+!�X[�|��"O�#��7d`��I�舺,ꢸ�p"O���mԉ>��0D��e�֡)"Oh��~����G�;Er��"O\�����PK�Lb��Y(2U�"O:��1�6{�� Q�cﺄ�q"O���"d��r����~~�2"O��ӣk�ŀ�$$Q!W8Dږ"Oj��S��-����M)x�
�2"Ofɲgd�5F�\M
W��d�(�1�"Od�'fQ�B�lӷD�<z'
I��"O���� bH&ȳ�CU�ij�x� "O�݃�,SB?^Q��b�)b��c"OV�;'   �P   �
  �  F  �!  �)  V2  �8  �>  8E  |K  NS  �Y  `  Hf  �l  �r  y  Q  `�   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl�lT+�:O$���'h4�l�r������UBJ���ާH_.`�ס�4b����Ì\U�H�"�CmݽrB̀�?�4��?u	�O�����
���U��e�qUJ%��GV����K�e9�#6f��u��ܠu��$�'�8��RG�C��!�\k��G�#7Vz`K�O�4:B	F��͉�঵0��]˟��	�D��ٟ�� ���v��iE��]0ei�eL��T���(;�T�ݴ��$�O�`i���>���O��C'C˨K�4tA%�!��iiì�Op�$�O����O�D�OꉺҮ~�X����<�G�R�e;�ڄK|�K�d
D�'R�V z�TC��Q*�1xEB�S �)jC�>��䣟�$�2���1�0���
R>w.��`�&�,(����Op�D�O@��OV���O�ʧ�yWǪS�!�͵c��C+��?9f�iD~6�L��! �O�)mZ�l�%��4X�0��}M�t��KĆrNN��!/��8|Q��Ɋ>P8M�5�|�Q?���!d��g΂�[(:�P $N�N�8�	v�Ay����̦�x�4bq��Ou��+W!�H���O�N,��{���Pcڙ7��6��r8���`
$��c�fV'�ؕI��M�,V�lZ	�M[e�i8Fݒ�l@���[��@�!&���0cC�9�vM��#]:%E6��צ��شkf�a�W���و1 ��	�@�y��ܢx�P�+\I���۴i�T�y�e��������i&�7m����e��9)�^�Heǘ�&Ц]q`Ϋ+������<���%Q/|���ڴu%��#�"W�`��%ʡ��A*9c���'��K��#����%��Q"�P��'l�O����O$H�������O�ll���ÖR��V��M�0%C��?I.On���Ol��;.�����J:wv���s�O�e���XQ�t��_z�@)�b$O�D�E�!5��
J]�"P����\~nP���l�|�j�Ɨ�5Bax2��%�?9�q��I�f�H�3�*Y&��cV��n��O��d;�)���<����F����&T(^� ����Ys��hO�I���I��+d�⵱��ۤ�j1�E�b	o�I�������b�O�h2���V50�it�F	PW�"O���ӮµlrHAt�Xk��1� "O�v�sD`١�*���J7"O.�0�	Ъ`��;rc"/����v"O`��¤�"@� �C���ZȊ]`�"O|�sA$ĀV����aCW(�v���'�����O��p�)L��{5��Q94	�����ҥ\ӂW(Q6��)�:D��3t&�5s{����aO=���g�9D�у^1�8�7�òB�f1�q�<D�tr���?l� ��!�F�b�I���/4�,[ġV�~�ٲ�Fw�\Tr6��)�����O����O��$����$�O|�Dτs����P�Ɇ{Q�@��$��BO�64%D����B�|���I�I��8@AC�*@T�`H)ZN���)\#y�����^ B\�&�݅l�AD{b�H!1�E�]�RZ�P�Z�q̖���T��#(ғ��>?� ���� P��[�62RȫQ��؟���R�(�S�i�Z�`$��/�L��	�M{�'���j�j�'P�$��7�iK��'�LJ爌,U��1����>��;��'� L�Y�2�'}�膶bs(T�Wj�9V��B������*N28�,��&m� ��ɸ��]��P�H/Z�ք�iK�+\(v! K~N���X9<���	ӭ�7`nl��wAY)^Q�|���O>�mڳ�M���f������cV���+����WNy��'�OQ>1� �#���xf�?��8��i$ړ�hO��m.B����]'�vى����%m�1�4��K����'E��'���,IV8��D)j %�e$W<�!���6wҙCq"�L2�ma�ױv�!�ޖTdhL�R��19����+P�%!��p	�@
/0/���R*ժ)!��#a��0&��CI�T���ظx�!�D�@U��A���%J?�pa��L_�7m*���J�(�	�O����O�˓*�"�Ei��[�]�d�C�a��an\�o�f1)��L*� ��@E���I nH�����i;ν��π/.HH�Ǉ�f+�)-�^��g�79�c>q��MK�d�2Q��$��@Q���47Muy"Ȉ��?a�����?y�9���+�C;=P�r�4W� �K�]�OHu�&KA&���մa�t�#v�'��m}Ӽ�ne�i>��ky���o���Q^�I�}ʥ��,)
^�7m�On�D�Op���is>��"��=�J�;���|g��B��Lm�\�Oj��x�)Ag��T�rH�>� @������E����O'���P�M<X����C���x�KC�e�4+B��
�B�0�A-LT�e����?���i�Y�p�	��_��P���UO��w���+n���"�:�ӆV>`uӃ�
6T�*�sb�_�r�H�O�e�bI����'��A�&N{ݽ��ڟ�+s���P����.�M��]�c���h��B���Ɵ��	�y����sU���{�? ~UJbN��	J�b$EәF�4�b�'��E�mX���k��RL���Z,G�>Ճ��uTH��A��0<�ǩ�ߟ@��4i�ɔo�e�L���`܋UE��:��?I	ߓH
��P���:��5�C.J9X�!����?�)OL�=ͧ1�ҏB�N�(���5��z7���?Y(O�EĎD��!�	������?=Y�M��D2U���E��᱁��1Y�pi{6�ޟ,���2x��.�(��D�O�ʧ��I�I��Pe�Mc��{��1B��)�,�`�H�q�D�xb��XՑ>��A�)+��e["��x�n٩�'?٦Dӟ��	6�Mk������a ��ܹD�ذY���'�|��'�ў��'1Tq�g�F)
����H����'k�±>�+O��S 8�\qq� � �"���Y�+��mZޟ�'�"���O~��'�rY��W+�Z@t!�L^V���ˢ�	a��\�����<��Z��|�<�&��=����d&e�x$�ć�yj�M����<���˛z\f��|�<�B��Y0D˕�@� �N �&��M;���?�6$щ�?a����D�O����O��q#N�}{Tq��.Z�*��+5�%D�TJ��Վ0�2�H%�D?xߠ���-�<1��I��M3���i��p� 4+���xv��?g`d�WM��{7���O���O����?)�����R.3>�}ɶ���� ��4DjX�8�'y6���K�9˜��1�ۦr�,D�D7�x�$K�:U"Y�qߠ\�x�z����6I����P,
GR$c��I�(xd��'����cfC�R��R�MV��4�M>�`�i,�'�,���d�L��OvHS�JV='a����m�K���a#��OD�d��%ٰ�$�O~瓬�$+�	^Y$U:��u��Q�P�5!���D�FB�h"1hGQ��{ ��.~g��E�8O�����'�P�O�u�c&D���X
Y*H�"O�]!I��(��h7������'V:��,e�|l1׉޳|�%�6D�C��'24D �dsӒ��O�˧1(B��h��(���UlB	Z�I.!*8Y���?ٵ��?�y*��>d�	�E�FT�%��$X�u�ظ�'��j���SҸ��͕A��a�ſ7b���
�I)��S�OF(�Ai�')6�Y�K�P~y��'`�0iQ��pK^UrW�˘wc��C��D�^�Oi�TJ�B	��h��&˓Z��i��'�r��U�<�T�':B�'�B;�xy��Ŏ6��k��qJ�laa�q��'�,�D�G�%��3ʓ���2j7V�2�O�}|��b��	�O�,P�@�0�3��&B,�q��t�d-�6��0��Xmڸ�M��\
��x��6W���I��upe�S�j�^��6)R,{�qZ���ן�R�Z\������DYV)Pf��79�(3C��u��')����$�O��	�O �,�B�1��p���J��K�켡#EݚI0�����?���?�%����d�O�����B�m�ë�$6��+ϭ~z=¤�/��QJ���;�8d#��8{Z��1�I/���/^ ���)�;AhZ���k��8��ݸ���9��jg�U��*7M\&,�0*�}�)K�N�i�FE:8�����w�����?a��i��^�P��s��M�Dq�DӸe�ʥ*"�E	s�XA!)O������,�i:�@�kת�� �V9l�'1���P�t��#N�`K1����a�t�i#��̐U�L25U4q���O˓�?���?��MK�U$ik�N�1!��'j��k�1|b�Q# ��1���>Jy�) �>��2f	,5
�VŐ��5`�%:&���G-ǐ�0<���A🠣ܴ�?	����Eb$�7����I�!������?i��?����И',�y��a�6j,k4-"���y���i>A��R��hSGM�S>�b������Iiyr���M>6-'��p>yl�͟�@�H-0�J�9'ћwָ�p�-�ȟT�ɞe�!Pd����8!b������gݎ4���O&"R)�a��?���~d�<S!�W�Iz�`�"Ko�O��峴�-#ƀ�2!�#"$���O�+��'�@6�Q��A��U�O"�h1�D�xih��J�Q]��O>����?���ԟ��S�b��2��YҠ:���C��	��T#�4Ae��|B_�?��ZG]�a0�oT�	~���
>Zy�?�g�'�h`p_�<AlxAPO�1�ZP��'��y�c�eJH�h�+:9�L��'Ș���xv �fˍ=/&p�
�'����/�!`���%%�p}��D&D�4ku'Y4et�+�B�j \��&"D��C�e/M����ԁ�3��I��ˡ<@a�x8�u�A*yB�Y&&��`2|�+f�;D�� r��!j�!ɚɉ&���DWx}�"OX�*�d��,�4�� /=�>�h�"O�D�pC	?=�@`���S�=�<�2"OL,(��g`����Ɣ�1�B��'N���'�&E�կ�t����7X����'� C�`�J��A%� ���
�'_�h���1v�X< �^�(�3
�'��Pۀ�Q�lX!�tl�#��a��'�!Zw�<F"���d;	���2�'78��4��t�8�	3-��4z���1�Q?	�,��k�`��`�?EDF�A�8D��!3i��>P4�������q�,D��ɀ��;:QH�˔�h�9���>D���$�L�j�ĘyD@Qg�R֫/D�<��Ӡkɐ\����$��`di,D�0��
!}d�
��1Utr$��`�OT�)��)�*�6�F&��lD� po������	�'����%Ўoڄ$�dG�X 	�'3����Ο��yjt+�x	���	�'��i��f�D����ushՓ�'�r@ʒ��C��prD��r� ��'����
���b#�̪b�L 
/O��ɕ�'�jAc���7^T.Hٵ�E�W����'rUX�ň5 ���o�VM.�'?t`���I7^ r5H�3=R��'FD����93���c��/�A��'�=lhl7 ��c�X�a���>���l?��G��~�$�Q�`��w xe�q��@�<�U㚂i��vmۦ���J	sH!�$� ���2��	��h��@ƲB4!��$#�`���oԎI��Eb�/L�w���2-�����%'<�n<���T��y�S 	b�)�;��=��@K�hO"�;����0��R�'Q,��!�E�y
�B䉜���H'�-j����#�<C��3��m��e
2]d:���/�=� C䉯�ε(���5o`hO	��B��SvI�T�W$nOP�y�Z�<��B�I1th�Cm�%4.Ze`�� e)��d	N+�"~��Kήs�!�Z�?ۨ������yR� Hl�sWaJ>>i4"$�w�<y�E�;_V���ؘ%��I���T�<!ҭվ�:|��ȼnM��f�TJ�<�B@�68aʉ�-�#���Z�)�m�<!�,�K{<))���|x�H�'�DyRK���p>J�!b�����&�xy�'�C�<�Eh��?��i�ÄYG)Q��@�<9�)� � �{Հ�Q@6�!SR�<aa�לL��%{r$KX�J���OP�<�T��N���0��@���|=�}"H��~�P�i�|Y��A�����`l�y��ķ;ư՘C�I�A����y� ߞp��+��{�X�٧E��y�V?D/�xѡÖn���W犚�y"C�4V��Q���m� �	���
ѳ��N�8�����n��G{�#����r}Zd�j ��3�N2]�T8��"O����Q�-w�P�Q+ߡI�@��"O��q!�9S��!�]�$�hJ�"Oj�H��^{	r4��+�\E��"O�������}���Ӽ�9�D"O𵹤̀�Vk�Qb���EA5�'%�%����6>��l:sL���RTs(
�g�9��^��{v#k���&E�ov����S�? �����]�}9�IR�@�U�ډ��"O>!Q��Ba}�O	�~�A�"O2es3G��YW�y!���d��"Onr�G�7W��1��C�|��;�X�HP�+7�O�(zq	\+T���� �^36]�Ɂ�"O¼��E��T��@��.�HE"O$����5T���]����雁37!�ɳI�(�`�e_7c�9+�*�-!�d�:k���k��_�zt h#©Ǫr�}2F�~�)EZ.�Ц�N�\���1�y����c��Lϋ�} �T�yBoD	kqbh��ʐ�i��d�*�y"镂K�2�b'�֗z�� uB� �y�ٽ�zM���R?z'�]�t-��y����9�l�!0@�q���"���'�hO����S*,��"N��~)���S̣;AB䉌YD��+s�]��Ɉa�C�ɥ`������Wp��{�n=C䉱X�Y�ao�lj���眶)�C�������?�dQ3ƣܠ,etC�0>�`�JB�w�T�C��[�M���$ީ&^�"~r@O�Q&�UX&N#M�H�Q��8�y���"+D�D0K/�:A����ym t8��J��CG�LȒ'kJ��yb,�g���l�#�JѺ�C��y2dČ$�с��>S^`�"���y���24_>�h3������b%����D/Mq�|��ԭJ��A�ÂնM6.-�g��y�E�@^��w�V�C��`����yb!��0��y����H��K��.�C��WC̹��bHq��J��
;lE�C�əm�Y��φ
A�<�L�j�����6��Q�f.@��ހYGB�3NN0aP!�D�f>��wS,d ���Ĳ;!�D
��0���P�ɫ��2d !��	8el�"f#�#�
U��NE8J!�_+c%x|���S��8�@P���!����"a���6��({�\�c�)�{�ў��N7�'Ua��4BڮR@NH8Q�#S�֐��T�Q�)'���+��6}5����U�Y�"f�=.����!ׯS�Ԩ�ȓE�y�dʁ�uQ�� �k+(`>l�ȓTg�p�����-�ҸP�H,\@��ȓSH���bO�t6lا�0_�z��I Q�#<E���՘?%ܜ{�ꌄQa���
W6�!�d�MM�y����, @L��NXG$!�d��qxnX
0h{E�h�dֺ	�d%��N* E��*�@*���U7wD�ȇ������@@�@�Bʑ�Z2^���ȓ6�.��R)2ڼm D"�2p�!�'[6�	�B�:�j�NS��d��&�,O����ȓq�"��& ��-q���&�ņȓ:���w�^�o�J1���Y"��ȓ?=&�I�Ь��-җ)�2,��*��H`4�ѩR�@T�ˈ.pH(��	7Q���	<=$()i�.�� aX��F%F�
C䉭<@F���,��H�`	B=QG�B�	�c��p�d�?��0��@� {&�B�A�r� đ$�T!��ӽc��B�x��)P����C�6��cmƅ<\C�a \�2I��7��̣t��@�=�ҭ��O2]�&���x��� ��z	�'>FC�#�L��a����zC�	�'�T V�E�C��(f �y�\����� �u Ч�"q��t�'a���$�d"O���q+O���*�IS9���Hc"O@���A÷(At�83�B9>�Y��'�ʁp���k�`���5���!T��'�2U�ȓy3����SR���� ǋ0�l�� ��H�1-$zU���ˬ6

ͅ����1�
�V@Z쐄�'��e��vd�����E5� � 'ʚ��ȓ$�A�Ӓb�|�ht!��I0���'�t(�YuĤI�� 4n�AY!n����@�ȓ`@��aQ�c3V@�j�7K�l��b�pY15&ÿZwR�CR�5�B�t�,U	� è" ^�#F@�?]�>B��5)熌Y��%r�Q��֑X�.��$	.'�D2sX�	Ck٥~I��:�i�L!��0ꪉ�D�H��i��I��!�Z5�H���`�>,2.���H��!��јoE����(*"�â�M�w�!�D��N�����N���EҽQ�!�N�4Y��5.V=��J�S�ўHy��2�F� ��\��4�3a!S=gi���C�j�Q�M 1~�ѨEn82ϸ=��`o�,z�)ʧzd
�P�E�hQD�ȓ*� ���͊N�Vtx��xR��ȓ/Y8��e���jҐ̈́�-�>Ɇ�"��1!����2��!�ʡ�ɒo�,#<E�D�ľj+������H'r��ő�j{!�dKQ�u;��C�/ļم�̩<`!��7oWh�%\ E�Bb�cB�<E!�䋆e�}ۖj��8���Qb�p7!�$	r>I1�C1�����܇}*��D�@x����3(︨yV�A�,<�Sh��?��A����oZ�8��0i� 꺻�m�����ߩ�!�&WR\��Хy�(�������@�������{�o�=�^����O�����?(��nҚc(��+��-�[�ǍT��#0K�>V���!�|�"[���?�������;�X���$Ӯ��`���HO�A���?q��D�J�O<�9�4iX�.��v�����3�O���U����}���=��,�'hp�UK�H8Ƌ�/tmฺba!j�"�'��4���'zVPq��'�v��U�ҟ��D.�<��aQ�*M��|T�b��ӟ�S��Q�RŒ����
���S���	2,����,Ӛ.Q���

��V+��80&�N4���:�'�(�c����k>����ܤG��iΓ%��������'���D�'�`5��ת2�<��n�at!�$X�%�	���3�(mBcA�`�ў�����7]jQ��͇?�N�`PJ�3D|$�'j�OX��>��ç�z���O��D��c��Vݮ�a�n;>�a� mź���qK�4�D`�p��=��,�����	Yx�eȔ[�
�9H8u�c]� bd�A�2�ةh��	ؐ)9!�G�$�$������:&�
��Ji�fĎk���\��ß$D{�1O}�$�B�>Z ��FT:K�[�"O��F/� ����_Ո�2��'�"=ͧ�?�y�e�����;P&�=4MR�b�1�?��A���Q�9>�4yj�m:t��?D��rDZ�BW�#�H] ��ȋ҂>D��@օ׷@8�����[4[wr$Y`�<D���'�XA�X0@@�9�P�Aԫ9D�ԛ��ںGp��&�7�j��TG:|O �Hv�>�%ߦk�YA ��6�5�%_o�<ɢC�+j�P����t
���@h�<�*�=U��a���T(�*���9�'�t��
L)m߰�ptF��/S����'�-`&/I6=\�zb�ԇ:p���'<�@�SM�H�b��38�p�S�����O�'I���)B���-�(��h	B&����n�:���c>5&r�Y4Y�0��T��^�Q���R�w� 5)��R�<� �@�D^+;Z�i��I�c8��  "O�AhG�,Q2l��cW�h4���"O�x���2x�����")f�R$-U��OZ�}�����Jր:����,?	�хȓ
v���Q��f)��:�h��+�4m��Ӌb_ �@�# r��$�����q'�7E�d�5��k����ȓ/��A��,�]����H�ȍ�ȓ<�i��L)E�$�"$G�;Q�I)`�>��$�E�0�U
S�<�&Aʧ焧g�!��$��E�~������^�B!�䚚!:����ǲU�\���J�:�!򄓛��`2�a��` ���S�!���P�d�;�i=l�6����<�џ#�Iey�'��Ƀ=6�L��� 2�z��ڱjf"�W9l�"�'�b�I&+�-�,�/WB�{'�V*Zv�`�;Ƣ�J�$	4p�l�Tgݝ��E|�$U	m�L��e�<8�2,�E��8sR�P���p�-H� �x2�+b�	-�"=y��O>��,�Ӂ[��t"1'����q�����V��0?)F�L�8PH���y��E��Gx��*OBԸ�P�k���� �IcKP��_���I͟h�����O6�T�@J���1�D많@!W� ��i�'e��}�e�I�|�R��A�W1���/�d���M�K<Y��/�ɜ�r<�����V8K���kc�Չ]� An�՟�
w	F�<q���۟����?����<�t��>�r�� D�6�T��mߚ	Q�t�۴�?i�F�.�?Q�'r����M�;io�s����y�j�o��p�3��InZ���?�����y��:�d�O\���O&�0�ũ��*�|��0��yf@l�sa�Z��'�%RW�'��3*o���u�I�~�V��~��*t!�"�V�ISʗן�wi�O��7�xy�O�r�'���'V�x�aI+&�޸s���\"]Q���O��j��'�r$җ3�1OԜ{fӟ�^wW��݀Cx@�#R)��7q�9@�M�
6-o�L��f�O4��]���ӟ��	�?�ᅕC۬)�7F�+k訸�%U�,�~h�L��ş$PZwH�4O����bퟢ6m�!,�֘3��V���R�lk�4�r/�O��I�)����OԈ[֔?U�Iן�1�A�tވ�(ݰ@�R�K&����Mˠn��yb(ъs���r��	�O����&%��$�;05�iL>����Ȝ!VZ��m� ����ry��'����O:� �oOR}�qb�Xy�!�"O�`��g��� ���xl�H��i�B�'P2�'��'�2�'�s����I(U�ҩ��%����׋j�>���O��D�O����O���O
��O(�kQBټi�%av&_� 5k�����'r_����z�_�D���1Y��c�G��+OP��M����s�n���`�?�����5*0�Ը2\����ɿN���M\7���EH�0B�/lHta�+Њ5Xݣ�cÅf"\C�	
X�xE	�C'%Q>m1"�9?4C�I4ez ���RQ'�Z'j[C�I:fI�����@ܙ�HFmC�I�~�^@��a�) ��5��hӶG�C��h�^��p�^6Ĝ� 'S�B�����R!؏B�v�Ip� C�㟸9�G,���q##F��Zl��!��1����"OB��� Ѫ���A_4o�bL:��d�����9厛�lp�2KIt�;A��]�I(ǒ�b�:h2%4y��cԁ��d])��+ �(O�3�O�'pq����V��)�#*E�L,�W���P5ԉ��j�6/��mKt(���JÎ��=SBO^�J��%��M����jso�.��zR2���O�H�!�ױm�(M�(\�2�v�C��Ib8�x�UAƩ4.yS6�P�A&���Q6D�h��L%?j� �M�&��E!g�)D�<r�-أ�P��N0U�$�I"�4D�D��	�/j�Z�K��X�{�3D��	mٛAK|�����#���+��$D���q�ƫ]8$�D.�6S���V�#D�h�tG�+��c���/����2�&D��{���!�P����XJLc��8D�#���;"���]�>�4���4D���HN��(�s�P�/�`���1D�<��hC�,V���7��S�<-S�:D�`����% 앁� ,�p,���7D�� ������hщ��>=���[�"Ot��b�/�tL��+��z��B"Oܤ�tk��c�hA��
gdT�r!"O��K�*-�D4J�h�tQ>��"O���"74�٩'��gJp�Ja"Ot$
����n�ܔ(b�7T��P"O�MPr�+u��I+�K�]�mQ�"OjHS�L�T�d���T� �d`E"OJ�i���Pr<��$�m솸�"Op�[#�O02�I�+�7���"Oਂ�
J�0,�Q�� ;�4�u"O��3�F*_�E;��[�~�U"O�u`PDX�{�^Yx�ɛ�y\�C�"O0���e,pYʖ� �<h�a��"O�5p��A$^��|��$�[n&9e"O~D)R�Y7rǤ�c���":�ȩ�"O�� 1C!Gò�b�Y&iSh�0"O,�0�FV�cp,l��ǌ�(x��"O�;S�P#q�8=C��-(�|#W"O�8)E�_
$�!���))`0�q"O��ڡ�=YS��۷w8���"O����8@�Z|�����9�4"O䑘�^5h<��`�*|S ��"Oʍ3`䞏0�D�a�K �3q"O�D�d@�!��I���[~|��"O��q3LI�!tꈘ��G�hX���"O(���Ƅ�e�� ��3���d"OF��k�;�x�p7E�I��Zp"O�@�q�ҊCg,�j��	4<�~���"OFe+��AD�Z�� ��>��Pq3"O�����B�:��!�2�Y�!�d�*uH>˔�գ^�!��7!�O+q��v��4����gH*!�W����x�K�	 @@8�f�*�!�$ٟ:�D�g�E�P�Q��#)�!�D�T�W��<��m��̗]!���;�b�#7I�4%��{�g�)�!�Ě���U`(��T8z��e!��C�Hc�h���ʋe��a#lގ_b!�ߝr�t�%�ts��H3�ŀ}!�Z�E�9���[�Ys�pɥ�b!�dW��N���&U�\e0|�%�š3{!�J!~�B��I;C)
�9��M�gb!�dF`�8\�W�2"*v	�vD�-=!�d҃0� I�$�0"��Ac��!�V�)'̍�lRj�x2�	�!�D��-�h�*�jX%"a�o��!�)I=X�A ֩)nh=Iq�V<a}!�@<v���z"DW�Whz<#��=9m!���8�J�{�#�]v���X�/.!���
Z�$#��g]x�afί�!�F6G>݋���SC���	�q!�$V� ���0A��?{#���TڴBE!�Z�\q�5�B��P"�5R.!�$�.�@��OP0s�x �E�� 5!�$�0?��X[�G	�	�*�:" #k�!�ĝT6��j#�@>9����`n�-�!���#Pnԓ���1	�B�4nd�!򤆸F��J �H�V1�@ź,!�$�^��}bEE�	�%:��[3O�!�d,?B�@���4y� �U1u�!�FJj�ŃEdE4}��k�e["}�!�T$)��P8u`C0�F(�GςU�!��8���ہ{�t���3 !�� �|���H�cz(s$.��t��Ӡ"O*����k{hi:v�S�ڨ�J`"O\���Ŗ��:|p�N �f���#�"O��ᄉ2'$��a�̐��N$c"O��h`�W:�EWaD'���"O�E"��z'XD(� ��B �"OH!��+��2()шT9e���v"O~-[��Y�G��X��(Z+��|��"O��E�>K:5�7^��T5"Ot�0 �)񜸣�LH�\��)w"Oq�C���R鱑僦L�R��2"O��sn�:@q�D�%�Oܴ�"�"OLh�=0�&�s�G�V��LIb"Ol`BpG9��D�+���Y�"OH��� I�8���_�_���"O�H���R�L׋U//�z���"Oԝ��k_w4��J۪8��i��"O��eB�a"`R���-��șb"O��9J�%m��K��!j�U�"ObD�L�,m���`P) ����v"Ox��"�����#Í�����c"O�����H�Ajt��D'������"O��ȇi��7w�i�ү��&�Zmb	�'��l0�a
t�D��ôM��I 
�'�4h���8<̞AӦ��*Gx4)�'{Xy�G�(?�4����	Dj���'@T ��`�?2Nu�am�CX�D��'nL��4���8�|���G>�!�'L(�Q��q7��pB��9Wnh�	�'aR
�$ԶN�\1P�G�4Q"|3�'y�H��L��t�4D����/olD@�'� �2�.G�1-l��#Ͽ_�"�'�n��E�[�"�� :S%|�z�'�ZD����$6����	l�x��'1,Qh�d\�J�e�I(\LxuH�'�Ъ��^�+0H�P�E�.A�Uz�'����S%�5A���q#���5���B�'6�p�/ʌ.,�ȸ�!�#��yQ	�'E�DH�OW�	���<��`#�'I"���)4'V������%��'ob5[��R)�����v(�C�'CH�C/C�!�2�)�jƵ���'���b��Ú,����ʍN�M�
�'�jt��k��̋��T3�� �
�'N���6�ۃ�@�i��'�hJ
�'����P��B�ʹ��H$TV��	�'��&�̎M�"�#g�Hi��H	�'�H��2)��W�Ni�OE;�	k�'�^5�q&q�����K&<�ra
�'ɚ�ʑ���$�8ر`'�a�:lr�'�>�!�!�9(�A�OU�ڈB�'���##��gu
yA�L�N6t��'aX�Ó��5[x��7o�W���z�'IR�RC�ݍU%��!�Nxq��'���+��_�o���R�A�6u��'˺����ÏL�&-Xƥ�/�@I�'	:)�v#.��{��,�MX�'�dE���ζq=����d�/w����'�KO)��݉�$��?�� �F$ R�<�@�|jд���L�=��m!b	�K�<ѳ,G�J�jA3 ��O��ÄJFb�<�p�F�@�"(PT@���%��:Kj�B�}�.0���Ku�-��a��<r�B�ɭ3\����X@���:F��xJ�B�)� ���M��?]0q2��<xӶ"O�)�s�̓HBh�����$���"O���A�z(l S�E$�8�u"Oʌh�3������ɐ\ZpR�"Ov<1W��G��Ԉ���3D��:�"Ol��ӈh\ �� �m�T]�"Ot�����q��}�Џ�X��9�"O��vh5~Y�Pa��C�6�(1�1"O������&k���$X6%����"Ov��E 5���q�uhU�C"O�h&"N0�Ca��ji�<�E"O`E��AZ�;�^0v 3Jǒm؆"O����Z�f����V �7=�x�I`"Ot�*Ԇ<|F��eN��j��8;S"O����	0q�M �K/o���B"O�y
�A1M�re� �\�0�X��"O�|�`�>d0�»BoN$�0"O����L�r���ĄX��X�"O|���T�O���8�mR.[H����"O쐁�#A���8pG�	1ʐk"O�5�`BΞX�F�8B&j`�x!"OZ���7�������H�a�"O����T�H�DYY5�RL� � "O���O?[$vQ�alRq��)�`"O��!��� ,���AƧ"�y�"O��j$�ּCv��Ӡ�_�~��v"O��˴+�<���H�[;�F	{"Or��V�V�? u㵯H�P�T`#"O\-i6�3Z�p��m�4`N��i4"O�(J�.ĚE65� ��#aD��(d"O�ų�*�=ҮY褅��3�|�u"O��j&�*9�$AӢ�;*�=K"O&E���
.C<�PСFG����d"O��
�mW�&� Æ����c"O�L�c�aG�E߼(ڄ��"O��"��zѠ��Ap6	au"O�X��cR�Yu$=Yq(��P�t"O�ЙbEeH~�cC�AY�Q�A"O���2�E�q����㘌=KA"O@ ��A�$�d��cY3�u�"O�91I�-��r�-٤?Z8s"O��;C%C�H��8R ��>:WL���"O�! %�Q�ֈڑKŧa>()�"O�ݘ�"S�|q��Y�K%�`R"O`�ʠg�>��3��T(/��m��"Ov�k�a�H'B���D��p�b�"O���P� bF�H�dݿ81B1y�"O�T�b*�f���܌[(� 6"O�[�dH�Sh�i �ɒ�!1�Af"Ol�Z��%&�~e���O~?V$H�"O>���ɑR���s�F� @�=��"O|T.�/����E	/&�p"O^��r�=*&Q�Ҧ/P{a"O���p=HRwAĐw��8��"ORT��$�!a��Y����~�V��"O���>Vf��P
ĭs���"Ol�9V/E,�0}���Ï1c^�0���ψ��Cc�ǡZi�`���o^�'yD]3�#��U�rX�V�F�(�
�'K�	A ϔ��,�t�V$
��
�'��0�#�Q�A�,`Pu
���@
�'p�3��
C&�� b"+)��@
�'3.LQ�(�*@~æ)�� 6|��'���8qI��UMMA֯ƃ\O蕚�'�
9�,�8/���b$�R�<�y	��� �8����i�`�cEBh�p"O��[�*6����3P���J�"Oz���ã�TYI�	�3K�.}y�"O(!P�MULϴ`�&��Ш"O�P�#��]èe"'�X�ɾ�H�"O�5�M�.
?dd;%�&g:IV"O�T��CI*xƩ=O
x#�"On ��'� � �� ^���4"O��Bf��<M$��K`a����"O��S��L$!A6=���T'9�p��"O`����.@��1AJMW�(���"Ol�9.Q�f��d�������0"O��"��"#�dz��.*�2"O���^���y�GZjL(�A"OL��J��C8���AЏ���3"O�)6��$`JH����"!��x�"O�m[g�o0|! �څn B\�C"O��Kc���
 i�w�"}k��е"O��j��Z<=�huP�Eϒb|YB�"O��DiћH�
��F�2S�yc�"OűDH�� �b��7�ڛaK��B"OBṄ/��Fd�1U��=?����"OĀ1	�';��2UJY�hX�w"Or�ɗMD�+tĄ iFv�l�ó"O��$������c�
<2B `�"O;��Q�m��E�w��A��Q!�"O��*���`��fڈU0�Q"Otp�-X�tHK����RM�"O(Ph�ޢ��|�@-�>��M* "Oxd�4��j"RM§�W�vC8!8Q"O�MZS�nIr�96a��M��"�"O��z�a�&� ��@-�y�fm�"O��W�=T��s��G l����"Oh����#��@���\����"O(�B5#��7��P��� T�`�"O��#��v2�eC1u��,p1"O<\0��5�9r�EV�1�E�s"O���D�_o������A'��"Oֈ����x�` ѲgǉD+�"Ox�� �*�-���3"��`�"O����E�)�0q�q%T W����"O^ȪJY�>��-�e�2jR
�8�"O)�W.�m���@�3(FJ�k0"OJ]�6"�<C�B���q�Rh��"O�8)s̃�\֎]Ã��?w�l�6"O`MQ��1x������0 tP���"O�J�m�<�6-��!B[ �h�"O�5�5��@��J�J��bݸ��"Or����I�2*�5����"OF�"᪝�Pu�Q�`kљ ��"O��� ��c�0��S �� #�"O��:��L���A��'�����"O��rq�놴ڦ� �)�jXcS"O�,A�ꌭ]����v%���N�в"O���@�_%E�"�����h���#"O�L* M�3x��y"s<(���"O ��b���!�4�WO��s�v�Q�"O0Y�	=Wވ)� U�2Y:G"O��#FHW�.�90ID�Uh�3�"OJM[ȈMfTYw(�wU�0{q"OF8��đ�T�D��T��U�jUV"O�i��H�.Gᘥ(�H&A�<���"O�(�&N��J�<�3á���~�;�"O����K��8ei���*�lp�"O� �=K&)Ȫ��tq�Q).( ��"O8����w�
��E#X�IsY"O�i P��\�ry[��B�5Wn���"O�@򕄑~�8��T�@�8��m�"O �f	~��*nYJ����"O��v�K�/�p4�Ջєl�8�pQ"O�I��E���W�2�*�"O��YV�Y:p `lW�2p�� "O�R��
;Y�D�,9z%` h�"O(�8��:U�2�;��R�2���Q"Op��v�3󈵢F��=���+�"OpI ��"��#�Z/GRVQb�"O6xڱ"S��B��P`5@��%C"O��YF)RBz���rHE"OT�"¯^�L��}���X	1H�Z�"O�u*&��f��1��;�\���"O�Xpg)ζz}@��hS c��t��"O����\<2G��zЎ��#�29��"O���"�P�~�rt�"�n��;A"OI+��Qq4Pa�,Q'lzĪD"O�ȇ$W�����J+ꨜa���<a��ȗ3։�R`
|7䑉�"C�<�(�&���i��ֺx�8^�<��L?�i��0y0Ű��P�<	�*�r�e(EO�`"U�R�v�<��;r��9` �e�t��"Jp�<�խ�!z9�e�j/(�3ԬL�<is��Ucj<irbۂv��kU��L�<I�I+ա�/4l~��k�N�H�<馇M3cCM���&���䀊ny2�G(
��OQ>���-kd�3���7"�۲�4D�Lb��A��D{�!W�Y�$���?}�,S�|3�JB�'��	��5��@��b�+������1 �X 2-|P3�ƞ�|�&@H��+_F��"��U<���[�rE�0bض)V��2��j�'�VD��%B�b��d+�v��	�∾^�&M��\�&�!�D�.W�
츖K�
�L0AV!�,�t�pa�Ю+9Dm���3$���)��� ��3' �j3�)s�bp&3D�*���M���z�@��^�����@��Mö�Ⱥ����G\�g�'�d�C�Ň]�(Q)e⟫k����S\\a�%	2֍c0�(-�H�d�ߊP��u��M<F���V1�Or�"g�1�,�`@��E+ ��F�dTZ��*PMފ#��X�ňX�s
�*tL3	(�����R�t�*܄ȓB�f8�7�ơ9�dpX���7�I�2��e����9.m�����<�#�-gc�Ѻ�NN���aamYr�<Q3����� �Ev�q�#��u����G�� �
�&A .�D�3_w��#>���B���c�L�
I��=��q؞�Z%a��gٞ�!��0j���UKN�;)v-�`�9.�.��D� 5�u��nP�
�!2��%�q��$d�@�>��,�{к@[6 �;�����ɦ�#o^�Z�"��q�p�Ys
=kJq��I�������H���\�/�V	���]�H�{���9,��D�V��H�VϓE�x@它�"I�`��a�n;���%09s�:*�ֽڅ���$S6�i�.xBCm͚;0Y�Ĩ���u��)�h�y��$ .��0D�,��E��I-M�t�˖�J�C��뢅O4Bq��@�͈	�aQ��U�n��E!�<�O��&�Y)J�(�S�c�=$,���f��U0W��{D���P ���";��r�8�0ђw�UȂ�E;Y�ԕ�����X���b������0 �2�'�6�1�P���t��yA˫g.��E�ō5�@�*W'ܚ�yRf�2W���u-M�=+t9(C�H�%�˓t�����b!����'~�9�Ŕ�q����`��������p�&���R�w֨�Go@�oh�f�+��x�i=��S�	&>ꦤ�Beܘ�����?�4�R!��Oʹtܨ��|�F��I}"py��ߜ5	��H���O�<� &��,�-n�
X'�>�^u� �Olp�P�
 xQ��O�>=ƨ�"q��\�'�͙-8�T���(D�tg��
Fx< �.:>�4<ڤ�$�M4�dh��	?0犐� i�&�jdآ#�*��B�k� �2CѶT��59�A�=��B䉵h�rq���W�8L�yt�
}�fC�ɾb�����=�&�a��&0��C�I+/�u�'`�<,� �����i��C�əiq���
7c��t뙤g|�C�	#a� $��!�HӜ���ʆ 8ߡ�$T�z��q��@� ����w��$�!�$S�P+��+�t�l��o�_�!�Dׅi�2��f�I�73��C1%��l�!�R2��A�Ԅ-X�Z�����+e!򄌚&}\�'��5:�z�r��	Y!򄛑eŰ�#!M��lG�Q�"ܬ{�!�$�( -��A�KE�{
��H�@�!��l-�ɻ��A�-_═��N�!�䉆X
5�'�T����b+!�d��}좸�6O&5.%y���!�d���,D�T_�/}6\��N�
#P!�d��U��1���ya��H%-C�cM!��'&)^D@���lI��%Z��!�D��M	ȀU�!�3$U}!�$!j��l�n�/"��Kp�;!�Ėo�L9��&
D�xU���_!�DY�+�p��@M�ip�5����e!�X�Xj�C�@��*x�g ��}!��.�n��n͞`Nʰ�f�7a!�D�7u�<���	��@&�%r��V�!�	;Hyx�Ӯ���F!y�����'��pӣ~��`Xw���m��
�'��x�'19ĄB�ҳZ ��'[�p�"�ȧI�\]�6�
X�y�'3���UmPa���m~,m#�'6Ĥ� 3j���lS�{�(M
�'V���M
}wVH�!� e�e��'.�@z`g��Va��{VS�.�����'�2��O�9�@�DcH#'��%2�'���6*�q�`9��DO##e|���'�h����@!\��*�����O6D�x�`8���B4%�1Nb��ʀ4D��a�L)��i2n�5�yC�3D�(��b\&%��}�C*��� �g�3D��ˣ'Q�0����DH�E����	3D�(��QO|"USOS�L�ј�`0D� ��[~�(cR;z^�`�M>D��
�	@����C�,�d����/D�h��'ݗ��x�kK�&U�њ/.D��s�%ڿc�����;c��ia�*D��(�ϗ��l�U�*
�~|���(D�8*��B�C �i��5C���)D��I]R�]��nĘDpt���#�y�/Z�W��h�`W�A�����	�yb[�6f����_�~��q�n��yϖ#4X�#��̈́s/�q�#n$�y�N�h+��PW��l���rs��y�� �J�$��בa����W/��yc
m���y��ۂI��G�Y�yb.G	Bo~E����t�0S��X��y��٥^F���
O�2#�И�L���':�L�f"^�.���3`�P&v8�K>�˗�#��y�i��c��	:&Cf�<1���c;�����P�� LQ��b�<�â�$G�Hɠ��=Zt�6n�Z�<� ����ߩn1.�'J�jM��"O�A�J[X�r�����>���"O���g.ƽYI��@�M|`|:$"O $�B��8f����Ah�В"Op�C�`ؼx��*Bo�%Kl!�"O�`p�R�T���Z��6k�$p�"OP�r�R>�RyӑO�f����b"O�D	)C�?F�db�̓�a�(��7"O��)�$�)c�f���l� m�Q�q"O�L��E?W�����XIT0"O\h��Ë+ẁD�S&6rq�"OD R��i�(��1�ڮ�4��"O�u��F�5�}{��Ëvi陵"O�����A	W�䠁�dXe󨝫V"O^աԩ�?���)Ń�0m���"O��7E_�Q
��B�ĝ(��e�"Opآw��"���@e��,�nQ �"O�A`Po��@����A�-�NP�E"O:�+c�שz�����U8B�С`"Oh@�����QR]��%�,U.�P&"O��ـM��IU��(��Hob�W"O�ej7)+5���(	�)[���"O�l"�gO<b�q��W��R"O0ꡥ	���`䥉��i@�"O:��A��S� �`���D�R"O�9�D�5qHJ�âd6V�ƨq�"OZ�p�(��'�ӥ�V�q���u"Ofu��D(��q�@�	N(��"Oas�G�J�����D)F��"O�T�6I�2E:f� `Z6J��"O�h{PN�5QX�@�AΑ�^7���D"OhL��c̏3he�n��k�ƽ�d"OD��BlCV�ޙ�a�M�佁�"O�$B�	�1�n4jl�9k����"OF��h]���9��,J>h��w"O�1�G	X������k�.���"OXӔOέ ����A?H�Dk"O��q�lʤR�R��<5���"O!�V��Yș�1��[��Q'"O��#揅�c�̐7�O�T�؈�""OX�ȵ#^0i�(�#��9{H���"O�������Iw�F�&dX4"O�H�󨅚^Ҩ���d�,��"O������d2��yЀ\��5@"O���w��%��͔>4� X�"O�1���qU,��EmR�O�� z�"O|�8�nм:j�y�Ҟn�.�*�"OX=�uځr�~pģ����"O��5nU�d'bi�c�`%"O�mw�S�%�V�����Kat|�"O\�1���6y�V�oɊt$Ze�g"O:�Z�%İ��r��%(�ր�V"O�\��#��@6!A��
����"O��e�WB���X(O*~li�"O$��	�:1
���tbƘm|<y�D"O�AY��ŠT~��cʇA[�!�$"O�QP"�\�5�x�p�d�,E$L=W"O�<��#ƘN�8���C�%7!$��"O,�:�&,��ʦ��8eu��P�"O��"�����2�"����a���3�"O��*AIGʑ��˷h�8�"O����f��^�9�+��X�("O����a� ���""lݴ#o�Ș�"O�;� M6��p�
	q2��c"O� �`I��V��pDj��
odI�"O8�c�^����Ol�:)
�"O0�̆84z��s5�Z�6�23C"O�cAI��X��Q �Y�u"O@�[��}� 8��"A!* ��S�"O�p� j���R���C�t�\{""O�h���+VxaiF�k��1"�"O�a�t��9"� q�b_�N�R"OQ��	kg,��a�!+��!"O(|�G�;;�`a�oФ;'�y�`"Ov)��LցV�|$s�[�&Ж��y"��;T��mD���`�L!�F�y���I����'@ăX�d� �N��y`�?H$MzŠ��J̙�"�Ϭ�y�*Y0ER��cζA�BL3񧛮�y�t�=C&�ٴ4Y���G��y�ؙ�������@
V�:E�X��y�eK�^b��Њ�>0�ȹrS��<�y"�ԋU�r�!��=2LB�!�'�y��2�h$d��1��ਃi�y�
L�9( 5�e
F�~��i0$�	�y��S=^m�
1E�vi�|ۗg��y�J��\?8�7�P�s�����kJ!�y��F�+L�2f̜:=�"���E�>�y2�Ǐ 5d���*>�����Dמ�yR%�3gVd�P$O�4�̹F)���y�'^/^E��1�|n݈-��y� �(X0����~�a�A'�y2d�:
PPQ���scfL�q�F:�y�� �L�a�*@�E���Ĭ�y�c4e\|��m-L��%��yR�B2**X�����*��)u�X�yr�˓az@��E;,�� ��yR�ÃT�V����;6~I�4A�'�yR ���z叁�.�\tR%���y��:2����Ƌ:x�8�o���yB�\�<�Vɐ��� �p�����y"�h��݉p ڱ8��I��F	�y" ��TA��x��C��lQ4���yH���q�$��0�P2s�1�y2��G;�q��I�-�1���y��.}��EB�o�	�\X�Œ��y��C�ܽ�ao�ڹ�p
�=�yBÛ�h������ƌ���GL�!���8(pm`�$�T� qQT�߽a!�6w�B��썔-�5Ja��z�!�dԧ�����:x�:�ҷ�$'�!�5�"�H�c����h�#ɗ�'�!���n�Háo+{(us��z�!��]) ڈ͂1��)Our̀1�G%Y�!�d��ʕKv.?Cf��`�H��B!���4K� �F��!)v|C��p�!��O6MH�Eg���'�P0����W�!��K�;�Ll)1�ݹla\t"��, !�H1V ��k"�O�.�Qm��+��_����(���V"�ӗ\���Z"O���4[�U��F�&V����v"Ozt�'(8xrL�5F��i��U��"O���f��/͊8c�.�4)��Q!�"O��C�N^�۪!��-ٴ^pԹa�"O�M��I��W�$Is��)W��`c"O0�@^q}�BQ��4VN1Cp"O�Aa��αQ!�R'��+�ļRp"O�Q�M�/[֨��TE�!�|�(%"O� ���&��v݆��$%�+w�� a�"O�=���',�(A�Cf1w��A��"Oҩ��Z8!�p��A��;� -�"O��$'�%xZv��QX(�I��"O�MP/�C��4՞z(�i�"O�lPc"MqJA����6�P��"O���C��('�:����2Fژ�j#"O�x`�b�o�:-���5[�l���"O,�'hM�G�d����>�"Aإ"O��Ⱨȁt ��o��z�8A��"O^!��OT2�Б����
�X�*Ob�f(�nG� �fIRxv3�'�� fGS�c�$�ۂK����
�'[�:���%Y��a�"dZ&I���	�'��K�!�M:�RG�)0D��'�����1p�Ly�BN��*�hY��'��5d��-V��y�2� �M�8�'���bT ހI�TB�lҍo. Z�'��P+񁋦*��ܣ��Ll��Y�'!��s��ĐF&�����Is�����'�\(z���9]x0À�+:t\��'� 
�"^͑�b[9$`�'�m��D\$z�pѐ�}�(��'u�%3��ǁx����=z�����'��������x�|dC�/��q�J%`�'�����_7�� �@�i�D��'R���!�yw��C�I�!O�Y��'m��ˆ��a @���.GXH�	�'� a����+dm�mzE T3Bݜ���'�zDXR�y�j�A��9(���y�ߚ;���g��#���6a��y���7�T��&�n��5��y�� �'�#�_�qVdse կ�y�	3���1D�������%���y�1|ƌ��E
v|�s�	
�y2MA�D�q��2����Bئ�y" O�Q�t�f�̘0T:�ZF�V1�y���#T>XãG..Q�$�Uc�yB�F���
�IR'�@�pU&���y2
Ӓ9I��Q`'�V�E�cI_��y2LI�W�B$j5l}���h�GX�y­\/>,Ƞ5K/g���	�&Ʉ�y��e޶	�bɇ)�\A����yr���6S�QR�aMF�a� #G��y�E>��ѱ�o�rc��cnO
�y�c�
�Z�[w+1nRP)K
�y��:0P ����3�L�7f��y�I 9��}��xh���-����'ˆ��u�M{i�t� 
7�p�'U%�u��'����D+�#%�"�	�'q��aT�P�>��=y䦖�r��m��'���)E!O&<ᓨ�0>~2�s�'���9���LC�!��]����y�'���X�Œ�������w5����'� �i-_]r\P&��!�	�'��ݩ�7p��P��<D��'�,9��T,A���[s�X�4���'?�e����-�!�2jլU�Xز�')ԁ��b�?��GݔI�����'��P���d���$U%G�t��	�'ިp#/��J٬��e�9q��"�'�t�� �W�� ��ԏ8�d���'M.ȳ��G�N�T�z#',�P�"�'y�YK��7hez�yt�� ɞ����� �Iq��X�/i�t!�H_Bn%��"O�a3�Yq�Hd�Շ�?	^��+"O�)q�BB!>^�yC��6-$�%A"O�eb�+]
f�fH���V���k1"O��KAʈ�I��a�à)8���q"O�e�#h	
Z�i��²"�^h;�"O.ْ1 �"|�M���т*�T�P"OJ`�w������1�k)����"O�Ҍ��
��}�uK!s�p���"O�=a��;Ӻ����=hF����"O��	֡E�`tʤ;�I"m@���"O��ô헁4�����ו{�|!j"O��k���{�mXK�WF�s�"O� -N7ahl�%Ϟ31��"O\P2�I�Af�0Y���l$G"OҨ�e�Ҕ�
) `��&y�ժ�"O�p���;K8�b�O�	�
�h&"O�L�%�G�D*�A�����!{�Z7"O0L�q/P�~��I�\�$8C�BH(�yB�
����̏�~w�r$��y��N&Ӕ�1��U�ET(<�v&*�y"JG�x��`g��q,��f� �yb�X� sUجc�\PV*�y�Q6�����\���A&̓�y�I�-�J�J1�^SC �(#�W��y�e�j�w�1J]Ç�X�y�i�mB���W�I�`����/��y��U:�8���H�v��ħ]<�yҦ.
���K���b%��P#$P�y���� ��ɛ�kޅ_ݘ8�G��-�y�B	1+ZabI�Zf�K@��y�`Mb0Z,�����~bb�ހ�yRg�*(�5.N�j�$�Ҕ��1�y"-�U��T�eO�aY�)�"֫�y.�	L!���C�˺Xj�<i0�Ğ�y�Ɂ�
�p�1
O�Jv53ۈ*v!�ąUJ$�x`��8}W����Nßi!�Ė�5�ȪV�5_�R2�$�UQ!�䆀ش��J 7�Y���
"e!��J�|� ��㑝/BBJ`N�HO!�䊜6�<�#u��3!P��]�!�D�:v �!���l<�%j�36!�d0
�����,�cDr�I ��HB!���Zrb�렮?��	\~@!�DԂF�6�Ȳ�7]22A�ч	�2!��P4�T�3��\?u#V9K��6=2!򄕖d60[��A,����z!�$�7R궅9�HuZ��1�` ,%�!�U�%0���.�4+`�@�/�# �!���,9��=��͂82��4����:?!���s�2�k���L�^x"@��?2$!��Ÿ�XTQ��V*��Р�2!�;��1���O;3�x��F@�-�!�f�
��el^�W�`C"`��[�!򤊏%)S,���\�0�L .�!�$�29~���E��: 8qa�P3�!�D��^ N9�f�C�,��JR���#�!�$�1�����4d*4�I��!�d�r�"A�F ��V L�Ө<&�!��S������T"�2��(0>�!��XI��K��\�|(YH�+!�ğE� �'��9Pֽ�EŔ�#!�%H����>D�l)6��8K�!���v�pI󈉕7��Z�Λ-=E!�� ��cM��x��l�4.�d��� �"Ol�� � �����^%�����"O�X`�dѭ]���HL���Xa`"O`4�ЏфI�m	3���0��	"O�{f&�\"�e9�h;��`�"O��٥T#���b$�'j%.��0"O���GaS�.���z��Jr4Y6"O�ab�Ŀl������< �h@"O��
��"�^l��F��6�2M�"O@ V'������S�}�"OT��j�����C�*k���"O<a�f�ף.�(%c+I1@Ū�!�"O�D��A ��x�G�(l��i�6"O$�����`�"�̀����"OrA�@x\I:TQr��]Y�"OΑ�A��]��1�#9�TE�"O�зJ��&P��G�-8��Hإ"O�x��&�?2ﶭ⑏ȸL� �'"O��P�Jx�%����PD��"OMui	-(�B��aJïJ���ɒ"O0�`��@��<�#I]>j1��"O\��Sd�8�b�Z1	�.-'ZJ�"O�h�B�H.Jj6u�B�7�8]�4"OH)����":������pM�+g"O|Tfa�(7|5AUn�ؕXb"OPlR�"���Pf�M�	�l���"O>�R�% OR�тD�-{h8R�"O���uE��/�PS(Y� �T8��"O���c`rc
R -ÕW�&�I1"O����Թ7�8i�w,�s�4�u"Ov���+��<�b�\0�z
�"O�3�\�����Y6?��rP"OZMB�:Je\��e�v�`�7"O6��p-�`�e�SD�&W��=P3"O�q"��J!"R�yB%�P,q��0#"O�P�D/�7J��n��?�`���"O2<I�>�ɛ$/.c�z��"O°� ��KF͖�=��E��"O�|`��H�(4�l�bk�%�����"O`�+Q��yer�b�	EvKz]y�"O���P��1Z����T/8���"OZ|�����mhĄ�)R!��X"O�x�wh�a�Y�!��#4��"O,������XuF��d;�fX:"O2���Ҋ<�ZA�17��0R�"OD)
V��v��D���ģF��\�D"O�ūah�5�&A
�,ιBE.�0�"O��饃ٚ_x�ث���0W7�t�a"O2�1�+��9�& ',�7C,.��q"O������Mk�5� �=1���"O�ui���|�~,�2�\�a��P"O�A�c3DT5^���`�7'T!�d�a�r��a�����qÃ#B!���t.�%�E;��ģ��MK!�D��dW��IB��Ye0���
P�q!�dZp4,�:�C�OM����C�	a!��Y��|P�J�14��,k!�dіFĬi�
�?f,*�c���o�!�^v�a����v)�UY`���'�!�D@���E(ûy�$���_�<�!��D�"���"G��4hP�gf̽g�!�$�?]�t�Ԅ�+,�ZL٠�@�)�!�dێ�`���ō�[�V= cIC�D�!�T�y�F(�֋�%��(���M�!�� D���N�$���$m�,c��5!P"O �J!�4`T��"4��|��"O`���a>N���]:cpx�"O�AHEOV�)XX�W�şm��Z�'��p"� �YԮ��T��,U��t��'Z\�J�iѪK&̨ыӭ� �"Op�Cj[8^��t����,P4T�g"Op����"fFDkD4��Ȱ"O
1V.P!R�b��#��$���"O����E�(|-�Cگ[�L٘A"O6����.~Z��&!��n�T-y"O�Yz����'J4IY��_'�:���"O𽠶�ܺxD��c.�S�YA�"O6�r���'9�����5:��@ѥ"O�k�KK�2�"��<��L�q"O4,��ʋ����/��mD@ "O |�GM_
6[Q-׸G,����"O\�j��*Y�Ƞ�e�a��  "On(�K�=$��ӶĄ�g#��aP"O��a&"�m�Х��&L%9����"O��K�0k`w�L�l�<�[!�-D��`�(��ڔh % �q�l��A�)D��1&�;p���T��X(���,D������9^D��e�(<ܱ�+)D��h�,�,y�<�ወ��t����"D�x�]�l��$�S� �6qbBK?D���5�lK����NYXDj�(*D��E^�r�ʐ�e�u<E�"�=D����\��B�k�д:X�h��>D��3'�EOp��؀J��м�"�;D�0�A�Ӝl�x��R/�����6D�(sG�)������&X�`5D���p��Т�IS�O��aS�!5D��Q@nޞ׾�&�[�b���3D��s�&C�w���W㝪W����A1D��JRi�)*���"q�8�e/D��3�k���rȁ瞅.�=���'D���FG�lK����j\�!����B8D��`6N
x
عcF��SvF�1�6D�bv�B:E�(�`��͹`�!��"D��QFkE�
�#��	��٫��*D��2�� 3t�Z�L��d�l\�C@)D�@�֌ٵZ�� 郆�9bt��;D���#�6id�eH�e]-GX�-#%D�0�@�&����Z�|�V�+El#D�t[4l1W�bX����x���J�#D���HZ?3�h�PR&�b��e(Q�=D���0���1�|٪3:-���;T�$IT�� ��E�ℛ|��J�"O>���"��[ش�B��-,Ի�"OBt��b��B7�a�_�'l0�W"O��J�Ă�j�֍�$Ɵ�LH��"O~����$DR�9RKJ�#�$��R"Ot�*�PR�[����e���p"O��ʤ�d��Y� �ӝ1b,p��"Oа"���^�TL*���
Zn�kP"O�B�.e@�<cEad�Z�"O��:�L"���BaH:�Ń�"Of��RG[�$]�$�:\'��Rt"O�q��&����kB���S�"O$!�RD�f�氰��'b9���"O�X6�FX�h �`��.���p"O&<��,Y�j
�1�@@�"l��["O� �t-�K�V̀#�C�8�M��"O� �Q�C��0v�,0��n��ZL:�"OD`0�n\J�FD�Q�
�.s"]*@"O�)*dڥ!��t)���.���""O����`�\�"��7���@��"�"Of�2E�W�V��@z`��1rU�������hL�Q���'Q��Z?����V#Q��U��a��c�i�N	i$�'�2�'��bh�oT|�Z��O�L��TɅ�|��#O�A�f���&Z�wa~*���F�'���a9d`A�P�/P�:ت$(v��0$�P��3��!%�dr�!��i̩
A�d��4�bLn�x�oZП�O�Bx��eQ�
rZ��1��)���Uh�Or��D���Hw<io��Y�}b
�9s�\�=9����'��6��Ǧ�m�*hʠ/˙e^R�tiؗw����M?H��ڴ�?����io�:�d�O�6-ƌJbB�"�'D�e��a8b��v �;	�Qs^�n���i���}���|����56��;�m�3�D�t���e���M���ʫ}�P�)��n��0�I6cv�Ze�M�����5���m�D��A�{6Lq���7�M#���� ��9���O���6�i��ղ���{~0D�B��WBn4��'cb�'��q�A�V�s.���+FM��4s��Ē�����4���Z^w�B%�/P������/�C��O��D��DcƩI���O`���O��dպS���MK��C�0И��`@�Xa�d挝_�0����0a���æX?�H��O� Dx�/N�<r�ё@��P�"3�R�:� h@�ɐ|�
ÈƮ�Y��bHs�i�L#"V�x��Z6S��q�WC�%	dP�A�>yĎKٟh���ē�?�����?#�ȑ��MQ�Z������B{Q����	&ml�(!@�_�(1t5� `*��i�6M7�D��H��<��e��jl����8�0c���-�e0���?q��?Q�s���ϟ��Ɏ7��H�#���6���抙zG}�AHӨ. �$�t�5:nB�db�-*�4]��$ʓ1.��ɇ�ϼN�u�S��=����k�i(f�qԽ|����Z�ZU���6aJ�#]���K�K��^F�(����Xb��$[�잯+۔A� ����M������O$�d�O�˓�?I�'*���Aj�?�p)0���3�!H���?y�"�>���:��"w�J	:&�A�'Rm�m����4�Zx�7�i"�'y���~��ë�2���3�DB�/8�t��,P58���'(�b?!�����M�8�0��ń�A,�ϧa�;r��%P��=��G���Ez� +1�Ρ�d�b�DA����:~&��3�y��5�W�Ѯ	����S�@�a���t�So�vm`��	�M�iv�\?�:"ˀc�H���#���!�HK��?я�'���'@����@m�t������8Mܤ��`c>�O��I˦imZ.u��5ð!Qf.����ݘ��I2���4�?y�����D p+f���O7�D�����cYp�-����H�Hp��KC�<(�O����|���ؾ�ԑ���8}8�@��BϚݛF�O�2�ɒ(A]����F��<E��4��!�!��ő�g^z.��&�i��Z��Lћ��z�R��"����8p׌�2��J��њ�ĺ�H�	uy2�'�x8P���	H�
��u��b'����{�8O"7�¦�%���OAڡ��Q�H�F��'Iʻ-p��-�,lOt�)p�  ��   �  }  �  	  .*  q5  �@  L  �W  b  �h  �s  �|  ͂  �  j�  ��  �  e�  ר  F�  ��  ۻ  0�  x�  ��  �  D�  ��  f�  �  ��  ��  � 4 D � M% �+ �1 8 o8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i�B�U��Q��f��?�^�Y��[}�p">�ܴĈ�,��*��Tɺ�k�I�DvN�s"O�X�T@�#�44�e
�>��U�OZ�<���O01�G/F}�F�;Q(�2�$-�SBH<��hU����(�)S�7���{e��ڦ%j�'R�BRIicMk6��$hnb�H�՘'�z�A�5ZV��F�j���d���(O�S�+�Q1@HS��
��A�?g��C�/�Z@�b��ܚ𑲆W�\P7-'�S��M���Q��M��!̅+�ny P�μ��<����W�.a��AOZ���A�,m!��+kE��2$ Ë O*�T��#a!�$U�f�U:�L�3@�&&G
6a|B�|bK?YX����EZ&�t�����'��zˏ�aN��Gۚ"X�4��̈́���'�ў�O������O
$�)�h�*���k�4�Px���+�i3��P�@�61���yb�)(4�����<N�`��>�y��D"J����M�2�*@��K�9�y�ᝓEx^�!�F�?5ę*�Λ��y2$W�!�pa���b�p��!�E�ў"~ΓH/���0@߀L���zz�L���Q%*�hm3.�Ib�A�>Q�x ��	�z�L �5��y�!
8#�>@���Xy£�!��X��(C��F!�
�y�T�#U�:�&0=����U�˔�yBfڍTs
eQf0!��*u!Ⱥ�y���U�9�R��5���� ���yB̑	LR���`U��`W
�y�@�(2�9AqW+q���bд���2�O�� ċTy6����:4"O�ݑu�@%}��p�j��à<��"Or��E�.[����/G�hF�p�"O՚C'�0AFH�(doYy+���"O�T�8Վ�2AF���) "O2ЉUc��f2
h󁋃�\�t���s����ӧ�
�1�S=![���g�A� {�C䉾!��#�$P%[IDd�t'2_��B�ɼ|���qi1
h>\�Sj�&D�vB�)� ��rPaF8]1���@��0��'3!�D��.K$H
�K?F�=k���(|!�$�Zhy��	Nդ��l�<1�!�D��+��I0&Vr��qCℚ`�!�Ӎ|(ʼYL��{h�CV!�<5!� �r-�@F2`��ڡ��U+�d"�S�O��D��+ɢ6�c��1~��ј�' ���c��<e���Ԩ��M�XI��O��I)-0ލ��bD�*��#�iѬ	q����>ᱮP�FC�qo!!Tf�YG��@��k{��с��A����,�X��}�Ɠ�ZU3�)V%@�;E��&2 ���'�""ΘB��e���P�m���~r�)�'�H1��ɵ2��H2��4��T���PfR�z� l����(x����hO�>i�Ki����Ǆ>Iiܭ��'~p�"��!gbv�y�j�"n}���O��0=�g
:�h��ňUo���
G��$�'��S�֯�`-�e�1����'f�x�"Q�4�p�K�L�!=p5��'~p��O�6n�ld
l��n`��
�'Pb��Xqu��ҷ���T�`%!'u���=E��4V Ͱ��W"�yp�H�$k��L�ȓ6� �����vs�YX��á-%���?)Є�(��1���&8r����k�r�<)��7*�[���*S���qen
F�<���L�S�䃃`�kF�4�d%D��`��3!΁G��
g��-�?D�d�D(�f�R�"g.n۴u��)D�����G?"��	�¯�-@�l���"D�Xx�1	��Ch	�����3�?D���B��+��]�%���}�d2D�@x�hԁ��Qj�S��i�e/D�P��������,1��P�.D��R��<<t�°LF�Nk 9D�?D��*C��	 (�	@�D�MS�7�<D�<SE�^�*6�й ���uF�`�!�;D��Ad�W�@m��O����×
'D�$�0K�?<�B�b�PQ�ы2D�� 2d��JZ�kTkH4_)t ���<D�3���3$R������rPO<D�tSs�	����k�*2"�0��.D��{�j�P�z$������C"O D��@��4)�ʱ�ʖ��p��D/+D�z�ʓ��U����bL��+(D��i���;`�p��P+Ҟ%eDq�L"D�@
Ti�&#�p��>"211�$"D������re`���([9��ؒ� ,D�tB�7RP��kY/� ��.D�T�ň��r4��k�9��u{�)D�hs��"2���Ʀ�/R�r@":D��a�!T:Qb�qS;@�x��a;D�D*�DԡM�z5Rf ��rR �۲�$D� +�A%oJ<�n�!@0��x�N!D�dꗭHzz$X�r@\�����*D�Ps�m�- �`A�&y��`l(D�\���_ )�����,rz�
&&*D����Ȭ� '��x,�Yr�j)D�0jf-N�M#�ぢI�d�� -D� ��ҩ2�I��F,�����+D����4<�ȥ,�-:�xD���%D�Lr!��^�vAx&o_2B.}p��#D��!�ҁr���(�G[�p[a�!D�4�nZ�|��(����<0�\�6�2D�� �� Wj���p��$D�Z��D"O��q�Di)����a�9��K�"O�ت��1��s��y���ʓ"O��p���_�@id�������"O�	X�B -9@F`vڜ�:��'i��'���'���' "�'�r�'g`,��o�H$�:Fg��u���'���'$��'���'��'��'�ƍ���U;i�����������'�B�'4��'QB�'_�'�b�'�H8�7�D�;��HjǄ�U��q���'�B�'b�'���'���'���'��=*F�,-J�Yҡ&�2�#K�<Y��?����?1��?���?���?)��'Ta��R�g�$�q��1�?y��?	��?!��?����?��?Q�a�+Lݼ̑��b:4!���W��?q��?����?����?����?���?�gf�G��1j��HRѲ����?���?����?a���?9��?����?��fӌ�R����{G�+�F���?����?a��?����?!���?y���?�6A�-.]z��­��i�n�<�?��?A���?9��?I���?���?i���U7h3@ߦ���� dM��?����?q���?����?����?����?���X<�T,#�FIH~Ģ����?���?����?9��?���?���?i����A����1��$L�����?!��?i���?����?q$�i���'������
�(����Ęyk~ [t@�<�����\JܴM�Vi��(�:��U.ٯ��9�C�V~"����s���	�:΁����"��P�F� �� �Iݟ�Ht�I��'y����?����]�D�ۢ�nl#w�(5~���$�O��h��d�ƃ��:��c��JQ�:�Eݦ��1�IY�'7���w�xb4��h�����O?4��	�"�'��7O��S�'	�nq�ܴ�y�MQd�����0}c �p��yb;O�	w/ў����z�I� Z�P����4+��RE�h��'}�'O07m�=1O�d���Ff���J&�.����.�	����O��Dh���'A`,����t
���͉�XZ!��O����+̊8J��?�?A�OL���/H��ܫ�G�m��@�<1*O���s�L2�-
B�L����>>�$pٕ�s��A�4'���'�6�,�i>���ML�I`��q�8)k��0�q���Iџ����RjMly~�?�8��S71��ʐ"�gb]+uL+h��$⒝|2\��ڟ�������I�\�w�Y�A
ڨ��&�&piP�#E!ILybjc��Z�J�On�D�Oޓ�h�Dր�i��LI9:k@�AI�0E�i�'���	 $�������0,��̀�&w^8BE��/?YNʓ,��	���O�dqK>))O�$��.M!�����19	�`T�O��$�O0�$�O�)�<�Z�u7-��?�bo�`ZF��t�F�0pd J��?A5�i��O�i�'�R�8�&mҖw�N,2WC\�,�܉H�n�m���mZh~2"U�	�]��B����w������x�9UB�G���k����<����?i���?���?!���FB`E�1p�%Z�5���7j��LhB�'V�kӖ� ��?�@�4��R	�x� f�28ur��UC�CTH�<������R��7-<?!���'8,��2 ��8(����C�9WF���B�ObY����D�<����?	���?ن��P�2H��KT:�4sׁK�?A����DȚ�������ߟ���?���J��ɨ%�
�sbne"T�j���IFy��'���|�O�B[t�x���O�a���C
Ө ��A�Ϝ@��V��p��?p�D!�$ AR܌z�雙4'M�7mթn|�d�O����O<�4�����O~˓&X��[Kfy�5&�Kܰ�u-��V�&���T�(��w�I؟ �'="喗r�^-Q�Rt `�u��<���'�8�%�i%�D�O��!�S%
�.��7�<�W/�|a�U�"/8Q#B�����<�/OF���O`�D�O(�$�O�˧?��|���Y�<[sn7e����i���(�'hr�'t�Oi�o���9y�TD���?����F<C\�D�Oj�O1�XkGljӴ�I(F��<�w��2�"�-�&6��3z�<%)c�O4���,���<ͧ��E�7W�@xԤ��
f�ɂ蒱�?����?���n#�5�M+��"����?T
֦X��lRG��J:�Ljf�����?a4Q�����D&�qBV�o"�$hš	=.��I��y��I�V2��z���Ѧ%�'$�D�UB?�h`xA�"V5,��� ǔ�����?���?���h���ąIV`�w,�1.L`d�>K6D��ݦ�٧�ş��I��M;��wnZ�AHR({XNa��aD���ə'���'2�E F�֛�\���~}��h��j���)t��-=�����D�j�V�'������'���'��'sX) Z5A�$��L��:�ZT����4X���?a�����<I���P}�3�x������E�������	O�)�ӏ��t���;��
�gQ�&�Qq��ͦY�(O�5�gh��~��|T��R�j���!L/T�� Hb��X��ɟL��ğ�SCy�p�F(Ў�O��  �E)&n��5�ݴtZ��b��O��n�Z����	����֟�CfE�Q�����:u�����<n�~"�C+d����ܧ�� �����mi��:'�ݔur")A2=O�D�O��$�O����O��?E��"R��(��$�+�c�埼���4��4g�"�ϧ�?!U�i��'�<�H�$	~�4��U:(,���ƞ|��'��O�:�S�i���;&�L���O�W���#F�G��i�OK���.��<����?����?ic�N4I݄�t�ޜpTQU._7�?a����\�P1���ß��O2��'�4E��@b\7cF,
�O(y�'���'yɧ�	��Cp��ҒF+,H�E�ؕqA4�8.p՛ơ�L��i>��%�'X0�&��z"h2e�ep��#(�܉H�p��ɟ���؟b>��'��6��7D%���'4(�`����(~�|��G��O����&��	�����O\!���K7�)�QQ(.�Xh��O��d�-}
65?���̲N�z�SHyR�Rc�J5���W~�8} 1�V��yB_� ��ȟ��I�t�I��O�&��:Pj����9��H��wӾ�S
�O0���O|��2�����^����g}>Z]�SF�p�X���I�Ş��Iz�4�y2�<
�B�ӥ�����!ǁ��y"(D2]~|��rU�'�	Uy2*P'r{f��!�S���M�3����0<��iZHd3��'���'˄�!��Q-V6�q��G �#��dD}��'�R�|���-_�F<�ć��c�`��� �����'w�^����q�j�$?�q�O���� ���GɝF��H"�F�=!�D\�0���a!�5��j��� k��dS֦ub&����I �M���w<�R��W�A�����\!�F��'��'��Z�C�Ɩ�x:�DH4�i/(\�Y�Ӊ�3'�A����dMĒO�˓�?)���?Y��?��Gd��
�o�*�퉵��.{4��-O��nZ2t��	�0�II��韰2r�j�U���vyY߳����O���+��iD�QX:�Z��:3|�5J�ӌS~,�� �@���O3�LQ���O�rH>Y)O(M ��@.���SDӂ.<�%�$��O����O��D�O��<�t�i��%�r�'�*�k�"h����˛��!�v�'��7�-�����$�O\���O���W(S7;�Ftr���(R)P�M�!��7M/?A��D6g���|�;#�B�q�¶��-�1�.�fDϓ�?���?���?1����O�t=(�
�xO�ysg˛	հUP��'�2�'p�6�Ά��i�OX�o�^��&z���6��$D��r�) �C��}&���	��S�6�Ul�p~���0<���Ғ�3C��Y�A�.����3D�|�\������������3A
e����E�ƛ ���ڰc����gy��f�0i1n�O:�d�Oz˧[�ܘ! ��� �cXi���'e���?)����S�$B�bZzIؤƆ!q�X�jp�D�� +����al0"�O��+�?1Df>�D�)ͮ4� vE�ԉ`Dy��d�O����O~���<q��i��m��^)N�lY0 gс~@�@�HF?Hb�'$7�(�������O,9#b��+����G�nx
���O4�D_?Q!V7�/?��
�v����0��۰R
tIZ�"�V��w!R��y�P�\��̟��I˟ ��ܟԔO%U��MT�����sA֔j��t�&=�q�O����OB����D�ܦ�;y[6���ӤD.�+0�� ^t,���ΟD&�b>��!��ܦA�6��5�uo� D�
(B�j�7"<�\�"�M�O"3I>�,ON�$�O��4eR�Aޠ`�GC1�0'�Ol��O~�ĺ<�W�i@^����'�"�'�Ȁ� �?Q	D��-@�S]"̨R��B}��'I2�|��_�"�h�'�6"����\�x`�O�}�GD�(1��6M)��Qa��O Ar4��j~Xhp��Jv�t�a��O��d�O��d�O(�}λ��\R� D�yj@�'ʙ\`���S'��Bڞ(]b�'{�7�4���O�� 1l2��HH��eH�~
���OP�d�O&� �t�n�9��a�)�?��ݴ/�\�����Q��cSIT�Iyy��'���'���'��'^.N]�8{E��;u����l��<]�	.�M�ä��?����?�O~��llP��(��@ 4K�h]>s���yRW���I⟈'�b>	�,?R�����,ՠG�u��C�g=�#�9?��a��*�p�D�3����D\s=���lG�	���d-���˓�?����?ͧ���˦]��A����c@�	
��e�'<��Q���� Yش��'#$��?���?�@�"����,�&?�!A��(�(��ش���mS�)p����O�����I��1C��=�����J��y��'\��'��'���IW�0I����G�(e�e��+�dEp�D�Od��Sͦ��h>�I�M�L>�����zsm�4�@Â�Y����?���|#�K:�M��O�i�b�׊{4� J�F��,<Tk���_tR����1mƓOV�S��<A�o��]�.5+��{���۵B*|MGx��`Ӡ�b1��OL�D�O˧9c�H�"��]�T���,��B���'����?����S���"{��tR�*B�C���Y�N�X�@A���^	�"�	0^��S�zFR&�j��بXq����%sS(�1HBNC���M+�E��w,��JXn����]��lQ��?I�i��OTX�'}R��|�
up.�.|`���W=	���'*�E�i��I�B]���۟��S�? XQ�l[�\bءFNX�Y7�y2O�˓�?���?A���?����	�>�� ��U�L����!C�nxYo�?N����I��P�	~�s�����Cd�Z��u1���94Ռ��(�	�?9���S�'3�xD@ܴ�yb��.m��9�4��g���3�����y�Iq��	?sA�'w�	Py��|p��[2|y "�ɚ�0<��ii��u�'FB�'�������7��&i�t�X��?��'H��?����w&
�ũOn=�R�+�i��9�'�zT��S���4����~��'g��rmVzªu��Q�H�*r�'�"�'B�'@�>���51��Ţ�(|ڼ��F���i�I��MÆ� �?A��Z{���4�0��̊7�@Q2�²G�܌b ?O���O$�ĕ��6�7?����2=����F��#�S���t�'5��I%�ؔ'S��'[��'���'k�B�ʟ"O���q!Ŭdf��6W��޴/�*!k���?A����'�?�1W3����aM�����ff��,���柌�	t�)�Su������4(|p�ʆn��?R��Q"Z����b4���O�a�N>�)OX�״p��eݦX��|�fH�;e�����Ox��O��4�n�*s���"^(b/��fp�. @;P �#��O��Je���8��O��D�<���<v� tH���4** ؁,�(>���rݴ��D�S�T�J�����D��̉0/^H(���� ���T���~����OZ���O,�D�O��d/�/���Z)�9i�o�1 �H�'�� `�>q�W:�n�^Ȧ	$���b˙�@���"�ڞ4Q�����[�����i>�2ͦI�u���Ġ��AL	$[� I��a�l 1�'���%�,�'m��'Z"�'��5qu H�g<n(�U-˧[���1��'.�R���l�+�?y���?Q.��x���9+��s$�0=�$p ј���O����Ob�O��P��Kw�	aSV��橑o�:�u�_?e�@��5?�' ��dJ���Y�(��D�	s�����$�"s��A����?9���?��S�'�����%ۄ�2�099)Ɣ#�ʴZ��[=V5�$�	ӟ���4��'X�ꓺ?�	 �IJ��`7KJ$Y�h<�!n�2�?���8��Ѻߴ��D��6$�Ɋ��N�2C��C.�:�뒆�yT���I��x��ß|�I��O�de��T>tR�AF<f7���s�r�y���O��d�O��?Qi���ӧ�J�Shts��]C�A�ӏQ�?����S�'t�Q�ٴ�yr�(P�� M~�$��C�;�y �����ɀ[;�'��i>��ɂ,���pn�'#�z����cr���Ɵ���ğ��'W^6-
�r�.���OD���zmR�Q���%)A� ;rk� ����x�O���>���4,汁q���u�D��Ɠ�O��G�(��!�� h��2I~�h�O�z��H��@�S�X�V���^�y Aj��?���?���h�L�[?���'#W�;�Nl�p�ȅ0��DH�3T��Hy��|ӈ��3n*� Шƺ"B�ڴ��k4
�	����'�z�#e�i��I�M��U��Ok�_�H��c胸Iz���f�>3��'x�	�8���p��П��(��`��I�'}|$�ň>��Ԗ'Ӭ7���m��ʓ�?�L~���x�B%�"&�b���6$[��RY���	̟(%�b>��W�T 
[�P�T��#cV��;�a׿D$T��EGy���]����uU�'�剩p��I�$oM�)Z��xeQ#l ��ǟ4��ğ��i>Ŕ'^�����"N��7e�q[�: ��F�U�P�� {� 㟤	�O����O���ˌw���"�̐�U�xEI��:��t�C)fӘ�v���"c��\�>q��v�4�;R�D�mR�tc塙�q=2���� �����Iҟ8��K��%�6���<zq*ċ_+VڰAx��?)��a���УK�ɚ�MKN>�g$��k�`�� /+�)Q����?��|�A@Ѱ�M#�O�n����p�RH�j�dᩗ�ݤ(�8H���O �L>i(O:�D�O��D�Ox�y�+E^���`��S�{v��ip��O<���<��i�r�ҥ�'�B�'\�S�W�XQӏ��0�&#� @�`�.�������?�O�a%�$���ga"?[8:�!̅ࠁ����9^�i>��V�'�\$�HR�-M���F�͙:�	yp$�쟘����\��ԟb>�'��7��2N�!M��3;l� ֌�� ��XZ�`�O��K˦��?�AS�4�I��	�bW@~B�
�$��t�	ܟH ��E��}�uGgWAy�$uyb��(4�=��.Y�{��@���
�yRS����ß�������	ҟ��O��A@K̑j'�%����(@*�`E�tӀi�@��O2���O���0��æ�ݙ>�Ԭ8,:p���-���*��ҟ�'�b>��PA�M̓'Ѱ��$Ac6�kQ��5�hEΓJrL�Xv#���%�$����'Y!�q��5Tx��ޗ,�4�x��'YB�'�RX�TP�4.[�8
.O��D�2~"%s�K���Aף�E�`�O��$IY}�'���|b�O/[R�<{R��9��!�"/Ǜ���?sĹಣN�2��������7�.�$W�5���h��	QV@A���Mh��D�O����O���3ڧ�?!ǡ�
^R<�"�V(	����W ؠ�?��ij�e�'�r�`����] s�:�a��]���%*�*t��	��0�'�
���i�I�]��RW�O�:� ƍ*�Ξ;���/ʎG*�PC5���<Y���?!��?���?���< ��V���6��г��Qڦ��3_|y2�'��O�ҩKx���K�+�S��	g�]����?����t��Z$�����	�*�*���9�����b��I�:��z��'9�5&��'[.�÷�.,��٠Ṃ+��̱��'Z2�'������T��r�4~3b����BL/r�k�	�4}�<�0@,�?a��i��O��':�]���L�4D�T4sR���b��$�`���VMt nk~�,0m,��$��Oew�HQ������O�Y����՜�y�'EB�'N"�'���)L�6s9P.C-8IV�˔E-v����?iw�ip��O�҄u�ΓOh��dc��3H�2P# �&��x
3�&�$�OT�4�=[F�~�f�Ӻcf�x�&�
��0Y `ep���x��(���%���O�ʓ�?Q���?��6' �b���瘝��JR�Ա���
ٴ�����r#D�̟��	埔�Oڄ���AA/�2m���a2�O��'���?M����,O�����AҚ!V���J��:�X�q��ۚ(����ԇ���x���|"��37ڨ��vj�U���;5�Q��x�.r� ���˰�N-�f�&���p� �p���d�O np��y��	ΟD�$��yi�U*4m�WI^��Ԁ\̟��	��qnZJ~�f^
m�]����d��3w�x�`��H9v
��#��<)���?����?)��?�,�� YDb�/|j�d��A8xf��0@٦��jMTy��'L�OrFf��.��<��c/�u�n�y$L�#�R���OF�O1�2�!fNb�������1��B��xsk�!P���	��̍qP�'�v='���'���'��#�NA Z�^��G)֬P��I��'��'��X�H2�4,���#���?����Չ�� �2Td@k��Pq��"�>�����'
���.B�Q)��X ��&x�����OPq��^%b�إ��I(�	ߥ�?��i�Ox��C�
�:IJQ�ƴP�\SSi�O`�D�OB���OV�}��Z#"9��ŝ0|�Y�qj�4j2 ����.ȲK7b�'�t6-'�i�(s�@�2�|�zT�Οs�J�� jk����ʟ��I8H|m�`~b眬R�<��S���L����(C�� �/JV��q�|bZ���П��������$(�C^�)tFp��&�8Cx���7��Sy�kӄ5ӡ-�O��D�O�����_�|�ȅ"���q���G�:��'1���I=v��p����Gc }p�M5�1�Չ%=�˓yH��d�O���L>�.O���ƍF�j�J2���i�E�O����O$���O�ɧ<�i�  ���'8�}ap	��qȴ��� a��T��'��6M/�	'���O�ʓ����)
:
����
R��(�"	�Ms�O*H�cD+���.�	��~�p��X7)�&�CC���KVd�h 2O����O����OD�d�O�?a�� Cbt���LΘ?�BA@������˟���4Z,U̧�?1b�i/�'u�%�4�H"m��L�9��\aЗ|�'��OZPXZ#�i��	pg eI���
��sA"O�l� ���D?�Ī<�'�?a���?���N,V/b|!@CM�[�Y�a �?�����$�ͦ)�V����	���O�&�fK�t�4���,эFɪ���O��'���'�ɧ�	�
pcH��w�	$t<���g/��5�A�}�"@�ɺ<�'s��]���]��@)]�n�`XZ�ɂ�Pk>A��{���HNvm�'��O�Fd�`E��X���'F�JgӤ�$�O��N{�ZK`�G�v�����J#k�����O��Cr�k���W���S-�?u�'�� x�b��d��@ 7��t�V횛'.�����	���I��d�Ia�T�V�8G�=�L�'s���P �7I67m�?i~���?H~
�3i��w�hS�)S?����#ʙ'F"E�2�'r�|��"�"<�V=Ord
G��)(�r�Z�D�)�f:Ox��K�,�~��|bS���Ɵ�9��
(t^}��*�8tP��
ܟ�	ӟ��~y�xӠ`b���<ٛwH�|��͍�!t<���/,!	��â>�����'Ƹ��Э�%1T��u�҂�رy�O`��v��,M-&�K��1��\��?a���O�s�ٱ3���:�C%(�0�ӡ�O����O���Oܢ}����(�	��KF��(p�m!p��t��v�П�'A�7�=�i�]2CA�O�ȹ[�*�?>R�c�c����۟���9C��o}~�ϟ�����9&�t	Q���X��padM̬'�'��i>M��ΟL������I;^u�GF>Y_���kX�x0�'�<7m�%}²�d�O��$>�	�O@	cd)�5OvH�r#B�@�Δ8m�v}B�'��O1��\�MS'>̰r��5s !0�݉��UY��<	���4q%��	������U�M�HxR��++�peS^Q>�d�O��d�O�4�"ʓS*��� (��Y�B2�A!��?xx�*R��; 0�E�����Op���Op��	 �ЈY����K�lu���^?>d�$KbӒ�2f�ҁ蟂�>5ӣوd���ID�ˬ9�rY:�[DJ�����NP�|�����Y�P�'ӂp���ŧ̢%��z��Ol�i����6񹳀�q%���(�=I��:iԒ >`������Ny�(�1�d�Y�ؿ!�1ؖǒ���<�3�S�#��-�3��E�ފPYFh���˔C쮭yŊļ(�4i�� <�ʤ�G=U��x�~�� ��B�B�P��\�Q؆�K&n
�ul�%�@3I/�E�E웺j����ug�:t� 9�pi�6�.M��� /�P�D�i#��'�bHO�*_�ꓶ���O��	`F�b�E��Y�4c��!�c� ��G�I����	̟Q�8� +��{9�P���MK�ԤRT_�x�'���|Zc�5�d 2I�`�dJ�O�ֹ/O�0�R�'$�Iߟ���埔�'�����T�KS8-P�`E��]�I�N득��O�O�$�O�T0�a�
SR"��s�G�0�|a"m���O���O���<1��N�A���dx���E�k���A.�8?Ǜ�\����G�͟���9"����I+<o���ADSq~�ؒD��h.Ź�OZ���O\��<)B��hX�ݟ�gOԒ/�YɧÎ�,E��'�
�MS�����?Y�`h<�����I�t
�t���:@3����4<7�O�D�<��:qJ��͟��	�?�H�@�Ot�q^�N�(r�RG�&�����8��m[�����&BZ�e�b���n�fy"K���6��O>�d�OT���V}Zc*l��̰p�*@��ƭn]\b�4�?��RR���2�I�
^��8��f`�q"���F��G�&7m�OJ�d�O��d}R�4�Ci@x9�K'N�(r-ó�M���Z���'�����0���O�*+m�ٰ�3�X|o����I�� �q9��d�<	���~��5'�ba�d�4ˠl4MS���'�&X؄�|"�'��'ל)�Q�I]h��FB�� 3"w�����5P��M�'$�	��<'����B�يv��p!$M/&�`���>�V���?	��?a/O�et�ە`���뵍�5�H��3��k�hP%���	��$����u!ڜ�^A �EʺrZ���!��M������O8���Oxʓ'��@[7�H	� ��L�zYHƋΘ?�A�@V�l�I� $�h����'� 9p�/,�����	�/}Ԝ�3O�>Y��?����$�[��&>U���ӟA���'��X1�)��M������4���d/��hӵF�e��E#ab�z�aΏ�M{�����On�`�ɺ|���?�����A}�"0AVǕ+h�<IxB�����|�'�P����0�G�RS�(1:2��:"�ybF^���ɓ����	����	��\yZw�V������a�10��Y�{��H��4�?9(O<!P�)�Ɍ�9N���M��i��흈z�G��'���'3��Y��'9@��l��<�D��D	ޢ-���Y�^�2��3�S�O�ժu�<wL���в}2�$c�-z�N���O�D��gM��S���>94��	d��|;d�_�%:�jA���቉��O�B�O��c��<	4� �Jf�q`�,��v�'Z@p"\���6⟴q`��KD"I�"�@0�b͝<�ē+��|�<�����d�O��Re���|	�҂�G0�����)V���?����'ZR�O��*����jN3F�N0;$�i���Y�O���O��d�<����M�|j��Lw^A�a*��.j ;��Yd}��'`r�'��I럄�O�BDFA8d*�k�
�����oT�fI��?�����On�iPA�|���!���^��-Yhԫh�J��#�iq�O���<���T�I;z��H 툡jJҐ:5�ùJ��6��O�d�<��!�IY�O"r��5�(�>I��@B��W'&�p�( Gր�����O��d7�9O��P�T�@�&╲bl�p�MCJ��&S��1��M3��?����]�֝G;�A�%Hu?��e[��Z7M�O���x��3��'��Xs�KS���\��3eB��Wa\6M�+Yh�Qo�ß��	؟������Ĥ<Y2��%�E�Z���H��66D0ڴ	�R�̓�?�.O��?���
H��aI�φ�.�&��-˓`ע���4�?���y҇4&<��ey��'_��鎬J�iL,i������G�^֛�R�4	"�c��?�����$Bd�"�棟�8�&�H���#�M������ W��'L�P��i�U��G^�I]ڸP�D�xH��>��-�w~��'G2�'U�W���Á�DdƜ8tmU�T�z,*��B�Ko�S�O���?�/O��D�Ob���t����0�,q�D����:�=Op��?���?�-OJB �|2���7yP��"�B��,��w���5�'uRP�0�I���ɔ���I�o��kP�Q@x�f��.<'9�4�?A���?���$�# !lp�ONRl��bJ���e��<�Q�J��7m�O���?���?��H��<�H�x�D��/wk�b��T�H��H{�����O�˓=�Tb�]?E����L��n��A@�4h�|�4�|��|�O����Oj�ĕl��D�O��$�O8����$��j� ��1��6M�<��K�]͛��'��'��$Ĺ>��wG�l�1�ܭ �LS6�M39;��oҟ��I#D����!��m�v`��I�t�j�� V�^��7m̅&�V=m�������,������<Q�C�0.-(����Y~���U��6-T4=��Ob˓��O�B�C�/NDѳ1+�#y����.D��6��Ov���Of,j��Q}2[�H��B?�A
�(8{�|��J��-��ǀ��'�D�y2�'G��'D�@�+z
����f�3YH�!3tB`�r�Dy�&��'/��� �'.Z� ��(�/C0f��<��g��G��t	2^�|��e�0�	Пp�I⟌�Icy�&�7]I�C!�)dh�4q`	�O�)��>+O\�D�<	���?y���[����h<���Ƽ(p�Ac+��<�.O����O��d�<��e
@��J)#�1��K�N��c�%���T����Wy��'g��'�.y��'H8�c�f7v���d�k�:!�`�r�����O��D�O�ʓ;�t�I����5�C]|�* cu�ƚ
Y��C��M#�����O����O�0OR�'����rM
^�^�!@�i1���4�?����N%m^�@�O}R�'���k��ZJ�J�	�?��m����VNd��?����?��x�T]�4�����ʖO�&YQ��ug܎{;,dn�py���;;:p6��O��d�O��I�N}Zw�P��A��e�*� ��ː��۴�?Y��%���:~�s��}�L91�F�ȡ�ЁS^q��(������M���?����R���'\ʥ���=O|��Xc�c�tA�Ĳ.�PpB)|����ty����O������u�٢D�i���c����)�	����	H*N��O�˓�?)�'�E����EDNH�S�V�ߴ�?�(Oj	j�<O�������@��VI�Xs`�|7M+�!���M��AG�(��_�X�'�R^�\�i�պլ�7^��Ի6Â�`j5�*�>1r
S�<���?����?����@&3Ft8��J��)5�Ľ�P�qDXS}�]���Ity��'$��'tR4h�I��]�*��Ca�0+s�\���.�yR\����џp�	qybg!Q�x��R����N�?��E�'M�89DT6ͣ<i������O����O��b�S��z��L�l����-V��+�DӐ���O6�D�O��ch��f\?�I2�Tm9�-�XWH]�UB�"m?t$r�4�?+O��Ov���;d���b?Òt��X��*F�)Z✢P������	؟��'�����'�~���y�'CJ���7�V�N�'Oߐti�]!F]�`�	����I>l>�G��'��I��F�TY	i�*,�����՛�X��PD��M���?Q���2�U��].?�0��6"ҷ"*�A1�AK4`k>6��OD���v\�-�$%�Ӗa��ѐ�mΐ-��s0��Z6�U�3s(�m� ���<����d�<q-AI�(Y��f�6�<5��BA�b�v�F��y��'2�'����ּHp�p��_]��
ɧ �0Xlٟ��	󟀛E%�����<	����d�1!�neR�LF &�u�Y
�M����� l��?��	�4��1!�p��s�T�f������9%R�rߴ�?�N�d ��ky��'������'2�� R�T��U�c��6Ύ�d).�Γ�?y���?Y���?�)O>���m�5d_.��$�;L2 �1�@�܆P�'��	ٟ@�'��'eB�¡ǅ�PJHI�2�*u�ƴc�F�=�y��'���'urQ>�ɓ'� ��O�j5�B
ѡ X$�DݱZ;�`�ڴ���O���?1���?�i��<	eL�6�
i:%�aE�,3���}A���'���'p�_���#�
��i�Ok��Z|ƙYW#̞/تi�A�T� T�F�'���ϟ �I���X��i��Od�8d�ߞC}"�HF,�=|���i�"�'��ɣ;�D�)����d�ON�钡ek��*Ԋـ*B�YK㩜#���'���'�!���y�\>��z� ���$�J�!A�(�Vـ�kGǦ5�'���ĥf�����OH���H�ԧu'�_���*.��.��F,�M���?Au��<�EP?�IB�'tj8Z� ���j�Ar�Dg�:Imڕy@pj۴�?9��?y�'2n�O8�Խ��դpN�H���H�	�.O�"�|����O`tI�
��2Lk�h�v�j��d	PѦY�	Ɵ\�I#
�.�1J<���?I�'p$���S Hkt�`�O� ּ��4��hvP�S���'���'��"���6��&l�3f�EQF�`�����t@%� �	՟�$�֘�z�j�{��Á6�|��wO�5i��<�� ���d�OF���O��[HP�b/Y�<46-2W�C�]'B=�Fc�T��'���'��'���'Z��4
�z���_}$��Q�I�c��X������`�IcyR�͹��SV��&�[=����mޘ2�z��?������?���^8`�)�[H�s*��r�^MҲ�ӎ	4؜�S����؟P�ILy��9I��윊B�
;9پE�G@�O�8@��˦���s�I̟��	�	���G�̢BB[�#j�TpрB:Qy���'�bT��#0&���'�?9�'��Y�tBЏ���B�]�$�x��1��O�Dд-o�?�$�?� R'~pza�&�֜�,���eӆʓ�pXP��i�X�'�?9�'y�Iq��)j�+B�Z+6�!��C
(�J6M�O~�$�51����}b�)G�C'���E �|���æ=��΄4�M����?����RQ��Gf����ƌ�F��8�WR���o0�j�	Y�w�'�?�D���2L��F֤{�lH �nݦa9�V�'�b�'�Z	ҴC'�I䟨�>��ps3A����ea���"*ݪ!lZ_�I�7!�QCH|"��?���<��X��	P�x�STR�'6F1���iB/S�wr�b�D��X�i�����2X$Ha��
Z�d�� �>�V���<�-O0�d�O��$�<q%K�+�Z�"VM'+��3�[�B+��p��x2�'��|"�'�B��]�j]��N+1��y�(�o;���'3�	��	�Ȕ'd��6�a>��Q�+q(��I�$� ��>���?�I>����?���Ŵ�?q� �t���=n��� ňO]�	BQ�����X�	Py"��2}�& s�n�4Z�`���Q>n�@��d�ئ��IH�	��ɾ5�8�	i�D�f ��6�ێ��F��?1p��'��P���aL���'�?)�'n ��YCJZBͣ!�%�ݑ�xR�'K�@�(i�O&���VY�D��'2h�Z��D�6 ��6�<��f�0x��fͨ~����B ��0�1h_���ٹqy@��Ḡ~6M�OJ�$P>n��D!�/�Ӈ ��Jk�L�y��J�T	N6�I�bh����O��d�O��<�O�Ƙ������B�=N�����>�"H�y���O⬎���(�8PAE�%J�6��O�D�O����B�[�	Ɵ���h?���N"X�	��W�t�v�:��Z؞���ޟ��ɝD���D��H� ᘔ�f�m��4�?�v�S `��On�:���8��L'�N�����#���Hd�Iɟ���ٟ�'(Z�qկ��jh2U�m��h9��,�W�Oh�D�O,�Oj�d�O��Rp��L�����Ị}�,��c�1O���O�˓�?)f"Z��k&#�,u[pd@n��TCc��M���?�������$���B�iu���@/y�\�ѶC��F�
-ڮO�1b'E(!���'�"}�%؋pi@ꐯa~�š��s�<Ʉ��L��� ��o�X!ae�r}b��)=�Dq8ӆ�-n�YB�M��pRP�2��9y��#$�.��S�	��?���c��=�P�r��:O���`�#L���8P��5mP}�7���Ta"t�	�����,cר)�S���!��hi��߽^�6�R��56!`4�N�	J���&��k.N�l�����$�O��d�;u���r�D.�� �MV�?WD�Z���ON�OF�g�'�}��>9�c�9��HB �E*�� �>Tz�;�?O?��F8T�4��%�.Cze�U�mElL��d�O�h��ʌ��'��`K�LUt}��D�v��0��'���8�sUvUjBNˤ\B,Iуĸi�<�Gxu�Xm�S�O0�$��47/��G�1i�H��'6��/s�b����'7"�'�Ga�u��ɟ�C��p�Ħޣ��A�aJ���?9�߅v��{ҊT�+���3ړ_� �W��H��Ò�Z�$f	�F�'�T��W�Ǹ����S��jF{�C�&S"�@7�܄<WW��~b���?q��hO�ʓO�=-$�5���N1����B C<q�m���d�
(/}������c�2(q�i>q��Qyr-��p6�	(�qV�����3K"J���O���O�����O���p>�JAl�D����T���Ӡ=�v-y�邾2�:<*6M`x�l ��O���+��Js: �e,@�^�h��i�d�Ptf�ٟ@R�Y<Q�y��O ��G<���ʰ��T���#���=q���/�5*��zdqC0bJ%|�ax���P�z����1ӼP�e�. +
�I��M����ٱ~8��O�"Y>q����=�L*TĉD��!Ҡ!s��m����	&%u:�Ht�Y����[GP��'_	@�s���9~��l��E���Ey��D�kf� ����Nr��>�H�h�ESL�ѡG��&{M��.*�Z�X���D�JA+�(Qy���rJ�!uy����^�<!��VN깠��T�
��hs'MVC�f��I��ēbH��e�S�Np�P3�%� !����	py��i��'��S+A��)��՟��I
U%l%�U�W(8�u����/���HG�����<��O sA�¿`Azu��eȝX�(��B�'�"<E��I�p��6oH�T)���e�4I���?������O">��ֵ�$s1�ڱW<\t�Ps>��O����K�!j��rb\#,����\*�hp��4���$�x�p�#�AB`&�9���#X���Ox$�A@�#!o,���O����O�=���?y��E�H��Q ^�"����v���2)�!�څ����]�)�֋';���)�b'_���$ix����K�iz�����9��p	��/T���őo�R�'��YPbT=}��d�e�L�/v���'ژ��bֆ@F�T"�=/?hycO2��|rI>�0��3e���د&K@M�EN1:ȝI�O��'���'G�!S��'2�'	P!8���2��5�۪�D�X͜�2#���������*A�az��i���LػK4�y�����9 ×:��qR�O16�lU 0��DyR
O��?��Q�.��f�:vn�`�S�ܱ�b�@��i�^����R�S�m�;��y���[�q� �eK��-��c�O�̝��Ϙ&
�l���iI�Y%^Xә'���ev�*� �])������O"�'6�F��G,�$n��U�č�/�D]��F��?����?�aOS���4�|*��%I�pc��]!�=ô�:�(O�
�O(	&4#}JEb�I��֎�%�X�q�A�'%�����?9��?�)���5-"IC�`���Q�B��b���O>�"~�S�? �!K�ŀ%�mr�(ҋ&�~3C�'n�O@�����f���)��2$�
���{x��0b�%1!���gG��6l���.D��Af���8���� 5~�\�!9D�L;pCќ8F�1Ԉ#m��z��<D�@!R`��]Ϟ��W��A�!�=D����� '���I5"�0(��h�*O>�fKV�8��I�V�"F�@��"O��At�L~퀸{�:A�y�%"O��C�	4D��h?����a"On!B�*�6��r%2_�<��"O^̓�
_7\(+�㖅T� ��"ON\k`� 8~�q��|�n�"�"O��?6I�4���M����E"OΩy�]P�y���j�e+�"O����)��c�:����$�< "OHM3Ň�t`����# ����!"O�M�D,Ǫ68��#䃟u�x��"OD�a�M�K6	�M�(_�T�&"O��H��X�l��9��,޽QC�� �"Oؔ`E	�M���1�!DC*0��C"O��`�V�zeT5D�͆T"9ID"Oάz�N�Wm��XjЫeR`���"O� 3 �ڂp��̂�I=r���"OL{Q
������'�]q�(Cr"O,���F�Q���u��5U6�K3"O*]S�F ��`@0� fmr )�"O����0E���$�ۀM^h���"Ozu��=��$h�3ESZ��"O����ϙk	�S�G�EGF}�"O^1�D�/����׆�#1�՘�"O�RV+]�l�LXb�/i���cs"O�K�K��V|�Qb!�s��<ñ"O^M�Cƅ�=��X��bȳ��`� "O}�#C+4$
��r��K��T"O�h��*�D^}�#�]���Hk�剶ƖH���N��Xq�t�Kb���#�ʑ�6Z!�Dʁ3}b�/(&��}��	��rY�<��c�%b�qO?��=n��̐�BY=%y��0�A!����ӈϞmf��rq�̥R��ĕ�Bt�Ls�@�T��-�u8�eY#K�}�����I�(��y��6O�@��F��b�Ƒ���J/u4�#"O\Dʡ!٬9��) �Q1��2�,KLd�!��"x�p�N�
�x$꓂èk�B�	�r�|h#F(<R5bd�@B�PID�hgʆ4f�r�"~�I��TJ�iy�Dh�@\�W��C�ɠ�3Ў �^cB�J� ۡ>1�OR����7��.%���[�l�)�!�DA�c[L�S�Cz@���~!�JѤ�t�?o_���H�>|!�D�Gp�a�̏<�z5�1��M�!��E-kV�B�ÕG�~CU�S�x�!���bc(���Cf�
��DhG
'�!�W ����Q��l���ǃ�k|!�Q�p���z6O��~X��C��3Ia!�$�(d���v��f�p�e��[!�ͮE�ֹ�^�4P�@c�ɞ T!�d� Ʀ��f�+C�ba�!��mm��
(�P�c��/>�!�T1���ZT�Fu �*5�!�ZP������b�ػ��W��č5�5��ɘWݦ ���V6��9�gZ�A�D��$S�m9�S�'��� ��%�7C�OZJYQ�'	tmc��Y�o��i�uN�/5E2u���$R�=dM#��� |
���kR�4�"m޾'v��"OLh�!G��ִ�a+A�{�0|H�Ą�zı���Oܑ���O1��'����D�
t%�}�U�1����	�'���
E�U���$�*R�z$q "���<7͑�9��`��8����2V���2�W�X��	5e���t�i[n����<I5C	d}PBʔ�d4��p��a�<�&H�+_ҥɃ@�*#�����'�_~����B��is�݉�H�i�OVly�!��G��1�n�8|T��'\p����^6f��4�G��<O*��F�A�E#�'�$����ҁ��Ϙ'��� �:<�n� �/Vp�� �'j� 1dӼPf�A�fK�^�L�+���%y�6��	
i���t.�k�OD���LR�w`���IP�`y f�DV$[n����M5k��%9!�{��k�Y�~��G�T��G	�>�aPNR����2F�&@�{Zw�lJ�>9Fh@�;�2H�`��0��!(�G�c�'e��'�4I���@�2��S:�=��� 5��E	�0W��E����OX x
T+�(^� ,2Z�ֽ��i��h��P�#�,%� U4�BB,��B�N��bTMC$  �b��@���3��B�^�8�2�f/x��i� CXp5����<�~�<O��@�0fC7�FJ1Ob�mM*�f!����
@�A�.V Q[֥ El�L?���|B��6裂hs(��O9h��D�8L��esre�RO2踒�^�_����0�*�kY�]����3G�Z��qᑢt�
�b�5P;Z%��j��Z��Z�(HeA�@�v] ��� g��Y1�LX��N�/(c����.,+��=iN�S��Q��8DG�� ��?) b��zys���J�r��V'�"b���^� ��F4e�l����'�ܙ�SJ.P^�E�;A��� �%�7�2�c��C�,M� ��|!4"�f.�8`������Yd��"P��e��ɢ"�';I�q�@�D?"%��[d>OBx����l��� T� �%&�Ƞ�|R�L�W�&5�e.��$��1�	�(u�U{�fB�_f�K�c��䓟�O�*�٦�-��8gm�9R�&�0��zh��g���� �e�*�hO��Gf�>�2Ұ��m9����+�T����|�#0E"T�±U�h��`�=� )�N^?!�G�)K`���Mͨ'I`��+A�hO�Z��٫���ϒ�ʑ#Fb�ӭ��Z螁�r�(f�,ҕ�{]jy�'`�@0�c��\�X��P�O�� �
�9t��6�D�qA��r��#Ñ�z�t�;O�:� |�����Y1=D�sN?�O�����İ3k�����;Hlna����OO��'o ���IG�Wt�<:5��:E��y���V�p@*�(�L/~my�C�#"��!kw�����Տm/�'�"|r�M-?N�\��<4]��
K(X����`�Z0�G� �.���1Et C�Ȋmɳ��3\	X�b�X�< �R6vLp$bU�B�'Ԫ�KQB�z�q�UF�.(�lQ��I�8�J�"�JO:��Jԝ~A��,b����l�� �T����QX�D~b�ť$#��D�����]�3���K�,�+4A��(O���	�dIB`��J4,Q���`�.�<���\p�T�) Bē6J&��j)#��\�I�L@����d���*w�@�z�N9�	H$rD�vD�-K�r�y�mW��"0�@�OlX �ރ��$W�-�ʧ��d	44���qㅽ���򉕏E��AA��M<7�^�4�',|-�;=�6����1<����؃B��.O�@���
#�
PJ �+�n6�aA@=.��s�K�lI�� ���O,	���3?��}�%����S��p�@���r�� _��Ժ�'�Ӻ�Z`����HA>D�;k��D-�*��%�nvB�06C��<	w�	�.��b/-#��|�|�'_��H��m���{S<��ၩ�:+O�dϻ2��/��X{� �vў��#�HQ�L���I#sgB}�O���dJ�'��9꫟!V�W4��)$?�v(H�qa`,p@,�6:��ф��.��6\Oz5�$�w�b�K�H��'�Y!�m�?\l��hf,��td9[t
�5R[���NL�&F���T>�������~��*Q� hU`�"��"�����(�R�iQ�V�ʰ�`S	4�01;��ŉ�Z��I�6�B� �3*^�ΧIr�<���X?x��!�c�${���1���<�S�2]����';+��5��*(��AE�ގu�"�� �Lx�BZR+����Z'��N����۠LYi����D� ��S�s��	.U	��i��x�2 C6�}�O�<�O�~Љ4'���	���F����A��\��^���2�b%*�-[1��К�C����dK�n��̣�{��~�Ar�����:F7,�����nxa��T+�XKtp���Q$�&!0)N��'"& r�!_���'�"ċ�O�� [h}����!e�<�4�Ս�y��އ(.�V��s���G��u����>3T���ƩS	�}��^�|x���/#�g?)1�K�ZB�%��a��p���v~2CZ�CBp�h[O?�1(�?�@)�ٱnA�P�"1H���O�=��7LO%bgZ�d@�1�b�5�(��F�������~BH��vr\q�=�S}&(4�'����w��y����B�,9>�H�����50s���$ǆqۈt%>� �T�H8]-
5�E��{�\0e��;��}r��$ұK&�	�/<��ff@64s����!�1xb��C�.�eA7��*K���#���^�1���'dԾE��i�>W��9+��<S(��dCl&xP�FFK
g��Z7�ٜY#6��b�%/�O�^��!c`ͼ'�f��;u�"��ɀ6�PW�ڀ�~���I�?L���~�#C#��lc���+�dʓ����k@d���Ar�R@�4��F��7t�)��P�A*l����,@HZG|��t����)X�-�ڝ� Y��y()r*X eg��MI0e!1d�"�P�&��%�iڐC6R��a(��l��6��-��xAI"#"��*�J��f�\�WĐ%0)�]Nl�D|bN�i\����C��~F�
�	ġXf�y���'ɐ��䚇s�	b$��?�~=�Y�Ȯx�ӓ;?�ͻS���qU��M�����1,�p���V�8��� /��5�en�?(8���	��PT"#?!��3c��C�!T��~��a���]�e�h4��P��Q�<@�@ �K=��a����
��1b�'h�	Γ5Ă��Qo�C��|�e��)7���'�����!�n1i��H�>��!��D�(Ѳ��-��"]���g��y��lː�E�n����7볟�=�	.5��E�R�J����m�\EQ�4j�@�p���[���Ę�'$]rNT�j�P0��t5���tJ�7`D�H�>��w�8�3�% �-6lC�����hp�'J8�1U��{L�T���F�UՐ}c����O��a��B%u�z����8k�!)Ŀi6���E�:�
IP�_�:@�	�o
��"R@��0}2�t�-Gh�"���q���03An�$��m��)���*s�E�2F�]��&�Й1*����T"L�
Fj�g�'>�,��4�??)�`ߎ��X�a�{J�KS��H�'Y`]�1��#\a+r)�4F`dQ��\����K
=X t�q�p�*�ʟN(.[�-�>l���:W�<E{RصP]�w���m/��D�a#N�i쨬;
�'x`�WM^.����L�(�J!�-O�!J�q��(�@� ^X�T���ɏ\���X4m���N���#ERt��DS'5�HpY䉁i:~�аl*U[Y
���_��xYG��B��P�큅 �~����uQ�PN��0�t@�@Kxc� 
D�5 �x�R��Ae�����	C�(ja$���TӿD!�Y�<k�t�KWR��Ă��8���˷._a<tt#1�Z�`ي��3?��-M4���8@$R��0�-D�<� ���p�B�M
�)HC6j
<�,C�p���EI��%	U8�0`�B?<sl�`D������:\OP��V=+���*q�|	U`��ܩ��g_t]���1$�闧�6Pdhԛ�j�L��mҴ�:D��r%o����C��/e�2��3�:D�����[.�ve+5EˌA���j=D��A��6V�ȣ��Md�M(SO;D�l�f�Bo�B-#E6 �B�:D������(,I#"��L�p4��8D�8�w�?2��u�J4%�2�&�#D�YGO�z'� m	-`
.�[��%D��i.��M� �D/H'7���0Ċ#D��i�fȿ?z��*b�
4���K#D���Pe�: ��p�TA� U�e��i"D��P��ͨw �� �
C�
��E �?D�xK��I%s��<	`e�+S28)�w�!D��;Т҃�6�aT�1=�f}��3D��sk��km����۲�h$(1D�p�F�¡=.��E�i!B�;�!/D���ď-�	�p5�|�*1e-D��h��W�~X+��,4@H%�)D� rd��=���,�
a�@g'D�D	0��P���I�$�8��`�$D��Z�l��J�^<��F݀@U:�L'D���6�=sJ��v���,�@T`�d"D��@�oGim�3d��{�*i2�2D��g�=g�TP#�Ҩ5�^9I��=D��2��^�3t�4c��B��0�Y��=D�X�a��:���a�D�9�&b?D�(���""�f`{2�� ;t� >D�D�q���n�0���*�~	��/D�� \���b��!:pou�@mɆ"O�ŋB��=Z�̂5��H��"ONݠ�"�1.�ఐ��I�{��a�"O�ɱ�_�@��A8��� e�2"O�T2�W9��:uU�
��"Oĭ�����Ġ\".j%N��yr���a�r1Hp�#ð�8�$5�!�d�-8<��fE��%x��hE�9�!��R�& �Ң�����X�![�A�!��дPX�r
�[NB9��S�$!���x���u2��ӆo��	!�Dο/A`Hr�J�0{\U�#O�� �!�$l 2�C�-*W�rqHC-���!��V&.@J͋������jW!�$��H@ �ړ'<�B�+D!��zް�RSe�B	�<B��	~S!�D�7j�y��)Kdu�բ��.g!��܀h��呱b�2(Yư����;�!��̘["��kE/�*M= �̈́�o�!�$�2T��
��Ϟe;¨�`�ѻQ�!��
b��]�F(�,�[K�V�!򄔻q�R�ɅN�e�(��!�<P�!�d��j�>}��	@�/D^��`��v�!�D� \�YF��[P`]�Go�6�!�䎰�i�H&d������& �!�dA�+f@!-�Wn���֤΀b�!�
�$�f�Z��P���%¢c1V�!�� +r��.M 21���ғ�!�[�,:��%�B-�Ȱ�DKơ0�!򄉢~�\`���}�ɒK�+-!��׆~y�Ua��'p� )��Iж0!�$�+S��e8g�O�+r�%ɂI�"=#!��ٱ����wg�oU�cб:~!��W��A��Ϫh۔�`��ձ,n!�D�0Ġ|(c��#6�������!��O�,���z����$��ň
L!򤑖@%�8�ďԤ͊e���4!�$]"�V%��oͣd0���7(!�8�V���Ƈ�|�Ԉ	�ˀ%!�3;�R4!���x�d���nBx!�O������@���U��˸_!�dǼ6��Y�v�R��,x�#R#�!��9�j�Sq�س1�ĥ���(o !�5y�|����-�2�0���8!��6$�`}�`�B�9�P�홢�!�� 6�*����,PD�Pk��UX!�DI/j�s"�a� b��U=-!���Ĺ3Ig�`��`�ڿ_!�$@,��0JR���HX���ʅA!�DR�ʤ���mJ�]<����V&�!�D@�2���2MX�p'���6#CIx!�M�o�0HS֏�m�\�� �� x!��n�����	&�İP�f[.Ci!�I�Q�b���O��V���͜J]!��Z�|�Bt��XI<TQU�Y9>!�dە����ֈ6�JX�%� &=!�$_"_;\ ����>P��t� �^�	0!�䕶V�rՊ0�J���O4@�!�$
/�� ���u��c"$gU!��[+Uń��'��=V��!1W0)D!��AJ�����'5�����-i9!�dF>3�0��� �P"5UN�y!�dB�%�D�(�J�m{0\�rk�W!��&|�x ��Qs������ !�� �`ĺc�*���,C���X�"Oĸ�'֠Bs�ID�Յ5���1b"Op�0c��{��y��۝��m@p"Ol�Tc�> �j�'h0�8�"O�K�cR2�c"f�{�>���"O�k���9~b�����3"��ȁ�"O��R#חkz��0�.�4`�Ʃ�"O8@���D�a��Pu��� R"O��8T�2� ����	�u�����"OhT�p�	�NCFU25I����u"OF� 6㏺of����J�j"$�s"O�m��E�(��X�1��t�rSsO@�䁇n�P�2�� %X<�{���x6!�_�E�Hȋ��ؐs� wj�b�!�dE SF@�����-�&<�3�>?Z!�d�
;
Xt��G�� ��X����2e!��+p�\2���az��0�\%9�!��I4��c�.��j��3�C�P�!�� [BU�&��L��ɓe��d�!�$�%g��}1�MV�z��h�%+� 	�!���*��C; �t����M�!���U鸄�ņ�F��$Hq@:y�!�$ s?l�9�g��D�L)�B�M$;�!��^�~X&h�J�3lm����A޽O2!�$FHL5���N�4?,��w1!�	��j�҉P�Q~�#!��[O!�U&}pF�S���0r��F>!�Ĉ�|Y�1�����o_;�<X�ȓp�0 �c$N�g�`mPu`�Y�tY�ȓ%D��q"UCx�a�KE
�U�ȓD�E�tI��ڀO6��$��oɐ&ǌp�P"č N@I��x��<���53/r�(Ç���轇�	Q�'y�MP��Li� �0��D�$��'��q˔?��ؚT"M�O��ȓ_f�z6��76�B ���+K��Ņ�\:�r�J�4:�qh#AL--��X��I˟$�dQ,?g���S��]%,��VO�<Ԭ��h�>D`��/���B���G8��FzRAׅX�<C�Q�����y"�ۢ����K��_��8S���y2��3+N���GH(m�@iYb�3�yR��0*R��%�_�s�XL�L���yB`�R,yi��(>��1���<�y2HZ�NB�L�l\�4tn ��L���ykK�A�Ƙ# Β1��0NԐ�y�b��n�Y�ծM"#��i�$��yb	��k>4�H��	�P��3�(��y�h,t�\y�X�zr����#D<�y2߇D����,p�z�1����yL��06q��k�^榸!����y�������S��R�!3b��yb+��x��X�m�D�
��C�B7�y�h�D��h3�G��f����рK�y¨�q����ō�*Y�aSaI���y�ŋ���h�ˊ<A���B���y2`�-,�"�A�8�Pl �&��y"��/wh@�CR!A*m (�Ԩ��yI�aLy���.A���Eܷ�y�
�4'���v&=�"�OV��yB�J�9d�m�D�F}VJ]�#A���y���0Y��q��nڈ	3��=�yb�7i]��[���1l)j���_��y�kC>Mz�X3cTc�xPa�?�y
� �%X�԰j�n�i�A�'����"OĈ�V�K�o���r�ʐZ�j���"O��!����Z"^,�ƥ�;���q�"O���$�[5fE(��&��"�"Oh񠔦҉h��ӰL�q�B���"OZ�"��4����_���V"O�A��1T>�:���jb�ѱ"O��y2@	�C�	r1GO� �,|��"OLd�f�L'$��[c��u�8��A"O�L{6%E�ar��+�)�+ێx�"O -d(�h9�`kŧ�����B"O�<b�
�*Bx�&-ܩN�z�x!"O�{eoC�$#���*ZV�L0�"O��ۅ���T�0�9�,N%W.��"O�1(R��J�)�b)��.h`eq"O"���!F�he���+kv@<��"OR�Q��I�U���=sgv]��"O����ʇ0���R�F]`X,@�"O<���@J��x�ÕVQyP"O"t���~�bЈ%�[9t8�"O8�vϗ5���Ґ�N�]�"O ��$Ǜ&J��ѧ�-6����g"O���m̹��hH�hM!,��"OYK��B���QI��L�%�s"O���N�Hߐ�R(ǽ;���p�'��'d\��eŪ.��X�U�
p�H��'�T�	F�?��,!��#}�t���'h:�K#���p۾�FG�s� [�'S���F����gVe�\�M<�����K-,&ؔڶ&�XN��#MR=P!�@�CP�h9�`�m���`��
4�!�D�����$MR�?����
�o!�$�/>����Ȁ��5�O*3	!��2d�b1�bC;?h(<�5�ʞ(�!�D܀>7<�r&�Yr�q�A�/
�!�$�"@��� ��i`����O�p�!��=>�U��
�!>A0�3�oR9@�!��
16^�`%F�<;l�cP� o���)�O$(
��[:B6����2U(F�c�"O��UR�4y灈&�$9�"OB�����;J�`
c��W!��"Oޱk�H5?l�Ip#�yb�f"Ofy�&J�f���"g!��=�HL	�"O�e{%��%��,*v l�z���"Oq��G�0q�,���1��t�"OB�K����]��(Aǅ#&����"OL�u@�sش��}��2B"O2���D�
��)�v��TxD�q"O������
>��7j`���#"O 钀��}�:�%Cc.�9Q"O��#�b�	����2C^��;c"O�A8�O[92��4�qb�Zd"O�$QF�O�j(�`��\Hy`"O�� ���(>��u��؞FB�"O�D��%�I@��p�� 3�%�B"O~�j�";��$ ��e�*r"Ov�����U�M�c�C�#� �Pg"Orݲ�>V��A�O)�p� �"Ob	�E��=D��۵-�	����F"O��wI�-��#t��+<Dtڣ"O��)c-��}�,A��.^+h�� �"O$U ��[1��KTo�2^8�v"ORP"��P�{2�pv�ճH�0�r�"O��k�$(�)����0X�"O� �q���Ք�D��� .���s�"O>4���Y�h[���D!I��"O8�$2z�`���i�=�C"O���CL�u�
�
.%3"O~��#�˶E�̅��������"OX���`�X9$�ȴ��;Y ��"O���ץ�F.p�d�ȣ���"OL��+V�s �	I��L{n��"O=Q4@��|����k��Ap�t�U"O`|@r
Lޚ�3K ���u B"O|e2���
?��er�����p8�'ŰQ��8<��+(�ȹ`Oh�<�e�}�:1S���j5L��d�<1R����q����>��P�%�F�<ɡ�L	~R�p�N�L����#RE�<q�iJ�-0��V#�<,0J	� �l�<�Q�_�T`�Y�R��h	f)]�<�FP�;�D9��	�pv�qW�<v�ŎH�}���A���K���K�<і� '\��![�O��5[��JI�<!� Ӟ:�Jy�f�	w6P���ZG�<)D�W�E��H�F����ٵjG�<�K\(���K ��=J�,�	��F�<ƋX"{�u;R��8L����X�<cX>@�rYP��kX}z�m�W�<�QL�@���x���p����@�Q�<���H����z�VA�
�ymIQ�<!�M�*�z0��!�F�|�YC	�r�<�u-�9�J�yc�߯WJ;�U�<a�LYYx> ��aO,b0Ĉb�C�j�<a�O�3|T6��FS���u��e�<�g/R�$�S�[S ����[�<��EG� �r���S;��|���[�<���g�vIKeQ!h�P\��o�<���R�/�ژ�F��g�<٢n�i�<y6a�Z백+A�̐i|(�&GM�<�'ǋ�|�����ǎ�����p�<�ҏҜX�LY�F���f`�ƺm�<х�E�H!�Y0c\;>�pH��o�<i�c�A%�sv
Ze�����l�<IA O�Ld<�Q󢒊,�� �Dl�<	V�5a�@�[�'uL`X��\|�<�'�z��40�kT�Z����!�x�<��O6L\̚�ǽ=�H�D/Ku�<Q�`�3lo(Ԩ�����8���p�<��
��9�����6w6Ѱ��h�<��%\�-�z�/0g��G�I�<���@�@3�ҁMȣv���)�k�<E�٬3v��BT� �z]�� �k�<�5��1+Ԫh����d�j@XU.r�<i'�J9p�t=8�OZ�5�`lP��j�<����N@��T}D$�R �d�<9��K�8����]�`��$��]�<�ǌ�Y��T�B
�����V�<yg�U;���ҤN��{�NYq�S�<ٓnӠ6O*�{�C+�ʄ�1AM�<�����P:� H�m�a��DM�<�e���lDY�7$��;8Q�KL�<QU"I}� �%j�-"��I�u�I�<�$cb��L(d$W)Cm����E�<	�jO\�
m��.C&a���4A�<12��S���ĩ��y$����˞|�<��� �r�X��ȿ{��MʒfGz�<�F&�=�&�k0��R����D�u�<� xU{�ß�;��4�&ی{�c�"O.�C��AH��p[$�/]>�Es"O�T��%(�����͍>�f���"O���Fj�������H����"OT})n��
⺁96�m ��2s"O��Z�MEM�]2&�� !��"O���C�S��q������"Or�;�I�_ 
�O�	*�P͸�*O��Ӏ��3�M3��O<q��h�'��i���
H(�x����:]�p�
�'O��xu�N ��9k���a�R���'W��feJ,o0T�@��=/]�q�'�� PL �������䍸�',t�:�(-%�,H�dڽj`6u�'B�hbJ�F���:6�[�8�"�"�'&,�Ƞ��7e����FR�4�b!��'�� ⁦ֆ!�����m^�"�L	�'�~|Q�R���ީarx��'�Nm��� �)��KT�U�(q�
�'���
�H�)"�{�KεR���
�'䄥hQe�=r�.��S�@]�@\J	�'T�{s�X�:�b�@V�G��Z�s	�'v\� ���/��)�el:3V8}��'`�A��S�x�I��z�.t�	�'x�ĸ$�ʭ�����o`����'��:���J��<��#�-mN��'��Q7͏4%8�0���3���'i�X*���!L̤4"pB�.��
�'hLx��Q57@�	,X<�@�2�'�P;0��,6>@������-"F��'�!`�������Ű+��B�'�b]���R8P7T  ��!)����'2R�Y�IR�$�2���N�,b�:
�'V �{� Bb`jɠ3��b����
�'��Y�m��)�
ɢN�4̃
�'�"���ӈWN&P�b'M�5��:�'x�B��S:R����PD�'��@��'1@�'m�#Hv���׮Ӈ"���8�'� ���� �PJ�@0ɚ�P}��'�К�	PvD��N��:A��'�0
��pJ��0�����Z�'P��k���?vi���޼s���'��"6��"z�j�1` ֆi��E��'����o��l�,�k������
�'��̉ӅŦMV&��q�[�g؁s
�'��j��8�t�R�P\\��a�'���H��%9m.��D^�XJ0�y	�'��%ӆ����E�Ύ9S�8j	�'�\���+K8��4���?d�	��'��R�N$z�ec)�2ҡh�'\���NV5U����A�A!1���:�'��ł��0)+��t,��.�,�'�<�!���+t :D&��+�1�'1�:����!p��JR����'� �3DX�Y�9p��]vE1�'AFѰ�C��\JjƥN���'s�@�!���$,�$�O4����'�Z�1��٢m�^Pď�>#x�	�'�^̺�'G=Pe���@�N��Y��'c�%J��	�x�N��F�QԹ�'}
 �Q.�&�h�F#�2�`P		�'->x2sI�(	z��k���(��J�'[��s
Dq���bI�W���'ݬh����ak�1R禘���� J���f	c��$�2�S���A�5"O�����M&ـAa!`�N�A"O�P��C�#eFY8��sx�k�|�)�ӝ[)���φ�D%��9�O�*:��B�ɩKz�	P�ȣ4.��r��^G���ݽ6����g�[
7֬��	D�P!�dA>;P2y�c������;1!��+�Qٱ�ܥb^DRqnݹ)-!�DԢ*TH<�q
�F[�\!BnQz�!�D�D0��aKT�41f��D�<���
�!bR��}8v���I�(�HC�I�0���zէ�LJF��VJ�`ZDC�Ɇ{����sHT|��X4�ˊf�C�I�+���˵	ߚR5��[��ȩl��B�ɔ4��� �O�#U��13��L�lC�	�h0q�'H�4co�0�%Жl��B�	w�%��@�(�����n�Q� G{J?��!5I�bف�oڪl.8!��'D�ԑ1O�*5AP�(�"حo�	2$#&D���Vi.��!Ud�>|eꌑ�A6D�H��ᛏu$�З��� Hw�4D�tqwJ��L����_�Έ�'%D���	9>B`�6DL��|@i�'"D�,�r ǼZ@a�`��B��3��C�	K;�t��c)j��HA�@>*��C�I.&|���B�K��ˁ	��x!x�d0�	u��~B��
�Ҽ'�'�Pź���y҆�+G�|E�g�++s0�ص.��y"ߦx�`����%��TiB�V��y�* �
� Ѐc�V�R|��
«˒�yrn�ze�D�d�6{"�%�"�̠��Or#~z��X!��d�84K�x03M�<qT�%N�t�(�	ȳ6�V���K�]�'ax�P�V.�����6`��܈3f@��y��J�.��Cp-�J$�Ղ���y�!^�\�Vђ X�8K�}ٷ���yB���#8�c�ٜ0Ԡ���(h�y�@Z��5Ar+�!�T�wL��yg�p�,����"N�*��Vf�6�y�V(]_�<�C�H݂1z#�2�?����䓢h����-:ΰ�RΎ�V�4�Q�_!�$��!�T�ʌ/{.|BF̑�y>!�$\+�u����Y������8!�d �,H2u��� �~}��㓀]!�D\Eq$�97�Ap���IS�{b�F:v;D��9Q�9�n��^4��'��O?�q'�
9�p�b�DŅ	^ք�1n�L�<��NC3\���Č���y֪
G�<��FC�.�,�B��/D|X�R IG�<��XJ�X(¡�Q�*�:KA��<y�TޒH2�ԇ$�����y�<�#!A%@�� �"L�\�����Ayx�LGx�del��ąq�4I��.��C�	=pv�\�P�0+d�гAޯTجC�� Z��@r�ԀlhZPj�HȎi�B�	7Qv$}b��C�P����e��lH�B䉁bF�M����9ӥaX��>B䉹cY�a�an�� �k�\�5k$B�I�B��.�:VV�q�c�#!I>C�Ik��B��ܰv�`��C�F=~B�	�s�@S�d�q(�q�$-�+�n�Oh˓�h���I�yIZ|�	ǉh� y��h��,!�dD�]X�pS2͓�e֊�[Em�9-�!�$$&l��c��)3�ܕ���`�!�� ��W	�ID][�ܹ&�bl�w"Oι2�΀eXfdQ�oǕ�hm*�"O[�+J�@��+n2�9���'��{Ѥ�w%ƕI(vH��	
9�D��I�RT�%(�	�	\�"��t��B�	
�����(�e�F ���^T�B䉟j�*��Â?	�8|� ˄@�B�	���,�T�,cr��7ϊ"TB�	���Q� hO���� ���qB�ɣ4�4��3��ʴI���L�Ԣ=!����'7�	E�w�e�d��(n؎<؆%��Be!�@$~KD���×:�XȊf���h2!�$J�9J��`j}��ǂL>z�!�dQ
G����2H�t���Y���p�!���H�Z��"��_ż E۔�!���uDB��������0� I�Q�!�$ǐ�*�u&�Ů:�bջ&\�'ia�$Ο*G,�pN��M�4sG����hOq��y+�'F�3�@�!k,1�aZr"OH��ͩo��jG&$�I�"O���"��?�pň�=�x�"Op1t�W'���������T��"Ob�O�1�bʑ&�p�l8'"OJq�1(K�'�%���["~�k���(ړ���H?Eװyy��F�#2nmӐN�E%��)�k��5c����@�e�3c>
��	�'~ ;��\�$PȤY��)V
�	�'�� n�.%�h���Q�;�|�C�'���8%��T�"CA I
L��?D�H!-��k'
) �( ����;D�@�)^~�K���Mv��5���O�⟘�<��h��_ټ�
1�[�N�\a��|�<Q�a�rJ�fD8 ���@$LQB�<��L7E��="·�\}b� ���c�<� ΋�]�����a욘��^�<�G��g܈�A�i"�(�`�<��FY�X!VI����a��`�q/\�<���9Z�L��fL �l8!�JT�<)q/ƀ����+ƲgW�����O�<	p䎱8��(�1jįh�D�K��I�<�D���SD�Avȅ*r#���"�AP�<�% *�����1q��l�'�A�<��'"L+'kŘB��1ge��<ID�ϯ�̉���/b���A�_|�<�$�+D`s�
����26�C��bI`��VeL�C|8A1���>O<�C�	?��B�NV
��Y�P�H�cM�C�ɞ3�z�S7��|*̵Z�B��C�ɳW���B��/;{�	#T�>YVnC�8;p�}���מ��x���
|hTC��,BD~�y%��3�\�a%
`8|B�	�Y��v"��ps�^�j�a��1D��XG���U��C��:%�AI1D���AK=(������Ԋ#��m;D�9��4`&x���.� ��8D��A�D*m~(��tZ�<7�%+��"D�$��D'k���#C�תҊ�i��?D��2�eQ�BA"�/�4)�D�i#<O�"<1�ЍIx�q鋃��IY��F�<A�(�V���B�2	� �&d��pD{��IV��L�ĭ�1L�0�P𪒩<L�B�	7��i��ז��LB)l�jB�ɡ�0��^�
\@Ң_�O�C�	'!|9�ڙ\��i��I#CRJC�)� �Ka�5q��!k�M�'<��!��'!�I-U*d�0��V�*���4�jB�ɩg�|�Fe�	�� !�e�K�"�Ĺ<�(O��}���(�!/�!Et�!��nY4��ȓ$�]
�NM(��y0"U�=o ���C `�N[��D�#�x;˄���4@���aH[�
<I`�+��LՅȓd!��eF"2��K�[�ȓV�@�A#!Y�}X� {�
�� d��ȓ0Cj�#U�M?�f���V�����?�ӓ��Fl{"I-:@j�j�'�!�D�G��P DQ���,B`����!��Q&N,�A�\9V�*d`�nי$�!�D��δ�u&�#b�r|H��	�`�{r���&r�5���y�(���	�0O$���E
j��#Q�W!`(����|��'���
��ɒ3�U�������K>)���i�=]���It��u�4���S�ht!�DI><v�����U"wBI"<�!��E&!nru���I
#���1��F�N�!�$�":���HFM�b�T��$�,t�!�ԩLF<�`���%�"�2 V��{b�$�&>�L�����V�2H �	��!�$F/�^	j��-D�Z�D!�3�!�$ �{>�$kPm�z��l����d�!򤚖BW�t��l�.6��cE��Ey!��]�ظQ2s J.F�@�����!�<o���f	9$<uѢJ�	v���8O���e�ZH%�P��B]�2s�p��\�E{r�I�b�2���U8����DzC䉓r`�,�|��}��I�P�C�IXH�b#�1�UH�`��>��B�I��F�h�I�|���q�q"O��b%�gբ4���ڊ?�H)�"O�=�T76�p@���J�P���"O�P挅_̈H����]�N�˵�'q�D�3�אt��D8eb߶�B-` -D�X`f���C�>xr]�s��p;*D�T#��;I��	�d�-�X2��4D�$�q*��Ps�M�AhI�P|�S�6D�`(�B�?c��=i.\7:�d�s�3D�ls4�]�	@²n�.�v��t�1D�����׶x��dA�&ĚwB�P�� �O��=E��K� 8X��ܤ"�4:`�%!�Dm�JaBf�ƣ?�<"4�%�!�[���uD�ą[�AX�_b�!�G4�Q�υ$LT�BcӍa�!���5O[�mȒ��I��Ͳ���.�!��Hm;��v� w�.a�A�5y#!�Q'
Q�#��dÔ=K���!�$E n��"Wl�J8�C�B�!�δ��#΃vxB0(P�Y�"�!�$��4��]a�,h�T {�!�SMCz�	�L��.�tʢkz}B��$^Z�5	��@���Jv��4��B�ɠ6�*(�NƖv���Q���j�B�7[� `vApG��)6@��@<C䉡`�`��L�I�{�XC�	G�d@S7̄i@6e�%J+V�B䉾 À �b���ItH	xBTB�I#dސ�hv
]>O�,��Ɔ5ZB�	K�V2Ƌ6L��0�B�ߨB�I> Q��cu�LN:��w#�J�|B�I�S<9(U䂶g}���+9�C�)� p{Rc�*lNL5�d�RT��[�"O�Ѩ��ޭF�6����6>b<Yq"O��p�À<=h�r�-ؕ	.R��7"O�cp��tG&� ��W�k@y$"O��	f@H�SS�H��#�hܨ��1"OrIZ��ƥZF�99���Y�v�2�"O����� ak4��`��Ԫs"O�D�+��� ����!����F�O�@ I򪉩xVJ!�7*�Tkܔ��'�\�I�)���T����J�D�֔3�'���@4 \��d�75��@�'�`��wf�2!c��[���4�����'�MCfO�\W�-�a�[ 3|�D��'�v�1pL�pj��1�n�.����'��|P3=b'�#�9�00��'F�#�� t��(q��8���'�Z9�1�ۀe2�i�`�Y�xW2H�'�t�IU(	�fy�WA��=>��8	�'d��S)��.2�:�D�#.�5	�'�|�QP�/�v܈V��S:4�X�'�f�c���.��0�fE��G�Pd!�'�0�]�p�t���DyH�q�'�D���醲FF1�����Q�'C�l m�J:pYгǏr`@��	�'��S�g.$bm� �+`��TB	�'q�렢Q�O�����!X ̀�'(�mՂW����ζ_��@�'i�9H����q��a���:�t�i�'$n�P�[�QB��*!��?}����
�')ʐq1hޙL�
0� K�L��S
�'� T�*P�O�Ą������<3�'�IR�J��E/��� c7xA�
�'֤t��d�>!5�]�i�,}�t��	�'r�z"\+?LTqI��+t���h	�'�i��G�s#U�w=�V5z�'*$ ��t����ug,*��}�<񀥗tji�PA�v����c�|�<y'�e���@C�>$((iB���5!�$�X
XI� ��O� 	����d!�D�8�t��R� �:�*��v_!�DV�&����n�.�.x:�H�F�!�rJҼ�ŋխb��yQ��u�!��?8�Z\A4�͖W�*�K6Fľ@#!��5~݊$��%����RD$2!�$.-D�E�dQ;�L�11�_;(O!�$Ő'�*��z���1�gٚ35!�D�g&�"w!9O�E ��ڈ+!��Y\.E�e��z=��6�Ռw�!�D�T�.��vO�;8�,��&R�2�!�A`�\�[D�Z���(�f�G!�d%]�,e�TƘ����� �9n!�d�u>�,z���^"�aڂs�!�$Z�J�:�nܪbD(�7+21.!�d;`�)`p%)Y,�1;7��]H!���yfM��iwܤ�p [A�!�D�M�8T�6E�#.(!�e@ڸf�!�fNBn�c�XO��fm!�Qw��J�GOO�03-�%�!�Bu����ġ��2z��J5�!�Ă�:�찕��6vO�!�K\�!�DX$i4�H�#Q�
M�eS�j�!�D�%x��u
!
�T�Z1cI�y�!򤗸Bj�B'��!2�`�rա�%:�!�D�'��u�d&"[�!���70�!�� ġy2�âi	v*��1`� cs�'Jў"~`(��K�V�ɣ-Fp�bB��y��Ļ#� eQ�\-4��ґL;�y�%ıyi���`��M��y"��o`,;��E�	U&1!�	G��y"aVM�$�p��<.��� m���y�˃�y $�ă�%4r�� �� �y2lU'iy]��eK5r�0c�@҇�y"M�=)l�+`���%���yR$�m(�4���	�@Y�����?���0?ŬD"�AY�͐�b��x6�Ux�<�f��0=�*xA ,I�EC����J�<���&$���Z!,�0*l�ѱY`�<�J@#�|<��G��z��"g�<��"Vg���kCd��cJ�ѐ'�J�<��P��l}Y�B�H�0��	A�<1Cљ^�$%��֙v����@��@�<�jH�Y2ڕ����+}�"��#�Ht�<�GС#\*�붬�#e&��1�o�<5G�dd�(�
���@�m�<�`��5��BR�5�7Ɇj�<�b/?�����َ8�X9�3)�K�<Ѷ�Ւ1�:@��3_b\u��$�C�<��V w�ȃ`-�.YLH��C�<QТ�`FDp�E_�?In�SH�i�<�eHޡi�i*e��'<�@��&h�d�<�FE_�tj�O�2rG�\y�<q��$;���,�qc�E�3d�{�<9J�!�|��&o���E
�w�<CL�>{@���F�ޞ��l�vE�v�<�`C�<�Z�B�J�VȜ�0�ȄJ�<qC���R�3��t�`�N�F�<a *��]܅Y'"��H�!;g
B�<AF,��-Nh��b���G�b�<��#�n�c煈�Tb���X�<	.<y�~%#��� Q������y�<�&L�/3RٱP��� �dor�<�3'R�};�e�S*�,�(A�r^m�<������4� `P%eݐ0,�`�<9@�w��������ٖm�`�<��̚k���B|����g&Se�<�E�1)��*�R�2��@R_�<af�I��@�`�*n�|�""�a�<��A.U��Ƨ�(~1BL�ρa��d�|ȉ�ǮG�=�p\b�nZ	!?��ȓe��`2�kܴ(2�kA�Ă?Y61�ȓ4���A�:!z�;��Ά���ȓ)�$�x%`N4I�<���T6pHń�K)�����2`��b D=<�n��ȓ5�����O� �քb�ƞNHZP�ȓ+^
����W
�X�GA���M"f)�v�G�G��������B�GZ�<�wɛW���Pk�6Jp����^�<��R�MF�b�J�0 Q�u�c&C�<�A!�
T�0(T��0ߊ���|�<Q���`}J��F�.t���x�<Q�H�6qX��1�B�9�����Ur�<A��^�i�@qy5�M�6!4D�� Jo�<i&���p%��Pp�H�{��<�.6D�,)�@Q�=�4AC֢�.}�H ��`3D��`4鞐c|�l�2%��q�jg�0D��8��!�4l;7I�:è�Q�/D�ȂU�K�z��HђG7dy�@3��-D����$^� 8�OG%NB¤�!d/D�� �1�atSt�{��5H!�'�H���Ӊ��M�U.���@piq�,D�ɷ�Ï]a�Q�/�.?j���*,D�xҨ��Q7�:RD��45f��J+D��*���kWl�P"'��|<��:#E*D� I�/A�d����è:)��C�&D����Z�1yBQ*�6p�d\���6D��j�6q����o��
<�Z�:ړ�0<��o�|����V��S�6t�S�~�<�E�TV��ꕪK$^1@foE�<��%^7	�*qp�,�G�����S}�<)f�]�@������A�*��as��O�<Y�CB����d@R��B�BHp�<�T�6�Z,!��Y*��WҌ$�����KV��Q�]��\�a��2�R�$��I6"n��36G�9_���U�.eX>C䉘{����t�dH��0�XB�	j��z��ʊ"|�|ӕ�{�BB�	�KN��ȴ�
W,`�9e��Xj.B䉩x��lGM͌�Kq���`B�<v�PR��	'�h��o��P�PB䉊c<VD��.�:t�(u�U�ϢO�F�$,�D(�S�ɐ�4%��)�R]�l��N!�$�+t��ӠoO�!i���A�I�7!�d�
{�@�J�I��AvTi�f�!�Ĝn���I�o��[^�H��KN�!�Dݷʲ-�&�_8OZ] Є-6�!��2m�!�:@KdQ(��B�z!�D�$4�`�p�L�8H��*�◜r$!�D��\�2-����5�:�A�p!�"6�<��ƞq�Xtp�@�)!�$��Ɛ]2��0mtR ʁꀎU�!�d�S�y1��>���;+�!�d<#��і���#B��RW(�: �!�$� J!T���+��?�6y��Qb�!�$�58� �*�/u�B��P�I�#�!���
$�(h0bϢ;�>��%��|!�d���8� �ϺR;V%�C�	x!�$!?��v�^8�E��H�!�$��+&��; �D�7Bµs���qp!�D��)p�,B]L��R�H!�!򄂔8�3��8L�aC'N�	 �!�Dʵ= �y���L�=�,�*�,�qp!�$/:1R˕%�u�jyS����-!�db�d �ԦP���U�TAƳ�!�Ą)�19�(FO_�]�j>�!��W?'B���̐�T5X
�'^��!��{��P8p��AE�گ!�Q� 8�F�B����m�	<�!�d�,M�m� �B�w���׫[�)�!�β2���!y*,L˕		M!��3��ã�'E��(�E n�!�ڢ0��D��(V���YAC���!�� kF܂�/��D6L����!���V���ؗo 6w5F8*�DV�i�!��R��!��KK^ĳ�#��6�!�.h��@�X&�0���#�!�$F��(��UHzw�i��� :!�D�'��MBsN�/]��WB !�$Ekf���֦֘$*��P@
!��	�:P�7��)]",��+W;R!򤇀-Ⱥ�{q�	84�"]y6�=&!��"&�L@�EM�<��a�V�.�!�$�QE��rG8}s&}A�	�4�!�� v�A���mn�0!��"��E�"O�,B2W�&d�H[P	�CK洈�"O����=u7�����J2���C"OR�C,�;�t�!�� /��"OJ��3���OZ���A3?���2"O�hQ&��1gȔ�E�)�%z3"O�)�FH�",�Xcg	�AlI�a"O��y�J�� Ձd,�7�2�@�"O0���O�3�|��$L�!k��0�S"O�0!���T��bD�_��lYV"OL%�FM�𠘡���%d���R"O�H:pl�9���5��1Xc8l�u"O sW�F#R`H�TI��G�I�"O���LG�	!Fi�d��Q�c�"O��á�,O�p��GN���!"OZ��7-#I���j���sgn�ҧ"O�)� ��ME�R�d �T�|1��"ON+6��,>j�RAS��6�"O֝�jՔh@NĀ�b�i�Z�ZC"O�mk��u
4�0���e+,X "Ov������J��(s���"K�x�+V"OL�9�G��>��/��G����"O����&
	E�]�&%D�;��݊Q"O�{&�L�tLDЁ��ˤz��bf"O��7�̈��Iꡦ�=�Мcg"O`�j!M��ciԎU-�­	�"O(�;W�Y�JJ,$�� B����@"Öi��kر�5)מH��5"�"O~�����%�����h� ͪ"O��!�����D+@
�,��`��"ODi��E-cX�ݘ#�C
@��U��"O]@b!L�	g����R������"O��2+Z�p�Y�OM� 8K�"O��B���2sHq:ƎC%w�>�Xp"O2���bɽcH���W2|jbp"O&�B�S�lP�?mBH3 iU� �!�$��]��E{3e�j�`���7j�!�䝜K�,�w([!3�5+ag�w2!�d�2d�"�K��Fe.]K�H�7)!�$@$
��,�d�6|�u��O$p!򄓢p����Ŋ���Г���!�D�G�~���/J��A'͖�e�!��
�&Yn,���E�EՑ#MWY,!�dEr�<�ŧP�yl��˂���!�$V6r�(���P�(_���.2
�!��
z�Đqaʒ�D�4�R_7{q!���R`��#:�w�	P�!��Άg�&A�$F^� ��B�_7_!�dX�/���"��1�**ƨʭ7�!򄊞@���a�*M2t*�(�|�!�ۖF�$��ħH�����!�ğ����6"
@,�I�f����!��3X	����Ǒf!҄�#I�!�!�䏻��8�
 ��B��%i�!�d��X���9�����Z���y��)�o�@�)�NFф,���B���
�'S���0��R(��D��
�R�[	�'Oؼ�ƈr,�bs�Exdu��'u: ï�:xtq*�B
�r���A�'���q�9I��0Ӳ#�T�l�
�'�z��Ъ���Ԡ��J&P�X��'JȹPqi�.�2չ���/�E��'pT4�(�Z�d��C�Sbq"�'0���/P����aE�S	XxPPs��� aH�зB+^��ᩞ�f�RŰ�"O��B�%,|Z���v�ؘ@gڔ*E"OrXi�,�&��Ț'
��*����"O�{�V^��#�x��}��"O�Y �^�~:�R�([>�n�c�"O����4_�����Ҍ@pHDy"O��!�_�&W��1d䉁Zg$9��"Oȡ�i�>@
z�St�[1����"O�I�m�kΤA��:@��ѳ�"Oڝ�V��=JL�Z�̅&� �bt"O��笐٘���4����3"O�d0�m �.�h�*p��_ �2E*OL������9P���  �'Vf�'ڦN�R!�f��~Lt,��'�,��GMC�<��l�e�ʀh����'x!�B�r1H��(��`�	�'V�ذ��	l���$��]�
	�'܊MP��
�X�È_h� �	�'L��	`�)T�����J�:Q��9	�'�4`cB)@�pJ�x $�[�H J<��'˪XXժP+ST|���W"H����'�j��
N�7|0�8nNBjd���'�\`��UO\�d���3j~��'�� �͘ M�t��%�;(���z�'�txEb)�����T�"��!��'O�9�#W�zL!"螹e�6���'bN�Xa�GN"�`�� ߳V�4H����hO?����ޞ5~���e\$E�����Xr�<1Q�J
&���Z��T9Jꚬ3Qa�B�<1�&�&���[���]��$ Q!J@�<��ʙ�`�
��U-
,`�.�`b�M{�<��c��n����,ݹ�Bo�<����6kl!��L�6]�ya�(�l�<q��3
R�WP�"��Ō`�<	�k�	e��$cТ�T�Αa���g�<�w�[T�!h�U=� �7.^e�<���}}���J�((N�Zԣ�_�<�b�B�r�e� 
��u�G��c�<�-��.��9�ȃ f�!�%�b�<aL�
/n�5�`�qC�1HF�]�<��AY�9c�<��d�?v�,���.�A�<��^%>|�#���2�$�3 X�<A���<e#a�</Rm���V\�<���\�pU�Ʒ/�`C���[�<��YA�A��7Az���s�<�s��l�6mblB0�����`�F�<�*��w��-!�Q��HH: l�{h<f���\5Y�[����cF�y�Dw�f���Q� ��e�E똉�yRh�%IrA�u-T.q�T!��h�y���T���(a��]�~�#t��4�y��ǆ��Q�j�Z|��	����y�v,�R�N	�N�R�R��?�y��G! �&2M9�`j��=�y�+�D����P']�Fj���M�-�y�ͽITnP`�C�L ��W�y2��up󴅪1�^"�J�'����C��	�6��QCX!d����'��iRÅ� RHщCoN�bGR)��'�r�����+p�9�0W�|Ԉ�'��+�'P���� �KH�t���'�uCs���� /B#�L�A�'�h��!-�����W���*]H-��'� ;�O�e�qq�gO;o�>���� ~���s&Y� �>m��h�@"O���`�0%����/�����"O ���A��@��#¥L��1�'"OzR�Ƌ3T�љ�eKn�Є�'(��zUɄd�|-����15hdl#�'Y��{4ET
[�*�`���ţPj�<٣`P�`vH}�"K�H m II`�<ai�av�w)�7�N����N[�<'N�:�xX'��j��X�La�<!��/Z} *VOѾ�NhX�TS�<�5D �D��`��6-X�yd`P�<1��X���8���P���;&�M�<�0#�9�LSfX�!\(�%�
p�<� �4e[��͕x`I�T��k�<�e�J�x�f�;(C�ZMR ��Sc�<�t��=V���@���ʔ]�<�*��	�>=ɶ��!l�}��g�Z�<9���Bw�2���)u`�� ��q�<y�	�4k��PbB*�#[#�5���R�<I�#�9L�v�f��p��H�ĀV�<9.AVh�l9�����`e�N�<LK�{����&��=�<<�%j�r�<��l�7$>���*��E�P�r�<I��[�^��襧�6Aݖ@�ơGq�<��� ���Ċ��< pp�)��@F�<��ǈ.,l8��v/�#!�)��+
B�<��
�8@�\L��d�4p��R��L{�<�b&�,�(���jxϜQ���v�<�����q%H�p�SCs�<�5d���@�dL8 �F�Q'��o�<	�CZ"Iщ0��
N�,�#)�o�<9d@�аS &�u�i�<YK�%���Y�iA՘���GJ�<����[�FXJo�����Jk�<a��=h��Z�Ξ
P��QIP�}�<�	�==��YpHR"�v�����p�<��KD���,���
��&A�I
n�<QU�'r�⹁t�س�aF�<�ݏ%BDpلoO�x����Y�<q3��)0�p�C��>���a9T��J��-q��,
1�tN*D���r��0�|2ÉEV��V &D����ѩIk�L2WF�yy���ƨ6D�P�D�j���V��R��2D��rkV�Wut�#t`յ~��(14m1D��V-���������
:q!�d�+X�ԛWK��B�Ƥ3'l�{e!�_3J=d4��,�0��NK�[?!򤎃~FȀ@oA�U`� &�,B!!��F�e#ye�?\Q�5�3cՃ+!�Ą�qs�2��g7�QBX�P�!�8<��Yԭ��d����%t�!�B G��d�f��o	p�h��]$!�dZ�pѶ�T�:��a�f��!��D�U'�I��_d�J%�� x�!�$��E�>�I�n�D)�! pB��Q�!�\�H�5�+lr�RƆ�7lt!�D�G�j�`ҁ�
-�R���"��!���N��a�` ���@aU"\�!�!��(*�V�X���� e�	9!�$�_Z�[�ρ�a���Q6�@�K�!�D	3I���3)Ͻ3�)�f���g�!�A�l�r�XBE�,�+&��E�!�$��N!���
	�iɊ�M�h�!�� ��Z�bPZ�j���)_�fQ;U"O><��F̯~z��XDH]���EC�"O�|��&=x���8s��18�6��q"O��O\���vl�-`��P!"O0�Q�.�$K��XS,�<q�D�"O�ъ ��<��Rk�h<T��"O��  d�5R��x�鑆W�ʙh�"Ov:�TB���ai�x.�`PU"Obx���c������h�
�:A"O
��f���6zaV����"O�EA��PqО�Y�b��H+��t"O�����:젣#���y�Iq'"O�ARR�O�]M գd ޯ!	�}�%"O���$)�}�H�p�K\� ᱷ"O2h�bD��b���:G"O��'';'��Ļ�E� N$�"OB���aUgNTs@�c����"O���Q�L9b^���/M�U��"O6|8`HU�h���Tb=/�y "ODP���՞0�<�3�fËXs�}B�"O��g!��tdU��|\H��4"ODp�/�⭪�d@#*)�"O�(��@_W�x�1B^-8�.���"O(���R�^��f; �^ѣ#"O�0���n�bђ �[�=TTR�"O8���ݪ�ְr��Y�m!.�3�"O�̈��$�����dX+�Ȣ"OlI�v ߥhE�UP6��PzQ�2"O��ca�׋"�nDQTL՝a;���`"O�YZ�hV�.�h�e+֥�Y�F"O�P����܄����d�>�a�"O>��j��,xA`�CԒ����"OD$�߃g/��� ��G��%�"O>iCve˙	�����X�@��6"O�XB�/@//D�x �͆;V���j�"O&i��,�zج�1GBF<�Y$"Or��4e�.>�A����c�8��"OX
��~��0�E�'(6���"O*��%փ2��B��]9kk j"O޽b��&2�R���DB(,MdD*B"O��!��	�`)#퉷"O�qr��	z�����I4���"OL����\�/DUCa �if��"4"O�AXQ�9u��kch��*z��"O��ς=��)G�'��y� "O���MG�O��	h����Rt�!�"O�=�� �4P���:�j��"O:�'�½{�N�y)�����Y""O*��FI�P��P��.l�p�"O�1I��]����c��*���"OTx��至D~0��#IX�Aӌ�г"O��x5JLH!"!��F:VD�H�"Oֈ�ׁ�rǌd�5��^3Rbp"O�3R��Vt���Qg�9p�G"O���A��>��D�W��l!�(B"O"ŲM�At�h����1[\PW"O�uBs�V5)���U�ʵl � �t"O�`BC���Xs W�2�:Tx�"O
�[���)Gh�@� �4I���"Or�@����S�O�_��dK�"O�Ɋ��O�`��������)r3"O��ː��8Y�Љ���Jr��2�*O��g��7>/J0�ը�5!~L��'7�`�&��@>Z8��,:`V}	��� �Q��έ&ؠB���,��Ī"O<���*a������޼��"O
�2��jXۖ��^�(���"Oab�������*zy*<!e"O ����99Pĉ`�f�<v��"O2P	��D1��@�F܁N>�UK"O���v��H	�惡*�<h�"O�Sp�Cqf.�IqhPs"rɐ"O�9c֡�O���F���9d"O0l�d>I%f���@<�q"O3ϘF��{�ǸVF|G"O�2w�.Uش}1��rT84�R"O�I9�B�,�:mx��خ=�����"O:�r�cQ�))��0	�vК�)�"O"��m�0"���)[ݴ�"Oz=yg�7t��@�,�1��"OdX�t�	;���JY~�i��"O0RFD�?i�D�[�ȓ�O(	@�"O���2��"@a���(~�K�"O�`R��ÄK\�g�g����"O�t��8n�h`��%�c�FN�<��Q$ͅ�3�Еb4�?
|h��"��G�7ܶ��#N�<Yn���ȓ#=��`���>���C!�Wu>���XZl���G3�l���NԷG��\��?��=Гb��(��{�G�C~jB�3@��\"��ځvF�]�gf[*1��B�I�'"�����f��#���)��B�I�x6���Ot�q�C��v��B�Ɂ$3.dgj��+r0tW�@�b��B�I�0ᚰ��GBpa��ʶƚB�d��9X�!ԃ.����� (7(B�I�{����ٲ5Bt�а ��0B��b�ʵ�d�J�8��焗2OnC�	�����ؒ5V�	��C	8�B�	:Z�XU�C��s��y˜!\͈B�ɿn�xG�& �����n�)b�B�ɿZA�ɻr<i"4 ��-�^!�B�I�g��T���]I[��� �B�I3��u!�2['  ڱ�(8��B�Im�t�2�s�����V>h�B�/TO�(�
M%E��k5���Si�B䉎=ތP�H�4��%�o9A\�C�	�v����j3(�^A�ә D�B�	qh�As�AW7�0���/n|�B�	�[��=�sϙ��@0a�ՀL��B�I�n�Az�F
�6h���a�C䉽@hy0J	��e+s��m��B�c~�����F/d�_�ٚӨ,D�0#��/���k�bѾw�:�v 5D� �֡Y�YA^���,~8QH0c4D�\Q�Ј �N�Ҋ�
K -
e'1D�$X���J�����Q!b>��Ԧ"D�4�Dn�bh+�Q'I��I*A&!D�h��!��T�`��Pm�+�p�SN>D�HrD�F/e89���WtP�<D��x�)P5T�\㠡C+]��Uڢ�8D����j�v8��N\�1��#�7D��*� �R��K�#{��=���(D�����
�uk:�
g�	���ɀ�%��0|�B�;�bHUCP�n��Dc�l
E�<q�^`5<�A0���H!���<����Y�-҃�U��R[�ē&�'jqOl��,>_ƌ�`�y��ʇ[��
�S�? "M�2
K��l *��ӱG�0�b����>����CNV8�To�w�D�B���KD!���5Ä��j�z��`H`�ɱ\C�d3�S�O���Sf W�C�E��π[dc	�'��YAf��C��0,�/0�y��~�9�.��rd+�0,�����U>�����I�<)s�b����Z�$�E�r�<��]���[���l�:�r���l�'??�+@��4$`�`S�:�`8D�쩱��al�Q@f�H����4D�8���NtH�@�1`��8W�.D�HyE�3����$%��bF�!D����@=���Ɵ��ȴ3U�>D�P�aI�5:��%y�c�GC��ZC�/D�<11��i�X����~�R�I��"LOP��٦��%w��10��#,^4#�. D�S�+N�6`�)`ש"n���c�>D�X:�
ɋؑ:��� ��vn*D����n3�qA�g��p���34��Or�=E�Č��R�
�S0�A�����hC	��}␟h��JO�1�A��Λ!���6�%D�����
�x�r1�ǨM)<))$�>�Ԟ|�U>!G��
 =(B�Ȇg�&u.��5�y�f� ����nB_�@@�M�����p>i��.�z��^.��C7�Kf؟Dh�'������|�}@5ߘ6�F,��'>���C��dD�t�n��B(LË�&�'4�)���)s��S@���'a~�9'؄�X K�
�2Ȩ����yҀƧ[�|P�B����${�⏳�y"
�8i"��X�d�	����bM��'Hўb>�s')��wM�l�/œ\ &l0c�#D�$�#$�-J��,[VM���8!a!D���$c� 0&5�S��r�B�0� D�D�6	΢�Z�iS��)(��k2D��1$�G��X�t��r��!� e2D�tp!�E9 �6a#�P�!e���D+D��[��7>����n�+?���@$*�D=�S�'�􀠡�W/L�������c�����O�$����s��� gɨl��,�?�ӓv�l�Fɝ�q��fX�a�~=�ȓ,����@�kafD��?B�H��d������%q�9����IY�K �8��M"\::��/Ӷ1�R�Gz��'�p9��@Ļn�ư@-��lzm��(�S�$�ןr��\)$�*�X��:f!�dE0}�V�:��H9&���jdO�:`1OZ�d6�IW�S�I��E%��U,�) (���$6?Y� 5�������D��Ў���4�'�ў�>���VY�H䈂�$��o>�Ĉ��6-�hV%�,��=��@�.��O���$� r8X��F�2�ʈi��Af���`fa� V�v�u�6ϝ�Z>��+���(�yC�3t$�l���9N����ς�ē�p>�U�]�N�{�O�~*���K�K�<٦*\�h:2d�MY48��x���K�<їoĀB�|}#��9z��d��AK�<&�C�8�!�γf��CA��<q��Dz�)I�鈡qt���b�5��l��Mv�ó(���UK
-D��2S}�<1a+f�Bm8c��1E���e��@���ē{�$6�$��|�C��$N�	�ɓ%١���h�}�G�^&���S�KE���OBFz��t.�4h��)�t��9(�]4�����O.�~� �(�$=p�ԋ�B�d�F4"R"O�H�B�<!��X&Q-r�0TB�"OF��U`N4
P�Y�KCz�JP�"O��iA̙3H��J�m���#"O򨉲EE&>�z����ϧl��8ȆO\m	b�]�Pss�%��%��
Xc�<a���_#&�SRr��`k��PiX�HFy�
�Z��,��$]J��5�y�a��bA��7!���$S�p=����#�pa����R#���d��!򤎑f�"Q� }pb�фc[�ڱO��%��D���8V��HX2�ٿD�d�V'�W�<�D'E[� $�E.D�I��a��/|�<1�
ĒC�5J���6ly�hʓ(L{�<�L�*0ҡϟp�L���Jx�<ɧ(�p�d�����p���oj�<	�	 p�8m����= U� ��\�<�A���޵KE+�I &)aA�DY�<�BP _�� s��65RT���X�<YQB�X��JE3PD�v�n�<�l�>>+��($N�Ay$Y�!$ZS�<9�G�6����w��0N]��#�R�<QO�9����ߓ}A�Re<��B���O��H#�ϕ�������j���K���'����W�:к���ܾ�ļsÓ�hO\:įX�OU4�A�@�R%� ��.�Ş\e��Z"���1��0(�;��1�'�ў"}�C��0;��y:��~Mje�b�\x�<qƊL=�f�����.b1�HVn�<�e��s���#��j`��h���<�'�ўb?բ��IK�@T�fطFIl�;uc:�OF�Or���N@41!KK�NP  "Ox�*@Ö>�p"W�@���1��=�S����y�@ߪW����B%]�M#N��-�S�O�$��a�֨!��L�H�.kG�d�!�$?�	D�V���`�[�j$x�� �4;0|�'�a~�D܆%G�D�712|P�I��y�8��:� B"bYMZ�b]�y̉�u�l1��W�a(v5	Ŋ��M+���s�j����'OJ8���R� �X-��"O4���C�ztd F	P'd�M��"O��yA!�)6 D�G�	)�*����	m����'$�t�ҩ
������Q)%�$��SF��G�&;h8���	hw�n�~ܓ�~���i���[�n�09rwk\��H��''��&�,�di�֥�P���'aX���B���(��D�*,X����DVs���)�.��t�^QD�փ0=M!���{��O�ca��J��1�`��)�矐����oD�, �,΄@�
#D���`(˜6���en2�ʆ7D�����FL<�(�a��S�9�2�2D���ąB�
!`<����)ͪI*qH1D�P�pL7u��-Yf� �v]R�W0D��/�l��-�:M8�(�&A���B� +@����:tp��V�_�Ma�C�	�Y�2Q�t�
Q�5@6��'B�B�Ia�A�Ő�#���&+�7l�C�I	���i���:R��5��M&�C�I�]Ab��eM\*g��G
��8�ZB��6U��!��:v͉3j�~6B�Ɍ*�A��N$C[Xa��G&!!&B�I1&P y{t,R0q~$+�'�B�I�����#�z!��8ń*~��C�)� ��RŌ�2�"��%gkd��"O�my�c�9���h�C�v[�l"Oh�8ǁƿ�T�P"�_3F`�X�"O�u �Ɖ�p��E�M9@;���"O��ʤ�G�LF�燷q9 9g"O����[J�T�@wEr*�-0e"Of �Ó�M�>��Gگ��Q$"O�Q��D(�����g�K0���f"Ov��Ă�ic�I{a&���B��"O`�ӎ��7�H���j��y��"O�5�Q��-U*^	Y%"O~�h�d��-/X�����1���z�"O���`��5A��:TG�ȼ�K�"O�x����#G� �0@F?v��h
�"O��a+)�U��B$�x�� "O����
5���d.�*�6("�"O�����H�K*�ac�]�9��L��"O���S�Ӗi�h�Ѣ��;�V�"O,��d �Kz!�hR�K:v�9"O�*�*JVq�],u�.�!��
�y"!Ս�JY�A��Z��zCh���y򡆂L���`DMf��QS�׋�y�B�7r����� p�0���yR�VR�n��@�\�^lF�Qd�D�y��	�H0Z'œ�Q���
�,]��y���*���:Ԇ�E�L�#����y�'+x�0ٸ(�B1V�L/�y�*� l��r���w��;%&G��yb��'EB�R&Ej���)���y�,u����5$����EC̜�y2�.XL,e��=W;����C��O,Z���p�h���W�,4�6"O���!�U6}: ��3��0c�"O�}��g�+&�(�	�a�� �<3U"OL���2B�Y*�a�'b���4"O\�T�5+�D� �ڵ4��p"O�T�`ߞW�r)*���(6�<��"O�$�6�!:�`�8 �Q#��x�%"O��2Ǫ"VX��,��k����"O��[�i��;�v�ʃ`��&C����"O�T��〕\;��U��JT�Pd"Ox��J3r! 2���j9��a"O���M	RA(\�e�юlq�]	a"O@���$Y�r��2�U��z�"O(��$�K7�P��Ꞃ(″�"O�@!1?m�E��,Q�I�"Ox5�3�R&�J�h��G>r�>��"O����Χ(�.���j.y�����"On`Z���8i+��J}�Iڀ�yB@�I�Ȧ /ؚ����3�y��לs��J���r�Z�� C��y�b�8L����1kp��Si��y��VZ�X�	(̌�cC�R��y�*]B��c����j���C�l2�y�,[q�؜�f�-6y�a�HJ��y���
9�Iq7���*��0�/�4�yR� �z¬�3�b^5�%�ȁ�y�-*1`�f7�x j�掇�y��I�W�V=�M�
����1����y�.
Dܫ��Uw�T��/_�f�P�!�}�S��y�!	�<I�+s�D�����y"��:qhv%H�kk0x'À��?���~ظ�u
%UM�0��UүAM�ф�	�G�)psa�;�R`T'�M��FH� ^��$I��y��щ��9��LW�C��B�I��'�ؙ)rAJ9C!�F�� �����غt���-�F��xBd"Ot��Q�%-�6��0L̲[����$�ǿ�hp��(3}�� �g}"�P*�"���'Z3�-�5�O��y�/�]��3aᇉ!�z�hɅ�MS���v)4�a�#|O֨���S��i�M�X��	� �'ﶵ�ӫ�6d���I!07[�Љ�����2Ǻ\�ȓ9 ��r%L�L���RN
XB�=�>�ǖ�~� �f�5�'l\���C�M>`T�����F�Amt�ȓ6�ҩ���Y�k*��+r�SO�4�C��]�:h���N�l ��Y�� 4��~�\�S�$2�V���G:D���D� 6hE�ĠU� �C�O�B���LX��D[F�\�'*�
(ɱ.H��a|�̎tCF�h��mX���]9\5(��4/65�ȓz�f��rF�U8h�[Q��?�@��s�"h��:�0��䨏j�,���aj.P��To��	��W���ȓ^�r��Lښp������Rm�Q��!ܑ��*1�<)���_�4B�ȓ7�R%�ŪK&
���I)}�͆�Z
���+�[T���MܨS><���JH���숈p�nQ�o)Gy���ȓق�{"D�b�� ��O�FxΡ��h�@���%n�i����`�6N��X\��"~ΓMP� p�`�)|����L	f���
i\�x�K�
/-NPk���`�1������ؒ�Du��K�H�CD$�ҍO=��룣5lO���'�C1v{~�J�I]d,��"9K�U�4� |&=��e�2(��I4=��xB�^,R벼��P�c�	!��e��sr�i�f�B��]�!'�1�O������iO4�9�Pc�m%�y�f*X����%V�G��kaM��Gi"�bA��8-Y`�k��@��,AH�&S���O�]>dx�"��O!pCH�B�I�=5Jx���wZac  K�={���#�D'k_��(�%�6����k�� ���( �OF!ɢ% =��\:�(ͧnI����'%�����X�>�Z��K�(/�4+��fÚ�&���0N����
C���Kv�Yn��h+���7
!b�ۘL|��P�'��{:���ɳ|�.��!L� hkRɱB�؈�ݮ;#ܜ��#�4���+s�G�QhZB�	�r��l��g�1JS�-Qe#N�ǌ�y|�d�aY�aҡŘq��`���D�d�)AU�P6p}"�RB_'v���x��"��:v��i	��S/E�i�-c�1h�D�`8�^,���356~4Ӗ���h���E��''`����:a�����G�=���{�l����.,=0�I�����!Z��[�T$T��¬^�R�Iae)qE�(����"��e
5\O�P�JsN�q��B�j����Oj�P�2D�&�tcd�d�-F����,�J?T�x��B�P;�T�R&R8�
�Cs╵j�y����%.g&�[	�vN�9���`��EyB�����I�4O�L!V
 �F ���sF���~���=gx��]�e�&91�C�Wr�ڶ`�_���D[�\X&dQ���O�Q�gG��%z�]�щ)J�Ac�a��{y�Ur�G�5����4 �6"�y�7|>Yۑ)�(N�q�z���[T�W=��`���T����u�I�2����7�U�'p.�����䋈�{�Z�f��I��5�ŭ�b����狼`�, �$j�X�0�2��+u��[���HOx}�wF�2q~H����-w��2&���{`*0C'�+��� 'I.c�^����a��O���¯�M�V/ДrÈ\ �`
!O^h��g	�E�K�gN �q�FM��H�&�X��GG�i%@�C�䁮H��!Rm}p�h�6B�EK����iB��Sn-P���.v���O��T��ja��$�Z���(��y21�p����@P�F@�\@NJ�MA%*C��I�JD�u�(�T�7J�Д��GA�	Q&!���ħ�M[m�1:�+��ء����D�B��4Y��2@�[�f(T��_�B�
i���;���AV\��)(�P�c�����9X��.m�̔np�1(;����g F�*��R�"5NAk���.��1�ѫ	*[�$r��4�?�O����U�!2@YC��.��C΋B`�ԱWa�?$z�c`��!m��tƈx������f�(���� T�E�������18^Ya���[t <i�(]�g�.�ɕ�b>�*c	��Y���s��3<g.�$�:|O�9��8B��:C)U9n��'�Õ#7��+^�v��%g��h��b�>7�Ul��N�r���'�T)ps�
�k<�eR&퀕E������ğ=���r��,�'mxj���H��ԛ&��L���W!6qnŇ�	�e�:�r��S[�a��!ׂGnQV��.&��"~�I�y�� Pa	��x^��'�T�o��B�)� � ���f�L${@R�/�T܊"O\��Pj�eq����\9Q�l�c""O���F���*����[}2DA�"OQI!��2A�(�C���`�^�)�"O�yc�	T�1+�y���+,2�C"O��y��p�0��F9p�8A�"O�q*&!A�7n\ij!�>e�tK"O ly#./���H�
H\xu�4"OR���M3�Y����2y@F�xT"O^�r�(Ͳa�tD���
:�4�"O䨩���
_$9�1����~dc�"O����hX'(ې�7h�V�"O�5��)��$ �`�*��@k�"O�h�AI�!f�$�� \�k��a�"O�a J>�.Eh㏜	崵��"O�!�uN�m3�X�U�W!;
���"O6=��@��4��� w�G*k<���"OD�2�7O���6�M��rhw"O�I���E?S�=y��̙O��ժ�"OT�B�']v�(�sr���.��e�'�~�@�K��qє����n�np������t�ȓ"����*�[���Bɖ��2�F|B��0VUar���l��v	�B�������Q�!�V%r����ȡ8ऍJ6)�&u��n��1Нr�Dӧ��Ru���:�|!1��	�N8Y3��#D��ȔƆ�
�)�G�8{������<���'��ͱ�?,Oh���
`���1@�*|Q�'~R�W�^�2���R���dC��IlĠ3 �aH<y��)}�6�a으ZmT��%�Ih�'�T�3����e	�~
w�Sx�*2H�T�9�a�`(<1��+P�j���٭U\����tY ��φ�h���:e�H���	M�O4�HYBoٮZ��(��d\�P<E���'�rźF��.'��'�|�Z�@ۄ]����ȔA���)Or���� VRTQ˓P:FʖÆ,o]�2`������'��a�w(@<kK*�O�ӓ
���2գ�-Wȉ�2)V��8��N�*4���bO�Q@i�="��C&��{I���ʛE��L ���CS��6,*yR �d�i�= ���@e���ukY?g;6IRV�1�O)8 FN�S�|���М2ʞ���Ó��5[�(G��9��9��M�O�t԰�DO�j/>�
�F�^ᓊ���>{���4�T-�ħ]|��DK&2
�V��/5fU��3e��ae�҉.�XA���>�8�'%�(3��\1^D�OQ>�b�-��fʔ!1!@G�:�P�$�y��N�Yo�$�D��3�����(��'"n��F!4>�ϸ'���)�d�T�ip��;���3	�����Q(ڌ6�BY;��rS��J�K]&���@34�O:(!P�s����녱f�J`�B�'����_�\.�'��=���ׂ��Ԩ��~���:�'޾��hʧaAV��ɕh*��M���*+(�qO��ݓ�$E�xg��PLôT�����"O�K$��*�b�����$����"Oj 	�d�k/�����
�f츠"O�@i��(S�f��U-� S�"�"O�|
P癌&2H��������)��"O���f�5x�P����j� |�F"O(@Xb�^~��qs�D>�Fd��"OX���SP��:"eW,Y&�1�r"ON���eӱ}��$_�83*��"ObM��ʂqZZ�I�M��:j� �"O�� �Ө>lU) KO��xh�"O��J$�D�|4��ዃc���"O�F�5�H��AΞ??�* h�"O���a�� r��ք�n��Yr�"Ob!���5�n���I8:��pT"O�:1�H_ HLJ�C�1־��b"O� <�ci�xdj�D�=�0�R�"O,Zvɟ�2�jI�֤^�_ZY��"O�t#�MŊx�1�q�˦k܈"O�@�0�ءPb���F��r ��"O�d`W M�#Z� r��cu@P@W"OT�rʙ����Z���j���X'*O� �D�����+��CE.���'�����K��F�X
�e�1<�T�	�'�er�m%�*�9�j�:
�q	�'���a��$S�����_ &~!�'GzE(����v���"g)Ա頭Q
�'�8�r�
U�P�2��qa���R2
�'��%Q�y{�<cc�X��	�'oʙ�"/$(~�<X��A�#���A	�'1�|	�)ߠ|	�,jܫ%�$�I	�'��4Η�eJ�kq&wL����'���j�)��7�~0(�.b�ޘ��"O�%PΙ��P��A�:s�BD�""O�͙��Eu�������p<��"O�4i#��� "�0eJ�,6�)�"O ��Q�H:*z�Jq��O� �x�"O�Aq/Ӣ9�t�6�K�5��ˡ"O��[� I�&�v��%������P�"O�5[ROIJi������+Є�y.ȏf��\JS�P�c�f08� C;�y"Ș�~�L��f^�:U��Z��y)��6�HDѓ��($b�R��
�yR��i�aa��M�����y��w{�̻2��E�|�6ꓥ�y�H�=6|�p��1h|�ƦZ
�y2��#�La��C+I����*�y� b�Hdi��}�D���yrfìS����M�(��x��O��y"1��\#��&�.@"" ���y���9E��{�fB�nV������y���Z|�u����r��{�-�<�yR,��k�|	B���v���p� �y�+��!Ѫ4B��~�H�Ϛ4�y2mݣ(�$�2"H�j�`w����yb�e�LA��eֻ~F2@��(���y�Ŷ)��}�1�R���}(��� �y2fZ��L{�E����Y3�T0�y�eG�@���bj|��T���L��y�K]�,߄�:B�L�D�<܁$���yM�.m-��CQo�6:}Ĭ�$�؋�y�G�d�<�GK�L7l����y�/~7Du:V+�
��d !�Л�yb��.��(�!Y�y��}��jF�y.����s|�*-)c��+�y����BbQ p��29kā( ���yR�E����1�c3�%PJ�5�yR�*&2��q-�[�<�w��y�)V�RS�+��WXJ',Վ�y�ޠ8�i���p��1�#���y�C�8�`����أ=���b�@�y�狂rF��:6���5���҂P9�y��<m��U�R%���,F�y 9���Ό�%��|Ҁԇ�yr�Y�C��8֨��.�*k��ז�yR�N
2����G��3q��(�.�-�y��[�b�M�1�[�E�d�(��y"�M�7�������<~��MJ,�y���1*�H"�B�)
B}�r��<p�	���H�S��y2D�#V�h�s�!�q�°�y
� ,�{��=���qc\PJE�g�'���#Aڸ6a|��,H�t��T>j�A�-Y��=���ͺ+R�=�w��O���՗}ɦ\�5�Oc? ���"O� +n�5T�00"�!. 쬒���	8��3�lD��h���PI�� �����`�6:����"O�,8�T�VC4qrƀ��O����K�eRPQe3}�E!�g}�%˂r��+�B�`�4:Qb�$�y2�a9�l�-\�H1�[����o�ڄ��E��+�{�g�?#L�q�h]�F@���@��=ن��D.�=��@�O�ȩ�c��H�(�3�ș�'"r�0&"O��r�)G�Pcn`{`��N��Q�d�8Lv<�
A��h�,��抍�!��e�a�
14����"O�
 D�/u5K͞u5�$$���(R*׻��?'�>�C��Rd��?q�(�ZW�R�]
f��f|ƽx�Қ)^!�A��$��P���V�*��"�Ub�P#w/ �M�	���Ϳ�����/�0>��%g7~��;����+���!���$*1�C��=���U?=\4����'
��xS�"O	Q5��x � h��Ow�5X�"O� ��S�[y$��7�ˈv
��Zb"O`�Sf@ªs;.�h@�J��""O�E��C�t�dh����X��"Ob�HT��'�z��f*X�jHa(�"O��ۄcS�LV��㷇K:z<P"O� KViښ7e�Vކ0ؒ�"O l�$a��HeIG�TXReS&"Odl��Y����!��"oN�ܣ�cF:]�}��{��9O6,w�S.:�2l�cL�&�P("O�P�P��4m.�Ց��I�6�ȆM�O���mſ80Z����#%��l�dS�^�V9h��+x1a{��+�,SUoF۟��5i��6#�H{7���l�2�rB&D���*E�<,�r�IQ2�Ѕ�$�ɔN&dIh�oɫ6Z�>��N�D�f��Ab��c�"��6%<D���-�+�H�h�e�9I��0k��?5�z��+L�$Ax���d(:J8Y�OD�_�1���X*�!��k*��ۦBB
%LDX��Ɗx��F�Ŕz�Jx�I����%��u��*À#�L��
3lOVq �ğ��Nu
��r���䂴Q�� ��m�'k�>��ȓy���QN�#(�T)�d�\x���>Ɂ��/��iG�&�'7O�Ub3��}�x}���F�q���ȓ���e@��l������!� ]�Q��(X n �N�F��OTa��MK�TU����:_&�`�
O�����Z��\��]�lgd��Wᑐ�\x�
���Э��>��T�CTR�@��^�_�FD��	6�r��JD�%��
$�O��Χ$J����&�}�0"O�Y����'1�r�ᄶ@)��*F�O>�I��ݡ �b���<�'u�$��6%�Qɰ������t��9��$t�qn�O��dZGD
�}��޷d��԰vFL�����/��5S�FG�5f0c>)S���7d����ɘ�)�!��P׆ܦL�|��s�N,�4�G����RL��6��\�RMI}�P�J�6��Ě(n�\�s���AQp�N?��'P�����J5qJ�	��f>@8Ab�L�O����!A�n耜C�($9�v����uY��*^��I�^�x���ՔMH�1!"�~�#ܔ9��4("�I�'�B%sC�<�b4���
7����ĊԳ4s4i�é��X�Si����IO%��'l������d���5{�-�f�I�L�0�P�K�FX��2q��\Oః��Śec��#�*M+�8�uD�9}�@�6f�>Q�а�'x���'(�X�z��/7�嘖d�-�|ٛѬL�=����
ߓ��ܹ�(Ȩ/;�͠F�R(�����	z����k��=�>�R�骟��s��Z ��1�T�MU�'>�@�3nr�P�r�W��\p�f�.JVt�Q���ʏ9�
�PE���=ح���Y�S�`(T�G�ן
� ���FUv�{FB��||j剐�O�$�2\1"���*`�F��i3SH�W�H� �b�RV�j�x-�a��pD"]>Aʕ��m�9B�O��	�+�6X&D���3bȼ�3����Y��´��>�$d5�����4lZ`M�ClI˟XӠ����U���8����,Ov��IF�Z
t��J���8ţr.N5d��{��=)��HsVƸ[����ý (���,O�u�,tQ��Ȋ;�@�Q�+�'.H��)� ��٬	�e��듇TT0���
g4j$	FBs�O�>XF)�s���S �'�H��'�Xĉ�P�8�8��'�t�8֪Ŝh̓�{���'`�	A�D;N�v��B#�<j��x[�'�XM1V ރo��8Pb`^�|zՉ�'�\���<����A���I+�'b\���ɗq�^U�����'��MҠjC-"?�L�c�S=D�%0�'�����*]V��r/�0�0q��'e��c�T�h��I��d�)P����'�:|[��*������LP�'�d!�BO����Fˊr��)
�'(�����l�$�W(j�&�	�'��ըD
����!K�� c�:`b	�'*�\�!�?'Ǣ1�4^غ�	�'Bڽ:�n4�P	d
Qj�8	�'���
�E�r0$��KIF~��'g*����8N����*�
B�h��'��5 ��m_�,8����i�R��	�'Ƅ�p��J�((�LQ�<��I��'_J���%ͰY.����P�|Yq�'|����/F/D�<)�3䊗I�z,��'�Je����MY�d(D�ۍF�r�'�م
Ns��x�`˴��I��tP�Qx�FW R�H�*w+;SN`ZueI�-��B�I�X!�#�MW5==6 ( fK���">�1��!r�ᢎ�d_�ERVxS��(��ș�� �y��4�x����E(\�t�(��
�?	+W�;JP��o'}��	
v�����+0 "�K���!��C�	,H�b� (��Xd0ʈ^G�˓U�n���`* v|��Ă�+FY�#l
��X�	��ýQ��}�D�T�4��A�C����bI�0r�Lq"݃S��4��KD��E�&Z�R��/�$@.�D{�b�T��Q��)s�'*<�lK%(
�/��I9��n� �b���� $����Iʸk��D���Xt�y"+�X����N��D����V�¡��j��{hr�P�ЛaxNM�T�^�S��|�MWn����"*.����	=��D���@��p����<��#�4kXӇC
����zy_6/Nh���^��?���'G�Y9�Y����&t�QYW`�+N 9�K5YY!�d�!y���CE��U�$���	�^�O�%��	�#��*��O�y�,$��0FIr%(��jbDq�ϖ�8���ӱ L1K `D�5'���E���^��E�H�AS��[�x➤E���צ�8�S��	f���Oյ��O&0�$o��I*�M|z��O�`�x0P2,�)�P�[�^�<��Y�N�ȁgF�Pkb��t��Tyb�ǟ�Z���Sm��S�i�$����V�+ -J�]�\��B�	&��0ӉJ�MA����aZX�pI�D�c�B�'�*�%?�(
�cސd�����ItX�1�M?�O�!"��^)H�Qb��R�%�<��c8COȉ�������?�$ܕput43��7$�	���p�����;��%��y�eRd:��[@)�Q5��� "D�Qb�̜R��;�NA-:��x��%}bF�7Xp\�=�:I�������ٽeE��D_Y�<��dJ�E����G�N�m�*@B�,Lr�<�s-ߊ��eHV�-.R.�����a�<����%<��ЦAT(�R��v�X�<A�! �}[��;#e֨l��SJPX�<�w��n�� *@�Qʃ!c�<��iá�%f^�8|"	ЧD�-&4$B�I�h�tĺu@�< \F��w��K.LB�I�j6ꔊ��B��Qa�aʴ5�B�I�7\\e�󣊒 Ɇݒ��H&$��B�	�Q�:�)xl��4H�5`s�C�I�iM�ȸ�d
 ̤��w��@��B�)� l�#$J5%(Z����>\�9�"O���c���el씁�FI�UЊ,RR"O���SJ�bjp���.�+"O�͘W�$T����^!!'�\�W"O�@Y��8n��eڠJg*��@"OT��F).@�OjŒ�"O���!�9A���J
M%"O����VY�މ8�kӸ*�����"O��c�	c������7��93'"O�DX�	H�y��Y�ȿewr���"Op��c���6Y>���OV8-""O�<h��H�J9�ě���5H�,X�"O�?����bhĮC�� C"OVt�V��r� �@R(�x��	��"OBy��)+���[��dX�e"O�"��n�$�Ó�@���]b�"O4]�3酆h��Da�怜U�D�K%"O��Q��,4�A�B�,����"O��ڐ"�D�TZw��+q�ҭ��"OXM�Uo܏d�F�i�;x*lC�"OzEcG(A jlX�f�9a�Hq"O|)֣RH�&�s$EV&Q�Ip"O�$"���>=���ㅅ�)H��[5"O�q
Ƙ˨�SF@�<��B"O��U�RfT�ņ����f"O� xrʘ	=�"PJ#c���� �&"O�Ǌ#��a�D5�b9�P"O�y��C9}n��Pd�_>~��3�"OԵ+ÉֳeG�%Zơ�*GQ$(
b"O����I�. ����_�F_���"O�԰ +UGh�J�W�Y�U+"O���h�$j���D��G���"O����ܜn�X1�B 7(��qi�"Oʰ�DK�e�.y\ �@���y��q?&ec%�qƢ"�ć+�y�"�������1gpBd��yB�ǉ[R�;��V�P���i��� �yNʇ>�8xPo���ea��͕�y�@H  �(���O��1��`����O�=����t�¥B��q[����"Of���I<Zk||+���)t#HT�p"O����(Ȏ{��)�"%_tj1"O�Ir�����P�fX/>`!"O�qQ�#w�R�����1"O�퀖�����g��K,)$�'J͢��i�kq�
�*��d�C��-|A)�{r��?��O�O�.���5Q{`�2���*�
 ɒ}� Ԧ����* �,�ɘ�Qz�9OR�ğ z� ����$�4 Q� V�왫�`�zL�'r�<�z�@�fŴ'f�H��#�{�05�%��$n�'��e�S�O3t��p�+Q�Q�0���Y�
ѪM<�rA~��E�O�F�q���<0U��k�X�L)��O慈��_z��&�"}�D��I��E�θO �#"�ۤM��l�ܴ"����Oa�� Z�2���F�j�x�#D�u��"�h޾���V�@G��Z�9�Z��@�	`� �z�n�<Ϩ���'ռ��+.'��K|���͙22�d��	7�r�aa�_"UiqOⴸ��*�(O���)|��Aeh�	[4쉀�Ggۖ�ҧ�]�$��M�n>ɫ�*��� ��~��hP!�<j����k��2��6�B�( �~�H?�X �@���f���6�Ƒ�a�	�aͮ���&���a�4#��u���3i �u ����L؇2����'��ч�7e�<褟b?	B���v��kpB��D�X��3b�>�7�ö!bע���zөJ��aH�Y/\��M�7�(59��Z�ǂ���b��M���ӣ��4��@o�����ۚOu�y���F	�l���J�|��	>'6H����)�d)��i(�r �+~Ҋ�ʂ�A���'��Ʌ%�4�ϸ'q�E
�,O���Gks�J�.�yrdI��(��!i�H8�����y
� V�8r�F?Yr�=G�@�5���v"O	�X�!A|�0G¹bv4(�"O�S�P#[2p���_=B`x�Qd"O�;!��i�� �%��"(�0KF"O��kJ�=a� 9��@�v,!�%"ONl����;��)Ⲯ�!`	t�sf"OX���D\F?�US�B��l����"O������D�V���盤�l�x�"O���e�����z� &�(3"O��(0 O��f�) ��V�2��4"O-+
G� (�Aw
Z�]�}�Q"O��h���F��hh_;P�В"Ofi0T��(k�(��T'�uK�A2�"O���!a� |����猁	Z�-A�"O������]����åU9f�{�"OT��BB�F�֡:�F��]�2	�"O|y"T�Y's!���&�L+��4"O�E��nDM=x�abc_��-�"O�0��-]}P1����C��j5"Ol]�u�A�q�X���]�N���k�"OX=�F��C�3w㛿4����"OrL��P2-��D�`�;�,T�a"O��&f� bf��A 8G��k@"O�y�Ղ[/y� Y0D��}�h��B"OT� ��:�"r�C��Ph�"O�3'� c�����ԋ
⪍�"O�D�� Ʊ\>�S`�=پ�"O�D8���$e��7�)&�$�h&"O
���D��������{E�ڇ"OJ�(�a��'	�D�0,ש4$C"O��v���8�c'KZ�3�j��#"O��f؞?K�C��D֚@�A"OB�ȍ2.�tp�
� 2��y�"O�e�kDn�!������(!6"O�u*Fa�/��y��S�a���7"O���`�8@�6�E%����"O�@PB�7;���l؀l��I �"O�!bv��.j�4�2k�"d�c"O�q9�-Fc0I�1/\��9g"O�a�I�[�Ќ+�#I�1� ��"O\)f Ha�];4�ϓ ��m�"Ol|Q�ʉ%���%��Rx�m�"O:���Y�#Z���S�a�!J�"O"�P�k� �&�[�+Y�ZH(E�"O�g� �������2�a "O�9��X�Iô�P����6=v@ȡ"O(=+����Q`D507]�q"OP|��h�PyV�eh͐3�]k�"O����'R�D��d�t���'(�Q�"O�����:V���@#F�7i���#"O(0Ȱhտ/��k�[�l�����"Oܠ��*Q�R^؀�D:A$��#"O�ar��B;{��!�e�<��9�"Ob�1�h';�<Y����C\4ia"ORY��N�\�8��ۙuT��E"O"�B֩������Z���mkF"O���+&����%U�+��]y�"O�	k�3�M#���'j�=q"O��3v���ts4��$qefm�W"OP�h�)�,b"DpE�:VG�y�"O t{-���%�Ҡ�m�
h�u"Oz��V%*z���J�$p�>9j"Oz��쐺A�2���h�5X#N��!"Oba�ƋS"3�b��GH׽r���"O� f1��%(��1��E(� !�"O�䚐�ьr��	gƷO��AQ"O�2 �$
�$�IĈ�,��"O��Ď$F��q֡C�
3�c "O.�tJ�a 0RKP v��Xe"OF]�q*/O�e�@��̉�"O��k����ǆ�9�(ehE"O�$J�`1[�t��g���3�赃T"OX(��h��Z�H\��A�.�*<�"O���p�āشYH�]�J�1R"OƬ	M�!%Tqᑋ��s�"O�"�K�{根���W!\rJ��r"O��#��̶(sj)�%G�mf���"O�����0�pad�ܰXR2���"Oڄ1�`�Qk�tTکZ�8"Ot�h��I�,���x�̉btT��"Or�C��B�g���У�"mI�3"O��%�1�i�P"�zl���"O���WH���yJ�k�[O$H�0"O��S�.ςn��p�!I*���"O��"��E�/��I�q@�8D�`ڴ"OJ��w���u(e@�#M*�Q0"O2{B�G[�"���S��M`�"O�� ���C�\|k�-��9 �"Ob��%+�*i3&�I��D��ڔQ"O��ȅ�*mlq爞�\� ��C"O����. �#J���XA[�"O���*�+��qóe%c*V���"OdU6*׎N��i�6"�c<tm1"O0�ш�hM�8�U�׬'PZ�"O���ŋo!�0pbD����zP"O�C��}����p�߹r׸Y�"O���׌ͰL3�����b��h"Of	�A�W�G�������!]y�|K�"O��Q�΀#oj�Y̜҇�] �zD"O�����5�f��w+�'r�4�iW"O0՛�	G��(\�f� @��8�"ObuSQ��W�Ĩ̀Kb}S�"Or��!�y��	2��(Z�5��"Oµh"}�꠩#c]V�6-��"O�8�厅'A��`�Á���0u"O��ЈI�Qov�҅����S�"O����g9V���4ċ�.2����"OD١e�1l<v9���D%%^�;"O���i�!�*��$̯,3��:"OBգ����8y@$;	v 5SD"O�JG�?%/�B��2N9��J!"O �h�$Xj�� �ee��K��1�0"Oh{Ah�4t�0E��B�vH<��s"O"���5��욳��'�����"O�+��#c(�9�s�̝C�`�B�"On�P�Ϫ����B�k�d)r"OB�3���3���X���&hȠ�"O�Aa�a<Xv�ie��m�]��"Odd �εTM�ठ8B9Ѐ�"Ora��/�й���X)���7"O��ӵ�I�a�X���Ɔ]R�x�"O�̙�d�f62�%D�@z���s"OJ�s�� �Y��aI�֯Ex̵�a"O6D��P�b}�l9�͙wԸX�"OVS�O�!�R�1�f��(��L��"O:i��䙅�4��c�Q�}�VMC�"O�˥L���J�f[;ou64Q�"O�(�p-Β]�<ԅ;t}
<S�"O� �S6gN�Q�^X�e�M�(X�"O��1r�8^���w�n&
���"O�X�$Bd����?wA�d�R"O��ի�Ss��	��E0 O�`��"OX��jG%���\�B��h�"O���4+��d�dQb� ��_tl8�"O>L�$N6cl�Cs��1܈�"O���5L�.@���鲍K ���)�"OH	Z`n�cX.�[�ꀆ`-�B�"O��M�uj�Đ�β1����"O@e�%��j�>4*dF
i\��7"O�B�a��j��t����e�L�Q"O0 FL����+eC_=%k|\��"O��P�lO0"�5 #� �h	 `"O�dA+F�x��4�VT�"O�ycl��C�a ��3�b��"O��ڵ�J�3`�E@��-C���"Of9��G��<����=G"A�G"O�8�Pϝ� ��ipn�F�|�a""O�`�Ua���@C̈́��8��"Ob0�j
(5[F����(s��Z
�'%>�ys�٩j�A�?0��Yx�'���R$^��05�L�YsP���'s�t�G�� N�6�w��XRn�y�'��|c3�4b����0�\�XɸH[�'P�m[D �$T� ���[W�D=��'+��؇'�A�xY�ʜQ���#�'Jmf�[��=R���>��Q�	�'{Z�c^'W���:QǼd
$(X
�'Q,А�ٚ��A�ȡbO�2�'R
C��5W��iK! D`�8��
�'J��@���$Hh����H��P��'&��A�Q7 �pm�s;���
�'Ƽٸd�1}L���(M�`�fY�	�'����� ݜj�R�駍� Y"�Pz�'&4L����/"դ�W�[+X��y��͕9!��h�O\r��Y �D�yR.ّ\�� .Ykh�Hx�Y8�y"k�z��C�Ů`�l��AiĊ�y�[*>L0Ѕb�Y��\S!ė��y/J�1�d�a��~ڐ,�@���yR��vЩ��Yc�(������y2mOOL	{4�9_���PM�y�N�,���3�㚼^x
����yZX��`
�� \
҆l�I��I�'1fy�r�&1[����Nx!Zy�'���5�O���ehr&�e	h���'�x2Ô�/��uoE�nS ��'�|l�!���A,Q���:n��p�'_ذ�c��n�xw� f�l�
�'������,JX��q!�X֮�{	�'O��:�GY�g��*q��b0\ĳ�'آM@�L��Sp��7�V혴+�'}t5���[�ɜLi��m1��'ղ�G�1d�����!gꌱ�'�¸G"��'H:����Y�>�i�'caK��ͧ3/2���+y2X��'��!G.�R����u�΀_���A�'��R��)g<2a�	O܀��'M^]��(� z�zYSw�\=@�0��'�B`���M�"�G�;D��b�'q�%��H�{�IA�b��.�Ȑ��'�p9Y�ê��%� �̉qP��'rհ1g��!q@�7��%]��p��� Ψp�陀�9��LK;�N@��"O�%�S�4Ejm0P�_%Qc�@"�"O�i���B"S�����&>T"D[�"O���5   �P   �
  �  X  �!  �(  1  Y7  �=  �C  1J  sP  �V  	]  Qc  �i  �o  v  ^|  j�   `� u�	����Zv)C�'ll\�0�Ez+�'N�Dl���32O$����' �
�eřq��退툅f�P��r�ޖ)�xR�h��

��@еh*���c�Q*w�W�?%��l��?�C�NǐM��8�M�Du>!Q��]�oy$`��l�=s.�ە���+b�Y�$����u�B�7~v���'@jG
���2 ����33X���X!c�\X1��O̔��lJ>�r���$Z��e����՟\�IݟT�IşxA"K*��8��
V�pՓ�#�џ��I��M#!�����O���e��b�dj����M�3dv�����L�\�5j�O��˴�<y�w�����'jLM���<��'	E<�1���]� �����O�x����/��M�bfˁG����X5�ș`"HP���F�'����\t"��ʟf���(X�1ɲCM>oB!$�'i��''��'�"�'�BQ>�ϻ#����e��IN6l�5J�r��I�M#a�iv7�Z��}�	��M�#HɆ�����b�ˠ42��ciC1o(xYn��E��"=����+�"��#�´o�<-�ح��+��L9�g!�/H�V�o	�MK��i5�4���r�R�\1����D�z���9�/^���)�'PN��M��#(� �5�"B��`�F:zP�e2�h�Vo �M�B�MV����=zF��H�OV���0``nט�n�c�i��7-U��Q��kL�{2�Q�PeG�T�:�s���4�V�	�` #iڌ�E��/R���9�i�' ��2�H��M;`�i��7���yv$�!|̎\�d��F��a�� U,C�-Bt�-�|P����I0B�k�E�\�y�����$��v	dȓѮM�)�L�B5b�i���D6�	ߟH�I��^���4��i"C��1�.��<e�U��O"U���	���ͧ����|�����&�ǟ���Hg��t)]�ZI�T�A�L30�ܼx���ٕM����m�	@��i��̃����v/�2	��xp��$��2U��'@(�g���@�6z��p"o̵o-�@�	�0��K�S�'�yb����N�I��5��T?��'�ў�S��M���ϐ9��ۢ
*7.h隒��6���DR�A��⟴�'��$c I�/N�=�D�p�]�ȓ&hm�N��N�-m�(6�� ��'?����w�~<���0��#�'�t%�#�4s8M� ��y�Ա�'�����i�6Fr�@a�4[����'�"H��FU�#cr��k��L�!
����Gx��I�2��L�c���!7li��P�\C�	($�b��E���f�6 ۺj� C��l��;1�T�v|*���Pz�C�<r�j$�KӳVɢ�����<��C��
;��O�Py�,���C�&tcؘ!�FI��t��n��:���Qo�ky��'j2W�`�O�	&�|q���_/d��+�A	y�<<2Qd(l��Q V�uxaz�� ��X�!M�/sa�p���N��Q��&�>)3���-��@���-�ў�[�̰
Q�B��[.V��D@M�M����F����ī<��Ov#eM�<n$5���~Sd�+3�'��y��A)n�.�;�O��1�eJ�b2�c�V���uߴ���0�o�ן�͓PE��]�t���/��/&���eyR�'��5�^�4�S�	�����4)r(\%KZ��J/2�]��
�7Wax�E��Y���/9N�L��5����īL9p���#լ��|��- ;� GyB�	2�?�ֳiu�7m�O��P�e�I�x�PN��T��Yar�<�����(�̰ؕ�3hm�dx!k�:G8�f���O$�}j��i���y�;����TH�c-���&|Ӛ�Of �q-��Fp�㟸��0,�@��\\p&E��,K
:~b8��"\��1GE0@	�i�� ryd D�<zQJZ�/�`���]�Z0z�a<D��:p��-W�����d\���R�6D����8E�<R�$ͱ57����$4D�`"@D�s� $[�-Μ]_*4�'
���$���a���?��IğD�	Ky"������.�	zU5ZC�B�YwjyQ�IQ�v�B�:0��	vU>�GxRJ��AM�1  $�:�~A ����\I0��U�37 ����T~J��ԭY�gn����l>(\�cC��+̌i���^��^ ��42��-�L��%��OT���OhhP1�[�1H�X�h�-�tmX#.<OJ�?�v(��r��$L4:�B7�ןX����M��i�ɧ��O��	yj�٪5䍉i�|*��= 0X1���-�M��?�����%��J%��E{�ޞ1cƴ�tJY�cN����խ.&mYa@@0y�Z��ܖ'��h�f�Aq L�;i�6��/̖F�sgV0�TlnڮH�2Q��剅��$2���Rr4�a�'�;�� � �OD�ncy��'O��'���'����Wl�};��$r�(�p�Z4b����7�I�<v��
"�Z�g�I	�b�W�~�O��n��'�T}�U�u�`��O��4c#�������S�XBń�O���E���$�O(�Ӳ!�r��-�)� ^@��-�kIR�;&��gdV�:#�'^��j��d�6]�]Q �_�{Wp5;�GG&!8ax�h��?�'�|��5���Ҩs*� F���y�#\*�DȢG��fJ��P����?�v�'��Po��+�p�rE���eL�K>�vj��aM���'TRQ>�c�gߟPX�+$y���':Z��ծ�ޟ��I+[R���m�S�L���@	�9I�:0e�OA�Bu�!K,?Y�L�F�����+�G'���V 3v�ŠԔ�$����O��'�"|r'&�.x�`a��,��"�N�<Q"�B�l�$02���?*V,j�v�'L�}uᛙ/�x�Ӳc�8W
Y�B��M���?�:��9�w%�7�?��?!��y��Y���G��\b}���_��t����?��[�+��q�,�Q��B�*ߓΎ�r���)���C+�3T��H�O��h��cf1�1O(1���y{.��r�΅t.��c�r�p�n�ޟ��c!˟h�T��,O���OC�$��l6.�<���8]h@�$�-V7�㟴��w�'i��O��uKxq8�J���.����?�@[��'k�O2X��Z����(���(=9�\8�#Y�Q����a˟��	͟��	��u�'�R�'��� �!�&!�0!IC�`�Ś�-��%�R�aE��T��tp��'�1)!�Hj�S��]� ���Gc�L�����̔x���	Y���CgACx�'2�㧯��P��|T���Q�:��#	7�?IP�i��b�$��l�'B�XJnßJis�*��-�������?�L~��y�		`���,�?{F�H;�D&��D�O�n�ٟ��'9�%lw���d�O�`���I�D�JD���&yDt��`�O���P�e�F���O����r�ҕXJ�&���"�`�e�p+üQ�f�����0�hA��%-OdK�-��vfH��/�9��m�=�]k���V�{��u]�ƒ(FQ��j� �Oz���ʦ)�	�e<��v�/�فE*oE��?q��O|1O��
Cf��u��MV���$��œ[���	ݟt�?�ON&�$��V`T��6�#Y�U�TO�7o
�Q�X�� Q��M��?9����(���?Y���a�6	�Cl��*��+�Ŷ�?�6�HH����>9t è�b���g���ȉdHS~��?�O>��`�H�B��A2_��H���3?yG$�hH>E�t� ��r�ߖ��yYҷ�yB���*�^�+����B`�"k4��OTD�4-Y�x>� ���Pzi9����WћF�|B)me���'��'U�	�h:r zn�6���,G6"x����l���)��l؂Ŏo���d7x��� �H�GI�P���`Ll}d�$X`9���yR`F�~� �?b]�L�IS�F��d�F��%���$T���gy��w�����8�,}���F��К��'&~p��D���#<Y�-�(�Ÿ�-W��A�ȅ矌��3��į<��������d�$Ѐ[�B��9��yj��N�D$��S#�������P��`yV>��'1�xX���q/l=��/O���Z�(��Ĺ��I�q^v�ytk��x~�a�&%r�0�$���t�摠��Z�r�Q�d�Nj�'�]�t��o0��נW�m�d ��N2�?)��3���'�����?)A�φ1���f�=_��Y�#����D:��ǘ'ba�fK�=��e!%N�!Tb��O>R��!7s��W���d��uG�'���̲p��uRwB�7\�pb�`B;j��Y�D��ßL�ɣ]���/ʍ6Ԓ��CH�<�!۩?��E��:��G��p����f�1*׌�؇�ҥnH͈�0tM�e��I�	����BO#ZbV�F��N �?�v�i{��'Ǣ�
6���Z��D�i]&\�b�'B�'O��'��OV1O�h��*G;>�TЖbPCD�x�5��.��|b��'���C�YV�d�G��*�H�����:qH�l�b���|��4�?����r�pCë�7�(M��oŜ�?���<�@`���c�VX�G��?�����#>��	�G`��K�>s�I� EX�IP>�+��ʚ�(����,+h��x�DEh�U�tg�\~Ү���?�S�i�6M�Oj"|RQ�3Q*� �lG:��
�+J[�I��t��Z����=Z�D�i���f�P�)dl��hO\�d��u��4��UM�|�B��&�F����h3�����WkґY���(O,t��<?�P���e@!�:��&"O���q�\�OV d�w�� �Dk"O,�&Ƽ~��-�7�J�~D h�"On�rM	"ZJ� &!u��	�"OB�	�+w�L�%��v��p��"OX@�1�V�ԁ�S%�Xp�T�Ш�/�O��Y0.�Oa�13��� �uY�"O� $�JD��B|(DT�Ϛy�@"O�ze�^2-�Hh�P"ƺ���G"O�Qc�	ݠ��Kw��b��s"OP�����tɚ���oB�?�J�7�']���'~>XR��Z&U�bM��_�h)q�'k(Ajw+�	�>���%l�аJ�'g8�����( _��2�ß_����'x|�y��U�s4�M1' d��'G�eH�ȟ��軴���p4.Ƞ�'5�X���X�(I���a��1���ą�W�Q?��
4$�h����Br@� 9D�زPk�'F�,�Ҩ��?��q�:D����i��R�����	�!^�9Ԏ7D�\JrG�f ~��0+Ȭ[��3�B8D�Dbf`�8�ґ{w
�$Q"�ل 3D�l*A'I�@U2����!:
<�Dg�Ol���)�$W���">E�,��bk��Qq`-�	�'���B7���b�����JME�	�'Q���f����4D�!�L�	�':^��$�7�U�\U$%x�'of�p�H�"e(smK<O��y��'���X�Aߔc_| ��x�Z�a.Op�
��'*�$���^_�1[��'2�i�'�*h�6��,L/QI���{T��'�b!���,E������/�xi�'`(�j��	A���Q8Bx��	�'��؀U(�"��YA3��6+��Ā
�T`9�3���Ȧ`@���p����3�t����Y�� ɱ
J�Y�(V�r�����ȱ�2&�d�X�EV�ܾ��ȓnR9BĆ44��T�%�3���ȓaڞ��я�2��u�"/�1\��5�ȓw'V� �K�,U��H/&}��G{� 6�����I	��D[��i2eC	�T�1�"O�`��"��-��
�cԹ.��t�"O	�քL�n�u�T��8;���`�"OrT��+� ��]Cb$H(���"O�=�D�X�n�*jVCV�{����"O���L8%�j̹�b��m�<�ȕ�'q6y����#9U��r#X�t�j��
�1��Յ�U����e��;��˶䖅/ez�ȓG��)`@�Z�
�*�� ���Z���5��[�G�d�n� �C��]�l��d4d	A+� �9@���Jv*$�ȓ/P\!�C��j˸i�L�|8(H�'�T�	�k<1E���5o�UQ�l�{��y�ȓm^�LS�n��8���0��}{�ԅ��T�!G�V�3���0b�Z��Ѕ�\庅h��F�PՊu/B�FP"��ȓnVrHR����;��]���raƕ��	��8�	�&	j�cjK(�����Cs�B��) H<�u*��l�΄��F?�rC�	�y[,p�j�N��(Q�Ϡ2�`C�ݤ�+4m^�w����M�+a^C�ɖIIBU dذa�j�G�X30C�I� N�d�9EF����T�=�#�Wy�O�ԉ�/҆nj6t��mZ�Fl�'�����э��Mt.mS�"O�,s�D"$܈aąi���'"OΕ�䬚���bԆ@,Y�޸��"O^!�"ȅ�HYRՂ\3�
�f"Oz�§����<9���m�8s�'���p���e� ��r�N���0��E�a��h�ȓ\�n2���H#�)�ƛ�F����S�? �b�ϯS���3�͘V�Zhpw"O��K��"i�ܓ��P�c�Q"OR��6�\3S��-h���`!c!"Ov�we��9�
�N�2p�t��FZ��ЗC$�O� ��E�SQ���歁�4�Vٕ"OH�0��6w�Yy�
�!>s�Q4"ONY� �����E#X�T<�P`"O�� �Y]�i[�l��6\�"O����OJ�� i�S&�R{^���'���j�'�r�:��T�١��9v.�q�'޵�e�]	͜U�A�Z9R ���'���R��s�L��#Ő(vv<�t"O�q���?	/��a1�3=gb�)#"OHD�4��6p�M�e�@�u2j�"O�q�v�}�Y	Q!�48��0�e�I>
#B�~�n
$H��a[�P �	z��b�<��j��*{�$W�:�^��Tj�<1`M�����"N�X�.�N�<)��m���s1jؖ:P�á@J�<��
C44 ��0i�[aU3�$�D�<���$��"�H�Dbhq��I����b#�S�O��aH���Jl40E�І,C�Y;�"O̘���[�%9�s�L�:4�S2"O�����H�#8̐��ʶ%|��C"O�q�)D>5�H����Cj��i�"O%c� �BN�m	��J#_�l��"Od�����]���Y�$R�x�]���T�"�Otٓ�d���Cc«UОx�4"OD�A��IlӶ(�F����"O�����ͯq��$#�E�(l	ja"O�T*Vi�\��<h₄�H��ܑ�"O���h�`\�X�O(<�&�u�'G��K�'h�U{�K2* �'��M
�j�'Q�C��& ��VDE6dH�'#�l��3/�2��E$�>��i"
�'�Y���O��ܺ�� 87:��
�'��2�Y�yI�W7@u�U�	�'6�yv/�,G����s���7��̠��dY�H�Q?Uh�F�`(\�g�K�~�ۂ�?D�8�`E���)���E�a0B�k+D�`�s���dy��e_�-3��f�.D�3�g�?@�Z���"�<i$�I�	.D��H��X:vQH�&I	���(��,D�<ʗE��s6=���œ8���s �O
���)�'=X�8i�׽�6ds@mN%"��1h�'2$�1cc�3�J��gJ��e֦D8
�'~����LTDF��gM*J���	�'��qx�d�)'|#�I�l�jE2	�'�fԢrK#utV�A#�������'R��*al@*P���hs�6MV|$�/O��Q��'��x#�&ӚNѠ͸��Z+L�Bt��'%X�Ar!љQa4��G�[����'�x�"3�Ȇ	<F��WG�'!��b�'���.P�NY��+���p�����'0`�5`ߩ_2ܩɖ���\Dm��#庐��qx���"Y�L��Y#3���[��$�ȓ'����`ҡX`���Q�ԝ�ȓ4����DD�a�43�U���������9�rYS/Ͽzn��ȓ<������t���Ґ��\P����>�H�iC���ej!����<E{k����@K?p�D]����=���G"O����&<�̤x%���*�ZIa"O�$����@\B�2�V�q^��"O� "����ܵY 2��4@Q�R�za"O���W!R�3,�R��҆NQ���"O 4�îK\�\�c��=���"�'D�:����U�U�R��:[F��	8NɅȓ
�4��ޱzp��JPM�<-1衅ȓ2���թHU6=q�:��M�ȓu��Ɨ�n3�U 'W2jm�Մ�Z�q��lȽOmJt[�
_��@�ȓ0N�6BdG*��X�t���'�n�R�r�¸�v�G�r*|�
RϚy��ȓ:�zA�SdX�nE6ț@�c� M�ȓ,�+��u�젛Cl��	������H܂>4ĥ ۗU�^ć� �^1ya�H7T����ƍC�dJ�����+�x��zʬ!��%LRQ(y�eHM�1�nB�	�{�%P�F3;]V1����oSB�	B���S�~D܈3Ea�;=��C䉷a����1O� �D��v��B�	�-�LY��bUdb���Ť"�xB�^neC�J�!�t��f���P�=���[h�O��H�6�*G~DE�WH�g�=�ʓT���"���MV���h� :�E�ȓ%���2��p��C��Z�y@<��,��Ɓ�b���b�kʁZ<X�ȓv�u��>!P�	 �D�p�-�ȓR�Qԉˏ'���S�G?bZ��ɪ?bF#<E�DŅ�W���& PEpF��1`��I�!�D�/D�2yC1��	u�u�,�d"O���GL@3��h:�h��Z�B�
@"OT��pn,n�>-Kê��%�`��"OT,b�B�,:z����)'޹�TOP�3�#U�șh��b���t��O�1��U���o٦�+4㝽(>�dNϺk��Z�aJ-b�����ʸ6�t��Ù/�?�֦ި�?����?a��G�^6J�Ǝ+������i�.�tr%�; P��.����O�1CG��-b�r�*�%(WcW�~:xX�̈�l@��Y&���1��9�)���(O��ɦ�'r�0bU#N4e,pi�ʹX�Խ�$V� ��ɂm��es���ܹ��g��v�Ol�=�'��8-x��x��)��T�@̘8�@��H�HGN����P���*r��)Mhx��U�U.p@)��n�D�[!Ʉ�g&>�Ƨ�l���ȓ?��m���Q�hDv�%�ӓ-6B�,;P�yc�N�0p���kɃu��B�I1�4pV Jd�=qe�̋ui�B䉴HGN`���M*|<U���L(I��p��	}��~��
�]8�:�H�7M�*�����y��5
hAr�U6K�.sj�'�yg(#c�ey�Dף7����!b�)�Py�\ ~��zG!?'��x+��Ij�<�qL��`I���(n���y�%D�|�Ԃ�;tM�Th'+�7���#q$�OfA� �'M��h�KX^�Mzoū�`��'d�ɚmI�����b�	s� Z�'��0�ve�Su����3T�\B�'���4C^i=�#�˝� ���'ty⠥�8I>V�1�8"�(��ߓgp|�Oh�B�ǟ)c�l�#!�6��p�e"O\e[áI2D����À�A��f"O��k�FB�� ��@�ո���9�"O�Y��Y�X)H� �W��a�"O*1��&t�͓r�i��QҔ"Oz<�r�Y/RT�%c�M�� @�e�$ʻwC��O�6T�Z�~]j�V5{�����'��qq�㖟�b�S(�)b�d�'�H@Y� ϡ�|��'cV�aj�Q��� D��B�ͫ�ț�E�"pȂ��"O����暈Zߘ�d��<�L��"O��@��԰A.�2�c��!S:M@gP��O�}�`��a` j����� þ���`�4Zb��I9`�s�ԙrr�Ԅȓ,O� �f�Ձm�:��c�E�s� p���>Q�P��L2T$J�Ղ�!�V�E�ҵ��bL�H&��&W 	!�d�j	��Tǜ�KӦla��.G�b �p?)3iDm���!�%�,f��yt�c�<	v��a�jwcO+$�(:��y�<�` �(D�hU�v�֎[ڈ�
�v�<QBf�4P�>$���P;����-�g�<1aD<}�����V���:!��b�'�L|�V�~ӄ��O�瓭Bo��L�Z��8p`@�oa��DQ�R���O���K<u��5�i>�d+J�+��%���T>tx%���(�>���D��g���t�ՉH�\��5�K��O�����'>�?��M���%[���yD���R"-D��ha�.<�H��5�N[̔��m5�O2i�'v������zBJ���kPW��,O����OB����Ob�g�Tdx�%FG�Lٳ�R"O�,؆�k�'4ܽq�g��H��@#���6C�����iG�'���|Z�.����/� �F��~~2B����:}*���_�uv��+у׭gz���q�n��uI��7?1��>�5��p��OR⓱��S�F�DH��%[:[��	��>�U�O��}Γ)��Q�҈W�܈��T`I[>�89�K�j��T�Dˢ^��W�Ӌ�P��I>95�p���)*\���(m��z_V�F���]2&������*yMڵ�`��́����ɶ���'�J6�CJM�����0`�IC��A$��	W�<�'�p"���L�b��&�*V�l=�iɶ%��ɖ7n�S��'�@ź�OFA1!��ű���T���rȍ�\\Nȳ+OV�S���ș�O�.�b.
��n!����<S�V�����~�H����?�	.~���"J�l��dB��*�EiU�K ��dF���?Q �=�sw�I�v�Jlbua�K�<��1��d�s*nl��5�NѦ���Z�	�����Ĕ�MCF$�;�h��gA�>	��IS��P}2�|"�~b�E�"0�)e D�dh��FK�<����]�,�C��
g`�*�k�F�<��)�(u\�(dG� f�Y ��z�<ᵣ[T�=-�d��p� FN�<A$.��Yx�ȫ���8���U�<i��Λa/z�wo��v��A��S�<q��un�hFGBsk�iG MN�<Y�D M�Hd�3���z��ჷi�H�<Y��L�����m@	]%RS�_�<��BPk����W��������U"O�E����&��%7��u2�����fI0�B���\�J�H��cȆ f��qQ�.Rl!�ڭ-i$��O��p��c(9�>Y��
GK���&�0a"1Z�,�cE$��tE�#t<0��`�+o��!$LV�|���AE�"���H�L%��Gg%�0B!��y�la�$��.e%�q�I
-Zȡ�"Q#N�!"1'�!z/�����|:�����%HL�3-ExQ$'7�#�;ODz �@�M/Eb��i_=6���y�͐o�^=qu/L������O�L�%�`��k MѦ���|����0�Ë�U5���c�(@��B�x�"/ek\H�R���$��x���� <Z��"'`�DɌ�MM��TسB�R��*���d��9��ΟPE��i�Î���i
�ϯz����'��;T��:�v��#C0yXR��%��|z��ɰJwv��D���a�ݬh�,�I�l��ɹ �Fe�/�.`-�$,�@� C�ɕaa�ؓ2Γ>>6�
$b�0��C�?`�L�B��j81�7�V�NC�I)+�2<�$%�3I"�i���@S�C�I	��Mh�c�(v�T
1�q��B�ɢ�x`�	�+�D�*ݧd�.B�ɗi%�q�����e���Z�P�M�TC�)� r$hoK���W�ÂQ��L
�"O�	���?W���
�䀌za�x�"O��Wf��P�v��ՊVF��xS"O�)G�Ý0���HW�!F�}�"O��õn� �`i��ٷW/�� "O�̲ `5��`1��JOL�{""O�IK@M������LJ�XZ*�i�"O�ĉ���F�P��W���9�\SA"O���#�82�j��g�ߪ).zq�"O:(q"�L�t���4��!$(���"O��1�����p������"O���6�Z"W:��a�Ϊx�LP��"O�lR/I^�t!Y��^�(�@`A"O���d��i֩�W�חop(��V"O���;q��H@T�*Vip��5"O��A�N��$�J4�s���Y�q#�"O����e2��mɖ:�6��f"Ot�����i��A�&@&(�0��"O�d��C�"` �ي[Ϊ�(�"O�
r�J�,Sbi�p �}`j�zp"O����Ю/�~)q�ω+YL��YA"O��ԑx�r�� #�婰"O��а˧:�P����s\J"OJ���Ʃm��m[�햄_�p��#"O��Q�jנ(D�#��O�,f �"O�5�o��hT�w)!
��z�"OȜxӌ��zTt�v�Y%0��!Z�"O��A�kB�oD��q�$B�"2"Ox��bB�w�hU)��^�V��x�%"O`p�`��{��VOA�+�}�`"OruQ6�Z�@�Z��'�O�.=0e"OX�ʰ��K" ����=Y�VD��"O8�˓�V~�4��T�^�@q"O��TH�v�����ǽ��q��"OrX��@\Ȏl����%e��"O�|$k�"kge@b.�wa�Aq"O�-��$j:%��X�J�X�"ObB�.\#�B	�]�"D�Rr"O�u�eE�(@�R]��e�#��x�"O:Y��,��̠�t$P6:���*OH�*���5y^���M�Y����'���(r��.qp"�|8����'�����0(W:���	�2��
�'�`�Gǝ6;p���+[�(,���	�'���*���<3qgɎV�|���'qLS���5sF���K�Y3	�'��h:��Tx�R4��#
0�:�'�r��6�03S8hk�..8v2�'S<�{c�\�Jd��R�H�S���'��u�U�S�4|�Y"ADT=�6��'z��@�B73\�k��^�7�Ҍ�	�'��M��KU*��	��22�U�'� �d�7UY���r΃fϪ�'��\���I7�U	��˽bIxM�'�=h3k�5	�� b�@,ZP��'K^��6h/z�lVGH9?���
�'���#F#@��頰)��*/���'�.�3��?2�<�&�M?q���A�',�](S�Ƥx���� �����'|Vi��/��R�p�e�DLڥS�'�z���֗��KU*Ա��'�,�3R
2���I��
��Z�'%�,9eDD�z���*0|l�=:�'������
��h�5k�m�h@���� X}�f�޾!@PX�c*|��{7"O�!��:T��sQ�:K��u�1"Ot	�����?�聒W�߾J甸ѳ"OR�+v��~Y��� Դ��"O��#\�T���!�ڼ)�#�"O��ѥ�L7k{d����k����"O`�:P�
7L��k!��os�D�"O�����;.��yH6�]`Bܑ#"O\�yQ&�6?؅��BU:�pW"Ot �B�Z7~Ea�����/��)�"On�{��0^�"����R"O����-�1Rt���d�'O䡚�"O�H�2 �v�p$[7|�zm�""Ov�	�O�1O8�{SM;��$(w"O���7"M�yg���P��m�8]"O*ifE�]@pÀ��q�^�(�"O4}��f��E��yY1�˂]���!u"O|0�ׄZ+~�2G�F�ı)�"O��k�V��>�sD�V�xphW"O�!�B���*(����=	@�A�"O��zc���Xɺ$L���q�"O|�꠪�f+@���-
	�ru0�"OT�EA�:\z��v-��3@!S'"O.,JuNؔ�����n՘W<\ ʡ"O�Ku/	�5麸��:6�jF"OJA#��z��N^�u/<�S�"O�YkF�2(���c���i3��3"O��(d/�4���@�^�4!��S�"O�:�׌d'�$"��Ž�@b�"O�Z�l�Rq�Ɖ�;T+IE"O�Q���=d��)���*D�s"O��@o��7��&�ǐ7o
�
#"O�1vN�9��5*�a��`�I+�"O���Ǌtka�@ߧ=�,8�"O�`5�P82F�Xsv,J!-���"O�lقaJ�z9��*O�b��q�4"OzĚq�@-@�2��h̖=���2�"O��(��B�s�~�Z�F�����#"OXA�̔9vS�iH������"O�x��^;:�2�{R�M{Ɏ|��"O���
\�RB�u3B8���``"O�$[��Q�Jظ���)y�"O�e�5�I�u�RI �cY�nq.X��"Ox���n�"wo��Aw�^!oX@$��"O�A��G@�Y5t-�@O�*6��qV"O4%�#��  �e�p΁-�P��"ON%�Dm�8t�16N˗�`�ä"O�YAB6~��j��P2��A�"O�I[�h���.����c��y{�"Od�yШƳj$��`&ӑ�4��"OZ8K L[)p>v,���F �%��"O���GE�M|20��� ����7"On �U��`w8I�rBB�%�p�$"O
9"+��#�.Ik�,��$��"OL�x��×|~�Ӱ��zir��p"OpI�ޯ7*�)��ɓGƌ!u"O`|J@M�X�\:�ʇR�HЫF"O�|3d�G�@��3s隰o`�"O.���~���*GG̃7@ �"O�(�	��1��Hk���3��H�"O�l2 �0v�S֮��o�Y�"OrXy����p��L޳k�*8Re"O���uG9*rul�OO�0q"O�1� mBr��q�ڭX!&H��"O� >�{d��4�@h�ˍ�C�fQ��"O��`lAaЈs��Z'E�QC�"Ot���+3�Isr*ܪp��s�"O&��'�X���i��z�~�'U��A�G�
z�Hp�נ�
a�'c�PKt@����� y�,��'�x�sL \��<Ȳ
t-�0��'���t+J�jj0Ahb��3;��'�(H����k�jt�A	)� ���'p�(�cP]�4 �G� �ʰ��'ZD1r���r(� Q�_9`j� �'GN�qp�'j66���8��q��'�x�(�\�n/49c�^�\eƝ��'�r`���B�}�:pP�� L��C�'��!��v�IJ��'|�z�0�'�Ɖ3��5?��S���m%�"O\`s�6u�V��b\�\���r"O���F�&��F�xP6e�e�u�<Q���t���3G��L�\��,r�<i`�[$2�)�)A��8@��H�<���H ":����;���H��N�<����"m�(�:V�:~��(��IHI�<i��A�m0��=(��[4�F�<��+P40�	�"]3*m3í�J�<Q!e�2G6]���.�8[���J�<��#ҚN͒,�1�؀m-С-	[��dD��c�6��q��29!�d ΢��6��|� ep��ЀR!���N®�(�i��f���2Č0�!�䜗j�XI�eT )�N$0D�X�!��P�؂K�5vQP�K�#�8�!�d27�Zq�ƃʋ8�8K�,,o!��ȓyn�ȹWɉ�,'����b?�!��E���ç^�<;�L���h�!�D�KC�$�aG�1!ҁ�'�)u!�D̂V����# �*]8�m�
q!�d��E�b䰇A�.z�:l��&�<^!�D� ����� � ��\UcÖu!� cIQ1��ԫ;����a�5`b!�ĳ(.h���֍O����jʵNC!�d�rm���$C��!�$��"8!�DS�@(-ؐã0���V�D0!�Ɓ�X	�C.��P��!I/!��L<d����P�2`��c!�G�Y��<��$	,PŴx��%��} !�$��v�P��I$�5��ڽtV!�dǏ|<�[
�Il�`�e�+GL!�k�|(� Ɏ�F�\��ۓf1!�$	1&^�D�b� }��5#R�'D!�D܁J3j�x��O!m^��Ô,�uX!�����s� �MF��T�N>U!�d^�K�i҅�bA�s���	�!�:��x�	�.h>��" �#�!�I&�*���g�,|<�Y�c�Ο�!��=7�Z��`M��v rQ�G�Y�!�$M�=~UcCc��������@D�!���KQ.�(S�X'�6���@0 g!��
&u:�Y�D�D�`	ǪV�!��^�;f�Y��K8�u

��!���Q~��↣C:���S �*Y�!��İK�lA#��F���`ΔV4!�$E
pP0I��EӬ�AsJ
!��*Z�\V+�q�����P0EȬ���� A�� eI�0I����$W������� �\�1pS��!�� r�hP�>�̴�$�4�MА"O��Z��ܶ.�(\�P̈�\֞-r�"O����ͷq�H00u(�-Ͱ�+6"O̝(��L�aD��l�%�A"O��Ig&_�n���r�ՁK����"O.��6� �z�2x�D�@��T��"OL�r#��/ܲ�gE�A`TQ�"OV1G"^��5�<� 4�V"O�t�����d�s̖�SՌ`ِ"O �(�$�66Ӵ�%�a�(M��"O�P3�\8!�l�� )똜�q"OF�3�Ē|��9��JF^�B "Oĭ�vɁ���P0�,�&\��s�"O�ݢ��߂6�:�* �f���"O�`K5��a+>��6�º!�!��"O����9�t��r�õ���V"Ov�R�ɐL_Ԕ@#+'}��|iG"O0�H���"xfBͰQDФx-"��"O�� ˸cu&q���2e	Թ��"O$!�`��\m
쀧�)}|e��"O@D��m��%���IZn���"O.��"I�9�t|Xr��4�zd�"Oj�E��G5�Ȣ$�3
�\h�`"O��)A�<�P��݌)��`��"O����I�C�*�H��C6Ǆ�"OXձ�'�r�Q�u���`%�Q0"O��*�IH�chB�rNZ�7F@�"O�m�e
<����"@�0i�"Ov�2���o��}Rj>{,a8�"O ��U#��?�XјԩɅ#Z``��"O0�8�����������xCN���"O��P`LԴ	��L�F�g�,�x2"O�eZ��K�e�h�CD�:g�=��"OdQ�o�4�&=��
!e�$%�d"O�4y%'�q��A�'# k���"O�S!&
FM�yiql� &��u�s"On��͢X;Q´HR- 5�*d"O���'�sg&<H�M�.0Uz P""OHE{����	q��J-��DKdaPe"O֜ڑbсf��x��,ߘBD���"O:Mb��Ҁ
�`|x���`�J�#"OP�Ô�LBI#��>���J�"O���⥏�,�G��/�$�#"O�|��	ڳOl��Ņ���Rȸ0"O*d8�L\�r�X����I�Jq�"O�qK����T1�MA E�f�6���"O`�����4��d�%#����V"OR}d�� z���C�ĳo�T�6"Oh��I�w
����L���ؚ�"OH��@���=��,(#䈓[���jq"O����ĝ~�����P�1H�q�"O�(����<@����/�����K�"O�,��E&Oɚ�pE�և����"O��Wᘏ"|T:`��E�["O��hf�̞�,��'��.�d�"O���UESA��=CpO|}`pX�"O:!*$�I�>5.�3���?sqʍ� "O��S�E�|Tl*0�ȃ �FYZ�"O��3�㍿(��4����=�x�x�"OV�h�̀+A�p�!�"P� ���["O6�3�j��y""�U�)��r�"ON��cQ��dH�d
)�x��"O�a�d�*jE0䍻B&��v"O:�:󩋽J�9zA�
�\��졀"O� <%s��g\2��Eo�8A�V��S"OB̫�>LD�`�L8;l���"O���A��"�|��EOB�#F,{�"O@���D4���Ȁ+�,�����"O���h��~��L�ҠIS�"O� �5Ot-���R0j>2p "Ob=�o�c�
`1�"�'J�KF"O�e� �3l �J0B�:�XQ"O�Es�`�%���R��P/~΀��"O*`C�%);yp���J^�?z�w"O$�pFA0S���)���3k�aJV"O�9CQi�4n�|�{�K�6cl]��"O*ъ��Mm��B5��$EtJ��"O�iұ)E>~+P��%@�GZH8�"O���ǧeϸ�%"V9d���"Oj��J� д B B�%"O%������q�B
@�0ӂ"O^�� Ս8;��홫zb�8�"O��������.��#��<B�"O �ʷC�U� `�u.�� �#�"O� �G�+��y�DC��6�4�P"O��*5o��n�H�6��u�+T��yR �� x��Ɵ6N˒e��yB�˭/m4D� )u���R�]�6K�B�ɖn ԑ�*��*��BeB�o��B䉞&漃�Ņ�W��YW���Zo�C�I |JB@�����	L�s�2'�C䉡�X;6k-��-�P녣=B�ɴ��Q;��T)o����􆏊�8C䉦1�U�'� -J2(b��x� C��*�h ���\�n���
B�OȪB�cL ��a��N�l��� �jC�	�te(I����*[T��љav:C�I$2��iB��90|MZvbQ�5�BB�	�}�P@������h���2B�	w��yeO߅[D
=��- 0tc�C�I"ɨP���T�ޱ"%[���B�5 ��q�/�~�(�'Ǉ~��B䉯�u)�h�)x����I�ՆB�ɞ5>.!���?������]��B�	�[���	��T=lQ
�B��_gbLC�	���o��w�5�5�[>6�(C䉾�b����O���"/�6��C�	W��=�_���3��5�85��"Oĉ`ᯚ�^�l���`L����s�"O�����+X�򽐐�M!@(��"O*�B��_�X{��
�5v���T"O*���DO� $�2l�P�L@R"O�iRD.x�"�ð�= ��z�"OX��Ռ�/\�P�;�'�m9�X��"Oн2�KF.U궡�P�W#I�!v"O����)M@�����KY����"Ov,��oT�}�
y�#�G}��Q��"Ot<ҡ�R�[��}+ �"fB"�#7"O����VU�VL��̌U����"O��SN�aJ
@�u�?jY�tQg"O�3ta^i:�0�9Tp])�"O�)�ǔL@�ak��7�D�J�"OJ�K��R#XxHQE�#k��Ųp"O� {G�"m�(Y��Id�U"O!ҧJ�:���{�Ǜ?}b�U��"O%c�a�v�@4 ��£ -iW"O���퉾k/�E��e��5hRV"O2\�2�{Z��� &���`"O� 2H�ЇƺI��lڢ���; D\P�"O^��2��<mnq,�Kh~�;�"O�0�bݸk� J\H-H��"O���wf�L�y���9�|�"O@����4%hX�X�%V�'4� ��"O��j��_�N���#d�d"J��w"O(�a���[Fd�Vj�=;�q��"O����?`�=���v*4=�w"O�	3�A_�{���5�N+�8�d"Ox�h��έ 1����<�\
u"O� ��2�T3�cB
��Yc�"Oh@h���b�,�-\YV�bg"ODd��)��7m-St�+�"OB�#� �Ak4�
�E�?NY��y"O"L�աQq�*�˦dQ�MP^ؚr"OXHa![ l��0����sE��"Oz�
@�
l���/͚t�{�"O�l��NJ Ne��DJ"!v.�rq"OL���(9���w�AfF�IV"O��0�ٌ 6�!��ݻ:}�0�"O�D��K1R@Q�Ud��.x؂"OB��N�#d~ a%�v{��`
d"O���M�9N���a'ݮ@���"O�p��@S2U� �O�+��=aT"O�����R�G����C�J�� &"O��hÁ��7��=B�Ȅ
�l�0"O(�s ���48L�s�A�M�TX�"O�!F���@L��S��7j����c"O�M�`C�1Op�y� �YK��z�"O�u��f�%����	�)x� ���"O�̙�#]W8���$he��̰6"O�|Ô��>t56�hE�"qd ��"Ob�����j�l���n�x7j��"O>��b�L��i!B�_3$M�W"O�ۥIܮ`��8B�Ùy$�:E"O��8�G���*
���40eJ�"O��9�G���!�����^J@�ۑ"O؊tc� FĹ�Sf�t��l1""O������A�֗\����"O�h���#Iv�u��*#��� f*O��[�o_�r9b�u/D�~V�Tc�'@X􃛵p����P�*6,��'fv�Qa�̈́:�<�;E�
#���y� _�R�Y�'ˏ+R���ZD�́�y���m��oO�]�@!(���*�yRFC!M�.];�L[�-l�e��O��y�B�4'd�m�%��R�AV�Ɉ�y����颥���߁&O5Q1Ȍ��y�V6z�t �e��\+2�����y�b�]��0�L�c�v���	�yN����Ө|�,�3�"ހfI!��0C�PI��.́�Rhs�4!�!�dV�Y�4a�+��q��P�3�=^5!�G#Y�"t���.Km�ST/H�x!�DƟj/�;�h�'a�4x���}!�d^H����WVj�T��6�ÅKM!�$ۜt���4��4B�
�$�*$!��^+(Q��IFp��paΆ�37!��]��ӓe��:]�.�3!!�d��w;�&�ʍU���Y��!�Dٕy�̕��/��P�0C��W�!�D
�8����M�`���aE#�!�$��
>��:�n��`2 �Z�Qr!��9p��p� �"DN҉�U
K!k!�� H��E�%
QT��Żs<��h�"O�0��3_���2-B4%T���W"O�Cf����L]5VH���WO(DFxPK�hɀ1�TUb��0<O�؉%%WR��H5B�����1"OP	 ��R.c�l�����F�,�"O~q�Ua�L^�V�� q*]��"O��bY+�� k��ܕbl(���"O՘U
C�p6��;��#N���r�"O��`J�H[��b�,J�%��ܸB"Ot���ORiN�A딚{C�=�"O���R�'��x��/]�S;��4"O�l��L� 8,q��c�P��"O�p�E#�%�H�CT���u9p"Ot�� =];J��Q� �j|�U"Ox�E�G�\)E���O�r��� "O�0���^�E��9��O!����e"O��V��_:�h��ԭ>V�yx�"O���eʈ8���d)Y���%x"O~�+�oT�g�R�BӇ� �`LѲ"Ox:A�S���3���N�b�y�"O
]�)A%PG6���KTL���x�"O.]ᗁ�;�|�Jre�(u�f��"O�,��.R�'�V��t�"O�0C���&>�d̂sÃ����"O: ru���hz'b��82VL�C"O�:&��K���	;"O|9E"O�<���A��Lx C�i#�T"Or02�i��ud̓�얓k�.��"O���Dҍ���C+A�2d�\a3"O�h�C�Ԋ]��������/  i2�"O!"��w�blڧ�}l�I�"O�����2q ���P�8 dѢ!"O�\���8�>�{5	U�(hC�"O���b`�F��V���=�Ñ"O���G�*�ΐxt
��uXx��"Oty�gaS�vX	�w�Q�jl�9A"O4hag���f�# L���:#"Oڡ��)0[l��n�/��H�"ON�:��Q�d���;����jɁ"O�`�� �	h8ĩ�I�'QР��E"O�`��u�����.@�qn�u 5"O�qC��P�J<��P�64> w"O. cu�;u��Iӎ�:b0�+a"O�=��)Z��n(@�+�8 �#"O�,c���3�m3t�W����"O���V\X�ԣ1fAl�\Ѣ�"OJ��r.+��L
�K@j
�`�"Oj���a��0�aqh�`��R�"O0Ѫ�F�\`��qU�K�q�6%8"O�͸f-�#k��E;''�' ӄ�H�"O��Xp��!���A��漳G"O��e$Ʈ>c�3�C3s�RPc�"O� Awc�0����e��V)�k�"OȽ{��:/V ��T#�!S�"OV�� #����0 A�%�qx"O2aZ$ �L��q�B#E��S�"O.�&f�8�+`�^�3��I� "O$�Ȝ�gPdp� �l8Ġ�"O�]3���҆�@�� q2���"OZ���I��)�D`3��\�%+�1+Q"O�tJ�͜\����1��?1�yw"OƨÂ��5#��Ӊ�d���"O�NTd�&���q��"OAc�aJ��cdR�R�x��"O� �A9�g��1e�A�%d¸u��df"O�(W�J���Qfa�f1��"O���g�R9���aN��(�
�
"O<���O�`��ْ�������f"O��)E�_�3�ĥ���^�,����'"O�$�d�����;ń�,f�0P"O@x(l�%�\�3�Ƕu�@e@%"O*|2���94�#'�5�b	2�"O�!��R�Լ# _)�j("O6�у"[&%*�9k�O 7.�8YX�"O���ZC�mQ%�ۊ�ʁ��"O.��_�n!jƮ�6]dXP���F��y�C�0D�Np��Y�>�>�:�Ȁ+�y�D�ybxTp238�d�"�Q��yҋ	t�tf�ͪG��%i�ID�yR�Qh�8�y�D�l[���'jܲ�y2���Ӓ|��昹h:�H��ٿ�y"
\7���A d�>["�X:�����y�T��-�0��O�h���#�y�KB�L�)��MܫFK���'���yr�T!k�R	ئ��8�f�1�K"�ybm&'j:`s
A@�������yb`
Qhb�����;�
8B$F\�yr�7Dȶ�h�G^*|�����k��y�G�EIH��l��$p����C?�y��;K����(��-�0�L�%�y"�
"}y�Q�P���P¾Y�PeY��y��h�b���mZ�F����Nż�yRAŮ&���"�>8��Y$�߻�y�瑒+z����Zp�Q�3nK:�yBI��'I�P6*��8�c߭�y�"λ!J�;Q�
-#�N��C�T5�yr��cEhA��m�v% ��(�y�/�\�h���ufv��`�&�y2�|�$+A͊0� �*�yBᑸ4�(k��Xzp��y�!��L1ag�Ԩ\��|���yb
��<�X[���=S5
��C�T��y��v��'�F�O�� yr�ѣ�yҋٟ���2�A7���l���yDR�&Z{@�N�"8�Yq�֮�yR�']3
� ��5��)�y��SZ��o�
��t�d���y���;|wk0f�c�0�j��yR
�+9鉓�Ida�4���Ň�yb[*�8}�bn��eʸ��j���yrƈ;by��j̏a7�Q�@�%�y��|�Nl�!Q�S��=*��y���=���i��T��g�^�y2a�5x�%iq*��p2,�8����y�툴x��K����ĕ����y&L��~���e\�ڀQI����y��v)�2���������y�L�g�\mKC,F�"u��S�y2�
�V���͊�Q�l������yr���t�u����'N?H\kW썐�y���~&�9A'Ȇ�>4���B���yR`��K	 � 6��@X�m���7�y��D��	�n�F�ű�J���D���Oٜ(qQ#O�&_����'�29����')�1��`˧hut�i�k�3[�!�'_Jpq�B[�G����@�4(���b�'
�������4q��92��
�'���g��hfK��dY�H�	��� �5��a
Jc�3vҫ$�HS"O~I;S��vt�*tA 7E���"OR�1�[< ����#@�;w�V٣""O��s%�l#��t�_�^x����"O��k3�94Ҁ(넪P*<qr�!R"O�e����S� 9�ԉYkbp���'k�Y�A	�X�6�K�C�y��9x�'��@�v�ԧUvP�/�u�`h��'����5��M@�:ԏJuv,0
�'<���<<��L�� ID�nɓ�'��\�q'Y�I6^pHZ�f*z���'*��s�Ļs}LdAG�	n�$��'&�����1;!�,RKMU��"�'����c$¡^�Z��Q�I4��M��'�Z͓��O���Hڹ2:؁�'h6� mĤI����T.��xE�`��%� �&P���\�^�ر��j�<�G�ɭG�\�s�
k�9��J�h�<����'-h0�ta�-4x�d��c�<���(�q*���0$cI��ЅȓW�A�2�P��@<�%#�dV���ȓ#*��2n�p1k��Bg�������C�f4:`YL]0�\���n��1��O�3.�x��E��(d��^�
}�N	�ޙPG��|�@t�ȓ}��Q��IC��R# ~}�ņȓ_�@y��g�8]��:�-�\���u��������b��:�٢1�+D�����>�l5��bD�u����l+D������ �X� ����%D���t�S�R�9�3��	a��C��6D�$�&Ꭰ���Sf!�?~�y�"D��BL�$|�Se�wȑ�s�<D��z'���n�\K.F(4&h���-D�����X��<Zp��%6DM9�A>D���-�JA��@33&>�s��;D�t[�F�Rw&��I'?�4�ؤk;D�ɒ�BD����X�F��qCa�&D�Px(S"��䡄�*҈q:Q�7D��c��|6)+�}d��7D�ڲ,�%\�bͩ�nZ$X�J��`4D�l�0�y�X ���+D+$��W'3D�8�#͐[�|�E� E�ȫ��2D��c��%���P�h�0eB�=��g5D��+¦Bk��+%`%zb<K�3D��i��L�S�)�Po��^,S�6D�XS%6t��i#�E��5q��Zu 5D��i���>2N�"�@	�#̍�R�6D����w肄����[��C��3D� ��Ҽ�h0�&� �7Ι%�4D�H���w�d�[���8+�t(�g?D�@��NU��<��F��>r�>�A��?D����,�i�:\�b��Q�N�y 	=D�Ի��E�~r��12FZ!!��R�G%D���Gг'�0����Y�P2ff$D��S#��V)��C��o;��V�6D�����T���B�E��� "�?D��iP<�9�O�M.�p;#d D�d��
"@3�XG-دU����=D�0x �̇YQ�}�͑�܉c�j0D�tH��ǽ�j躳���p��ѣ�c.D��� h��m:�6`�V����6j!D��æ.V�aڂ��2�V}��B�?D�4�W�ˁ�v�6 �<���ď8D�� ��a	ty�q�A�2�B�b�"O���	O*�A���gի�"OH�1��ɑ]���9E)���2"O�}(���P���D0�i�"O�ͱ�ƣ+4pA�)�e�|�"O�a���N�vE���-L߈�J%"Oi�S�[7 |�`FȄȄ�"OX��5��	R�@	c�_�Dx�"O�ę�苮������)J�M�$"O�(@�W�5\l�Y0��'@hd"Oԭ 兂(i[dX����$_Ɛ)8�"OHy
�&�Lg$�C�K��n��4"O���C@��4��e�1DֱqrVHu"O���C%E6*�`�S��ˊyL����"O� :Q�܃~�U��"T��8��"O�]z4o':�Q���֓!���@"O�􁄄���b����$��]q�"O��@�VÚ�� )_*H����"O�Pqʝ�h~QY���e��Ś�"OnJH�^3�h��������"O��C���LI�Ϛ�17,S�"O����e�;�%Bu�-~�	�E"O�[�EO�	�p'K�)=�8���"OV�ٗ�O0
<h�%�� u�~0P"O ��6)ɐA��ء�ОD `��"O��#�P)%Ÿ郥�]�J��G"O�$[q	�>l)hV��1[�i�0"OP�Xe�	Aqƈ���U�=�ެ!�"O�%PW�H�^,�k��϶4��"O���1J��
n`�f�K�����g"O��Bj�v�+b
�%;�����"O���Mɦ��1��[5#�L1K�"OhK�kJ�}�ተO�RĨ�"O��c���
y���J�͗)%� @0"O(�ӣ�&�ly�B�5��ͫ�"OdI��NŬAn��������`0"O�\;sF�#gd&���֪:M�U�C"O>�ö���9ż��‘�n4����"Om�U
�kF<�d�8/ܙ��"OVQ��ăq��H5�3�!��"O$�֤�\��4H�BQ"��͂�*Oj����"+�
Q���J8�t�'��0yW@��O�|�EDNs�$i�'Z����V��0{u��E�T��'�dux$$R>(�tO�6;V�B
�'<c�I�����GJ  ��'�6�S�@D�\�\94�Yza����'�K��ϗ=�d4z3�ԡn��(�'�1)�o�=�!��g�h�>���'�ΨзJ��YP�b�N�4w[�T[�'I��B���*@0�շi0�@�'�����I/ռ�0r�@"U] 0��'����%�mv��ġN� Z�}��'�>Pa�#�WY���T� o۞�y�J�-��&��B�:�')Õ�y2��)�d0@��A�3���d��:�y�F�+��1��1���N��y��VN��!LI8:n5����=�y��,_��22�F ����f$E��y�6>���D�Ћ�t�����yR�	�r�<!XS�[��D�q���7�y���i�:�9n¼Gn9���y�$Tİ@!��"�\�`�#	8�yrH� �P0`��:x]��gC)�y
� �١O׉y4T
�B�k�,��"O��r�_�"���q_�q�dT�!"OΌ�Ui�#u���V S�w#X%j"OF(���Q�K��3�(��2�,� "O|I*�!�We���r������P"O@��P�]Ϯ��%&�
	�a[��	i�O~QpD��Vd�QK��zH|��'p���$&IΝ��H��t���:�'�B�@xA���?
��'�TUb� �+$!`YqP-K���s�'q.�z�+��
�z������n�V��	�'�R��6g��OlaQ`惑#�|{�'�"�2Jڥ�d��W��> ~N�j�'_J�)���  M|�I�Q�_+�t�<�B��2I�5�d��N~��p�<I���;!�=�d�Ɂr��=�lUi�<!�N��y)|isFY�\^� �d�e�<��߸d����A�QA�2�I-S_�<��IP�vdnP�`�Ը+æ��Ǭ�Z�<��c�v���2 ӵH4��R"�j�<�@��^&���aֱVu�����L�<�7J5m*�Z$n��n�0Pˠ%L�<I�H�H~A㲅32�83��H�<U��@F��#׈ψ+j@8P)�L�<�1�R�iqvР2���v2���D�D�<���4-�{U��:�t��,�J�<蚷3�hH� �P8��H`��C�<y�D'K�tAKQ$��0�3�&~�<�B�ְXN�%���+ ����[w�<�U-ַD_��aq!S
'��l�aa�u�<q�n��P_DI����!8
@;bng�<� I�-^�� �� L���`*v��`�<�C��
�l��lI4x��2�F�Y�<�Os㖤�FV��lQ�a��y2�ϊ(Y��K#G�u7��#���yb�A�e�r�2��i�f]��Ѡ�y�E��t��� �(d�@D�aG�>�yBb���1�E`W�\�X	��]��y����d��hb�M�}W ɋP�A��y�l^1t*С!�K�+�La"�bĈ�y��Q-T]t��b�2}xF���c^�y��~G�9���w��B0ő�y(߲`�|[�hwk�=��� �y�k�8�ΝrG^+N�s�"ڀ�y����q6F`@@@�^�閭��yB�PC��m�Rm�(v*�l;����y����;��]�4"gJ. @5�:�y�� ,l��,�✪W��m�i���y���j{V���&��̙��J��yҥ���<dÀ&��1�^4��@��y���GE���ņ�%<8��M\�y�(>T�A ��*�81�W߼�yb�0w�&Y3B�+��m�5����y��Da���X�%V������	ܯ�y"d��[jD�)ѷ����D��y"���/�D�����.���A�ذ�yr�,dx�� !�U8��F�y"c�>���1Bļш	���^�yBӠ�J����f�P7����yR*[O|R��Aŀ~E�R�@��y�hW=2=L�xQ
E:}E��P�y [�0+R��5��#RQi���y!�`�����ąH!����ć��yB%f�&�.��V"��hr`�*�y
� n��� 
�iv��	'���K�l��"O �"�F��)�д`��=��8�"O`��Ñ7��8��B�i�T���"OFd�w�P�b�2=��H��)�Pa�"O\�k�Ā+Q �I�չb�tj�"O iK�\j�1��I�R���B"O�`Q^Xe˄�Try$��dI*|�!���82�
�;@nO�>v�]b���K1!�DD�/"4H�c�=5�&hs����;2!��V3G^V�akS/ߦ�)3,M!!��0$ò��C�B4y$m݄N{!���I�m0��Q�{d�d{��)On!����@a�f<����HU!�DӰ6�������1mJZ��L�wB!�Ğ3���pv`ͣk9�m��쌪1A!�$�4~�̰3Oѱ38���I�	o.!�d�+m�|�D ßW6z��+V2I!�d#"��G�X�tTM�s��5YT!�$��tX^�J'C̡=���a[[!�d׬Z��e�(��8�W(�LF!��F#4��a#�]�3�V�� ��B(!�D�$��lRR�ߕ�0�tB�0m�!�D��Ͳ<�g,ƖpZx��fBM�!��4w����f� OXk��G:r�!�d˔]����Ô`@�H�E�D!!��$�LC�CC1V�"���#!��u��Y���o\�1`Lˎjj!��ԭi�>����!+����E�$g!�U&��z���L
ؕ�a���!�d�#Ĭ�3�m�"���+@EU�A8!�D��^���Q��� h�h�"�-!�$aE����Fw�D�!�%�O,�ȇ�iR�Av+�w�U9�@��Aâ0��t��XNF9H�BX�%Ƃ��`�ȓ3}�=y�؇AE��z��SYp��ȓ+��a��ă5p0BD�D�]�HՅ�D
��u#��(�q�jD8?T@]��@�屃��8#D�(�i�Jb���h�^�/��2�ȋvnV����K�<��(I;b���@����&�X��BN�<y�J\=&�mȴ&��`�]0�#@M�<�%*ЊwHZ�)vnnef}��F�G�<�ӧ\�xҚ�(��Y�D%��kơ]F�<�u]�ތ�%�H6�����)�<)�b3I�vU��9 2 ��AIPx�<��/	��]!#�6Z���wo=T�l+a�$U�|t�0�.6�\���5D��KD��G���Z�G�;:�}�3d5D�,V���C�떢L��B1D�0�uGZ9��`���+�����i0D��C$T�.E�T����:�.D�(*�'[7�~�9�dP^��QqRO-D����OE�FXc%M�0��@2G-D��Ń"M�8�⋮��1Q�f5D�8��@�hF��`�H�}f���W�4D��K��̃p�`a�s�R.+�}�23D�ܩseT'0�q�T�4�	)C�<D�D)�ˌ?.z��/Ґzh� f(D������� v�Y����08�8!S��8D��ˣ��;GR|#L��skR�(��7D����W�3�hyB�)�Q:Rᰱ�'D���b��������,X�<0$0D�����^�Q����[���xT�-D�P:�c�3��7� 	}�|uy�9D�� N0w@�c��� ��<T�"Oؽy�#�7IȬ] sn��$�d5"O�{��O<$�����BR�!�T	r�"O�(Ca��)2^�����#q8��"O����9�Pc5�@0�"O2�3�e�v�@ ���.��V"OluC% �<!ZL�$�8r
��e"O�Z��U9Ga �!�A� [n��"OF٠W�c=0iJ� T0n< ��"O�P�D�)^M`��Eo
l8d���"O�52���#b,ʍR���Z��u��)�O2�sc�X��MìO?�I�i�8�voO
5����f/��Q����cF�R���Y�N�\֦5�%P?j�>!����0�w�_$Dg�P
���]JU�i�PM���Ęj�I𥟯}�ʉC�s��B��~���2��%�-�Q�wӒ1��'�7MC�����s��M�5��"77���v��|�|k�ɔv?����$0,Oΐ2�K Ek)�g 9zĴ$i3�䦑yڴ��+m"�)]w0��c�,ֱ�E��
d�}���<�&a"���'��9#!�F�ȡ[��ɨp\��2h�"�4PQ�Q�w�<�������Ɇ�O�hg���q����U��(��@E�&E3*�
&,QIچ1*�G�!=5�(�O�����.����M
<fb��	��H�Ƞ��HʟD`�4J��gyR�O���9MҘ�	3+T#��a[Fo4�C�ɀx��P ��ɋ'�
����7 d p��il�7�)�d��B�)�<���]	���{���+������b.�y�'Ͼ��<���1�l ���6T'V�A�90+&Q32Ϟ�(u�t!b���D*PD��0#?����'����
�)� ,�e�R|��0AF��g�&�0���L%�5;���D�ҽi2�aЁ[�$��C
M�'u� �d�G���	ey�'*�'�����x�,ĊW2�hЕ�~���"O~0ذ�]�@�$�����P���O��oښ�M-OZy���������I�ӓY-X�4&IS~���7��P��}�v�D��,�� ��N���>���󒂄�D�%���&(�j@鉒'&�YSDD���3C�u�҉Q�O���S�z�p�;��յC9>={����2cӐYo���O�F8V�	�h,��+���84��O�˓����O������gԓr�ˋ\ $0��'����uӜ61'��X�P��/z �:�eY�������o��0����_>˓��8����j�{2ck�(ʱ���2)�#I�Z�:X��C��+ʒ ��i��Ɍ"1��`�0B�$�Nd� ���MK��Ux����#[�x�<q3��E��|�1y�������xa��[֎�
O�D�n�yC��d�Eݴ�?����i&. :s�_�Ah(Yg�՝0���'�Q�h��C�S�4�ѰBq������$���ڀ�E �(ON`l��M��;`���'���N��Ȇ9
@�Sf�S!�|C�gy��Z7K�6-;,OjC�YVh���0`����e	�vE `@�"�R���e^j��5h�|+W'�	Ff�c��R�e�@DBÄ/A8�r��8B���je�J�F�����v�dȭt�R��
ѹo�l9�f	��� W�����O �$���	Ɵx�'J��H��+�D��%~�Xh�>iv�S�3?�����bΨ�2�Ӥu�����i`6-8�4�@��?��jӊɕ�  �    r	  �  r  �   $  b*  �/   Ĵ���	����Zv	L�l�H3R�PΓ���qe"O��r��<���*�a.�s�"O��Ѷ-��cU��`ȋ�}E<x�� �h�(�BVZ���y�E� ��)�&rq�X0͎�imlآ@#
�t�t�x7
Y_���A�^,(~
�D̈�I�x�P�+�'&�ĕ""&�DФh9�Rs�z����[&<VZ���Ϗ�U�u�㑘B�y��e�?7F�e�N֊'D�q���8�:�mC��?)���?�����*D������;<L��1�C�I�� �I���y�&�6,����bܘ ��3�%ҹZ2O��V�J�W$�8�S�P�%�Ԭ�p�T�g�:!q�Fx����5a�\&���r��o$~e� Ī�����<��e�ɟ���w�'���;:Ǌ�;�m	�X��J3��n�!�ű��)1E����A�L�!~S� l��HO��O�ʓlC�#�$K 3��#hH�op�b3��;=\����?���?AT��z��O���U��%����cf����rn����[t��9�`ݤ|�����#Cm�ʣ���j9zQo�#@� r��Q�z%����>&���oZ(-%��)��bѢ��5@gHe�%d�"5���ѐA��e�n��M���D�O��擓\#@����ǯE��Y⒂٧&�((P��D�O���2�i���Wc<n+��4���8%w�V�dҦ��Iry�DQ>U	�6��O\�d�OkLR�Er��r�nͳP/�����g����.]b��'7�[�y��Y�6��W�b�'��� uI��9�J��%��9D�+�ў �O�	 i�����/c��	/I���"0-���+f��/c���ʦ��ٴ�?y�O��8��ƈ!d������'deK�498�����?-O�έ?�K7"j�d�(@�`���|��L�Ă*,b�'�ў�8��$�f����LK	uDb���̏j�`�'�&Hh1�`�����O��d��48�a�Or�D�
@*zu8@��0�\H� ��w�@lګ'nޔ0ii�%+b���O/�S_?���
�m� =X!��T�6e����L�uiޞ,�<�_���|��
�X���Q�	�%�$���@�$i,Q�u��X�z��һ?�r��)����Ƛ�'Iq0���A	Y@�'�<\Pr���D�O��d-�S�>Xyؓ*x�����Nufb� ��"���<I,��8�0�_�+��_�v]d|j��ʦa��џĊV���}��ҟ�I���\w��@ ,r�,p�%��;��P��> >��6 ��ɖZ�]���A��a��A�+;"�Y�E��I�S���d�i�zm*6����R`�Q�Ɋ�0=���6d~�h@�D�$z��P�
o�<�$�=Xy��8�%�? ~�|b��Ԧ�K��4���Op�d�=aϴ}ːN�1Gv�i����.��<��l�O2�D�O�d�Ӻ����?��O+d|{��h����B!V%X�.��fC#�M�&5�O��e�O>ݑ��;F�RA�BF�#KE�����'B����m�P��>�� a1&�,EF>�9V"O ��(U�b���
���}8ำ�"OD� �$_�4D�Ȋfm�C)8K�R�X��4��j�p���i���'J�	Ь���)����%Çl��q�C�<.r�'�2�ƻoU��ԟ�=��S�U�*R�'_ ���ɒJ�`�~�J �v�@��v7hٓ�E�'p�"��5�>�:4�!ɖ}� �5/���3D�H�&�>xS��3���w@v���-�O~�'\���PG�+,nb'b_�3&`��O�X`s�+1�8��3���a�!�	U�F�с���HJ�Y��
�H�B�Is�\���$�h*�l�S
V�p��C�	�U�6�Pv%'^tJ�7+�a�C��%a�
��'n�,e>�a ��V1�C�	Y�IF��'y ̏��rB䉞^g� ѶG�:���*�D�XB��-$r�@�k%*IcUHP*}�C�	;6qf�kcc��B\�Q
�nyC��5C%�|���O9 �&`��I��ͅ�B�0��-7a1��7Xp��>(������}�. ���Ba��ȓa�<�Ã�����b�Q��ȓƬ�"Ȋ�dy�Hn�N�cXXA��`]���6,GI�!"�jm���i~����>_^��A�� Y�����7
01� �̐<��m����>MPɄȓ�,�+�l��X��LI!h�9|Z.݆�cWve�0m!�YBA�23���c���T�Q�B�-`r�Sg<>���S�? �-��E��p b��M�'^���"O,`��g�����'%C�+�"O
��V�A�"\2aP�`ŀ`�"e{B"O��;�	Zl�*�+E��2]��?�yr������EY2A�����/�y뛪H\��Â��@�f��'���yO�K3��Y�	|lK��˭�yR
xi	�#�?0��&F�hk\!�ȓ}m!3#��JӦi-Iђ�$"D�DbɃ�g����D��vE���!D����G
3��lC���F�vٛc&/D�@X#�"�($B��O�;�YqP�-D��ѵLӜSO�A�!jZ\X�젔�)D��R��>�T@���8t`��Q )D�|��.@�����K�w��ZO7D��#�To}0H���:?ޅ:�E4D��r���,Ӯ�	�ٓF���2D�$�ǆV�  7&�[JT��4D�h�e)ӥ]��}�gD�_� 0qql>D����%�Jyf�-i	����yKY�Uq����iǁ}G�M���R��y��*T��&���Z����'�yB��:�Ȕ+��1Hì���yB]1_����@�7�6,�i��y����W~t�����*C�4Є�[��y�/�	�Fԩ��Q�+ �E=�y҄
�3�ʍ�i�%Q̉c��Y��y""ށ]�� ���]&V�llX�� �y-\�t4��D�� �����چ�yB�Q�̱p���R��EK��yR���,���^U{`�ǎ�y��ܣ����(�xA,��#ѫ�yr�L�B,��� ���mº�q�$��y"FL�� 8�� d�tQ������yb�EYҕ��(ר15�]b�,R��yrD�>]��P1� ��([���v���y�H�/?��Xrc�B�(tڱK�+N+�y�B�J ��0�ޣ&���C����yb�)uH�Ha·#����JN	�ye��5N�i �:Uvv��L���y�H����1��@K�B}�����y2b�8\���C�76���IRo�,�y�U�X0���1/�* ׀����̊�yBϡmZ2���ˈ�@PF�B���$�Py��σc��(G��:� ĝt�<����*�!�T�U��L��MKo�!�$��V2�����)!6���e�2uo!�?V�)��7O� �'eσ�!�����c4l6(@�0`劊�_f!�d9=��)�#E�*�Ԡ�	ŽE�!�d���h|�D��3 "�A J	0%!�-�`�Z2FDiyDs׉;6m!�D�3"$�ҭ	2{���!�!�ȕ%�ec�Ɔm���n�9K�!���(����D.&4H��ǟD�!�G�+Z�C���~*��B��J\!�ҞMtm1��'f"�ReS!(�!��B�SԊ�ztk�/�����G�O�!�D�/N�Ԥ��R�\�h����ʵ�!�Dˌ5�z�To��&��e�� f�!�D�a��A�Ǥ��|`R&���!�D�:MƎ%ضKΡ3xDY�bW�`!�d(Jn:�`�+& ؊$C՜|}!�dl�jfn8@7�X�d�ȹC����� ��KÆ�P�ܕPvO6~z(!�"O�$`�G��M�Qd^���bO2D��o4b~|�#��ܖ����?D�H�D&Iֱ��m�"f�h!�O<D��P���7c��!����5�4���;D�4!w�؈Y���{��ՙ2\Ġy��;D�t�'.F[KЂj���K�#D�BS�Ŵ�%1A�T*���6D�Th�	5�6=���o:�<[�/D���D�,측I��گ6褒�/,D��J!F c� ���Ư��d)D�<�D� _)�܉�.X�I.�2�d3D���r�	(dw�] �7�(��Fb?D�$1cc�3"Y'T'�9 �'D��Yq� tJ��"A��5UR��!�'D�|���4p���R�� u��I*D�`��Q�L<<Րe�!(�4�h`	=D�p�Ŋ��3?F4���<j�Q��(D���#��L"^9���B.���(D����=<6��̜0���B��t��Q�k�Mx�hʗ�X�^�d�e[$�n�z��/lO�mi�L����	;=�l�B�ĜP� Pf�*��B�I�4b�Ol�<)�[p�Agk!�"yD�CccQ�W�bD�D�H64Gd��䫆�\�\�2�'ݚ�y�
�vԨ�ʐ �[�8t�1/��kC�Z�L��ɓN��#|�'wx�'��.e|ȩ�Ǎ�&f�1��'�@���G�O�2����8����K�~E��!�:K�:���''PyB"��"^�8��@�>zh}a
�ż�s�Ǒ*d������
H*��t�LL�H��ulB�_w���"O�\8��0�����]4e8e�>Y3c�(Jp�qa��K�� �/�'S�X1�0��P�aA��yl�%�a��NT^����ER�U��nNY�L1�@�e-��4I��3�q��'{f8�Q�..���ׯCyĥQ	�'�f9�U���PJ�0 �6�0E�X�N�	��� C��p�i+��y�e�A�|Ё�ۥMnP���J ��0<I��._.lp��������	Ā#� ��\,�Yc'ĝO�՛���qh<y��БP���r��4��q	V~B�	H� i
w�(l>8bc��̄��NLo<p�"Lx��w"O¥*`�xjʄ�!½�H@s L�BFp����\�l�"�y5��$t�1�"�O��pu��?	���e,f�T�O��rq&�nN�m6���y�dȊE=&�	��,˦ �Hٙ�E������d3-�Q�P�p���t��x��WJ�4A�ƅW�'��h���#� }3��ͺ;wʜq#�$d�ՅȓC�<�9��\�=_Ĵ�5KņwyBQ�O��k�c��Mo�v���u�����I�'R��3Ed�/����nM�$�!�d˭Fۦ	I!r��uƙǶ�h�e��Q� �O��}��&���xs��D-r���^�	(Fd�ȓ���{���E�n�)w.ܰl&�lZ�<�����-}e΄��I�|D6�A(!��U��?l���ĝ ��z�/���?9�$M%�8���L7M>��B�F�<QS�V�O7|m9G;<t��C��B�z�� ��j��*6�|D���_F@8A�* �j52$W�M��y"B6j��yY«�d[���F��h��a��"�w�	��H��ɨ1i�i�P�݈ ]���W)	m5:B�ɢ{�:�h/G4��b���'}bL�	�Vq"!���!KN��� 느o�j2�D2L
�C�Im�� H\#&�j!ڡ���vB�I����a ��BOF�5.\#Wf�C�Ɂ�v�р�G`���f�a�hB�ɔ6
Ta[�aS�8y���� �K%�B�I�7�ޑr��L9V�4��c��=%��C�	�i��9��&Q7Z�*�� ��qϜC�I-�. �p�H�>��� �־"zB�	�{G��Ze��!H��\jd�վ�4B�)� ����.V�<
��8�n� r�29;�"O*\Af�Y\�iC�o-z�A"Ol(vLT4R.d��oߧ+p��"O"�A�Z�V��n�6jE"�[g"Oj��cO��eA��W�Q�dhY3�"Or,QE�&s�8���`X� E��+�"O8uS`� �7H����7\W.��1"OnŒ�e�zo�(��1 �N@�"O>8*tǄ1�ֽ�$�)�L ` "OT�#(̌J_Z$�&+�"��T !"O<�##�+H�HT�)��MS'"O��d��U�0Z�	�6��1)�"O2�)X -GIc��K�o�}�"O,� �NF�q:z@`v�2R��iJ�"Oƨ��L��0D�H�m���Q�"O�Q2�0�*5��|�RH�r"O���r��?�R@����L�n�8�"Ox�1����(F�.d֖ɀ�"OT�/�5;9<y�v�#t�
�9a"O����I� Βq %���X�d"O��!�L�7��C�` S�<�@q"O65����#R��) E�A�<&�8h2"Ol��뙳[j��8�N@1*:��6"O��	��oЧ�b���"O�Y�C鄦H#>0�ǣ�%[}>�1"O"!H� �|x�K��&���"O���߲x�I���/Z�|,��"O��kT"T� O��K4H�
�P5"O��s��[�:��΍��h$"OƘ`܀.�e �9Qxn��s"O ��ׄm.y[ 
R@�<u"O�EP�e�f�1��@F��v �1"O�e#��I�2FD����Y��2��"O����h)�խ��J[�"O����cA�Jw���e��,�:� �"O��"g��*��̐�n���F!�"O
鉥,�/t�aHTmR:֩f"O��&K�/@a���2KU'}>>(*'"O��!�mke,� �=�29�p�<I��p��(�F�E�[I�C���r�<�7�����֋ʔ�r,i�NE�<��!�Wyb�21�.s�eR�J�@�<I�f�T� )���%OD,r�B[�<q���G�fp�s 
�}��)�#��P�<YW��X:�����:gr�H�b�<���R�!2
�i�!�TG�T0�ɉt�<)�n�.L,�7g��al�<���U�px44K�O
\�;�Hr�<9¨�#����-����S�Fx}��.N�h!f�N�RuB`V�Ձ�HO�\�WH6r�y�������f"O�)���Ȣ-R��y��۽}��\y3"O��0Dِ[�*�z�T<y��Y�"O�Л�V��be<`9���"O
A�� ����0$[�#4ژr"O�X�`�^]��H֣N�|�:��2"ON咣N�#���0M�-Sb��#"O�K�	�,F�J�+ÂԝYR�`"O��3�W5q0�2��&k�����"O�ѻ�l[�A� Ȼ H|� x
g"O��B箏�]9�1�&_^�j��"O�dq���g������]�uҶ"O�L�R���,4�X�%C�=r�p��E"O�љ��W=e���)�B*���"O����k�"Ty�+�H;��7"O� �y��B+v����OD6 Ȁ��"Ojȃ�Čl}0����I.v	��"O Q��哳8"�S�$�+�dh+7"OIcW%Y��-�w㓠=|�Jg"OT����k�z��peL�1"O�ŸL"8�"�+��R�Q�"O�Kt�9R�����Л8t���"OĹ��Ɠ�o��*���,��Q"O@-yC,
A�Y��Z ^�lA�"O��[W	�����(V���y� �3"O�i-	�4��b)�~��3�T��yT Q� �����P�^L���
�yBU-�b��@U��:�	���y2��fr�i3�/B=�.4��%��y2&�~궝2%���Hq�:�yb��|*��x�"DqP퇾�y���=H��7�m��ز���y"�ӿ;�8�����"g]l� �����y2�	�_VE9��ƶ^�D	��N��yReȹ���)J ���a޷�yb��w�%��ǉ'��l�D���y���%)J���fW���%@�����yB�{�^=��* �XMd���y��֘�%Q������c��ybn߇&��R6�*~{���,�y2���lA���G`��`U��yҧ��:��`� ��h}~\yDK��y��<=��hPoD�4Rވx�φ=�y�1M����*�3a\� I+�yE8P>p0fR�/;F�	��ǰ�y"c�/N���;"��7+��d��j���y���a���c��6c:�c��ޅ�yrl�	?����J͈3��ז�y��'0�J��D�\�J\`3E��y"Kם1�p1B T��<P����yBi��B�+3�A��J��y"&p���c�	t����ݍ�yON���{���9mu�%�yBL�<�,P6���,P��B�K4�y�D˖6����p�Q$Ehrr�ӏ�yr@^�tw�Ju���
CB��y��E+*yh�kD�9�&��J��y��S�uz���ҡN�p�*��y"lA%��['�K�I|�(@����y"F�f��� �<��,�4+Q�LK��Y�����é�� qSd��Qڒ�!D���!V�nw�ș'�#3�H���bl���B
�Q��d ɿ0�9h�/_�7� 8��	���K� ��&'�0@vt0�"�� #���ȓp��i��j9~�RP4�#K9�	�ȓ>�0�0��v���[д�ȓ[
R����%V,5x��u�D��ȓ+��[�Õcu�h�lX�*�ц�	���키f�̉���-���ȓ@
���w�ٺ�v��m�%>e>)�ȓ7�������,Ё`��z"�ȓǶE)�Y�RĲ�� D)J�pe�ȓ*<.H�1��LɃdL�����#�> (��F
3DIrƇJ�&�ȓ��c��U�]��x�f E��1�ȓUz��be��	"����,�����(:1�޴|��ѳ�V��0��}ʤ�X�����2ˀ�IL����m���F�Z�4h3A�<�����S�? (�B�n�=I��	��ŌicNi��"O����V�_���B-6x��qf"OL�Jd�A�s�:��Ȳkc�y��"Ola�GD�0����Q��"Od�
@m�~Ӕ���9�x  �"O�����.�5#�DAz0<�u"O,X&&@	Mxj9�bIƺm�XBS"O�M�q%d/�] $���+$"O���KM*Z΅�5�٫>�d	��"OYq�kݓHcf�`�㉁�L�X�"O�qAƄ���@u`N�H�v\�"OV�1a�[�8 8�BMJ$n�̜rv"Or	#R,N"��<�ұ"��+�v�<�a!Ӷ��%����-���I��p�<�!'�QՂ��سp������n�<ᇠ��I���1�E���P+�i�<��N�J:I!���-X�6Eq��e�<`�R:5�biQr/�P%��(6L�<��K�4� q�	ĺkw�-C�J�]�<a����,�R��3]�0Ȳ�#R�<I��ĭ<h���1c(T��ÍT�<��԰��i��ݧy�TU��`^N�<�, 6�j��1���E;�t��eGS�<IA�.Zt�)e.W�I����S�RO�<�4�Z�!hYЗ�ȿ4��!	�O�<9a ��(�Ń���e!�Us�<�w	O��L�a��8��@bWJ�<y��bh�`&
Y��m��cD}�<�Pb�_�əŃ0�z4��z�<ѕ� .�����<b�D�(���z�<!�j&:DhY�j �68@#jO�<�F�C�0�����T<��9d&�R�<i�ԑ�\�ۦ"��,.T����x�<�P��18�3����r};�ě[�<�cպ$Kz��f?)�UK�BK|�<95HI3%�J�J2f�9't��#��u�<9'��')��x��CN��7��u�<�p��1@�L�ج�F"�E�<�S��[0 ����N���  �@�<9���U�8(v���3�@M����D�<��U��*�*u��^}�KJF�<�D��	_���m��c�^53rZ�<�C�J�mv��@%�rv{�L@W�<�5�ޠ ��Ȑ��F�A��mǥQ�<��#�`bL�+-[vm/a�PB� KY۱oT9�օ��`� B�ɨ?z� Yfo"�@��X� �4C�ɢ�"��
I2<���*�!U$t�C�I7,�(=h��ޟM��d�l�U�>B�I%�|�[��*�ુ��a�C�I�Kmh)�S(�"�X0�EM���C�	6_�t��ɦ%��� �Ǫh(�B�I2d� �8�Աg���0G�c0C��.dc<�r%ɗ
i2�\J��C
yC䉘����fG���3���B�	�q&<9�2C"V�J憔4I�C�ɊVB@�� ��N
T)q�־9#8C�I�
���@�l{�d)��� C��[|2e�F���g�������Qu4C�	�1���`�N��� ���C䉇'���!��(L��4C�¦
�B��*	+��R��x���c��VvB�ɮ|mL�8Κ�:#�1u�ιS$�C�I0&{Py����6z��f�!X�B�)� �`G��6�l�L�,NDP kq"O�ՓVj*B����L�o�
��u"O~DV�X�]�˱a��9�8,X�"O��r��<�"�2���=ۢ8p"O0��u������NP�(`PR�"O(�s�חe0�<{%�
\��t"On�<O)J��G�
�nK@%�O�:�y�8CVQ;6��;צ��GlY�yrc��&�&�H7��6�\�w䋣�yb�R+I�ZT�� YS��Fό,U�!���m5���ՅB
q�Sn[.o~��dB]�Vp17�2������
�yR!��S��HE��#�x�g�V�yS� �0!�4hό��PBi�,�y�/�JD�c��*q1�6j���y���/�F�"��z��E���y��I�~��Am��nvH6g±�y�nκZ_�p���Z�%��K��yBa߬!G���b��T�Re��MR��y��di�0f$��yr�{  ��y�@JyڝSF���:<���y���!�0�cE�66���Snی�y��H�2n�qs��(�S#kR�yr#X�v�-�vDO�Mni���yr�ێm6����U'DĨ�(�-J��y"lR�	���@��@>�iZ�u�
�'�x�@N r�&�CBş/�R��'��(�d\��>�H!n�7"3��p
�'�`��5	�lD�;��د�h
�'ֈ�b�T#c�ɫ>~�̭�'�H�I%%�$i���%JZ�^�2�K�'�8țB�>1$����BxtQ�'�ة�e!�r��)�A��}��9��'�
��`i�'d�<�Rb�̝p���9�'��*��V���Q
���f�l2�'�HaB`CP�~��4sR\�U��'��M{f@��$�TŨ6+�?�m��'`n\R%e�	��A�D]�LD���'����âW��CPn��Um\���'��zс�h(�yʏSR�#	�'ќوAg�8K�������>B��@�'�~�Qdn�2��-ӦõLB�s�'ܸluh��-�Vm8�lʑSʜK�'�����S��#c�טR�� �'�&Hkj}7>Hp��Y�Hm�Q�ʓw*̭�gИ� ���H,Nb1��M���8�/�m=Xd�7gP�S�d���e��QR�ڔ��A2J������ȓG20`Q�h C!��V�*�H0��F�̈xg�
�n�i�@K� "���M	�oN$-�l��m�$�X��ȓ'B��ZQ&�XJD�{��C5~�u�ȓKi
��P��X��̱&di��Md"� � @�?   {   Ĵ���	��Z�ztI
)ʜ�cd�<��k٥���qe�H�4͒6R64<��c�^F�Vn\�c�5��Aߦ#���y�r�7m
����4Tr�Ī<a�O�6-n��)�䈞$�p!��ʂ�#25a��8�D��ג"�qO��N<q�Ւ\�p��4�p�ض�U�
�ǁJ�d�j6�7?�d�Gk*�8λ<)T�A�9lPJ�"�<��+��D���A���a1�N�$yb�E�9�����O��C�H��U"�ݚ9�Z�I/�8]�ÏJ2���/��!j���휐U0謻L��I�; ��cGmT?�'5iR٣1��vv6-D�����%)��R�� l�$*c~q��׼����3�Љ�"(k�`�:��@�D!	�B7����s��-�qF0L�a2�c+��u6��83Dԣ�yC�"ܙ�<�8����O���������ď6;"D��"��%���,ya�>I�� �)h�(�s'b<��`��&��ry�a��$��Oj�s�A�jdZ&��5�X�ƥ��N��OFpю��߈���I�Wz:$@�E�x����t�ʽnL��~�ܺp����6S�5���;�d�Y6G4DE�9���D���O��j��L�i��fڏ2�@���X�t�x�<9�k'�
g�O~H'�7i�]в�~����i?��2M#�O* �<�1&�$3R5��o�WG�-r,܌�~b�^�~��B���ʼ���N�M��Y0 ,�ta�������q���s�/�4#<��&}b�եRbܱXfK˞mv���!؟��dڲ�O"L���$È1�����T ��R�)�2N!�D�<z �  �x�F�Q�(�����;�B��凐7*���2�3�$��^�A`Ώ�s���,�)�!�$��)^�CS�G�i��Źv��b���S���t�z�b�L�+W8�"b�'u��:d�V(M0�@�5ޜ$�`��{5Bh�Z�Qp�%k@Ӝz\\�t
�O���q�
N�H6���ݶ��xr㄀QPH:!I� 벭�� ������ �ɲ��#�J�:%h�#T�����ǝR<]j*��j�@�t����yJ$N����틁y�(x{�KΥG dA���ȰH[�n%/�rȻ��4�#�D*u�� ��([����j�o+��J
5R�D���<
# ]��� nG4�{3�X��Pȡ4
�%x 	�rL#<O��3�菃J=�Y9P�;ZM+��I��*��b�P�sn<Ej1�*cl�%��IзY��!�/=�\��%"و��x�b�k�1����-�!Z@d����BXv�]:�`����Z�*ֺ/L���t��2N_@����:,�d��`ż�y�o�3�KAl�Quؼ�s�R(|&�5럑TD��Q��y�(Ă���y�fƒZ���F��I�L�Y�x�nֲ�QZ�'�
33.\��iH*+N���h�e���27�ҕ-���ӓQ�v�p���:s>X	a�ƇZ=�i��	s?�ʘ�O5z��2�ɮ�H��t��E����E��1}t4�;�'�A��ρ 7-�)��'#>�b�}"�٨O.XAj͞GQ>Uz���4=5]��)�b����D�!D��aDE ;�hL�R'P��8�H��SP�T���t���G����A_L -�T��ǯ��:�Di	�'�L���c�	0gF��R%Ѳ9Z�@ɔ9*�ƜwnĘo��{��J�@n4T��4]�������=���t6� ��'��S�*��Dk�К�ۤ&�����'��);�f֞bI�|��/�:Gej����\-Z�~�b��h
l�gdK+_Q֠+b�QH�<�A�I�o�`�� �է4bE����A�<Iwƚy�ě�� �v�2c'�]�<��ʗ=v؊X���
w�¹��hC�<�GɦJjh��hG-�ν� ��A�<q0GK1@������a����6%	u�<����Q�uK���*"�(�`� �J�<���Q�R1�o�#d�����P�<�T��ȩ;e�?ez|8Y��b�<s���Q�\� ��9<��`��SU�<A�
^��b��dB5j� 0�#z�<���N<;p=�dɌ�=��|��gMt�<�1��-v�ӃO�7cl�!��r�<�uO�(#�Uؑ�ڇ[�`:F�M�<)Am��P9����េ~TF����S�<颋�mV\���Qp��s�&T��8��Qm����LE�3�a�C�*D��س��u�"�ރb���!$��S�<�A Dz"\t�w	�I�L�(�m�<a̅2���if�X����Fa�r�<Yu�͌Z�u	Ι,Rn҂�y
� ��Q��E74�&�S�
J��ȹ""O"HK�H}�=�bjW1E�~�u"OJQ��H T��х��)3��"O� ���D�Z�D@�l��Q�U"O��4�Mc����v蚌���z�"O>���!^�9�vm�oT�o# �k�"O� C� N#�>L��nR�"n.��"O�Fe 0]����ZI7���"O,Kю�p����!���"O }��aٕr��;A��7!����"O�p��ԑ~`�ux�(�2�A��"O��c��:Rj68����M���"O:�+!@ƞy� 	s'��'����"O@�!Jɬf�hI�S��'p��"O`��6��� ��e# ��%b+4���"O���F�JT%b�
�3Nv�EHv"O����`3}݈1�e`O(Z� ��"O�\���	y�(�ᬕy����"O����I����G
01̡� "OF��
�!fh=���65�`-
�"Oj���2
ܑk�C$d6	Z"Oq���3i��0QvC7S�
2�"O$�۔$TJ��Y�C� ���"OX�9��7�r����H2R�TH�G"O&1@��@��Ӆ G�B��Y�"Oh\��K�}N�\c��� ��y%"O��9$Ws�Ƭ�-�<4��3"O��"��<?r�ڰ��	2���"O�=�¬�-���8U�ϼ$t���s"O@����=1b
	� &C��}H�"O�y0�K^�<\3�MJ��0K5"OV!p�吐ZH<4����h5V���"O0t�(*W�pA��>=R80�"O�� ՌD�k9(%ig�%1�ԁ�"O�-�W-�:dxB�C�E��W"O^D��8�X��S�P�$0�"O&�!5�^',A��P�ʼ4�D�A�'x�M9AnN?�0t���:>:x`�0C\�C�I�Y}����	X�]-�P"�m
�4C�ɥ6��@�T�˳R)�izf耷G��B�	�l�2�)��s1�1{�N�1'y��DE�L��!/��c�<Q:Pj�IQ!�Č�kj\��Cσ&�@W_�RJ!�dE�8��@*���v\� ��
/!�$�20�H��-�=\RT��RĐ�w%!�dI*B�.1㭆�,:ޔQ���$q!��O+���)�r�ĴHc�B"G!�D���;F�������"O@yqU�ֹew���f�b��"OuK������r ^�_��1"O�ǃؤ~ �|�T/��5��LI�"ON )QK#o���a�ę5����"O,=���T49d0�� �P��Ji;�"O0�!�B�=;YT��c�4d;���t"O�t�Da�-9!3Đ.v���b"O^�{ �R������=
�` "O�zb�_�%7��i���r��=��"O<��*t$��`K�V�5[�"O !�A�R~�2�Bǌq�`��"O�9����	�d�қ� m��"O��TkB�W�=Ӈ�Q'{�pD�g"O�tB���7��-؆�TS�p�8g"ON�a�:"�:-�R��9 �� )T"O���L])�+pdC�����"O� �X��hD�+Q��0
O@�i�"O�)���yI������*S��{�"O��x@��dd��C-Ou,�ۓ"O2d��-D�b�s�� h����"O��y�m�+m)�$���ّP���"OԐ˕�^�@%��;Lf�	q"O��ꒁ'{\5)ٕk��L��"O��0�ДvXđ�#�,y.Y+R"O8Tb�"�3[%X�
�rY"�C"ODa��9n�HXB*��/�̐��"O��)F24^t��#�KOb1�"OFt�uIݰ$��B� ?8��"O� a�]=d-f���@�cI�%��"OBP�"���t�{��R(*8sE"OX����62% � Sh
/)�h�"O�<�Ɩ0�dg�_/3?���C"O����
�T,�@U�A	�"O�}#�#;��C�+C�/�`�"O !h�)ة��hh���#��Tڴ"O\ðE�KP�� �Q���:"Oj�3�9�`I���1�"��0"O��bqn?P$.		�,�%b��B�"OF]��O�fz�h�s���X.6I�w"O^%Ia""8��-Q�67��s$"O�XZ僗6'�$�O�Ũ��"O&`�� ��`�r�r�D4PDp0G"O��5cNppP���wF T��"Otȉ�F03���u��4Z��c�"O@�,��`���0�n�!MQ��2Q"O�Q���W�m��H"��J�P�&L�q"Ov0�%IT�WfZH��,K�jJ�P"O2�Q���KY�5�k_�yL칑"O���ݍ#�~�p�
�*/H��"O�h��'�-b���p��82t�U"Oʕ�f��A���{7�]+.�Z�"O�X���P�衙FMm><�6"O4y�$L�eR��
�琔��r�"O��s���E��
���8?�]�&"O��J����f��#C2���4"O��k�N$]hI��JA�E� "O"�{�@)z�A	�0_���B"O8q��J�P��Q)ب6XZܩ1"O�����K�QXR�N�E��"ORP۷��4lp����FG/C�)۔"O�$�QJ�F{�,� �i.�� P"Of�g`��4�ȡ�)�]`<��"O���`��>3��y�)�4n��)�"O�d9��� o� �a��/Zt>�c�"O<@S'Nt�����%S�"O^-��@ݢN8�Mip)Bj��kc"Od���*M!$��|��I�a���i�"O���H6��A9#�ʝ:`|X�t"O��8R+�";��1�O2gJ�݁b"O9�S�T�2oV}� i��Y1�ġ�"O|��㣉7�<�b�Q�Q@f�E"O�I��XQ���s��5(���6"O���' �qv�E*s�C�Ov����"O��@	��-�6� �%P�8e@qKc"OQ�ЉCB��%�Y�t��"O�S6%�	 P���k�"O�ps�C#�4`[V� #�F\��"O�yRUnH�:������w�I��"OT�a���5&�f"G�I�XQC�"OP�`o#Qq�0�BшT���ZT"O� �d�դ�"�L�"�d�6�{u"O�4À�D3n����3-�rܰs"Oȝ�5b�rB�#N��!� �i�"O>��� ��Ǯ�����;\��p"O����57x�Ƌ�"3�P)"O|I�t�A�)��b��]*��Rs"O��A`@�'�Z��&i�
R���"O, ��e��S�J�����r���"O0�*�#�.E�lF� �V<ʒ"O�fBҙ^~<e	A+[4!TM�c"O4dq�������"��rxx\��"O�9��R.Ȣ�RT��8gH-�r"Od��t%��~Y7�·vf�l(e"O�%�ɤR��2o!CE��C"O�H2U�[8%�� �$. �v8~}� "O���\�9���Z�N�x/bɈ�"O��Y�1�F�܈R! ��'"O�LJrhբŋV�q
�!*7"O��sZ�u�F���x��cc"OVL�1�J�17�t`�@)7�jh�t"O���R�AD�"��͓g� y�"O���՞�2AXd��6��"O�e`&M4���-�S���"O�Pe��?�b�cKx�+�"O@�bDK�;0$�@dĜ)[��+r"O�������@�����*q���+�剢"�a���:3�������b~��F�K=�y�0K2��3�I�R9�0)���<�?I���%m4I��^�W�6�Y�i`�U�ȓ:-�=�ba�>�$��vb�����'^����F�U/��p���h⅑�n�d�@�'��ȫFA�2'�T�dXj�,i@�'0����� �V�R���7-vxEa�'��!;�"$�l�� ��#3��10�'���0w舦w���XS	��+�6`��'Y�1� )=���d��%Q�A�':*�`an_25瞭�A�٠�0��'�BmX�/מuq��"`��>4x��'��*G��h���S��V�?5`���'�p<�� 84��P�U�8�����'�@�X���PU�T�!!F�i	�'
Ҝ���YÊ�ԏ�������'|}�#H��&�}'mג<|a��'\��v	y�2]�n��R�N��'��%є�W�r�Θ�)�#<��+�'"jMbp<��![� ��0�d�'�pQ���v֦8��E!��!R�'��P��-.v\#mMml��p�'����T%*���Z#f�j)�
�'�P�C�)^��%�"FZ3N�K
�'+�e��j�
�.u9�"�ZfBX�	�'�F�6f��\��9)Mc.}��'���')���n���Mh�
a�'��%ص[��
@���_��9!�'���H���%z��gJ�(Q�~0�
�'O��#w���-�ɛ'\~^�
�'�N����`5Ƶ������	�'�&ػ�w\@���J̆|ݲ���'�%Z�q�ʑ ����|�8Z�'���	���(��������np�'��t�F�����V�
|�P]X�'�0����� l@�Y5
J3qq���'��@�u�?L��1h��c
$��'�*)�cY�v2� X�ιiϼ��	��� ,���1Z�t��Azq�2""O&T" L���2Y� f�/\E��"O&�1KV	Gp�������RZ5"O�@hvj�&x�)�c0�^��%"O����
�70ѳA��k}����"OȌ@3�U;��m��@:�4��"O�T�'n'<<�%/������s"O9����(���L�~�>L* "O���IJ���Y�K�c��!a�"O~��FB�I�2�20�X*A��9�"O:š���eC��ꠋ�R�Px"O��"�.s�~-ȵ��?H��p��"O�)��u�͚�Ȗ4N�B��F"O�q)��N1%��X�ٛ3����A"O�����n��K�fR$%�b��"OX��F@�w��-�Ce��I�f��"O���e��rX�!vD�W?2���"O�m$�Kkn-�0�b�|�B"O8�sCD�7�����O4.��+�"OZ�����^U�A#��U�r��upc"OPeBcIυ8�X	�`� X��m�"O�c���Z�`m�@���"O����EՓ�����O�jg�Dk�"O)���$o�J!x$O�*i?���"O��8	�9yղ�s�Oޒ:P�"OȹV�@=&��$�� =� ���"O&��)�P�9s���$��hD"OR!��Ɓ�@b�(2� ����ð"OppX®�+X�b��d�G#+�AC6D��;'�h�$X��F�]�b��U,6D�D�k�;^\�a�gƄ�zt	6	7D�@�Ri�!wd��ABqaV,���4D��*���6Z,�}�G���00��1D�!p ��em�бa�����1��-D�АB�U$@��E�$-�;Ǭ5���*D�SBI2jn��ȳ���x%��`'&*D����R12�IZ��"-�����)D�����(sO�qh`�=X^ġ �.'D����1�$|��!�T������#D�瘛.{�X����2h�<$�6D�D�&&W*Y���Ԥ�'aPЄ6D�Hڣ.   �P   �
  5  �  L!  )  �1  �7   >  zD  �J  �R  �X  ?_  �e  �k  r  Gx  �~  ��   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl���q�6O$���'h4�lE� �]��P��v�J�hJz��u�iЛA���!2B�Xu	pݍ �'�?�"��?�[�O��A�� 
"T��'��>+�kJ�+��93�!�eglUٰ/�'�uW�ǒqC�T�'Q�� �cS?H�PU�㫍=d�өɅQzT�4��O$5�'�͓Obf��R��%QS(H��$�I��D����X� LX؂y+����IK! �П���l@��
0!Gey�'��ٲ�O�r�'& pv/@��feQb'��DxZ�:�'�"�'t��'/r�',���u�i���df���
�Q6�x����|p�H�b�%�OX手^^>�e!Z<Z�
��-cP��O<���PV���Е?�q�D�-�ؽX���Gi+ၴ�?1��?���?���?����	dޕr�(q7�`JG�t5��r!�O��L㦩��4h����'&p�ݐVj����4o�\H������CN	�潚��
�3�>����V���y�Q?9��R"[�A8 + �c��R0Ԯ]z@Pj��9�<�rf/[ᦡ��4|��F�O��A�!0d��FR,5��Q�NP�c� ��$sU&7M)iӂ��e�ˋD��d�I/]j���&-�*[�J�lښ�M���i��}2f��pƊ	�Ҧ�;@�<!���H�c�
h��.x7��禕#�4Oؾ���&c���Q�.�3�g�V��M&T&�ɣM��t�"�id��  ��dv�i�7-���ջ�a4#y0�0�.L�4^�y�M�C�ʰ���ijV��	 �ܴcq|=�vh���JEǈ�@Ũ�#�'��O��!pH׽>����C)�=!���Ot�$��֟�y��/�Ms̟�4����%��0IM#(xF��W�'�����	�|r�/�S���Ш�'�4��I><��(�2#S�c��8Dh��gjL��	)�R��e-��{�̼�0Lßt(f� �D���)`N��c�"2O����'!2�<�D,R�q��b�`�Yx4��7�Aޟ��I���?�|��'���嫃)(|QĊK;~p���b�i>�*ߴx�U(A���Rf� bh�1v[b��q�i�O��ȣ�$���?�$E�As�M1���)�����"T�T;�i,�S�������ȗ�<D��b-�G�tY��[k��� 7@-D�Pz֨]0X�L�/[���d�a'D���Bl�2b���ا.4�L�B�&D��[�̇ \�̈d��KB� �T`�O���O?�(�K�a���j���-0
U��F�<���L�+'�X�����*L�<�2*�y �s�K�	�^��b@L�<����6+Rx��$)s��ⓠ�l�<��aϕ�ӪF p� ��c��c���D�Dl M0M�T�P�	0�(=����P��~�'�"�'X���'r�'s��qAc�"�rq��� �/��@2�K�Xk<� r�^��0���%<O�PA1�ץ#\0����-�T	��m�9Z7�Y�bEH�b:ˎ�K�Vi�%6*�ў`��e��h����CG�x.�k K�5(8�H����<��O�CK:R�:UCUh�)�p� ��'�!�����쐘 �@�nfm�C�ԵW���o�����a�4��ȨnFθnZߟ�ϓC����'��a���YT2��	]yR�'_b<�&}x���q"������@��L�,�T�� ��ju��4�ˊO1X����>�jͪ���:7����؍_*��
�ì�b��"LX���q�'R�`(��?�Խi��
��vѳ��M��(��@��-���ڟX�?E���ӭ{F�A:ӈ�3K��tX���(��'�퓻�M[!i�2��3�_/7�0�֏"��v�|���D��0�����䐵�C2s��#0o��JA�(P��yrb�?]������^���)gC��y�͓.n?@���*��_�jtpc����yB��WWN���U�O�J�����ydK'I!�E��`�
�:I{T�T$�yR�+V�n��%وv:���bM�_]���|�'��2���'���'n�	�1쎁�W�ԒZϦ�t�^�m�IգG%����.n"2��F��^���I) hD`��ߥ;�T��)��N_.��&J_2���Fc�"��&$.�V��!��OX����¸��9Bi��Ni�Lp��uӺq�'��u����?q���?i���),�U1�	ƙEi:��6N���<1���ԏ~>�����¨^H�3���G3B�'B6-��'����?�'^�*�,ͻ8ł��7��CFP�5"��%��6M�OD���Odʓ��'��p�d+J�|��w䂺`�P!R�@�-��7�N�M+�2�?�DQ�@O�d�$8�eT%$��@0ǌ8�z$A'�΋X2�ɇ�ɜj=H���	M���Q��n���p}i���O��m�yy��'R�'���'��S��>� �e�?�l����X��8B�	3xR�	j��ѻ1V�(g�H�k�,�O�lo�џ�'vx��#eyӚ�d�O89{�-B��(�:"�����Ob���!y����O��Ӂu�B�D.�)� x�t�^/q�}��A1N4��J`�'��9ʍ�d˸/��j� �y@����P�o?axb�U��?Af�|R
�/:Ӧ 1Cŀ� ����T7�y���
#����+F�eO`���F��?�d�'�D�ْ`�/\?�@@aM�od���J>��kg�&�'�_>ps*�ԟX�vi
51���B���+W��bB�����.]��r������Or�'��*y���xB@-/�h��x�"�{1�q��3z�x�C�ӡ�h�^ è[$|�F%�ЖzCv8a3���R0d�OV�lڐ��O��6�m�gd�!nÞy�m��C��H4�'��'�	 ��S,V l5�E�ƢW���=���;>��vy�9��rv.M5"�X<���R��m���z����O��C!
�(1��l�O����O��fޕ�A(փjjv�@O
,a0P}��'��� ���` J�?��M/.�H�2�]�^�p�,�:|���q�شq��ǔ/ ^-ˏ��y�II�=���Y	�l���Π�?���i����A��Y�����ID�z���df��!#L�x�G{��	������Ù�:��'�?z��`w�П4��'����<a*���$�<P+@}��K+��G�2�[����ib�A��B?�?A���?)�D|�n�O���q>��B�-QX�%���ض��� ()�C�ɼf4E)��'���zDǉ�*���a#e3�X	�#P6`�!Ъ�p�h��2/S :�dAU���ȡ-bߊ�փ��/�р��8D����B�a�tÄ��Eo�H���*�DE��%�8���M����?�"��<w��U��d��>TRI��!�*�?���)ɨ����?�O������'<���&~���.ʷ2�}�	Ó.��aFxr�ٽ;�a㢋C�,�Ό:�(�0<v�֟D�N>�GD��.��Y��b^� �)���`�<�H֊�0�
�C����բ�Z��T���V���ȗZ ��W���|2�U%����f��M���?!+���)���O�@j�7Q6���q��)m��c��O����)����+�|�OP�q�%�q�x�ީly�Ñ�8��2�S�OH�`	�bGbS��ˠ6W�EP�O��:��'��O>�®8/@�<J2m�3=��ÄB9D��z�� >��<�L�4��+��8�-��>U���L;#ߪݩ��$&����	Ŧ��I某�I�)�D�c��ڟ`�	��D��Ӽ�`�5J��h�E�O�9�G�����f�P� D�ER�g�gV��� )6t�^�����3{u�M>1�	[���|�<a5C	=:� !a���'��ҟ@��������䟼�|�'<�.��=�ī[5"�ik��.!����>6Ѹ���fZ`�" �O��C����ٟ��'��*4�E?>�.X
���Y�*���ɩ`�\6��O��d�O�˓��'v��"5�(c�p��Č�C��#�i���b�'��Q��E�:06$IkQ�y^a�+Z1f5ve
�M���9��a;,On��g]�k�\�1��A�-bjH�jE e]��'��6�OB˓�?���B@R���%�P*�>!����%����L�	v�D(�� N_��ͳT��
:��'l� �>�*ON(rU�ڦ�I�<!�I�V�ĉ�Q��[x]��B�ڟl�'!b�'���AD�Tp�ғl7�!�6O�(!��R�<Q�M�H$|?9b��'��a�ai�s�u�� Ow|6�M&CF$p���j���]�Ȑ�Ó������M����?9����F�t�R(,�P\��-�?����?���?!O~z�y�J��HA҅%��"71s���'Lў�ӕ�?���4MHJ�HTj̏(������'΀q���l�J��|�٦��I4>6��&�6Gh�}p@��J�(��I�$���5�~=��.0_l��	r�'NT<I5��#�����,`x(��O΁P4�
H�&�1C�J���dF�D�ğ4�	��#F��ur�Ի��0Z�	��Ms��i1�S�-�t��,H7B.�R;֘cSc&���O���&�S���^$P�	�F�ͨ\y�WI�'�iuӚ�oU�I�I;rY	�Bрl���%���	/jnE�?�g�'T�`&c��a�\,˴`DM�f�`�'m����B��1�D�L#����'�"�z0(�1s�,��n��J	���
�'�0��*X�L���sgC/F/|Db	�'8��@�Ro�a���AdQ��'p�}C@�W�<P>�S6'	�H�6��/O���'ۦ�ѷ�>\������������ �̩g�R�cΙ�Cօ�JA�G"O`�����r��1q�♐�l�`R"O����^u�գP�@�e�$��"O�5�E�Q&)9� �3�k2�r��'��(��'? P�pÀ��bUA�k�'[���'&<�r!@W9+�0A� �P$��'dn�B��"ܗZ�zHä�y��P�7��i���L8A3����y�FE�N�X(� ں�0��U	�,�y¡T9A�h�M��,n����hO��Ӣ�ӹF�T�ƌ�Z��9Y���P8C�ɽj�:����~�5+Ӌ
A�fC�I�2@D@ūS�lwR�㇨QG��C䉹B�:��W�Ǜ�>lR�P
#�C�I#e\�P��Gy�.T�)o+�B��;$�V�04.L/
� @�+F́��?��,G����V����}�@k�J\ol�`m&D�cW���,�N(�C·38���1D�I�GZ��q"'29�����1D��Y��3���6Co�M�T�-D��1AOU!4N�d9�i�7!��S-'D������7�^���$JP���<�f��{8��7!ݤL6>�sE��o2�'�#D� 2u�V�=�*<�
�)ap���?D�� eb^�C6���͋�0�u�c?D�$�,����يS�H9=� �n:D��a�;|E�JKkY��X�5�O]��O�Ͱcf�9�����.(2Ub�"Ob���ʌh�v���.F�4�h"ON�Q���E�a0��ˉC�*��"O���5L֓Y�d��b�����F"O ب�V�Ͱ�9!�P@Ir"O�|��-�jj�����.c��A��ɠD`�~ꅉ�		lbw��F)0�%�IX�<�&+C�}� ��(��q$����H�W�<��	Q�K��X+MH���sS�P�<���H!k[�U !K�I3�h[ ��H�<�c�� ~��Z�.M�;f�1[!�B�<)0D�2i�>D�l�8�T�؟�h1<�S�O�0{`�Hz�=��G4";he��"O���Q��1>�.}(''_k`�ȥ"O���"U�w���	`�p!��"O2���CҚ� ��  �R�R��"O�����^gj�A�&E�1"O��y�ㅍPG��t���g�:�(�S��b0�,�O� �Q�t��N�8
�+�"O�-�AH�:����b�9O�)��"O��DGȋH�Ay�B#5�<\9A"O6bw��W�$,���+FOV8Y"O���#�B�@N�{q�҅^4��r��'�HY��'0bA
%+�M/d|a��[�Z��X�'Ɩu��*�P�Ra[rML��(0�'5��*@��.?��Y1%.�I]�-�'[��)'��!ʮt�tCP�6P��0�'B�a[�L!�
����46���'�Tq���~F*T�U��'z��8���*#Q?=�3,�Or�0����![���0�.D��:1�	8t2Q�a��]L���*D��(�DW�cqTȫ]�?�. +�o)D� �F� �5�:�rt�M O��1�%D�<�� yd��׮�V���b�0D����bT6o8((8�`�W��-��@�O��q�)�Q��Ac� @%���)X�c�Z�C
�'�f1*5�ϫ)$d�Sd\+pF�yx��� ����Ȁ�h�QH�D��D�4�@"O�s��1�5�t�� ��a�"O@�8�A�����?=:(�"Ol* ��dZBI�VE۴b"\]9�]�����%�O����!�~��Ӯ�5&�9�V*OJ�Rä]e������T��r�'� �:p�������A� �̙��'�l�r �P��T��`\�k\��K�'	6D�D��2+���p&�)j�	9�OpԑU�O�}�U!�*6ZQ$�u�\��"OX�q�Ӟ[#�<�� ӥ��}б"O���F�<�J�F�ʘ`j�"O6��EG'�:=j"�>�� �!"O*�R�H�&g�h�Ȕ �N��q��"ORu�㍞;2?$�⒡�&��X)d�I+b�~��F�)x�0U�FԄ/B�J�(Tt�<�VlIz���b�
_���q@�i�<��Ă*��2!K�����qA�k�<Y� ;F���Q� X$��a2��f�<	�D��Hw�@A,��#jjxQ��a�<���U:y� 쒁�./���3��WןXh`�=�S�O�pAM�c�2c���<��X4"O����O��v\����0Ö٣�"O ,2Ui\�4U�e�bͳ9�nT;�"O�x�(u �(�6j��{T"OҽA���;�2�2�� 
��S�"O\�����a!�z�䖐0#�^�x��"�O���@�K��� ��)Y%$0�"O�5�1��I&zXc��U5� �"O�(�#E�c�����x�! "Oz@c �-��pڰ^;EJ2F"O8թwn�3hʸ��NX�{�\R��'�(���'t�����UP5�6�W)L\�q�'!�]�G�Q�}ZȌqv�1�Ĉ�'�.P2���#p�F����|�0�'MR�� K��\;��.wp��
�'X\�&I�?\�`��Y��Y�	�'��j�K|���h!��PPH��Ě�zQ?݉e �?Z�M�b%��7y<�!ҩ$D��b�іeh�BB�c����#$D�T��Ş8�,�H��N; �e/D��gl#A���[E^�w����.!D��цޕYU�5:A�ϳ�X����9D���En�κik#HN:1X��#��O�ͳ�)�	����a��6e�0��E��"O} �V�d!اA�,Q�r��#"O��E*�ҤpT�\�Xm�"O�m2�#7Q��#A/��c�����"OF����дl>��C A����"O��&ED�><y��ݲ[Ԙ=�PU� >�OZ����K7z�ر��($6]J�2d"OF����97�� su�֘KK�`;�"O���Q%�%]dI�3��?�m��"O���3���	���Fϋ?@���"OƠfi�0H:ĚF.,�f�'����'��h#���W��$���ۢ�x�'N�������k6UI̎�VR�1�
�', d��i�I����Tj�1a@ <��'h�IP�E͈I��d ý�L-��'�|�D�Q�S��p�cb��}��|r�'�\�$���D��l�C�)u� ��䉃(�Q?e��
�8�"���I2*&���ӧ'D����Ѭ-cNqba��27q�y��$D����؊}X����됹��) �� D�� R]C�G�B1����KG��X�"O�)��H��n,B��ٯ���2r"Ozq ����$ <j�h�V�'nD�����;;�2D��
��O�}�S
Y�Z�pЇ��P�Dځ`S�)3�[�t(@U��n~0H�Q��w�t�b��/����{tj���LĨ#4�TBtG	!'Ji�ȓ'Nl�0e�1,����B��M����ȓ";�auFE$0����E	�@L�'��m;�*��hZ���hj��*�(<J���H��ɁG|�j$F�"@������[��F�L�^Tв��OE��ȓf$��P��)K:PH�%O+�p���+ �@���.J0VlzS��Co�؇�I�<��I*Bqp�J��i�p���-�E[ B�n�$B��_�ZXf���/3L�C䉽/BȜ���5�@L�ᆐ�Y��C�ɪYҪ��p���w��Gg�C�
q/�ˢ*ƿP���ѕ�W,F�HC�I�@\ָ
��xT`څ��C%F�=�b��h�O�F�y�Ҋ
�ҝb���w���c�'��x�F2a���J7�C����'�S�?HF�q��`F;�|�
�'�p��������h�`ԂJv�#
�'�6��#ػ�)�r�� ��-K	�'>�A���ڄ� b�D�~`8\{���T�Gx���[����L���S�#�^B�ɿ'�6���
$��Tb��E6�LB� ~`d`�A�X�/���ru"�m$FB�I�2\���&ƊX�j�+�E�l
�B䉚Y7��������H-����?tPB�I7Z��	�蝈VY������c}f=�	�Aq�	 Bv6��,^ߢ�a �K^wk��O}��H��m׮�zѳqS\���'˜�Ӷ�'�2�']by�GJ�#}�b|2��]�KZ�	lz>��� �!`�,e�g�G�c��e)�}�8X�
Q���hA��ЎMɴ�v!� tR����!�7m!	�킈L�FXh��DQ�%:��'"1��X�6+���!U+��k4ո�
KAyr�'a|�B\Xm���\�/�֥�q�D��>1�^��ꐫ��&s:�v�?3���Bi�<q%+��?q�ך�?*����+����G�-�b� �J1�����=C���$��iu������]RwN���ʧ��O�T�H�Ds>@�;g̳i���қ'��yŉ7��Eʒ0
��?5i �=�Ta�IL�KFvyI'm��ȣH�O��$1?%?��'���1�� ޠ���̕�TC�ԉ�'M^X�S`9>��h1r�R!:o�I��Ċl�O}��8���4K0,DI�OR'oBP�OW0\$2�'#�lA�Aj���'�?����?9���D��nL �a!��5 :m�q��$\&�@��΃&��0�+G��D'=2���R�7PЁ���_�a��q���	N����P�P rt�Q�e�g`6pF�?�ҏ}���<�Q'���(����!a�����\�t�'kў�͓3�v�I�-Gl���/�����[���P$h�D��r�*��-
=�	��HO�)�O�c��`T�<������K���O�0H7�'Фx�r�ͦ>g	��ZUTT�R�'I�`�#��*�Ԝ(4��c����	�'7�@�oŸY�ìɥ^�Vd��'X`�P��q��{�Qk�,�
�'OR� ,K�M>LU�3i��eǘ�
ߓDl��O�yآ�.�T�X�М=�T���"O��Җ�B#���B2���9�"O�|�Ԃ��^m�CW�,�T�XT"OȌ�EJZ�`2,ٻM9at^Q�"O����3)>�9��шq���"O�؛c�PB����1�=i7�dX��O9�\'$>�fuk�%ly(���'e��!��n9h��։3�5��'^`�r%��{��tمd�1�Re���� ���+F�X��-QFA�LhBX�"OP�H�L�Ԑ�j�l��q�"O�I�初<4�yx���5��@[�)G�O΢}��s��&J_x]��
=j�t)���nTy�GS�I!�eq�A�<$E���ȓ[�E3n��R�D����=n;``��fx=��ꑈ��q�7�_7Z�ޤ��,�"��a����1�EjN	I`���b
�E��_?���F\���	�'����(M�M�W�a�W����B䉿p�ZDE��+6T�5��D�Q��B䉞[�j%��$@v�cr�@� -B�I�k�P����>3=����6lQ�B�I�
�*U�u̶}�䌳�+=tlN�?Q2�ڜ0ڛ��'��9�����+~��C��*6�V����'�",�Q�'^��'�Jh���'1O󩇑>�6�Q��A7\��$���I�8�'b�@I�D�?�� ��ڤ��$G|2�(�?���)� ��bU���J-F�Y�E�(%�!���>9B�����Q�f�(�# eJ{��}�<A���4A�(�W̞;s��*�K�iy��'��[��O�Қ?�'/�%M�x���ǎ`��e�2�%�,��>�(��{L��똜O��3�(�	���$���U��4�1�$��([8ł5������|6��Oe�x�p;u��O����Du�� F#��Q�؀�T)��ꦭґ⛘]ҬlZԟ(PuC��xϓ��M���]�����D�yp��V�H'jQhO
<#���?�u�!��'.�N�O<�$�����d���r�
�ws���D��8xVL@jAɑ-&V��O������O�扜tr�s��n�K�ta[�L	H��E�:�l���G��?QP�����@�f����~�d�O��9Ox8@�B�4� � �Y�5(���şTs��Ot��^�fV>�dv�4� �?7��h��/��B�@R��M��OO�O0$�n�<�2@�ß��I$P��'�?����S*�,]b�#D+��"�Q�m�)y�dtٝ'�TM����?I���p��p�\�g��?nڮ1;��h5�
$s+�)4	�<����s���$r��O�O���E*gs�ST���V�̼z��G���4�P�̧f��l��4V-�U�'�����?����?a�'�:IњO/�<�GQ�a�&� �/�
&Ĥ�ڴ�i����'��韄�)�>���	d���c>[|"4��|�<i/��oJ��s�QF�Rv��i�	ԟh�	Пp�	�D�I�l��56�I�O�͢��Ƕ"Z������M����?����?i���?!��?���?��i�(?ư���� 2\���%Q�m���V�$��fyr�''�gy�X ��D,����q� �y�7� �S��MK��ۢedܝ��b[��>u�a�No}��'v�Z��K -vy��J۱-��!��'`ɪ����4�����%r�`�
�'R}�q艇V�l(�0��>7|��'��eM�J[d� ��2m�,��'I,��,G'c��r��BJ�ea�' E��]"B�*Z��#�%�y�)�""�B�yG�3N�`[�F�y��*9F����"SL0�M��L;�(O0D
�'t�Q���Ҫ,v8J0$E����ȓb��9a��7�H�����>k�Pe�>����3V���E3��Ԣ�#�H�m���Ku�i��.�
+rL����
W�l�[���P���@p��  ��L���0	�6(�>C��a��kݜx����d���:�B�='R�l��MNf�)R��I?����0�0X�藊T<�;�U%7&��S��|��?b|��k�/%#$4��enO�u��B��^�`$�]�"}�l�EϦmRB䉷W��h���HW�X6f�+hB�ɇ`���pt~mI)�H�JB�I�7�����D#$�Xaq�`G>U�>B�?�&��Q��>9�4�[��B�I��ٚ$�H�;g�A!�,`/�C�	=$��ᯓ;JĠ��4; �C䉕#�� ���G�f=�%9�� ��C䉾?�H�Ҷ&�0{G\�]Fr`C��U����Q)}��K\<X`C���V9��b��=����}{�B�Ɉq�,ݛ��&֨Đ��(vp*C�)� �p�O����� �텲9�V���"O�E��K�=�1���4pA�xH�"O�񪃾R6Y�g*V�cP쵂�"Ol�҇'M���I�1��cMj�q�"O��rvO�FȾH��;"N��R"O����e�D�\m �MI�����"O�HbP�h��u��M�U�� "O )���0<Az��b̒�Y
L  "O>���1\Q.�a�� !�@��"O�#Ҙ#���"�>Y<иk�"O�p�
Ѧ,EإKP�T�h�X��5"OF�Q(J�,�D�󄃿]��¦"Ob��#�J�7f��#�#?�a"OʱRO\�r58�E��K+f�Zc"O�"�\90�䨱C��&��ӵ"O����e6|��kc��!{�\j�"O\`�&eȖU�������X�SF"O�xY�)#�`I��C"ߤ�4"O��TD��h�l�@�>#5��+�"O�;�jY��ꕳ���4||�B�"O�T a�-����S�3�^��%"O�q��*��� �e[�}� � �"O&aJŎ�4&6��F��}����"On�Q딻iNl�P��1�$���"OL|�c��o�nh����?|��![�"O4$�'��<��p�թO�V�ic"O�5j'k�@M�lIt�����؄"O�i�;#I�y���Q�lp�3A"O&1�FE1~�6\�7HO�*���"O���O�h�d���P�� )t"O��t�"��Q�aG\Q�����"O"Ȣ��zjA� @�C��x�b"O��K�C�����L�pz��J"O	��!��^���i�9�6T	t"Oh�s��;|�:��G�q�l�T"OĤ����f�ld��F{B�`a"O����hD�D���ӆZ��-h�"O�8��Ņ�|I���QE���NXk�"O8�C�!IJ��G#P�uh�v"O��t-�NP��DB��DB4�"O�P`��.;F��G�\�)c���"O��@J�)H�.�bS@��&o>�u"O��(Dj��i�~����p���$"O�ZAǉs^���)�H��"O"xC����/�y{�I�l�����"O*xC(A�5����+V�JQ"Or�ڇ凊0�\�$%	��� �"O�s�NQ��ZD�6�>L�j�"O^�`b@�l�9�g���00M�B"O	Bwn��r����?�Bق�"Oր�FnV	6Lq��W�^��MP"O(m�ᬍ	��`9�k��E��;!"OhA	�i����5@��G�]5�y8�"O��0 ϯW�8��(L�Ѯ�H�"O��z#J3-�0+DGW�Y�����"O��8P��F��*�[�6d$�"O\t[Eg�D`�A,�j�2��B"O�Ii���15&!��	�@F�X"O�(��K�`CL�z��Ύ0
���"O(T;&�&YX�:���.Y!T��"O�A�G+�k�= `O�Hx�cv"O����&w(��+�\	���s"ObHR�f��6b�P��*{b����"O�x8��Ѕ-+(\[&�B:�1@"O� �T�� �W��L���D$:�X۶"O�x�@͝8J�@��q�7!�M��"OJy��_�2t)x�D�*[┸"�"O�Hi��4.���s��;Z�2a� "O�� I�$�*�qe��+��,�S"OL���; *���Jݗ%��L{ "O@h�`�γ=��(�J	p�ԨS�"O
$�0LA�+nl�ôn��*�i"O.᷄��08�%���>g���y�"O"8�0���5�gΓ!�*���"O����z�ԩz�g�U[Xh2�"O� 7IW={k ��֫ЌF��j�"O&���n�D�|T���=%7����"O�UH��U�X e�{%�kw"O\q�r���Dx���7,����"O��*s�ExM
����!:�4"O�-��M��0��S�(Zu21@C"O,:�Ĝ�!���b�O�rp�s"O���8,3����kY�`@�x"O�8+f��S�.�(pKB63=6"OZ5��bCkHD�F �l(F��$"Or\�����s�|}zq/�F���"O01�$��nr0If�ȼN�D�
6"O���"@�,����)4����"O�	�JL;Ib4t"�eP��f�B"O� �����^8qJ/ǜ]c"ON0���ګ̤�cHB� ��QR�"O���b 1;��T�6�X
S�^8p�"O4�	�NՋkWzka� =�F<R�"Oh�c��x��Y�$Ň,~�� "O���.��e1M1CT�Zh,I3"OL)k�{4��ro6I<M�T"O�8�ѥ�<+�葁�g�/8@`"O̠�6!�K�N�#�=.��4"OBl��䍵=t��W/�%q`x�'"O.Yp��B0K�������'����@1:x,Ro]�
C�i�	�'���!oZ4¥�^+4낭Iw�E�<�B^�?�&'� |�Mѡ��\�<���X�l�M�r�ޚ~������O�<����w9�ըAg�"�w�PN�<Y&	�=�(�"���aT��%�FT�<Q�G��^�\Pd^�p�|�DÖM�<	cjN�F��0PՈD %���`�q�<q��.!.9��Օr�e ��C�<i��9p�MЅAQ�6���DD�~�<yD� v����@. ;t��Go�w�<A��B��M�K� ��5��,�o�<AkMR�` Q�vU|M�7�Wn�<)�^z��D|JA�`��<q6M��pD9�ܽV��(�+�{�<Y��4U2Ҁc��ɺ|�0Hq拆{�<��T��x�Ҥӷm��Xï�y�<�CI8l<����1
�|l8��w�<ٷ/��u.�kuc�*&2��!t�<y�gU]JH��S�[o�i9QF�w�<)���_����C��V�����q�<��u1�R��Ǽ
j@���[p�<�`,ݩ~�Ĉ���X�=K#FD�<IU����qBȞLO~�rc��K�<�m���`�H?+$,�J���p�<�'�z�^�rT)��O�����Gv�<��T�i�<v�w{Dr4��I�<���\g���s�@S�0��i�!�Jn�<� �̀3$��b�����X�����"OJȹJ_���qI��$|���U"OjP�P)�	~.���CP#�l�I�"O�a�4�P+Z-lu������u��"O|�⦀��lX�6L�$B�y�v"Oj��.�Q�R	3��ސKB�J�"Oء�á+9��|(�l�?H|��S"Om��ᓵX�* Q����C0�h��"O��*��΅�yj�ɯ��"�"O�Y�p�6&��*֩Ε}��a�"O @ӧ6��9SI+2���"O������(&�y�(�9Tm<|��"OdR��S
7H0`��$����""O<PsČj�� Z I R���{�"O�Yc  ��%��E�����q�"O��K���5&a�a�>�B)�"O�-�sȗ�\X���.� 
�Դ��"O4�7��C��
��\�i�>Q��"O��S!cP
*J�Ǣ�����"O���c8\���&˘�0�Yq"O(�5(�1g����C�U	^ԋ�"OY��R��L���T'?YRy�7"O��P�(������_Sm��"OPq
�\;K"*�OT�!U<�y"O�l��N8y!�t{�.Y�~\���"O��+�n8xN �@�ѸP��	�"O�lBr��)T� t��d����"O:<��)^@��c�O��H�"O���w��|�\�W�˹�"�+ "O�L�SL�`2`�M�T�2�c7"O���B��$ԁLP���b�"O� ř%T�������Y�"O2%�"�^q�\fㄉ���bd"Op�B��%v3|Q�t��4y�Q��'$���+6�HH#�8E�m9
�'E�$ʴ��=#�����G����'��Q�ą�?m��0�ۗ>�0���'(Ш�5G�N��,���ރ7��@�'N`�:!pH��U��|����'alp*%	s�)R�,:"I:�'��t��оa����#D�z��-C�'��ܺr��'[w�T�E����
�'��(�C�C�Te
�%�[6ke�	�'���cT'ԀI*�YR�nC�1?DX��'�|y�a�YO\��Q�_��^�z	�'�`Y:b-!3�<�P�+.b� 	�'%l8ل O<+=��{����*�LS	�'[j=�@�U��rph3�ŋ6�P	�'ބX*.�u���:v�I�'	T��� V+���b*Y�����'
f��Çe���JJ�`9
�'딤���4{=�I�%�[�<��q�'�~Q������mYj-$m0�'�Y���Y!!���k� Xqp�y�'I����H!�0�EO�=jg��j�'�(��� �)�X��o	.p0�'pѰ���R�\)�Tl }�Yq�{��.$�,������'/����Nɴ�������2qA�J�{���8l�E��[2� ��m܍O`dB�I2ވ�Y�7JR�x�D�/�B�IV2���Ъ߄]�.}�M�33�B䉤P�X�c���E�9���/�~B�I�jǸ�3Vy��CfI�#y`$C䉾,���ɋA[���h��cJC�)� NQ�.�n!9�B>^>���"O�J�C�5E�x�*�#X�p+09��"O��٣�Q�I� �͝R�TU!�"OС�4�7����A����"O&��kҀv�4�!r`]�!�$M�e"O�䢁
�"w�|�䆖' �J1zE"OL5#�HɊ4�L��SƄ��0��B"O"<aQ�U�rt��&�$t���;�"O�<���T�H�s�/Y���E��"O�Њ�/ݾ�b�@���ض"O��J�c�`Dɳ@�Ǆ�4Yy�"ON�8PmֵYD���"�g�=� "O�D�Dٛ#��89�C� ��(�"Ol�,���B#�81kZ�"O���G��g�~��`_":���Q�"O��Q��ft	��'үV9�0�"O�jJ�F����%g	�4���u"O^��"(͸0`�E���� C�"O,�x�aσ`py�떷C�VQ�E"O��e*�f��z���1Ѳ�&"O�i��/ÇD���� Q�>T*R"OHl�P �c!j ���z�r�"O ���.�
��Ɋc�nq~P�'"O�P5ʭH���K ��$Z�����"O�LH�*ڡn��ps⚑�h+"OJ��P�EbU
��]2��9�䞴�yBC� *2D�DF�j��A�X�y���dk!�Q�
f��@�[!�y�ϱB<�P@�Z�h� N�+�yRK�{@ ��K�&%0���y�p��E�>��+D)�/*��Ĳ�'�L�32d{��c���7�L,��'$��&D�/fY"�-d�B3���yr�R �P�
�g�6�M��n
�yB���_�5��B��,�@��3�y��3F���Dݑw��S5Iֽ�y��
i��|�!�@/��d�dĆ��yR��40iʵ��F��Q�`4�yrf	l"��(1�]>6mDɧ�y���/o�T1�,�3)OP8��Fş�y�h�i�p����
�h ��Ա�y��Yo"�yj���&)#�y�'ɕ3g��[��I7�tL3�M��yRd��b�:@R%�$�hq)��yBN�5 �(�*��2a�HYw.�'�ybEM�FD��xפ�T�4d#�d�)�y⯀�p$�6l�Gj�T��	�yR�ԍI%jT�!�؛vʀ#��Q�y����Z�C����D�zd!Fm��yb��n^4hW�ECW�L�FGJz�<���	�(Q���NL=Ei\%�KUB�<���9K�%H"߼fw0�X� H@�<I�˞�B�<��ID�3��<����Q�<	u��^m�X��_�OE�`SBj�<I�̏�4jj� �D9�N��1+o�<ɵ�ƨYh��R�8#/�Ð�i�<V�	D��3 � �@��<����g�<!�HQ�t�d$Y���LFh6d�<I�ꀴX�@(n�I�1X��+5b�c�<A�� �:e앪�ޭ	L����y�<)D&
0����?8?�)�B�_�<�!�A��)b4U6`qe��W�<)���%�F�Wڵ	v���B�p `B�!�����B]�B�)� t�P�@����x���̶*���W"O0��#�R� �*i��I��}2iJ�"O����c�0�T@C�\+R�t"O�X�©�5 K�]Q�a��O�V�B"OҀ+3 7s~`(
�-K~�Qp"O*����Y,l�ZG	�-"D��"O����Έ�A}���D-�::\�s�"O���+�h�b��lJ�q:�"O�ĸp+L#5�nN�\I�G&D�((����7��	)L�� ��kT&1D��{���&-y�,�'1j�,R`�;D�t�!G��zm��kA�k�̸Zh&D� �'"���պEn�04�XL;�$D��2�N$	Ut��Uc�� �>���!D�*�˘'+�=��D�412$�dG/D�:����&߱dt�H�Oe]�B�I�d?�ث�� �`Ț�bI�kZ�C�ɴ
���CB0��Y��WC�I O���"�
~��Qd�U-t�C�	�?�*�f�%mvt�s���-k�C�	3&w�Ĳ��7kEN�ɖF�u��C�	�w�6�k���* U.�"Q_�f�~C�q�%� �Ѷ�̣��ǅq��B䉘����@�0'��k� E�h�~C䉛S�bT�H����\PqH�k�4C�	6VrH�#��!Y�8{3�a2$C�	�Ox���F���z���m@�j� C�	9{��:g��D�� -��C�I�d��B�g�#�nY�`�Y�(-C�I�i=Jᱣ�&9PQi�JǗ���J�B���I�9+��)�)U~�M�QI�Z�!���A��>K��8�g��\t�<Ĝs6��4��<�@j)���G&��~�R,K�*�Z���PC�'�u�5�V A 隵�M�s�T}*�dK��hB�I�#E��3g��BĦȡC��Z�D#=�!�ұb����Rb"�1�J������r=�f�����p�"O�q*@)X�|0bI��̞�tQ�Z�"�B���+��:L�XKm��"~��H���t�ڐYa2��L�K�B�IR 
x���ŕn��2��ƇI�E#�4qֹ�vɝ�&t��4!��|F|r�^3���I���8���U�5�0>@DԈ"�s���k��)�iX6RZ��i'�Q�O��%���˺���Ą#���H�&!�¨����41B�O���"N�)Y��ە����S5�~�@�G'f,����<<�@���Wj�<���hL��jа(�T�񏀏a�`��ɔ
,	��Z�Y�D��;Or���<L�\��cC:�&�p�"O����[��m�%��C`Y�f�ަa3d#H�:�!v \KZL�݈�O�,�nV�sy��@lP�ތ���'��h�ȋ19�[ �7}��SW�Y�ZKJȊ�^�8�0|ѳ�A5e�����A��(��3�y8�w�ON����$Vt:S���4�z���i�,t2,KL�-��t9!��5A�a�]j��gg/�^Q`!8Q��d�	K�<�&�l:�'Br�d+F#$�R�#XD����\�F]!��C�4D&����)B��U��#0><5n�_��"A�I�*^�y �wݥ#��$ޙoh.y[�È�Z��U)�'ʈ}��{�aL�2����3#ι/�
h���;L��3t&ȉfe�(�t�P�v[����Ԙh��,�d\���Ij�U�3�i��Q��&*̴�{�n��� �~b�������"�=���B�`�d�<�&,����g˽fd��&Ϳ�~r�|��4!g���MG��'P���R,K�[�12@��$N��b�'�`�+���Dx^�k&AM6 9@��<yE��$I�6��5��bf�	BMJ��P.(�2`��끑�p?yd섹&��)Bt2L0Ѕ ]3%|� `�q"C�	�$W���댎U�|�+L[F#>���Z�B�~�ӵ�J`�'���J���nء��@�<E����S�? |�KqŒ�{��RTX$%����OD���ć�z@"�O�>(F��j���¨ƙY7H03�<D���5�����F�8P�	��j<�
1 8���ɚ*�Ɖ	�1�X��2�dU��,բ\C'�P'1�j�Y�Z���o[��i珉7 ����& &�؄ȓ>=�5�vː�zd���ܛIDzԄ�a�F������s��סkR(�7"O�������K#�D��k�� U�XY�"O���m��IҨ��S(�+aq��"O��;��ؗ�>�X�OhL"�3t"O�	S1˖6�R,3��e��T��"O�����8�hP�R�H�+}���"O�!�	=Q�r��#^,rP$`#"O�����W.Lx��3R0%X�<b�"O�U�v(��I���O'u@�	u"OB=�q ��tస�Q�<e��p�"O��%+�x8��b�����"O��"�d4\A��㥇�
���"O�l4m�#K#L��B�;u���C"O��A��O�6Y�u�K�G�T{f"O��A� ۝$W�����E�s�b��c"Oz�0D�\�zw<!щ'˄�I�"O8��%E˓Lv� ��#M2��y"ONAS��ˤ�.@��ͷ&��@F"Oؑ���C2X|�2Ph#mo��:F"O���G�N�B�3���b��k""O���ԍS�Lb���ŃXI<yhT"O�(#/��$���Q �A�C
�"O�dB�-@$X��తҹw�n�b�"O*Z5%]&�hRb���庁"O�(p&
ǟ/}"�zt��j8V=��"O���%U��2�FH� H��a�"OFp*#J�N��$EV3r�j!t"O�+@�L.1��)�C�ɍ�~j�"O(� �[�6 �:�QZ�t��"O.D���R7&�TH�%�@QnT�"O mCL�M�q�A�9J���1"O�]��O��Næ�
�C����81"O�<�2��x��;v��2r����"Oȝ�1kӹ}�����l��l<,�"O�@pe��5�<��0,���F��"O� e��[�6��,�T�R1ۤ"O�`��֓窠;�$��3�ZXC"O4 ���I-S���kQ;9p�0�"O2���B�J�qj�a4tq��"O��;#d�
��6�۾\�ˇ�y�C�Ty��p&iIJ�~���L#�yCG��ЉV!7G�j���"�y��R$Y�h� 5��N��HX��6�y� ����i�L��H�L��y2e�?~ �Wg֬i��;�eû�y�M@ p~H��B͒�Qbf� �y�
�r!2��/��˵��y2�ȶ(��Y�p,��	�r���H��yb��.�:���)�(o�����yr�ܠ"�"���H�0�
�*����y�%�d��ܠ�Q���q�V����y2�J1>Z����,a�)y�"	��y���!wZ���C�
 �
��Ѹ�yo�+P�)���.�h
$��θ'M���7X+ށ�EHQ85���YM>aT��k�$倐��i�re�Is�<�ǃ�e^A��I�H�֕
U Rl�<yq�˭4D��(�2ct
*�'�d�<� ��ɴl�(����M�n�T`��"Or=��i'���(��N>�&Xw"ON��F�јFH23�iGJ�@�"O2<X1�2� 4��o�"�К�"O�q����p��H6�?8<L�W"O@ݨf������	�):��!"OĹ#rJN-�� �( �mj"ժ�"Op�0��ɈS����R��+/���"O��E`Z�C�6���-@�-����"Ov��&ƓXϢ��LZ8�T(qt"OU	��A'����A���Z�PQ"O���
Q�a}̸s�޹ �j- �"OL�h�'�L-D����=�c"O��;�ʠk���q��X��l��"O��kf8ܜ�R���!K�i�"O���Se]�(�(r$��:1f|���"O*�2�I N���$��
d�<"O���'�I j��4BXtb�x"�"O��x�(Or�dA���	V�>�r"O���`�
6f(��kY�o�e�s"O��ؗ'Y[�y 7M��p���"O��s�M>(ޡ UM�f(%��"O�)S��.�f���	dZ$��r"O�q�� �(��8����f��"O6�� ��:���3*��6p�#"O��U�]Z�E�ǆF�6� cU"O^53vd��_�lt��K؀7{@1X"O�u�V�)\�r���Rv�&"OfC��݆`�<AI� 9se(�sd"O�l	B+	&��|y@�ϗ2a0i[p"O��ч�֜W��y[qM� V<\��"O���7K*�fe��m܃CN���C"O恀���<76=)�N�g�n��@"O����/Uns����K��.�� ��"O.���'�{B�dA�%8ٌ� �"ON��g�k|pp��WC�"�0�"OF��d��1$� $�T�dHa"O��TgH�aQ�mᕋ�4n5�u"O$��nZd	�y�d쎵e��d�"OPx:�Ǐ@����勞�$�,��"O����n�n��`��r\�U"OX�aԠ��T���W�Y07���E"O��Ѵa�2R����"h�Chd0y�"O�;TT�J��dqHE5fTJ��"O�����e��iR���AE����"O���p��C�T( ���w*()�"O��Q�c[8U��B���78h�Ic"OB5ٖOA���Ro�?a����d"O���Ȁ�U�bTJ��E9,�Z)�"O�j��T'�$ۤ'�4f^�H�"O�yrqo�
S7�Q�#u��a�"O��0��	n�̄H���7HI��"Oi��JEpr"�jUBEz2@��"O�����R����E���˧�[�<yS��6h�r�͸	�#b[�<)""	�[�Dt��m�+��a�$.A�<��m¡� I�P��-�:䫰D�T�<�pjͶ c$�S �ީc�<i��R�<ACnĝ1�]���P?����`K�<��R�E(� hq�E?6,�Q��L�<��
V�u��0��<Kuf$�U�2T���� =6��h��)	��؉�6D��9 �	�:M{b(0V�H��g6D��s�=�ݛ�E�`�`�!'D�� zE�#�R.sՐ�I��N�"��"O�{b� )� 1`��g�h�u"O*,cf���o~l�3�/x� i;�"O�h0V�n͈��nC���Dj"O(E�����0��G�ۘ\ZeH�"OD�Ц�@=E�r��jS���my`"OhDB��Ո,RB�xb�C8f�P��"O�5K�.�\b�)��nԠ*�` 0"On20��A4�#N
�X���Q�"OB�3�\�q���ʤ暟6�H�*%"O��8��ǋ7�y�˒-mu�5�"O&L*WZ:4�q��ꔠG��y�"O:��B�q�Ġ`�L�(T3�I�1"O�(��V�2�q*wl�p��	�t"O��jb�)�Q�b���9���"D�h��E�iV8y��҉>+&sc$D� 0��\2�)C���{S�YW+%D����
y!r�I��Ȩ6��R@�6D��	��ֆgm 9"��4�a���/D�t�,&x��Cl���XJ�B�I5
���Q�C��C�����f�9V�C�	=�L��b�G�Xx件c0s�$B�	�}"5p�QDbD�P#�[g�B�Ɂ
�*�;��30�-q���8�B��?ZA��16��=|-H'�*alzB�I�,�:8�m�A\q�R�ߵp^�C��S��U�w%X����!&^/��C�	2m����'@�$��ց�+�^B�	�p���i4B��$Š�@Э@g~B�	VR`H�	��8�ɉ*�vB�I	-Q�x��&W>b�&�2rcܜ�,C�I9]�dU��5D�N!���T�:C�$1f������SF	1C�Q�*C䉁R��ٶ�� ���W�:R��B�ɔav�bv�S�J�
]{u
ΡZ��B�ɴh�PБ`�e�@T-� j�� "O 3�o� Cn�&UH(ؤ"Oh�H��wB5j��ڣ6�3!"OH��_�/!�ɛ�( �.)��"ON�+u���$�<1!�Ύ T$�4#"O�Q�1ěՀ�j��W���!"O؈CKL�uB>�#%�e40�!"O�U3�-��+u` �nW-����u"Ot5y7)�4DM�I��P���	@"OfH��MJx�y84��:~):�ȃ"Oh�V����O-I�|U���LY�<Ib � _�`��1bŴ���Q�<��
a�J	ZP� If���OXx�<irI_ L_R Cg
�_�0���Dr�<�qjԁ�$�r2d�Bd�@1El�c�<`n�]�����Z�i�r���,�u�<i  ͒}'��ҧKN�I��C���m�<��Ԩ�����˓6eB��t��C��D{�*S+H�0��+ԒΕE���\�C䉴F��H 7�L.������(l��C�ɣ�����[�gܚ�kQ$��V�C�ɅV�1+��{C4��F �H1�B��5l�f��Q
M"wL�)�0�_{��B���ؽX%��o~tIdE��]�B��
M3Da������2�?3�JB�	���	&�3f-���Z�B�ɢt`�Y;�h�-)D�+�H$;GC�I"s%�����(��(�0|��C�ɖӒ��tְ)RX|���ǝv�C�)� `���
#�P�f���T�^)�p"O�}�aؾj�0I��t�0��"O���ț8Z_� $Q�W>�q "O0(��J e��䣠і�Ⱐ�"O��V�A^�re��#�)4"O
��'��]P�y�m�:�2���"O�4띞}���(G�o��b"O��ٓ,ܘ-jv5�A�(k�T�"O���N2���KN
1R�Ԉc"O�� H�b�V�*��g;�9"1"O������	E�t��l��b	cG"O���W������K*9��a "Oę���Gqk��Ӗ`ɛM+���"O����!�%T�� ��#
`]��"O��P�F@`~�0��֞U�p"O\�!TdVP�j�N�!B� �r"OF\� �U.)_ʵ�@���4�*lY0"O��37�μ%Fh4���O�:[�\�ȓTԶ�0A�X�M`2ՊS˄k3N���L��@�aU@�|��ۦY5� ��y8B(�q�Y�\񓠅�C9>�ȓzP���̖&X�z��	[pa��aH�5�Ĝr2�Y��<>�8�ȓb"2ʰ��i,R\	��ϓ|?��ȓ (����,Obth��̩��W�S�Y�ka�`ơ�5����ȓK�|�2��;|L�K�m0b<0��I�dĢr�2S�$��T3%|t���H��Y��Ό�s
��cC[)Y��������I�l���E� u�Nɇȓ�|H��b�'�ͩӪ�|u��ȓn�\��U��a:�	)*@}�XͅȓH�^-���	2��x:�A�*���ȓ\6��� #\6��LJU%Ӥ���7��"�B�"z��·O@,-ɸԆ�T�؀0Љ���E��愩c��M��xiҜ���9Md����Q�|��ȓ`ݘ`����QI<�r* �{3�M��o��9����u?zH*b��(u�ȓK���y���o�6�y�`ڶ_a�ȓ��ѩ���0�T��2���4u2�ȓ#}����K��<��Q���$i���h�h��\�6�"��b�P�7J9��s�}�v%����x�#�;�P��S\�c���<��Y U�G�H��5�ȓ��i�R��,`������lV
!�ȓɨ�X�@B+B�`��Ӂɵ$Ь0�ȓv@͡"iV�qy�w鋧[t�ȓ#�<1ƥۊ���bO̟ L �ȓiu�Q�ej�ΘC�_$V�zY��U�,j�O9n�@󤢕���A��nFX1��f�<X�9�@�MD�����TBÁE�v��i�'��<,�ȓ.�(8�@�4M�hfŇw�
��ȓUȕ�2&��P8���Ϯ�"O�Q�w����)x$��S�U6"O��&Ó�_v�����_��ِ"OX�:�m >��Sr��/��=�#"O,������f�q�oߠ�摳1"Oj�cr��e*"���HC(�%x�"O ��H�?|�y�'��]i"O���N� r(D���,�n �"O@�Z���bմi���G��0���"O|LKF)��f�����a� @'"O� ��33�Н��VC��y[&y�"O��s'MN,1Ρ���:A����"O`�`\�l�J��(%��z�"OL�����:},=)�F"7�@�"Ȏ��n�]����%�˷h���"O�pbv_&�����	���T��"O:X�S��(g�H�qv�T<��@"O*UY�ᕊG�ĉ�&�[�f�N���"O4�C��|�H�
�*a�6�&"O�����?G��yb�D&�x$�3"O��R�2��y�VjS$?Ȥ�ۣ"O�����X���prϟ�A�\��$"O���lJ�<,,i5�âg���[d"O�030G]un\y�.g�h�9�"O���r�Ȯm�`H�!K)x�B�0 "Op=��˦|�̈ˁ���{��m�F"O���	O�Yr6��8kr�q�"O�]�T�20�m�ׇ�2[4N�*�"O���p
�%T�dI�#!�"�Ah1"O�,
VIπ,����`�.#�l�"O-��%ՉO�X]J���ڡ�s"O��QVG4:��X���~T��`"O��[���.s�1z��ؾ��"O�Q��mA|�:p.��tъ��"O.`�ƄƋ�qS�Ӡk.��c�"O���@��\�P4�_�3&� �&"O��i��+��<�di-L]��"OH�;�(�=NM�Ǘ % [�"Ob�ر"�7��a���O	.�9�"Ov�!"�E'y2
�z愔�a�S�"O�(pI���ٲ"��%hH6x'"O&Q&kN�TF��1���af���"Oh)Rs'�Q^���E���HL`�"Ol1:P@��8���`��KJ�C"O�hS��^�M�����t��0�"O,!�T4Dp]Y&+H+uքe0�"O"�k��#�d����[0 ��8�"O�-��cF,$*Y�R����F"O�}a��
=8*D�.��;��0"O��{���
-.�2q��\��"Ov�B�Õ�FV��'E�*1�����"Ol�B������%�6	i�@�"O�	!�N�3;�0`��$�_���"Oȱ�.��1(�Qi��04"O04����J̽��N,Xò=*C"O±��M��
�X���4����""O��ړ͞7Kd��O�$�����"O�y�SOW*t�xE"0�V�� 5��"O*�'�S���m^�p��c�m���y�P�w��#��n�&�0��6�y�C\��̐a7b8R��b��˝�yR���x�i`�;O�n��rC�'�y� N7$&Iy��X�@����VJ���y��E�\���Ɯ*���1�]��yBҗ��T�t�į �i�(��PyRBO�]Di5fQ�z��<Z�\@�<iVE�`9�E9���5D׀1
R�z�<�c~��1�kל'M$l3��u�<��%]&�	�����KQJ9D�TQ��3��  �Ǘb�a��.8D�̈%JI��MbV ��G'ځ�6
5D��2
\=5�������J*��:C(/D�Q��]�`��f�3Z,^�$3D�\Y��)U~Q�]�&� �3%�<D�� �M�������b	�i�(�q "Ot)
5�h%H�!�8p��ct"Oi���(Jv	Sᗥ.�,���"O��0L��N�s0 ^�i.X���"O���'fB:fK$@��(׃#1B"O �8c!\hH��Q��%Ib��"O�����L,�}I�ѐ{�&�H�"OD����O�����O�x�Re8"O��y�GP�`wJ݉�̴g��l�"O�Ũ��.ql�G�~�K���y�g �1����e�%��aH>�yZ�d��D�2<@�3B*���NU:�'8z	�U-ձ	SL(
B&��M�y8�'K�*��E./�u(4-�(K/J@�'
�3��!#F�����I�����'�| P�����#�1���*�'�@��q&�7	�8�`ۀw�@q�'m5��G������E]�tJ@�
�'��Y�!�6L��R�#�7=h4�`	�'� X�@ǦJ��\���%R^8��'+�0����#ɚ���
ʈEI�'xj�;P���fQ��@�K.S�'�h��F+I�l�H,�t@^�_��d��'�f��A&\�9l���a��U��y��'�,���DK,VBt�G�y��e��'�<P`

��6�բR�.�$"O��]���� ��]�JΦlk�"O q��͓P߄��Ӧ\^���"O[��R�=�F<suC��Q���"O考V�ۣA�1؅"R�5���B�"O"�̃�7nh�����c�����"O�u�␄\��i�
J5���r"O
xǉ�b#H��'�Qr"Z�{�"O�Q��26K�?DjnE�`o$�y�jL�<hv����$7\T� �)�y��F�aİX6�˾!s�<�7@�y��G�PǨ�X��V�����֬���y"�P�n9$%�M�~X:�����ybh
}�=��e�g��\i�,�*�y��B���2���s<�U�v���y�>dM��(Ze��Lȳmۖ�y�a�74ʌ��
�t�*�$�yΈkkn��3`lB��2�Ȕ�y��>J���r(\��`08M/�y��K�{h�
����7�@� ���yR�#��Q�C?)�@My��=�y"�:$K�0���ɷD��V���ȓF��E�0�R�Q����gkJ�[��\�������O�3+R�Q�Ң>���ȓ,ϒ���˱f�-�����(��8�ȓ~�����/n<|a��22�Ʉ�i���l	�K����D�e�1��0��c\�&��1@�ܟ\X���P9Ʃ۾mnIi�Q6�x�ȓ)	d�P��95@4�i4F�+��Y��,:�-Q�c�@�^�'�S��ȓ7-��kv��$[j��n�=u����ȓ)R�,�%O�xdc��X�]<���ȓ-�^!;u.�۬���
R�@!��/&�*
�|a�A1$��4pT��ȓ/�B�b%�T�4}\$���h�⽇�B��AаOI3/i����%�� ���r�Q�j�3KY��x���
a�2 ���4-��8:4�X ���af2D�� ����ņs�"Aٶ. �m�� "O��ۡAׯ]�`���"�=!e"O�-��@�?E�\ �M�^Ҝ��"O���פ��:X�uF8I�0yi3"O����0&AbWg�6�p�R�"O� ��c��j�}���a��1�"OX�RC��PH��W�B	�R"OJ�ʐ���k<� ���
 ,,S�"O�I2��%s��R'��@��y�w"O
��Tk�y�r"�۾I�؜�"O��W�	:r�*�B�V��&"OK�N2mc�� ���
D��yr�@�ɨw��$M�k	� �y��72l�CiM�mqX�9����y���f�T�J����V��k��y̘�D�����$<�ʭC���y�J�jR()�����@�UJ�4�y��G� �#�$���	�y��í$�.���4|�H�$���y�䓨J��5�nɥ&>�! �I���y�FS
!�*q����!��mi��©�y��L&
��Q�I"i<H�H��yRO��P�4�Ҏ;Q��ݳ7��$�y�!��E>D���9I������ �y�R�"!�TIR%+IlJT!Ǯ�0�y�F��t����� WkD�2v���yr�Q.��IS�H<fDJ��.�y��!%Cr�؅u�r�ig���y2�X��L�7H� �s�#�'�yR�P�׀[~ChRPgJ��y�\Yc������{:ޔ�gˀ��yrP8X����EXrI(��wA�	�yBc_�����رq�r��Ǭ�/�y	G uz��J��T�J�C7(P�y�/P���0����H��j����y\E��2�/�:F��x�!����y�O?�TY�ؖ;�E��mR��y�B��\;xQ����Gm65�`� �y���jB��hs팙VAtk�A[�y����|�XR�c��˗d��y���E,�X���D5U��Rw�N��y2G_(![d\���#JL�x�����y�A>�F���.�J���0�yR�ЏD���	Rm�G0�qw�'�yR�O� ��m�B��B�8?.��
�'�a���fIe�G���J���	�'����aa�w �iQ��I�
�I�'������T�����{S.��'z� 6H��@��l����F�,���'�>��Y5<b�ȗ΁,x�TQ�;D���v	ۊK�h0Y�K4[���B	:D��Q�A-c�����im�ˇB7D����Ʊt���雺NH�1AI"D�p�`B"1Φ�CD�Z^pzV�!D�����D聢��
,`�S	!D��HA� �)Y�Ԑ���
<ҡM)D��r�D����ئ�+7,qZbh%D��i���9��R� $�$����'D�dY�`�W�S���:w[��J�"'D�$I˔��U��	.���8D���PB�^bR�"dZ� v���p5D��S!��p���v&ؒY����62D�:���>\"���dU#U<�D��1D�0�T�PɴlN�a|���4�<��B�)� v�gI�
\JQ�����y�6Y�S"Opib��\cv`:tΕb��;"O]{��М�M�cH�|�u"O�!	�	�k�4��"`�|��8 �"O�|bg��v��5�EC'9���R��IԟDQ�攊���'��Y?�*��Q�R\(�&�ܝ$^\0S�OS�e�TH��?A��]��=K`��m|��	%!R &0����~>�b��'h���F�~�<�І#.�=��I"l)���a�$~��bB N$� ,��%Z�h3�,+e�}^�� �k2B�T��O@oڳ�M+����	��8��� �h�?+"d��Z�eX���IF�S��?I�W�j�@u��g�BݛtCP��,�	�M;׸i�����9��ɪ��W?l�H\)鐓�~�'Y�e�����'F�Z>E� ʟ�I�����l˽,l�%.�2l�j���䝏s�nX2�Ƃ�d��a�%�8 )yT��?ŖO�d��|�!(ó�v=�o�� < Կis��1�f���+1F=�0�W�]Ss�U�Q�z�����#Ԫ?~X~a����.Kb�	1�i�Xu��՛�jrӂ�d?��qfN�?� �0�)�?���be㨟��	AX�@�e�T"!Y(�s'!
.mH���/3ʓ ܛ��xӀ�O���vݽj�ϛ�� D��A&Mx��ϫ�?1��l�VU�����	�t�I�0r��J7MǶ:��9��4+�����\���`Q5|�m`��D�+n6���G��?�) �/F
��iF)C,[|Az��:�0��W恅f�6@�U�]&%ܳ�~�Vڶ
��=i��<I���h��M��
���IFIS�4}除
���z������ʟ�'�V����h�V�R�f�%6x0;�'/0pD�K `k�"*��������[�4����������lpT�.̈́�1��6
����i֝K����O6�d�O�%SN�O�D�O����T �Fu#+�/`j�����>��0��֙,�HP�����ZKH�����ЕQ؎�(D�T�o$4��ѫ��a]���'|�pfd�")�8yh��j�@a`C�Z߸'�4�1��M� ��Is0qC�0žu�s��bjO��$Ʌ�����|��m�^ۖmc�l�K8(��I	I�<�pMJ���p�#�Ӂe \P!��G?�b�iS&7��<�3�$~�v�'T�Y?��疊���&I�g��X��d��RO������?q��p�p�L,��<�%��e��KT�l>��DG2V6}(���p��)>�a�X�3�%ݰ=����7��	�U����#peP<+��X�2�K�BqA5��35$�a2�{���?)��Q�O,�vL<$��df�P/:�2�d����5�)*�}Z0�q���o{|�Q���83����H����}�N6T�%�j�����3\$���fƮ~���Ÿ}d��n�ڟ���L���P:Ig��'i�fe�n�8�&I�=V�`k���xV��GěW�&h���6\r5�$BĊ��4[>q�����L=E�D�ٚe�&��ExR��9s�L��P�W;�\"G!��*T�3�i�� }��{�ODU���)��E�`�@=iՎ�ʦ�`���O��lZ%�M[������F� }��p��	$]Ό�aBK��~��'R�'\��P�~���*+�]3��$v�
=(�,F�'1���f�B�O��'0�ChL,
��ՙ����×|��'��ј� ��   z   Ĵ���	��Z�JwIJ(ʜ�cd�<��k٥���qe�H�4��S66<���]�f��->(p��o�!9�0��o��gZ7mæ�‫��y���<�a�	M���$a6v|�,/ff��K��J�➨�U�xr ��4�f`�`�i}����!p5�q"�
�8�|B�O&�!q䆨?vt�-O^]ڗg�]��(Oԅ
�IN�����$	�o�Y��Nш4鴰i`��9�<Op��mR�m����|�"��+?��!ywn1D`���)�5OqN�:�L��1 s�ނ"�~�2�O�l�'"��Agc�>�`�%d������@��6����A���&\dx�oИ��DP�X�D�8A]��3�\��Qn�{rt�r�Y.(]S!Ɯ=v��G"�I�D�$hf�X�H���.ڊb�d�BB	 �O�)����ն���	�g��P�g�"n�vI[�$�:?�:�b"<�Dg$�����8p�1�0)>�6���O����$���j����r.����JN� 劶�d��OF�y�Od�r��A3 Z12�� �e3�T�|k5�ɳoR�O�𙥪؂5�P'����Ѐ[�-�ODd�����?�m@Ȋ�B)��H�d��q�~��#<9�/.�$��O��`�������1�ߧa���Od�N<�c_���!�H@��hk5��-9��y7�O��Y��i�J�EG0�?A�CQ?ͧ�~rq���R�H�ؽXTh�u5��gJt�E�d#<��/}B`Q4)��1�s�!A�4 �΁;��d^�Ot�s���	�?e
M�'��,j�\ٻP��K!�d�? �  ��u�r!ʯUi\q�9/��$�O���Oa:���O��$�O^Acc�r��i�a_�T�ԕagJ�)p���Bgo�uZe*� C��s4m��C�Q��/�e¹+wa�:���
�� R^���݉k��#Ӥ���
��#%�9�MɅ� c�9���^�
 f�,�ȸP6�ɪH5���հ�M����$ӼR����]�|��fƇt���Y��ٽo5 E2f�`�'aayR�N�r>�c���f�T�T�ܪ4e����6Iܘ�lɟ!��r�`L��u��'�"�S���;bR��U΅�f���	0%\u(����'�2�'BX�����O�MۦɅ�v�<$�!Bk���@/#�T�s�F9E1|@���@�h�<i��J63��i�r�1sT���    �  �  �  .  q#  �)  a.   Ĵ���	����ZviL����0R�PΓ���q�']�ڕK߼=���똁{h���'ꌝI4�\�s(� �WO܀nE8�`7��B~�Y��C�H��]�|���I%Ř�aܜ`�Mيzmha����^,64����%�щ�6�pA�L�+ߒ��CGR�0����ND��3��#@LE�P��"�FЁ��K�7�L��B�B�[SdI�����Q�	Z�=�4S�B�:a0���؟P�I����ɒ�u��'Btb�È7ts��c)۷l�����u�z�$N�������l��`ɑo�!� �5���Yi(})�j-�L!n��Ǵ�Z�,�I��(OP�	F���B��1P���!�D�i��HY8���'|��gy"�'d�$̆�2���όeWx��䯏�~m�O��=���?����t9�𰴩��2=�h�g�Am�f��>!+O~��O��Q���R�W8�����k�f�j�F٘���hT����<�	������u��'B�'a�ӕ萌c��)�+�>�&�#�	C�4Z j&&,�O����8ҺTQ���d�z�;��%�8Cai�(�UL+<O�4C��'.]�(�;e������vj�<���h�@-�>���ܨO�q���G�J�419B� �#�($#��x��'�V�4Gy�(����G@�;c��0�����M���cl���'�剠'��k�4�?y���?�1zP@)��GдC֨)���(/o� l ��$��������'�x��	b�S"�.:Hh����	Ğ��e�c�'Ȗ��)��`F\x�Z� �2�K�[:uў�����O�F�T�^-�D�q�^7V�
��t����y�JVx�V+Y�S� y��Tΰ>�����a�V2�x��PHQ�"������>Q�ꌉF��f�'"R\>�R��������[�|�"RgT��LS� �X�	�4S4<+�阧��D.0����)��x����&y�+��O?�+g�[�pd�8'A�S�(�K�Nٟ�*��O '�"~�%��7.�,H6�^f�>�pG�L��y"��Fn��z��7W`T`�HON]D�����p���j��gݘ�X��8[r�6�O��d$R۬��`k�O����O�Ďٺ���CĀ�&����q䊣5��O[yjˊ�p>)��@N����a��!2�w%Ny�&��p>���Y�6�r�B�[\m���sy�C
�?1��'���p�:4���9��K�V4�yR.μ.�2��C�9l^�a���Mc �i>�%�$#���<.���Cs���d�T�h#����b%�����I̟p�	��uW�'�5���:D�'�����I��"өFԛ�m:�O�h���O����b	r����d�
�Ry���'�Zy�� *♊$M:Ch:�k�&�L���Z�"Oz	Hb��4[�$U��Q2"O$8���([�0dc��$���Y�$�ٴ��
���K0K&�U7��P"�p��i"j��/�b�����S�Jh�Y�'�
����"{a4,�F�/U��E�	�'U	��@�m"�!6���Y���r�'#�0Vd[���]�L�$Yq�<H�'�\y`A�����b%.�,S����ȓ<)"�q�H�e�&�GJߪ,6du��kg�A`���<�fI�əM��ԇ�DJ���p*D3Y�	��k.H>؅ȓ%�H�F�J>l�R I"�G�4@�}�ʓ:r8��3���1e��h����D�bB�ɺm*����"��mdA#��X�*B�	�G�h�a2�H�l�`����1Q�B�	9|�,�P��-��!h�@ܰ6>�B�I4)$�(�2@��5S�A��_�:�C��=)��y��-�%n�P��#{��C�I�E[1��B+��(�7Y lB�ɼ)�8t��6e�XD�"%Ƶ׀C�I�^��1r�(y�l���)S"B�ɀ`�%��@$��駏��B�	�p�20pG"�!9x1�ć�o�B�I$8A�KtB��A�*�CvA�C-B�I�OJ���w�E2�: �aI-	B�	B��P�d#�:�p)qDA<K$B�ɓ*���"��9�r e�ϗ"[@B䉼D�,@�f�F�Dt�F��KB�)� \Pɴ��p���4 � ���a"O<-z�%W�f?4�0�Iѐ�8Ӗ"O -�OD�r�*ڜ$�t�B"O�Ay�b:W����c�j����"O>�'�#��ǣM������"OH�H��ϲ!z@u��B�R0�6"O�8�%�߻|��;��=����4"O�4:eo��~)\���8d����"O��q�a&M�"]� H4^�Z�*"O�-�5@�?}��U���aT����"OlD�"B�[� $c?�x��G"O޵a4��2e��As��k��Hr�"O~L�#Ε�]�') C�|�
e"OL�K�'��x<9�O�!7p�$"OrR�� ��5+�n��7(�kE"O&*6�_r���3��A;k!��2F"O�0�뚥x����Fئ-�L���"O�p��\��
��E�2���Z�"O�����<7p�ah7Ý��tЛ�"O�|9�N]���%��#Nl�qJ "Or1R�M0u�8�ʕ��b�:��a"Oڕ�M��噷&�p�r�8G"OB�!D��,���҅D�,q�"O�M�ʞ�kSJl�3(�m@<��"OF Y&��g�P��bm1Wl�0�"OD��0o�2vEDE�!��y�j"O�P
t��&\�Z��֮�3w�H�F"Oɠ K.	)��)s�֘j�<uRr"O!���op�����Y��훤"OB0��ֆz���J��}��"O�eP��L�b��P��rP����"O\���i�>$zU�0f�1]$��f"O�i�Q�)lp�1��N��[/�eK�"O��#v��O�<��&� Z{yQ"O�� )�1��}��d�V-rs"O,\���է1^���dǝ�Ҙ�"O�y���ȞK��4ȋYא��"O���oۢ4�0�Q�/��6�M�!"O�A�%��%��d�5�9%���ғ"O���$XC��Y�Ŭ� n�"O�Ԣ�LPl\�x�$#в R�i�"O� ���"�h��r!�0��If"O�L�� ҥkf��#�٫D��:�"O�%!�$�>8;�Ё�Ɗ�gxa�"Ot@i�a؇2�b쐠��P�.a
4"O&y���86eL�� M��Q1"OZIq�C6���1�`k<�Z�"OV��sa�1 i�XS���-i:���"O��c���/Xk:�q�nF�+��"O�E!f�<i|��"vM�e24i�"O
�KN��B��J��8H�"OH�������#�_ 9�dI�"Ot9�������B�ׇ]Z��E"O���H_�X�E�@�S�W�DXa"O��B��]�$- )r����^�<ໆ"O$�x�D/m<�AfB��k���"Oi �8F
�"�O�o�2��`"O�iP3���P�c���H=���"O���W���7��E#bg�
Nt���"O:�Bg���.:
��a�ڢ(RL�r"Ox�i5�-�t� ��������"O�90�EX#ܮ$HU����i"O$q5��&�V�� �Y�	��a
7"O(��HI�8B�倗�0s�� �"O� nU�r�O���!��������"O�hF�[�|� �B1�T�w��[�"O��0E�]�| APLQ�~��"O\9�v.��*��	��D���S"OԽ�S�؟\���
X�@����"O���� �f+��_� �ȝ0"O*]�ŤDÞ�:"����as"O*!�CPpg�)��
RL��"�"O�x�f��aj�=b5�Z/5+�e�"OLذB��	̐4�S�G�V�:r"O���4�@��e�7�(K�"O� {@�_�7�P�ڇ�מ5�͛T�I�9jTG��
�>|¬A��)޺+�z�K�5�yr�Wp��%A��W^�R�g�"^� yso�q���H��I�]Rґ�`A;%�ݒ5M�!��B�	��.0Z�Ł y���P���rN��85���	��!�A��D���Au��S@�Ƭa��wJ1<O��QD�֌!d��sBAԟ���w��	ښ6*8����2D��B5Ä�,ѦLaE���i��I��>�7kS��Fѝ(f���-*�'cސ)I�o�  ������>�~��bc�
��L2e�1b�n}�!2Q�@��U�(c�FM�ǥߡ����^�¤��"�&-�x[�͔L�&��/��tP \���xP��J�0!��H�A����姘'5��EC�1LOx���ʛ+A�8q�
œ:� �Cd�'^\�����������aC��U4������ ��Ё���y�4%� (0��9i8�d��b���d 	3Rp�˂��&D_ࡒ�� �C��?��N޶� ���d-��F9D�����AO��1d]�C2��qk�.1��ɰ[Ûv�S&7�n�$?�IM>�U�ĩO�py��9&���tMLD��D�Q�ԉ_zy#�d	=:-�L�6�#ވ��Q��˖ѡ���$,S<�3ϓ,����X$@�9�#��X�F㏻"�\����LNbx�s � A0JM��c͹f
� +��-��u���$4��w�RD6&-�q/�.�j8�≼<���֝T4�����2��\��	���?���P�b���{c�Bq�4d�� D�`�rN���E�P�p��H	0e;����"�QȦr����Oy�Oxi	�Bڠ), �c%Fʫw���SOxh�j�2|s&��i�! ]����^��)�3o��p(�!�azʛ)[KRd8�@��K'�0<Y�*�8 |�����8�	�ń�PXFr҆ڳ[���X?I�
��ȓ��]cEdS?;5�Pɵ�m�6|�Oj�	�-j6}�Uf��6�|Z�`*_�a�U�B
kI<�q���X�<ّ�m�@8����,;�)�		�]��P�"�#��d��>�F��]BV��3u*�	d +�\���y:4�S��K/$#�-�(��in�&:
�t+��_�$$�{ � pŘ�Ä��-��PV����p=a�i��hԀ� �[����!OȲ4��m둯��}٠�Z##4D��D��8:�9Čն9-P���0�I+�b@1@�y�O�~8���<+��Se傽:JVE3�'�B�/EB.YKud�-cn@��"(�	4y�O��}��s3���a���N�T<�5ʅ���q���\t�@؃ &���0�ȓ�]�+�>T�xc��\�L�9�ȓL��L�a`�Iż�9B/��B�D�<1"��'��{qD#M���0��Nz�<qv+��;-b����(8r>����w�<�qgՔ"�r�@D/ �Eu��Q6��z�<�K�% X��#נU�5��L�A�x�<�F��
?K��b���~V��7cRn�<9�)x� ��%�<��𣊉S�<��cr!�x��U�P��n�<�aDY�`���t�U1hTL�W)�S�<a�S�\{����Цe�<AgQ�Om.�T�^r+zeH��KV�<	��ͣBxR�PC�^�ȉ`�Uv�<� ��%Q�x(b����*�~��"OL��a��4<rLYg�.X��\Y�"Ot�q�.�	{V�ZV
�A� �"Oؑr!"M�m��q�}fp�B"OF�zreI Zw���C4s��a`"O�D��$�t��q��T+z�X\�"O�(u ��\��I� L�)>���ё"O�8p��$�S�Z2����"O��S'oќB<������|6d��"Ol�qE$oH�c�dF�x`�v"Or�C3c��(2`kM2!��"O��q2ΐ�L&$TR���%^\�b"O�U���8$��a�6�ѭ Ɖ�g"O����&�maj�XT	_�W$!*q"O4�p�/0�&��d��.FQ(���"OL+��G�^�{ �%E�@u�"O^ȤG�z@���ކ76����4"OZ���\��	��	z�܁!c"O��!�/S#���@4����@���y�iЗ@�Y����$�<R7*���y��ؖJ�L��7�<&T�j�5�y"O*6@ˤ��>@�)a��F��y2��dÂ顠�!��#�.��y2�"3�H1W
-W-����ث�yBȆ�D��� yF Ԑ�'��y�H�s"�5�Y�h����� 
��y��X�F�y���J�JN����y�*���R���7�r�ꧤ,�yR���0t�Qط�;�P5ۂ¸�yR�¢4���d��ݫ��(�y����d�Zu"&�K�Tj�y�уK��y�
��t�����_Pf��i�B��yB�[�n�i[�+ߴ��@6mF��y2�Ա]/�ࠕ@8�[�	��y��+Һ�J'U�<{i�g���yB� h���Ѭ�8:S^u�-���y�.��QHpe�?�� ��y"h�t��I�<���;� ��y��\�������..=v<� ��y�b�-;��0���	3�&�J#,���y�'
yX�%�&v� k"fO�y¨��Qy����hQf�U�v�Ҥ�y"� n�x X5FF�5	L�yN����O�p��Ⱥr�Hb�ƣP��ՐֵiK��[�ˁ�ю����&?�H�#�'i��x�OU*-��R���8)Z��'~亃�X�Й*���.����'H�ͨS�߈-{�0� F��u��'���6�	_C���Ǭ����'�d�a��7�E ׈�'x��b	�'�,�����'WX>��&OG��hX�'��	��͞pCA#Em͝9L�!�'@���a �>-�*��k��8�b���'�� IB�B6n)*�� �_-�D�
�'��d�@&�gǇ0�����'
�И�J	T5j+H1/�}��'XB�i0ab��� ����6\��'���d��B��%�Щ]�	��H��'(n�+�,��-A:�*0�۾.-0X��'����M�;k�9IFFX/ � ��'�� ANR n`b�����l��'t�}�C.�hO"\�uN�I
rm��'�B�����y�v� F�@�|��'��e2��ZH���0�^;)��h��'���ZC0/���`��#�A���� ���tX�!$��ѐ��>�l�"Oؤ �L�5��t�� �c��+E"O:��H�8?.yP��U��4B�"O��1�YӦ}9d��9ז\	�"Ox�gj��3d�iE⅃�t=j"OL���I��l��� ���-�t(��"O��BGE� ���bZ>C�`@�"O��#C'J�>%�(Z�.�=V;Ĩ�f"Ov̒�^�ʰ�-o-���p"O��k��#���Y���J�(s�"O�x�b��P��y�Ɨ�H�p�""Ob�y���<S(��0#D9kM����"O�	����U�@Ђ2n �����F"Oz� w�^�P�D����X��-)6"O(�K���C�Q��L��(��`r"O�Y���}�zÓK�:h��Ѥ"O��e%L�f-�tH�a�\��t"OT��́u�0bh�6$�`���"O�X�EZ���`�蒉Bj�a�"O�BAL�9#���f��B�p@ f"O �$: *�"b'R��"OPݰ��$E|l�pvFZ�]�Z`�"O�-�FM�l۞0�gc�#���Q�"O��[6��,��\Z�g��sTt�u"O.ٹ7�ʮ0���gɘ�����"OEq0��)�𴪴IJH� �$"O�t�0n�(v�4��Ν�j؂��""O�s!��2k��࠮��!�2���"O�0d��#��R���x
�"O�d�PD10��.#�VU3"O��J!����Hݴ�9�"Ob��O	�m�J�h4lTj�*`�%"O�����X�P�\��fj�I�Xl�A"O4�b�,��q4��DcV�W��P�"O��9%�I����q��Q�:�,X�"O�!r�2V� �u*ڽ*y2S"O i����T��	��i��@'e�D"O�a��
Q�J��"�ɟ�x	�H�"O2h+����QS�'��
�,�!�"O.H�uiM�1����U*uU�C�"O��pw@��A�(�#F�F|E<pg"O�Z��	�?�L�����A�"O"�p#�M�3�T9�l�Nix�� "O ��o0\X�I%m��cU���""O0��R@<-�r���E�vIW"OJ<yf"�4�����ޘBX9a"O�T���U�wW,��*ώN9r��b"OУg�d���ٗ
���(2V"O��j�l�%�T�RT��B�u��"OȌ!WO�	k`M��F�#|���"O�Pk��=ÚM8uey+��i1"ObD;�HԊP�II�aN�<�q�3"OȽ�G.�$n���bQ�ܔo���(0"O��P�2�b�)�I�=B�8�"O��cLI'R����3S,�h�"O�p�@ǜ�`�2����3U<��S@"O����E�B�������_�X��"Ou"!/I�hD	��<��:�"OF�Q�'X�Q�>8[�NO���"O"M�p	�&d�A��
D�"O��s��2�I"N��1y,�p�"O���P`�h(�@�'�|n��RQ"O��`��$t0� u�<���"O:��&-��*������B��M�&"O� �D11�՝o]|�c�Z\�l%;6"O�̑���:h*py���-��qI�"O�y)�&��D/1�B���0YP"O,�D�η�Px!�� bf�\PG"O�U���:iH���N+8Uk�"Ol��F7S6��C	�$9��ݰ�"O�y�Rm�1zd����jR0BH��g"Oʐ�C���Z���I6H��xKd"O~\x�(�6e�$��iU�&%P�"O�yA�V2F/4YX��Q�;�}��"Oș�Ǎ�%���aP��+���2"O2,0T�Z_u�yj���z�A�"OtS��1n�F�@Doŉ
�"p"O�ĺ��ĨL�Q+����"O
�Z����m:��M��=w"O�|�a�H8fJ�!�@�o��2�"O<M��&){�\ds� :�N ��"O^�r��K�^0�� �fT
N�""ON਒��\��kW��86�Lp"O4I*D�� �h�?�,-�T"OBE	�ʏ'}��K��7J�Z���"O��k'A� o��ŀ�~=����yrK�t��P��Xh���!�yB�Rj�3�b	���Sw[h�ȓlZ�̀Q���U�tY���	j*0������"�\�o��e�p���sr �ȓ6 �p���Z�g����bҽ��D�ȓMETܛ.ZU΀hI釣=�pȅȓ�����ӃP���X���gF���oc��FָA�&a�L���T�ȓ�*� c*R�g�J�p���z�Fx�ȓv! �3m��j��ڜq"�E��w? )��p{�ɬVn<��"O�x"�1n������7B�����Oru���$r�v�S��SL��Qt��X����w�d�%$�0�c�^L�T[s _?1�!��U�6ؼ�ᦣ˿� A&e��h��Cy���遲#ސH�`��%k��� Z�!�$�5U�F��S��G5�p���i!��@� ��a�d?(2�91"CIR!�7#�6���R%���C�Y�!򄟽8�"�pao�1bn���-@	�!�E�؆C��̧_j���ؑ-8!�D�R�`�لcL�tx�A�Љ)�!�Dy6�YwiO/T4��"���9�!򤎀!����/f	 ]�W'�i�!��4F�r�ƞI�DM��0&!��Ie �聉�vEdM±� !��F!x�~$ !�B4�H�d��#+!�= +D�qlܐ{�b$�%��e!�V��+���-��e�$�R`!��E:Ɲ��吃)�ld6$ÎsJ!��0>���!�4��u愖�9�!�$� LN�G��'{Q��P֢B7��/h��ph�pMي�y2�B�Ḡ� P�њ�C��T��y2�J�KH�:'�̇S����N7�yrJW=���"�Y�A�B)�y��`,�� ,!e��f,^�yr� �e�2Ejϛ=2�0$XF*R9�y�L�;V�l���ơ5�N�	&	��y�Ε�Mi����W*��\���H�yrhǯW  �@�5��-b�N'�y�m��ِ��o1�H6�y
� f=�$e45&�k�"u�Zx�0"O>������ɲ�������"O�ˢG..Rag�"����G"OVI�!ꄔs��:��S�E�^�:�"O�i(BL�FPNQP�E��6务C�"OPH �@\��ƴ���ۘs4"O*��e��]�QgC���"O��RPG�$Qٞ�zঃ(L`"Ot3b�&d��А�ńu��	�`"O�j�&�?�=3�
�v��"O01�k�=�p)#�
�_L�2�"O ��'���d㖫T/�X�b#"O�u�q䈍H����i,a"OTYP3+�&qfAz�	��g�MiG"OeQ&��-o��2�C�UZa��"O��R �<O`m!A&�J���P"O���1�	�NNn��$��`�$�5"O\�iG�8[F��FM ⊹��"O\h��HfZ�)Ȃ��2�N$"�"O�����Cdi%��5nPCb"Oh�W��,/X�3"G�,�-kB"O���Y!^��EX��XP�`"OD����@�9u��-uț�<D���'̀8k�>��V�	MXP�;�M;D�؃ n[)&-`&��%vz���8D�z�̇��a*�L�e;Ŧ1D�4qQʔ9eZĴ7"���
V%D����I��@���XP׼�Q��8D��k�d�:�X����?�v�+s�7D��0�D= l��k4oҸ*���c�!D����cR&_D�A+1y<M$�"D�3�aۗd��`⧊�,�x��,D��i C���B��̚���3 0D��2Bi��.m��AFMIT#��2D����"Q� a��	n@�w�-D� jƥaa�OAq���q1�pW�B�I���	�b���yz�,��'�s~B�	6
L��W.�'3P���NZ�w��B�Ix� ���O(>z�ARO3�B�I*s����s�3#�@�����o��B�>��1cd�L6��4
�ē58�,C�ɔ$H�a@o�:���(��;�@B��1B���ъ� p�"Gi��\�2B�	#�Y�ő�u+B��S�P�U�
B�I�1E�4D�]{�cP�d�C䉊~�F�hOx[���C�I�\��`6�$LF�v�˧E�C�I�<s� P  �   {   Ĵ���	��Z�tIJ(ʜ�cd�<��k٥���qe�H�4��S66<9V��2]����dY\�.R�	X�S�	)�6����ܴz
�<1�O6-l�,�@��`�@�-�';6��:�n,d�\�s� V�]�qO"8�O<Q!��! �h���4nE<�F�N�r=�I�EG
�'�4�B d�?Z����'^\����,��'� 9s揑\����GK��~+�%�rX�a�Y�4R�&i�'"�4+��_}��l>Q�E[)�^�჉��%��c���p�T�� e�'!�1ٔυ�&�n�ͧ�?�������;�����Z��Q��c֊j��y�!���~��Q-fP�
C����$9y�q�E-L�C��"#Č�wM��z�#��/bF�`�!Kլ|)d����2��01^3wh��Cw��*:.� 3ͅ��OX���d���d�%颐P�տ|�����:v�� �v"<�� ��;ZϺ��U�ؗpZZ����7F�O����g��!a�$Ϡj����TD�
Qo��kw��˛�O�u��OD��G�=I�ZH��	���keV�0i��I&��O����։pz]@�J��t��9��R��OlQ�����?! %����#k� /����U̓P��#<��!�D�;I���F�Jhd��ҳbC�$R�O�DRL<��#ޟ��F�?�����9V���b��O��bW�i𨍁R'ո�?�F�Jt?�'�~�-{�E�Cn�&k���eNS�}�I�qOI���#<!@�.}¨��E���[V��&$}��k���D�2�O
i�����1/ܼ<K�ˊ�D�(]��"�3H!�D�� �  ���!8��9ňA5��#f"OF��pC��4G�M:���f�Y�4"O���P��5|Pܩ�AP�s�� �"OdP�#�Q;Sr$ŨS-WR�@#�"OD�C�����[#��X��mK�"O0�5DF7�Z�r��	�(�����"O~�`"��1L���˧Z9�D��"O@L�F$�61F�Шg�-#<P�b"OV��Q�3����속Q"��'"O��9���SX� !.Z����"O�='��Xe �̋<~h8e"O�E1�)�*f�IR)��~V�D�"O�Z@�\�sx<���fB��s�"O��A��6*��qg��8e9�PXd"O��&��q���1W.Ʊ4z�`�"OfdXC��x<I��=gr���"O���֬ў3�    �  �  �  ,  o#  �)  b.   Ĵ���	����Zv	L����0R�PΓ���q�'��}�@ _\�iPt���0�L {�'�*�Aǝ9k����шz[���D�Wh����H%4�Hw$	�D�`��+N�k��Ԃns�(��Kļ����nY�1� *j���KD�L ЀU#d:�A2 ��E�l{ �BzQ��">7:X9HC����k0����;c|(���$�\���q�g�&�:i4
�W����Iɟl�I՟��_w`�7/��8"��*\v����JW��^7M�O�U3�M�a�}��ɝMVԴ	��G=a��U���
}j����AƦ�t�R$:���ȢM�i���D�D8:�u"7B�@�;ӧ�%����'�J��F�'���|�'�2�OJ�cdڎiG�l�U�PC�ц�D?��?��SF�a��L�lFr�
���xA4�Ƿi\J���$_���'���%:��V*�`��.KO��	�m�gR]�	ޟ��I۟�)^w[R�'Y�gB�~�&���P��P7N�:�@��PF0&z��d�+HU��Af-�*��1@$��P�(�G*R�H�"+Ո7*,����*R��E�10��E�C�_Mf�mC�Ig�7�G쓓?i��$�+ZI�qFZ$��vƅ�a�'Gb�'��IZ�'�Ѐ�ub�4;J��B H�~���ߴ�?a��i��Q�hp� �
�M����?9���M�Q���ɓ̝;?2޹���⦩�B��՟����p{�̖ӟ\�<����qI��`a*�H�c�9d��F{��ߨ�h�s���D���7�
�5�R^fў��%�O�F���<k8͊���?}/�����y�C(� �0Kպ|��@�Pb�>��>yӞ�L{� ���J ��-&�U�c%�>�umD��V�'�T>��	��p�	�����3$ޜs��E�7��yr�4_�^�Y�㘧��d�XY�m�	}�:m�B�ݯf5e؊�O?]�GG/*�ᐬA�N�������삲N�O
&�"~��O�-*��ݢ���H�j����yBȋ?U���iW9z�d�$�1�HOvTD�4��0#J�[a��p��Ѻe !��6�O��DW�Y�\Ę���OR���OT��A캻���G�/ڮpq��ϼI�$�+O6�@�'T�H��O;4:��q&̿?P"DJ*O�l���'��9 o'vk|[!H%"��p�,Oֽ�e�'����	a����q�*�*�����-7g!�$wd\�r��
B��t��e�a3��|zN>Y��se��g�ևK�d����ֱ2�<�7k�
�?���?��l3���O��~>y1��O��T�#u^�I�,��`Et �sqx�������dD_E���Ȅ�ã(����F9�O��ӕ�'��m�3m� �
����@<m��J7D�8f� R�z����N%hـ�4D��I�ՙv��h���"�j�@�>)b�i��'�НhU������*Xf�}�*F��4/�l(�3J�N����� D���@�RV��� D���"'�!D����ʈWzx=t&AkH�;�k#D��bg7� m8��M.h������#D��;d��
��(��Ʒ&ƶ��0	"D��ЅdRW�@�[ ��m=V���4D���ѩM�0�ĉ�«%fŀ�1D��z"ĭH�"s�K^�	�T����"D��ٓJ�/g�f����h��A�"D�(�0b�7.V��hf��-Y&��Ƃ"D��sƈC���0�<��i[P�/D�H�G���s%]1d�~��B/D�㑉�
QG�EM�'�j�Zb:D�DH������˅�ظB�>ј�`%D����i�h�քIV�Ĭ.� %A�#D�4�M�xٺ|R��]2a��`A�%D�� l�1�8;t,�6Y��%D����)��IV��� �%g�H��'$D�D�d)e�h�qbM�`��0J#D� �#$B>r��T���?!������#D� �a��)����gKɩha���6D�X�G�Tk5��C�F�����1D���蒐Bvn�R
V:��D ?D�����ʨ/X�� cߪ=¨!$&;D�@ʓ陼W�Hxs��@B�@�;D�� ��c��?D�	��wx{"O��X'N��(�H�6�ĩhqP�"O�m��!��F(]�d�D6h]���"O<9S�+Ͱ�����T-LaP-v"O�-�` 'd��/Ȥ:z�{"O`{�K  c0ei��Z�~AU�A"O�Q����9t"�
3�:tr$"OXS�� 2W�h�$��n��y�"O �Q*Vjvl���S�����"O�1�7@� b�u���0D� �g"O�yCG޻:�T(zģ˧3Ӿ5A�"O�h�#Y%5�J�q��ZM�"O�Â��7��x�@& HD"O���D(U��Y�&�2,r4RB"O��0T���xX|l���%C+���"OR�aQ�֡{�Z�a�4��B"O�E+�n��Qgt�� �_�y�"O%+"o�_�����'ɨh0ؒ4"O�
C��_r�Ha��8@�%�"O�<��FL�AY������$hU �9�"OXTyv&�'hI�tPw�� ��U؆"OAA���mI����9��H:�"O>�8��2�Zm�H2J����"O��2��G*��5a�ʙ)T�N$*�"O�y�G te| s�"��D��s�"O��*���q��va��f�h��"O^\���2	��H2���g�����*OP���X�T�Z�ɂ
�%| \�'�,�˥bݶ3/�\���~ ����'bx,Ɂ�P# R��Ǭr
��y�'0J�� �)z�lȋH�p$e�'�V�"�]�F�� D�D�AI��
�'�a#���j�	����s��`��'>,p@�5T4�� ؜Y^]��'�Tm�-��~u
ՠ�#�� d�'&����-�����JQLLi�'2z4�0�,��|�3�Юi� 9�'8���錕]�J�rc�Q); ��'7���Gk���������,��'fBm�3�J�)����� %p�k�'��(���I�>�u2©��^�(��''~�I���*"e�]�%I�1Vռ�[	�'3��:|�Ш��	I ���'B0�i�O��K��1HR�7z ��)
�'#FU�#��0� h ���=D�����'��P�-�1�����-�6A�
���'x�t�T�ٚ�lH'�F#~Φ-��'~���%[�d�ʑ
�:~y����'=�!	��U}�}!A_�t���b�'E���3�6E�
�A���i<V�x�'O8]�u�O>�&YBh�f�<+�'�҈��\=A���"�1�NHC
�'��Ya�$�@�1�Ѧ	����'� �;Q�Fx���1���j�H�'iV�(s'F$X��H���:ǘX��'��yXU�٢-�Q��8�*�K�'�:� �^�M����v�R7"i�
�'1���a�H�h}f� j�`��'[�4�S4FDvu��d�&T�P�'�����L��@¸�qM�6v&��'E����	)]�A10A�0�L�y�'Ʈ�b���`d����?�����'�Y��T��Dµ�\6�d���'��@�眡P��mٔƅ�F�@��� ��0�=���n�6v��$"O�!���!x1)vηh����D"O��	 ��&��5�PM6��԰'"O �����F&�P�c��x�H��'"O�0;���f��#�L$p��U0�"O���l/�n����>l蚵"O�� e�U+1:��F�B�,q��F"O2t��MZ:pPAk���@U䤛!"O�P⋆�mp��	�$����"O%����	����H�z���[�"O�ס�,���n۟l�8I`"O�(iD_�fmR,
��L�8� ����	$R�ҴG��AΡf|:}�SD�5~����IF�yB�/G4�kG/qG\H󀅈-tH�p@��]��H���44�V�A0�ؾK]�y��I>��B�I)� ������QQ��7_l�ԑ� R�`x�'Py���f	��|X�e�!d��j����$-1<O�d�%l��*z��� %�ϟd,�3$���ɖeǾ[��"��>D���q.RY=^8��lA�<�� ��8�$ɢV�F$�E�ݑR��Dh'�7ʧYH�	�->�
 �e�'钄����E�7�A�F����-QY��s��M$>��c�mӾ$�$c�����>�>�3�!�.4,5���$@��Ɇ��܈ǅ��0Ұ8JԂ��4@��"­8܈	'�������B3LO*�)D�R�����1L7�0�9��'�4�Ѧ�!�`���ߡ���q�����cG��b��s磚��yRj�co��/쒵i�C�x:���O�%i�
�>qt95��8G�9I#�?�����E�0�(ad�of�w�"D��!��r��Pp����Y����Q�L�)3(���o��.z��y����c1��@$oD���W"����U��yd�B�P<d�*(j�.�k�����@ A�X3`���Vo⹳r�	�1@�0<O�}@e�(W�4XT��W��2b��� \|:�hA&�\�X�	3�PؚX�B-G42T�y3-"��4�	�'S<9�P�&z�|,���v
���/O����C&z��(JS��4�,:����O���kAo-����F��6^4(�'�,]K�N&`��sP+�t{��H7�$j�UbnIݦ%��fߒWi�O�j�O� �1f
)k�6�u�9PD�O��5n)�@Ur
�mѶ-��l^� `����DQ�A�e˂LMaz���%�X:X?4$	��6��ԅ�i�g$�_����wF���9Ãoр�����&Ǡ+�d�X�O�/@�C��H��=���j@�"�z���'���::M�L���ϓm1Q>�7�C3>f���E�B�\�Ӧ�%D�p �D�@T<`�`/�~��iA'r��h@��Ov�	$�H��ɆRZN�Ѝ�=]��D
�cG2j�B�F���g��pŔ���=�7�O�`��#����=�BȔ@�xE��ϋ.�h��Ŕ�����8xa3�g�O6���Rm��b��W��z�"Ox]R��  �u�W�C�3_vU�W��ܷ��T�qm8�'��=1�n�s	`�Y�I*�栅��E	��N�@�$4��#џU�C�E@���'f�>�ɘ`��E�@�Êd<�xBr���U��B�I�D3̕�Ƒ�V|R%�A���b��C�>������<�FEa�菣y��C䉕Tp���L��/��h����C�ɘ:�#����2�T�SR��.G�C��"8F`Y5K�4*p����V1?�C�7�p%�ub�2 ^��W-V���C�ɛ��S�cY�"�X�I�#|�|B�	s�l��/D�@D��0��G2�0C�	�	�&�ba�V.1w��
�"h�PB�I�c�ï��2#�I���@"(�C�
6:~��ʩ?�E���0 �B�I%FThfN�˞`R��:"�B�I#o���e�!(���q2�C�~�C䉟YĄ;�(S�,]JiYV�D+$�C�)� ,mi��ʡ�޽��J�4 �kU"Or�� ��-8bQ����%k��y&"O0�5
Ο'�J�HE��$Z����"OZD�ClηN ��$K� �N]��"O�mAE�0;��덧<��|`"O��`�]3M'ư0��!x�����"O.�iV���!�`�hu�BO��L��"O�0\�(!ar�F�Ab4刐�D�<q"� ��J�C��J�� eV�<�&��)2&���,��f�S�f�<�@kX-.{��'���=�ɋ��z�<�D�u�tr��5�h4��Kt�<��6V�2��3%0BfޥP�G�p�<���_�Yb��pΚ�-K4�pe�p�<i1f7�Hq��L�2��	�Jq�<�sΎ�p@B��bG8���q"cXI�<QfNވwr���qe�V����Rk�<1vO:ZG�3�	�f�=S���c�<��8�x�8qğ��
���C~�<9V��{�̉�f��v �Iz�!T������z�g�ϲ5��,�';D��0m�9h=b@���6�J�I�-D���
�U�8��b��7e���7D��12�1RZ�ţ�bC]4��4D�8�AI�$d�L�W�#p�8�Ѫ%D���0	Nbx����G�!k��q#D��3�XS�>]릃O�9��ZpI/D���BԔ*�.�pmY����0*,D�ĺ,^r t����*?�zQg+D�\�(��2{���@�G`���6D�|Yw��{`�-��-C�˗�>D���h])|@��A�)��*@�=D�0x��VKԤ�#�R�J<��K�=D�P�����
�+4S�V� w	>D�0h4�Nl9���'-��g4�{��=D����)}��T@�e�$6�p�A�5D�� P%��k����O�f�����(D�p�^�܉	(zS�Q�}�B�Ʌ~�mZsH�2�� s'D�+�B�ɖ;ps$A�*�����&fC�B��&�];�`J4s,��b��R��B�8D`y�SZ�hܳwÅ*��B�	�m���P�by>���8f��"?A�I�
5������p>F1Rv��榙	�$M�=�r�cu��	{ꞰbF D�����4tov9rP��s<ٚ&�!D�����ٯ>�P��@"��tn?D�8{d��s��8�H�&U�F�Zu>D�(*�cRu�� bҫKu
��V�?D����*r0���ME�>2`n<D��ce%�[D���F����3b:D��Y�Iز�Z��k+Ks�ʐC9D��Za�&�l��Pe��X
���)D�\h��Y���`&%ǬS9�As"a(D�dba�ʪ;tdwN�g�ر' 3D��Z@��8\�5"�)�����['2D�PEKd��s�;��,��-D�� ���4r�ؠA祙�8���0V�)D��
1o�9�P�w!��|��)�AO&D�t#q��w0��pղ[� ���E%D�H���2|������_;$��R3o=D��9�&�SC��s7o\���&D�r2
Oc�ֈ��� 5nx��[P�%D����!� 1&T����C0w����a#D���ī�Yn�L�a*�& .9;��?D�� �P� lYG6x�Z�oʱ)�d�"O����O�-ahb��J"t :�"Ot�c儌t�H�D�:$ k "O�5���C �y!� �~����"O��)�$J -�h9W�����R�"O ���Μ�~M��HÍ�F�;�"O8�p��6Xth�x��D� "Ob���+�w��kAhI>2��ہ"O�t06$�68@�U��K#ּm��"O,{��z�!&,�-c$h�vCï�yB�OP�ځk�m�s����@�*�y���F�z�����5��ū�ˏ��yrH���
�RQ�4�r8qP����y�lFT��@�:�h@�g"ޗ�y���+�m���)i/�P�l��yBܟ?�^��%
�N�#�FC�y�(Ւ�32� ���
>�y���JRrbu.��`e�`p�GY�yBa��?�E��bJ+[ -��7�yB�F�:��0� � ��𠰅ȧ�yB��)���)]�x��s�gԵ�yR�A+62�xRG��&��`�U��y���Bj�p�ǒ!���@R&�y"��:���ȧ疬�\�Pm��y�͞>g��t����0}���y� �0`�~��G�� �:�	U(Ε�y� s�+�Hxk�;1oU��y�L�3F�DJ�np�3�H�y��Rr�eRA��
_��e��O��y��\�p�@��l��S��� �Ԍ�y�ڋȢ�pP��Jݬ�
�E�>�y�
;Ң�I�.�*�2�,��y�厓r�H�95��4jX8T�̞�yB�O�{�"�Q�C�#����K�7�y�S;!a��1"J���{+G��y�C\#0d���B�B���D��yHV8 (L�ǰ �t�
@�K�yhI!.���Ն�}H�p�A^�yR��=�v�g�Z�����V�yr�A��PYp� J�"�N��yR�
�(襤!!�ü|��}�ч(�y�a�i@�5*b�j�d����0�y2JQ3Y>"�l��e=TI�6�y2/Y�P�W���]�x��ӓ�y��=M�2�����P�
J���.�y2I9h��XB1E ��妜�y"�|z*LAp,�@Rj��CA/�y��'�� �G��G��s�'��y2���q16	H��;���t��5�y⡏.ZHl� �l
u��ecE��y�j��W�|d��.nR@��A.�y)��$��xP�U�F��5F���y-ʦo�1�@J��]{��ȧ�y�	�lN&X��GE�&\q'+���yBIU_/�-�"b�Ns�0��.�y���O�J�����v��T�7ǘ��yҨݦ4�JэN�t�`���;�ybb�t�*�4��Bc�?���q�'h�E��lG+H��D�Q+@�"��u3
�'dY��9B�hz 9-*D��'Nh������%X���#�����'�V�+� ʕ:
�h�t�"kO(���'�n@���X�*gtkD��i�0��'Z�d�C�͑!�p$ī�/�x[��� ��Q4�v�Z�JP F�`m�MX�"O\m��@4��A��-RIL��r"O8�����^�v��ŌY7v�^���"O()���I�{),Q%,�9�bP"Oy�p�;h(x	&!��=m�]B7"O��P���#�vD[�@�43l eiA"O�qk�J�&�XLqeO�+j��"Ov@
S�L�@\����o�py�"Op�`n��8%X��X
?a~1zb"O6L�rE�9?,
`�uO�*Jl�ə�*OI��؜KC筏�1�,��'�b�JҊ�_qR�W�4�l	h�'��@����+�|%ۗ)�$3,���'E��p��9Wz�����DJ�'����m��~�����<bE��'HZ-)��İI�FpP�hR=���c�'���s���?H@����8�P�(�'*�����#�<�`-���\���'��z�/����ᔘpT��'���e@ovL�cS��~��:�'�@Z�f��l�� Sn]�t�1�'ۚse�~޶����B�~��A�'Ϝ��îѻd��D��F̀~�����'FQ�G �x����ð��-n�<�0e�K��A��c�tE[D  h�<	3h~+ ZP�N�&����m�b�<QE��=0�6��!(�}�&1�$�a�<Q2�/A,�'o�
%jZ�:�KU�<���N-[D���OǛxE�����E�<1'�J��;0g�=[F}����A�<��V�u
ą��/��,al@�<A��.�|Er��2�X��h�e�<QPa27?<IxA��j�j�1�ė]�<�rH�,R�����Q7 ��FX?y��'����3�I�
�(�؄%�(H�L�	�.��x�9���)(��p��^�
����h��!S�^��0�B�Vt	��Fyb�*�S�D�P�O�XA��/,ԕ�r��9�yb��"zHd�K�,�@�"M���y�@��T�#�O:3�΁z���y�gy ���
}� e�jN�y�!e�X�Z���L��4���y�H�=7� `N[�M޾d�ĩ���yB�	?<QR�B:T��d�!�Ӊ�y��J�*ِ�P�ʃ7G�!a�yr@P@�� �r��
d { h��y��?Z�@��@���2cN��y�L�Yft(S�S>�0�Q���y�g;<����~b|���D��y�E�	��A�Ѐ�"nRR��V�y�掶c�B��M�hh�����yB��5�L( A�pYv�h'L��y�+B9TR ��C�_�g� �+�U4�y��Vm���Iwg�x!��	��yϞ�a뎠"L?l�,b�hV��y҇J�FzU���M1d!~��.���yR%]�Z�r͉��rg<�h h\��yb� �ѓ���3u<xY%�C�y�B��yX� ]�B�.tS%��y� ��]�8@�G�8���YC�	�yr�S�4���
�i׻;G�DH�����yRm�k���+�iڟ2ȝY�5�y�*6N����0���d��y"m��x��9����9�dj���?�y
� Ը�&c@y�ACq��8V�|��"O`�!�D�,{�e�oǚڢ��"O���P%l(�P ��1��"O�}��d��R ҬpKUR�1"O����ˆ��@���ĤXMD�1�"O���N�̻�l�|>�{�"O|ڒ�B794�r�KP9gW�e�"OJ�rE �?N���+�.Q�Y��"O4��$��I��X��22E�m �"O��a/;�f�ɗ<+;�ˣ"O�y���̉�4�ːɅ3&<-�g"O ���F+1�`���A
~�ʵ�C"O�y�1�Ԡ33l����@�=Q�s%"O������T���U;a܂�	�"OT�!1j_�p��B�ޠ2q<�S"OJTs�&\�qzfI��G��]<��sV"OtP��Ƕ��$l�>����"Ob����S
I�v�[�KQ(1b�"O0t�ʇ�(4x�eh� lH�"O������6jeM�4cO���"O�x�ƌ�0D�+́�t<�y�7"O��+m�;4�hRv��P�c2"OXu����.{�E�C��Q�H�"O�����)�~��2�����(�6"O`jK�4Ƙ���^�r��P"O��$F�Z��G�Ǽ^��1�"O�hj��a�Z�s,��xuʣ"O�D��emҽ�1KC�f(��"O�ix��٧/��i���N�����"O�%�B���]2���CM.#�f��"O�Z��� ��S����ϐ��"O�)R�,O�5
1�։���e+$"O����I�\�,�+$(֓E�<��6"O�G�U6C`�@��Ɠ-���RA"O�䙖��B��8�V�T-f���'"O4X�A�ʝhMB��sǊ���piD"O�RQ B�D]�u2��@��@��"Ob��DW�� Ch_�v��ܑ@"O aP�#�4f�H�@�'T��P�"O�а���cB�p��NW2��5s�"Od�bۍH�.iaFIP��i��"O���4�ΟS��4�e�/llz�"OxY�f%M|0 L��� ���Ѓ"O(�Z��<+�p0 �(W+y����w"OL����ݰQh�('��kh��˗"O��9�g���B���^&V��#U"O��ʢ��`'& ���A�KT$��"O0���
  �   }   Ĵ���	��Z��vI
)ʜ�cd�<��k٥���qe�H�4͒6R64<��c�S�VN�7(�;�(R���R�D��6�æ}��4D��d�<�O�7�m�H:f.�A��l�@��+_Ҝذw�E<C�U�g�0qO��yL<��)�1'�TH�40I�-;��_,m���E$!C��-�'�3K0B��=�'Ԍ�CvD�"<N��'������^�����B�-ziԸ�R�GIuy2�k��CEcAT~b���(���FoΊr�Ԕ���P7�M�������!L�<Iu�h%��%��iY &O�a#�Ov�BpLL�?�H0�aT�u�c�a����	�b�Nh� �<A�(E5`�l8��^�����C���!"�+@*Ԑ&gH��y��I�]"$��{2�Q�'4f�I2��*JSP "� �<jL�!�A�#<�&Ƚ>	2'\�)��I�h�PS�0H$O�H��΂�O�ѡ�{B&7Wd�޷8hXB�˂y��Yl�W�����&sܢLr��0G���O��f�<<�I,����Ȑ��X��[��,�gG�"
L$��
�<I'H!�8��⟴����/8��ؐD��
ne�EȔ���X��h���)-��Իv;��RZ$�bۺ�p��yrmE�'A��$��!a�T�\�4Т�C�o�&��6N���W�#�')8�k�$m�M�ԏ5�8�e#Y���5�>=�6͜^~8�iw��ɩO9�妟 z�ih<�&	��:%�u1�B�5G��K�{��e�'��	�O�M�ǎ�,��`
Rϊ�}}�G\��$�I;S|�x��.>R���&�;�
��U�3D�@G�   �'_Pĩ�7"O$��ɉ!bJʐ��ŝM^`�*c"O�u�掅$VŐ��F��ʅ"O�hp����y{�������u**da�"O�1����(t��5���\|�"ODC�*P>�~I2"��K��E:"OʤQ� �c׈XY�j޲'���kT"O\!h�J]L6]J�)�#w��)9�"O�|3�*�c��"�">/m���"Op}�bi\���UƠ�i�"O��K'���C��6m�@�"O&��s��@$��c&�ٖ�`JQ"O8+$���YHv(�!����ؓ"Oތ�F/U2@�J��tcϗ~$Mk�"Oظ	�]����b�Ѐ;J��3F"O(a��M��yv�_�2g��b�"O���7g�69��d���ԝT    	  I  �  �  *"  z(  -   Ĵ���	����Zv)����0R�P��
O�ظ
�X|���.='.�|�d. �h�0�ȓ'���RÈ�H���"�`�22/��3��x�.\ j9Z`����.)��hZ�ꏊZ۪�BW �0Y�,��i��l�n��zn���J��+�d�z�śK�N�$��"�,�Y�U�]�v�%k��V6$��H��?�4%���>\�	4�˃��͉sўVr C��� |���!Ҭ@�D���g�O����O*�޺���l�E�T�Bo�v�c⒢Tx��D��?��NZ4&����|��2�'�Nš�Ƙ/2�npZq$���ʴ�P+�j�u�mD'\�x��O@s��o�/"貸$�����3r��H�D&1A��F�<���ڟ��ڴv��OR����p�&Q`�f��̎7p b�X�G�>����?YJ>E�#Q�X�P3���w ޜaGT3��6��u}P�۫����<!�$X�*����åU�9�r#7T�dSf���?Q��?��uq��O����OT%3��#h��5♘f9$k� �.<ԡp�ݣdBz���F��¡��)B$D�D���⃍�h��IK!@���kHE؞l!$��O8	��é�VXh �(1�.�J�k�	!��n�ʟH�'���������g���u�Z�/|��{eO��2<Zٚ���Mkj
�hO��<1�5� �x��S<e�I��Ʀ��I��M�����ɕ2�hloZ����ԟ�؏c��8� �3e�p30
�/�,6M��a� ��OD�dX)���g*O#|
$����O���*RIg���i�BK�p��=	�`��n�ku��9�Q�i��1cÞ$"�Ub"��8C/Pa�'*�-u�.�Gy��8�?��3O�F�'���vp �i�H�M*p�3�H_�p��F�'u�O��,�4q��E�1*7�}��Γ�n/�n�4��y�S�&�>	���w���B��H��)� �|��c�u��iR�'���O��Y)5�'���(X�P�᥈�'�z��?\��7��wRt��3�|�>�׌L=B�Yq�A�(ЭѢf��X���4�S�OHb��<;��zS�E�YinH���',�����s�ɧ��V �e
�0Cb���v ֒u����n;D����M�|�VL�ŧ�2Z���?�I�?�a#G��ni��Hՙ@đ���A�M���?� �5f�t< ��?����?aǷ���ƒ�#���q�| ��ƅ=\��W����j;�O~�����{�||�fE�'px�	5P���2K6�Oޠk�ET�[�ㆸIfd��7U�L!��O6ԅ�E���d	 \�	��Y�r�B�ɥ�J=�Q�\}��i@��=?�6��V���D�|�ʯ1�HEX����)�N��O:y09"C!��%���'SB�'42�]�����|�ԟ@�2��C,���p;;Ǣ�C�kJ���>yV�G~?�A��b�ٴ�Ja�^p�b�Qx�l�b,�O>4�� Š-@Y@�Ԛ)D5��a�a�<9��%3�l��Q�L$�^U*V-If�<� D+>��tP���r#���1LJd}�H|�(�O´�M�(U���!5��?�$D��il�bs  �r`��mV!bZ�	�'��݃@
Yn���+aN�4-Bh��'@�H`"�;W��+!��5a�
��'^�r��mzd�+%M
:j���' ��i1�B���i�dlJv�lmi�'�d����[۸�B�H�%?4�J�'�x�(�,A[Fii��"�����'���E)�G���	�D�v�
�'��#��G�!�B���&��u�����'�,(@�f�@ˢh;`~�`�'| A��Su퐝9��J<C>��R�'A��sI�ZD(@S�;u��K	�')B��j�!H��,�%l܀g���y�'�ҙ`��B -F�m"�F�b+b���'���gL���Y��M�OX��'.��2�YFT�	E`��'@�'~0H�D�L�����_��d��'^&��י/n�H0�]�?�d��'A��)ᅆ2��qu`��+J���'�B0�@*:������ҮM#B�y	�'�bX�5�ɲ'g��X�gW/L�D�:�']�d[��b�0�2�cH��C�'��c`�g,$��&\�Ee��j�'��I+���\A���A+F{�����'34��4c_��Y�&K��n[P��� \pQƌ��q*p ���T0V"O�� w�W�7��!#�CQ;~{$I�4"O�3�"��P�T9��<uW" �p"O�1b�}�T+���GX�23"O�	����P��֠@'S�l8BE"O�R��L�^Ȑjp`�8^Y��"O\��*��Q���J?s���"O>��)�D1��ܻ<�$x��"O�qZ JHs7�e���@"�R�E"OѪ��ܩ;����j�Y�R�r�"Of�iך+Fz�.֤a�J�4"O�)z�
[�`+V�;�k=o<B�*�"O�E���?./�{W �B�譐�"O�}h�(ʹM��٣�4M�j��"OBM���cV�9�"�ǫ7��p*�"O�����b��T�D�q<�p��"On=r�K�%=Na��D!]N(�"OrДAM�P82�0��å
��[�"OH�:V�+��q3bb�3� u�S"Or�+0�̎[m~Tq�.��U�d"OΠʖ�!m��� ��4<$��"O�P��� y,\�q��V����"O���#MÓC�!Pe/Q+���[�"O�p��)��A���7$J3]L<�i�"O��M��$�D��������f"O �s"��>^��1��5�$�	�'c�1��ٓVN|���dD�ar�C�'6�9�`E�~�N�Pg�4'!�		�'s��s��5�$ѐR�P}x\�	�'�\ X��� b��ѓg� L�:	�'(đB��7N�F$C/:@���'oШ�"��[�vL�&-�"��'nЬ�`EUY�D"A���p�'�t$�G㛊-�<ZW"@� �H�Q	�'� i��HZ�Z���O�4:��4��'����5A�I\s�`�92@
�'ᨐ�aE�-x����Ƃ�!k�0�'B���« =��T��B�S����'�\�Cq��� 1b�bԬx�صk�'�~��Um��v���a�\]R�'����bR�;ʹ�V�_��9�'�DK�ZLfpF�C�;����'�2��Ư�6 �����k�S�i�'}�%	E��^ �T�d���`2�B�'��B"��G-���K1
3�"�'�l���]?p�D�[t!���>�[�'��=�w͕�X�ї��L��	�'��� 4�$vFѣ�I����	�'+@���`I�360q���S�k7:�1�'¶Mru^]E���G�O�e����'i���C�L�(�W
�.�����'0lD�<�lsb
��.���M�.�	���Y�'j�Z���"O�㣅:L"^�R�)�;�2�:�"O �p� �k�a�V�>$��4"O��U��?�Z&�
>q�h�4"O4�i�-�S�~���!�7|�.��"OldbrF¯^��� "�䈐�"O�9�� ��xzDЛt�I(�L �"O�����$\�L��d�v#�D��"O*�P��R�� `'��+7�9�"Of�8ǎ�4U�����ӲR17�0D�@��</���SԈ�v)~�R1D���&B�4Yx� ��! (�W�0D�� ���t*A8:�����12� �q"O>�hu���Y�-��]r���"Op��wDX?e>@]�R�] <{�)�"O�hbǙ )�f��ꅪB��8�"OXx궢���j�)�7NS�Q�"O�q�I�5I�����)X� Qf|b�"O��j�웇8z(�Д*��Ba�h "O�� ��֣=tn�ѕI�9Y�Y"O��-6a�2DF�z��͂rݏl8!��6x�ܹIٿ�䴣���f!�ě-'�L� �O��-�h��#�ыy!��еD�6�0 Y�Mmމ(`D��~!�$ޚ�<�K�M�(\4�h�-ִ$a!�D
�A�s��� `l��D!򄘉+�h�D�'K�r���� 9/M!򄉉cN4=� ��u��sdg�!�M�;��%��fKC������ɺ>�!�����#&d�?e�
Y��)Y�!�$�9n�,i���4V2��h"5�!�䔍\N����W�Ze3.��-!�$2¢i�E�T€"b�CN�!�D	��l�ҲjD#=�
M���	q�!�dٸP�*tk���f��W��8!�DB>Z&!��
29�*�����iT!�$�4E\@b� �'�L���b.8�!��p�9
�H)m�~�FL�! !��ڀg��eb��Q#�5x�t!�D?nô����K +�� �k��1r!�d�fU�/U}*�u�R�D�!�߂m>౰�B7w*���4�I�KN!�S$S�$)g���5�t�0��tB!�dE�,ܪ-����Y�$��׊$�!�M�o\¼���%Fc
|Jt�f!��@�Q>�]��BX�w���L"i!�$n�XQY�HIT`P�B-B�!��r,%RE` �V�����ʝ'w!��<N�(���K2D��}�a(J�1h!��ޘ#�N���[�JJ�n�/L!��N&:`b��.Ny�Q�.
�"�!�D]�����7�'��#��U!�$�!]�兄�L�x��L��PX!�d�@Q�`p���7��ʆaʡ1�!�ĕ+8:rKB��%��3���7R?!�$�16�,%*�阎@���GA�B!��X0p�8��@_(匁0��LF!��2I��m*L�4�X�T%�!�ߜ2�V��΍� �v���gT��!�$�@Q���Te�;i�R8�@l�)�!�
�-��M3D�6b�.�XG��5F9!���g����0��Iq�)��n!���XZ�*��I i/|8�p�Z�]y!�M�l�����HϦ-z�AG-D�e!�D�>#spx��M�p�J;��I!�D�=k���e��*��+�o��!��Y�$�R���	%�H0�� .!��4g��y���"	x��F��PyhŰ2�Ը�@��e���(B���y�Nt�VL1���3����u��=�y X�,�x%Q�,��
v!( gɄ�y�M53����āwL|ysf\�yb��'� �0��=`�x����*�y�[Xk|�3eîg�h�"�
�y�ʅ)�Ι�P�Ȥ&8��¢l��y"O���d��J�$d���!�0�y
� �=ڶ(V�a�ѳ|���8�"O����^Έ[�A=S��84"O @���M��A��(�h��uy""Od��E�<Ut�jwϯF��(F"O�P�$�&&�X�C�	�:Y�l�3C"O�v剆~� �1�6p>Q"O؁2FdңDj�\$�5��[3"O(-��I��=2J	���I�*C~��@"O(3�J�{^�|�1(U���A�v"O�l@V��:�R=���x���:W"O�Y����7*{n�i�����,`a"O�m�=��݀�9%�PM1T"O�+R`R�3���Ƅ��m��ԉ"O�̩7"�%Z=� 𡑎L�x�d"OvZ�J�Y�8P�ߞ$�*��"OB	w-��v	�1�#,.��Q�#"O6Q���pY2��+S�=�x�"O��Q���ݘa���j#��´"O�a�'�,��`#�:L��L[Q"O���S��)��
��;p��)��"O��Kp X�,8�CA%v��J�"Oڸ���W�Jr�d� Zl�Z"O̡��J�7>@��aL�O���"O@�Ip��<C�QK����8��f"O����ER�k��
k@�/�z�"O.�KC��^�����L�-��z�"O�(�I�2l�Q��a�1^�8�"O��Z�*S�`���R#`����a�0"Ox��)�!h�mć��a�̰��"O.�+��QmÎ�ۆ�B��
�CC"O�Ms'"�s���#e�f�B:"Ov̛"뉤A����vM�=Q�<pc"Od�%�ܱi�n#4\"%֮hhD"O
�K���l�@�fM
�%����yr�5r�:��bd���)��ݯ�y��	:)��Q�rI߄L�h�k�Jͻ�y�hD9��B3��>���P����y��/=G���Qd�9U&0�� !;�yb,�_(�<��ʵE�R�S��*�yr	ߵi���۷��E���+�(���yRC��4�!�l@�2�[F_*�y���f� 2�zy�A�vK��yBa͎E
�p�(�d�̈"G�X���O�l)Pd��g!�%�fB)Z�Je���iʠ(z5옃j�ԙ*�FKQ�e"�'0ã�-U�E��)Uep�	�'���҇�Y�&AQY�$�8I�z�Z	�'=��K#�h��s�h�
I��X�ǉ$D����N޲��g�XY7����"D��S��F������8bc�����5D�xW���P���ZeH�`8D�pJ����[�u(��
2qj08��)D�Ȩ��A�EZJt{ף��Xq*���O'D��ba��t�VЈ���m��`�+(D�x1� ��Qx��òN	ZRHɂ��'D��a���l�"�c��C2����7D��{p@��.�١da�&=
���6D�@c�E�G)��Ҕ��4���u�/D�41��1g��1[���!Q����"D�̠#��;�2��¦&+ش{b-?D���7�*V"p��2F�O�h�q *D��;��F�;J���-8O@P��1 >D�2WLO/'�d�IQ �B�4����<D������al�yv!��&8��M(D�<�F��.��I�Q�P�])#2D�� �uIrCX!�d�2��C�X|�R"O2u�V�,&83愖�+�B�"O�a�p����J�7��~v���"O���U+1W���˝Ws4��$"Oj����F!xF�*�?_Y���"O^5�#C#vP�e���Y�Y��"O�	��E� ��{���!f~iY7"O�]��FS(�@��2C�UcrA�"O����*Ac� !��</j1(F"O�-2e�8���$-E#U9��3�"Oʭ(�]\4��Ŭ�(;9�Y�t"O�!iݿ��M�0�ґoPd��F"O*�*��P�C�4���M�oG�Ź$"O�$�D���/�N�
�m��~CX̓�"O�e)B�֜,|����B�D2�̹�"O��� C#Dx��9��d���S�"O l���o��d��^�?���"O�yB�@�i�q��v�P#E*OlE3���:S�Ԕ�%�QeB��'�@���$�H���|��u
�'��*�6Od��r	� >D֬*�'9�4��ҁ_o���Q�Q�4`�}�
�'᠘bVh� ^9�� L�1�*�
�'�t9a͢ 26��K$��p�	�'}�he�\�m�s%�C>T�	�'������Ȑp�Z-��N�>��u��'��(!���$8�LB5bE-7��s�'�d�0&�mN\<���1�ZHc�'��A�K��p6D)���5^�!�'!2�� �g�A�'�+o�\;�'��y����<V�0AD� '(��'Ɗx�&�MT�t	���Y�nb	R�'�T���e��;�ƕ	�jٍ�D�'oF�aҤM3�I�
�/Y�~q!	�'^& ��牋2�(�Kdl��d|
�R�'��  ïUf�D
��Ոp�t�;�'˦� G$[���aB@�ڪr�Q��'�4��x�#�<�W����y�GY<kHz��$O��	n1y&9�y�P?r����Թ+u��p�eA)�yr瓽 ��p�띊+δ���&��y"H��ho�k�B-(-��Z����yBBBd�8��ˍ����g�?�yR��5@ibT����d��F�$�y�e��\{$���[��@�gF�y� 7K�*@���W�UM*-@�U=�ybF�*6���2e�ȰO9����yү�1w�LЁN��;F�`��/�y��S�2 -"���/�R�Q��y�G�P8>��sŔ�Vr�"R�J��y���m��ǆ�KϬ8(����y��=���mF�H�1pL/�y�S8>�LT�����>����+���y�%h��	�n�-/ez�@!�;�y�� n���O.�8LH���y���"(ߺ�S�a4BͲ���5�y2%O�4{lz�(��&�
���g��y򮊈B6����C]��"�*�y��Is��yQo[�
-����g�?�y�GG	PЍ�t�����F��y�nJ�$�T;f�Y�4�nd�d�M)�y�.DL�3� X�}�^����y"O��>�8��#C��4���Ҽ�y2��9��|qDm�en� �����y
� ��)��+�8��
78�s�"Oz��g��c�(y{+��o�`�s"O�92��;ͪV��-r�Z4�1"O�
l�
kfƼ���D�
���!A"O�ٺ�⓸J�e2���,5���"OXH�t�W>a�<�{j�R����r"Oص��C�	e4�H#H�K��$��"O
AE�Y�'�0�ČO3h���"�"O
!������3�]&]���&"O�zɒ�f,��dO��P�8""Oz�P�F�Z�w��]}�[b"O���)�Y�4�hG$C;F�-�"O.�0,H"'���"�U�.[Pt3�"O����J�2�P�Ru"��$!�3"OF�K'���3�Z��%⃶,��(�"O��B��pJ�8Ro2��i"O�4�Ug�"_�t�!���Z"Oh1#��,������B��X�'"Oj2��"��"rNF�a;긣�"O�hroǠ$�x�k�=%4V��f"O@�R҅R�e ��{4jĚc!���U"O<�g\�:4*��i�4#�P���"O:�1g&ňN�*� �J��O�$\�W"OT	B����+�#�}�""O`0h�D֖��I������"Oc]���A�Ẃ�k�tQ��"O�m�z� ��t��CG�	!��ǖ�h@Mٵ'@���fÀ�^!��U@pІ����l�Gȑ�i�!�d	�C4�8�%��)�B��w�!��1W��QDX .<����ҪL�!��A)RX���$�˱�%/��xێ��s��cB��jX �v�]?F�4�� j0D��Ӷ"G�4���)\m�ޤhЭ�>��4�tMr�b
�O��&!	>:V܇�ɛ��	�4�\�4��lT�A#V&��v;�C�	�"Ϝ��ԉD.�*�@���C�ɸ=������=���D�����-D�(�G�����`�(7��e�'D�x�&��e!�ȓAM�Z4 ��%D�x��$<M��u��ɻy@��M$D� 1��"C/P����Ąd����<D����Ԯ	�|y��1*��e`1m;D�x0$I��x@#�?[R�$ 7D�@;���%�"u��`��6!F���4D��	0kT��#M�(��-��E6D��kC����p�:E�I�t�&D��9�D�i
�d�%�C.W�<���'D�d��ł�P�6$�L�:/����#D������mVs!�G�6��ĺ��,D�$y� 5I�|`	fX�o~ ��p�<D�H[�K p$>�ۧ*�0ҕn9D�[Tυ,r���Cgj;_�Ҭ��!"D��&%I3�9ӧ%ՒF��t)�  D�0��_-jZ�[$$##�TQ��:D�(A��6�����'@q�`
�#7D����[� I��$]�x�s"�"D�<	%o�wz�*Ϯ}DT�A!D� a�$��*J�) �ԁ@� D�X����jӂa�&Z|�,�c��8D��ҦE��'�le�FO��\���.7D�`K&a�5E�8�paO�&1�<d ��7D�D�ՆE:�&�y�L-?B���9D�|rd�^5v��çT��)�m+D�� 4��1l�/ǰ�	�ađ2ͬ`Sw"O�;�"�I�N�˗�%�Լp"O*���N� )L��0�LC.C�zX�6"Or�`,H�ry���J�A���"O�)��%2p,E��I
�G���3"O@�x�f̘�<Xu(IP��MB�"O�x1u��c�TKҩ��>�,Li"OCP���}2)+GbV�[�`TRw"O�U�F�i������֐F�i$"O.Ly�FԸ3�<`��A#n2���"Oڡs��m�$���ι�L�{�"O`FE��M?ʈ�#��\�TsU"O)QJ���t3�C�^�8)��"O����d��n�3g�D���"Ox	��0e��A�]x!
M	�"O�x{����1��uS�G؅j�S�"O��#�!8~��}`w��b�Bu+7"Oи¶$�oN8�0�EA���,
�"Ot q�@A;�`�ᑣGi^vTj�"Ofe�栊�"56�hfh�\R�Q�"O�\!�MG�Q�\�艣l��`T"O��0��;$I�q���D��"O���jQ>x��@sN�-vt�,-�!��I-�i"��m�t��&��2[�!�������l�B=���ؤq�!���T��\����x̦�a!��Y�!�d	�[�XI�BZ�O����&���!�Г5�~��޼Y�q@֍S'LfC�	%o��B�e��u�^��FS�adC�)e|��8n�V!���:#�C�I:;�����aD��Ri̥ 3�B�:Z�F)�N=.��}1nޗ}��C�	?}u�4�s�D5q�9����:!C�	�Z��lh$e��z�A
@G�0Z��B�IwV��Y���^
H���f]!��B�I(nS��Auj��5#h���Y8/d�B�ɗzL��P���30BM	ń��T�JC�	{U���C%RPqVm=}4�B��?�>�y愊%2B�Ѧ�--�PB�ɫkJ���	¦t(C��69�C�	;
�*EA���/^��P��%=B��^k>hp�4���c��_��C��,��T[��ӯ\�� ��V-i�C䉈xv��M�5$�~�Rdʙ���C�I�5)L���� (�X�4�ĞITvB�	�76cƫ�yT	��_(C�II����u�PuRG9F�*B�I�J� P  �   ~   Ĵ���	��Z[v�J�(ʜ�cd�<��i*<ac�ʄ��i�%m�lhx��ǔ	��6m��e��9�����N28��J1�<o��M��i7���Xy�Y�o��<�����|��<z4#��H����4`d����G��#F'z� ��x�L��*���i�^}�3��wfhj l��wh�2�Ox	�&�,�z@�`y��	&��S��UyR�K�Ը��� ǰp�4�E���p�lt���ۿ�Mӆ���yRɀ�\3�u�'_\��i]�Ɂ�� ���6�8x��1[�� 8P<6��\�paS�;�n�0䑟�Z�K�>�������%�¸ͰW�Z�D�ji��a韌z7�;��{5-�<�r��	 ^\݂¯�5��dV�1��q��� � @i���	�8qZ�L��`���J�{�B�O�'1ZlK�IE)if��"��P۠�2�j1/�"<y�%�>QP��xD�M���Bg�����h����O^@�{�k't��$
�vh�ٷB���M��d1�^�b#<I�-�j@�!wJ4KGL�ZI���>�B)���7
0�hf�V-Ke�ibᮉ)|�J��'J,iFx�DIZ���9!�ʔ���p�����&M��#�V��#<aê�Op�Z�F^,<k\�P�	R��,�s��M(�O¼�J<A��_4`w�#��W�vtk���a?A�7��OD�#Ep��n�R5��gnҮ1�5�`�'����i��E�ũ��M���E}�'�~�gn�Y8��T}<�Y��Y!dC ���R�^��#<���-}� x��t!�*8�ޝI���1��D��O0�ډ�K ѦMk�$�
SԔ�L,!�՞ � �  �tтqÈ�x��%�"O���`NΦ)�T�E%E=��ɐ"OdM��ٖ"
 ���?^���D"O� ��v�|=K�ذm�.���"O��� ��������ױ-�|��@"OԵ0�Q�+��@c�]5�����"O40��킠.� +#KQ�l��@� "O0Ar��1��A�䩈�"��Pb"O L�S!ˁ�dc����Z�"OH�z%	׬P�ĹB���azG"O��!%�	�\�f����KR�Z�"O���0BD S��x!�
�FLU"Oa��1]����#�m!,�8�"O*���D��e�dⅡ1#h!�!"O��Q@��!�d: @J)g�T��"O`�i%���u$�%�i�j�"Ou�����8R�2i8��"O�iVȁ1���Ҏ �Ln�m�0"O(����>&`�g�C� xb�"O��BO
z!ҽi���Pm�P�p"OiK�lXV�`i��h�Qxt��"O0$� ��\� G�n�af"O��ѡ�SgC
��Q�M$Yx]k�"O�|E	3~D�f�ͳ2>J�C�"Oa��fB#ז����h��	�"O�`�u��_x��x�����A"O��{�CS�~b��B

�(�FPe"O��Y��W�6��b%��o�$T�$"O�iH���K��-�j��q"OF���T�| ��!��h��R�"Ol1����j�}Z���R�j1
0"O<Ԫ�+[��`KDj�ٰ���"O|��
S�R�~����_�jqK"O�Ȫ�L��p8�X��,�8�R���"O<`A�'ð���`2F���"O�$�ٯ���!R�]=���"O�x�@��5�JM��I�O/�,�@"O���v'ģ~��G;	�X}��"O
�g҃0~X(ö�yIf]��"O-p��w:�x4G� B!���"Op书KŅ�Q0V�?d���P�"O�a
Ul�Px�����j�8�9S"ON�1�3 Z�}9�hR4Tp��y�"O���T��$9A��-�,@�"O�5`ㄹ-�q�2�� f2�ۄ"Of�ZP��
O��ëƱp�����"O �2��L��% M~�"H�"O��1'៰DY6�n kâ�"O@1 �B
��v��v�(X�X�Q�"O� *EX3B��H��}�w����"�"O���,ҹ;,a˲I�>�h}c�"O&d�7-X#9�mYa�Ҳ-_]�U"O���@�ؤiݖ͉W��"_ �!�"O�;N+r�(���	ƞjAn��r"Ov4���.C��Y:��҈1����"O�ܪt���fQ�]	Ř<|�Q�e"OH��4gI]�~e���416e�U"Ot��A��1g�|��vO��Hl��"O�8����N�eR��M"�p�У"O6P���B8�<�'�*l�^p��"O�hR��N�7��l�u̗�^��t�s"OD�Z���}�z!Z�M�=fv�Ȫ"OZX�F�[�&5��
��D1����"O`�Cu���B$@𲗊K Ojh�³"O�A9ݞ.:D��0jʋz�Lh�"O�X1���L󦴙`C�-(�,{D"O�� �+�M��ܓ�A�';�
`""O<\� CP/�p�"��3?�5�"O�,Z�U ����ܭ&��p�T"OD�ȏ��p��ga��~��m��"O�0��화�����8�jq$"O�u:gD\6 ;�@�U#��2�����"O�<!!�	=�Fa;EɃ�ؘ��"O:"�(٥����J�+�٪�"OPC&R/�ĉ��ł%}r���&"O~jai�3�HI��٤uU�i�1"O>!Ȓ ]#0s�h���2Sp �g"O�|@�� \lH1�t$�e��F"O�P��(׮cYZ���,��_��"O>�Ke���@�٥�	2eH8��T"O���A�xz��q��D�G���"O��3��Q/6��!sƭ��=���v"O���ťl`�t����A��Y�@"O�p�Hϋ%"���vH��"O�$o�ٶ��¤K�}� ��"O إ!G��Eq�C� ��h�"O��*p틎+�ԱH׃	�F�,�b"O�ER�n�R�S�?Zӄa�"O�s���>殡#Ǉ���Mjr"Oԥ�$��)jƃU==x�"O�Ő�E5j�R͓�䗜/�ȸd"O�hA�bv��UAQ�-.�E��"OEz��Zg`mi�j�34?ZP�V"O<�����Vu�ӊ�e/jeB"O�h��ǅ(dH�1Xg	V*E�|��"O�({g�٥s�9�'c	o�V]33"O�3�	U���=�A�-�h�3"O�(Q�#��L���+e�
�5����"O�U�� �ZW���'���nԘ�"O���`Y�4��H�,V1��K�"O(|����pA�$�� olS�"O�p�7+ GW��2�)ϰjaԔ��"OVpCFc��N����1L�Q@"O��O�C��'εKݐ�i"O>�$M�4*Jy��2o$>�Z�"O$�hS��Lh`���I�6h��jR"O�i���N�,�Z��!�N�7"O��k�IO7���+Y{�IR�"O���wK��k� �l_:.@C"Onp���%f����6K\5r6l�"OX\��N�1Vᚁ��&��P6"O����C�<	I��׷d�t�'"O0�РhE�5\:�G�rq�};�"O� �M�dKڜl��9����-{Q�1��"O���e�>`��+��23���"OZ@��^FԸk�g3���U"Ox����;�n�[U�g�@�P"O�H��� ��M�W��%a�5�"O��jY�1@�e`��O�1A���"O�A)�
��p{�͔x0�:7"Ol8�Z���� ��u�@�"O~�G�8IS���J�\
ViS"O,���"��~I	Ā#�8]2"O| �Lk��b4CSA��(�"O��ؗ�F-0~ c!�>���{w"O�Ç$�#n��(��@Z�UJ�	jF"O��!��  �   p   Ĵ���	��Z�JwIJ(ʜ�cd�<��k٥���qe�H�4��S66<���EO�f b����Ɗ_)2$���Ϙ^86�����I"�y��D�<!ĊɠH�hp"� Y&:�`�<W�0��D�c�㞤IR�ɼ4��˒*W6�����;qz� �m�=���V�(�`[���D:vVuR���d��(4�ġ��$F�ar�L&[�B!�!a���M[T�Ĕ0�����(�Sߟڝ�aa�!RЁg�\}���G�bU	4����e�cc�!�O�p\9��u~��o�|�R!8����q%�,r^R(�u �!0�m�R�O2� ��<�y��]��3�gÉG�
��Ł~}b�+S���ӨU�j�Qv"�&Gdh��g��>�rq�=IG�8�<��Gj��נ-	4���,h����c
��[�S�x���س.H#!Z)28 SPa!}��K�'-���=Aw����4]�Q�G�VX�v����b�	"Y��\@ԤWDxF�b��f�lyh��� Z*b�|j�ቌO�I1`,��E+_F��6��2X��˓i��#<�0M*�I6���ņ�h��k��7GD♀�����r��'�2���)L/���ˎ�ZH1�y2�NV�'��$&�4�rĕ�N����k ��5�V������I1C�'*v���cbpiTh_�@��Ct�r@�m��Ss��y��YR��'�8�-O뮼�h�_c��Ya�%�8wJ�ko߄|��y���]>�O�3H�(�4� �D8z��cn�!�nt��&�>9�8�;Ǆ#<���L�]�M���;J#� 1B�d�<��h�= 2  �"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  z  �    �*  h6  B  �M  fY  �d  o  8w  T�  ��  �  R�  ��  �  )�  j�  ��  �  e�  ��  �  r�  ��  ?�  ��  ��  v�    � t P  �* �5 �C `N �V �\ c �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����O��=���Y�+�F���eIq���JK\�<1!( )�%p@�ř'#�ܙ�TW�'w|��I�E�J�����{�)"�/�F��B�IX��-Iӯ�7�ة5�Jba�u�	�'XJXw�
P��-��I[� �l��
��� ��{�*\">d 0� o9f�:�"O8����e����!(�"R �R"O
=�kZ�t�:f�C(kA@B2"O���1aT�l��yj'&�8l��u��"O�"3�	K�,@A�˽\u���%�'�剁IQ,h�A� 
��T@* �L���'!`5MV�+�z�i�ݕ.G�P"��HO���Q��cD������z-�"O�܂���u�0"
]�8�Z���	��0<��	XX���0��r;�}k�c�F�<	E/�����b��B���t��E�<��NʭZ� �被�������j�<�R�)����ɀr����F�e�<IcY�n��,��%�T$IUF�M�<QCK�@�������Ip��EB�<�e'��%�!A�*Q�)�THX�@�<Y�!]2yΈ��� �I/�P����p�<٤H�<��y��фk���Bn�<�1�D|L��a��=�m0�yB�E�`+X����I��A��y���':�kQ��h����y�+�F,|��Z�0�i���Z��yRE�!���h2ԋ+
����y"��;(?�h��c�!T��	i���yB�N4�M(���M��9�����M��'7��b)Ÿ4w\��!��=L`����'@9{�`4Lb�,`�թQ���'���(6�Ӿ�x�J!��:����'*=�� �g�H0�- <PMz�'y�0�q��.)(�� ,׃
��"�'n�؋��O�7G��\�*T����'>ys����?ڔp��o֜��C�)��<Y퉟:��|�go�)r)l����b�<!cn�/@���bd��u�*E`B��x�<!2悑D�\)��D�2�svMIu���p�{�cY>/QB��e��0"U𥣗�y򥟏=Ҧ` ��Ns�X���=��'+ўb>i��C��0���2���?� 	 �M7D����ǔ` <2A��c�� �V����xB�Zv�L$��,Ωw��TI2KK��y���c�:|�!K�>̨)�d0-M�=�'9P�	Ǆؑ0��H�Pm�;R��

ד��'��a)�A	>#�����9!�>D�
�'�����I�O��� 䌑�q ��'p��˲d̩��,�@f�Յ�;�yRK��|��� ��wI���V���y2���q�h���F�.#Z|XƬȻ�y���L�\�c.M�%�������yRdհg_�Tٗ"�>�IEfނ�y2��^r�9�%�/�0�0e`Å�ybOڪQ�n��T��"��Q�տ�y�gS�+�T�sdo�3_04Aլ��y� �?/l��nK� Jǝ2�ў"~Γ�j��q��	���[�
�)|R��ȓEA�y�h5T����Mȇd������?9g/�r_8��֎ط1�@PgDx�<�U�ъl��fS4+�8 d�r�<!�B>p� K�V� �z`��$F{���Ŕ<M\�0�	��j�d%��7�6C�	����b�)u-&�:��]5C��/}����LϪm'��9�Fߟ6 D����<Q��-se��#�_>v���z�<�N�	s��L8'U��hS��t�'#�?�hd/� d,��7\�xiSp�7D�� >}6�ͫP�D��#�շc�`��e=O��Dz��IG	�������������D�Q�!�$�]�X�k$">n�R(@'.�&F�Ї牑I�I�@̙ �`쏨V�C䉪&D$![a�!��E�	��B�	�N�@�0s�E�$$K�	��(�pB��Z�Vi*R���N���F��C�I�q[�0�*��Y�0�I=��B�ɷ)�b}�r*K��
�ę3�ZB��8Z���B���Y�&�Q2,6�_8��?a�@ăD�X�@'�!&^�vc�}؞� �Z��j�41��p���-VH=��<���ȓTZBmqB��*J�����i�&�m�/1�	[�Ok�̸��&Ze�πri�	�'~l���G�E]y`D�B'T�
�'R�}Q��8k1�X#��)3���	�'3ġaǦR��jY�ťܱ|���	�'2\q�Y�&S�$T�BvRt1	ϓ�O���#f;�6���F	{eܩ9�"O��x��Ž��,Jc�ךw}�!㗟|"�i�2��>}ȱ�U?Eɴ���Δ��@�1�Cz�<�gC� 8�`�_'/��I��u��u�p�$�>��O�X��̙ƌ�(1�q��2F�zC�^�C��R�z���!@ǐdJ˓�y��S�\T�d�����C�G�q�:C䉸:��br�ʄ0�l��G��dC�əZ�*!h����`�H7cǚd��B�	�>x֤b����R6� Aj��(��B�	!g��F�P�(��q�M�(��B�<6e��b�D<h�p,�y�B�	e�̉����<>�Xt���J�CƲB�I�Y�X�;��ݡc� �;e<]�B�ɈZ<��4�T�����$�B�	�Qiڹ�R�D6U8���_�K�ZC�ɐ_�Ȭ�JK�QT��wR -�"C�ɷ8e��X��F��Ԫ��"6C�Ie9he��Ԍ��ȉ���3lg2C�I�6��$��CT�P���:�%�7^`�B�ɶId�h� z��L�< ��B�I
T-� 
���d(fp(@��F��C�����
�/"�bV!.��C�	�	i����S���t��&��nz�C�	)��4��J� `��f��6B��.�����A*b���ʒ�n4�C�lR9
$�I�T�شk��B�	�+� � �BO25h�!�5N��Fk�B�I�jhy����8 �!�*Ћ�C�9S4�@��4&��p@�*W��B�ɑ�H�CA�u���+�d9�6B�ɹ!hآ�R�tȐ`��=s_>C�	�~���'*�=;*�P�`*T�-QJB䉠6]D�jt�9:,�T�k�?t�(B�	8Y=��Q�N}�,��lN_#�C��"�*Hs@�C�l#����L�4/�C�� X�@Y�cƇH��<�Gi-�C�I�<�Mp4!��F/�dA�f?\e!��� s.�IeD$-,��GŚ�@/!�ă�C�5@3l�})r�⣍:i'!��%	�4Xg@\*&$X�c\��!�DΛcT	�m��.���!@\�!��]e���ZP���J}rS���0z!��P��[���;w��P�Cτ:f`!��6�$)B��.�:�P��<w!�d7%6���bސ����v�Mb!�� BQ2Vk��48u#��5[����"O����(ð��4���Gߴ @"O�X��/ݷ���ÖHڤ6����"OAQ͆�a)��PDʜ�_Q.eS"O�Ժ�坎z	��;��k ���'r�'���'�b�'��'a2�' ,x��u \aZ��S�+GT8h��'q��'C2�'B�'b"�'���'�T��!�	�ȼRm	%xmF����'��'�r�'���'�2�'g�'�&�Z���=7Й��)�
	���/�?���?���?����?	��?a���?��E�)���Eo͕v.�����?	��?���?��?����?Y���?aAO�+P`�|8�LN�n��p�KR:�?I��?	���?a��?!���?���?y�$�3X��[��[dd�Q)`D�/�?A��?)���?���?Q���?���?�� ȣn�$s�[�S�t0��Y3�?���?	��?Y��?���?a��?��׏������[Z�*��D�L$�?����?���?9���?���?����?���C.8b��"t���b�S��?���?����?��?q��?���?Y�f�L�� ���)O�z��TL�3�?9���?)��?i��?���?���?I�e�N����ݰ\��	��%L)�?���?���?����?����?���?ač��d�4�j��@�^��,r!�E��?���?1���?����?������'�B�Q;`@ah� ��0�%�m��B�˓�?�.O1��	(�MӒ��5m-��*�.I�$-gAOuL�X�'��7M<�i>��@����/�v��,� V4ȡ1�����I״�o�b~R:���SD�)��[���f�G�E�TC���]�1O��ĸ<ɏ�)�$Eڐ!��J�
)��͈î:�%n�N?^c���Jt��yg ׂg�H�Ok��ږ��cF"�'���>�|�D�@%�M��'��ف4i&�bT[�&@G-��'�����Pa�i>�	/��l��冲s���ȕ*_�O�0�vy��|B�a�����_�>��#�㐈Tt��M�t~���Y�O���O^�Iz}bO}x�� �Ds�q�U�Q����O�A��*�#4l1��E���4l��d�i<�#W���h����fZ;���D�O?�I�(�&Q��!̫e�8�ףހ8���Ɏ�M��MXg~��o�t��%�Lx�Uɀ=%$�iRb�%u(Z����I؟̘�!�����'m�)]�?-31�<6K�D	W�2@%aH;a�ў�Ry2����X�*�������4������Ȧ](S�2�I~��f���$�H�sn��;& ���
�R����០���'�?i�^i.=+��F�( �AЗ.C�,!8�rnߧ-�j�'�U	��Is�B#T������	0%�9т�P�H�"�9%v.�d�<I)O,�O�lZ�f�͓U�iˤ"4��ʳ�C�2y�X͓J�V�4��$�OJ���O���Y;�
�#	 �(�3GB�J 6�f�ts�ğ!6�O����8(��H��s⍍EB�Y�#f?��)��<q���d�<E�4j�6g�����'�6g6Q���\��'H 7�~��	�MKJ>�0 \�<��1���.��j3�� �yB_���	̟���3��m��<i���?��Ѱ.�J\�`AV�Wnn��2�o�����hO�ɵ<��hD8Z��	̽k!b�
"j�����5q�&
���'E哜T�l�N�5e&ֽ#sM��2��m�������	�<9O|z�A��x�t��X\}ٱ�$G�.����#!Ƭ���s~2�'B@����g:�'M�<��ؼ-r�r�%�X5&4�5�'���']��Oe���M��$�2� !=��\ʁ��2$�=�(O��nN�9��I��M#ɝ*����)�� �Q����mZɟd��#�a��?a0O\�G��1�1(b~Ϙ!Qhlp�V�%%��Ώ�yBU�����$��ڟx�Iϟ@�O6�����]�Jl�a�(U*,� `���ʦk�O��D�O>����DΦ��3���ӂ�A�<|;`�Ө;`
��4h_��0O�Ş5���ٴ�y"0a��Y{�H!n���Zc虅�y�/��E� P���ݠ5��'��i>����F �$%�%x�bI)�V�DS�I�	�����ğH�'.7�F�|� ��O��$Ux�(4#���1��yH�i�$#P���O()o��M�'�ɝ��J�
�"t��)9e�G�3�
�����B'b�P�$@:«"?1��8�٩\w����v��	X�K��~�*rf��Y
���O����O���|*1@�N���'��EL�Zy��e��&)�hX �'�"6-�T�(�
z���4�������ej@r2��FX���?OXHl��M��'P�-�ߴ�yR�'f�<A� Ly(�I����Jq�9ᤍD��De�a�pN�'��i>��	����	��4�	��lpbQ�s����߼X]�'��7M[�q���D�O��<�9OVj�x�D�(v��!�v��>j�NU�'�R7-MЦ���ħ����$#hX��(a�J����߮�
$;s�9qQ���'dEj��'A��n�p��Vy2C]T~0�$O�@���D�@
��'r��'��O1�I��MkA��?9��������8��2��33�����&�'Q�'���?��4�?!FA
4r�^<�E�6�2X�IS4��۴�y2�TK�29H���Z�:���_wo�]�q�? D�S��@+b��r�M��g0j�;b3O��O��$�O8�D�O��?����K�̄iA��-PRP�92L̟\�Iڟt��4q�m�)O�lf�	�������U�u`�!N������mٴ�?9�gE	�MC�'$FY��ě-�=j���t�"���ϙx$x�G!ۧ4.|aJg�xR/�<�'�?1��?�ģM,R~��c@Y7U��!i�4�?����A⦱S ��8��蟀�O7���c
���t�u���m�n؀�O\��'3~6�����̓��'�*�ʋ)���z�N�tq��K�j���82��q�t��'���'�h���Tz�K>���G�\8U=&eX�j
{=����ܟ���ǟ��)�SWy qӨ��n��DWD�J�]3#��Rt�C�|���t���\s}s�,yID�ӭ�Ha���&=`��4$�զ���1�|lZ�<���J�}�3��H�(��'-�)X!i$q�h��J�)WI��'��	럠�I؟����L��F��Q�&��mٖĆ>a����6)�,7MX0:ږ�D�O���;�9Oȩoz�M���5�p�@d�5�V�ː ɬ�M���i��>ͧ���XL����4�y�
�*��5�` 
�R�= Y�<��e�2`�!�U�+�N�M>�)O�I�O�E3�Kb�89S׈��a�����O��d�O`�d�<Q"�i��c$�'4��'��d���œsvJ����g=�Uɴ�$Fy��'#��2O��
]�	�M.v{^#`N�ϥ%w�x�	�=����q`��V$R���d�­�u���O�պ��˼$=
�Ci�訃'�O&���O����O*�}��
ܜ*�%N�s�-e$ѫ{D����fD�v)�)e��	��M[��w@�)&�>N���UH�;MnԘ��'�X7�������Gq@nZ�<���FJ�x���V��Sq%�C�6��C&75�m�#D��䓷�4�����Oz���O��ēz`���B�!:c����52Д�z����7(��	ϟ@�3��$K�dɥ��j&�]"` �7��I&�M�'�i���3ҧQcF� �G��tG2��`�4�a*A�E7z���'8hH�t��ʟ���|bP� �R%�1Frh�(E�b"F=;�+Xğ���ş������]y��{Ӕy�l�OX�Ǆ��!�|`$ӕg�f�ْ�OB7'�	���O�6m�O������Q:$���E�.Վh���\��7M5?y�M'?h,�	0���56�۫w_��U��&
`ޡ�D�֊�y��'j��'��'��	κ��e����<#�HZ`��/2"��D�Ov��E⦗�#�	|�po�J�I=4� I3�
M�#�CV��$�ϓ����٦���|"4�8�M��O����E+�\���x��"@*M������x�O��|���?���i���pd�K�h����
�F�����?�.OF�o�/0�Zd�I��`��b�d�'\�A#	B34k���2�����O}2�r��o��<��d#A `�9�L�
~�"��d>r!d
\:/?�]+�O�)P8�?�WH!�dB9`Y*is �ya��s�4r�����O����O���ɶ<��i��5��ゾcG���ra� yD�8E��i=�	٦��?ٰT��ߴ^�"�J3�]<ob��5�
D,����i)�'�y��8O����(����'?���C�B�c6�R�.�\a�f ^�"��zy��'�"�'���'�i>Ї��4�(����^����D�T��M{�ɋ��?y���?)H~j�'���wG|yK�ʎ���A��� Ö4*t�w��m�<)�O1�b,� g�*�Ʌ@�D�C�M�B�(� G@4��I>��|!��''4D'�x�����'L\��
X6\��FR�
��iR��'�r�'
"_�$�޴cV�|K��?���r���kA�E#�9v�݂P��!9��J�>鰻iKB6x�@�'4�Z��2C�aB���"A�����O�4Ò�M�:������	9�?���O�$CD��pT���p�� ��#��O8���Of���Of�}���#��Z�5:�xH���w��4Y��F�܆j�����?�;i���~^�AP��V!VXHΓ?���Kk�Z�Ā��Z6M2?)���GV��� '�b��]C��G�X805^l{J>/O�I�O���Od���O�	�aTuT�t��@�i���`ζ<�b�i2�pZ�V���	]�'=uT�q£Ĥ:�jt��e��+�����U����4}\�5O�"}�F���D��U�>���D⚯b���ñ-�}~�ą_��=���{��'��	�>i��8R�N2D|x���/S���Q�	ɟt�����i>ŕ'��6��h�6�$ �(o�i� ���p��6$���f�⟄�(O��{�[o��L$���+ ��)*��A&
Hhź�1(��H�Z%����>1Yc�>�{�g����dׁ���!�'~��'Q��'���'��H3D8���ذdC{��s�g�OD���Or8m��lm�d�'�V�|���( 	�u�[��f���I�'����c�4�?��l��M��'�r�7(9���4�:pD�D�0x� ß�Q�|�P��ş���֟P����X�*L���	<fw4�V�͟\�	]y2By��x��O����O�')��Yp.G�s�0����y����'�*��?ܴ�yb����Oަ5��� 0=�!�ei�B�T#E��ԉR1�؁�O��i��?A$�2�dƀ>NT�u�C�\g�c��;I���d�O��d�O���<週i�$GH��7�̰�A���<�*����*p��������^�	:��D�֦}P@Mڱa5���C�X��(��(�M���{C`���4�y��'Ɇ�{�(��?�c�O� ީB�G�66��:A`ċQ|���66O<��?���?Q���?����i�+Ό#5*�5z��`؛*R*lڍ~�D��	�0���?���~��y�չsۼ���c�;")��Q-0�X7m�֦�̓��4���)�O��h��i�T� �N98��3���d�C��8O�rퟌ�?���)�Ŀ<ͧ�?��L.#� ��ş�V2��@�R��?i���?���d��XkLПL�I矴����~�^��� ȴ[����A$j��z����MK�i��d�>!"�Kb8$b�)�i7�!�aÊH~B�S���5C2�F٘O��)��YE�%*#���r�R`NL!#(�QB�'���'���ן0X ��@��ȋ��?*x�p�`E�����4)�*���OH6M/�i���f�-��ղ��a�j,��`�Бش:����'��Ң��=��d�04��q��jD��:���,a����Gi+�37�:�$�<ͧ�?����?����?� ��7�~�;��
!��(�FNO��$�П0˰��<����O�`�L;s�.m�2)!����>�A�iS7��q�i>���?�
W�L�b���(Do�
_zPE)H+�k��$gb�IU��<
Q�'���$�8�'��s&oڋ$nIЀc�/n�"`� �'���'m2���DZ��ݴ]�Y ���Hu�P�P���Z���3��)��M[�R�<����Mk��R��*tʝ*�f��U����D��M��OF���.A������`����K:M��H�8���,A��$�O��d�O��D�O��;�S<C7z��A@�0E�\"E`�*��ɗ'7"�w�v�*�>�d��Ӧ�&��8D��Ti(ŀ�ʎ%��l�F���<Y�Ov%mڦ�M�'`��,B�4����!2�(ɺ�+�Op��(ãК&PH�Ycf��n/8��'��i>A�	����I C���Z�-��-=�e02�Z%~������h�'��7-ߦg��˓�?�,�B��A�`���QoٶAt�=�Ӕ��OB0l�MS�'ñ��5p@�q�ij @��_Z���e�[f��P������i>�I�'$�'��{�k�ab��i4��'~��������Iȟ��I�b>i�'��6�=kƆȡ�⏋Bx�@C�F�~��Ku,(?��4��'U�����Q�ExJe �<-Av�b��8M7��Ϧu����A��?Y�ժd��	���D�m����G��^Y,xBp��N��d�<���?y���?����?�-�T��p�§�F�!�C�`B�dQ"�@ݦ!��韸�	ޟ�$?��	�M�;+�$k��4�,Ԑ�)�#0�Ʋi�:6--�4�����O��F�u�|�	([�N$)��9)������{ْ�ɐ"Z�Q�"�'Y�t&�@���D�'t>q��C�h5�Qb�;=���ҁ�'l��'��]��ڴ<��	����?!�� �p8��˙o(9�!��b�l-A���>�@�i6f���' ܙ �J��lա�� 9H�yÞ'�b�V�:c|�H�n�=��������oHB�$F�3�$�!��_]ȈWD�:W��$�O ���O��D!�缛��]�6d��[��'`X��"ʸ�?	�is$��$��m�P�ӼS ��"	{�E�'�:)6�T��<��i�.7�O�����u�6���papE�))��tc�j��"��/hq���U�_��'�`���$�';��'f��'Ӭԁ�'Oa��H5���K�l �^�Ęߴy��Y:��?�����<���h���%U�~xΙ��e��\��	��M�Էi��:�)��N��N�qKr	�򁕓u�d��;%X���e샠?����w����'W�&� �'�p�ڒd(eܤ(�g`��N	��J��'*r�'^"��DQ��A�41��!���KJ��SS�� ]M���+��&N q��M��b��>�W�i-�6-�O��[R��x�� 1D�t$��'�\�	��i_��O�A@�$W��r���ӣ�5��Ө>��	Vi;c�$�I
/�y��'�2�'���'�R�Ɍ��|�Eg̢i�h)�aJ�`!�ʓ�?��ihP�ɟސn�f�I�B)I��:�L<���WN�r}����O07=�j��dh�l�H��)Z���΂{!:]n�2�fB�]k��$�1����4�����O��$W�TkT�Q GD�i�Ɖ��;d���D�O�ʓp����95�2�'�r\>�8ï�2	rh;qW�
�1��*1?��P����4Dn���|ʟ��@B�K��y��C�@ΩP�A���~H#���s��i>%���'�T-&�8��Vx�n����8^�ppH&���	����՟b>ɖ'��6M� xW&l!u��h�v�����?�$��e�Ol�֦��?�QW�ȱߴUꂹ�fCA!-F.y��EK	
{5Z��i���ΰH�V��h���P�"����~:ƀ,B�:I"���8U�hH8�AN�<),OV���O����O��$�O@˧=���ƄZBB [�(���L���i�hm"rS� �	_�S�<I���#c�^) �ޭy�R�
A�$jC(%�$|��Ij}���bI2-l�3O�H���$|��UB�@�;��m�7>O�I���?��N>�Ļ<�'�?��K��>�A�D� .�~d��L��?q��?y��� ¦ik3' ß ���g �6np��v
]�Y��J�d�^�[���>�M�d�ir�>�,���Ȣ�!Q�uP%z�.Ec~�!CB�hq�5@����O�jm�I��C�1-�|؃EV:JG$T*5��4Sab�'��'���s�-�����r	�%j+`t CH���"��Z����':�f�4�\�a�iA* j$x�=p���9W��d�ꦝ0۴p�mӏZ���0O���3�X��'	�� �BQ͎l��hZ�e��r���+&�D�<����?����?����?��E<g�.�S��s��B$,����9�pc�������%?�I	q�����+�7PVA���2;B�h.O��DkӞ��s�O��Ȑ��N�zI1�҆H�ظi�%ղ{_�<h�O��q�&*�?a��=��<i!+(?9���1-B@6L��?����?y���?�'��$�ͦM�Q��˟�0�oJ<�(� �B�6-8�c壟\m�J��4x�ן�m�ȟ�1��͑x��a��S'WV�A��UU�
�n�^~���W]J=��k�'=�k,JKPB�� l
��}{�O�
���O���O@���O��� �S�he�`�AL'u#�A�ӂS����	ןD�ɮ�M�"�Ԛ���x�|�OL�
�$�#s� �pq��h���t�0�'�6�Ȧ���N�~�l��<��W�-y�\Tܹ�ȏo��e���
��'��$�t�����'q��'�x���E1f5���2�$��-"�'2V����40D��i���?y�����\�(by�FB�_�Xbe@ J��	������4�y�iFU� �B�"����ĝ��vdAFŗa$b(:Q���ӧ1�B�Q�ZAȬ�r��!
(JԹGK�����P������)�SIy�u�ذ�������1C�ln� N������O8�m�W�E�	%�M��ٶ
��)��$(��3ŧS!"��'1�Ұ�i`��O<��AD����x���J3n�##�ȿ&?�y.i�0�'���'�'�"�'
��1I��A"7�E�]ghY�N�mJ�K�4@x�����?���g?�����2#Աux�!��@c�<�4�
/7·i�d�<%?�84��'iT�ɼ(a"�G�K<�ڝ�f�=R��Iz��|���'J&�%�x�����'^$!e�*gRHQwD�0x����'�2�'�U���ߴy�:�k���?1�;qB 
�.P6��E`�
�N����>	��i46Mv���'[���酮0��8#ӯ�y�ƨj�O6�qP �G�
�I��ID�?Q�K�Oh=�3�R<J¥��H7���rw��O���O"���O£}��o���� �O�?V�����VX����v(���:O7'�iށ���ݐ!��1W��d�(q�Jh���4����'��S��B'��dT2�4s�'_�x9���WU�]+��ӰKŚa�7��<ͧ�?����?���?i��ū[f����QuO.=�C-&��D���	���Qܟl����$?e��<0��$�Ѳu�0	7h�_b8Y��O�oz�޴�yR�S23K�T�AŢ$rz��h>��(f�T�o9t�*���@,�O4�RL>�(O��Q�;t����7jZ4�Zщ�O �D�OF�d�O�<i@�i�F!�4�'
����E_�c�.���2W�'՛���~}`nӬ�oß�����	A�����,A��Kݕy3@�o��<!��]��i���'?���r�z�Ε)�Q@�)�F6�B�J}����֟l����4�	۟|�
��V��
��#�x�Z�� ���O�oڮh����<��4��'��L��a@�d� !1d���&�F�A�'��	�Mkg����@��-1�����uJ���թ$��#Q�jؚs��\���#a�'�<&�������'y��'�X�j�$�B��ؠQ�H�U*\�(��'�\���4sU�"��?����	�"	,:���L
O)�@a�HZ)9��I��D�馡@�4�yB�)^��qJ��.��Y�v'��U�G_�t��q���6*��w�	�Zb�*�2HN�t[�&BD����|�	��)�Scy�cg�� w��+[^E[�'՜g������V�j��MˏRj�>�ŷiT!p�h�0	jd���(Dj���@Cq��䟇1�7#?�E��$1j�)0����Rgf\Y��Y�Z�Ԋc,U�ybV�`���h��̟X�	ӟ��OT<p1�*�Є��&�:0��+�b��q:���O����O����t����AWXp��OtP�r���0H5o��MÛ'��)��3�:m��<����9��Y"��َv�.�2�O�<�3I�%3X�����䓳�4�����m���`M	�3B�`;d���<j���O���O<ʓ}��6�	�!3��'9RJ�p��q&�Ӭd���fζg�R�|҆�>)��i�>7q�x�'A���ub	� q�x��-b �3�'w2%�8W�ꡊ�
�6��d럪�{�|���$�7B���7x����rbF_�B���O����O��:�'�?���پ2�� ���$�z!8�F9�?a�iZ �2��'���xӖ��ݴZ2H���DG@sTQZ燑� ���ɘ�Mk0�i����7wn�F��lZ�Q8!���į�>�Q_ux��R��'f����|B]��ϟt��柸�	����k�`�޼����S$��ᰍ�ey�y�xxY��O"�d�O����|Γm]Bz"ߋs-Z��ϝ�?"�&W�p�4�0O��:���O�rЎ�@��T�'&c��q�T�����l8Ƃ��BQh�Iiy���*m���|��ٲw�H�M2�'	��'��Of� �M��ˆ��?Q�	�<�V5��;� bC��W?Y�4��'u��5����n��\�U�V�@p(�0h�ޔ�G�],rj�4#G�r�.�	П��Eb�0����0?��p+k�X3��=hU(�h��''�,f\���O���O��$�O��=���s'�H@��2^uR`ƀ��H�`��˟�I��MdZ��dr�P�OF|���-�`���H�*�ͱ5�d�0�'������Bp�������g1� �py�O�-��f/"�{B�O�?�C@,���<ͧ�?9���?)KE≮Dc� v�M��͒)�?����?9�8�d����?Y���?1���4A�2�h�W`�>c->�C������$iy��'���On���JQ\Tx�$��)7���'�OϨ� %��D3��O���R
�?�2�&�C$V�J7�D��|0B��X5�����O��d�O��<���i� �����t�n(��Zi�&�0]�*��I��)�?�g]�P�4RX��Ʀ�$.��U*yP�a#��i�R!��G����pcSeR����~jÀB8CO�5�F�2���� �b�4j�%[`h�QC@�<"�Ȱa�I�hgʕ���8��`c�	J���a�X��py��nG����K��+�VE�Ў�e�ND�`kJ��h��S�� �h'M@���d1h�1<���o�`�g��<�BgO�5���`�6eQ��L�!b��A�b��t5N�Se��LH��L�!��a!e�'?�@*�/�"�� $0 >�xв�	�<��!���B;n�У�`�3��j-�>�r�s�'
:4��X�HS�q�	�FƜq��@�a]�)HD�NЦI��؟��	�?yJ<�'XuN�� 
�*�����Q�|�F���`��'��G�s�T��Q�E��AҰj��,�����V� �޴�?��?q%�_�I������'���͗s�zl��i!SV,ŉW*3O��IWy�����'���'�b���X�0��
!z�rjeE�.�7��O^�pWo�N�i>��I��\�'�X�02��`�VR�lÉP��@�x�b�D˶<�1O0��O���<"b��Q���%��,�t�ӱ�84]r�XR�x��')��'���ϟ��ɾ:qFX�#M��@��@�ֈƷ,&�eC"�&�I��,�	�'�L0aci>�9�G�Į�(����")�`�&�>1���?QI>9.Ob�afX���2�� ;
L	d�B�@�Rq٣c�>���?q����d���<P$>�b�ˉ��dR�KV� ���Єk[��M����?�,O�D�Of����	�7+�4r�I�dϐ�+��Z#9�lZȟ��Iry�������k�ּ[�(����T��!�G�%k�'��ɧ1�,#|��O�fbѫ#�4Q[F�3@�^(�۴���-�,n����i�O|��`~���3o.&��f��.b�ԡ
��A��Ms��?�A&
���4�@����'͎��:H>�����W�'�F���4U��s2�i��'e��O� O�I�j����"J�$�`��#�4ja��mZ�Q�����D;�9O��<;~6h����<O"�b�v��%Lh�N���O ��P0M�T%��S��2;���"�K�iµJ�=�6Q�']�I�T�c���I�L�	�4�>��4
Y1"{*�8�`N�C�����4�?��#�dd���D�'��P���+�	��*��T�"iڂ���M��Z����<���?��� ���X�	�7f/�� ������S�j�N�	����Id�'���'��!s��
]��1pP�C�1Rx�&>��'!��'��Y��Bg"��T�>�$8�����0k��ݲ��?i��䓦�Վ	�ɷ4{:����-o(v���t&���?���?9)OXE��N��of �NM�&�1aI���ٴ�?y������O���RvP��^��H�M�&AC���7H)D�9b�iG��'I�	�EDjL|����1C�`�8&'M�c��<�wʇe$�%���'�ȵ���)�?�J�ؠbf�Q"���S��I�Q j�`ʓlȘ"A�iQ��'�?I�'f��I�8df����ɑo��h����1�d6��<����L~ʟғ���m�	:�v�4�03�q��̝��M�`�����']B�'M�4M3�4��avFI�W����O�	_�U�����C��5?y/O������O�P�n�x�8D�!���<dT��N���}�Işp����-���D�'k��O�PYC)I�`YuӥƓ�2jp � D�j�6�,hכ�D�'0��ORM�M�L�gü>!��	`�i��M݀\��	�I���=Aƍ��Z�xG͛�/�z ���}bmT9o!
�O���Onʓ�?!����AH�8�A(ɺT��$`JJ��ݑ,O@�d�O��D0�	���a��~j��a���1.g�5�Eї*���P�5?���?i)O�����Q������$m��d��|ʒ�c��_ ;�6��O��d�O4⟨��=$�4@(� `�T��Fm��>���;�d�C?�As�R�H�Iӟ`�'��c��z���T�6퉰1F<a��+���typV���M���'��a̎��A)J<�i�Uq��(X�%���	���Ijy"�'F�t��Z>!�I՟�Ӯ	�b𪇂Ίqe�Aa��(2�"%�	�<������b��' p�1���c\8�3��X� ��'5�#�5�"�'��'P�$^�֝�~\>��F)QS��҄�|M�{�O*˓kl)GxJ|�����U�b�rAP�%Eb�P����!7͝ß��	�����?}���d�'#�s�	@"����JV�B�F�Y"w�"�x��]
I�1O>��	4 ��4�S�-��Hr%j׏3J��`ݴ�?����?���	��4�&���O\���s=��!�$I�&�2]�lu��y��Cd��f���O���5��0;ƬݠQ�θ`��� vTx�R�
��,O����O��D1�uR�����h�:�a����szJ�#�JM�!F�\~��'r�Q����f%VH� �D�F�t(;CC��3�E�py2�'e2�'��O�d
=V�!�����!J"�E.����Z�6����8�	yy��'�mi�ܟ� �ܢ�!��fKb�G��Йٵ�i���'�"���O���FH�6�Y��e^1_ںe���\�����O��d�<��qN�#.����N�(��[)�JL|��E� t&�n����?��*�<�F�h�I!�������5x^�sfF��27��O4˓�?q�D���)�O������9�-�jcBy��٢[#�A ��m��?Ydk�-?+Tp�<�Ouԙ����~J��"��)Lh�O*������O����O��	�<��L��Ҁ@�m��:GLk|���'���0o�ƥ�y���J���R�*ч�<�^�	Q듓�M���*�?I���?1��J,O���O>�X�l�<3kr�2�EZ�L��9�3B��r'�Jc�"|j���~)j�b�:q�
Di�bW>E�N��лi���'���U�i>1���\�g8� @��HD(2���(r܀Ȋq�D�>y�~5%>1�	՟��E����&Q��iU�_�B)��l�����sy��'���'�qO���uI�:R���@�ԭ`�W���&OU�%Z���?������O0�d�B��j����Zs'�.H<˓�?���?q��'�4�牖�7���R���W���	ʵNa����O,���ON��?��ž���ɂ
 ��ᇁ^���S+�;�M���?����'B�M^*ٹݴ`+�P`��2[��@���&@+ND�'9��'��ٟܰ��]���'`(��!�b����G��-�m�!�h���:��ߟ�bm�&WHOVM�1�R��Y�́�LRH�h1�iU�`��#T&��O��'b��b�zf,�h���T���G(�8�c���IJ�eJL:�~
 ���C�`��į�1$�F�b4�Ds}�'�v<��'uB�'���O��i݉z��b�����!�|u�d�>���#K�A�DTw�S�n�*d!�I
,�Q�T!E��mچR�0�����D�Iܟl�Ky�Oy�#K �N!�"�؋D�A�R�S�|6m��N"��f��S��:ՎX1WRx��h�R���v�׭�M����?���!��2-O��O��Ķ�0�f��f����=:����CҌ��'��q���-���O�$���D��'�:�A��"o2���lӺ���<8�ʓ�?����?��{�$ �M*x��eL�Y(�Q0�f�����S�"5������I�|�IEy�I6��ġe�ݴn��y����z$iC�-�d�O���*�D�O����W�H�YդƸq[`�R Fo*
��N�O��D�O��D�O��D�O6�D�S+�	nڭ9���y�DL*��ؒ��06�\�N<�����?�2B �=/|�JB��I�9#1�Q7Hƴu�i���'1R�'�剞_��1��P���.�6�i��0L2`�E��o�ޟ��'�R�'{�A�	�yr�'��$O>��yS��!d��I$�������'p�\�������)�O��� �PB��:��9��LJ n�T��jZg}��'S��'S:P��'��	5k��@���E��M[
��U�`�ۊLz�\n�cyMF�;(P6��O�d�Or�	�J}Zw[�$9Ue�~	��H��4�?���r�Z���?Q*O��>��@b��(q��WƐ��HE�u�i�*УE�ܦ�������I�?遫O����)�G��e������!��0;�i�b�`�'�"T�����p4�@"�$��ch�����7��ղiE��'r��[\6��Or�D�O��d�O��B�)�*9P�G�
kh�k��^�X*�F�'��	�29��)z��?��)ߚ�o�/x���QM�ĳi�r�/�6M�O��$�O����V�T�OH�'	?u��9�Q�Ǚ":(��[�P;�$j� �'���'.T���J�s��X�pa��]�Z�q�cʏ
��*�O���?a-O��$�O���Z)7�C��;T��M�w��5v`�5X�1O���O�����O����<������I;E��Tb�f��6z��$R�R�&X�0��by2�'���'\��!�'��ј���l��8�5*�-%���?8�I�_����IΟ��'l��+�D�~��D�T�Ϥ[z���	�-5t��E�iBZ���	� �I.b���̟����m��ar�*8z5>`<��n�����	Ey"�T;0�'�?I���)N  ?���R,[o�0M9���8���֟|����`���h�p%����
���*L!~�`V��V�f�nayR�%2��7M�O��OZ��x}Zw�t�%%Տf���a�Z�g�x%��4�?��l !� ��S0Oz��}�����0sT�BkN7��Q*�C����*rCN��M����?���g[���'�D���˰y�m�Ձ��B"s��D�ہ1O2�O��?u�� ,�֍Z�lX�WV���lȍpA���4�?����?�q��b��I\y��'��$@0�:�js�ȬoD����M�."��f�'l�	�r� �)2��?���0��$`��	i�����,͈�ã�i����Qش���d�O�˓�?�1=s!�o�=0��`��0�Ҵ�'K\$;�'���'���'@�Z�$zu�[�$�"qC�X�R�������S�O�ʓ�?�.O����O�����<���TJ)6Ͳ�"�ѵ;�}�s2O��d�Oh�D�O$�D�<)k����
q��2���:��"!CB(5��^�P��My��'gR�'��C���WȘ6d�N��w�(J�h4�i��'�"�'��i��с@^?���B�����I6n��E�����n��dZܴ�?Y.O���O�������O4�$��~�3wlT��`X�&�S��<x���O��$�<a�
�T���Οt�	�?E1� Z�h'��.���qE	V�&�-��T�������I,_����?%Ac`��uc�X�&��T�>�c��s��gġJñi���'b"�O�>�Ӻ�r���U��J�m��\�G!�������h{�(`�43���=�ӁCM����LW�k͚�k�J@���7�ϭx*�n埘���P�S;��ĵ<���)�n��V�U�����Ձ�O��?��I�{���۪n��Y�*�lq��ܴ�?���?��D#���jy2�'��E1A&�h��ȣJ�h��fA���V�'�剧L�)���?	��1A��!OE�6�c�'G�8���Ÿi0�G�/`4�Oj���OJ�Ok,����ː�T�e\� i�	���"�L���EyB�'���$�Ag �8�f�J�Vys�,R3p�*��i0��O��1�$�O���90j�:$�C
^"�ز�*$#�Bh+��6���O*���O<ʓx^&�K�=���qV�����.5��)�N�H}��'�_������ �	�"��r4��фdN�6��YB@�Γ\�
��'v��'nBX���܆�ħ/hH0��@#`�h	��R�3��a׶iq�|��'pbB�yr�>1f`C���K��H�̌�`ud�ئ�I��'�XM:0O<���O��iA8WM<�9$�O�T"�&D�0�:}%���	ȟ�X! ���%�p�'j��CmH0 T��f�=F=F�n�Py�0��7�Gl�t�'O�$�>?)�N�*xdT9ʴ�E9tv~�{gdTЦm��꟠�̇ϟ�&���}�g�8_r�Z� �2�r%H�C���W�K��MS��?1��*�x2�'�`���h�7_Flx�*
h����r�α �7O\�O�?����q@e[�oϲ�B��ڨ�F��۴�?I���?��N���O����|0�b\�\�%I�!P1(� dz�Z�O !�E�t�SƟ��I֟�w�G(R{�Ih��B4�ڵ3%γ�M�EJd]h��d�O8�Ok�W�C�h�ô�ث0gܠ���ܓHH�ɐ%�p�IDy�'wB�'�ɟr�ق�݆Y����<a�@�1g���ē�?�������O����OF�J�ə!9;8%�穁�4��2�&�l��<����?L~j�	˛(C�I�� �~�P'��?eF>�����-%�������Py�'���'��й��'BR���F�9�2�+���`Ѧ�qK�>����?�����/5d�%>	�QM_��.]�5KG�'�`���+�M#�����?)�^.�� �����~���͕!��x!ĕr2���iH��'��I�!b@�N|���B��Ϻhx�hAƁ�L�n��P�H�W�'���'<��K4�'�ɧ�)�7/��[�H	�|mlY�/�=SO��V����҇�M��T?=���?���ONh@Jɡv�v�`�K�H�u���i)��'�Jp��'�'�q��ِ�K~�U��n��� !����/W��7m�O��D�Oj��Iq��˟P���H4B�@ Q�S�B��˕�^��MS�l���'����R.V�;�%}�tRT�FHG
�m�ៀ��ß���H���?a��~rK #����܉t`$���#���MSL>A(��K��O��'�҈��L��8yTGA��M�c.).�7��O:���B�r�i>qGy��3���q����Tnl��sT����Y',�t�D�<a���?A����DZ-��e
�˙#_DJe�v��E�< ��f�IןE{r�O�A��I��J��k'�P-sBց)��i��'�r�'cB�'j員k��	NȌ�񶅏5��b� �f��M�޴����O�O����O�)�!�]����
@ �T��,�y����%��&��D�O��$�O4˓zv>����4��$x�M��Pf��� 2��)�7��O>�d4�ɠ~6�c?m�g�Ƅ[Y�4;1��'�hȚ7�p�<��O��d�O�@hA��O����O���L�`���Q����G@&���B`��П��������&�~�iaҕ(���Q���0�j�mZR~b&�^��v��~����"2��@���§�irA|q`��i�����O�i%�)���b:���+K�D~�B��ǯn�`���	z�6��O���O4�IPV����7G�4Q�\B�mD�C!����̘�M�q��_���F��Se��Qd-Y
J� �S.�l�� ����@H���<�ē�?����~���x레zf�	��T�h)ބ��'�j�+�y��'��'��y �G�.>�:C�":\���.q���ā uf�&����۟0'��� �R԰B&!p2�`�n�`��H�ܜ�<9��?�������n�٨5,�<D����J%�A�v�;���O���<���O���E����a�9r	,�K2F]�=J���D�O���Ob�(4�O���c�Mx��� �5�D��O����O �O����OT �U���r�F�Z����,ϕRC��SD�>����?!+O����6YQ��ӟ���j	��޸q%k�_�n���9�M������M��	��xL�~;����`�SM`�`�쑿�M����?	(OF�����ϟL��~춬�gl�9D���Z��U��� pL<�-O�����B���N�Aq ,ҐlX>+jpEc/H��ݕ'�x![�Az���O��O��8M\訧��3y��Cq�,uܐo�Kyrh��O���abУЕ'�bJ2B��2\��rP�iR�l�R�|����O�D��'�<����� .p���]3�%�f �gl^��ijBx����۟����Y*��z��% �1#$J��Mc��?��^�x,qלxR�'���O�)�i�p�\�#  �
�����$TK1O��D�O8��צ ���bl_{��H�f���"��n�ן,�������?Y����r��oQ����D	=>Զ��j�^}r���'r�'�]�Q��.=�qBd��n��y�)B4R��K<����?�J>�L� �a��X5�`@�=iIŬ+��ɟ����8�'y�iCE�k>��,�Z�
`ـ�'}�B��N�>A��?iO>I.OH0��R���W
߽5�p�2Q���5`�ɓg�>��?����S�'��&>���m�<z��r@�ހT\������M����䓾p<��)59>4�$��!2�n@J�`��]�Iӟ��'5���g&��O��)�A��d��:��Q�����'����IƺA�a�������1j7�<����64�&��~����Ԑ�̙��R�
��1�Î�s� ����`��B�	;:R��TO�x-�V���_�7��"M��Do�ʟ��I�����+���?���@<�z6�ך~���J2#_�_�a�'�x��!.��)�$���	l�8�p�l�$�Oz���N�&���	ߟd��)���ucR�d�Z�I!�V6H�Bh��؟T��۟0�1	���t�f˷>��3�gB�M���Thi��?�CT?��w�I��X\��F�D�`� �۽:)���O"��][g.�@"N�W�l�OBL�a��Tq�y�ᅩ	?l��'�~0jk67�28�'@���[��dI�g�uC�(�1{	��J!`ٵ<�Vd�6�ֱ\3l�jU��l}6m0p�T>� �kt@��@���h��p+[dUA��ݧpkܘ����X��q��[��-���Yc��q k_��Ja1"��,���WJ��d�ҽB�/�->��`��
�C���n�)Â� р��,����Dr3�̈�̈����ipoڞ
8="'�'���'�Qcf^8bLL���%?�|���WE���׋*C"�� ҿ%���T�A�'d�Y"�%b%�Ӧ��d�	P�B��-��Po��l��1R��; c��P'm�E�'�p]����?���d��>	�B��׉f���q&/���y��'��"�,�l�S��B�gD�;� �'� t#"l�0Ft���c�7����'�Xȑ3D�>�����\�D�P���O��$�0p���HƢ�,uwc��"NRIz�H�n���qn�G^� ��|����O�����b�nE�����m��T�D&A� �5"�>h �Y�𧈟�	 zl��1 �+������ ����'3"����F�O���Q!&u٪l��aѠ5�l�XR"O��Y�$�2Z��Y��Vp�i��I��HO�>y��c��q��%����8���I�����@ ���	۟���͟0�]w���'n��r����D�ѻ�B�MM����Oxu뇨��{��t���U'�������h=��E��'�R")׺H��4�I>o��� 1��8�������$UgP�%8a�X7E�v\PV�M�%���	C���'[ўt�'~ 
d��Z��#�߹���`�?D��b�⊽Gi
$�����(��]*����HO�DyB��~�X7M�6}b,�qK��k�F�C�O��D�OZ�d�Op�Hm�OT��y>�cW,Z����Pӻ:��be�� ��d"�LB�6��9� / xx�$[�k���$�ˁ��O2E0t���|\T�ck��X��M���]x�H�ck�O��$ƟzK<�&�#F|��4%�,{ �=��D�m� E0�	�c�\����@� �!��< ����+Ȍc��S�#��'��d�d}_���5Nɬ����Ot˧u1�p��<�>	�ucO�w�&}Y�#��?	���?��^bT���r��-4�􁡵�b��S�C���s#��5�Bp��T�+簢<!@H��u�dB a�/8���$�~���CPc8�Phɛ$z���UH�'�V���Fb���0���9@�O�#p����q`S'w��	Ɵ������qxPc�#tm␰�f�	AC���d[J�I|*��P�
R8 ߪ�P��`����1M�|��ڴ�?����)�1U���O��d!0�D%"���?reQe�D��1���;+
}c�9?�O�1�2�γfh݂�%R'�,�k� ױo�z�u&Z�;(b}뢙�"~�	�>�H�P��4N�*��(Xv���'���H۴}䛖�'�?�D�.*"�Q 6���NnB�����;���O���W1;؍�qM+)VljT�T�rn�l��V8cnr�$-x����HK�^��8Qr�Z=I��d�O�qqSY�����O(��O�<�O���X a��EJQ�,YNv@3&���d��#�z�+"I4��!���n�ذ��+,h�l�sd4.n���C�)��]�G+�
 #��r�?�=�tX&KS��y�Nگ>���Z��J��?�$�	��?!�iUV6ݟ�̟��'�2x���*B�����$��YX
�'��`xR$)����LL�	-|Lj�D3ғVe�IlyR����=� l`� ����iRƊ�8�@y��O����O����{�b���O��S�aF��Oz�r5ކ}T:��G*Ck���;5�'n�k)O�́�b�3AV)	)9f{��"T�'����?���@��kFǘ5N�	#�a����?1�������8ax�x�v��	GΘy)C�=(!�$Sw�"hp��E��07gNd���]y}2[�|ʰ/9��D�O�ʧ@A�4��,�18�;bHC?+d����U��?i���?���[=O����/Y8 Ro�#��0uD�Yv�ڕ,�>-�qM�zQ�����!�8e�ԏ,����B�?	ҡBO�7N� ;t(�DN�M1� ʓ0� h�I�M#��	�����K !ն*�^���KZ�$�OZ��$H� �� ����*��Ȃѫ�G�a|"�)�D݁N�x��M�z���L�'	��'��Q�'��\>	���Tݟ���,��nD2�0�A �1
(�W�ՆY���!2�5k��"�D�	�?�O81�2��, 4�e��i-
��+��LCq{���	�F|�1ǉ.E!����O�99����E�C +Ɏ4�aYr���$���,O�O ��U�� �%��/�z���Jns#�/D���b��^�)��ο{`~�s�g(�I��X���$������%t,TX ch��2F�4��.#Vm^,��˟��s�K�r �I�����ɟ�������A�\h�&@�~F�l:�!IL,�d
f�<��Iui4 S<�8�sK��E]L�	r�&Lq
�7VΘ�LX�6aҪK�!�
�z�S������?��S�'x�V��p�f��I�9�A�T;�Ҝ��g D��[�F�5x�(c��%'���3�B�HO��n~��}��f�ͫO�N����lw�!�A�S��'�r�'��U2��'��<�6���'�)H�r�:xPqk�wH�1cV��5�p>15
Thy��
J3����G18_t��+�#�p>)�����3�xU�`�Ȅ̰���[��C�0{�$ep ֔=���Y����4�pC�I./�F�PKA�,��h"ą�(\#��I���'φ57�f���D�O�˧tQ*��ddN�zY)� ��(x(�HM�
�?����?	�c�V�,�b
�8ոٱ2Ƃ��(th��a a߿swT��D�*0�<�R��1t�pP#Ö�D��׫����T$8h���)�F-0Z̄Ey�AL��?Y����ڨ0s��izh%��@�a&!�à6����ѵDwt����A6p�a|R:�dI�t��D��6\�\ ��۰T�1O���K�%��BT(��^T"s���>Q�!�䃃y������J�\��`�	��!�D�D���ؐ��$M�zP�Ԉ� o!���9����Ee�Tֈ��(��B!���:��pP�F��*���S!G!����0<�IU�ړ8�$[��6]!��0V��B���6�dE B��!�D�6 㺀qSʙ0/�ơ��G�!�Ą�4K��ӂMGu
�K$A_�2�!�dI�~h�J�ǝ� �r\1q�ݯL�!�D�W4:��`!�)(ơ���!��P2}fq�"�vhq��!�d��~Qб8�L�$�5�'M�T�!�H�N]�D��2�5��'5!�G��pqS�m5 ׎HB�	x!�dƊ7�����
Ia@�Y��li!�9r{ YB���(Q8��%D�Q�!���g���K/U�����K!�DԟwM�H�&�ՄIM�eBd���&�!�d�V���1@�Rx�bcX�{�!��^b �`��B�lXc��)Is!��QwDm`��&����"k� qb!�D's��ai�k؇P�F�yf�`!��{� b/E%{E�H;#h¥8q!�$�H�hYj��)�~q���me!�(p���f�ػ��`PAfB^U!�*D�pz!�>1L|�s�J<X^!���7���!F���r՘'/�[U!��OJ���kƄt�8�"��	Q<!�� ���DA�A���h���Ls"O�6�G�6bf�OF/5fx�'"O���C*#|ެ����U)@�I�"O�e�tWt*)�����lHsQ"O �ɴ
ӎjByX�n�!?�9�"O��b��3m�@�wn�"k�<#E�'�̵	ϙ-
���'R�Q�R	s����� \�l)h��
�'X���넏DĄږM�Y�d��O���%�^3|��0��Fś��X�N�H7�إIYv�ȓ�>ԓ�*�"]�i&E<uX0y��S������rZ�Q�'Ҵ�Q��c�
��\���d�>w�FII��X<a����N]�4 ��(a�̏}ˎ���o3�����
�?ٱ� �A ^|�0���4�
%)�4<�F�;J�n�J4�:O(H���P~_�PPq��<Ʌ�ޝ`�$*�_;zk�A7攜<Hh�
�HY�r�~���
!��<i��V&]q=��
�03���GW~��
O�v�Y`͟0n�Ɏ6h��ڷf�%_�85�r'�<&g�=�v`�&p[%$zӾ̄ƓeB���Q�׉dhjTP��"l���DL�qm�5�k��I����s��OD��
E!?y��@ܘ���
0�(����-v!���S�бC$.��f�\�Rv�����h�+d�BYk��]�\�DϺ&8���&��&l\�g~�Q��&)���د{2�H��N �0<i2A�fG~ܑEL�6r �B� ӧx�,��vK�AS��8P�_�C��Ê�PX2)Q�cu~4;
�[��!(�Wb-
��,B�"��'���X�LDzccD�R�R�%i�����L�v�P@�^�: 8��X#CD <�LݽfH��f��A��jA k��h�@ �PI0c���j/���)D�1
��	#Iz@��f�i�D ���nN�Y�rd� ����֧Ջm�!�d^�`���$1p��=�S<qDN���eԾQr�O�3p�<�A�ܼ^����,0=�< �#�d��I�mK�j�)}&� ��
�X�ax�eK�S�M�7�}��İ0�и`��E��*ܤ���׷p�"�U"�;L���'�T9O�|��'֒�e��%��x�G��3� Ȁ�Ov��2�>� ��J�4|�7l�<+���,h�H�
c}���G���j�;���*��䂅Y�>8��b��6@�e�D�Y�>Y��ⓓz��+wU�U���sӾ�d�@�a�U��Լ6T�C���dLY	�Y�F��Im�0��
�s��+ ��z~��S�q�┡UJ�S?�O�5�׎G]�a����A��=�B��,g� 7��x�Pt��D��{I�}����c`ax���d��	F��~$�]�=6^�+ ��X��tzF!V$u�x���딚F�j!��Y�'�bDPc�'�^�)$�7�i>9[�3��[�aZ�_c̔{4N+?��Ӕv7ֹk�`�6'k�U�fk��?� m����Ė$b���C�3B� 8p'@��zFl�Ȣ8,��>E�����E���C��J2�,�slT0YY@@�4^�����O��-�wdD+�y�eR+&�|��1�Cq�����8��d�?���ɷ	-�M��D�r�V�P���"�&���c'�+=�m�kJ�d�t���
�"/���ݤZ���oZ�Wv�(äL�&V�Q�vK�	����UX�0@��9�$��=v���i�i�COP�*��?R%Y����V�I3�ՎB��!8��'�+ea=�i>U��L�^��=��I�{m�4a��9�j���b1�u���f�8���M(.[��(���2C��V�հg���/p�є-N�>�j4 T@W)y ��;Y���w�V#�t䓖�o�p�)§"��D�� \�{�\�A��-+��	��CL�ÑM�?=.~�+%F
����'�\�jSB�4N��y�Hχ7�AsW��3����c��1��>�g��Y�}z�뛮=��� �!K�1
�T8�-<�yBi��f>�hR5ɍ�(����q� �HO h�0�F_�4�|�[9�����)ђI�1F�Dn�<!�͗US$8����?��T�����b�$W�%�"~n�Y��`��_��*RMU��B�I	A�LM�-Q''��T��JR���(	:8K�����p=1pk��^V^�{E]/<������xX���-S1�n6M��	�Lq�
�	����C���!��%<�P$~���8C#
(]đ�� ��I�>}��,D�x!�v�J�8�c�6D��!��3!:,xX"(N�	��TA���O�1��2�O���5	
xyb�
`9�X�6�c�̫ dJ+-�!�̈0Gh�	��noJ��$J!`y�I �~B[�h���O~qyW����I�C���;��4m�p�dΘ�0?1cD��?�'�	_�`a0�Y|( �#�	��r��'�8��G	�<A���O[h�#��v�X�b�af~	��i�h�+7�	�y
� (Y�@'��H{b���"/-d��ض���L�"����'�桳�g1F�X0q0��{�Xb�'�Va��x��4��Ƅ�R��q�韾*������;�8H�v��]��c�܍l�r��	�'E�ّ�d�lV8��˄gr�9�4{Ґ-a��i��r%͈�=e^5��G�a�y��gO���N`��g�s�(�iP�]$L9C�'���#t�'(@q���S4#y�lp쉟r]���od,eqo�EO��kS�.��)��|�6:�x���L���AeA!�^��Ҫ���OR�;�A!}R&[�V^�6��@c�탶d�8^�m�5J[;���J���<lC!�c��^���A�'�m*@A�*0BB��Z�d�ѝ'�ā �>٧��%��J�N��ū;sda�6�DA�Fe�T����}�&�W�VH<9@hN���1���#>�n�j�]����j���M�p���_��X���=J�r���J���5Y�\b�;E������`E��0?!S����?�'�D�B��X�#��	C��{:^h�� �!�Ψs�� GP@�O`-	�F�1��<�b@(g�Z�%,*��X�&f��D|�ON,He�"���i�0�Q� �#�x��blIe=>M"A� |p"�F*Ά�V�Ҷ��<i�J�l�bW�,�qqao�A��$˖�e�>0�M
ț���; H�b��,�v���%�b)�Э�Uh|�蜨L�B�
�'2��J���b��Fa\k"Ԕk�4鴰b��ic�pZ�
1�J�&+�4�"���Ne��Ƥ ���l_�t!���+�8,���'����$}˞�i4�X3�,d����G�1A0�؞Bۜ!%�S���a:D@ K��SV*,e���;�D�3TG���A�ԫ	��S��S�JL��s�☓9���x��'J�qR�y�@<!Sm�~V�25�8�����̍6�F��a�-W����Q�X�[�ay��U?l�&x��bA0B�n�I�mВ�?�bc���!����,���EߟX�Db@2F�~�	mѐn�HՃ6!N����!��=�D��E���B�9P�)�aE��|}����?a�7%��DÂk^L�t/]9w� `ÛGq$�f�I�����^HC�"�0#Q�ِ6��f�|d���'M&��&��+)X��T� >\@��/Ոv4te�T�	��-�CŻ
sB�*�KV�J}z��P�O�@��'Ũ��X\�B��
�Y�
}�1,ՎW�d,Ez"k"l.F��GЌ �b׋�ybbU�ܥ��U9k0�7	A0q�\�e�J��1�ۄ	�bX��P�*�*ᚑ�J6?�xM�O�pKĩ�Y)��c��'PT�R��'�:���K27�98�M��"Q.� ���`�ɞ&��h�	"��xO �S�LF�,^�z&�!�M��� =
����Z�TG4b 	�:&
,�'h��|
�D�#��1)�x`hfl�0(���P��"b��?����Q@^�/Z�����O9��9'��Fa*����^W<�Y���,iD�����_X��1E��S�	�@��Y9"j��6��� �@�#<!`�Jl�vL�2K�<"��h}�b
�>lԋW�"�ޥ�2�9+�!���G�|�pAj�\((���	˓��M�pM� �SF���Q]��XD'�NW$	R�O�%��(�m_n}�I��{��	c�N��*sb��m��kQ�4��$���ֹ;1_� <����HLC�h��l����=���e�b�`�E�;kI@��u`�">\�A�'��y�*�G3У��29P��&���`(�i��㊣>8``�K8/4����=�O�x�%'�Xg�Y��-�A`����  y��mrF_�%���X���L��!�3��G���[.O"=�@�3���nX�44�� �8**:0;�k��M&��U.�g�':�D��	�4�DU"��kM��'��7�|�d�BpI�+T��U�1+����|�+O@�R�ƮV
 �r	:]� |Rf�Ĕ7�>�I��R�&E� K�L}L�s��R� W�i1aC�I2����?O>���I��mХ��:���	W��%7De����/NP9C�G\�-�\�CU�Nbآ4 4lO���EH=/.`� S�fl�j&(��IQ��mڧ�~b�V�"
��,5��X:ua;Gb-��5v��[}J�i��P�6��IǶ�8��Dm�kJ�8����C<BK�A��F�u�ʨ#ԁ��@���a0��$�~�S����(O��iM�rjT" "� 1x,��߅���;`吒G�$���s�'��x�D̝O�$�1���e$��sӀ�m��%����Ê�F������O(X�~�YVQ��B�4;�pM��fX�9$v��0��*qU���W�gW��ҠL�]fX�S�;�xzrm�MJ�m�a�u���9��|�&K�0-d�!%J]�?ƈh!QJI�	I�U�r�L$����匉�����^-O���d�H�=zbd�7� ]�w�]�*)�Ȃ0���<1��~��E�j�L�:�d�S?0|��䬟��LՈ�bz(��"�L�;*`a1�'�j�S5�a�2T!���'�^��@�Z����o��d�� 9��J��d	`��	!~�KR��c0N��S�D���Pbg�� �!{6��i�$@�l����ח�OT���k�]���6
Y0f &���<��HM	EHP�+�ϹfW���g,�(}�ԕR������)�	�8N"��GI\+�@�i���[�X��\��BЯ(&�͋ �ψ����%��K���fjΜH0��*��'��,3�O�RQ��ʐ:\�<��J���`��O��Q�揍?C��
0S��M��V����G� ���#g�>w��)r��v�b?Ak��W�`��3��R�����*D��%@M�/��q١���HI��X��U�����?�$杴d���T��M>�w�@�� }��E�����#�\��$�+>�
�b��D��Q4��ai����`V�C�f��
�����<� TX)R�	�N=B!v�B#6>���I�g�:�
�l�K�I�T�^<U֊�7��N߈�B��V{d����f!�M�YD�A-6C�u���U!4�!�$Y�6��vnƅ+(t(`l4`w!�d̑�j�I�k�;%����&|!�$��Wa�A�VO�|Pa �Vq!�䊭a�U��(�-2h �V�P�bY!�$��� ���NT2���i[Fo!�D]'F��Q�YG��1؄8W!�$Iڬh�D��;T�xd��� %2�!�T�e��:�NL�@�L�A�R109!�$M�H�tMr�iÿF0�ѣ�տY8!�DćPOf�R,R�b|���.��$X!�@�it����4�^�Qg.k�!�d��de��Z�l�{��i:��:�!�HW�}b�-�T�����o�_�!�AJ�q����6i5+G��?W!��� �ni��/�,6���nK!��#+� 8�D�;l*tL�+ԣY.!�X�z%�I��/�@�|SD�T*�!�V�v��]�&m�"���|�!��8���@�${�(;�KQ�T�!�D_�7�4 #�a.Ĺ��.&�!��N�,�j0��ͩU�N�y`A͍^�!��ȱQj�"��"?,��k�x�!���B@�U/h�QB�GW"!�$B�}�TLB�eS�Y�BA�]�E�!�D��B:h�2���zH��mD	!�d@"Z|�9�2��|���,��!�P6~MV��(��/r�(sbl�s�!�J�vQ��ҀŁ�<YdMZ�@J"8!��H���)��'�� O� ��!�䇡O�	�`P�h/�)NQ$u�!���&N�8!�f�W�*'���4b�{�!�ͿIʜ<�� g	 ���U�" +�''<���A[���P���<��'�<,zd��[TT�;��Z�{�4u0�'�H�20�βZ��$sw�$!��Q��'h���cG ]��A`��b ̰��'��i�d��r�Y��Ȇ�,�x���'���"W��W�%qgǗ� |	��'��@�!�?��K�H�D`�4!
�'�X�����>�L�h7j^$R���	�'!*Il.jXV���,�mu��		�'��x#tIM�1+?8>�;�'�d��/�l���;�K@�1,p��'cx�!BE����Y��TX���'�~��f�*-�H�$��4Q8�I��'�~�Wᑈ~�ؽ�F�6L�K�'"ZŢ ��wFik�
�>�$�����!K��	f�+�@0Q7���<Y�O̭:W�u�L�EW� ��g�<��A�I���H���7rx��3iz�<i��N�$\|ŀ��R�Y��!���x�<���7x��ido�t�l��'�n�<�'���!���#�F���gMi�<�7*��@Ȃ�"]=�l�E�l�<AD�\�D�j�����6;��c�F�e�<I5�Ft���W�U|����K�<����B���
#��3�]'�o�<�P�"U-�s���)(8�����j�<ѱ'Q�tn&�aA�>sf�P"G�e�<	r�Xx�L|X�(��_��E�b��_�<١���v�5X�U�k�^�<� J\هDw ��#b��)���X�"O(��K=si�D�t,�^�T���"O�����J!c��g���ZE"Oح�g�/=@ �A�U�D|����"O�ب�R%f�2�gJ��r� �"OY�$�͝n�0�Ce��b��T)r"O@|Aa�/(J��H�-��0�(���"OV���Z�M_|��R+�g�>���"O.����ȕX���k�	J��<E{�"O��A�G���M��(��=��ړ"O��(�냄:�ЈHP��ʼ-�G"O�H�/���J�x�Oڈɲ�z�"O�� �AG�����2D�a��"O4��ᜧ@���f�;���"ON�0d�]|a��lB
	���"O���RNO2�2u�F���业"O��y4gȾB�Rd��}�A8�"Oʐs�M�a�6�"�Ci��� "O��Wɛ�M���CCX�`���"Ol�W-�"Y18(�@A+-��R�"ONMc���4"�,jc��cĨ���"O�*a���$����C��[↩;$"O|����a�@\94I?W~��S"O�\��F��2i��:#�fc"ea�"O�U�6AH*11e13�޵FX�,�C"O��e�"uߢ(���2r>^X�$"OH��GA�_�`��aW��n(� "OrM��.kk ڕ�Fb�|�j�"Ol<� g��i�H��@�U�Xta"O�eؗKX,��񐁁�N"�&�X����¯��ª�ha��QbB�Z�N�y�/��fB��{�G[�Y1�تe�@�y���vŚ� �.&Z�u"B ��>Y���y�ٌ_.����$m(�R� ��y2f��Q����!`
>$S�텨���hO����{%�5�@0W U�}~м��"O&(H�ㅑg�p���ȸ_j֬2�iR�"=E��4��uɅ�)T���	(ڐ�ȓ[V����1�t����Y�H�ȓJ�,L�t�]>�:Y	s�\&E_�y�ȓ[uz�rj$j�ɡ%`Z�(��A�ȓnӼ}R�˅�Ff�Ճ�{��|��f��ĺs�R�"`0S��-n� (���T�"��1H> ��V'm����	J<1���5QJ PR�J��,=��/�I�<d�K���	��TmZ�)Q�_�<�F�kאհ0mOd|ht�ǬE�<1p��#Iܡ c��V�"�� F�J�<9�K�M2�� ͘3
p��O�<y���$�c!��@؂�0GN�<ac�X6F��i�hQ�W���h��Q�<�QBԉc'�A�N�>�x����EN�<a�b�2�T�   D M�*�K�<�4GӒ@�"��<�2����JD�<i��`E�TrS(6Y�9�&Ɠ�dD{����2�H�P��E%X	�}Fl�<i,bB�E�^����4w�L3W�4T@B䉚3�&|SK��a.�)l�$gf��d;�2}=
9��dV�/��zŵ9wrC䉣��qv��9?|\��T#ˁUg�B�I�DV�sp	Q�g��{�C\h�B�	(`tN���偽Z9>�Ae�,GfB�	�	C�9*��	�?l��.S�@uBB�	(�z=2�-��y�ޤ�#�15�B�)� X�VL�$`hb�m�x�ɇ"O�q����fH�x�߾
�>)!�"O y�'�ؠv���b�۪J��L��"OT1��t&�P� ��O�HD�"O�!(w��*�M��ΪOj�L�"O,�#�L���ҨًlNv�0�"O�5K� ��-8���^� %"O��R��1Q�ps!/F�8`�8��"O�@S`�
� ����G��-I�m��"OX�xvD�Xf 0���V�0�ح	T"ON�K�fU�U$ht�*H�5�	"��'��$I54��7ɼ#�`aRc'ʯ_t!��P�N.�ء���x�^�0l��yX!򤖻�0��3\^6�`21�!x�!�d]��\ ��͛�_�|�ðI
v�!��
j(�K���aCG���P!����֡(�JD#�Vl��g�y�!��Z1��*���N�p9��%�� [!򤜬6:�Xr��Ž(�~�B���
q=!��WL���%&ڧ:��a"��V��Py��CP�`����Õhq��`��Y=�yrJR:*F��pAL�V�jprS���y��%$�A��k
�<�\ѓ�� �yB�\�9"E��%؛��P���y��ъ=h�����"���7�0�yB	�{�DX��+	u�RG��yҫ�	
��S��w���aq���y���t�"�@F��A-jY1F
�y q ��ECE�b��� ��M���	V���O^�|Cv�>3�:����ߺkL.�i�'z��֣��'�Υ���7_�0�
�'��!���&	�ԡ�@�Y>����'���d��l��j�L�<M�����'������F�y���<G����'���yW���/��"B��̸ ��'AY���-t(����V��$R�'3�ej���_�:��ČD�U:�K�'B I١�O�cJ���ҡ�W�`�"���8����NZ�>�6\``D̤��h1"O~]����w�˅��w��PQ�"O0�"�IÒ���:%��/��``"O$�*3��m�P����ȓj��u"O�Tp�Q�&l����,U�;���v"O�8�­�/c�X���AO�w��9�2"Of ��B��C�n��ӆ6�h��7"O$���f�ԤHunT+g�L�["OUTl�j���� M�q�v!�"Ohש�!F�� 6 ڑx�"O���sG��Y�`��D.v��#�"O���最$�|�ȦG�t����"OXf��0{o��1T��:�k�"O�a�g��%�6�pF�(Q8��"O^y�"C�&kC�\b4�ć��"W"Op����<!�"�u��M�@"OB�zuÑ3�8��゗	����"OL���@H-C�Zd�V^"�K#"O�)"Bf�>�(-��BP�*�a2�"O X����82��!��kg"O�X��@o/`yJ��5|g��A"Or�k�M��8�0�J$�q*�"Oh"��P�_Gd�AAK<]��1:3��8��	�es�U���7Ga@��*N?1�NB䉯ApU�v��e�z�ڣoN�7"0B�I�-���B�	)QlԺb��$nC�)� �\u /��}D��??��q;�"Otɤ��)S-
p��ѵ��Di�"OʔH㤛�U���!1�2���*OD=
c'YP��j�ʷ_q
�'z�a ۙv�I�c��[	��@	�'�y�ӪV��3�ν&�P�X�'��[��I<y8�j�hA=���'<t|��FN��$Er��)"��� �'��c��'�~����IC��T�<Y)�J�������4_�Tu����b�<)��Y%!FRp��ʔ�6���ɏf�<)�Є ~ ���(�ԁY�<ɕ� (X^v|R�'��[�8�!� ~�<!��.�XكO�v�6���x�<�0�
6��	���J�4�CAQp�<���� *�@ �1OK9i/�貧�v�<a#G�56�x�ȍ25�v�
�B�n�<FK�8.��)ub�3�����
LP�<�e������V/%'����j�b�<)���h�fWJS/�x�D
�]�<�T�U9A�
���M�N���+���b�<JK�#�ԙx�΄����8��UV�<�ʋ6����T�((�x��2@h�<!���mMp�J!�C�3� �$�l�<!b�ک7W�t���%"`T�5 �a�<A3�%g ٠1�
���R��a�<� ��,ۼ�1�K�!-��i���[�<YcS�=T�a	�-��Y��	p�<�4�E�;Y�Q� ���R���Aէ�u�<�`GZ�T�L4�R�4=�
�ea�s�<���	��ֽ�'���U\A�Yn�<��h�,��i��2m���l�<Q.�$<�y:AmD>��-ZP��e�<�I>N�NxC0+�(M�	z��y�<	�c٭�T4�qf�Y��L�ԣ@\�<���!x�� �GjXFEre@XY�<�DK�6��UB�ԓq���HY�<q���J|��%�H�4��Ĺ5��S�<y�%!M�y��Nӄ:�0d�C�Y�<qq�Ԕ(������?�xIQ�MW�<1SoP7-FV��aM?}����AG{�<Y��9$*R���=-����b@{�<��H���9 T���*�k�<	� j�M �O�o�=����_�<�e�R�D傸XЃ
ABb�K�"�T�<��F��C(Q���
=na�$K1.�R�<���=Xr�H�4}6`}�q�H�<�P�U��(ATL�0u�0#�Y�<Q2-U�cJ����-�.~)s4��Q�<��$'h��s%�<Ğ�Z5�^f�<q1fF�~E����Ś�J����GH]h�<T��!1�D�b��K�N���4��n�<	G ��>$gN��.�j׉�m�<1c��$e@�9Q'�	� ��s�<A'-�/�Z�#�_ƸZ҈�r�<����&U�1��E�>i�PHQI�<9��~v9c'�[78P�<��fLp�<�̚,�r��/ݵr��Y壃p�<av�Q�
����CK�W�R<J5��m�<Y �[�o����A)2�d�1ħ�f�<ᠤP��0��IȤ~�����e�a�<Y��\�J�"�� �*L٨�����[�<i`χ�O���sW�$\����1�CZ�<I"źi�ZԐ�gG�r�H�J�<� D����"�.�)R!	#B�`1P�"O̸����3���`���-eɚ�7"O0�
5"��00�⃩[�8�;E"O�5C�Ő�"�A�g:qW!3F"O(�2�c	>���`ԼL��h&"O"�
+�=!U�E�@"S� 2�D2"O�R`�V07
��ȅk (o"�x�"O>�в(��G�}0"離- R`0"O~l)"��e���8�WOZ䊑"ODU��e؟���"��NKJ�C"O^9ȰoD2W�f0;�BX�A]�9�7"O�f�Z�;ش���Х&Gܕh�"Ohd!)�=6�	��nqV�y��"O4(B�!�<^M���@S�"U�4K�"Ox���B�u���2�, �xP �r�"O�ks<��5H�F�P�5Y�"Op;VD�<:�8�`׀'A���"O����R�e	�<S�6J�}i�"Of�b�K�0h�ޙ�U�͙zG@L;""O:����J <���G6nG�2�"O8r�e�)	�8��CV:=Lqr7"O�,�SK�4Q�!�LR'W$�i��"O�4�ߟ?��@3@�[~\�"O�8x����Qi��I�	dظ��"O�e��_?&�B��!�J�V0�f"O���%2�2=( �� �
�d"O*1Y�S�}�h��aJ��(I�"O�X��NHT"X�F�$h���"O6��D��{О�)e�i.>Ԫ"Ol�S���]օʷC��u�H�4"O���#�H
j[�i�rȆ�Z�C"OH�s坵+c��EgM�	B�8�"O���,�@�>��Q�@9m<LH�3"OR�s��u��Jd�?��"E"OnDcs䝱{1�upG�+3h�K "Ol�jpn޲��@#�K�[>AZ2"O	��W�;�D)���R��QY""O�u�!fK�X{�(��@
�Q����q"Orؘ��X(3 �C����"O(�3���?T-��RIZ!w*Z�"O((oL;��0R�HH����QS"O ��D�@</H�Cg��`��}�"O��CEҜWj�)r��Y��d[%"O�ܨ1

#^\5����Wed{D"OZL��	Tn@�yWJF1J~q�U"OJ}�@ o�,;�)9q+<Dq�"O2�kYm�VA�.E�ܫG��d�!��D7 � i�#/���͉�-B!򄏡�l<�e^�n�� ̖	=!�%^*���%!�o�}Ѓ�ǀ�!���`<�p�ƪ��}�p��	�?7i!�D[9j�Lq��
3 ��1-�!�D���#t�3l�>Y)"��.<z!�źX����,�z�t؀ǟ�i !�J�g���Ü6ܢ����\��!�D���a\�1:ȁ�U��.�!�D�DZ�N/4#�<���҂/�!���+�>	�B&"g���rڮd�!�Ĝ%U���qr��>�I���δ^!�Ē�`��9���H�"�� �79!��BN��$�Ō�
s�괹��!��F)k�yA��-'
�8�'	�y�!�D� D(�UJ-;�r�Jd(�4-�!�՜I�0���P"씱8�˄|�!�� ��iA�ٙNCVp�FP5_|l�8�"O
��W��H����4#@�`�3"O�� ��� .ɾ�0��+]'Ya�"O��;ס���D\�n�m{V�a�"OR��U���
�:m�-C
	��"O�� �C7-���G��{�6���"O�h@$�Zy��1�l�&�fq� "Ox�r�+YjB� �H�d��|""O Q+"V2f$a��@-a����"O&�5��sL��,]!p� �R"Ox�XDIV^U�E%�n �"O���(O�#����}���J"O���QB�7��lz��
%����D"O šq��(����AX6Iy����"O��'�J��a�� ^v�<�3�"O0jr��
������#�R���"ODPF��>O���o�&5zDܺ"O� `�K�&<ȡ�s�G��:�HW"O�A�b�=q�\D�Ň8��0��"OZ,ɑNޏu=�<�瑳"o�`�"Od�[T��8Q���r�e[B�)""O`t�����0�K�kSPL��"O���숧F��pz$k !S�N�С"O��:A�[�i"�A��@\m1��0*On�r�ME킽 p��4�$�	�'�P	�nDU�<��6L�a��	�'.& ��Q A�ɋ
4V@`�'&}�fK��՜a�6\�����'�z��㑶~[�(Zs�0�K�'����⭉/R��[�`вd�X<��'��ª��R�岴��&WT���':0����?��ꖯ.P℈�'f�q�7"lX;V��7�l��'IFPq& F���<8a�+�, *�'kЈ5Y)��P��r�����'$��(�/I�a"���ƫ,_�`	�'�`��b��]�����
!A�T��'��QD�.Gg�)���� MV���'�X�T���I���# �xɒA��o�<�>)G䰻�J�R��"� �j�<9&���,�l��d�MF��Q�oE{�<QPpf�9 ��Bi�a�<ф��� @�����>�j@�v˞s�<�J
w  \x��b����v%q�<�b��  �3CJ��BDol�<y�f���4�S�HRT����m�j�<	�瞲!Ҫ�*LR�T���f�i�<����-z��ɒ$�G!X�.u�4cPd�<��_��L�KR��(�8���^�<)��%	� ����p��`r�M�]�<I"��#�y4@�>s
�m�� o�<Q��J��4IҺ/4Й(c-Vt�<	��71�ؐ$��h��i�S�\q�<��Q �$�Rp[�Fv1 �c�i�<��k�j�h��c� E:Reg�<A%�Y�pi"(��fQ�PP E�K�<�0*2T���d�v�D��@
�b�<����FFK�U�;!l�
���^�<QU�K?S}F��%T��Q)&D�<���&z���V	�1�����h�<��e ^�ܜ���ѡfY���7"O̓��+�5�rS�N��z�"O4�����	n�x�D�B (B�t8�"ON��㎶��ɹ0!R�656�H�"O� �sf$#���Au�ҁ'p��D"O�){�G�.��{��;!�!�0"O��aP��T���0aE�<r"��"O*=����Kj�Z�C�P����"Ob�@�%PN�`�`��NW���"O:<;�� &[�pT��A*H2��e"O��p�.ΰ~Jp��G�[+бiP"O���mK�?F|�k��ԇ{�HA"O.8#� ��bQ��B�K	cX<�"O�yY1��;_�H4�#J�+|��p�"O��X�.O�AK�m!��0E����'G&@{.��X�`���4�l���'g"�I¤Sj��|ˢ�і+���ʓ<Yp�S��2�f�1r蝚T�Ru��652@�a��byވq�ܘoΜ��ȓ�p��7^m�ޡ�A��(�*�"O�8�G��*:��0��:B` "OD`J�,����2�`Q#N4r"OH`:�O���,�h�iބc��"O���cPjptHΡh��m�p"O	�Ӫ�eOL9�b��- ��X��"ONm(0EP�jj���e�0���;p"O�=��� Q @I��M�6K%"O�2G��(h��A�7/}DT)�"O�-�A'@P �S�Ϛdy��9�"O:)���G��q2�2�@�`�'4��" o@�@|D��e
m�
�'l�P'�	"!�F���V��	�'<���"*E'[�hp��ゾTxVA��'K汢ק	�9vx���� N�H��	�'Ӵ<�G�	w�ЈS�I�t�B�'"4��iٿ}�HIq!o�Q��%��'�:A;QeW<Zi\�I ؝N����'и3"+�(�I!�*�)����'(�Bfʄ�*6�@ke����'�f�!a�ö&lA�fއ~vT\k�'�6�*&ڔwI,���ĺ���'S��;��нb�js.J�7�!��'T �0��P> zjX�ۭ|
���'$�б��	~�@�:��ǭr;�8��'y�����J�b9�G\�`���'Z�����B?L�☚�*��N�,m��'�H�*AA.o��A��j�M��1�'2���f��4,�:3�;J(�+�',�YAp`�;%g��Rr��B�� `�'��\��K�Z5<����6r�Q�'���̈́�l�x��V�X���K�';��Hr�_"S6��pӂծ^C�z�'����E��>#�0�q�.��q�'�Q�CCݰ(b^�
R��-*�H2�'����@(	���C6��S�5��'�MCn[�Y?(���kǘ��
�'2�ö&?@��$i�(Zi�ъ
�'�n؛Sb�����G�73�F�	�'�tc�]�ot)�7�]��-��'1��ӓ���i��胆�қ_C~xY�'�nѪ�"��h����E�C;0�
�'���
!S�����V/=7����'�D��7�~�ҕ�'�#2�4�p�'Lt�s�&��Cd`���'Wh�q�'�l�;��#5Ǌ�1!��T����'���C��4_�,��DµJ'f5��'	<A.�$mG_�x�DX�'j�i�d�_K�����ާ��	���� ��r``�$K�ؘS��I���@$"O0���@�� �ds�c�7��p�"O4
���=R��'A?u����"O��R���<R(Հذ+���h%"Ol|�-;.���O�2�����"OLX�Q	�S��C<p"��t"O,9�,C5I��@a�+�ZL��"O��
1fM7R�dS#,_�P���"O^l���K0A�PjD+T�?Ҥe��^�xE{��I^%�:-�#�\?C�^����ƻ7!�$��N�0����C��U( ��"m�!�dF�a�,Z��D<1)^��-�!�$
�.n���T�h��sjʽ'!��"2K��b�Իwt�U�E*ɫ*!�DX������4`V~x�%����'�����Ɛ8�\ S��H6�|RH>y���)�	�t��]Z��G ?9���D�;L�LB�I,{"�D����Gаq�0�R-j%�B�I�Z�Blk���%@�@]X ���i��B䉧|���qƀ�a|�QWC΋_[�B䉴"W����#�L9AS��ǐB���ީ!�.R�,A,��/��w*R�`F{J?�Q�N-��(s��]�#�^Yx���<���?q���?����l�����V PJ�B�H%;�!�'A�Αs�F�S=����^�5t!��l� ���5{�`x��(Ğ�!��'y
, �D��=��E@
n!��ӑx�~i�fK�2M�09��EM35!�^h�T��Gy�	s��!�d+�:Y#S��?s���
�@��!��9�>�2C�A�sPԫ��J"�!�$�!��؂�C7 =��SՌY�B�!�Ğ�F�`:��  �m�gč<�!��E�=0��Z��ԍ��wkQ��!򤗕f���h��znX�۲J�	O!�Q?J�,ذ��(_aH��R)G41!�$��b%�}i�D�z�i�-�?:R!�$�5
ūj�&�=S��5_���ȓ����o�b�f3`��\0���l���ʻcP4��rI{��$��n5|�vj�00�8����9H����(�(ā2ČX@\�0��x݅ȓJp�Q�F�&�tL1P�V/�t�� ���j!�@<f<�KnFuEb�S�B�bz�P<����B�"GnC�ɉkF$���A��B���Å�VC�	6B�� Svk#]�ٻ$��C�f@,�Rb��"m��Mj�%]6wVC�>1T���$�:E�бi M�%" :B�	�l��q�1Qw�=˄ǎ4:c�B�I+e�z{#ɓ�Q���2�f��'���?��hOzZ��t���W.\2*�X���)D�@�	�|ވщ��UB�ɧg)D�J�'�=���A�A	"���-'D�| �ܛF(��|�[��L
�LB�I�xI�0ДoZ}�z�xÄ�T�!��U�H�jN�=K�l�I%�$N!�$�@��(�G��%�=�g��
 4��)�U��us�"�2�4�Ї�Β鎰�'��4����-f �`CG�@�m��'n�҅X�R� �J�M�����'�5;�g�6�4����܆PN�'��y�'ID�(�;�M�#^��
�'���`�!F�]:rJ�<=���
��� ��Sd�X(2R��%NO� c�բ��$�O��}��"##2��;,W��P�u���ȓe|�ꊱ4  �7�N�f����ȓp5��3�,��>��&�5$p��ȓ�h����w~q�`O�.P�����0T�DJ�G5>���@H�7����_~�p�6�K?��88EM�(q[z��ȓ?���Rc�+Ym����!D�v���Iu�''f��c��'9d��F�/	�f��'������	o
 ���M�yD8Y{�'�@q'�H)ڊ8Z�Ț�p��!��'.��i�Jގ	���jѿa��M��'��q2D��Sy�Ѐ$茒1�d	��'���)��/*�x�R-I�V2vi��'��il M� �("��<Q��	�'Y�݊Ġ�:(pbJ �]&̻�'�p��D�Ua2XK�	��g$B��	�'�0ԋ���.-�|����S�rh	�'0�3`��#Q���j�H:���'[D]h�jY
���'<_�4x�'�x��O?�$�"�%N��'�n�ʂ�L�4n�k�������$�'~F��#i�}gl��',#y��ȓU�~CQd��b�A+Yt��ȓZ�2 QwbQ�q��#����ȕ�ȓy�(Lz�`�<T�fe���=E����L��K��J�]��s���8'��!�ȓxm���6�07(��� `X��ȓe��\�����P���	&Qq�X�ȓ5X���):��X$͝i�:���9�@d)D�����X�g�>ö!��P��D�)4�V�y��= ���u
l�iKC�ʁI��ـ:�zi�ȓ!�N�j"�A�>��f B:h�>���i�B�9�a�zYT���Ǎ�W����ȓQ�B����0Zn��sa_�_b��ȓ1��Q�!A�Y��bI��{Ⱥ��ȓ^�-��M�s�DyQ!��x��y���.�9��#�xQ��� �a�ȓ[ά���ȿ+CLM����;ô���()hJ5`ΌL�(�����Ar�̅�Z
@�XP�#E#0�y��EVD�ȓ6%򠢁Ł9Z(�pbN9����:3���m���F�������t�$��J�;t� �"�G��N���_� D�6�9n��*7.�48�ȓW��XK��l���8��_�t?X�ȓcA���Q^
�@�Q�*�zمȓu��1:�	�b�"d[�٥a��U�ȓr�$C7+���VpZ!�S�?B���u�nu风К��,
5hA��e��fS��Є�ݝ?/��r��M)D��ȓY<�0K�RU���؟��Іȓ[�|� ��H�*��T�K�N���@���0A &��Ю8`ڜ��E���Ԃ�g�J�JT��)y����q�Z��AF"+����٣|��D�ȓ7�WcQ�W��0#N*\7\��ȓ|�����1w���'�l��i�ȓS�$`��v1��k��P�i�x���cs*u��&��i�b�{�(�%`�L�ȓgO��%j�1a�mӄ ߚ]����ȓg��)~}���`W<!�ԙ��i�VyX�E6�DLռ�f���S�? �z�FވP��ĉvC�Q�v\ʱ"O`Hue�+����S�b�t)2"Of�Q�Hˉqq�G�{fz@!"O��i����P���3B�_C�`�"OVm3�Fd�>�p�A��+=0�"O�ɺ�@L����C�ʜ�]/V}�C"O����M�_L. :��+Or��"OxE:��_�+G>ڕ��9M�M "OXXcu��Y�x0#	`��D�"O��#g�M��ݒ7K�29���k�"O.��vn�!OG��1
��f�0�1"O��$B�4�*=����'b��"O��oK�r��u����΂��4xJ!�䃍Rx�
6����| Ӆ"hC!���'2���`�)$׀T�P���	3!�D d�TH�Wg�N��鍪$!�D�.4�h���@]�x����2I��!�� .�K��Q��EhO�>��9�'�X�񂀬�ҡadJ�7�:���'%"���G8Bv����3z�4��'�N��4�P<jϠQi�`�w�J���'Z��S͞�TW�i�0&�j6�	�'88 f)��b�x�)#j���B�'�,80�"��c�X=ۇgC+b�$��'����A�4G���[�!��o��p�'t��KcG�(�"(�F��<�̙�'`za���54#hl��M�/x�	��'ۨ9�!��-!x���䃤+�����'��DZ� �-��0��]����C�'��l0�"�w4��װ�!��'Ϛ�+�
8/�!�hU~�ze��'N�Kvi��X�v�i�+�,z�(S�'.�!A�F��ū�D��RL��'�).��}�n-�Cȹ
�����'v`� A�Z~� c#�
^\���xR�V�?���ד,��=Zज़��y���`)i��+�A�����y*:�pX��!)0֙��N��y,��6T�1`mϔVlB��pd��y��csJh��/?5:ѩ �]��yb\�J�f��d�	:�������y���$H��������s��C�I�e�qɒl;F�H�!�U"oc�B�I�X�Ҭ˳�1=T� ����vh�B��(܈��F6*�̙���QG�B�I�M�A�0'  �Y�'�ilB�I�K��T�ϵZ�-�2B�I�l�!)�4��EH˔e�
B�ɵY���P��
�U2��Y�`�6q�C��%c��ա���K�e&cEI@�C�I	��ж���>�bģ�ÂZ�C�	�V���J���D�cn<r܎C�ɣBIܭ2�(^�.�L��7aPC�	�op�5�����dl����dǷp4lC�?HȦ#��W�+L�����I�4ZC�ɏ4}49��R�����\�c�bB�Iu�<� �e�H8�&��&8B�ɾ @���(h�4xpg�!
UB�	:#�ԋeڰy��`�͈�q�C�<P���Q�~���J#I��B�Ix��`sjѲ6	|��&*H$3XlB�	1%9���vF��e�!�i�SU`���Ob�Or�}�0�-b�	�,s���&��Y��Ԇ�m�@=#���!��P�"�6�`��S�? �� ���:����N~jh P"OH�{J۩j~l!�ʳo���8V"O@���'_3V�n��"O 8����2"OX uBh`��N6�*���"O��)�C5t��@{�ᅮ4���Q'V�h�'�ў�O�$���H�YlH�K�x^(�[�'��a�Ga�6��C�	Ԥl5��K�'��r���wb}���^^@�Y�'�V1��/2�Z��m�Sshp�	�'O����eN��0��R@���{	�'���RJ&IG
�s�'L|�	�'V�D�K�m��̣S�H*���	�'��Q��\�h����&�C�Vps/O�=�����x�\;
�^�x�cPK�98TJ�y�G>D�D�!��|"|����;���J�!D�D1�G�_���r&F��`���@2?D�<a���!6�M�7��*�j��)D�lr��p�<pG�$hl2,�r�$D�LC��P�x&Q���CGc �+.D�0[�̡�N� �&��kb/'�����虛-�%��0妄� �~��"O��`�b�[Y��Z� cg~�R"O^�#Yq"$���Tk�z��{�<�nݒ#�=AW�,F�@6�[P�<�  J�o��AJ�+��`��x�<I��B�n�����5̒@l�p�<�t���̙�Bj�
��p�R*g�<!a��q���t��	d|����c�<��458�aE��^�.#6G@b�<) N@
#�0x+�,�|�d$�w�<)BD������bJ�t,�x�M~�<��PjМQ󂀁�.<�zT�ph<��dF��`K�O4H����Ƨ̙��On"~[� �N�2M�eS�B�d2�1��y�@���o��EZ��S&=��ȓ0t���	QW���`�%x�|m�ȓW�7n�EF�!Fl�$l6@���*��'i�8 aaP�d����yy ��:1Nm�V�C�/0���ȓ�|5X1�K�HȢ �6�ت"=>���Q�|-`4���B�u*��˭.��ȓp����/��%¬��CX3��ȓXLlp��ӡX	ʡy!֭K�lU��=0>͚����zfi���i�n4�ȓz�A���9˰$�R ��0[�%�ȓ2pF#��@W'j���(�+CLH��N���1g��(i��1�b�}�f��ȓW#�i�F�Z�{��S��/F�0���ė'��d��Dx̬za'F�?�����D�&�!��7R�6yړ$��:�0}r�,�}�!�dB.<�̑����T�ȁ�7	-�!��G�ڀ�v� )�[�M��!�	< ��m����(�>�s��	�!��/'��ڱ��2g�@�� �Ȟ>!�D��nU�qC�1dwb���G�|e�y��	6Iq�A�[:8����E�ͼB�	�,l������;�:6J@�a��B�	��$*��m�H\�� "�B�	�^��� ��E<��1oF�B�I�D�:��dP[�H�!�#7-hC�I�r,�����A�!LD���J�nɘ�Gr�q;��An�YzΉ�a���R�C�<5®��EM0w%�@����C䉜
��sD.��g�x����7��B�)� x�Z���"��]��!Ex�U"�"O&y@/��!�p`���݉2�N@"O�Yx�OA�$!����%pj.P�`"O,�PB�AAڇ��Ҩ�"O81#"B�GX��!$��%P��#�"O��Ԇ�(&����ҖX����"O`U ��X�"9�a�J�<T���"O�z��;v{0���ƼQ<�L*�"O T&▍C��2�mX��A`a"O�M2��R)�f�b���`e"O�T�c$��4�j�r�k���RV"ODڧ$ۼ4A����ʚ� �:���"O�����:fu�(��	o��m�"OVxbE҂tE�适ʗ\���BE"Ol�sU�� (����+[�(����"O�푣��/���CL)�Q	�"O�ͨdlx��r��ZR�I"O��D�Q���ȶf[|��-J�"O: � Qń�Ƅ�E��aӶ"OXEr"�3i$�i�Af�6s��pk�"O��BnK[�^�u�I9�l��"O��Qr��9��m�fDL�y�&,i"Oz����ר>T�Ӧ$z��I�"O��Ѩ��x�Y7#��T0F�S�"O8���'�{���S��Î^+�	��"O�h�`�LL�1� �)�@<IP"O�Q���,9����ےWZ�(D"Ot�F�.?J�4sq��u��D"O��ǣ��y�0�9�B��iRF �&"O���!�%M�0����!)M@�Yb"O,��6m���5�ۼdAv���"OR�� �\�D��B��F�]1\Q�"O��FIZ:�d��/@�)�� �"OBGj����tNӭw�~$W"O����I�Ti���M
&�h�y6"OĈrD�
�Vi�G-�l|�5 D"OF8{u/��0�5)v�N�GSp��"O�%���LX��k6�]�"O���	!;˶�*�%�A-���t"O6x���I����`2��A�u"OX��RnΗd�����S"ODD	�n��,G��!�`݌S�Z}P�"O����^d��Cb
�N�R��v"O��K���#T�zeaQ�T��D�d"O4���H�1C�Y��iX"d���f"OBP��OK�:)�Aà�����,�J�<�u��2I��0	��hy��b`�Hy��)�'|�� jt� ��0��ȝ^���{�&ݛ# S�V"@-�ǂU�(J���q�D���MI3����bpC^��ȓ-(��!PB^J2��y$`ԕ+ڈ��{�Ycn�Y9ʬ��NP�7�]��,�P=���)}`���~� Іȓ)µ�wa_J%x���I�H��ȓP���α1�
1B���3�t��BY񑔡
x%�R��_"��E��wB6���W�h�r��V�%�~ ��@l�J�Kι ��r���'D�p��fe<�1��Q�k��%���ĜF� ܇ȓ@;�x��D=ypν��eƀ,̰�ȓP�,4cF�r�|�1׆�uiP���sy2�'��	ly2��˕�L�Mb& ?o 虲�f�4\�!��0'��Db(�XK�H��� !�$Ϊfͱ�̅�|�䈀�P`�!�� r  F�Жt	���w�X�2"O��R�Ȍ4@Uh�3k��й4"O�᩠,B�G.��pa	�]��Y��'�ў"~R��/P8�L�/u<D��b�,���0>�լ��1��rЭ�:"�� �Ly�<���ЄAO��Z���&���d��I�<�s��l?z4�eȞ�dV�iA��B�<٣B�D�D��BN�&4\iG�A�<��k�넕"�,T�BäX��.N@�<�P��~d���~��ܸ��Zw�<� j�Q3T�bc+_� I��P��Ο��ʟ`$�"~2�^�c0\  B*��9��戰�y�N*N68S�i #��g���yBM�*�r�Z��Z(�*��$��7�y���sR$	(0nBAL�RĊ���y���3l��L�f�\�,�,L
�M��yB�D�kY�9��Q�$^\�r�Ʊ�yB��f�����l&l��ř9�hO���I�X��Q	���-/�-���X,d!��(��|{��{�8�W�,�!�@]=2�XB/8D_�USBK��.�!����(�8��.�`Xl`�!K��`�!��	��BE>|���`�O
H�!� D�@��@M��4s��v�'�2�)���S�D�I�R�*��i��*����O���$�'
�D�ӗM�00�єҁ>�!��>vO�����Vz�AjV��8!�D�\��#�ݾcl��Ȅ�҈N�!�$�3F:����܂i����	�Rt!�$�?I��ٱ�ڏ_Y��ʶJ��=r!�$�Q�����5YYA����#�!�dͪ=Zx��!A8?(l��a@?a!��E� �qF��N!b�q�K�,K!�d� 9���9��>r�P�[�l�!K2!�ա/�f����:U�5�TKG!�d]ff�H���~ƾ�SViю5!�Ě�W	��AFi�S�-�
b���ȓC+��p�n��+*lC���*�~��ȓIBT���Ǿix�M�d͠cVP1F{R�'�&(��$%��
�cY�M�����' X\�F/�ER�U��(Tn��'�l��Bჵ5ܒH����YN]�
�'�}h���;����UL� (J�ā	�'�8س�.4R�e1`��-�� ��'L��c��&;[�p�D�\������'���j�@Q�]�XPt��@�ZH>(O ��I�,s��'�� P���Z�*!�$X�=��c �n��S��0h!�d�_ Rq��g��v6U�E�ƤpX!�Ğ\��0���A=T�����\}P!�d�����6�ꘪ�f�n�!���-)����ΊTڸLBe��U�!�D�h�FHR�JZ�9�8�i�BG�L �'3r��7�Ʌhf��F�	�T!�K9'B�	�jk���E��F�r {��'��C䉁3`m��Q=���t�N�y�xB�IҤ+1��+#dڱ�勽sAC�^9 ���nΨ;������T C�ɺ_o⹊�؅X'bB��"��B�ɟO��4��b���t�0���}�BY��@y�'�ў�O�0��Jh1��ksƈ�R�R�'7�A*GE�I�����47Ʊ
�'e�\"�¯O���h��34pI�'i�z���L�L�сǬ#������ �C�e�)�� !�oP�v@�tp�"O� �'O3l���^2n�Р""O�AH���7�PQ'HJYh�6�|Q�@��ӧj��0��#,$m�S�K* o�B䉰c���H.P���sԪ�}��B�	� cB����D�#���ȀbO�z��C��&�^H`v��	lV��o�	�C�ɩ@�"��ՠ� �z��F��#+D�B�	:L�v�	S�w)��(P;R�B��2 �{UO��	�^Y�`M�V�B�	#|1�,;�E�>>,���/aшB��3\ܩ`l�`�(pa�%+�C��eQ�]�s�Y X� U���P�\\C�	��$K�C�U� ł�f��^�C�I�"�ͣ 
�Z��iy��F:ve�C�	�x���wa�UX�Z 	�2��C�I�5dvU�I�(Qi��6�O�T$���D����� |��j������;�""D��	�b��W�H�ďͪ=��4S�>D�Jg�:Ot9�����-����@�)D�� `�݃:�L@􏙆^�b�pC�%D����$�����
]3��ԠF!�B&��\��$*��)gbX�!�Ac.
����k�*%� o͔?pў���K
ņ	mE:�D�*'��B䉱V�a8�E�9Nֈ!��*��B�I<�RpuI�����H;��B䉼/^�e�Ԅ��`�l0�u	�'dj�s�@�5Kȕ`�DG' (�
�'�)"'�j
�1Z�K��U�3
�'�ŚgiF+�*��G�|���'�(��C�8���!/M�V�Zz�'(��x�dʴFߺ�+�M�2a�'Hd���k��|���B��܋N��h�'�`����?R�V83�t��'d
T��$@�2�JQ��H�'Y�)
eN޽	(���?��XK�'	��+�O�e�����˳u̘d�'���sFI�0?����uL�r�'�:����O��&dShNt	�'*lT��-]>A���"��>Ø)�'����3N�W��x�#/� Z}��'���35e�Cc~`24��%C ���'/<�����+w0���g��x�� �'DLq⑪�IaH��rcD�q��<��'�Pb�"�.���+�ۚ|c�x1�'��i�Bf��c����F�yJ%[�'�NU�B*L&��T�V�r^� ��'�"X"��~�42�����
�'�];P��5<�0z`ƥf/L݃�'���1V�M�x5:P�8X�P���'�c�gE(���G���d�q	�'h�q�bB�b��7�a�k�'���뷃șcݒd���O4JN,x
�'�fSa��T�9Ч�>NL:�	
�'�&4x��B�t�XtϏ�G����'ڦQcD΂#�M��Hŋ7V���"Oؠ:�V ����h��1�p��2"O�F,F�!*�颷�ڜ��7"O�5���W�����O4VP&e�5"O �p��ִx�@����{瘨h6"O��1G��~ʦu��-���"O�PA@����
Ԏ߾N��H��"Oș�d
�] ���$��n���S"O� P�c�4'Ȏ� b�
�B=K�"O�"�k�)�쨠b�Y�!6�Q"O�`�c��<E�qQ���
b>y
�"O�q����*a,�����Y�?�u"�"O\��4OҾ�\h1O��_'I�5"O��
ư}[~�u�T�j&^��3"O4��C$�u!b$ݞ	����"OD%Z��.�6L8�r��Ѱ7"O��P/J)^�ڴBI-��e�"O���2���2��ź�@ڿp���"OA���!>=����׌Y�&��b"O&@��Ǒ h�̌�$��n����c"O����0���C�S;8�j���"O��̹B�<{wBٯ_f��0"O���"a�g@�~^��"O(�@`[�E��(2�	+kh�E��"O
�J���_�F��4��"_P��Q�"O4Q���\8&(T9N���R"O���P�Y�&,�����'G~��"OjP�FΧ���Ƈ<l|�6"O���*�z�Z����0��0�"O���ŮwjԸxe�F^gҴ��"O��sR�/b�r%�ʣ'`��s�"O�-����4�����
�+QlH�"O �'*+�Tv�G+�6���"O*DK�C&}p�X7�H�*��"O�؊�CG}�2hR*�$*e`"O�D���
��U�刏�f�=AB"O �bvb�R�JӍȳG�h��"Oi�Q�(�6��$gӚs�T�*g"O���PT%]�\�qc�j��5�"O\�q��fF� 	.@hU%T��y��e���W��l)(���NW�yb�)4Fa�'�<W�mSW�Y��y�����U]4;�<dw(_��y�["XȦ�bUK��7ߺ�ba�C��y,�n����E.ؒG�Y�𥑄�y�3�D�S"ͣD!�us��X��y���0x|ZQZ�+��Bp���Q�׷�yb��(|D��"�]/V-�JG��y�+��j>`������$��<s��I��y�6'0T��ϗ�#9R�aЊ2�y��yT����n�/�����^�yr)D������)��(ͨ�(��ߎ�y�,V 4p���%�)3�
V�ybE =O��|�S��P�%k��R��y"f%F(�b�0�iʇ%�:�y�h\(���t�08�N�*�!��y���`t��!����3I�E�Ō���yBl�/p� R�
��x~��"�j��y"@�Z�h		R��4Z���R#���y�DD���Hk�U @����c�^��y����[����#��
<��\k�'�9�y��O�Ԅ��e�F���0�jA�yb��ri�=DER������y2h��>��;��W�<^l�P)���yb�?AY�QRNߘ-(�5B��X�y��Y'1��p�7V8n���N��y�]�`�:Q��|ڎIc�OP8�y�J�N��I�d�.tP�����	�yb��y�v�R�oY�sx����Y<�yß :�|��$f�o��M �S�y�kа ��ɹ�>R5*���yr��:�}rMK��|��b7�y
� R�����~���#���MG�y)C"O���[�&|�C=!��I�"OB�{D��Q�`��e֡x���"O��"�L�ef��4�8�:y�"O��*Z[���q�^�0޴�G"O��`��M#��)ŭɟ����u"O�(B@�O+t��@���<<����0"O���OYN�:t�w X��%cZ��y�iQ3��)�bKL7h�&��ΐ�y�cL~%c��8KЎ��'�ý�yR��Z]��i!4Q)	��Y�',4  g���� J�Hz�:Y��'���q�#ӆ8��[��2L��	�'�B�����7"a�d��m�0Q�
�'��	�0OX!'��-�R�$O�X�	�'ќ9bs �t�A@b�0A,$��'~��q�J�L��ZfO�<�����'������*�qau�̞4o�5��'��ұ��3+�N��D�3-r�Aj�'U(E�FT��~]�р�%x8J�'gp+0��� iE�t��`
�'P�uS��-uZV�y��G�p�j��	�'�Rq���8X6(����rO>�K	�'L��"2nP?ݰQ �gvv�2�'(H���B q����L�&o�~M��'U$h#�
�S������a!�	�'g�1+G�
'���BAO�ia#�'ŀT�f
'+ :ABUIJ���E �'�T0sU�4v�|�!eBү#d�1�'�pi� ��j30lID�Źq7"���'��-��c�,Q��{�$P���Q�'l�'$2Ѥ˦,�&� ���'.Z�С̅J��9�V��8�
�'|�,KsT�5��3.�D�gϛS�<�ą�8f��d�Ô^2�`��R�<����]OR�h���Vi%h���d�<Y�Ր_v�pp�Cх7T��)	`�<�!. :�t����<HxZ��4Ϟ[�<)���8���(�*
�T ��p [[�<��ƌ����=�|x�TŋT�<��Q��Kg�W���z��]k�<���O���q�ܖ5�z=���N�<I"�UY��ag!�"��4Z�	�s�<q�e,U�D�bDf� WYfuh�S�<�B-P(@C5b�H Lg����M�<�+S��>�;���"<�p@($C^�<u+� bv�q�t�)GQr���c�<�V�^>;�,�������p��� \�<a��[�c4��Hbڭ:�\��*r�<�m�[����(I�]�P��Do�B�<�G#N)Q�����mm�JF�<Q��˭	%b���O�>|.���$�<q˂�k��)&lQ>WJ��Z#��}�<�E)Z�C�����h�f�����U�<y��lg��F �,8�	�J�P�<���3vL����Ȓ& ��2�LGI�<� �')�b�ʄ�]b,q
�j�B�<� &]�u��̂SF���1�T��A�<��.?G@�5���DqY�I!@z�<e
�d\Dn��@�a�2�yr(ښ3�<91��.=n0����y���x�3�]�7��,��IS'�y��ܭ>	�	C��YfA�fX�y��������@��V�T�3�݈�y
� $u�E�=A��<@�#YTmHP"O��5N��>|u!���V�tP��"O,�a��]�_~@E���E.�Y1�"Obl���ʡw��ZqnM7���A"OVk�K3P�tM��#~<zS"O$��69S�9��?2G"O���*i��"�t�s`"���x�<��˅k|ne�G��~��}�x�<QҊ�:��\ٱ�ދ>�v\���H�<)���.�f��� ��H�D�G�<����*u��Ը5,�1�� ��Ai�<Q%��
)謴�R j���
b��h�<)V��5	�|г�53�VX*���o�<AɺNK�@$Iǧ|�Iz��l�<��-%��)��)�#C�8-*gE�p�<��+�F 4R� �^����3G\p�<A���7'�QSCF�8���W�<���Ҋzt�����]�
�P͊A�RG�<qW�J,Q|��$��p��գ�<�d�ӕG"�ש� a�E�"cV�<�C�ݯ��Jf��m=����GZ�<�&ǟY�}��D��*�4 �P��<�ݞG������l� ɱ�DD�<)
ɷ? ��u �x��p 	k�<�F�AB�p�/��#tf��B��j�<��H�3F&��vX�ln����@�<t�V
�����Vr���B�<i�H�BS�$�fn�>bC Y1@�Z�<��Z�F�-y(��u�YY��M�<Ac�9�0�%��+R%&�8f(LJ؞�=�a}���J�E^�B*dH���E�<A�փSI"qٕ��.+�r���NJ�<If�'հ�iiԳ7�F�I�n�P�<��A�nf��e�ƭ��}��N̓�~R�~���Ĝ1hf����F���k���K�<1J�,*���`l��h!��ǬGJ�<���[�t���K��	�l�yp�SC�<�����c�΁���X���H�<)�AL
TP�N�fĄ�E�'�ў|�' I tTq��B��U*M��'�:p3d�D�g�(�j �ԍt���	�'�"�:��)��(��v����'g04�s���Ȱ5ywA�g���p�')��`���� ��� ga2_Ɯ"
�'GtⅯ@�Z��J�[�7-JUI �&D���挙pXIJb��A܈t#��#D�0��l��=�R�,�/c�| �D�"D�0с͋��x���o/^h������'O��Y���$J�4��xi0��'J�B|� qӒC�I~4dYBW����!̃�}��D�B��<��O4�@Q3lgd���K_�jx\Z��'��'*P��kv�Y����&=�<��y��'B��	,�'^��QT�\y�[W�޶Ʊ��	2!��O������ `��O(Ԧ8��'�ў"~��O�s�ję��t_Z�Z��'5Z0��M۟'��)�i�/K"� �tL��l�r�m	���c8��o��F�����Ԑ��F\9Uh�}�'�ĉ�a� ��~��~⨚�g��P .�e�ȁR��-��>��O�����D�f`H��ŀV��ը�U����ɿRd\ �S�D�F1z�J� %O�~����?�"��9]Y�� ��i�d�T�<�f@Ihdś��T�_�ty��Oh�<ѕdȱD8�u��C�PX(U��H�<q�^+�0�� K�1�ِ&Mߺ1`��m�L��t�S�? "��b��o
�9��
-���ku"O,詡��_�`�3����U����C�'��OpE� �*qu
v֨;�~L0�O���ъ}�̊5B�* f�h�^�!�$�"骍�&&�8N��U��O�!�(qy8�@-"��䐗f�	E�!�d�5Kd�Q���X�ct��^�!�dܖ?�Հh�iڒ�!���={ar�ON�`j���T\�C�=��{R�	�<���	J?a>d���� w�:9P�)ךz�!��?���u�H�x��Hպ-�!�#x�z�L�6kA,��g�^�!�䓊;%�S4�Ɠ.h��g�/w7�'y�|�e��%�l�K&EK�?J�����y����2 �Ā�����Ԃ�<�yb���I��:.
�ܻ�
	���M+����Y�>�H�ǃI��dM!��"R
�i#�P��r����&!�d�i0]9�BX�w:8�!��U��	�'����I^?+O��a�D"L� �� �E��)�l54���7��@8@�{0a_`jF͛�A6D��hA,�rn�{���G�%�&�7D��Q�Ex��
�%�v��P��6D�|[SD�),X[BHDb�t7")D�4
A�3R�"�����H"�Q�s�,D�����/,��s　�q�`�2�&D� � �1��a�iD�N�j�Cw�"D�@���"QzR4S��5kAXeBRm"D������p4���+@CF�xSsI"D�t�C��y�⠚%�ߞ�@!�S�*�d-�OPa�`^1;��K�.�*���T"O�HY҅�#]1�\w���t^�m��"O~�0A�]+?��9	��S�R4��X�G{��閅=���B"`�5vLM�c�֩bs�<�ߓd��xgCWm���w��.? ���IJ�+�91O� ���ᕿ� ��k54�%��2��BwL�w�i�'V��?i����@	�(Kq�z�H�H�ġʲ"O,8�7i��q/2�F׫n�c3"OF(���,o� k4��V��y�"O����߯;
t:���O]�����$4\O� (t�T(D���B��BURUhg"O�P! (R�Z��b��HT
�"O�x��F�l	�	h��y�"O�r��L&'�|u)�A� Q���`"O�Z5��v.B�W@�LGt�A"O~E9��N�!�����(� -�t��	h���	D+*k�p�酁Yk���N�"e!��m�Q ��)��Y�'(V�G�!�K��m&�� B���3%�$<�a}��>�B*�6`04��"�����A�<����'5���B�cneF�^����?1�fWg�h	��b^NT����,Xz�<Y�l�x�&*���.m���r1��Z�'	���O���1�E�l1���Ύ�]O(��'��.�0��I�Jn��A�6�y�C�΂X����(O@��DL��yRo^
/~��1�S�n�I�ui��n���$L�$bn�[UIЗZ�P��%���!��.za$Jr�،���W	�!�V�8��8�A1��� � �#�����?�H?	`�dN��x� P>n�񘶤0D�p�#�	!��`�cBZ%}8>e� �,D��"0�B�y0��p�3r]M1d�.D�� ��)Ѩ�v�љ��S~8�C#��0�S�S�y�h�vܲj�X@��@7ekbC�g[h�ZU�]�.�
Q^�E��xx�'űO?�n�H��a�'>����n�.i��O�':�O��	�1�KQ�^��`#*�� 6"OH5BPk�!����#�5Zٚh���|��`~B9OL�� -ǯ^�TI�1!>t�kB�'"�'6<���)�_;h0�����@��d%��HejS���RSn�Kv.N:�B�ȓo��T�N�>:,^H���[Æ%�'��'��)�Y�:&�'aP����33����1�O�d/��>hJ�H���&�Y�@ٺ�E�'�,���p=ɀ��*E��m���Bh��cFf؞��=с���S���BU��}��T@8T�d�D&\���ز�+�l��U�r�,�È�$q>��nڸlPV���Ο��Ԡ�iU6\C���FX�6�8g��U�#k ��������Y����G:+���s�Pr�'鑞�ce��B������%m�*���9?qF%!�O�ɐ�X0���Ha�՟| "s �>���)�S͒0�A�
鲉�ta���ʙE"O�1U���m��`���vd��X�ϓ"qO�#<�Lޟ+9��y��%WR�P�*�Y<Q�֟�f�����V� %�hX�~r�E�ȓ��9LZR��d:1)�>L,D���o���B'D�,2>tݣ���;0�ְ�ȓ0�@-�qOZ�,��5��a[ 8Ol���{1��a��G� ��a���R ���ȓ&��Ljf'��9�U`kZj��`�ȓ<?��MT(�l����&&�2��ȓa�fHq�e�X����7Ț��ȓ;���3N�56�=CV�1�XĆȓ�P���	n��S�(_�fE��l������;�]81��*E
nH���<��`I\��pb5��9����ȓ2�f��%�|���+Tfƥ�ȓ��b2 �M.�:�#�	pپ0��+}��E�д\cu2�,�t���ȓl���@�\-�`� G��!8�4��ȓ�,{��?<����M��Ņȓ]8����J�X\x�d��K՚؇�Bh<y�0d߷n��5�P��9,6���R��E{CQ-v��!G�,�xT�ȓ��k�, �*8�D��s�Շ�:�}�0Iy�̄*�EJ)L�fi�ȓf����ǂ�\` ,���ʝ,�\І�&:rY�S#�7"�ԩ��^�~'PɆȓt��|i0ڶ,ji�a��?"�\��_hN�!Ƨ�
oij���^�+�̴���<8"'[�9�ڸ�(�5J�!��%Լ���B�&�8��y�HC�I����aޢ4q$�xb�O6*��C��WR̄
7�:(���F���Z��C�I�b˼�)'�˓.mF��t��"��C�I/6���e��X���HʷTp�C�n�!�ѷ]\
X`Q,�k�jC�ɅC*��q�E\)�1C�V�@C�ɪ7%8Ey��8#K�.�s3D=D������eJZ�#��3�6%���0D��"U�H�y	x��N���Kcl-D�0�O�$e�v�q&*�6�ؔ�E�+D�� +�1�8�a���S��cc)D��㓦UL�N���e>5����V�g�H���]Ux�+���/n
f��cF4�d�Y	w!,np-�a	l��m��S�? 8k��'8x�A�eʫ":~�ɴ"OL$�r����Ph�Uf�c�A0�"O�I�@L �F��d��K|�D�G"O�ik��?~ո�S�Ǝ�O~8��"O���f���:��sD�0�x��v"Of��W�~����<_�v(�g"O�uB�Ƅ�2�UY�fɎ��%��"O�8�F����Q�.��s�"O�!��C�+N �H΃�ԭ!�"O��a��A�:��2��F�8��V"OZPs��ԃQ*���bݭ&TD�p"O�x`�%��r�X%�[�94H���"O��(�ߜ��XX�o'D�4���"O��#�=Ԯm���Y�b�ԁ26"O�PqV�K�Ah���a��]��ce"O��$����A��.h��(c"OLIS�I�qĤ�QH�qh$yP"O�Q
�-�|i���r�V�O`�#�"On�K�Ƃ���lO '}�M�1"Oƽ����1/��I�.˂����'��Y���{��=w��y"tm1L�I��c��C�ɖ+Al�i��߯HJ�L뇏W�V��'��Ё�o�/�6��Ӥm��ͣ��ǇK���%7�pB䉢m�-��]��+�P{��=�F���<��кS ��'+�"��Y��3���3fn�+!8����V�2���!3�mx��1�ŭb垨�W��=	�	4�'F��\1e�G�~AP�����Ab�ɱ��	YO�zE�4��'��g��H�#/�W�|�T8�2���Cb��X^��їEN* j�]�O%܀�ƈ���X��w�� [s��E�͘o�"��!��6�{���0�+�wr�\�宆�8�uy*��j��]8��M�Y�z�C��|�&Kut�@��9�ט�X�v؀��O+e��=r�w�B�I�KxP�2%,��"ޒ����9[ �=�Ǖ�S�Z@bm�@���E�Z#H~X�2<O��A`��^,�睑;H�A�weC�m�"ʖm�*��D�S�:HS��I� ̢Dz6n]<<��*��ǲ^�f���c�%d��ͻ�ˈ �?�E�95�p��>8�� :�{��I�����+,��pz5���O��� CD4I�L1m\PU��\�nt��B�&H���3fS�&YLP�� �<t!�x�`K�;i �02��	4ȇ�	�h��1 f��w�|Ĺ�IڙBY~	��i,�7��}���yWi��=�t�1O��B0���YB�LH�.���4 3D��`ToҲ%�Q2MBŸXR5GЈB�*1["K�"�4�@�$Vp�0ԏr�f=J��/�Y��O��IR�L�)iF�l �#UM�di�ff��� ��v�'���겍�9&�-p��L	m�hP1S�W�~�~�:��c(������2�r�ҷW(0���a6��h�zD	#ϗ�}�t�
�O��	pG�Ҽ��b-4K���B�5~TdY�����!�Y�5�[�k8�P�we�:	�K��&v����ϖ�L�)��OU37��@:��_~�j�ɔ.�n�P1�'0�Ջņ;bK�/o� cs�
5i�`��"��/�\��6��12�J� &�h/L��b���m�$3Ӭ�1`�L�F�U�*��mB�^"ⵥZ��ֹ�/]���}"���!_Z��|�H�0��@�3�I!-�� #�H�8*���g%�
� ���M30�ν�B������$�B�̳1�ڝ����z^\�����!/�֘{���O�H$c��WZ\`����c\��
�2��OrTq1!�E�XťQ�׾őwJ	Q���ȗ���?T ����Z�|���X�{������
а�ɷ��	Q��Ĉg���`q���!C�^����*��.ؽZ%�"=!���Y*J�gN��b�'L��Y-�%��Jp�h���}��H��19Kd8�T�V�0����h�`�  �ㄆ�Oh�CN
x��`�JC0;Hb4�d`s�4��É���n��V	['�5!�Γ=?��XV�x��4
$�-qW.��:��cЈh����𢚒p�u����Ib�*T'�~�����[�
lH��ԁ�.Cvh@�A�ٻ(�m�&T�(Oh};�˅:�H=��S�\,���ip�����漴�`ʚ"\b����W
.���nJ���Nɔ��=��iF:�<%0�c�+�D��LJY�|�ɓ�R�@:`qD}�l@(˴@���ƞ8rr8Dk�D�&t���C&(�h����D�ơid��z\:l��v���`b�3�jm�"��Ǧ��UoWJ=1,�2Dpd�g@jX�D"8K�B;�"��c�6ĈT���M�QɓcE\<+!�� P�`�RXj#��V�+bghU��5,8�m�"	jd��R�F�S�D��X�n+����Z)fn%8m@�=���d	#
^�T{WC4T�  !Q�;;M��`�4v7��:On Aw��C�ؑ�n�k��!@�"ь�� *�↦H�8���f��n.��Q��e'xD�MC)Og਱F����,Jf�ǤL�2��DF��~B��}M���$�ֈka2`�2V��o� �aMOT�ѓ"�
4��Q�邬��d����;+��H�o��BOJȹ�$��x���@�%��g�~d{d���L^y��,�fX�R�o��FG�i�%�U�{6�j��ԸJ����KOV�41��	t�N��d�]=Z��p9u�h�� 
1�Q*w�.����,� qB���
�)�@���hc�K�Z�
q"�R;C��1��J7�ʓH�3 �Ѭ,:�4���"��Ď1�5����.$&!��X�j�����eS0���bS���-�'l��BDdP6��b�R����Ǎ�?&X�eB�-!I#�e�2AR19 +�B,4#D�4Yh��d����"�O뮄�[�2a�d , t�p���B�\X� ��3��@��d��Go����$ؼ2�(H�K����ef��ZD��s3쁀�p(ۑ+ۄEh������I���Z�9 �b�P�S-bAI��r����# �,��ju�֕9 U�f�۹38����R/x})���i����4��m���`莟*���1N��MY(�f������ ͙�%�?��ċ>B:`�;D�r�a��Y�	0-
x��x�&$�1�s1���ޔ����5iJ�=3A�N8\�=X�m���X���ܲ�@.��&��2��U�,*u%N+��+R� ����W�}�����'
��G�Ǻ����,*�^l� E�H���3�HI{�т�ŷYx���o>!����a�/-�@@�P�֛K���k��	ڼ�ˌ2�(��e�ؾ�#�ȟ,c ��
_�|HQ��OH��&X��I�6m��,��,5���ʕ�� Nx�\�V��{�.���⏬Z9�tGʦlLi�7M�;"����!��L}�L�v�Еy� �s�*�IƲ,�V`�	�#���'k�Ob0��*�P!���!b���zP�1�M�@�D�4B ��/փR 6�h��O!z�5[N
�<�DКR'�;a���H2g��6�l��pGM�e���P"�I�V���S�넑qutCA�V�0�B r�JL�A�\<y��V3ql9�L� W���k�KD�ptt	k!V�2�HR���>�U�C�F�|1���V�aF��@�\�;�f�1˓U�"���u6l�J5��mR�0cN΂R��x'c��VԸ��2��8ݴ�h� ��Z7�y�F� �2��w�hX��d�� ��!�U+ש�`��]�ĺ#3� ��v
@<@QphIpg֪*����-A�k�
�#d��uz��r�^�������BW~tq g��/����Aٟ|I�ە����Xb�I�-:�9Ӥma��ۗ���䖍[j�iۓ[A#����B%]�Y�Q�վ��g��t$0I�OZ�`��/s�D��`g"� 0B�`0#}#V�2�N�eF^�ml�`0/E�V��A+1̉)5
t��q���R� 5nv
 c�W䘅h@@K
"TRvFI:A�2`iu����G�D�P%I��&x�\ʶ��Ph�D���M�7	�n�!I�U>)��IߧR��A{�d��x�2'�U����GυS��	"�D3�OXa;4F�j\�P��,ç.j@�0`O-���A5�^�o�,H�f��l�*ۙQ����&�"�W�uz@"ϛW��X�$љ`Q>t�%��iUo�<��e� o���#fT�:�� )���	WH9�f�O0]�2eAR�Q	P��+4���� ������M#1@�{�����l2x@h@�)bM�,X�Ǒr雦-F��S�lțD�B�\
!�p��`��W���Q�DO#0�ԝ`�F,����._�%lv����[��MH	ߓY�E��n�(��`��QTL�T@�%0T(M�B ZbfH��M6Pb�e��(	��HЦ��SZT��`�5X>e��@ۏ�5�D[�В��6��+z\�a��_��O���k	7-�=	�9�?���>C��@��� '�*`*�'П=��vlé[\��C%Etɡ�n�c�:�.,����9���aw�U1��䊌|��iȢ�s�:���+�`���W���(�< ,g�B��1Tl�#��O�y�T�_�H�R��r��!X�j�s*�$5l$���ݏ
)xݪU�V�:��]b�F��U@��,P~Ն�I�aND�� �b �S3�ĀL���ɗh4-k�$ bL|Cb�k>9C��Y�&bAf%;�b߈T,ܴh��!}9�<�q��|��h��-,Op<Qr��.��cA�DBS�ĩ�,�%|/�t�'�4M��)T�
(�
P��K�/tHY�4a�DZ���r�'~)�d�ڴk�,��J;�D]r�¨u*� �끼1A���?��;x|b��4jO�U�Xb�O@�髓+�5�.5�ѥS�I�.��Ҩ�='��S�)R"U*����C8-� �c�4�(9��œ<H�(���X?�	*4��@bΏa�f�`��S�C<Э
0#,��x&o�O8�*�]�4��P0"��`�b�hЄӪB=��݂/w����#�;�b��&ϵ#J%�ɉJ8��cP�W�'a�|���B�'�������O��Ar���-G����K����d@�":�����ШA��y��H*H���E���`Y�US}�� 2ÿU/BT�IADcayRL�|�L���� *�����N�W-�I0�-<�fى��/��PQ�b1��DV*̀����P!�y �	�%=R,���ٽSȵ�"���+�qOX|��̕�Q�>��0B�/��� N��J�^M9%�r��b�k�����C�c���J䡔� �pM��̭:H.�Fn��"~Γ3�8���_�?W8��V�5�h�.�8I��5��eS�l��M�7�4��ԙ��`��y�����jD�QY��P�FcU��~rC�9���0��6�uF�B#H�]y�fX��9��\s�8P@r��m��(1a2J��A	��!M�AA���
�MKf)}ݝ�$!т#�-c�����^�~�����:<��Ҋ�D�6xg���cy1j���_Y���$��`�9 ��7���$H�*{B���@H���rQy��@���.0��� (��T?1��>N�C#DN1XB���G1�d�`�����b�B3�#�I7co��q�뉛y)�4J�C�T���B^���%ɥ(�m���I< ,�S��ے]��S�O�ҵ�qI�YP"H8rc�g��Ę�g������e�B�"4,1�zzʝ�����٦=7��ͻ(�H����w�RId �O��O�
��@���<1%�,mԨ�k �E��E��FW�cRB�i��!�Y��$�z�K�3,�jI��m�/$�M�=���:`�t;�ㄸp4�3�b
[X���&��t�r0�NĖ5���p�*b	Z�KdD�t8������Rr�j6��9AL��z��_Z���h�U2Dؐ�އ<�p`��B>�d=~�ɘEĿw�*��
���@GY�)WN�;�gѨ|����ЄT�1�G�R��ȓ7�¹�HV�gle�ĉb���(#�]�i�t=�A��0R�Z�`6���1�ҥ�6�|*A�3u?�N�7jc��ːa9��X�R3B!�Z�zlB �w*F?ȎIɠꇂ,5��GfE3y�f��3Lؕ�z$�"c��xiL ��jǛ;���������Uh�(��0��!e�&<O�YH�ȋ�4��l��+��@7`��Z�];���8t.<�Q�
w�P�ժP7'�f�[��'@ԁ`�,�ki�8��CC�q�ഒJ>��#C2s�b��G��5���O�6 K���+DЅ`ĥ@%P�x�*2�+!*�q������y
� t����N� 1�j�E��"�>��T��I���0�)&^�)�ҫOxd�����}�D$�S��杭6�*��a+�-48cL��TΒO6<s5���O�x� �P/fN���@|��z2�N6#r��q�(]	&6-�=PL���6�Π]?"�KA�8���η w ��`�&	CR�B���/!�x�yB/.2e���dU(&���R��$����'��a��M�Ca��q��A�A�h���\*��Df��5/�4�'��y�Ow�q)O�)�L�fEB���>Y ����Q��I�x�\�a�*���H���-J�X����%[�Y�RJ�˟�	ׅ�?�|M�&�ƛ_/��(���p]����mW�l�b�ѵ�
�~���74T:}:���(l�\�PV��_�&A�ҥ�����D�`������50\*]�B(�u�"�,�l)Üw�*I�U��;	۞�*P.	9m�Kd@��䗀vA8�)3DXc��{r�҅^�nt*R�P5xU'Q)�r��#
G$ 1qQ�Gе0r���o�;�zXB�c�0pA#c�-�l����'!\�xz�$\�Ϭ��woM ��`sS%M&5L�Fy�\!Ǹ�؇�L#��tC�̤0ڐ�ї�?�(u��l�>
��bmH�y�����S�k��A��+-ӊ�ѷ >�,e�,�;���D��@�w��0^gZQ�o�g����'�Ƞ��o�	� 	�Ԛk��pK�)/��M�P�S�V��F%M>w2`B�G�"����&F�;S��[G�V"j A��A�kd\�E�~��~B��:/R0l���&u��

�N���Ń'y�X�a�5k�x��+T�)^$L�W�	 a#0����y� 5[���!E���8�۷�ȧ
4Y��	��Qlh8�A�:{ǚ\b�g�'6A��)K4�2v)� '�BDq�@��� @�Ꭱa��<p2�q�+�)
 1�,r���%�\tY�l ���4xCE�{�X1��mT##�|��f��9_Ѐ�w�s�'��A�F��h.EC�gY�+aT�C��<e��CfAF�9x�����j��֠Y?a|X���-���q]<g ��sv�F$>r�����?���D{���1�gD&r�N�il+}rF�N��"�蘗p�h����57l����+5��Ea��'u��Џ��� ��ʮ�xg���s����g�������%w�?U�# �w�
��t���W�����a��y5(� qnN�8�nR���+0��#������!����;ZV�����rU�H!���F=$�i��;{ɬdA�e���;DCٺK���ݩH���j6`�$I	�Ѱ$�� &K҄�d(J�d�\����I�X҄M�I���r M��uW�a� 	�*"/J�!���	 żT�X9S���5$�-<ڕD~�
�y�ȝn�Q@�)���J�cJ�!{�� }��-�sd0� ��ٲe���k_�>CQIc!dC�vG]�}��!�cT>�QaG�K|n��eb�a;d9�*��ŎW	R����P�e�F\�Q��r̩a@�� @j�a��eQ?i�m���n8�&j]��Y��+!�&tlX�ૐ	��� v�8}R��!���	�z�&����c�p�c�oGUٓ&O-Ĉ5m��(�Q�b�#ը�!��1��OL�);�&%`$��'W`\��'�JpRUE:"GX"�!@�_�(�����A*��"eSd�O�([�k��Dx�h��!g�����I�^�ڠy欟:e������$D:#Ni��i�uB�7@ڃ�y2��%#~Xq�Y	{�~�[�\+��Qb �����O�"~�	�7�x��{��dA�Z��|C�I�z*�h"�M�
��H%C�5&2˓I,`c5lO\u��IH�h%jSǁ�AM>{u"O�@	�B �BF1c��##�87"O�@�%��/��Ӏ�(CR"O��CC��G�d�@���V=���"OD��*�,@A��UO	�+^DA��"O|� �!W��`	�ΞpC�B�"O& �s��'C���3pÍ� ��I�"O���p΍8kI��y�%M�J��I�"O�i��Uy�!�vi;�0�B�"O���Ǩ� ��iR�)�[U�Yr�"O��� %��Ra
#fʒC�hi��"O��¢nUH��Z�%	_�R ڦ"O4<��KI�]�N���ܛta����"O�hP�c��<��c]�_�%#�"O�e"e�6.�U��9/<��q"O&�
�h��2@8\'>�B%"OZ(K��ħY@���d S�.'�a)�"O:P��"�,f#и����(���"O, ��Ȇ<G��`��/T����D"OT�A��r`kql��O�2 �"OLD���%I�H1��aƧZ�����"O�����O@�m Ǡ��AS$�+V"O��`6���� ����&@8��a"O.�3p���$g���CY�ycP-�"O`䩀�H�Kj���኶z��'"O��U�ܒKf���K[���CV"O܀�`T0�|x)�W�
�"O� x{�"̈�H�c��Y�"�13"O�H�-!��!�m4�f!�!"O�|ի��`���XĖHٚe��"OX��p'E�;�@�Q2@�.?��l�!"O�-�Ixi��:0ԃ
�nD�"O��+Qm�&w�p��_���� "O�ђ�f�7�F�
%�{�pJ�"O<�($�F�-n!��cL|TJ��"O�q�tE½0�p�z �/G�5"�"Ov�C ���
$�]r���F,Hap�"O��km�FWBD� ,�34��#"O&1`�kH?��]��J(9��)7"O$�F Y�O�n-◀��u�,�8�"ON�ʂ'D(	���U�F�t�1��"O�Iz��?���i�Bi�N�@�"O��䮕��M0�R�e��,�7�7D�DC� �4���3��)<�1���4D�(�u�O�I|ѐÄvz�	D%1D���G���d��NT�HT!W�,D��yAՎl�A'��}0�@�'D���/���@�
,Ej Z�H"D�L�������WŃ�Q>a�Ӏ D�RE@\�q�(��LL���	#=D�L�lF�j�&t�K�<D�U���8<O$p	$�4�����Y��e�`LX�R1L9LH��S�B�V�G%2I���3?�4��O2l��߫f}a�'k���b'˭J]M򃠕�uN2��
ڵDQ�_ed��μ`=
�;��  �yB��&n��+�Cо
�>�G��y��ъ]ʨ��F�H&�h�Fh<��>�f(˼s���` 3d��1��-Մq���Y�D�j cFL�:�P˓9®1 ���1|H�"<��k=2�xɪ5M67R��R,�s�'��u�e-^�d�j�ڦ��*_|I9���k���
|����լ'�z�MN;gx�}��G~RZ��d�Ǡ���I�/P�9i�lC�j�p�0葮mC����e��>��O����ĉ,W�-I�,C���͖:

x�����Z�҄[��v�<"F�b�Z�q�F�Rt���+4%;p���>�|�p�Ǎ,�JMCR�F/c�\�I�V|�Բ�����&=_�h�Ŏzt|5�'dE�Գ�<%�<dÐKʂ7�^C��(.�V����ЩZ��%@�	1�z��"�'8��U� 1�D4 ��|�{�F�++D��UW��~4��A��O8dʔm̠RN��C+C-.�(FC&O�� j�`��V���Sn��R�HMscA��}Q���޿:��mkU.��p=1$&��F��t3@��4 �=�E
Ba�D+�i	�Ze�����[P�|f	5G��x0�5�5D2v���H�n���:D:�Y�ȓ/������:L� ӈ ���"�p��lI�Jᶐ���ӈ���ܦ)i���P:PJ�`�����E�uw`�CK�;Moԅb��B]`8Jg'&,Oڤ#�H��8���(4�#i�!�D��"q��KF�F3	pt���Iv�-rA��;g`(Ӡ'��&c��4'آw��c&����T����5�B}1
�qa^����S��*I��=9N�.�r4(c�v���ԯ�&��&�@�N���ʁ�z���YAӸm.~}XĪ�^���ʘYy�!ѫ�p����%���^�"@�H�FbI> �mQf&؂i���`��
�l,��;q��ge�1��ߌ'J�h��B�<
�Mi6��k��\��b�*F���ፆ\j�)慉�+,r�m2��2ˏ���g��Fѡt`ӌ+���@�>l��ԝH ���Z=���3v�`���K4՘�A�?	,p�۱cƋ�Jͩe�D!�X�袂ٿ��{��ی^\4QrN�/(џ�2l��l4te@�D�Y�LL�anۯY4�� e	�@���%i%����cȍU�ĠX�遈X�BP��X4��p��
D���U�ǆEَ}��&N.3���a��#k��I��#n�4PY#g\�h��$��03,��A؂6W
�X�'P[��aaG��"�HE��6|&�PU��y,�"a� 5R �p��ҌQ_��I1�-#�PsJR�ف%�̆+�::��eͩC��ܪ!���r�oZ�Ү�q�(О^9�L���up��!͊�QF�����S�C�8�B�ꉍ7V��H���	h4�dӮ���(Ӆ�
BA����&]�'\fH�h�g�q(e�[ "�:��4 *}+1��!�HtTĒ&yb��*�bQ��X��
�4�uǉޘ,����٬c>f��@��ms����֑���ZFc�w��>�'��x�|5�q��F'���.����a�.�%q�n��<�0���W.(��rL�A%����0
��qղiS�z�HD�>LH8�0��T<�<+Ç�+9�0ř��D�&:�� ���hTQf�o����t���<X�eC$
��0T��9x�,Qc�_6>q�*��@��$��'��$1*|�գR%��4(+��<s� �c�Z<*y�@C��3!ˇJ �@��P:Б���7�\�T����y̓<P��&�� ��V��*� \x��F�-[�	���Ԗ!�����%�t�2�>�Xy)��^(z�<�b��(P�%�S��IpO�=]�����`��v(�CSX���_%�$�d����I`H�+p%H̓t`߄I"T� '����R8��azூ���<1e-D�g���*�	��d�����I
V�R�9�H�,S��k�*);��q坟�2�u�'�%��� �]9V�Q_D�p'��p���+#���aT��Dۃs��n:xb2�Ӣ,�"��\c0�5@�4�Ç&9*Ǡ�WG�	*���
7Uj��袩�xrH��R�iy��˧I���y�b˯{��[E0��`�$��F��Eb��gf�sr U�[p��(@hE�Y/��!�f\1$N����P��U"�dc�!� ՜]��x�(�_"� ���4N�2) gGƿ�J�H��Y"9İT��i ut�a��ȟ�]�/�2A�����N
A��c��(�B\�UՊ����$o��{A����	Cu�
)�L@�F�:ӓ#;t�D}s"�%�|��g�><*�K�4^��CQ
F�)t��ІC�8F���S3�]���4(l��@�_+P��h��Z�=ohl����
����¥"�&�*�k�?�6�"(��[%bPlӭt��̡S�/%�&Dڵ �<�B/O�$�P�W�G�֝�?`q2q˷*��d�s�@�a��l������L�M9�XV���;j}*!�˵/��P���A�d��X�qC���^$*�Z�g�|}����\��-���Ġf'�Yh�O^qC�#]C�DT���OU�4�5P8�8�MDLM|��5���C�\U#��B�L ɔDV/Z]�bT(ԶU2�0��D�KFv��w�bE��폩`l��;�具G$�� ��)����Fظ"Z\ҧ������"Y'^�� ���X�����������X�AQkT�=�T�A�+�)�P���R��#�����2�Y�M3��� ���EXG��M!���s�˰�jm�bF�&d��Uha��{6�����(g�pZ6�ۆ��)�M��x̙'�]+(�ؔ�UJL$$�D�Hz�ȑ���^��,ir�,ғpu"Q��*�%��h�E9L��Ig��=��,9��+_��$�X$qv*E���ȑ&��t��P8N��]"''S���2��]�,��̓��9`Gq��((G�5�2�'w�X��n�,$�w'X#o�%@$ggjT����"~u�	�&�i����lM���DO3@�*c�8�r��@���-��^�%@��'�|�C� ��4�3���C`|ق�$Z�]u.�`D���9���D&�,JO����G@�u�CiL�@epź��ZY:�(�@ڇ�?�G'Y8}�n]����(�pvG�|�'v ���9y�~}�F�ß�8�0�G�>��kdf���4�Q�f�0��Al��韰aA���;�f�Z�'D�:�bT72�d��#�)�~	j�4^�P�҆bG�)�jlbeB٭E"����+h-r4�r/�$����/b�9���5��ʰ*T$���k4�P#)�:ą�I��z��$��[D@�P�h��&ڀ�p��4@p�5��e�^�)Bm�|��`�%�BAǈu?a���]0����bN����S@X�n�8UZp�V�}s�ٙ��������lզ�|d�ׇ^@~e!0	�-�LY�щF�~x��E}-��Ph�ǃ�yA ���k��y��_!q>���'6�U�"jx����3�_Ert�r���6)�T�	�,(�.X��
�� 1.u� �[t�>$���iWZ	7 �e��T��*�8�!@��Z��L���e�Z��gG � �h+�CV��ƀ���Ԋ|{ `0��4%7|E�`o�2X���*[2\9�+��G[���u��^��{���]�fxȕ��}ڴ���ƈ���Xs��%q�b<�'��,f�P���5fVnlZ����}߾���FH���|#%�'t�z����PQ���:M�ӌ����\B�ɘJˊ�ҎU&>x��' ���,Y�&�By��سv�ֹ@���D|��	g�Y.%�	7�܈r�$k�G[rr�]�rB��r�g��1G{��� i�
�<8��2Ԩ�$��+a��g����(A���1�,uP�'�\9RԎW��#�J��D�[�\��|K�F+�>�X+�O����]~�� #���RT �Óp^�����;!���Pg�+���d��	x�͇=�\-x��,[N\HfN�Z�`��q���BEŇdclU	��Om�0�R��``v�UX�HyPe 7�8)�`�/Ҧ��te�7���8V,OO���1��+HR�Ma#܌a���!�d�?޴���%��3����i%�����UX�T`�{ �Cq��)ΰ@�ł��0�Jf	 G�&T�ҟ̸P��1Lo>!�>))Q0A�5.�\���� ���r��E���'l89"�P�(*] a��~�e���q"�.��i��GU
(YX,JF�޲+X�2���NxR����Ţe��	�Qb�.��a��g�
)[Z �;���3�L=D�ht�Љm�t���0�ȑ���%Fz���M���O�-W�;��:@+V*f���$��qt��˱�Z,�x�2��?M��t�[�
��W�a�ԋ�o��u}&��`��ʝ����9S�P�nӬ�
��dU-q��)�T��\�����L<d 9ĕ�S�Ö��>z,��ّ�F�!CX����m���g"3|)b�5���ɒt�vN����8xu����
=8�(��7צg��S��?S��Ջ�̓�������B(mc�c
��b��3�0H~�S4s4�pR�����?E��'P!4��"EJ3d�\
.�&YB^>��SO� ��2�Ŗz�:#�b 8��O�"Ub�wST��P_(������B�1�'���r1�%a���hUJi�'��#���'g(�q�HM����;u��Er�B&S�����	�M���h[�d/�i:�47�>�'B�[D�ӎH�yö��=�p&�t�>倌�D�ET�st�����c҄�u��*CdI2U����Hg�O%�ܑjTa�&P�8(���*ڃ�ɡu�YȵY��(c����(� `U hҰ	� �.�&����ӯ7	>u��e͗X�TL
H,�R��s١F�}����Dǟ�8���1S�d�	�xBr�aa�#	��S�O!hd �J�0*(�C��3��ZT��V���K�"18wD���/FpL@�����i�!�1�;/�����)~X@1�d�t�v��O���B@���<Q������d��pWP`�$˽D��uY1�	)H<rUY�M���m���´�����'�RP9�	T�j1��f�,f�!���j�"�匫^3��J�TX!B���8�_�m�C�a�^�1Ė	���P�Q�>�"��D�m�(�±�F�MQ ��4�F^�'��TXs)��4��#m^$_:p�p7iˆ0�<��A«<���y1��5I��P��*/]H�s D�`���  �ݚ��S�4� ᧮_�CV6C���,hy:�s�*@�{��=0$��2�өE􉣟w{�uk��ք*'��r�ɪr�V���'�^<�ul�6G� ������$����!�Z�|es�����Y�+]-(�-�l�4B����� 8��t.R�>��m��,	
n��It�'��}�,j���y4샨N�lux�غ0!�+���Y��kֆ���k��ѹ����ד6�fLa�Yk��E�r��|$����M�q��`X��7�A���uU��`�H��4�dL1��F�aÆ(�dkت@V� 瀝t�<A�C��KN����"�ܥ�v���&=N,���;H*(z�)+h���JL�ӻU����w�h��VEP�R����sě;XQ�X O>�c�;�E�I�=����c�%1�u�ƦS<?��mY��ߛ=6b�IrcǦ}�ק:,/��C�'ƭ?Mh��`���di�nߚ?2�%C6 ����uV�Q���2e�Q� � �8;YЁ	 ���d��={v.�/O�  ��
%`<��0��E�����T�K�0��D*�cʌkX��N.�����R�i>Ia��D�F>�a����|��3?9����)��/Y�*��h�� �4�!��^�l�i��x�敩�Q�=��96`�$�~���l�{���#kߑ`�@r �O?���^�6X��Q�(k)�p¦(św"�Q(s �����&�O'k�J�Y�_�2T��q���	ڠd�[ 	�!��a۷I�J�ǧV�o��ضU�Ԃ�?:�|lX+�qO�	�p.�Qk\�d�M�"����G��my�F��H�,T��I�`l��� �TfF����C�O�,��!F���Q��0;F�jB�W%<� R�DY�o"02���)�(OJ�J2��':�2dD�0i2bS�J'Q6r����G/:��Ȼ�C?*�XB�#�(j��S�ȾO<���Ү$P6v�����/8������˿��d���=cD=Rd��D�Z���c����;7���2s!��?��h��g*B��#(��2nX���5_|���M0 �	1,�J�li���ؐ2���cS�d�jV�z��	���O�Z�eK�xa�h� �H0b5���P�O�@P��g&�<k��M	��<"D�ʝ|f�d� ���`3����:�<M�f8xs�4#f��13�H�o�_jp��G�N1flPa㣛�P�����S�\o���_D�^�@��,dEb=(��Y���y`Tn�2]*�
��� 7Ê���ބ@�P�`��R�"S�d�^��� Ș\=�q	`ɚ�%�����)3���#�W�'�����FLx`&!�B��Њ]�M�^1r�m�
$�y�q �.��A���T!R��ұ0�! �,��m�t"T��8�!��ӻ[��5�^�v2���cmS_���'�`���'-��YG�;%6��un�_~�M�Bks����Q��7H����YZH\�����(�(S��ӄa�%ĄY�*�q�#��E?i@���?G�TbFg�	T�Q��:a���SdH$esF���%��'*ީ+����;@�Dzf7��I�"]��[��_p�^���f^�khѤE�<G��	)7�.a�����AHS�կ���O�$"F�ч�4u��6D�N�P*��b�iX��S&M��pc�D1�,2v��0}�\w��Sᬃ� ���*�HSg𨅀��Ղ�T��0
S�~�$�XF�H�'��(�J�Ħ��W��gh�ab��\�K�2� �������_'��ٛ���0E�������^g�E`���M�6�`dX�~�响#�ⅈ'͆�ܠ8`t��M9v�?�7b^�} |� Q�{0��U�+xڐh��F.u�P�/D�
Wȹ��I7L�t�����&�H4�P��;�H���iHTHx��W3qb�B��Ë>J�'g�̈��ǟ�Z M	�	��>Mr�*�z�)��J��������Y���.3�`@�0�_8|������DӟH�R�AV+U� K��cS�L�	�d�V����Tz�MG�;�1����	v�ݨ�'Ѳ�pS	�'^���#��OB:��B+��q��^7
�`k玪M��p�~�R���2R�S7z�t�
��Tx�<bA�]�ֽB��.Y�^|��ʴ! ��e�Uʼ�O?��ń&��p���ܠ�Z�+�!�dJH�&��r�\(�nU!
�4l��5r[�ĲE�':QJ��5�a��
Ue�L�	�' 8;�i�7m��q�Ռ�-D���:�'�bm1�%^�Z��;�C��U��P�'���ZGg�0�dBX4F���'��`��8d.X�Kƾ_*�;�'a:�zvJ�@ʎy[E�E�Q�Pi�	�'�$-��nȷ�q����Nբ��	�'c���'�ޛS4�]�F���8��[	�'�j�0��	e*�eAvmV
DĜM��' �A�5n�9J�D�ҀY)U��5��'%Y;R*@5p��V�K���'5*q�Ɓ��x���.N��{�'ru����>93�+��,+ T0�'Q���dW�~V��S��$��,H�'�<D��E��1��YӢ�\�w3��[�'��X��k�L�1ė�cn�� �'w�)�.<a�Ը�VꉿQ��;�'e���@�X�%֤HUŔ:Rܨ��	�'�u�M�4<��`��ױJ�P�	�'���?rƜJR&�)Eܜ�	�'Y$�[1��$;��a�Q�X�?�xH�'� �'%�$|�q��Հ&����'���{C�:7L*�*E?�^�
��� �=sd�7]!C�C��L�e"O��K�˙�d!���UJ�
'L*��""O�1R��ث�vY��AL#0��"O.-�E�޹x.����̚='�i��"OJL��A*_9f�!�sL��W"O<	c�D"�d�kݬR�.ub"O�չt䐼X�Q��:0�iٵ9O��@a����{�[Z������8W<6�p�͏�6Ÿ�D��]"�{�CC�w��l�<%>i�a!� ]�6@�'C��% w�Z����� �J4̙;4)��M���=��(G�ƹ�0|Z�ܙ¤%: H��t��SK��M3#c�4Dm��s{h���_y�O������X���3�J�|���	���L[r���Ό�3�V���Ȏ�0|b�ӿ�bDɳ۱M�82#��F�2�c�<ڲ��ȣ!2�ͅᓤ |RXs`�¥r�MZD�����L�ŵG(X"'Θ$E�ʜ�k-����Ռ�9f��m�7=�����\�J�K�A��x�C�Y>*�a����	{�i��S��(Y7LRT�2���߆H�:���O��ᓙF�|�+��&An�@���a���=Y�0�?牠^�@5�׭d��Pg�ٶ`�jO�ñ�H�<�b���D�F�d��-P�lUBeI҉()5�Ec�(WX�
�4J�.M2�'5du���(�'����=��(����l�,Ĺ�D^,�?Ѳ�����f�[I��R
�',�jpR!�R>�d��hM�pF�����O(�[!lV�Z���	M�'���>S�ͻ��֦^\@�Z0�<,�R6 9y�T�ҬO^�ˢ*%�'�N�]Jt�͉ra�u�Д��>gx!�Tg�>y��� 0���0��OX29�B�F3O�����V|�O��s�$�0O�����h�OY07�@<�����u��	�<E�@�K�<>�P���p���)�'W��c�f�� �7lO�Tl*��geɻa14U`��M��҆�I>�M�_�E��X5Barh�d%B!p�0���?)�JW ��)�5 ���8�̀	THBEI&�.� \P�Ο�H�d#��"�O#�DcddU�+��[$mQ#[D��#B���n��s�MS��Vy ��j����f*�9p����J�i'�-��'�����^ ,N��fB�r�ϥOu*jE��JJoB�d 7�Q
	mV��'`�1���8F(&�Q��9OY����	����Z�3|��	�"O�i��O	�d̜���0T�<�"O&��7�N{9J1��m�gm.�"Oz��F+���j��*d�0Ӈ"O�@3�	uQ���;0ǂ�8P"Of�
��@OZ�T��J�´"O`���@�M��BR�+�Y��"OĈ�%h�xpi���Ă�d�"O�-�`D-��|Qf@J�^�x"O2*2��#A�̼z�	�u(i��"O�(��KƉ>RxEP�ko�a�Q"O H��N8�Ȅ�u)WsQp�Q&"O(�K��D�.���H�t�4��"O}I�o�?i/�Y˒���j�A�"OF����
Z:x��q�M�p���6"On<�u�JJ�`��R�H��$�� "O���@��Li���O]$(.t�&"O@D��l�-d��ٸ�`��?/�+�"O6�`��c2��r2��7(t��%"O��w.̉]����n��U�J�"O��9���5s����4-��f8�I
s"O,D�Մ��Qj�q�,WI�*���"OMj� *3?�㦡�M�̠{�"O�i�g�{@�%kg D�HP�"O��pAcؖ*Ұ�xRO8�&2G"O�P���
?�:��1X&f!��"O����#ަ81VA3E��0�&�
�"O���� ��8
���0�M���2%"O�c�P;>�6,����~��Y)�"O��Sff�=_�FK���@�V�2""OZP�di��
:x�8��-^N|��"O�9sfLU�l982DÃ4H���"O:�k��֕<jĔb��ǄJ߸��u"O恁���$K>�=[功�~���c"O� T�Ұ�K2C(�Q�	�e���(`"O��"�lC3	�A ��Jg.4��"Ox��&��N���@���^t5Q"O&��T�-�h|��AĝK"Vٴ"O���b�U��pӳ�ʳ	�I�"O8A2�Z<-1� ��`�5�U"O4��!�X8>��Y%ݛ%1��8�"O�M���	�� x�U;m�a"Oƅ�BџX~+
� 4	~��3"O�!��B	m��B��z�t�s"O��y�lŗ'6ت3oʄJ`F�0!"O&�����6Q�`�^XWT��"O.�+@a� 4�]�SM�:H0-�U"O��"%��6`�e���(K���"O���*�O����r��{��L��"O>�B뚹�q�q�K
j�졩c"O�RB��3����֫Fs���"O&� �Y�b����t'ىP��ə�"O����D���<��f^u{�(RE"O��	sP�/��ePr�����D"O&���*��j��l��$i��IھAc!�$��\��Eb ������m!��J:
X�<��	����b��ȯQ!�8S@��J6(ɐ@h@ �'�Ac6!�D֙lb�1�"͘�	�ry:���("!�Ď"r����f�r��i!�䊘�\9�W!:�R|��!�$l�!��Q�nYn�:�)�z���z� E�!���Jr�1�k�W�f|b��۝v�!������!�銀j���:Vn'�!�È�ʬ��X69*"N�
!��+�"�*7���<����O�2b!�dͣ_d81���V�0i:�oT�/!�D�A�@iyeKȨ1���)þ>!�d�n �NЛ 'b��d��{�!�$�='��Zg�]<�pt: 	�2�!���|�&�#�D�Zn�c�O"V�!�B�0e4��(�^Z��#���' �!�˰K��]�?X�Xf`Ǭy	!�NQ��,�)�nqR�«+�!�E�3C�H	�͌��h�ĥX�f&!򄄟c�aѠH�=.��ADT!򤋓}�
�b�E�����d��!-!�
8d۔=���#��c��S>`!��Q.���C�S�	ᜉ�$f�!�J��;��S�����`"�z"!�Q�aԄ)RC�@#�`U�W,O��!�d�<v�4]a�@�[<��p��� w�!�8$|(��
�d9б�@~!�� ¾`k� �6Z�
=#ȹ�!���!A��oL��+�/K����'�4ŋ�Ė8����f.ȭ�i�'������Y��
	F9� ��'���Y�(֕�(@��� �>!�9	�'g:���B�9�bQ�Dk5
��lx�'0`�I�-W9S�Xq���D\5��'�:�c�Q'!���� �ؔL��%p	�'Q��2��#A�(�F�ːW���r�'� "�)�T��4�T��M���	�'�v��!C��6-��b�"R�K���
�'hx|�T�jġ� �·U��A	�'�lzV���viF%����r�	�'W,�����!d[G�
pf�y�'`BP��\�W��f!�ؙJ��� ؃�"^�����K�*zjܰ"O6�{���vL�ö��
R0!�"Oԭ�) ]<Pi�f�hj���"O�C��A&i&�҅�S��ɓ�"O$�h�-�Te�ҥϢa�M��"ON�`D��=�&��t1,���"OP�g��6~.�}�b��5NJ���"O|h��l�^D 5�G�����S�"O�y�����m� �I����"O|�a5����6�s]H�"On��֤y���vf�,m���%"O
5I��]2E |B�ޔ+Vnl�W"O�,p����S� ��a۞_>��@�"O�U�N����Q�A+d0�e�3"O�斑q7jxtA�~wH{�"O�u9u��3���A�@I��c"O�1H&��c& ����97�2��"Oڸ!��X���!��+u�!��"Oʵ�t�ەN�=B��P:>�R"O A����42�u2��Q-$10��"O��@�	�vY�P ��R6|�a@�"O^���T-M~����,ͮ8�v�C"O�5�`dGN8t �޷TC����"OBlB��� �\H�a�ɡ+MvԳ"O ����8+�H��bgǁ疴I�"O���˴f��Բ��	�.��"O���gX%7�"|����>��ՉW"Or1���M�ԜxF O"&{���%"O��C���Yd������$�$�g"Oy1 %w���Q�-�"WR�Ra"OBa��;h��ip'׏pLx`�"O0U��&˩;Fܲ#�B�>/��D"OB��L�z�8pe-P�}z���"O$hҗ�	���uaDQ�z��!�d"O4�Q�-��Q�X}h��ԉ*^ܨ��"O@���ҫn���eޒ%�|�Y%"O��;��N�r�Nɨ ��t��ɲ""O�PB����M*���%�"%�G�,D����^�5���C��?�(����)D�pJ3�ՒX�xH�Ȑ4��}ï)D��"���=d(P]���Y/V��U�&D�X!牨O*$�j��D�*ef�!��"���%l�$Ŷ}S�Ա!�Ĝ�sx ��5�xE�7� 6�!��7$������>{(�PX�!��Ћj���Ì�9,q�h��L��!��,���� ��	�2�z��J�K�!�dE?8�r-�Ť�6e��a#P!̀8�!��/	��`��P �m�3aD
"�!�Q8Ȟ��^>�j�O?Ne!���N����c���p𰤘
(�!�d�>t�`jg�739�y�lF�|�!�$�S��@��!N
G�y3P��0e�!�X><8�YL�9)2�C�)N6D�!�D\6�Z�
��N�c������$f�!��z( IQ,�b�5�/�Xo!���� 	� Ǉ�b�8�Q�d�!�Dͳ���+����DN*c�!�Éy�~��oX%:��Q�N# �!�Dŕ^~T��blV�;����� ւ0!򤐒A����FZ�i�R���`�7 !�>v��d�/�~L{���-O�!�D�6��Z�GPU��+�م^�!�$ۗ(в����H�ShD���>!�� � `�
VT��Ա��RZ�έҷ"O1!�4�dL)��I���DB"OF0h���9Ѻ��q���,�r9˖"O��HWA��~�ܸc 92�(�"O
�:��*<,AS*�7����w"O �j"`W[�Kթ�AP5y�"O`�ڳ���R��]
��� X�֔�'"O���e�o��)�RƞS{PA"O�,xQ	K|���AO�:gvtp�"O�y*���9�|5��"dm���1"OV�I��� k�X���P�R^�A`"O�T"�cе4��#��� /N���$"O��iٗ"����"�ɓG.�M�w"O��f��^Jx���@�&����"O.�����>0�92������"O@90v�֑[p��,|�\A�"O�8dD[�T�p7Q�)#P�3W�2D�Pq�@�I�V�B�l
�-jz �o2D�8ʤ��c�T��aL?F�@Dc�'$D���k�N��� %j�  ���/D���bف$�
�K	"D�hZ�.D�`E	K�c@v�����V�bp�*D�p�r���W�hu8���nQ��/)D�0ku�W��e��iQ�?�VM�S�:D��d��"�9����B�@E� �5D���%�5r�� �.4)�q���2D�8�2�+)l�l�����Pݰ�d3D������$sC������'s���0D�Цg�Yp�!�R�;�dP`�G4D� j��m�H��AK���|���3D���F�0�Z*��9�b�L3D��I��N�G(Q�蜾���E�1D�l�G�l@б�aY�I�qǇ+D��� ��WD^�wGٕ){�T!�i+D�T��
¿9� U0�F� ���)D��rs$˩b�2��R���E/(D��Z�   ��   �  �      (*  u5  A  �L  �W  �^  #i  s  Gy  �  �  ,�  p�  ט  A�  ��  ��  >�  ��  ¾  �  I�  ��  ��  ��  H�  ��  ^�  I�  � �  � l! �' �- �.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i���$�>Q��ۑeK,āc��/:TR	еO�'���,�r@k�� c�x�x�iY+bB䉇KxHA�ׄӏO�jM�6��TK��	��'"�>�Ɍ[���zA&��D�Hq�2BQ<S?P̐�'��L)��?z�(�4[0�`��ٴ8!!�4��'�
*m�������q)�{��d��\���䚀r�V�+�;<��{��)Z��K���ѲBKG�,�4��� @�<��B_y�NtCD៙n���S��զqE{���i����j� ��i�1B\�#
ϓ�O�zP@C!p��2�"��yv>(��3O�E{��I;Z7��@'�4r}c�N�W<!��6
�\������椚�2.�P<">�J>yPmS�e�f��N�(3�v q4��H��p=�!`�=Ԝ�J9$���� ]��hO�'
Cn�HRJ��Y<��'A����mM(<�p��=�q��ǹh�����Z�<	���y�>�1�L�8`�B W�<�ЄJ�H�m2w#��x-�%��P�<�ތ��̀�ʘ.f� TO�N�<�#�	n��(�%�֢$Xd���$�"�hO?牝��A4'��Hh;@�*`u�C�	"���(P�"xyv�[J�Db��n~���O�Н(���O�^,
c�Z{��AI���dE'�2x�%
H�ض�ʵ����'?���'��x���7:R��g�'Kn`��d��?q�'ȰY쎄 ��G��n`��'ή����D�p�!Q�P�v4� �'�H�b3�Țe ApQ�\��{5"O�M3`+�`� � �^�4��g��Ȅ�ɖ;��2�.�2ye<Lڔ̒�7sF��d!}��<-.YS�%Ԁ	��l��L��y"��!!X0�Tc[O�2e0�N@��y"G�:?���D��I���RD��y�hHP�m��ȈF��Y�#E��y2���}qx�b��R�����'��?�����1Vj<CƦ��?��0�2,7D�dhAAڒ ��@I����Nx�	D�3D��9��4WS�ț���	2���A1D�� �YCu���~ۘ�!��t���zA�'�!�d�j$�8��1���c��sp!�$���`���ݙ^�&P�&IҮ,T!�%d��]��a
R�J����[�QF!�dZG ����]!���&@�>!�V?�N�؅	���H�-��O��8�S�Oavu��䎘���N2b���8�'-����<2��:�'��M�~("�O���I��<����O�7k�ڔ��0���>A�`ٽ����]�c��p�uj�ޟH���vx���F��:|ʢk�rΔA��F~���]8�E�C��c�P�*�'��
^C���i���9�A��T �~��)ڧ&�q����1��P�W,�4F����ȓ2�\LA`�W��<ё$O�<��)���hO�>�xe`��5���s�H�s��p�6D�\�r�H�<��u��؁B��g4?ɫO����!V���sЖ�hA��:��~�T�l2��Az�y��'ա77 ��%F0�IA�����&��@�y�&�U$j{�dA�d/D�P����� <Y��(TZ���A�?�IS�az�h],8T"(A D�?e�Y�B)�M����s��x{�f^&�~�*���?Z�ZY��"O�X�T�L�.AV�ZG�Α����1OH���df���5K@��B��Z�k!�$/Ei�M;�䂅}��0XUfܢ_!!����AsE�e����߅!�ѵ
]f�ȕl����3/�!�e�V�
�M
+����B�"�!��ǟHH4Pɱ@D�d���QQ@�y!�Ȗy�~��VA�tI�'mӳ>f!���1L�0a��3J��(���k�!�E 1<�v�τW0(��ѳV�!��$pӀ�b#��K�pl�-���!��%~�H3�M�&�N� Q��I�!�D�"Ap�<i��+p��aaqO@#\�!��³m��x�pk�.vV�)���x�!�d��00b���J=nY����U0�!��6C���l� �� ���$�!�d��"-�ixk�<���ʅ��+	�!�d���̺��
X�����CJ�"}!�d��G�U��}����-�!���o{�e�$]�d���1�wb!�� ��2�2R�`D�m;�]-@_!�Ę�D~�1�t$Ϋ �>�{�Ãw[!����Mp��>#�
<i2%°l�!�����`��7�$0� ��2t�!�ć���2*�B�l}"� �,�!��=F��n��Ҷ׊F�!�$ӽSq6�x�%%au|�o\/X�!���
s�� X�nQ�� ��-�#!�D��;.��q�#�4����"W!!��͏��+S�P�|��кBQ%R7!�d�����A�m�{�ݻ`��&!��rC��C"J�j^6ps��6`6!��@���5 )�����K�y�!�Dޙr*���&�m}h�����!
�!�-u��ar�[5:>���d�D$]	!򤘩~��l��`�!����7��!�!��~�8á,I�x(q�G#�!�D�y�hcB�ޅc��	b3 �4�!�$=�4�x��$�B�N-i�!�D�E�!���E����2�R�7�!�dB� ]Ri��GC�4 UB��K�h�!�� ��aY�X����H5� �10"O���A,M�x�x�O��2�v���"O��W�	-m���^i�N�2"O �bQȃcY˃��gf�x�"O����T*�^�5�`T� �'��'or�'}�'��'	��'@&�y�@8� U�
O��N���'8"�'���'o��'�R�'��'jMe�L�0��o��K[�� ��'���'���'f��'r��'W�'���N�.@~��p�6�#V�'��'���'��'��'d��'��t�$��hk� K���-~Pሳ�'U�'���'"�'_�'R�'g.�B�_�^��A��49�ae�'��'�R�'�b�'��'*�'���Ӽ�ⱡw�k��S�'_b�'�b�'u��'�R�'FB�'jV�1!N�vw��I6��+��lSd�'���'c�'S��'S��'���'�V ��Dޮ�B��0�̈O�e��'���'x"�'�"�'R�'��'������.-np
�G+Q���2�' �'c��'�R�';��'���'.d�P��C�k�Y�0�*$�"3�'3��'xb�'�b�'$R�'���'=����"
�{r�@)�ǎ%I~A���'2��'b��'Or�'d��'C"�'<�e�B�K�%���M 2 � 1Q�'���'�R�'"��'M"�m�����OR��DR&��q��#0Pt�u'Mxy��'��)�3?iU�i6�RE�!)0b@��EL�`r��7� �����Ӧ��?��<��O�a05d �|���PA����˞����	%��l�m~�;��Q��]��߿:U�r-S9l��q���G�1O��$�<���i��
Þ�Җ�ބ<�4rWmǚo��oډ^��b�(��f��y���0b+��%@�&�I�5/�7:��'g�>�|:1S �M#�'d6=jU�ǻ�`�h�愙	����'��$�Ο����i>��I�8�<!��v�1z@"ߝ� �SyҘ|2�lӰ̳�D�_2�AR�$J
IH��0�U�چ�!�OF�$�Ob�i}R�ƌD�jx�����H�T�^����ObP�fnA=>a1�bT���>ah��Q�P���������#L6LJ˓��$�O?�	�	T��Ҡ�5{�
f(��0V��=�MC@|~��g����S#6���u��1f3�I���R.(���������R���1�'��iJ�?=8g�W�~d3S�[$n�����C��'��i>Q���`�	�\��(Y(��!M�	BS�Tk���'m�7���2��O@�d%�)�O�D;d�=uej�7�J7Z5��
}R�'��O1��8���8���8��I�+�|�Q��p������<����=�����䓖�Ԩ��D�H�8�>�Ktϒ'Lza|"Mt�|p���O��2D�	�L�2{GMK�Z���ڇ��O^�nZe�!���Ο�i�rH�*F�|!�fMՂ(ꎉ�4�L(o�@ToZU~2�Ӹ3T��'��'��K�O�+��
�@> ���h��<Y���?���?Q���?����	�:@�R(��w�+�o�;t�2�'�"��O �JϟؐlZT�	ZìaA@탐&��5AG����c�4��ry�Nʲț���U��r#nx��J���a� �+��9g�'�Ԅ&��'�r�'���'(diq��_4�P��
ɿA�T����'"R��b�4k�.<���?����iN�	��8�0�D�	
���A !�$�O��'�2�'Cɧ����a�ǳcw |��HXOLi���4�M[4��^`D��|���Ol�YK>!��ہ"��yY�DY5�	��b�?����?����?�|,O��lZc۪ � �ҷX���{�d�+B��떉
�x���M#�2�>	��)�p4���J���#;�Ȉ�.OB��gm���GS4�P	���`�)OP! ��@���P��kG�z T���>O��?9���?Y���?����� ����X0�	<|�8�P��l�!!f�0�	<�I@�S�!�����DY�\���M�Q�P �(���?A���S�'��l�ٴ�y���1���$�!Q������y2ᐢC�������4���ě�/^T�X�H�8I%���b��7+v��D�O*��Oʓkb�V`R4S2�'��C¨4S�L�d����[��Ȅd?�Ol��'��'��'���@���?_ �� ��yt�k�O�@�@�نW��g�阆�?�g��OH��%���"y�H;c@I�+�H�g-�O2���O��$�Ot�}
��nuX�+	�b�:��QA��K_�+�B��V��7:b�'�x6�0�i��Cc���k��h��d}�1�5�u���Iߟ�	�7��uoZ{~R,Yl|�/������@�F�h�f��,���%�|�V��Sҟ��Iߟ��I��P� �ҏT�m��4MP�c��R}yb�d� �p�O����O0����Ā�#�$����^�;�`v䆚�֭�'4���̉�Jm6�
�g�`Ū�.֋!B*hXrmئb�>�X/����O�a�J>�(O�A(��,<T�fm�J1R 'L�O��$�O:�D�O�	�<�"�i*����'vd�J4'[�R5ڵN�.�~ECu�'��7�?�ɟ��d�O�d�O���ʥ[*T��IB�~��id@~V�6m<?a��`}v��7���� �=�vP�jTH���(�Y���S?O���O����O��$�O�?-�`!��9�����^��F�ӟ��	�� ��4K_���'�?	�i��'����ʶY7Б���+6 ����|��'��O�ֱi�I;|$�@�����P��6 �Qؔ"sŇ!?Y��>���<���?���?yGF%�&,@����%7MAcX �?�����ݦyHԇܟ���џ��O�4)� ��</�Kƭ��!@z�1�O���'�"�'
ɧ���,XκA˂ ��&�ZA��"ۑx1J�R�V4{2�:2��<ͧS�������ڦ$`�H�	(=�}z-Q�"������?q���?��Ş���abe�݂l�Gɐ�j�4�aG�l �5����0��4���?�P]�@��r�b��/�K�<�R��H��m�	��(Z�$ ͦ��'������c
)OR�igb� r��:���^/D��G=O.��?��?����?�����iǗ_�>� �ϝ"Y��%rf�S�Z��dl�	����I��\��O���ā���Sc`]uE,$qDBӧN���K��9�?Q���T+��M'��0O:4�w�Z?n�I9�b#S���U0O��S���?�n9��<Q��?a`�1jJdh�UH��E�.h� ���?����?!����æP�l�� ��şx{Wi&=ܢE�3$�	m}`�Z�Cw��#��	ƟD��K�	�h��|q�,��hH!c�:.��Y&Ɖ���%^\���|R�B�O�����4p]�6G$g��D�1�)y�̆ȓ!~�a2#J1�M&Wcj$x������S�&'��'��6- �i�݁��UUlPåm"kc8ف7����	՟(�I� l%l�Q~���Nb��'h�ś*{�.��C%>l�;K>�-O����O����OB�$�O�l�V��B�>i�0U�?�yQ�O�<�Ʊi�d�`��'U"�'��OT*Ѕvv�ʇR�,w�5�CQ�jMX��?����ŞP�f�! ����b¨[���Y��,=+*O
��ğ��?	�!��<���P)�ı-��#U���#
Ò�?����?1���?ͧ��d�Ħ�KVG��8 bA���:܂Ā^5g�,�Ukb� �ٴ��'%6��?A��?A3lG�T�AM;6y��i�!A��Ma¾i�	#'ڜ���}x �#w���!d�#G��jm���	5W��BUb�=dHp��˙s��D�I�X�I�M{§YW�t�j�"�OH����
1,D�`�����"}���4���O"�4� ���}��R�n񻦤كN�Hyk���R��á��cK��	I��pyR�'���'�2�T3u�8p����L���f��1'dB�'��Ɋ�M���Ѻ���O�ʧ
�2�YF�&WӖ�"A&���\8�'C���?�����S�$���5]�	1v���'��J�&L��Y㡜/O���!�O�I9�?CJ#�dM��0`%�_�juP�c@�� ���O����O8��ɳ<�c�iF��P�JX�$��R��0Ұ50c�GR�'47�:�I�����OPy�%���6�#�I��+D)n��d�O0�#"�r�^�t<��z`/����O�Z�:�(	-b�(tI��E����'��埀�I�����ϟ���Y�ԃS�R��tS��9ɠ��Q,'p�7�NH����O��'���OPnzޕ�d�'"Z�x�'�.,�� !��C�p�	I�)�:6=�l�<q��R*>��fǀ<��ن^�<�C�ˀft�������d�O����Eh�Q?f�0�A��=��$�O��D�O��no��ҕ3q����<#���&A�H��eIձ<s�1e�r��Kk�������s�	'#4[r��><D��׎ӚY��t}$�r��O��Ms��t�G_?��'����Gʊ|�����Bۨv�=����?1���?Q��h��.Wr�p�TKЋQ~p׋ڑj]�������V5:��'�6�$���O�N6y��`����!f1�}�E)X�d�O��d�O"<� ~���}��Q��G�?P&^ ���C�^*�eR5E�S�Ry��'�b�'m��'iR�K8`�(P{��	A8�s�D���	��Mk��ӝ�?9���?�N~2��$иɹ�O��h B����#�T}r�'���|���⋊;��H3%�L�@��`�ܣ0���+@N������oaP]�iM��OZ˓��P{
ĸ���Sb��<��K(O���O��4�P˓���Y�v,�P�ym,��
�l���g�=lO�(e�X㟄!�Oh���O����������|�Ճ��J�Gwm��I���+�vݙp��8�>a�]yvvH����[� yQÊ�d���ԟ���֟���˟��	S��f{%�'�+&D9�p�Y�
��mK��?��,a�"�(����'�6�+��ɝ���6K�2�v�`���>{�1O����<i&�/�M��O�܉��������W�Y�I�� �@�5/D���{U�O
ʓ��'xv}:�c��;����3�O8e#�ˈ��ЦA2&�Hϟ�������O���`G_�X{�	�"��4t���O,]�'{"�'tɧ��� 5e�"���D�X��3��&�BZ
)���ī��4�.a���ؒO�5;IS/�ʡ��o�'v��Oh-n71O��k;��)�E��)-j��˗��ϟ(�Ɋ�MS�b̷>��y��(KqA�#>$�a[�i� f`jx����?�e��(�MK�OT\P�M���DX�� �-ڑ��G00|�L ��Pb�7O�ʓ�?����?���?����IX �5v���p�Hi&A�Bvo�y�̅�����r�S韐C���ӷe�9�hY8���=�����E�?�����S�':�
�	�4�y�j��@^081�兪{Ac
��y�3HZ���4��'N�{y�L�!ky�����r�04��GF��0<��iuf�)w�'~2�'�4U��D�|�pfC�;����Ě}}��'�B�|�`�Rb�G�,M����֬��$��y��y��s�t%?)��O��s2nqX (I�d
`�Q/՛�0��O��D�O��#ڧ�?�u�1ц)��7Z� ��5$��?�s�i@N���'��Em����]�%�ԅ��Ƀi�d� CCT�k?*�I�<��̟�����ʦ�'2�����N��۶WT9�`b�	�D�	
Σ�䓈���O �$�O\���O��$�<M�\�i��Ì'$�B�Ƃ�$2˓)u�&�7��'������'�r$��0%���:c�'.fm�F��>)��?9H>�|bAf�2$�iᷨԔ^���,�>���C"\l~X�7k��ɺX��'h�	�kp�zVř>$�Q�˩h�������՟��i>�'�6�"���DՁG��1gAY��"y�2�UT�V�EȦ1�?)�P�D�I˟���K���i�bR,xڎ�k�׋G���J�¦��'-q ��?��}"�;fYB�Ƃ�|�֜:B#�r�U��?����?!��?���O0�xp��\$/~ܽň�<DAD�'	2�'�d7�ڷ��	�O@oZp�I�*�|��D��i$M9�b�%�|$���	ן�8���oZ^~Zw��0��aZ�$���
*ck"�
�B͆q��	@�	Fy�'���'1Ax���P�"Q8��H�wH,��'?�&�Ms��M��?���?�.�*(�R�Y1=���^�|����P@�Of���O��O�0w"d4y��H�i�ڱh.أ��s'G�'l��h�F� ?�'E�R�ę���(�Ƹ@ �K�=N5�ç�+#�Fԁ��?q��?��Ş����q�'��M�R,:5����i��I?bE��⟀1�4��'�V��?a��� "�x� D] 	�P�u�?�?a���Ԑ�ڴ����,	4U[���.��9�V]؇��4�XY8���4�y\����џ8����������O��`���n�6�B�Ȼw��X���咋n���'|B���'�F7=��a ��7C~lX�PO[ 7L�8��!�O8��'��XA{R6m~�$�v�Y/W x���#7�P8�A`��r�g���)�ġ<�'�?�b Y�s���/d���k���"�?���?����d�Ǧ!�A����4�Iߟ� f�C�D߆q,�#�2e22BI�:k�I۟��?����R��q�r 3B�0���kTy~2��+f<D���)\�O2@���(�ʔ>"��-&��0s��G	ޤ
���'^��'����ꟘJ�m@���c�3`�Is��^���۴N0�%���?YB�it�O�؇s�@�s��=H�����-ڙ-���O�˓8,yܴ���؋1۶���'q������l���$�^�j+Li���'�ľ<����?!��?���'`H�R&�ī>��9���<&�3eW��Qش6y|�A��?y���䧺?9�KQ����rV韔
U�9@b�\%���۟���R�)�S�}s�t����x�	�R��T��#L}�,�'nJ��B$�ޟ��#�|T�x����8M&�1�Ⱦw�x���f�ޟ��Iԟx���py2)uӆ�s!��O� �-՜πy[wb�+kf�@;O�xm�p��Rs������	ПD³�7ȥ�iD�\��-�'�U&+��l�C~�̞=W��<�SOܧɿ��@�f�4A`� �w��z%�D�<i���?���?!��?�����]RW^-�UgJ0���E'=�"�'xB�w�ZL��7����ߦ}&������Zڎ��ê]��X��Z�Iȟ��i>�IЅKĦ�u��@�y�LqK���:Rg�ߘ;I6x�S"^������|R�`�I��L��ş|�7�\#&d�=X��\+f���:��M����IDy�/tӪ��T��O.���Of˧v>� xF@j``��̞f����'9���?i�ʟ�ШP�ϱ#J���U$��	8ؙ9���5�9�D,^���|�$�Or�N>i�@�� O���	�h�T}`!LL7�?���?	���?�|�/O ,m�B�T �ϋ��P�Ճ�?:��p��Oğ��	��M���M�>���9)�I���� `��ɉ�ł�C XE����?�,\��M+�O��� j��������$�`��zvLW'�mx�hB�|9�Ġ<���?!��?9��?q(�
�X4f�-_�t S�P�l�U��ߦ��6mRΟ�	��0$?��M�;�يR쀍m�@@��$�ȵB���?�N>�|j�Ɣ�M3�'_DQ�Q푵\�U0�'T:>����\�Y������4�����sc�m���D K��i
�S�d��Of�$�OBʓJ�����6O�2�'?��W2%ń��@�����cA�L��'�h�>)��?)H>� �Xm�B�L�=�Nx�7Z@~�ĕ�/���qg�6uQ�O?���	4u"nͺN�h�0�+�"uK`LH�=�"�'>��'�b����p'��U��]��-��L�1�P�M̟jߴ�6!����?�6�i��O�nS-\�ؠHǠ�^���j��=6���O��M|��4��d��-�|�K��^�� ���L+K���b���-䘁��D#�$�<����?y��?y��?�e��{)nt*d�2?�y������)�P�ߟh�	��8&?e�ɳ�894��)����p�^��O$�$0�)�ӂ�H�;�*;m�B@���.8��y��ٟ3�䑖'�� A�֟��מ|BQ�x{ �H�D]�49��7t`���H�����֟��Iݟ�y�&e�28s�B�O��%#[F��z��/\���2� �O�tl�}�Q0�	ܔ'{@��M�&
���@���O܎p*C�m�����t;vk@����|�S�����4S��y3FQ;�
�E�k�D��՟���ޟ��������U�M��:�JN�w�^�i�7�?A��?I��i+�y�O!�!p�D�O�`2�F3{��u���0AUDX��-���O��4��U��i���Ӻ��P1��a����h.}��-H�z�(������/�F`"%�\+'�\��t�_�$��#Xf�SH�V���A��A�R5�*�z���Ϗf��z��[�k�P��O�#�x�a4��!i��q'퍸'�1O+��JٮQ$��Yֆ�z���3�~A��ʒA� 󅍙(?9�<��m#FØ|��`9I��YR�@ɜ'�.�S/M�D���c�M���b��
���	�z4��U3�paP�(B�p�����
/�#��	�ZT�aMQ���3A�S�.��@CY�Gpdd�J3e�񦈝%1J��I��Ʀ��	����?�� c�xѬ�S�lҁ��<�"�_����?q�z�f���ܟ48��HڲZT%Q��1hBj�C���DΓ$�mɟp��ǟh��1����Ƒs��Ǒku�����2�����ib�'�TA0��']1Oq�T �b��~�|����YH�5h`�i��Q�#p�(���O�$���	�'�	���������;�ܡ�Ψݴ
�d8h���I�O���@34�5#�nZ�h0
	���%�	��H�I+�=��O���?a�'��i�/�9�����g��#y�]j�4��|���Ԙ��'�"�'B��A�C��@N\�@SB�Q����|�|��L%i�e�'n����8'�֘�EOF�P�p�y�G}zpg\�\`c+���`�'���'��Y������{q���v��L[�W���J��z}�[�@��`����D���P=�H�G�4��bJ��\�%XC�Iޟ ��ϟ �'��8j�+h>u�RB�!F�\�S�.0@��@�
y�@ʓ�?iL>Y��?�槂��~R�7]��%
`B�:�������$�OH�d�O>ʓV�ltW?m�I7]��R�凨i'@`�5錐9��Ѻݴ�?	L>���?��V���'_��P$-�`�PUU,@55J�ݴ�?	����y�%�O���'T�@��S�~�;@o��ng�X�E���RO��D�O.��b�;��x��Sl*Z���o�he3����e�'��:GD{ӈ���OX����eק5�$��2,|Q�rE�7#����@۴�?��>	�(����	�m��-rrcƟR*�$Q��\-<D���U-E�h6��O�D�O2�)�M�i>esu�(F����!j�8i���M��?Q����S��'2�ѱ|��z��̠1�4 �@���]�\6��O����OȘ���LK�i>���Y?�$j�Qq��&��
�0���"������X�ɓ��9ON���O��D,qJ����R6J��-�㤏�oZ�����L���|����u���2����F0 ���b����ē�?L>�*��D�O��֩�EHeH��Z+�)q%�I�@����?!����'���O�%��oE�7�lH$#�T5:9"��iHP��y�'x�	����Qa�@�^�sڂ�Y N�}A���Q������	��L�?����dX�t��vHM5��<�d�
<��ˣˑ��ē�?	.O(��;	�T�'�?��F\�W�*�5F�#oм�ŉ�Dg����O�˓\�.A&�������wm��##��9�Vd��v�n���<1�,�p�S/��d�O ��ƒ��c�0n��Y���zl��貐x2�'�剢$�z"<�;]֜�i�
�!3sFh�n/�|�'1��� tjR�'�b�'c��V�������u-��0�F�ҵ�)dU�6-�O��B:��DxJ|Z���9R"	�?ĐSH�צ�r@$����	ޟ �I�?M��������ᚯ_�n(X��M?�����Q� с�>�Ş�?�A��d�"�b�}�j����\�F�'��'�8]�E#�4���d�O
y� �K5�1(Hoƨ�A
�ئ��	���'<��'��i�O��IKx�@EBː��T���j7-�O��bB�<IU[?��?�ÀޱR�̀�
5�.�*�c�'�n���OH���OH��<��	ʏk��!�Qa�l���J�5%���xr�'*��'<�͟���W �6 ��5!�4�R�M�<��n�ʟ�'UB�'y�[�0��c���ם1berKߧ���cȝ�3+7��<������Ol���O��W3O48��ɗ:R2j�(Ə�w?�+���^}��'A2�'��I�s��X
����䗺K(�1�,���rM�bo+q�b�m���(�'��'�
��y�'2�J�
g�@1�S�n�4�����Er�V�'p�]�$�Q�[?����Of�$��
�q���2v�#�$E�w�0{�a�\}��'(��'���ϟT������>{>0� B'G�Z���?�M�/O�xI�
V�����4�I�?!�O�΅o7�� c(st,8�7Q����'a��X���Ļ<)��ԁ�:�^��+5����G��M�G*���f�'nB�'w��m�>1+O,�� �"��{��D�a��#|�1оi� ���'?�Iٟ����*^���S�Ըj=H���U6*�ey��ij��'��J_*,������O�		 @��(�.Xcj���4K�7��O�� !�S���'��'!@%�A�P(����&C�?F��B"�tӊ����vҔ��'��	ٟd�'�Zc�0�XÇ�G1R5ʗ-�^iZ�O�-��9Ol˓�?���?�-O��Z ���F��L�&�ٟ/�l��`��%��'��	ןx�'�r�']�.� zJ��p녩9��t)D��5=���<���?���?a�����K{��ϧz� �۲��6t�L�i�6�4Amfyr�'m�I����џ�g�>�G��o�>��gB��L����Φ����H�	��|�'\�:!&�~��v[v��M�9
��k �5c�鐿i�V���	ǟ��I(),��I[��4�����[+8�}r�G�,%���l�����	ry2#]va��'�?�������9na⬺ �Q�0�\aa�	�1��ş��I㟀��"0���)X+Y�4�p��A��Y�ӮS��Mc-O:L)�/�ߦ�	�0�I�?E�O�NׂK� ��րҕO�p r����2��f�'���yb�~�θO�����À0�2�atÒ�(VE��4q(8x�%�iZ"�'"�OE����d �p"��W%ȟQLa+g
�xf�ll�:D��Ii�I[�'�?�Q�^hZW
�'���sB���'���'�Dac�>Y/O<������@�Ax�,����r���V�}��$�<!B`_�<�O�r�'�@Q-o)r�8P���"�^(4�D��7�OJU�G�
K}BY��IQyR��5F\ =?�1�!CI_f��S�����D�R}�$�<���?����$��0�D�B0�G;;30u��(՚P�J8 �Oo}Y��Iry�'�R�'w^�{E�ײ0�dT&
�bi�d#u�Z$�y��'g�'FrZ>�I�@�J}��O���L�`M�!X���F~TP�4��$�ONʓ�?I��?I�)S�<Y3 ��"�q�`j�zAr�J$ɛ��'���'y2P��"b����	�OkL�m"�8Е�؁]���
c�߶x����'��	؟�����f
/��'�<8�t*<q�5A!�-���ܴ�?y����OLy�ODR�'l�䥓>{N���غt�0�١�õe�2��?����?9�+��<a*��Ĵ?�j�I�=���;�/��#��![7nm�:˓�NQ�i�R�'��O���ӺS�m��Ր�a��@<fw,���+�Ѧ	�I��[*c��1��� |�N:��F�a����ЦG�\6��cr�l�����0�S�?��	��I�Sa�môdÃEz�9IMۚ5cZ�ڴ>���p����P�����'�0�22NہS�I�����|��V�{�F��O0�dI���t�'S�ʟ���$�ph �3C���bci�-�d�'��Iq����|Z��?��ڸ�ʓ,i�h����w�2��`��˦}�	-Q����O�˓�?a+O���ƒh�,�'�!��"L�a wQ�)bn�`����\��؟З�yRAХ]�U`3*w
�@�@
�_��EO�>I(O���<A��?��m�<�[�K�~CL�𢌟p�����.
�<����?����?I�����G���ϧ3���!*3��Q��Έ�S"�msy�'U�I�@�	�(��k�,f�;7�B���3��5:�!ٺ����O����O�˓N�(1#�P?���;7�H�@-Ľ �>�Ӈ�"g���4�?!/O�D�O��$Ʊp�D�Op�d�V�|$+p�AdD�5 â��_�m�ǟ���y�#;X֔�'�?����r�R�7HhIJ@�=O*�{&�ЄQ�	|�����c-z�0��y�П@��Q�0R��Sc������E�i�I�r���cܴ�?Y��?)����iݭ��*4�q��/�)K�P� 5�b�����O��ڗ8O�T��y��	Q�-I����à?�AA�Ɲ=	��%��7M�O��d�O�i�c}�^��IbƋ���#U苹n;��rJ���MS�.�<9����7��ӟ�ZHߠr
�3�]a�����Q�M���?��� J8JTP���'`��Ov�R%��2fFQ;`��~�� ��i�BV����h��'�?Q��?Y�R�3#�EA�(SY�)��`׾U�f�'H�`���>�(OR�$�<���{$��>vHd�'�_�ʵ�Յ�P}� (�y^��������Ixy�cٰl���a�c?_Μ$�$g�$Zl�d�>1.Ov�D�<9���?��UF�q�acE�'Y��s&*\jќŲ֌�<I���?i���?Y���F�G�|8�'H#�<�W��0;��$B�g��poUy��'��I՟��	H1A�w�LyTgL,�4�a��޳�e�Q#�M����?���?a,O�)�F�G�s�M��ޝ}���ac�&�`< �u��� �$�O���7#ln��1}���z}�*�o� �2aO�*�MS���?�+O<�E�}��8���zzH�0 ��R�ˊ���L<	��?����<K>)�OJ���4���J�0Хb����ڴ��$�3zX�o��I�O����~��G�D��iS���"���fW��nڟl�	�.��V��^ܧ�4s@ހo_\����Ol4�in��U� �4�?���?Q�'\�'����\d`�掎jq��#���.p�b6M:P����.��,����\����c<Ru��<6 �#G���Ms��?����r� C�x�'TR�O�h�d�?#^�S��\Z'�i��'A�y�N0��O����O>���(�<��|�f�@glU@�OBڦ��	�\�.��I<����?�I>�q�? �`1��ԤD�$ER�)DV����7X�j��x���'���'��Z�Xɣ ��e?�x�"U|0�y���nG��AN<����?yK>���?iT���v^�rf �X���a,� [�^)̓��$�OF�$�O��B����<�~u����.]�2�IF��]�����[���	꟬&���I�D3�$�>�!,Œ;�:��uoڛ ����E�m}��'��'��I���`K|B�D�)=����ȏ� �V-��
�K���'0�'���'/"p�'�||��A�Y6~dA��ِX��<n������lyBl�>V������\�Iu/�'y ؐ��AnC4 !��c�ß�I5ܦ�IZ�I[j􊛑T��VE�w��x���ݦu�'�z���{����O+��O0��^�"L��Q�J�
0�2��Z	�lğ<�	�}�"�IU�	A�'�`5���%r�>�R��*B���o��(��٩�4�?9���?��'G��'�r�Y<9���6��_���4��7��,����#�D ����P���z��Y�܉n(hrR�]��M+���?�]ے���xb�'��O��:GȈ> !'�VR�~,���i��'��e��G1��O����O�R�
O�9�Z���.J<��e�ڦ��I�hL��Í}��'�ɧ5���z��C��g�t��i$��C��&�$�<���?Y���G,��UlؑoȄ���
��{vsc�[�Iß ��_�	ß��8X����E��'c��h%�WC�p����]�ҟ��	֟��'&�ˁ@|>��p��
K�a�N�M�Jeg;�d�O��O��D�OH]����O̵IQ��U�L����ƻT��M �.]u}R�'R]����"�ԔO�R�=��H+%�P�ԕ���(nT�7��O��O����<�PA[r�	w"\�Ƀ` ��i`�ѻ��7M�O8��<rJ�;e��O��O2\�+ǊԒ�<d�B �p��عo6��O���D�#tf��[��?/���Z�KN�J���^��R��֠�MTY?����?���O(��F��8E�&`��m?�rV�i2��'G����Ƃ�J���Rd��/6T���4b��\�f�i�2�'mB�O!*O���J.4��4��lQ���	�,N��@�m&Y&#<Y����'t��GH�"V��`�!HC#m�6p�Kj�B�D�O��ָY��S�D��) fH�����l���І��,��<9��ځnG�O����ѫ>�b�ɓ@�(�RU�5'�i �G/9Q�B��&G��M��O��hc��J'�B���� �P��"���AB�&�& ��*A���	A�A:��@��t}�u	�8HqP%�8v�Z���<m�h����9)�M��/�)F�X5 �[`
��T.�4׊H��	R���D%U�X�z-P�,�#R��`Ё@�]:���+��B��J��`N���F
.p�\L�U���'Y@��'���'a���'��'���9���&?nx���,��0{Ǔ'!zh��Զu�V ��j��z��RV��0&�O8p�/�xb��"�?�����I�-Z��R��A8\G��B�U�LQ��韠��i���OW@I{�wۨ0�AdF�8�r�#
�'�f7M��W������;����@ (k-�$m�sy���� R���Iz�$j�B��<�v���_�]X�y������'�XY{�,iB���)��T>��OTD�yw'ϡEC�<:�n\'�.T�K�l 7��y0�ũ�#�	�2xD���Չ6���hL%� (�Tb���	Jb���OV�}��O �(ڴ/�D>Ȩ��,|���qh�E�F��!�JѠF�R8z�椚��4�R,Gz2ɛ�Ҭ�l2�@0y�b#|��6��O����OthclFVZ�$�O���O�n�m
U�KH���*�7T�jq�Q=�l��ɫݰ�2fJ;�3�$X�#%���`�!�p�Y���o\�8�FF�fb:��	�b逖���w֞�ڙ'����ꈁ
r�Jҭ��c�����'����V��4�\�=�%��!`u6`�2n��f[\A�FJ�^�<i�[�0.���T��=|e�d�<Y��0z����ޟ �'?☋���� JƵz�K���6B!�'���'�Z�u7�'��?��`0�$ԲV��\y0�S5k��W����pV��/w�H�G�'���㴆��]�u2�kԯ`7h�kC�Z�zt٠Vi�cԄ��d@.��Y2Ҁ�xE��
b>;� ���'?��]�0�h�VHH�lqD(��#td�̈́ȓs�Vl�$Æ`i��1�&�KT��<�4�i��_����&�M���?pA�6u�H�dٜ)�\(Z���?���Y�f����?��O��Y����?X����A��=�Ѡ��Q(����	�-���� e��T g��*K� e�!O;O��R3�'�2Q��84`&@k@��R�cn�*~�d�	��p�?E�CM�D���ԥ�*�ԅH3W��x�r���J�' j��ҕ"�!	S�c���O��g�����i�b�'��38����	8M��#g胐|@�mB�e��)�t����HQ�"R:{�#I>�O��S�z�5��n�C�+#��	���'�ꈨA�-eɧ�π X��3φ� H��P�h�.� E�>��������	���	E�'3��}K��]�r9J�b ���>�0%�<����<�  FAشq*��B���NM�����:,ܬ�����c��؛'�
h\�oZ�����؟$zdk��8��m��۟��I���
v����(;{%b�d$	� uaW,S:X�T�	"  jݓ��J�$�dۺdͦ$��%	�Ex�!�V
�&�l)J�	-^Hd)�᝚n�΄Y��I�-i (�h�'~z�Z�!�%u,��j�#.�0��C�'Ғ7��OL�sĥ�Oq��Iן�	�Du�<H����hʆ����W���'�!�F�]�|�ˆ
��Lg��1vr�����M�Ĺiv�'���Bp�O���)_��X1�)Űao� �%�>3�C�I�~�H��RB1�X�@�K �J�B�I�Zf4�S��jhi�b�	?�B�ɾs�@ݑ!Ϙ4!.Xxê.L��B�/"�;U�s(��t��'^B�	7R�N�H�r��MH��k�XB��:8��q�G�4fNy��'>_�|C䉧+�%+!�׃|"<���5�PC�I�3�X"ugϛ�[C�U�FbC�I�A����B�4ƚ�J��C9�B�+ nh��C�]��%��㈏#C��l\)�爮pΦ�
6�H�>X�B�I�������*�KŃ+��B�	+ɤ� �OɣA�Jc��D�*D�B�		D$#w꒱L�j�Ӑ��ge�B�	9)����>mV����Ζh�6C��"qc���R��'pp��,�5v�B�ɒC78��R	#WT����̍85"�B䉷y��t'���6�R�G��`7�B�	�U��M�FIϥb�qӤ��!�tB��,xBvբ�͎l���:�N�3j?�C䉩@��Pu��'Iz�P1%�+BJC��9��q�V!\��.���rB�I7k�1 r68z��xk�,�8B�I8eu�d��喼<H=Z�5_WVB�	�Vp��[��Z[(���@%�B�	�ar.��Бfخ��*Z�Q�B�	 o�B4���h���b!�7S�B�	u�����BFr?���r�Zz�~B��}V���TA�&P�j!�EZ�]~pB�I <�M��,ި�D�zB�V�n��C�%�-��'3���-ֈZ��B�ɩ � ���NW!T���m�5>��B�	�ZY�'L�=\��<Ja��Z?bB�	���P��Q�N5�&��b�P�	�{R@�g ���$�+f�6)��R�"��:s,J y}���1Lz��KBo
i@,0դ�<\`�R$�޿�xb��u�2d�!�F��A��ȯ�p<�E��\c���K�1h�R��T�1A�.D����W�<^n�1Ǐ�U�3%?}�b�]��%�=�"�IP3H�$�c�d��c/@S$Uv�<Q"-G�t(tP"Y�UE�1�TGrܓ&�|�# 8O����Nف9�ꕢ��0G)�y8�
Of�8��Є@�Z�e�ڋH]�,���1r0mH�'�(̫���5<��q�j��u
�Y�Ә'	&T�W�q�9���C�A�	��'�0��'�׎#c��RɊ D�H3�'��Š��E'kc ]���@G���'c���&�^��CLrr��
�'nJt b�6( �a�N�G��
�'h�8�S�/�PeK�	^��h�	�'�Hz�`ZA�F1K�f��}>V�h	�'�xy�F�Q�X�8Mbi�v��N�B�I ��y���yBܜ:����C䉘qTّ�$ ?ʎ���E5d;�C�)� uy3�7K�-���S92�9q"O�i�jY���	��
�'HV�a�"O�p��j��1�.4:�G0KK��c�"O~xi� f��d�ƣ'e�-��'����&�	�B�����̑J�8�'(
e�B�ɦmA-�P#�e���Ʉ�g��'�=3	l�S�'FzJ5Y��Bl��0p���)_��A��`����5j�)PZ�%ȴ��#9X֘�=�v�(c\��ʰI��ZԀ&Q�0�\*��|�l\<2)�l��<��Tv�J<59b�s5'Ȟ9��5��IG<��|;.p3��ް:�\�ѡ`�'�� �p�f|��P��O�^ �p��%�J4�%M����I��'����!.qxx}Z�"��]x ݐ�Č<�b�l�K�L�24;O?牙.��|�� �.;(�=�b�G �C�	�zڄ@+��� �֕�fɿ9��	�j�q	�i�����\U��
6�ލ�n<��f�%{iNhY�f(�O,�IwJ�"�MK��0"LQQU��%�T�!��G��!c�5��Z�
�0=��X"�n���eX��6L��x���O������H�'2nl��(Ll�������I����hI���Tt ɫt�X�9��������?���#}�,��?�1;N������IWHE���X�z¦��ȓV�d,X�@�9�t}zQ�ռDU�I̓u�THӣI&��m�$��=Q�a�n���v ,Zk�vk#u����	N8.������'7�1�g�D���IO�C	��Q��48�@��V��&n�v �}�^���	�rWj�� ɝ���i*�ɖ2I��H�vp:�Z���ص�\2�x�K>�I~:�J��M{0cJ� ~DC�f��p��nע�j��Q$�|�t�79iv,8�{*�r� ��g�M`S��0���q�M�l�DPJaB�O�	��[;W~��D�T�6�3���S��5cpR���G F���*�:61OF���"�v��P1/ŏ+pbM?�I2vhh�bd/�,�6}�Eh!VL@6�h��O�d���,h*�O��@�b
�;��ћp��V� 1aD#?���	�I��ku3��L>iɟx�C��Z�����( "msŞ|  b�lq��/�4[� ����'~n��R$�yT�)bcb�4OK`���8i���K>����Of%+$,L
S�:�F25c�cF�B¥2��C!+t� Q�{*�12�*wޭ(�-��X����"�R^�C�C�O���������$�_� hu��-�y
ײ��c�xǒRK��(�m����҆�~Γ^lu�UnL+���x#f#��I_#��z+(&����F'N�ֱ a���A^���E��/�e� `+R���������r$$@�|&���Ov���&�L�0�(��K��pI>)ł[7]K� r�h��o��ː�h��bT	�̷Pq� ��B#���Ct'V�P�}%��E��'���b ��G�h{$�g���v��i��izЇ���q�=�O�΁�A5�6Qjt�7yAӅ�X��`�&�in���.�(:����*e�X����'9�D��n�b�D��f/A���P��%*�q���:Yb� B �R����4!�a��yB �H���0)�!uj��!�X�,�[F`K7(��Q!tMP4Ҍ�St�B�%��u��'������
j�ʧ#H����L|h%`�ނ��N>a�	΢U���D��̕�c�Fb�#)���j��:��|�(��z��0��H1<+��u��-��#<ї��0�~���FP�5Z�[#
=� ��
i��X�%�)Z'����O��z���*E���~��I2}�H�Ӣ���썆�ľ�c �Ҩ[�.�xVLN	~��<yRD^)?���E��F�(�>�ɚ;J��:�H)/�@e����@��X	o<@d����T�@���LY�l# C!� �^���$�8?<&%�2j T�A�!�O���51���D�O��=3V&����I���_{� �T�|��O?;% �P��#��h��'�4ٸ'�� �Ι6	N�zʔ><�-��A@m�h�'�x�Y�S>IFx2��7|���È��"(�J�=C�|��ΰ?��I�5%�b�S�I��5޴_z�,!���g,x| �7n���/�22�^pz�G��,���7���:sjӟ@��Ls2
�L̓ t�Mq68�)��S����!G�!?���,�%s��0��[i����)Ű_}�x
��/m�	Ra��B�A�5,�8�	�h] ��{�I������62�R�c% թ��ILzH�q���XY6ქ��9|�����d:�1j��W=:�����'`es��}��03�����b��e	FW�>��d����D$�.��I�O���4y�,�n�������a��j�Z�7K����	i:I���6c��H�P�,-�t���2(x�h1�N���6i]7)��,��o�6 NI�T�M�Vu��kLQH�rqx��� UT95iV=�1OT8	1aF>����O�~�:RJ�2�\@�� �<P���'�t(2C��N���{?)�O�)"� �>� jt"�L@�W�j����?ji�t"��VBH�'��@.3��?T���O���T�H�pռp���M@�Y����~�[���yC��R�����*Y��H �BC��6F�Pcج�qD��Dp.�"0�O����ϸ'���"5N�#0�"1�'{��h����<T(����r�}E}bC��N!���G�O?�� S�f��$m��\��Q0/�n@0�e6��pH�D��拄z��y���6I���ɒH˧!%fL-5'zY�<)5k��zXY�c+�'�R�q �=^��Uj%�Ё�VP�'����
W�6r��G`��8���4pq�
m���*O��y(VզG��k���o�����'�g}��O���O(6�9�g?� O�,~���5�*;���Pd��p�	�Q���
���B#��g�'��T!��ڻm1
���(7_ظ�se[5X����@�	�p񅅛��=��I�[*���-SN2y����4��T;` \,~`�1�(+�A*K�C\�C�������O�My%?TJM���Z���8�'��Q+1͚�+�����[�W�I�A��r,��4�u��ћi"6!� �2jqå�^)]튈ӎy��N	m���"j�0b�0�+����'��]�UdeW�%Zv愚k B%{�9�aPt�S��Ω� ,L�gp�\�Ul6%׼$���(�Q�2��)����[�)� �
�m��(�J\�.�ax�wt��ʲ�
gP��%O�[��G�g�v�@���PtdH�d�@)a"��;D�� Ǐ.����!o�wY���$�<:D����Q,^e �
�1~����.^\�L3�Y��>"��O]8�p�7�<&�j�� ���>y���N+2v�#� �-�� a�l5ړu,=�ю��[��-v�a��)Y��ʳ{�@�P,Gxj�I�̜-�С�y�Č#m��ѣ�TJ5��p��ָ��'xX��F�K�QHX�*1"�7̹�'J�C�F\�1���#th�|��e���d�D��?}b.Ϲ��� O�CP.�`7A�Xf��1���; �/�0=�C+m��P�v�.$+rG��p���n�P� $hq�Z�b�ayB- �h����*�9�L��7	�9`T�ę��P�g����Er��ۂkٰ�z�n�(D��(˓EW�`���pш��͚i�<@�'+�()p���e͗�v�R���18�����J�5S"x�u�0Y.�q�S�lpA!��C�'d�<s��!��]��B�
Y"��Oޘ��@�e�p���)P����#�DG8��3�/ȡrKl�ʁ#� �1d���`�p]dpy'	�mu���H��V��M�70�RϞ\�Ӂ$B0=T! T.�6��J�-�]�"�K" e�!i�(��D]�x&hB =���%"�D;�$��%�򰂊���(k|R�yB��`�^�ql��a.���L�V�x8���%p\�K��w@�MIA'c����bՉ]fZ�d�� �ՊS;�c���OZ�`/ͤ ��W�@�)AX�1įY |���;��	0z�
4-+t�4	��??��	�B�V$� eQ�������Z��h�dU2O�d��g.nH��K��(���ݬ=�4[�kɑwa�e
V�D��Q�U=�{�L� �L%���͌}0�)�S
i޴��,A7�����O 9���6'��`��a}�Ҕ�'~Jl���������
� �D��Զ�
��W'��k+�	 eA���4��s�F�h�<���
&�2	�$c�>�p>� @��ߝ� ��p��y���֨;���Y��TL�80
3Ď79�hb��3���]/��B�A@U��,U�">q���h��& �*�>��³?ZÏǭF��`��'(�u��!*D��p�DO	_�bl��EM�ZFN� ����xk[�m�R�0vb P%l9E�����L����hF�`Q��YDA��y�A�X�h�����M9�=�S�N��y2Fʍ!
<\j%l��E�DD���y��!M">iR�!�*M�G�L��ybV2����2e���؃Wh��y"�V/	�*LI�I ~li�֊A��y�`FI�'-J8@�J�ڔ+�(�y�۬,*1$3m0�an�y�$����.1�P���T�i\I�!"O$��@a�R�5'+1&���"O��{ƍ�}	�skS��= �"Od4(��^!yP@*��:�f�;t"O^�#nB��<c�OH�CKv=��"O��)��Z�ty�i;Sn1s/z�s�"O�xP���"�(��N��@M�c"O��cE~��{��P�|L֕A"O~��F+�y�B���윀[d\��A"ONБ��y��$X�=lT#�"O��1��K�OZ���`�|-�q�"O�)bw��z����!��QE���"O�Z��@R�O��d��m`�$�+U�!�� R�2�O���r6nƆA�ѱ�"Oh�+bܡCqz	�7G�;o����!"O4BW�ө@��b�%[<�J0��"Ohh`�f5�f�G��7����"O �q�s�rA���!\�����"O��bp"�*��Dq��C�4���i�"O��cW���8�
��r�Οf-�q��"O����" +#Zn� %BY:%,��j"O���R�n�=�s �G��8�"Oi���ރ)vJA�GNP�_�r�	"O����Pcx82�����2"O�yZf��s���ɰ��$PA��f"O`�(�I#\�`�Q��تF0�K�"O0�2T��� ]1W��> v��r"O0q���ђ$��m5*�c\��"O�s���4+�� i�"lK��Q�"O�	��ĚwPqY�ED.�ҍʃ"OB$i3�[/Qĭ�����x(�"Oz�a%��e`G(�B�z��1"O��yE惉/x�V����N�s�"OU ��I���S���\���"O�a",E�7 ġ ��5_p�H`g"OP)��f��l����Ŗ�xjȐ��"O�m�T�/:�jz��K�g4,X�P"O|�Se�ܫd��I@��+����"O]�ku`�(�,�'l�ع�"O�wE4|(��S&r��"O�����1I����j��t��"O�E�7K�p��9�3�N��)#�"O��s4G�<Q�\r��Ӏk{3�"O ��T��h�|����zbN!�"O�P���<K�仅i� ]XU�"O:�FI$[xZ�h���%PBu��"O 0 Ћ�:X8��E'ԼJ���0"Oص���~���!��C�q�"OTy���=;��% GS8"��p"O�8yǼ0�x��΀�ZLM�"Ob��1)U���8���P'�Bذs"O��+v��*٤���D@�G�P-�"On�K�oA�6��afH�{�j�A
�'¬�q7�9{rtA�El��Z9���
�'�l���ʅ�"Z8�JW�&�t	9
�'t�y�&@�8H9p猈�#ir]�	�'�nuS�o�;5Y�8*6�%�FX��'y<@�U�7$��ta�]�w.m(�'��pB*#Xx a�s������'�p!�
ح/�~(i�_�����'xJA৘�s�\t�r�7Rd��'n�W��M� |2���$��e@�'������SJ�}��f��Tx��'�F���|���i�EsK�e�<�U�6_�b���G
����d�<�2���_���g��9��à�x�<yTc�>[����Ac��+ H��Ջ�K�<�$���T	��G}ܥr0�D�<�q��lgT��׭ 1$
򈂡 YC�<	�k�3D��MsĦ�,U�\�!�K�h�<!�˂� �<�ѧ&x >H9��L�<���_�_J�����"��!��SL�<I�n�)	��7V�|��J�<9�/S�0a���:Ԥ��M�<q��/Y��F)ǉY�2H`�DK�<q4��M� ���@Aa�4�d͝J�<�EDO�c�.���ק{"a���YH�<� 2��
f��Wh��GF�uHq"O���BJL�Pk�!B)��aV"O�	S�N�v��� ʇ4��,p�"O|Y��E��Q����o]��}�4"Oz��\�R"�8�$�\/5T�["O�QГ �ʁ�$�T9~�P���"O�A���;?�9ŃЂCx��"O|�8�-X�.�"�BB�<e�X� �"O`�6����vU�X�"3L#5+!򤙻_�$R�l��"=�`HumT�,,!�+��cՋ� ?�(�����d!�$�Pe9`@)|�p�b'!��+�L�k��ל �(˗n��[$!��ސg�ћ�;@(Ds2ă�!�D^�A,�b���a�����R+7�!��C�yԡ�fn��05�Q�P	E%�!��A�mBܴP�d�p(n��苲'm!���>P���φh��Q:c�A	J!��H�H:��D'�4"������!�ֻGa�(sB�PH��C�&t.� D{ʟfQZu��C��	 ��3l��W"Ovu{Q
��}Nl��@^�6!"O<ppe�70�)�%�B!;�>d"R"O� C���3C��rd�P� ��x�"O�]۱f+[���'G69ny3b"O�{��P�B���ZAe�!m$�|�"O&]�@h�.�&˄�lH�"OZ�"�/)KlmZ�dK��ݳ�"O���Ժ#2�%8��'?� ���"O�}��K5&ix%O�G�z9��"Ox!9���H_f�XE��Y-�й�"OX ��HD��� Rw#DPa5"O�DI�m|�����{��ɗ"O @`n�.~F�SR�h��P�""O�m�$��qqTnĪP�pHV"O̡C�������"�	t�6P"O��s��Ճ(0X����+^�<�I�"O� �v���Wa���*ϐL�
���"O����ҋW����X?Cq|+"O�d����66$�p�B�8�t���"O��Q$�9}���f��0�d�1�S��yb��m�d48Ԡ=5�8�(��yRG-X�n�rsh�ֵ�� R��y"�>��d�-~p�(ԀV�yrG��d�0܁r(�J���	�N���hOB��	�(R�3� �9��eQT!��F*!�d�/uVu��ʀ)#&p��m�cH&G{���'�
���Ȑ.��S5��;a�y�	�'~^��e�@U|�4��\o�P	�'N�t��`����$X��'f���Β&V%QFA�q�H=��'�"����M%�.�K�ahN�,�
�'�h�F��l=P�c2�M�s�B��	�'X,Jfl�~i�)�n�o�	S�'�d�a�;��1q!!;Z&ī�'��D��휂'-hyR��I�A�����'�XP�V�N�&]�#O�7���',΍�VJ̴o�T!3��[0�-�'�\@����Y����2�ƋG`��1�'[�@3Aߜ<�s
M�8�F@+
�'tT��L 6^4�r�:,�
 z�'�\ɩEK^�.0(%"Ҧ��?H Y�'���"�=%ΰ)�4@ɘ=�8��'6p�f�':�4LpT��:�x����� ��� j#@t`�*׈(lV؃�"O�xc� �v��r�Ӟ5L(���"O:qB�'� �r����Є=�Pq�@"O�,Sq��	S��r4o�.$��%"O��bo�oZ���H$F�NeC"Ob�U�B:cnUr�N�(o����"Or�2�C�jbZ50�NZ����"O�TZ@��GCt\�P�[�"^�82"O|�9B�D+!1�p9���)a0�3�"O<h6��.�\�#E�^��ݣ�"O �"t��
���!2��6"O�T���~%�`U$������U"OnMJB-�kЬɉ�B�7 f��B"OУ��l����aa��m���"OvP�2��=��]x�@S/���b�"O�E�0�1)̚!8`���|�z;�"OvJ��;(]�O��^�^���"Od�b㬄�]��OK5e� �"O~�;�!Ӄ}���Bk	5aK(��S"On�B��F�2n� k�kdt�"OJ�q@�_�ta\�@�� x�*i٧"ON��4��)�|�q@�G�/���"O�q�ZT�Xp�c�Rk]8E"O��g��2|F�	P�"gT��"O�L�l�'O �L��	\�I4<ڣ"O�\��/�:Q� ���8S�N��c"O��p㇒>R8����8'(��@�"OPi1	�/P�x�7P�~2��g"O<@��cZѸ�dG��>�d"O���j�U��Iٸ/�nuС"O<��-�?@�h�8��\p���"O�P'�LC5D��woL�Od�	�"Oą�w*�D��i2��fP�8H��>)���IU�-Fi�p/խM�h0�#R�]�!�d@:���ȇ��>����Ł��!��4W�@�N<P����	-@�!�D�)w@����B�a�jm�T�Z�7���y���&F",��� �%.����k8D��J3�V�5�깛���7� �S�5D����W�\����I��{ւ)D�L3�Ƀ%K&d}(�
Ш�l鴉&D����A�c=A�rB�$xl�S
:D�|�#��VO2����ǏJPTc�,7D�,�ԥ
/ �޵)�) v1�L�6D���� �K�ɒ`ߕ�>�fi?O�#=�&��4A��h�D��/1��<�4,[x�<!��ίQ� �ʕ�گ1�h��,J_�<9#
g���a�ѳ-a�`
�HB�<��#�
�h����
8v��u	Y{�<Q+� �Y3l�]Ny��JFO�<�`Bɜ2��A6`N�n`��^q�<�D��¼�4�=\Z�V�C�C�5ARBiA�e�(H~�W*ǭx��C�ɴ��l�f�7+����V-r�C�I����	�,��s���*pC�"�z,x�$�N��A�B�L� v�C䉹K4�ٻ�aґS�l�{���T NB�I�9d��q3�I9?���HH;?�HB�I5I�^y�M�>I�ذ�CC$A4B�I�[R,��3bH�.b��i���(5CPC�I&��%���F�����ӾU�HC�ɳfS`��1�׎!Ղ���0�C�	R�x�z�'��?�pز.OX08B�	�z�!)��]+H�N4ز�Q�L��C�)� ���1j�h�h�@F�yq����"O�Q��@��n($Wa�%f��r�"O36�G<�8}�� ��tX�"O����#F_�}�4]$j}�`W"O�xѧ�j.�툢&$m���Q"O��f�YWp���rDu2�"OV2��ѝ��HÁ�+��$"O��#��9�d-!$NV�f ��"OұI�'R�I\�-HB�̲�}f"O������u�BK� ��C"O���ҵ�v��B�L)@�V�2 "O��vHP
11�ʳ��7E�����"O��Z�N�S/�8��$P1����"O^�3���-�ޥAB��Fd��w"O�$CƎ;XXDh�,d��C�"O��s���3Mf�y�m����Qe"OB�JQC�*n�:�е�+~�����"O>�I@H�t��MH�,�Ħ���"ORM�4��,]/���
ӓh"�]�a"Od�U���)���r$��S
�i�"O�EA2)�+#6�ܠ�'����b"O>� /�2�rA�@!m����"O"�ᔏI[�����G��ؤ�"O�����2@�Q�Ǌ�|��4�"OpqB�-}�K���N�v�˂"O�Q�6&�
%M�`˱#�bt�Q�"O��9�oB�G�d��X�j\�P�"OLY��� R
� h�jV��X%"O$�9�m�',��C�-�cIb���"O`�a�.ҒA]"�"��-�(`�"OF��$�IV{����J݋/�~H9D"O�U��J�s��b���D��g"O��pP���
�,��ĤU�� "OT�g�؁$�zy�eԓ\�PQ"O�m!E�T�#��1tmU+ª|c"O2q��c��o=��P�����.�q"O��j�oHu}���J�����"O��6e��KF�Hb��0��Lc�"O.���J�3k#l�j�FPU�ܐ"OB��C�xND
���`�`�"O�(���KR�S*�%Y��"O�t�W��j��%��I�@p�|@�"OP�𣄍e�"�k7�:���"O�{��ӢH�H�3�E�qӆ� $"O���Wf�6~%A 씜Ѣ%��"O��J�<,�pY���3��9�"O�|��#��a�5��ْ]�8��"O��+����X��Z�*�v�8["Ox���H�t�l���ޫ<z"O���%�>o�Bt�g�M�:iB��6"O@ Y���9Nc@�z�	N?s�1R6"O����A�7e��y�өݎ>u��x`"Of��gÂ�I0
}�3'�_�|b�"O8���
Y'�DY�QBBq��"O �h%hD�W.�F�I�=h�JE"O�墅k�_�lH0�f*.|`�"O�� B�-�f����Y�iN��"O<��K�� &»2�!"OF522f�D�N����N�w�j�)r"O������ZjXҐ�����jp"O�5�uh�%HW,mr�,����"O�kR�:tdH��%5�r�*"O�A0���B��MSeN�1bi�x�S"Or��/ٚ=^,��*U�5c��	��� �B���Y��HPѯ	"I�H��3"O�@ �\\@��׿6�iq"O�U�rc��e���V(.�R�v"O�}Ql��X��@�|��!g"OX(8v W�@/H]��A�.xpT�@W"O&@A�Q	z�@�F�hH
�"O�Y2�Ο�A����{@\�"O���b���b�)q dj|Lk"O�����r�
Ģ�%KDU��"O���!�D�d{C\gB���R"O�$y�␘t�ܘCb�4n19A�"O`����M+	B�!bsK��dkB"O�-2e�H�I�X1j�*JQ\�	!"O��Z�'�I�4�H#˂R����"O��.u�H�Fm� ��UZ����y⅀�H܉�F
��i��a���y¦ݽ��Em�;	Z�����:�yrCE	P����J(P[v	�4�G��y)_�XڲXiÌӬD?h�҄���yFV��$I��=�I�m�?�yrf�+��1�e�Ϧ;$������&�y�%�<$U�\���y@�`�Ƌ��y2��Na��AV��0��I;�y"��7V���B
ճ?k�P���y�-Q��De9'��h
�i!����y�͞�kNT�#�k��Z�4�Ⅼ���y�kf��A'�
K0�2�n �yB�%z,��ÍS���3%��y��4��H�k�Qg�!�FMT2�y#��C��pՇ�7�r{�BU��y�B�����ͣ..�(�n��y�aɯK$���Ŝ�"j��qb���y�)I$J�!�>�6����Q�y��_��i�EYd`�EO(�ybaC' �2��6eP�*��܊�y��F7|��0���f�%���]��yb��y)VU� jQ���b�y�\�"}��bc� p����T��y�b	 ����A�`����*Z��y2�]�O���p��Qy^�� ��y2@E�MQ�TYt�N+L��U�um���y"KҴwlH�ql�E���%�y#P�*>��Ë�evH)뤫X��y"��0a� !B�٫K�,!���Y3�y�:w��aC)Q�FSv=p����y��ߋLLqi�f߰P&`p�l4�y��[�D�l1�GKV�=�fDऎ'�y��ƀ?��$#��/�����<�y"懏~��T"^�&�L�IP��3�yr�6Gƪ���gGM�,Zgʀ��y£� _.t��@mPt�Anײ�yL�#�!���gM���sg�4�y�-W�L~�y�3b�&L�*���K��y��X�I���bnǮH�%1B���y�KT8M{�i�ظ>��iQ�E��yR/.�����ܰ9�Ne�p�E��yB��mԬSrHU�6=��`횁�y"g�H��|����y
@����y���U	:���qe���v#��yRƒ���b单<��
��G��y�DM�B#�h�Te�d�l�Z'�J��yr������I
e���p��8�y҇��
��xI��ݢcp~�9�)B��yr��:�PB�R(g%�����ώ�y
� `}�P�p����0��4�U"O��1U��(,4�k�N�eZa3"ODA��J\��z�B��H�%"O �G��.�ʒ�J��y2�$	>��a���ȗ�yrBI�`�Hw�)&���Q	��y��2h��XT�+J|�����yb���$�
ͪa`�7�L��%�*�ym�9�4@h�Ö�1XRd��䊃�y���/�|�#��R3(4t9 ��!�y�G��!#fϋK��r����d*�O���%{8�dʕgI��<��"O4q����e�؁�E�;V�F�T"O��+U�ͤ<K8��w�8[���"O"�H6*809�cb�4����"O�yPD	��f���Q��R%/�*��"O�-X��	<�^����9a�<xa�"O�i�"
�湘��\�}�]���I@>�z���"�hUB�ξ. lyD�#D���&�}�:�R�ON�cE4u�A=D��Áh��@uN���-��j�'D�P9CZ
7��dd���r
���D"D�T�D Z�0��YK	�VԪa���=D�X�d
�S\����)R8�ۂ�%D�4ʗ	R2PIL��*I'J"�r�A$�D!�O�9�q��6n��x�:�1��"O��q�n�2iS/�.���*�"O]�5��$ �h؈c��?G���"O��+@��)Xv�+/�V��p"O�YoF�jW"\�RJ� [c�!��N/D�`A�f��jt�`��C4	P�8u-D�2 ��40F�+�@ʗy����M)D�x�eL�+T�t�Y0bG�R���h&�O��dVٺ!v�ڐ	]h�Ҍ>�C��$BP\���jl����K2pŖC�	�I��U��62p��C�x�C�	(Qo\��/DVt(3&��_�bC�I��0����&r�@r� �%l��3Z���	@�\�R��tR�#m�ў���I,K>�u�%@�2���;PhY�.���$|���:n!�e0dN(
�U�#5D���U#�Q/`it
��MB�p��3D��C�()�60 #O50ܝH��$D��{ǌ'$f,�I
/y|��V%$D����3~ܓPK�r�H)��� D�9!��e�:�Ȇl	61���`*D���NK&�=A4+��jUX�3�%(�OT���7�|�z�%Y7>�P�mT�|�d:��rRD�4ae����$�>'���0	0D�0(t�1.ĲA�r��3 c��Cv*-D� ��Z�}�ʹ�e�BS�i�t)+D��H� V3��3 �7"�b���*D����a��UHU12L��l��R&�<����ӹ|(D|�G�T�;P�A����9��q�IP<���ϾX���S�%ЅrEj�<���	8���4M�%�b�O�h�<��B�&�,	���X�p�j��\�<!n8�(��L��
Y�-���X�<	!JW�.l��Ah9v��A&UO�<y��=2��<�V��=2�Sc��˟�G{�����ꐁ��9Q-N(���	XKxC��5�v��2�l��)P�c�bC�I�t���aaH�%g�Z��a�@�Q�^C�	=O�$00�̌"E�pJgΜ�L�BC�)� ���%��L�Ը��l
I����"Ob�Q���2Y6=
�fM�c����"O���Q�]�v���#B�f4qI�"Oz��ƥ�$l����d�q�(���'��%R����iV�.P�93�$���v����N{#ص`3'� ��)V[i�<�*@7�T��Rm�Y��$)p��c�<qǢ��y@����O�q>�C��]�<Y�K�t^ (�CZ�b���d N�<y%l�"j^Y�d$V������<�/��!4�U��O�Bᚱ�@G�	g���ԗ�lH!�H"{$�p�'��9L�A��?D����LZ��`���T�&�Ԫ=D�|�֭�
Q�9�L�1x�͋�B<D������)���&吞�rL9�:D�x*�F��Ѡ�4%DDx�7D���.�.l:�P�&E.��� T �O�Ojq�2L׮MF#%dN3w��㟀��{��~2�B�3�J*# ��!���#���y�C��%���-�-U��i3��y�d�1�����I+aun@fK6�y2���쀸�ZE�KB��y�I�Yn�=)0a��U�<uِi��yF)`���)PO\ك�B�yb]/M��-:@kM���$FW.��'�azb�N�~r5H���8
��쌎��0�O�l�BMX��8��B7,J�ɋ�"O`=! ���uQ� @<vN�H��"Oq �&A?T���&�3<>
���"ON�
`�R�T����ZN��"O�CVf@>��! �	���%�\���>��O^�H
�4~��lg��*���ɤ�|��'�^����F*Z���xը��$�#"O�A��oͯ���+��\�U��x��"O�q{bn�8W�`�2 1��q�"OF���P�'�@d��fܡ��0"OJ C1b,�u� &[�:0�!"O�\ђ]�R����ݺX�0��'	���m=2�c�G�T ִ�P̝j��0?��Ŷ6�.�q�`�r�1q��z�<�刏�G���C1��D�%�ԡ�N�<i�	���\`�tJʧJK��@��C�<�eś?
X���&�hHX��I{�<I�P��|�sV�S!$x��PC�v�<��Nз)�2��
$��x0��Sm�<y��W�!���i�m� 1���3��Lb�<���A��݅sy�4dNu�<�  ���2s�ہ,p~X����p�<��������J����[�%Jn�<I�ɒ�{��+��Q�v�,�"�f�<A�FBD4]�b�G�J�d���^x�<�G	jDhJ��_�0�
!�ՉP`�<����8����)00�1��^�<1D�35� ��N	�U�x%(��_V�<ɐ˒a��p
�A,���FU�<q@A�,5j}��k�����kF�N�<c+�	I�|�&�5O ��JG�<�R#SCyr��
�.��{u,@G�<qsN�5I:	0T�S�w	�b�E�<�tm	K�Cz������m�<i 	�hMn\�)��}��mP�� Q�<�f�ݾU��|iČ�j-f)���J�<��� �c $�y;FMQ��b�<Q�H�_üds�"���x��*Qy�<� ����G�%�z�&˔*)3��"Or`� �$�����קh �T�'Zў"~r@υ�����#�N&�k�/��xRfI54 \�Z�DL8����8d!��\�MV����&�'[Q@�h��	�[�!�B�YhB�)on<�Ї�	�!��۟{´���� G�M�F�}�!��E�\jWI<?�B%R$�w�!�$0B�$�2U�3���2��D�j��'�ў�>�bQI�#��$�bk�k���0&�1�O��D)KUVicfP:3���r���30���0?�AD���ң͔6Q\����d�<qD,����8�/0��{��a�<�1���a*\j'�Dގز�oI\�<yG� �����ʐB~f���M�<�sL�=p[~x���nGF���J�<qE動Q���`CBįE�4�r�Bx�\�'nh���:dP�0�oQ+"'fl;�'�F"��d�5���"�ЉH
�'|� #I?4��qViT�2��
�'Q��1�NY�'.`�Iu�I&=��
�'��t�v��*�֌g�C,ON�=E���J3|Yց
-R�L@�sQ��
��'!�Ojc>-[��͘X�~�¥�Q�N� �xbc*D�P����D~�t�R��j�ZS�Ƚ<Q	�(��i �L��!��S�p����1[@���enC����T��Q�����Ĭ)�� Kb��vl��ȓ,���C�-U��"�J'!�nj|`��b�=D	։z�� B�"�xh��'9ў�|�')��j�\4�wY�A�1���j�<�&H!���Y�cP�e�n<��_�<��]�>�pti
L�t<���\�<q�̔}�|��!�Q�dY���P�V�<�`�Y�$��X�� Y�Q�T)���y�<�U:[AXG,�4jP�	e�q������xR�� E���0�ŐF"�S�'/!�!:�2�7�H�a�̻o!�$H��h
�5^�~db�ϋ%X!�$��BZL�@�� Gւ�hg�g9!�\��
qYF˒�VT�i�L�5(!�Đ<���@ve)��ɐfG'P0!��$ >DJ��R�1,c�& /1.!�Ĭ��]ِ�
2'"�}��e�9D-R�)�](���j���K��-_���'"L���N���0 ���,N���'@��@��^�r�����B�ۮ�@	�'��k�j�"}Dȡp�ˊ�?�P:	�'1��B圊E"�r�lּ�'�F�g����I+Q�ۛI�~���'�Bm��dKL��l�`@�=g����"O��ൄ��}~tɲ��l��&"O2P� �,XŨ�� npb8(�"O�2�J�3"<	���ߌ3���B"O�m�"��`��C�����""O�]H�
د<'�!�w��4yt]�"Ox�$��X`�h�p@]Qt����"O��J
�6B��s���:����@"O8a�'��-@Tb=����r݂�"O䌛'@ �'���Rk@��X�"O��(Z�y|2�C�͗lհ��#"OؑH�(X(6�ڠX�Ѯ)\��H�"Oj󡗫g���Q�#�W �I�"ON���`�������!֯W�"U[�"O� b	��!�<cG�Xs�� ;G�>�"�"O��H�/�	z��M��΍$;�L��"O�ū�NP�z�@s�G�$�ָ+�"Ob�S� W�BT6�+��;%:��"O���0OhXK3��&ʾX)�"O�X�$ᒺ�(K���^���Y�"O�!K�.=���F�^�+m2M#"O��J���B�)3��+TW.iBu"O�H�fS�31���ɚ)NB�"OP�
F�Zu�c�U�X>T]{�"O�KN��F�(\K�J(A�V�A�"O`�@'�=�~��D��'%͆E[�"O~%r��ԑj:f�RLQ�t�b��%"O v+/7�!�ga_(+��d"O��H��Z5�������zh��@�"O>�r��{F%����,h�!�"O��BS Θ,�ѪO	]0�1�"O�B�IV���j��*K�:;W"O��f������I^���I2"O�,B�c�Y�4Ȓ�H]
����"O>���?Q��}�'��� �>�pD"O�� ��5���C�>dp0�"O`-+AA3��k�bL�\AB7"O���ˑ�^3���U�/�,pc@"O8��! �z�zhK���g�{�"O䕓��	�&����p>�q�"O�pb�	9brV`S���98ඌS�"OB�SvF
�q;TpZb�;`��R�"O(9�R�Y�:����@�����R"O<S��C�̺7�ך{|�T3�"O<Xfh�#OD�%�BL~�θ��"O:� 7�G�L��5K!� m@���"O䭋$_�t쩫 �U-8TZ��B"O9���_�������CQH�	'"OeJ��B�Y^�TM".2��q"O�`�%�O7Fº�ʗF��'6��"Of�2F.N�%`8�@V�
|;�բ&"O�m{�B��;�L]Kf�˝d~�! �"O��3֬T�*}�A�w2�S�"Oj0�gEȻ@2���-ĉGW���"OT\yfI�!�LlcU�$�6�G"O$q�tmP+Rh �#�R)дU�0"O�)bB�J�0���1 ���Р"O@�k�Q��!�5��H��,P�"Oxa� ���H��x�N��"O\��q�U�*d���b���}sJI��"O����Y2<8�c�ǐ�5e"pyp"O�i�d!K.\H9(�NWҘjP"Od��tg�!�|}��fJ�vv�9�c"O�X�cnU�e��ӄ�2VD��q"O*�ZsT�WHXYc��57(�q"O�=����/�RR�L�n��uB�"O������dlrmJ�@���("O�Q"�K�u���TFB�MB^}�7"O�ʄO�F��3�0B��iK�"O�06%ӿ��1��wt�)�"O���d,0�JE��X	TW�1��"O� �`�J�� iA'�	A�9�"O�����B!��V35 ��d"O(��Q�N�O��uhgd�.�X97"O�| ��6f����$�� �QV"O65{���bl*���R�l�|j�"O� V�xj2u�'��74���u"O�p����i�K�~o* @�"O� ��X ����0�¤J�XknM22"O�H��L��K�5r��ϘR�m��"Ot@82�$��TbH�tj���"O�II!H� V���J@�3�X�p�"O� +bE,k��ICŪ�6����c"O�P��L�K*�P�&���b�2"O�4���r��� �ʇ%R�p3"OV4�2O�Pre�TI��B�V`�"O�3SM(I6�
��I�{ޮ�)�"O�m�vbOj���H��ș=�y"OJ�G.�5p��eX�^E�^�8�"O���E^�|v̬��*[\���"OҘ�+&>����!])Ԝ��3"O���iΊ[ԌP���!�J�"OBA3S�ϩD;�%��(�^��u:"Om�R�����f�WE��e�'�����A�,46͙�B<�Zě�'��t����mi Ū��&�|�!�'����ĎZ@������a�'��U��H�(����gbű b���''�L��%�CT6���c�<t$��r�'��u��D�#Rɞ�C#O�ڀ���'�\pf�! ���RE�\#��{�',��B"̀W	ȥ�l&�RD)�'���Ar1�]�m����k�HC�Iu��ip� �1جZ��ݫ\WJB�I�Y5�x�p�Կ,vt����'4�C�	�o��C�n@�i�JLKg�Z�y C䉼:8ʩ�s+҃�$p����2A��C�	�-	����� �1��QB�g�PLB�	�(�賵�F���p�n�'^I B�IQ�  ��� L��Up��8��C��8`璄�Sퟃ>������Z� B�5L�<IB���0Y�����%4�C�>s����LPD)سH %g�C�	=%�d<:TN�
\�3�K:�hC�	L���!oa� �R��Tj%/8D� ��DlƼ��M��h:ը(D��9��O�a*L�Be(E=���'�$D�����O��b!Z��2JIH|z�j"D�4�C/F�I�.eMJ�u D��@�D��E(-�`I�.r��Bo<D��ka8t�H�X�$��lPf�5D���mM�C&0!�P�Ϟ9� \�@3D��@S���s�b�Z[�1�e�%D�����Y$���h�C�E����$D�$�b��L{�܊�M�����l$D��� ��F��Mࠏ�=<J 4l(D��������p�ț}�4�A�A,D�l�SiO%P���k6�!z 8��D?D�8�""��";�kGA�&r ����<D�$���9"��(�#&Z&t(T8V;D�<(	��>5��� Z-j��p�t�.D���c�E�H�`�C`��9r`���(D�x����>[��b�� �H)��1D�����O+-t�C�Ŷ;R"���/D��(!!��D���m��bm$l���.D���a/YfCԈ�v�ª-���pR�-D�R%��� �����C��+D���.}Քy�3�^Vɒ�(DJ=D���g�k��)IF��e6�9 �5D���@˞=?Q�4
=���4-.D�,9��[��k�! �v�铤>D��8@(��� 	�M�> 1�>D�� ���a�.j�d�3cV�b��{"O�5��IT��HS�٪ 2��"O`�i�߽#.��s���n��F"O�	"�+�'2���ТCۊl$��"O�Ȑ�g�g2�DI�bC�[����%"O���!ԉ���#�y��<�"Olܡ%J�����R��X�"O<l���-%vĲǟ�F�ʸ"O�thDɉ-�Jp1�F�-�:���"O��`0m�]�&�R�B��^�2Yw"O��"�;m{�(Y��B\�l�ٱ"O(���-^�̤!��b»4��Qc�"O�e�f��D�풠�ҭ�NIZ�"O0�f$G�7��`8��A6tbd:"OTLu�X6����
G>v��"O>Q���R�
,�Č͑02li�"OV����y	$�"���4K(�S�"O�g��0w��� b Ƙm5-`!�dC�>���a�c�v���#5��8H!�D��R�����
~��7��/1D!�$�S����%�`&l�@]�*�!�$����&�êQP2![�nA?L!�$� \���c��Lٌ1��-�TP!�D�9C�pl��IFŒ��t
�g!�dC�I��"�S9%I |�t�E�!�䞚DҺ 8VI�!)����B�{ۡ�$R;_@Аk �,|8`R�,B��y�� $��UrH��#v���b�"�y�jP��,TS1����������y�;.��l��˘�c� ����y�K�_m,��?~oXOY��yb��j\�Qkx�BU��?�yR�	ds��s�x� v�B���,�@�f��lT��G���]�ȓ:p��Ce}��H��
�5g���mЪ�a0S�l!�=�5ϒ)��$��k�b13����#���ArR�]WЌ�ȓIN`�S]��R�y�!��"<��ȓg"�QP�_{�:��Z c|�I��1����퀘tʌ�9EÑ$"�����Z7D�j2 �=��q�s�I�І�#�0��4���)���1tx����0D��`�(!3�Ͱh|� ��b\B)h�C̈q�hە1�Hu�ȓ)�>��������%�ټ ��:�p:�̕!o1�!Y%Ǝ5u�ȆȓGt�x����i�е8v��"@۲H��O��ii'�\9kMvp��Z��)��r(�H��M۟
�n����.�֥�ȓt���V@�/tM�=�J.u����&��)�=u#�l�T M$>P��dU��*�.\/�g��b�
D��`|�"+�-��]he�y�<�f股K��	tF�5A|H,@A�<I�n	;a��	
���_�x�˰�z�<���K�#6P�Q�N�G��ܪ��B{�<�ե��W�zh�m@�RZ���M�y�<��-�X�|H�hN�	J�J�n�w�<y�f�Lw�$H��ցT�n<x����<Q��Y25���-]RXa6�}�<�� }���S���!�T���T}�<��FG�8�Э@V���S��x�D�<yĠ@�U0p1�LK�&r���<a�G�
l���F�M<����@W�<� Ș�%O�1�2��J�d!�J�"O�a�Gh �+� �a�+ڳ��}34"OT��(I�� ��^ %���"Ob�Q��OO���*��|�"O8�H���:�-$Q|�)�Q"O,A�s�'5��p��ߔs�ժ "O����P��JLQC���}~ $A�"Or-�� ;P^�%Z�BP���H�"OF��E¤(#�T��∳o(tP�"O�B ΍�(X ��--��a��"O��i�e@>�P�ӄ�ө?���"O�mk�/��Ц�`D�U��Ȉ'"Oм�2���q�V,!MM(� �#%"Ot���Ҍ9.��� M݅�.�V"O&����NB�}`�KӱQ��,X"O�̻ �FN��@i4��
V��$�"OhAe-^;]E��t�\2a��8�$"O�(j��F�u�d�����H�����"OL�Q��
1S���t%�@�v"O�`��K�\�����?Z6��"OD6&@_&�q�&a�J�ހA�#D������$H�"�ڒ�Ûl���;ä#D�@��'0~�f��s퀷&��A��,D�䋒�,��xsi��|��L*D��{�~gAb��s���@�(D�x@]J�}�%�L�K�z5sQ�$D����(�$�֠���?q�P�t�5D�q*^�$�f\��F�[�H��W@4D� �6��8r<$��çM�F��c%-D��(0 �aH�|[�MI.Q�U%-D��IB厖V�(b�߉$d:ժ D�آ��sְ�ꈵ+���g?D�(�'&4.*�A���7H;U�t�=D�$���B�f8�p��Ɂ1��<H��%D�s�K��A@���AӖr�L<��#D�$�q A�9qj\��A�:El���� D�@@�)
�*��%����
5U8���<D���1蛫^؆u�����u��!@�<D�ㅣԵam"�R���Z���P�K7D�xa1
E�/�l�֢u0dU)�+D��ؖ��?TO�U ���[�Ny��
(D� �Ue��3{ X�A�T1/{	�*D� ����|���
վW4�;�J)D� �f��5DO�:�T�XvB�D2!�(rWl�C��S
I8h�����]!!����iBU@���E�(!�#4��n�8o0>C�II+�!�dG�SӬ<ڲ�I����Ʌ*X�!�ՖC�p���Xjl�8r^)>�!�d�I�Ҩcゅ2Y2�R�Q�o{!�D�#������t���:A�!�B�{��#�OF-
�1X���"4�!�D�0�|̠�΋�h�X2�L<�!�D)(*<��V���a�vZ0�h�!�D�d`�!�CP?���Psk��!�d1lոA@D��:R���� 	!�D�;�d5���Z|X��l���!�ͧ&	���!�Ѝ �N}!�+Q"P�!�D�3��QP'�"�.��b˔2|!�D�<�����`���Dv���"�"O��F� #�$91*�����iq"O(�&�9W�6�3��D?�bq"OxL�'���j�n�����ڭ�p"O�Ik�'��(.��᧋�c ����"O� 4���@����hg��]���s"ON`��K�X��ĉ �0���"OL\`6�'@*�e�%��$wl��"OD�d�(_"P���>c���#"O&8Q��.JF��$@+5Q�ؑ�"O$��j�.Y��
��F-R�b|�"O���Aa&dBҏ,_�V,��"Oh����\������6&��Zp"OX����Prʅvm��
��h�"O� ���$Qܙ.�&���QB"O�ty�D�5. d`�M�5C��"O���� �=P��m�v�� ��!R"O�����*��]	@�X�M "O\r@HW�!����E,[��"O�!j�:2j4�s��  ��`"O����7rY�P���?��80"ON8�U$ȇ����� ��w�֘"W"O�ph�o[��|��c��(v�|��"O�$�Њ��Ȗ(�*c�� {�"O�٘�*� ���P�f���4"O�}:�㊕*%v�K�O�z��]14"O�������Ua�)��.Diu"O�����W����`_�^�M,�y�I�.J�@E��뙰�2�;o�	�y"l�12j�A "l12�\��y2�Q�t'D���8o��� ���y�Y�
��8��gP"T���AA!J��yR��;,W��IR�No��%�߬�y����fĘ�, �o�d1�C��y҇�
d�ܨ��R%c0���ı�yBƏN�D}3��C�]�0d���8�yB
�~
��P���=_���Y�$�,�y��V�aH�9o�.T�*4�����yS�1�a�rO��4�VP�ް�y�AM�/���F��d�
����y�h�c�tDH��Ԙnv:���@Ώ�yጡ
���(��<>�
q���� �yKҷ�(Z�́:^p���Q�y���K? ��a�.3�J�A"O��y��JK�,����1{@�2!�\��y�G�最�, d�ە�	�yr*Z�N�V�O=u�,��*
�y®H�&�6P�qeڜvK�2ׄL��yb��*O �C뚆o�\�#v\��y�/��w�1Z`�G*�L�5m^�y�M.���Q��0�R��4"E�y���;Au��xà�p��R�Ø�yb YQ�h�򯓓�^%c"�?�y2��0h|�L[7f�D}n<)g��y"eܵU:�Q��(-Q��:�^7�y��� ���!�դ{PB��rNI<�y2� �,8XE����,$ I2A*�yRN�$k���ă;o���TϘ��y��2(��X��6����cѼ�yj_�I����h �b���cT`�y��ש0����@�˜T#�I�⪒)�y�%��>�����l${@h���܍�y�&�S<��O�v���J�ܛ�y�*� �V���g?�=��M%�y�&ŮB�`T��L7M�����y���1�>��8�6�	�+�y"�T74��g��DP�� �y"n?+��� �3]y��B�T�y��01tˢ�ЇV�8q�ᅒ�y
� �u�V�@2�Y
��2�h��"Od��q�ހ(��a�������b"OXT�>j��S������#"O�yw�[�2��p�������R�"O�9�1f�*T�h]�e�O�}�)�"O��4O�2�H5��D�~CҔ�U"Ox����77;�-�#Џ��sF"OXٙ��
��E�r#R4av���4"O9h3� ���{e,x�Ó"OU�) n]ʬ��j�7Q^>u"O�țǊk����iج`Dz]�"O�:�(ׇH&2		q��/:@�%PQ"OX��'۠#(v�2	Vn-H�h�"O�<�U�E6N3�"F/a� ��"O�}`&�ʧ �����_�
}
%k�"Oh����`�ڨQb�,zw
��6"O>a��e�	jE`\��c�xm�T�D"O�)��&%)�U���Fp����"O�i��*�H|`$�G��h��"O�=��M-��zfB>�t�"r"O���H�3jkjܰa�#c�L�+b"Ov(C�/55�L��AW�@*�"O��r����ry�c�� ;{�1�b"O�D��I�%O�b]"5F�l�ݐ!"Ov!�6@۫d ����m��欤�"O2���ꍥ4:�qM�E����	�'�RTːՖX���[�R�!*� ��'��9rԉ,�%D�j���'���ՀԄ 
�TJ �[��i[�'�T������:��$�#̒B�)�
�'�� �֬Y"�8\X���<�,��
�'�P�����,0d	��'f���'�v���b�*Q�ޘzC�9)n���'�������(6�X��M[=��'��8�G �0]�"PMl�}��'�$���Ʌ?;*�B�!�8>:8�'
F�G�� ���ѡ� 6�d�
�'�ĈU�+*��ʡ�E,|�
�'\<a�"�#h�$��ԃ=��r
�'���C�>�Q0h���1��'�h�`W@ �),~(�4l�.�xx)�'D��i�N}3jQa �,0NRb	�'0D���V�%K00�&��l��'���2�Y�,^$�����͈�'g�)wcY@�� �G��s^���'���"� H�,	�9)�AKJDx�
�'�x����/,x>�m�9Yo0\�
�'���bWBՍ�^;�fƋO��	`�'����D'P4�X�E\+Ա�'yJXc�	2G�$�CG�Q�j�Z�'�h8�nU�n\z$�OؖYI��'(�Li�EK�kf�9)2āS�p��'�ҍ�B�4����f%}�$8�
�'��`q!�1}���r�
ͷr��z�'�z��񮕔_�,U����*8�\��'.��&�[�3�� ���.-+v!*�'d����˒�,�$���k�
&�(��'CX���#s9���M��z%��'�I[�b�M]�ڡC����@8
�'(Rq���ڤ��@t[ Ubt�B�'Ð)��oŉ�5��.�Z���',��� �:�.���Q7<�Q�'��jp�N!3��{���JW PA�'�z5Ί�MhZ�Q�/�J�hѲ
��� 2��7?�=a&���}��"O
�'&
0?(��ӭ�)i�h@"O���(Ϸ4�A�4�B�Ѕȓ9Ѫ���K,fѰ�{�$t����ȓ�S��=8U�n*/K�}�ȓ.�ƽ�Dh_�3�X$2��D(`�b���J�2	a�E�UHLHz���"y�@�ȓm'���քxUډV�˜'"8�ȓ��%��`=��	�lR�7#2��ȓsH���a�\�T,�vEY����)ā��T�����yj0P��S.���	�'}��p�`��� �x�ȓ~��"4�I'D~H̸����"4�ȓ!�����*� @��q+�4�F���$VBG)��p� 'X�B�ȇ��\����ܱ�B�xիRLV�1��l��4`�:R������A=֡���Z�9d��C�
9�"�ŧ�z���tp�
'�L�O�6���� =6u�ȓ@��=з�ٹL/V��"��G��Ѕȓk@
��e��e`3�G^�Đ�':B�ѡc��{Sv@j���.e�q�'^(р6�O-�hE�Җy�"!B�'ܽ@-�<��i��G�w�`�'��x����$IG���n\�m���C�'�TԈ�H�mNJ��@S��uS�'��$[u'S)q[B��!��@W�l��'4��2J�xhz��V�=����
�'Ɍ�is�	%"VѰ׎�HlDI�'BtZf⑻p��zB�Qdԓ
�'�nѹ0��5D,�phG��>	L`0j
�'|��:��ɼ�#�������
�'r8<Id%� e�]I�9����	�'���iCǐ�=߈���C������'^��X�3z�iks��2y�Xh`�'hw��!\�#��C�s�vJ�'��%���N/3�	�u(�
!g�e��'Ÿ�{c�W#�i�.F�1�'��C�H�)`$HE� �
�'o�Y�L�%�:��9�\ݱ	�'B�h�T�* �ZC���.�V��'��M�����%�T�{&��]Nm��',yէ�	m��2�F�
� ��'���6lM ��)G�"q4`�h�'�������U��0�V���- ��'�� j��|�~U*a�� �����'j$�*���8����@S�l/��H�'x�|a�X�{+�����
�7��'���Ґ�$T�<I�wJ\<'�x�	�'�R�`/ءR�:ˣg�?zUJ�'\dp��P� hұ�"��236L��'�0��@£#}�l�w�T��)��'�������_Ԋ,+6JP�E�^y"�'��E�Ul��k�z`��/�Dp����'�N�j�#@W��`iS()��C�'n���B\�N(x�F/+�����'�@A��i�NK�Y���
���
�'�V%��e��}��4�iA0E0�	�'z�9BT��9{�l���;g�b]��'%�A�a�+`d8�è�X��ai	�'j����)P.�P�I�R�;�8�+�'(|YGAJ�4$��)��H,	�Ā�'���8q*� ��͒���Pْ���'��:⦂SI���"H������� v���k܉H�H9 �J�0qM��"O2��PAˈ̸���AQ�t5��"O\0��W�K�0&�)���8""O2�S��Y��D�gj�u�օ�c"O�	�eA��V�fщը߆HF���"O�h"����,ܖ�`��*K�	��"O~t���FA�Y�G�Y�p!��"O�!R6iB�>��pC�|����"O�(���1�8`rFٳ���Z�"O�0BC�k�*@��M���|B"O6��7��G�����m�3~��P�t"Oޠ��A:eȶ�:�k<<���"O,�0�#!8��T!/0���*`"O<:��Z.m�B���픝�FԲ�"Oh��/!
FĨMҺy�:M��"OBD�!S2A���Ԋ�[��lZ�"O���&��,�B] H��~j|X�"O�I9",^'g���3FgN�4u:�h�"Oz8�W���}����Ca�2�`�"O�����N�P�µ���'�!A�"O:�( �;�XP'�۞-�ȑ5"O\�I�!'`�TbtC�1��AD"OdM��JD�h�H�A���~��Y�$"OnIh�#��7���� ����0�q"O����E߿��
Fc�x ��"O��RVHQhJصz�B��	�0-�"O�I��g^,��%AǸ� L��"O��i s�,iÃ����~�"O4"���H���.�
~��JS"O�]��꛰tGT�pȖ�)w@��"Oh��5F�.7$Y0(�$Vp�}��"O�9w��1��BW��ɻ�"OZYIŉ��#����D�Y�X�B�"O�I��l�9���q' P�֑w"OJ��j�,Ř�K��Hi�&8a�"O��zs�U.s��1�o�1=|��A�"ON���T�G�����LT��B�"O���Ub�$~M�&��:J�z3"O\Yg[p����L��=5�a�"O���� �&#VH�h�D�gO�$�7"O��CԬ�� �P�"a�?k4��a"Ox,��/��w��Ȑ�[�F��+"Oʩ�7Vc���V��1W"O2IZ�.�~���[e�������"O`t�'G�	3����`�«l�v"O$�3&�U�ilD{�� �E�4��"Of�����}Dذ�d�(��	�"O�U ����R��[�S�&�`A"O d�V���+E(�����}����"OҬ@��,s`�!�W��R���"O
� ,����Ƭ��qa"Oj��"!9WN*\����23ú5�'"O�-eE��l�A�h�87��`�"O����B��R�z���#)���V"Ob,��ݘ'�)�Qg�i�x�y"O�%�P�&��(0����R�F�I6"O��jf���>��Y�K�,Ǯ��u"O���3��m�E���p���9"O*�㖯׵)F>tQ�"B'x4hb"O� "���.S��hW�@�x,��U"O()�P�h�VAS��:V˜�#�"O�-(�ǌ�d�"�Q�^�Q�"D�&�8�v,J��;vQ�B.?D���D��W�l�R��[�z}H�u�<D�� �Q!�%[�${"����O9�����"Oz���T=o��]J���4C��h�c"O�0vY�f����Ă+��@u"O����F}�� I�8
�)q�d%LOX�x#=N�X�f*q�mr�"O8��¥J/y���$�v�R��B�44������;U����3
������>1��d\���'߼U�PAY&(�T���k�*F�a��'�,D�O�J�]��,�X�Jl�H<a�O����3l��sBA�%&�Ls�
!}�!�DN8/Jr��p@�N$̻�j�
����6@�c!O�sH(3gǒ
���d0�IzVX�ӗoA%v
��ڶ��
��7D�|#���'�"��䬟�b��s� �	u����Q��+G!��S�ĉ�C�R��C�/�ݘ-�`s��%eΣ=	�2�nuX@�4Y{�D�Ru��XH
a# �Q-XEr����w0���eF��_*��q�l�� ӄ0��83�Y�f��l�6�QP���nh�ȓ4U05��ߝq�l��@��\]�ȓ�N�x$'	�X�J�̹<��̇�$*&y��An,qJ�h7(q~�̓�hO?�hǃ�4.Z�� mS7V��i��*D�(!@.��z_�T�q�0p���)D��b��O >�N��U��G���U�(4� 0GA�}��I���]�)sÀ�e�<ap'\?m
�;�m*5��!kCOM_�J���O!�`�!X��ʁ��D� ��
�'��R5����p��`��2w�����4u��'���~�'���"�Bko�� ��3G9�hBד+�qOL��Ӎ�M��ˢ�
\m��"O�bW%�1"����t�	y�dID���Q���'V}�,�#���t$����L�����Jtĥ�񈆙_�B蒁�Z<mm��E{bR�LExRJO�6`06�θm����-N(=!�͙Q��|�g4�qa��>\'!��	!B1��Y��B�"\��!�_�%�Fu�͆�}�T+��Q��I\x��j6�ϩ��a"���m `}�"�!D���!<������-t�x�[�A!D����˕aF ��Q���Pxb)���=D�t+�eN�?k�@�"l��A8�<*�.D�LJ蟓iW��󡇋d��4��K-D��x��ۚ0�$���J�'>=�Ё��,D����� #p���h�R��Uc5��<��D%L��eKȟ,_�a�E�^2�b����m~�S�2�Ⱥ1�	�250����yҍ��~m,� �Nx4�)vD�0�yr��+�ز3���^�胵쐆�y�BB+��)Q�=b�6��A�O��y��)��n?�S+e,���ň+6���X���B�<ID�
 ,V�:�+j�� H�%�̓���8�SZ��F'�H�S�E%t�>��%�IE�h&�� DeV�(t�؀��~��P#� ?9����'7�O(��AX(�ꠉ"ς<_Վ��ҟ|��|�>=��|P�⟮���R"��<PӺ˓�0?����R�^��E���%��| lx�'/�<)�R>�"1�ΐa��q&�۠V���#�7D�� �S0*9��	��13�}Hg��O���$E�`4���	ԋB��P#^+Da{��$��w򬹗˸J��=��BX�3!���(�M)�&L�y��m�g��4!�$?;j�Y��
�[*�(�c`\	�!�� 6�b���,p\�ݡ�@U�` )[R�'ў�sd�/*B��7mAs¶C��-D�\r���<���K��]������>��hO��b�b�i���	��������*7����:?��5;G�y뱉1 �]z5��̦Y��'qO?7�2��(���Xb���H�,y�ў���ӟJV`���(��ɺ�ꂞK�˓��} -[���6��8sw��`��HO$��DG9Q��#Ȫ_4��Q Dw!�P!5�b	c�@�R�������(0�!�$�4,�����P�l:��!��d_DD�`�Q�W�D�z%��h�!򤈷5$�dI��ɟt������-9���4F{���̢��2LF|����1�1:�"OH��K̉[ټ=0r 9K-�+��i�ў"~n/]l��4F�\Šd�����E"O��X��Z�:`��4#��j�Xa$�OҹEz����Q���a�
��$ҲAS#3L!�DD�{���`���Cz4�e�S-$?r^�HcI>������A�֝ ���@+�Z�!��!��E�lR��^6x%��#��ݍ?�!�$�	m��l�
�4�l�����!��( �ᆏS�[8�@VM8%�!�d�����saô82<�*`��3�"O��ԧX�NZ�`hݧ�x$"O�"��@r�e�FO�1��1��"O����@�1���#����� �"O$�
��HaH^�qF�ڜT�\= �"O�4jD�܎���SP���:͒TA�"O�Eޗ>A���"�DM����s"OP9����`�gX��Z�j���Ą�	%Y�~ ��HX>s��LPӦ���Z�Ir�����ղV9{�@�V��4����1�S��y���v����E�,t��@u��4���=�O��z� G��&HS3D ���pӵi����,+r6�J�cV�"���%W�/@!��h^���R'��x��	�׊U ?ax��	&=����vo������ȗ�xU���p?7�Ґ9�f\��l/�ڈ2�Ms~��)�'45\�.v6(�b%G�x�XH�#6D������X|��pk�c' a$)!�D;�O�Q��� ud�$ΙO�<����?�O�O���$ɄQ̌�#e�,;��#?OJ�=��X�'X�ي���ނ$�&E]�|[R���'��6l�:\>nܳM�*~��'l��F�+:��q #.Կ~�����'���k�e�=f����P��46�-�o7D��c.�=M0�t(qHL�u�eQQL7D�����6b3���KH=5�p1��1D��"BƦf\� b�K����4k0�D�<|����3�أ&˪,1w%H�}���CoW�Bw!�Ʋl����!�4��	#��8zF��<y�)1J�V-P"K�"�z1�QyL��ȓ��@�0a��:�Ё�hǔs����c�&ģC�c�Z��d� ޾��=a��'}��aCH�7.��3UWn�~�	�'2Ƙ`�K� ��鱧$@\C���E�<�H���y(M�� �6�r/M@�<��EƄV�5S��ȿL��7 JA�<A��~t�İre��%�v��S�DX�<!aKɧm����2,>���
X�<����)B�P&��\��|#G
T�<a���g�fy��)DBlB��K�N�<����*9�a���0{b=A!�� ��àU&J���ɘ8����"O��u�]"��"ZHЬ�
�"O���V�C;�xIC�VQTv-��"O�\4��c��4`(IV���"O&�ڷ�H�,p�Pf�:�:q"O��
�G�x��fdI7�f� "Ol+��K�%�$�`�)[
��"O�`��qk�X2r�6���A"Ox	��7{���'��C��Ss"O�L"��҉Q����D��(+(�+�"Ol� �A��9\���$+�Hsg"O8u	 Fn�x0�Cٔ0��H
!"Of�[1�L�I�M��a�6���"O�$j��ߺ<�4ـ�[��^���"O*�̃�PQJ@ G+㠨)�"O�<rq��j���hB�W8ZA��9�"O���Cg��g�b���E5�E:'"O�4c���>S�d�г�H5ܪ%�5"O���r�(op�E2�#�`�!g"OxLѓ!�1;,r�ɐ���1RxA�"O���ٗu�z�
�c�&&�u�`"O.H؄;%�Y��BU�O@��p"O4�#���"�@;�JƸ�\�P�"O&�@D�Aɬt�J]"4��"O�b�dߩ'4��*JJ�W0�3"O,�
�^�P5�IT��e�E"O��[� �}�2���v�� ��"OԤ�3V��0Y�2g|��9�"OH�S�oD�l��Hz���.0�2t"OnP4���d����S�	�Q�T"O�D��2R�V��T�A nBn$�5"O��5�^)#�x���:6@�+W"O��;���M(��6kH�h? M�w"O��8��ސom8:Eɕ*=�V8�y��3S� ��B�/9�԰�����yB�k���ua�(/ͼ|�QOQ�y���H;\!u��5.�(��!���y��[:o��D�֥;Q�>T����yb�#z� �T.ZA�c�S��y�b�!R��� ��O�=�rC� �y��pI�9J�}eK��,w�(C�ɻ��-�d���m���Q�ɀI�lB�-#�|���CnP�weC��?��\����
mą��CA�f�^B��*h��-�"o��-����)�B�ɩ3мk���	P� ԉ�)�
I�C�	c��U���D�F�(1��%qM�B�I�G�>!�e\�8�\����5^ϦC�ɨA����ٗ �`!"�I
b�XC�ɒ�p����]:���P��F�"C�	�$N���,_��`���-JW�B��)D}� �?$X;��O��B�ɥuc�Pcի)`W�Hb��B�	�R��D��� 8��dy��X� C�Ɋ)�6�cw&��y�(�rG�=o�C�I�A5�xY��M�b�2�a%P�B�r��UB��¢k�l���V7sb�B�I�x�98&@��v�1�G�gg�B�	*ْM�g�F�A#6���R>RՔB�	�P�64��3ȴ(�d��7<�B�I�?����L3mxމ�Qn��-LrB��7Ns�\P��*hm�Mq�](Y8>B��`�H	�G܈g�j�)�-�(S�B�ɑI��u�зy(�A�
�B�)� ��å׏4�P��ֱ���0"O���a� 2U	$`:��!G ��@O���A���G��c���@@ۀ��� 	�'���@�Ph��փ"zi�0��D�'JRT�ak;�S�9 �X۳
,**| ���p�nB䉫~8�#%�>��A���	G8T�(���P�d�#�LҧH�x���ŝ�*mJ�4%������"O�q��"��S�:��'E�	?�2,���?}��
�t�M')���޺?��Җ�zB �@J@�ga�lB�psN�J牜�Q�%�%�[#E
R]Z���q��!����F](UxvB�(��e���U�,'T"?�IB�}�hFn+��_�]'�I#W��3>��enJ�I!�D]�A�x{�d�?�3�6j
�I#%�<�� ���S�O-:)$n	 R�Ј�d��+
a��'k��C���)O�գԮG�r�)���>�i]��c���}��̓l.��2��-5,֭�����?�����6�0L��]<�s�,��~�sC�S.�����ݹE�b5�.��v�XKP J.�џ<�� �;~�5�|��V=5U�ٱ@5~�2��"�Q�<��C 8�$�j
R;	E���q�d~�B��w��=E�ԋ��l���A_&ma�����y�N�&<��GÈ0ds�}�� ũ�y���#�����fӖY"1�ސ�y"(g*(��3 �4$����h[��y���Pɺk��\�,*�	��L4�yB��61ʨu�Cj�� TeP��yRL��nd��Z�gʈ�cJנ�y�I��@�"�!ɴ98���K]8�ycO=t\��M6̈b&W��yre�*��a�+.0�u)����xb%U*��f���vZ
��W��b�N_k(<����
�z�����4v8��`&�z�'v,��Q��3_�1�N�@�c�^}zWLQQ\uRa"OȁC@������l�)+(����V��ؗ�U�d@MQ�?O)��	_K���C@_�yoN�tk
>o!��ݩfJ��	�H�1AH�px���<Og�7m�1=��I
� �ڇi,��d��'F�Vˀv\`Z'�ŜVa�`
�zC��b�ܭ�� G�Fjh����>+�ꘅ��:I��������*�*�%MQ�"?	E�7�h؀�m5��ٛedT$S�o6W ̳4*M�B"Onѵ��5�PQ�S��*f�NP��P�����˟$�B-3T�>E�D˗!(e��!P���;����yr���z�2�SJ��r�b�ot�/?�źe�2!���''�W�:m��I�D`�?Ԧl��
:�OZI�m��th��ٶ��u-���D�Q�zp2<s�����?�S�Ìq��K�َ ��a0`Cp�'2�s���p��c�C�N�'d/",�Y�$���jp����"O䅓� ʞ)�P�3砜�4�0��j�8+���2,E;r��览���q��lH�[� ��Ӯ 6J�(�ȓ^�ꘋ�%P�K�ʤ� ��w�����i]
���.L;>	�i>y)�R�1���?)؅�9��ܐ�
ύ	��Q�6LOl@h�GF�B� �7�A�QyC�;
����� �]p��.t���0��\. ��E' ^y�O~z�П|RC̱Wj�;���	1�9�!��I+f�C���#G
r�i��c��_�F��(Lu��CNU�uW����/�.6 0$�|��#uj��f��	ay�H��q�hhش��N��ɲ��ӦP�qxN>6�<[�`��J!�
����>��֟<�{�a="d0����l�&H�e3�~�)��UG�yx�#2	��(�Nj��'�X�r1��=�\?m���!r�):)���/V��!��],o5�y9��d+8�dp����q���pf%L��uI�9ʞ6e�	^9b�\#eg�N��@Q� S��=��|
��)�O^��GB^oc���/�MS�U��Q&�6GX�����䅀��~j��*#���-P)T6. tnB�i��(* .��R��I q}{e��say2
^�H9�%��7���WN_�Vi�0�U/T�"^��F0w��ٛP�&���Jd�h?q��FBsk�G�� ���E8}��/n����idő .G�(�=c���h;�0�V"�j컂��3'�Z�����q��~Z�:��*� �@��l�%2q+�̖U����I�3��`d���Y;\�
/�p`hN S�I;�쐺���:�3O��a%\�3��ېI�<�'r��<L>�e
��
-
l���K�(�B-��Oy�-϶,��4:�H̺?Q>����)Y��q���6��Т�g\Z��키�>�e�O�3���L#Mt}³gŞ>fֽ�`�A��OԵ�0M��1�1O��#C/�" y�5E��.�����
O晱'��?m�^�QD��">�@�/�%:�.���'��<�1�J�����a$�h��A�	�'��XX���\�]�aa��M/�y�˜�hq�A��z��飲�Z��y���w�q9�O�|�)��H��y�Ɠ��A�q�Nw���H6f���y�Ei<������2��� R�/�yb☂DYX'D�-�������yr�Q70��q�l_Jة�$U/�y�f �m4R���l(fMw㛃��/�RȒ�&<O�Hg`\����,��n����'�lqڳ&��x�3q�_��2��BQ}r�����Wy(<�6I��Ǯ|%k
�u5�ak�gI�'�J|���^�aS���%�z�S#J�,�ۂ�ݼ!;�LCE���4B�	,c�(�`��z����G�<Bu��j���`����~߭>�
���O��RѤ��0��
�,Ǩ�"�"Ov�0F@5r��LX��V�����W��P;g/��v.bi��n��yt��	E��IIe�D	�@��_5����$�"}��� $�� x�I��(���ٞ�의$S���I��H��dk�G��6ű6"�$!`�0.$Α��n�0"�I���#KF�OP҄�U囉=��`�6e��Q���	�'<~a)�p��e�3L���W�1���Yg`�"_��-�T,��h�F扽6@�@s�̏�"�b�@S�*B��i�%#�H�7"�YQ��X� N"x�&��2��]k���#�C`�⟪)G{��5r���*��s��	��>��=1ׯߑm���#e&W6�Х��n�%���곩e-����N\��H@��j?�O.̑��I�i�`�����V�0x��D�-U�|ȓ!Lݶ��CeA?��qટ( ��nI12Xɂ�o�7�<�`a"O�aA�� ���5�ޫh�4M��N�69� .F�t�z¯ԶT���z�M+�'�y)ƣ��F��,�&%k�-xEB䉃r�F����o�X�f#�78�,H�T�U���f��k:$U�K�D�ɉ�$�- �0O�vZ ��@� �Q���i��,�ɝ˸	$Mc������_C:hT�R_�<�#���	�,���� D�a}B�ڀ���d�u&� ���M5�� �=N�ɒ=B>Ɉ��=�.y��)�"5�[�yW �oH"M�G�)hۜ ����y"��� ���Y㯏6s��1"҈����e ��Z2��P[W)��!�V ��� ���a�O�q�����ɐ)P0>�����7!"t�Pao��x3BB�|p�갹i��e��G���A��Z��\7K��0D�)X�M��	������K�t\�9�f���4����W��O:h�Aj�㶨c,O�Y����*MYh���A�6u\eYt��Cs�4�bꙫRlLqs���0?!W�͓T��8��C#N�t� G�pB�1�K�<�Ɇ挴Y���7z�i�Y?�̻,p8P N�i�0�Y���$A�`D�ȓgf��¥E�#��h��g�-I�p�	+(YJH@2*�|$�'Q������.8���Da�(}f�Z�d�:��`�g�'J��ც�$~�Lm�n_������O򒭈�a�}�O�!S+����<q#CW�:��/��U�j�;aHF��r%������6#}Rp�D�'l}�Յ��%D�>�B�I6
�V`S��?�8�b���yz�`���E�G^T	%�"~�g׌���*@&�Aa�%!j1��ȓ`��I���E 0�	Y��D%{1�-�� o(�Ot���^�\�lx�۩��x��"O��b4�G�O�t`펇�`P
�"O�	��cD3�Ne�a�ư"�Hѣ�"O��K�B�C���C	ӺWȄ ��"O������B��3G�1U"��W"O����M�;�bQ�'ƫ)^գ�"O$h��A8X��K�'ܲb:�a�"O��s��_�g��Tf����"O� ٠��2Z��L�5�ؐz"O՚�Q�~q,�h�#��AD��"O� �A�uY,M�RB�%A�l��"Ou�C-�����`�R2/:���'�����2n���D�ײ��"O:�IRg�Vݤ\�PgM�0�N���"O>Ŋ��4e��L�Uf�B��5�0"O��T �<p�,�rFU��`uJ"O�M m��Q���)��łH2�M@S"O�|��U�qƽ�q�>,�A��"O<�5	Y�L��DI����ld:�"Oĸ��V(�TyZu)�&f�pA�"O.l��F�[d��������Ba�"Oz�yw.� ?�FI8 '�G�4�!�"O�I�P�ѓ8cp�1�� ��92U"O^x!@�Rsď�g�n�J&"O�0�mZ�O��-3ӮY�yx�s�"O�Uӥj��p�|`���"�r���"OV� ��	v�*\@ʒ7�쑒�"Oֹ·9�<��R��)TАy"O!I
�8C����mB�C��"O����.o"@T0$��n���)�"O��C�@�+U�.X�H�~cn��"OAĝ>8���!ǥ��|���0c"O���K��r_Z����
�e� ��"O�s"/EF^d#!����A��"O��ؐe��&�.,�S��:0�4���"O�8aL���
�xq	�b��y�"Oz��B�ٝH}V$#�8�i�v"Ox�Eǒ�l�z1��B��ȱ�"O�U��!��|z���gRLtι��"OP��C&�8a_�\)PfΘV
2���"O��z0Jr���3��ĜG*�;%"Oh��!�͌ZU2u�T�ӭ!�l峧"OTh�1K��N��z�	ƾJ���"O�XGG��Y����UN�I�.]b�"OZiB��B�D&��H���Q�3�!�NZjYC�� B�,@`G�0<�!�$΂/d�`��#���20�;�!�D��e(e�S�5�"�z�k�#�!�d՟S���#�N8o���Q)
�!�M:QV�}��� P<T��HN%O�!��P-Qw�pT
��O2�Ibeʊk�!�8R� �?-dճ��#�!�$��z� ��ŝChT9bʲ)�!�D� !0T;�H�<O��m`D���:�!���<�4L��b��&�v����g!�dV�>^Re[�Θ�{�-:C,
<�!�dF����襣R�)n����
	�!�dI>G�$ܫq��+TL��
dI�s�!�$��q��I��\_ �rUjw�!�0 �F�{G�R=��;��S�M�!�^�
�ak�eϖV�~�F�ĒT�!��8c�uig.Sx��0�痹 �!�D['A�\dc$@X�r�]�I%!��9a���` *O��Ȗ !�$�9��Ԍ�:�墡�8.!�$�>bynD�s	Вt��KBǋv�!�$/�
8��X�Yi��Y9P�!�_�-H@G��i�D+�	AF!��ɂf�T ��Pr��9�g�T!��w���b�˓s�S��m!�,<� b'A �v @�L�P�!�Dזtx<+�+�)~�ԝ���ڗ]�!�� �
�DĴ
G��ɑL�{��)��"O�M�3�i L�2��	u�B}`2"O�=16$֋	�,��._4[�^��"OU�� ��:�څ��m�&L�,x8F"O��d�
o!fL1�kȩj��U�"OtP���B�w���W+�*[+H�x�OvX��" @����)��� }�4��86�	�'�4=�]�R4��I���$����OlMx`�5,-&c>��T/<R�|��ݔb� ����?D��k@��PuԼ:Ԃ�i����2F�>��FU �>T�W/}�����9��ɀ��TP8b˜�!�F�q砘Q���#
���J�ɋ3<�d�'rY�5Hc~f��Oޡ8�K�*_�� �&��4���';j��h�@^�]��D�8&�ID����X�[u���*�o�+d������2RI��&�N:p��ԍ]���pp''B��(�L\�rȥ�`"OzE�Ū�$  `i���Ζ@a��� Q�)qZ�jx�"3�>E��dɡ�h��uF��f;B	r��O�yR�͓S�t1��
0
���X�-�%|��a4}��Z�H����'U��C�Y� �d	k�48�Š<B�δ�r`�D��cɆYF!H�1��Tcq'�O�`h�ذ RX @ƌ�������c�\I�@Ys�' ����H8y勛94��Յ�Q�(q��)hv� t��0m���'���a�g�S�O�@l��l��6� �a|���
�'����4P�8ٲ��%f�n�<��LK�j<�KG!��V��<Z��Nj�<)B˗O䖨B�ٍ_m�"�X�<�1�:2����O��G� 3�M,D�d���J�L�\���C�d�j�0��,D�`s��";Hp� �*2�a7�-D�<ҲeĔ2�^�RP�C#(��(D�h�pJ�=�XI���=h6�c#D�Xy���S�ܠ��]�%:����-�\i����tT��ru/]~$b̓���b� [W
OH3���N�.�"`��? ��59�I��0�����i̧I�����c[=!�f !E�%B28H�ȓ2�����Z$�1c�S|u�'q��1mH U���O�>��Td�/dlrXc��Үy�n�B#�8D��Я5-‫T��
;��i��q��
~qR��h�3������R� M'C�������dU�;��Ï�`1Ǎ�U2d�����9�洉	��/߼�R)4;��E12k��_X>�E~�m@�O��-D�%?M�A茍n
X"W82
DZ�"(D���A$�,1`~�xb�ǥ;��IZD`�>��F=16���2}��)���	��b�4%:��$N	5M!�$M�7Wxȥa«*A��"aO@a9��'W�,���.�z��O~�ǅ�X����&$��1��'���qo�L�~-� �0q`h '�:#���Ĭ�R����U�	)����g�
�~(�� �2ʓ}$��u�+����G�*�ӿ-\�����\�r� w'Z�-D���ԧ\�-<�����֬(P��UJ9Ky����CH�y�nŚ�O?�	�e����1*Ad4J�c�!3o(B�	�o�q� ���1�&�1Pϖ�)���V ���m1�����4�$@���?��韠�@�Ȟ�wh�.�ّ�'�̐�@�`���xB�dӶ8%�NQD�Tő(����8O��DŀOX�k�<ͧ4AhI>���1��`��ZP�\�tN�]��7�����	�=o,�#s6�d�8.p�t�g�}��i��h���<
�F�3hN���F�u%ѩ4����d۬(��-"�|	�L͸+�v�-זa� ���lӒ�9'eW/����ҁ��(��)K�G�����]
��U�Ҁڐf�aXT�'�2V��>ޢič�����-5��[D� ��ӵ�Vd�R�~�f�-p,dA��۝5
�E�Y���Oġ����k}�8H�/��c�IjZw�2@`��O�^+�#(5R�zt��7Z�̚b�!>��xE觟��/�iT�xRG�>�4�Z�횟6��1	H���$7ht�`�DY'&w��i���1JG��c^M�? ���oE��~`yf�?� �����J?1��K1U���XV�=,O ���t}�@Z�Hz�Te�6IQ�mfj%i�'k����Z�j�6j�M�.#��p��'�BM��OH
LBs��9��X��큤pj�K�� �O%���\�PE�r�'H��H(AL���<�E��+�Ze�

�~"�I,��i����W���I��ԮA�e��)�3m7�M:��d�Q��-��
'ʰٔO�t�3����h"�����~B�M(�')\��f�>K:H�7T��ӈ.�(%�<�f�9\����c�=��m���<Ɇ��2�6���I�(������7T���'?V,�b�&f8H��L��H@���L�azR	ܚ-�Y��_�$%FYr��۝E��'$BIZ�ۜĘϘ'ʌ����5��XiA��8B�x�'G��6�5-4�i��w��4��`��T���.O�#�ǵ+r���홶Ko`M��UF4iZ7#Q4FF  P 瓭��H�ȓ�.�d��Hn��k����W�����#�j�@�j5G��#[�%6ތ�ȓJѺ�Q���$ֵI��ìA��фȓb�xD��0���/4��ȓh���cA�*>���P�X&>d~��EGr���ʎ�2q;�P�*�0��N6��ؗ�\���H䧐�)!�5��ڦJ�F� � �"�"S	D��ȓ=�(99�A��k�2y�`�4���ȓ�6�����6%�����(݆ȓw�pm ��L�H�S�T�dr����hO��т��D���!*��Z�n���dK�m���@q�<uzf�ȓry����\(�X���;�T��2)ֹ�"�'m͡��gl��ȓm����o�,u
�0����&4l]�ȓh��|��
\��Ѫ�)�,�ȓos�d����n�)A� �u��%�ȓ qFh�@Bа^���
[�^���=�mY.K����b��I�D�S� ���n�&N�!�dR�Jȼ⡊�k�P! R�W$e�'��p�𙟠S�+��a@�=s���$��rm B�	��\��*=9*^�Z��ϡq |��<�~Ń��'"~�A���4�Z\��ƈ�C�p��V|�$���@�
�<�0�� tw��ZdM�k�$���*�|Q����r�!�l�G��'�	�,�A�܋���5�훔�� d1v`ƨo;��C䉴�nT�E�&Dr�3�B��ˠt;P���	�U>�q��OVAɲ�݅Z[j@C ��07B$���	�:�RI٢�SG&:�(��ܬ=<м����cޔ[₊d������'�p5N��-� � ���x6���U�H�r�|*��X���V�.�O�X��Vj�����I�k~ژ��"O� ��bΐ\��d8���u�m�w�'/��5��� MJ|aG�zҢ�O���J|��g��b.(�ȟ$"m<x�C��t��@���8��U��ihT��KA�IW�S� �I�!FJ��'�a�� 藇R�qU��Ƥ�
��d��6�	.d��"o�$N�>��B��K���%��h+����%R�*&���@9�O�p�aJR��5��L~n�5ӡh��:uh���C�1�g?G�I%c&�%dܶ� ���%PW�<��C��1��]�mte��HП��
�n<�Y�f�'��IjA��%����ȻF��(
ߓ`4��;+��"��7m@	Gp����GӠ1���`̓�3!���|�H��4��7�h�#MA�G'�O�!��įx��P���I
t��b��C?J�P�M��!�$��t)zת 6]*�9ÎR
� T0��ףu��O?�IF+��'ĝCX.��U	)z^C�	�w�r�$�wc�JW*YlQ~�	�%s4��'��P�LޚK���:GhZ�n��'�2�DK�a�Zĸ���QBP�C�'�("��M,B����{�"�h�'�H�T͒p��� 5�KA���	��� X���\�cbb��
	�~o4�P%"OT��!g
e'\��� o�4;�"Oν	PC�d�FA�$�A�dr5�5"O�R�H�P60l�(^�sGԔ#�"O�t��Z������H?e3~18�"Ox��I,3��q+��̝7!���"O�K��ˍ���&��:l,�P;�"Ob X�����c��[�KL��S�"O�����2Yk��AU�џj���v"O��$�F�0�
$].n4��1"O���OD�$e����	1Evmg"OD���ʙf��1x�%*����"Oؔ;���U�87R�0��	�"OPE�WΑ�Z�nı׆�����CA"O|�ʵg-P�L@Z��9Ddc�"O�I3q䀛8W��j��p���B�"O�-kB���Y9�1p!B�4�l��V"O��F��;�4AS�D3�q��"O"=H'͘S{a)U#G�0���b�"O�=��c�#}�< �n���>D�v��	H��J~��`�9},�C�	%d�2aD�_Z������]-��C�ɥC/��t��'����r�Dd� B䉹:ila �0Q�MJ�F��{�C䉞"�֜�Y�E�	�L.�C�Iy�l�$ 	`����3�B��:Z��UP�m��5VvI8�eJ�Wr,C�	6x T��Lԩ,m��	�h�C䉓s�H)� ".Haz��`i��@�C�Il&x|�!�ɮpRf�Hr�D&Y�B�ɽ\a���V�B�S��:6jG:&��C�	;:�N�5�ڒ[ ����GI��C�	`B�,1����j
jyH�GE/g+�C�ɗt����!`����� ��C䉮5�D�����nw���B@�5��C��_@.�)�Q�0W4 0�E�@-�C�	�H:Z�C�8z�-@B��?gŠC�	m�	�cV�|OB<C��.&O�C��;=6�����F2F�0�̜F�C䉙r\!!2-�3���7��3L�FC�	�	�APP#˟Q{�Y�E�GY��2FIX�Y�G`S�I�r��!�!�$�/L���0�ܾm���7��3p!��?l� �g�"E�4y���;f�!�:[��Sf�G7H���۬X�!򄗏_�V�{1e�zC���B�2P!�$܍ *�9�@0?tyJ��&R�!�[?IJ�x2�iƔd�H�a3o�!��!88بw��0x���"��=i!�$� P�reA��7��<2��B!�$�X�}��N�D�@[����^�!�A I"��c'~D���ʵ�qO�APb�:�)�i���^ �a�~;BESu�_��!�t�������2�ȭ��mc�XYy�N��v��P��o����'��+VG�S��r��	�.�G�t�)�kA>3�HO�d��(O�O��9��L�q�Z��F�3���"L<q�.�S�"���;gV�S,D{�͕���(�'��Fy����y�r�R��ͮ9����V�F�o�6oN��g�?�H3N�=008�`I['D����I�(t����><���Q�F�-I�L��"��v:c���2�]H�Ş�y*@a��6Ĺ��+��f�|��M�qc��اH�\H��jC���5��C�h-�=*��:�4��-�����/�O�2����&��E��Bw�����D�+$�U`��S�}P�]!dX
�JpnZ>
Ry�O*�gyE,��U����5A��)�ꛓ�y�l5�?D�|��� (I�3e8��C�ɟB�t$�6��$:R�"}�&6��U�F�L�*c�����X�m�\,�3�D۽����I۔E�)���,B�@%�AoޛF�'�4�Bࣞ|�S�^v�sD4_b�D:$�:4b��'Ӣ�s� ��ѥO��O�F�̡;�I[:��y����K�|BǝǪ[�}��ī%z��ɕ- }~�A֠���yBf0g��S
w�6��B�y�/K4�ٰt!�\~�u��G��y2B�+O���'a�v(���yҁ�>޴M�V�Q�[�$�!�K��y��=�2!s���[F�)z�J��y���]���P�!�ebr�cM �y҆WM�������LvrQ��oV�yR�'^�rP���?��`X�'C��y�iB�E���#��^:RP��J�yb.Q�!�&Q�BI�}���GL��y��B�4�/��5B����~B�!:��ZA)���!��l�32qPB�I�l-�H�HƳ�L}�S38B�	J�ʨcğJ�RXBIط��C�/�2�)B��-,�T�10EW�B�C�I& B*�02M��t�2���+уH�B�	���I��������l���zB�&[���&����da��nSNB�d[�+L�h,9;v���)VB�I�W���
#U�D��@B�I�Q���[8t�81�N�b�C䉥L��d��$5a�X�ZԪ�	"�C�I#-OH�b�G�X>j��*x��C��<�>�i��۸�B<��e͚Jj�C�I�\�4�X`*V� ����֫�	��C�ɔFF~��t������xLXC� ��|�G��1K���'���š�d
*b�`1�s��!fb,�(��L:!򤟻I�i2u�M�I�ۑ�!)!�DF8v��`H2F̰LaW(��!���>pHLB�A��"����9{�!�dz��uj�jԸa>�Rb���]�!�d��v��M�+�y�tx�Aؽ�!�]$G�X�3�ޖ|�`YY�e��!��<T�X��TG�����Bb!�d��e6J��E��;D,,)�'�1�!�ԛVZ��2�n�
h5�<�7-�#�!�A ZЫ��
a�}�!lM��!򤂕Y��uF	;�<�c�W1	E!�$ �T3�PBA�щ��d���$=!��<U�l�����%��p	��N�s}!򤉬?&"�P�/�� �բ��	�!�]��p!Zr˔z�xh#Aa��7�!�$�qj"'�Lq��9ÆY��PyB�"-�
��%�Ĵ�2�*�y�!=���9"�D
!���e���y��� ^���r&
�8�b�`"���yba�>]Ǥ���:WWE�aN_��y���
��4�4aغ��ܽ�y���b<��YD!�p�h�J��y�ġQ(�d�#�=n�J�`�OZ�y"��.pNt��* g �DI�%�2�y"jϚ�F�� D��k[�0g���yҌR�8U��@A��]-�	�m��y�bX��PF�	�anP�PWnX�yr��,f��q��*��#��ަ�y��ďc�xp�O��9��4��P7�y�"o)@�!ף@���I��[�> ���S�? |�u��!����Aa��k�p��w"Oz��C�! !�o�Tk�aY7"O@��'�?8���fɓ64PK�"O.�I��]4D�d���ƍ�{�d��E"OdX����yt������j��qh�"Ot|H�n�jYx :�a��O�,�`"O �ڤ�$S/n-b	f
\�#7"O��Pt�@�&g8q`��͑��kP"OL��e-R�X"рוR� ��&"O0lY�׀B*-1��o�� ��"O�-���Ԙ>f��@aa	�[��)��"Oh0��	�Z%�o��^^�qrF"O���H� �
p�%��!����"O���"��WdTj]����*�7�yrm��s�h��p5\EKt�٫�y��\�42	#4\:�>��ј�ybOI�&��=��K (�������y�A�;(����/O�\�Sj܎�y��N�p!�.ǄqڲQ3H���y�.C;h�&���'�Y��U�����y�CԨb������M[U:�X�yR ^�?���H2ʇ�Q~�����Pybm[�8RphA�NI��>�"��QE�<���"#�J�J�n*��jW�|�<�En�$t�!��m
�QbHU�Bb�<E��.�����վ{H�-���[�<�`G�O�:�P bҽv����0���<AD�h��k�!���"��2�@�<��	��@�!�t�ӧSy�<��o�U+:I��B��o^Z	���q�<��b"fx�sdH۶b��(⇤f�<�GhC=_��1`C��G��t�Sj]_�<��F˳fyp�C�	��|�j0� G_�<�p*�+��e���C�5�d����t�<��iE4��i����@���H�Hs�<q'�ÓN���k"�	9L�Ċ��Z�< !�,A�ȑr���D�Ē!!�Y�<�������h]'2(,{�}�<���5c����\�~�� �y�<�G�rɐ�)�I�Qv\��C��{�<1a�V�g]�1B��^��PZ��O�<�7�\���i��N3l��� �I�<�/�I��vA�|Պ	3��V[�<���'�T�#�G�w���R2�^�<�L�}h�Y*֨o�L٪�LF�<�#@Q�$
)�$��:~mX ��AC^�<�"EB�a/���%�׾HN�d���s�<����>,���q
�(n�2'�r�<����D�S��27_6�H��n�<���%��!a��.w4��
�*QD�<��k'�Z55���B�B��$g�<��s	Ɣ��A�?6���w�AG�<I`��-4:�Q���Sl�X���*DA�<9���n���R��%HF��
�C�q�<i�B����wo�u�"��e	Dv�<ɐ�ѳQ��)YR���@K�i���p�<��۳:��g���n��"��OB�<!�/��G<@p��/UU&��L�@�<A�E��j]D��a� � k�ʝR�<� #V�4&��5j?|\H�NGz�<ѣ��H���HS��=6d��Vlw�<�EG�,��E���ٺl
Ћ3. n�<����=c���׷Y	F�fR�<y��S�u<����W�� D�N�<� ���Ml�mk�d�;E4<lyp"O�4�T	B��pI�7%K�0�M�p"Orl�$��d�T*6e�/�cp"O�@�f�T�T7�8Av��gܠf"O�j�.U6b��Yq�Ϡ;�8�#"OI���ėJ�����],5�"O]�2�S#���ȇH�~1�"Oh����.=��4� �Z<s~�-��"O�(1��&�%@��2s�`9#w"O,(�Ɋ*9Q���.=î\��"O 񻃧�5~�:Ȼ�A_�JtZ�"O����H�!^��&P:!?���E"OR,�A���vѠ̸��#p�n�9V"O@ b�J�Z��L��&�2���G"O�a a��vBFQN�$	�"O�D0�	?w5�4���E8�C"O�D�ri�	c\,�g�ߊ�dH:�"O��"���7���z�9q�8�*OļP���o�9�-�eJ���'���Q��� _���K�GX��b�'pJ�6��W� a�NˀA��!�
�'�:@�*Q�'�T�����).��P��'HD�2��ƭK�v���%F�,���'TFX� ��.�>� ����?�y��N,+���``Ӷrj�Ȇm���y��2ᆌ���W����h���yb��"3� p� J.Uf,-����
�yb�+$?X�hg/�M��t�΂�y�N& �.����>L�� P�'�!�y� XF0���F�?vΈr�剅�y��pf�P��2��їM��y�� �����$��`e���yR^�h�4�ퟵ�ba��Ղ�yB�Ü-3���	�."f�࠮��yB�/E\@��ʺ'�Dq��A��y���5��@�w��2&� ac�,�y���*2��4c�g��������y"��!Qè=S�"H�vu��B�6�yb�N�	UY�E���$t�Q����y"� 3XzP��H���pCM��y�oR%���*(� piP��y�a7Aj�,{��Vn��������ybH�5 �jA�R
�N��"�؊�y�	<[Zr��V	JUu�|������y�ŏ�m�$hBF叝P�����y2�Kg(j�OX?|���ЁAN��y��Ƙi�P����w��L	�����y�*4��,3d� u^4郠����y�惗3����"�zIV��dW�y� w�"P���\Zj����ª�y�Ɛj����r��bv~��5����yB��+K�4Dq��I`T��kd�]��y�D�$J:|�B�Tx���SΏ9�yr-Q�V`��*P�����y�����8���(G)���.��yBb1ъ���k���i�-�y"��b�x-�-^4(����y�+I�*��Bҩ̕TFUi3�1�y���HA %X5�:G(��#�
��y�F�7��4�dF���Bqd���y­I$Bt �炵k`���`/���y"��/�8$DG]d�8{�G��yB��{=� �$f�F �JU��y�Э$�|a-'����S%E��y
� ������)�d|��n3'V��H�"OH��q��r��{7�^�=��HQ"O�,q�%� ˀ4�$��t�"O��BiW�w� ;����x�"O����؍o@��Ƣ��H`�q3�"Oz\P��^���5���݂���"O�p�@!X[��K	�%��`)�"O\�se�$g�x�"'>E\�Ċ�"O`����`U���R�Ԝ]>N5��"Oԭ@f��p�t�Y7ޢS2"O�mȤ    ��   �  �  �  �  Z*  �5  [A  �L  �X  �c  >o  �z  e�  Ջ  5�  Λ  �  w�  ��  ��  T�  ��  A�  ��  ��  5�  ��  �  t�  ��  ��  � C � % � �' j. 46 @> CE �K �Q SV  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j���/S&0��$+|Op����� r���1N�gM�|�
OP7	�04��T(|���"�E��U�!�t���ው=g��1�1eG�#�ax�a,ғ/��J�(�i�t@ؒ��v1�D�ȓR��3 鄏e�xA��X8-h��O��=�
֪Ӧ]vq�w��6l���$�Q�<��L6p%�h*��3?*�Y�dJtܓͰ=�5�	+ʁ ��
4����Y����>�C���
����)?h��`�T�<���R�Tjt���uc���S�I�HO����ܝ��X�gD
�-�b��"O�t���/dv�3��'�Bm���]o��`��"������^>��)�-$�:&iT�K"���� E����2.:�yb%�1����.UP����%����'Aq�j��d| %�Rȇ�>y�	1���H�!�d��x���� S"l���(v�!�$.Yb��t  �h��e���T�!�1oE��8���W8DqpGP�q)�'�ў�>���-�h�a��I�n4��*%<O�ul�V��`0Х�&갨hՍ��$=ة��j�x�7͸%��90r
�D����<7�>�Ş�@5�d��1XxR�{�<�&�ȓ`˪����?,~�1��Kd��=�:���؀�bq��2`���$/_!t���Qϲ���"�:휥a���){JUnZW(<��%]17����\�z����n`�<���ł|�x]`���A�Ԩ�qYw�<�W�F+d��p'i8o¼yU�q�<)�m��L�T��������)�a�n�<�J=٦,r�m�Xg�A!�Sd�<)�bD�6�QҎ�����0�W�<	��ƛV�򅁗Q�8��A��+M\�<i1�ق&���� �ޗRk�hsn�Z�<Q*�OYꔀ�M�VK(h`��@`�<I��K�0"m���3@�dt���[�<���\�*9l�4j
�rΈ#BG�W�<��Mά=�������K���JDS�<7i�"CӪu��쉐W�����Q�<i2��y�\��w铣&�ȕ���^C�<i��T�]��h�' L ��eF�~�<�HY:^y�X�ܙ1������Hx�<��l��N��Z�ˁ.E5"fDn�<��� k��`�$�>`��8a�f�<��+]'B�b��_�n��6#�h�<Y+X�@��x�Sd�wo izT'�`�<�fe�R�V���J
N%l�{� v�<�ED��t�V�� O�b2�%�ӆp�<asė�;Y�xW��	a��e�<y�GR�+�^�Pf��L��.�c�<Q�T�Y�T �,^	:5��b��6T�� ��h���)T�L�5c�')��Ab"OB��&(�F�Hx�sK�5
n�s�"O�eQ�D�y�I��G8o�h�""ObI��`WZ��c�$�a�"Oz � 5
)�I!�m
�ll�7"O��3׭�J�H���+!/M�Z"OdDjƫA,@�QV�K�a>"�	�"O�4i�b3�H&À�ULH 2"On����Ogc�1#!,�\�e�"O�tCj�<��  skί7��"O!�i�."�P�h��m$r�0"O8����!7T�+�gA�@���G"Ob��0B�$6]���(�y�R�A�"O(�i"�1�hmQB�?"��"O�����>¾�����6���R"OT�a�iD�!Za
�oC.:����"O���5��@1�aI?F�n\"Oph2�`O�36�b��L�"�F��"O������(��C��	�h::m��"O����$�d��5��J@)�"O`(����(���{���Ć�y���VZ6� ��mU^)Q��I��y�m��7�m�U�]S�%2E�Ԧ�y��Z�����-�as���q����y2��%?:�9w. R�"�1��<�y�)��\�b�_�>��vQ�y�!C5=�r e	OM�i���y§�9�`�����VcFa�T8�yL��Qi1���\4ѷ�R>�y2�ٓPO�%"���O�(� �'3�y҆['p�(X���œ��|��y��I����VJ�#V\@��!�y�[�g��]I5+�*)�L:�cY�y2nS�W�f1i���|�~IX�h%�y��B3�>������yLt�؆�yҠ܇~'lT;�Ͻ �H+&NS��yBB؅v�Ƀ֝zWN-���yRΔL�ՙg��)fZ&]K�%I�yb" 1^5��*4�(mӴ�����yB�E%i�|A��P�:x:3�ԍ�y"�Y.y֩��^p&���A�%�y�)V�n�@���[��Yp�>�y��9$v�!7i�<~aD\�@��yb&B1g�%	���|�x��"hJ/�y��-�d��P���Fx)C���yҢF-V'X�H��	�'�fP�&��y¯�,|"���r%0uʸ�a��9�y��K�t���#Mp�p��#b@�y���
��g��s��x;�Z)�y�)߼|��R���
\J��D;�y"���)�K� p�!d���yr��@���;}g"ݩ��ݘ�y�ϑ�R)@�!��u�&su���y��(Y�:5
�E�3p)�a +��y¥Q<���)�i׊i���'JT��y«�Zp�k��/P��f��y��Zc� 1��@��Üi`�e
�y½J�eГ�
99 �UŉW�&B�I�G��w�P	Hd�M��MOF�0B�ɋG~����eey��ʎBbDC�ɯ.H =S'�ʍs��l�C�<h��B�	�2>�)�cM� �� �/9DfC�	%y̲#�P4�D+�X��bC�k�*HQ �-n.~���0C�)� �`��S�|U�S�ćW�@�b�"O�	�jÚ,dؼ�'o
,>x<�2"O:Iȓ,�0��1��7c]�y�Q"O��K I��&T��g��%H�-1�"O�Hر�>�H��Q!f����'���'uB�'���'���'��'�
�� �&*��4E�-ޜ���'���'HR�'�b�'�R�'Z��'��d��S68N� �m ,N�\���'`2�'���'uR�'xB�'��'nJx�ɖy"�@��2;-@��r�'���'���'p2�'c��''��'��J�d�4zN}!�o�6�qcC�'72�'�"�'�r�' ��'���'9}�Î�;&�� $ ���ZUz2�'���'�'h�'B�'�R�'$�$sp/K9Z�B�0G�el$�p�'��'K��'���'���'F��'�`�	Ã2u;�M;C�c��P��'k��'@b�'|2�'	R�'�B�'+*-(A_8��@'�D"wЙ��'���'%��'�"�'���'��'����AӬd��#�*�R��Y�R�'��'�R�'"2�'���'���'��p �+Z��p���2�p��'8�'���'6��'���'���'6F�;狄�e�n���̰%)�XkD�'���'���'�B�'���'#��'�Ƶ���͂~��y�S�ގpU
*��'r�'.�'�"�'D��~�*�$�O���B#Fˈ����_�,L����ay��'u�)�3?Q�i�⽨��LT�v\�f��B��1�����Ȧ��?��<��Jh������ʐ�壝�6����?��Q��M�O�S"�bO?у�C�f�P�`U���|H)i�e*����,�'^�>u)�N��-<�i���\�"����G��MsQ�|���Oؾ6=�-���A;���K$�Z1��jr��O���l�lէ�Om@Ȓ@�i���_c	:��/�gL|S#!W�Z$�$r�4���5p�=�'�?��$ǂAhx1���C$�Y��M\�<,O�O�am���b��zTK��eS����l�6j3�P�a�j��������<Q�O���Gi��er���H�\A�1b[~��'۠��a��ߘOۢ��ɴ__"K*y�bE0f� ����D���_��XyR�����ȥ88�ȆNH/7�� �h��w��Ĉ�����#?aŹiG�O�#U�A*�B�*
�I�@$2m��O$�d�O�%�V�d����$��nTa�ĕ#R��)Pt�²/]��H�����4� �D�O��D�Op���D���q��0y�x��ē���d����b��Gş��I���$?�	!h�+k("��ӵI��=6�J�f�>1�i7f�)��g�`���O#:��H��Ӧ+��5�7N��m��)�ɂtW<u�"�^x�1��|��'���`�j���Fɵ(��ɂ� 0H�2��?i��?Q��|�+OtAn�4�J�Ɇ�%fE 2�Iqe��;���:O��lZv�-�I�|�Ʉ�M`�O�fѲ�X��,$����Ğ9	ݴ���Ë'�.���'ƸO�m
^�>�ðo��p!��+�yB�'���'�b�'�r��F{�D�r/[�%�{Q"��I�l���O���G��u��{>�I�M�I>YE|V���Ż:�%��M�Tx%��+�4K��O �i��i���	.?�T��!��"�N��x��rC�<B)Ro�	Cy�OJ��'(r��6ň��p�2�-�Uf�4 %�'"�I��M� ��?)���?q+���L7wr%(�fҜm��A���D�O�Hm��MC��xʟ��8*J��m�4��'��-� 		���$��I0�i>) �'�`�&��sH�d��A�).S�4�hf����	՟��Işb>q�'�<6͎"�R���/Y�U���G�ݲJcL}ҥO�<�նi��O���'&<7��� } �B?���!�E�WR`=m��M[PiX-�M[�O:u��&���rI?qI�mP�
(09̌j�����l�$�'2��'|��'l�'_��3 >.�9d��/l�vQ����% ���4nA������?����'�?����ygI�t��9gG�SR�MSr�Ċ��7�Jڦ�AI<�|�S-��Mc�'@dz��!0^��T�ǭB|#�'��4҂����z1�|�R��S˟cf �$L]�I��b͗����B�����I����yy�uӂቶ&�O����O.d�4���<�����5��U:�."�	 ���Ӧ		�4D�'�Xt��!�C�Y�ѝ�ܜ��O
-j ś�3ܺ�i7�iX�?97L�O�0j�f�%�GǺs��`j�!�O��D�ON���OĢ}��P���&�2bx��7ĉ�<���Z�\X��,�����'Hx76�iޙ���#c�� �@-ߍ@ɲY*�t�89�4D��cp��t��h�l���d{d�쟶����9O�j�����7.P<{�������4�r���O����O����/U����r��%��xdL�����hN���c���'Cr���'b.|��!NH�� .Z[z�	���>A��i`�7M�O�)���Wʡ,Єh:��ʻH����Ԯ�8��5R�O��3�	���?9�(:���<��F_2(<���$�J\��%	�?����?a���?ͧ��D���t�ߟ�@&OO�X�,���̐SG.����̟X��4��'�b�a��*g�p(oڟ[�86��ʳrM�,��9�A��^��6��4:V�Z���i��� `��Ä Ă�;w��y_�01O����O����O ��O��?i���^K1)��~.شX�$_�� ��џ�a޴ �`�ϧ�?!�iw�'d�����^�j�hSn_=]l8c�9�X��1���|2�&V7�M��O�(���
.�1x��ڈ+�*(� 
9.�����ꨓO���|����?��yHn�4�4x���K��ѰZ"����?�-O¨m�5_�������J�$�V�i��`PC�>j��s��F ���[t}��'R�O��2D݀E�]�ys$4�r&S#y�@� �C��wq�i�g'Xay�O����ɜ`��'��䱡@S �B�;���(2 ��'K��'{2���O;�	=�M���3B�2e��(�EĘq��9g:�?��7ϛ���qyb�i���U��D�K�L��NO�uA�.~ӚUo��ZE�tm�S~⬚�D�	�o���c[�� �bڟ-�B���k�8aT��<��?����?����?�(�`����?AN�[v����	������zg �ȟp�	ן�$?y�ɯ�M�;2�B큵��-o��U���ԸKϊ� �����O0�*g�i��$3uhD2��P�Bz�BaG�%7�F$H(���vƓO��?���:��i)��U`y�	(��PD?�Ȉ���?!���?A.O�`o�
���	���I"s �7�O�a��9���H��x�?ɃP���I��M<���s� d�PL��En�H �e~R��q�d�1C���O �p�I�#bM�$%~���j�dl��A��L����'�b�'��S��,���̴=��;R��>��M#����dZڴ09�p���?�i��O��Qsx5��O69�΄�u/,l���O�7��5C���䦁�'l@��F���?��-Ȟk�u$���;��	���*��'��i>]�	֟�������ɋsn��)���7�$��tLEr`��'�6�8E+,���O���)�9O�Q���/�0��� �;��x#�R}��'2�;���-�F�
��fl�,b)@�,�ʄ�Ӡ){��((�Tj��'\�$'��'.�!Q���6� ��@C��e|�3�'*b�')����DS���ߴ"s��i��e3r���i:FʑJ���:8�L!�z������g}��'�2Lf�4����.�^��rI���(R�l�>;9�7!?�
32�I*��ߍkǜazLг2%��e-�� �%e�����������IƟ����I}�XA���`�8��7�߰�?����?9��ik^@�[�H�ڴ��Q3��a�e	;L�,�aL��^�j�R�|r�'ӛ�O粌F�ih�I��Ш�ԡ+���w�@�0�ޞN�YP�_y�O��'-�e�2#p|�%��~~���㌅]E��'� �M+�K֑�?����?a.��O̧��4 5��R]��@���2�O��D#�)�@k�5@�b�*Q�ZC� Id��	�
XS��'բ�r.O�P�?���0�D0���JĨh����V�Ab�$�O��$�O*��i�<q�il41�v�ϟ ���D�6M���sA�m���1�M;���>!�	jj����Y���!�qy\y�/O�Y���v���,N����/��X-OPI�gL/�lkej�M2�d�U7O���?����?����?q���,��бw�X�I���Pr�S�]�\lچA�l��џX�	G�Sџ����{��ʶG>]�A�7G��u`�'���?����Gܷ7M�6O��k���ubjR�ڛyr ��:O��f�!�?�'G(�d�<���?gS�<�~)ZtK��
 ������П�	�P�'�7��^���OJ���y}�H@%u�p�Y�IG�e�D�H��O��l��M�u�x�MY�V�q��@�p��1�������M��UK�#܁2-1��Ys��7-:�$�.)0eq���;`J(S����Y��d�O���Or�D5ڧ�?���"��3K�LEN1�k��?0�ik���Y�`+ܴ���y���%,�-�s�M%|EaU,X��y��zӎ�m�MS5��/�M[�O2�RƊ�0�℥��h���d m*�p
Eϑ%L�ؒO���|��?y���?)��0)����:f�jp ��/V�k)O 9n�tLz���˟���r�˟�À�Ƥ���'� ���*b���D�O@�b>�Cg���A�:d�E;I��:��á��t��~y"��& ���.��'�剂g�8�}���h�àQ>���I�������L�i>��'O�6�#����"\�:1�6��L�G`�;G�������?��P����vyr΃� �>hٴ�O�
����������"�iH�I
jjF���O_6M%?���~86YR�c�b �bE!݁/2����p���P�Iߟ�IN�'$��1e'�=H�ԍŸ9�Ҭ[*O���[��MyFB}>�����M�N>�"S�S�����׺V�3�6) �'���'m��R]1��3OL�$K�aݾ�g��>d���FdE-gɶ�9��-�?�C�8�d�<�'�?)��?�4�=�:�aq�^�8�J�e ��?����ۦ��"��֟���퟼�O��x�L76ۊYs� ��Gʪ�@�Of8�'��6�Rߦ�K<�O.^��r��&,r��!⓻;�B5�╭+ 
�0Ю���4�8h�]�F�Op(�hFf?����:'_n%����O&��O����O1���:��F�G�B^�"���\�j��q�]�$���AaT�T�ٴ��'�j��?G(��v�,5cH�~�h�����@��j7m"?aD T1��)���� 򑡕��<IL��Ԉ��=�����6O�ʓ�?a��?���?I����IV
������{HJ�b��c���m�a�����ɟ���n�s�����s�M`1�v���dq�`'Gܛ`Ӿ�$�b>m� �ݦ=�N*���t�QPu�4SC/՛wK��I�U�u��OL�qO>�-O�)�O�cP�)N���#J�C� �8���Of�$�O^�$�<�#�i�r$��'��'�d�!I\?��??��;��B!��'��i��6�o��&���Ӊs�r+�P-l��IQ�-+?1V��o�� b�b�'l��$�"�?��/^%k�V-�С̠pyR�愝�?Y��?�������0�-Ôj�����Z\��KMßtHٴuL\����?y׶i�O��\8/`T���˅_��e��e��C���y��4[�fovA��i��ɾ-�h+@�OT<lI3ծ8�(:��4q��h���V�	uy�O���'���'jJ�Q�<���@��J9�d ��V�剔�M�3��?���?�H~��tݠ���f�;<�\�"�P&h}�}`]��"شL��/��i BT�)�BL�B�d]9��B5d�>����̟'��	�jSdR�'E��%��'3���ui�]�Z(�H�NV�3�'�R�'����Z��ݴ<\��n��c�#ѐ�s-#M̡Q�@4���O}"�'��	�ҎD@��5�xhJ�ƌJ\�(�u�צ�ϓ�?CIMM)������D�*�.�[�|�m1Y�t�3H�1):��O��d�O����O���4��]�"����;!��XB@�M�2�|��I؟���4�M�#���|�I���|�'�!���̚!���&��'e^�-�$�md~�',��dh�)�`�Ѵ�ئV�P�)�៌rq�|�Y����ҟD�I럌�eIT�������9u0։��� ��oy�l~ӎ0q7��Ot���O˧#�:`'",�ՁF*	�,���'�.��?9�ʟ��Yc�ɬ�@��'
�g9.4��
J�.&�U#�靻}q���|�v-�O��	M>vF�3�$���I@7��y`��F��?a���?����?�'�?�����զ���Q�*��( ��гl�Dq��'��U�I���柬�'B\����2�Ԑ���J׬��pi\�u}`<������E� ����?�!)׫��Ya�AҸ�򄑙O��̠V���'"��T�
5�<)���?���?����?�)��ȃ�t[�ق��S6?�����n�ǦQ�ga���h�	՟($?m��-�Mϻ@u�e�5#R�8ݦ���� %�b�
w�i�b6-�w�i>��S�?9r��Ʀ�͓^��,���Q�L�ܝ�"N2C��,~(� �,�O�${I>,O�I�OD!!��<s�U*`Y�Ǿu��O���O����<)t�i(��G^���Ii-av��"+z����b� *�Zp�?Q�U�8�	զ��O<!�㟂(����ҽX��%`4Ir~R���{A�<��m���O]� ���e��A���bO��E��X1�òO��'���'����Ɵ���%_�f\�ۢ�ӵ�V��¢��,�ߴ0��x���?�2�i��O�nv�`���#��I�y����x���O�u�ġݴ���S�С��t��:���Q>]�DHS�]����(�$�<)���?!���?���?����f�(��d,�� f̣a���'+�7MQ�b���O��d,�ӎX�Yp�FB�Y0h9&��a��LӭOB�D�O�	'�b>�pх�&)v�쩇��s�%K�oQ�o��8���0?Q���"3�����!�䓲���Lx0te�4/@4�f�*j�$�Op���O��4�Hʓ5��G��d�6n��Qy��V����[<!�%��D�y}�Ik�d�l��M�Cg_�9+�]����TA�-s	�L���3�4��d�%1�����'��OpGC��K�0�0th̯e�U��U��y��'���'��'���IR9I2�ɡ��.'���:YF"���O�d�����dy҆dӈ�O�B��>�����(�P��ԩ�a�	�� �i>iBD�Ǧ��'~�q"̈́�"
�1�&�I�)r�eH�X�H�ɐh��'��i>���럌�Ʉ|Lx���0j��`��h��͟8�'H6M�5:?d�D�O����|��A�7���@�w���2i�E~�O�>���������l|�����Z\T���ѭ'(mpǧ�
;�"���H�<ͧ})���֣��tϰū��	�HȧeZ�B��	b��?9���?1�S�'������/�-"?�y
��Z����\��	џ<0ٴ��'�Z�;���
]�>�*,���A.q~v�ڐ�̊3��7-�Ŧ��e��ɦ!�'�.@�F���?����PC�m��Y� ��Q��`ܖ��b6Oʓ�?Y��?1��?�����t=ڄ���X1�d���H�9���lZ+Hr ��͟<�	G�͟������F��������m��0�y���B��?����D�O�f>O�����\+�`)(b���|/
��5Oȵ�`�?���)�D�<i���?@�ΑfF���4/�w89c���?����?������ݦe��Í̟���ӟ4��#�7w1��{G�M�L�����Q����ן��I��ēNx�p`N��*�0Ma�a��|�%�'VH!�r�_��!Ҋ��̟4҂�'��,�W4F����d̔.bY��r�'��'�2�'��>��I *��Z��P�f�j,rW�Ä[�2(�I��MK���$�צ��?�;89ƹj�d �4q�� �\��ϓ�?q�����=U+�֗�PX ƍ/w�d�5� �\cd�foH�ó���b�<�B7�/��<ͧ�?���?����?��-�`'���L�D�hYB2!�6��Dۦ���ҟ�����$?��əBz���ɝ!N��Erf+N..�D=r�OL�$�Oby%�b>��`l��?
�}9��>k���bJ�&&���'?���pO�D����dLq�� � �an\�f߻I�����O~�$�O��4��ʓ*���úDg" �/O��]z��3'�p�h��<kb~Ӳ�xگOl��<� ��(����`�Y2�� �
�;2`�i�4���P+g�2�I��9y��� �.�(��K�Ď�@���T�!����O|���O��D�O<��&�S(d�x������(h��S�I�Vz��I��(��+�M�bd���ą֦�&��Hg��8��X JׂZДɲ�A�ē�?���|J���MK�Ol��ߴ����((]t�+hV)�$�{�'f�&������'C��'�l��lё,�p�`u+��O+V�˦�'�2X����4�١��?����iN��L�f+� `�֌O��Ɏ����O��$MD�i>���4��� L�D�yۖ�H�u^�1@�ds|�J��#?���5�������-^��K�C,�EoC���9���?���?��S�'��KǦ}Y ���q�V�9po)i
 ��e�ܥ:���'@�7�-�	*����OR���� w�F�AR�D�~�k%+�O~	l�)t�x�n�r~�K �h��<��|���{1.�2JK.ӬīdE���<����?1���?���?I+��t�$B�M_�m"�I� +���DjE˦�js�K��`��ܟ�%?�ɥ�Mϻ5ܘ�1 ���"��W
S,��9Z���?Y@�x����6`���5O&l!�D�6���(_(G͔Y�8OF��cC�*�?	�l9�Ľ<�'�?�G�	�̢ hUqk�M��ㆰ�?a���?��������2R%���������3eZ�E
�c�M�&\��D��o�C��I��M��io�O��Po�@Z+����R`�5���*�C�.�4-�r8�/��⟬�pM�	���V�K�,��{pf�ʟ��ϟ0����D���'����bÒ9��R��ܣ<�xPF�'kV6-�j�˓}���4�z}z󅊬
��3�/9s|� )F<O(���OҘo1`yoc~�Ɯ->m� ���/-Htq��#Z�Fd:G��I��QŒ|bS��ןX��ݟ`�I۟��#&��{F�ȡ��2[���e��Zy&a�hkħ�O����OT���p��RNh�D2�͓X��'��'�O�I�O��)��Rv���#�K���c[�#ݐ@��9;��	�b�y1v�'s�&�p�'�@�C��/T���c�V�zP�'+r�'�����W���4@�9H��f!���T*���Ӧ��g<p̓o䛦���{}�'"�}ӂ8H@�Db�`�쁊-�0{fFʦHŀ6-g�p�	f��Ta��O�����P`�`F*�/�Tl6�ٖ--�y͓�?���?���?���Oq��B`�16nD�W��)�H�x"�'��'Q�6��-N��o<���|¦X	}�`Ȳ�Z�A�^Y���D/ld�O6��O��]�6*?yS���+W�2�AV̖0B��r�>R%�O$iM>*O�I�OB�$�OR,ZebƼn��i�2%ƬQ*Ha9Ҍ�O��ķ<A��i\�;��'���'�哌��	��*M?9r��#@73UH�
y�Iן���"���|B�9���[���]�a0U���8�v@B�@�!��e�f!�r~��OUL��	�e��'x�p#Pʎ������4}b���'���'[b�O�	�M����U�~��2���b�x�D�B�blB-Oإm�w�b�Iٟ0��-P&[_ʀ��T�y��F��D�ݴ
ˮ�
�4��D�e�I������kM�ճ�IU	j5[`��'Tl�}y��'yr�'���'�RV>ysaI���xrr�է3�\��F�$�MSGEH��?���?�N~����w��@�gLG�R�Ԕ��h!V�a���'�o-��I��
��6�h�8ص`C�Yh>�+^3U�u�bq���%�����G��dy�ON�D��Q��`��g׀ �F�B�)NR�'-�'t�I&�M�B�	��?���?�3
�,v��l�94ZL��m ��'4�˓�?I�45�'���2t']�>��"��ɯzh���O1�F�'o�T�'�)��?�'�OP�m�`K
�;���fϜ�2 ��O��D�O��$�O6�}r����tLH8X���c-�V�4Xy��o���G)v��	��Mˎ�w6��5o͝z�Hr7IY"=c�M{�'3��'��7m4wH�6M,?��,��;ˬ��H�$4h"��</,�`��L�|#�AJ>q+O��O����O��$�OfU��������ㄒ
��%D�<9Դi�L�ɤ�'�b�'��O�B[ˆ\�%/�5�04P��@*P,���?������O�R�(�Xh�l�qh�pf@�T�O�a�O�� ��(�?�0�>���<a���/�j`�2��`���
��?���?9���?�'��d����V��㟴A��	+VJ�rF�5s��d�a�۟@��4��'x��{盖�f��$o�=�� *�A͎d֝��ѡYN�,�%�B����'�fQx3��?M�}���E�e�gC�Rb��s����?a��?9���?�����OhEy�B�(Y��O83��a ��'+r�'Þ6�F�:e�I�O�np�I��%�@̓�-�Z�qhsʸ��I>y���M�'T	�4��DD�+�� ���!Z"Ҡ2cfn�@�B�?�%-�D�<ͧ�?A���?�ŇR��4,�&�E}��)��'�?����$QQ��ǟ|�I���O�x=r�.�$ݬ�`�J�:�@C�Ojt�'�B��?1I�)��l��䲧ㆂe�����T��2��5��{?�	���dN��� ��|�L�8�IRE��oAf�Sb!��'��'��$U����4jD�Iȥ��j�L<��ƀ�� u! Kք�?���ig���d[}B�'���ZF^N�|�����ȰIC3V�4F�UĦ��'`�=�t���?i�X���c�-���U�fI��Sb`�ܖ'���'lr�'B�'*�-�Ah��ؠ#p8�D������4rH��?����䧰?�T��yg�K�rvW��(apA�O��X�����I<�|�C���M�'��=�@iL�g�i�WL���
�'��Ly�P���0�|�_���,��;�n�v�,��%�������	��	xy2Kg�X��D��O��$�OB̋�Cۿ�������i�B�cf�$�I��D�O�� yg��JI�rAJ5*v�,҇�5?��%�G9ɠ����@;����?�����>���0k��N ��`��M��?!���?1�����ݟ���V�%ҨA	F4{��Q��ɟ���4	��Ũ��?!��i��O󎖡�ڽ�e[!$.6u𧗲O���O��Y&�iٴ��DS�n!��'�@�,.�tqI�9��ш���Li�'��	ڟ����(�I�\�I�K�����ܳy�"�yS�_�bՖ'��7�\�v���O��D9���OH\�@�ήɨ�h���5��UP��W}BOg�,�n?��Şi�"5)�� +9jiʗ!¡i�.m3R��H���'�h5�v��3�|"U��ڤD��v(�{�lY��8���B�'���'��O�	�MkP.��?����Z~\��e�4���G��<��i��Obh�'��W��x�N�>@j�`a��zɮ|K񈍡Yy@9n�T~�-E.6-���ӛ@{�O%�揻�,���O�~��ث�M��y�'�R�'���'�"��s\Fh!D���!ش���N����O��Ҧ���YyR�g�,�O�0�LQ\��(Ӓk���a�#��c��⟬�i>�����Ħ��'v�zVϸ!��ʮSî�U�TR%T��I#yq�'!�i>U�	����	���1pe�<M������/�6��I˟��'P�6-�>�\���OV�Ģ|z&`�	\����a���0��aҴLW~B��>ѐ�iO 6Vo�)
�����`����"a��Ć8r�zQX�;:��d��G�埐�&�|BE]w��`�(�-6��c���pz��'���'����Z�`��4C�X㜫Pr%(bB�F�`S�#�5��$�ʦ��?IR��l����A��*������O�K\��rش �f@�YU����� ��+��T�~c�D�O3\ "��t����<�,Od�$�O����O����O�ʧsAdX � w?��c�d���,Y�i|�� ��'�"�'��O��}��.	�^�L�٣�P	g�RA�o�'B�Ym���M{t�x��t��{v��3O&���)v��yBG@г:����=O(!�C�_��?�).�Ŀ<ͧ�?����&���I�l�9���`G�3�?����?y�����u+�ӟ(�I�@kbBO����)5��%%��Z�[u�-��I�x���ēs���*��.^TLBF
Y�OB8T�'���)�/�d0���h��p0f�' ����[+@����4�V�z�L����'O��'�"�'q�>��I$la�A��OR3a4 ���H�3h�h���M�*K���$���q�?�;�����͉`s�8S�Y�@��?	�1����-+_�V����w�٩G	�d��qJ^�ʒm��@0i���4V��&�x���$�'�'wr�'Mjy�'�]�9v|}yW�Q=KK�d��V��pܴJHXB���?�����O4r=�" ��t��mb�h�.-�9��M�>��i+�7]v�)�S �rSF�	�ڭJ��� *�`��O�1o��Rb����O��9I>�(O�-�Q� ��8�J\�U=l���E�O����O����O�ɬ<�i�N���'ǎ���/
�	0U@�=�p��'R.6�!��.���ڦ��ݴgś�DE�{���k��Q�"��0Zp�@�J`�i���5h��QI��O(q���N���^U�D��8���a֥ާ{����Ox���O��$�O<��%�Sn����-)��a���.����	������M�II����K֦Q%�(�Ý7a| �wK��!C*�pT�����B��qӲ�i�0U�6-f�,�ɣy�ܝ;�a܂i�ڑY�IV9R����(�>r�]Y�y�O�b�'������ `��O��R�n�u[B�'��ɨ�M{�C��?����?9/���r��Z�����3 @,�����x�O@��1�)2�O�[t$��?Wh�Îʇ#����17�6��)O�	���?���/��:lؙ7 �	�0h�Pl^�P����O����O���I�<	��i5n<a!���{�XPQ�P>V>�X� ^,��ɂ�Ms�2�>I!�i�F-+c�n�y�a=V�d�@-tӼm�)s�n�_~���(n�e���i�=E�@�V8u�dͰDj]���D�<���?a���?Y��?�.���Y�iU"7ά�"͟%��p���Ѧ�a�Yy��'��ԉlz��p��7.1
`���8�s�ʾ�M��i�O�����霘��7�p�� �@�����@���	ѹ�� �3O Q�ժ�9�?9P�)�$�<�'�?�`��m�d
��M#��IբR
�?y���?�����dTɦ�J�Q̟��Iԟ$�eaF�mWz8K��	9?�@`�jOp�|G�I��Ms��i|�O���b�ƶ�2�â�݅1������p�7L�hY"��O.擗i^�Oҟ�ӦG�X=��.:����¡< ����O���ON��4ڧ�?i-�:$�	�B54��܉�D�"�?�A�iZ8����'pRJ{�p��]1}����ό�pM�p�ej��-
D�I�Ms1�iTl7��"iՌ6�7?�b�ǚ%X��Z`�F<K'ɇ�2�<-Qj?=��N>A)O���Op���ON���O�zwE8�D��F�^K�,���<q�iĂ��V�'�2�'���y�	�y�(�3�/�>cMZ�hϬh6�꓿?i��Dy���O�y8���M�Ya��Oc�f����g�HI�O�������?���#��<I���PcXP�$I.Z�̸Zg����?���?���?�'���򦭉�n]��t���M�()�@�3^���rw�o���4��')6��?�)OP����M;Y80�ǩA�:�	���"!��7:?����*��� ��'��{��<a����w�$|}��´a��<��?!���?���?I���-E>�l �hA6�m ��9���'���~ӺDR4��<1��izɧ�6���Z��i5�K+mM�)�ġ���?!��|JG���Ms�OEB�:tt��PkN\�ȡĬY�G2�?�PK.�d�<�'�?Q���?�fF�kјkd��#��0��M��?Q����d^��-h�gKzy��'��qI١(ԗm�:�B�E�%\���[��Il����S�t-��]A��w��?{�����d�y�5��)\��a�O� �?��J/����qR4أ�"L�tv�i ��" ���O��$�O���)�<�#�iO\4���<J:�)Fa�4jmpM(;��=�M���a�>���p�pih3�F�\d�تpT=,0����2Q��'�,@��f����B&U+3`�T�~���L��daE��>u�;�ƈ�<�,O��D�O����O����O��'l(�z�m\�V���[����l-���i�d9b��'-��'��O,��t���F�������D�v���g��u���d�OX�%�b>���̈́উ�7wuz�ɞ�C������2��D��LI��)�O� #K>�,O��O����(̅Ex<3���$~��b+�O��$�O���<�p�i�`�Ҵ�'Y��'�Y`F�R�?���z�NY�I(ؙF��y}B�'x�OD|�eCА!��|��ɿ$W�Ie����$\�*����r��Z�S�+�"��ȟH��mV�$S��뗥��f�xa`��������	ş G��'Y�����J{�&ڰ{�}8&�'oL6�3T�ʓX �V�4�4�а�3<��JvA�z �`0�0O�$�O �mZ�M� DlJ~2`L)r4�Ӈ}�����)� t!�ə��_,RL�8yЙ|�[�������I��|����H𤂏%ܠ�!C��y�ԕ���pyB�a��`z���O����Oړ�����"?62]+��C�Md�j�MN }���'�"�'zO1��I���ߒ�(���qp�̍x��������)�&��R�\y�[�C�V��3AF
�l��d�:!��'R��'G�O�� �M/����ɮG|�������	\�i=`���M�����<���M�ոi�Mɖn��?x�7��1
��ca��cd�&<O>�$IX,2ȳ�����?9��OYNu�r�Jsm�E�W+P�?b�	ǟ��	П�Iӟt�	O�����G"��eva#+T(� ]����?9�Q�����|���}���|��ۈN�~a���G�;��1��qp�Or�d�O�I=D�6�4?��-O�?G��
7ν Z Q�+
�-�yCS��O��H>Y+O�i�O��D�O���o�	�.hr�b�-5����B�OD��<qp�iB�l��'F��'F��w�Ф��	�X�B��vb��T��	��\�I8��S�$,��6Qj����T��37X�
�2@`a��x� ��O�I��|��!��X��ɂW�՝@*���͕�5�������sr�]:�*�G�4i��ʤ  @�gf٢=�z�tϞ��D�kB��G~�{P,
�{���9H?����a*˞���2�O]��X��l�����a [�̢B2c�<8z��/j�R��w�/Q�Ψ��߈uEܹP�k�"7����i��7��=8�F�/��X����.E���p�ԞYlAm�8�B\3n�9*�UaW`��=�>�چ��&��4���㖿+�f�z��!"����W�Z_�926]����aI � ����ǒ%N�V��%S9$�$E�\���Ke��?�K>�,O��x��e��PQi9ve��Kv	F:1O����O<��<�ɐ1PW���4�.2�2���F	>�	П��I�IP~B�S}�Ҷ�Hyz�oÄo�ʄ�@���d�O@�d�O��#ji�ǝ��� �F6�� �bG|�Y�h�6��7��OV�O�˓jP}�>�����%c&��W��������i�I����'C�e�P�<��O6����\�R)Y#}8*�D��W�0%&�P�'bR  ��T?MS�BT�X���W �J��CW.|�Xʓz�xT���i���'�?i�'��	�S,,-:��"s�x��f^P��7��<��h���OMZySf	�,�:��
q5� Bߴv��{��i���'�2�O�b�S�e^�gX�X���%E�.����M{V��F���\��ƳG(J%�O&�}��%\��qo�ş�����āvoZ����?����?��� ��a�����1L��W�dx%�Q56�1OD���Oj��	�����&�#	r5�Ѹ{VB�lZҟ���A�ē�?)��������J��)��L�d�D�E��K}��Ø'���'V��aR	��8r����h��̐�%����BH<����?�L>�)O�m�"��4�(c��~���CE
M�1O����O����<��IX){�	*��Lh-�?�����mX�H�'��|�R�x��E�>�W��0_bX�a�;b�P1S̄P}2�'��''�I6[�",iO|�ć�/Tj(URn§������L	A���'J�'��x���l���8�c�;`�H�p5����M;��?y/O*4�A�v�Sϟ���lʨ���
H� ��ap*G�A���sM<��)�tC,Y0Li ,��<�l�,�I. H���ן8�'��$�'_Zc&�#��Ƀ8��A�
:7Zڌ��4�?q(O.D*%�)��7k`Zј�Kc��j0%P1M���LW���'��'��4Q�0�O���p�
��M ��:]�کA$(�>Y���^���O� ʘۼ�h�Q5#À1˗�Z�P��6�O(�$�O�0���O2��|���~�<M������XU6��"h��#<����t�'��'�4�T&��$R� @7�Q��t�{��>��	H����<�����2q2tBR
 �\32��6gx{s�x�����O���O��p4zY��F6QRx9E{F�:A`��AM��xyb�'��'�r�'��쳗'�3�~��dV'@az`"��tpb���y�'���'w�I2V�ɨ�Oh��A� L�PMR5�⑭#���4���O*�OP���O����������JX�afҬMܦy+F�>����?I���D\K"A�Od���#����!�^c��í!��7��O"�O����M���m�_��� ���ln�QA�/�(H�@Do��$�	~y��C$z�'�?A��b�c��z�̍��*�x+4��[�VD`N<���?)� ���'�I�;6 ��;�Dͬf�X����ڍ	���V�T���Ջ�M���?1���:�X��X�+���"���u��{$F��{�T6��O<��Q����`�}�A%ϫI�"��l�+�t5!� ��QNݳ�Ms��?A���:@[��'H^��KF,n�+�Ůz}�x�e�{�n���d%��l�'�?y%˼:T���-9!��0�eI�Yśv�'2�'n���Ǹ>(O����l�R�_�Lv����S�$����6�IN	"�'���Iʟ��	2l�8 ��X�ty#��6Lx�ݩܴ�?���.��\y�'5ɧ5#��'C��ض�G�S����P>��d�7M^�O����O$��<Q���Xk�r��!{?8�`�ώ>e��ȃV�̗'���|��'���G'9��Ab��F����i�1��0r�|��'%"�'%��Ĵ��OQ�˛'Y�0�����8"��x�ܴ���O��O>�$�Oz������R�NK�U�w�[<5���@�>9���?q����䗕1�~q�O!B�N�0X����D:���Ȧ�V��6��Oʓ�?���?��d
�?)��Tq}B��O�F@�� w��^��M���?�,O���Ig�t�'�R�OZ>����:K�FUA'j���|E1�$�d�O��DT�G78⟼���
�᧪�ZW͛��F�O �oayR/^
>�d7�����'��4&6?!$�!!���f�݁]�^hzA���і'�db�'���ؓ��V�B���bR�r���$��.�MCcH[�GP���'$��'X�tf*�4�0�����@����/1�e�`ɦ}��,П���~yҞ��'�r�A�E^`h�e�?�j%Zqb��6��O����O.�"b@�i>]�	x?�|zn@st��fe���������My�ML�b���<)��?y��\L�����>L�6�S"��&��!C�i��jU�y�BO�	�OB�O�NN�u��0qΆ�}��,���$f��	�_�0]��U�	����'�2bJ7b�!�F�����p�5���1V�h�Iҟ\�?A��?��ߐQI �P�(SiD��䥊%g�F��b�Mw~��'���'���;..�ȟOZ�u �aeN�QE�w)�t}b�' �|rW�83Ġ�ܟ� 
�k�X\i!��b�l1/�����O��D�O�˓/0� e��D�Ti�җ.* q����:Ȫ6�O��d�<I���?qҢQ�?�L?�1$�U�IF�;]O�M��CkӤ�$�<q�{��,�����O����| ��>&0������xr�'�ίJ��eX�y��(�R��j���E�
(  ���i��2SB�4����������'w8��Ң�2�7 ���6�<����?����Ԑ�ܴt����@��e�b����5X��m�^9jD�IߟP��ӟP�tyʟ���G���p�V�a�J$I�A������K�	5Ks>b�"~����/i� �� !pv�%0'�P�7��O��D�O���&�<�O/�M	�L��8J�JqGS,U����'��ڄ:�$>I�I��	 $Ɛ�㭌^���SG���Yڴ�?Q�+�W~�����'�ɧugfŭ`�&����I���DH��� x��$!���OH��?�ӉH6f�(�q�ףjx��W-K�C��`k.O����O�㟸���08� \�+TOD�A�Qpiݎx�T�r�(_'=
�y�'�B�'/"X������4��[�46_ v�L��Bջ����O��:���<Y����?s�P&r�&�!��A�]��F9�����p�	�̕'tRPA5E:��6WO2�:�c�|D���Y)y;�DlZ֟ &�D�'- Y�'��CL�xY͜�\�\ ����lN>l�ޟ��'�r%�&J�͟<���?�FL� �&@5ʑ/�;7O*��OJh�4l�;1O��5N�Rl �"E�`�6%L ?�7�<I�0Eb�6�'���'9�$'�>��0�����T,hF�2�,\
B�8nZ�����0#�V�I՟̗'�q�4	 E�?���2w�H?Jŷi�ĔHqj�Z���OD�������'�	/(ef�8dF-I�y4b��m�d��޴�f���?Y-Ol�?i���#�਱�h�}��	�fE%WiJ��4�?����?���
�B���NyB�'���	�"u4���R6Tj��Y6&���v�' �	�m���)���?��"unm�pI{�A��R:�����i"������d�O�˓�?��6�,E� ��9V���M�'S�TQ�'�hʚ'����X��͟@�'�F���[���ȁ�fM�v��9@��P��등��O��?����?�Q%<N���ʈ/we�� �.S��̓�?y�#�\�{��?�(O�K���|P�718���> Z�ؗgYԦq�'��S�t�Iǟ\�	�%f�i��G���(����
[�8к���>9�"�2�?!����K�RM�OpR���k�\�h�*�Uk�p�$
�*EA6-�Ot˓�?��?)���<-���K�<:9"�$�2t �(@M�&�M���?�+O��1�h�]�$�';�O��D!w »J�z�3F�J�V��9�K�>!���?��w��Y��������Ew�U��)m�Е���Ţ�Ms*O^�떾�6-�O����O����e}ZwC��y��ѥi�] C��=��4�?��X����?�+O�>Qɑ�ɅKHJMz�@V�K��L�2*xӠ��bi���	����	�?�)�O�˓pL�- ��.p4� �&lN[�4�лi^졂�'��Y���r�h�0p�F�ӆ,�>0I��%���պi��'h�ᇧXE\듬�D�O��Ɇ0��Y
D�K���Εt7M�OD�l���S���'���'��9Ѝ�~ ��p	�)Ao ��tӸ�ğ��,�'�����'�Zc�K�5U�|��m�����NayO�<,O���O��D�<	T��@�j�%���OHP��N��_�n�ʓY�\�'��V�X����|�I� HBu�L�ܑ9eL@
o@�P@t���Iٟ@���@�	Jy��݁B(�ӹ@eD�2���7pf潙�"](�(6��<9����O2���Oj��G7O҈p�(��>���g	�I)�q�C�Y��M�I�����<�'�����~:�I:P(G�5T"$s'�P�Ƭ�3�iD�W���	ߟ��h(��i��(F��(���H�ma��u��6�'�]����'��I�Od���8�uKA$l�2��e���3F���S!U^}��'U2�'>̡���'��I %}�c�D�y��#�JM^a��T���d�݄�Mc���?i��Z�Z�֝�h58�3��\�Km<52��d�Z7��O��D��PT��Ol���O�&�X��֨6E:}�#"ΕR����4Y����i���'���O��ꓫ��Ú[�H�Ks� '�Uc$�\	f0o�9-f�I|��I���?�pN���$1�E۴3"U��5f�'.��'���f,�>1)O
�������Ux�F��E�CXz��2��x��D�<�CM��<�O�R�':�	�(Ю���#
Z�M������'D�H���>)OJ��<���ի�]F��*�A=K�h�P@}�AP�y��'�B�'*�P>�I'&�t����g��wo�y��اEI���Ħ<)�����Oj���O�bSb�28����N�"�rl �B�	D��O����o���$�O��{�0MS�>���R���z��!e	!!��������O�ʓ�?����?��*O�<�RhőMM�0Ձ�1_������>*���'���'jR�Hz��<��)�O05i�#��k�<]�LV�-��)�b	OȦ��Icy2�'y�'����'���O��CO��?P`P��W�O���J��i,��'��	�L�E�������O��)=�NĀuC҂P�&<�`DL�cn@�'�"�'c�+�!�y��'�Ɉ1N4�i�{E0-Jł��.?���f�<ԛf_�Pi��M��M��?A���dQ���"P^�" ��T�0�� �j7-�O@�$3p}�Vm��'�q����Ǝӓ.!��8s#S�vgJ����iNT�r�Id�N���O$����Ƅ$�\��7v���a��ؗrB�����,\�dp�4�ܜ�������O���(�BER`��L`\۳!��bwd7m�O���O��B�Ql�I؟(��g?IF� j��=�'��	�����ҦE$��[��h��'�?1���?�  �%uQ�xIv@J�AZ=�P+[�@���'9�ԡ�'+�	֟�%���gT)1"���5�Pm�ƥA����/Y^$�����D�O���O�ʓ{�h�z�J1=iFyq 	ADl�� 4i�x�O��� �$�O��d7��e)���1A�u@���.hs7�d�Ol���O,�=B\��=���Dˏ�u���faء#q u3��x"�'V��������$��x� ��� �a�`* e �jc��=����O����O���L�����h�<Q�R��A�8̐U$K�;Q�6-�O�O���Ob�a4O�ҧ� �A���8i�� �a/�@ɢ�i/��'W�	3ns���M|z����K��X��V���'�d��n���'N��'�6Dz�'��'-�IR7@��IX3lĞ��:4��"��X��D�
�M�#X?��I�?A��O6��	�77�U�2��
���"�i���'���c�']�'Tq����t�B��	��虁X}����i�\-�pu����O������&�@�I�K�V8���V#qeb�j���0N�2l��4A���c�����O@�i��/#4j�.`n=;B� �,ho�ȟ�����)t ����?����~���o�l�z�f�-�5i�\��MJ>��K44ɉOQ��'PR��r"�W�q�N=��H�~��e0ǰi���R>'��b���	g�i�y�Ə�>{����J�1P�Dü>�p��<�)O����O ��<aË[Y�xx��܋cDڀ)p�˻�dAP��O��O�$�Oh�(��;'(��R2
��)�s.ҳz��<����?�M~�����<��IW<%N��
C�Z�y]^���\���	؟�F{2[��I'b��C1�(I��]�3	�7UZRŠ�O,���O���<�7�ܺ�O�P{�!�����q�L�"�&-85�lӰ�=�*O,�2}��£<�P�wʉ�� ��4d�<�Mc��?���?�Ŧ؅��ɲ<���Oy��[&�[VPbqJ�i���`��x��'��	�@�#<�;i��T W�b@��%��2'���l�^y"�[�	��7��O����O����r}Zc{���`�\��� ;'�!Vi� �K<���hO�'O`1blѕ#
�hG�-G��@Qܴ�)����?��?��'�?1���	�� �n�V�,cE,�{V솷Tݬ��'9��Ѝ����O���KX0YJ��0�j���b̘ڦ�IП��.;��H�O���?i�'D +4b�)N��9
s��u�,�j�OL˓k,���D�'z2�'�
�X�'RvZR�k aV/5������y���D�a���'Q����'PZc|���3l!�zt��C�`�#�O���"2Ol���O��$�O*��<ᔁ�= �I��(r��i?*���4R���'5Y����ݟ���,%$�0�R@�L(����G"�QD�c�L�'7B�'��O>xa��(q>�g/YU�b5R�^:P��DH�Fn��˓�?a,O����O@�$؀P���: "h�A���_�lY��7m�O ���O����<Q2�ƯxD����ؽJtĝ�%��8�Z$hue�m��6��O���?���?��G��<����?Y�aX)3��@�"�Pt���x�:��?�(O@x�3KL���'��OBfh��Ɉd���:�T�p����ͻ>���?��)�T���ɧ>)���� ��5�TAH��x����
�
_�7-�<i� ��1T�6�'�B�'����>��P)`�!�.�"J�2E����uoZ̟`�	$���#��9O4�>�c���pEJ	2�C�8 6��	Dt����Ο����ϟ�	�?(�Olʓ`�+
��Bp�{q�#���� Φ1��*g�|%�����;����$���|�h�
�"�;�$�;�i�"�'@roY�~�z�����O��	4<�#�dR�hG:�JQ��A�@7��O����8�S���'v��'���hՆC�Yi1eõh�y)�cp��d��4,Va�'4�ޟ��'5Zc�J�B8�G� '6�`� �O,h�;O4��?)��?�,Ob��G�h�H�[6�η�,�A�AXɌY�'��ПT�'~r�'BR+�x���0��G�;HNl��aL@���y2�'�B�'�削(.)��O����@ɕ:�lݨ'±~zA@�4����O�˓�?����?I�<	C�K�U���1������A�M�#���<~�����ݟ�'����S�~r�U���@.9w3�LK'͂�A�Y��iz�_���������0R�"�O��V�W'��ш�+�x���ٰ%ۛ��'ir�'0�)'.��̟���?=:�NO�9��eb��*� #�ē�?)��gcR�Dx�؟Z���!��)�$�����<{�\��[���� \(�j7��$�(-0�e�G"�#����dNQ�G�!�D[�-_�ؘ�dQ. ��UCӨ%����Ŋ	aX0�@B!�6S)��ҨX=}�H�ǆ:(����A֦9��ep����&�zc�.��Vb� DܟC�iˁ-�+@�Z9:!��|\���䭒�
��h�+��~2�u/׸�~x��eZIr:�i�!�^���	E#�uy� �(D�R��O���O��d��{��?���o�
�A� X�.���
�+[�NLM��0d^���*>�p��g�'�tx�/7A����JB�Q�2Y��	�O�̲�ơA���sw�ޝ�����@�?TT�3�@6:t���O߁~���^�$'"�'�ў �'���27,UB�e$��'F�& �'u~8Ѝ�)ci�<I6H��<!$9�8��|����	�u���n�?��ii�D��޾����/
xH���ٟ����xx刔͟����|:v��`�a�phR�evL���D*6�fa;��7��S5AJ��<�Q
T� �^Mb6C�W�1$Ck(mK�M7'8Ds��M���<q�M����	 8 U-ږ(�BP�p��h�l�D{��I?�0�pF��>?1,L#��ԏ`5��!�r��4�#L��gX:�$KL]��ϓF=���'��4�P<ꭟh��|�q��A.�`jGl� ������O�o�Б����?q��qX&�U�1~H�T�J� �*�� H���kZ)xJŎC�GѴL���ɠ^���Չ�Jd��C�N�֟�åk[�\��L�	�T0ʣ�_"��J���,u���O0�?�IG�P�T�Y��^��jx�\����`"�g�U-o��-�׋�%+���hO�A�ɏs`�	d�8��g� �V�I�s�����4�?����	A!��$�O��J:��k�A�3l|`�+�70��
2���|8�J���T>1�|�	�y��|�H 69���B�FW�&;"`�̇��Dܢ �V0	�)���*�Ũ2�ČW���(+QN�.1P�Iğ���'��B��<�BI��3'^7-x�ȓr�V��&ő%ɪ`ˁ�ëU��IGxB�-��|"��x�W�X=Ti�fh $J+�����?�S���y�A���?���?�v��<��O� f@̣B�,��׌�r�nӇ�O���$�'\��v)�,���!5k�0I�'���y�x�ȔC'�7]�����S�4}��"����[������-&&^x��)V3?lX���+D�iS�$tR 5���5����AH.�HO�)2���2h��mZ3
���`�E\15�~�#g�؂$��t��Ɵ<�	����6&�(���|��	��]��.�lWx��'ݶb�:�`���4�N�e�'���d`��,�Q�G��B.A��&�"<I:�(E�B�Ev��ĉ���'0f�����.K&}�6�Q1Nh9�E�@�'�x�Bυ5�"(�ì-Tx��[�'�� ��܊y<z�$߯au8x�'�06��OʓYTB����iB�'F���l� l�M��jg�Ԣbϰ��ņ͟�	��l�D�Yz�X�̉�FM6��S�t�ےK����%���0��)�_�(OVYy�A�j�V�¤��(�B�o�+� �RQn�1'Nx��@�\`�<�1�� :�Q��C*�O|��#�)�OP�4&HF}�ه�	h��I�O��"~ΓLֺM��b�w�P���<����'-ў擣��T��;DI��j2�ແ��?��M�<�ꍠ6�i3�'��S������П ��&]�e0��E�Y�-��a�S�P-·f�M��<��O��h��(�攻w��3FP)��Y8������O�9����]��$��W?���ce�� .����OB��?�F��D�%:�"�w�\Hhp�8�ϓ�?��C�� �����74�k"N�q�'�:"=�O.��$E�x9���0����"&�'j��؉"j���'N"�'"�wݕ��Пؐ�W�}�l�p��2��������?AŊȠ7�H��Ŷj�n�3ړABTq�!D�H�9�ň	�kBl��b�'K�Bb��i��P�5B�fF{�+N��P(� Д6by��f��~B�B��?���?���U>�Qf��O�ޥ�f��v�l]r2�0D��z@HZ�ʹ���	:\z�P-��HO�	�Ofʓ	�0a�i��C�Kˑ>��Ջ`,�=1@p�Q�'���'��e��	��'�rLħ9+n)B��F'G䶬��g��Bd\P��*] 
M4��]������=F*��7tSS���/�\�DH�u0�J4i��p�F�O
�DE�v�D���N�F���fݞsS�8l蟘�'���4������v�B�S�N��̒�+��N��!�I�6Q4չF[�S�1x$���ئ��ܴ��'�r�|�N���Fg��Zj��4�y���s�jP�$�Ƚz��Ǣ�<�y�m@�udXMRCǗ��p�#����y�-4L"��������.O�y�MC%���0􄄧KP�S��y"��$k]6��v�Q�r�ra�t��yR�j��̓r,϶zn4��!�:�y�!7l�9BU�t⨐B�LV%�y)�q1d��ыH�r�J��#i��ym�erb������x%^$)�W;�y�`	�W����Ǒ�hp�t����yA�8���[�,�d��wcM�y�GC�&�d�;AndZ��8�.��y2L���� "� �i�V�n���!򤄓Ay���C���8�T+��t�!�@�n�7�k�H- ��Վm�\B䉁X��y`���m<ZW��r\.B�ID�z]���
�g� ��D�E���C�	�^�3v�p��D!*�,7�B�)� ^}���E37Y���$:<�T�G"O�d��.��T-���!4"O�(:4K�-)��P�TA�!,�t��"OR����/��]q堛�u��+G"O쬈�aE�1����҅�+H�DX�"O�k�偞8�|�{���5w� #�"O�ѫfHʹX��l����=qP �"O,$`EfH�z��qBoB�$��9�3"O�����L�ck���L\�tנن"O���s�f�D�gLYP/<%y2"O0�g㘉TYJ��m�;�"O���a.�:K 
��!nthb"O�͌+qBɣ�R+5��;D"O�:3��=v��EB��Ci튤Y�"O�%�m�CO�(�Ge�3}J��'"O\���c�3�d͟^5����"O�q��T�2����E����Xj�<OX�i���X���`��"~Z�$�?�<�SE�W�	o����n�<����,\O�g'��"3l��Ëe~��OMv����0<9$C�)}�̙
�
J�'�hh`2��H��Ypg�#�^ �ȴgd��c�-x�A�t+�
�B�	�vi��K��	+��!�K-o:#>aS.�}��aabD}̧3�|�%yn�@��EӚS�.D��D�Pk`	�=�J�J���ky��͓���èūp���秈�Ft �ė�&� � I%��L���'7VT@s�� `������ߙ&v�y��0Kj�zo��9d�����I,���Ň�9猼�gدBF�?QpjN\��[!���e��V����է��	0D�0 HH(��C<9� #&�:��@�5|x5ؤ��uy��B�t��'O�8 D�Qe?�|2�뇠)�a�􇀨G�x�1� ]�<y!��F�0E�y����e�<!t'�
Wl.�	4��T>���`�|~"G���r6�/L�i�-[��?Q�G�%��Aw�K>e��T9E2�T���b�>9e�˓ :�A&�n�D+!_�`���K+<�t`�5i3�x=��3���>�BkӤl-����Īw�~�Z�m٨P�,�hĥ
�8�P����@��A�����X6�}j�19Y�ٕ'Rr��w�Xb}�Ȗ5,���S�',�q����(02�Ȋ���ąȓ�2A���W�N�}s�GQR &�\3sG	Yay�D�����ү{;02�΁��?Y��@��#K�A�ܩBW	I;1sv@"� !$��+B�U�w��D"�`�2B��Ȣ�&'��S��R��1��� ��9�5J�~p"q�L3*�H�D��#�~"�,v5f���? ��R���DJb`�X@H���5���`L����%��'g*�;���.q��@���&�y�#�?y�Ik���U�tS���5�~bDJ�DF<��3���IF�`'?��7���	��ӟf�rA#�	�$gvlD�kMV�DB�ɝb�bx��ǂ0�5X0H�?��x�E�s���Ѣ�5g�?/��I`pF'��4���L=,����e�j��)��	�V�2���)�䎇��Y�"
DJ�-Jf ��B��yZ��Ӭ8v�)�(J�P�F|"K���4��=t�$���1ᰋD;���7�  ܁�"O(M!���?Tݢ7� :��:O`���K�:ZPĩ�n�a�ā�7.��a+�E�� 0�F�y�IX;B��4k�j�C��R�l��w�����dY�$��'�N���OjLy��Q���]A�B���M�1�'m&КSk�+%�^�R&�.G�H��B_([7����%�����ɫf�Y3�	�f�.���OִI��#>yф+ 5Մ�X���O.�!
��V�J5K��R�(�J�'x�lJ��F�|�@iӓK�t����ن4Jnu��/	!6<��G8+��m�S��ߡYegOTt��a��׫G�Hm�U�;D�Ĩ��ű	ZL��3a:'TXŊUU�d�4Ψ���O�p�AF��?a��'��H4�q�� Ku�K�&�ƕ��yr�[�fƔÔa����O�š��ڸ:x��3�Z�x1 L>~���y��G}pP02w�E��ģ��Č8 ��!6 �-yX���C	K��h�8"��">�!۝!6x�S�? \�G(@?j�=�p.�:Q�x��U�y���.OD��d$�\��V)�c-�@�=�:��=y����O� p�4}�� /L2�gM��R�ܐ �)��<�3Ɗ87%�8�%	�9���dE�!N�ĉ!AU9u(b�IB�� 1Ve�x&�:CI�˪OT�Q�*��T�D8	;�щ@i[-{��s�,�z)�`��>��
I6MtR��
Cz�(l���1OL%*3�H/,F��G�_�C��I+$�]��D��f�O��:����&zL$(7�X4o�F��C��ަI}½��� �3HV��!#G2S�l��/̛�
8�Z��O��h͟����g�:��1;�O�� 8W�ޅj�v�����;$�WPa���U,̜iyz�0GN
zM�B��2OfL�ѯH�2��j�@:_�t�o�N���A�+��YՀ��\I���䅮Y��h�F@�dz`�r�G����S&�ӲgD��j�\�Uh�ɷE�<r� X�F�P�����˦I���	�'.�(�d:u�x H�j
 #�ْ(����s̓hh���"T����qB�,�<ySo�F7Υٶ��-0B��C��VAiv�T��M�J`Ctq+���Hn�I�eK]ܓBBy �mZ 2A��@L�v	)�(�'2Y� ��-4A�Є�Io�~E�&BC�|RVX��H��G��y�u�O���!i�e8���Ņ�|!�Y"�%
���c�#,O�(�F�%+
���Ð'}8�q9u(G;f�6� �[b����:���ف��L1��8���4�� 5/O��Z� �$Z�՘c��� R�&�Mn0`#���6�G�Y��EiҨ
�)� �@���.�c��/U:�`��O�o�:�b���H�@9�� {F�9�<�W�߽ (���-�d��J�$V�Xu|�ɿ,I�%�D-G
fq"ĩ��N T�"<Y���1�xI��Ğ�s@�yȀlL�U�
aD��J��">qvX�?�_�Mq�S5A:y�����$����P�8R���,`���D��}�Y
&�T:������S7@�4�'�d6��] ���*�s�֝&I{�d!�Iب]/�͋���"����J$lOڠ�Q,ƒC\����C�"�Q�A�X�@����Z|� :�#។��dӼ]m?{ ��V��y�gd>˓P$UQ��+��	����G�pe�>i%���2A�PM�<�W�擾9����2�F��d��j#8:6MF3�f�*���O\� f�'8 �J��[��p��9�hd��R�t@s�����S�	D�W���b�w���+����G��a�_�#3�f�^H<Ѱ��?L�Q{C��%F8�Y�@�K��	�w$JX`�'m�iZ����Z�4^����ӌ�7 �(�+��pg<���I�t��9�!ϟ��w,@�qO��B����ܤH��!�>y��'nF�0pf�t+���e[��R�Ez�
�3w#~F����4~8�=B$�M%�HԳ"�Ǹ�yb^S�,��LU�*-mbRDF6�~Ro��O�>yYgH�d�����ԧ"Pp��B/8D����/� ]�$]�T�s�\4�rI+D�X��.Ѐ��l�?XM��(D��J���b��]l�57����"D�<�����:l8�+�4A�l�D@,D��X$�.(��dƊ �{
����?D���ѡ�:�m��L�*G� �k=D�Љ'@N%�V����Au���!��7��@q��z"��we0	F�R%{�$)�C����=��M���?9���s��*��Ѓ%H�&.���b���'u��v�0\��5`	#C*8y��dI#��,e�>պD`(��yx0O7".C�I<z�rG^J��=CRb�NGV��ӡ�O�U�K�<���Oָ������D��#������"O�1��(�AS�� e�4C��'��-���'6�I��'6x�� ��z��0aN�x=F��ߓ����y&X�@K�q���լ��Np�ɶ��y�#�0��p�l�6
��;3nҌ��Ol�p�<�'p�&��!䙀Iϴt#�j�H��ȓi7�A��t�����<d1p	�'�]x���Ӑ$�*L��4v{�S���#�HB�I��qR`�O�B�qW�'k:�OR�1�-LOĴ�7K�Z�d�9V I;V~�lsc�'Ԕ��K�t�|����ɲ+���GD#!��͡��Q���O ����F]�\Bax���7�OV�� �V5TR�����*CP~�;C"O @Q��68�mԋQ <5\x "O
(SH	� �~U�u�ֺ\@��"Od�A�T1�\`�藸y�n��"O� ����l}:D�"��"OԽ�EX�|�bm���8	��(!g"O^���&l��,x���-Ѵ(��"O���Z#dl5K�c@cD3"O���d�	{����ȡB�rq�'"O��2rVH��}�6�W�}�,X�>�pmŭJ�O���C�g�l�b�A�N�����"O��8'BR/#\�Dģ�,�F�ɤ��FX+�DÓ�����*�����D����y�襋JF�b��=�s� "i���A�R�|�tB���i�ڈ�*?z�����ˆ
�f��d�\���Z�yү\%_�03�L3a��:����y"IJ�y6IÑ�ә#3��
�b����ɥ7Ovȑ����E~�R�B x.@i�h��NU!�C�Pc�X�L(����\d@qO�X9�
0�0<�+
�F驡	�a����a�P(<����@��0,ԑXQh4�:�D�p�%�0��O51��Ra(ڗW���� O��`BJ���'���"��>�~TǨA�Vݜ1��'$�h[nQ YyV�@���P���I<�F�9��O���Q�%���4�h2�:8�:��3"O��A5�B�*V��b!XG"O������)'�,���
�И�"O�U��
�	9��Sˍ.9�4x��"O&���#�-c�� L�w��1��"Ohu�tgY�\^B�ʐ-G�.���"O�	�c�B�&��\��BZ��̊�"Oa�e�҅O,�0�ϥ0��	'"O�}�#�6u4��p�uH8��B"OX][�9��ћQ�-F�`��"O�M�EC�>V-R�0��ɳ*�h�# "O\D��Ct!���,W4`���"O��hS�&i�VJQ�<t0��"O �ۢ�>Zp�ꌘT:<�r�"O2��a�$���GI$Y,*���"O��ѱ� �%tux��B�I-��"O6����M�,r��b�Je�`"OV�۔�Z5
d���%2|�Z�"O`�� N0�p$cRgН,!s"O�2o˸¦a+����P�j ��"OJ|��؊%2��n���ٱ�"OBU�E"�LT`vm_4X�� 9e"O���D�_&\���A�H5$�JА�"O,�cG� .D��y���'zRE��"O��#գˈ;��cFC�h>!1E*O�u���09a*`I0��E��'s�H���V qS��c�z	��'8i�@b�5�p��R�Ba�&i��'�(ț1��)G �7H!p��I�'�<���Oܮ�D��F�'}G\�z�'�b$xp�D]�ٸ�fR�G�@��'�������<@�
�����5R,t�'���� �^�^A0�"K4a<e�'%�,[	�!�H���
%hd�a�'v���ǐ�omչP��p �� �'v^Mѕ��H��1{��VBB�C
�'vXd)Vm\?`����F��P�9��'e!rEY��ɋ��ݻL�~Hc	�'N�ZS��"t�j���m6��@z�'#�h�Ik)$S�T
9��yJ�'��!6 �is���F�
E.���'� ������w>5I@/Q̔B�'h(�����^��K��(JW��p
�'8fU{0�S���\�协j��uQ	��� �	�2�̐8,٫2E�4h�vQ��"O�3���#��`���(.�"O4�ЍN��ؕ(T��s5ք3�"OB)����W� Ir�#j��H�"Ozkv���u� �0
�6U.ر�"Oh�k2m��4�|��"J� X�=3"O���DBy�@f	����"O�Xh��ɪD˒��֧<f(Yj�"O�C�G.e�⹀�)Z�P2���"OL�ٶ��`�X�H�h��	�b�rc"O���⊁g%'([JtX�@�"Oؙ��+�����i ]!�D�6F���@*��yjl���[�P!��H�!*���v�<Nf\�a�F]I!���ޱZW� 8,H�9���x-!�d�K�|ݙ�ޔ _��`�c�#1!�"��Q ���n@P%����y!�dB-�@I�l�((�z0B�r!�Ă��p�"L%�B�����&&^!�DS=8
�kq��ȩ0Bоu\!�DHb��=�1IE�`@t�V�;O!�@�HDS%LK7w����@K:S!�D��CJL����� )��5�`_�^�!�D�Fhbx�P#Vؘ�X�/Y;!�*����x!�`�� ,�!�� 5rPa���j␴#)̬
g!�$B9��ݣv$�IzЍy%GQ'gX!�D�v@����=1��a��f�<u!��Ȕ(]���de�D�$��Ȇv]!��9W�H���3t��!&�ۑ?X!� �_������ْ{g��v��?:!��f�9ULжE9֨P�G*!��Į	u���������&(�� $!�Ė"e��೤��C�x�r,OQ!��U� ӊ�3���Jm��KR!�䜎?��X����"L ���CB�!�$����hZ��Y+�$�UB��u�!�ۙ{�	��n��r+���!�xD!�-��=˄�C�����@�=\a!�$�;I��� ���!�sN�,`!�-:�"̲q"~zxL���˪s!��;x��g��xڞ���-�<r!��<5����wH�?^󠍜���~�P��4�ЇK0:h2����y��7D�肐"�67�Z��F��-!�@���+D��"Ѩ�`��'LK��#��5D��J�b�h4;q�ĉ*6`|�q�=D�d�5A�I+�ڴ�OVl�{��;D���v��,z�L�1�Ωmr��2�E:D��R�5�(��̔�И铫9D����(Y�yqh���M'�C�H6D�T vC�9Y�q�#͖<G���c�2D����V-�&�X�@ʓf�@= ")%D�0�S����%!o�!S�6�Р&>D�X��aP&r��v,��rq��6D������q"tC�@�	J��� � D���ǥ
,�Q�a��wڪi�b:D����D
;�r��P�@��!Hb�4D� `�d�'V7lk�iA1jr���N1D���@�E�e�~���[�H�$�lp�h��I}1`D��	�)Ǯu���j	C�	
7*�PЇ!�.Q�u	��F�0��B�I�@C$��mZ�s��je"E���B�? ��5b�M&a���Yk��"��C�)� �Q�.�5.s̱sы 3e�"O.4Z �VN�ig��9P���"Oޑ����Vl!')�ɳ6"O�a�u��a��c��S��l!C"O��a�j�4.�#+�Ȃb��)�y2�Bv.B�%M��d��↛�y2 �R-���TEP��8t��M���yBCS�g'Ty���Dt��ި��%�O )�-O�pߘ�x��]�V>�s"O�h �.��j�t#��!n$>i�"O�`�Ŏ�>D��-�"� 	�˗�	n���)�[�bI��,]A �;���"z!�� ��Tj�B'e �ы��L�<�!�$�Rv��K!�4_F4)�$>]x!�d�x(�0�䤞?J �l�B�->q��=E��'��|����.�v=�����	��]�	�'�Z���	j���J0V�	�'�h�k�/ȏPppa��`~�X+�O��=E�$��+iQ����ɡ+��ً� ��y�\j���O�)7O
ɸ��L���IGX�`3u)�+]�r\���
�XǼh�J;D����حR�69ٰ�&������:D�laG���^lz�	V���L� !�8D�d��ݒ7��8���2dj��D3D��B΍�	�M`w%��6"i4D�` ���[�̈�6O
�aN&M��*&D�̃�+�HB>����/Z
m[�nȼ�hO?��[+�0�I��! �T��lܪ|&a~�Y�dS�F�d�N��쐈1|��8D����5�N8y7nPsRhaE7D��ʡF�7�@i��?�T���*)D�� ˝9���&��yB`<�Q�1D����7��0�M�P�^h!1=D��h&��n���X�E_�,�bq�0D�����֠G��y��F �C��D�b�,D�d���(tF���3 ��4 ���>D��h�f�z�H;t��>z�a�n*D�X %D�c T��BH�F���{��3D� ��#�\���I�#|�ޭ`-1D������"�؁�E�!0)�:�)D�8�C�!�>�8bL��e����w�2D� � ���`��@����Δs�@1D��0'k�38�3�.�f�}��$"D��!T�Q �5Z�NO�$�ne�G?D�D�T�O�(�����Ad�(�b`>D�H��䝻e�<��/�t�"�
�;D�����N�/��|#��t96�E�9D��z%�!#!�%j�n
�%~4�b��6D�p�ص}9Q/M
�6)��5D��z6fќ&�4�KS��T�����0D���ˆ.x6dA�`jקS9�`B�(�O��<ЊȪ�ꭚ�)X5!i���Z^*m0 $;�N,#���'!@���]��t��X �1C��1�L�ȓ�Fm�u�-i��IH��*��ȓ4���h�NZN�)���ҽ 7nԆȓ?����"&I�~���Xw�5a��1�ȓ)�8�[y8 �&�_�(�h��ȓ�~x6�D�e�*)�s��H�L�ȓH�D�:�b�/EV��n�[�Y�ȓjl����	f�6P�3�ݎC�d��r��x�gW�L:�%Au�B|⮰��tgh�����:�XI���
C����ȓ�]U�O�L0ݸ�e[؄�S�? 
�`S��M�Ј*d`�8o�"�ٱ"O�����U�Py�u�I�H�s�"O���0c�7co���c�o��b�"O�1X��b�8�C:u�.�"�"OHM�*�%�<D�Ԙ5���"O��HT��;G�`���7J�`�"O\ D�z� ��&��D��iR�"O����\ l�$���ۚ8���ا"O�XJ��X.A�5����/��E�"O�,1�(ZK׺-J�×�k4���D"O&�(�k�L R�I�o�y(�"O�`(q0I1���q_�E	A"O�������U����!�PG�]�5"ObH��bϝG�$}�T�#v( "Or%Ӆe�*|��Ĳ�+��U0�"O�m��� a�ܩ���A4G�z Y�"OJa	�(2$x����;��Ih�"O�(�G�@ &lZ�E�3q�ڰ�"O�X�NM$.`�����-z:A""OX��r�\?�.e &��=9�Uj�"O$�+��E�\�"e&F�",���"O��#�g�
+� Y�J�5 ���C"Ov@���O'd9�E�HY� ���1F"O0�1D���N|3�,�7Y���*�"O,҇͘�2wZ��k�-wv"��c"O��K�W,�1)��=-o���"ON��֪߿03p	sQ�5}m��'"O�(���Jt-�R��.KZɉ�"ON�Ѓ��\|��o H-nG"O�0�bk�/TT�a�K�o*�H$"O���W�]�Ҍ��E�fun(Y�"O�i 0�v��p��	 `{����"O�s~�M��'�z�J��%��`�<Q�Z�\����g���&��"�EO_�<�Cg�h��8��f̳����`H�Y�<�u�L�8@�<AU��8N�a�Q�<	q��]C��X�*�,�Ġ3I�T�<avo.l���H�k�&O�PШ�ES�<�w�ϯ<P�@x�'�#m5��q�!�K�<!g �%z.I�
@(~���P5C�I�<�`�u�P�Rs�-Z�����M�<Q#�D�j����؄G(&1�ee�<�R+��"�9���[�>����c�<U,�j� �����d{��v��e�<9�B�9(��u�A��kJ�;��d�<1���m��T�v#Rlś�K^`�<��P  ߸���l��;p"d�c�<�A���V�"=��� 
�&�SU�Js�<�"�R�W�1�g���k2&I��+�m�<����U|&���G2
J`���Op�<i�M3[��|Iv�P���R�ʁa�<��^;�`�h�ā)@����+]`�<q���f�����f=?+@+N�C�j�R�3���]
���D�P�2C�P� ��ݐ0��h-DfC�˖�ӣx�^h�G�Y�FI�C�I
!�X�͕11e 4N¶^��C�I�0a�="F�Z�����L��
�|C�ɞh�@�������;��A0 �FC�I8�41�'o�:h�h�F��0��B�	�
mh=�p�L�p,�]�7(�#��B�	"�ح�BխCZ���p"
�96�B�I7l�@`س'�S}rȧ���*B�	)^��a�@�c�2�����+VB�)� �<Zp[VFy1��2O#����"O �n�PC�@��ܩ$r�D@�"ObhJW
ܺ/DxR���$i�tp#"O=iӃP�D�jG(ZJQ̠�"O� �e ���"��T�4!�s"O|�9%�S.;YJ� ������y�"O�4�7`ؕ1�\�2�᎓2 �4�"O��j���1rL�󧁈�1�D�̓"�4��R��#�M@���F�<��)ߐ��P��� h.ua��6X;ȓT`�(Ǭ$��X����'(�����+@�x�Sp��"s'3@VD�ȓK����4�=C2� (u��x�B�ȓP"b	�h�"	V���)��Z�ȓ'-�!�3R2��D�0�^�ȓ<��i���7(k�АƏ�	�	�ȓ`+�)�p��SNB��Ubߚ2�|��c1@1n�3,��ŤU<�^0�ȓ$$���EDV�����:@nA�ȓbd�4
��ɃU#.�y��<�Ņ�I�~�	H o�j%y���]0��ȓB�(tMU�*9�P��
�e}4фȓ8p"���]Z
9�Ы�
D⪔�ȓO�YQ��a�@h��i�=��4��Os-Be^�k�X��ЅèT��ɇȓoex`�D��
$3��3,�	b9)�ȓ5T$�"QOG��6���+y�tx�ȓC���Cު2����-V�e�A��6 rTXU�QU�j%�ԢB'R@�ȓh��}�f�_H�U0�h�$rDr܇�|(p��S�f��% �W�.X��ER� bД��ys4#��@���ȓx��P�X�0��p��&�$,l��;LIx���l��U��.X�I後��;�0�#T �)3�.���X <����NI)�f�%����oʳB4lцȓH(���I$W$�����
~-��b,�J��5,U�f'�Fژ �� �q�����Z��rh���.�ȓA��J�4m�l�j4���/��ń��B'�6q4$`��M5�ꍚe/�G�<��*O�r��2��+�����\{�<�A�D&[	ZYIQ-G>J(�����q�<�����B�1���3D^���k�<�7�J�αRS�ڬJ儸�b�i�<��D�π=�fȌ-j 2���A\o�<�Ł_�h=2!x�@1,�Вt�F�<�����Wk��pf�
�<��t�r�JX�<G�	��Å�ͪd@hB��V�<��B�2��Y a��	T�<I2�&�Bx�FKz/�x�%�S�<����b��i©̚$a�(�d�P�<�0E �uP�{!	[\����"L�<���w?�٣��n��j��J�<eΛ*#d���@�U�	�I�<Q�.L:Q �b(��o[����%HE�<����)�L"7bD'=HP@(�u�<�0�fP`�M:�"	3�i�r�<��C\�jb|C DV�E4��t�<���6�%���	�_w��)e/�s�<�fa��T
������4�x!��z�<Y%F�R����� y�cPw�<��d�"q�41˵.0fqq��N�<��Ə�
�9��~�|�ڕ�Ea�<� ̈� �]�u%�)�$�-u�C�"O@8j��F8w��K�)D�hc���S"O�pjc.�^����ɴH}���"O6!2/�2z�M"�4n ���"O�4�!@	&;B�I��;�np�"O�e�P�3z�y{F	/dߜУT"Ot��d^!5�$k&�M�x�z)Ѥ"O0�$Bo�p�h��uР��"O���L٭�~(�A�ȧZ6�W"O������O�@ "��!P"O衢ϯA������H����"OZ�0�_�~�8(k��֩zY��8�'#l�c��ER$Jw�P�9��1�ȓ�ձtM^�3�~�9ԏ�	p��q��=O�B�M�O��Py"o�,8�Ć�����Pk۰v�$A�$㙩H�ȓ;'Bq����.u��(M-*���ȓt@`0d�p�hY8"�̭_��ЄȓkrR�� v3N�c�ʛ-6ˠ���m��͐� �4��k"�_-~H2x��B&�-۶�
9o�tm�0�Ʌȓr&������<���L�l-�\�ȓJ�\�%���	��s�!��. �U�ȓh�~qZ�Lۆ�l��V��H���ȓ"VJE���0G���j��\/m����ȓ��[�x�ਠ'���v��ȓ!�>B��7!@{'���t,��:�b�sƥ�.ah2=�#�O:�U��HQ�xk���2�~�A�\%n)�ȓI�y�vA��*DS&��Cx��ȓpS�5�@�]N�s�"P�L�v$��e����֖huP�JG�ǌ/v��ȓj�f!a�!6��mz�GN�,gJ]�ȓ�~}(�;k��Pj��A+~�ȓi���� �5tOf1�BC�&n$���$�t�&k�� L z0I������V�:����)�D艒n43� ��nv�d��.��a��/R��H��C�����)X�-�r|��C�o��}���Pm"�l����9�
�+T����ȓS��q����^<��i�^(H���ȓ'�BAi����+�؍���Q�`�Jфȓ6�ʸ����%1���J���%�,Ąȓ\� �����[e����&��L��n���SlߝZ�B���nR��ι��2?�x`�&E�V�q�KǱr�8X��x��rN�T�C"�18"ࡇȓ2m@` &J˻,�Pl�G�ѩ#�:�����p�G
�@���%^,���i�(����"a��ۧ�� QrX��+K <� ��:E%rQ�
��O��ȓL?5�¨�$A����be�t��-�1Ɇ+��k�"Pe�l��ȓwhx3A������\�&��E{��O5 �5 �o��U��_�v?�h��'��E��H�8��!(M��k�B����0OD\R�b�-�0v�(�b�HB"O��(�e(�T�A(WL(	�d"O�\a�D9>�8��P�V�j���"O$�a1m�B��(��Ј�`% �"O�}����=�<�cc�.l���b�$�O����O #|�,O4���K@&��ÚJ�<a�8[[�lSm�
��BѦʟF{��	\���hڰOF�M'D���T�05 B�)� ~l)���Ĵ�� �Q50��"O|8wϓ�apָ�AȬ,PB�"OXh��]�ȡ��N��A���"O��[�j�� �Hɣ��ˣ�8��w"O���w�'�D�2-G�N�q�&"O,�s��{P�\X��!n����"OPd��U�@�1�$m�5{w�J�"O4ݪ�뛤>i�9!�M+FZl���"O��@�Q�1�0�̙<R��a"O~��M�5ui�=c׫K	qG���U"O09���v��YF��>|8���w"O�	S�%5*���P30��a"O�ES�ЗR�D,�p��,�T"O�P�eb��(7�m+�!2����"O2���2  ��*�@�((�S"O��S0��G�i�W�֣>�T�"O"9�eʔ{��l�0��M�F5+T"O��A�ߺ&~]C��T]������4�S�I��l�(�8S��!l������ͺ�!��[>�^�3V#PW'X1�� � �!�DD�P��͓1� *4!����[�!�$��!,2�Kʗ�rT	g�Ɵl�!�$ٯK��m��n�����oM�	�!�$"/K��i��[�@�!D�V'�!�dFZ�`��%�Hh�BV2�!򄜗sLd�0��,bf��B�o!���g�ę�� "_4J���-<!�$_�($4y�I�q0����!�D�#%(y�
BG�Z` "�Թm!�䁦A#(�"�Į\0�#��<!�R�!+��"/����ވ.��'9ў�>��6/H�x�D��e�B�w3H�R��*�O�扙p..5X4&�,S2��P�v��B�I�8�,@��%^
F ʢ��:3�B�3�117�M ]�4<��T� C�I�3�X5�+��n(	�6�TC�ɜ��R" 0Tˊ;T��u{(C�It<QVe�GZ�IR��.*��$|��AQ�/`�z�����6�<).O��=���!b&�J�]4)C���c�!s�"O�� 1*��H��գ�c?DS�T��"O�� �_��9Um� ��Ubt"O>)�B��6�^l����4dF, "O���A��)AA m�/,t��+�"O@U�$�ޱ����D�S������"O�Бr���0�IT�G"qzM�5�	f>ə��e�H!˵X*��Qf0D�D#vş6e���� s֬��`"D�0`��G�0e���e|����%�<�	�?���N wtyR&gF�+j��w�6����T�u��ʎ9�u��X�����#ϔN6����ϋ0�����a����8񀠤A)`h9!�(�m�e�0D��(�M,\]�U����.[<�@���"�	Y����''I����
A&,0#t-ȦC�$B�ɭI���ywe��.6��c脂	c�C䉍a�֭Ѥ�� ����+9
�C��O��ْ��-Ez�fĸS��B�I/."�x��g0�E���_���%��D{��DGT�wa�P�V�:&��``$�?��'����w����1⬋�v���8I>A����5_`�����=5�0�!͓S!��� �z1�5C�"�5H��]�!�$�J�"����¹p2l���J¶d�!�� PT�EM-p\��b�C�-�q�@"OTruc�/�:x���4O1���|�P����W�R�!�ߛ:�<�%G�;Oz�B�I�{fh�z��T�d �`��4	�<��D{J?B�J�c��
��Io.��B��&D���Bm�_d�����E
�4�&�.D�P���4��%"��C%�8h��:D�(�'ި����g�ޅ*��h!VA>D�슳�W\ 
M�p� ~�x|+��;�O��m	~e�#��$v��* 	��
T:��ȓ>�b��Vn�����=�}�ȓX��$����5x�6�PѯȪ{�����l~�׍\�*)���T��m��&�/�yB(J�xz�h+�Lj$L8q"�y��hb�$�Rn�P%���a���y��@�S��E�d��M�d����\"��?��'^N-�Q��%�F�A�	=�\��'�x�2�M�$=��y�Cg�(N꬝��'�ы���3Ȯ����
�E�����'�J%�u���vY�N�JK�5r�'� z���D�d�@�E��5��'�9�uC&QB�"�g2&�db�'r�p�k�/)æ�+��  �~%���*�	ӟ(�	�!�����(?�~����?uri�ȓ0`��A(8��u�Q ����ȓ&öP�D���24�'�"B��؇�	�<	�J	�����p�M�u�<��VNMLpp�!�1f�,���K�o�<�o\��V����n�K	o�<�a�_#f<&�:b��-	3BY�Q�p�<i���-%�X�h��*ܑ�D�We�<1a"�3*���;�|�aU)c�<a'�}����v%��ssR`��lΓHEX�HL�.LI��EL~ P�IP(<�g�Q�U�N��L/i~� � d8D��PB��W���(g�)v�P��u�5D��Y��_y9(���-t��B�e(�O|�"����eU�t\ҥ��NO#wf�˓��'�ў�sdJǯ;3�&�4h�d\�dPH�<����v&�P��8	Q>��b$VJx���'ptѩ&��g;�8"�(Y��6]�	�'Ƞ��'I���,cG6��qO]H�<���
T���k� �7�jbq�Ah<!� ͔g�>����}�)�tm���x�����iÄ��y���
�ўD�	w�O��� ��®`b‖+szƬ
�'�p����/JO��F��r6b	��'C�܀�I��L~�P�u��g����
�'��b�O�XG:9Y&ɟa�|
�'��2Gʖ�GH蜠⇀*m�<Y{�'[�E���S�
p��QJZ3e��Y+�'Bݩ�E��
�h���̞-
(�'q� ҷ�:|[ Y3p�S�TS
�'&^h���O	8~pu�F�L\4^q
�'�`TX�g� <�L����YclL
�'-��	`E%n(� eV�Z�x��	�'����]9Dt��g&Z�&+~��
�'�.�	S*S��5 @�˔0��	�' ҹ��d #�`��'<�L4@�'Ū}�P�ä��i��*�34�T���'��C�(m�.�9t�A�/(��p�'���+Dh�;%�bx��ŭ||
���'e��ƈ!x��5����hh���'�X�1����� �b�c�F����� ��9b�\;
�����*Y�&��%"O��AW��_��I�aJ-d���7"O�����xin��6�ˋ*oV�Ѥ"O� ���Kn��t�21;�p"OL�:B헭T�� e�dG
�I�"O&|����R����4$Ƽ>�b"O���-��J�UR��G#�I�"O���oG;U9Dx����K����!"O~e+ �(B(�=�B�_$gDB�r�"O����Ў:����ąC�{B<�"Ǫ�Teئd�����#D�P�Y�"O����V�'�tY�d�
ƈ[F"Oy��b0%�m�e�"=��%��"O|��aH���t��ȄNZ��["O�L0�OOb�T�B��޻!H$�"Ol	�r�GO:����	��$=��ڳ"O����	D'1jy�'"6���s"O�8�朂)&�� �
fr$!0�"Ox��@[y��ա����6˪�a"O�D�#��,u�z)CW阠p�4�ӡ"O(uh�Q%�&�q$��)!{LU@ �'����%�� ����F?� HZR�.D��;�&3# mz�OʓJ\���
?D����c�z`0�[ �`7��;�&=D�r�0t�⹡hRX���0D9D�8�G��+Jb��i�g��uh��2D�$�&��73����MޔP�a0D��ARe�&[����$L��X$�./<O#<���f���s�%C n���" ��X�<YF�+g�Y���سSnPt���X�<��ˇh@R�$bް"�\��S�<�W��&#��H�k̓E��`�G�^y�<��ƅ	�(���� i,����y�<Y�oA/�J���U�#ZX�1'c�w�<�֥)/�P�;��&���� Mt�<q֤�$b�QG�>p���ɔH�<ih��?��(�E�^��J�C�<QR���6�ȅFO>cZUQ��Mf�	t���O��З�0,I�;R�F,&z� ��'����f$�n���j��
z
�'����E�Bl�>�Ȑ#.1����	�'�6|ye�7dt
P"ޑ+���A	�'�@a�4�/���C-)�}��'Ϟ�����$�DM� �2&r��0�'�!ԅN�N=sqe�m�>`Q�'���&�ZlH��E�0yZn�P
�'�.��C�ˆ���9���	u��@�'Ԝp��
l���CAcS�斐{
�'�bĳ�i���x�1��U�訙"
�'5�ui���j疉����hwx�0	�'-�mV
I V���kSN�R�����'��D+$���jP��SB�F���	�'��<� �68�ICh�-��:�'/����V��\6�T�.?(��"O�,;+�1mb�s�A&X�$�s7"O�� ��$}N��G�mn E�q"O�[0�D��8"�F02�t��b"O��9��_�e��9�d$��X�$ݙ1"ONi��N@5L����E] 	:���"O0qis���+�
��ópж���"O
I#g��8/}�� ��t��*�"O��Y���&@v�[�#_�z,��"O�����'L.�THp���Ј�e"O<�"'�L�p��a�4��:�ΑR�"O� �\0@d�)@CJD#7��=H�@Ăf"O@�3�����l���B;�30"O��q���8���+���X*d�
�"Oz��!��Y�Z����[�\|�2"O�!1�(A�iH���W��=��X{�"O@L�a��:O�*���G���.!�"ODAs�fJ�R��7��)��}�V"O�����I�ho��1�o���h�"OH�C"DӘ2y�!1@v�ȅY5"O
h8�
&�$ě�KΏ�>��"O�p�R !}��BK�*�@<�f"O�8�t���Kĭ�S@˓p|�P��"O�0Ó)�%����a.��#o "O�He��h���3EM�{ZbL"O649�c��3#���� sI�m9�"O�d��`�'!�ʨ�f���_1x4��"OV$��lF6fH�|h�")!�"O�q�����?d�hYdW4� "O,%�v��*z�zlrCc�,ZƜ�"O��Y dT�M���b�D��"Ox��*�cJJ��䀅)�x�p�*O8���ʗ��ȗ�*o�i
�'�T�-�l�t$j��?kz:
�'�N<CՉT`�L�"'̍8a9�y�,{�>����٨Z��qr��D��y�lc�t{b\�H�r�È��yR탵t¤9�@Qqa��pA�y2E!��`����iƎls@�̚�yb��7r۰� ��$[[nl) �u��ȓRO���P$W�n`�%�#͒�;7Z4��f�F��L ~5p��oO 
D�4�ȓN:v�R�k�3ʺ�325}$��ȓOO�yh0�� ��ō. VRp�ȓr+^8Q"�n,�A�[1	K.-��t�R��ங����TrU��0s�໡bP�����n�t
*i�ȓP�<`ꂧ c��C ErM�4�ȓ	M:i���ɚ�!F��,� ��ȓ>P���An��2����uʐ?PF����4�+w��������P n��A�ȓb�d����J��j�)���0��=��Tc���F�8XΖ0�5D�*#�d@��� ��%��0#�NY)����6�����J���� �H�*X�8��B���ՇȓE���
7aзl}`��v!,Їȓ@D���W�Vi�<�EΒ
�D��3�M�Uȟ7Jxs�(F�	����.�������a�v�CэJ;������D~Çt�ةR�dJ>�P�z�)T�yRϋo\�c�A�?�=�V�I�y�l�8�(U�f�P�#���V�6�y���)f+�(�5D�/#���2�A��y�-��(�H\�smO��L̳�K��y2 00��ˋ�u.8�š�)�y�c�0V�@t��U���ˁ��y�"Z!W{PX�0O�F�Q"H���y�	ϣd��g�O����Q�����y2�ʔ_�,�[��ݥe��RP�E��y2�ǰZ>d9�̴N�Z9`Eϣ�y⍇��"�i��ڞL>>� "lD�yBb�{G���)�?-	Z�yA ���yK֒\��@Gń�^d[QhD��y�h˻L�"����*=Q�0�N��y�� $Q��M/�.�I�����y
� ���� ��$�ŋ��2�����"O�9��@Q<��5S��J�i��"Ol�z���,���Ђ�Z�4��3 "OXC�^�]���n��І���"O����%�.�WÁ/�X$���'��$q�G�[t&4�v�	Sn���A=D��P�i	�84�r1#� G�L���<D��AGh�)��Py�/A�vR��z@/D��!�+OE��r��12�R�rm1D����'ӨuK�L@d���X���h0D� �p�^j��!�]�{.�e/.D�T�A'ǥ]�|!�%��j�7�-D�p�f  ����J'��0�6D��	�IY���4��f��{��tK�!5D��Ť0unf抩O)�Y1�6D����̶[�d��U�V��|m�b�3D�D����v Kq�_9'�N����/D��*�f1p��ҏ-,n��QG/D�pKV���G������L�:)L,�֮+D�x�d,�`<��JU��'�p�$�,D�\�T���:���@��1/�A��(D�4��!�9/PaK�!j�mp �'D���c�4Q��M�eC�l� �$D����<G픥�c�M�"����6D��ҕǇ\0�x#�o�CYxu8�,3D��c��ńP@�4"׬L!&�Hu�$�.D� K��.m�~�CU�2ve媶O D�� u _�=lh���ʋ���D�=D����N�|3%���F���8��<D�� g	H�?y�q�� �bi�%��5D�L�B��>u�1O��,b5�#M2D���k�"TٮD����@eD�@֏#D�)E垕6�=IV��c��*6� D���u�ފmA@ #��^��h�"h:D�T�`��F�Mk�j���|�f�=D��'&ߐyQ
��U��$Ttܔ <D���oC<T��D��K�;P�� ��8D�(�	$BI�D�D,�s�ܠ�a8D�<�Ǭ�_l���ɘ1x��4D��#��,;**L`A*%bP��2D����T�,���r��Go*��0D�l�P���u.��xԥ�}��Q���9D��$�Q.,X@c�!$���
u+;D� ���vA*��匀U	�����4D��)�bT;��ف��Ы	,��8��0D��ȕk �b�J`�Ϧ��i"�*D���!MΘY����J��u��2��5D�\�7���F��ŋ��2��\�uN(D�D��_"=&,tj0J�?e��|���$�O(�y^��+���<\�`���,߄V����{��sw�ӹ�� �����ȓ�b�I" �Z3^|�� 4����nJNP�V!�qC����%��,������x��ϡ.T�3�|C<t�ȓ#�P6G_0�hw���z�Ή�ȓWT$9�7 �`��������X�����Pyb?O2�iE�N�eܤ`���H�q����|��)�S��B��c��&(`�!�
�vRB��,z�JT�H�	��́1�,|.B�P~�0��m��a��Y`0AA�8�B��)Vry��R�=`XYa_�GD������x�Оf*������l�!"O�@x��˼h=��j"��k���Cs�'R��'��	mD����	���;��8(��hG{J?� �ԩ�%ӌZ{��kѵ�X]�"OxЊ��o�4���+zʾ���"O���FZ:}@��s!�36��(��"O(�q!�!L�LA�A��h�PI��"OR�*���V�� 2!�S��`c�"OъF��D�$�#�4t�9K�"O.`I�']%4x����|� L��'=0����C��L�i�
R�M��'��%��*�$�0ه��L���:�'��ѭL3%r`p'�ц7���
�'�x`b�Ù�Hl$@w(�~�i�'+b�P£En����B4q�x��	�'�FM�g�ɝh� i��ƕ7��a�"O�űAm���2ck@�s�$�r"O��J[�����	c�|I��z?�'�ў��<�k)%D����.Yb$�I�c]J�<��dLn���S�"3B
e	qÓ|�<q�K�1>H��7#�/����p%�s�<�t)��E��A��݃+��h	D�s�<�?;��(��P����D�Xx�Dx�CW=}���r&��/_a \�0�1��;�S�O�0�窝�	�>9Eo �~۔���'� �C��K0��)≂�(DP	�'��Y�E��,��	@�ϕ;��Q(	�'F2ŀ��@O�~a{�*�)7'����'��D:�a��jIp�,^�.y*T`�'�8={Ae� �������$��� ��O�P��J6$bųcj��Hc򜑤"Ođ�J#Y?f]��"I
^�M���$�O^�}�WV�D��� uwpQ���l�0��B,t�2�
a����ҍ\�H�ȓ��A�������@	G.,u�ȓo� 4;���.��e ʜsg!��
��薉a�t�7%Į1VĆ�H̓G�p8[�8]+���(۩F� E&��E{r�dГ*S<� Z)^ũ!�	c�!�S< V��QD]� �J � s!��Z��ء�H뤅���hm!򄀝du<��6<�V��&�>kd!��>k�h����;<�i��\�kc!�$L�4bLO��
�\|W�1y!�$�hL����h�#Y�Е�bހI���`��ğ���O�b�� -b*��R.��9A"O��頫�NŦ�:�*ȋ7ల�"O�����N-M��4`� ~H���"Of�Q�J�.Ը���.���,�"O�X�Ul�$�`�F�ߡ^��[�"Od���Li&v��LV�Ss��!"O�l���X�o�Q�ËWYd�H "O�{����I��@�oCbD{U"O�y$i،mE�$�ֆM+���	�'6�����!~�����Z��r3�'��<[����~*�+(�/yr0��'v�Ȃ�M4w@�8���s�F�s�'�
�Ai��$����!���)��aS2Y���	6����/TA���Sc��z��B�I*�^���{��U$Y�����O\��B͖lN�C��׶)J9R��&D��ID&$4HL\C7�2{�@�h#D�l�#�A�W:	��.0|HE
f#D��_�B|�H�ĖAmbQ��!D��HED�H��̒F��<.���C?D����gʩtXf hTʏ/>>2E�S��<1����(��
�i�2ҴeQt�3/���3"O� �(f�ۃ��YK�@��q�"O�a �E�=�B���_>0lb�[�"O���@�M��J��A�ȡQ�X�[�"O4@��a��Vg����\#!�|�s"O.ͻ�ꄵp�h!�+��#�% 6"O�<�7(�
>Cah7��%)S����^�|E{��;f�cf�z�z$^�!��
+��!�`��nf����F5�!�d�,1^�gi޺8o�1j4O^;Y�!�Ę2��,c�J�M�
�P�H�6�!�D�(T�h�䊄&�<4��'[�@�!�䍇m��P���{�XypG� ��'ў�>�˵�c����
�J���
���O�=E�A��аi�@��UX����!�D�:��`��(r���
�4.B!�d�G�Zq��䂈;/����	�!2!��vj�(v�ѪHX0s����.!�d�/.�U��ȉ-4l���j	�F?!��


K���լ�8�$�Jg���==!�$���y	c!�$	�l=c&���U!�ę/ٺ�1�� �R� 2�ۄO<!��[�BUI�M�g��X� N�!�$[�7����荼YUv[�$i�!��Ѯp��{�O��(��'MP�>!!���k
�Y� �߆ӈI�N.!�V7���Iঘ�h�\1�kRv!��q֔d��L\�hľ��%*�-H!�Dn����QAϜ:�|	�G�r�!�Jh�F�R� �<�@P���;,!�ΝI`��92J�����	Tϙ+l�!��=#|�k��ɑ*���	3Y�!�䆺"cz09P��-!��PU��*8!�䈷2��cԅ�z�5��,i*�'a|�c�n}�(�)��]��r�mײ�y2�X9@�8\�cW'׎�X���yb�Z=�Y#�
�ڤ��Q�Ѥ�yrG�pX��v�K�V�ٹ!�T�yR �,�d�*௓$QY�� �#��y�%@11�TX�ToV'X���8`���yr�c�x�#r�!�J�b'���D+�O��6mךhO\���e/`�	v^�p�?	�������uD�DDf���՗6N���"OF� SDE
K�J�re�E5��"V"O�@��S�	�(�H�d��E(��"O��6��7<> ]��I��-h��"OT-
�Z5dD �񩒇7�@A�V"O��q(%{7 Ԩ�Yh�.���"O�5�b/��W�Q
�	ވ�H����|��|��'>�q#l풉Aì�>6�=A.)D�$k$#���ƌ4����@�#D����/��|���1$×>�fX��`7D� c�Me\1�qg: ^L;�:D�<��V���{��P�B�3D�P���?(��KZ�A4�Ԩ�j$D��#�f��t���ْ��4(h�*'@.������I/ Ǡ�����	v�
�'��u��웚-%f����1�25#�'
ʄ	��#�*��枭l�$�2�'{t����g�\�Cf�zS��#$"OvЂ3��#F��(��J�(�H�3"Ol˒��)[HY��
"t�(A(D"O�a��.Խih��0�ށ��U"O iSe" %�h�V���4$�%"O%K�n��\�n�3��W�+���!"O� t��SƽS���:6�>c����"O��X@L�G����M�[��a�"O��P���,H� �V�NHYG"OR|y�Ҏhx�� 7�K�Rz�I"OЄ�S����pq�
�
���1����� E����CA���`R5d �����y���}R�@�c�.|��X�9�yrNѥ4h�ʑ<V��1�ב�y�H��8��!�
5+�d	&+Ҧ�y�MQ5i�D�it��	}N�H`�C��yD�!Fm�|���m�>���e���y&�e�x(���k���c����<���_�K��z��L8!�8t�	Ø"U!�A�#�̹�O�Fb4R�1O!�$��ѓ�Z�H6�]0�|C!�ԄeP�%p�b߃9���[t+�>!�V�J_���WǑ%ߎ��D��7!��ѐDr��O�U�Xx��(�6!�D�{dtD���&�d Q��ՓJ,!�dC����㊂[thb��!���ioܭ{1&S>u>��"��< !�ę�Bm���^�5y��Cm!򄑊�(���� �Er �S�_U!�^
 O�}���ʪ{[�h����DT!�D�#%�ͺG�nekP���!��#A�@�V�UÒ�ӊQ�ў����/l5����ͫ8�\p�̞�Z��B�ɱ���VB<v�D����	�C�	���)YŤ�������'!1�B�	�o��p5"��@bT�!aiۨ��B�	�1~��@$�W�II h ��׬eZ�C�Ʉ|[��A�"_8����BYպB�;��z� �}��y�`��3)�B�	: t�hk�k��d�$�ՅKcZB�I�Fh9�PF�
}�<I�tj�y�NB�	�$ a ��@/*m %	��PC)BB�ɽR�t��4'{]-��$�o�$B��#b�, є"�
vX�!���VR�C��zK�UZ4�8��|ieE&w_�C��:2�,�#�>e�xHcMļB��*}�H�x���-�ՙ1-V��C�ɕx`���5�Z�܀s��.g��C�I������M)S(��B�K�z�C��1<�.H�fJ�o��y!�J�.j�B䉙71�������r=�զS!��B�ɯl\���eBI�FиTbR���B��
�8P��V5u���a��',;HC䉶=�*`;U���?"��p��>RW�B�	�)q�(wJVY��S�;��B�	�jE�X#�A����hPa�R2&jPB�ɼz`�MH�$�,ߚe*�"�2&fB�ɐ^�f5)�oƃX�X	�,��M��C䉲t�p�U 
26�n�2@J�{��Oj����" �M8%K�d���	��G�ўć�S�>��p���!��8�#�	`4�C䉚.�����. ��Ȧ)B�o��B�58�m�#�j���8QlR'	�B�IG�.):,�0A7Ψ�e�2|a�B�	?z�p}���e� ��M
�FC䉔��@9@�
	���b�D >'3:�d:��0LO
�*�d-�I)saP�C�D���*O�A�v���)P*���@Y4U�Z���'t�V\�[�z���e^�<H��'��D��� �\�4YR��� �U
 H�Q9�UA�^~��R4"O�����"^8�(D�Ӧ��R�"O������"#�z��:A�.I8"�'.��'��Eh$�N?G�6y���f�tU�	�',^�	A�$x:QR��+bFM��'��ݱ�!Y.m7xus6b�+R�ְ��'@Tt�Vt^�����PP���'8K� ��k��p� ȴ
����'[L��ホR�f��ĭs5��'j�y��TU��z$eA�jm���'���G�L|RX��s�E9��0��'?�d
��_X{��cG�p�B��	�'4�!q� �40 h����~li�	�'�,`02��2s0ѹ����P	�	�'j�L���`�\d@�m�
�j	�'���-8;Ѡ� �Nǹw����	�'�P��� ��, �G���p�'%��0c�ա`���aC����	�'����!��As�ݩq�������'ÌI�@L��r:��*HX�'���Q��/;�R���鑦"{,��'�.���l�:=�Rq�ܢ ����'$T�2Un�UɆ����T �>]��'kXAy��
LD��I�4�x�'l��i�8C��]�ToV��9�
�'��pPV�V,�������"A4���'�PԨ�� �iE`媳ᛈzx���'�� ��MK�j�����*�.K�d;	�' H+��[�>�i���b�t���'E����]��\*�c�"qX����'�JiAe�f�$q7LZ�ev����'Ȗt���Q�X�f(�T�Z���H�'���ʕB�7M�>H0�N�f���
�'$��@[�{(z��ۣ0w��c�'C�� �J-i����L܌R\ƙ8�'�0ɘP�:A�zT!AEB�M5��'S� ���%_�:0�p�#>u*��'��y�:l]4�G`C,H�@��'�"�:�S�~uBD����<�4��
�'J�z�E�oa����6F ���'0xxA����*�dlՄ?-�8u��'�,	@C��=�qow�:pv�<�� �1򘝐�
E�kH��k�@�M�<�c��e%��	�k�a�ԡ�ǥ�I�<�fg��N	�u��;bz���Ǎ�m�<�E$ňf������L;Yz��jRj�<yg��'<��Y��X8�r�Bf,g�<��I�R�2�3d�:Q��Ӊ�n�< �\-\P��b��9B��A��$�y�"�81;*����q��ؑ��e�<)��ɚ���"/͠,f�+�a	B�<��%ɱw/������%C@��Bh�z�<A��O���B�/ٕU�� !P��N�<a#�ͭwN�bg�Ԑ)��`"$�N�<q���(-s l6`�
>�(��ĚD�<��Ι9��qAU�VRZF�C�<!��?clNh�4KH�:�m���YY�<�6x}�I0�\K@�@U�<���^�j�;s.Đ6��Yr2��j�<�U*1º}��e�I�=R���a�<��R=ՂS���"B�r�	��H_�<�� ��W� ����	�fVD�1��]�<��E��4I��$B������[�<��V�N4����ٗQ��A�GC�[�<� 1�kö8:��hG/W��ӆ"OZ8�Vf��8oF�����B��Qg"O��ض��|�.E��<U��+�"O-���	��D�B�
S>E �"O�,�F)�)f��4a̛FQ̼z�"O>Y��)����q%�Q0z5�!'"O4��	�^���(�C�4j�Kv"O~U'�U�\8,�0�b�8%�Lz"Oj٪��ZҨ�a�!�l=�W"O������m�C��*���"O8��7K�5pգ\<t ��@��y��|�N\�@Q�i�|q����y��	�"(d=���Q�f������y�ψ(�H�S�E�W���F��y�#[1)LY�@i<M�\H�u���y��%����C(D�pU혿�y������ ��h:|
�� :�y�o�0i5(�"DG�cf �Dlŷ�y�+�(r�8\���2V_"��SM
�y�*�,�Ъ3Y��M��-�y�
	F@����ּNhp҃Ģ�y2�Q
l<^IiF���D2*�3F�y��ˊMlP��t�D\� J���y�
����x�f����S���yF !
���N�b��b"�ߋ�y�(ɑ.ݦq�b�ۦ�1B�O�y�
̰>
���1hX�\S�#�ybj	��k$,�Y��3�y�F(q(���=�J$P�LN6�y�#I�+W  �fЮ<4B�����y�KM 2B��S�a�Hؗ���y"IL
`0�q# �`:��i�g��y"$<Zu�E���X���Wƅ��y�<P�LA;O@	W��Ű"���yLd�u�!I�fnb�ڡ�I��y�N�&�n�)�h���j���y�g0{�)���4����T�1�y�$[��������x֨%�c�Ũ�y��&����Ώ�x��Х�(�y��%ڨ�ʖ�Ҟk&�� ����yrƏ�(�(TT+��^=�Y���$�yFʌ'm�%�7̩l���`���y"n�:ê�C����b�\�a�'�yb�T�c�\�E��F���mП�ybM��	�����
]�y
�eV5�y"�W[�,`bD�L� ����1/C��yb�ƢF.@�����p����AŃ�y"�L�0U�6�ʱr�^��p�[�y���;�*���NI�j�PH�o���y¬�����e+<�S�j���y҄��k9���EԞrk�%"$P��y�σ�r �6.������1kԣ�yR�%��	�U��@���y"B��H!F�W�<�0���y�,b���S:�(��@�ۆ�y2M��)D�åR7/F�!�LN�y-��m�h�p� ��xD#q�M�y�	Wu\�b�)x���@,�y�I�xR����m>�=�Q���y�#I3z���kO'a���
O��yB�У,O4}Å��T��䒓i�*�y2�_-X��k�Rs$�Ht��y�&��s��h�d�=ISvt�ù�y���<2���q׾H��X�)ʺ�y
� �Ds�3Z�fM�Dh[Y*���"O|�8��/�� �FfK_���ɦ"Ov�x�G� Q5<��pe�0��6*1D���!D8�������� ��.D�!�B�$&Ƥ��eJ*N��|#7�7D��A!�J�<j��
$����`�g*OXH��<h�mt�E�z󚙹�"OdՒ# �b�,<1�3��d{�"O�g�	%T�0���Ė��@"O�x����6�$
�焰S��y`P"O¬���	^���֨;M�
��"O�ɳWB�9�~��;C֖��v"O� ��.����#'a�@_��2�"O�#E���j2b���@��*T�PG"O`͓�h�D|lKa���N�y�"O�h�"����=)M��<��Q��"O�l��ٽ%d�{KE�k��:�y�K;X�1�U�G�����y�U�G0��=MlL�5�;�y I�=Z��f�A(.��i���F��y�HP�zA!$;�uB���yRX$�ԡ:$H)�d��Ñ�y�	?��p%�q��a���y"��-,�h���"�>o��y��a�yb�ݗ���˔f�.14	x!Һ�yR�S$6���0୍.Z:U��ȁ�y�ÿL���`�E+i^�k��G��y�#�)Pb>����צ��*�+�y�f�xk���D�*:<Ÿ�)��y2���	=��IuLԧivz��2-���y�L_�
�TEe&0�f��A�O��y�oJY���hW�"(���@ ��y���@�f�Y�h뀊D
�y�c޸�Jpa�(w\���� ��y���Bx���mg�#{PBlC�'��E8eB���y���N�n2��
�'(��4g�>������{���9�'�2\ q
Ӈ}��U�5J��yqT�x�'=ў"~JB���K��`$�\'X��#�"�l�<��@9<Ƹ1�aID)l!R��5b[���D+�O�-s���A�,�)G��)<��Ğ�<��	/x� A�$�N�o<tk�C]�y����D�<y��O�~��03h����7ޣ�y��˩n�f�	D �y����F��&�Px�(�L�$'�@qZ���^��~եO*�=�zS�	x�!�c@�.�fU�� c8��Ez-�"^R���[ �1XD�Q9�y�H��<8ི�d�#N]�ruA����Β�~Ҝ|ʟ�R�x�b���>��S�V�������n�N�%�w��!cB�t�Q�u���>�G��4K���G�z�<�C��;$7č���V�g�1OOF�?�*�'Y 
���'cj]`n�i�OR(Fz���mZ�%���y4dB�6i:a@���d4���t�D[��`qyF	!~���ԍA�!�=Y�~�,�H�
J�?�P��-Ov�/�i>	�<aC�� a�T=��x��
�q�<	1S�@�r��P�D0q�IX�hFy2-V"57����I���ί�yBLϨ|욦�<��9pTD�y�ǜ�M����I�H���B��N�y2`��~�P��9WOKQ�2��P�!B���c"\�т� 0�j��ȓh��I�/ɜ�Pً3�Y����UB\0��E�ML>	����l����S�? �d{`M��}�h�ȶ�T%^C�,j�"O�)AvJ�2YbB�`�E�����"ODkGl
��>��2" �bm�@P$"O���%N�/Z� �@�^dҭ�"O����@�	J@ޑ@UȒ��x��)�S�V�D�S&�H"�Pi�Ʋ,ȆC�ɢ=\���%�X,3�ha���yrc�t���-5D����ߠX+���5l�-�2C�>-�8h�E �"���r�H]�._��'vў�?��ۆK��Xk!�ɲ]&���j?D���4dێo4����z��囁�>D��� i�.�T��6��� ���"�)D��`Ɯ�:;�\b�*���m@�E$D�Xh�l�4]�`�p��`��'D�x
PFL�t �1Sc�2���bC�+D���n�^�.ŲpF����")D���@�LD�<z��G��#f4D��3$A3��\"�+@�YI�(Ö&D��ХW�\p�֠�f�����j"D� ����h�\m��a�b���I!,O��<q��O6I��h6�$��t�Q�v�<i����&�f��3�]*oI ����n�'�qO �'d.�4�@Jܹ�d-�6I� �4]��E�>X�AK�Ƥ�EL�G�2�ȓK�a�D�4<�� �CHPێ���iW�,�S��)8�ZQ�C�6]T`�Γ�hO?� �[l�qZ%_/q0����/�O�2� �K����jH] �,�Aᘡ�ȓ%\جS��loN���K������XQ*�-3V�0�S��Aڊ	�ȓ:����2g	�\�F'�c����'�ў"}J�F�-q!�u���x,"$���]e�<ia'F�v�K��0kVM�G�Qk��"�Q�t9�y���@��q�b� �Ѳ��ߒ�x2�'#����Ή
���s�@՚0�f����'M �x'�H$ ֐���@�36 �)�'{�Q�T<^�� 2F��5������6}��)�=�FAj�G͍\Sh1��ʼj_RC�	|��D؇ʉ0f�&O^7�C�I%� a���$�`���Z�h�̣?�D�����!"�ܸ7B�Q�e��(��a�O4��l�(�x-�bB��o�mzvC�N�<�u�&V�1uDP�Gp��{�K�J�<�La���:��,N�>����S_?��g=�S�O4	(2k�%5�9�4�[7y���[�'��9�E�	$�p�FG�8u�M�J<	7�'�����*ݸn���25�G�#(�<�L>��O�#}��O'���t�E3�f��%K��R�'R�\P�l�J���ݖ'5�90�r�'wP�aRnӣK.���l������'��PJ�/���I��ќ	]�$��'����Ux@H	D���,>̹�u�)�S��?��D���L�����3�l�5�T�<�wN��� �^�CnVqhcAڦMne�'�Q��P���	 Y���ԫ;�>���@+D��Z�B>V����Eϝ�d� F�<���<�����[U�|�t�ޗ{̀L��� �Q�!��
=9O�y�e�I�t���ri��o&H6�'�S��yߢD}�1fM�A�F�P$@׌�y2�U�QY�M�@�,eJ��0�y���/o�!�앦Yqx�������0?�.O�!�Aj�Kնy��)R��6�3�"O�U�j�W����(��lܪd"O��P
�lcb4it�����"O� pu���%%T�� HI����O6�=E����Ψ� B��>)$�� �L��yra�=_-���S��#�N�(E:��6����a2[�c��c��;0MۨF_!���Ħ)(ȋ	O��@UA��T�V�x��?D����8Dj�9  дY�<�Ȇ�=D��JS��s����ժ�$K��8�'D�\ڤ˕�C�
�K�O�+�4�� %D�����$Q�@a���
�H��<��%!�X�ΕE��D�
	��;K�+#`&�8�����'Fl���C�puc���];�(զR�'�D]"ef�>O�<���'����i�>H������(��ʆ#3��9��'�$�2A%_��I#��E�0ך���O�U�L>�rg@��u7��^�XT��|�@9�3�&�p?9�O��Z�"��mi�.��@�a0Ƒ��G{���&����r��qCP�+%�4!��;ЖT���R:|��0b"F�z��'\����ɴ8(�(Cŕ.i����'2�=�çHL��'�C���d���m(����aPNL#�c��\�X��ˆ_�\M��e������c��$Z$�Ĩŝ>��M�$�,�O���On�Ӥ ��YA0܉��#ކl0�"O|�Xf�4&���� �$&�	���'�ў�ڐAӼ3�x�kck����L���!D��'�ǲ@���!�@���i� >��2�SܧP�|�T�֨L����&�	�$k�i�ȓX���`���U����mO�9B��oZH̓�0=��̸+�­�4��6���Opx��Gxb"�?8@�*��g�ҵ�݂�y�	�'b,�
�F��W;�,�GB��p>	K<qw�ԖH��\�u	�-3�H�
T%�d�<��������PENS?-u��pO@�<���S��Y��M:�4�e��g,jC�6�l�6��.<���K4E��t���Zz��4A��f[�,s��ҚjH���v��[���;lg��g%��	`B ��cl� �J��x��$2&��8�0 ������H�	���0��b�PCҁ��-<�C�ɥkf�CW��&ø�C���6P�bOf7�,�S�')��= U-�g�mY���2{V��Po��p�m�
^Iҩ[cD2�� �ȓqF�����@Y�n�(-1���ȓH#�|3Մ�sr�D�7��#k�8݇ȓH��B��:�(� �^°��V�kg$�2��p���_j�ՄȓQF���!�m�R@C���nyJ9�ȓ :3Å�k�a0ժR�5C��ȓ7¦�Z��$��=`�Q�2�M��O��b�IR����X�a��?`}Ys��dh�Y�/\�p�ȓR	���cǾuDTKS�_��ȓkkl�2$�-�cV�T�d#z�ȓZ�h`�P�K�4�p�
 H�0��;ֲ�"SFI<��[v)�+�B�Ir�XQ�� ق�A�T&��C�I�������TlH��J�C��!4*��)� =v0�Pge�&�fC��,>�$"�ŕ7MV���"	6l��C�	0%]Ph贀ש:&��d��6s�C�	*;9�]��Ѵu��Q��/ռ �C�Ɉ/��@�Jh`r�q�ޏ?��B��)�"���Α� -�(;1JQ�B�	�XQ�a�!B�P�3@\lg�B��--S�A8��=a��T��ǟ�/�B�)� ��r�R�/%�U��c�R��)pQ"O�h+��L���#��:Ш!��"Oq1�L�PT R�a03�����"Ot��#�P�&��)�B�Y�e|R���"O~���f^�U� �K�j��
IҠ�g"O�(�(�ap�J-TH�!�!"O6� SlٸM)����'�@h���"O�#hS0Qj\�����Z���U"O�(cA��S5���%j�֮}p��b#��JG>x�Z���"6a"�	:0*��j]�f�>r ��K�B䉔Arė4tN�(�j��1�� ��"O,�����J�	nz�P��"O>��p*�	}�Zx�v��(9u��"O
�QcC�'45A��(���2"O�u@ꔜ2�T�$�]�f}d��B"O�Eb�`�"Uv
�m�1ʤ��"O����@ Gޕ@"���3ʸi87"ON�[t�[��4Z��Vb��ѓ"O\���a�wBx���	���"O� �C��E$�b"�D A�<���"Or݊�)��}?n5R��
�0�V�c"O<�Y%�q����-i��!p�"O̩�� QRn��eZ+(���r�"O���qJG�j�tQ�1�)�JX�"O�u��.СK�KҠ+z*A D"Ob`y��J5Ө�K��;���b�"Ob���\3�X):q �.0p4�)�"OV�9��(yVѓ���<s�$h�"O��p'��������ʇvh���F"O�TR��B�!��� U����"Ox����fM����&L6gc� "O�T��Ę?%��S�Z��x��"O��!o� a�ݠs��5^҆:t"O��*���4�ȥ��W�v�R "O�p�B�� Pgl��-�/i�M[v"On��lת\l��g-�%^��1&"O������W���フ�1�V5"OT4�����;A��h��ܦ@��Yʡ"Oʰ�f,�tT�J��B%,��`"Ob����נ{ˈ��F�_�i����""O�4�Ȟ9�^��@lW31�D�r�"O�0��4?����q���>l�,�c"O.EJ�i�%�B�;��sK0�t"O��Y���-P=i�$H�R4m&"O�}��	�'^�ء�NL��@�"OH��b�X���-�g�� $�S��'�!`ebP6�&J�2������+O�UL<��E���p=��M7S�Zq��J�f�	��Mv�'آi{�mT�W�k�Q����'x���{���'1�hԂ�׋�HC�	A�RSe.E�u�@�y���w�n7��
c�¹P�.����$���@�S��\c�����`�<^���(N�lM��'G�x83!��.x1a�E�A�����'�NH��+��  ^
�Oҁ����'���:�)K"!.8���a����O�0+�k�_�(�v�-m�L���)��T	@���2?��������])���)��h\�� P��hOZB�J$'wđ��O�� �NԊNA*p���P|�8m��l��{��E1�',�v%֏-4]V�E=wĤ��4b۠�qG!(ŮO�M�����:��{�2TS���(8�~AB@"Ofhf�\hx�Q򨐢"���_��h��@� 	���'�q�G�B�V����#���Щ�
 ������� @f�7y�f�h��W��@��;4���@�,2��p,<����d�=7�z#=����% Pp��w�#����>$�o�=mhj��U)H��2C�	" �r�I�Y�bK5����P7́�S�2�!A����)��� �w���?߲��CH�v>4	�`"O�82�����ۣ(��1j�P�_���c��#Z�@��I�n\��ssތY3`5������s��Tx���&��k�nȼ^ r��㧗%�!�֌H`*�XE��K������[�W�!�$�5n�X������?d�"��b
!�D��=G�
5~�`z��uS!��^�b�
�#���K�ب�� �{\!�dߠL�̔�P�H�g�j�ŏ_�t�!��<2;�<@�ߤn���GnL�qH!�D�*�u�A`��e~�u��5f!�� �*��f]#$XpC�?*�!���i��|���M?� ez�

�D����B��(��I�o�Z����w�ޕ�"�-.�$B�	�:֌0�r�ũdf�H6B+E׊�C��*tX�Zv�'"� ����Ά�k��$JDF��
Ǔ�f4v/E�A�.	��k���_9!W��W �X"O)D� �˛o����盋*��1Cd��3R��	,]|����/_�FE~lZ��O:�.�z&`H!�Z�BJ�Rᘕ*�"OP��CcH��$Y�J_�&��	�ş:6�H  ?O�H�M]�#��n" ̛��)�)8|A���Z�B�r��>�(O���iW����,b*T%�Xwa4�5��tӸ�d�� �P��b����7,�6j��c@�-�a{"��=,�Z��vl�H���R(��!s���m��dGn�[wZ��ؼL�0�wEЙG��1v~: ��ӥ.9��r6�r8�ȓε�q�E��l+�4c��иq��:�P�;aAJ�7x�mk����¥��>�x;7����;F㲅xR��F|:uY���y*"��ɗW=P��"�D�f*S�4��c%�F�����*�qa�?:�1H�ɔ�mU��XwgH|8�`os➬��C�\Ʊ@��D�GF�l��O%��o��8ѣ�`���D�EB���/h ���B39e�Xa��� �j9�����8��F��3���!��S��x	���'ĭX3�U-"j��h�C tA���������[PkS�
�B��'J�3NL�sO�����;�h�/^���u�R�U#Ҩ�"O�XB�(E�W�� �G�:n���'�X�!k\�sJ���J,g�xz�ER��!P��z�1~�x#�L�#?�xi��5����O�C4:��`0�M���yLm����f��y��U2/W���� ��)*��A�n��yzH'>1�=ա
�bI��.���4H���a�K?J�ztJúbc>�24
ú:�����d�Lx�k%p�\u�ӀR�<��Ѣ�&J5�U�뉘�LX���:t}�h�c�'�����E�n%N�'�L��j�H�`�(>�����0k,׋,*�{2m�*U�DT���A!�$�+XJ)J@�M�F�)�'kg;9T#��ZD�Px�f�[��*ZD1r0AͯG�1�V�Q��ܷ`AL!;׀��9���'�'^��1tU�9R�X�hP�0R	K({ڲd�%ˎ ����F��������[��b>c���v�O2I(�i�%��X �/�Oz�ZCI��?��Q�cb�7��l3�I6S2vUY#�=@"4P������m#5�'�",r���f#�=+�a��?�d������~Qx�$[�7�@D[*�1x��09�z��a�� ]�착2H���5"O�����ƽk����
80�����"K�
�b���M�<���#H�?,��G��2���w��]�\�G)`x���q"O깸e'��}�{�
�c���)���[u
�(qGιS�X%��R��D�I�0R�x)R�W���P_ i���$Q
��5�0���Mc�OO�aU��p�j[e�PS&�|�<i�CM;H�� ,0�J���}������'ds�"}�$Np䐴�%k���3�Ig�<�U�J���p�r�Z��τ]b��P���|*铈h���H$*h�# "�'h �$�59!�$A��%	��H}$��O�4 <�P��%�5���RПD�A�O�=I��� ���Qe��k�y�CN��%��{�f�6<�j�j�TϦ�QgĽ=�� �flK4c�ܹ��Eܟw�N���jò��27�"iuF�_0��$ƙ���<#�\�fjjA��u�vܡGM1F���q�:����̠9�tH��
Ǎ~ĪC��5}���,M�&�PᗙG��0��ھI�|�+A8Ov�!�Afv�ų�����!�J Z��	�P�Y�.Ġ
"O^Be��T`�o���v��5ԢQ��i�q���8q%�g~O�vL�<��	$A".� c` 2�yb�	:Т�억;�*h�5��QT���m?$�`M��S�? ���5jE�����Vg��`9�%��':��!@���iL��I�j^�m�@��\q�b�B����C�I	�a�Ci�"I�$���ŋK�c��`���E&0"ڠ�ٗp�BD��@��H�l��va�g�<Q�� �`�R��1��� ���.E`�<A�U'u�j����_VD	c�OK�'�Х��S�sfzQE�?��*��J��\�eH�In�,h�!D�����%rF�h��h��uyǩ�>��U�Hk��:L�j����9�V�[p"CA�
��́b�<��h�O�hl�2D��B��Sf܆x����'�D0�pʔ?>`�q���O�u"QJE�b��(��cٻ h=#��'̀ipw��+r߶q�#8���hV��`�m�-z(���'N������H�ãg�{�����J=I��Qo=:v���go�~�"�9Y���sf�M,0h��Ed�<�+��\��񱢆��ࠁ�gMg?�%m3�L�8���=m�6mˍ��[ 2Ѽ�9�+%X ��j0q+!�dӵc1022�ؒhu��q篏##�.mkf#�#"�%�&Gq��$b�ߟ#=A�-�4|�\Tˠ�J�:ZR�;�t����b��Z���'�]�F��E�A>�q(GG�X2�a�u/E�.D\D�>R���f�R��$�ӂ�R(W<f�?�*G-{�$y�-$E%�QX��$R�z������ �&����8"��܇ȓdw�)�a�5BA2�y��۴Ha��j�M�fAD�ӛeo�Y�DƜ,�H�`�#9��ҩK��H�%
�*P�,B��!}����@/�
]�*n���B!|��ை	[׺����ъ.�.�	?�h�uxf`��J�#Q����-|Oʅ��L�1��T��4fr1����o����P�*��8��e�~�[6h
)
�`ȡ�3N�\��?q���~�$�p�,0�'%��rрL�=i�E,���ȓ{Y�|��ȏ�`lF<��ʚ4dL��ENI��(�>����O�j���%��K�D�:+Pۇ"Oz�!�Ύ#7eL�u��YL`��'��,B#��Z�L��I6A����1�N�:�x�I���.l���ןWXȈaF7�MK��T,r\�S���*d_"�'�B�<񕀜RN8��HV�Nn>�b�v�xD�&���<��"}�Ë X���n� <��|��Qv�<Y�C�2 h$��d�c#�q�]79�����ML铵h��D�@&��RiNLVD9 ��T3#!�$�%�v��5�ɣEB�າ�
K*��׻[o�
T��n؞#tl�6v��{4OI;R�B���B#|O��un�	J 83�47��������O��xA	�Vy��ȓL�PقV�
xz�-¶�YIN��?Ai	<�Z��%�8ҧ�l�R#&��E��&	v锱�ȓAHH��"C�ЂpKr���D0O5�):L>E��'G�U�g��Rb�|QƞM�8�k�'v\HY���CͶq1c�Bàd��'��z���Y�L;r�ļ�xt���ވB|���6D����d
'���pJ9&Z�#��(D��D-U��.�cS�ʴ �\i�2�)D�Lၡ�"T&�3�g&N::��$`;D��ԯR
@#8���������B��;D��p���\��t��*�&�`��v�2D������)]�Q�� à�j\�A3D����&��8��o�-~�&� ��7D�d��d�-��]r��t����4D�|1�#�YJ��&��/2����6D���C�H�,��Q�NA5F�����&D�0Si�М��" ]�/���@A�&D� �Z�'�Q��ٮUԌc�g8D�8����#1�NH�cT-e�8��#D�$�	<ŪT@f��X�+� D����
_f�@���pˆ��w!D����a�1	��p�� N4����3D�!���&%�ȧaM���d�+D��I'�^t���!��1M��l)��:D�� ��p� 
W��S��';�m@�"O4�ڵI	��p�[�e��˅"O*�s��� �n�r�V.�$\;T"OL\jCĎPb��`)��-s"O$�d�Qf)(�҂[6���"O�ҁcɗg�����@�<��pj�"O~���Ea戋�ɕh`�R�"O�`�7
��(|2�X��w���"OJ`��,D8kS�L��Z��|p�"O�U��a�	R�1*���%n^N<8�"O�Iw�Og݄�QХ�u��4yg"O�y�LR�~\�j��p��C�"O�u��$��>�,<��d�7���11"O��3��$ݹe�/��À"O��ȁ��0�!A���xx���"O2ܩ�l�@����d�]yJ��u"O���Dɝ4v�����$��H{b��a"OB�b1b^6�j,�wb�,E��e*�"O�M�wk̻r�\,;p�B�g�F(�W"O^��f�ü2ha���i}���"O��iV�+Z_J�;�
�md�x�b"O�d 傎?4� �2#2B���"O��6j��~H"@�dh�n$�#"OXǎ�i t(��Θ�N��}r�"O�)�o�::h�z��;#��,��"O��"so�X��,��U�z$�"O��գ��j\R�'N��:�"O҉�C��3�4�� �#j�p\��"Oܥ���͙�%�Ld�t���])�y����a4��6S�,$�Sh@��yi?C�𹳲�T:c<��T�ƕ�y��V�fU�⭞�2AB� ��Z��yr��(��)*9^��6e�7�yrI�!
v)� �-x�t)�녙�y�� 	��:I
�j�=���ں�y҇]�-KSc�붸�0Q��0�y��iX�yT�]�f�z%��CS�Py�#� #���/Z-�]8��_M�<�b&ڧ�� �"�D�6:��ICO�<с��P�\ܐ��Y4e���4@Ml�<Ɂ�E�R�ȼ�榍�K�l$��n�<�rc:^v�;�'	O$<�F�P�<)�غ����K� u@���%�f�<i��]�3�$,� W�P�2�*Q#�c�<%b��s����4i�6`nHݘ�P\�<��MC�p1���N7 ��H��N�u�<QC�g �8�'hF,k��u��$�O�<i��ñp�搻� @(#�q�QJ�<5L��RHvĲ�/K)f
��af�F�<)P`�]�)I�g̩2��T:KJ���eŁ�F<@e�
Ъ8r�
�1x�e��#D����e��A�����ܜ}!3�?�~��a������DljGjl��k�ڜ\x�: "O&Dx%��6Th����<~eK�i�@e1�f�Z����O?7��JтR��U��<�R_�v�!�M�C��i�"NC5~�p9��ֺr��	s��3%kI(M��y�M\͸񐔌E�JΘ`B�	�7�>��Ɠi���Ы��$Z�}6@Z�a���2U�_-U�>B㉩u�Q:�C�-86e`1L�c�
#=�(T�<�0��q�6��xa@�H�ኬv*ő���!-��B�	�I
",C���1R�!�n��v�6fi0ep��+��)����.�.ޤ}���S�I���A".D�̓�l��&�A� ǒ�,��@Q�-�>���B?��L�7D*<O��qC x:ʰBd%No���u�'�
Sk�?E?d� ��H��]���ǌ*���3.?4��Ke�/�9�WL�B'���!ғA�Ғ�����?�I�H�$*�8�!挙�����+D�ԓV�C�ki�@p��аQL5�E�k�Hq �M�H|N�"~n�-d���K��F���3!�%�BB�	�sB<�#V�`�}�g��kǒ�X�������0=yC��r̪̉ ��#P�6 2%�H����vFDX@�Xf��)E���c:�c�ՑN=!򤈌?BP"�0C�> ���
�U!�d�3��(�E�/�6�p��{�B�ɊMW~6��5(���F��C�	�A��qq��R$���@�%~C�ɏ5���%!V�x����O�+ԬB�"*)����BѲ,�2��,V_"�B�ɚYB�t�!�b��I'�ȩQjB�	=w���:W�!��[4AI��B�I�� YP�bҬv��U�6� R�B��%)��T�s�O�Vh��g"�2_P�C�Io ��` ��4G44����:��C䉺gO�(����p���)d9
C��P�j=���{���H�M��B�	*pz����㜪`���3"	�%��B�ɐx��D@*S�*��ɋS��9l�B�
���ф� Y���뇫_(0C�	�'�p}���'a�0���<	����&#~�΍�Gg�EYAd�H�P%���@u�<�#Ӷm�" @�K�1Zn��vm�>|2:y�f�����S��y�#׀=V5��JV��t�#.�(�y�$	��t�EB�H�2�K%�?�-��B Td�4lO�[���9�2(&�^�F�d����'p�]*t
�?)��o�[��rg�Ŏ{�:������.�C�I�5Ȕ�9�ٻ$� �eN�3-�����D�zg�5�S��;��q2�]�cv �U`�N�vB��$�,�IQIQ�v�b�g�:8j�X�qO���yO�E��'��A1˄�2AcH1�l�h�'�
-2�B���x��,e�H����!v$L���<���T/<rb���B83��/<t�{B�27�Ղ#t�2K$�[:�8j���
V�,����,D�L�����p$��c����y�-$���#j���6��4��>9�Bhְ{����%��L�6�$D�h�!LK�*�Ψ;F+X�
i�\�F�6ƾ��2��z�)��<A�`�Q��U)ҭ��]�9D�BA�<Q��Ҏ �<\ru�jVD���IIv?�ġ�z�����S?Kr��K�-��qkPE�b�H�Rl!�ğ�W\�p�`�߫|"�bnֵW2!�䄈"�Y#f�����I��|�Q"ϓ'Jn��E%�2�����o��Q#R���{��p�1`�$B�LhB�@��$Fx(SF�<u�P��i�\�`Gأ+��=;QJ�x�C�?z��OH e�j�xQiы}��+�Gס��ZN��E��'GJe��,S�UT!�G) �8�����'���$�[�vh�4;݌�Z�MV�� a)�J7����Bx-� ���v�dd��Ðaj�{"�9v(<I�&�ݦ���J�t ���Iһ\���F-D�����	"U���1Oܖ����'?�I�}���K�	N�F��>�zR _:u>8�� �00�T���;D��;� ο��mAD/��'L���!�8P�̋PK����e��~2��"\hh�ԬMl��A�f,���y��+OU��Q �>ol���/��MR��T�O H:�ѳ��O��'NQ��EybK�jla�"�4j`�ȥ���=I��F_��U�@kt��[��Q$�f����ǒv�D R�!�0Q����)Za|��P�Z��-y�b[<j�BI�e���O�}���A�"�6�d�}�ʙ��ۅ{����k�f���N�a'.����P<S�!�D� u�HAEn��l�8R ��L�TBɔU���N� �h��$�D�v�Q>�� *���"�(h�'/��8�"�I"O���'�!M�� ;��p#�حx�8J�����J,�g~�+�4v3l ��Ԧ"E�y!akR��ybiD-Xy���'��QBT�P �q�L��%g�)|�X�	�uּ��1��;"����e�ڮ���	�j)n��ƋC�~"�V�A�Z�
s ڬ���0�S��yR���u�v�bP-�x�X T�˯��'���+��ȟ����_�`=z9���x���d"O�`�2dL�M�l{�iI�C��i��"Oz�#HMi�J��7�W�
��� D�� 4_��;q�__w.��O�,�j�͐�� � ��~4�d��'�n��$�4SH�HӤڣi%��O���"�$�Y�(އ����1���x�h,�DI�F~��z"OjD
��z;^��£'Z��E�A��H����/9&m��H>�g�M�P���P7LV��"��`%��	<Z$-�ֆu8,�+'c˨��9��X�Zpu'�C�v4����I�Fv�Q���)iP�J[��;d#-�Cx�1t V�cH�*�Կ����%?%>�I�)��:��c�K'�!��#}���)C���jQ��1T�]�s��d�	�Lh��G�L�2��U�1�'fy��[`�n�\l��ꈭ�,���}O��:g��"�N�0U�]�s�>��7�J/qU�(:�H�V��Uj��I���d
�*C⠒&��? �%��H�P�a|�n�F?ʕʷ�ڗ$�\H鶨݌W��;t�oq������k���H�+)�O�����91���bv&�?#Z>(�O���?6%)W�1V��������6�� �b�NE�<�+rf!�dM5��؈c��? L�,b�A3Hd�L���<`��+�dK"4% �DF-�'�y�EB�7�"�2���/#,h� a��y�#֘u	$!B"
>U���#?f�AǠ�$(�����ӕ|��A*���O�x��#r�n��MW�=颙��'�~�SΛ:%N�poZ�k�x��\�P�]@#���]spB��nߚ���oͭ(�I��KXp�z� �r�_�Ъ)!7�z䌴z g�Wrb�A�l�&u��C�,wa�u��S�H��5pi�9"V�B��ޕt2e�L��F��'�,�!�CZ!b�� �� sJY*	�'�\[��B�{�H��p�ɪZ̡�%&��WoD�����Ͱ@�I �iő.bɒ���\$�{f-]�N9�%�M�h�F.Dy���K.k� 駦?D�P��XA�b@s���O���xq�:�I(�i�M0��>��`��e��3׎�7(���G�;D�����
�v�ik��D� �&��LS�<���	��ڷ��	f��~�*����!g��v\XE>�y�b��`i��Bǹ,M68@D�X��?	P�4z!l��$#lO(@��eK�O��A��-�%/Qh���'��@��ŗ9L HmڪN�$BC��4��y� O�DB�I4�L�h�kBTeh,X5m�}�d�h��/_-?o������,� =)�l^�w�d-b���o�C�	%J�z���K�4~iQ���^�zU��ǩL���'�"~Γ?�13�G�+z�p��v#�f��C�I5BIl}0RW�����g+u:�ɑk��-X��'�"UQ�N˹};tXJ6�-O �0�'I�IA4fÌ[�"H@�f�$/���
�'3�=�(�9)��ak� f��d�	�'�"��x��pT�[�f?��:	�'�(jqئ!�$i��l��\K����'hİ �O	��dx�f�,X� ��'�������kI�9��7u� h�'$z�����{��]��Ɏ�kL��z�'x��ǌ$yy���A�"3װ�(
�'��v��{��U�f"�,5��	��'F��;ժ�f�(�!���,fժ��
�'6a��/�Qm�h�G ,]�4�'Oڌ���s�%:�L�?-�I��'P4�kӎк==$5���Q�^-�'��4;P��J�.:���e��s��� \h�	�$'~�1+ϫN���"OT��!%��l���*��P�Ӏ��4"OP`[�@=j�б�$ӟ�� "O@0���?�PV�-4�V �"O,�ä�"��{�C��7�\��V"ObĹ!���W��qeD^�_dL`��"O��z�"�"MN�<c�����Q�%D�lX���0nF� 0C���Vގ�)�"!D��D�P'V�l� %�ȡPB0؁��>D�p�1+̐x��ekU�S�6���4�<D������#Y4��)�̣��=D��h�d�Y�8k���$Fā�w`7D�LA��G�����jT�r�Ѕ�#)D�d
�	��R��;#G��<>�1k��$D��C�M�5��L�!�,b�d����0D���5kѤ/�� ���0��(E.D�;�B���I�� F��<���.�g�Lt:A�� Z0� *�͓ꈌBW�A��D\��f�?�u�ȓ�bb7��5)]�53#	!��l��i�$���W�vB��V-A�I �ȓ?)��C�L�1;�}��ׅ'����B���㔌HSP����
ǪhXlp��eN�1C�ŏ)����B(�7o���=)�h�7S���A�Z�@}c��9$��I�P�B1N��IsI�����,�*�'zC��v�ɊZ��JF��9�T5��n6���Uk^j�)�'!�����옪o��x� �a��X��#�/Kˌ��i��<&�i�|��}�S��I��gH���� @������Vs.O�zbH39��>�|�h�	u�Xx7��wA�l����d�w@�h���T?y�;�L�pKØk�1����9�,}�'�H9j	�Y�S�O�<5��&Ŕ�C`bZ�k�e �'�*�iBl�|�	�ʈ�`�K�&Qudͣ6�O�8Ɯa�,F9DhqX�O�=�h����>	�O'8p�b(W���L�%���0� �:d9�'�v7m���>ɂş�Rg*)h�Ȥ>4\�B��5[Y�F���O?�����<!1��r�	#w��Y�k�<��ύ&4�p��� 6��HF	H{�<�R�"v�
�Ξ�TY�`���C]X�h�O}��nOb���"��M8����""O��Sa��?M���B��
�2]�@"O�y�̒8rk����B=g��uq"OxP�A �CWȥ��؞{�4y�4"O�%� 9o�2�Jw�L 9�RQ9"O؄soGE�������K��H��"Od�[���,.̒d�w�_q�h ��"O�$���)ʊ�j�O�&��Uâ"O�1���(,��)�$!(��5�G"O���OB9��:ƨ��|
l��"O^H8�I�9(9x,����4t����6"O����r��=%k�C�rH�t"O���mCP��K���<�RЛu"O�	�C��W}N�S��� ��"O�i@g�,zA�1C��!]����"OLŉ$瀼m!�	@�T ��Q��"ON}��E�'��t"�+݌>q�0c"O��ڕ�I2O��`J�eR��k�"O�A)a��"7?b��U�B�~5nxؕ"O����jm��;�D��;N�m �"O(��B���]�8��GC��48`P��"O:u��ɗg�:$Y�#c��;"O��@�E�7i$֝Ya@�  >q��"O���LQ�^@ 0`��E(Y���A"OT�2��C�)�2icG�XsU����"OJ9�t,.}M�\��gY1;�0�F"O�0!G	�e.��ԇ��$9��07"O�!�®\X)��Q*.�y0�"O� �8kcł�E��4&#��"O��t*f�B�e�="�3U"O:���%t�x�	$����MP�"O�u��g�=?PQ9t#	,sN9�"Ou�s�t�����<l�TJ$"OM��P�+���@���QjE"O�����.X�pjB̒&��('"O����悎8��Cl�#J��j�"O��z��%	q<�3Kհ	D��%"O�hR6�V0Fs�m�-�(9�Ր�"OV�7�
<���R�V4b���7"O���j�5=��`�,z��	�"O��8�/� Tz:*s*Z))ܹ��"O|<�H��<jL����Qx�#F"On�	�i�h������7pݐ�"O��H��2x�^U�EMXG�|U�"O��o�W^��2�D0a��4�"OxM��D��-�\�'���U�R0��"Of,���"UM�Y����j}���"O�yY�g+K�(!#M k���"O,�r�Ê�$���FJ �����"O;�k�&U<}�PI
V����"O`M��'�"e�dI����^�:m��"O
\���KL���I����D����"O�qP�7<>�X ���%�L�W"Oʵ����k�����5�<�
R"Ov1�����" :a���4p(]Г"O�	6�Ѡq���t&~]N���"O(@�D��x�z��@j-?T�q"O�U��K"r�zX��* J�̛1"O�}�3aնX,1�*Ŧu18� a"O���m��,�\�S�@�N��=��"O`A���M;N�V��)?1����""Oj(�d
R QrL�`����m"C"O��� jD� .�ݠPi��̺��"O��+t���J��0�'�8f-�r"O���V��?<Į�9���[H	s"O �����h��ubeG	H��arS"O�0!�Ȓ�$A���))�`C"O<t+F�1k�f���D�8�Aӂ"O�`��ҼqD<]��qn���b"O��07A�wh���mߙA����"Op�j�ʌ�%����]��P��"O���b�6��$b���.i.���"O�T�C
�@� �a0�-	s0:s"O� R�����p�!$P-$Uj��"O�uA�La�$�if��;aG���"Od1v]�n`�ac��p���2"O�|��ኇy��4�2F6Y��T��"OV ���G0XPsw�o�pi"O�!`��1ح�����7���"O�
7��an����
�x��ȥ"O��sU��
p�Ȃ�͟fž ��"O�0gJ̶1Z�Uڗ([���!"OQWD� x���WAφe��)!"O�y1" 52��)����/O�E"O����ʶU�j倲/Y�D4(B"O�h��D�@����Ѝ�k��R�"O��'�L��1��M�R����"O|}���ͨf䙻5l�&[���SF"O��Y��(�Bm�R��q[��&"Ob$ZD�$8R=6�ZY���"On�eJݑ.Y�e��{�H|�d"O���sΔO]4��s�/ �8���"O� x���H��C��DAF�҃S�ڕ "O�Yy���nf�h�������"Ot �k˕xtv�@�`����C"O���5���vu��)S+sDH,8D"O��� �lː�I����hA"O�xy J�%DJYZq��@��"O! ��l�
��eCK3gsZE:"O(��q�G�5'��; `�3F
fl��"O�{���[h��n��8ڤ"Oνb��@���Y6��3�l"V"O��YR@��id�{tɻ��XYC"O*H��İ�p�t�T�&�A"Oҙ�%��2���֯ۃ	�n�� "O��2QZ-�|)BTO?�H8��"OZD�u���BeY( B�
�%j�!��2I��U0�%�-N�!�N���!�D�p�*=[��T(I`��֣��5�!�[\ƌ��W���!��'���Z�!�D��U\� �F"��1��jU�_�P�!�$��4�-b�,ֹJV�Z �dY�'.pI����8�����χ%��Q�'u�
��	�l0w��&gN��
�'�\�x��܊(����N�E2 �
�'Ƹ�Q��*�l�v"޿0^��
�'[$I�!�yW��f��z��
�'�����/c=��3� R&$0�xA�'��i�-/�DH���ӠO�-Z
�'B��S�BR�~r�kgȄ'��T�	�'K�96��޾�a�Q�t���'��}�"٬�a��#���#�'VZ��cm��B��l� =+nf���'��k>]��K�Z�����'�ls��(d���nO3���2�'T�Q@�MB�~h�Y1�ض��'xؖG�l��pC/1�p@��'�<�"���l�>iR�aU1}pA�'�T�����K�2�`���8
�'8.��£�+53@i1� Z!6��
�'`Bٸ��X_l1�0�C�;�A�	�'�8��Oъ��D1�8>�Y�'�"�J�KB�z�t�(!���7����'(��l��9:�x�F�0/����'�)���W#�,�A���'�f�*�'���ЭȲ5��/��T6�8
�'�nH�e�p�ɅZ1vՁ�ƞ��y2���C��ǐ�b�d9w�ݟ�y@��=J�)P�H|���Y���ȓ��ZkT'M�,�Dn�
?0,$��O�La��ٌ(&�B�i� �B��� �� #�C�S��s�)/^�����7��{t�]�!����V�]�L��ȓ-v0p��@6$v\ ��.���ȓ}�5@%��V��:��U$x�)�����!UڥU���6�X	1�N]��e�04SSJ^���e@���M�l�ȓ%�X�JB֑TR�iY2�������pf��xB�	�1$����"0	�l�� O��i`���@�}�e ���̤�ȓ|�*�Q�!u��<���O�Ah����(��-b� /t�Ni�
uW�<��N�][CJQ�q���a��-HŌp�ȓ#z�$�ªJ$)A��9��gu���;,���Q��&h�a��K(9r��ȓoy\%�vj�Z�P	b�i�y�\���S�? �|3" 
!A��a�� N+=L��w"Oػ&�}D�X��
 ��S"OAj��،Wd��S`��;���	"O��y�@L*ע�C  ^![^���"Onu���2_��	��I�$ �x��"O��Xϻ�9��OO���z�"OD0.�Rh듇�>O�����A�3�!��M��ूIX'q������^��!�7"�����͝Cg|�b�ƕ	Y!�$�34�Z�����?EG 8�$�(D!�$D�[��\x'�ͦ#�bFa�W>!�$�~]�)�g��-U�8�f`1qM!��֛|�5@�-�	3E��,@!�$
Z��*�1�,��AV�L
!�E�@M��3V	��f��K�a���!�d��XK� }����n�%,E!� �G��#7��u�=X m!�D3Bւ�r�,E�h��h���"!��҂{��#ԙ9�0����;�!�D�dfB/I�*��P悭9�!�G�L�`E+%@��Lz��A�V U�!�D�)ۊl���*o��	��?m�!��ݫD�ޠ ��=�������'Nw!��2%u�%���ҴH��c¤Z_!�DN
4Ѝ�g&C�yX�D�#�k2!�ܒ��ꂠ��tG.�(�۸K!�$��~�@s�S�u=�̻�/�?v�!�$�tN�4ض�#,�i3��9%�!�$�X��8q�I,8H>@3Nv�!���p�X2�\
h�\h�J/@�!�R����S%Dsƨ��)] `�!�ė�@�BȺ�-}S�k�Ζ��!�D�26}z0۲�
R�Fpm��Xs!�$�gZ�-�nO�}�&����Q!�d�[?���G�%6�=xt�@�"!��5VR�����랥��o!�d�:)
����a��{�f]4��!�D΀ �ڕ���R��.��@��7�!�Ĕ�>K- `�9�D�$�L��P"OzP#��	��9x�m��m=���2"Obٻ月2��Y�l�X&<X�"Ov�§�!^ Z@	�,+�tXz�"Op-��̘DrL`ć̽@�P��"OT)9����8y6�/����"O��(��"��`q�)ݭ"��%hD"O�icՉ��j�ECN��X9J�"O���q
 
  ��   �  �      .*  {5  "A  �L  �W  �^  �i  s  Zy  �  ��  @�  ��  �  T�  ȥ  	�  M�  ��  Ҿ  �  W�  ��  ��  ��  V�  ��  @�  �  P � � � @! �' �- �.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i���$�>Q��ۑeK,āc��/:TR	еO�'���,�r@k�� c�x�x�iY+bB䉇KxHA�ׄӏO�jM�6��TK��	��'"�>�Ɍ[���zA&��D�Hq�2BQ<S?P̐�'��L)��?z�(�4[0�`��ٴ8!!�4��'�
*m�������q)�{��d��\���䚀r�V�+�;<��{��)Z��K���ѲBKG�,�4��� @�<��B_y�NtCD៙n���S��զqE{���i����j� ��i�1B\�#
ϓ�O�zP@C!p��2�"��yv>(��3O�E{��I;Z7��@'�4r}c�N�W<!��6
�\������椚�2.�P<">�J>yPmS�e�f��N�(3�v q4��H��p=�!`�=Ԝ�J9$���� ]��hO�'
Cn�HRJ��Y<��'A����mM(<�p��=�q��ǹh�����Z�<	���y�>�1�L�8`�B W�<�ЄJ�H�m2w#��x-�%��P�<�ތ��̀�ʘ.f� TO�N�<�#�	n��(�%�֢$Xd���$�"�hO?牝��A4'��Hh;@�*`u�C�	"���(P�"xyv�[J�Db��n~���O�Н(���O�^,
c�Z{��AI���dE'�2x�%
H�ض�ʵ����'?���'��x���7:R��g�'Kn`��d��?q�'ȰY쎄 ��G��n`��'ή����D�p�!Q�P�v4� �'�H�b3�Țe ApQ�\��{5"O�M3`+�`� � �^�4��g��Ȅ�ɖ;��2�.�2ye<Lڔ̒�7sF��d!}��<-.YS�%Ԁ	��l��L��y"��!!X0�Tc[O�2e0�N@��y"G�:?���D��I���RD��y�hHP�m��ȈF��Y�#E��y2���}qx�b��R�����'��?�����1Vj<CƦ��?��0�2,7D�dhAAڒ ��@I����Nx�	D�3D��9��4WS�ț���	2���A1D�� �YCu���~ۘ�!��t���zA�'�!�d�j$�8��1���c��sp!�$���`���ݙ^�&P�&IҮ,T!�%d��]��a
R�J����[�QF!�dZG ����]!���&@�>!�V?�N�؅	���H�-��O��8�S�Oavu��䎘���N2b���8�'-����<2��:�'��M�~("�O���I��<����O�7k�ڔ��0���>A�`ٽ����]�c��p�uj�ޟH���vx���F��:|ʢk�rΔA��F~���]8�E�C��c�P�*�'��
^C���i���9�A��T �~��)ڧ&�q����1��P�W,�4F����ȓ2�\LA`�W��<ё$O�<��)���hO�>�xe`��5���s�H�s��p�6D�\�r�H�<��u��؁B��g4?ɫO����!V���sЖ�hA��:��~�T�l2��Az�y��'ա77 ��%F0�IA�����&��@�y�&�U$j{�dA�d/D�P����� <Y��(TZ���A�?�IS�az�h],8T"(A D�?e�Y�B)�M����s��x{�f^&�~�*���?Z�ZY��"O�X�T�L�.AV�ZG�Α����1OH���df���5K@��B��Z�k!�$/Ei�M;�䂅}��0XUfܢ_!!����AsE�e����߅!�ѵ
]f�ȕl����3/�!�e�V�
�M
+����B�"�!��ǟHH4Pɱ@D�d���QQ@�y!�Ȗy�~��VA�tI�'mӳ>f!���1L�0a��3J��(���k�!�E 1<�v�τW0(��ѳV�!��$pӀ�b#��K�pl�-���!��%~�H3�M�&�N� Q��I�!�D�"Ap�<i��+p��aaqO@#\�!��³m��x�pk�.vV�)���x�!�d��00b���J=nY����U0�!��6C���l� �� ���$�!�d��"-�ixk�<���ʅ��+	�!�d���̺��
X�����CJ�"}!�d��G�U��}����-�!���o{�e�$]�d���1�wb!�� ��2�2R�`D�m;�]-@_!�Ę�D~�1�t$Ϋ �>�{�Ãw[!����Mp��>#�
<i2%°l�!�����`��7�$0� ��2t�!�ć���2*�B�l}"� �,�!��=F��n��Ҷ׊F�!�$ӽSq6�x�%%au|�o\/X�!���
s�� X�nQ�� ��-�#!�D��;.��q�#�4����"W!!��͏��+S�P�|��кBQ%R7!�d�����A�m�{�ݻ`��&!��rC��C"J�j^6ps��6`6!��@���5 )�����K�y�!�Dޙr*���&�m}h�����!
�!�-u��ar�[5:>���d�D$]	!򤘩~��l��`�!����7��!�!��~�8á,I�x(q�G#�!�D�y�hcB�ޅc��	b3 �4�!�$=�4�x��$�B�N-i�!�D�E�!���E����2�R�7�!�dB� ]Ri��GC�4 UB��K�h�!�� ��aY�X����H5� �10"O���A,M�x�x�O��2�v���"O��W�	-m���^i�N�2"O �bQȃcY˃��gf�x�"O����T*�^�5�`T� �'��'or�'}�'��'	��'@&�y�@8� U�
O��N���'8"�'���'o��'�R�'��'jMe�L�0��o��K[�� ��'���'���'f��'r��'W�'���N�.@~��p�6�#V�'��'���'��'��'d��'��t�$��hk� K���-~Pሳ�'U�'���'"�'_�'R�'g.�B�_�^��A��49�ae�'��'�R�'�b�'��'*�'���Ӽ�ⱡw�k��S�'_b�'�b�'u��'�R�'FB�'jV�1!N�vw��I6��+��lSd�'���'c�'S��'S��'���'�V ��Dޮ�B��0�̈O�e��'���'x"�'�"�'R�'��'������.-np
�G+Q���2�' �'c��'�R�';��'���'.d�P��C�k�Y�0�*$�"3�'3��'xb�'�b�'$R�'���'=����"
�{r�@)�ǎ%I~A���'2��'b��'Or�'d��'C"�'<�e�B�K�%���M 2 � 1Q�'���'�R�'"��'M"�m�����OR��DR&��q��#0Pt�u'Mxy��'��)�3?a��ibA��ӄv ���������;��$K˦A�?��<��#E<W��	At�����-,b�3��?y�k �M��O��ӝ��M?��7�O}�C�ޱc �B�� ��Ė'7�>)����80P b*-'�:���)���MS�@F̓��O�B7=J��̌�A�� -�&�#�f�O��dz�֧�O�l@�V�i	��ܔt�x�*Ħ�A�8��-�J�v�,�(��=�'�?�R��" Sх�%h,��:���<�(O��O��l��0:.c�Hz�
[|y�"R�%���$��d��?��	ڟx�	�<ɭO�!LT;i�j���|������dM8�*擁dL��ݟ���ê1e�]�f�/��X��Hyb]���)��<��� i3�,��"�sxiqF��<���i &���O�(n�g��|򥅖nP�<*$�L�8m�t+��<����?!�K0)2ܴ��m>т��ZRȕ*�E	)���Ӆ�<�ީf�<��<ͧ�?����?a���?��-ƴ͠i�V�t�)�/����]צ�tN��\��̟�&?Y�	�1b =���S-:L�3NHWw�TȪO*�d)�)�����R�>t�xf��JU���3�H�( 2��'!*�	�B�����0�|�R�L�S`Iv
@��&ɏ>\���;�L%�OlQnZf�VX���s��Y`�&B�%����t@�P��@��&�Mk����>���?ͻl2A#�E#F��[o��_e���'o�<�M[�O|��/A���D����w��� c�G�@u:��Ee[2�B�Q�'��'w�'���'V�X��=RI�ht�޷~lL�A�J�O����O|�o�3X����|B��c'����O� G:m��ɇ��'�X�L"�'�צ��'���9�kRho�� TH�4)��$;V�
j�"��B��'��I����ԟ ��~����`M�l(+A�X/}�!�	⟈�'�46����O���|�QCaߖ�p��a�|a����<I�Z�I�����r�)���
�t��Ui��k���U_�x�0���P4����,O���?Y�:�$P�a.<:!B�V�q�"팹*?j���OH���O���	�<iV�i��-xဆw�T���Xa�<�8���72�'��7-2�I���d�O6�z�A��8DV��IyT��Jvm�<����M��O�	:B$T��Gű<�3-�3�������4�^�!T��<�)O��$�O��D�O:���O2˧a�4���x��AX���0� x4�in!�%�'
��'��O�{��.�s�l�$��-I��H�e^:�R���O(�O1���up�&�8~#J��!�/>5l��
�����ɹ|.��c�O��Of��|��rYP� G'o�,p)����!����?I���?�)O�pmZ�j�X�I͟��	��,%�$	��l�v(#���6�68�?�uU�$����'���P)50x�b����"�X��-?q��[	9�!2��B�'8��č��?a ,00#S*^9��8�+ˁ�?����?���?���)�Oz$`�j�<0�\y�3ɊA+�/�O��l��1좕����ٴ���y�)�$��Q7�#���f�2��������ןh�v������'^�iYTl��?eҀF��O��K���9+d)9�" �hi�'�i>��I��Iß��I��60���yťIH+�����wyrcp��3��O��D�O�����$�l}:4
��
.N�l���QXS@��'�r��P:��B�7\,�FA��9�^�*�nԬVV�ʓa�`3A�OPY�I>))O�T�4��<�F�P����qp�?rr�'8�'��Ok�I+�Mt�[9�?Ie	ÛC�.���ݤc��5��P9�?Q��i:�OM�'���'�r��+oXa���G*AOI�c 
 Y�j����i�	(Pd͠��ORq�B�� h���O���&�#'��d
��I=O��d�O����O"�d�Ol�?e"����^�~��&Ҙ<��yC�����	͟���4s%<��'�?�նi/�'5��KC�(2'����Ԥ\����u�|��'0�Oc�	�@�i�	���$�)B<����"8�*ч���5���<y��?����?y�����7�փ#��|3&:�?A����D��Y`W(
ß���ҟ�O�r�C!I�_xN��שȅm����O�u�'O��'ɧ�)�*V6��C'�X�j������a{`e�jN�xѕ��<ͧpm��V6��c��BE�(&9b0k�F��q����?����?I�Ş��d����g���`�$�V}lD	2��+LW�����A�4���?	 S�<�I�e�`Ӳ�ĕZ�b��t �<��������HǕΦ��'۴�81��m�+OB(^R2��"S�X8^��y�Y�l�	��I�����֟P�O�8��gn��Q�Z���e�����M�x��f��Q���'������'ZL7=��Am��OӾihר$Pi��E��O6�b>�ib!@ڦ��t��g�H<%�\����ۖQ&�E͓y���+�m�O�mQO>*O����O�@���Q�F��9��CK�A@r]Zqc�O@���O����<a׿i�tU�a�'���'X�%�IO]��C�d\����D�M}��'R�|2��M4�A�Ԍ��"�P�85ϛ<���9{E੊�o�7|1���y����:n�t�Y���9\�	��F#!�$D�W� ��g΢h��DHF�K�sZ���ma/[ܟ|�	��Mc��w�D �0�8�@`�m� Q��'#��'�©�_����h�%��G��i�Ds�5:��ƃw]��T%o
��O�ʓ�?����?y��?��sK.��툓M�A���~��H.O�o7������x�Ig������W~z��G��%Qeh�ZģU����On��5��*���C���z4a %�>A��I���=1l�˓:��M�e�Oа�M>�/Ohm����8R�
9Ip..�,����O����O���O��<!�iP��s�'R�:�e�18:�;��5UN�7�'�R6-'�	�����O*�d�Oְ�����.�"��ȯz�lӐոe�6M=?9��F62-�|j��<��?Tj
}8P��
W��Y1Mx�$��I怹��.;' �!�
&iQZq�	����	��M���k��Fdӈ�Ox]�	��[Ԓ�r`�G=0����7�d�O0�4�^��Iz���^<Dj0%�6+�C�(���ZZ��$RZ�Ip�IFy�'?��'2�J�+lJ)q���V�LP£���B�'�剱�McFF���?����?A,���SHQ�
��i; j�)Kf8��G����O8���O�O���.(���g�ZY�L@�
U�q��]�2��f��]�5�&?�';�
�$��pq��Q�m��2x ��������?����?9�S�'��Uצ�%�?O7���1� c��x�)Q>�����<��4��'����?� oًqxx��!�`��q9�GL��?9��P�iܴ���v�Jk�'���-U,4�a���6{���r��3&���I_y��'�R�'X��'�^>��`ߐf�屴� 1*��9���M����?��?!K~�tݛ�w�R��ro�YT�GlB�Z��F�'7��|��D��v�V:OL��QL�{���a���
��]2�:O0-`�N\��?�p�1�d�<y���?y�������z��"�	��?a���?q���L��&)Mß�	�����J	5Ym*����.�8�@��Q_��Rr�	����F�I=.ȝ�+�_6r1Bϧm�� �0�2�b��Mc��� l?���[��I��ӷ�4�¡�K�`�|B���?a��?����h��܈5�ѣr@�u��1kgo�1|���D�����lT�������M;L>I�Ӽ���� �"j��Z8��S���<	���?1�]�FpCش��� ���(��On���w������j�8n�&� s�|"Z���	ԟ��I�(�I������>9���a��-d�z5����QyB`�8�1���O����O�����Dʺ_�������v��4�� T�E�'���'rɧ�O^�$�����Na���(/!�&�6�h���O:�@���?��,�d�<�S����M�ō�8�J\�Qh����O���O�<�`�i�l����'|0��ɛ)^|�yAF�S��+��'�7�*��%����O����Ops�eB�&�ޡG⒓i��$ˣoRH9�62?1���>ݔ��(����!3��Pp�d�!A*A�5��8�Ek����ԟ�	��l���������1#�<�0`ע�Х��j�?���?ْ�i,�Y��Oc�)gӦ�O��`�`S(b������dZ����O����L`ݴ����m�D�e��k�����]GP��e͔�?��a �$�<�b��1
5����S5u`��b"�1�O�4l�.�*��I˟���I��ߚ!�0�e㚛;�@�NG����V{}��'~"�|ʟN���[	�^��'�_���\#�������2fO׏{ul��|JF*�O���O>i����{�F]a�B��Ta�~<	t�i��]iǁ�4%���`ЂB^>\�פv2�'�r7�*�I�����O�V�\Vz!S1A�(vn�A��$���?���pA�d�۴��d��~�|���Y�� ���rΧ
ɢ�Zti�]'�dCd6O���?q��?���?�����	ǧoI���T;0�y� (��"��n;[بP�I��	L���`�����GJ��`p�*L�c~�!��1�?����ŞdY���ٴ�y���i+U��3p๘B�F+�y���R7�E�	�)}�'1�	_yB �(0�@����%<��Y�MX��0<�c�iך�Y��'���'�|�@I0P-�`�%E)��z���SW}B�'���|��--����	W3�F!��Ǯ����F��2�|�'?QQ�O���Z���Snݥ%�ʠP���*,���d�O��D�OX�D=�'�?�o݄�`F�Y�C�j�5��4�?ɓ�i�P�c$�'��x����]
'4��c��˒��0%������ܟ,��ʟ�s�)_ܦu�'*LIA"�b����I���� �}��6O؟�����OZ�d�O����O����)1�E۔ �CJ$���BEH�ě�"٠(�'����'�0�%!׆"+�d����pđ�7@�>Y���?�K>�|Z#e�|>`(�0oÍ w�h�@)_�4�����CG[~R�R�p~���	�6�'}�ɥS�%Qi�vÌu�'�O<vV����ڟ�I韨�i>͕'�7M��*��B1~,����B�r�ܐkS�>B�*�d�צq�?�TV����ןD�	���Hb�E\���¦��A h$�ǩO��-�'5���G�?1�}�����5:�CY W�E�q�!�N��?q��?���?1���O0����+r� ��� Z�����'���'��7M[([\�)�O
�n�`�9%�\k�� !I޵�cތYp�`$�4���擄V��lb~Zw��@G�G�\`��,[�	a��1��uS��s�	Ny��'���'¦�<_�.H`���lH�9���G�~"�'��I��M�f��/�?���?a,��$��� Z����l#`��US����O0���OF�O�S�9�.�ya텅a�N��ɞ�4����s�(\�>(8?��"�'��%�P��(�.2>�q�ˇ-���w�D埘�Iǟ�I͟b>}�'��6���"F2E+���g58� �l"1AqD�OD�D�ͦm�?�P�D�I�s�܀�{�� �#NԪ{RR�'h���.�����-�Z2�)�9���ࢄ�Q�"!1���E�ľ<���?����?����?A/�:(C��?@1�*�;X�.�#�ʦ����_y��'�Ob���Y�����Ү��n>,�5�^ ZJ��$�OʓO1���B#p�Z�	�4rBi�t+�`k�`�_���'�<e
�!Z?�H>�(O���OPjҭ�9t~���!8j����gn�OT���O���<1G�i�:���'@��'�"���߸[RhW4{���7�D�}}��'��Oha{�n�:+� �@6�i6�� ��D��o�!�<�(���"���^�T�d�1��e�w��QX��A^����Iݟ4�����G�$�'��yУ���$�ڼ �Y;.������'� 7m�1p��O�Do�e�Ӽ+&�.V�LE�B˸d|�Đ���<a����D�(�J7�;?AƧN<2�).�����8$������)bE�K>�-O����O����O~���O�|�$%P�_'2�	�ʒ�W.j	�a)�<��i���{�'[��'�OZB���@[%`[;R!�y��L�Q�N��?	����S�'/���UDڜs�ݱQ�ɣ_n�[`k��E�Qx-O&|isN-�?�F�<��<9ӭ��|��@J���zAB�K��B6�?����?����?�'��SۦX@ٟx)f(I?s<9r�0	�j�����ן�"ڴ��'9���?����?iS�Ƥy7�Ը��Ζ$��͒Q��2+H���4��dF�hD������Oo7왺��t����)�ꑀ�y��''��'���'��iZ06V���C&�%G��@���F���O��Ŧ%��L`>��	 �M�M>��N8DͲ���mR�Z$yɄ	<�䓮?���|Z�[9�M��O�NE�	�&eh�-b���fC�=��P��O6hL>9(O���O���Ox��1���=�n	�ч�|��e����Ov�$�<AU�i������'���'��	��4���G\�DXDo�����J���ß��?�O��h�g�Y�T�a2 ;Ą:#������HU���i>Ợ�'`V&��0D//񃧇��s�F�k�%�����I���	��b>I�'nT7��p
b!��.�x����c�@��!�O������?��^�����5��cÂ;_�b�v$]Ey�������Ҧ9�u�Ƃ>^���$]@y"��Yc���q ��eܕ�JD�y"V����|�	ԟh��͟��O��l���_�h1�m£Lf0��mlӂZ�K�O����O2�����Ȧ�A��{wf7$��i�-�<{���I�P'�b>�� ߦ5�=Y�խ��Ig�ds�bC)]�đ�^�vh�dƬ��&�p����'�:̒�oNg�����G��9z��'�b�'�[�,��4;��I#��?�����1L�?���"�k[�0PI>y��.2���x�Is�I/Q�P�")��
WZY`����\���6���ͽ*�x�O~��i�Ol��RO\��c	�b7�}�!
)�$����?����?y��h�D��ِ~�
Q�d�܈�<)��Q�S��������0�	��MK��wό�����H)�P�	I�\=a�'KRW� ҩDڦ��'�I�D���?��� ��r�g�8/���Z�f<�!�%��<a��?���?����?!QO���Rd�6�B�9Ƹ��B�>���禽�i�ޟ��͟x'?�	�!�r}1��@.���i6u��e˫O���(�)�<)M�a[���Q"fd�%%"�:���e��'�� ��lʟ`ל|�\� CD��{�T$�B�_#"��2�E�����矬�I��SEyrm���0�x>iA�1� ���K�SD�u���O�l�B�&:�	�Д'yz< &D��F���R�)
K�&m�T�� `(����,�ԂӜ
�4��d������3#��������-K��*rNr��Iן����I����U�_4M4��&��AZ �� (� �?Q��?)f�i��i�Oc�(jӞ�O��K ,`&���=xI��G8���O4�4���ĤaӞ�Ӻ��V��B��
5d����a�uF��cM[x�މ��o�Ym8p9dY�5`�l��T�.���YB�u��/�I�b��3��%ymJ�[��
**�����D�sA.7���F�a��ɩ�B�]%1OXx��c�-�~Ї4kpy���(=��JA�Ƃx$�qˆ!�~_r )B��D|(���z,:�A6� �<��y/�<�4�c��<L����ŃQ�j!j��&hn�bg�Lvl��)���0"&�*`B��aE���E��ݸ")'U|�:�荛i�^��a�S����b�h�,P@%L
0I��a��iAR�'�"�O�Ũ`�
0xM �N��x���Q3+&�$�OT��Q"Yb����s�X5��8��rf
F3'D�m�ayB�S��6��O���O���DX}Zcm� �c��#�
X�CC��������Id��Ix�S�'c|��Ϟ�G��1
j8�m��j�����4�?!��?���|��Ixy��C� ��4���Ӫ3�v�0.���Żi>��0��8��ǟ���+��8�����T�aG:�MS��?	�*�@��U�<�'�2�O�5"�NW�B��m��"��dQ"�J�i��'3⁲�'��O^���OʩC�dPo>���H?�Z���
�	��;��8��O����7�5����@q���4D��M{P��1w�lM)�W��xBM���0�'B�'�X�����X&3G�9�v��vx�@��ˌE)�O�ʓ�?�K>I��?�����W��(���zQ!����6�jM>���?����D
(��ϧqjK�`�,d�����fUuiҝo�byB�'��'�R�'�,����O\�I��R�z(��M#'p�P�\�T����ByR�ƚ�맇?A�@A�NL�t��5}���N�rś6�'��'�"�'�6�Z��dŁ�4x�q��'iN�P�R)d؛�'o2]����������O��գ�`�)*��ؚ�D8� Y+F�	r�Iɟ�Ɏ-�(�?y�O@zu��:����im�����MS+O�eؑ��E��۟����?]�Okl*jtܽ!�J��:�>�9w,�5g��V�'�b�Ձ��O��>����ǚ8��Q�wØ"5Vn��o��@�g������՟����?M"O<�'M?\� 'c��S�h)�(^)�>����i���'�2�|ʟ�D�O���1� k��M�4G
1S�)��&Qܦ}������ɚRdڄ�K<ͧ�?�'�ภ�̏;L]j�
\*]����ٴ�?�I>��S?�I�x���4��#.�h%���!���$&��M��FB�P��x�O���|�%f�4Kt�Нs��U���ӇY4�O���,��|Γ�?���B�l�"Ƒ7&�n0aQHI�@T!(O����O�㟔�Ip?�0��+�:��$��B] ��T�����m#���L�'��f�	d��)Р�Jqr��^>�@xV�Jڛ��'�����O�ʓ5%��mZ�(b�ˀf^8#Z��#��0w$pO,�$�<�P���*�|�dCTNJ���/(�R٫5�#`���my���?)/O�$Px2C�k��
D�<r2�q�끺�Ms����OD��0l�|R��?Q��%�X�ϼ|�G�Rb�KP�5� O*�ĵ<�a�L��u�cļTg���gG�.�
Af厖���O"�F(�O��$�Of�$���Ӻ��F�Q���±�
.�"�Z�/]�����Ry�.�O�O~�i	$D��@v~��;�4U�������?����?�'��?�i�E�$fT`ɡ"UJ/�t�K���䔱jV�b>A�	$¾���!�/<B9��I�`F0@�4�?����?)�"&v+���D�'�2�҆�,����T~`�$�D1iҐ7M�O���<�\?��O:�O���7I�/J��Ĺ�![_u�`�P�i���8V�	����+�I�I�~Y��G��	����7,S� ���O<y��Y~r�'���'��O��,	�!�#JN����[o���&�(���?A���?)+Of�$�?U���T�q^d�h��|�CfDeӀ���<���?���򄕃C�\�̧ ���2�L�C�,����נGZ`@lZsyr�'��	��������a�(+�
A�l�ޥ!gi��*c�ǖ���O&�$�O�ʓd�`� ]?I�	�l��4FjL�Ajܠi�Ώw����4�?1.O|�D�O���W�Kz��O �	j���q"��c󀽲QD�5:b7�O��D�<)P	5 ��S���I�?�v�Q����̀�
OR�
����O���Oj��C�?5�'o��7]���/@�y��=U^��S�tz�H�M����?����
�W��#��)�%N�&��i�P#ѥU
�6�O��D��2H�Ifyr���'uD��@�J�N�
��f�23\�6����Z7��O����Of�i�k}R]�H#
� �9�P�F;�N@�rk��M���p7�i�vi��'T�I�P����� *��	!=�z]a�o;r@}A��i<"�'�bKC8/�V�����O�I�$F&�!�NיU�xzD�Z���ܴ�?q/O��0�4O�S矀�I��$I^�j�@Ð��~t��0$C�MC�pp$P�_�䕧oZNy���5FKS(�K�:7G����H>Gr(��'��1��'��	�(�	ߟ��'�|�V�P4g�%�1�r���ʀʀjM���$�O���?���?y��X3F�1*V��m!��ƣi:���?����?��?i.Oॠ�h�|"g�8Rd6 �h��`��d������'��Q����Ɵ����?�l�<n	�ƀ�N�`�2V�k�J�lZ���	����	IyBJ@7xXD�'�?�%`� y���Ae� �0�\R5!&h�6�'����D�����Oi����M�q)ÐT��S�4�����ͦ9��ğ�'�����~r���?1��C6��C�S�s4�уD�������R���I�<�I���"<��O������>A����$գ���Ѧ��'eR�c��~���$�O�������קu7��е	6IY. ]RҥX3�M{��?� ��<q&^?��L�'
]�����%���2�]8��<o� 6Ri��4�?)���?��'qx�I{y#��< `�!�׶xBhl�� &|^7�T�(w�$(�d$�Sџ؁�(S%n%0�s�㎫;���;�k�,�M��?y��/��P2S���'Z��O�=�VL�"��x�HƯs��=�i�RT����x���?����?�V�; ���bHB$�E�����ش�?��n
$ez�IKy��'��	˟�Ohą�%c�&�H:c!�:'���6�����$�O<���O&�d�^t+şR�L����IeeVu�#�M=���dyR�'i���,�	ş\;Q��/^y��F3��z��/����ǟ��	�<��h��'%Np�e�f>��3oI��x��*P:k��@դy����?�-O����O��d�1l���*�(AQc�O>P��j���&�oZ埄�	̟���Dy2Ƕ'��꧌?��<��� �M��ic�����Q~�o���'���'�b��,��	����)�P��M�6��Q�v�!2�yӤ��O$�}��p��P?i�	����Ӣ��Uq�֚ ���숀Q�Tyr�O��$�O���*%��ĭ|Γ��t��[�5����=+�XqӀ̂�M�*O&IP�^ۦ���ן0���?1p�O�nC=<�����_ds���/ӛ��'�2#�,�y�c�~Γ�OH�P�G �<����&��
 T�{ݴ&��b��i���'���Ot���'B�'��Q�ҧ�9t��`��"@X �Bf�uӶŊm�O˓���t�ߟܨF��̠�p`#�7\}��PQ V��M����?���7����T���'��O�MZ6,�|Jp�zfk��[\ ��X��'��x�O���O���O���/�$~�r]���W<��C�������I�_!T���O8��?�+O:��ƞq��*
:b��i����Zq��[�,�wFd�$��ğ�I�����y��Ӆ&�"Q�6�U�ڇ>�vQCA�>	.O��<��?q�m���2��^�b�,��D���IjƘ{1��<��?Q���?!���d� �A̧9~�M���=��[���1#G�}o�syb�'������ş(Ѵ�g� �4kKo�t��L�o��PQ%�'����O���O>�EʁI�]?Q�	oZ�`�ph�
Il��!N�F�6`"޴�?�)O��$�Op���=ZY�$�O6���^�[���70#^]�d-�����n�ß���ky�l����'�?����Qo����P
b;V)QElT�v��	������t�W�j���y�ޟZ!!w��b&ʸh�f���T���i��	�z�=�ݴ�?i��?�����i�-`eΡ1�t�b�0B�Z�I�Cj�.��O>�9OpH��y"���P������:-���(W2�6��W<�7��O���O���x}"X�h�E�k���q"�d������M�gA��<I����d4��џ����W�"-X҉ �,^H���k!�M����?)��_9���3T�,�'���O��y�B�nՐ�bU�V%6����i��]� �p�c���?���?q�Z�w#bQ�JN?_0Pě�!��C���'����gd�>y,O��iU���"�heAPE˃w�h��w V�#���HĨl�����O�d�Oʓ�$$a�޶J�n̋��$��l
:(�InyB�'g�	�t�Iş|��_�u��_.TMVi���Z��������蟔��ٟh�':r�� �v>�[�/A9�0��A)�%|Lx��g��˓�?1(O��d�O���)7���^�����>@�ZHX��	/Ѻ�l�ݟ��I؟��	wy��שY�"�k�Ι���)�H �*�&� נٿ2�&�'��'*2�'l<��G�'��,b�����@�E����,A?��\l���d�IXyB/ʟ1'��������[C���!��i�~�L���_}�����	�~՜��x��ʕ�Ȇ%���Bɋ�Q��m�Ӧ�'�0� �fӨ<�O���OJn�W$p�gŏY$̹Hpʦ��ğ$ �,a��&���}�$"��N�@DA6��
�Д8q�AȦ���k�$�M����?A��R�x��'��T񴪕�!ܴ�0��n�6�P�o|��{���O��OT�?��	�V�L�B�kC�Ec��6��'H6��޴�?���?�����l׉'�2�'���E��~Y��^��.8SC�HǛ��|���6����$�O���C*,?�0x���5N:*�"$ɹ�-n�П��kG���?!����� �YB�oD�t-N���M�k�`��U����v�P�'���'�R]���5L��dM���AK�5r;|��Ǔ2/�xQN<����?yJ>���?iu�]�FŸi���α���j�p ��͓��D�O��d�O�ʓg��@02�l�!4��8sD.\���=`����$P����ПD'����П���%�>��/B���� %�*#gB���{}��'��'���.BK�dKM|��P�5�ib�!P����+���%q����'��'���'���'d�P$����0�1���1*^n�՟H�IFy�m�(�v�.�$�����O��0鈩�ա�֑ɰ�\�	�I�K��-�Ip�I~2����XAb!�J��V)Z��U�'��Y2l�"E�Op��O���4���{�%�z�h�P��PEto�ߟ��I/[��O�IMܧT��H�qN	* ��H;�jT'@Cp�nf�eZ�4�?��?���0��'9�G�6����˿<�6$�Տ�Z(�7�O�*G��4��&��˟,��i�(brvE��h�RS`�i��V��Mk��?��]en�j��x��'���Ob-�t�@!E4�L�2�@0 "A@��i��'c����)���Ob��O"]@!	ǹY�>�(Ď�/��t�Ԧ�Ŧ���B�ڱۋ}b�'�ɧ5��!$�4T�"$�&�a�� ���-*���<	��?������	<@��L��嘃a�2G�v4����T���h��}����l�ɚG06e��l�M6͇kĎd(�τ����?���?�.Oްy����|2Rk�=�ˡ��f�B��,���O`�O���O��)� �O� �@�]�Uop`�R��h�U��}B�'��V���ɳ~on�O\���C[�����u���°A��eĚ7M�OV�O��d�<���y�I1|�N�#�.S!4��:r�J`Y��i���'�剫}�� M|:���w���c+h�y��˖5?pEq,�d��'j��'��) V�����RB�(/U)ݴ��� �'�\Mm���i�O��
T~���j,���B��N�RO���Mk��p?Y���3X�0���"��.�0�)��ʦ� �Oӳ�M����?������x�'�!9wm�4.W�� ���
�a��g����	u���?Y����
6iz���q���O�� ����'���'��{S��'�?�O� ��A&ƺd�L��f���h��-�	�I�,��J|2�d£O�R�!D2O�ŪB�� d,�5���$.�h�� "O���C���6�J�N�R��F�'İŸ� �0a�9�g� k��� �f]3h�B��%ϒZ�vӇJZS��c��B|���d�U5w��Q@udX9|���J� Ąv����L�G�J�A��Y8�@���х1�6Yu/�^U�us���cF7J� ��5�*��d�Ѝ�F��$:L�an�.�Ԓ7hG�A�r���ES��q�'�RjنP��'x"�y��|Γ?a.H��q�,!,�h)�p<9�H��'�H0�G�W�wcP!��%-z���@�td��c�V$��񄃅S���'ɖ�C��jw��=
�fE#�\&PVj����t�	R����O1b]���Er��ݫ�A��D����'�D7-�(#^
c�J�AJp���86�Pm�Fy�	R#���?	(�p3d#�Ov丢�O�xm�\I�8w+#ˢ�?���3̑���Õ&I�s�e�<8�*�Dʧ=�2ZS��3�z���*4o�lѥO�I��o�=x�bY���\�v#}��%����D�쉎V�,���WM�D�r�'G�>���$st�19k�9�R�{dL!qC䉐:�΍j�ʜ�J�zUx�&����E{�O\$"=��"@#Yx���V-D�-��L�ą[1_��6�'��'�����!ҽF�r�';���y'�%1��e�vΐ�8�.�����u<�RKR=]����'$ap�[6�|���%pm��f��.�J�KR���NTD��$�kh���=.�\z��T�Sf�������°}#&4���Y�������ą�(�O�ўx���*]lh����n�x��j2D���%�
�2��EW���֮k�D�	��HO��OZ�z�rX�G��Q��h���� K��U�@l���?A���?�G��F��OP��c!>T��E\�a�iZ�2����#���>x*(a�����=Q'��V[�9y�
��/P�;Q�� mJ�V�X�d�����'�l[��+s�l�٢D
�Izg!�"�?����hO�� c��ޯ<Ȣ)�'�
�SH�Y�0D��b�cV1CB��� �]��$P��.�	��MC���Q�_�m�ß��I�,�U�fX�%�"� f�K�H��h�I�4�"�ɟ����|
�`���$�� 'ϩ�,��L�L�n0�W�,Ox�33��DE�h��-4_�Lɑ�#=o}�x����?a���򤀡V�1��G�'��ac$�@y�D�Ol�=�)§1�dQ�4(M�a
B}0"��93�j���N�6������2h5@��f�غ"S����ߡ�M��?�-�|t����OT�h��7v���@f���������O���H�8������d�|B*��U�ꉬpV=0���
�j4�ԝ>��j�E5�i�O>�� �D8�̎�\_��I�!�#��Pub:}�U��?A��?�����O��]ó��e�dѠJ��j�ļڎyR�'��y�̝�S�:�ٵ��<Qx��խ��0<�#�Ɉ]Gn���K�4`��v,I�ި�ݴ�?���?ِ��M"|����?Q���?�;G���rF˗�h��ٻ�>��@§��P�|�8�{- ��Щƿ��	:�ɾ=<��c2l��u��it�,gk�X�Pe�#��=�!ךwdܣ�f$��3<S �j5O�и���"NN0�ⵍ",7&�@�d�O�nZ柈R��F���>��?I��U�
S����ʶB�X��!���=�I>�d�\E�Q���hT�`j�F�<���c؛^\��|��
i��P������/g���hX�t�bV	>D��"� � `�@+Tj$u�NȨ�I)D��j���o�<(hV�N���ѩV�'D��H,'�  ���Ez�5C%D����._�'�[�I�fCx�#��>D�<�T�X���qG�ŪF}p��'>D�����#X|�4$�hL��D$(D������@k�`��/>o���w� D��q��(jүd��d�V?D�hX�S��rED���rUn=D��K�Ė�i�,�A�#A��Yx��<D��J�Y-�!�;-� �(.D�T�e	p݆<Y&�#��(jw�/D�\p�j�F܎U�a�ùg���3��9D���&�ۓ/�$1"��Ý���ZP3D�4�V�Q��lZrI�5W� l�41D��x2ϔ$>��$p�f��p�� *��:D�0:d�ؼ m�X8c"��D<D�L����0(����	�� ���<D��R���q��qM��<J���8D�ܳ���Kc�\� ��q��dm8D���Am� b��4y���=`C��d�04RŤ�=&�h��s�"C�ɪ(M������4d�͖�U�C�ɛj;��AE� 6��WA�>J)�C䉇S|��Y�$�/��y@ Z�dC�I(GՖ�
)��L��xv���B��8u��+�kR1���ħܯKV6B�I����!�&�|(C��+B�I�d�>��!��/,4�Ц��#<�C��1,\՚k��c�āZ�M�C�Ɍ^K�E��K�8=�U��$��y��C�ɯI&a�+�%��ђ4�fB��04H�cȪ_��1�6�C�	�C���L�〽!% *i㞰R��p<)6$C�R����,��`�h�](<Y!ϏM+�<yg �}!jX��E��t��ܘ4b/��k�B�)��d��JC�y�P�$�0O��k�)��'4��;"@Q']n�u� ��}�&]�
�'��Up�'�_�h�)�,$qmF��J��2� X<L�qO��%٥�Ђ#䖘�!��׶Px�"O���Ζ�Cw��ف!�,tj��[T�D81A���>�!j0�Z20�&�ܖksj<��� �8ፈ�.K�<�	�=1@�Yڶ�^�֘B��0\��%�О
��x�ȝ3q� ���<�I3R�� 	�̓�~��A�[�O��B�		^����>l<!3�!&/�B䉂 � �J
��r�ܠ�S( ��B��>Նܹ��g��6� �yҋ�������]���&�u�<��eȣA�H�V��z�؀��e�<a���Y��@i�E�=��E2��^�<B0���B#1�y6&Z�<y���N��1m_<F�Ay&�QW�<��[*y�
���8b�0=)$�R�<� �	 iH&D�R �_�,B,���"OF\ T��%-�!���#L1�#"O>�k)�	�I� ��l�z�"O�I��T�4�eJ֎ۙ���D�'IN�)8�	� ,����B� ix�!�R��cC�I�3�����GY�g�yfϗ")��:⋉�?��f��c�l�)�矠C�lL�X��� .��G��HƎ+D�hK&M� Kk�q)��cfL*�Gk�����Ba��,��M��H���q�X�U�ȑK1(0��&D�B����A%t���4u�H-!�iÒV�(�CcB�e�2عd��F�&B��$s�naD@
 D�))��A7y�"<�"G� 	fV6�- ]����J<u=&)��&� ��&ބ�y2G�	H�D ��!؀ע]�y�ę� EЦ�r�4���s�(�/%0cT80��ő:Szl�� <D���CY86|b!��4xp1��}��a�/F1"i�f�*.���i%�!�-E�7�4�ٵ��
�ꔇ��&c�d��W�ik�0ڰCV��X`A���<���2@j�	3t����v�^�;�+H�R��- R�Q�k1�UExr%��jmJ��I�:�������g~� �n�~1�L���,�y��[�+Ӳ����Tp	�`��ܼ�6%�~�ӺK�e[���5�͏V�܊V�a�y��f�y2��>*&P����A,O�(I�FՂ�yb
�k����?��큣��'��D��e�,�Y$��w�
"�Y��PR��2���K���L��{�V>�[uJ�=�Ƞ{���pG�Ի��f�N貃J94o�XB��ٱ:7�ܲ�R>��>�%�ƖU�۵e��J�#�ّxrH��m�%u�'��OK�>�M�u,��>�!k4��6�� e����]�2 h0��>vl�!aၧ�����N;�dB\c� ���$u�d:�J ,������IP�FƁ�?�փ�m� S͗,�9��$*��=�x������bǸ,�<ٕ扎"G�-I h�d�ģ��/��'.��2�Ɣ7�t������fKN8W��Mgg_zT|��ț�q�䄕O���R��ZFؐ�O�I���/&Qtۦ�J�'9d���i�H�`MW�-:��{�K
��L>yΟ�rD`}6��!�ճ	�ع�Gp}B�WqnL���_b 8 \?zl���d�
�8	y��?O/$�*D혜���������'���Q:$��k�$�U��.����vm��TD�����:5�����/.W�xJA�;�|¥ȫQ�j�!d^%6�&��s =E�0��%D_��?awcҿy���Q�'��0��;�~�:�����'6�FlҕC�-\h`��NB!�y��H�B#�`������ʕf�9OV�S�\�
��3X�T�(tlb����ʐh� �"�<��A͌ћ$]��:�Q��kOl#���苓�j�����`��2*N�9{�V�/ZЩ�v>�O��'R=�;�)O1���s�	/~hD�'9
�aG��W�hy�E/�^Ȝꐫ ?6�qO�%H"�
�urmc�i)Y)ΐ`JK�db�A�T�|��	2��hJ�@5EiJ)���9v�� Vʒ�Dj�QP���l�`�ac��!%qO�	Խ��;$�X`���ͪf9~�v�8 &�ym+LSԵ[�$׏��v�&�j��
C�I6=)�$ˢqܐ�#
y��c���'(9�Չ�lób�q��D�43�19��)h� t�w�[�
�y��	(; u�s�K�J��Hq4kv�ah��C1�t��b�+��@e��<��'k\�B��򄊎@Z�'{�\�D��3���⴯�x3���L>ᰧ�78���� ��%T*=�t!Lܓ13f���ND�S��(#%�(�j�7k��XjD�{���2+��#<�$E�(���[��L�~;Ph�`mN��R剖�Șu+���5�)�de^���1�cB�u���(�Λ
y�)�DiPC�&�Y#�Ϩ"i���I=P�&i(fŘ /����� S�]Zu�<��C��tqg��"֌�>牁&Q*B��Q;,�*A9�FI�����AlE*@;�N?	|�j���7R��B� }�$����A?���z'�	T�p�#�O��JQ?��$w�1�O�<���aF�_3� ӡ*t�a�r�|�
4��`�v���f��1�ݸ'y�������?��ذ&�BMNL�O�����'���$Z>�Gx���������)G-v���%[�`���?]_��p�j�H�S�)K(�5޴a�:8�a%��^�0�#+Y�v�b���X�R���Ui��8b��ʼdc|)	���Qf�@n�M���Df.�)b���W���g�A�/�^�ʅ�.�~�p�x����)Ƿ(�d��I7��Iۆ6��L���� @�q(FD�� �lj�{"MG����o�%E%�W�S��I�Hq���`,F^��1�U�'"��d�?MFb���ujp �I�2�����'��豈�"oZZ}�Sn�~	t-�ÇP�^�)�ŗ{ev8�Hǒ����O����	��!:��9�	�ʺE��b �0�0����#��!+���S�.Q&�!%Ï(��$�4	EwD�m�;���`��\�OP��t�Pt�S�\c?ppA�9?���	�gS���{�y�o6
���=�|2���8̤�gN'�hu�T�	?gpht���d.�3zq�� "I0��<LݰI�aQ�p(�,�$cY�%��R�)�ӂB�"��OB�a�"�M���Z�I�B+ě�~�gڷ7�(DE7���I2cSZ�9PAڈc��	 ��8Rw�$12�վC���:��OƐ����O�s��Z�J��'ٽCό8��-q5�P���T�=�Q��9�Ę�^\"QS�O6\��e*C|}�7#�#m/�ܚ�f������ fܖ���gVZ�4�Ѐ�[�
�l���� ��*#�� E���('8���fiPV M	��Z^�@
�&h�	�?tz5zŋ"i��I�R�P��W���)GD�{�,M)Y�3&@U;:Ѫ�p�H�wHҕ�'*�Ћ��$ό��xc*h�� �8L�AG�<UL-�3����sdB���fb)Fx��

|����A�~7��W�)J��ď^l��sܮp�쑰�g�'y��j����O�&l9�ɀ7y*��B��DН1}4}c�n��.�7/��8��cݭyƒ�YU H�AU�I�57�I�nE�`�T�nZú����yo�(�B��8��M*`,9}�b��<)d$
=(bܒ󮛒k�ȃ' �D̓>l���Fc���"����ş��'��2���jf�� �6��t�H��s�����Y�<xe�`䀨
>��KBЩ>L���'�G�O����+8O��
_d�}K�-�PLV�QȀ�1�,�nښ/ɾ����
�
�1Na>#>	�'ћ�U��(p����`8�|�Ra/�1O�!V�\�x�8dC �S�$d�n	�p<���r�L������U�qꚫ��Q��ҝR��)y�j�X���+�b��G-f��u⊋Z�D���Ի"o�	x⫗�1%
 �<y棇�q�
��A�>@�)�Ί`̓z[\�`��Q��ɡ �=j�Ԙ�?�C%�:Su��(�ɀ-&#���GPB���1��#���:����D�%��''bH��7 �n�az2�81q��C|o����
�FCވ���37�>%��n���X�}�z��,�N������Zm�d�=Y�`�����ɑNlx�� ͏%-q�,���F�����'���[rܧGt��/P��j�'ȄJ��+!�����Pۓ9� %�����mD�yٜ$p�Lt�����63�\#<�b���s�8K��<nh ]�1��A~b�D,\7Z-����gS� )q�A��'�.9
eʎ�8n�X���N��N�0��a�X	��b�.:I=SA�x�&���Ț6n2�A�l�U��������BӅ^^�0x����x�gYt��T�1��'^أǓ�>�y�J��
�|!
0n� 6�"w�����9�*�����(5��+S.�L[���p��<�^�Pۓ:���/���1E�H�gE�̐��1I� �#5?�%/�g���<����+�:T�]e��hp���R	Y������=�k L��q�-n��Y(%#�1U5�͓[�����1��2��ܨ�r���*1!X��A�h��ɍ7�Q>�	�)��`F)8��i�Ԍ~Ű�I 6�d���ɿ�@��S�iK��S�'�����.<��lQ$ƅl�I��_p�;Bo�`�.�b��'�p䃧��;d�S�\4�0�aW8:�����Q�}���CDk����4���� ��)_�Pu;Pn'&�!��9�p>���C�߁+$�b>����R�V
��܀Ҙ@#��_�_/(b��3�	�s @L8Ğ�KD��K7�^��#>aw�Ig�ّs���4i�p�C�?�kw���,�PiҀ@�8-�� D�xp��l��`�XE5ٕ���Xj`+�$+��(Ơَt��F��������
�x�JE�v�X,�y����s5Z�
W��;^�$7��y��
`�t(7�J���Cm\��y��f~�Y�'(C(C�<�Q���2�y�"�#"���˅'6�� ���yR��4���"���hq�T�y�B�?�� ��B�b�1p�!?�y��΃wڔ�T+Pz}!�n��yRd��|N��TM��&��32����y�	�1x���%%�XQ� n��y2GM�?dƽ8� 4J	�W��yrKE%tG��2 g� YƨqT�1�yb,�&���� ��F%;�y�O�7w%��r �Z�~U��+�_�y�]�q�����DD:@qSe�ٟ�y���<��P+1BN�;���'J=�yb�_�V�B��*O8����ą��y�"X5'}��C�m�0�޹����y� Aky2��q�L�+�J��(��y���b�ɐ Ā7r6�l�`.��yr.K�(�rį!g�:E���y
� 8��A4��p��ͨa�JQ�"O��0!�.R�x3c�����d"O2$����1@��Ua7!@�'�h %"O`��և	�gx*��m�����"O�QYW�]��D��u�.�`��v"O�(���&?*�+�e�G��9�"O��y��p,������)d�`���"O0��[�I0�,���,ζT"O��xn��@�4�:�އE��R�"O�9񶃒837\���΅�D̖�!�"O0�k�2K2��4.�>����"O.|��$�턔�K��"	��"O��	q�Z7.�T�{`��	T
4�W"O�ؚ0k";.4iA�\=B�\�ɢ"O�ܫr�@<<$��r#ـ8� �x�"O�!Z%%��|����S��E��\��"O���$��7�IFk�5D̎���"OT���F+<'�u"��ڮd��M��"OR×�Ԝ�U����G����AJY�<�2�P.ɸD{!�4&D�@I^o�<�4�^�,�B�+��L�?�����B�<�dΈpI�`��.K�/.&=�ψ@�<9�`��="�sq��y� -�G�q�<��K�7݂��DK[O"��F��o�<S��>q��X
4@V�蕈2b�h�<��h�c�
9�C�]PB�T��e�<���\�@��$�w%�u�䓷�F�<񐮋�A5DQ⏂�L�ZX{�@�<�5�D�f�%z5BJ�I��|�aj�B�<�N�4w���(+M厹�n�c�<і��	i��H��c��{� H�A*�j�<�G�D>�
ؑ� �<N^)��	j�<)F�\V��B�I¡]甅�r��k�<� l�
1�&Jm�vyJҁh�<��A�|s�)�"��2���d�<�w�B�������X�����\�<I3.�0T�|�I�,�C`@Q ΏU�<yAJ�EY�`MA'h�
U����O�<�aN�6b��HXp��#�♩w�N�<�u�T+_etY34	T.5� �3G�K�<�F�*bFLі@�!Ƥ�Ȣ��H�<q�e/?֖�[F�ܢ<��40��B�<q�i�:8d���*T)���B��~�<� ��"oX �N�"��T�ǡ]E�<qb��[���y� �"����/_K�<Q���#��вNȈ��qH	E�<�V*E#"y��Ë��I�<��AO�U�<I�.ܷ/-|���%Q��ږDO�<�t�ՅjX���ܷU�>�{�E�f�<W�So��I������ @C�X�<� �,1r QR�Kd��h��U�<i�k^�mTr�S	I(֜ s,�|�<�q�+5)�b���mX$T���s�<�d�X�mLu1���&0�-���{�<Y`F۵j0�j�/H�d�0��D�x�<�h��L��q��86�ب�"j�<Aĥɟ+0A;�� o*��!�d�<�q�S�R��U�# ��2Zh�bE�z�<)�*�RYp�LP.[yY��K�<Qs! ��"4�E#^17.e!DH�<���	1B�l��Ů��H������L�<P�����ӣ��		>���l�<aA/@�<�$ c2n˓} ��/�@�<W��6��5�#��GH�����<� �b��B1cJ��Ҳ� �4��b�"O"M� �H�IXތ����5v��(J�"O�1�
= |�а#�)i�P�"OIЅ��0l���$M�Y�r��"Ox	�	6O��@eŇ?�:�Q�"O�}3d��~b8���Ē&��1��"O��1��ĥ)�������g��p�"O�����߃3�t!LW�1	��"O�|A!bL�y�.�ö)�\��(�"O���a�Nwی̫�G�d����""OPY0�ӭf%Zd��*�`�2�"OJ#to�`t�\1pBN�4���[g"O���H&"�pu�v��X�J�h�"O6d��f+�Ԩ��A?m�4Ȓ"O��2t�ӝP�ZU;E����$(� "O�D��O��&�:��I�(����"O,�q(#@�n� ���3��9s"O�9�ߺD?d<�������]�3"O�TK'J����+@�;
�h9�`"O�m:�N_�w�9#�%�%U�i�w�~����Һ)5���E�2L`Xb��Z�n�!�D����	s�:BX����BR�c�!�dI�3h��H��sYp��X�x�!�DݦV���U"Y�^����vE͊e�!�$��Yu<�!��#��Q�MO#�!��u��eb�U�V���Hb�_e!��n1�0��&Y�� �,��:�!�W�.��@%͵|�Es4Y3H�!��Q��B$�l�¡�d��!�M2(�����)O8!@��W�:^�!���y%"x9�n"S[��qU���^�!�_���tE��kN
l���گV�!�ċ� {Q�([1�lepT��	�!�䋯��'���Y7�DZs�Hd!��QYQx�Xw��(Ҋ�qc/��!�@0|�����9V���C%�N��!�d�./za[0�}��!��lˏ$�!��Y�t�De�(ٗ��pᶫ�?=
!�N$4Ǿ�X)��}�bJ��C'���,����k2�� #D�%�ȓy� ){���L������'T"�"���s���"��?���"F�d�t��*3D�T*&�Иt>��O�MK`�Xu�2D�|�(Uv d�b�@�g���U	1D�H�5F�)�́R���*.3���*ړ�0|:�(L�K�,Tt�����#�pB�	�r�,8�	��
@��"ܵv��ʌ���O��0W ��z^:I��ǒb*���q"O�����! �̬e�@�,Z��@"O�h;�L�6M@(�хI/H��UW"O.�aD�E�����ҸQ� ��"O�(Ձ����dBJ��XH�"O8 ��㊆�Jq��H��0��"ONm�J�x8h�qc�{�@�� "Or���LV�L��5!��K�%���i@"OX�HcIZ"R)nAQN�
ǶLR�"Ob�r�o�*��\PC��6
����"O2)��E�G�|�ӫ��II�@�&"O��ED�v�*��L,���w"O �� ��:��j��z����"O�Xk�&���,��T�W.tp��"OrjB&P85�d�:ak�h@fL�"O�I�u�7�8(Bq�\2VI�q"O
Pbd�.<:^4���7.��%�"O� ��ᤉ38MR�$����*�X"O��(���Z"T��!�E9(��}�"O��R��_1��6��[�N�@"O�x��솩j��R�-����"O|͙�,b�)�%ŏ�\s~�K�"Oj��b�Ǻk䜼)���z{�tb"O�� �A�"#�́�ȇ,���I$"OV�;B��g���h��G!Ј��"O��c�	Veʁ�a��|�x���"O�aCoԵMt�˂�ͤd��mA�"O:����`Ů��vFH0U�����"O�´�^Zp���z�(;�"Ot�h�'�:{�9
���z�w"O�����	"��htę����A�"O&x�Qb�t���q��9}��H""O8t�`�! �9�@�N�.�r��"O��� �S-v�� �&�?	�v�Ò"O����n0Cmh�AS�V�w>^���"O|�F�?7�D�����gF]�"O`����/��	3��[�d��"O0P�C����� ��\�j��d��"O�Y�ĝ�Ӿ��vnĉ/�1�"OlD9��9���ђ��  r���"O�Qp/5mDkЧ��.����"O��y��٪XJ-�F¬s���7"O"�PE�(lP�3k�[Aʬ��"Oz����s� �Q���p0�X"O��JA Z��L�!r�ɟ!���"O��6�>x/|t��( Y|5��"Ox�I��X�Li��P�P�H�|k�"O|�gDG1`�@�!�I����@�"O&)�`'q1�	����%�L�v"O����d�5��.�r���F�>�����S�@�@Č'LF,M[ ���7	!�d+�`@��	�dKfհrN�'!�䒦3�P�2f�,�vt��j\�S�!�D�^qh�a�;O�$�'gK��IM�����EGmt�i��O;D��"6_-v=��b�^4�339D�p95n��Rt���t��h0ܢsM6D�8��[N<��#uf�W-�ͪ2k1D�X�eOBpX"(x�P1( ���0D�\S
B�0E�`�E.�&7��eI��0T���5�� ~CʘS6HЀ�(9��"O���S��	<��12��h�E	#�'Α�Jbȅ& 0��Ra�!1����0D��Su�̴q�ܐVE�:_���aAj3D�\8S�ݨr�h�H�%ڵ>�^� �H1D�`eÝ0&H�����;05Y$C1D��B��Q�e6��q�)/�Ż��"D�(��Z�TI�H=x���� ,D����M ��n�[�0!���!�a/D�(��L�*��e�:`HѠ2O9D�,yp�>h��peCO�D�Q�T�5D���c��m�±G� }'��44D��dC�MeL�#剭f���#g 2D�l�� ���������PF.D��K��R�y�ހj�kʨ$Er� a./D���sW�9QZ�$K }�F@!��)D��XT��3V�TmhRFJ4 ς�c�<D� �7�ʘN��ip�\=S5̨��>D�(A��	�<�xS���1����>D��r�혬Or��nK#h�@�	7D��*�$K5���a�ȼL�2�0�4D�� Չ���I6\}���[
�����"Oi����K��0�S�E�C�X�1�"Oԅ��=f� ј��_"q����"Op�ESh!��rRMC�U���H�"O(�MB�@<��:�k9)�  �"O~��b V�Uߦ�B�ȜB�$�$"OT!)��� �0� �(X�s\43�"O���GF�+, �F��2��2�"Ora+qb�9m8��ׅ�4����w"O������p�GoԞC�6�0�"O�cA�
>�n�2���e
R"O�! Ҥ��Lgh���Ѳ#J
922"O4�)��>?��Y�b�x0�Dsr"OT�'�H�W"������{p��F"O������%8Y����u>48F"O�L�bK^)(r�����PPr���"O*�B�˘|n0#��DJ`�bB"Ol�!���+�Q�"ՅH����"O�-�&�m�4�Q"O�8>dv"O�*#�dܚـ��'�H8�"O�93S��@JxCA��ƥca"O���͐�9�x�p���,1�L�1"Od������t��ఓ��b{��y�"O\�#���6lxCD���wg.1Z�"O*Y�ժW`��L炠LT�l�1"O�Q��O@�T~\8�c�Ƅ��#�"OƝ"�?[��rD��n��"OL�ju`��*�ǣu�b1Z�"O���C
�+t�l�"C���B`"O��+s�Z�h-��q��?J��4i�"O�p�1�[� � (ـ"O$��n��M�b��OO�Xd`La$"O��P&A�
[����.>^ܰ��"O�"�Z%l0��C�ϣNN��zV"O�(@s�ƾXl$4�6Β�f�e"O<��eI"6��3͆�L(,8��"O�;G��O�Z(�Q�\F�	Pg"Ojm����]�~ /t�qE��e�!�dZ4 �(��Gȗ6M�fe�p��b�!��A�y/��g$ȽS��xgM+�!�P9 P$��v���"$�91��p�!��W�_9�|��×�?7䛵��0�!�d�=���P�|/&K4K]�"�!���9b�\�W`�,&s�J@/S�!�oԊ�q��O�4�u��T!�䊻	������/��M�T`\ WO!��Ҋ,����k� a���Z6R�R�!�DO�d�ꙣpc�%�~Q�*�F�!�D�<����)�(q�:�'��!�!�d������&H}�a����$�!�$�%w.D
s��$%Tf`ȥɉ"�!�DĴ&z�M�xIz�3��@�zR!��%@�vd c808��QF"��y[!�Q�D$�B��,n�n1���E7mO!�$�u8@���&Q�.��p���kF!򄑏MEN�Ҵ�!=�b���`W�!9!��̸+w��Z�o��_���U&y�!�d��"�ˢ��J�9�DI#s�!򤌎GA�Li�φ1B�Ed,[!�$ԝ�,zǊJ�*#�\�CL	.[�!�L��С "�a-*�@��X{�!���u��9��PI�*ek!�dɌa��|Ԫ�	jM�A��>�!��[���b$�!�� �CL�*!�� ʤ��M��$L�)PX�m� 8	�"O��p%�6Mڶ|� .�0<�.��"O�I�A��(氐W'k����"O4�� ��>| l����R�^�@T"O|���.u� ���5;�M�a"O�8i��޵[!~��d��y�v�ҥ"O�t!]�bӪl�TI��>ڎ`�e"Or���LL�H�P��j���T"O0���L\,^�9�@�տ:��p�r"O����m�5:���$��e�v� �"O�����9��xS$"�"Z���
"O�Њ4��'���@`&��b����"O �[Jԓ|�xD��D�w�plI"ODD��)����0�D�j��ط"O$���]�%`���~YP`�b"Of� '�X�d	P�!D&hc��ɰN0D��;#ϺI�=�Sa�<���6�9D���Ŋ#�4ݸq �u�����9D�t`���?_4\�ꀷ
�ε4�7D�d��j��?&�8���R�}]f�#�o3D��a��ȡN(����l�`�i��2D�r� ^
I����a/Z�}�<iTk1D�|z�!O�vT�ъAA˯ml
��C��
`�4,� $(oxP�#�@���B�	�r(�4�s�ȣ3�x]3��HM�B��	kt�����N�`z�/�MyBB�I}�5�䉙�u=�c�(S�B䉶p��SPmU��9"s�Vd�C��A� a;ᅏeXdy��?G.B䉔{ \u*����Z�{�'�#� B�I�>��"��͍FG�!�k̸^5�C���kTE�ogځ�@e��H��C�I ��P�_�]A�T;�˗O[VC䉏F��Q(�

Q�|��	�'��B�	3mHnmk�na
-��fՎ@�C�I��Li�dɋ�]<�R�Э�B䉉R�Y6ɀ	�(Q ��RM�.C�ɢ\��pM��:�
5��00z�B�%H�$|�/�1-�(��e ���C�	��X�s�j�/�t'� �D@�B��*t�(���ճ����Ph_�:0B�	t>E�� R��H�%�.&�C�	�77���V&`Nz��L��tF\C�I���i3ց�v�`�cf�J"�B䉋b���NX�y�2蔱!�DC�	�#���(�"� A��\"cᔩ<z�B�ɺr�P��e�Ǟ�"��j,�B�+d{ 5��'s��h衉�\�NB�I/\r��hE�x�U�S�]\*B䉺h��	�� �H��t�O�ge�C�ɔg:AQ��4?z�*��\��C�k �Mb���B%z��5��C�	&t欥�V���R��`� h]�jpC�I
L����G��	�A8��r�B�I�:`LA��(;���Į��C䉗qa`���%�Oj��@�  I6�C�ɱm?~�k2D֑7f��T��%&��C�I�+�bP�v�RLA4ap3%��X��B�	�%)�i��h�]����ةhf�B�	%*Ѐ%P��A����*f��B�	6,�J%��%��q��ÇK
/A��C�	�vu`�B�*Uh2���b���!g&C�	+%�,}��-Y "���I�/�]�B�ɡj>�1p�A8F��H��\3ӄC�)� ����j����`!dY3m����*O왺�MQ-��+QZ3E@�|��'��v$ƭ��x�q��!��m��'ߺi&�(��y1ɒ�{����'D�8�$��c���0(�q4L���'(�D@��ͿC�x�'�+l%��	�'
�+�I.-��]v�ůw���'`�%�b��2��5�H�GV͑�'v$L�t���X�k��h*p��'��l q-��%�^����	Sl����'�tC��H�Q.��a&���N��i(O$���̓x>��(�9)^�i`NԲ0�!�d����#'EʲLF�Z1螑�!��#+��i�)%��IB逐�!��NP5N�	B�'M�uq�S�@�!�W,R�H�� :[�B��d�51k!�L�kS�Ƅ�� 3;#XAR1�+D���
T�8�X�G:d@�����5ړ�0|��DA�(.��H��(S�\y{��\f�<yRJ-S��}ׁ��G�<��t�JJ�<!����nG���G��hϊ	G�N�<��kʞ�v��T�K�n�ـf.M�<���2Uu���7��B��8QN�F�<�b���L�|5 �A��?�0|�q�C�<!D��3�^JA�Fi�D�z� �j�T��9��RJ��Y��H�k^uՄ%D����Dy~N=Q$�E*R�&1�f/9D����kѠI��		�m�����Sb�p�<��'SR�@SO�K�5��Tm�<1�cP�1y"�i��ݨN���I�DHf�<��e���5��4(�IfI\M�<95Ǘ�nޠQ2A_b�X��a�<!͢\� q��D�1���WGQ�����8>/DRf��i?�Q96BI�}dD�ȓ5`�b$,/��(�gΦ̈����2�ɵ}b�m�t�]�ږ�ȓ/N4�1  &d I�b��*�^)�ȓWr���.^V��qn�o&���>��D�D���m@��rFQ"J�E{b�'��(!��5�`��h�vW�+	���y�#�$ke��2fϴ�h2� �yr�kڽ�g䈰Z^N�p��Y��y��?���PÃ�;DB���UC3�y�A�-
Y��@��G�7�z������y(Ɨ����(>!%����$ 7�yR�++�l�eIJ;��Tꖥ�y"ko��L�bǝ�~{���ǘ%��?��Y�����"Cv1l�R'L�6���y��xRA��g0*�
�蔫j��=�3'T�y�Ͼ+��Y���=e�đ3L��y85f x��8M4Qg�?�yr%����5��Z�J�\���a���y�ܥ.�h��\�?�Ȥ�3
����2�S�Oa
���wL6��ʏ?W�ey�'!��#G��8����bo�����^'�!�䜯s#Ni�&!�33m\L�� H�Q!��2�^]a@+G�vg8U��ϛ��!�d@>G�Dy�pNZ�(���� �!�_9^��	��!-6��	Г�K	u*!�ѻ~�����S:�TT��b�<d���)�'p�Jq	��2*���#�
څ��'Y���*�f�� @�/I���(x�'��Yh�JU�P�F����D<$ƚ,��'B��x��	�77z��d��'\=��� :rqi]%[������\�*�1"O����Wf��R��*{�6��0"OBЈ���mi�ep! +t�3�"O�%̔j�*�3�E�����y��'(�$V�$l38oe$vGm2�M����t�T�<�޸"#f=]~y���"D�$�Mǯ=�(�e�3W��aV�-D������$� R��F�lgz����=D���E�1_bX�aF��t��88t�:D��@FY�s�$ՠ�m�O�a -D�,*�.I) �2��⁚,Ĺ3C�&��'��|��O^�� h��1(`�4�:�ZQ�"O���aH�	����؂Ԭ���"ON0q���P��y�-���Y��"O�X�մUm�샱+Z
5�"O6\�⢄�UuJU����$=*�"OT�k7O�j�����R�e ��3�'���ܓ0@@��
yę�!]$��O��$;�g?16�"*j�L*�[�i'��xA�q�<ဤ�-^
�K�Jн}����k�<i��(oC��)qG�=\O|�R��c�<Vi͜4��P�=Aѐ�J�nCi�<�A�ܲH��@U���h�
ezu�i�<��O�F}�@"��z�*Q}�<�E��g���d�M
�#�x��0=�S�В����a>x`�8���Yy��'O`q%���\h���(���
�'��P��' Rh��.Cd*�
�'B�[g10 �<#���6�RE��'=�AHK�K�J�
P�^!11BX�'�Z�{�@	�e5�t�G�U�0Qԑ�����C(s��	
�Ś/��j���0]��'��{�L�E6�a�RK�a��يp�ܱ)�!�D́!(Zɒ��v��4y�CR
17!��{���I�$�x�������:y	!�Rf���U������GJ��!�Mm2b(8�C��Y��	/;�!��֭L�x�� CՎ;3��s(�;k��}����aţԏ��a�Ǣ;��9�l�<!	�-�,��&��_�]�@S��5�ȓ[rf�����W�>�EC�#0\ꬅȓ@e�3���Zm6);��_/�Ʉ�G�*`Ӆ�ۉ<>�p��Q}�a�ȓ\$2$;q&Ǹo���� ��*̆�.��MK�_'�雳uL��:J<��@��*_a�`fA�d��$�����R�E^�f�&����͆o~���ȓ\ϖ S#h>�Z�� Aʙ5��d��\'�d�����F�����<#^d��,��8I�O�}�(����a��$�ȓl{Lh�l	�$�Z$�s-��q����*Mn�xV� |HH2W��
t��$�ȓa��դD1/������	M+8i��,2,I ��
eF��ȇ�k���ȓ?z��k�OG��V`E`B�nc��������a�ˢj��x��ʓ�2��-�ȓUV�!L�bd	�#� T��<���p�� ��@���CA.�Q��0�ȓP����fYA��i#��C�=z��#@*�ك�($���"V��7O���ȓ5�`�t��*)f�� h��7>�E�ȓt��u2��ޠ��l�Ʉ�9�ظ��-^��3�@�_,�3�P�tN����r��P�����Y�Q-<b ����S�? .<����\��Fg�O�DH�W"O`+��Px������	�@�'�ў"~z�Ӈ!j����T/J�́�ơT���x�b��6�ĵ3Q"$P���RP �!�䁗9ᖁY�BX,%{Vл�J��t�!��G5L	B�х(�Ph�d
�p�!�+I��#R�֊�(�srdA�w!�d	,�h9�R<B��L�Κ^Z!�ĝ#��˥T�2~��J�"�8��'cў�>e��خ3=Z�:�aO�%�	)�-4�O���u<4]��*�) xԀ���u� ��0?�!�
�9�|0�bI�`�	���F�<��Q�b�U����+G(�H�$]y�<���\�k�Y3я�$s��T�W�Ms�<y���oЪ���H�f�Pq0n�<���s��JA�m9jh��"O�	��
k?��A���?VN��	����L +�R��F
Z�9]vi%��N�!�D[�X��	�,��sB4#�J;�!��,V2$���;�i�o!�@J.�d���1`� �  	�W^!��ބJ�(�����=_t�U��({>��P��(� �K�㗡,{@�9S�H�>���V��0�IŖ	�6I�BXV3�!�����q�\�ȓ�X+#ʓ�b֢Y���lɜ��'�a~�dL- Ȃ:���&�jpZ��H��y��_�Y��C�"��^l��B��y�IN��,�2�,ܜ�q�[��y���1|Yk�/]1u�2-�  X;�yR(Q(Pb��B�� Y��C����d(�S�O^��Q ������!#�hȀ
�'�Y�Ŏ����IGa�#X�}��'�R ��H�@��逖S���
�'�6)1�##<|~pL��G=��
�'c��H�йbq�<zSC�56���b�'��p%�]���x�U�+���	�r�|�ᓯaaF��e�Y:_����m\�a���0�Trg��0ڥ�[�O*��R�3D��'�ִ��+D�ĆA~��&i-D�|1�⒇U��H��ĒQ���"�(D�|�0��F��m�B+A�C�P���'D�>��ᗯ�6��M�%��(n�C�I�w�F1Z2F�֘(�(0gU�C�3�N`�#_̀�1v�H"58�$!�S�O'�k��>0h)�%�������"O����(P�(���j�%�q&��'"O���W"~Ђ��Dͷ(���W"O�I�w$���x�@���Ӹ>L�B䉷q�XT�e�P8_��YSf��Mq�B䉠�^����� d��Y�@پ"��B��3C*p���	|�W'0��q�ȓB��H�%$l�" ��A�M��=
��+��}NRi�ec��E�(�ȓ ���ŭpNf�*�%� ���ȓ-(�����}�tjW���mB��V/NE�D'��<� 5����mfj݄ȓ��1�j�7�̼��f_�>�tфȓJ�����L\�԰��MTy��-�<8���&�z�2C(��N^r��ȓ}��03a�ƣi��g�ߏu����IR5+F��c�d9R���dI�ȓ	�p�D�*
,�b� 0�(I��hN,	v��'(⠻kU�0�ȓF�4�6���Na�c�� �X��S�? �ف�m�%9X��� M���(��1"O��,L��8LIfK0�X�3�"O,�¥N�)T��� �M�v�BA�d"O$lS�e�����|Nލ"4"O��[�e�(ڑ��V�B�M*E"O��A����d�>�x%I>=:v�S"Oa��C��i���'m̽,@u�B"O`p��KN�BP�����D�W"O�zbL� �3�cT�=��"O��[&��D����R�ܮ*y���5"O|Q�jJ"��̩�@���a�"On�! �Z�	�V]��a�g���"OT4��	Ļ���f!ύJ�"��'"O��4(�2����v�V2m��Q"O
�F�6�|�1�0'��uC&"O���ĢG�B�ؕ0�bAd�q"O|m`P	�?m�����	�$Ez�QT"OB���-"�xvg��B����"O���BX� ��=a�E�7l�H �"O��k!���vOx�b�������4"Of��"��TL:P�N,?����"Oi�t�"d�s��.85�@h"O0��(�&0�hƺ,$ �f"O�YYS�L�fWv$����6��"O xCc��ix��p&�"��h�"O����Gږo"�K��F�"��S"O��d4M4�cg��m����`"Of�+��M�i�3/έ%�0L[@"O���ѡ��wR|T�@B�����"O^���N	Bx�aO����"O�D�C�ش!Ӟܨ0�B�\p67�!D��"�'8E���q΅�z��\s�c?D�0Rg�=x}��h��а1��"0��C�I�<$|H*��A2�0�A����C�ɺm]����')�ղV@0}&�B䉫K^�<b�L��X�#Mq�B�I?DA)p��(?��4��sg�B�I-]�"%qrOZ�H!�U��$L?C��B䉽{�p�T]?Yc��@�Șf{�B�p�N���[�G3N�y1�E6)�B�	oE�РgoS=�ꄸçY~��B䉭i� m�FM7X�%�%L]2��C�I5�y#tՋ�)�V� C��B�	
<v��E-A�t�Q�� !j[�B�ɗ%� y��V�DeI�.����"O�-�T���\T��)�&G�tL@�"Ox�z�v p�P���);�֔H�"O�=k�-M��|!��*-P��]�e"O
�ЄEM���Q!�GR�4m��"OD ��V�,��Y�O�� �TY"OQ 򤕾[ d�Bo��R(�P"O���aj��-��24��Q�.H�T"O�e�$aI�*
1�F��"B�ŋ1"O䅺7��s�`K��T�[B��#"O��3�F�=	��ԉ�'ے�"O�<��S��v�z��*M�� ��"O��ar�B0'q�h�����(���"O
i8E�I$S��	��g�"N��)�"O8�s�E<K���3�H�(:L��"O>�S��Հ8j�Q�01�M�u"ODh�TXȅ�vc�%*�9a"O�h%1D5(娃�1)hx��"Oh �3�/z�p-��y8ڔ`�"O�Y�B�d[�lq�e_�$��
�"O� :�ȧI�<m*]�5�76{v��"O�-��d�81Q띃l�lYBR"O���`B9Z6�-C����cq�I�"O�djuE
�<%&�9�(�Kh�V"OL�ғ���urRx(�b�\���
�"O��ce	ʰ�p�@C��`&"Ox!2�Z�$1 ݑrG�$%��{R"O�[���&wmV��vɴ��UG"O�tzac��{A��.9b���4"O�`P��3�|$;b�� h:��f"O�=�7)�d�������c �U	�"O�!�1,ʬ�J9K�i͟/�~�`"O)��o׎���(w�b�B�"O<I!rCHd�Ix�#¡l�ʨ+�"O�	ff̉;���:�m�N�+�"O����A�)��j�09��!e"O���v�W;S+�=��A�l�:4��"O�y!/8P�������\ S�"O29�焤n��t���e�(��e"Oh���M�R2%[E�^�m�:�G"O�<Z�kW��<�AG�mR8��"O�i�ޡ`��u1!�,[>Y��"OV�SRÀ�:��TPad�#=��p�"O}ۢn#>��PQD�<�콹r"O&eIf�_9rXd��"N�[vJ��"Of�!e� !NԊs��&J|*��!"O�]��Ya�e��;�t=� "Or�xb'Z�
��h
��O�`=��"OV�zŬ
�V��)���9�J4�Q"O8M���	3C�����,Ӗcl����"Opœ���;q�lɦ�S�<z��"OX�*@)P�dS��Z�L[c���Q"O.a�U�S$D�j����V5J�"O�l:�(F�� `"��I^��t"OXxr�'7MFNYb@C6B>I�p"O�<yDI�J(�)SϏ-��"O�)��	%'l��&N�4]�2H�"O�q��ݿv�x��jF�}�P�""O>1���<]�>T��)�mkԡ�"O�H`$'��0�<̓�(D	�f��"O��v�Aֺ-8�"��{�U�s"O�	ȅΝ	*�ȴbU�na���"O���A�5xPi�`�G-[=��3e"O"y�a))��8��1o'p"O��*����V�%)\�*&"O��Q
I;FF�
��Fy30-� "Ozr7&��q�X ��&J�O)�%�@"O�m�􋀺�uz��4<����"OB4�b΃�qh������$I���%"O��&��/Z��4�4Fi=�5;�"O6h��7zf�\)�/
+\+�\�"O�ڦo�V֮�x��(�ij�"Oxl����_Rt�g��s,��6"O> �@�Ǳ"���ǐ��D��G"O� P�f�|�"�F�S�:���3�"O�A����Dy
�ɴF�j�NY(�"O�ٶE��EԠkq�:o�J�q�"O���󻤈y�! d�-M(�y���#9R�4�2"��N�Zd`��қ�y/��QI�P-L��X4���y�d�!_���:b�הI:�d�_�y��\=>LK0���Bo>0��)��yr�*q�5y�2e�@���,�y2�ݲuB�0���12�H,�݆�y
� ���ӭN�����T�˝(8�c�"Oz���*B��,T�� ��|���R�"O�X@Qȗ�u�!��!�!�ĸ��"O��0/�������9u��i1"Ol9��E[�2��y����G�l�"OL��T�!Ȩ�����b�<��b"Oб!aG�u0��,�G�lyyg"O�C2�Ӯ7Da�aƍ�p���qT"OV��Uf^�`��D��!S5�@s "O�$P���:(�����K�.�C�"OX� U� K���P��ޖ~C&X@"Orx�Cg\0C��������1"O�����#��Y�eD|�  �6"O҉3��>�Z�'T�F�"O�I�uf�N=� �S%c� ���"O4ԋ%������Dm�F�d	A"O�0Q�#D�S��O2ޘ�"O�zf��zΖt���̙a�eR�"Oڵ8�K��Y��+��|�P&"O�X�6e�"V���P$�`���"O0�3�"A�D���ߥXr��!"O��x�?c�ҍ��lSLT|��V"OڭRa-�&28�� @J�:�"O��@�	Nd�h9�jN"d5sS"O����	Գ!Iu2����|b�"ON�H�WW�i�)�S����"O���᪟�X�����)�
ў "O0=����bB� �犰9��6"OZ-:U牻7[�I:�� �z���7"ONX�D�Q�Z�V��+V9ʘ�W"Ovi��_�?.
m �%S�=&rI	"Ox�rp�2/��S�n�!
�x� "O�0"�N��di���/�#�	�c"O�"��;P��M�c�G)7�6iP�"O���د}�xq	F�ˋ9�F��"O����I�:��2�0��=R#"O�`�#- 
f=��M!����"Ol@���7y���O�$��{�"Opٵ�Z�jW*�i���tR!t"O0Ш�n�4�D���P�X&"OB\ �$H�O���X%̹SM�Lж"O��8�N�1~�mIE��,TVPU!"O�A�R/��'*"h�\Ｙ��"Oz���E�I�V {����n���G"O�4!�!�5�����S�N<�0"O�����ZT�V�h�+	,���&"O� 
��,f��d�'	��l��d!'"O�X1�(Ω�b����ȔQ�
�`�"O��W#�2�pU����| p�"O@i�s�̭��(��,�{���K�"O
�tLӧ\x�
���l~p��b"O��б�N[���1��|ڮxA#"O���[���� ��b}S"O�7
Mm�
�8�Ėv�
��"O�@ �nۀD����䂾}��	r""OjM�� �(k�m��b�!�ȸSw"OH�q���3\n�����i��t;`"O0��u�	�Vj�K�J�1g�NiB�"Ov镫��B����#
�˴H��"O@)�F.C�S�a��(��(�9J�"O�P`�-ôg��=Iw� �p��"O���v(��o���!�gE
n��Y`�"O(��a��.��� �?�D5r4"OBIP�,͗:����k�1ɖ,X�"O� 0}�`�\�4�����i�b,�d"O8-�/� o�r8Vh�
}�lr�"O�l�:�nx�� � oh|��"O$���F7Xa��j�o٭-�2m��"O����POآ,�1Owj� �f"OhQ��nN��L�N��8c���G"O((c��	�@o�D5.&�|5r"O�}(� �:�Ф����/����"OFT�aΘ�~4��� �4��"O�8Jᩖ1'ƺ�b!d�8$�r@�$"O*\{��	�,�0�$�s�T�4"OA!d������ �N�$Nā�"O2l2���1T�(�z�Hˠ59؝��"Od�����R(��Ң�Ԅ4��"�"O܈bC�<d,��;@�W��D`�"O>4�Cյ5qt��2�#Ḍ`T"O�|x�C�����SaN4��@X"O|쩡*X�m#�DSrG�F˞9�$"OB�)���Y"���G�N� �H�"O��* B��TR�p%T�t89
�'��=ѶR�a[�i0E��:Q��'
����i*k4��5iSa[�'JY��.�-zRe���ۧ
��M�
�'���COF
萨Ğ|�\Ղ
�'ML�3�����닑zs���	�'�8L��h^�{D�(����c����'��i��&	�	�4��,�����'~��A��B���H�ǋ:%O0�P�'i�5ʔ�&w�Pʵ/J�1��(�'�`�ٕ	�!Հ5�q�Q�]����'G6���/0�HB���j@���'�$0
fK��+��1�ώil|��'�by�C�L�{�A�0
[�p�-s�'Y�%���^,l�{M=�$U��' �Z⌉ZG���q��h3.�	�'���[dc�/,!ny�!�P���A�'bT��i��D�Ht�ڧC��c�'��h;BF�q����Ӥ�;���b�'lQ���-cܰ�G".8��9	�'U2T�wJU�~�$l��`�4}�x��'t��IC�ܴ��AjZteV�1�'��\+�@	��*��_"f���'[��Cp@T�,R�,��#�"Fv`�
�'����M�++�MPդ��-c��:	�'a���4�˞�*-Ig�:7���(�'x���vղPr)����5V�x(�'��y�Ț'e���u�?%c��
�'�,��_�%��Y�t�ӹ2��	�'�V������kT����ʓs:����ک}N`x�k��E`ه� <^���jR8wv�2! [	<7�D�ȓU.pa�EeI7$�ڽdT�L�bP��L���Eć9�ބ� ���m�����9_`D[V��sw\M���pu���xT�c�H	�N(Kv�� z���
�����(2f�����u�чȓ���A��*e< �
��	
(��k��	ɢ�ˮb�րrpJ݋uF���<��"iX=1b��0�24a�������)rP���i�?dr��ȓ~��,Pe�?ٶM�ť44� ��bkP<� !@=�87.C�Po�ą�
��h��*�5��X#�Ϋ'>�ȓ���Ə�?"�F@�ZY�tĄ�S�? -���
�/7��3 V>����"OF Z���?6�ZQR@��챰`"O�}[�\�,��� ��/�\�t"O�(�Ad�f6h�vnV=��=��"OR����l^6	��HA�>��3"O���G:s�I��L�r�:�aT"O���W�4��Xb�؁J�
�p�"OdL�`��QU�Xi�
GS�6A�t"O~�h�O6��-%�Zr���k�"Ou�aL"<�`+Y����t�<a�䆠W@�8�\�%�ꨪf�Y~�<��偮Q��� ��"F�ݒ0�Tt�<����,D�`�¢ÛZj��
�!e�<1gNN�D2J1��.��$;Q*��u�<av _� �n�Pr�Z�_��=J�M�|�<��B\�&��ѓ2�(K�b�� �u�<1��Y����'P&q��!H�n�<�����^(�Eͪ�=)'��g�<��Ӻn���P���� ���hY�<� ��#J�|@���'Zs8,�r
T{�<Y��C�6�*�GeD'.=hC�}�<I�FY6)������.�@�(��SO�<�w@�>�%��c�]�5`���I�<!A	M�b��V	3���i�E�<��@�U)���KѠ�&h�rf@�<����8�:0��*��I��]*�(L~�<���<$­)*w�dP��.JV�<��oI�d*��r���|B�KL�<�"ń"I��B"	E�[Bڌ�vf�`�<�w�0B+����~Ŕ"���G�<i��۰o���
@D�b6�x��GB�<A�IV,Ă�9E��O7��{��\A�<���?<�i��/�s���҇�A�<�$��.@'�-�P��R�,P���RR�<a�f��<�|�%�W�#� !��W�<Q��ǝ�H��D�7e*�WbBP�<1�G˒j��A��*�|�"|Z���c�<�7�!]�r�N�R�8�а��J�<	�"p�v�(�L�m<kD�SE�<aFFv�~!�6��I�V����
C�<��	G e��ip�CZ�T���CT�B�<�q��\G>hs�#Z/˚�@TB�<�1��MҨdif�ݪ<��hv�D�<��4oށ���Q&n{�@X��z�<� c�f�� � �H#0j�:D�w�<ᠲ�,X��̀9�L���G�0�>B�O�q0!��:X�0f���[��C��>�pn��9�$��V�2B�\��ȓw���QÛ�K:J�1É0;�~��ȓl(p�j�,�\Lm�ċ�-]^��ȓa�����@�H��m�`��\J<|�ȓ#�n�J%H�?��Y(�〣.�~-�ȓ4E��� 8N�jHH�a��P�ȓ*���{B�,�"�B �̅@���?X����ʦN��<�$�M�@��}�ȓ8^
�҇*\�W��H��} �x��=b�%��{ւx8t%�aUv��ȓF�Xd��G$=*|�C�
�at*��ȓ2b���֦ɱ8q���d�doL��=z\=J"
�@~rB�Ńub�ȓ��bE�Q+v\����=-�L���Z����!����� �3}�Ȇ�q�Tk@hǛg�H19�!ٷ+��l��A��y"�U08����#��0O�6��S�? ]��E�k�6A�aȦc"dl�d"OBL�ȭK�����M �3�"OґZ���-����������"O 4�u+$&��dESv�� "O����|j���������u"O�S���&�(@�$v���0U"O|��C���^]"U ��D<-�@e�v"Obt����"�6bv��G�ʥ`"O�0��MÝJ��rI��l����"Od��B��lb��nD,�z��"O����LD)%�h�b�ڂ8�&��"O��e��L	�Q汲�!bCi�<�3F�)e��!���-"؎\�0$d�<���&]w\��4��l�e���b�<q��_:��h4�T�o�j)"��W�<�u�V>+����'�;gX�y௓R�<ѳNA�Z��U���Ĝ	6Th�G�<�a��1{j��GK�-?l���BCA�<����eҙ�I�\jl �z�<���َj�4��C,\ Zk��#��s�<ivA�W���10酸"�|D�U�<�T��8�2�閇¶]���m�S�<y�h;F�xPe	zEh= рZ�<a�Y�uZ�]��S��
w�V�<Q0"�,T��1c��
uM��F�Q�<��	C4��hq���H�,��F)XP�<!F�K�:$4�l�>%(̐*&��F�<�Q >~H�f��=P��0�6\D�<q��§v����6�l�Yfa��<�V�J�p��-���O6u����|�<�v���Y�d%�H��l��D�<)'�T:��iʮK�
��E���<��J[7UԲyq�k^+r��EVF�<9��O�g� :Ц�U�|��D�E�<�kL�S�ΐ�s�Qq�z�puj�D�<�v ��1!d=����/�����Ng�<���[����35 =��'A}�<I��{�(��ԫI�E5`���Hz�<��K�5(B�+�nրg�ʄiY@�<�"�X&ƹ�H=Jz�s��z�<QT	S�3��-�膺H눤q��^�<i�� $꼙p�6n�^�8u��Y�<�«Ќ_�
�%�[�b�����'�S�<��R�f�t��e-_��\���Q�<9���!�������'T�峁GJT�<i�H��PD��ʔ�]�\'X	K�L@Z�<%�̗bF5 ���>Ax f�U�<i��?�T��Qs<R�s@��F�<��l9^%���I�	��+0L�Z�<�� Ŭ@e4��c���v�Ƅ���[�<��Y�v8B�a0�Y:d$Fh#��ZW�<y���[`��868[��z�<i�,��f��K'n1^'�	a��r�<���?�hK'�E) 7R��a͒q�<�S�եN��-�%G���D��m�<����@]�Y��HP"	��L���]c�<��ᄢd�>4��i��^L���d�<aqd޹ފQG�ٖ
��8c�a�<���<5�j�b��a;4�b �\�<��̎wD�!���l	0�"�T�<�q�B�*��1�
79�V�� �Q�<����O�L��@JPL��ip'Es�<q�j��`^51�ғk�ܥ�Qm�<��+I��Л���'4���Oo�<� >���EO�%��"��M� xӴ"OT�a�2'XRܻ�U�K�p@�"O�-��N�6���#Юވ9���"O.�*��3�JT Q��T���q5"OH!@āهR�`�S��ҫ=��1��"Ov�b�Z�z.���
�)d�$��d"O��8a-צ��a��:o�Z�K�"OB0K�ID�LؠT��A�*V���C�"O9��ܞB��+�oʸa��Q;B"O� �fŅ#�b�2 X�.���sE"O�9�	65�\T�ծ�9�(���"O��]%$�Du�S��?j�!�"O�E��%�yQ\�Ó���]��"O��Y��[�,���*ROY�b�LɈ"O� �D�ŉR�JP��8Al���&"On����]Zj���	d���C"OJ%���� �LI6��hU�"O��#��ܧ{���\�dl��q"O�P�aN�B;FD����*"THr�"O�mk���|�Ɛ��L�Q�jX��"O�i #(�c�.��ލ?����q"O���5*�]?�ءf��4�(a"O�A�#i$h2Bd��	�^ʄ@ "Ov����{�X��Ƅ�=RT�``�"O.`�G�L��x��7Ê�FCd`J#"Ot��� �*,����=0ZE"O1@5a�[��*�B�<N5���"O�P�B�\-�ԡ)c�K+.@h�"O΍rW�V��܉���9
.�qf"O�0c� 'W_<�� ��nx ��"O�\���ب��A���ȋmn&IP"O "*E�0"�*cG:��0�d"OV�p��H�Rq��ˀ��� ��"O�|24�4�fXxvf� N����"O�1͏�X�v�r7���jXqb"O�⇣�/x����AѤ/�Ti�"OX\�g�!����!�Bf@�7"O`�x�eO�&���P�L�qd�}8�"O��Ad(Α8paawl�#af��D"OhY[��<R���a�vI0�""O<\�����d�q�� =�`�"O�Un!B=q�N�	`4:eb�"O2B��>�@����$||!�"O���Si�J~H�iǌř[��z�"O�]3%��$Gu �1ׄG�O�WLw�<�Wh\E�~]i5�͒P�~#�Up�<A��_0jJĳ�M��ZsX�
b��h�<�*Ψ,>4�b�l5�j�
���i�<9���:�J�3$�V�%A(����O�<��'/jZ�Y�F	LH>���E�<����W��E���'����_l�<)*ܲ-?�}�ь l��AH��RS�<A�4��%(B�йf�lQS�nR�<�Ռ
�-&�y����}iz #�	�c�<ae��zܨp������@���B�	�L�6��q�,`��2C�
 ��C��b�4qsT!ɤQ�ĝ���H� �B��8o��)i��;b7LP ���Jp�B�I�+-(T��U�TXJ���.:C��|�`p��_%�lQp�^�-�C�Ibq�ʅ���2�&8��HY�1��B�. FY�#�D��0��0��B�ɑ`,��ᴀ�C��M��3OĘB�ɞ=��\���?K��c��E�n�lB�)� Θ�SE�bj`��cQ�&�ta�"O���k�4����� >�Qf"O
=�Cmʠ}J����λm[<��"O
x{��2�@�i��P7W�x��"OFԳU�Q!_��`�8/&|��"O$qɗ%��(Yc �!� ��"O����՞H�4@�+I�.�m��"Oj92���r�x%�f�+�`	�"O0ly�+F8e(f( 6d��	Fi�"O�!��%�1�íqc`2"O�����ÔD��=Us��x�"O�}H�E�N,��"EA�B��A"O��!��y�8|۠ꇄt]par"O��)�`Q/*[�a���h=6<�r"O`	�f'R0x�\��	�,Q3��a�"O�X�fF�e)(}�R(�
'�m
$"OD��դ�)��JR��`��ZD"Od��AM�JxF��E���p$��"ODL��cê7����a�X�����"O���#�_
=+��A�an�;1"O�Ȫ5kP �Q���$4��Ip"O,$�
��e� \����D�6�j "O�+�+u���4F�l᠜��"O���M59D�)��X7�=["O"@�V��9�	�1�T�`�D�ؐ"Ob�I����B(�E�0�L��'"ODhH��B�x]��`�?���7"O�1:���-w\Z2��
S��%+�"O�8{�E%(���.On�D��"O2i	��P=��(�J�;}8��"O<����6aB4Bi�,t���"O���Ќ;�.���!�H_��2"O:�k�˴�4l�p �cJf�"OTx(�!�����^0iv�(�"OJu�$iM����KH>#B��I�c)D����C�F��)��D}��U�:D����CtmxP�Q��m���N7D�\��&үM�Qҷ��;����)6D���uˀ��!����L���U@3D�XX�E)�X�r����G����>D�,��ʀ	%*1Q���
l!�!1D�гÏS������-LZR�A��.D����Dt���A�B�\q��-D�H3�[�i�j�J�_�G�H��,D�x�U�O;Nk��Ȣ��Pt	!B>D��B�J�o�X���)~Fj�;D�\cg��)ꐌxb��)�2�{�A-D�ܳ6�@�W�X᳣���<[ju�ծ*D�|8#@�4��R�D9/��xQB;D�d8�G�3e����������m=D��c���5> �A���~���Qn<D���!�;�vi�������9��,D�d��E]��؅��1A����7D����2 ��� ��Y�"�֠:D�(A�Җ._\,���Ѝ�T@EO:D������nN9�T.M"�4I��$D�@+ph@����A�O�]1�4�q�"D�H���O�����76�6�I�";D��(5�B�(��e��h�n���8D�\�$�^32J�c�mY3H=�M���5D�`j��M ����S�2��u҆�/T�H
e-]�|c�u��N���<��"O��#��״hƪL�+�,Jʸ̈C"O^���;�Ztj�(
B��(�"O� �`P���i�4I%!��^����"OI�R��)|K�Ǝ�2C�Ȁ9�"O�P�6b\�tT�=���K�'��E��"O���N϶�C ����8���D:LOL�'�)UG&L��@�jĄ��"O88�U�D%h&n�(�jL-
��@r�$4��0*�Q��ɇ���Eo��gF�>I���.��'"٪����k�$�"I�Ce����'��x�����؅�A��7A���K<ѪO���DG�4(��S�V	+!�Y7&ւ	x!��7Uf� ���7�l��b�?#q����F�(d��E��b��������e�tM���qܓ���Y�Aִ|x@ ݪ%<�	�'�h�����("`�	b�0��r�)�$m@��|S��F>~@5�2&��yrF]�u����%\�y�VT �hW �hO\��$͂P�TBFB�:��5�2F�3|!��G�*X��#� >�J��w$��
 !�$��ԥR��8,H�*A�2�!�D��7�N8#�L^-c��Ӈ�T?!�$CB����q�M�2F��g	6	:!�$�$`y�s�S 3r��GG�<�!��ӻi���"�m�y�&[���D1�S�O~@�P5댄Z��8�ck�cx��'��,pr�	�(��ux�'j��܀�'�
�S���5W�2p@���Ԙ@�'��a��(Y�:���Ay)���"O�}0$l�(Z&���m�7[�X�t�|��)�*#���a��ӌp2�U��%& �B��w���$�Z��A��(d��6mU�Ity�	?�B���C@�w-<�f �!����_�"��Y/ƪFM5`נގ[�tԅ�QY��;'١?���`\#��>yU�)�I��b����ߣ0�:��B�K;!�������M�~N %YW��n�ў�'��а�����.�!��&kh�0�:D��%�μ���+"�Z�<�V �S�7D��+�g/zQ3$ŋ2e�;q&5D� `�C�B�2X*�e� vA���/5?��d�|�b�{��$񆅗
@�\��t%�x�`VI%��ht�[��P���|���acB�o������������As𤟓wb,�X����}e��ȓ|����� �&f���g�11���ȓi�z�ae��9���@��;;X�e�ȓ>�Vܲ��6TD�cwOT4e�D �'Ya~�jW%0�`����&l߈����0��>	�OJ���;!��eIcJڍn����"O���We�09���@��ӷ3����&"Oj(�h�>�D�U8m�J�e"O�%Y���#V�$9֨ <��ر@5O��=�~��'Ð���mǇ40`=i�%{-���	�'��
gJ�2m���'��= � �y�V��G{�OO4u�s�̮/f��p�DB�<^D�

���> ) �@'8]S�i
��'T���$��5^�ޑkq��.p�x�3��vL�O�O�#~R�4�$x��Y�a|����]|y��'�8�@��-Ƞ, B��U�Ɏ�D�r�'Tt�'3�\���n�r����$�-K��-�ȓV�R�����Wm�qE��|�taie*�j�	c������[�u�����	Υu��[��%lO��pP�mڣBB�pj�� �Zs�ՙ�"D��z�ʏ�N�H��6� �~���9��!D����3E��!��*Uġ�"�3D�� �y����5ҊAsU��
7����'=ўD�"܂�6(�w��zͤ݊��*D�����I�����aD1?x���<ʓ�hO�ӓ<��EmH<6��lc���$�����%?�N� M��`�%Z�	#n���nH���'wqO?7M��;�d����'�����9lў����'�L��X::����`Ah�M��}�%��}�!A��[3����NÛ�HOT��sI0ƫ����;a�S�h�c�'0�xb�B���ԌQE���'6b%�ǧ����{��Z�xC�z	�'Ĕe�2Ɛ&1Z�su���p�2̨�'��]i$�j~��!U��>V��p���9�S��oͿl#����C���@�]��y�Ŋ:h�aG%��+F��`-J�M���s��9Ӫ��y��0��� ?�`,:6"On�hB��#7s���iG;�P��U�O��Dz����� P��sG�� �͡�ޤ�!򄝎8 Xע�X\H ��_k�Q��SH>��Wj�Zɔ@	���􁆃$L!�D�����cf��V�XР��K�T1!��$�~4�'B>_�,�{u�Qt,!�߶$pb4�`@�#�8��H�"�!�$C"�)�5�^8'��Y`�5|!򄕂��4�%}N^5kS�L�L��C�	�y��3���7z�=�Х�J�C�I�
� q0�
f̎M�W�օkhRC�ɢR�N�s�U�W��p*�ȑ-L>C䉜��١s��\T�)Ad�3Y�C�r`�a��׀db�[��Ƌ2�RC�I75`�p��o�^8"*X�f���>Y�b
%tE�����.B���K0N �<	���Ӄ6E�u���8d:u�3C6J�҅E{��9O*L	SFE�4�t�g�~U4�R��4��I�P�(�=� �'�H�lj6-'���!��x_mLn��9��9D�| U�X�	��Y0(I�I�٠`f1Oj�=)F@7��!�d��M�����^}b�'!�� �'	G�ΌQ"%!Kj 	�O��=E��dH��zā.�"�L��$϶�y�m��B" D��ՑkTX�����0>��Q+0�,|au�[�Cg�ģ����p>�H<�wbM,��!Q�O���v��<1���O��I�B�<!(�(N:m9���B�5D���� 
�H���e(0J�\E���5D�8��4��)����S>�P'-?$�܀��W�Sw��G��
K������y��_)���Ra���J*�1x�hF1�yr���3͌��**l��i�'j4D�k复�Q��x���%lXp	a��1�@+ؠ��3����f��� 2ͅ2j���j'k Z�!�&{9$@��O��m� e�a!ڤlS��<�
ߓ?�e�%�.����!�)������|Q��*��4ȠBA)
����ȓ*f� ��IIQ~�c���<����=a��'�*�Y��)i�!��ѭB�^Q{�'���'�jH�lx ��^`j-)Q$�L�<���b��A;ێ�8`d�<Aӏ�� ��d��ί�^t %i�Y�<��G43���P�XO2fUHQ�[k�<A��~4B���� ;8�fx��O@�<y��֨g0Q�VN�34�.�� a�<Yr,ٯ2! �h�`��,4�M�b�Y�<rL�Z�F-f)��!i�y����<� ��3��vHxJ�K�'Kt�q"O��3@"�5:K�(hce��f��"O
�A��K=Ap����)�p@��"Of��d�;�P\��v�h�"O�m�'�8S����D�|�b0�"O�l���E�@���C5~�v��"O�ui����q����H�=^��E�"O���fkXA���Ӱ�,g��&"O�����B/Q���@@L�L<|��"O��(�e��7g$и�/ʿ۠�I�"OhD��-�P������J b��{�"O<���#�Z$G���m����"O\,)���R��#��ςC����'"OR��gIF:@����F�&' ��"O���"l�;y�T��F��#Z�b�"O0�!p�]�]X�g�8�D�"O����3P�@��S
2���Q"O*I�U�є�B=�'� &|A "ON��`��O&A ��?�����"O�P��	��,i  [;l�"O*����8����CQ�}��qa"Oܕ[��d��8C�&dv��:�"O��a@)��2UnH��Bе;v�e�v"Oj�y���1����7)C�� �"O�����&h��!v�J6F���1"O8���ē���-x���&3A��� "O�y��d��E���GI�z�v��p"O�D�T��:�.0��h�,^~2T[s"O�y�Ɖ�b�֤�e�-^�k�"O�[����dj!	�.S�� "Ob遗���i��``�H�v��x!�"O{s/ٙ��Ɂhɯi�X���"O2y���
}�603�h��	�`�e"O��
��̮Q?�8s'Æ4�`(�"OH�6�Y�X�6�1�*�
囲"OȘ
W*+����V<r�v�Zv"O<`:��Z�Z��Y��$�2ɾ��"O т�B݊$�@I�FԸ#�V�9"O*�5�.r��x������"O4�(��;P/D��%�T�R�F���'O$� �^(0��.P�s �H�'�l=1��[�F���ꍣb/��C�'��M�d/>Cr�I�Q��6R�i��'��M�򇋺6#X��1	U�S�h`0�'Fֹq�I<\H	p��M�|
�'���@7���Q�(�ehI�D��͈	�'�8�k�p��A��a�)4v����'^8�)K��
U��' x1�'غ��f��O������Z�haj�'�*hqkY����'�a�t�[�'��XCD��	d0��1K�3A]�Ņȓ!X����I$NL<��N�0���R�TE�!��[4��Vm\?[f:Y�ȓ�$Brl�D`|�1��֭ ��ȓ_op��`�Z�?���sM�B~X�ȓ3���+'��@���!I!G�v݅�Pdz]�EąI�6HpK
e>���6�� j���9X:x ���]�8�ɇ�Q�Azwe\8V�P���r�<l�ȓ7����FcAb�{ �Q�	�jq��%$��"�?V��K�o��#Ct�ȓy�������w2���ү5�����m+�钋 X��p����l�t�<��&�]���0��Iwpj���. s�<� N��3�  �M�g�.ȫ�"Ox���DĔ{��(��=�@X�Oz����0H���q����,�H]�!&��+xL��'�PZ���8�Đ���Q/m��Z��D�>H3�|3c�/�)i�x��'�Y�a8�HB�(��VC�IJ�:�6��>r�v)(��[� #8�y����ƫ��N�PӧH���B& �3cG���4����6"O��吰T�օ2˅�W�� (b!}B�
A�Pu0�$���M.-��25-�!2�"�:eHZ�`a2B�YV"��r�!7`��#��: X�p�Q"�-�F��I�C���b�́�&pȒ#�>w��#?�'̔�i���6��X�4C�Q
kӂRp��C��ўp�!�D��:�{!��1lh18�`�Q��I�+��\�5�I�"}
�ʕ�i�P����2���KVn�<��eD�r^NtiCJԎ*��,��/̤��	�S	�Gޙ��g�~� �U�7�U�w(µk*l��	�L�(4j�Z	-��a�wn��+���Oؤ����'����5S1z=ʉ�����F)��WN����/�SW����/.W��P�aB�#M"C�&]"�A��-莜
�n��(���nY�)5�=�)�'&�v�C��ԕz���uG(-�5�ȓx�J��QKG�p��t�pDA+q4�\��#��`�2�>A�q��!)����/�uA�KHJ��y�E��Re��"�"�����n����eNNF��`���������	A#P�h����}�B����D�,y�IЋ
q��U�r�r��޷;F>���B 	����ȓA���uE��X�H����Zq�.��ȓR����s��v�.����S����R��ѓ�Ⴃ<#h�傀 �B�FɆ7H,Bቆ-�4d֎~�dx�ȍ�5�v�?�[>�1J��4�
�]�N8�Cf��V�h�bR+�y"$��0Θ$V5K����C+����"��E����y�ff΍D�Ԯ�"E>T3!lR�H���C˦�y�-��f��s�I�Qx z�띶&ܛ��\�Vu�9QJCE%f�㖔�4���s� $���J�|N�:t�Pu<U��	'�q(pǊ�m*����S����	?{���F�ҪN�>��kK�R�����H<Z��'�<uZ`�Y�h��E~bB3*і��	S
��U;���l!T	�L��=as�]�wp����0A����i���ȋE	��sBͣ{���]� b�͟8f
�;T ��n�6Az��������$��2������Z��-C�O3�y2���
�eҮ[���2Ơ�h�a	�� _6��E��-c�l��OW��X�\����>�1,ǩ^�-��c��"�̰�Gi�_؟��c��P��h�׊�F� Yz��?F��b�ȗ}���P�ѧ����r�
ͬ��O+�V
,��p��f���Qz�+[�'�ָ���
-��d��&���M:3k�x4~��� V0��toC�g���Ңӕ5ۼB%3�O�X֩�"^jb�`%����E��g�<�W �d9p!��KX� )��[`p�Pu ����w;dU+`�ٌe��i��`@>Jl���'������	AJLpB4�w&zl��-�(Oy6�@4��%C�\Y'�ǖ��$A�&!45
`7��6�)K��k���h�,���է%���yZ��Q��R�i���G�ig����NH�4�i
���=�$A�6fY�_�ȃ�C��6F�a��I��u�旺#�*�8g��Q�	%I����gO�+��H�D��	E��'V0��IF�9�,��IV�W��i�K�f��!�2M�h� �I�?$Tqt���>k���f��5z�P��cF��æ�=l�ay2���+�@ F皮k�D���s�q�ҋ��cq�7M*��MBWN��[|�X���7^ܼ�RH�?y������IR|v���SJ�+o�����5�D��$�h8蠳�Jκ�$�DjC�\A���'|��@`D�M�O�aU�]�|*��
�#}��� N�2��T�Q#E�XU ���8�j��'R�@� M2�=&�
7?�`�g$~�n��&��*߬xo�Qଠ��]�]�-a5b��"�ᰅ	L����M<�G�P�3��-`PH�6x�,�!э�qy� � t����E4_���	ĪLp�&ϗ$8"��R6M#W�A�s��,��˅�̍2���P*�8����]�Z��S<,O6��e��p�H�1�_���`Z�%R�hVL\(�t�B����KŮx�MK
�T�*@C����j#)�?)��ѩ
�8���Ӏa��9pJ��p?A�dO!BwJ]	wMүp�jq�ԍ�M�I�g��r� ��Kپ\�Լi_�ڪ�ly�̟���b� V�htB
50���fګ$�Z 9��I	+v��tck��tb)��es4`M}SX�:���Y�D"1OԈ�GE��Snb�.�� �	̾(/V�b�|�/H�r���	�t�&��1i�����¤j����JF�,��?�lZ0��:שפO��@��-K;p���kp�_<�x�,��	2�!LO�m��� ˒��e�@�c�D��%�;����a�N��ț�T(���O,� ��K@���C�i�t���'Hi�֌ÎmZ�E�7	�$H��
�dG�i�<���D9�dᆚ6��5e4f�8��b����`��p k�g7.mꩇ�c�P�8�!U�Y���B%�.4<rD��v��%�"Q�RW�	��'"$���g|b@ Pބ0H��j@�V�l��T\�9p'��Թ	Ü ����ȓ}W�0��iFx���!
f�����y��8J�@�>Ulyk�kڃ4�����r�`lK�L�Xf��D�&�!�'��D�@$�s2Y�.K*:H\���'��2u�ә ����l��:�����'�"�0��	-qV"Yp�Ό�7t쌃�'��%��Y4l4"%����,Yz�']�8s�^� .�������!	�'�%Z�%��	m$	S�ɀ+�����'1	��ŕEE���Oݒ�m�'M��Z�'~ݠ���bL�	�'�đ�7�ݾ7]�A�oʗH�R 	�'���c�QP�T'[F��ƁG�<)���)-xSxً���h�<�2�){+���#�8r��;bBNgܓTP�!�3���WɅ.߶��T�9$��la5"OF��� � T�D��w���4��9"���B�O�1��3?Q��* ���ge]�+8:%R��_h<Y�aX�!��Ҁ�104��`��	,7��"�
ˡ����$��F���S�:��aˡc�F�y�`Ә>��I���OY}2���2ٌu{d�˘W�r�j̎�y�n�ArN�UFBYN���s ����XK��볠-�#��e�#v�^��EF�2y؈���F�<y��0�F�+@X�21p�H�d=`�����>���I$����	=t]�"j�W,��%b��У<� O�<v�}�%��*�|D*��1yy��0�LmG怂�N�&q�>���P:nh��c4n�,�pp�	���֦�Y>�O哏{֨����@�Id�IEz��'���g��|�'�_LBC�I�_qJ��RdZr�z̰��"�r����/C�9W-�Y�4���'��	���O���s�MѪ ��!�5͂�Dº�ߓY� ���Z���6�͌"�|������]����2fY����'��Y2d\>�z��p5�_�d�|�acs���?�3.Q9$���*(ҧ/`8Q%�R�ɂ�����X�b��WX��ɝ>x��χDr8]��GH(qblȡA�@(��hXL��D��'����sb� ��5z��7&��p��'���[�	_$.sJ����2	�����m��'U)�N���T5DU)��UmU�q{O_��{r���c�0��u,����˅��1�x"�d�7J�99�J6D�P�ua��;[Vy��_�%�ޙ�L5��;2t����+�0v�>=[T��S]RĻg��1M����i9D��C�S�(�V	����(��{��8%M:q�R-�p�)��<��FS� j��J���:��E�]o�<����Q0
��N�-��ar*m?�q(ذwt���DO�j;r�IQc�w\�C�Y�]�!��/N������W'����@�f}!�d	.%
-C��B�4�I��@
$Y!�$��^ظiʄe�;ځ�N��J0!��9=^�x%H�6F��Ip[77!��Q�[L�0Rd��~�zu&,^�$!��݃��!��n�%�hI��)��!�$�/��-K���7�:�R�\6]�!�� �Zdє<H�q�Ԇ\�F���"Op����W�F6|���-� �Ű�"O�!���*a���+�Ip���"OD�c)
�7�*�hADR�u!""O��9� C;yTH�a�J4(��G"O� ��NK#g�L��&M�80�b�p�"Ox����ZoǜXxT&�|��XyQ"Oĵ�w���0U�	�K�|`h"OP��v�Ò5""���D�)K|*�0�"O�0!ЂT'}�01CI)89���3"O�{�M}a��B7l?��YR"��y�!�$���@�+�c�Rt�&�S�!��U�aW��/�ddr�	&��5	!�$Ѕ{Y��a��;Npj�q��,#�!�$�5| �����>{�$;'�*K�!��{���"[�0b���C���!�Dω!Z��STOI�aP��
�Â��!�D�&& ђ�̶3�x�x'!�7�!�$�%R�`t8q�$����G+`z!�d6D� ��2*C� ��ԃ�'E�Y!�ɑ����h�U��Ir�JB!�$��;��yh3*��fypQ�J
�52!�dӧG��e;���Jh�˖I�!��B�!�H�3 �͊rB��P���r�!� �
4B�K� �2DM:dA%���!��V�$����rS�-Or���j��?�!�&s�����.�->��Z5��(T!�$F1:tuk�H�;< ;6f�;7M!�ѱt�N�u�K�q�Q��O��,!�$G�e�21����#N� -�"x!�D[63�L��S*KW�pp쒑n!�-�\dQ�eƦP�
*
o�!�D��# >��GO�8nLX:1��Z�!�D�1�R	Bo�q��"��L�!�l3x0i�o��<�(g��9`�`C�	�sр��匯&�m��,B�nlC�I&;�xPG��5��pˡ�.	>B䉮p;D1��P<l�<⯜:��C�ɂ^�aQ�m
�dB��Ã�� �C�;]V�1A2X.��Q�Y�C�ɋ5�h�Q�	�A�\9�A_"+rC��/r�n�[#���M��xY�d��iG�C��1YD�|�0�9�I��e�C�I�-�z�(Ӡ1)�a���BlB�	?���6.��D���M̡q�C�ɬP�^��$��("Z�0�U`�-c܀C��9p�#�O�:��=%��C䉽GMNI8v�;�`���li�C�*+�A�1/�&9bX��GJ
j�bC�I
z��,s OY� �j����F(&>~C�ɾ-�� )�O7T�(���<1�B��:?m 9�U�|'��$�TG�B�G�0y@��a�ѱ�ո�hB�	�p���(�N���q���ռ0}RB�	��P0U�V44���!@g����C䉯'ax}@�A'2l�
@!�%7ߨC��b��B�Nڽ
l�� (��!U�B�Ig7�Ɉ��+zR4y��ݑ9ߊB�I!9m D�k$;=��0�ۀ`^C�I�NF���\�e�h���[�T�C�ɺ۞,�q�Ǒ�� ����]�C�ɇ�!�o�>/I��,d�EP�,D�8��@�+*�B�iV$K��w�*D���eS,�lQ���Bբ�Y��4D�� D� �� �f�.9��Τ%H:=;e"O�MS�'�#�4�sR�R�125"�"ODR��8El�@���u30��"O�(SL��HWN�벢%.��S�"O��$��JCB�sÆ�'&� �"OƄ�G�?xz�9�B��D�
�'b�����9W: �f�μ�a:�eS�}T���� ��όA(����IGJ
YD��1[�в�	V�0¦�p��?qP�y��\=4
!�D�>V�p��L6K���Oއ+�I�e�E�@��~��S�O� �x���a��`#a�[����'5�H ���ĕ-Q��h�p�>1�c�)^�n�ᢑ��}��D9O�t����[�����?��C�t��)�D�4-��Pr/�&p��2v��H!����Ǝ B( Ŧ�}����ZΑ�92��1����5��$A]\A&i��B�_���{s拄�yB�NI�%1�l�Il���
��d�d�vx��KT��)�'I�d|�X�Bn��쏐S�
��}�$��O8ZY�tJ�S�mBH������%��y�L|�>���Mk�v=��N5<ih��c�^؟t��7��ѕ�Цt�����>���")\h�RN�3p!��QP��=1� �g����O�F����b>�U�:�<���xi��!��)D��`���=g{����$!0�,�3b'?	��H@b�"|"q��y^�8�&�؅�r%�4��|�<y����?PtQ���͢|�'`�~�<���ϝ7x>i�L�@B$����z�<� �H*-���V�G�\���t�<��BD1v�<`�ñ4R�p���\�<�G�ѭ|*
��R�4U��	�c�\�<�L�Qc�}
��,m� BJ[�<�Eφ�i}�ae� ��a)rEHT�<��L�,r#�i�r/�b8,հsNU�<idh�κ�Hg'�Ut��$�TL<aD(��^O����%�:Q*܎f�@zM�B�	�g���1�+E�'�Nt���9yc�?�FT/ܖ<3��D��my>�rd�o������L�<I�c��1�n��F��Y0~`��NCO}b�7I��Բ�C�D��\���g�%Ixm���fC��7P�����+]QP��.S�\E�O&� �<X�f�&>c�d�A�
-/�,�O��EĪL//�aB$��X���T�|����7*{Z9���8':4�*�O�{O�0hRI���
�!H(tx��Iz4�9S
S$6W�Oa�\����$W�a�%�Or
��'�ʈ�@ĉ�c�v�E��-2<A��O�3�Q,*��y�I�"}&�Ж`RXU��/)����$�T�<����f�)��Ɛ�4�r��!�)��	!aoz��1C����g�zy, ��U�Rf�Ւ�W
N��ԇ�ɝ{��D8��ѝk�j9C�l�RF �q���@ɩ��'t҈���������H& �Q���䐥nvր����}�𬣌�4��>YK�`A��zJ,M觌�&�y2E�+;����̖9Y6(�чJP�eR0���m�_�h��EÂY?E��'&�+�D�9(*����w��(�']X�"��2^E�Y3�͢v�25`Х+��<���4qn���|�L��k��ӧ�R�� ^!��ǻB�D�� �D}���{�C r*�XP�b^��M#q���_������'gZ�B�-��<��ꑪhzL\["&E���4���QM)�D�9���0vC�-/.����
!I�[8ZTw��A�8X��GW���S�*�(]����i���!�i\��/??J`�V�O��`S B�t��	��B��C#N��.ő�DݤS� mո<8����i3���$�ہ.��*_ky���'�L�S�t�`��	s��b�n�+A24���) �O�m"�Mұ <y)�&B.�L0ab%�� ���'��c�� b�$�$�Ǝ0�:Cĥ�6\ ���'�`џt���7�@y�f�E��!�����:S�0L�:���R�a�)c�'G*���B�L5>m�`�	P?ͧ{BM.R�'lRD�l�[ښ�YvnQRn�Œ)Oj}Sf�غCCP�����$�M?�Z�n�0%6�� ��H����3���!B�hK#hQQ?I�'#Y:�%)�;,ODc��2I�2 [��,5U���2"�
8�4c�f飥"ǢLz�8F$��`�uP�';}��O� q�F�P)��;�1�j]�L0�O�,+d�/WW����
�:� �3V����%��Dm��!�~RF֩��i���'|��d���d�q*�F۱^������� ^�GiP�o�~ݖOݤ�����5�ԁ�
��;���H�'y<sïc�:��S_��S>t$��&�����JU��##
T t��hz�H�<y�.�Sމ3�����(�\(�"��8��pZv�~�d������x�N��01�_�3az�kL=��p��Hc\�3Ac�g��'bX�Ý�Ϙ'@n<bT�Qٚ��炒!>���
�'69��$��(��@ݺ#0Zi�'��_N�e���I)�)�Fͅ�td.��'���ȓ�y������S�="'M��C���'?'�6q�¡9G��P�ȓ�L��6��9J�Lre�T9�I���p""g�����z� ���4��:�&�5�ћV�`�W�]�!�(�ȓ-��x�F�Q���S��[�P=��H��#�g4��C�/�I),�ȓe�Zy�wÔ�=ô�;�d�~�:���r��}�'+��oZ�X'F�f:�5�ȓ~)�3���g~�1��/L�	��8���0�Dӟ&���JdC/�t\�ȓn���s�
 �B|�ī�qF&���l��	qDÝ<�vb���GB]�ȓ-gX �%иN�^<Z��2)���h.���J=��0Ď�x @���@���O`� H�΍'W H��Tp�8�	{�p���C�RGR��,�f�S�
�&u$D3�GGoJ�ȓhF���m�4�>ȳ@frn���ȓK���a�Ď!50��\[�T�=i��̮,U����[2zw8�Um����!oU!�s�r�PWjD�:����G��8gS��
'��^8eV>�)��l"u�:Ɏ�ʵ�� ����M!���|���Ӓ*[�8 AQ�Q,�Ia��'�O� sɋIǖ�mIT3��zv�'Ş�襽U#	j}r閩,&2��0�A9M"�pJ��yR��L���rw�A1jR`��P��� o\H�pk�04"*A�@z"H� [���ŖA�<� �P6��"���H�t��UE�,Jm)ő>awK
����&]ܝ��A��h�����Ɖ0h٪�<���
&_ޣ}b���2��;��؀U,̱��J`Aө�: و��$
<>�k�CT{�r-����6F���cAû:F�O�Ss�e�HO�4��������b޴a:�,ȳj��Q͌B��!]�D��D;w����FJq t�dԜ"_N�K���m�*�(g�G���	މO���Z����G��{�ޡx�f4
	ߓ6]�=�'-G���6mS v�f�9��Jf���P�!t�d�O�( �3?�p�\!�Rh&��*�"��r�Ao�5[`�ea;?G`#}���8�(I�s�0��o��Q�t������0?�8"d ��N@�C��és|D�k�Ǔ���h����$1����*DM`1�ȋ�!�d�z��h ��ô	Uc���Im&��v@~؞��uf61��t�7���j��s�E4|O�Z!�>"QHѱ�47!�-@��ɱ!���K��?�H���K.<�+�ļI�İ!�ׂSÀ��?QPʘ��R` w�?ҧW��)9э�Ss���ff^�cll��6 5�C&F7�\�/1"�V�hC��8ajyK>E��'�`�	�㉏`��Iҧ�ӌg�"���'p��"�LJ#p��H�&��/���'S.�Sz��%�HP>^q*F�^�nA.̫�	<D�@X'�*:�<�p�`&
D��c<D�[B��.��p
]'HǞ�U�(D������L��Ʀ�B�
&D�� "����L�DU\dӒ���"O�TqΏX[�A9��I"g��A��"O��HP� c ��E��~{zh��Y���aT�ܢ"Ez]��˰8�2y�ȓ>����ԗE��3�L�nX�ȓU�"�ˣ�F�q^HC5,�m@�q�ȓx��Ma�iI�wd�@@ &֫hcF��;�2�p�-G�dU��ʁ������ȓD9���ŃN�А�$͜1shP��|պ$�un*^nz�:���z�Ҁ��+򜼉qA UD���@MI,���ȓl��h�D�A�x���;U|����e�Ȇ�Lm&���0'�;9�6���v׆,ꗫX�(-�SF*Dw�A��8����Z����@�P	
:�Q��<N6e�pmB�L����s$x��u��KZ�ZuHB������C�e�I�<��jB�1�x� �+����gF�_�<	d�սN�:`sb��8=��M@O�Z�<�Tf�"$�@q���3R4���#�m�<Y2ŕ�?�A���}��3dQ�<�doD�,�"l�P/Д���&��R�<���n�>Dh0���wji���d�<A�0����U��'��l�FOf�<I��y(-��f�T�<��gÙ`�<�f�>~Ԫ�Qa!Rk�.P��o�D�<����,�;A+�'cNy@��@�<Q7�8m�i���ޞSB��7��v�<�v�4)"��`F�m��@�T�<�	@?&z,\���V��Q�G�U�<��뀋1'ax�R�i ��Hz�<Ya�ձQ�� .�h�FpP �Zv�<�rEJ�8��iH�'�2AW�}@��Lz�<i�M��<���X �P� d{�<Q��]%F\�p�gO�/YJ�Y�&r�<��Y�8ܒI�v��|�����o�<���Ć7r�M�&�6���6�~�<a�CA�\ш�g�_0�J��2�G�<��ϳ?]�pJ�������B�<�W��L�=;À�+y�Y[�.z�<�Cb��ʬ!��Bً%R�[�w�<�D�Z~$�!->sn����J�<��C�5R�l�T+��^�؝�����<�gN��Y|\G+�9/L0�R�PC�<1�H8�"Q��5"΀���a�<QH@}��I@�H4R (D�V�<9��U(#��#u�Kd����Nv�<�a,�Ă
"�ҹ�4'EW�<I��ݱu�
�b�,�M���nNw�<��]l� �@�R�38�J�<P�B]F����,|U�e{���k��p��J ��	;�Q'��!�l�FW�C0�(�I#+��%�?%?]�6��7}#L�j��!
�d8��&}ѻB�O1��	�RnV:�H�K/k��i1��d��@ �$���O�� �{J|:QE��\�]"��R/� 2s�	C���2t�)�IRa>t�9#�}�T�P��^�&S�'�p�Dy���L�#p�V�01��	P�	2�J����	�(O�>�k�<d2LY���^��x�7�k�bɘ��N8�_|Rى3���C�k��I�K{T4�bI�
�0|Pb·l(�j I��
���@��	v�
���H���ą�-�ldzrB\�/=�����E*�yB�F&'&������S5Wh�a��U�:���닦iDH��ّ�\a�C�z?)R��k⓺A���4�>A�\4&Ujy3H�G^T�q���P�AkB��1����˪5����Y���BG���ӊN("���U�a�T(��O�&�"~� �P8�H�7&iЦ'\�.C��ʑ�K#��"}0��4��B�OՊ���$L|�f,�I�޺�
ç#������XnU�L�`��]� �'�H���?�qO����"��6���+�ဗ\bȐ��S����f���S�>�g?��ܙ�E ��KN��b�*A�@6�|r�H�@ b��>��gʛp� �	���#�tt��#D����H���H4A ���7�!D��h!cɢ(y���D�d2x��?D�$�쒗��%�B�O��P��C<D�
gƛY~�{�C�r^( sS9D���l�#=�R�U!F2i��2�6D��S-II�رX	��i�y�s�9D�t��������O�"(>��BT(8D�`i�$�k��ո1�-p�,rr�6D�|����&\��� 
[�'=�PD�4D����8p���e�3'U��� %D�|��D�jK�LÃ,�561�<�a$D�����JJ�m���B?H)��&k#D���d(&N, ���4p	�P�&�"D�x��P�]NT�{�&ʝY�|$�7,!D�Ԉĩ�!f�<�'�%uy$�C^�y�{��8�֕(m�%���&�y2Ɩ�Y0�mC�#=x�tC��+�y�hW�_A�Y�/ �N�R��G��y�b'Ƅ��Y;�XPU&R �yrO�,����g��^\��D)Ӓ�y����&���@�� P�d��yR.�K�(��W��9
�������yB�ь+�8P��˔�uܜ����y��ןL�zM� �F�f� B��P>�y��NWL\x��\jNɹA��.�y���5���H RN�۵)��y��?<����ꕣ>�6��4����y��+sL�W#6�J��tΚ#�y/z)pr��lЊT�R�Z�W�j���8e��c�qTD�ed�4�lL��^�M����&�e��\:"��ȓ	Er���٤94f�8�C K�h��\�^MҢ��kf�HC
�-"����M9>�RQ��/�����-k�R ��Ftj��� =i����F)oވ��a��`�C����=�t'�.T1&�ȓ:�ڨ�4�_+r\��S��.T+���~��Is�E6tQ��iGc�$6X�\��?@�ı�MD�7�\�9��"] >5��4�t�p�c�+R�µg� t�`��FI��
��þw�j<���#x�hi��AJ��"�Ɉ\����2@TI|����M��9����Ri^�y��C�RՅȓAav12bQ(V(,��.�6{�lT�ȓ*�Z�I���f;E�.G�V�E��Ne� ����q���$���EѠ���9�)��Vnl蘤BA���ȓH:D�j/r	�E�Z (�J�ȓ/� iv+L�wG�9�I_:W�لȓr�4����A��2b�6*<��ȓy/*��Be�P^y��a�)���ȓ�����1���3���A��y�ȓ
�(҃١;�:�c�G/R���ȓ �$�%��$��Ÿ�D�O񊄇�a��P0L�-5>b���G��Z�d���}k��@T�U�,Ő��2_�Tl���e hi��ف�����Y G�D!��'�n� 
%B��u���9Bg�ͅ�S�? 2�����2>R��FX�<v����"O�]�$��
J^h� �!H�}Z�"O&8{7�Q�Z�5c��ӶM+Vu�"O^Y"g�[Ac6�yV��&!$4��"O�h �ŵ~�h�%�I/@���"O���*�B���)�癬T2Bq�$"O��02�F�"�H-p�� �"O�!��	�6�"�ig�C�k�k�"OŘĂK�:��j���g���E"O�(�I�\�h-���C.G>a�"O�Q*�� �P��q�]�1��a�"O\�2��6`[��VH�����"O@���*H�A��@37gףF���"OL�˂�ڄ��i:���eg�=��"O��+@OXK� `P�^�7b$ͩ1"ON��a���Vڸ�bu,A�w�}�"O>��&�+����\�, S"OT`1צT93��(BI�nb���"O�]JF�͚A���#@b�M�V"O&�pCR�4��qIw����HD��"O��'FASV����U�,Z���&"OdX� ��5:̪�G'N�t8z���"O��p�5q|<���fѷ˦AK�"OL�d捚 X�h���'L����"O�	Sm��IE�sM�m!�3�"Ǫ2uÓ<�ѫ;,�֨�d"OА�@�u|��Ib`=��"O��cÉ�<f����fp�;�"OB�ò�W�>�)@��;bS�"O��aAJ��9�W�r�6t��"O�ٛgV�8�n�h��a�l��"O�S��%��$�t��#��0��"Ox�1�G;I�p!���ߪԺ�"O�����$�=���L=T��&"O���� �� �d�I�O���T"Op)CE]lw�8��q��f�>�y���%g����Vk�,���0F�Ԁ�y�#ڿG�i:0k�!qa�Q'�c�<yu���#�&kD�3o:������X�<9�(��7�*i��L�d
Δ���X�<��M")Z�T�DHH�Ms��uAW�<��M�J�2!`E�:�Z��w�R�<�"$�5����,�0�"hB0CXw�<�A"|dN0r��-J<\J�AVj�<�Q*g�t]r$��N}j�h���9�y�Fd��Y��O?���`t�P��y�F�`{�\�@�*2����+��y���3*��,#�*[��l2U٘�y�!&�� ���M;��Q3����y�K�?�e��ݚ%Й*$K �yr��[}h��FM�# �a�GF"�y�+�?h�pa��O�)IfQ��Ͳ�y,��y��&A���� 6�	��y�P�ri8�p���F�
��eh��y��'����Ĉ�,�*}�u���y�ğ)J����1+߇���lJ��y�i�/P�����`ȪX�yB���y2����iŘN��9��b܈�y��b.4Ţr��-J�iEI �y"��/F�)�UC�G�h��E�3�y��?0��*�iR-9wb��d.�<�yb�]�vp��3)E5"���5�'�y"�ܴ ��'��� ����yRf��8�y�D��-¬���J��y
� �I�1�Wd,�ԡ!eƎJ��l0�"O{���`�u|
�2�ϝ2Z�ܡ�ȓPb�њa	đ MX]�$��:%b>�ȓ��p��E���KӎP8]%��ȓ{�r%#�,i�H��H[�9׺��ȓ/����� �c1H���E7.���ȓD&f  H�5H><X�#Oɰ/V`�ȓ(�$��e9s�! $h��5"�ȓ|FF��+�36'�0����'Py�8��o��H��4MT<ii�,*Tt��s=f`�Vŕ>��� �>�ń�=�,e3e]�8�F��b�� nl�P��?��1��AH7�����]k�̄�/�v�@$��eL"HK$ꟊ5��e��nB�rb������fϭp�0�ȓV��;RI��~	ĥAcT�o6���0�}�O��J�fE���B������"��6U�ByyG��MGPu�� �V`;��Ÿg]����c��΀P�ȓ��xPD�۫hh �*�?�A�ȓv��4P�&\~�p���g����ȓ�V�h����0j�rU,�;,�e��ah8�k�l�#vdzԇ;� �ȓe���*q��_A��a��?t5��ȓO����Â7d�fQ���8+�؅ȓV����
�i$�����F�^<ⵅȓ/d��B�?�x%���H-�H���o���N��]|�#��Ϭ-����T�� �3���V����D΂��݅ȓ/�P���"Y>������m��E��I�i���X%y24�E���W�N��ȓĢA86,GJ)��F��}T��2�\�U�}�|a����2�Ȅȓ&> �	 ��!
����1��M��p:����13tLB"�G.bP��e�~a���f��udb?b+@��ȓZ���	`�T�A��'��3#� ܄ȓH"�3q �Px������Y
���ȓ9�MI�KѤnRqB�!�r�p%�ȓ]�r���o�#@1"W(N�%�r���:��BF+R�wZ�IP�ߛ+pԅ�#8æ��
Ϥ�8En��V��Ʌȓ,�mM�t
	�jH	5h`�ȓ`'FQH����0�4P�&=�l\�ȓ.�PJ!���c� 8S��:��=��s��1 4���#�BF��D��rzj�
R�G$���J��T���
y��-	�&��T+���c3 ͅ�G- ��  �,��5�B��g,�-�ʓGpH����>`v��ٱ�[�@��B��4pƌ��hIm-���j%�B�	h�y"�nL�mk
�,�(l�B�	� ! ��[�%5�`�d�D�'cxB䉨��	����3Mk���#�0�&B�I$"qVe�te�5j����ã�cM*B�	�(6䑫m^=;.��n���B�Ih�t�X$)n��8�'U�B�I>���w#Z�<�!��/vFBC�ɤnJ���c�x�8�'�&z�C��| @���u[�(kqK�^�DB�=Gc��ۧ�* ���X�NdB�ZcRڞ1.|M!��C�_��C�	06��MB0$t���j��>	
�C�	'w��X��ϓA�P5[��\�g��C�)� &�`�dN�?(e&,Da�A�"O s�ʞJd��Rk`%�DE"O�Ի�I������^��8ȃ"O\+��C�_�����'!�����"O̅�D���qa\I�,�&D���@"O��;�I��U�P���$�.<��x�V"O�ܢ�K�a>�}	 �+�f�"O<,c��U�(V�Y`�Sk�ڵ�T"On�#$��%�����/�*ͩ"O4͹'.��i��l�a�ք72e��"O�u�   ���%��H��k�a���ç �\�<�2��*�L��(� �&�cg(^�<q��(4`�l\���`�e�Rx��Gx��
	N�`
a��j� ��5ㆳ��'^(�EyJ?�ІI͂X*q{ C�5,2@���'D�p���;a�h��A�&3d�ͩ3G2D����iZ27R�1��e�'����.D��(W�Ϩ��A!���(A4�IqE���`��	b}��K�kD��i��̠:�D���eգ�p=ٴ��C�:a�T�\*͂��D�CB����	�'��rF�U���j@	�[$�� �{��']�O�Oe�A��M�G�&��ӳ����'�ў�}� �0�FF'����k��W�L!��O~c�h�㉄�\���@��}2u#����k���'�a}Re�"~"��@K�J��A�W$bU����ɾ���m::MbGh �Szn�c�S�azR�D[�ux�%DYT zQBgeQ;aY!�d�>@��xt�[<0�a�I�u�����'����`F�;֢	*��E�ՂA,D���O\6���n��e��,rgJ?D��!#C��f\ک0��0JR�l��2$��SF�]"'�ZE��Y��)3cݨ�yↈ%O�BIzv�[J����ع�y�[�V�P1K�*B�%��5�&OO��y2m��p������]6 ����Eo��'+ўb>ّ0���%.E��)69MR��I6D����#�
T�^Mj��H��&���2D�p��(k�d�ree	�� 0� 3D�܈SB�#5s�#��G1sư�ٗ�2D�x,���Xf�p|�����I>����+�Yվ� 	��b�� oI*��B��+w��9�P.(�4��&p��b� E{J|:���J�i��!��/�r��W�<��]�V�L*SLU�.^-�T�S�<��E�E�̝
�B�/YY��()M�<�Ơ#q'~Pv˨V��H��
OH<���֑.�*ԀR�\U#&��S��%��{R��Y2�[g�R:�}j��	�>a{b�'(��R�k��'w[(�kÎ;) 2`���\1�cg] _�	@���3J/��G}�ŕj�O�� ���Y��A,^o�`k��d?O�4��O ,�ظO�"Z��h�u^��F{Zw5�O̔��"R�.((Ԩݭ4�93�"O�y�+�_���Z��ع"�!4T������9��xFz���7�����m� T����?��D֏&˖�G	ؐЮM�TNON�<qwo�;8T���l�O��ts��G�<a�y$��!U��#L��רM��y"�ށ)�J��K���W�Q��yBF��v��TIU)�1I_ ��!�3�?I	�'p����I�;��1�H^�d�L�+ÓJ���35�4#�SJ J(y�'O6D�8S�&O��d�$R� 	];��3?��)§8�����֫=eH��� Qf��|��&0&	#c�!j|�`��M��VV���hO�>�� &��A�D(%�"�i$"D��$�I�^�F����5�`<hu <D� �1���;�(��
Æjv���q�:D��	�j��o �H�� ��'`:4��l-D���@�7َ��4�ʒ��x�Nl�p��ɋ3����N�(W{� ��K"X���Dv�"o �A�D�[��F2F���[+yh<�c,A0 =���"���.��d�D�<Y�a%�!�ËYzպtZ7�Bx�<1��I<i�i�7@�����qx�|�'�\̀dW�E�����(�¸��'���C�]7`�r@�$�s��̓�'N�H�j�0
�fd)�kxTh��'u�s@M�4q�z���=n���'"LQh��/@�$�*ci	N y��'���)W��L�jS����W����D#�O,$��k�61��!����5@D0qr�'��D�E!�?`����%Ќ7.j�&#*D��Kr�&t��m�6!س�Z ���-D��F釋r-�XY����t�9t�%D�8R]jD�6h�@N� �	�$�0��)� 2����A ��)$)2+ �H�"O\3�ɕ�v��eqVH���;�"O���*I�N�,pڐHX�~� d�@"O���h@� w8��&�'���s�"O
	X�o�9�H����ڤ��'��Dy��)_�a�R��R��/&��a� ,,OТ<yu��2t�pie�J2+9�D�"�	X�<�O|(�G�T�]�<����LSGv�r��d`�<�>ͧO.�	�\qh-�G��~�@�a�6�j���'Ԝ��N6p���'�Ÿ}���{�\�4G{�'Y>\�ǫ�;�>p���6�@݇�#n�t��O;�A�$ь�6��=9�4�O�O��iQw�ό2���t.��4�I�'�����5Z�F�RD��4>!�PY��-O�9 !��i���)c�74a×"O�E��dƄ`��4¦�=r�ڴ*�"O�}p�ю#R�0E��i�J���"O�$��^�p��!�Ժq"H���"O�h��ЩNZ���a�/�֭�R"O�41W��)A���� �?b���z�"Ov8)��V(<M����F�!x��P��>	�$��	�׸>%|���R��p)��	Xy"m�.��ܚ��afN�z�$��y�Ǘ`
��ۂ��UK��˄K[��yr�	.��v�F�S�
YiA�2D�dC�������6��d�(�a�$D�DS���3?^lm�E-]TƐ,C@$D�,��/IVy��Kچ��3��"D���f�P+o���eM��o��<�%;D�l��[�+��A �S>��S�+#D��h׬'�J܀pi,IE����5D��0�F��A	�ϰ���7�2D�@a$̒�(Q��`�*��f����h,D�hg#�ʞ��G��N��k��*D��4Lܢ@̢-25��Eeʸ�s�&D��7-�9]䠸q'CX& �0�DA%D��૆#a�RD	���>]�V@y!"D�`����<x�ajw�W�8-�p�m>D��1��N�x��v�փ;7ꔱ(;D�d:��ڮCU�AB㇖g��<�Ҡ9D�(�UJ�1 Hp���3��#� 9D�l��'ȤP�~�!a�S�q!����9D���ϰW��()V�����r�8D��q�ŀ8���bm�	�*��c�*D�y֪��@�Y�a�I!5�2Qivf'D��P�c�|���Z&R�N�/%D���Ʀ
�@:����@�1Mbd%yF*Op���݁�8 ��]���0��"O�I��ī.�>-ȗ!��6�$YK�"O�� �O�,G ��U�]���K�"OFaa˚+"�
V�[zte��*O$�ʢ���Z���L��I�A�'vtH�AU0U��Th�� 5,cl���'�-�t�%o�~�@Q.�l���'�J��h!1N�Y���!N��S�'R�kW�̣n��(Z��O#}eJEp�'M<ƕ�B��ƛ�E���'� %u�%}"i`�Z<�"t�	�'΀� QHU8�U�4�8�	�'��TBЋA$D�
QJ$E� (�����'l=
��?N��\
$g�'�nԓ�'���Q��X-�:�`@-\��R�'n��� �1Q:���C�-n$59�'#�-C$J0_�d��2�_��d
��� �Xʆ�D�L�"-�D�q��,��? \�
�'I-0$!!ATvńȓOHX��F���n��X����Fώ��"@@���	��`K�=Ilv���c�nY��� v>�X&�Q�@����ןt�I�0�I�h�Iϟ��	ԟ���{��` ��
4xJi!VK�s����ǟ��	֟����� �	ǟ��I��	��>�s��� f�8ԀP����I�����۟�����������ӟ�	5Yg<�k�FE��r ����+�d �I쟰���<��۟��	ӟ��ߟ�	�6�!��;((�2������<�IʟD�	�������������Iǟ��Ɂ&Ⱦ|��X6{=���B��<~����ҟ��I�	��������I�����:V<���A�tV�2�J�1�F���П��	�����џl�Iʟ ��şX���	�F 3B
�1t�8�Q�|�%�	�X������	����I蟬������ɱ,:�SD��U?(yr�,_!������X�	�4��ӟ���������d���i����#AqB^��^�f�����$�	Ɵ��	�����ПT�	ݟ��	;0ӈ�8g�[ht̤��$�*鸩����������I����ܟ|�	ҟ��	+�TԚ��+�`�Aq��|�����$�Iٟ$���������������	�����*�#H����4��iʑ�����IßL������I̟$��4�?)��<$d,K�@�-�t�(�E�T��i�UR�L�	Wy���O$�m,keH���A�(R�B��7���|��f�$?I�i9�O�9O��d�0K�~����>6\�P�L�=9��D�O���wGt�����ԡ�(�O[l��F���9��r�*�=6��y�y��'�IA�O�(' |�d���_�.���1Phh���8�D6�S��M�;J��LY����"�h�ئ&>I\^أ���?��'h�)�S�pR}l��<��b��RJ̩���#c���5
Q�<I�'<�D�/�hO��O���Fhŗ�8��G�k���(U5OTʓ���FD���'Č�a�5�@���H̘J~*hjR��NJ}��'��9OV�Ũ
T,�}��ͨ`�.��<�'�bR�>��1��d+ן�1g�'$$~�ؤ�3�Ig.��2k��i%�ly"�����dT"�V��p�����F�5H��Sʦ��Q�7?Q�i��O�	�� ���'/�h����+��D�O��O��I7�m�*������ �k�mV*�.	x�@�0��`j5����4���D�O^���O�$N;'�A �R%ԕ;�\<�L�Sg�&�R��B�'�r���'�n}��(\V�%����)��yj�o�>�ݦi��d�)�Ӟ=����Q p j��!��U�|�<�"���S�O�y�N>�+ODP
pj�D褥�2fA'h�.Hz��'=�7���L��k}� U�A�e躁�!+΢����XϦ�?iP�t�I�����J���֩ߟJN5�ȕ%N�rplA~�4WX��ӭ69�O� G;&ȴyV�O�DT���,˓�y��'���'�r�'���Ƀ7|��P*�bt�	`��1"q4���O�Ҧ]a.�i��'|�yB�߆�x �rC��1|Zp:�|r�'��O��a�������<<���
Y�U�ѪG9IPT������V�&��\�������O
���O|�Ĉ,{ �����r���2K�-f�.5G��O�����=��'	�O}W�����i�D�0kӀ��j�y��'b
듥?)��O�2'3�z)�`��AnݔBA����L�:��=x�U� �Ӥ2t��D�	 |x^��f�SI� <�4&V#q�\�I���I���)r��?��Ė���@��"2%ɗ�]�Y��8Rk�/�<�'[(7m�O|��?�0[�����y,����*���`��a�t�Iԟ�
q�Tڦ���?!-V~�i��$S�t�.�`⌢a��r�#W�Ģ<����?A���?���?Y.�:H6i�"٨I�&O�kL��n֦MH������	��D$?�I��Mϻf)���&T:l-��:p���j��?AI>�|�uG�8u��Qϓ-X�xW�''ux�l��o֤��w�pB��O��N>	*O�S.pTEҕ[,(�1�r��[�F�����E������	���� ��e��'�qڂ|�v�C����ş���R�	�n�B,[�GM2|�T��snB~`��e����Z�ԈL~��I�O��R�|ٰ�P��>u��p�(R����?���?����h���ĞR���%�{~X��#d#Q6���ݦ%y���ky�OlӺ���E��]��,˷�����l��t�f��ş|�Iݟ<��f��E�*�:��Mj����L���_�R6��TE�v�<ة���
������D*�MK@kL��jB�ʍS���M��D@�?q���?���D.O�r��8�V�ǵ�k��9t���?i���S�'_����K�?P_�����8��0�M��^�옴��W{�$4��<�𠝠B0�XC��D	q���u�S7�?����?I��?�'���_�QZ���ş�*���&9�r(�f
]A���bhW�|r�4��'����?��Ӽ3��.�Bb`��>P��m���0E+|t�b.{~b���a����ӪBD�O�� : ��]�8A�N�oX&%��:O.�D�OF�d�O����O�?e�+0��H[�zCfMZ�C��X�����ݴY�l�,O��o�n�c8���!��,���s��H6�$���	����K���jP�&?�a�D�j� C*��Tn�����E'Y���1�/�O�YCM>9,O���O��$�O�� Ƅ�LU�!9%� �j5�7G�OD�ķ<t�i�hj�'���'�哚(ϫ��*P���R�:xbE*�O&��'��'rɧ��,0�tt�@�	���Q#�&ѯ?q���2	�)kn�Z��	S��~�� 87��
� �zZ.�(V�L!�v��	����	ןx�)��CyRCgӊː�B��P��*\1q�*��q�ѭ#�(�r�����]q}��'�l��߀k�č��\�{�j��a�O@�D�y?�1������0nW;1��ԟ~��� ��1�A� �l�Q����<))O��OZ��O����O>�'�Ƅ8QOѡ6B p�tiI�.��` �i�Q3�V�D�	L�S�P9���;#��7&�H����w	��jތ�?a���S�'��M��j��<Y�'m���E'X
d�Ѧ���<نa�>X,�מ����4�B�DN�|�&xr��Z�3�������I��$�OZ���O0ʓԛ�/ȔU���'D��]�\D^Aq׮ �N�ks%=r�'�R*�>!���?9L>)7}����D�7��`pA���<���4J��S�
�j-O���ø�?y��O%0��
5��k�n�ia�\:�"Od���ծF7�,˄�_,}F� ����O4�oZ6�r��	ܟ�2�4���yGd�C` LY��؃W��iF����y�'H��'[&���i��ɂ" ��a�ޟ,! �= �Z&J�S�J�a5
)�d�<I��?!��?���?I���Z�h�Y��_�=�t���9���-"D�X��t�I�(%?�I�UÔ�H��اIy��u�Ԕx��1��O����O��O1�t��� �$$��{�#��j�j�!i����9Ҕ�ЪQA��a-���s�	Syr�
?O�^,�΁7Ƕ�����0>��i�z}�$�'DTcWB�	&Ď��el��7b����' �6�8�I
����O��D�O�t�v����y����d2:A
��5b3H7�<?�)�8����s���-`�^�Ҕ:�d2 9jՓ�s���	�|�	��p�Iџ�&?���n���B�ys��$=�p��oI��)�<^���O!m��"��'��6��OZʓ	5�UJ�*� B6�Xe.�d���<Y��?��X.2q0�4�y��'j�4��[����ѢI�k{���^�x8�I*d�'��IY��.�EzRfE�W������hlHGxr.h�b�i�O0�d�O��'l���P�g�
�����Jm����'���?����S��_�yv�Ö��
p��aA�e݆S������֔Bq*�H$[�據[T�"�~��)(��\��J��pI�P�L-!����<��ɟd�)��]yIc��U0�-��!4i{PF�.�p�R�Lؤʓb���ćW}��'���Kߖ�xQ�"ˤ]�"^����	�5+́�2I:?���͋t��)3�4c�Id �Mtu�ȱE�:�y"P����ԟ���̟ ��џȔO���юB�^��a��DX"4`�D�pӪ�«�O����Op����d�ɦ�]�N����G&;����!����H��?�L>�|�6 �; `͓Oظ%��}��Y�Od�H�C��y�	n�`Q[CI�(N�T��NU�\_f%�E��?(�$i�O�U���taX���O��Wy�=��䑆z$�Wלe����g#�:�M鵄ZX6��Dy"��
,�
 �`�1M�� �ţD����˵~�<����W��R��G	�K7MP/ V���Дo����*z��#�Ȼ.�:�T�Z9Q|d��n*d�hlJ1)ܢ�@E���4F�>��6
š��}Z׍Q/}$��˷�ǥ	�x�RE)�]� -Q�r�R:@b�d� A���6��q�Ĩ��<<\9�!-v����OU�tBA&n���Ȣ1�Ĳm�Φ-�	|y��'���'WB�ZsT>�cu�UРZ����k]��7�Ҧu�	��'f��#��~����?q�'e���S�I]�B�
���֛H��ʄ�xR�'2"ˎ�E��O4�&,/δ���I�i��|�b�*Ɣ7ͥ<agL�'kP�&�'*��'D��a�>�1x~��1�	a|y�ք�6EO��n����I�(�:X�?����ɏ3x�#�-�>%�P&��+�M;��F�����'-��'�����>A)O��%藊zr�x��M]ql�A%����	�u�ߟ&�������7�(��B]��4k���Y���'U��'E���G�>�*O������D�q����q�wl���	|��Oi���x�������蟔)���;q���F�6%�hS%(��M{��W�Z���V�Ĕ'.��|ZcU��#T��K�X��a	7D҅H�O`|�$�O��$�O�˓`	�q��I�3A.l�"��h~���[7N_��Ny��'��'���'*����͞�Jzv��'�ߛBhQ�T��9�BQ���I��IEy#G
Kv�-aT���(�_����f@:~l7��<������?���,H��'���3'OǕ}���C�}�d@ȯO���O��$�<�c��V��Sş�3�!�A�`x���&^���`ߛ�Ms�����?y�||F�"����	_T����!Vt$��߽|�"7��O���<��!�/^��ԟ����?�A�	�&��QݱJ�K.�%���ݟ��ẘ���d��^�j�!�
�p��Ӆ��MK-O��Z�KHߦ�������T�姀 $Ii`�ƇwW��c$�	#pI6��A�i��'���'���$�|n�:�=�U�H�!,�i���:Q�B6m�	-�m@����L����|���ŗ]��b`J���L�@	ǝ���'}��'�R�L��y��'U� �T�؀sF��۳�"L �	�n�X���O����
 ��%��S՟��Ic�(���_�`���cWI��!�&3�4�?A����Y��V>Q��M�C*U"S�&Ip��Y+]*Dڰ�M���ɠ8^=�'w�'��'�AH�Ç�ʈ�hM�:!1��%I�1Ox�$�<��7]�HIV
Y�[�vqr(U�}��K�����O��=�	�����j�>l�A�	@��IցQ��ȹm8R����?!���?�*O(��R�A�|�'Ɨ&4�|�[2��8+�补�Z}��'m2�',�	�ORI�|��9����R���˴�ڠ.-���?����?a)O촲A�KU���vb�J@U�Q�\`��V-c�	ڴ�?�J>*O���O0�O��[��4LN���ɐ�_�2��4�?�����$,��&>��I�?ט��^�i3��p���阯 �@6M�<���?q���?�L~��CU`+[����J�1[+ԝ�æ��'�ڌS��tӨ1�O���O�N�S�0�I���*b���y�Fؼ �@nZƟ��	�����ɭ<.�����F�����냱*�^����8�M{𮛟�?���?q����(O��F0F!#֦�%� �#b���4���#�O�����)�'sĄ��T��_c6؁���!a,P�f�i�R�'<"E@�*��)�H�(	գ�B|:��e�� 1�ZIF-�O�4'>�������	�j�`�BA�"[6� �C"��,�ܴ�?�Vˁ&a���4�'��S��BA�����9+D-�4ߦ�M)O���<	���?�����dǬ�N��U�8c��ixU`G�"t�҃��|�IΟ�	S�	NyZwA(8"j�&E�1p�\��Ԃڴ�?�M>I������OzAW��?}��Cְ �:�B��n�(��j�H��O����	qy����M��N�� Șb�9 ^���ZL}��'B�'��	� .�:����d��T��N�a&�t�� Gw���l�؟d�'8��'cr)��y��>�v��&Bʰ�g��#9�4�S�����	����'%�}2D-�~
���?��'��x���rB<\0�K�&Aᰠ)�Z����ɟ�	�L�X�	����'����4+>�quB�FVd�������vU�(�o��M����?y��r�[��7e��E��	R�R �pd��B'�6�O2��A�{��DT��'�q��|��#�I��0s!�΍E��TI�icD!1�ct����O��d퟊��'�剂�HC�*��dxd��Ei�>�b$�ܴ5��̓��$�O��?��� e�����ެ-(� ��ċ�"�(#ܴ�?����?Q��M���ly��'!�Ā�4>QSC
ʌWvy*��B�����'k�	�Z}��)���?q�OJb�X�r�Ǟ���{B �9{u���'�����>�/O��$�<����5	�2�4�p�ǘ�uE�R#Z��50�	ݟ�Iܟ���Z��'��hK�1}�N�X�H�����0��%d����D�O��?����?�E��-�\p�P/��;c�@Ã�٧%9����?����?���?�(O�m�i��|����tBH�dK"����ԎZǦՕ':T�������I"0��牝���Cb�0�-���J�`z�� ش�?���?����Dڝ>�F��O>"I#�$;P.�.A猬Hv���4]�7-�O���?���?IG���<�/OB= ��� ~����!���R���������'�R��t�~���?�������dT�6P�\s�]��<8�Z���I؟���%wQ���'?�DP�r�@<f����� Z)t�L�n�Hy�ċ�L7��OV���O2��Pi}Zw��I(,��j��U�Ks(`s�4�?��Ԩ�ϓ�?!(OF�>iQ���v�ht���8(�X!�&g��x��ͦI�I������?ᣩO��!p�*� �7���cW�w�2��im8���'c�^��b� 
�{��0~�r!� �s�h��p�i�B�'�rX>�H�����O��	�-�t�U
+#&�slӱG�D6��O˓W����S�d�'�b�'��k��*_ ^ �6J�`�0uGb���ٶD$�,�I(%���&�����P+JD񭏧0+*�M�ĸ�<���?9����V�H�b�+߈CQr�f*H&S��ࠏ�j��?i.Op��O��df$|�C� 	Sg�H��k_�;�օP�b�O��?���?)(O���co��|�a��}8��]>�n��c*�B}��'�b�|��'�B�_�~�dH�Y}6T)A#�?s �6)˷(��ꓘ?a��?A-O80ɷ`A�S�a<�7�6c8���9�-�ߴ�?�K>Q��?�"+�<	J��R�[*nCX\���֩=�N�BB�oӊ�D�O�ʓ|j�q�Н���'��T�[�O.�!3F��p�P�V%��2b�xb�'�"�O��>=����e�"Ll��5;�6M�<	3���6ʪ~����g��P��Z�,H��B�*���bW�mӢ���O�$o�D"�D%�S���5�u�ЦZ�D�3̛ R�6M��%�Bn�����՟(�S��ē�?Y�N�6w4<�i��i��sƬW;)��V�_��yB�|����O������	p-�@��JԾj~z!��馩��ן��I�89:�}��'��� ��%���X�29X5	��%��ٛ�i��'Q,��$�/��O��D�Oh�xW���K$%B�ZF`]&*�ڦ�	Iئ�3M<1���?�O>��2�d�Я*gMMBdJ��O�D��'��%s��'���������'�l�9���69&��Vnc|�̙ԁ@
d�O����O�O����OX���_����&TP@�Qo܀��d�<��?�����@
4� �'n�����A2�X����}2�$����e�I럈�'w}��ɣ?���&��/Ԇ�҂oǱ;M�ۨO0���O���<����+Y�O��y��A� 7F���GB�[����}����*�$�O������J��<}P$>� @M�6wU��0� ϟ�Mk���?�.O��,�$>��	�?�%�*O��*�],�i;2���ē�?���c��[������EG�J���L,�q���\�Mc*O�,�O�Ϧ�Ю�V�d�4��'Wj ��Q���P�� ;r��4�?���>��i������O��\�#�L!q�^T����kc
"�4T���y�i���'��O��c�D��Z t>̈2һP�xP6!��MK����?QO>���'4�IJqIQ7!��bԊ��ujΔp�d�l���OX�DF�4��>���~�b�n?��y��\@l,�چό�M�K>�T�Җ5�O\��'t��Y#�Ӌ�,)�Όp���K�$6M�OJ�q7�
Y�i>�Gy��rM����Q������?Y(O����O��D�<A�'�1C��U���O�(9����T�*s3�x��'dў��hHXu!REZ�7�,e��H�4x5��o�埔�'K��'�B�'�"�K�����uB|��6�R�<�Z����Dݛ��'���'A�'��Q�!�t������;>��1"�,�l)At]�����X�IbyB�V�F,��b5��Ĝ��S��I�$�X�j1G��	ٟ4�?qf�O�'d(<(r�b��&Z؄����!$�o���X�I۟����$1Pp������I�����Epm[ x�J��ќ8>ܱ�M<����d�����!Dc6$э�z�&ZEFW�)�N��?s&���?���?��������d�J�hrh�S��)sաQ�M�����Fqr����e+F�Ә�b*k02y�f�iе�5z�����O��$���L'�\�	,[s��`-ƫ �:�UnB�d�����?Q�,��p���������J��`��&�'��'� 䊓C7�	�����q>��ǪGE�Q��EA�>��Ն������x��g"$,Xl�!͑�#enѺF��Mc��Y%�=2E�x��'�R�|Zcy�0kd���w�.p	S�_M
@��O�쒦�$�O,���O��"��(&��A�T!��"����J����'-��'-�',��'�BH�QAؑ4%�$[�AĘh�F@rt�L+��']��cׁ,�2�HCӮ;iv��'��b4�	�ݔ<f�0e�!2�:Q�ɲ	)�щ!��~<��@��>:gp:�%��O.�5hʢx1\� "8��ǮUX�*
n�C���X�a9��G�/��\a�a�;z��0(ի�*}�(���_���B&Ԯ2ݜ���'2�9P%����]��J�<$ |K��П{H
՛Ђ�=�L��2��{�ʌȴ�� �]A��V/��y�/΍B١�ҙaK�MS��M����G��� t,��h�!�	?(�|}�e��+oY�����Ρ�D���ϟ�rdCԢi����SKM���)j�E��?�Oc$۴�J�,��v�Ե%ݶ�H�̲`�[�\kd�
��@�R�
��eǋ#����M?��W P&,$���¯�p|Q�!}2ə��?i��h������0�p��%�5S,4a*b��,!�D� X�r5�t͟	2d�8�GaxbD>�74�q�%nU� {�<��C�?�D{C[�X��䟬�����T���ID��ޟ��=,�J� 楎�GG�U�7EȲS��e�W?��(6D![��>�3��ם$��4�H��FĹS_�[q�EH#�Ř��$���d���L>	�/�' ��E�a�]�4Shq`����?��O������d�I#s�:A�� ֽ5�d���w�C�	�{�0�sc���I����!���P� l���'��D�/4���$�T>
��}k���E#
<���,2j���O����O���;�?i�����B(�8�P�*N�aS�H(��(hw���?�Nm��2lO.��6�]��*؃ 'g�ŋ���*z��
pl��.����!T�8�E��3��+���L�-HD�O.�d,ړ��'9�e��C	9kV%3!��x3z�K�'xT�䍀!�1�'�� ��y�ȥ>!(O��v�k}"�'��3�ju-b�{G ��tW4����'�R�ńwr�'��i�O���y��?R&�-��2��#ElQ�G��d�T9���	%r��}C����C���'�lx�E�ߝM4���a
�'c{XU�
�|t6M�	�$�'"jmS��&+v}�d�[�Љ�y��'��H�mT�U�`m8u�TV�>���'^z7-fJ-��B�8�\�Z!+8i��<�5@
+`�Iꟼ�O������G\6�t��c�~a k%͂�i�b�'-6DA��ݪF����	_}*���'2u�W�Z(.$��K�Ʉ�B,X��O�zbI�02S@�z�π 6����	O�$4{G����LsQ�>QƎ���h�IJ�O�I;+iڵ�#燵�)��[�y���#�X31�����/�0<�鉾�L*�D��(������Y���ҭOT���O�p9�DM�����O ���O�n�3)`&�j�i�3�H�.� v4��@������c�t�XA'�3��'���7�ݘO��`�
M���ٲ�_, ]��=y�!�W��|"�y����0��dL�!���m��7Mwy�!�?�'����DL`p�9�nD}*��"���yRT=��Q$�� Mi��	��D��'E*���D�*�$S��k3�q�$ۢ����`��i
���O��D�OF �;�?�������h�|ՈQ�˿E������?!(L�E+ڔ�l4r(Ô�0=��G/GҺq��KQ�HU�d�i�W$�Xs�kX�����CCk�����2cG���V�G�b<��F$kW��D�x�4��'�b?���'..���l����pk�E,D��8�K�}�R�ېBҳNh�d�0�	����<aaO��c�&�'B+_{~\Đ�ɦH��"d`�����'����4�'�:��x�D�'��'�*Y�cN�y5l�3�
9}���>E�?٥.��scFd��\�:@=�%�m8��9���O(�Of�`�A�9�4a�'�Z+M�I��"O�t)d�J%J ��K��׳i>a�O�n�?"�~���N�9+F8���yX>b�t2O�*�M���?�.��y���O������"�R4�7!�T��#��O��$��Mz�D1�|�'�@p@�D/Vq\4)P�C�a~"��O���&8�S�'-f���u#��)}>)�"�W����>}�g�"�?��y����$Ĩ�����L_yc�,W��y�ћ�F���=Hܢ�Y�
X��0<���ɗdT�	0H�#t��PΗ�6�BxA�4�?9��?ф�U�?I֩����?��?ͻ7�%�ӎ��M����0NгW_Z�q�yB�ݨ��<����q��ڡd#D���Cց�_ܓz&���I� W*}�##�]��e`�b�T�<!%����L>1��A<�1qcLVZ�HE�R�<�A��&>�L��"��`8���E~Ҫ!�S�O���`�fӖ%��	00<�PԠ��L4�Z��'R�'��Fsݑ��ǟ�'1o&E�tk�%BH�����;��ǫ_m<����n�p�)���7���k��J�q��!��m�pH*�!��v�� i�$,�<� n�埌��	 +�zQ���6n~̠sPI��LX�B�I�*�XՄϰit����11�db��}r� �,�7��O\�� K��	hqn�*�Z�B�
�34�$�O�1e��O��D>���ON�O����I�68̽�'�����&�'�P�b�X!�d�8�-A7G�ʨ ���-�p<�a���$&����5�X8r�78�e��h5D��[D"�/��|`t � 'J�1�>�H�۴>�8L!�ϏPѮ-)L�/p3nM�<�`蓮p2�f�'�Y>�d�ݟ�auF��)i�H�Łˍ@��T�KUߟ��� xs`L�	e�S��O���G�K�,��D�h����>a��EP���O^�-�B#M=d���b(D��9��ɳ=_��:�)���M�"$������X`��ʽ4<B�	��h%�'���H؂��S���F������B�'�.u@�K��(�1��h߬L���̲>q��?�0�)E��!����?Q���?�; @��˜9�F�FJL�4@Rb�E&y�I��Nk��xa@�U?��|b%U56�Pia�&�4�Z�22W�N9��+�,.�l�e4xQ����|r��9Y6�t�w�D�w�p��H�)�"����W�O�i�O��P�t!Łp|K&)�JdQs-D� ��F#h�H8��MѦP����`*?���)
-O�Q��Z3<�P��@]]��}j�A@:2�1yd-�O����O$������?1�O��x�wąB����&�ط ־�c� ʛ�x�ɞdc��c5 @�d�)���eS��k�'d��[B�͉+tS�	A/3�2����¢�?�
�@�����cH@�Hb@͆ �@Ņ�k4�0���4=�����P�y%��<Y`�K�4��'���"Y�.�2fE�D<�m��8"�'#D�S��'�R6��i���I&���Q"��ē���i�zTYu$[�x�*<
�Z,�p<qc#�Z�����
�X�dʣ@���I� ��R]�*R�-b���C<R�'z�)� b� P
h��snÌT��X����O����(��A��&p�P��M͡q�!�AצIDEF$y���c�Z�z'��� oo� �'q���Q�c�2�d�OB�'j����A��]h��&*�쉩�+G��TA���?!�/���?y�y*����[��$��GG���`x�aH-<��'n������)�� ��4�S=!/j$80�;;�yF^���H�S�'TG�Ի�I>TZT��0���ȓ6�dn��~�<�׷x�l��	��HO��ť��0(����r^��p+N����П��I${���hC�Ο<����i���,�*G�d�3f�^	,Tt8��@̓5���$�O~D��Ll�<PQ�eɚt�qO.,I	�	W~�hG�e��� �֪�������ҭUm����?��9��G��"����l��y��'�D��p�����ɂ"� Z���OʸDzʟVʓA�|��ԇ��a����*0�̥J4��\��	���?����?�ķ����O��)4^\"Cɢȴ��s�A�`�c)�@[�a�`FС���y�4�Y�i�a��B�	b��'�E�ʝ��ӣA�����h�O����J�8�
�`B�AvTԈ'HȹC}!�D�66@r��ղSU�Ȃ��z1OM�>y��^�B���Ο@1�I�.�84��.˹"�ބsd΋ş��I�y���I���ͧ����'��R��ώs�R��VMW:H��Q)M�:H���#�p<�У'��h���I2P�����k;00h�Ԧ~S|���&@� W���D�|?A������d�0%��(K�_��x�6�V�X]1O����dA~�9��_�H��Y@�D(W!��j�DK.8��з�z��[�\9�ĵ<D���o����'�b[>9�$�՟X��bʻj��Ā�!�kҠ(aT$�Ɵ<�I	o��uK�R�S��O�y�f��3C$t[��ȠW�����>��!I�w���?�
���o:���f�
0��� "}���<�?����䧔�'?]�SU�IZֹS��(q�<1����<���J���F`W��`��$+]}� ȏ�Ø��X�5�N*4�*1r� �V�:��'��'IXiyG��ND"�'����y瀈�O�����gٍ|��U:�_-z`D��6+S$y6\Y�D�^�v$m���i�~�dC�fߨ��$d���7Ā@��j�)����K�N�����y'��f�D
%��})�(D%Yx4CR�E(���*?Q��Hß�q�'^��i��)�|���ĩ$��0�'���Apˈ�����q��f�����O�Dzʟ˓S�n�+Q���"4�Eo�06z�)
A�,>�v�p���?����?!A�����O��Ӕ5�$��`�@�>m0 ��O��t@�
O`��$�U���q�F� 4Ҩ�r`f��PxR���xZmR+N�	td��4B�*pJ����?�H>������~�e��4�M'k��-PЊ�N�F�<�ਜ਼
(:��3Z-&�!��|̓%��IIyb�PZI�7-�O��ّ@�ʽ�$2D����W,����OR ����O�$}>�aV��O��O��p�kz4�W���3�TW	q8��e�-�I!�X���g��2R�(ԺN���G�1��|���t�l���
�	��yr�N�>�b0��sK�#`N���x�q�H�ZbZO7��	���$��(w��E�*���'�bV>y��^꟰q�IW�PR�(4#ڊT:D�[؟��I�c\|I�f�:�hapԭZ��?�O哋!�VtPE���]�So�D$��'u���ES3����2��Xv�>���S�9�86	�mJ*@dk$}�?Y��i�l#}"�'CAB����F�J��`9橛b����'�v���	�Ԥ�E�6b����������ķA\26�����:~��F�'i��';be���@��B�'x��'��#,��Y[�߷[�t���'�4�<��~x��ST��&2����&j�t����1�ɛb����_(c��IP'*T�J��D���w��c���D�Oq��'K�a�1JJ6z*f�0w*�Z�ȸ�'^Z"&נz�����-�i0�O@�Ez���Ƽm����"�Ch�Ia�A�&e�D� J:B-
���O�lZ؟ ����a>U�Sm��rҔ�"�J9=C��2A�Hu��2�O��+��0
��(!U� \l��0\lE���(�h#t�('� ܰ�m�ş��IΟ���ay��')�O� F��� ^?UN��4]�Y��@�"O�S�D�	3�i�F�i��AAA�~}W��[��ÿ�Ms���? �Bj�9�����`��q��鞵�?!��9jt�R���?�OSH������B(<�y����P�$�Kv#�PH���	�-���H�ViB��tE�����A�K,Ot��U�'n�'�z��A$� �N-
G䀖��Y
�':az��[�9���6���>��	�'��6-�{�������#
��Th��)�1O�I��E�	�I�� �OH�4�'"�ܚ�b�#9���`X�P����'ObI��mi�T>�O����c�'=�L+�jٶ7]F��OF���)��3 �`�����U�8mvB���&�'��q������O�:�Zg����=��o�SRF�'�6���E�~�����I��<��HiÓё�� ��3��� b�P�h8#�,D��!���_�z�8cՈx��S�0D���"�[���Qoئ�rUz<D���%6-o m��LL �J��-;D�겎M�[�\�#U�y� LӇ#$D�tٴ�R�#�)S�Q�U@���#D�4#׍ȻA.ni(�@�4 �����L D�\"g�ř6l�����ƠL�-(�G>D��Y�gG0��$B@_�l�����0D��*��v$�3r�^�.��� w�/D������O��Ix�5Kn�kWJ,D��K@a�"c}~��V�9)jD*�d)D���A���|3"�8I�b�xi'D�`C�G݌[GL�i�HU�
�L|�t%D�0����	u�J�ؐ���f�H��M(D��rk�&��yp�Z�h�@��&D�tTB�rGء@ę�IR~���#D��
�.k��u���$�|$�a
!D�p"�l�$:φ��Ud��!l�t�c�?D�$3���4L�H�
�b�l�8q�>D�Dy'��#�X�^���awm2D�\����A�*�W!��'"�iR�*D��'ͩuŞ��ӈ�l�ֈ2��%D�H����z���2�ْ@�h�*)D���v �0i��B⍖�1�Rjr�'D��+5�sĞ�@V5&="a0�8D��5�K�L���=3߮�P�6D�T�R�ĪTe����Q��@Y��6D�0��f��)��	��ʑ�@98	�c-4��A���#������'���$�<m�:�B��Z�D�00�I��<��C$[�D8E�#ct|��,�\�'Pz�����E��B��rx�!9�O$,XP
f�������?�W��W.�:<8�Ņ�#y�i ��OmDr��§ӣ3�\i8��'�B�8�!�I�z���B�(>��� ���%�)�'y`�}B"�µE��%����f}4ݐN�d�ax�'�-LTp4����	�3��|�Q��в;6N�I��?}�`GA�'��%q�G�Q�0LkG�
�"~��9�FǗl��q�P�$�,\$U�4�j,����@;]���<�TD��N#,���H?r��!ȡ@�v�'Z6S`��(K?0=և�:�r)�'�B�x�H�/���3�28�P���'ԮG
Ġ��9}3\!���O����OW���+��NbDɜj���y�^=��h���h�rAO�g��E}��eh�a�Ft��iZ�a� #!���6�(O�>�kT���`V��	%U������zHb�1!L�8���4�J1�r_ɼ�B�L>X۴%�D�V�N80�F��@=��=�ÆܪcfB���-a�������'��T[F��G<� �DE�w����I� 	���{J�|8a�ڥJ�\�3��*<O�}:e�ʅ
9\�1���0Hhd�ՠ­(���ȇ�"k: ��ɭ>�3Vtl[�	���2�hT�Ft�'�BY��/� u��#�ʒ��<T)��D��j�����O����{���*GnR�b'�*O��I0A��3X��p��OT���|�9K0C'	� ���U�$ք�6/��D�tp�� �	/�\tiD��օ�2'e�=�iX�:
`�VF�V Ś4a2��!eN�*��B�]�* ����P����2mH(����O�;2T��q b�ɱm*?q��ȴ(b��īK�*1�Ą�Wy"����'��$�/�i`��;LĦ� ���R)1���i�I�o���q#�I	o�1���v��Ba:w�ax���N�����)Z�O� " g����I��?@�6)+�����G6�>��JqΕ}j��R�+�:A/����@�Tg�}�Hc�7��UE:�`9Lp���13*ISQ��@��� �?��?��?q���>��������ѐ���	��b���'��`��dD��Sm�K�`,¢��E�8c�h#�O�����F�=�,ԁ� �O��'@���gAy���ip,V�9�^�9�'Zɹ��FGbԛW��C������%���k@��<�l�S��*�SV��F�h���F!11>���(O��Ҁ1�pm���ӑ$�:p�%
)��'\h��G�������R��=���ȆG�:�bh�C�/;R���'�p�Ey���)޼��?��,H��;n
L�3G��y��]���ޢ\a����O�
M�7O��S��&l��!
�����`&��Y�$ߥ��	�O��Ez� Ҟy�zIإ
)Y�8��D��'�����EQ�}s���C62-���?�I��9RP��X0:@�"�̃f�����*���D|�4nB�=jңX,D��[��7�Xi�� P�
sFX�1���8W����Qìp焴��w-�O�h�cL8Z�)����:?-�(2��H���'
L! Va�]`h�x���v�C�b��d�[�A*V�V+"F��1� ֹȖp��0�I/$�8��?���$`R B�W	6T$�*�$�=��M "�4�z�b���7M;�'�xaÖ条g켪���$J�� U�,���u��˟L��Rkoy����a�\ m���f� �Dy��K�Q���~��+�>Q����_�iB@h�0�[�m�F�~р���O�)�@���l>x� ��u����aM]ش`d��w�dӺ�O�Q7v�X�� Ns$Mj���`�ʍ�P.�$e�*�
�D�ğ��̈Le�IP2��@�뮉��hO��c�Γ!��
ާ^�>���|�2O>��$� z��=�!�1O�����އd��D2`��b��X�f���|J�?LO,U��w�- ��̽:�L�ޞv%�KƎ�"0��ݩ������k�2ݟ02����`i�m�X7�<B���iĆ����Q���q��1D��]i��
p�~�ᇮZ
�>A�`˵&�0���׬Q�~騡��џh���V$M�+E�&Ww��+$��?�A9S�mpI>��O�!�S@�;fn4]�R�O���k�(>m~���Ȏ�Z��N#��D{j0���hO��"2P�[����/˸2qx�{�V�l�ɽ(����q�:9?����7�s����p,�+My���g�0X�0��P�ϛMG��А�?O`���"S��svƄ-Պ r, uΤ	���,g�`M�V��!bGb��2q��p�����d�R`�E�'o�?n��5eˌB7�����	pC"�3�Q���aN���ä��<O
ꡯ�RU�@�m�Q��� �^z�Z���JT��
U���C�9{�����ꈳY�Ь�Q�ig��j����cNf4@�jV�X��D�YPb���v���=�ܐSu�қi�%�թ�O���O8�I��C)pS����'��y��ٍzF� S@&�=�̤h������� 6����?QD.�}e̥j_�M#c�QcG@�!E͆�3�J:�F!�� ��<yc�_��y���3��5��nX"s�jћBa�5��'�(���u�TT%?��XH`�NA�:H]�P�R���Dz"��+�$�y�(\=d�Q*��Z	���!p�:����@.�$�+�!X0+n æ�HNe�OVݤO�U���� ����mA�iU�O?��17,Ҥ'�*6��mh<����0uf�D��LM%���� S4A�$!��Y�Z�%�Ĥ�O0D�O��IB�Y"�����'�d��w��] �-`�@ v��r�AV�=w����C�����t{,�a�'�I��.ծW��AA1�>&���K��Q=~kR�D|�b�h���X��q,3Go�Y dJJ�к �1`0�DZ�VP�!ʱ`�2�>���� ��a���#]�u�Uf]o�'=b!�'�$q���X7!�n�[�'K:T#&�?D|���]�=H	���S"�>���A�e~bS>��$��MoB��EB�?e�&��U�<���5pp4⢋�O�i[���#lL`�In:(d��>��n~bE�8H�P;U��N�|�s0h=�?�����갪���G&ѡdM�l*S�%�	@'>�ˡ$G7x]µ+�è��a pꃞ\�ru�'#f����x�M	]�F���W2@��ñV��yK�玧@x�1�+S t�8iA玗4��y�����ywo
�	��m�p
��r�f�y�A�9C����4��6� �j3�i>�;c��6\�V���O�ӄ�vA����NwB	i�cT�x�8DD��B��ɈPy�P�j�&�����!����u+
�=g��c�P[��aX��x~_?A&��7���w�\^�E8�>q`2�<s�ԋF�r�d���I�4-���'�?�7OY�(� �MҠl���)��3hP��pN�8<v< �	�B��0���#���g��,%��g�;�L�t��Y��B���vF�x��,�p�!�� 4�H kc,��{L�p�	��M�|ڱ�۰"�$�S׈��t�Z5�a$�'"�)FAR5X(H��'i�q���T���b˕�F	
`���^:gj�}BA!��?i������R>Sl���?)É��g2�qYt��Qk���,A<)ǁ��C�0�MP�VӶ��h�M�
8���zQb���uk1e� ]�\� ��?�J�-'E~ٰUj҇j��=a�3O�9+�Ö�>U����Gp$ؒ� �(����E�e�SOƓR?��ҕ�'o��)UlI&xud=+�L��)�*��O�I� �gް �ˏ7[�h	�A�>aEF�?/6h����I�d����;��Y� ��BI�w¥7�@)x�hѫ6C	����u/L:1�
���I�1),�j�B��$���B/�Lc�$���R1oJ���&_ �D��|2��O�<I��胪f�dJ�	)H���'<H�U�B�~� �ފZ�(�a��is�6m�?t�������J��{��?7��b;�T��mSN������P��t����'
q�GWo�pŎ�igL�MA<0�k��vMjAS�|?	�葡[T�iVb>��.�F��R��%��nޡ�9� ٦}����'�"�q�PR��|�Ɇ=e��)qH�����#�T�d��m�o=x	0��O:N��BaA���=�'Y�)��Xp'դ7��h�W��x̓w �i��<␤�V�ܠE�RL��M����D��!�� +2��	<-~C���CD�:��Z�nHK�䕉>��M�dM�O���eN��T�^���#̤
V$�I�fh'?�8���Fw@����[�xaDؕ,�����&V?��x��	g
��t�:���:.� `S�8]n�AS�-N���i vU�`����|F|҈A!hJP棑7���@���~RJ�_4�S�:[�(�� I��s��2�Lßl�p�J:+��P�яP�g�<���ٶOw������ڰ>��N!�x�"[�C�\��z5��O�ĉ4l��<��^U*x�&K\��:���gV�#�\�VF_++K܉��'n�퉐�?|� ��DL������h�j۴#َ�)�ЈB�ҙ��
�����RP�*`'����D��,� �X�B-7 .QSL��4�<��d  Y+2A��Ѕ@�
�P����� ��j�\|�8���I�
�"4	Чhö����'��q� �P |�24��9��d#D~��Ѭ�*e�E�Ӆ/��G�a�HԢB�=�\�na���0������K�^�a ��v<m�ƣݸ8u\� ���][(<cC��/�ڌ�W�%�O�a3����s���`�J�A�a�)�G,��M3$m�P���L�O�x&>��w���^(�Pƌ��,�
f��p?9G��vİPb�DIu�8�0fhR�Sv� �ԭ%6DQE��CƦe:g�x���L�p�0�����"8)�O�3f%�dō,E�`���<aǈ��`�%Wr�(��F[#��4�V�J$ry4�#7�7o|Pxr�>1Cf�//^,�����YJP�@&�F��8�.���	Đ�pcCG%`��ئO��aƇ�* r4�ĵ`0<0�&��[�l� $O3��\
�0eY��2�ժV��@���C�R��	Q�-�1\�h��'�l�إ�H�����v�#��޼=�L�������C��"��֬�̩�>�ݚI��Q	�"��-B��.t�*C�ɦd��c���n�@Ys�Ťu-`z`�B+|��<���A�����	kZ%��(�>sVu",RzC��+��Z)q���&�-O�-���ݕ+%� f�v��	�`C��0n��v��'�A1uJG�?	G�,7| ! 4't�bK�N�'j�m�����vNp��Y&�ȂI����)F2L�Kݔ7�1sЦ�)��� L������U�D��$�ڊr�@�{w/��o*p[��'	�T4��V����Mʜdz��^�s*(c��;O\�� �Xd�'����2�ҭ��Hx��`��T�PQG
O�I��m�_|��:%͚;�ڬ���
Tf�Dx���X?�AqZ�u���[c�5�~b^�KPd8���D�m������а<1�a΋���8).�2uC��.�{C,�Tn����O4�+���wD��C�� �0q�I �l���ı% �W���	&��䓂RGf���ON%7f&��PP#b�bDj�M_	�` u�S-jX��f!V�F]���� 9,��qSq��N�- ��*���,X�I#�)��Q�����V0|���`f�)N.�C�Ɋ9�,��1i_()h�S�*�����=I�O�ر��'o`*V��'>mª�����
�'�tP6M$b��p����l\��6,I'%S�A���=!�@	�͆�;ϖTS��M1���Ė�{O�c��;���o읣�$��%~0h�7D�8س�/d�lQE��:>�6+9D��"r)�ɨvET5�6�F�7D�$a��M�t�(R���8 �,�A(D��Pd�����̲:��aB�8D�(Ю��mG�Hsu(�:�٠�,D�@;�N3��\�'A�!��{� 8D�x�1%Q�&@�4+2Z�+���jm5D�L
փI��(��K̪D���c�3D�|YC̾Kw輹C��R궱�7D�8Ctkz,���
.�@	�� 6D�L#6V�P����2V5*�`�#2D�t���<'�α`""��dm�%qGh0D�� �i(�Ŏ@�r��2����8��"O.���Bĳ]|�pJE�I߶�"O��ge�:}�����4SĜ5�"O�x�Wf�5tx c
��_TNC�"O^�9tLr�I��nɍuk�B"O=z�l� O�@�,Q~���Y�"O��qd#���(M(���$p��uZ�"OB ��
��b�u��	�(���"Ob��^�i��b�ׁ%ʥ��"O�а���ְ���A�a8� �"O��愝&lnxa�́>��� "O��H�(%�q:$�]&9��7"O�Há�^-	��H��ݺc�.��"O~�2�ŚeV�0�� �v�j�"O�˧CW�za�Q� �͒�%D�T��#V���9q!���HF*DH�j(D��c��	�"9��、='p �B�!D�tv���&X���-_���c4D�Ȳ��[o�>��6�D�y���E�1D����"t�壵急VE �w:D�܂KצB� �Ġُh=���c�:D��1@���;��h��X�u^H�둨9D�hSe�N�O �T��DW�*�y���7D���tL�{�:��)��	��"D��	��Nl�����X*�Ua�L#D����)�SH"�b��ޡ�n�q6`!D���C#�U��,
��� d~�� # D���ՠ@+�̹K"��	�P�( �>D�d�W�I�F	`H�A�"<PH$R�f!D�<�AW
FX]��eS�xkx8c�<D��Q��Ţ.	b�����4	߂%�Qe%D�t�fd�[��ɚdȐ>��p�$D�(�D�G�I�>�ɁkN&��U�� $D� XA)�R*$��GA�(+�0�@� D�08Sf��?]v�br��$���!�
#D�4+��_2 
����:y����=D��b�'ډ~N��CVm� v|d���:D�8���0�]J�]�3�c�!���+")�u�Ѭ�Je*АE`:�!��SC����#�Q���z�.P��!�$@�i�5yo�w� �$L_6�!�$N�Z�*@ �� ����$�{�!���l����.V��uhp�>Y�!�d7SԞ@3%S<�d���&
>:"!�M�i�eی?D�%Rˑb�!�Em�e����	*���Ū� !�OQ��׃� �=zI��V!��:,��<0ƪ�-�� ��;ء��@1��#H
5� ��1JL/l(^B�	�JYJ�k�հ"�Ha��K�*B�I'��@ජ�/}VdS�e�n��C�?k��d.�<$&:�CĎ�U��C�IF�����A���)��C�	��Ė�A�FIHE�ϋI�p
�"OI3F�^2G9La�� x�p�e�'�ў"~"�Ӕ�8V�� hY�G ttB�Ia�>�𱄐b��k���-igf��$h�9q���U��`����g�yҌ�8_WB ��C�%w'δY�@��yr��1�aO���TEO��Px��i�$51�P�H<���r�]�a�.���'4"Mba�A�F>�)�*Y�,�:��2�S���J�Fl ��.���,�����)�y���K��cC'EA����"��P���π ���e���i�X8��A�X�$�a�"O��Ʃ_�c� �d�H���ב|R�'��}���ٳp]:���%Z�@,i��'kN�h��ܸv�e�v
ȳI�ڜ'yў"~*pEZ7�F� �dQ.)����N�<�Fԓ)�@:p�Q�Q�%����s�<�AH�0JJ�s�)\�L���R�HF{��i�#Ŋ}��i)H�.I��m�C�$s�F�2��H+�5�7�Ԙ�C�I�)�V�7�ܝR��D��:�8C�	�OZF��ǭ� 7�2p9%�@4xL2C�	�Z�"L��-	�\B
�9�+��I�0��hO�>U�%�"@��0;���d�T$#d�3D�Z�޺4� �͜�Gd<��2o1��6�O�q)��ÍE����� ?~`bh{0"O~勔MM�{: ����ގ,W�q��'E��X怅)@(�/�ًu�L�y�!�dܵg��k�eХ/�����+g!����ykq/D�jsc�;wR�F{ʟ0Y:��ա'�.���៛V��"O$�R/��$k�D-'���8Z�<���'��9i��׼O�dkF냩Vt�����$\�%�h���ű)'~���D�/&!��=v��@��+q
i�$$�8G!�%B,�;�E�8
<�.	��U`�'��|XB���)#E	�E��>Tp�'����#�l� �[�`M����'ȼ�S0��l���1�" �zX�B�'5��tה*%~ŉ�SHX��'�5"bٿ+�+�usTUk�'+$R�B6NNȀ�,�>|l�	�'�J	��V2� ��-�j(B
�'�y�E*ˢPl�!�J<� ��'5r\�@��2Kezy�P$P#����'��	�jM/Q��Q��3�6Ѐ�'{H��Z7�.��S  =(
މ��'vt�`TMNX�t� ئT6�H��'f��1�(�P4���R�U:�������OOe��M�b!R�M%�H��gh�Т�-h��UB6�T-r7�,�ȓuxPb�/��!F��+iݖ`��hC�P+�R"���פb�>F{��'�a�E��v�����R;/���2�'�����*S�#��%YUI�"W�Uq�'(.lkV�T�`��]���!u*�Qx���'J�(#!X�F_Z��c	��*kh�	�'\�q�جE+^iqs���)���')���ƿ{�34bPB�6)C≝F8���a��d�z��j�n٠B�	? �~)XV枎K�N���PS�B�I�C��Bd� T@�FR$V�C�I8tĨd�׋M:]��)ϓ��B䉀/�}�A"��	��*��B�	:fjyHw���/��$�a˚s�P#?�����T���pF��+T≡�2�!���,'[�H��ː�N;�0�p�O 	�!�#(�ؤ�s��'9X:��	0K!�d�O��� ���R�|0:�)�H���[��'`ў �q��/I�$4ʱ.M$za�2&�OP�	�$��cr�I*\���yU�@ bB䉝@�45���*2 �Fcɛxd.B�4C����tg@�o��&��'�C�_@�,�T/�9X���w�NX&�C�?*LD]�Vxx`�K�\��B�)� :h��/� j8&�s��',N&�+E"O e	q@̂Q���	��y9Tq�B"O.�Q�ʝ
M&DNH {e"O�@�Pc	�(�M�'jStE�D"O�d���2w,P(h�ڵ|�:(��"OU���+8��jv�T�u@\� �"O���Ǫ�9bq���2�4 $Z�"O��Ƃ)(�a�B+�� ��rR"OhY1� B6���k��,@��"O��2t[6?T6���U��k�"OP��u�J/Yv��$�Q6�&�8�"O8) 7��*E_�� �q�T��"OXe)Rhޟ>V���L>B�ȼ��"O�[R	���%�Ǝ[Ep�uk�'
2Hɠ�5f�$��3c�)B�8��'�T%��[g���b�ʞ'�d���'uf8�b�V�I2��Z���좍}��)�)<5��m`e�ʹ71��bW#]1�!�$6�\���j\�t��A�Uc���!� �G0"E�rl~�yC��ŝ3�a}��>�Uē�>xF��+��ET�]�Ga	b�<yG�l<\�S)B��H��VJH�<sg^�.����1�ér?P�A��Sk�<!��ʰFXus���+&Y6�AD�R?����S�dR>���됷J/�(a��޶o�fB��+N���srJ5 <��AE^�(B�	�XH<�	���P�(a�ri�iT�C�	, ��4�T
ɾh���"q"��#��C�-�����c��c;�5�C�0K�jB�	�H�ểW&6H�5��DR�.>$C�����+�&�3y�jek �Q.p�B���@a1F%�24c(M�B�O�8!�B�I�<���I &��TՀ����B�I�i�,!�D�i	,U�g*�1{��C�ɿ6�����R�*��#��o�!�Đ����˰nVdӰY��ˋ�����	�T~�u�2+]"92T�&۳z
6B�	�~H�J�	M.x�VP��ډvhC�ɓ"�j�����bxhd��r'�C�I�nI��x2�^�-�L��F#w�C�ɛ���0tkW9���H`����C�8sJP��U@rFv�Aa��!� B�	�j�.�`�Ȧqe��ŝ���C�	����B�� )����[�O[�C�I!,D>tV�E+
�n�����C�I4�2p2%��9 9B�c̽��C�ɶ0�1	�	ȝ=k�HvA�� C��J%�#��7:�A�����i5 C䉪bVNh�#��c��M۰�ߏZ��B�I�&4ѣ���)z�h��S� :�B�	�h^h#R2&q2e� H\p�C�I�lZ@�҆�qD��׫� J��C�	�IYz��-�(�LӅ㗳FX�B�	#�����jJ ll���-��+��B�	%h&��(��̋#��E�c�V3=$2B�	�PҎ��i�fε��ּme&B�	��>���,�P�|}ؕb o"B�I���)c��*�N��b��V;B�ɜi�0�� l�:�`��^VC�q�8H���:hY���,F�B��*uV�1I��.b���+�Ç��C�I�&I*xP�ҏu^찰&f'��C�ɌK �qR��6B�̨�g�^�JψC�	"D:���be�5!��8�C�9M�B�)� JD��O�={&��u��X,*���"O��+��ϣ	m�!a��FrF۔"O�e8Ĉ[4��eJ���*>g���"O��!-C7D@ �+�t0�"O�� B��mQ����
�} ��"O� ��m�TY��2�+�!0\�a5"O�R�mڔ\' ����R���@�"OV�!�~�0܀P!�#�L�ba"Oj5HRh��+�TԐDʋ����S`"O����6%fQ�I�5M}l�"OV�(��j����D�!e˦x�1"OB�㥇����2h�J����"O� !�-�� ,^̀��x!����Nx!򄂾�t1aG�#g��gZ�j!�D=����R�:STy�E	�5h!���N�p!ё��V�F��31Ns!��N���gζD�Z��M�p!�N���i�jMG��l�B�A�}g!�A;PƠd1�O�K��A%	^�UI!�dP�5�\���e�r�ZH�Q#!�QR`y9g刪xp�<�#ǾU!�d�'*Ɏ(��.l�@$r�(5�!�Dء8G$iy�0 ��=�ԋ_9A�!�ُ��LK��!x?
 #�M�z!�d#(_�⢎�9.�ԩ���	%ij!��̣E�rq䕮?���� �@D�!�[�f9�|*�=8OLa�tKZ�"�!�-&���g�#D�a�$kJW!��%}�����X(r�(�ů"�!�d�s{���h����1fȚQ�!�J,�����1&2�����f!�oMl�1A-�1����#A�q=!�> g8P�H
�n˦(�A�^"[!�$֥5����'Hb��(�6A��H!�X{6��a¤߿Lú������!����&�)��0�Z���!R�H�!�$��������c�TiT�IE�!�$�9�l�J'Ø�]�\0�'.�!�$�"4na2�g *`��<�!�D@>>�p3���
�����7�!�D �{3`��	\��E�H��&�!��S�5?�y�@�W�hq�$��w�!�$W�HŞ�"�&	 Q� �@��ƌQ�!�Dϵ��#n}@m��,G� C�ɑcXhl�s��'Ob0*�b�z�B��<Wl�`�����ar0<��	A�w��C�I�w��a'ܗ5BzT��z�C�ɺDP�1i!�7:�X�3hE ]��B�I�6��H#���8�k!��86~~B�ɒI^�c��[6�aa�DIh�C�Ik���ҁ /$��y��G!w�B�ɏ'e��ZSg�g?�q`"�.Q(�B䉑k�R�r��ʕ��E�2)A�ɆB�A
�`��N@�� �o]<�hB�	�<l�x��e��)z�CAV&#�B�I 4�ָ8���j�ڒ���;�B�ɳw��$��/;0!�Q����C�ɥ2`h� �
=*];gH׳4��C�	�T���5�]�<�cB��9/�B�	y�Tl��	�r�q���B�ɼp��2��9��(s�
4h�B䉬1����˅�y�����E�j�B䉗V�4�p�Hm�4�ؓ��'WZ�B�8+��{$���&P�˙�
�B�)� ���$h�p�RQ���a�
)�"O��G�O�
���gՂ�"�	&"O� ҀגO~�T:dG�<-�dQ��"O:y�d���؋r%�r�N�$"O��J�N�?��<��*	�^k�,�r"O�,y��ä�$e
��\�؄��"O^�cb�I�k��q5(K�"��J�"O ,��$ͻ?z����Us��� �"O\Qq!c
d{4X�e�� #BX#�"O�E��iA
w��X/�\y��u�!�D*Z���&ְY<h�	'�Z�!��/#�N�E��+)7|�A��N�kf!���*5�r.�"%V����M'J!��4e�Ш���X�R	p�ڲ�w/!�d�a� �a�)-rX��
�E{!�I1>um �M��A�ZeQ��Q
H]!�DH�6c�J��u�P�ϼJJ!�^<N��IxU�K�P��@�#D?!�$�9Z�\�I�b���L��`�?E!�Dߵ[~@JE�1(8�җ!�$�7\��`(��ϸT������'�!���d|���)�)WJ
�#���!t�!�$�mY�\h��Q�I%đQ'�އ$�!�D�d�z]Ip����Q�8j�!�D�6J�hܲM<*e#Vd�!���$B�����L�bqڌr���!��O�#����dA:Lk@��'W=t�!�d��X�����ā�)S4��6N��!�ě>v��-��Z��Ҵ,3H_!��ӑ���z�$�>Zp�&� $�!�D��w�"II%哷 �����$/�!�dI�Lvԁ# Ȃ�T���#g�@ �!�V9Qn����k�I!�g!�D�	l����Ȅ=Va\[cB�`!�$�7w�~0�P���y#�mX�o�!��[�[�t�˧�H3
����m�Q�!�Dϗ"���q�&ӹ0�PJ�/a~!��ʨw[d��IO�mޔ���
�rj!��|��<��ΏP0�f�G�^/!�D��A��o·-�Xԑ�*̳Gq!�䓣n�L����8o�
9%+=Xo!�M=��e���7QH1�D�ʂ9k!��ԍ-��`sG8'b$ӫ�a!�� a�Z�s��^���ܱVkŰ)�!�̪k��X$�.�� [�*l�!��%;R���F̶1����@j!򄊮@�m���½g�"��t#�jE!�$͕���WM�j�r��٨@!��)K	NEz�E�`:|r0�58!��`46Ļ�c�=dY~,&Ač)!�D7]y҄�0 Qf!�@��!��]�+B8h��#����(��g�!�R�~�=�b W:��i����-H�!���Z�.��3I�4��I�֠�=�!���T�0`)F����xA���v�!�DG�VBֵ97`EA�b�Rf�, !�ٻ[L2�ȉ�b �����ٴ>!�$ �e������92~���A�m�!�D81���/W#FL4r���	P�!�d�5'�J��劰;�����K�7&V!���5�ms��]�C��|����Py��g~��r0��m^d��aϔ��y#ַ	�3�nU)`̦a�񀇣�y"�$CB�EPr���VW��[A��y
� 0�F�G;E�s	ѨT-�y"O���Q̒�1)
=ks"�5����"O�iP�M��F|h`��FL�7�!؂"Op�؆,�d�9�N�aH�}��"O�	9�mK?w��㔃	 aH,��"O��i�Ǒ��-�!\0��t"OF���O=9������R;(���5"O�+T"( �t�	�)��'��Yg"O����̓t4ftx'	��K��T��"OPt[��}`�YrAgN(_��x��"Oty�V��<�����*_�`��"OL�AG
��D���F!�Υ��"O�H�X��ӸhH"���-�!5!���Yx�q c�-&����H���V-�v�p&�A<����M��ybٿPv��H�哹dq�,a���9�y�P�k",�P��/d���&��y�в^�T���$��T?�����#�y�ID?T`~���g� 6k$�17&��y��U"�����5�� �Lޝ�yR�[�24Ș9FI�-�����㎛�y�Q�hl��M�$�0�r�f2�y���*S��k�Q���Ԫ�&۾�y�1��ȩQ��bBl���[�y�MV�k� X���B 6 ��U�W:�yR��{�2p�d��*�ܼ�$!	8�y��\��3%���S��E����+�y�kY4F!�q:MD�Z������6�y�L�%n�zȳ�D*��		�T��y��(Z�^�	�-U%AEz�� �D&�y��IV��$�$˶"��3����y �E��4���� g���
���yb�]�>���2fVl=�́��0�yRB +�x˱�)h��$�C��y��S7{������c�	ek�;�yHUTQ�p�.Z�)��E��y2�[�*�d��W-O}4@qe�y2fJmު���#��5G�bR�M��yb�0J���G�"*m�������y��ݯ(��P1�ߖ%:R 1@;�y���9��š�C��G1���Ѕ��yBfR����k]�*�(|ۧQ��y�o��Hcj�*b��(r���D.�y�����$�"�>I ��8�C�I�f=���'�u���U�JC�I'��!��29���o�x"\B�I���E�^j���H��G���0e>D��g��6&*6�`w�K��x�1�1D��˲ȯ5��]�g��C�� p3a5D�1�C=v��`	����2�D2D��#Ŀo�XQq�/E+0�D"¨1D�hڇ�H?1�����϶[��Q���0D����� S�𝢖 @�=,�:B�I'?�*�RC�$1讕S��ڙ[#�C�ɫS�9Ŏ!Y�PUB��^(#WdC�	>9B�Ӈa�0"��`/T�8C䉗;F�d1"j��.�M�2��2/@C�	.a:8`��ݘJ��P�0 �D�x��0?FH�K����  ���ū��]m�<�wfF|���� !�U�qg��j�<q�C!�-�re�}h��WL�<Y'�U$2I�(�V��GJTE�<�t�ƯC�n�5��P3vy���C�<م"�y�B��#G�j��y��Z}�<� ��5d�r�x0
�*i�L�@"ONmx3J_�mN�)���/����"O��"�n��E8xd{�0-��U#D"O�dN�D5�X�v�F�Ov����"OP�H�;c0݁�-�*a�O<�y���fy�̸%�C�YX���Z"�y�EƬw�����m,��Y oQ,�yB��
XY��6@����c=�yB�U�T"8�����< "�@�!�yOՋ���!!�A<���a��S��y�bH�;
���$7G�m��yR�WuD�	Üw>�i���y2�K�g�1`5�9XcX���ޫ�yrg�!	ۼT�2��IjF�I�C��y��@��$ZRh�42A���/=�y��[#�i�s/D%+ ���%L�y�o�))��|:7$@3&j�T�ŀ���y"�RJ�T�S��$�ZM���"�y2�C?R��i�ꏣ劑x���y'̉#����D*A�~;^=K��Z=�yBA 
ryα�fU�o�9������y���?VMc��
k����"ض�yb��T�����O,X-����$��Py�Dݤn|��pD X�+y���RU�<	���:��d�'�,Hc�e\�<��I�<E`���")�95�B�NS�<i�����
C٣���ц�W�<9�K���L��u'^%KJHr2K�T�<Y��X�Qyg�ܞ�L�	�Ex�<@�P�)���P)�<�y�&��<�%�
�9j� �"VL��Nq�<�a"Jj4��cI	�-�s��e�<afa�	7��y:eeI8~�s�dx�<���˖*�jt����OE�0�b^_�<��/�,Z"��S��{��P�g�Z�<@^�j�Hp �B�$t��N�K�<��eə-�BpJ4�&dfzЛ�"K�<I2U�v:�1���N��@�H�<���ֈc� �ae��7��P��k�<�d�E �0�;�4j��<!���c�<Y�^���54g(��c�<��fA��0���H�c(�:R��t�<��A^�x�
�{#)�
*I�]RC.�l�<�����!k���"CI�$��q�<��j��U����T�� LZ�X���l�<A����yl�Qs#�<A$UX���i�<��i�K�D]ȳ���=[�ݫ`�i�<Yg��;/���(P�
?M���3�(}�<�6o��R��#T�����C��]�<Q4k$^�ᓁ��F��؀INA�<a�Jعp&(q��^1v�N�`amd�<�5��)jߦ�0D���'�`� ��YZ�<�������,��ǔզ-��a�<�`���ɫgE̚QH }���^�<��%��=�SFeΏAB.�G�R�<am�>Rb��������i�n�D�<��^�>����v.TA�HA�<�$AZ�9�<��= _�yAF�}�<1u���:`�+�� ��1�S��z�<I����\��CK�P��,����x�<�ޔWRm����s6ڭI��?�y�B��B�f�A3n�	hۦ9��-�yT�S�~�b��bcb��1���y��l�\ rf�O�S��Hb��?�y
� ���$U�
%.���ڍ[.�Q�T"O�h���]!%t���	ҹ?8>�i�"OČ��0�EI0�Ч"O�`���CL���nV>0��p"O�@��˳&L�$[�Ku�P���"O�[��>5.J�"�H�O`¤/!�d�k`Rђ�!��͹�eQw!��ViV␒TI �|��Sc�X�!��G�@��KG.+2���� �!�䂅M��h�׌�6b>j�h�M=7�!�dG�)��yʥ��~�X���J�!�^�o/�ٳC"ֶ%�M�0���!��߷3�)��G�5"����i3(�!��7T��y6K�6�FpGf^�xn!�¿-޴����)�`<3�g�J�!�� 9lvD���lۼ�zЀ�0"�!��J6AJ&���
����E�#�!�ܓ���㍲;<+)�Ꝇ�Y���y���7S��E��t_^�ȓy�|�E��>]5ި) $T�V�ȓNFPAFO:a�Lɷd�fI6u��4��l�5	ʖ!��� ր%�ȓo1L8҆�,Go�7����y�
�'����P( �������.�(���'Pa9���o�~TI�$�3-R�h�' 5r�+��}���(��	�'�d���넥P��P/��ٔ���'# �J�[���+A�d<K�'%V�3�-F7}��-�&W�Q2q��'x4y�	�=��K���W/4�'y�,Z&Y�z���c[�WCJe	�'����v��Ÿ4�җM�U��"O~=҂�ݳG'R�A�&�&P7���r"O��)g�ۥg�	�V旺3)�a[�"O�A
q���9~PႆC��#7"Oty�d�Hg�M	q���Y)�"Ov�
gϓs@�3�5;(�a"O9��B]�� #5i\	�:�a�"O  �ˍb����ITX�"0�!"O`Iˁ"5-��]X]���@I�l�<�0 S�1u�|�7�чG��R�H a�<)G���߆�����-�P̲7hD�<�#I�x��s�"�[���j�A�<#g�d�D�R ���[��@��jD�<��a�0%O@M Q""|9bvnB�<A����{O��jƚ5��ip��S�<��2m�"�Q�X�|ji�2��M�<ǋ�m.�4�#O��E�%p�G�<�CXw&��#2/ˡ:���D�@�<�\伤# ���l�s"�z�<� �T�<��1d��|�Pc��s�<A4�7�A��B�*������f�<�DI�1^\��O)	��E2�Db�<)RK��6�Xi��Թ;ʄ��׋�S�<!�'ݺo�.��G���p3�pId�S�<!�$ߗ.�d����0g|]��`�M�<��"՝	���Jâ-�.y룏�R�<yPⅆ"mdL�!�ȧC���X���Z�<a�N�T��E#Sˋ&!�|�w�X�<Qw�ʇ���h��=b��
0b�[�<i?��]�gjҩM���	 �X�<���"jNqS`���<q1��{�<�ѡwS�P��sajTQv�x�<i%�=��I���.)XH�&�D~�<� ���ff~�TE�d��=�� J�"O�dZ��א9�} ���M{Rț@"ORT(��OR4dX��lΗ`o4���"O��q#o�9V�e���/$i�@+"O����gV����2�ͣ+7t��G"O���ݶU�l`G�:H��Kt"OV�bF�S�Rhb�����jd쫢"O�P��$��L� U���"O��YBԼv�f�6�0d!rT�A"O��H�/וe̌ B��&{JY��"O� ��ޮF������I1}�,��"O��+�f��`�HX�޶Z˾��"OȊS�3N$8�㬘:q�P|�"O��kEF�2ּ<�k�=���T"O1�c��J�d�u+EiqLdv"Olp�J����x��,[_x�
""O8O]%7GFd!6��! �,��"O���"��
G��F�h� �"OJ%�D(��f�&�H  P��"O�[�4	�D�X��IZ��}[�"Ov�Dɇe�����R�?� �[G"O�=�Q	$l�f�bF2����@"Op���C_�ՎL�e��}��H "Od��4��� �c�,�}b"Od�x�"׾�ֈ#
x���CB"OX̹d�!4e��H�#2I�6Q:!"O��[�]�X[��hF�ҪP����""O�+��)nV�c��2n
P���"O*e��f*N"���#��-��z�"O`MqF_�X����J�8њ,�A"O��T�J�P��:%J�-(�L�ҥ"O $��F�=w��I�FÒ�f�ZŃB"O~�`q��
��� �3gR0 &"Ol
�l�z�p��M�X#�*�*O�H �Ni�PR�
��qh	�'#��sg�3�2��pG[�<e2��'i�����ɲiL��
�NС6JF�3�'l����*�X���*���p
�'�v� Sb	4N4(�x�A1%%��'\�Dɰb�)�nu�YØ�	�'Ć[����,��*_1���{�'͸5��y��ժDf<
��
�'<�g�/�K�8z!@�a�f�<��C�H�9fCO2Q,.�3vDn�<�C�Q�t�B(X1=���9C�
l�<I�ҺH�s��V/N��I����R�<�Q��D���,nqw��I�<�I��W�:���)�~t��8抐l�<�2 O���!���H|�hM�$�_O�<���!n��-��ʀFj=H�IO�<A4j�6L+��
:t�8�e�J�<�gN߅I ��*�X q�`p '��L�<�!�Z`��A�Q"�|5`��F�<��)1+�T���3.V4\Xs*�~�<�	S;[�3o��\���x�<q��3��	��++0^�2-y�<y@F�;$ʤk�� ��X!T�Gw�<q��-S�
M!,���(��
h�<y��$H�	����jL�� 'e�<�ȏ6-�̠�f�Ҫp_8���`�<Q�*nb�q
��% #�t ���Q�<y2@ϙҼ�J�(;͠�6�_J�<A���>D��-�9_��b�}�<���*�8���c-8j�U��D�<� �9�J��(�K�h�J��q�"O��i�O�n�����Q	��q"O�=���.���EU����`"O<���n9�&)�*��U���+e"O�D)# �0+7BL3t'Ɯ`3�!a�"On����W�$�4�T��z�5�!"O�i�`%�aN����'���a"OJ�A�6]���3dĹ5�BA�"O��󈚡���q%��R��h�"O$E"�g�4�D�Dg�
IUnY!��'������G�w�.��3ϊv�(�B!8D���$�ݳ7"��`:qz|�ʔ,7D����OnYk��8�T���8D��(�(�w\�x곁��)���-2D�8���!BY�e��D��=I�1D�X҃��)`�$A�$�‵0��9D�ܹ�*Y�
�I�I ��n%�p�"D�,IW�� J�L��g�@�p�+D���bMeբb�$ɟ&��6h-D����e��D���m�.���j��-D���c �I�~L���Ůhf̐2�.D��*�O�?\��  6h����0D�)�B��gb6����ϕ���"k*D���I�3Z�0�c�F�?Kbz��j'D����ϙ0�L�	W�ȱ~ �=���#D�$C6mȍZ�8�ZT4|��?D�d������[�J)o��BE<D�d��M�S��0��A�6�Bp,9D���!�\%:vY+��s!�ݹ~�xC�%#�Z�q��	:����<=:C�ɢR���g+E�8 @�8e��f��B�1x�$a.IB89�b�xٞB�	]H���O�o�` �*N�5B6B��6���2ec��l�PD��ڱx��B��I,Lu��F;?8*�p�%�?�B��k�N��$g�=oiD6fѮ4VB�	��q�w�>'m��C!~�XB�	�:pT����F
Df��R��$RLB�I�&�|���R�|��W��&{�B䉛 3�x���_�M�T�a�	�\��B�ɥBT����52�8(�DS�|��B䉘VpP\�ӒAГ�U	"4�B��=Y�t�"�N-s��i���T�D�B��+:�<���A�&�^���-ѡ�d�9WQl@���$,&d�2&;M5�y�
-�lqK���'0�����Ԛ
�B䉽"�)�*f%H��g��X�nB�ɒ<�T4o�&C����g'04B��>\���A��:
 , B�0L�^C�Y98��Dm�@ۡ Ѯ&�C�ɪ2ҠܘU��9`�έb�̋^vC�	�TӚY)@�Kf{���w�L(@*B�I�N��̫t����!�4ΈD��D�O J#�6���p�d;L ,�Q�4D�|av(��`.Hxp�Ćq�4Ġ��?D�t�1/1r�(�I��ǺgCZ���>D�,Kt!BJX��*@B�e!�Y�c�<D�p�ři�`��� ����CS/;D���"R4CF ��w(Y�_�>��eH:D�|Ys�>B�`�"A�Y ���$4�(zA�{�EI�E_S��H�ek�B�<� �DN��n��J���3j�W�<���1k��1#��p�"H���J�<���V؀�(���s�`\�DSD�<� �A�C�܁R�41��&F�`��"Ov���b�-|�n�QRF�MV���"O|�)�h�	9W����O�N� �(�"O `HU�W�̢�0�DK�M��� �"O�1z�j�#w'�-�$iW�5�e"O②�������Ǥ@�xځ"O�AHtN\AlP�x��n�,�r"Oz1��cj%��R�l�Z�"O��"BeLw�����\	[ɘ�q�"O:1Ǯ@�>���A�D��θ "O�4�E�A�1��C�f�hHk4"Oȓ�ǒ�R�>�`"�70�J\��"O�Aqd@%n>��"A�J��ju"O�L�R��"<�v)!gO�j>`6"O�Ń��=5�p��@��4o\2d��"O81`DE��""l:UkESx�&"OHIR��6o�Ȇ������`"O0�ᣌ�d��5��X�����"Oޥ�6�^�Q0"��j��~�°"O�p ��X�W�L����|�`�k�"O`19�c��4
 ����7!��C�"O`���D�=Q�d�L�����"OAR3�K�j\��`C #\�yBa%W��h0��Ww�p�*�kD��y"�Őo;��i�.�5$hR	[�Џ�y��H�Nl�!
�+9�� K��y���4C'~���,	��z��[��yR�p�r�C)�du��ER>}I>�*	�'v|Aҷ%G:��'�G6bxH�1�'��m�b�J5Q"��g�F�`f�Lj�'�R@g�p �����ф)d��k
�'A^t�!����b���ux�Ű	�'[5@��
�]%Z��Q扲>�l���'>�t@��ݿX9ЄK!�66*�	�'��@�B���4`!B��T$-��t	�'� �10�T��#rl�(.�my�'�|u���)�>!���+�!�
�'�] F �,w��D��+��G�B��'��`�!�8��⇄�5P(���'�H�����?Q�0��i�>�p��'��ۆ�H�A��2lڞ݄���'kf���>]{�����B�~�zq`	�'�T����gKެ��T�r�t��'` qir�:-���d�q څY�';���1KƞlV�����1q��	�'����b�c��8��K<���'/T�2S����9@��۝.�� ��'�����[����3�\:"�>��'�p�p§�EMfpÍ���՚�'N�5j$N��صs-G��^���'���F�F9'�fȈdmƖN�Ij�'�T�P&�U�,�ZʓH��8�
�'#�E��d�N�s��D�R��
�'
��持G�(��FjH���̰
�'��HO[�|+��ƂD(P����	�'=<LhVb���@�Y��ֵ^�L�	�'� �īX8fr�*&d��[y�8�	�'�&�b$J#V�Q(�'Q�ZJh;�'�
����H�J��%JI�W9`h�
�'�P��f��g=�����C�=n�qc�'��X�S�ۧF# !%��5&��	�'~�\���*<s�9�T&�ZT4��']�0���?`�M���	(Ω	�'T��p
L.e8�x1a�P(|���� \��$�=pvH����$!����v"O.�+�$D�F��*�2,.5�q"O��80,�:��� H?<d�RE"O�!qL��uU���q�֜L�����"O��A�C�=��XQ^d���c�"O�݈���E�h��Y5z�ు"O<� EE�]���R�I)m�+�"O$��P
͑e�A��P�C�a��"O�PapĒ1.��;P� `U�,�"O$RTE�>�<�a�L�GC�\K�"O&����ar�D����	&(��(�"O���F@+2V�{l�v��C"O��!�I����D�K�C�ur%"O<	���$)q��R��V�|:f"OD0x7f��lx��DFЮl��ȹ"O�aYƢ�"?��,y�ߛ��p�v"Ob� ���3��Ya�CX��6$��"O��S��JhEء�Q�er�"O�l�3��S���Q ���Km��3""O
<2�"ʏV�`]����^-��"O�}�6M��$��D���nY�Q��"O�ݘ���S��9�5�YQdxѤ"O%0�i�c>d��
�
pc��pQ"O����I�,�|�U��U����"OLPR&�7�����" �%Z�"O��3-B&&������*-)"O�"�^@b�����*#�Ƞ�d"O��Sף�*�����/�2QZ6"O�0&�B���,	�DE.��`��"O�4B�J�8	/b�;�$KEņ$�"Or�'��%��<�DM�N��Q"O��(�Ň�f傦�L3W����"O�=p ��\6T�ô�?�Ԙ	�"O����$G n��C�A�+8����"O~��EG�"$Ȱ�K5c�ޘ��"O�,Cpa��o�:țV��nD��"O��S̉5r�T��Ƌ-}�;R"ORu�v�J�d���Fd�.}�1�"O��1ר�?K}X5;�$�>'`��"O��@ԈA-$NLI��I�ް�3"O)��Sd5$ ��E����i�D"O��:�V�7C0�)!�J�p]Â"O�*���E=0�xP��3� �y�"O��k�ǎM��DoV�R���h�"Oj�����b� �����ɠ"Ohݫ�j�-�� �.J�ge 4h�"O��8�*�(���:��8To��2"O����)^�
RF�ƍ*���"O�a��`�'J"|�K�a�T��@��"OzL#�eO�IE�t�� ��h5R0"Ozty�řEt$t �����a"O�}� Δ��B���.ب�����"O^h����JG�1���;�N��3"Or@
�O�<p�޵%˂A���P�"O�s�JR�U+�����i���"b"O^�����'\����J��@�"OB\�%�;��l�DU+��=H0"Oڵ�5��h��qd��{���E"O��i��&+�2��ƀ�"e�A	#"OP�K�aQ� }��@O_ 8�"O�쒁)��Ws��2f�Ur��`s"O:���H�	�dтn�2}�<H@"O�
���kp���B^�e�D��A"O�CᏛ'N��SF �da��"O� L IA�g�(�(!FZ������"O�L�!�>3(����eK�1�Ԁ�"O�Q�1�ʏE�ll�'ע7u昁�"O�R%�K�"������,a�Z "O�1#���
�
��QFߙRI���"O4�����-��@Hp��;�&�"OΤ aѢ:͊什�A� ��QX�"O搉��¡6��<s�,�p}*Ux�"O�U��L	�?j ���ڹ�`�6"O�� S�k��HKf�(a�肣"O�\���
T��(!�
T��� �b"O�I�wFJ�u%�@bA�(
��;�"O�m��h�7Ah���"��%G�
��q"O�]���Vo����FV f�2�Ѵ"O��Z��?u��x�bO�c��	��"O�M�fB��������&E���'��'��)�3}��O�jz�hE㏸�Փdf��y�y���*HV�lsS� �F���Q�'i�I���3(BY*c�E�U���`�'IR���G"o�Ʊ��-@ L����
�'=�|�ҍ�1Ch�YJ�Du�
�'X�`�r�(+�x��f!�5{|\��'�l�����-<#��ic��w#(d)-O�˓�0=!��DuC�ѫ����:�� Pe�]�<��	-Hy��� �R����P�<q� c�F�0��	:�ZP	�F�<)ѩW�ys�e�GME�7�� d�A�<���(��C�@��e��C���<�` �xR���[�i�X��d�V�<�e��>?�X��.I���E���V��p=y�'��H�F��w$��Ժ�a�4D�l�!�v�PQ��)�kf��6�1D�����Cl�Z�I�:Oj4ղ1;D��p )�("�t���W v�\"U�9D���S�H����	r����Om�<)P�E:vD��$��nj��υ]�<y`%ӲBhX�i��_S®6�N��?qJ>	/O1��R4j��F�4�B�k&LݛI~9�ȓPj4q� �χ> xA �Ř'�.ńȓ�F�j��ں3{�К�ƁP~ ؇�nU�t���Oޮ̢s��1ymF@�ȓBr��9VfΜ*��yé�~? $�ȓIN5"!��.��01�R�<$��ȓ�VLK���j݆��芏8��e�?�ӓ:��}1$*&ހ��GA.�$U��abL����7"�Q���^ԁ��Co�Dc�ùz��9��͇6X�D���8;�]X�K�8R�H.C0K���ȓi�A��G8��4j�H�5b���ȓL��8�@�mֈ�p�(M}�܇�*A^m�U"Y��t��1h��?��Q%���'�ax��q����'"�"~\8Y4O���y"�K�4�����A=,��]hԦ��y���Y�ɰw�N�����E�y�P.(�=#a�K::4�Ҕ�H��y�J.ZAn̈P��n�x�P�	��y��8$��y�e�U76���2�y��7z��S6�߱z%�xҗ���y��^H��Ew�*����/�yr�
,"4����EN6�b�d�3�y���'ZRyB�ǆ+�.U�&폏�yr��3�D�੍�#kƄ�"��3�yR���c�����)��S��y����E�,�Z���'��Ųa,O��y
� ls'��Eh6ؐ�Aԫ	����3"Od�9��E"`�0�Ѣ��D��"O�陖/�"LY����ϛ�V��ѵ"O4�ҧ�Bx�p�A��25w>��"O4�A�� Hn�P���d����*O�|�vυ(X3��S�n51�T��	�'� 9w�L6A��d�6N�(����'��qf�*B��L"6��$_���'�J�1ש��'���#���b`���'t�{�  `�r4�gʍ�n��x�'�Ĺ�
ٵoB����̂���'���2��Ҁ,6��#r E3�`��	�'U�P($c@�AJ�Ժ��U�{���'���JV�Ѝe#쬒 )YkpE
�'�6yy�D�N��+`�E�}q��
�'��}	Ө@�?*�"�` �� �
�'$@%z��V��X�s�'��iA
�'f�)�_���$��e�<&���	�'�0�F�[�%b�X�͎6�Bej�'�*M��L�^A��9��R $0,Б�'�qf�G���WC�.���'�(H�CŰ
6*��6OȆ}M�M�'��XBp�Z�&`j��2�&v�����'�$�q/�f!�¤A:_�,qk�'���#�[- -�6e �S TX��'d�i���ʔ;��s�DAԠ��',e�k� �S�l�j�:���'5���`D�/j�$Lː�Q�d���b�'��Q�M�6t��A{%��0^^��p�'.ZL���>"�N���~9�
�'��e�e�\U%X�:���8���'���S�W7 ,�ȲEV/34ݓ�'"t]j1V/8	���D)ո��1�'~z}0K&_� ���&���p�'�*���e��L�^�����k#��
�'�Fa1�KGz\t�Q�E�\�,UH
�'`` �*�\Z𪗒y����'���"*|��PbeP���y�C�'M��tatjةx�(q"@[;�y���O7B���!�&d�K���&�y�-��md��+��u���X �G��yB�<H)��'mh3ز��A��y���0�(x��/(=�h�t�T�y��D� Ȝ���ǁ�Cp�뀆H��y@$T�J=�q��/?��hC�̨�y�#� ��`q� '8�T�rW�U��y��_�� yEA��(��yxV��y�F:N��xs��/<���Fm��y�)�-~Ȯ\�Ba� "9�)�e_�y��O�(�`��+1�5Qi��y2ɘ��j9���
�8��QG��y�?�B9��̓.a\��P���y�;.ܱ���D
{ڤ1�I �yR�H/} ��B�ˋs�����,"�y��-����g�f} 'f��yb��h81`�ő��T�!��y�l�d�X�惇�X�j�x�@�yR
݅Ki6�s��
�I�^�Sь�y`�<4u����j!v1	$gT6�y�n[��&D��/.l��tT �*�yF�Q%@��qkbT�*�J�y�iA
j�(PYD�/H��s�S��y2Â�Q؞��h�}z��ڰ�y"�ۊ:N��� �f�6L
��y
� J�땪/v��t�Փ1=�6"OPx*�#�0OR��v�0V�0 "O�!%�	��N����� $�l:"O��Ҧ�w�~���g�/7���F"O�7L�$R�C�B|��""O�MW��.4ʕ�f�öGf�͉R"O�-`D�G:�����lZ�cT�"OFr�aȞqK��Ic��2Q"��2"Ofm���U�Wbf(�ǯ_-Q�a("O�m����mբUB�.ՙ0� pc"O>��ue˔u�½kw#,_�t"O��vO�dz�S��H� D�d"O]�ݥv2�%b� �6Ry�V"Ot١� 0��1�!k��X@�"OB�( ���(�0�D�(oۘ��W"OX�C��#��y�'��/gR��"O��Pq���%(�Pe���Z�U94"O,�B��)-^x0��ЖSl�]��"O�9�.����2�FO4w")��"O��ǔ,d1����� w6�%"O(x���1KHݐ�N��A|@�[�"O4�+��-:��g�V�7[:���"O��Ѓ��*��h`W������"O���3���
�h��,��w��-�a"OP�:BW�C���(BFǆ "te��"OĨa�eғ5|�����T�D��I"ON��'�E>Q}|��A�	j^�!�"Op,�QǛ4|�-
��݊Dn�T{�"O�A��9~&<̘�.=[�j13&"O�=	����Z�"1�V�N1ȶ"O�0sm��f��Y��߲x~V\"O��`�IG,&\ �Y$lJ�vtTHe"O���+�%\ a�L�:+Z��c"O�Tz����yX"�R�A�%�U(�"O4���Ƴ}�8єJ\>d��=2�"O|��E*E�	���bp�^���"Ol1���(8�Af�� �|��"O���F&v�Q�� >�\}85"ONE��Z)E���Į��t���"OjS�A_u�)��cU�`
ԣR"O��Ys�żN�"A[8HM�p�"O��cuh+Jb`)B�P�<�$��"O����`D�+����nϺls��*�"O�mbs��Y4�x��Y�'[�ۑ"Ox��#IΪb�2�c�!J���P"O�ث�/4$ӄc���#�JA3"O���&�?"\��7��v�t=�'"OV�`F�h����!�ء�.�D"OV\0p��	~e���� ��$3v"O>0�0�гV˺�#�"���D5��"O ����"%������b�Mb�"O���$�ɒLd����:<�5 �"O��33��2�qb�ʕ�E�<�Q�"OJ��$��qpx�RDQ�Z�9"$"O����DX�"@��It"O0�Cq�Q�$H�!T֒�d��y"cN*`�8�� >�4ȖL��yB�C�{3P�e���2������^��yڌm���@G%�"^ RC˘�!�_=o��iƪ��^� �RHZ�U�!����b�:���y>@Y�΅�!�DQ�����*uZ�]"�����!�d��fn�+�l��uK�	ZE��2!򤝘G�\4rC��RB�u/�zN!�� ���֗_Ʀ���D�e�RTx�"O�]�h�(l2�D��+ɸА�"OJ�%C�7����s�D,���"O]�%�%-ߘ*@�F��f %D�hӤ#�!z���k�oۄ%;+��!D����c�6I��NZ3d�x-[VB?D��dA�>i��#��+5���>D��$�
Rdj�ɣO�*�Q:Ï>D� �&nA)-�.X�F�J����Ջ D�P�Dӡj.�����Sﺠ*� D�q NW1%���CN�i3�X��B>D�(��)����Pr� �#Rr"�җ*>D���	�I΂#��F�,�ˢ�=D� @�h�԰a� ��*�$�qe<D�$BU�θn�le6*�;-�gJ7D��Ue�r�-��n�c5a��f)D�1K���4�ŠW+�ʕq��9D�4�w��J U�1U��M�j9D�(���� j��@N�b/l���A7D�P���
�`�!�"m�!�*7D���E-��Ś}��뢼���5D���ӰxPb��CVc�Ջ�*Ot���A_S��m�,Ԫ���"O��v
9@��`YsM�\�����"O��� ׄ�
�B&�/��љ�"O4j�o�(�hͫ"_3k�)��"O�a"����h��\7\0 )�"OX�;���	�$Äቸ	r@Z3"O�Z@T�l6��[�����&�ybӝ(�������q��Xw����yrf� R�M���	�b�ALB��y"��&���٤��_�:U饍�(�yR&���]Q�^G�ׯ�y�J�n���C�W(Q�+ˈ|&C�	�O��ѱ�_�PD��ǅ'[��B�I�8�*������9�<=z�"��F��B�I�m�r��"gY%$`Łň�B��B�ɰ_��Q�E�
 �zBI�%'�C�*f\��c�đZ��hj�DTm�B�	�a��eQ䓔r�мR�h�<E��C�	&C%���䂈2���T�
,��B�	^�ەȇ�`�,��
0j�B�I�nF���	;A��b'�7��B�I�BT�@Pjش�� G�ˡ�DŦ3e������-�Rص,�{H!�$ ��p���� ��Ȓ�6T7!�D

�`hV��8���j��I�!�d��L��u9U.O3G�*�oMj!�D,Ow�sU��:m�ݳ��Ãt,!��ݽh��dz"M�E���P�Z�!���2wf�<S�:Y2<U3bbڇ%!�d�"��QAգ� &>�����mH!��L��p�`3~9��	V�[0!�\;f�\�
���(ΐ�ըO�y�!�d�<j�xsHS(!��S�Z:I�!�d��m��yw=�脠b��!�̷xθi���ҎY��HA�H#!��Z�p5$�� �I�A�V�{#S4p)!�d	[*
�ǼFo��5n]J�!�d7�"-�7���3Qe;n�Z!��Z.���h�GџMY(	�#� -!�d�4Ť��3��Jt%1�j�!�Ĝ8mv�S��'@&�:� U�A!���5[��<;���'%d|2�TD�!�� r)S���?)IR��n�=ܰ���"O��G�L��t{��.4�P���"O���b�B7�DK�`��j����"O�IT�R�H��a�ک�F"OJU������ԉ����
Z&8Tڧ"Od��#�<_N��@ĈQ�&�!�	[�O�fc����#x���DE�'��8��'�\��g�8(�]��X�2��'�~8��ė=�3��S"G�������*�' ��Q�.	kv����H
I#xX�ȓ:��Y� �Qd�r�b
P�)���ढEE�Th��Ĉ>Ivt�ȓG��4
5� �la�8�8"#��=�
����ĀU9v��Ǯ۲%��p��M� 'W�V$zt�[�Z���BFq�<Q���$t�I���w�|�4�Pp�<YT��`�5���J�w�@��d��w�<AV�$kW�	�K�������Xw�<�0mF �*��S#ցITBG�Rv�<	4h�-SP*8ؔF�N�y�c�p���<R�[8����G
?�aI)�b�<QSH�=F];u��&y$
T��U���O�4y��:>^���\���.�y��ǔA��,R�`�2�R`ŗ,��d-�O��f�U>��l	S%J7|�i��'��	l����t��>�F��k_�"�lC�ɲ[�,,�h��t�p�ȃ�,b�<����:����2q4-��$'HJRh'��*�`B�I�v04-�P+��E�n��C�=,)Bb�$��p<Y��4aζ��֪��W�l\�'��x�'>�?QQ�b�4���P���|-�� �l>D�H+G��1��ʴ��e�$���E=LO���&�D�����S�z�� �釀~��^��H���K2䛂�Ez�$b�����	a�Oㄕ�Lk�>�!ꇳ>$Z��H<1
ߓs@$0*#���,�H�+J�\r�Yưi(�𤖝3�F�Cc�.��D+��K�Q���(�|�S宔�:�N!r���"`������2\O4@��+X�G{Eʑd��6��<�C�i�Fy���i��,"��D�p�\)��&[zJ�4P$�)��<�  W�un�rEŖ:.6,iS��b�<����%c�� �+_�{զ�<�	�]����%��f�����ǟ�n�����hO?��r&Z�T��dr*J�e���+D�p�bd�I|Yd�T�wv�H�K>?����=�7��&�8�h!��((�P�+w"^w�<��\	�Z����S�3㨸��v~��'���� c��QҲh�O*�	�'�X`⍄=딁��K@�|����'<"L�cLL2�P,����
L�Z	�'ݞ�K�!?���c��3:�5B�'O�H["��6:~!*�ć�,>q�ߴ�hO?7�W:+�D�3HA�~��ӬNW!��#:H����L8�b����]7\!�D�]�^M��oW
@���؇+B�%&� D�H#97�pS.�/v,��`O��yrF��t��x��+K��c"��y
�?�$ s���Q3����,��y�K_)Q���	�E%���˴J#�䓾0>a�#F.S��:�+��z������`�<ɓfːG޸�c�ؿk�ұ���Be�<��h�t�"� 7n~e6��"�F��E{"NT��M�iA�D�ivL�V/!���Ms�|8Ci�.L̹ ̛�,���hO>� ^����TSpR �q��;l���c�"O���s'ź^���� �O<\�Y�"O$-�u@F�y6���$�+�lHC0"On)�� �,[��RB"��c$�m�"O�9p#%Smfm�� ܱK!�=��O�=E�D��.6�vM�K��	9�MkP% ��y*�}��<�d,�/| �S�Æ�y��iό��=�����'��X��I�d
�"E5^�nT��"O`�a'��5�Z<�#��:.Q�e\��D{��I�;#�8E�5ĚO�Tju����!��
n|q�b�C�����FLÞk��'���$͘
vt�1��:d<�+��?��h��(�@����A�l)�ˠ&�jhKt"O�t�RD���h鐨�P���������E��ȁ��
�G1;@�q�"^�y2��(��S�"Ҕg�b��s�"��OT#J�Ȇ5�F�dK p�,�`�Br�<р͟K-4\��L��,�'"AC�<�!HT58��$��3Q>�Bl�{�'4ў�p����A���͠ ��6�E��H��Y��
ޒKCĭȰ�@�K����S����,h ң��k^��	���-Ğ���j3D�p+�KԹ�p)���j��� �;D�,��lX����Ȕ3f4(pZ`�7D���u`���P5������B#D�B���?y��K%�J�M2���'D�t��h�1A)�=���bPHS��$D�L
��<�t�6o�!f��=� #D�<�֫����s3��9{�Y���<D� �X��}h%"�*��GE�<0�O �=%>�yS
L���!�NO�,( f�9D� ����Q��#��ҊFe`H+��#D����ƫe���z�$��d���3*#D���B	�_�0��e*ɤd��P+�!D���'�K�)�����	�#^��3� D�8���8`2�D
=PZ�Y��&=D���` ֙oɜ��R�
1^�y�n:D�� %,�;T?Ν ͽY,y�V�5D�������,���A2Y41�w�1D�d��.�%��GA?�8��*D� 2�_�E\�3��^17=��:gh*D�i��Ĥ)�He�[/�|�-#D�л��W��B��!W�%��AR��,D�`ae�Z�->J ��aڇ�r���
*D�4����8��q&*�
�\E�7E)D�H0"��r?�� D�+Ft�t�3D�<AwjIr�+��@ʤ�$���hO��hm���]T|q*��D�kZq��"O�a(�� n�-鳡�E0��c�IG�'
�I�4h�+�G׀w\�1@c#��C�ɡ\��Ђ��K/�E�7M3��N<�/O��=ͧC�Y��bH�����j�t� 4�ȓVe�lt(
,44�sF������ȓ�����"\^�h����J�����I e���$KZ���'��U�(�6)��k�NB�ɰ4�$�4��%����?+�#=��|<��݆.�vj�O�X+R�ee�JN!�$�d}��Q ��F��g��r��O�=�� q��!TM
��DD6]�`#�"O||"��� fѰ�n��*t���+�S��y����V^�	�g i8�J��yO�@�xlj��*����iF�yr�͐
(�k4u�x�(�+�yRow<:Q�*_g�LDkB�@&�y
� ��)E�3|bL��C��++�\�Q"O̱�h��W|쵭/
�A@��y�<	�D* �Ta�P呠2  u�w}¬7�O2]krŜ�n;L�2gɣA�`1�U"OPq0҈��fh�3���"O&0ȕ!ܔ �A�)$g�,����4�S�S�����LI1tx�f��Q�,C�d;�0`��K���I�4��2M�=Q�V����O1)�ส�!ڂ3�h�ȓY�X�WD.V������rĥ�'�&�c%_!��C~�ԡ	�'�(I�2,L�@��1���
ļ�	�'u�s�O�%����W={͸a��'�x�!����(�H-"+7�t��'�t�Dkʨb�u�u�����
�'>�P��3g�<�����9^rpR
�'x���H��v�M@n�C4"��'(�9���iv(!���¡;P��c�'��!ĈPZ��O��~˶���'YʈX���}Uށ�w���s'��R�'zm�*�{m�� ��p���:�'�$�a �14�}��do��'`�Yc��ǲ!(��3��|� ���'�N�����9DQ^h6���hvb�'��-@�!��N�R<(�����'�4	@A�����A���<t�]��'���Z���8ږ�Z���s�tMh�'�m�B�TYE����тqll���'�%���ì#��tRB�5p�H�j�'X�@��d�+ ����%ѕdYAy�'�J�a��_+{�M���κ��'5 �;1gLX�4��cK�=𲱉�'�xyYӎ�:�F��V�k`-�
�'�n:EG�|��tb!,7�x
�'x�����<pN�9��C�{�f���' �R��Zp u24��:c=|y�'P|Ap�k�t=.��#��-�'(N����n?2�����
LVe��'�B-Ç��f�������00�'J:���
�}� 2T�`�'��]�Q�vD����	$�K�'誵ʗR��4���6HE��qN�({&n�Y苰"T�ӓQ����M�'6���[CKQs���N�^13'�@) ]{C�ݕ}}���Rf�)�K�-���z�*�_�.��g���QE	E�i8�O�����ȓl���؅Ԩ j�pG�q�1�ȓj�����L!ޔ�P�D�D���8�#��5l� �S�m��P��b&�}�T��&��xrc���p�P�ȓ|	�)��`R�F'2�qDȑ�[t���6�qoB& ���3	גfa���ȓk�j�B4E��[d�(��
�$�$��ȓ<�@Ph�`JS����-��D��d�\�zPdߗ����2�ϬM|1��W�Μ�����Sŀ)^ӢЅ�s�z<ra�2Me�%��g�Q�i���fśs �I9���C%(�HM��o9�4c�m��<���B��,y�u��DF����0<�`ѱ�������xM���=� �'Ö��vB��:k�,�2s��3Q�L�s�R
7��B�-'��Y�H�6B]� Qd$Q�C䉷��P;�C���M:��Q�Q��C�)� ��17��v�0Qrn���4"O��`�24�b����P�1"O��)�/:!ȁH��_�"�x��"On��r�U�(W��UH	d)>���"O�\4��N�P%���
66�k�"O��)��9P6����049�"OpI��ʑ�%ٔ}�F��*�Z8�f"O��O 7%��89��;F����"OJ��A���g�a�����h���w"O(T�A�IDl�oB� ֪���"O��#��_�V���I$.��]���K$"O��HG���&����P;�ȅy�"O��Q�C
�e&za��Fl��0�V"O�x����+��iA!��N >�a"OбC$�@*(vys��C����([��P�䋯4��1�On�ȓ� �r��:�p�i�g� �H��ȓ}��Xxf��V�,�QE�̂0fơ��\I�@h��meLhq7fO|���
B*�rf(Eز�A#DY&X���ȓDV���~U���g�8L����\��kȕ�p���7s�y�ȓhY�t���7E��kg�L�a����ȓg�PhB�N �&8����9��h��\�:�!J�*!F��J������CiKSh��mؾeuu��r}^)CrT�$��p����4=b���*���q��O�Ψ+F���ȓhb�H#�H<j��,�9��Y������7�͎;C�1�7�]WW��ȓ"py�^�A�e�T&P�z�`І�}:���"�;� ��V�ӪB\�ȓH�%��V�R�`=���%5d���!�)8�g҆;�� H٪N����?Q��>~@
�[���'YPL����n�as�@�z�!�B�|�xR��	q�,���F#q�" �w �&GZ�'�#}�'���2B��V(���D�BWvQ�'RfɢD�«5��ɰr�U�5�Ѐs%E�HB �bS��)X���5i��P!�F']P����j��z�@�64Uiရ�֛VÜ7O�X{�cȲH���B��y"��L�����=BN� I`�
���'U�8���o�b|���ӓ
dB�����38���j\W��C�IV`jA���N6�z3k%%=� �&ח|wN��,O����Y��i2(�
[��؁F��@qƥ�Ǭ*D��ru�ȋ;Ć�	�N
�1IN�{�X	Rb�'�Â>lOXb�,�D
�DBH�8�h(���'��C�"�f�CU�i0��k�Β� l��"$S7>��� �҇R��d�G��g��C��㑡z���rnP�ڸ'�zQ	Gȇ�=�*g�:
i��i��O&B����a�E/i�N���F��7*�'�J#}�'d�<��$Skd���א]��"K��Q"��>�&�)��	ՔQ�'����/���z,c�3U�́��j] ����AG��0>�����b�P��!�Ah�4tG@�ޟ8�JŨ���q���@P�y"I�l� \Z'�P�|*�,�n�ij�����dBQ�GV�<�H�'z��@�&@6��t�dc�
�Xe���ui2���H:^��`�g���yW��!ΐqxs�ۆp_d a3J*�y2�@�g��4�r�Z�q,����j\8	y8	&�-}�5*�B�O���f������E�A`��y��A�eO����\�N�{Ҥ\�����A�Ҧ���m٭X���`P$CQ��tc�oޫ[ܘ��N��@6���ݨ�P)��������%Ը��O��"���W?��B��(4��	��J�r��ӿ5>�p��8�zH���˟nLB�	�,$�mj4��y6x��冗4����ߥ@�fm���X^d`q�0.&��?�ϻ%Ҷ�E�ӥ8�����Y�<����9)B�	�,��Տ�8P�u  iY�"`X� p̓]����?1	"�%�-�
��q�P0e'xa���6f�E��I]p[&�%,��� �%k5,�#Z��"��~�T���'��)��nX����ڴ6ِؒ%(?V}8g�,�复�U�O5�h����s����ɩ����C�EP"O�=��O�,n-b�s���4g��i������������O쥉7	��w1L��'l]XL@��"O�0qO� d���fIQ"�5�=Obf�츧������]0t!���$���Zg"O����ϗW�TD�N�Y0t�0V��CQeӻ<bń�	<[݀���bQ,X�Y"��G�?�����Uy`��n�EČZ�=���jË�l�����''b��U�K<P�āiu���b�Z��գ9V�zV����O���O4):�ܓեL�,K�%��'����VEO��D���
;&'�A�۴Pդ��#���Pӧ���k4@���A��[|�\2�@z=�����Z~�T:�O��3'�ݱt�B����$v(�x�U��f�6Q��<�c�'�&��3`�j<���'�??�����y�g��=����a���ނ�ݏ]N�Q�E%8|(pC�Ыn�U酆�
��x�ƌL�X8��W�H������fd��4�%}�K ���1i	d'��'(��,��$��{
�3R'� AK�B�Ir
:��T��	$r���PI�7[�:� ǀ��O�d�Xb�����I2����.�s�L9HFQ�Jl��-�c<x
��'n��e��f6p�'�n���л7��ă�'I�>-*O��C�*�&��dƛE4��i2��1X����S��\R�,�t�+5��m��V5!�$FE4^��Շk���t �$UZ��$"Oʡ$�&u���c.��CA�9A#}�2�3}2�A�8��t�>E(ع�d�)\jx����34��@b@
�l�0 U��(�a�(& �HA���a}�ù4�dq�S�H,8-�1-÷��<�s ��K+65�mC7�y��� E�F���i�?<����f�lC�	D$�Eb���T9�d@�*m��1֕|�D��(h����ʢ� 5D�����-0x�h�(��-<-0�+U9�y��L�\�Nd�K�<��bN?|���JD��Pd��M(����L<Q$��.D3l����7(j��q��\xH<��Бy�ah�Ë���@GAR����%�0�p��9�p=�C�7E���5�̤D+�59FRW8����-0���V��,KXr� �M�J�֡k�+˵5�X��DeF9!!��ݢ1H�0H�p�I��φ��`������
�!leZaàY7#|�Mk�th+�'�7`A��q�\�<�'��!B@���)Ǫ?"���C��y	5rtU~�t��#A�	;Ľ�|�K>1��a��(�C'ӡB(r}�s	}<9 b�@"�=��H�n�L��^v���ƨ�!�
|8d���\/�d���{x��[�"?���mF�>��QKU�7�v��+�k5��D��M�;[�\�РnE�pZ6p#!l�+g`�ē�FْP��D�Y_�D��jZ��Ț�세c��I�T���%EW.a+�!e�[�+J�QC���ǱR��X�56�"���x!�$�2I�����˛n����)�Vmj��m�(���ٶ�!	���:e�~r��u�	c��*��;d�|��"��_Ê���ױ!�qs󠓶;���b�`T�Xqr҂��2*M�c�,pR����&,�y����k��h؃�؞{�1��N���O���ˏ�;����߁$�`�Ii{�Ç��P�ǎ�x&*pɒG!$�8 q��#2��iXAe��z.��(���ٕ- �K�O"BK�x���[�<��~��L�
ݪ�l�k�T)ȑa�J�<��$]��x���� 4:��hB�U���$|1ё�A�6��ܤ�z��c!�d4�Ȑ�X�,nNt�4g�!5�~B�ȌzĐ��R#R`|� CX�c=��y�F�^�"-u&�
3C�UA�^UjaybB��t3XAI��tF栣�H�,�O�bWc�g|Jhi7�N�(���r��@,wY��� ��odnDbw�/�la��9$�,�EH�r�ʬ��ߛ@F8 �G��>Qt��.r��*�=����dջAc^��~2�d�SKt���DK`b��EkUg�<Y��R'. =��͇ "⌘rfDG%$�(y����)�p"�)fGp\&?2�x�J���Z$�0��	WD��G���y"*�?Z���-��*��`AVH
��?-H ��m�(��pQF�'�$aKR ��o�ژzAG���T\��DQ	V� iC��T�YU�P�C?ym���a���y
� X)"P�c��zӠ[+��0�`"O�ٰA��T�X�HQ7<9#�"O��Sf�+�D����{�!@"O@�ѷ	U��ؤG�&Ci����"Oi������E�Z*q��"O�yB2B�WG"�;ҏ�#dP<��"OpRǫ ��)2��?�"�"O:���޹>36����ǳ|s����"OƠ�P��Jzpx�TfX��ٰ�"O�}���];B�q0b�rn(���"O���&�\�Q[���ЈC�"9%��"OB(4]nZ�BD��r� `�"O���Ğy�%1��A�<�B5"O�T1��#[*z-���}�mhg"O�Yu �?ID�7L٭qh0aS"O����喃.�tH�CkιP��*�"O�(s��4�ʴ9��x���g�J�<�T@j���em,jL@�#ɏD�<��R�K06tYBL�M�4嫢BX]�<�#)	�.mU�@�z	�]�VDF[�<a�#Y1:O4���&F�e��Hs4�T�<����va�ŪG�M
K%�ٕ@�N�<��]�ZTt���R ���0�C�<�cN��qz���_Zv���O�}�<q�A8TJN��\<a�Z`z%m�t�<Ѱ��[m����>&@�BFx�<YR�ٳs�QR4�&�"$���A�<�6��L]�M��+��;d�=����~�<��of���ўo��A-Z% L!�D_��N���N�C,ess- �!�D�+|�q� S��#D�Tl!򄌲 E 4��.{	>��pB}C!��j.Z�I#*� �.����3�!��X6v�h�)L�)��Y�d`�	U�!�D�6t��� م�G�6�!��ű0��;a&

����,�x�!�$]5l�ȕ�$�_�v T�᥋TLV!�H	8��Ӈ)��@��t� K,{S!�Ј4( �q��;ژ�X ��h�!�$ױy},McuK�9;���G���%�!��� t2��q��dϰ(�����-!��zB@�q�
y�1�P�#2.!��BNH<T/,W"4ӑFϯ�!�$�w��4���0M��q"�L�A!�DP` 40�	ÚO��p�@T�|�!��( ��p��%O�RL$�1�!��_�Q*͒��ԙn<ĳ�lXV�!�Dԕs�8��e�\�}r���"!֫q�!�Ě4\�X�ŭW+sP��"C��<!�H�@�r,2��lT�lQ?(!��ǭr-¸�6/�8s�}� �T)Q!��!o�U
��]�9t�ST�k\!򤛁".�bզ-xzq��N0A�!��7r�@���9l�v����k`!�Ą*^���*^��IR����a9!�D�(h����S>4�����f��v!�ď"9u���eϓ�{�a�7OΙiy!�ʉL���d&թEk��3a*x!��'}x�S��	S�m)V�L"k!��a��s@B�d�8(HӍ�0!!�D>9��l{1��{�d��˷e/!򤚣�������+ngv���(!�d�$�`!��_�������p!򄆞:��Aa�*K�a��T����)�!�� i@����bڎ�c���5W�X�"OJ�$�ӒB	\}�'B�*	�	!�"OJ|zǦE
/�9AbE�`:)��"Ob�e� ��$�獈�a�"OА0�^5p,�`c��12�V1r3"O���T����Pl�֮D*�"O�l���<�v����!_`"@�r"O��u��#i��U1�S&m[D�"O��p�m�Z�Er�[� 3����"O���sm�,�  L� ���"OXi�@I�i=n������)s�"O�
��n]���,ܜ;Mҭ�"O�0֨I�*qL��᫉ 0���R"O(��s��3kb�SVLޞs˞u�3"Oh�1e��1��ɴ.��x���c�"O����ŭ:,��LɉT3 P��"O�����Ԍ~pZp�'jBl4X��F"O��0�. -0n�H�`@Ts�\%��"O�d�%I�f����1QR�s�"Ol)P7�փۊĘaK�*��豀"O�� ���5��бl��G
P� T"O.%Ѧ��xu�j9p�6��"O\�X�/��5�М*�
U�����"O.���#Ú�c�H�<HT�9��"O��[����U��G	������"OPT�h2]\�5�R�� .��u�w"O�p�'�-cH�1e�>0��8�&"O���RI@�jst�P%���$��"O^�����q��Q�&\9�
��`"O��������hU���*=:�"O���%WrQ����?���R"OR�K8ER���Oj��E�B"ON �M��bapE�R8'�1�`"O9��&V1}��ʓ*_	̩��"Ox4��D{
�%�u��jmHe��"O�	A�G<V��ʄ`L4�\�1"O�)K�C3
�X��R�|�"OY�%��J�2�q%N�>r���Q��ޜU=�(�Fk:�a�"�t�#[���CJ�]u���ȓhE��PE��!mش败�8P������W�V(J��3��Y��
��V/n�d��-$ݸ�#��)D�4󖫉{D��6�t��q˥`F�o������8ju:(C�ƀ�b e
=o�X����t�N���	���Iy�l�W"XoZ�]���#�g�F}-�p
T?�C�	zSt��rAQ�S�Ȉ�c�νF�z�Й1�_ I1���ңMU�O�D@��#$.�Q�V��`�	�'7L|��;�-��_����C	��`��<qW�'�gy�L�)�r`�,���akǽ�y���sB�6�q�C!'U�8EסE3iO�шA'!lOL����� ���b��1(��F�' (�؄#��D�	ѿi�����k���ۀB�$"� ��reG�d���f���KV�H9���jp���'EZ!��O�(�� 3��Ӕ1 ���Ra���Цx��\1S�ވ|�'��"}�'޵�E�Tq� `쓗ꊿTL�hP�bVPM�Q�O�4�}���
�UO��ɏFSr40f���1����A�_\�`�ǂ`at 3��1�O��{VO�Fnx1���� �'�p	{D�"��@��[f/w�x����� 41��ѥdήh��ϐJ�V��T"Op`��JOQ!��z��]>1Rx	�FG�	��X!E"���;Sņ�&gd|���imޭ�\K+�8q��?[f�[��-D�l[�¬3`�Yx�he"�oR��Ń�z0��0bC[�?u���C�'{��G��1N�p�hQ��^ܑ�Y��8�mD�J~7�3z�I��F��m��q�3��+� ��Ǚ7a0t��'��",��p�C+o�;��Qq�`vJ����G/\��5U�pA�@����i��15Bˑ3��t����
�y
� �\�Ҏ7���`�&�$6GƉ���)� p!KΟLr#�\:یH����{�혅m@ ���YTޙC���%"7D����	�1vޝ���_&^AN���aY:���0�\�8�u�'��I�	2~Q��I�*��8��<�@�Cb^����+|O�`D�+���A�4=)��S�Ŀ
x@�AF�*_�8���<�H����'���Ԡ�?+u��ِ��O�H���d�)s�\��!�'S4Kf��t̓s��h�P�ȓA��5�����Rƙ#��΋1�q*ܓh�.�=E���!�����|������[ */�D�ȓg.�R��mͬ�a�gQ5�Z�ϓ wZ5���*�)�<�@�4��/��1r)�贅ȓ^ ��HF�9_+�e2h��;�<�'�x��ƭȡaz���2+�\Z� �gU|��'�%��>��^�II�Y{s���v��1$�x�H}0-��r4B㉧k״�pC/G�(��� Y�P�4"=��ӷnPD��a�7�S�}��$ۥlX�'����e���C�P�E�� �0a���b�5*�7M�0+� �q��S���)�禅�lԇA���,
�Mg���� 8\O�9��-S���̥]`���b^_7�y�S;|�������q�
�"��y��O:{��p牿�6�;���$՘'�2�� �%T[q��	y��)+v�%p�Lۜ7`�a)��%��Jǌ��xr�'.�I!�+�S�n���\�6piʂ�=}��W�*n��d�9*�v�'W�条U8	�$ϿP�
8C��K��B㉇x�YW�J�!�q��QPi�t�ǁ�7w�pN���I;n��q�v�<�s�������ɳG ȋ2NI�G�'��㇠Ɉ5DA�'��lpt�_�0��:g(��()�)O� fHܠ^FH��On
���U��&[��)s��'/��'��y�"�$*����~�։� ?;�)��Ҽ(6Hq�%�����K�b�^�<����Fs\혗 �-,�t���mQ�Y�d4A�>��A[�����ɮ�<9k��d*n��5 1xT�B�I�O�XDc����iBt%K�[\H۔��63��)zP�'�N��T�X�_�P��SbF�ClMH�_�Z��#��2An�:�Q!"�'4$�Y7j���ȓ6�H`t͘5����U-IV��<�u�D�}L^�`��I�9���{a�%
f�QI�(P�!�6Z����
eWF<�c�"\�L`�E�$���(��ɵ�൒��qǸ��KR/�$C�I%w*F$yu���)��d��U�yn�B�ɑ@��4�q�<NX������v|�B�I?n���e���d=�P���&<r�B�	&	 �haF&_(u3�r��4��B䉳'0|pz&k�ь�B�n�#jw�B�	f��p� ȫIYZɰ�۳s>jB�Il���w�-h8����,)�BB��;���p�!��q��Q�[rnB�I�u���R)I��| ��	R
@�?��
٤%w.b?�"$0 	��Ď�Id4�:T0�!�D�P��y��I-Wݢ1��R���-I`�r�VM�)ҧ�f�QO�^�yi���a��Ȅ�NBD�+�$Xl�i���F��T��XC �zc̋�W�-��*�Ԇ�W̓n��a��Q�h��`�eY�l^����	h9��'�ɔD2���L�5_!���L�Y��Ti3O6Q�E"��J����䆈0:H��qBRGz<"�)C�#�Q�� ��U�+0yX��'�6 	�F�3?4`	!�0b$���m����CVH<a&
�*F8ac�^;]��=�/s?!��[u���ꇯ�O�!#�&���!��D�<1@a��G�~ æ�Z �yҮ����&
� ���pjچ�?A��K8m��
b��	������RF&�%��Q�
7*4�a�Ad�H��/�O����/şS|�|�GY�PE�uA�Ж5ܔ�Bg�6�?D��E� �-,Ol��H[.ZnU���W�
Q�@ؐ�	?`����!$m2EȅUt�C�W�eS`h� f�`�p�r����Y���p��@��*�#Ohz �'�ڐ�-T��D��|�8��)���O��� �C�=�F��fhK" �b\��'�U�F��`�,|i�KNEFQ!��i& $8F/B�d���qD���'f��O� ��he�&n�tC0��1�]�P@�ȓ:p"ɥ@��<�HÁ�%�'���Q�����y�K�%,���r�n�$$]XĊ�p?	�"X.t����f���n^v��e1j��pc0D� ��S5�2��F�J�$�{��1D��ŭ��B�n A �H�.�8Ċp	/D�ȹ7!\$��a�gㆥ�����h9D��۠-L.y����	܄��3D��"�ڍ=DT4���� ��3�)$D��P$��9&ʝ�Fj�)jpn&D�ȁE+�e���EyH��#e�2D��"�
�5�vKƍ��GȰ����7D���PbI�^��|�s�;,`d/>D���t���J[r�@.Mf@	C:D���'��w�|�2��@�Q2��7 9D���FbBA� ��۔>� �2�d6D�r0� 	(D�{A�/o�8�:T�2D���0bI�b� 8���$��-Y1�/D����Ձ!�`js���y�D%��7D����b	# �iv����#P��yB߽o�A��h�8�c`��y2�Ͱ�v�����ݢ�F\��y���]�|��! Aj�t{��J��y��<C��B�-˟Dݘ`�휨�ybm&�P�Fʀ�1g��`�@�3�y���{�p0�q��!����W���y�J��β$C ��t��'�0�y�c��b����A�RT��CN�%�y«�7tn"��@�[6����Gȿ�y��7Q��#��h��vh˒�y��^��N��&�3�)�E�(�y�F�X�d]�A��k��3N� �y
�S�v�(�JW��Rd�f�Ѧ�y�*�x!���ɒ�L�8��.�yr+P!!��M��H=mLp���yr��(J�`�	W�2pڊU�f�2�y"i�&ߨ���(����= �@K	�yRX;��-0tmo�D���*L��y�(��gP$\���W�2��\��'ٞ�y*� �6��E��F햙��g?�yR�1��ᬚ96�X�sWA��y�D�U/.m�+�*����N4�yoR�n�Y�l�	EFO�e�X�R�' �����іI�������3
�'�ZD�R&�9{%�9���ׇznX���'�
Þ�J�x\)�.��{Z"�:�' ���܃&`��).E�t�L���'��I����/"D8qF9��5��'�,I�@%���F�*;s�4q�'$�ya��Q8F�0�5I�"ff`��"qT�4��V�����SB��	/A��y���*� ����U
N�:T|EFx����1i���x�f��Y]�5��H�H�!�䆲y�^��ɘH6�,��d��g/��%�S�O^`�se�@�b�@��1$d���'�0<�!uf�P��eD5C�>!��IÉ��9�5�*^������L&D�4��O�ӧ���L�閱(Q���.�-R1Ξ���A������ݻćٸ*��`EW8>=#Ճ��e���#�'Pv����O�)�\�"}���J�xI�˝�?�l��7ʂ/atܨ�O���v����?ӧ�)�)Y�lU%���=P\ �O�&s����<��߶�y2��m�OA���B�N6~e��0c�ߥp��`�Ĺ<�2���y��:�g?�����N��	�V(�;��(�O�t~�p���=�O�剱舘b�k�jEq��$;���ɩ�D7�3�)�'�a��h:.k2!8�X 2K0$�qkQ���뢖x�O���G�� �x{0C�xȄ� ���:omԉ�����0/�p}�f݈M@a��@���4��'Ǡ/ۜpp��!A�=�Z�x���Ó,�&>	֧�i�����֭lcJ$:Să�gy�듿~���3��E��'�{�Γ�>%S��"�3�'�>�����%	�t�h��9!�/^�J*�ĉBj������D��R��񢴂(����0|���ޡ3F$�
tɈ%;��lх�A-_j�2sd2?Ѳ+��0|��i1;Vi0�KA�q�4ܑb심K���CՆ�M�%.�;S�y�ç3�b] &cC�`N�u�'I�$f�h�2�	���M���;N�&͘�LP���Tl�F�Oܤu��OE�Y8�-K%�$3W�9��m�~�V`��c�2TC�E:cߓ�~��I�Sm,	p�P�\q��re�K��v��# �O�?�("K[�>��m���K�A��ݠ���"���Dכ��	V�,[�{%"��9�!��0� x{�Z,=B��3o��#�!�dM71���&Mn&u�G-�'|�!�$��q6�l�!g�2v<�L�1I�:�!��:����"P"4A�
S�O|!�p%�yG([4p����f�-_!�$M
-�������B�U
b�}��"O`]����a�L��3LE��W"O���L٤_�.m!�+A
[2� B�"O��A��n�.AYGJ�8dya��"Oȝ��ξl�<`:S�J�>i��cf"O쀨f�0D��`i���iM6��"O̥bC�M5��	e<5R"(T"O���&˂Pbia�x)*-�"O��3��=Tnd����Zj�Pkg"O �"��F�^ł�@�lK����"Oj�Q�$ѐw�(�8�"�iK���"O�ȵ/�4C3���a�'	=fh�"OlF�=N8�a��ю|~��"OZ�+q�Z�)�&,�2_d�9V"Ox�ÑÍ�j�Bc��4{:J�kF"O:刁ɘ;8,���*�8.Xd�g"Oѣ��^�fq�p��	^]HM��"OE��9�T��&�Z�unD �"O�KRB�$w�jh���ڴS�|��c"OZ�K����{�8�'�,%�ػ�"O��
��l!�s�עt8�p"OP����͉&��rR�Ξl� ��"ORHñ�߷JŨ�5Ér�&@�$"O�9�`Ӫ�ʁ�s���q1�"OԽ�f���L��QQ0�� Rč��"O�Q*�%pJ����� �BP"O@�j��M�r��i�.V�%v��"O��q�a  2�vĊ`�M�2SPm� "O��BCQ��8�V@]�&�*�г"O:���A�/��
wE�{vظ�"O�-8��[�[�����hR� a ]��"O6�Y�f��B�@�;BN�\�p�G"OPk����b��
��%�"O�چ�U�*�����&��=�R"O�Ȋ����^N�18u�V'M��`"O��K�oK����Z!c�'Z���"O����� O��bV�U�E"Od�r�x�����L�I��l�c"O�L�t�߀`�Āh���p� l�E"Od��Q��V&PCB�?��X�e"O�z��:I�l�C�J�UAV�zv"O�4��+I�;��ĥ��u>b43"O��1�O�{Ylu���U?`��"O��rI�h��Y��A�K7��:�"On��*����;K�	eSP\��"O��˞�jO��T)	"
;�ɂU"O ��d�"qrNH�C��-�H��e"O� `D���R�A)�A���Y�"OLMːN��qARɠ"� �9]耹�"O�l��	�7mRp�u�Y�GD�5��"OBE���6�����'8B��iv"O��K���G��Q�3HJ�C�%�S"ON�ò�>P����D'O'l��["O~�@�DI�E4�GC�@��4Y&"O~�D�Ρ:`Ѐ	��R��h��"OЁ�҄Yz�%���J�]C�$�G"O�� W��]0+��0+��b"O��z� ݫ%(��4�_4\N�B"O&	���J����C皭�!�"O�a��T�Vt�G��$�x��"O5[�h��65�u�� :T�
�"OP��pj6�\qA��ȸT���q"O�	�:�X�*V�F�U�����"O���#��(+g0���F���ģ"O�l2F�+H�(9" \?��t"O���vD-��Ts���)�d�C�"O6�!�@���FDg4���"Oz�#���υ�A��ɓ��'O!�Y�D�����H��H�s����!�H r����Ո1����c �;=�!���3\K��[�Eot��(�
"!��B��q2�Ot�l�3�eS�!�$�$/J.ͩ���/�N���%	!��.mL��b���E�Ā�4�!�[&]��I��o�;I�z���.ہ?�!��F� �gkC�laf���,ݰ�!򄂑o����'�F�d'�Q��K�*_k!�$_�w- �׫|�>�[�j	�^�!�U"Zw.����߭b��!:���&�!�d�)��P�B��e��L�]�!�$V�
+j�a�|4�D�'K�!��>F�r8��֟/o�%!s�S�p�!��(:&X�SE@%[���$Ι1�!�$' CԡgulN0���?L�!��Q"��"W'fQ�4q"JBK�!���������j9P��U�	�cs!�d�%�&h��#�o)p�
�B�6!�Z>J��uc���/=�ȫŌ��R1!��X�� ǥ	*��a�X0.!�ďM� yZ���Z-�SeѾ*!�D�GP��x��W�O�(Uy�dX�g�!�D��Q����j�=�Zz�i��	�!���$7~��'�/:�=K�E^6n�!��w8��GJ�L
m�EF��!�ڭh*R�#�ǊZ�P��
�!��*D4z��A�C+��c�\�Z�!�䖬_���6�ؾ`�nUAw��n!�$B��� Jve��w>R8��
;!�i�2���D��8'8�C��4!��Kg���P�Hq)���C�<�Pyr�-�{�.���x���]:�y���#,&��t�sj_)���'q(��&�^h���BfA.e�u��'��-�5JϚ��EЕ�a :���'y�,s&)
�r� ����ӌ���'*�#&Oȉb� �JӢ��D����'������P�l�0����N�Q!�'�tC����4#pBwy��z�'TƤ��"	�+~�����l}�ժ�'^��C2��U�)�ի�6?�e��'�h��iW+'&VyXT�F겸���� �`x����$-�=	��1�p"O�D���H��T���~b��""O@���ψ�S�% we��mk�|�"O��竑'���Z�@�
�$`�0"O��	p%ى�xzuC
�SS*���"O�(�V�L:xS�q5�A66�p"OD�ca���J���Eoɺ2RՓ$"O��e@V�g>`놏!nC>�a"O�j��Y�8��XNK*(8"��2"O�maem޽|vP@쎳'��D"Ob�"�A�`��z��֐�"O�E��:WJ1��	ݮA@"OH(�� A_����� ���3"O^!Ja<_�Ly��HH�l�(a�B"O~��gQ�漹�̗(�
���"OƔySj��m��:�	!�n��5"O 肂��g\A��^	�δ��"O �J�%��x{*RDS:	��'"O�E��c�	R��8k��Ƣ�4M(�"O�Aɷ�e5�5�u ·.���Z�"O��� �R?��Iwo�m�*��"O��H!�ݷ_�XK���
��5"Oz��4L�:J�D�C�M�<4&|0۴"O�Mcŋ�4cѾYG� (_�$iU"O0��J�Ex�� !L�x .剗"O.��v�K�>o>y��T�� ��"O�5D�5Y�b]qJGw�H��u"O��0���0DDK���e5~��"Of�C��  �&�kD�ʒ (���r"O6�R-�8j�d�;���r�"O�d겉�sJ4���R kK�\�"O�Ik��&?��ȳV��q���#"Od5Z�*C>J�����7E`P5�B"OPC�`q���BFA@���"O��K�N�_�,FS-U�"O� BQ�B�,ct��E��##"�!�"O��gB�2�2	����;#4���"O٣���,�4��FØ�v���{�'fX0PTmcY�}�Q� �g����'@����J�A�P��9-F
�ʓnHpV(�Wp�p&�94zԅȓw�Ղ3���h�Sp�X�(�t�ȓ	������}�ҹ��j��.�R �ȓ{z�Y+@���[�J
���W����ȓ��Ѹe��*AϚ)��o�A�� �ȓ~�a��:+�TE���L�0��X����'G�=1*�s�LW	#o(pa4D�x�7"�!Ҟ#�Δ�V� D���,D� rEH/`��]�5%Ѡt�mk#*D��!.-Ʃ��&�8�v\�p'&D��hש|�r$��,�o�yرe)D���e���/X*�4�I�l���c�%D���C+��Q3.!�6჏WA��(a�$D��R��ϰ)�,41B�α�p��$D����
�2Ek�Xi#l�7'H�L<D�@��pm�tS7��!;tY�A�4D�T���Ϡ_&�Q�
�%x�AhT�2D���Dd�
�=S`-J�D����3D�@)�"h=��%Up�4Bu�;D�(2�e2m��F&��5K�,D��J%�G�[��JFe�6�
}z�-*D��"�D�2�dY
Y�e�0a<D�t@ K�b��#�Hؓvx�z�<D�<����
�"�"�=FL���,-D�� 6��f��0���˲i׊��5"O�L��G�>zܪU��.Α#i0��U"O���A�,<��dR7q2�h�"O$���+K%>�[��g����@"O�$���Ġ-��QrA�f�J�x5"O�-x'ܺ,�PI��gD44yd���"O`)�LG�1�&�as��ah�U�2"Orm� ��8
~�0Zá��[�"OF�i���8$��IRAO(TP���"O"dĦ	�|��/�"<-��"O���e@�!>^�X-�"8�A"f"O�L� ��!eln�"Gl�k �X�#"O����g�3��`�u��=�*��P"O�!(����]P���T 9L�0�"O���cH>w+͌K)8��d@O�<A�   ��   K  �  w  �  <+  �6  A  0J  FS  �\  -i  �q  �w  [~  ��  �  *�  n�  ��  �  ;�  ��  ̶  �  a�  ��  ��  5�  	�  ��  ��  l�  8�  { �	 � Y � �% �+  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,͓�hO?�zP'���|��6E%V�ၖN'D��At��j��KC !sx��rh8D�@+�-�65b��@��B��`8D��S�;���!%�*��u���6򓑨�E�3#νw;@R$��Kv��U�'މ'<�m��.[&�9�BM�3�ڴ��'@�X1/�U��yk�H�+Y�8仈��?�S�T�ݚ���t��e/��� �(O��d��%۰��w��
K����d�ҢB�䛿�X⟢}�wi٪M,�Ad`�,M�<Xq��N�<I-�� �J��	f[p�Ё.D/����#�HOP��x0��0*��`�2准N��A�!8�O��hG��:�޽`�y�fC�<f���?��� �S��H�eB��B�2Q��!̟C��0E���3W\��"j^.ܤ�r�S���ĉ�t�f\:%m�8/���J�#��xb�Ob�>7M1?�cɓ�%��H��k�a���ç �\�<�2��*�L��(� �&�cg(^�<q��(4`�l\���`�e�Rx��Gx��
	N�`
a��j� ��5ㆳ��'^(�EyJ?�ІI͂X*q{ C�5,2@���'D�p���;a�h��A�&3d�ͩ3G2D����iZ27R�1��e�'����.D��(W�Ϩ��A!���(A4�IqE���`��	b}��K�kD��i��̠:�D���eգ�p=ٴ��C�:a�T�\*͂��D�CB����	�'��rF�U���j@	�[$�� �{��']�O�Oe�A��M�G�&��ӳ����'�ў�}� �0�FF'����k��W�L!��O~c�h�㉄�\���@��}2u#����k���'�a}Re�"~"��@K�J��A�W$bU����ɾ���m::MbGh �Szn�c�S�azR�D[�ux�%DYT zQBgeQ;aY!�d�>@��xt�[<0�a�I�u�����'����`F�;֢	*��E�ՂA,D���O\6���n��e��,rgJ?D��!#C��f\ک0��0JR�l��2$��SF�]"'�ZE��Y��)3cݨ�yↈ%O�BIzv�[J����ع�y�[�V�P1K�*B�%��5�&OO��y2m��p������]6 ����Eo��'+ўb>ّ0���%.E��)69MR��I6D����#�
T�^Mj��H��&���2D�p��(k�d�ree	�� 0� 3D�܈SB�#5s�#��G1sư�ٗ�2D�x,���Xf�p|�����I>����+�Yվ� 	��b�� oI*��B��+w��9�P.(�4��&p��b� E{J|:���J�i��!��/�r��W�<��]�V�L*SLU�.^-�T�S�<��E�E�̝
�B�/YY��()M�<�Ơ#q'~Pv˨V��H��
OH<���֑.�*ԀR�\U#&��S��%��{R��Y2�[g�R:�}j��	�>a{b�'(��R�k��'w[(�kÎ;) 2`���\1�cg] _�	@���3J/��G}�ŕj�O�� ���Y��A,^o�`k��d?O�4��O ,�ظO�"Z��h�u^��F{Zw5�O̔��"R�.((Ԩݭ4�93�"O�y�+�_���Z��ع"�!4T������9��xFz���7�����m� T����?��D֏&˖�G	ؐЮM�TNON�<qwo�;8T���l�O��ts��G�<a�y$��!U��#L��רM��y"�ށ)�J��K���W�Q��yBF��v��TIU)�1I_ ��!�3�?I	�'p����I�;��1�H^�d�L�+ÓJ���35�4#�SJ J(y�'O6D�8S�&O��d�$R� 	];��3?��)§8�����֫=eH��� Qf��|��&0&	#c�!j|�`��M��VV���hO�>�� &��A�D(%�"�i$"D��$�I�^�F����5�`<hu <D� �1���;�(��
Æjv���q�:D��	�j��o �H�� ��'`:4��l-D���@�7َ��4�ʒ��x�Nl�p��ɋ3����N�(W{� ��K"X���Dv�"o �A�D�[��F2F���[+yh<�c,A0 =���"���.��d�D�<Y�a%�!�ËYzպtZ7�Bx�<1��I<i�i�7@�����qx�|�'�\̀dW�E�����(�¸��'���C�]7`�r@�$�s��̓�'N�H�j�0
�fd)�kxTh��'u�s@M�4q�z���=n���'"LQh��/@�$�*ci	N y��'���)W��L�jS����W����D#�O,$��k�61��!����5@D0qr�'��D�E!�?`����%Ќ7.j�&#*D��Kr�&t��m�6!س�Z ���-D��F釋r-�XY����t�9t�%D�8R]jD�6h�@N� �	�$�0��)� 2����A ��)$)2+ �H�"O\3�ɕ�v��eqVH���;�"O���*I�N�,pڐHX�~� d�@"O���h@� w8��&�'���s�"O
	X�o�9�H����ڤ��'��Dy��)_�a�R��R��/&��a� ,,OТ<yu��2t�pie�J2+9�D�"�	X�<�O|(�G�T�]�<����LSGv�r��d`�<�>ͧO.�	�\qh-�G��~�@�a�6�j���'Ԝ��N6p���'�Ÿ}���{�\�4G{�'Y>\�ǫ�;�>p���6�@݇�#n�t��O;�A�$ь�6��=9�4�O�O��iQw�ό2���t.��4�I�'�����5Z�F�RD��4>!�PY��-O�9 !��i���)c�74a×��_���O�l�S#N��k ��`��S�	�t���'4R=�B�I	\�r8��j.Nl����",O4����@e1��k1��:-��82"O`��A��I�*$C�E=e�htqs"O��A��&a��CT%��88�F"OX��=W�f<If�ّ�0�Y��>I	�d� �[fM��(0���S�P�����py"�Y�`�{���2f�� �&/^��y� ݤ:��A#��S��<B�R��y�d��g�Bs`�}v�9�
�y�k  <�B�!�L��8[�%в�y��E�w{��@�	#qJ]�T-�-�y�Ǌ$�N���*���� D��<�yB�LTn�P�I�H�q��Bĳ�yb`p$Fu�B�G�;�<@����/�y��O�6�ԧǈ,���R�E2�y"�Q-ntt����Qu^�:B�Q��y�
�(мu�Q�БG��y�Q !�yn[6�& P�m�?��Y�����y�̿BL����[)g�P0�r!�'T4�����7C�=��&��F�A�
�'TH�pB�/��@"�l����<��gӲv�
|H��և[} uI�O�<YG鄊}���z��G\����T�<y&+3j�I�,��|0���q��f�<�a���jŇD�K;�l�3�]�<YQ
�|�f<!䪀~1���Ä@Z�<�&�G15��hD�ėo^�.'T���d��"u�44"��I2R_Π���,D�p���^��R&!�3%vR��)D�0�.R3n�>�x��C�&w�#t.(D��97�eZ,$���L��0�R*D����/�����c�%
�C.���:D� *�&�څ?.n�I2�Z�is�C�I�,1��8��9cf���p&�C��(C!6q��'���c�TC�IVڝ�BEpE�V6��#�"Ojt���mTh� b����!��"O<�;�"\�� `���r�~��"OF�3a?9+�	�P�+j�HM	�"O����$������J	D���"OD�5�i�"�1t�ܱ(nHt"Op�[����th���$�gꢄv"O>m����(�h��e��?b2tP�"O�� !$9p�3c8{�T4��"O�!�#��/b������
��}C""O���QA����12���2�"Ol�CkŅ �'+�!��A	3"O�1S���(7:Id ���>Y{�"O� �!bq�F�&(������j�ӥ"O~�y�۵*D���4n�
����"O�P`7�?_��\y@�E
��� "O��Qf���@����\24^8��"O(t�vnÖhPJ�b���$8 �8��'���'1��'6b�'o��'U��'��4)6o	(<@�R�o��Ix���'���'��'���'���'���'�h!�UA�(n ��r�g/�P��' �'*B�'3B�';��'a��'-&!��-��BIZ��� cwf!��'��'w��'Y��'�R�'jR�'��L)���d��LɁ���y���RQ�'�B�'J��'q2�'���'���'�H�r%M^1D���ځfÍ��%�S�'��'<�'i��'��'�2�'� ��'~� ���d	
�'���'��'��'g��'���'�v�s�\|ݒ|Y��]S�]�s�'���'���'N�'���'"�'�\c���2����ō�/@$HE���'��'�B�'���'@��'���'D��2ō�c������H���$�'���'Ur�'ub�'u��'���'��݊C�]�:>j��AI�� -�!�'2�'+��'e��'b�'���'��*� ~'$�b3b
)a�� %�' ��'8�'�R�'1R�'���'.�;���	q�M*�š5,��8��'��'b��'R�'�b*e�����O�-!��rP@���״&��H���Ry�'��)�3?�C�i���늣s�~��u��)gU�5`U�'���ʦQ�?��<)�)�@�9QM�/�x	��+���Ȓ��?a��Ǡ�M�O|擰��J?͹4��>R���E��:Di�B6����'��>i��ƚ=}bI)�`76�q���
�Msv.@a̓��O6=�6��t���CIHak�e��L�U�vh�O��$v� ֧�O����'�i��$�;,�ˑ�T\F)	��\W��Dc�B� �ȣ=�'�?��Ҝ*�4�0�ϒRu�my�N�<�*OH�OʸnZ
G�b����[�7K4C��Ɠ���	u@Q���I�4���<1�O��F�����A�"�j�	ӗ����<Z�4�+擼["�K�@��h^��B��3w��AQ�DTy"P���)��<�M�?�战$�<0Ѽ�4e��<y�i��؉�O(qn�S��|r�a�C-T����M�u�h�bR&��<9��?��j[>��ٴ��D~>��'qԎLs���;E�2E�7��P����O�A��1OX��|j�'�?����?���h
����(Ĳ4�h|��h�.{4��,O��oZ2h�t��	���	�?���zy�L.T�C���>]!�!N�f����?)����|����?�3"�q��Z��U��P�'�W=g�l@����f~�O��z�D��I�Mj�'��I�r�� ��%F��l�yL�7����d�禍���K��4X ��A�$1 �j�Wb#VCf9��8�MK�Rk�>Y��?a��0�!��^�hLk���g�D<�%h^��M��O�q�������>�	��H���7x���0��$&�J�c5O����Ov���O����O��?��BIҘq� �;���6sv$`��Nퟀ�����ڴxX<��O��6� �$�'u��P%ĄJ�4��/��B���O��$�O󉂅4 T7--?�;X�Fܡ�A'.f�#£ö \(}��mF��?!�B/��<���?q��?���,E�u;祙p��|��ڲdΔ0����	צ
OV�t���������ec��0���+J��V�p0�5w���	�����Or����)�	7�9��nےq0T� �I�_����ě�y���'����ӟ�ç�|ro̅ǀMj�)ʅ�h8�U] �"�'��'�ʟ�B��<16�i��
GL)Xn̩:�A��U�x�
f
J?p���'�d6m�ON˓�?� P���ɡ��{��ֽ6�r�bB�T�;��I��L��OO�Γ�?Y���~o��)T��򄂮0b�����#ZM2Z�`�۟'��	��y�� ֟�I��t��ß�ӡG�lD(�C.�-�&i��]1��ݴy[hu����?�����'�����;[�b�i� �&=��t26a��q�Z0�I��H&��SџT��/��dm��<�f�Rpn����L�.|R��A�<	�捍Hz��d�����?�P`�ݑ���� ���@��DkM$O�<lZEa�H������I�tĶ���-D,z���v� BP�?�6T�4�I���'�"�Z�q�GV<i�R���Gy��y�ܥH�����0�J~����O�0���>L}#r%Z�*�yX�T�5 �?����?Q��?H~�pj���?��J����6����OS|�,��j���P�r�'�|R�yG�(��-�U啉K��mz�)T;vr�'���'%F�J#�ir��Ozk���(vk�Y�\-R����0
�R�@j�alX��O>Q)O�?��(\�E͋>J�,e�u��S~r�|�H,����OF���Oz�?�+�`8�\�ڥ&��b�!t�[)��$�O���/��ɞ o�pY��C\�R��i�v�!%,d���x�8��'9>( L?O>(O���ڟTQb���\�RR��O����O����O�)�<���iu|l ��'=��qL&4ޞ؂�䔚eUx���'��6M;�I3��$�O����O$��#��4A�����B��������3,X6�;?��+�C���	�?��ɿ� r�*�A\'I�p0�I�c�X,�0O��D�O8���O��D�On��&���V(!yE`�f
(��$9�� �
�O>��ΦQsv�_y�,`�h�O���� ��U�ƁٴF�y�<б%+�D�OT���O��ڂ�nӐ�ǟ@1U��U�0a�ej��hЧ	,�R��'\P��I�nw���jy�O_���'��J̪zG����&�W�Ԁ{C�8(���'=�I��M{����?���?9)��k�T4�De�����3OJ�D�U}��'Қ|�OIr��M�H�Ҧ:D�A�(��8pش��Xy�[�Op��ԇ�?A�*�O��x&>O�cv�Bv���s�ܸT��8��O��D�O���O��OpY�%�<!6�i�4�b
�`�B*Ef�4����vE
�/����M+L>��4���͟��s�Q�?=T� )��^򽲃a��H�ɺ��o��<�N�&����'[�|����P���N6yf<��'�	���
#�ş��	ԟD�����ӭH����V�.̱C�y��
�4Z2��4���?���*���?�����wC�=��)�L���Ųq<�7�'�|�O���'��M�g�i��d�.�4�QB"D�"��=�7̟�t��dS?$Z�
�~���O\��|J��dY�^�k��R�Y�ԭ����?����?q,O��l�J~ȍ�	���I�,�c���	[���p�P�G�f�%���I�����ON��?��S'p*�uh�R�NqSSJ��P	�$�Or!��K�)v��Y���<��'j���$�
�?YH��F��`�m�2?�;�(�k�<�E
��2�ܭ���V�?рM��mP��?��i��"��'Tb.|Ө��]��rP`�a���c�l,��؟��	��p1`M���i�'�D�Yv'[@n��/��	I�ˑh���;wc����6���Hp�Q�̓C�(i�a�C ���'�\7�"6��Ob�D0���+،8�����{LX�"mJ[�Ԑ�O����O��O1�P�A�a�F�B����$<lV��K�8Vā9�(�<I�+@,><����"����dL�D \�x���(M�h��]�ma|�D}Ӻ$����O�Y�f�S�G]r�C�{.��+�O�qm�l�I���\����L�UG@N��a�����Y��{j�%lY~�g��?Gx��'��)���Vī-��,�#τ>r�b�I�,f�x�z��+�X�a�%H��9����1݂��̃0ZX)"tK��U��\�sDT�~�v	���#r^���Iv��d�S$T�k�[��P�@ΘDc�l�PLǁe�!A��Z"�\�u�����WMc�e�aCɒPK����NI��A`qNP R��Q� 
��%���ڤl�<U��	�X��s+��S���!�LUN��p�	��1��H�%��4��%Ad*ǰ0�������E&R��˔�������<�I�8_t�ɯO���?i�'��j�I��i���tL�BٴD�ݴ��Ca�x�H>���?y��k@O�(�lx�`��'�mAԫ�m���/B�x�O ˓�?�K>��2��Z"��jh"�Y�EO:4H���'�J��0�|��'�r�'{剃S�h���NV�u�!��d#(Q�D�F����<�����?mdӲɳ���1���!t���
e@�W��O����O���<���UX���4p��PQ�Q�}�|�S��ן;�V^���Iz��ʟ��	�|*�I�u����ƃT�dk���N�#H�R�ةOj���OZ���<)��#��̟��g�-�ޑ
C��U&���V�ҍ�M������?��=�p�����gz��2�%	�J���	���\�7m�O���<�wM�3IB����,�	�?i	R	�yo�� ����0�r��lƛ�ē�?9�1���Ex�֟�����	�c�$�&ɖ(8��ұi�剡0����4�?���?1���i���G#�2r�V(
��y��z�}�j���O�����O~�O��>U@�.WJ|A�E燥Sɤ��v�y�Hx0�J_撚�I��	�?��O�˓r�M��@k���p@��;Q��ɩV�if �{r�D$�S���P�ℹJ�R�P��xy��t!	��M���?���r�� ��T�̔'dr�O���C�4<�̪�#�P�d�s�i��'a���e&��O����O�-�3hZ�t:,��L
r�]�悙��I��%(��Z�O���?IL>�1;5Pe"C le��BS�í)��'τ9냖|��'�b�'�	6f��+��$qJ���N;���7�H�ē�?1���?�,O���?���� &�j����1���1�Ai�N�Ļ<!��?������G�%ͧ:���ȣɔ�(�Dȗ��xb��'���'�S����C���'�fx�X�M�JTJ���
}ڞqI�h�>	��?������#`(y$>� &˚�`�V��W	^�xo( 1�#E��M���?A(O0�D�|*����S	�.� ���NB�(���=D/6��O�˓�?��@@��	�Ob���k,��Hw
ݓ3�>n��h��01�'�"V��A�!�Ӻ��L$kE�d"v��R@�TB}��'p-�p�'��'��O��i��:�ϋ� �*�e-G�1��}�Z�D�<��hW^��ħ"� ��o��q��� ��|�2�o�U���*��6��O4�韶%��s��Y�Ƒ/#.�a�X"����F|Ӵ���O����O����9O��$P��YS���>ۂ����1kO��m����П�k3�I����|���~R"�mҪ�M��aǦ�C�j�8�M�����f8�s��������m�*a0��ۚ?���$Y�a�t\�޴�?�B�7I������'�Y�d0� ,� �MD�j�& VK"��3�i��	����'���'��V�в�������1�Z(%�*I<	��?!�����O��S�Y��d+%�ڎE�bܣ�>�F7m�O>ʓ�?Y�����O�H��ÿ?Y0֨�%�8p°�Y��EjZ�M����?Q�"�'k剄A�r6�D_ y҄[�t��hQ����U��'�BX�$��'!���O��苁9l�a����z�@5�bA�$ �6�%�Iȟ��'&��[M<)����v�
�H�BF�g�.�f���=��ҟ̔'�*@�S-;��O�������#,V��-% �⤻i5�	����`��\�s��X
%aP����H�t��/��47�<q!
��L�~���j����8�O��+�6��$Ԁ[��+��~����O����Oj��O��	f�ܴ>$4�BNN4���H�"_�xdo�4aw�=��Ɵ��Iɟ��Syʟ46JE�vX�D`���k߸hz㋚q}�ݤ�O1���M�<ĬЉЄ��/��j����̑զ5�	͟,���Iː٩�Oxʓ�?)�'EhmytU$/��4bB��0^L��c۴��g�T!�S�D�'��'Z3CE�/j�$�1G�0�1��`Ӫ�d]��-�'d��|�'eZc0�� �hCr���ũ`����O��X�?OF���O�$�O��D�<�1�B�x���d�(�Ra�fl�~�@��W�d�'j�\�`������I�]jt{��0nN���P�U��-	"�f������	ß��yR�T�s���%4u�BA"LC��3g�6ͣ<y������O*���O�� Q;O,h����7k:y���
W^��#�L{}B�'���'e�I�ڝY�������X��Y�R�B�׼�X�J�>^�Yo��'��'��	����Mcc#�]縸)G���{l��a������ßP�'e@鸑l�~����?i���z�h�F���B�a
�h��I��Z��I�D�ɾz�Db>�E*k��1c T)��N-,����ꦉ�'_�-c�"m�&�D�O"��柪�էu��G�{��1�fD�v�رF��M���?A����<���d$��K��!�����Ol�7-�(�N�o���\�I۟�ӗ���<��O�y�d툱@ %zLqɰAN㛶�J��y��'�	|���?�eiN4n�聕��/`m�}3Ń_jǛ��'��'ζ�b�>�-O^�䧟�E�x��]Xd� 
�8H%�wӤʓ�?��#�<�O/2�' �E�	&�2H �o�~�0��h�4Z�D7�O"�����R}�Y����{y���5�'�(T��(s�z�ص�����\�Ÿ'q�'�S� IQ�<�٢rOށ@Jʄ���I3��P۫O��?9.O��OZ�$� ��Lz4ʛ5�؝qSH?�Q�;O����OV�d�O��<ѴI�+2�B�<UH�9�Ж=Hh�`%���W�h�IBy�'��'a�|8�'r�������]��S�Ȗ
���
 $z�R�$�O����O������RT?-�	��p#5n�+t|p&�YR8*�޴�?9*Ox���M���d̓��iyr�!�hS�2������IA*�Bݴ�?����dٵ	8%>����?�!���a��50$��:��)�	�OZ���O�!����A�*�3��5�2�Z���P��T���'�<<	�z�.��O��OX��Bh�eK� <��C�Y�(8�nȟ���?�:<��G�Ib���OZ��j��f���D&-Ω�R�i���"�w�����O�������&�|���U�L�	����K.�X��&�W�	�}����t��^���?!FΫK��j�Kì&A�E��+@G���'���'�J)x��(��Od�$��x�N�e�H7��[�:��@Jl�ғO�a�4O��ş|�I៸�1��	(U� h2����N �!,�5�M�2�=Xxb�'y��|Zc �L����dI"G�ľk���Y�O�́q���OV���O�˓qꜹ��̕��<lȕl�����5�ԫϱO��'���O��
���1�SR8u�x��3������ ;O.��?9��?�,O�5;2*R�|ZV/�	?(b��D����N}�'y2�|�'x�n�yb�D*����NY�F
�Jծ��H��?����?�.O�u��H\A�S�0S�4H0��)��(�w�����A�4�?�M>)���?i��Y��?�H�����I�j�뤣�"D�="�Igӆ�D�OvʓJm�E�Ԕ��'���Ɖ�i:}�#E[�*��Q�%�>Q�rO��d�Ov�Ik�O��O>�� 8Qf�
G#ۮ3ل$yH
7BZv6�<�V�+)Q��d�~����R%��sԏ�:��E��'R  �jPJ"d���D�OJt� G�OF�O��>9;eo�;���ے�P��<�a��1�g���e���@�	�?UB�}o�'�8p�Ǜ&�HY����V6$D�~��"�<�ԟ`S�#V��W	��5�IӣK��Ms��?��]-he�@�d�O��BP@����s� {ǥ�G �7m#�ăy�B�'>���ȟ$�I5��B�A�${���n��v����4�?� ��d=�O��$;����h����v�@"��:�H��\�x:�	Mҟ��'
��'WW����Ĉ5k��T�!�@�  Q-W����N<���?�I>����?��ѭD=�d2��I.��x�o ��}C����O@�d�OʓS&�1P:�����ud�8G�\�4�[�xb�'��'�r�'`�d"��'vz�  �B�iB1*�a����;�p� QX���I��X�IHy� ^l��Riz A����š�L� -*2��~y���'��'���'�� h��'A�`B�A�ǠˌZcH|�+
kVl���IIyb��!&�����kLL������-�*� c�J�-�O���?�ZwN��fN͕b���ϛ�V���4��~F�l������O��iII~�I�/��`X��P�.�LT�@M�>��$�<q�����')	�TaR"Y�63�M	w%�`}0�lZ!l�Jt�	������4��sy�Z>��"�׋e@dH�Cl��yڊx�*�����ա��b>e�	�e�.���KJo���S��K�f���4�?���?��,$�����'Xr�W�v��TCv���H�ř�LJ���c��Ɗ$�I��p�	��������׫�&�4�j6b����"5\���O���?�M>	S� �슂�����
�R�'�؍��O�D�O���?�-;���K[=���e 3z������?�+O*��%��O(�I�^; E��a�]e�1���2�P6���"�Oj���O��$�<��U+󩙘\���.QB̩�΋l��	����Iy�I����=97�Q.U�I ����o�
d���i}B�'���'1�	�ERP�J|b��BC
9�D�QK�p����7?�v�'��'nb�	�$�L�9v��s�F��"��;�6��O��$�<�@l&��ϵ޴��e��p��Q[��CsF��Qhѻω'%��'�6�ˉ�T?�:�1j��e㖆@?d��h��t�X�:�T%+��ivN��?���~���*W3ąZ��l�!�Ei�A�7M�O���֑;��b?)a+R"��\�uo�V��8�Ӎ�8�4��		�_�~H��� +�*x�R(��d�W�T|Q ��Kw�Ѥ<�<1��U ��Ձ.D����IŚ_BJ`�BCA��ԫ�d�|��%�" <4�!�OR��0�wK��Kj�H�@F6��U��p�,�K1f�#����7NL�H��E�Fd�r�*�0�P�E6}\�
�d��`�shP�CHD�F��
_^�1df�ti(�@wEZ�*n�wo��`�DD����ʟ���֟��I��u��'s�3�"���S�$�'�'>7��q���~�"�0�ML:dP̫�eT���E~���H+6	k�6Mgrj��Y�6
D$�8qG\A�g�
���v�:|D�#=bOܰb��IK'������	M���	���E{�]�p,���}�,�rAŊ�^)!����hT��5=J�@��޵HD1O�\�'��I�Pf�l��4�?���h|2a� o�~�0�DK��H� ���?�wً�?y���t@�?aI>�7���w�Hś$=@"�" �J8�,Z��>V>0ٳEZ~����6��|+P��$Ri�|Zp��6DH��Ȍ�Ix�)#�'���1�Q�R5�p�u��	N̍p
�'kd7��D�t Q$3��yY��Ә*1O�}QS��x}B�'���T��I=C�4Z�F�>u->�R�ꑖ412��I����%dM�b�^�x�
!t���|�*�NܓF�Ą.��Q�恷��Ӛ>�Q ��XMx�6��L�Q?eP��� '@j�J�G�*Cv�h0&�2}�d���?A���h�>�$؛.G�=��=wk����
ν2k!�D�1g�y1Nՠs����B��ax�"4ғ�� ���|`��E�77���Q�S�|�	� )Hɰ���	����	֟�2>� H�x����.1�:�� �I�c_��;B�Z�q�c9�3�D�W�Ҵ��F7[0T��0:H{t	�����H�}|ZI!��L>!t�m((�J��Q�8�a_�?A�O�d+ ������b�"#�&��RE�_5;�B�'$�=�V���=4q��F� � ����'��D��D�leqU�N m���@�5W�A�g��)u����O���One���?a�����,�fyC(l��чE��|°����pV$$�!�!lO�ɺpa�"Zj����>D��q���(~�!ScJ-k�e��� 3d΁Qj5j��ѡ�߂���C��OB�d;ړ��'v���LC�c��|�3�+[���"�'�ٸ�*��?j�A˳�WN�.᪏yB%�>�/O�t�c�p}2�'�xb`r@b�A��zpT��'��#0��'��)֍E�~�sȲLi4l~ӄEb� ��a�"|����'T���pf�L�.墷@�'W囖�c�p�k �ޘ�C5b]��p<	P�A���xڴe��ɷV�t�5�� +aR�Vp�b�@��Gx�D9�h�$�hAѓ��s�(�8V�8���ߴ���%��b�bIӰ�S;6���Γ��D�2	�\T�'MbY>����Ɵ`q�Njj����X�x֙�bO����)�R�*p�ё
/����<�Og�&Rxĳ�m�z�N�z�C	���'�!C�
2}��gL��h��s3*	~R8�臭,�̵�a�>!�'ڟ8p�4�>��!T���*T�w���F�+T���S�? D-��AK�.�J�W�� d�'��#=!u�]�!��B�A4
8�iK����R���'@��'/���G��pI��'t��'�0�]1w�a� �D��P3LT(���<i��YMx�@�$ʐ�H��Є�Ȍ��a���7�r�x��$�/*���m�$&�/&��Y��Ę��L>!�e��i���o˥ ��@�J�`�<�Ӧ��B`�V!`> =P��`~r/=�S�O�|�Y���=ʬ{��ը����6+� `�'���'��~�i�����̧Ax��(M]�bYǩ�C�ܡ(T-�n<�0� 'k����p��>u� X�i��5�~����h��!`�숗O�pU3P�2jH��Q��ßT��I2?���;BM\�z(�T�C��90JB��H�3��GiR��e��"MjBb�XX�}��́/�6-�O4�$G�->cbO��F�����ſb����O�г��OH��d>	���O��OD"�i׶> �cqHΖ}�U ��'�$�!�b�@�	��	1�gAQ$�� տ�p<9f�Tޟt%��w E6V�$�,i�.�9u�{�<�6��+2A� .قZ�����M<	��iU�a�`��~䊩A��w@�yEvB6��O����|�*ސ�?�ІׅA���
ʅ@�d�'E�'�?�@�~�9�����Dj��@����3i�N�#��0}bj�O���H/A�3���U!N����+v�>aW�BݟP�<��T��B�p<r4�>.t�����H�<��jPs����2�߫j2]��KFA�d���E�W���B�к���GǇ�,�R0m�ԟ��Iҟ(���fԮH���t�����1f�:�@�욇\|)�gLD$���<ɕ�IZx�(���	,���x7����piaL:H0p����,�h��DSR�_�aZ��$�DY�a��L>����.���" �R��Rƣz�<�KS*!3e��dQ
����a�y~""6�S�O|`,�s���%�Z@+q�M�B��.�4�H\[��'���'�b��~�������q�F�9�隌���3kM��x��m@(�JY��ɣ5^���B�G�vB�EZ�1�'lG�`��X�2�'L�a���T�����~b4A U�?����?������O~�h١(�T�ڠ!�bˊ\��)�i(D�L*��1�L�!͝�� ��!�ɹ��$�<!���=z��I��\`�h��%���K�	ǅ^��$H�C^ϟ���.P`pl�	��t�'�0Uc� C�m�J�aF�5�&02Ǎ�<vdx�1C
7<�t�{��:O~p�A2�<<��HͬQ� �"dM��O|$x��������F��p<ɡ�Uʟ`��By"�B�=���nL�~�8�e�2�'k��'z�IT�ǋB�Ԕ+c�#D"��1�'��6-[7v0p����.6P��2CG��i�$�<�����)ߛ&�'bP>���,����W�p�y	�Ɔ�[7A�G�I��@��C���Id�S��Ob�B��$]�P ��e�1і>��`Zb���O=���RG�;2u���6��/�ajJ�da���ONc��?�c�h,�����hӎ0i�(D���B �1!鸄�Ȁ��Q�l)O�qFzB���`�L��ai_�o�h)�ɽbvj��?��v��X���X��?����?��Ӽ�Ҡ]&�IA�
?C��IÇj�'k��@ah��p^6�&P����u�|2�]�:���jU�%��)4O�U,�x�
_Śqlڗ�8Y����|��,$D����ñ&�~���LD�E����:��O�)�O��ș�S�k5��2dF(�ʽh�/D�������3p02嘇��K�H,?���)�-O��"�!ЇD� 0�:*��#0�G�iI@y�GD�O����O^��ǺK��?a�OVx�@ ��`�� �S?s��"" 
�xrĘ*d�x�sA��?���;�".v4�0�'c�x���}'���'$�	2�� �?���k��A$��72���фNE o�����l�E��]:��"@0 3�h�<A���P?	�R�o�џ��I���e����j<�S��:���Iҟh`�ɓ����	�|��i��'��� ��-z݃��R���Q��G9O0l����J�dT�x�D��&�i�OH���xr�ݒ�?�����d���E��'
�4!(���/��d�O���2�)�'ʂ9T`�uƍt���R���l5�� t�p���)>��q� HD,��,f2O,�TF�R��i1"�'��Ӓ%5L��I�.Si��
V�g�A8�*?����ޟ�B�Iݟ��<����Y!z=Q/�@v�1d���E��(�4�Gx��d �4x�� W� =[t������	<Bz��4�)�S)�\����_��P�mS�*&�B䉢oi�Tz��˫`=x R��/Ж��DT�'t����ٙK�Ġ�@dL 7p��J�a�>���?�5^����C��?!���?ͻ81JMaB���x"Cʼmf|a�p�P�8-�R,ğ!bz�� .����	���7eO� .~��4
]'Qd��#L��E?.�c�$ڧM��9��R�g�	V�!� ����U��������g~B,����C�'>v��(�1$��J�
��39�C䉘�diF�w�̽jS���\�Z�f���'��$L�&� �(���lx�Z�h��Lȏ>����O&���O$����?)����$삨������"
�a;�oƵ%=�T�Bb��*��Š��Hq�7m�0A@�
ƥZ\�����'���(T���Z�!G�D����?������?�����'H*<�2��.7G\��V�F+J��b�'�>x��A�����D�G�J�"���y�O�>-O�%iDI�p}��'R��z�CC�^���gH�=3ʶP��',M/|���'I�/Y�jҰ�wī[o�xql@�J�(���ͭ%C�u���4��I�����h�O�'e&L9��&>�T��>Z��p��=	KR������O����'��S����,@�v����a�j49V�9�Ij��  �S�
�M	K-;f~��'
7���ߴR �H����0F!M��S�DU͓���1|^N�o��P��f����*��%_�W�f�5,Z	)w�(�b�SQ�'�$�'!1O�3?���I�'� � �E]�H�%bQ~�DD��(O�cW`\�L[�t"�o��.�`zǞ>�d��x��p�S|��"	��8R싥FE�"��J��c�d�	Yx�����B*'i�р�Z--�	�8O��Fz��׊.����8f� ��þUj~7��O��$�O�y6�n]�d�O��D�O�NP�&�F�X���ٹ�-� ~r�c���U�6<O�����=%,��p���N�"��C�$�<U��y��H�)���1�/�K�y�K�.3B1Oi�S�����(E�(adK�1���͝�c�Թ�ȓ+�<���*L���Jg<���'g�"=E��m� l��iÆ7��`����b��;��(K�"�'���'�]�|���|��	����PHq�
x�6�,<�vUPPN�,��I���<A���<l`� ���#Ha񫆲/-�e�� \#��0����<�� �l��h3��9j�f@ukĲA��	2�M�p�i�O\�~�A��	PdxU���-|*m�@��`�<�f�װ v�� nI�b��TH�OF]��InyB!_�$86M�O��d\�i�T%���r�~D�uϋ&e�J�D�O(؛���O���x>9���Oj�O�4j�/w�<�Qpk�<��	���'�Ӌң�>7�P���l��i���C�"Z��p<y���\&�|��W-(����/S�����5D�$��-d��$�	�<��u���3��;ܴG�8�g��L44hֱ ��q�<9BO< ����'RS>eZ�����H0H�A�X�`�	�\NƤ��N�ǟ����-wV\��cJ�S��O|� ��&5j�����%eNʰ�>9��K
y|�O񟢬��$�M�ʁ�q$��a�t���>	����I۟ �Ix��W��0WF٬6x�q�֤Զ�(��<�����<�s
<e��:��3�QQ��L������g[Ή�Ѕ��*ЧP4�m��<�����rB�.~8����������_�5Y�� "�BX;K��2|���<�͕Ux���"ݠ��t�B ����y�h&A�t��۱LmP�A�MiЈ̱qI�<3�c�Бq��Oq��'ItS� ݃]�����ճ��'�!�� :���1r���|lb�OȄDz��i�#&���de��ޭ]،X"O�)�Bl!+��T8���#$FZa*�"OJ���	V�2-$�Y%��i(0�x!"O��1�@�?@���)�E�>O� l(6"O
��"�s�"=�����e��"O�h�S���1�ER%'B�=����C"O� .���E�%z)D��=G�<p�1"OZ�*�hW5r�P0�!5Y���"Of�7�I#.VZ�۠nߨxThȨt"OfH�q�����f#R>T"��"Oĭå�P$Q���c�|��z�"O��s�_�bKl)ؖ��c����"O �*�kѫ;�����N�	�
Q��"O�D�S�H4/dސ� CЛx�V	ؕ"O`�1R��c� �.WH���"O��'�]�XW:Xp��8�||	�"O�Y� b|8�N�<��pA�"O�����iD�AT� `�x��"O�,;�DA�������_p H"OfHr��a�2l�%-�q��@�"O�SCk@�C?<��v��F!�Ua�"O��Q�Y��}ےF0�ܚW"O���6'9MA�8a����A�Ы"Oar�kԂ2q�!`��ْ�Cq"O�����N��� ��EǾ���"Oޭ�WC�$�D+�w�r�i$"O�<	�>�x �OZ�y9f"O���qB�?/%x0���A�tl3�"O�4 ��T�v`=8�	�/|�� SP���� >�<��
\a?I��$]#B���&P$1�<�(�,[�iO�8�D�'���e\�Az�%����D�����逮���(�ɘ|�g$��]�L)h6�ӵ~�t�J#�J�~���DG�t������]�_�S�c�3� d���Q.Y�|���c1}�mC�'��d�~-0�@ל �С�6��X^�dt�P�yw<��>!Pj�=O��@��4Jbx˗����9O8�0AE�f;�h�Dݴ3:R!�v���LQ��ɮp�6PA3圮���I,I�L�r�n���@k t6DÖ,ڤn�X@�a�:A4q#��?�<��)	��˥�F�s�y����0s��ސ�l�8�)��^�1b�	I Q��h؍]������2��t���	��?�a�.�S�O8�q���SӾ�#�d*!뵉SQG��Db��06��P���g޽RÈ�a�*�#%��$YH���)}BB�S؞0�J�*�������\�f8Q�#�0�ا�+� DQ�6I(�*���a�O��'�,��F�W�Q8���%<@�2	ϓ?��P:���|�@�0���M*��D1|𐘑�횃w�0Hp��˄rJ��9	Y�8z��d8����+��Bd��d*��>�R/$"�e(���a������!	qqO�}�䏜:rM�@C7\e���'	~Ȩ��(�T��ͻj�� �� L,D!�;�i�12A�-�R"�<���@�ّC�"=�;#�[�w�v�ٖ�}&4�!�* ����dK0d�"<ѥg�=p=`b�P�?��QW�A�'aJ�!�C߬�:�x��Z�`����*On�hCgˮ�p˱��%�m2Go�<y�%���O��*�e�:|���͆.L�� �"T/%0���V
v�l���� !�B� U
��P�l�b��''��Y#�D��c N��gK�x#N<Y�'O���B�Ը{���"�`~�[���y�oI�P���&��X�`�|x�X��)B*ͻ+���Ce%O�=�pɁ�H�b$ҽ�f����GzZw�z����{��
sw�H�m� 9�9��Ej�'�����¾i���2A51����C��=�}����9���3 �40�����?�s�(��&�
K d��'߃Ƽ���X $K�v�'��<��o� 0�(��.�IbxM*e�ԥ,|�arH�=���� �Ǆ�J\���Q?f�����?�<���\�1�ˁ�F���ǂ��c�h㵨T�%�6ep5�o��OrMѶ���\xı���G1f0��*���ʁ�)�J-��|�B�`sC�@NY��?`���&�.v�h��$��?Y������
�ub*��-J�8q��(��$r�j��'�ֈ��r[��&�O*��; �A�i�c��c�h
�,��l�n��),�p���O��'�TKG��r��q���0/p���'�̑��	�h�| ��
.XTI���0.�z$��6�%�1E+!I*��J����k��N�Y�ıl��Q��)B1[]Cd���?I�SG�O))�O��IZ�HElt#$����'���k��B��xI����x�D���G�f�,�c �U�Kl�'�JѬ��(�W[h�tcS+6t��BC)1
}r��F��6�D{Ҋ?!��Ҝwh��kb� ����ʠ �� �O�p�3h����I�1���"NB#�(��Ŝ ��e �	�H�����ӫA3�aY�n�$m����� ��6����I�{���
6�&hY�$���� �Őy4� l�9� ��$WJ����V���j�}*��Q⇘*�����F�p Y���	�\��E���!�\���U}2'B?� +�*L��u���349�"<���ި)�0��'M�/WLr<�r�Ni��<�t�^-�쌘��O��p�'m��̓f:^�)we��\!�R���T1�tj�녺2����	ۓ�yW O�Ѫ"�IC�e�:*�0 ��-�j�`��I.V@��P �����a�B��uN�V��+����o~<erπ_�'g�akAf����OUB���bZe�q��B��7�rH�W!o�UQ$����S��'�`�z7��a�]x%L������}f���FE52P�����flD���t�����/�I*uHA��#"��o�9%�P,�A���hr������;�O�E�����'�
���	(������M�ִ���&/�IH�Cϧ$O��dی�$%_=ReK�u-$奟>��u��9�'؂��h��+<&�p3㋣N��,:�'�xM��>�tE+��h�8�B
=�@�H�JO�"����֮�$�"s	��@������ g��_�/ӊ	r����Z`�(!D��#�'ŷ)E��g���#ͧ�Z�Y�JH�"P{��ǅJ7�i�ơ̯a�(�$���
g��%�.U�5G�?Æ#�6 H�aW/�A��AU�m�p%���rl��4���(*�3��'�kE�G`C�(���Z�<yQ$����3`.�y�h�S(�lcM���g�@$���'?O��
�o*0���^uƘeJ�*h��mZ�D��#��l���@�i��I�\j�0ɐb��ݍ)�EJ�-U�{�|Aq%��
)�ܚ��J�4^R��㉌f��I8�w�$)B2J[�C�2ubN1}jxh�J�2�4�8�'���Q���o$(@6B�~�����d@!W� `gQ����ɍ+ўT�еm����K�f�p@p�BԡaE�]r!A@+*���bÒ>f'���Kw҄���cɨK���Ln�+z��jt� ��t(Y2q�x��B�
/;w��k��
��MK"��P�(\�a�5�4Yt�@Ҧ��_D�\�c���Y�'�N��i��G�t�#�L�#
����H�@��Áo�	��g�	�o�x��1)�ȽxB��j.� ��B��W�.�`�ԛ�-����~�Od^=#�aW�k�iP�5�4��+�:t��^�h��,M*��4��N8�Px�] �y��@9=�XatB�<�@�@0��Ck��ҁJi�0�!�d�|�2�ڟ��$C|�0^ce���� %:�8�w��q����%ғ&�Hqi�=�@��ژN�ZIh���f ꤘF'S%B#�@ "�D�.;��Q�V�	��uc�����S�4�hd�Fl\5H�$���mW8y*��Z�3k��A���<��u��
0�nI>Y�ܹ��1O�`��J�s��G̕�\_Nt��V��Ö��+��Pf�G�e�X���ޟ̲G�/e�h�BH��qz��Ò��?)qC��:��$�H�,M{ L�A'��� �q��X��M��m�i|h$�4�"}Zw� M�E/��U�1�ℎg�Ԍi�ň&h��qP+��8+N�z�AݸfތiP��>��O�[�wy�e����y�""�� �&���oN	:�'��Ls+ߞd S�O�X���$m�VL�3j�����]�@\NM��5�)E8�@�@?��bÄ3���$Ʊ]��كR��;hʄ��"u�b�q`�?,�� ��O�ʧǐ�CW.̀O���O��Y(�1x� y�f
�dO:��'F���U�tZ��GMb@�)f�qH�Ә)7�X"iũ4yN� �C}�X ��ӟ�H���+0�8�sP�%rИ<#a�~2�}�Ɗ�2���+�F�;����MS�N?�Ή�fo�OB��e�5e�P�S�}��nI��u��/Bڨcn��[H��A�O-m"GN�f`h��L_$�Մ�	�Tw`�i�C�X���H�ȷTZ�Kq־� t�eLͦ�r�Zk���>��?	�dB4hN$#w�ʼ-�=��c��$�V�P�f���"�������dfɺ�Ȁ3�I�uao����V�fȸ�ؠ3����?�2�I�>���a\�q�J��'�.O�����V(`j�YQJy�L��,�_kJ��B���]���ǹC���D I��7��k�0�:s�J**?�3����ɶ��:�ʤ`FC�u���j�Kń�"Y��;gI��`YV���|�'��m2�P;�"ؑ��;`NQB���ch ��e ��]��{��^1b�z���^p*Dƃ^	�D�+V�w�h1�qW��`=�Y�����w0�X�`F�J^Y�Ԫ���Q�
�'��Y��h�;H�V��'��I����]���I
:2��Ц��=p���'(�>������ 2&.�6��t� 'OFm2���'p�zGZ�%dL����^'�I����7��Dքx��(�q�$���@���'��A���-q��;d`ЬB��`��O��s�Ѐ������u�a��?D�� Ctَj���w�޾�z [@B��2�?'�{�#�-d��ӫ�7/?��J��E���'���H��g����F� x=Zx�.����Gm$��f��5T����ƾ	`$u����$�"�GOS���b�-w�9XR'�П�2q� O���p�a��e��	�S�'b���p'��,C���m��VJ�b`�t�pL#Pd�vyb�G�H�4uj�&S.���`�ܔQ|���''vm0�jJ�H��L�O4�����֨	u.O�P%��k�A�(��I�!J��$�0U��0%?�$����t� 1U���捱G� ���V�f�S�� ��~�\7*ď�>��A���T�ũ�|��e0�y�LX���?ႝw<��H���7\��\y��Q~��	�S���W����+�J˟t�z��dG]!TS�t̓F���	�4t�)�bZ��?����{a����|jeaؘ*���G��4��Q�4��qJ�HD|RMɹap�╎*v�اF=�?
� �L����-y��e��.V1;6$�2�ܔ8/rO�kb�gK��o�����(O���&�ͣ��5l��X12?O:���J�0X�R�5cs���"����yBjS�%zn��tÒ� �U��I�o$6X��V�
�,���I�`�@�P��/t�(h �)v;�B�*Uj扢Fr#<��yG�(I�
T`�!�6/d��i���0?�t˛E@H`䪗�K���z�N֗+�`\kQ,l�'Er���W<r#��5���=�MZ����)V����	v��e
��5������iE {ڜbS�M�@�^L�	�WW��c��
�F��4dH
}{P�'P�k$��4Vz��B��Z�4�4]C��d�����g�h躵j�(��	�+F�qc�*2��A�DP0z�^!�� -��u�j`!�F�&�6��g��Jv:9Y��6B�i@Dam��غ�
=��QFc�2��g���K) @�7�1\�T sf+B�x>����J	H�Ft���c4Ldr��9[!��Z+�5�Wiۆ:?��ui�?5.:( d�Y!��O6���g�k��s�IO
ة�-��w�d�K�Iݨ~���g���0<q��L
bV��ND�|3����ݛ7T�����,m@ř���K�<�'Z��7�?zx�Z1||���D�^��|�G�\�v��#��3`h�əNe�8x�O��'@�	�у �OtH���Ƌ���|\k�=c	lxW�F�jz��A6����c�'��	K�m:&�PT�V�Jp�� �Ǐ�Z&�aU5-ո�A��N�'h4�E2�N����E�� �b��fRrQ�ON��uc��@ZL���B	�XPl��N�3_���I��$�0y	����2,1&�ڲˍ*'>��^%X��$������På�f�xbj��R�&,�K�:4��S�xxE�`�(U*`��"7��H��B"(b �B�Bv)p�ыӈ'�[]��#U�^Az5����2m�%%��*��)���G�)z��`�J��նW�M�"��MC0m ��_�^� &�˔n2Q��[* �IDB܅E�YQ�	��P�d�OQ���&#����dC�y	H����O�OaR��P�X�a�r��n	#_8$�'p\F�5}�d�ҡl��+�n8���5��~&�2�j�9�L@�@ψ�;�2���%9$�� ��46��$r�O�  >�˧��Ha��'4>ak�K��PGh�S�gجu��Z�+!��x�J?�$�KJR�A��[;B
�-��M'�!�D	�j��t%�	^ܵ��	���'�ܴ�����P�#EB�)S�0I��"Ph?=�!�d�	�<��K�E�A�󡗞x�!�d��K�A0%)	]A�<iSCP�F�!��I(R?:q�+#���DR,2x!�_�|������x�F�fƝ.Ij!�D�12�yk��RB̼�3�:Q!�$�	}�`p�J�G��h!�@Ѿ+�!�D�*)v����@��\q'i!�!�DV�C�h��P�mS+̭C X���'��aC�T>$,��Q	!9'�E��'�
M�w�I2&k��;�E�77�Ԭy�'�D\K�ǅ�V �7�Z.z����'�ԉb"H��.�̐���=|����	�'d�H`�O�
].T��"s�VA��'c� !�
�U��̀������'��P�I7|�ܑ�"ꑑqrp4��'�ZMɁ�U:W��X e� 0r+�!��'���i�;1S�#�+�jM �	�'�h��
�m����P<T���	�'��`�eEE�g�����a�;K��(�'����c((5\l	v��J)�I��'�RTsƚ.w3h�0���?;�Az�'|�U�Cb[������g�10-P�H�'D0dcB낮m8*���^�SbJ-y�'���ЬĦ+�ew˕���'r��Jp �Ee��J�>
���#�'E�x��C�?��X!��"�|}��'�hD���
(8��X �S�*�V� 
�'	d�b�4c�x0%@��\�I��'�v�q0�L8O;�`5,�#�.$"�'�6��Oנj���C���C�=A�'��T`�N� خ���ݱ:���R��� �Tj��?=r�����BKT"O���WcߒP��U:T�\3	|3�"Oဵ͂a�ܙ���
���0F"O��RwCF1e������Km���"O�7O)M�L�r�P�@X|��"O(a�'! 6���bCc�5Pd�m"@"O�b�+�C���`b������"Ox	�#�:�@۷�1�z-��"Od=`u��	��q"C�֩MN��u"O���#=}B��q��6-j
{S"O�0����8��7V�1�`��"Ot�p�H-
֔i`�f¾bq:�	�"O\�a��q�A3� �WZ�,�4"O�ي���(8� �w�MSr��7"Ob��Tk�$Ynl�`�� g`����"Oδ���A�x���T��"O��1T._�H��y�ŃuO\�F"O(��̜#TJ�R7�HD���"O6��� 
5(n �s*	�\7&�c"Ol�����)*�t�q)�}���"O4�2v�i�<�5iO�ؠ��"OHВvל�ހ:�R�R{V틷"O���)��d�h�'#yf�@:2"O�đej�D}dq��&��"��("O�𪰩��$֎�q!��K��-�F"O.HBC��3&DaC��*vԀ���"O�,�^7C�N�3!AU����"O �X�m@�~@ֽ� ���C�, w"O�P�7�=gB7@�0vo�� ��'��*D�3r�>tC�Ğ���<Zu*.D�HY�G�%#>�|)����#q\m�F�-D�l�s�� =*� Y�,���
��,D�8�%��Znpi0̓�o����=D���P�S	yXDpw�ªJ$~L���:D�آ�Ĉ�C�V�1�( �&�)���6D��1u�E1e`��f�8G������<A�1�x0[��:���bKٶu��Q�ȓ99dPa���a%t��4���X��|F"�S(�t}�G�TB��L�&X�@zC�	�tG\��@,٤lK��'
��^�hC�I8v�P�0�a�5?E�18� �E����$;�u��ԉ��T�(�+�K
&H`R���R[��ݖ�IXĴkNQ���1���s�	AB����I���gO�u�t�/D���+Ħ� ��6Տi�:	K�I2�	n؞���AX
qz� 2ѦԮ
�2pJ3�O��	Y�*iKWj]%	�|̓W/'I��B�	�ٶ!Yb�ſpFl�yfj�s��B䉈o�|�(@ό)(6@����l�����>ٓ���'튄�G�@�Yx��@�{�<�qn���0E+G#F j����k�u�<Q�A�U����"�!^�q�Lyb�'�Z5��b�ug�,!dI�� �艠	�'�0-B�ӥ{�j�I�⎦`'7"O�iH��쑢5fZ�O�}h�"OPI�Da\-�,(�G[#B[4��"O:,+E�E8n����0�����x"�'�
���7������6Ś���y��UP�N!��ݗ/><���п�y��ŷ1�"��l��(�z��R�y��Z��r,�C�Y'^z�k�����'5ў�OO��"���S�$�ba���&x��'��� ʻI�4J����$(U��'���g�6�����ƣg��r'�)��<� �-R�-���y��@
>�^@82�'���'�eŁ�<�1H��%I I��'a���Ŏ�eE���ME�Q��ӈ��&�'
/^X[���#u��$H��F!f!~Y�ȓo�>��)]��+�H�y�����,�1���tR��oR�E��U��!7P�`���9
�=j����t����Y[�qr���"�4"6-�:k+���ȓOO�l��'�>!94�Q$��4tOFt��c�Z�Ђ-G8;�4�����P���0�@���Z-�@H&�ӽ �=��W亸Zѭ�a��((&		x[�ȓ@R��J$k�s������7!����eq�XI��1f�X�j�`Z���Մ�Id�u��<�ڐR��ּY�-�ȓxB�RmFTD� ͔�)ЖЇȓR��ר�W �hR5|i�u�ȓ#� ��FX	'|�(F�U�F�v��ȓ����x�����,S�h��ȓ6ؘ="P���Z����b�*��|�ȓ��E�q���|1V@CPI�>jxM�ȓss�t(��1a�P��Ap�}�ȓ
�̬
���'4\�ʃi~.0��Iy<Q"i�!n9np����>&�X2���z�<Id
Q"cC.0�};XE��p�<q�.�)#�}kQ�� �fy�e�h�'�a��C��=� )�@@���_ �y�ǲXz� �r�ϤY�
D$�'�p=��}2n�8vR��E���g�b4�����y� $_�l��#�I�ju �� ?�y�L1{D,J��U9��"h_$�y� 6��h�@/Ǆ+��h��Z��y��=^~��Պ��$d��hĂQ��yBH)U�]� ��+IDbA��b�5�yR�Čd��D�@PL���a����*�S�Ozf4C��+@�����U9pQ��'�uC!,U=T�:	��ǴT � ��'8���DjL�U��� : ���hO�a;"�ŲRx��!W�C�Z�=��"OF	�7��׬�9ũ� Ec7��a�O���	��ܛi�l9�T��$r.�ES
�'�zɕ 6z��1a�ꛧ4��1Y�'��9�"
PY�Q��TT�͡�'�Йs倀& ׸%�q�E? �y�'xdW�E� h 7;�A��'�80%�+�>� p'��tl��'�Z��d�K�Y�6p�WLZ��,�j�'�*DruI�>	�8@�OU����:�'���c�T�r��¾'�l�*�'Ò�A�LU�b1IPAH�"B1X�'�E��o]Z��Հ ��6qe�� �'������MD����e]"��t9�'�P#�G?��4c�D �v����'���K&E��I�ǅ��d-��'6����_0��S4K�l:
�'��m;0�"Y��r̚�Z`F��	�'�d!�W�	$%����>O��x@�'�T]
ȱ`p��X`��A.�)�'�zQ"U�[N=��G�N�h�De��'�vȊ$k�=G���׈H�8�\\i�'�r1��윁S�D�8��$����'e���N�9�V�ˇA���m���d-O�4@� �H�F؃퍽'����"O��+mW�x_V�׬�;�Ab�"O� Hyy�L+n	���̛6w�.�I�V���	Ǌ;���u%��P�CJ��.!���u����反��;p.�=!��*Eg���F��%P�t�E ��lb!�W;��8a�Y��I�.\O铜�>���IA���p����3R�l˵S�<��G�b�����!z"%��lL�<1�O�i�T�@���30�@�'iLE�<A��ә0
}��bL>s7J$
�.�zh<Q ��Jx�jɠ7k~ٺ�A�$H(|C��7�<�6�ȺQ�X�YD�o�C�	�7��@�Q������c�Q)F\�B�I�<1���U-�&9�vA�v���f��B�	�R=:3/�,��0*^�hQ�B�
T��-s��[$�޸Pg� z�B�&W��@�N*ꀁJ!kZ�V0B�=M�Q��7B�lу���n��1�ƓH֞�p��RS�`�^�VO�$��E��=��kW�������|�B��ȓ9�fPHu�Ɗ��	2G�-V�lЄȓf���D�U���( ��#���ȓ2��q2c�/��1�Q(ذ[m�l��M������$� ћ�%-=ĭ�ȓ������F������,��ؠ��q�Y�Fᆇq�E�	��d�ȓ(T�#aр_�~e�Ԭ��5!e��h6\���`Q3y� ��O�
0�*����}1�(,�|Us�"w
4��[j<|ۧ�J+j
<�3 �5;B�h�ȓO�j$�Sd�x� {+��ިD�ȓbќ9j����F�J�`J8k�  �ȓK�N�+�!��ع	�퉷2�J��i�"�c���z�t��H5/9(��ȓa?t�#(�(o@B��7�U�<� �ȓ}������͠z���̑A�P���!Rv��qg��x�YA�`v22=�ȓ5HVu�BJ�&���� ��l��QSha�ĚJL�2��]~�̄ȓ�2�� ӿ3��=��ǚ�y���v@��Ɗ�*�0��� )>7�i��s���bۣ�X���$'a�~T�ȓ:Xf�P%��*r$!�lǩz)ȝ�ȓEWLP���:;�:u�L˽3A=�ȓU��T{IܶImR��E��a(]�ȓ5�\��e�JBy�"�<H�D@��-�I�t��%��S!W�SO$ ��|���c0Y�"��@`���6U�")��/�\�fÌ�f�N% ���4����L'(�B i���Z!` -@�L�
y��_Q���0eT�]�>@�PCS�I~����:E-�%F�j\��{�A�FH��'�R�kELȏ��s�l��B� XA�'��� &�Ȯw�,0�k:3bQ�'E@$���y��elΦ7�8�{�'Wf��Q���/�n�c��09"8�'��(�t���o!�٨��͛#
8U��'�p]ҲKْIV����$J���'���ˆ��q���K���H�'�v��eEd@�mK �)vcB%��'��0 ˗,�Ht1g��0o����'\H1+N��l��Kf(R�h�b�[�'.Lç�I�T�j�:�,\N���'`��˶�F�voD�[��܎P'�C�'jn��# �5�U����LO�$���� �(�Q!ϴ4��c`��a~��ر"O�c'�ǭ� Y�g�B?q���1v"OT�
@�n2�E04�Z(n��"O6�Bg�(LeMKC�Sio��I"O��@VH#Xe�BꟂ"�q�'"Ob����aH,
�$#��Ac�"O.m���Q�<I|y��Vr�ҹA�"O��8ϑ1r��H���D�r+��[�"O�� �*l��r��g8��"OF�S��xa�Q�l�/f��4"O"y[��]�	�f\���۹%֬�W"O4Q��뒼PP�́�ϐ*Bt�E*O���A�D/]���2�``��'�����/�4�JS�X*x0�'��S��1f/�\j�A�3����'`lA�!m6*�����a�*���:�'�Ұ��N�*R�Z��I:�n�B�'����d�x|VS3B"���'V�p块lv�����${(�c�'kN�+�ɓ�A�:IJ�,l�P��'���b�Cظ 
�Ш�=\���'�x��%�W�E|�p��*�S�<��#	 ����	б��)��[R�<1�# �g-��h՘[�tQ�uo�Q�<i��ԴQ5�<�qEB�p�*s��E�<�BZ�J����A+��k�
a�$�Wf�<�D̦?����PmY�F8�w��K�<a�Ds����V��%G��1ɞa�<��
;N5�b�@ޙtP@��M�`�<�m��)�Ԉiw���U2���I
R�<y��ZMێ`�#�پ9b�|rӯWt�<v͎ <R��*���ʅ2��As�<	�B�>��(�k�,jؘw�p�<i�!Hh��\i &� Lv�h��XU�<�D�^5VFe�ʖ�+�r�b�J�<!a�	�}S.�� hE�m��B��A^�<ٖ#B͂�  	#=.Ʃ:PMX�<Y�jۇf��	#��*-_�a���S�<Y�jX?�bX4"E�(�/��ftB�ɿ}:�A�MU3q�*Pӊz�@B�IcƢ{��Z�f�f����ϗ;]B���X5#�a�A�f<��4�(B�ɈDo�=�i��`MN`y��<��C��)1����AhS�O�$i׏�eِB�	�30�(r1�Ud�P�[D��K�B�	Y�6d�`�@�訨��vQXB��,�:aBQk�<��|��J�]�DB䉩{-H��J�� �� ���-TPB��/:�.@)�ػq��	�FK?�.B��lɒ);����tE[s�^�D$B�ɦu�<P��1�^��BFʼZ��C�I:�*��8-+2�F�/u��C�I�y�Y8�`
P0Y9
5k��C�'��b'�Ȗ.�+. 3(� �'�	3,ƞR�ș�	�U<�e��'o��A@d�?���ʓj�T�\���'��M��: x\2G��P��'Eȼ�4"��5t�x S>s��r�'�Ldc��֩4K,`���d��X��'*؉Ȁ�D�4���'�^���	�''�聓��4�Й�T�H1>�S�'*�U��+�T���� Y�-�`���'θi1g?ntL��+ĝMe�<��'6��p�I3�LUD�&@����� ݓpG�\�(���i�"O�u[����t����.YBXq�"O�щ`jZ<'���rQ���@VVmZ�"OL��d�$ �}r�le_V|JS"O:�#`���y����+;�� u"On�cV����13�h:mx�"O�!#c��:��Dy��ѹ~�6&"O�a#/K��V�(�#Ě�#�"O>��R�ܦ4��Y�u'C�2Ӳ��"O�p�2l�<!=h��4' ɲE�"O���V�S�4��I���F0´q��"O��ĝ#��E�A�4GK��:"O�d�E7P"��pR��#N@�ْ�"Ỏ�7	G4Qj�M�� �rE��� "O��Zv+�;,��ز�ϖQ��"O��3 +�:K�X��PdK�m��"OԹw��$�T�5���6H�=�#"O6(���:��)��I�i�h5"O5h���߸��nTG
Iq4"O�e�r@[��6��QC��y�"O�,���ԴT�:Pn߳pU��'"OQ(ҜO���צǪ=��mR'"Ox)�D��q��5h��2"kh�""O��I��5�t�sD)MS$�r"O��rn,Ai�A�c;)6�P�"O�ڣ�C�z�F��F	�8����"Onp4IBs���fa�8���"O�����s�D��p�&�ʣ"Oh���7E�]��F�&[l��9a"O�+F*(�F�۠��+(����6"OPe;bn��?�*��%cժf��h��"O Lx�F$Zʐ	"ʍ	�d! "OF ����(�����a?U��$�"Ov���ҵH���#�ТF�>p�"O���II��AhJzD�E"O�\p�82��<3�@��7n��i"O������*Cۘ��&DP�9�"O8�$`I�r�8b.�:f�$��"O�{ƢԧS��!QqE�X��i	""O��J��˹�B� SE�y��L��"Oj�k!�QKA��!��[1����0"Oj��D�)5b�HH�,	l�*��b"O�Y+@OB.^E�}A���.�2��b*O�\Y1��0wI=�Eݹtk����+rP�*g�F<J�8��㏅8l9Z��ȓ��%�ɒE���㡎	7n��ȅ�Wf�(�bW~Z6���0
�R؄�.��L�R ��]��hB"Bo��E��|�E8t�&��d�sMAإ�ȓ�h1Ï�}1F���O^?ZX���*�>���	U#{N�R�&��Nt�ȓ^o�L��({3��C#�7`������� ��ʑN��93�$�
9^�͆ȓX�Jm��U�p�*I�`�W�Nihd�ȓ�qB���%�F�H�I������!!,]�6f��<�A�!I�c�|�ȓtW4��@N�Iǚ!���6�\��ȓ�YS[�}� @��p��;�Q����/2�-�5�C.�(�ȓ��I;%"�h��m@�*E��ȓr�tdX Ʌr�J|�_�lvlh�ȓzCF�1�$��qW�!��o�ui���<l�!Z��\p�n�/�dцȓq�|1`5�ݧ� �ʲI�,��l��S�? .4:��S�F.Hi��Ȱ9(�bp"O]p5�΍F��M���+QE)�"O��S@J
YhP�Po̯TA<(�P"O�81diκds�,���ţ "OP��͎F�0x��8q�Pn$D�|ġA ��l#6�:$x�@I%�;D�0� �8$>�`�m�gt�P�&B9D�h���B�q�bѱC �?���j'�"D�����mA��	P��=���²I#D�$��$�
F��!Ɩ�n:�܋1e?D�l�5�˷&��j4U*)�*1m<D�����
/rgz��pf� Sm~0Fk:D�x:Q
*A�����<H6g%D�8��j��,�JXQ ��q��%D��JT�÷R�b�#qb>�i�c+#D����::�Ha�NٗRծ�p�6D��k���*e�x��]�܁	��4D�L �χ6Ud���B��Sr�B�4D����ˌ�|>\��i�W=f1�8D��t�Q�G�4v*D�TL"i�;D�D`���������3��c0�:D�h�s��%�v�#j8�~%��);D�;q�
U�v1AV�[���y��:D�P�'+����b��Y3`2�Ь8D���e���4B����F)��
8D��r�h�3JX`���7����Ю6D�����9-�.�ui�R����1D�4��Κ	+�5p���n�@� �3D���%ö��ht��:`A(�"��/D��!���F�z�E$�/g,(p�R�+D���E�ҸB���r���&� D��J+D��ä�(N
��u�֎o�iX�&(D���p���w�^�Ci7X�0���8D����
M�XT�jcK�b�$��6D����!�c�D)�ÀG�J�Q*D���C�(�M��蚄-�Q�F�z�<Q��>)z� r$A��I�EOu�<�c�	g��H�R͡o���*�c\X�<�����ҋ����j�{�<�B�9f2���99���E�WR�<I6�m�0�Ñ#�j���X�<�a�ih�Q�	J�6�hG��x�<����>R�:4XEeˠi�r� I�s�<A�jB<:��]��mѱ�8u�@R{�<�d�ݜ�D�*E,fPH�gZzx�\�'ynb&��3!��9�t��p�8�'R��r�ٯt��{�C	d6̔��'>j���ꕤd+F��C��WZ���'���5$��;�`��Q�f$i�'�zܳ"*�H��#�,H�K[����'[0��t�Ϻv+ش�`�%BH^�#�'�P���-�w���AP�@�MO�]C�'�@hڕ��(���4�<j��9�ȓZT�:$�Y�=�(I�U���.��)��7 FhX�W�m:��h���%$����cXf�1�#�4�����(�<1��/�ԃb$�9:Z4�"�'�`���ȓ
�D����>��p2bۋ'D�q�ȓU�Fmp$����4�%��9ʈɆ�],��� ۗLH���`��Kd��ȓ`q��˔F��$��a۰�[}�X��ȓ^*cІ�1z��3ӥc���ȓVT�x�w�Q�%��6�F9Z��ޠd@J �-�~��P�ɚ�^���S�? �|��	��d	'��Ds��
Q"O�q�G�(;�\9�2���:��$"O:Y)�L��l�,��3�+�ܭr"O*���W^];0��	8x7"OT{F�
��9�C�q��$Z"O�}!NT�!o��P��ɝa5^A�"O���G&1���`��PDb��7"O�Q�ʗ!4�:�V�,| @�"O����u���#s%�%��"O� iAj)Hn���6eە>���g"O�)A�Ofp�y#D�1��2"OT|��jÿ$��u1���>��x�"O�5уl	C�`P�僇$;#���"Ov1p �ԈcטT w�A5`o�=�Q"O*�F��!H��e��u�e��"O��`$V96�j��e�H����"O��*g������S�e�\�Z4"O�Ԁ׍{��;`�\e鶩��"O�Ӓ
��f�֐�+A��zq�"O��ag��R�sce׀n�
��"O��wY?P��բ4.س?�@"�"OJ��s���轠4�V�m��aQ#"O�a��ϴ?�:� 
�N��g"O�!4�
$m	~\��<f���"O.�z�$�,���� �ObL���"O:
A��T
YC�.�-� P`"Ol��ƌ�\n����
z�����"Ouа(�59��c�bø~��0R�"O�	k�J��:�� ��%)�N8 W"O�y ��9|r�xBX�3��t#�"O � U�ͷc``�p�ǀ!K�5��"O�pR����4�$���NZ����"Od\���2GI���4C��<��""Oe`7�ZzV	�`��*K:���"O`�C��ғ��&��(A�]k"O2ȳ�ށl~� �K�73�y��"O&����tfLaY���!QD���Q"O8QP�Ꙓ;wp��nH:D�4Q�"O��B�Q�
��A��[G��"c"O
ثv�ca����{�<��dD�*�!�Ď.o�L	�MX.$��:�a�#�!�$�F��Q��D�b�L�Ғ�Á}!��u�~|��!���T̺w@�{�!�D��C<������%Y�d�)q���!�,�`��M$q�X�*u��O�!�Q+6th:A�_�-r��\�6-!�ׁ~�$�
�iHE����D49 !��@2%�aŤ =B�0-��|���'v���J��Z���f� ��'�2TiD�WF�p)3b�h�����'o� ���C(>���뗯,p*�[�'�4�	��|%Ҝ��/�?Rڴ��'�A��c�4@q�)3 žC���S�')�0إD�i��#^8etK	�'�n$2r�W�?#L��$)x�	�'8fQ#���,Q�-���κ ����'�V���+�8jR�������'���ņCy�P�DM���h��'�zؐ�À�+5��Yv�U�H�<�a�'� u� `�n@���G�Pm@�'T�(H���m�` kV*�(�|��'� X�7#��0k��ɠ�h��
�'B�[q�؀!��yt��zhx2	�'���c�HhF 8�*�(lߚ�@���  ��`e@�}�PDy�e�q�L��"O��@�*͉%�i*�!n���k"Ov����	�&B�9��h�7;���""O4�0�CE;���æ�ق��h�!"O��J�>$��g��-�>�+�"O��)2O�;6F�(��(Ѻ,�#"O<%Y�䓶-a(THɞ�l��V"O0$��Ô\���ذG�x*%"O����Z�j��}3Ђ�	f��%Yc"Op�ժҲ�`��Ql��:�rp"O��"���<R���WR	��"O ���n�[�ŀF�	5�	�5"O�Y2�H \��գ�@ �8E�"O~���	�"�ԑJ!�D���"O���2� gԔ���� ��su"O��CȌ\"���&O
=TJ��2"OĈK��Y�*=�r�D>tGh�i7"O�]��-�2n�L�4��-�8�"O\y(��	;<A�����w�b�Ps"OD��W!ARf����J�9[>�X��"On��#'Z�T@����dWq$R��&"OX́�%�?(�Ys�)G�	RN"D�H�F�U<�йWN߆=���[�i D��)���3W'��{3�+K�9���<D��H�oLhr@��%�}k�*��;D����(W���2U�Z	CF��ڑ�;D���cK�|��	��b�?u��͐�D/D�<s�ï��LKX��Zɡe�.D�с�_8~?"�����Z�v�1�h D�@Ҕ���/��hQ�����x��=D������0k�,b2g��CX�p(�N:D�P�*.*i!Dʑ"I���9D� ��W�c�0�yt̱O<<�t�,D�\�5��?\�t2C$�;2����*D�D#g�~,��Yg��pL���6!5D��` H�P�
��i�v�(P��0D�\��I)ܹ{�E�g�P�%�"D�pc�͋��"�����A�L,h�/ D� ��I�g���e��S�&���/>D���+�0Zx�b�,O4D�<a� N;D�t8�c�*:�F�z#��G�01y�.9D��(񌁠nu�� �סMc�TA��7D�<8����+1z�y��I�tQ���*D�lx$��v	�|rb'�~�����<D�$yWTIv�8F�8*�}�P.D��ȱ킲\����`��B���B�I�����S�Iy�HT%C��B�6|Dfm�m��p�
��Y�Qw�C�&[v��A��(g���K�npC�ɾ�dI@���/T��h��'*B䉃y��q�0����y��e�P$*B�IG)X�)�$�'Zѩ�,�%8C�E�����O�kXV!Je�PHB�I�q���眷)�ൌY.�
B�ɂg�=�ՊS2���Hw�)t:C�	�A!��0a/�
>���#�?y$�B�ɯL	|D�a��
w 1Tƚ���B�I~�� ��'D���,�9X�B�	V�v1��L�	{|� ɡ1[jC�I�P�x�CgMW�%eR��c�\�|B�9&��(�#�B<*g�x��ٌn�jB�	��"��֩�&͠=ba��<�HB�ɽi�ЎU�JQ2�Т��
B�I�]��8��۾���� ��C�)� �xz2ᅏ��0M-&���"O������"n��!�LQS3�Q8"OP���/!EN �B1L�"����"OBԸŇƬ~�ڂKN	)-���f"O*s���j"d���5	4��"O���'��:
`���W�Z�X�
�"O��*.�=_bz �W�,�)�!�$��l����T'FD�iᨚ5!�DE�g�j�ⵇZ-��#�<!�D����xg�Y����6��_!�1n&R9����\�|
��o�!��(D�K��@�@D`c��2�!�Ā-3��9�v���O�&XJc��YZ!��3�zl������|	���F!򄋤j<0���.��m�feC�86!����8`I�$ӝ#�`�H��_�
6!���k��iB������w��9!�!�ݑ9����jJ�n�6� 2Iݡ1P!��1`� �`�2�`��إW!�d��?�~-ʖd�j��V��EQ!��L�d� ��O�&x�&��?}B!�N7��UӦh�h��Pc(�B"Oh�	ݿ8������r��c"O^a)NB	&k̀C���<R��-:D"Of����*F��1fi��C7��z�"ON C��x�Jsf�+A �lK�"O��1Á�7�,I���C�J���3"O�!��
�"��V�Z�u�԰8�"O"t C@�[�Ny�g
�%V�h@Xg"Oԩ��Х:GZ-
���Y2�0`"O~���`� ���A��X*�N4��"O��k��C�F_�7'���"O�iHS�Zo��=",6sT�2�"Od ´�ٸ4����+�3 \р�"O���q	�k��pRQ@^�FȖPsv"O�Z1�ȶΰ�y�� ��f��d"O��;�"]�;���X-q^2q��"O8,�Ќ��;���a�J�85A"O�i� �!�|:3��^|��1R"O�8�*�!��X��N@vP��5"O|h�<����d@���2"O�z�AmCΐS��-)��j�"ONQIABھpKV #�W�u�q�"O�,�Q���.a΍�T.�[��yX"O`-�W�C�I.�X��ԷP�X}P"O�$�Cؔc[�(�aI�Fjy�r"O�,A��߳c�����T/_� �"O&4bwj��F �v��"�PU@�"O��2Ҡ
�uK
5�RF��-��b�"O&�)V���(�$���њ#��`D"Of��⎁#4j� )��!Ύ�$"O�A���̋z���UeP�V咹"O�A�4�����X��B53��I�%"O����ɝ9@~<����2���"O> ��o�Ml�8���V�|B�)�S��i	�'2\���TO�B䉂~*�YZ���Jh95NQ��C�1*Qı#AD��Z�,Щ��͉Q�B��JO{p�=^t�}R�̬z�B�I.K��"uO�wF�����K|�pB��:A��a2W�P�T��
G�ɼ�TB�ɽQQ~���A�d� ��D	w^:B�	"1B� �K��l�A�ψq�4B��8)?	Id�ցIk]x�(��nL4B�)� �uk׀�'_�b�KA<5k�ig"O$ i3��2�����FO$j@�"O&;r��*7c�}�q�&y����"O��S!%��\Z��aD@�n����"O�e�0��/-�T��elO> �J�qf"O�-9R��=P�])Pb�5r�(Y:W"O��A�Q�x⡪#7�T @"ORH��/��G�F�8`��=��X��"OL]�����>E1$�lT� �"O�h[�kْ,��HЭmQ��1"O�\�s��+S��p�u��m0"O`��#J�y��dG��-8�Z�P"O�O�)K��(���Q@v�e84"O
��抃! ��8aƬA�l�f!� "O���v��/��9a�h�Fr��P�"OTp�J.oH��J�I�"O�p�ȇ
�LddN>����"O��2d�v�*�5-ǝ �8c"O�Ua�R.J�����鏖芀�!"O�C�,ڸm��� ��@}ٶ��"O�T[Ѐ�]��u[塘�OԚ��"O��R���f�!���7����"O�ATnN0d��,1b����%h�"O�@�Q$MI0�SC��T"�!�"O$]��Ht��R��7@l+�"Ǒ���/^��ɢ��$�R\ip�|"�)�(oG2\���Y[��%k@Q67�nB�S/���I�+k����O
%�`B�I�ɉ�N�M��UJ�(fL~C�I0(<p�U��8�z���֤�|C��9�5	v-�c���1*�'�<C䉋]�:4�#gɍ0N���`jؔ@*�B�=P��%0��	5Tx<�Pm6�B�I�U i�F�	*�MP�(]~���?�����L�2�"��I��)�ER���[�"O�%���G8@
��[����"Oڥ���O��Tq��+^�"O(0��4<`�#'F	Sl��"O�����j�qD[1)mr��"Oġ�R	B�� ��BL?N�4��"O8��r�S��IQaҰ�|dp�'q��J�
K5QA�G LG�f�)G�'D���sn�U���B�\M$0�!D��aM��RZv�b���
gRı8��>D��i`�� �FI��,Z b��ec��/D� PU�B*M
�Ќ���@w/D�H鱡M9��� # �����*O�4Ia��l�.q�2
�-_��;5"O�ab'�s���2��;zдz7"O����8el �Hp�O�Qj�9ڥ"O�M���\@ĕ����XW��"OT��Eb��C�~����
)�n�r�'C:��`�K"�ؓ��'DCRL*�'�z)�J!�t�b�f�@�D��'|
}���ʶ����[�7���0�'=j�M�!P� 5$�ߣ4�|Tb�'��\��o=Q\ �R��"`?����'(���lO7z�z(��L�Vİ�
�'�^�{���0-��'�A�#�D��'��(��,�![):�#�.( �R��
�'g�Ms�&фK���P ��i
�'Ü�sO�.B�"�NY/f�0�'RX,U:Q�u ��c��H�@�Ow�<�����H�
��e*KAdH=a�ǉo�<� h�k�LW�"/�,�"��O���"O���W�05��wa��d���"O8��i�B����.v�(+3"O~��Qc�G|H���M�,���"O�xa�ҝ6��`�V�,֠x�5"O0�
2�?*D`��#��1�$}�P"OpXöƘ�>L�ؑ�-]�A=�,��"O����s
����E6�a�"OpH�� I�T*}Ӓ�˨,��"OB��!�YH9[��\��<r��*D�Ta�kI
A!�!�ٚ��MY�k)D��QED��o�=�q�V$6@H	I�*=D�(yu��4/s�ar�T=+@TT���-D�$�A�w��4��Jm�L���?D�TC��T ��|6lLGx�(��:D��ч�B?b@��8�dگl�͈T 8D��
��ٺe)XH�H�'n D������s+ ��3���=W|eh�9D��3�9K��ɂ�E �h�r���l#D��2�	�TÊh�`d�vzFU�U�4D��0%�JY�fg_��8ez2�2D��1���
��Qⱦ�md&��j1D� d�9%���!/P(3E�{�0D����22��ݣĩ Ә��H"D�d�w��nnƩQB�P!t��BQ/"D�\
��Zm�����ۀa�&�Z��?D����3���Д瘷��шfC?D�*QH ~(�hC��j�vrG�!D�X@f)C�N�*p�ѯ�41�Fdx7�>D���q4EP��3i�HIzx�S�9D�xB�x�HУǏ�\l�+��*D� 0+E��Ѕ��	ϩ0Z2�<D� za�JQ��c�͘3C�䠒o&D�$������T��dX�TZ�((
!�$�<)��������u�x���(~�!��� R������Qf����G0T�!�D�.~o���!�jH�cQ��K�!��%(��s0��)2*� ��Bl_!�>X�]k��7(���S���!�H?.Fd�A���r��tc�3m!��$]8��Bu�ɔ B�a���4�!�$@�<ڈh���{�Q�Wi[.,�!�K	t�r8jv�@�R��h
�0tl!�$�w�X\���Z5�4�2�HG,|!��T-� �/ɝ1�����D<zs!�Ą�yw�71��xѲ`F�^q!��k��RsKZ6��ib�O��_V!�dK����p�D\���X�"A!��Ȫ��2vިW8X�5�!*!��̱b�L�p#Pq\n��vKQ	hB!���E���ƩX^�YJ�J�!�ĉ�\�P�hUH�:d�����߰�!��5?�}k�o�;X�I�j��C�!�̡+ǂy醣��}��(R�� ��!�ƃ<N�k�&"&��u���%�!�dY�y0�1.ǈH�� �ć,�!��$g��XprZP8pʆ̾L�!�$�8
�q��/	д%KB@�!��M2H�}1�-Ǡ)˅��1Sh!�$K�n���J�=^�H��3Q!�d��sM�}���s��P�KK$ k!��Uڎ`��N�: _��x��21�!�d4r1� ����(NrD�E�É_?!�ԮM%D�'N�t�p�y��Ͻ�!�� 8�Z&'R�8�*�Gߨ�
w"O&���^]{��b��]�nYA4"O����@&������ƥ95p���"O���	��%������Κ/��"O��pl��I�:��w�2n��j�"O�Y���ns�9s�ɹ�|݈�"O�a�їtxr<�Íӿ]��9
�"O��[e��>"ܪ4��*>�N �$"O���%Յo��Ը��Q0/��y��"O����`�,;�$2 ]����"O�9+�"nr>iSD�/[`Ƹ�"OYڔK�� ��xqt�Ԟ>'�Ms"Odh����-:����Q쌢4�4��$"Ofe��듫|��U�r�(��"O�T��U6e�����X�W�I��"Ol8k������J�3�>�:�"O���d��e�p�l?����5"O28 R!f����zQ /�u�<���	W���w��,��]�үF�<�u�D�H��R"��j�A�<�T�x�����Ѝd�|�2��}�<��"��Uda.Wt��+�O�<Y�e�9w����GѼCsl��o�I�<�GED�D������ <���,�D�<����)$��p��`�T�q�i�<�d^�8U�t�%
8r;"���WOy"�'��U[â�;m�$��V�C�,Q�	�'��Cv`�^���"ր13��Y	�'&`�Ja���1��Ų��Xc�%�	�'�Eq��)��U�T�3W,@l#�'�IZfo�5O�.���ץe:~�+�'�����¯{� �lY,n�'^0x��� ��J��5a����'ﲬ[�K:'.��tʀ�+Q8q�
�'�P�W,�^#��Y�E� )�q��'m���B.��rx�)
*�+7(A��;�:a8��$?RT4�D��%"�t�ȓ3:��p*O�1eb�YG�թb�.�ȓv�~��g(R,�r��aN�E�Ȇȓ*DHprJ�2Nb"g�,C���ȓ��@�3�['e�:��N%(X��ȓ 㺌�"CCIX*PQ���3�%�ȓz^0D��L��;5$V�t�`���b��	�d��d��q�A��&Nr��?��m��cٯB��;�"��o'�ȓq�kQJ�:=1�Y`R��$y¥��D��LI��1_��ՂPŚ�>)f��?���3?� 
���$r�۫#(~10&N�N�<I���?7)����+i��a6T�(��/Ȫ��C�B��b{̵���$D������$�Π�FΦl���n#D����'�D��0:7#�c{F{7�4D�p��b��� �� �7x�j��U�3D�����z�e�7,J�z�R���O6��)�	g�'�� �� 1�j4��ab�|`�'Ӹ����F��YAH�Y<� �'=�!i'�C6R@Ep�bAe��؉�'0M���H�Z;6��(��pŨy�
�'� h�E��*���q��l/r�
�'VX��`��M�&-���٠Y�Z��
�'n|m8Q&A6Mք
0��K��%��'�j٨5�&u(����
\h�'�JT@d,]Q�A�N�a=>�	�'c*y�t!K1xrR���h�W�>P*��� *1��B.&C��ه�Ґ_��:�"O���0�ך:P���/��=���#"O�%�����C=�A��A���Q�"O΅���#^�J];uϟ�w�~X(�"O�e@GíX�`�s��)M�q�s"O�A⁓6NǼ}bANH�14JM��"O��ST���U� ^����"O4�X��R.?F��2FF	�o�H*�"O�Y��.
CJ�����η5��"O^���n�"2��䑺6�bI�C"O�YS#�	�A��Ԃ�n�	s"Ol5����ik��n�G܌��"O��Z"OZB8}됣�'<��!zr"O�5%��<z��B�'�F� ��"O�刐��;�l	G�2'Y��"O숊t��7�����F�4XZ��"O&�+r�Zג"�˨3��ѣ��*�y�N�"���6��*=�v*%����)�O���� }B���gѡ��A�"Oh�xq$��Y%z5J�%��>z�I�"O��!���	�E[�D�q<d�"�"OL�Ј	��c�'6.�1 "O.��#�âG� B� �v>T��"O���VA�N*|��"T�o� H��"O���(���Ή�������$"O��2!͏O��􇒖t{���"O�QB@E�yk���CЄ0k�L��"OH����-��u`K�juk�"O�x	`�_#��}�6�� �X�E"O%[��	�D3�B�G�<���ȗ"O�Y#q�� dEb�fL0�x�Yp"OrTs���$�L�`TCW�k�88Rg"O�Q	��ƥ�mi���5:�h�s"O���Ǌ=�l���	!?��<@�"O�Y��Ŝ;������V���"OB`�Qc@�D~q:#��`��R"O������<�p#4$�E����W"O`2�JE�����>O;�p��"OD�%��(gS�Y3�@=xTA@�"O�wGq��%���2[_F,["O@����ǊS�`�a+�6K�cc"O(���؟(}�$S'!��ML4��t"ORH�vDY�/.D���NGK8��D"O�TC2��L���p��MJh��5"OM�L�9/���m�<��R"O�����#p1���I�
g��1�"O��C"��+#�I�+
���� "O����J�]"ir�iZ"|U�"O:�8��YY�̓�J��K��qF"Ot�ve�3S
q/�� "O����;F̋#�+$B���"O.��7�A6+�Ɛ�4!��	��"O�����+B���@���d�ҥ"O�aQOP�r��)�7��
��"O�Hc�Ȏ�sY��3�� � v����"OL�҈;j�VHs�jO�CIB�"O����N;8�Y*V*K!@�4�%"O�P���ќ?;Ȉäi�~��1P"O��C�6V�3�.� �3�"O�{�PC1���1���p��\{"O`��'���]���8�"O���˜@�B���2=Ǫ���"On�(�d��4�:�����X=s�"O.� !��'=~v�ѱ�f���"O�  u"��ۯ"��83�Ąs�f1��"O���cM�~1��H�A˃Ad�-p6"O�����*������M�zNP�0f"Ot�Ua��M��`z��JH\c�"O��h�G��ݔȓ��ՌR4��h"O�L
p-��k�%���Z;>d�%"O�� �j'I��9��)=��ɫ�"O��IP���D*��+պ%N���"O��eb�Ri2(x����Y�dP��"Of��!�J`���Y8��)H"O
$Д(�
M��SM�jS�#"Ox2AV3gmN;�.���� c�"OP�	�Дrj��aw��/i�p�J�"O"5�"�5.b�`X�lċv�6�JA"Od=I��M(n���P��,y�H�:d"O�,��o�"z�"QA
U-�����y�Âa\�U:�/V)BDXI!�gE��ybA�L먱���4:L;��C��y"h�����j,}��)S���y�⋳8	����,m�pUZ�K$�y�/�-A�[�L��l>���(���ybϜ�0p$h@I"j��#�A+�y�m�UL��R�j�d��$�y���yO*]���R�_�l5I򂌎�ybI�XJ�9�E �3�z ��f��y���`u�ă6`��z�� ����yb�ʿ�. *0$��F4Ԭk����y�F��.��x��l]?V���r���y�L���	a���:7D� ՎB��y���(b��2uo�,�	�tm��y�� K1�DJĆ]�#s��o!�yH�9p2d	'�L�x;�G��yR��?&�N���S3����Ri���yb�P�kF�����Ѧ-�0٥�C?�y�C��#D�`�/= ��(0b'�y��<C�5��fZlJ.�Q�ל�y��p5�	���N�\?��b�Kߒ�y2���0�"dzqO&	��cV���yrF�x;b�E L4D\�p���y�)� ��i��̗ Vh	�$��$�y"ì�v؋�σ�
�q�1n�+�y2�E�bY豥�}_ �Q�˜��y��ѹ/��J�EI�o�m0qH��yb!�_��d��`ئ|:���p���yrc�2J���&�q%Q!�A3�y�D�2;/�g��f���n�/�y�B��|��P�++fN4"֧���yb�t�(yp+���ӥa��y�æ2���Z0.�J�`�L�$�y2�!�����LQ	dHb�#��y"c�7j� ɱI��~�
1K��:�y�l�x����i\n��(���X#�y�ʀ�@����Ł�.|C�F?�y���$�`��E��%�&�H)���yr�Z/Q��dl�3\֘����y/]�eW�ŘȂ��8�.W#�y�	��x�Ҥ�߸]K���Ȏ�yB�ۍ_Uj%�B�9M.�9#D�:�y  �y�Fy�t�HQ�UASd��y�H�5�<y����y�uX����yR.S�T�6`�t��t�:�R�(�y��uLt��J
Uw�d��?�y�)�
g0Z�2��'���a��ó�y�kWG. Xs�D�-���z����y
� ��I@O��q��Hv�;Ԏ���"O�|@�Ǝ;����d��H���k2"O����޴b7*p�3�Z�M:�"O��*pN8dQ���'F,��((�"Orh���M�}4A�'�0�H�"0"O�qH�B�*$\#�&�mڰ�Ӵ"O��b�/7��p����j�B�S`"O0i�!M�X�n ���-7����"O�%Xd�>M�ܥ� j˓:�D�C"O�yj����1�5��LH"Oj]�1�S�)~�3G����"O�8H�,Ȋ�:\��,]�9i��V"OH�K�d^��\9��מgWB;�"O��r�΁�k��Xwa�U���k"O���jí$��: ����"D��"O��t��)�>T�4�ՇOi�1k�"O�܀v
�*|U���cǆ^��@�"O �ᷯF:w�f �DF�o���b"O� ԍ !|��r��C�(5��"O�H���R7%�U0��K*O����"O1Ȅ+��0`0��hWo2���B"O<�����^�j���!(hh:d"O@�D��[��Ɖ�}"<��"Oĸ󁄛;��9$���#�m�"O�m!�9p#���D�J�@��"O���lʙR��]�M��HD�<����%�ʡ)@��
�N��E�<�E�9p4$�'�-/o��P��y�<�ѣ��9 蒬'��@cn~�<��Q,e�tdj��B,i����'�`�<aqϊ&B� ��\�
n�,[W��B�<A0hE�f6@�ӕ� ���yB��~�<��� ] �4�J$
D�"5K�x�<9�#�kD�z#��$6``Hrơ�u�<��?_ˊl���B�IR�Eb1��f�<�U�
(S��Zs��%Gl�K��Oy�<�4.���x���3�S-�~�<�)�7@Ӧ(��P���iaj |�<�!I\�a`��K�(�%� ��E�m�<�e+�47��H�PDd=ɵ"�r�<i�!F�`T.����k�v�+@��f�<��M�
0O>���E�EY�;���`�<����t�b5 Ek�3���b޸�y�슑%���ZcȨ{���@�KD�yR��t�� x��r�tiDϜ��y�Ę�!@���*p_���PaN�yR��.%TLc�Aň3!\��P��y��� O|�����/�T�7F��y"B�a����:WV��(E��y���0EhV��!��:3�б({B�����ْ��%<,��Ԣ��LlF؅ȓm�dpy�h��D�&��VO	�;-�؅ȓs�PD��@^!=Z$���Np{�a�ȓ{d���.��r i��M�a���9-.ћC�ѭ+$ЬxA��6m�9��Sq�U`�&ƉxH�����X)I���ȓ3�>���
�N ��31,�(u�2��O$�Y��ψc����'.�(؅�c�X�sΘl��hܡS�@�ȓ7�؀�g�<k=@-0¦òT{���b��iӒ)P�j^Dä�M5���ȓn>F��e��F�����G���t�ȓ]�򘚗G>�6!�WJ���d��=��0�Os�d�2�ؼw6��S�? )��
��X
�8i8�c%"O8�$N7v�	��BL��"OD����љ#e��s�'�dhBiX"O�<�%J�Q\́Ғ��}��)�0"O@k"��`���&��4��T�%"O\�At
^)��X �W���z�"OP�A����~���"0,\=]	|� �"O���lh�hDk˨h��8��"O��R�_4I�Ps j��Q:�("O�U�5�ˀ�H�H����"O i��fK�>@x�W&)�t�W"O�`�E��R�p�jk��v� �"O<���7BL����ҁ�"Of|�"�C2VȄ�T�8
q�c�"OB��w��(J��Hp��/�l��"OX�9��`U�&Ʊfs1"O� �A�����#"��0�1t"O:]�# �����e�S#���"OD��ǈP�[�z��O��d�=�s"O5hh������n�/C�xP"OH��A-A}*0�P�LP�$�(y�"O�Y W��B�)�!%" S�"OH�µ�R�~����Lw
��c"Ot@TS�
�� ��p�ȕ��"O�,٠
�>����q�ɗaq��c�"O¥*"Ǝ;�	AU�S�jh"O:-�l��h QA��c��9�C"ObT��
I�2$Z�� �T�m�8s�"O�hөU�M�v�qၘ�PӾ�@"OL!`��!u�3�\ l�����'�����Q�{-f�� c��`���z�'�A��U�]��WLV�Vgf�3	�'Ѹ-�sJ(�tt��ǆ�L�N1i�'=t���a>������E�����'�,��#������;`��9	�[�'h��Q!JşpJd�7G�6�la��'����j_%�}��i	0y`���'�.K�N�f�b@ҕ!���&�J�'�"ѡ� �y�L!(Ua�j�"�k�'���R`��bWB��,��/&,
�'��ԣРݠ+`��v�U!����'F�@�Qe�MPD��E�ړ�����oq��dA�m�tM0�͛!@|���
�D�q�T80�y���5�j1�ȓ��K�a�0�X�C��iJ�(U�t�<��Q1-���Ӳ�9;7~�u�<�î��<�X]CU1	��	���Ot�<i�&T�f�8����-+���J�<��NC��¡�JȤ<9�!q�<	r�F&?��x�)�2O,���y�<�0#�:E���%#0�@<�d�vy2�)�'5:H05'S��x��fi9r��Y�ʓR��M �o�[�D"S�:�\C�I,U�x@���=;v�{�$�v�z��hO�>9��ϑ\X�(�)����7D�t��'��
~���儝�@C�,2�2D��a�B	�R7BV s��"sͭ$���p�`A+d�ˀT���ᷥ_ 5��%"OF� �X+��K.��<��E���'Ց�,
�.�!	X�I�o<@.�;��"D��J2�A�.b�4����z�^h�$D� s���2/��cʤae��k�"D���&�"U��Ac暛�X��Uk>D�@�ׇ�8�2ujQ�[�G3y�;D�� ���
�2���J���,�l!H��d:�S��V�6u#��5�2${&�M!���@J�����?� ���M��].�O
���v������}n�U�B�CI�}R��:���Q�fM�ʍ!s��x�� &D�� ֪Z R�Q��9jR�DJ�&ړ�0|�	X��XɆĞ�6{B��s�GX���O|��B�<���#`�!3�j���鉂�hO�i�?�������D �r�Z��!��O��h H2M�f�s�1�,��i��Y'�vqiq�G��C�֊���!�S�O͊T[������qŌ�*�L��'��a��΃�.`zt��X�X=�y�'��O1�Z���c 28�������#O���ŕxb�'+B�z#�P�5��b��2ͤP	�'ўb?��c����pnǘp�l�ѳR�K�,��I���=ٖ�Z�*3��`�CژWpN�H�#I�<�Q��'�()��
I*`�>�	"%�y?�'6�OQ>��$ [�ʵ��T�x5"��.���y�D̴"���Qc��s�>�������Ą���>1cO�$@2��K��4'��<a��1x8�I�Ɂ
���Xa�L,�옇�IT�	.=�Z숕���<n�ţaŒ�h��C�2���riކTB��M������>�!�K���
Vȉ� �z�;P��u����I䟰7Ǎ��jx�r�_E@�����8D�p��g�:Z�{Em^&]�+�P�a~RW����ՙ3� ��j]�5Fp �RF7D�@��c��1��L�T<K@p<���'D�D����	vbn]⯁�k� �C��)D�����!۰���o
�0y�ƨ*D�$�&mЃ��KCn�4\(\v�+D�PSs�G�  �"b.ƷJ�+�b�>)��Z����tHs��<��ϕ�)P���)τmq�d�8���"5L�G��A��bﺁ�e�݄w�Jc N�Ti�1̓�hO?�3
��?
�@�[�$Ѡ�:D�d�a	�d	��K�'~� E@4D���p�W�Z��)15�_�=�<��1�/�OZ�	�>��z�N�����Ip�Кl�"B��?h3��9����P�8CWKP�w��C�	�Zx(�0qI�2��6�O<�C��.�~�JӀO[Щ��ͶT�t��hO>):�	+r��,Bt�[<fn��G2LO��9!��:!��UH�)9P��I0�v���{K�	2P�yQ�/%ULq�ժ-D��@����pK�,i�D� ��,D���%��6h�@a02k	:A(	:G6D���C.+�(��aD��.*iؒ�5D�( ��ǞW�j\�4�CH�:�d4}��'�ܐ:!��u��!�"/�z��㓱ybT�t�Gn֧j�4����t�4��!�<����'�Dxr��1-�Ȉ�%���l2T�35�=D��@����`!�1� �G�+�Ju�>��(�O�!��D�>��;`�����25�'�F�����5�%@)J>x�G�B�p�!�D\\L0�cmC�B>�d�_���'Na|�'��]���{�-��-~�Ԅ�.�y"!D�-����D�@��d����{Ӓ#<E�͙� �ճ� �7�� �G��y&� |!��qUbʌ2��T���~��)�')�^�q'�[=J��I�J4>�ȓ(�܌�B��9��,�,�!#<p�ȓ\� �9E`�A5��zQ�y 5����s�� �4���1)B��iD�1H��H5"O�����-��$P�"[0v��W����I�sb�y ��Px�a��_�C�ɻY�Tb%A�+ lV�a���LB��l��UBJ>Mi�}cac�S,B�	9]�� �j�&;��q� �{9�C�Ɋ?'���8������0wU�C��&G�f���o,��P1�&]%}�C��9ah�h*e#C�UG\0"�ܻSVDB�	�����eJ�/�>$8g�[�~[FB�ɑE�T��B�۠\+�D�b6,"=ǓN���1��6��`��m��1���ȓ쒅yUb�.~p�jBT�e�ȓp����G�54�`����H���|��6��yC (~�R�Nӓ�d��O���#��.��4�e��	ʘԅȓS�~M�CE��Q%4�c7�'nⅅ�=x����ʀ~'�M÷�)#x�,��}�9ka��Fo��R$��(b7�ĄȓD�N	�H֦D�vJ#5L,�ȓ���q"�+Y��,ڤ�_˖��u��y���9&��ɗ���4L��}?�-��	�R/�hy�(طA��ԇȓ\���#��{���oQ2'A�Շ�D�I�la�f�d�0%8d����0�p�g��[%��&�3?Ў��ȓ��h��
��9s
�����_z0��2E0�P���7-�ȍ�#LM6����>1�jI��ȱ� f��m��]I��)�'�|��c�6�ȸҡWOh�(�ܴ�(O~�=ͧ3
�"��)�|�΃9@Ȯh��	x�ßd:c��01\��FLݱ�<)��{��F{��	�4�b-^�-�4��>�!��(�P�z�g�`��ȉm�S�!��?<"�I:`ŉ�:�h\k��7j�ў����S�y�D�9�Ry�.��/��C�ɇy�����%M3�Y� T.-��7MC�	1�~���ig�Epa��1h@j	:$M�FX��r�'Z�gͲu`( �C��9�	@��D9O��sEI؟�l*��rY4�
5"O���3,��ŢԂ�FU� E���';O���>K*D�!�ޡxT:���ď48�!��-�R����p���)�!��U�&lǄ_�R@��b�@�r!��şi�4̰2�"I����]d!��_�f6��Ǉ�<-����n#C^!�L�6�U	��Qx�a�.��@a}�6?YR�K��ı���)��,ے��t�<�5��eU��s/�L���%�r�<� ��Bj �gi?5��dsRq�<ae㔕T�\�PfA,J$�b0�ND�'�x"'��^����-|M�p���y2B߹U�" +ƈ�?J�9釩)�?a�'��<B$�M�y[R�2u�ڔ(5�:�'�>L���[�V[|eK3`K�`\��'R�]Z��5.���s�ƏDu�D�
�'��$����~�ʜ���<�Z��'�A�e�����zg�:�^u�
�'�4���"�zs��Ѥ�ڃ?�r���9���j�S����!��-�� �ȓJ�^��J�|ݑ�#E	+���D
�)pT�Ҥ[u���=Q^4��d$ biX@.<5A6JI-��ȓ֘��Ӯ� ML��G�S��Ʊ��S�? :9�R�&y���X�O�5�Ɓ��"OٓX*,t��0I�:`�@�"O:H�璟�<ћ�ꁰ&����"OX�J��ߋd� ��I��m�Sw"O����nӺZ��b��N�rdx�"O��ǩ�ܔ�%�A8��)�"O�-`��ג%�'%��8�A�3"ONQo��2f�Z<ba
�W ڨ��"O���#�
a��-z��4;{`1U"O��ffک�Vtke�[�lf¨G"O����I�?
d�;�ϔF�J\�"Oh����+P=.s�	9T�Za"Od�`��$o�N�;wE
&M|���"ON�j��W[�@�1E6l�6��p"O`��šΐ?�i�jU>�*`�p"O6��4GQR����J6h��a��"OFIqB�(X��X��J��*H�"O�=��%f��X���D �2�"O6m�2��=,uz�.�& ���"OA���C�й��
�=H���"OD|Q"d�'%�Xss�W��͚E"O�h�I�.=�Vx+��C�V;x]�G"O���W�۵~3 �p��({#N�q"O&y����e�<�*�y)⼉"O�Zw�	��� 	�/h]��"Ope��J�/o��2�i^�&С�"O�h	W��='�~])�h�M��L[V"OH���F�_����d���9�"O��`�n�|:�u��$�]�"O�\j��W�M{b{l�%"O����aB:k�*�8�nV�}Yth3"Oҍ��'�4ʶ%B��\	|j�""OK�Zl���Gh)e�Z	Z��	��yrM�x�\���f����'�yb�D=no������:XK����Ԍ�y�_�h�T�(����+D"���A���y�m�;w��8���
/�dy�q'R"�yn]?/Y��QA��.T�4�z�����y"��.[�^!!uD��BC��0�	�yB^�+,�H) i�MܒI;A"F�y2N!'�hL3��%v���I��@�y�,�(>�My��/uz��m ��y�H 5�(��Tū}N����yR"�<e�P�"�9gŦlse��:�y� K�E��I� o�����׶�y���K-l��F�J&fո8�����y"�E:ypX�F�� [ �+G���yb�O�F��x0�L���D��y��Λfg�[�`ը8:���p���y�B:;Y �&�L�i��a����y�g��XḄ[��n= p�N��y��+8Fx�*1@ҲW��!���3�y��M�dے�y�!O1����kǛ�y�m�{eeA7�C2�¨$�$�ybMǧp� �D���s@t%��D��y� �H��"���U(�R!�yr��N��ЮҺ�Z�G���yB"���1e+���쩁�����yb�R��|�K��ɚ�ǃ��y"��J�Fd��;pw p�!��y��0N��l!Bk�l��1s�-��y��в#k��� �,a4�ٛE��y���!�j���,M�f��:再��y���5i8�1@�Q�c��ͲԮ��y
� "	Z��Qb�^�CfkK���=�"O0�S��%�A:�9fݒe�"O�|�b�	�r,�glǹx�XM�`"O�4٢�\�.H顴�[./ɚ!c!"O��ƕ3Z�d�D��D�"O腂,�6]�����*�^,D�4"O����_��ɲ/�h-8�"O�A���\��墁M��,al ��"O��۲ꒀ�����NW���"O�t2�

_rx��p�٪WA�E{0"O�`r��_�
	՘���|L���"O��w��;SY�̳cA�n3L�
p"O&}*�o��@�&|��B �=��j�"O�9�da�=Q	�R�A^�6p\r"Oژc,XD(as1B�rvL�'��1�6�U�|2����̾L똈�Ι&� ���3D���g�R"s`���Ή�1y�]�G�p�.Tj�N-�k�(|O^Q�����"�ʍ�"쀲Q�H��	�s&��̆&�ZUlZ�'mf� ��gXF�!��s=��'����FW�r�y �H�-����{"$Z�c��]�e�͞6��>�8G�;�x��Wfd�p� ,D��y���]��;T�A"b#�u���H�a�$m�U�й��+�(���zKFH�NM�4��=pP@�-�vB�	7H(���j�2PC��`ꙶ�Dp��"�
Z�~c�����=Y�+�?Rm��ր׿+��Q�0�Ca��<ȅ��z�2�� �E��õ	�+�,}[�Lܹcg6�4���3��DE��x��d:h6�J�h)�$bQ�A/��'I��Q��8�,8���iO?��Ū2C:LOĩ��B�����D,*2Ԭˌy��,+0ШGz2�>��q��E�jx���a/�'#E��x��eYX�H��֝�<��Q�%E�h{���q�Ok̕^"���\>�����0����K%=��L���'��L��P$ @j1�D����4)��#aJD�H*N���c��p����2��8�BP���[8 ��9��E�T qøe 6A��!�t��'0!0��ox�����\��.e9��8�%P{8XnE��P�H֣΍!eju�A���9Oj8�hҩ�y�h�8vx���V�. ���yA̐�0?)#H�F�ʑ�eHK�P��z���[t�h(0��X���bu.N $L�O��?����.GRR�Gg0#�r�PꎑJ�� �S��h�&�D|R�Y/D�y�)\� vpb���&C��.p���Q�
.H�
�<*j>��Rg�+��I�"�O:й�LJk�&yA@�K�R}���'ɠ�ƈ�� ���TԅO�"������?qi0�M�Fa��9�2��F�!�\3�ǎgƀ�"O.,+����0x���n`hE�����G���p0�������֕,k>4��O�6h��kkpu�6���(��6nYH!�1u���l�Tx����{(S�J��-B ��B-8p��F� ��S "��:Ȫ#�'n�%9@�0'V)Dx��1[/���Ц�f��L�ԥ:�hO���!,։`j0��*(0&]�Ί��u7jӸ'��is�MVA��S'���MׄV�o�a*����ڦHX�zP��A���bC(��	-l����aԞZ�)q���;���ʶ؟����1��T��;p�<�U��1	0��H�R�!�l��%"��r-�C�JR+^���FΏZ'H�2��N8�6���/���K�Y\$����q����L����M��ɤ��U�E%��NA�L� DܻP���X7��\RN!��dM�Hʥ#EJH����I�vO�Ղć�6w e�Dk0�^�
 ��H�_�촘�&N�.�l��h�����G*[P��wEM�h�V���e�*\O���+��&��� ї�؜�g7O` rbo؏2 ]9�jM(zr����D��(zs�����7T���#�%K���PHMkS!�
/�TS `âQ6MX�'\�FN��0�b��(�ᓅf~�YY�$��(�L{ @#}�i�){�E��*r�8 �
��%�}[�~"�d��<��I!�Z=����b���_��ja��{B�8N�4�+&�:b>7� �x	Da�6��!B.L p�d����C j��c9RQb �'��S(4nm�Wb��\�j��HI�&���
�*��FO���D.!�%03O�5���q��3?Y�!��=-Z8c?�K� I�dY4G�"�j��V
�*����JWq��D�/1�� ��Џ� =�3��8I�~�.o`�8~��d�-7��(�@�0}bipމ@��E:�Uas
[.T�e@/4��U��'V^�1��.�?>�<����ڡQ@pj�݀,�>��K� ���		���|nڞv�j)S�K��5��Ȇ0^�Z����6�4���1��� V���gS�6 ��&L�zt�ÓQ���P� �7f���#�'-e�Kt���Be..� ͲL>���,(�8劄"0�S�C�lMBqh�a�2,���8UT8��f���-�(�ȓ�:�0�T�r�&�0&���� �B���aI~u#c��v��=�;-tEjr�}�Z�EOc�j��ƓIq(�b��5�ԁ��H�|ӂ(JEg�/@�h�h=�O�p�5Ȇ7uPX��hŚ^D(\G�'X@�(D�ZB T�'�B4 �.˃9�d�2#G'.z��'�dUД�I��1Z �B�F�:O>Q4��A�H�օ͈������L=(�X�b�
=�2��"O5��Gϯn>�kԣLd](�,�Y��O*�W�3?��FЛ:�������`����Uz�<�6�ZCv�(��ŔSy���Ү�0o"���$�L��@S�G�=BJ�]�%잭+
D���9D�H�D�[�4�|x+��>ͰѤ5D�غTB�g�2��R���?'H�+�,D�8�Q UM*�	�':(DV�8"�*D���s�z1lIKDC�.��)�b)D���j��C���y5�S��4+$D�(�F�#b9 �K�9�.��@/D��BGኌ �0�V����m���8D�l����9rH�,��CY�J�*MP�=D����捙js�����	p.>�Q��<P�NS%�㞢|�&6\̻`�$9�����AG}�<9T@h�Go�lBy�g�yS�O��Bo^5����W�:<�9EL������-��7��~���\>��P(�X��ͫC*�)��Au��	��t��R�E�O/LO�i�2ɘ�] ")[�E M�����	&)��Q�� �W]�Y[��}��ȪVเ�`ٟ[Mt@p�@ȉ��B�4Erx`F/�$+LP�A�J�9?����x.2iB��HWL�!>2,�ǲ��Oz�ac�Ls9;�BCv����'&�IC��L7`��$Pqhі2��q0���TSF���
QI��Z��S-&�PБ �:B�����E�� �!�q 6�Ob���F�*.^���ϿP7���Dɖv �M�E�
�?%��I��DQW�>,O��`֯���I�Ə3zξ	���d����Q�nb�L[�^���0�o�]�Mہ��
���)��!��_�ΙJ��J�*���wg�����uV�M��?9�:�D�.@�T�0�E���O_XY��׳=���(R)�)`���'���$cضe(�Bl%q��X���M6�MF���,�hD:m�5��'!_��$�X�`�^�Th�(�OE��q�&�OjP�@�T�n��Y-��x�x tEG�z��] �'(ы�㘡(?Ї��hݼ�p���8'-zx)�N#'������OS�T��� �b �͑�	U�+��tt(F B�I.h��	��*�xZH��؍<��>��jl� "|Z���d;p5(��o.��*�h�y�<�K(v�&�@�fŁ[bR�hKz�<I�ßM�@�!�D�U&��I��v�<1��_�`F�V/:.�4)ԭ�yr��(�e(���;6D���L���y� NN0T�t���#���j��y"�6AU���ǖ���[#���y2�C�"�2�!#~H��C��M��y�m_�ar�xfA
)]��e�*�yR�٣cV�pk�j��V<���`��6�y�M\�[:� �AE���r���y��B!�#�F�*�,�G��y�%O�w�� S`Q�`X�k7%���y���+|��1x܉ք�	�y���|Ռ��v��q���󣑖�y���y�#� Y�z���lT��y�Έ���q���2���ˍ�y��|�h���ٓY�|pJ	�y+�i����a�9����y�! U$�Wn]�p���"��y
� �T�!�WV�I�
۾��6"O�D�W&ԛRg2�J���~���C"O0�jT�;��IU�L�	�U"Oތb�A�b.�$Q3�QUn�e	�"O�!�Ҥ�-꜔R"�O9*�L��3"O�s�$��))t� �#W4'���"O���ՙf$�q���/g�t�2�"O��ӕ�7f�����Aݞ#� y�"O0hK��X>Z��@�$^8��"O� H��ގ���yth�#��s"O@ՂD%��g�&���I�j����"O4i��L.>=�Ȫ�m^����"O m�d�P�V���[ k�@�@�Ȗ"O4$�D�j֪�2E*[�3T��V"OJ������i�|�(�>Z�JD��"O �IŃY-Q_v�R�Y

���Aa"O��c�ާ,;8M��cъ���)�"Or�sU"��b/�|�#�3����"O�i�Am�V�Apԁ�M�ɸ�"O��z��:,F�Aa�6���2"Ou��b�K: |(����$�"OV=���.���%��{פ("O�̸B�D�n��AJR�q�c"Oj��hA���M��X��v=�V"O����%M(�P���	��E�7"OF]CQ��)N�8�0�Ʌ6�q t"O
E�.Ğr�05��#���@�"O"h���%>)S L�u�yw"Ol<�����@)a1��?-� ْ"O����f�'\�feΎ
�m��"O:[&Ì�u<ܝ��� 6���@4"O ��R�T��}A�hXn9 �"O"؉֏F~��՛`���-[�A��"O�I��W;D~�u�0G���V"O����G
wi���(e�*�y$"O� ����9(�
�{ �4n}� @�"O2�-�-	��0 ̹Fv��	!"O���ևӞGK��u�	���`�>D���b��7"0�(��x���H�+D�l06��Oܮ�q��?��H���'D����@�?B�0��0 ��~�@"�C"D���@�*
�+d>�Zg�
�y���`g��g�q�105o܅�yR�љ;��yHeO����������y2KlX�ƒ.z�](1�� �y�.N�_&��K����~�0��&] �yʍ<9yr�/W<p��0�"�y�����%Pq�ְwjN��uC9�yri\*ne���iֈSz���ecI�y�e��*'<-�0l��OLѸ%����yB$� S�%#c�� m�yȅ�*�y��ٱ;����u%K�g�F�A$�yB��;۞`y5��N���;�#��y"�ʶ�0ē `�@��]�`e��y
So#@�@� A�:Q�f����ybN�$h��Q���U��pv-���y��:U��ZWo�A&-��N��y���4�hr�+9��hX� ^��y�MN��}HĮ�I|$ɠ�
��yr`�r�\|���;B�j���R��y�!XzbY��'0����� ]��y� �|�f��TMY�{�x� W�ص�yB�F`3Pb���h༰!i�(�y�p��z�� �p2� ���y
� ����D/�lt��b��*�~�P�"O�$�Qo5�"Кf
ΐa�6� �"O����$�b�u R膙b��x{�"O4}�d��=6]
��$���'y��sd"O������h��C�Q=Ch8M�B"O��:��1}�r��w�-Ze��B "O�,!�/������;;��e�"O�����$k��\x��S�\�l��S"OlJ���|W�K�m��6K�"Oʩ1��T@��%���J��}p"O2} �I֔% ���@ *uxHX�"O�h$�F#V�0y��n�3`ԕ�3"O�Y�D�V.=ERչB��Mr`�j�"O��{4ɝ�x
r\"2'JR}��"O*��&N��8�0��J�� J�-2"O�1���v���D�
�@��Q"Orܨ��;1�yE@�]�n��B"O(��b慌\N	��>ry�(�e"OXI�S`�y�]Cw xP�}2��4:b����|������8|�F�v������!D��:��yc�d��
[��p��o|��`sόn�C��,�R����O E�̣G#;\O0I�s倐*�����Lx�ԉ$ժvN��W�C%D�q�"O��"���|����$AJ�$!�d&��D�#["}a�,4P8��^t�$�HᤜT�<A7�E�z�����ƈa7V}b�C�q�B��
��.��	�9Q>˓Nb��k禝8&�|� �E�dy
X��z[���#�(�3FE�.h|�j����J�:aa{r�S/^K��h6,�-:\��b���p=�"k��/�����E�<�M{@�S$XP򯁝r'�!���T�<qg��*d����$����h4NFd�T�vJ�c9n�D1��Ɇ$��h����]OVD�UȔ+D�h�@aB^O��h��ē�g�����`;�Ȇ��:#�0�!f�z؄�'�`G�,O��`�a	E�zH��B>cnC�i�><��H_(��|"$�
V�]p��<ڨu�e�MS�*�=	+tU��`{�(r
�4���Z�ݦi+�ő����m�71d�@j�+��q�4Ig -��=�0ʓsت�'8�V���MF�h���V(D���hА��t4Od XU/I(���9���ئ���,N`z!��.Yq\4z�"O��ya[���fi�Y}��"4)]����1� b�2�	�@��!���R�u�~첑G��G��X�3�-|O �I��
7;{� B�4,xT*V�ۡ!Qv�;�cь =���E�g�-Jbŗ{��c�U����#�C=,�E�&�Ig�|�p o%/ E�5[�b,6+��|��(ź7��Qz�O���Qp ���y2/e�yx�@5��� �%vN�2!$U��$ʺsVp��.��O�m����&��n{�E����E!��3°q�DAv�|��\�V�� [ql�Oi�1�l؟�{��O��m��቞]P����M�s�d��D��0Y����<N�~ �uꁟ�M���S�8�Q�����iZ���'B��q�U��h�zp��	XL�է��n/tu�DH�3�����#&ո��9�B�Ov}�d���	�<c"�0A�.��!�%]j�!�d�	m����d�^�;������ޤ��f�O��O?�	8>V�=а�D6;l����R?,6�C�	�F�����:�ƼJ�NB,�D�������$�'8��z%�%d|}��I�Y��$)�'TZ�sa�NJ��	!�愆i���r�O��bM��p=��&��1��Q�G���@F�dx�� 拥KoV�`�B� l��e��ա�N-q0��[�<	��-r�x���"g�D@���_X�'��A�F�l8��E�d�[�O^�3��]Y�<ٷ�.�����3-@�y��ئ�1 Z'1�� W�>E�ܴu۞�	wf�z��b�D��9R�����p�Z�$U%��ɪY��F��%��y� ���&B[�djN�,�'��}6�Kv�'a�m�r��'��w+ݹ yTIcH�%T�(�b04�� 
 V�׾���iĢ��z`�1v
@cG|�Ob�vJ�gIf��p�8}"Lt���4��Z�\H�眽dzŻu�54������<xd�����3��,k�+/H��s�;*xF((K�����s^�b>7�Vt]dt��P\�D��a�$Fa�y�I�X�l���d}�(+z]DT�w�КM5��H5�ȼ����<I��p����*��<q��g�t$�v�X�fb�ƭ�U��!av����Kq��EÆAʊ&��MOٰ9�ǧC�@^��؁�=D�ȧF�o�%�,_�'��ݐ��z`j��N���QK������3�i��rc��U!Hi���t `)[�O#4� �6&�h{")܂��̺ �ؼbFtX�@7%�a}2B��3��y���4}�~���\��<��G�6x�j��Q�>iE���y\�����|U�h���Q�<��B$_*%3��"-Θ���C[R�I",˔����`�?ek��A�*�J�r3D�|�6hH��:D�<�'��
^\���%��1W�"Mtv'��!�?�g~���&c���1m�+� 0��hS	�yj�1M#ZD;E�[�!�-�����m�����4�0?��C�y-dA(�-
4_��d��K�<ǌ��}U�,2L*chh@�{�<��[(�:�l
�R��\b`��x�<��k��R,RTؑ+U"+e��Za^a�<�5 ?4� %�c��_|b,p�Gk�<-E5dQ�GfښXA�P���ۇf5�C�I�����&%�E��$stȘ�J�C��+�8A#��A>��#`�1 vB�	LAt�Z��e�@�K��fk0B�I�D8*�s�S��@�cF�2��˓LW8@B#)/�)ʧ VP�8��W�R2T�K�87e�ȓP/tx�d�b�hs!��7qBX%����F�wk怄�	�XD59R��6^.ŠP!��B����$V0|)�Ɂa�t���E?>�L)˅���@�'-��9F
n��K��D	I>�� �J S_-���7�8B��1�����2Y�rc����s]\+��턤�A�|�F���5-R|�$�G$[�����G�W2��09,�b�dF}:.�/�Y*�����OY�������� �2�h������'fqq�B�a�ƭ�O	4S�F<,�Ji�)q�Ȭ �` 2��S8W��%�TI�����%�Z!Y�.��?�O����4FC��Kmhv:���Ɇt"H����?�6G	g�D�g",O.��f�@mD�x��.xw"����:j���QtFU�E�R�Ү+U0�������(A%�&(��i��$Fd���H�~-k�o�7B�Ĺ��)9����}q�	ZU.Ϳ*ZN��]�W����[ ��O2�M e�+m� ҫ��K�h@��'� �PpB�} ���C˭KP��#X!�wAû8�Ȓ��A��ħs5x|%�|��%ԑ�rzvN)X\1Ia� �O
t��e�e�%���a�� F�>A4��'�<y8���3�����#hI�D���ŕK����T�����ʪN�Uk�ƔW���� �q[��H3&E4W�hB�	-W�(��j
>tA�`ϝ"�f�>�W��x��"|�`l�%�N�꧉ͅ[�@=�0�ZS�<iVA	�m���q��^�29| �uh�t�<w��$/;�Us����6�����u�<)#��<���6F�/올�ENv�<Ѧ�ah���P�}�$hk'�Qs�<q�f���:z8��뤈��2�HC��00��Ո����cl�B�օ�:C��TGt��F�lQ��R�W�]}C�ɷz(�p��	/}?F� $��j�B�I=HCl�`�Ύ!dz$ٕNJ"�<C�I�Cj��c�C�Gq"pS��ˌ'5�B�	��$ c��QS��yv���g��B�	3}�PT�!N4-��!9����C"O�����A�i`�(A΂�pT��"O�����RtձF�;q�$�d"ON����<8D2�M��qH�#�"O� �]�c*9$Vq��-/bsv��c"O��j� �>�6��@�N�PV��y�"OLax%��Y��pI���-^ ��c"O�1���� ��da����xuha"OF�
�)Bռ�2 ��p�I�"O
1 ҅/�����ED�f��?D�����H<Q{��P-Z#����&!D�����ڔ> 4�k#��0�0X� <D�X7A�?T���
��a���s$*O",R1'ܳ'����B�q�x�U"Od�!�M�$�bݩ� �8e���Z"O�����v�����A�i��J%"O�acoͺp�2=0s/��+W�8�"O@I@�R0�1J' �*zI�=A�"O��f�W*C�x�\#D��"O�`�$
P@0�ae˘�y�@0""O�a� ΀B貜 d���w��$��"O��a�nݲJx4�1a/����"O8u2�-/x�В쑝G���
�"O��:v�L�_����ƋD�A��"O^�R�g�;-,$�$͐�V�� "O5�aa�S ia�lÖI\D��"O�98aƪ2��A�CŃ�$B��"O
�B��-�8�DޝG h��"O���wN�-����E�ɤ[�2L�4"O0�0AO/n$�(b�o�� QA"O �c��Ú~otq��A�R��0�"O�]�r�%װ��BG��FM��c"O�b$`պJp�ٓPf��9b�h"O|���H�~�r��Q�EłU��"Oր����3#�Պ��$JM�`��ɣ�~��iY!`{<HW��4_n%C!D%qV1Ol!K1�'��LQ2��#1<r�S��Bs��[
�';t9��֖A�a�?bZ��O���dΞR=N�LH:3+*U)��@}��G�*�q�V�N�m>8`�hB[:��'�铺0|�!<��R؆6�q$�M?�I�D{2��<���N=/5�4�'eX�YDAR�+X�	,�y��i��С��P�O��,x��*KG�0Ӕ�C+A^ܴ�Z�\2Ҧ�f?y�.�?�J�g}�U>a@��)_O\0�O' �t9��tl�������TJR%���2��߂>��X�#�Y�
�&�	�S���f�(��i�|Q�P��H�&d���7@��~ꛆ�0��$�?�F�I~�S���D�(��_�x2�FA���'��	�{K�?M24fP�Tl�q[2jA��8	�(?�D�¦Q�=�'�zX��5i�H 蘪�o�
�h��q�T���)���H<�O
�O��Lz�k�	-�ȼK�a���������$W�T�lZw�<��'~a���gF(�
TU� 0,��!1n:Hyv��)@$�D�>E����a�%k����$��ض�81����[� ��(�����$!���v���xa�ܲPa˩�H{cb�����-�d`+Q��	aw�m�O|��cMJ?Uy(X���1n���:צ�[��µ]l�姨��I3������`�?P��b��#�PR��� �??1J~
u��4˭T��d�M�CɈ����2��B��6A��	�E]^�ᓉĂ���͛�`� qb�>/�:��P�� )R�q!t���#���Bp�I;�.X��	5,��P�Y����ʶO�eQ@Ʋ�0|��A��1B��#�~hۖ�����Q V��"}��37�v��"'�bu`�����c�<	��H3d�<Ak�k�#��R `�<������ڗ���L3<M�@IT�<�&�"lJb|S��o!���5�h�<	"C�,c���7/J�woҍ��~�<�eF8t����vȇ�Nݶ耳N�w�<����B�tkG�Q�M�.|h�ML�<��z���I` ������ TR�<!���?����F�Q�1�K�<� h�:�H�4"D����J" ��)�"O��r& ��~�~ �M�L��2"O��C�تX��ao[*=��Q$"O$���E�h*�q��G�;<���"O�� R�7��`#� ��v�R"O�)[�$�!k��Xx�n�53j���"O:0��Q�P�y:�Q:h�`#"OlQP3�D�	�
Ysǅ�s�Dв"O����e'x=�E
y�贉�"O0A�"LX�%`t���-��]�P"O��"0�G1�ܠ��$Ƈ#�L9@"O �ȶd(�@��,o���y�"OhX;Gm�9^%�3���h-P��"On��'�;<9�-�<&Ȍ�[e"O>��� �`�,a(���"O�PS���
j����d��:d"O&�ȆA׎8i��!	�^,��"O����Ԯ0�8���Μ#jڮ�"1"O�	P��^&p�eYn�	n8AJ�"Ou�R)Rx?���>M��pp"O�K2�!�N�@�_"K�D	�d"O�rE�!�P�Ј�P}����"Ol���
�,�N��h]2#n����"O���\>q��T��mW"�"O�@0T���M>�|hƈ>"&��"O^y�S&�����1�R��"O p�r�H�|�< ���r��� "O=�l����pi�� �r��"O1'�	/_�`�E
�3pܒr"O��B ػu���aS�D�S�Z"O6�"�T2�1���3%A�i9Q"O.1�P��kPb��fJR�
^�H"Opqwh(!ht�ںHָ�;7"O���B�*Q8	iץ��dpt"O��3�(��͙��ĪU�-��"O�-3C�� �VIj`G���d�T"O���I�����ďΩ��E1�"O��֡��q�� ��뒘Y�����"O<���@r>�E��I���@q�"O29��h�:	�x�jti��6�Y(�"O̍ӪP�H�1��k��I{"Oj��&�*>��l���)�Ƽ"�"O蠹�<8@lcWM����ʷ"O��I6ef����+����i"O�	�A��c�na���%��"O�j�(�>ݩI�c�xr#"O4�b!X9rڤ�bh�IP\��"O��d썂H-:4"%��>X;ʙ��"O�e��*�)錍k�׼e*$�b�"O��!0 ���!�*U>�@:"O�(���*i�����͵'�ԓt"O �"v�FU�������
��"OAPTŘVh��X�iؾ ���"Oj	sj�
M�tpZ�*^�A�lu�f"O�y�#F]s�WJ6db�8t"O��Gi�<}�-%(�s؛"One�U�ѡj�x��(M:3YL]8s"O6���O������Ŕ(FD��"OD�a�Q�N�Nx��ŐN	���"O>,y� N�HR�)�t�͝f l"�"O6�!b��ql��Y #����"Oԙ��e��Q4B�y%��= VТ�"OH%ʆƐ�M�X$ˣ��"y4��"O�A�����s���:s�i@�"O� �����8O�� `A
�u�q�D"O!Q� P���yX���"b�"O00�tHR ��(֮����AX2"O�� �Z���Q��'�D3�"Ođ��C#eo�8Bgڮc�<;v"OX�Y�G��a�A+��f�H�v"O�Y���]�«��Dȶ!�6"O�Y:4D(H�B09�!J�!���15"OhըEV3y�����?:Ĳ�s�"OJ}9g$�6%9!Ś!Z�|��$"O2l��`��TV�iRF�'��̲Q"O:}+PFбk���{�Hԗ�x�B�"O.H�Ĉ:K���Q(�
>���� "Od�d�ҟx����!� �,:V"O�M��<z�ܡ�a\�Xi��"O�iA��4�<d;U�!Pip�v"Ot��O�'�t-��P�Da��"O��CeɍX�� &���&���b"O�q��f�'<��R��åb9��b"O��
f�U?,.8:&�W"k%"O2�!�
��e`��H�SN��0�"O�5�PlǑe�L؊�bZ$�T3�"O�d�B3Vހ!#��E#3x�m�T"OX��2��/��ƩN���"O8�	z�.���Ea�V5��"Ot���a�_�n����+}��4�6"O:� g���g��}��횙&���b�"O����M��^�	Lo�6�A�"O��!n����J�."�nUc7"O�cf�5ܔ��1 �c�(�k�"O���-I#<�8�E�5o��tx$"O����L�XwN�3�Z���B"O�фi�8&�]V'��tބ	�&"O͡�)%��S�' + ��k�"OV����2���1CFH�\-i�"Oha��)�n^�ZA�?q@, �"OͪA╁$��M��hE�q/�X"O&��Å���.@����# &�8�"OT��%��<���Au� *$1�s"O:,���U��
E 7����"O�"P]���7n�'��l�6"O�������kzPMs����b��d"Ob��7l\�qv<D���<�<<2c"O����P5[��Y�!&�-d|�u�s"O�Q�F�E0�0ğ�gj*�1�"O�}���bg`��"�'<�@1"O"��$��)���خ#b���"O�$��*����5㕈�>�G"OztA�	[5�i��g�,i��):4"O����N/����AG̞3nX���"O����-����LRa1�0�3"OZ���PG=T��
�1Cr�(H7"O�٢4e�>RN��J�	K_X`'"O| W�U-��\H��<2���"O,X)�FT�%n���MP�{Ll�"O�0s�B�eG-�vkƓ#Q��R�"O��)sㄬ�X���
�N8��"O��C�J��Y�Xc�ށj"�$�"O
�:�cL9 �aB��F9�pT"O8������,��Ǡƫr�$�"O�	�N�
�݋6�"I�j1;g"O"����\56I�H/(e�����"O@% 2��NR�PЮ!G��0�6"Oh����>���dMS*=o
��"O� ���!G].9����N�H^�싄"O dqs	��W��<�d����؃�"O��p`��5�C�H&<��a�d"O���Ra]H� Qf�(� "O�#E��[��s�l1bG�Q�p"O�DF<�t��@�C5�LA�S"OF���Cؑ��a��P�Z�T1{�"O ���@�T�T�
R&~�T�$"O �5��4'���dS�3�4��b"O��9b� ����{���
E�@�"O(����I�C%,�����X�n�QD"O�ya����P�)4!� ���"OXջPC�7_�u`7b�]�|�1"O.�)���{I�`�"I�z�%b�"O8|X��B1�U(�'2Ԉ1�u"O�(����B�L��К0�Te�5"O ��U�&� iG�CԼ��&"O\�6"�(t�����%�14��e�s"O��1���di���DA�O��q&"O�9�ḣ'ک����K�ļ��"O��aleo.���BU�~�Dy�b"O���#���~x��҃S�n &a�"O�}���D"Z����!��e�� Z "O�qM%R_�R jT�v�*dk�"O4�"����dړ��­ �"O�|B��	~ς�@��Un&� %"O�@`F�2	�P\�7)�n��T��"O���2�R�C�t!(GaE�x�	c"O�ۧ)�n�{�m��q_����"Ozqg,^�Dо1[g�I�0NJ��@"O��R�6z`�"C1VZ��A"O�Ya�.N����(��ko0��"O�[�a]��Z��[�PN�) �"O"]NjG&��		C���C"O�3�J����lE$r4��"ORT�w)K���j����`�*�"O4�si��]���B��O�f1v=��"O�*�e�
R���p�O�����j"O��r#��9�F=��n\�,a6"O1�V����0����ZR��1"O��7�C�p�}ɕ��W��xAB"Oh���h�J�J���D�&��u"OE���Q|ȩ�lY���h�b"O,��ƎN/j�����Ϫ9���"O�S�NH�X�$�*��Ǜ��Pc
�'f��X�e��4��A�Z�z���' .��#y���7�P=U�����'$j%AjֈUPp�$̞�]/&���',Ա�>1�<J�P�Q��	�'~��	��f��bǮZ�I^`}��'E`�aDℽf�I`���:���'�f\�P#G}�hǀ�:�����'��q�`��t����%=+*M�
�'2���������테V��e)
�'��(A@ªv�n8��+_5Sd�=

�'���6�_G���CBN�1R����	�'�X!`v��~v��dC�N�B��'�¸{S+�S�l� B8F�D1A	�'R�1aG�~TI�u�
FN~]��'Bt�z  ���   �  C  �  �  �*  G6  �A  �M  JY  d  |o  �z  7�  ��  ��  $�  z�  �  l�  ��  ��  @�  ��  ��  X�  ��  �  e�  ��  R�  � $	 h � � b# ?* �4 e= �C 9L �T �[ �a 2h rl  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�h���%k�2�8�!#$>=�B��PX
`���*�M���y�' $HBR��,�O�o�b-��'�2P�&�����dΧ)����~�D��	[�\�2f$�*�B�Yé�]��?Q+On�}�2aX�n�<�ah��nY>jE��+�V�R?��'P���nzޑ�R��
ks8D贀E*b����!	ٟ��	�<��O1�XYل&mӐ�I�&]��T�c�>@�0`�n�L���<1��'��F{�O�bH_18���T��t���b���yr\�8$�x2޴n�>��<!�&	��TME�>`t�9r�����'�듰?���y*���Q�(��Bu�X80�̈́51�9����I��Z$Zch9�S�rhY��H"��^'*�L�"��>L�b��dyX�H�)��<�����m# +$:�!�PE�<�c�i|8�k�Ot=m�_��|2��-!����ӥW*;]S�#S�<���?��
�p��4���m>����L���  �U�v�KE�D�^�4���@*��<ͧ�?y���?q���?�2阊x�n�  iX�r���r�>��$����d%�Ty��'���A��:� #�B�%j��0j��n}�h{�4n����|��'��N� d@�܈#S)w!t�8p��/9�X��d���?!b�� v��n���ug.�dPy�&�1?�n䠢�ƅ~C �5�_YS2�'���'j�O����M�"��,�?�ELW�E����ɐ;d6���Q���<)��i^�O!�'Hb6M���:޴6����B�V|�0��%N05��\��O��M��'Ѱ�	��P�+y|yxc�:Z�B�OO����w}�
�	R�}`<�jФ�<]�"��'���'��'%b�'8�<��� +�� o�xAVDa��O���O`�mږGi.y�'N�7M6��O>��lK��E�H���0Í7r���'�n���M��'vk�Y�ٴ�y��'|�Q�d4TL��V'�dI��K:XTT�	O��	)�M�*O���O��d�O��Je��1�� �S"��h�O��d�<��i������')2�' 哿0�[0'���q�Z�	��M�I,�M��i�O�� �`��A��g��(i��=?56�h��3?�Izv�=?��������V��Ӽ�d��S�(�0�C (�4p� "�?����?���?�|j+O��n��^$�-X��O.?d@
�P¨�^By�lh���<
�OԈm�<$A,D�e�F��6$0�)F�$K��Kڴ����L��;Od�$�/37��x��K1��E/��r�g�Q�P������8P�Y�4����O,�D�O�$�O���|��ē�kԄB���M��@�'r���VP���'yB���'76=�
�CU����tψ�W>h�Y�Ɗ�E�B�'��O1�vHju�o��$�J���b�u�$�KSʁd ��ix��P'�'���''�7�<ͧ�?i�+$���uʃ�;��}�0
�;�?���?����$Ǧ5�Se�Py��'N	2�@`|�c��):��ع��d^}��'��d=�7�Jd3���Ea����f��.T��O��Fӆ���R���	]w�4h�I�j\B���=>�ɋ��7S�൰���3Rb�'���''�S>]�0"+:�J��<�2���r��@ܹ�<��� ��f�B�創�Mc��w����#���2�b��C�ӟd[^ ��'M�&f��|n~�HynZ�<y�2�^${���D���,_/lF�-��	ӳF��5ӂd!����=�����'��'b�'ޕ���σYe`�� Q�f{�1�RT��@ܴU�1�+O���,�әr��7�,b]S���=L���8�O`=lڕ�M���x�O����O�x��&�Z�ff����b�&��t�������c�O��iD���?	��<��i�I�eS Y�FgT�n���D�@�y����͟��	��i>��'�Z���5#wr*Cˌ��/�<(L�&T��yR�h���3*O*�t�JIl��r�@p��A@,:�,�#O;-�|��A)�����?����l���@~Rjk���=� B$ے�NG@�j��~���f2O����O����Ov��O��?%���]�?5���ShA$,| �D�F����ڟ0��4R����'�?	��i�'� } ��֓G�����_�)`.�鷟|�fӸDl���L����	�+���h��]{��`��Q�$�P�&�_?��K��Oʦ'�\".O����O��d�O@�Rkb�xR�_��B�(�O��ĭ<�ƻi!���V�'k�'��	?��U�����E �c��[�;���#�Iğ��Id�)�Q,?�d�+�L?Q���;��U�b��sc�x����TƆ�3�|�%�t�у��4��'hѾE���'uR�'����T�ߴHi:8�D����(-J�j�Ku�ʓ����y�?�X�$�	�Ne�ň��E���ܰE�3^��q��ٟ�'�ʦ���?�)��p���_i~R�9Z�N�scl��!4�]��鐟�yb_���I�,������	ȟ��OƆ$��@/��(���Q��y�io�؜r�e�O����O������Iܦ�]�m�S��Ȋ_26�P��R��.T�� �Io�����pB�nq�:�ɎJ����"V�>��ysďw�0��+<�b��S�'N��%���'r��'a�	"��I$4|r�gO	O`((��'Wb9���'m2W�ȳ[wUzqz�V�T������Ar�oVJ8��S�h& �?�0]�R�4X��x�K�2�X�{��7��09�e3�yr�'��xsnͳBAf�gT����>7�¬�ßP1�ɖ�z�jӡ�Q	i� e&RП��I��(�I՟�E�4�'�Hȑ&��@0X��"MF'���K��'�,7��_Y��d�O��l�r�ӼCG�M#nF,�G*  D�u[��D�<�@�i9L��h��5ey��F�t��a��4���G1!zD�*'N>(�3�?�䓎�$�OH���O����O>�D$/�,Y`�+V0[�V�h�꓊7��t��61W���'�R�Ʌ�d�����Z#|���0����ؐ�'V��'ɧ���'B�EJ�Ҥ`GG�1T��!��$�Q��imx�&�8xHP ���%�0�'0��bJ1|��EIW01A�@�P�'�b�'�2���t^��ڴ-DrH���_6�8�	�-�D�R��ۗ=�������M|}��';�w4��I�� r�qIdm;0��8��Z�PV6O�d�pVv�s�O��	�?����Fu82l'Kp�<��ɫ>)��	ǟ��I��`�������t�''_��r�)~O�m�#�IF�c*O��� ¦���?�մi�'��(eI��qD��(B��$Nې�|B�'�B�'H��0w�i����O^͛R���G>��a!��&
\�A�T�lR����O���|����?q�yfr�i3!P�`~h9��L�5�����?i,O�ToZ�]��`�������?��ӊ��pr&��i��Tٷ�X�_��N��I矬�	f�i>	���_�<�ȶ���x,��Ƀ�7�J��e�C"yv�x� �"?���L���υ���Q���ؑD�>X��k��a���?���?��S�'��d�ʦ�Ʈ
3���@ů�J�H�@�M�<僧�	̟���4��'=(�8{����	/�m���=�z%t��2�7M��y������?Y�n¿y}��ɘ���D�h���xǃ�6��<C�gX��<����?����?���?9+�P��p 4>��}j��� @q.X�`%����]��h�	ǟ�$?a�I�M�;`��$�}R�]k��Й=�>� 1�iR��*�4���	���t���k�p�	�L�l��"��;6��7 ��<����7��풓�'�%���'F��'w2�B�+�QNa�f��%��T�'���'w�[���4 ���+Ot��6��D�V���aN��SD΢!#���H�OLnZ-�?�O<�"i،T�)%㟩o�����c~J�SGx���#ƨ�O\r��	�PR��UD��7&�9�2}Ɂ�O��B�'B�'���S�����e��ni�׆P�0�<B�%������&
��'��7m%�i�M�#.��i�e�fE�<A�(��G{���������:B�>�n�<���z��)�B���%�G,�A #$�B�0J�]���1����4�t�D�O����O����dj�h)���Ȭ�Gڛi���v����8�"�'z���'>ƭ�6+ �������T�x��E��'�>���i�L7MRt�i>����?�Zr�a�^!���N�����HV�8@,���%?!%��,
r��䘋����I�<D]��@9T�B�8�`Q#����OX���O��4�.˓'�e\(H�L�1fh d��aŴY\���C��B`�8��+�d@}�'o�"`�	�]ZV����}�2-�	]>|�`đ,`�nZ�<y���p�L㟔��.O�i��TD��GSf�#��_�=��B�3Ox���O����O���O��?�rz�HBF�"j�4��&B៰�I�Pcߴ,�@̧�?���i��'�*1�Ǹ^�N�jC\= ��阷!1�$|�,�o��?m�E���Γ�?��hE�,�d��B��K��x��9�"`#2��O`��N>*O���O.���O�� sj̻V `a��"��B������O����<9ŷi�8�1�'�"�'�哲:'lIц
�N��r{�h�1��	����	v����)޼b�@��T�&V������x���kr)�VĦ`�qͲ<a��q2F�Dǵ�'�
MPa��$�����ɑ��0[���?���?!�Ş��DW������P�r�y ,]صA�!,������$�K�O���'�6mM�9��ta�cĵ~��U:��)[���nZ��MքG��Mk�'�"��%:���S;��� ��a��k_��B� ���0:O��?Q���?!��?�����<tD�Ӂ�>R�H}��lF�g}�,o��P8��I���	D�s��9���cЗ R����d�1qj��� kF �lj�(5%����?�S%e}��lZ�<aQMʉ#t�0�m�7)�����
�<1"�.ؘ���!�䓯�4� �D��1��KBK�c�0`�p�@d�p�d�O����O>�A���#w&��'���E��F��vi�%j�8���BN�h��O���'dr�'��'_t���׬hOfӒ+!"r���'C2f%-,N�P�eY���$�z�*�����d 8��͑'�(R���4�Ѐ\�����O��d�Oz�d2ڧ�?��CNu�<��� ��4�C�9�?�u�i��*Q�'R�g�f��ݜyB��w�
�P0�[U�T�B]X��P�	�<��Ц	�u���(B_����{��@x�Ye\Z7;,��Oʓ�?����?����?��G�*�Sv��>[�<9Ҍʞk^-.Oޥl�8x}�L�����l�S��b��]5�)я�;
Q�Q�����O ��(�4�����O2� �g��k:0\2vh� X0@4a��K=Xd6mTy2��wU��������$^�cR���
�36��h�r��]L��d�Ol�d�O�4�$�	"��"ʤ&���Ҟ����`�Q�g����&�Ѐx��m���(j�O��D�O�NG��tHG-�.8�Di�kœL��vHkӪ�I��xr�_�*��)�<������h�'0N��� �^=�x����<q��?9��?���?���Z4{ F�rK� ;H�9�g,*�B�'���{����V�<��i�'����7e�W�l=jt�ب��*a��'wd7�V�M���w��io�<���g���{3��h��LA���$a
.wGXՁ6�'n��%�ؕ����'��'�.���X�9$�D�  X(r&�(��'[�W��X�4$������?I�����"��q���7U��;7�������������Z�4dމ��)�=L*%ppL:T���eK�&}H��d�!��Q����,E���Z��4@%�9��%6�ε�U�U$T/��I���I⟈�)��oy�w�xL���5pkȨ�����NiK�@��4ʓ =�V�d�O}B�'��ĸe��i��	�fl�(W�*�Q��'���V��2O��^��vA;�'T��	�b)8!_OY���q"��M�v�	By��' ��'�'�"P>�g��N4���:c�����`�Ms��?I��?AJ~����w��"�#�$(V02B-i:
D��']"�|�Oo��'� �aǰi#�D\"y�`AQ'��y�H@�ꜷ8��D]2�L����̓O���|�����|;��&/�`x�"/V�0J��?Q��?�,ORl��{h�	��	%*Ol,��DψGҵ�)ԅ,�`�?�S����П�$���'���_���@�1��ِ�x�\�	Q�Qj3'R yԊ�����O���$�,�*����
�H[b�V�*T����?Q��?����h���$ 
�d���YU���H��&u��DŦ!��V]y2I`����$uF,z3��!!�>���"J�x�<��
�M{3�i��7�[0Ed46Mt���	�n�� ���OF"p$N�;g�4�Ђ�+m�"�ëa�	ky�O��'���'��.]/F���lE!y�ǫ��I��Mk�m���?���?N~�0G��Xs"��~�z�B�:x	neQT�tk�49���o!�4������]k�⍡'����U�&��b��3��*"��d1uE�g�D�@��IyrFY֌��.�!�x%"V�(1A�'���'U�O��	(�M�����?��	W�8	.�9C�~ �	�#*�<���id�O�$�'#�i�<7��<w�qy��E;$֨�PI�L�l���b}Ӱ��ϟ<C#@U�^~�T*;?Q�'ƿKu���y�`�uH�f&�����<q��?���?����?!��!�%R��Ax&��g�D��N����'��Ns�vtk��<E�i��'KҘku�\�0M��j�*L4EM���d-��	ئ�j��?���ݦ��'OҸiEi��p��S�7����sf*@��$��+9��'��I��T�	ȟp��!
^����ʟyI$\���4K*����'�l6-̬.�L���O��ĺ|:��S�Ҡ��QoH�pP�UyGƖ[~b�>y`�ig6�:�?m2A�>7()���Q�BY:EB��'<Jղ�B�[�4����jBȟ�{@�|"NI�7�}��-�M~�����Y���'�2�'8��$P���4yk�ԁab�{��4R,�#Y�� p6��?����$p}�&x�|\�qŗ?!w�Љ�.~ׂ�c��V����ߴa�T�#�4�y��'��)��$��?ͻ�X�h��,�{��p�cZ!����2�~��'�r�'���'�'�y+l����]%���@^�: ��Q޴I,D�����?������<�w��yG㕾Ȏs���(A>h���	���'�ɧ�$�'��oVX��;OX���@�Xx�����V�
�Y�2O�
����?9� ���<�'�?9��P�H��X 3m�����̀�?i���?1�����˦�⁬�����	��p�H^�s�@ؚ��T:^^m���f��l��I����z�ɠ5�$M@�[�9q�Ar�7b��	ן(��!Q��ڄoڿ��$��)��'��kN6:(�Q�#s3X8Pg9y���'i��'Ib�sޅi҅��O��p���3��A��oڟ�8�4Rl��+OF<m�I�Ӽ#�K(&|ࣔ�L4 �c"�V�<����?	��0j�]"�4�yBџ��2��?� �]�@�~�T��ه�$��l7�$�<����?9��?���?ɠ�M�FH���J�:(Ov��'�0���妡�#!N����	���:�h_2N��d�S�_�BX�ޡR�����|�	`�i>U���xz���4h�+�	�o�����%Ա,��HnZ��d��aY�'��'��I�
����i6rx�E�*Q�p��؟��	����i>)�'�r7m:NL�D�6B�Ёi�טo�<���E�nK0�$�ئ��?V����4G؛){�J�1��D.@��	i�ɛ5"�DE�#��_�6M#?9�s�I1���A�Ȉ�^�f�ZiX�X7E�y2�'�'
��'���i��>&��YE
�1H�@ؠ�Y��O��d�O�)o-n4��'R�7M>��I�q��y``�J*g�h�6�� ��&����4!��OҬ��S�i����O����Ei�f�3' ۰zs|S�	MC�j��v��Ob��|R��?)�] (�3�5.�hE�)R�c��?a*O�m)D�Y��ҟ���J���Y? ڞ];#�  �"������d�j}�+|Ӵ9�Is�i>y��R&�9�H5b�J��!iS�	$ԩ*媁�`=�A"V�Xy��O����2)�'�<��D��Kuf�9A+5\���R��'rb�'����O���0�MK�W6}�p)^I�hTނ7"���O�������?�bP��;�4ilؑ�d�W7���ApK��{�R�Ӷi�(6툶E~�6mu����%
7����O}T��'���[&�aK�x����
7*���'��I�x�����	ן4�IO��L���X�P��+0.h����	Y��6�
��D�O���9�	�O2Tlz�E��Y�2��@���֔�D�R�M��'���t�O���dK�#�F1O�X	� �;R*��H� �'Y�!�1Oj�c�"��?	�E4���<��?�ǂʔ"ᤤa�bN:[4ACl���?	���?�����G��咠̟����\�3K,P�p���\)qrr�Z�́T��~��	̟���i�aش����Y&.�A �i�)��	�X�d\&p\l� ����&�K�'�"c��D�b����R��rŦ]eR�'D��'I��͟TG��3yJ$�3$ą=t���b��XR޴DMԀ���?�4�i��O��̆?���O.e�����DO2p��=Γ�?���?��Z��M��'���B�w���SrjXdk�N��w��|����%>�q$�h�'�'�"�'�R�' ]����U�E�ȕ�:^u#T�PIߴ{�N�I��?	����O��p���,\5J(�ā�+1�R|ӂ��>���?�O>ͧ�?��_���S�&Y�̒3��14�J���M۠_�����'�d6�Ĩ<9R
\:9f�AH@�=�h������?���?y��?ͧ����妑�n]џ����4_�2�c�2�V��|�t��4��'�|��?���?�f3"S4��]�N�=���^��sش�y2�'���F)��?A �OF�I��AZ����"�����!D�_|� =O��O��$�O��D�O�?�Y�L]T��h�/�.!��I��!ݟ���̟���4ud�`�+O��m�x��^*��k���Z(q
��-G||$����ԟ���"4�$�n��<�����0�"0j��<�nO!*<�Ŋ �!
(��$̓����4���D�O^�D���ӀF "�({�gw���D�OD�$���G�r�'�V>AS�l�Ӧȸ�"E.ȨԨ&?�S[�H�	ܟ�&��n!nlR@�V)-x�8�3�%���&<�.���'�C~�On�I�ɘ|�'�-��O�[7�9�'/�?'�ؐ��'���'�2�O�剖�M5�����/�8r̍yEIܲ}n���)OTml�i�t��֟�J1A��r�0}C3�O>^�^��!Lğ�I�"��n�k~B��5L�Ҙ�St�IS8�$%�"�{T���a�t���<Y���?q��?Y���?y*��L��CI"w�@�)��)<�	���ꦉ����؟8���8%?�	��MϻP��\*��س�ꬋ(Ԁ*��	���?yH>�'�?��=��u�ش�yR�45����P���"���c��A�y"i���	;f��'��i>A�ɑ4���{���w�\�p�Cś��E�����	�'�n6�_,z/�$�O4�dM�(��sW"M<�h� T%U���$)�D�e}��x� )n2�ēHS���M�O$�у@�����̓�?�E��*�p� -m~B�ON����8Z����7?4z�ˇ͜Z}Ip�N:�'���'���ß�P	�1�$���+!dL��!^ʟX�ڴ��k-O��n�W�Ӽ�aL�A� �rR��nfZ�b�nS�<��i�H7�٦��\ئ��'���PU��?��Cg�'rY�4I���)p�%��_u�'�i>���|��ҟ��I�(��4`ѩ+��k�N�H�2 �'��6�ΤD�N���O��������<�Dm������.�*�\�Hை�h������nZ ���?q�S�?�6��A~ K�c\e���_�H����7?q�iE�m���$�������8b*�b�&őn-ب������D�O~���Ol�4��қ�j��z�r ���場�Ǔp8���6�y��~��⟰��O�yl��M{#�i�\T"���8���jÞFd<�A�N?��?O����|�൐�'4p�I�?��]B6��aף�^VP�qG�?���Iݟ��	����Iן���X�'U1� ���&8�7a��J��?���:���"�Z����M�K>�%�A=y�H:�K4�� � -[��'��7-Pæ瓝}2T�np~�K���� �������RݡPɂ��|CRJ�)�?��	5�$�<ͧ�?���?�c�X���	�D&s� �p�?���?i�_��|R��Y��?�+��!oz>�a�!��c^~x��摴��!�G�4?�T_����4!N�&�8�4����3o����F��+��N��J��0+�Ô:��p����� (r��P^�80�j���(����q��∙4Ӛ������I��)�by�k���r��]R���ɭ%�SDG�&ʓ��V���m}��c�6����q�	�'(��T<L��I�	�شr�X���4�y��'�4,���P�?��`U�4�ś�=� � '~b����$r��'���'ER�'N��'a�S�YB�\bu���
� �G4&�B���}"@����	Ɵ%?�I��M�;=: �Qt�ܛ_�T�i�,��?ިЄ�ij��$4�4���i����� e��	j� �q0oϣr������Ρm/���{�H'�'�8'�X�'�r�'8��C���#�\{��J�$�k��'�B�'��Z��s�4p	��3���?���K��ڔρEy�V�"A�T��2�3�	���d�����ē�P�s2�ʵH@���T�B�8Mϓ�?��9>��Fj����d�����NR��MVc��IM%I|�!ys�[�q����O��$�O��.�缓�Ɉ?zD�᠕2���8g���?�r�i@f��'�ooӴ��]�i�00�vɿ{������+1L�	�����x��K��eΓ���_+3��B�dI�'��%c[�0�b (H���O���?��?A���?a��]q�Ѡ��;:���&)$j.M9-OZtoZ�W�"	������]��$� Aߟv��)fc�$��2�ɂ����O@�$0�4�\���O�1�dj�	#B�i�������I���0��7MTzy��͙Dh
���䓵���v׊��6L�dm�MS�����N��O|�$�O��4��x��Q�����,�r�3.^��!���)P�Rlg����)O���g�l��&��+Ck�	Jёe-G�>w.U��O�)Γ�?Yևݥ=N(���B~��Oa�&�D�&U2Ft���aC��y��'+"�'TB�'�R��'���k�]�������(�$�O��D����:c�}>��I �M�M>���X��J�(T�s�d�2�+�3z\�'g�7���/l�r�nk~���l��4	�";{�MIB̯}wB���ҟ ���|"X��ڟ����)vn��Gh��%��-��*BJԟ\��dy��o�rm���O.���OD�'��9:��H'k=��4Bų�8��'�~�C��f�p�9%���?���� *f�SEd�"euv�dę�=�z���'UN���@��O�YL>Ԉ�P�P�ޑca���BW1�?���?A��?�|�/O��n��`�4\R�Ά>b�AC���X2Kקw(��O�mS��&h���MK�"�Nxɫ0d�p.��D�0M(�F�i�xMl�D�I�`rB ���i4?ѣ�^����@��m�$PK��<1(O����OL�D�O����O��'�V<��τ�?n^�IK  XXE�2�i<�=���'m��'�Y>����Mϻ&e��ۗ)Ĕ<w0e����`ъ�k���?�K>�'�?�L ���4�yb�Ę>�|��e��!Gdq1�J �yr�G�\�(��������Of��^NR��]� PLx�� /n�^�d�Oj�d�O��I|�n�(�'���O�qΌ̡�텈iGjĻ��D�F�Oz��'���'D�'^@e0��1�����0�p�'����q�~H@�io,��B���|��\�&h�#✥=i����#k3� �	����I؟��IZ�O1��vV��37�M͖mh2�F�(Gb�y�V�H�)�Ob�ā�=�?ͻd*Z�kÇ"��I��hw��̓2��fq�hn.��n��<���$�@&���D�sV,�>O3j!��)VzLMp��Ԍ������OX�D�O4���Oh���F�(|b# �5�* ዟo!�ʓ8�V��[��'Ғ��'0�u�2@N�w�Ӆ�ľv�v��#ǻ>)��i�H�$7�4��������a�#��&Q[p$�g�^��L�n`�,Aq�<Y���kQ����)����5Ct��)�� ��8��:�z���O*���O\�4���r�&�ܝX�r*��6H�oL�(�+���j�*�g�F���F}b�s�VL�����h�J�.
�d�o
2m�8m0瀕�Q��aor~���!V(Ѕ�S�$��O4&�J�|�A񉅯� ��D���yR�'���'��'�2�iK�xx�Ze%V�yD��zd/�Uw��d�Op����E� ��Vy2�a��O*%kN�/�ؒq�B
�͂��2���O��d�O*M��JmӬ�Ix��%�\)3pgG[#b�I��FT��I�'r�'���ܟ���˟D�	�'�*���A/1�"h�(N%x����۟�'̐7-
:�����O���|��	����h�dG6ѡ-�M~"g�<���?!H>�S�?щ&`R&1`������k\����ƍh�&}���0X6�x�'3�4,Nɟ��r�|%
�U�b|�ae��N�p��b��2�'x�'J���X� H۴Iq�ٛ��T��|�CcÔd��dٽ�?Y��42�F�dL}2�'�ʇCA]�
�A �2/�La��'⧒*a�F>O���]������թ��"I�2��Л��X��y[�X���`������	����O�X�Z���C����ˍ<\��5kҌr�X)xg��Ox�d�O"�)�|�]�wtrp�"�[�~�Qc�8Z�$qxAcg�֬m�����|����:&�A��Ms��� ��[�b�8<�DSU�o��̂�<O�7B�i�BM�Z�	^y�O�ү��8���ZZr-"��ׅu���'2�'�I0�MӅkD-�?����?��*)h`���
�ehCh�7��'!�9j�F�q�j�%�䡡�
�-�X�w�{"0�k�8��)}�<�Y�.����OF����?���Ov!B��ߙK�<H�B�j�P�{�&�O��D�O�D�OH�}��/�\x�g�,�D�O�d�R����H���E���'�7M�O�O�|���EAāoq��`�fSMJ��P��*ش"6��M� _�0O�����KiI���y��-�Bg�`�2�h�fTMr�)f�<�$�<�'�?��?��?��)6"д�o�1Vz�B�����d[�	YdϔRy�'���`[ҧU)M'���a�ު?G֭�%ʄv}�'5�|�O�b�'jq���S�O�x�/�=B#�P�>��O��4f���?i�#�Ġ<��S�"#xI�����+�D��?i��?���?ͧ���	ɦy�3���4� E<!��a�D���q��o�ӟ��4��'����?��Ӽ�THT ^��XQ��e��M[�k�)LP8ܰ޴�y�'r�0�h-O$����T�+s�P�v�8�{��ݑ;��d:�7O���O����O8���OT�?m�Uj�G�X�&�);.�	�����������sڴSKf��.O�Io�����'��Z�AV�f�ʤ�D�1u�\�u�|B�'���'8P{E�i�?�[t��2���(
I��A�"�7 ͊H��������O����O��׶TIS�c�`Ӥ�S9�a{���?y)O�lڈr6*<��ʟL�IK�t��K���gN�i���(p��-���Z}r�'�r�|�ORj�"�LԱ��#X���zfB*^�fy*�4oA�#�<�'��	p�
J<�ݺD��?6:$B"hT"9^��I�������,�)�ey2�u���HW(4���\�� �6�	�b���O��lZ��C ��3�M�C�ц���8��${���E�^�_��֠~��p�1ks���΅� 埒�O�PU���0Z�����*�)6��"�'����D�������0�I^�D�NMH�
S�թ&}X;���58��7-Ġ]`����O��$2�9O<oz�]pP���& �ǧHk��"��M{!�'����O����iA�d�uXL+3.WΈ��Ś�	��D��v�H�	��WX>�O@��?���4xL�y�ِzh:�$���Yj�4:���?����?�/O��oچg���I����I;�l�ah%Y�*L/�l���?�]���I�&�`�6Y�H@$��� ���{d�`� �I�H�rb�G�A�'m���ʟ�"��'h�-�t^�)��FC�}�T-���'���''��'&�>���vp�yv��*VM�u%�_Ξq�	��M3$���?A��
�6�4��a�թ�V���o\,���"2O��n��M�7�i�ؑ+b�i��d�O��r%����!�^�`V�߼eI�oޚz �O���?����?q���?���ho9��'l� 0k�
#4Ԥ�,O�nZ�:��I埴��w�s���P/�&c��Ĭ֡������O/����O��>�4�Z�D�OD-r�`�)�(%�fcPt���t�W�lrԀ�"��9���*V�2EHe�Ijy������sB#D+��pV�
-L��'q��'��O��I�?Y6fKן��ׅ�'��I*#g��!�f�ʴ�i�@�ٴ��'�x��?����?���+ei&A˃☉X�l��O�:����ݴ�y��'���q��?e��O����lXjd�ϑc[@���t��j�2O��d�O4��O���O��?��A'\����wK!	�p��&�ޟ`����h�4N
�@̧�?Iտi��'����ND[�5�l,,�,� �|��'Ib�'�H�҅�i��?rKU7mk.�P����vW�E�ĝ�v�V}�����$�O���O0�$ԛ\��i��)
�Rm�Ö�!���d�O6˓w�K��I��'��[>�1a�C�
%�0M�xp���W+#?Y4Q���	���%��ȟ�{�I4S��T2�i�:Xd�0�$��w�T\�A�B8S�t��2�#�O0�ZO>�C- �c��1$iC�Dp����ӿ�?����?��?�|*(OZ�o�a�,����{i��k�m��EH�)���ß�ɪ�Mۊ���>Q��?d<����}!g�@AB�j���?�4$���M˜'�	���ry ݰN��<b�A_�%��� -�=�y�X�@�I��P���4��˟�Oy��9�$U"R娽,J@�O͎F �6M%P�����O���/�9Op�mz��1V A[S�p`�-�b�Af��͟4��G�i>Y��ϟT��VƦ��~w�a`thL�}bĉ��$��D\�5̓G���7�� '�З'���'bf(!pb�/-��@��'4E ���'w�'(2T����4N�Ta��?Q��{�590�I�BNR|�!����E����&��I��0�	l�@r�r�h�bѐԣݢ_'B����8��#�P%�����Qy��OJ���	�#LV��͸�!EznZ5N��}��'^B�'�b��Ο$�T�+41�EB ET%4:$�@%�П؃ڴ~�������?Y��i��O�N�+5��w+�=f�X�!�C�7��ަ�K�46�V���F;OB��	\r�',5(�{bdA�@��%XS^�꒮;�$�<����?���?	��?AG�Ԃ1`�����:��������DŦ!�s��EyB�'9�O�r�	�_��P`��B(u��l�w�[����&�OO1��y[r� ���E�.+�j�CA@ƈ~舜�@@�)���#��"��O�l[I>�*O����oZ�W��ġ�[�M�>H�f.�O��$�O��d�O�	�<��i�X�;�'��]hS���q�E��.;(�aV�'��6�5�	�����O��4��Ѳ���WBl��󣍿Ef���>4'86m8?��:v�(����ߩ S�����Hr�$Ed�ڝ
u�n�,���X���$��ߟ���֥#0F)�@MW�w�0��A���?���?��i��0]�H��4�� HleC�Kэr|8���/�9$��mJ>���?ͧ-�X��ܴ����ek����W�E�f� hg0���ِs����z�xy��'���'��#�"](�(��+9Tn���(ǘ��':�ɵ�M�qkL��?����?i,�����Nj�Y�c�_�H�
���8��O��d�Ol�O�S�L�8�DJ�]CbxêQ�Q��(ʴ�S5�zdn���4��e��'�'v�� p���]5~@
�D�����'���'�2���O��ɋ�M��NAK��x��n]?C����"�9g�� �,O�an�V��F�����MK���$@,�ѫVf����'��t���e�V�i�b�F.��cf�����O���� ��;X(���+	AI�'�	�p�I��x�Işt�	C�t�8y�ڴC��JA�xb'#W�_�7�D���D�Or�d6�	�O���w��la��D�DD�-8�r����5dl�Иl��S�'p>���4�y���s?�ap��T�oFE�g@I��y��� 'SL9��&x�'P�i>y�	?�.�Qǭ�B�y�Sa�4Y^���ٟ��	��h�'?�7m�62����O���KG [ӳ��� ���yw����O��nZ'�M@�xBd�(����LۦB���i��y��'�(ď[4���A�O����7�?���OdQ:�-��e&DI�E �0��]����O����O@�D�O$�}��� %�-)T�_�&VT8Ҥ
�F`Uk�hM�V�
E�ɀ�M��w����'� Mjjd�� ނ;H%1�'22�',"�ۻ<��7O��d�-1^�b����yȳ����N�)a���8!��>���<ͧ�?1���?��?9�ួ�*q�`���Sm՗���Ӧ����ޟ��ȟ�$?牫� ��qFT*�:�2*�}�ΰ[�O���O�O���O���K�~mh�ݼz��a�''Z�f��X��ǆ��ɴ@�*!�d�'إ'�4�'�|A�Y�}$ �U��I�Z@��v���
B�K�B�v����
&rtq�b�"��m���hr�O��$�OB�D�~)��T�5>����G��2�TI�$a�^���Ȩs��?�'?��ݑcq�h�J
+�\ +C������@�� ��
�Q�DQ.W���2�ӟX�	ҟ��ܴDf�4�OP6<���B$���^I�H�
�U�̓O���O��6��6m!?��u$���ȑ!v�𪱧ԦCm��G`ڎ�~�|b]�|�?A��A �Q!T
�����S�';�6�(KG�$�O:�d�|�bL*�bᱶ�H�(��e�R~B)�>	���?�J>�OPX=�tb!J�p]P�m]0��1�U8J<�!J��i+&��|�QN��h'�t�B>��"bL�21�"L�o#���4a㐔�+U5�P(��Ȅm. <��-��?A�w)�����J}��'��P�V��jh�r�(�7|n؊'�'�J΅����֝�jj��'��D	h��];S*R�6gJ(���U��ľ<!	�q`�3tė�h�b�/(>� \ۅ�i��\���'nR�'��|�nz�a�D�<���jFG3*��PE�Ɵ�In�)�8-�(�nZ�<y�+��uxk#�8w����EO�<!QG��3Cj��|�Xy"_�����t�N@�6��z4Q�N>OL@ow��}��՟4�I9�be�H�2b
< �b�@ޑ�?)!X�d���0$�p�A!\�������6���d�)?)rA��p38Uy�4g�O�dx���?1cC4[X`)��nP=��(3l�p�<��G �_xd�ie��5~8h��-]�?9�i��&�'P2Io����]-+����g)�PM����+�j�	ҟ��Iݟ���JϦA�u'�A���iїX�UC �ܥ��d�����O�ʓ��O�y��a�0��]��Ć�n i�ǟ�dz�4'� ���?Q����O�%�U�Z&;���r&b��0K�>���?�H>�|����<m�=�Ĉ�w��R��	�~&����44�I7!��;q�O��O�˓,�X��VNU(:�X��J��o�F����M;uH���?iu�Ȇw=0�3�!�\���
�	��?!��i�O���'8�'�B�ߚk� 4���)/d��gNB�f|Pw�i��ɟ9-��֟����əG� 5�",�Q��:T�$2�OB��A��t�E��-L��ꗤ�O���O(=n�<KԐ�'_�V�|���wI�k̨&J�����'F�����)^0�ƚ�֝�wA����P)f�e��@+x_�Q!�YA?�N>q*O��H�ߌY�,�ӠIL�1[h}!�5����b��~7��'l�U>e��.��hd �a	� l��8� ?&S�$�I���%��g�? �Ȇw�h�����$8�*a�V�P>����g�PQ����N�v?�N>i�crѺ:PD�U�0k$d�P<�D�i�ig��#%O̔*��&��D�6�ݜq���'��7�5��!��d�Oΰؔ�_�[�A�O_5P�x́f��O��M��6%?��l�E	�Ot�n�� �I��h휝Sh]	(�d�I@yb�'aB�'EB�'��P>5�$A\���)֧1�e�����M��
U��?��?!H~��m���w�<H�Iڽ\����bA.5�L�[7`�r@�	Y�)擶T�X,m��<6�#��ɻ�*�,� �r���<q�J�<e����ý����D�O�$��*#Hl{#N�SrR=I�GM����O����O,ʓ����9��'Qrl��~��Am�/�b|�  S1R��O�l�'>�7�R̟�$����J,*�FMI'J
�Π�4�4?��N�% �9�K	��' >�dJ��?��A�a�X�Hr'�f،��q% .�?q��?	��?��	�O`8���.��a�4o����(�O4nڌ x6��I���a�4���yW�T_�j9��BŪ�N����C0�y��'K��'�.�0Q�i?�i��r��pRV�'CW���u@�$���)U�����D�O����O���O��$�IW���tAΥ5Հ8c��ٿ��ʓ���^m���'O�����'�Y(�̩I �͋&�_K�a���>��?AJ>�|Z %�:V�8���%�,6�,c�E��p%���4{P��+.,�#1�O2�O��p��`$L#x'��0�E�$_���ɧ�M3&d��?�A�)I��,�#�W� �c��ز�?Ɇ�i}�O6i�'���'pr�ͅo#n�J�	A4I��0g�!'$�x��i��I�f��sSџ�����n�<�$�#��j�A�ԬŸ,3�d"�O�T� n�Q�"�	r��Gǐ����O"��Oz�l�
5�)}�ƛ|� ��Z��=ůDv;�h�����'[����9o�֖���Z�,KcZ�%���QBcI�V>A��p?�O>Y.O��іF9o�`��<�z�q��#����������u�4���&��k�J�`%<��A�Þ�	�����O��$)��?�a��+E��se�{�\Y0���&&<a�R�Hۦ��+O�I��~�|bGQ1��,��d��A?��(^��x�Bv� �B��_2H��)�@ ZE0f� 6 _�`����O4=l�L�l�	ޟ�I�*���ҋ��p�i��F ����Ɇ ���m�^~Zw��9��۟$ʓE��E�;EXl��&�ے�����O����O����O��D�|��� [>NI)�@1a���焰e���g�)G�'-���'c�6=���0�(�	�"}a�+_�Vt�!�L�OR��2����%dX6�i�$��ɂ	/tz�	T�`}}���z����DG$7�r��G��dy�O ��%`���䝨C�H�T,��`��'��'��I�M�#���?���?�DH��]<� hfiz���T����'�Nꓝ?i���}�}�7���3�~���1��d�'et�S�m�:p�������L�������'Avr	�9�ҙ�"�g�2����'���'p�'�>�	�9�l�xrBn�M�MK&�8�	��M�1�^����Aܦ��?ͻa���b@Ҋ0�ΝRr"6����?	��?��DZ��M��O����������J`Y"��}�,@��C�/jΒO(��|����?����?y��{\�,A��-���Ճ�d�`�y-O�Tl�;pt(��럼��C�s���6�L�:Κpڴ��t<+ `
�����O~�d9���P#^a��q*�w#N�⁚�)0i���&��5]R8��'7L@%�0�'�Z���@�h���P���\r��A�'r�'�����T����48�~$��m�ޙs�)�6@Ap*Ύ	q�p����D�f}��'���'���ǮO�R�
����]r������Zv�F�����*q��4���窱���e����b�JP�:OR��O���O�$�O��?��7eA24;K�Ɯ�(�0f��8�I�HشAz�-OW������+ƶX˺%��!�F���I>����?ͧl�>�S�4���F�Dr�$ |0�J"'@W[h�ɰ�9�?�G 3���<ͧ�?I���?��
��`a�G�ۗ^��`�H ��?����Z��3-�ݟ��I�8�O��s1��`��Xh�%	?."���OvY�'�2�'�ɧ��'�lX�R�@�Y y����n����6G2��5���i2kRC�I�z�r���Q�l�<[�iK�R��I��ޟ(�	�� �)��`y¨y�D=;3A@6J�ʰ����!ᬼ�eF� ʓ1f�F�$Y}"�'�,u҉ɽ{(�4Q�n|���'��oޤjp�6��lbr��8H�$�~�U��#S���3!k@�f>a$��
hP�kFm�8�>d�`P>� ����x�|s�iE�z,N񡥂�|3 )��柚O�p��	]9&�&X �*�,&Xd��6����2� f�J�h×
P,��Qb*Z�=�L���	;+�-��Fܢ]c`�f*����O������0��� P.�dK@�Fޕ�@�m0�hU	D�#�*�[QU�X�:{�a(C�a��Ô��*E��/q���/M�1Z�B���B�H���1f!r���<�� �W�z�B	@�@Fo1�RԪ9��-�U�?��\iDKq����O����$�>s І6($�CJГ(����p.�?�����K���֟`A	� ���rlK���2��UK�2m���i`r�'�b��0-[�O���O���
(z.%��ą c��(K�+�-U�c�X:��;�	����I�����˗q޼�j�^V��5�Ď��M���`�(ԫ��x��'AR�|ZcJ�	�/ն>#��[���w���b�O���B��O��D�O��q�~������f�։��$�P�:�!��)܉'���'r�'��	!Ȱ�E �
�8���#�;R����@&������ǟl�'����r>�����:-�R��w���2k��>����?YJ>�,Oj�iX�xx���
I'Ǒ'  �h��ʧ>���?�����u�45&>!õ#N�E��dj2�ͫ+[�MrS"Z�M��������1>a�O^���A�bdX�c�1W��X�i���'
�I'jWјH|2���������Ȗ3!��R1
�&��S���'��l;ȟ�i>7�[(Z�l.e�����뺩�ڴ�����T�lZ&����O��I�K~,�5A��,�O#_��I�'��=�M�.O�ё3�)�� �D��6(N�H�Z�`��A+�7�ЍHպ(n��$��˟��S����?i%�E�P��T�у/�$U8�Ξ�`ܛf�O>��	%`�̀s�XmR@��n�.~H���4�?a��?�aoE	[��O`�Ĳ�4X�,� R�D�BC��� �7�I�whb���	�X�	�/LN��Q�� $ŚYB��NjH���ݴ�?�73/+�'�2�'~ɧ56�D:"U;��=h�mz�G�%��O��D�O��D�<i��\Y�3H���[��X�Jqƛx��'0�|��>�ʅ���p���E�5(ɀRBDm��?���?Q+O.�zUB��|�%�R�$	�T����hR�t�")���M�'��|r�'B�G�^n��@�fθ�BeAA="��Z4��	�d��̟Ԕ'00��&�~��f����&ƛdJY�d�\ p!��i���|R�'��hP�/qO�I�@�O��x����l����Ӿi_��'��	�1�ݻ��~��O�����HB��!3>\����4 ��x'�x�I��U.�U������cB.��o���E�뜻�M{(O<	"����������?}ȬOk�*1�� h��+؄��ӧ	(Л6�'�L�!txR�|B��D
U�qe�#W���S(J6Ǜ��J��6��O����Op���U}V��R�G�	��i��=:Q�����M���
%�?J>)����'x�y�"�;��u��A�[%<�z��a�j���O���.h1�'��	�\� �T��SM�%k�p�QӁR/4����>7G���?���?Y�
	�y\���I;z6��W%D5e�&�'G �[�+�>�(O���3���:�{p\��Ř�ȏ�EPB�;�R�t@���ޟ�'?��'(�_�\��O�".�.���'I+;T�њ�)Te t	��OP��?	K>����?���,U|��%b�=}u�huiP�#�&Y�����D�O�D�O����y�:���[���t�zq�����-�$�i��IԟP$���	ԟ��A���Ba��æ�� E�0I&˒N�����O&���O<�[����!V?i�Ɉ+qRs!�r�ny�"��4-+��ߴ�?�M>	��?Ya�M8��'^��"A��!���R!3,�,[�4�?����dL�p/�X�O���'{��J�L��� �ޚ'x `�ɸ*t6O*��O(�ze/��]:T��>%���[��E�e̒Y�ч��Y�'�UjF�z�`X�O���O���(\|Ai�C�Ʀq��dD`�a۴����Ov��[��w�s�N�����NG�j���a���qԴi�,E�Ѓh�D�D�O�$���%��S�F�>��U�Qy��+~r2�
�4%������?i-O�����O�����/{���Kd��|�d�	঩�	��x��B��L<�'�?1�'�ɸ!"�*^иi���7a|	��4�?Y-O�|�ČF��'B��'-2�>8XXL�R/Q'a��Ȃ�K�`@6-�O:IV#QR�i>u��b�i�ո׍@R R�b�)�ڣ΢>1���?H>����d�Oja���΅A�P4��'
<���cAU��ʓ�?�����'s��'�T3��>Y��Q�A�v�ЅcP�\�.�ҁ�yR�'��	ɟ̣e�eb�N��{r�a'O�(n=>d�aNF����ßL�?y��?1D�K�ffYl�-I�TɆ�
�TBJi G�j�TO��D�<A�x	f�*�.�$ �ŀ6A��}|�;D!D+gp�ne���?���w�	��z≞I�}�w�ǜ3� ���ߤkS7��O���?�a��$���O��d�k솉wz�D��O&��}(#��m�''B�'��Ly��+����	�+� =�v�N�B=�c���Ca������͙П�Iӟ4�I�?��u''�/d���Y�X&h
���U��M����?����'=F�L�<�~2c<��}��P$u�z	)ר�٦�Xg��M;��?������x�O��;�V>cܥJ6mΏ0?r��a�lӊ4sR��O��ħ<�J~�'`�A��-F&�C��I;�h�h�v���O���ďF��S�T�>�����YA���i�&��US��Gw1O&Iz�B�c�S���	��5��-Ȱ8E�4{������M��"��e���x�O2�|rgKM��:ą�d����@� h���z�j-J����?).O��ęW�? �TK�d+ư5b.R��`���5��D�On�$?�����ɠ,*��q o�$s\�ax�a!w��ACjΡxHc���Iuy��'�d!�֟4(����%�JX*�@�W�,���i���'��O����O����Y�r5��`\K��1q�� �a�ʱAۃ����O��$�O�2Ul@����Bl���������aW:-��7��O��O���6�p�����LJTA^,L��
$�S/2�|7M�O���<�T*F
x`�O����5FdA	��� .]Q�!2a�������sB�d"�i�?�J�f�,+R�����u���W.s��ʓ O�ݦ�ʬ�R�$�x��'mu�6f�!���"R�N�}�T(j�4�򤞷0,���T[�m�s�rQ��N"3!�$��BC:�pPK�iwfUJ��'"�'[��OZ�)��N a��!�������x��+W��N4��+�y��i�O�13r!؍JiL�iCb&����KԦ���������~���OL˓�?��'s@=��*�,. ̕�S�Ed��H�4��ew���S���'���'&4P��*N�Bu�&�έu�@��n�B�Č:$�t��'9������'8Zc��I�B��H�`L�}���X�Of혀�����ʟ �	��p�'�>P���y/���`J��tH�!�Z�8&����d�Ojʓ�?I��?a#	�/{mj��ǂ��<XBP��rѼD���$�O���OJ�x��i =��9i�x�lA�J*]��T�ļie�I⟤�'d�'�B��7�y��0�ʹ�EC0F�2��>-�$6m�O����Oj���<���MW������*G��5n�"pn�<H�t��Ɠ��M�����O����O��>O<�$����/֙Z��a��=0���k5{�p���O"�y�ꌳ [?e�I������X f�Cb�0��uE��52B��O����O���&K�d�O�ʓ��tO�����J
�!���"$��M)O� �'�֦a��ʟ��I�?UڪO�n�P��V�П=B�u��n�.���'��n�����<���T�?xJN�i fI�^`8#�7�M�냉k�6�'���'�����>q.O��{d@�(fJ�%��16�yh�ȑ�=�AH`�'�$���fSa��U~�v#�Cª[Q2P���iB�'�B�j�2�����Ov�	�H�����77z� 3,�']�6-�O ʓ>���S���'PR�'���5v�J,��I�d���lӴ�d�:/�Ȥ�'���ܕ'Zc�l���s�fX�@Y'3`�A�O����5O��$�OD�D�O��d�<�퀍ao$d��(�;��D�פ���V���'}�R���������,����L�q�N�{` H:")j��7La����������H�INy"N�瓻%!88�s�I��E�Z8��7M�<!����d�O����OrA�e7OPp�r��z�A:�ۓl��]B@������������'�I���~z��C[҅+��^
��3Ċ(Ac,ɫйi$S��	ş��I! ���	a��[�B��Հ�/\H�;�f�����'��U�����R�����O��������T2���ƉE�=���Vb}��'-��'E��O^ʓ���N\��L���Ԑ.?�@s�W��M�,OYP�%Aئm�	�H���?��O�NN(�Z�P��@7D'v��6�R ����'��nG��y2�'�r�'�q�"�`d����UTf��C�i�65x@/`��d�O��D��'���h[z����.	X�Jd��V��*ڴU�Bm�����O��+ �Uе�@6��8i�j,oZş������hq�_3��d�<���~����t��qV�]4=4�I��o �M[��?a��'"&�S���'|��'��E#��� )�����H�H�@Hw�f�$ǌv�.5�'��	֟�'�Zcgj�
m@�	K�pa	#o�l��O��T>O���O���Or��<��a�>�x��CxL�sfgP�644%�q\���'�R�����4�I)���Qs�Й)�\ġ�/�>5�2��a�a���'���'\V��
C5���N��(V>���i_�[N0��J��M�(O ��<����?��z�^͓QF9&DՍvWDqF��}IVY�V�i�B�'��'��I�:�8������cf��S��YE�I��N
�2Ul���x�'S��'��-��y�>�*�7H���
�)�2G�P�G
���	П��'���~���?Q�������^�N�"�Y ^�.x_���I�����Z~#<�O�:X-`��ׄS p�Иp5���M�*O���Q�m��ן��	�?�q�O��=y�ܻu�T�3� ��,�+oq�6�'��H����D�<!���-M)n�(T��fB#TSν�C�M#s�U�<��f�'��'��(�>y-O:q�G�U7�\�č>���Z�ʜΦA�W`��$������uݐ�HV헃5.��z��.7�> "�i�2�'nb���D\Dꓵ���O��I4g�%�M�-W��*@Ǘ�0�(6-�O��[e�I�S��'���'��2��E������d/	`���`(b���d(U�ha�'��ȟ��'�Zc�|���B�${�:a����"�X�X�4�?����<-O:�d�O8�d�<��g[�-E�P6A%"�>���I�s�aeT�0�'�[�4��͟��/}��d�Q(��F�|�ƄO:�B�p�On���'B�'�Z�H�ķ��T�2G`'I[?6A��7���M.O8���<	��?��-���'����Q�_��ۧjJq��1޴�?����?q����Sg��OgZ� ���@�KTM
��Pn�:%����i}�[��������	&5В�I_�ď����	�t�^eD�	أ �?8�&7��O����<	���0�O��O��9�0!Ʃx@��c�)t���;!2���OT��Z�_$��/�d�?y�"�,����.a ��y�nn�&��3v�i���'�?��'T�	�*i���V�ظ,�Xe�#(ɬ7@�6�O��d@�F9�D(��0�*� �P OH>���ʊ'xݢ6���<Rm�꟬�I��T�S4���?�ᎶX.�p�/��Oo �2q�F5\$��ˎ>/|���O<y�FĀ�a#����]��uФJNݦU�	����ɕk�V)��}b�'���)����o�kZ�E���޿V���|"�ڟM�2P�H��Ο��i��
�$O&~$|iUa��Z,!�tӐ�����%�4����'pZc:��I���=��Tɠ��=?
䝈�O�����O���?���?�/OJ+ ���X�k�肻T�&�	��K� "��>�����?����"�!�숄冀p���-lT��$��<�(O���Oz�ģ<�iZ�;��	'�D�DH����#V�2{�������s�����	�s�z�	y�>Y��K�c��S7nO7u�A�O���O��Ĩ<i�.��N|�`叓p$�^�V����.W�Aƛ�'��'��'�`U�'����

pW�e���O.j�]n�̟@�	|y�� �������.���:� �޹e�p!��_�����IE^fm�	F�e�c��	O08�V
�B#�SD����'V�)|�9�Ob�O���k84�
��:b���IZ:��5n�柘��	��M��v�	[�'#�E�P'�.Zsl����bt"-n�=TP� �ݴ�?1��?��'x��O�E@�KH%�ty��!�2��G�	XQ�v��'�����3�F�S�ꅬ�
 Z�m[ +jX�� �i~�'�b��Q�BOT���O��I:y�(��aH�An�K��Įy6m<�$'T�.4$>������9-���0�ؽ+����u�BE쭓ߴ�?�'U�H��O��0���x9*���2*����J�58�l�^��;��C��ԕ'���'�BW�t v$ �8K�DiM.{�0�p o�h �K<����hOx�	�q&�,�c/\�!�ۣ��_�n7�O�˓�?����?!/O�T��K�|����q�hy7�R�x$�}��N}R�'�ў\�'��a	:yHp1rcH�|�顧��:p��?����?y��?�����I�O ���C�*�A���ԨA b�æ���r����'��asK<Qf͆P;�4;"EC�P|\�C�Jզ��I؟l�'adp��-'�I�O�Ʉ�N�̂w��	%z���	�vV�mU�O�6LD����Mk7�D(�,]�����2������֦������	ҟ��	ȟH�I�?i��5&	B2;92|h��b^�Ը����MC���D+���f�-Ȯa�Lє$��m���#o?��a��LM�7M�O����O��p}�_���R�J*p{��`G-�ܥ�퓦�M+�BU�<�I>Q���'��i�J^&F�|k�-�7�x�r#v�����O��$��E[���'��	ڟp��8j����D�"t���p�R2t���oן,�I�t�d�~��?Q��?�B�ʉ?���&zE��eNߛ��'�Hp���>)O���<	������ ��'���a�x5[ w}��;�y��'�r�'���'�剉5*�0� �x��!�BM.ob�����=���<!����$�Op���O&U��	8�$r�L>����M>>��؟��ݟ��Dyr`�l����A?��S��[�}]�!zG[=R�7�<�������O����OL��]�ȣF�F,L�xx�'�c�y�Iy�
���O����O:�����$^?Y�i�%�	���(` B��N��iv�����<����?���0Ӵt���ihj ,Q2[eN��	��f�ܴ�?)���$�7*�8�O���'!�����*͂ �/�JJi,�F$���>����?��e���̓��9O��ӬTKV� 2/�	�~(��dO&Q>�7M�<��Xx�6�'A"�'���d�>�;:5� �E��^�D�1���g�P4oן��	�f��Iȟx��ʟ$�}Z��G�ָ"�fv��"ꦕi�-]��Mk��?I���j�Z���'�Ђ�n�Z��_�{pڠ�bw�D�18O��D�<����'ഀd��f����vJ��J:x�P�~���D�OL�D��2˾�'���ҟ0�xZ�p7i݈���
��#�9o韨�I�<qfDi��'�?���?a���gK꽳�KW(T����wmL>���'����>�+O�d�<����� C���A�45�s	���)����$�I����֟L�O`�ć�ܪ֕�=0(Р��!D���I����I���_�	��R�^)�A�P>Z��=�ElQq���m�˶��?����?),O���	��|*��D�B�2�G1n��%	�jJq}"�']��'R�OJ��f[?��Rg��{Ж�z��ւ-[z�#�k�>����?y���?��<F�<A(�p�$Δ%��qb� >�(d���#�^qmğ�%���IDy��L��ēZ�q���W�+O�� c��&`�>\B&���'��>�I�Ag
9�f�:�%�d�O�b�C�	/r�<C2h	j���Q�KL�E�6�Bp�	2 ���vm���;7��*
k�P���z��!q����m�f\��,� �HӦ投�,�r�ɟg*5�&�)WF�h�����rL�� _f�x�%���,"L(�2?����	�#C6�01���i^�`@����C�h�+\j����͗:KX$p�iR`�b
ť�O��d�O�$Ϻ#DO7/�xH9���e�ҭ{��5u��P�!ʎ4����'U �+��4�0}��@�]Ҭy3@@�t9R��U�c��4ʃ�m�9��#((�};���.��(�v�	�I	`q1Ge
(���7E�$Og�)��[~b���?ͧ�hO�(EE�F|�8�`R�Q#�"O"�HGo�'0Ŏm��"T%z� y���� ���?�'�ƄD˅I�i��'X����A���t�����'kr�'�b{�9��ޟ�ϧNu:]@O̞�|L�
A��0qH�ͅ�#��PHj�,v�a{r��Z�u����Ref]/K�Fe���78�zyS�ڔCa{r�P�4�b�퉚�)P �N�t�"yq��?I���!��t��h��P&�ΰÎM3^�B䉕Q��EB�#�	M��R�o�
p��b� ��O�ʓ@�*IPRU���	�'+��Y'η뎌z�-Ǳ
N���ܟ��e��\�I�|�Յ��hx�pK􏎭4k��_�oՈ�4�X�6	���#ܛ��x���5W��cm�@���"M����(Q���r��1�R���D�[���'��	�{o�@����/l�h�;$.�<v�b���	�B�
h��O�x�,���Q�Z�&B��2�M�j�H�A� g�p}"�%M�<I,OLD���Lw}��'�#`�b��I�~�p���o�u�7f���J��	ߟ@ �N���I���|�*�2�����L��u*6�w��4`�>i���-�^	XæE�Q?��e��P����)���"��:}BJ��?I��h�`��#M�-8�"�
��i0��� YW!�H�KM\]���i��1�V
=g?ax=�V�L7�ƿ�\��� ��N��a]����ԟ��EG��v����	��������y��	al.	��c�l�}cY��L� �4Y������ UN�g�	,R��� 2m��9�C�0b��|�"�9���J��kQ�Z��.�3�Ā�1nĜ����h���0Dh�xPh�*?Q��؟�SX�'Q@Đ+V+��eK�*�'R��	
�'�|��mÒK,�	
eΕ(0��O��Dzʟ4ʓ!�^�´/�]�l"DK�x/����'&T а���?���?ᦷ�t���O���-���"@ɜ5��C��EK6����a��%fԜpP�]� 5�(�W�'�H$HgKon@� ́(��&�qQh|��0�΀�gLN8�X����n�\�4B^	ލ)�@��[Jb�d����`�4��'6Xb?�J#�O10�*Ł��,��M�n'D��qI�$~��P�Y���?��)��Ľ<�w ^�q̛��'�򩚛^��L�EƏ�vB�Y���Q	D�2�'�Ldi��'RR�'�P���JIV7LYzv��r��H�.��-Y��L+z�n�����p<I5Ù�˨af�f>��3� E?&���Q�G�.P�� Zs��7q>���	:=����OV�o���Y4-]�_�(�h��
/f�<����_y��'��O>�Z'�C�dW=��,I�(�y���Rk�����Xo"����U���[#��'L�:(6 �Id�'�ў��R+�}�z�y7Ί0ef1@�@"D��1�NT,#��!9B�X�VnR{�'Ӱiz�.N�A�]C��;`36�z�'Q���FfO�54A��%=+�2p��'iXM�A�5ʎ��"N^���'B)�!M�C5��Í!<�A��'c�}JD�(�eS��֗	�����'\T��)�LR��a�^N���B�'��|�1J��C�½�Ѩ��G!2M��'ÌQ�D��'iB0���H�+h��'�H�Bq���y`�	ăC�v��2�'M��V�X+�ZH�Cb۫ aZh
�'�F<c ̑�)�u��J��,قp(
�'e��㡣H4<�])bfC/A2��	�'@�+q1vH�	F�+t$�	�'��	;6΀�i�2	[�B�18�s	�'P�H���<p���i+ŜWENT		�'�L�P��XH��2d��L�h5��'��d���)��c�
m�9��'����t�E�kzpػ�g�l��!��'��)+�e[BT��C�)�Z�pq�'�P���=D �2�)U�@,q��� �0v�J���C@����"O�ũ�� ��r�_�eoL!x�"O��7.M !��m�b��+ISޑIt"O�t��ڃ^L�FN==Cm�&"O�����ߔ+hHC1n
�|<�1�A"O�M�蓌)�zm�f�;5�PP�"Oz�x�慦j���Wo܎C���ˁ"Obѫ���*7��y�-�;<�p���"Ob���D�z(�h���1�@�k�"O������w��P�Ѹ^
0yA"O�e{҂�7�V�&�Kg`��s�"O@|ZR�D)�r��gԬ^�`�"O�D�@�� 	�ݨ�!"r��}��"O�H4�ڽm��0 Gʚ�KQ"Ovm���+��9+%��(�z�AR"O��'�'Tcl-9D��6��lX�"O|�f�G�P}�pd�ҖAZ*�q4"O�a�E�z,
9+�*
s2�P5"O�8�#��8J0� P�k�����"O�HCr�ʕK�� �D6@*c"O �	U@�&_$�00J',�!��"O��/\����Ԡҝe�����"O��ă\3B�~��gBʘč�$"O�L���ʯ`]Ҥ8��'��q8B"O�1!���2ƌīR�5/�Xp3"O =�f%�ل����!o�pe"O��`ü���B-Ĩc4���y���'m��2b�
>�����:�y��FNJqq�k�7�xlIv�Q��y2��2C�&���V �k�CY�y�I�W�\�ƵE���T�ћ�y�jM�}U�,z�"Q#o�h���*���y�`��y����wY�_�@2����y"A�"��c�ީ'$��dǎ%�y�!J�a��tmT�%ܴA�!��yr"�W-(����!k��2L��yAR ��؊�	(*�~�g���y�I0&���jD��+O��p�+��ybd	�h<�����^V�};ƀ��y��U�+8 ����E4�\Ce�М�y2���%���i�㈁I�AB��yB��#<�|3�&��������y����5y�M���H,
��0`�S��y�1*J���� 0�ț�H�yⅉ��⍃��'���# <�yI߻�ȱa&��2��X�dM��ylߩE�V�k��D�1�L8�Y!�yRm��*�,�q%<,`y�ȃ*�y�BW%����&	�7h�Qq$��y�&�,-c�b#҈d0R������y�DJ7st�#��ПD�<��t�X&kF�Ts���;�g?IC�Ycb�0�Ye[$4�$�t�<��CXm��;7\�&���v ^*9a}�d
�+���mͬtގm�3P��=	g�ٴ9+�X��$2��
�N(+����U��'��}
��["i�j�*��:e*#�ҧM'fP��E��/�Ո����!�"l!���z�<��CDANY���D8	�O[?I��W��h���zeL���b4H�*5>��"OD:i;�� �6(��*��>�%�-��=�%Q�
H��c����Y01��G��,�ca�Ԧ}�&���=ٱ� �2�K�o%D���F٧c�ʹ�t*Ax�� ���;Ka�]z��=?A�&½�~ʟƹ����ӓ�X�aH:�h�N?"����z�<� �4��7���p͛.q�F-	��N!(��Ʌ��$ݘ_�7�����S�D�Z-/ 24:P)W�0�a��J��0=I����v������<7�C�C��17$x�mCq�pл��
D�13cQ��'��'����F�I&ƀ�e�B��ڍy��F�КŁ[����yZw?�T������S�@���Y�'��r���	UA����%2���X��H�<�@Ѭ^;A�yb�HI���8~���|
��@�\�ݰB��K)���0/A�$���t�;\00���8���Q"�	��(�05Y(4�S��.k9 ua����<Q��Z\U�鱐(}ʟ}�PBYB��!A����6Aj�'쀀�eT�]�0�H�'�e���G��Tl��a���<�#CH���ɦF�֟��u������lH�H�IZ�n���zg�U�E����<9�T�A��̓dK�O���6��ڨ-���%��A��i@�cJ�B���@XR��$\O�`޻l��`I�L�rCܘ[��3��V���q7��?��ң�DK@*�ȕ�eNjd�	�Mb��YB��?A!�L�#	!�$�s&B8�v�a��%��!��*�2q�"��o�< S"�G�؂m�D"�"����4$�Dc>�#0$��X8��zkϪIAlJ� 6LOz�5gԦ$	&"�;O\�#��?�.��D�)Y$z|�d�]
p ���
��M3!�\�/Pl�>�O���>S�Ht9�� s)Dٷ��"w!T8�7�K2E�Q>�^�C�xS^nH��Ab@�5`�8-�'P`��(F,�p=)�DZ���a!���@�(ɋ��MX����NJ#A�P���?z�؁K�L�U��[q��d��&��y"L�9����u`���0���!��w��`q��[R��*1���(��d�����7ԙ�!�Y4cK�`��"OH顲`'l<9�@�4���P��.J�Fp!����y�� O���(Į� �!T�q"�[A!\u'���R�"��Ս_K����j>&&��+bӺ�g�I�^ތ�דG�И�����x�"4K�:ʞ)���L�j)y��	֦I����c|�����`���8��,D�`B���8\x�Ra��t�#�(D���PcJ25�ҭ�f(����"D� �B�RBq� *L��9:1$,D�H����r��J�0��Q��*D�(��̙3v�>!�Q�GN�����y�Nڇ�T(u��I���Z�@���yR���4cԙ1���<V� �`����yr��-6u2�+�M��ap���2�yb&X->xU��̞3[�0D��@7�y�ϡR ���G�%B������y�څ�X�C�!�F���B��y��֣*�\Q�#ܷ�L �D���y���8J���f؈Q>%��P�y�Hۍk�H�&�R$��Z�Ȭ�yb�U Y(use�E.[�8	ă�,�y�lعg+�Dc�G���C&e�-�y� T�;h�Z`��3L��l�@+L �y"�¦�b	����J�Dle��~�KI�^v��$�5��y�D�1J'�E��i@(4N�|��ߤ�����_��A��Xб���E�C��$�՚g�ґ^��!Ѡ���r�<)�*� �Q?��R�̞ �����"o�>����)D��"AO2"�a �Tr]Q��H),�a����O�ZvaG9Z�P�A�H)Z���"OV�yG�A�?BlK�D�'&1�$�R��Q�#9�O@ʤ���[��-h��m.�$�'"O�<zP�+�8�Ec� {n0x3"O��J0ː ;���ʉl����"Ox�A�S�(l���gʰ�F�C�Q���V#%�S�O�0}B��H�`�.	���^&]�e�'��P�![�M7��
�"�2IU��O>IV"�0�0=���`��Ԑ�M�,fdpf�	_�����L��I�E�sn�z���s�m��G��e�uNGQnez)M	4��F	�;e>Őc-ӧ8eR�[�$��7u�����1D����٠��)ԥ���T���B�<��Q����(�� 2P���هV�yp����:�pIV"Oba��$'���0��K�2�p%ȡ�|�J�6�az2�t��<��8��h]8�p>�cJ�q頬���w� `��7\�T2aO�C�bB�	/F�Q@A�Sb� 1�,̳$�<��B-B�#~2"��7����ѡē�z�B�c�^�<95�C�14fU�F�H*!�E�ѵS;(�[�cWG�S��?�B$؀*K� 3 ��RQ|���
�K�<�%��<�zx���n[���̌q?U�ZK�`��$،n����
B�1$FP���~Y�|�A���E�w�@�jc�3R]������g�z`��!��!����s/�%pfD�v�Dy�`%��F�D�۞��U˒�$�U�3��8�y��1#�x�ʰ(�}E��l��h��9s��F������R&Rb ��QG�yL������y�����\����u��y��L��~bʌV8���1&�xcŁ?������Y�l���$�>�(͓\�n�҆��5$ʹAӑ
V�-�f��HJѬ])wp@�4�o���ȓxP.��g+`7�)[W��2�|��oU�q��d�.>t8�5ߡT\�x�ȓ��[�eœ����s�ܨYY� ���Dp2��
mk��$æ!�ȓpEVݺ��#A�����lw|�ȓV��e�� ����S��l=�3"O�����4$#���֜P��1p�"O2-��,E�7g�!����/l�H�) "O�`yƉ֦}��d�5�V)Ku"O�%�Uҩ7j�!�T
�Si9t"O��$!�'<�aˠE�*PT�V"O�!J�!/�Xp��]T�@H�"O�5Ru���/G������,P$��"O��'HF�F��pí�?(� <0"O�}��������3f��4�*\`Q"O��z���r�l{���),䶆"O��
0��$.�V����ε4z���"O4�I����m�t�Y�-�+I%ش"O@�:�B�2e8����Ŀ;���	"OJ�wN�#�d�j�+���}�"O2�Ė�p9���Q�b����"O�-� ] %�.�x�	V7U��Yx�"O�p�!��x�e�1�Em���u"O�Q !��<L�"
�*�.��$"O�\j��
��h:�������"OV� T��^���A��2�h"O����J+ӈhH�V/l���"O���B�u>�y�ȥeԆh�&"OLĹ��a~l�bJ¹<�<5�"O(dj�A1:�4���^�^��"O���"�V)+Gp��l�;_ʶɘ�"O�)����p���2�X�QƝS"Ov�H�A�^�a�ơ Ej�e�"O��1��ާUf�Ҥ�S�W A�$"O
�!�.HN��K҅Y悕�"O0](��؄%�@j�+ؙ�ҐHv"O����(M482H����H�n�  "O>d+cA�&9D�vO�>��E)F"Odx�d$�
a�F��.C"��"O�8�Q�r�n�#7K F�PKf"OB@�BPep���k3Q֐���"O�$����|�H�y�ʐ�St��s"O�s1a;��Yc Ģ6j���f"Ob�*cŞ�C��I�d\\��x�"Ot<�A Tk��t�F��UX��,�y
� h�YW搷[|�%k���1�"O���v�G�y �m��j������"O�� �%Q_��9sO�$p{paie"O��@�˟�8�&PY�6
��ۡ"O��(!&٥|X�ɢPjŜ/��$	�"OH��s��ѹ�^~�`��"Or|
���>2謹0h�{	��0T"O��*E$(j`���W�*(�"O�r4n�7���Y�
�%��s#"O2%�b�͌H�F|�VJʦ{
ڰ�"Of����;Z���f\�^� 8�"O6� �D�"��@�\:�N$0�"O,@#0�J-vg�:3KE�p����$,\O�9�Рӳ(�J�*R
JWZ�[0"O�a9�n�	=�F����]�&;
x3"O��ktn/>���۱��--5D��"O����Z� Q��Z�l�0# �h��"ORة��%2Ơ�aj̜��a"O��rD��,��Y�W�n�0f"O9xt#Ɉ3ha�.Ҭ�w"Ob��QGI�6�^\�@.�fEP'"O�0S� �M�p��`��Q�x�"O�djֆ@�(�l  Qn�G����"OR�� �_?Ӗh���D*Y:|�"O�jW�C�E����,P�X@B�"O(yT��Y&�𰠋�n�n1QB"O�y��O/]t6���l���� 5"Ox�5�� g�Dʐ�ǡ{��i*�"ODd�vl.R�����k҄�6aX�"O�)�f��D�X����mb���"O0�K�f\唰���EpO���u"O4<�@$Z%���ZЈ�`�
5��"O�x3�)��H�0Y�FH�I���"O&Tz�B
_����Bvv(��|��'lfA��<^��.�0*�Q0�'y���a�ۇ$;�	��J�*n���'=Z��F�ܰ/q�C#D?�0�
�'D�dső&�|5#M֖Q�=�	�'=\ĪfL�zz�a�cQ�b�N)�
�'���8��8�Ux6��D�$�8�'_����%�$ c�EEL���'����4V�8�^��Q��!4�|��'�l+�q�l�� hk�X���M���R�Yc�j  �F�Z���"O�ЕB-x� �r�O=C�:���"O��ʄ�S�,�����#��{#"O<��6�K*I)�s�B�Q�J���"O*�s��c�$q���G�C9��h�"O���)Ǿ�P< ��+��<�F"O�<��$�z���I��9/���1�"O��ip��_,���S�\��"O,)E�ݢ��Q�ńПR��B"O@�V&
�nyK���kh����"O|L�c.���x��ā�u+\��"O�8�Ƈ�;^��@�\}���w"O�)ǥV  ���F,��8�S"ObQ���mXצH\{D��q"O��K��$x<J����Wy�0`�"O�E��e�?|�̢7oԣ����"Ori���\�|�*k���t).�h�"O Qsao��\R�Q0"�Y�$��cV"Otɘ%`�5Vd0��b+T
[�I �P�\G{��)X,n@J�[6��Z�D!3U�,�!�$D,<K�Jw	��Ll��	$���%�!�� �����ô^�dL��[�V�zC"O����J3%క
TnU#��u��"O�Ӣ�L"�t���b���	�"Or0!2�� Bb �5-��fo�YJA"O��9�
���(��˒WV¤J�"Ol�`��ˁ�:  %��.8B\Z�"O���Wώ4+,�1��zĴ)9�"O6�N�?x��(C��P;L��l��"OP̪��H]��K��ͨ�E"O���!����Q�&ZbD��A"O��)�鈳0��D�BA�W�H�!"O�*$N2c���@�ɛf�<��r"O\�Fn�V��LS���!n岗"O`i;Uc��jx��ǧ�� v��"Olu����S������Ȣi�T��"O��Z�Ɛw[�ĳB�9d�u�U"Oy;fL�nd�8Ea� .����"O���t�߈Z갡��	~E�%�0�'m�dE�P
���Ѫv��`�DCR�O�!�D��M."�K���Dꊬ����,C!�d�7j:�jd��=�3.**!���Nb"ܒ�j�'d�!
����!#!���#M��sa��~J�P@X�7!򤋁py���"�/A-&y8į�4!�%@�b��'T���y-!�$������q4r��3B�!�D*9�rq�
��} �����<u�!�$�����h�6���5'��!��A����쎴D�詆���!�dD]�XԢ�NR���F�V5E!�sy؅�S���\���5��s�!�'Y+��"�$݉D�T�dL�n�!�$P�x�A$G �
G�)�G�2- !�DUq$��$��&��i��� s�!����]B ��-����B;U!�DڡA�Ƹ3Ge�L���B��%7!�$��G�,]��C�%j���LDG.!�D%2T�X�j��\�I��Ȥb�!��4�`��
G�#V����ݹ�!�P��
���F
A.��p�M�y!�_5�j�˲�
�%&#�o��$ !��Ck�Ꝼ�NY#qR�T�!��صL�T��3#G�ETj8�0�x�!�7�j �""�"E��p3*Y�t�!�$��,�P%4}��mjd	E�a�!�DE7R��yX�D��p��p��'�!�K0��a��δg�l�s��PrU!���W�(��B D�X�&j��Z$K!�D�4h� �o�<&p�UQ&R�F2!��3�  d#�%�����Gu,!�d�X�ڝ��a .�d��$+!��Ȼ9�T�`��5c6�}#�=E%!��ψe=`ڵf�)C4]Y`J& !�	�"C�`��,j����t�7}!�!wL(I�N�U|"�����kc!�^�G����B� ev���	F!�DZD�$���pp4��&#�!�䀓K"���l%=�4�jI�V%!��[�6O�`i��� H�b��w�!���&��`yrm��J!�$�7�p����3���lMqJ!������ �[�Z��	ِK�j5!��Q61��(W�@�>��j�F�!��t��5+��Y|�l����~t!�� �)qhM$	7񀅫Ҥ���r�"O���r�S4j%���I��c�`�r"O�}�fc?6�z|YF��Xl���"O����ā7<?T��Ei�y�J��yR�W.7YP��Wn�{��� r"ˉ�y�G��&�~�{��� �:�[!	Bs�<�3�B�
��ܫaHM8ـL��[U�'Ta�t��(K����=5�� 0p���y�합m"�uQ���*��1�l���y��;sth�BS75���M� �yrN)����D���L��4�y���2����-���3v�Q��y�候%�����ɼVn�A+��0��-�O~ + e�% ��b��]!�"OИ�G�:�`q�a�Ɋ7��%"O�ZG�ҭO�0m�0�ߒb넉���IwX��I���;d2	0��Y�-C���3�>D��J��<�r`�2iY:;���Ã!1D�P�S���-�0��p��vAx���a.D�����/�����3ih!��C+D���fA�$w�.��$cյQҀ@h�h$D����D�/!�g./2>R�)/$D�|����_��M)Ư��`u:��$D�X�H�5p��r��M-0
x1���!D�4�3d�Tň�����<���M>D������ 
���hi(:� �<D����B�"�*Dc��ǾR4U��m5D�4z��'t2�J7!nz�s�,2D��sAeʰ;��P��V+s�D��.D��K�U5[@ (,���z�-D�8��A��6��J�5�(PW.D��#uȳI^�A�.�{��\���(D��rӠ^�w�J�y��جWV��3�9D�T���.���+����XpE��B*D� �ʗ�B��[�)]:|5
%[Wg)D�D�_=T�(�s���٠%3D�<�G�ل%צʕiC1;$��	�+D��n�!vM\� ��kɆ���7D�H��MBxU����>?�2�`7D��Q���+8�)R��l�n��"D�����2<)�WnO`��d !D�p)Р΋��hF�|YX�?D�@��D^,�����B�1��+D� ��휪)�<q+w$Υ_�,1A�i?D�XY���� K4c��8�8�7D����
G���`��.��s����3D�,�E�8sO�|�6!S��l鳇&D��0���)<���`��f�t��R�8D�(��Ä\d�
X*B��0���1D�@��f��<�L�J O�zXk�/D�<�š��}��`�S�͛B�tls��.D�pC��v)��&�>n�Zhc#'7D�����//���-�8��C��3D��� ���C8�l����[�����&T��p�H�3�:{&֔X��)��"O�,��BF23�ZX�B ّ\���	�"O�����,/���a��(�� Q"O\��i�
��y���.�F�:"O�@P�E�[il)��'3Fkf���"OR�:u�]�)�y4hG�TK�d��"O�i�5%�!p� :s���:���s"O41�` �5�:���O`Y��)�"Oر����;l�����^�)ߊ`�"O�Q�g��iҌ53�DռGh���"O�  �#�N2)���cO�co�d{"O�7�K.�;��
.Q|T��"O�����;l<H04`��#{0�s�"O��i���4�x�1�� ^r`m "O�l����4�>�D�F8\e���"O��[Q��J/�]x����>*�$9"O��Ò�Ƈ�Xic��yq�|�s"O�D���@�Ф�p�=M�\le"O�AC���)6N�����$Ja"O@L�a��0��  �� �LiC�"O�T�'�=j��� �a�+T٤�p7"O��cUG�3a_��1N� Mm�Бc"O4�2�΍�-�\�"�_�xXx�21"O:� �J�~��w���x;D�� "Oj��&�p2��aR��1)^aS"O.Q��/Q���A�D�-N�Ҁ��"Ol)�� !�`]+�HAה�B"O,��d��H��)8�C5.��"O�|(Q T�z�Zm�^�[Ղh:�"O.��#���"y+�Μ3u����S"O`��RlV�������X$�"O�*�K.m�y!������"O�M����54((��.�L��yJG"O �y��ݽ����֮�g�&�P"O�x1#�?j���u5�� [�"O�%�v�:/�9z�"��1R�"O�<:�	5?U8�P1�:�!��"O�Q#�%=
,�Q��(|����"O����Q�@<"E�F�5�����"O.1�U瑁��p��eid܁�"O0!z�C�;�����خ	VޑA"O�Y��Z'���#`��'��T	"Or�a��[�FjZ9�r���\�{�"O��[u,X7?dDtcq��H����Q"OL�Z4��	� ��p�@!�����"OVē �Yh,��
��8kC"O�|H����L>���$J�n���"O�t���)9}(��Rr�� �"O���kZJf�@� ;M��D0"O΀�G��n3�pk�K�I�hX�"O�9R�M+{v���XEC$aC�"O~x��ޯ1�&��4�	;+V�I`�"O�B��X��铱��!M�n�:a"Oj�`�CH5w��p�+�g�r@)C"O<�"i�3�-!#�)ʶ���q"Ox%��H�c�$Q�C'�!C�4b1"O�9x�d��7-v�a��<�,=�"OR�3�a.������#tD���"O���Dƀ{�� P ��;n�A��"O����
��KM����kʁ�y2J�?LJTp�O��t�TX�e��y�jI�P�p���	l]���!��(�yB��9PpjXE�Ҿ\;�+��y��ޱ!�E� ���~�*��ɐ��y⡙� Ҏ��Ì�e�z�"����y�%�jx8a�ʟL�`D:F�+�yr� #.y�bK�>�� ���y�G>i�l�D��v^-�w'A��y,[�X�6 �#��*f 	����y�n�e��������,�����	�y��<�rIR�#�80� �&��/�yB�׻pb,���"�D�(	+�y"O�!o��Q��m�(�~D҄
]&�y�)_A��5���ݯ
c�9%�U4�y
� �)����08��+��ւ/�|@�"O:x��-�.(�}�#�L-)t�"Ox��o߶�|H9mũ)�P���"O�P�#	�B�ܰj�+٫nʮ���"Ox��l�NG��qM]!%�2��"Ou��C&��R��Ƴwgz�Ӓ"O,��*�B�\ ����&TcЁ��"O:�@��9*x�4q*�*j�T�� "O��`qDF�{z������5��h��"O�E���]�^T {Vnݰ�F�@"O�0��Z�E)���2M��W��|�"O��b	-�,i8�Ič/��"O,2w�H!"ǖ ��)*��"O���!��"�F��	�h��� �"O���n�d�2�C��5!�*��"O�\���B����["�X� %"O�jW
A�q����"_a����d"O�,K��y�� �ЫD���s"OH�g%�%#z�œ��U���}R"Oz�HN"qI6 ��f�-u� �ȱ"ON��1[�SNa���8ozR4��"O��Adj�� f舁�؜NL�a20"O0�2�ѓum�d�H��:`����"O �@e-��2���b���n~�:"OT�zF�1_�R�TK>5a�ɢ�"O��Z� ]R���j2h2OV��r"OH(����/՚�;�l�CH&	р"O�)�"�ӨA��-r%S'!>�	�"OԜ!�N_Z�4W�I,5���"O���i�$6�^qҕ�H��.�"O��KR#ׯ&$�O2k3�"O(��mI*Z�C2n�6S�t�@"Ot�zR�I�	���v.���3�"O칋�f׈f)S!-�,r��Ӕ"O��ф��)f�����TXi.���"O>l��6}�����d��@�ʇ"O����D�)Q8uy�aC�h�6��"O�L!�NF�T8.܀d���`�'�.�ˡ B3��%��!�!{�@���'�v�(��8p.�*�dؾ����'|^�aRI��ZLT�&�Q04�`�1�'�
XA�/���P�G�"0����'ǲXۅ�Z"=���0��QJZ�h�'��͒���p��9b�U=�Z���'_X��`�@v�9T���U��'�Ę#CCW�����"�M��'v�Aq��]�f}�T/��|1����'��i�b��x-���Dd�_���'g>�:l���P��̜L����
�'��D�$��- �Lu����(F?lH�'ъ�0%E�*]����.F7��Ur�'�PR�D��>`�!��X�$q�'�Fu*nѱ�����2O�R��'���ӗn�e����]$J*�(�'zP��Û�R,JQkG��9W� 	9	�'.�}�W�54��IR"BH�1�'&B�KT?�A3�h;>��q	�'x����mƈ��H����3�p��'�:Q��MΈ9@�0u�� '�I�,Of���L�A�JD	�l�X�Yp��
�!��D��fͰ��ظwD�Qg��tq!���f��4(Q�	1T�
�@'!��H�s�j������$���;E�!�U�Y�&�D-f༭#�����!�O� �)�s�[�-���x���cD"OxuJ��]�#��4��Gӈ$��i�Z�P��N��X�lؖ%�@ɢ&�5]-𴀅c�<q��0>A�FM�NT��ӻ�H���^�<qB��3�����h
�3Z�僗$�O�<���*	0�d�W�E�	��$�H�<���Z|�M��"Ǆ{��CL�jyb�'�0�P�J͚q���9h�a�����'�*�b GU�#�D%���6a�4`K>i���(�I�P���C(�&�,%�~��ʓ�0?9����A^�;�RE��V�<�0O�/_^���7n¤])B��M�<-,�X��h^ �����Q�Մ�5�h����=!rmٌ`rx�'ja~2� ;(�x����&��zT�P���<�����'�tIK[qSR�B띃?@�Њ�'��H��cP�{餑"���	3�X���'���{��I�]ٺ<r�M
�
�'�������%P�yHIʞ���'p����Ξ9-:� Q�?{�(���'�h�$"����E�m�h��'~�	@mג#z�x�v�Jl�<DA	��'�kՃΊ|�\��O�mʩ	�'�q	��J��\K׋�5bHQ�'80�1ӥJ�^�h�[���X���P
�'E:=B�����s����B)t���r����E_T���dΞd!Z��ȓs,�8�w�G+�p���F�����7s�� ���:2+�!хͭb���ȓg���1��7! Mկ)n����ȓ�vtJfh�}8�d�d��(#�=��b�N�qu�֡;��Y@��
ȴ��ȓd�����/Ղ�~)�"��Zh��ȓ��;&��c�x3�@QC ���Dg8��2�KW��[Rn, ����ȓ�,i����,!2EN��%��KԖ!w�ǲ|%���'m
t��ȓO��y`a��RF�4Q��:���ȓ?!LtCU �j�eBI�fz����N�H�Å���g6!�� ?M����ft��Ca�$��E;<h����
l�q��������R�2Rh��4�t��A�.H'L�Sd��>����ᄠY���H���CD���>��D{r��o\�0ƥeu��Q L�f�X4�ȓP)�aqE�[��e��/B��h��{����	�EO�a�*[ p��J�n�B1��+2�l�u��%
	�����r��9" ��P�M�Y"���>���P.�=}Xf��sl�-��@��e��[v�W/<g.�p���j�$��{,��X�	��qojt� />�ԓ��x��W���g�2��c�,�>�y�G��2�1��׃|4e�M��y@�=ezn�A�,��x�-F��y҄ǯqk�l#wa��&`���Ć�yb�۶ T��p#ٙ�VE`��O���6�S�O1�a��މ8Ӽ����`f�D��'̺X�6LL�z�
�#�l��ZѠ5+�'0�� ��{>���C0Z�4i8�'M�����\����ri��Q;�H�
�'��`�,.A��e�R ��Y�H���'�,���#� �.��
Kh��'@��+0g�Mϒ��0d��o�<�x��� ������5�>�ڠ��C�P�y2"O�mi2�������To�N��P"OP �� �>
��A(vډb=�(�"O��A��6�Utl�p�
]� S�<�L�B����ːp FKAM�<	�L��4�C���i��(��KM�<Y��"p�L�'͘�$l���CS~�'�a��!����H�f�"���A�Ș�y��y��A3� �({�h��Wmƍ�yB����@�I�m��)�'���y"eۄT=��{"�B;drl�iW��Py*S�՞C�
/)6��2�m�<A4�#$�H��M�)n�F�:R%j�<��,L�!�Vt�#)�;�����d��hO�'n
5�f�R���a���0R��� |��y2n��X�<�1��$����z���Z=D^��4"�S�m9WD#D��ivŗ4�&�{pÇ�.�T��!D���q��#,�܈R���1��<:�	%D����7|�i��<=���C6D���$	�c���j�E�:=e�1b��2D������rH:���#��m�h$�O���-UV���HZ\G�$	v�O������s��$��!�2�1s��`C!�D%`%:��",�j�>�S�.Z1!�@�QF���.�]�|�8��T'!�=��c��6�\��D��]�!��+M"�점kܥD�n��� TY !�ֲ'�dh�MZ���G��B��ӭs��M
�9(a�&ܞ~�Hʓ�0?�2L��M�.��bAG{FL]{���D�<���""^q�1�^�j�[�fk�<�� ���4\rB㟋tRX��A�m�<���������Ѓ3Ԭ�5��U�<�ѭ�%MF,�A+�8+f{�<92͆�U��Ȓ;�B�R��M�<I�+�&$8�q��䐌q��0	G�<6�[�Dު��0����q��ȓ@�<YW
J�{�,!��ΠW� ����<q$l�U�uAt쐙d��W
�}�<Iҍ��on���3u�aY�GD�<	�Ɲ==8��0�L�8$��F�GX��4�Iq~�l,��b�%�����?�yB&��2P��3�S�h?���P�yB���3T�mxGWv��31��yJJ�`�T�X�`?i��R��	�yBh(O�IT	ޠQCvQ��"�=�y"!ߣ!@�$Lƕ:��<����y�B_�IbJ�9��A���=�yr L�L>D���
Ֆ$L�� �=�y�U�R{�]CjW,�j Z�c���y���+)�0��2��@��V- �y�A�/���+e޷Z^�e��Ɲ$�y�#���%a"�Xj��ɻp��)�y2	�uh����fD_˦i 0h���x"(;���]$J���H�n_�q�!�d�}�dlSeό�l�HirMиT�!� ;7��r�Y02����tm��_!��U?ϔ�#�H�V�@��%��wZ!�� 0p�r��&��)e�^���I�?!�D��$d��A�)�6��D��dO!��A;B�'���ӊ�6=!��̻Z��T�7�ُclH8B�K�NJ!�$�Y ٵ-o��4��T9!�� DIB���R�z)
��Ǐ}��Z"O�m��� �bXa�KkH;�"O�h%��M�j|p�N�-T��C"O�����0#"�@�c�]�����"O�X�$.,$y�Ƣ:x�t��B"Op6��V�\��O�h�R [U"O�hC�?F״D�6��6�8 S"Ov���E�F��铥(y��U�"O<m!���j�-rS��	<�(Y*"O*�!�D�Gb\c1�%k�b%!"O*���C%B&�Trq���q���"O���E��=+�!t��25��R"O�xٕ	S�cX�a� oV�q=�"O$S�$I	Xqr)0ahM�y��c�"OrrM�VA�4�v��2����b"Op�h�%����8�̡�N��y+̪�&lA�/ )L�%k���yR,E�Mn�Ap5�,����n�*�yro�� ���B�O2[�䣴�
��y���H` %��l`� :�$B/�y�Y�>caj��]гg΅��d7�O�y�D��{Hj� %#�wc��xV"O~�Ѱ�
?�m�⋓)�֜��"O����AŌ��4��=�p�ID"O\ ;�Ԕ2mX��¨��=~�ܛ"O��ϑ�&���R��By�ږ"O\����;$����kG�fR2)b�O�����@x���:(�ҁ��ù<����&�I�{�^�ad��e���"�C�'4$B�	�/NBh�!�7N;T(�%'i2C�	�8�zY��
�H�+3F��2�\C�)��L��I�N�>p�(^Ex�C�I+#��9�G'��?L\q�M��bC��@�����͉�(��^�2sFC�I�
��P�Z(Y]�d��E\�6�����bx�h�<���fYH���+҂�f�
3��z�<�M��-K�qJ ��"�
�Ԩ�K�<����@� m�Q�,��xф H�<�@ŎV�$qej#Y�X���E�<QS
"s���3�DR�
�u�p�TC��( � ��%퟊^�Tйa�,c2�C�I�Z�����JK��m�/%��C䉮k�y06k�.E��Q��+�7%)�C䉧]%�<٦,î��� �iߏwq6C�I�I`�i$�ԭs��M�A�[�C�	�� x�s����J�IV�L�C��,U��)tcY�@q
��Â�6 �B�I�nB�(���6o;	��F�1Q��C�9��1���|�i�!��c��D-�Iu��~��mV<�8Vn��8��b��5��d(�Ox��Rf��Ys.`#է�4G�%�"O@4��oX@�=�t&�"fR<  "O~�[NU-p�ְj���>�<�"O�ձ�/N>vivEBD��`�%"OV� d��2�Y	2�K=�~42v"O*�ye�)pS��P ��

ޡp���Z���D�3W�%ZD���Q+�
?D����U8x���i�=�;!�=D���ȺI��p�D�`�0�$%:D�����E#31���ũ�6C�����2D�����T^vvP+V甓\�$���*D�����3Q1Q{��R�TZ�I,D�x�1g��Z��(i��U��ړ�,D�ؚ��	�:ka�R*�462=PC'%D�� �5�áG�*#��ڳ��W2dQ�v"OV����J�|���ۧaƶ7�E��"Ohq��/�4[���p��	'���"O4y.��f��[��߫}����"O�����&�>mI�ݷx�D�Y�"O�!�@�
(�j�!�̀
y�H�[A"Oʁ��Ya�||��m���|���"LOVK��B�v��,߮K�H�ie"O�ȴ�ںȥ�IV�$Y�!�-�y�	Z�l��Թ�-L�E��	9����y���@Sf�\�3Ѷ �&k��y�e�:f�^QS�ء+�����)�y�͇;|P��`h��!�4��f��?��'\r�R%쉺'�X]�bB�@T���
�'k<��6�Ӧ)2h���U�1����'���B*����9QlP#�ۦ�y"�P �T���b��A��aP�ٗ�y��I&�����ِL��AIǋ�yR�ѵ]�б�t#�@�~�BWg���y�� 3�T����+{Θ9����>��O�x ���G�� JI�{e "O�i�#O�>!Vn��	," �ц"O�5�CJ��GϤ�&��
��V"O����Ul��D(aȎ
�|,d�'��Cu>�4�$�N��F�ɻl��� �~�Z�%XM�@�I�&�Bq�ȓK�v�G��LZ�h��ݰ8���ȓSҶP�Ƌ�i�Za�D���"\��:P�ۂ(!T�j�d
m��h��gT���W�P;'��`��	�Ec���ȓ#,�ɢ�։`�rq�h ���I�t�]<�d%�␐?�"�J�r�<���"50�[8\px�ڇ�]l����<a��{��Y!	@4L�Gl�<��5:檝�'�0	n��Qp�<a�*݇hD>��Ʊq��U��-���y�4Y�0�TXE��PĎ8�y��ՅI�T����clE8u ���y���Z��U�ʋF��jDc���y�g@&MQ��"�/��D�8m�s��y��R5�����E��;�QѢ��	�y�`��!z�iS�k �V�IRjN&�y"�S�T�+���S�>�i�!ս�y"�l��%�A�D��+��Y��y��sq6M$��6,�\|)1���y�/�l"B}A�,� ���w�
6��'�ў�OP�Ds�+� <Ƅ@t �$0���'�>���&9)ְ�K �#j�0�',��0�J(ѐ�B�Ԯ)��C
�'����SJ�{�x�¢�S5ޅ�	�'v��ł[4vXɢ$G��R@�'fj�AA��E�`I�B�H&hmS�'�h�*e�T��)`�0}��q�|�U������ �j�
dĹ�RȎ�\q C�	�W"���O�J�أ�ά=�JB�I'f�$T�q� -�jM�RiL�&$B�	"WAʔ8��
f�R�b�"
�!qB�	BC,X��@�#�"������ C�I	_z�4s�P��FdA��\h<yUA���=97�!u��R��K�<9�'�;x]17aEgߌ�4M}�<!W�I��n���Լx��@����c�<���^�;p9`��:��˅�Sa�<9�KH��j�[�I( �H����	a�<� ��)��\�;}��
S�@О,�"O>�ء�܆6��|	�HZ�3��a"O�4[Ү�:�a`d�Jx:B"O=��M�&=xJ��Ԝy�"O��c��O�r�6P��0}>}+���p�O��)�V��e�Hõ�U�M
(�	�'� �:��T#G�-�a�,��<��'d��{�$
-C{�	�M	3(g�W�<�R�Z�(�6]�)�8	CrȰ�,�i��@�<��S;7%�	6�J�4<`�ȃ_M�<	�C�t<�X��דzа���H�<iu�G�\�!a�l��\�0 ��
B�<�p��*ĸ
�.U88�P ��}�<g+���[�C3;t��[Gɕn�<�7F\�My����ְp���BO�<�V�>f¬�M�2m�0��
I�<��R5�>�I��\4=4�)�e�Zn�<I`�]�3)0�!ФM<�
�g�<���J�,(���f��P�%_�<1���=[����}L��e�47O!�!�"�hI '��è]7@!�@-L,MR4`�5#Z<�AI��!�D�z��f$9���$�X�_g!�W%r�;�'D�l��b,�T=!��;9F�-��+ESL~t�2H�I)ў�����ahh��d?Juq+�6B�I�Y�<XA3���I�!0� �*i<lC䉵*P4�lK';���FV�2'rB�>B�D���	(^�] ��/B-TB�I�J���C��*a�|E)ь�sA,B�	p���bG�X�"
Y��M�5"OLT1�kJ���]r�&�~q�B�"O^X!$H�lAZ���ڡ t�ъ�"Or�I$��."�Hqp��M#s��`�"O��;q�[t ���yQāHv"O2��VG�yL.%X��%IZ&Żq"ON� )����"��,��s�'>��f��@HG�[�	�"���$�/[nB��/X�҉ �,�QTA��i�O B剡�`�&��	�Z��gَ4�!�$��YL��	�*ӆ���;�gU%�!�DC�e�!C�@�8Y1V�˕��	X�!�7��1���9 �A��b!!��k����[
\���"�;f�}����P�e�8b���!��[�G�:��Ԅ!D�X �睁I,�bS`�*$7� �� =D�#vh�lܺ��B#��S9֜���<D�h���$��,Yc��$C����" D����.THD�hW ҂�0e��� D��q�f�8��9e��'w�Ε��;D�8��d�J�Fr �������.D�|���2E^�����5]|t��-,D��9f,ԑa玅Y�M\=vb��c7D�T2��;6�$MJ�Ě��R-��5D����L
e���S`W��
�f.D����Ҙ� �Y/`�ċǄ-D����ݯI�llic�V�^˼�i�)-D�t�TDL�������!Y�|�!D���(ȩ z8�A�iNpt��4D�\��L�-5ĪMC�߿�>����$D�(���/x���7N�,Q�ލ�BJ!D�`���)!$Q���M�Yw�	��>D���d�U:cY4TKSh�d�i��n<D��2ТԖWZP�2&���F����0D�� L%�p�C8;��)���F��q""O$ !j�<���mY�8��$��T� �'�ў�OH��[��׷~:��愔Y�IS	�'�4�`c�D�d��&��$La4ȫ�'��S�c�w\�B��_�q��((	�'˒m���տV��	�eLK�g����xgU���̙`/�Q�BY�V�� �y��t�!H�c�"����	��y��qp�4
��"ȂHau��y�X><h6�PנF#d؜��(�y��R{�YYaA� h,e�Ǐ��y��Q�� ����o�43�+���'�ў�ON"1H8M���h9+�v�2	�'_�� �C&��a��"4HN�j�'k���@��<�U���(�N�)���*�u�dsV#,p��*�"Oq>.I�ȓ!�1���TD�1�A���T��X�\թpgƹ+��`#R&ca�Ԅ�2��X '�F��R�#H�-��q�͚�57�*�0& H� R`q�ȓls�cN�֞A�"�R��ȓ-E:��m��Y�I�~����Z�'�C�ɬTz��a��S()�����'ޝK׎M�K�I�QZ�U���'=�9S��4�r�j�Aa����'c."�#$c�$��a��Q2��	�'�j��.Q��Y+���?Q*��
�'�h��Lc~i�ș#D��	�'RȈ�B�w����k��-*	�'�d9%��L��v�F�Y���y���d=�Sܧq��P�]�.�KW��(?
!�ȓ?Ĥ��dǊ�*�^ �Guh��kD,�R`�:q�@��`a0D�	!#�&f�r� �  ք�S!�)D�`b)�P;rx�S^�L�H5N;D�ph�*ы~;��b�N�ERL�rDk:ړ��$5§�lYa�ǝ�بAF�� bd��ӟ�����U�\-m�U�~�T��`��b@B�I�s�H0A��n�P��A�VB䉔X_����6Y~=�uG�A�fB�	�%�~�����v�LA�f�Y�,B�I.7�n%�V��WN�a��։�C�3�8KcKσ.�&���������&?�R (�\�	$N7Fp]G{��'��hT�^����:��<gq�']�`��
�36�|5�S�׾c؄���'L�M⳧�y0|��K�W���s�'���E6D1�VKW�K<S	�'����ּkm����-WUȝ�	�'�Z���JE�Wъz�
�`�����'>�uPp�Фs��ԩEH�����'����!u5�����qh�Q��'�ܼ�@�2H�@e�c�ĉ��'i:�*5M�����Ɗ/F�|��'��2w�Ģ'���*pŚu��	�
�'��,���כas,AЧ@̬D����
�'�Й�%�G�j�b-�WF�C:����@���^&P�\E�@�H7Gm>|�ȓ&��P5EȩO��\H�����T�ȓ܄i�dM.s��x���/;�~�ȓ�3��w��DҰG
�,�Pe�ȓ ��N7z$²�Q�,,�t��(�|�p��s˖@��ė�#X�ȓ:��&�A��p�{�n��%Y�ل�S�? R����lv&,��+�"�0a�|b�)�� mK��c��L$�q��+��B�ɨE��k� ^�'� �i%I�)��B�ɠ%� 8c!ˑ�M��)c.�J|�B�I5*�V�QQ1d��D�P��;��B䉍�0���S�h�)�b���B䉬V��`8bo�`[�I���ݗD%�B��8*�Fh2"��j��U�ড়
�B�I�j����&�!g:����� �PB��|�6��fU�*��YA��;s�Z��d7?���Nf��*�
�Z)p �Ci�<�IL<�0�&!�$!�ȫ#��@�<��k�3<�l��	�bxx����Q�<)���W�
Պ�M�.r`��AFV�<�Ti
��)���x�z��@P���I^�S�OLpD��K�*0��u��_�T^>,R�"O�I�6���(�"���SG��Z@�'ў"~�!#��;(��T�Ez�!󁨑��y2�#!� �!&͊g�ܤ���
�y����Z<�Lu�d��C��7�yrE��h��<a�؊b;�Tj�d�$�y���Q��Y{�*�,+g6���P��hO�Obʓ�?9�f�-4v�6��"0Ra���ۓ��x�G-)].`q�P�M��D/ŉ���1�	矌�E�ȓ�� ����4U~Z��ȓrǲ�1&�аW�6�h�L3�\�ȓU�VxQ�Н-���IP�/"Ɇ�:fVehv"Kdl@,jV
 z��,�ȓQ4��T�+2��i�*Ŗ/�杇�I�\��mL�PYJ}��E,,a�$�'L�=X�
ԟZV��H�_6*i��Xg��)LOL��'����,t��ː9E�Iz�"O�Yq0c��K&�9#mߚ'���g"O8 X��X�B��I�T4R�)J"O��V%Ԭ.�t��� PL��"On���^�VӠ��PIY�aE�Kc�'h��'c%��`fi��i_�؉�BY�f?!��!=# �����ppH�r�A�"EG�Oz�����tI�!���B1�wMX�T�!�d�4e�\y�k������;s�!�D׻,�J@g@��'��H�&L3�!�DK_����C F��f9*�*A�)�!�$K� -��X��H��Г�(��!򤃝8��0�C�x�RY�ʓ-a�!�d�Fu��h���V��ԣ���!�((Qp��Q���m��EF��!�D�2c'~=�b�0p^"@
��
j�!�dH�h����V��Kʩ�R��=C!�l��l�1-6�ɰ�<)!��-u~p�V�"r���!j�;!�D�?X�pP�! KH�B���S<1[�{���ޜ.��5�e�Z����Qr�9,!�$�7�Y)b"T#hP)a#d�g)!��<��"\�To�}���U _!�Ϟj%(��ǩ�Yv
� �»m!�$��bؼԩ�*M�e��i%�!�D��A(��!���+}DKd�B�y!�$ ?�}���
b6��DN�L�}����0h�=W&F�#���}�Ă"D���e)��Z&}�'A� Q�u�Ql5D�@�$�Gk���� �E4dТ�ɷ9D��9W�C^��6d�<,.c�Lg�<A��8Qհ-�d��gFL�ZE�}�<١� }?f�ҷ�W	*�Ƞ��Qq�<� 2��۵�����#Żh�� "O֍s�5G��@����.=����b"O�X0ҁ�'�`!:�+���U��"O�`��zL��"B�קj����"OȈSn��,<�XH!�HY:���"O�źsF��� �Bc �)b���"OqI�)�8-�<@���Zu(X�"O��A!$L���@f=(�#g�'21O�BT�������?n���"O����� e���0̈U�, "OD��T�1��t�U�Ns�I�"O֕��g�Ly6�;E�G�on��p�"Of�SG�$h�Oր%�\1�"O��s�+�����e9��܀�"O��r��++y*���)K� i��'�ɊM%� ����,u�U�;��B�	�5w����(�+ޮ�� ��5h�C䉓B��Yҧ$D�4�Q�+�6�hC�	�1β���dD�y��ճ�*C��%G�JQ3�eE�1^x(��ӯ#}�B�IvGDa���	Oa�<��퐠{�B�	,lA^䰑FS{و0YC�ϲ$����$�O��ɀR���'�^�;(�L���kf@ʓ��<��O:�yqeݳU@�#��~�����"O���G��i�$PϣA1���s"O�ë�t��++I@�t@7"OftZ�&ٯ.^I�� ]B��"O6�p��1B��i9��';��V"OT��C� Җ8�b��G4T���'���X]���qCΗx&A�F�8f��'>a~� �q4��N��Am�XQj��D&�O��)���-�~eTfX�ƍi""O�h$��0tL
تpdE�6��d"O��bG,T8aQhHZ�K�_Ւ�w"On�p�RH)�g�M ҆e;"OL���TY:X��
������V��d�O7�]����\��<��58��#��'�2�'��Մ�^B<� ��,Bs������?�	�(�=
G�a��X3b�d�6X�ȓZ�l!�����j�8����_�*(��
�|���� s��]�5��?Z�p��d��3�k��V�^
�nC�	�c�P@A�H�yS�H�v�F�)Gv�FR�'>u('�	����ͯIJ�)���O���d%?A�땻I�H1�r�s5.i��(�ޟ����^WD���Փ3!����!(�ޕ���f�`�j�;<���əi����ȓT����M�}�Uf%�@%��'���
s�$I�uNZ7�\��ȓ<5z�2�P3 N��w�t�Ih�'��IDy�U�n�.q3qo�|h>���c��D�!�� SG4I؂σ�KZ��@ݓQ�!�Ƭ`���F�&`�"q`7�Y�y�!�d!qH�x��>ax^��MF0-!�d�&�����29e�!qP�ĸ%!�-Jhu�2f�/)J�|;DD�c�}���(�d@��
���;7*��T`��j%|Ob���&o	�Y���H4AN���5H#D��x`�.}��F�H?5���H#D�̲ �X�C��ak�JLByF&D�P0',�c���F(�$б#(D�� B��#F����,sNtp�i&D�
`F�F��`FD�y�0���d#|O2b���!�	V|]y��ߩGv
<iO#D�� &��k�FF���ߩaG��0G�'��B������TN{(��`Ƚ!�_�� 5�7��\���7@��!��݈+	�B��!���s#��V:!�$~������Dm��(��չq9!�d:?���ڢI@�&l�K�/ !��G�N2�@A%�x~�����~.!���@K�͐:j6��U%.!��Vd�H��f��Mal=�A��72!�d�&�!s��\�7���Cf�.!��� f�bi�Wp�R��!����
d��@ ���'G�M����L�!�)Tq�b�ʘ���hϔcT!��	!v4�1heNɺ.o>(!'A2?!���*�t\P���#P�H�V&�-!�$��5U��2CCJ�u�j��g뇘S|!�D��Q�p	�7*g�NX7��"�!�$C,�D|�c���,Eh1���!�!�D
8р��f b�fd��.�>ek!�D�/�*	���'"gٱ� _.<�!�DՄQ\d
�a��HRމ�n��!�dM=z�`㯖wI�T�v$�"zD!�$�̈-d�Ӯ3i��E�ظb>!�DЦm�pMZ�eo�@*���W&!��,,*�"e�Ȧ��a �\$7�!��K�[ٺ��n��p^8A��?�!��J�
�Ip��.RD�JFސM�!��;bt� �[/U�~%�s��<�!�$�9��j�I�!C("h���!(�!�d�+�KA�<�6u*���"G$ T��'Ȣ���º!�S�N�On�E�	�'Ȁ�J����m�+C<��x�'�l��%�8b�z��7'W2gݲ��'F�T��G�rMF�����5f�L,"
�'�h���
��]�rǃ�S;�*�'1X��,O�W3��t㙇J\M	�'�
���$�w�
Q�A�Q5� P��'fm�Uoԋ0�#6FƏ2l���'���0���=G���0�t�&�	�'�6Ȃ7�R�#�	�	i�����'ht�� ��\�����6e���
�'@0�H�j��I&���^H0	�'����L.J#�t9�K^1\J�M�	�'�j|Yt�kB)�e�UD��
�'�> Y��הi�b@���8���:�'׈Y�*�0j�.�g`59 ���'e����f�;�Az��V�298,�	�'�q3���80��w� �=!	�'�"q�OI8XrwG�7e��i�'�j1@ �������O2x%�t��'U�шA%�,*�H� f%U�v:x5��'��A�$	�)��mإ�Wg	�'^��rc���`�����\���	
�'?bXꇇ[.�h��C0Z8��	�'Rtb�"��y��a�D�M�Kw��	�'�Qk�#OCLqѣ���B[8��	�'|V\H�)�1Y4(rjU7= ��	�'��crH�`�$�ZA���G��9
�'K�JP�,#bhR��X����	�'�4-������n���!�N��'dJpY�,�%v�N�`�gM2M��� �'ⲬCf�@"����f�X�N`ځ�'�X(���"@�XBG��YU`�
�'6:�� �� ���ЄVo�Q"��� b��+L�fb4-��K�l�X��"OV��'��."�;�J0��h��"O��`���W;8�NIc�Z�: "O������w��x�W�Φ���P"OV}�r��m�a�f�S�%+~�"O�9p��0� �Q�A�~l� �"O�ĲD�+ǈbC��.Hl$�"O����ؽaM��2�,�v���*4"O@@ؔ��6mXp�˰!M�]�zQi"O�-��,;FR"��A��x`@0�"ON�	ţ�)0�mi�J�>Q�p�w"On�	BD�*�9��	�O�j��"Oڌh�$�|��̺!jՍ�"��r"Of�ӗL܁�
����X��V,�4"O��iu̎�m"�Ā3 \��eB�"O������"����Œ%`��"O�e��c�,�䨂���U��"O�pYc'�j��k�2�$ k""O�tHҌ�"m�׉Ģg�0=R�"O� �t,�=C�^�Ӓ(�Q�~��"OZ��Aʑ!mP�RA���m�l�
�"Opq���U9D�⑫`NE�L�V�:%"O�P����GL���P u�\�Kt"O�݈�� <0���/�8+�\`��"O�H�]�� �����zb�H�"O��j�ϲ-�$q��B�$V�x�"O� ��+YK�dA
��"4m����"O85󁭋���I� ;�t��c"OJ� �i@9-��=��ŏ$QJ R�"Ox�4��mNp���A�=�JI��"O�A#�	�P��ɫs�ټ����"O��x��!U�vnV)!��T�R"OZ�c�Ȇ?s�ݹ֫A�p�}��"O�@�!��{����ӖG���"O&Q��#�ox���9ry�S"O��P<ZqhX����&<�Ǆ#D�Đ1Ϟ�@�0|ړ�=@����q�6D�h���J%;��0+����T�����i6D����_+�lA�M�M�xْC7D�`A�땲G KH�8�蚲�3D��q��:2�������%Y��$�-D�d��NK	s����a΅)��� �/D��z���&�*�K"j�66�ʽ�v�.D����R#��`"�ʃ�X p$�)D��`�e�S�<��ȶ �~ &D������=��y�gұ]`�I��"D�ljAkF= Ԅ;�IP���i3D��C��X6���q��3�~H*&�;D�XB6Xc\N��p��k��5�ƃ;D�t� ���GU�(�*X�0�l��CI;D��PtkR��B�����-�<퐁�<D��aN�3n#Th��D<Q�qG�:D�<�Th�sS��iǅY%M͔M*�9D��a急X󌘒�۴�����#5D����"�'F�iA4�2QM��1D��q��93��flNzΐ��¨/D�����l0()9q"��`��,D��J	#2XV�����M��jP�+D�����	{/�P27Iݶ6p���+D��9!(Ӳ&d���o�x��0�*D���b�sI�m��Ę%n����@N)D���7
R):���c�L#��ic`H-D�lb@D�/�H`�EOI�!�iK/-D����8.�h,2p�(9>��R$b)D�� �5i@�Y�:���ȕ<$��m�t"OTx@�%ˇMɊ�(SN�R�a"O�oB+6Tz�ᇈ�m�p���"O���`�Iל@h�HߛM��!�"Oj�p�$� ~�@yŧ)m�N��#"O IP*ИZ�$��s�(o��PX"Oƴ�BK���m��ߦr)�("OB4ȴ�B P���p�ŶFl�3"ON�!�dA��̰Ŋ��p.�)""O��p���"[9Α��C�;6��u"O @xČ�s���!c�Ҿ��p"OF�*�(L�XD� ��c��&"O�%O~ 4Rg�%.�tx��"O�|AUi̬Pc�������b"O܀cq"/�l�!Um��]�(�"O�9�����y9��ӿM+@q�"OLҧK��gnn���N��x'��8�"O ����c��imO� hh�"O�AIE.H�.|K6@?GWv`��"O��C�D�y��Y2�U�"�"�Y""OB��h�M�[�BN�N���Z�"O0x���t޶X�F����>$��"O���l�#S;.$cە�*��v"O
��_%��RW�	]tl�B�V]�<	�+	8�iq���Kb�scNId�<i���\�ȣG�[���c-�\�<��c��?r�����?m�H�U�<i2�J�.�]���0C<(��	�N�<�i����42`��,N/�A�K�<IV�ӱhx��a�;uAI�<q突�f3|�
'ܽw6R(�0OB�<qQ&�.6��qZ�a��_4K�)|�<)�O�;>z�)E/��\�r�rR�w�<�dD@69*���5H�N��ҫn�<y��9vuKpEW0
|�BRm�<Y���2 k��13�C$�4(����M~�d��<y�y�����P���'N�}H��Y��M�*3!�F	?��q+���qA�(I!��
�'ıO��P
�������/��� 0,�NZ!�"f&P�3��Vt�Lp�'���I$>I1d�l<a��L��v�.^x^k��\y8�`��4��'�T��H>,,l	B�S�Z��Q�'���"ѩȩ
����#��Wr��IO�l������-��3S�����Ӡj�1�!��ЋE��1O�e��E�� 2v�qO>����6R����jJ?u� �se�@|��}r����b��*���!B�+a&Ɲ��1D�X�D�֦Q�u���2i�=�1*ړ�0|�u��,���x��
����BQ�<���.�Vl�U��!X�N��e�s����?�c-�Q�TT+�Ah�~I��3T��S��Hj0���e��yLe{F�1�	X}R��c��QN��F�&}���2D�(��KD*M��}a�&ãe*J�&2D�����&�T��:w�u�Q�0D���a�����,H�j�&A�a�/D���'�ݜ^V,\�3Aπ\7�yt+D��;��{�TS�'�0D���eH(D� zg	(%�N�JaIwR�B�*OF	"Ьʋ�4E�R$<�59�"O�0(q�V3s��%��ȺQT��"O��!t�?׬��'�"��e�A"O�ْ��G8{�d�s4�R�y��P:�"O&)��@ՇP��L��lN*f�zi�r"O� 0Yrj��6$���մYlz�"O�9���7Zk��i�*�88P�E��"O�pt��l�V��RJ��uQ�ف"O�y���$<� �B�؈[�� "O0��d�Od�=Ґ��s����"O�$Ak_"�aH���Pv؜K'"O&�RF� <j�Xs@"��)�y)�"O�y	 CզG�1�G��#�	�2"OdY�G��	R'�Pg��T%s�"O�M����>EU��%D�0�*ͺ�"O��
[���hg%��hgh��##��(O?�I�y�RMi2��~��k�(*&nB�ɕD#&�QD�2p*���A�L-,C�I<6^��閭&: �x��ފK[�C� "\ �f�<���a��'�C�Iz��z��Ó4��J��;%vJ�<��T>�b .M�W�zx�Rg:Tl9�b7D�:e	� phL�*uG�b]�"�7D����Zy��ya�@�!+���0D�����(j��؟Y�R����-D���"I
��@��3��|0=��B-�O�˓nR(!pցM6P����	��&|^���-�<�'��
b&>ԡ���V͜@��(n9��Z�e�揁+�\��q��	*�D	�`"X9��ġ1�8��{�,�h�Û�x(� )��U�+kv��W4�	7J"lA�G�2t�p�'%B6T�C�	 .�\�P`��3�pD��J���<A��T>�R���n�ȓ*B�n2�7D����$�K	�`�2��=1�h�b�9�(Or�}�+�a�a�8�$��f�!9�TF}���6$��p���1$*�eL� XV�p�a~��ҥs��Q�EA�Y�r���형���&��|j�|���)�����ɮB!�$aE�ސ�y",�J�f��0�XU�|�w�@����~7O�c��'kR��Bg����L����;Xt���DU`�K��&fj�d)ӇѴZB� ��g��h���&a��h����Hn��c�k���ay���N�qB����߳X�zIqG��)Q�=�N<1�N�>E��'�{�(^kXm��T5FY����'�,����!;�9��E>��@���'ay"/T�ΌL�ҥ�,�RT���A����HO�l�@�|")�HT�ȫ�-X�xS�Ԃӧ�y����hG�:x��xqc'����y��4�SJ�c�TC�}9w�>�<B�ɭ2�T]��f޸�J��)��?)�C�I�z^��(6��%N#�<Q�W�3�����\�q���xz��̭'a
|���K�yB:�8R5��=�O|b���Y�Z��wF '�r�iU�	5F��O���:W����Rɝ-r�t��+28�2C��<E��1��ب2P"�8Ǩ�m7�4�@?�Ob��Mkc���o�ڭ�u�ơ>���1bE�<1�̥D�<����E&[$�Kg�N�<I���������'@�X+N���̜y�,IQ"O����@ڗZ�*��f����uY��d"|O���Nۍ&d)1k�m�t��R0O�����.K���7F�z�ơxAF$��z"�^h̓O[ܫ�	YU�@Z!��~3���	@���H�d#W���8`e2*�>IJ�(D�āX''Vdc �A���J"*¿�y��-tJRBh^  (�P��I=��D=�S�OD�I�P���6�	���<�����' L�C��Ui8�,���ڎ��{�'m��)ɉ}��]*�&)������� �aܬ]h�z��RD�0�k"O^���[�:��t8���I�~�%O��Ⱥ<K (Y�%�7m���Q�+���Z�'�1O�3p	T���˅�N9(�a
�֢���}��~��	�t�Z���l�-��$����z�f�	��p?�q�ƨ��� �{�\����R?��g����'����.�~p��)Rd�?\}F���'�O8y	�O&�+�<?��u�ö0���)�S��y2nQ��4���@?
����+N��(O��)ů2�':�^}o!,J��x+�Aӄ;�LQ��x�Z�l��:��$����d�ȓCev��&�0B�Nu����bE꽅�2�D�N� 5�!r3C4CZ���>q�����lJ�LT�ZQ��-�����S��y�&E1@��cp�̮Zv~��Q�ϼ�HO��T�>�R'���S�(U�t#ϴ!!�d�,��Pr'�0'�z�s��[�!��P>8l��H��uZ�����N�Q�,D{*����M��$���Vg�
��r��3�-�O\�#�nH�_��Z���5vޠ�zȅb��H�:�	i_r��*f�v Z���;?B��6�̙��!z���c�T[!�$�'ўp�G-wb�� hƳO��(I�eA�<��_,H�D��tK̬[=�u0"��@}��|�C �g}�mW*]	�T�5�Q, t�1e
ߥ�yR�P�2Ƽ�h��X�t��IMX��P�)l��w#�"K")U>D� �#/͔5�7�у4�<9vi0D��h����*[�1v�Д`nV�Q��-D��a��E�U�6��@�(�@S�6D�x!w,��5�^��y,���a5D�,Ӣ+K�S.Ĩ�%��nF$�!��>�L��==蜹ca�ϗ&�,uB����Љ�Ɠg2��J!%�!�DR�O@>e9@����K��/|"1����� ���:\s�܅�#��� N?=,m���0K���ȓh���함V'�lQ)��!�T�<���\+v�:#���MF� \Q�<ѵ�Z
.d8|S�lј1	d�`�K�<i �IM0�q�ԩ�J|�Y���
}�<9w�]) [��ÀɊ3*��Y2�"]}�<q	�o6�IAMɯq�K@�`$B�	=V膕8��F�`�d��B�Z;(B������V�y,D��sၻ��B�I�
	�0�� ��wjjY�ƍ� ��B䉕r㎭ҡ�#�
Y$)��l��B�I�Nf�0�V��,e���W��5B�ɯ<�&�,� X��Pa���-�&B䉅zD��m��-�p�R�%	�O��C�	�/NH�@R$�"yz�h�k�kۘC䉛p� RB���A5������	1��C�	$Z_$�*�̝q���v�,/��B�I�#��-bdK�3.���㊝F��B�I�z��h�@̰�(��R�F'�"O�,����P�`���_)GSXm�"O�䀵�_3(���/:58�@�"O@��䘳n��@�.Q/Ք|q�"OfM	��M�U�@IM,l��(s6"O�m��T�"��,)�
M�|h�"Of�ց�.��<�g(ɒ�D�!"O�)�qAS`^ij��OS���"O�XI++|r]���X�D�%)%"O�؀�*�b���@�
Z=�Uà"On���A6}c�	���++D~�"O� ��r�Q�wl��qƝ�E� �"O�hg�m�r]@ф$"���q�"O�4k�]2e�����,�q�P� %"O���K�}����G���P��Q"O�A�qLի%��d���	�l���"O�KQ�'y)��_�婦���l�1O���VJWk��!3�ڤ~&��s��77�T�s\�7H̃p[C�	�Q ��ŗ���$áȳ?pXB�	)T1˰���~ a�N�PC�	�K�>Y�f
��9�J��/��2C�@`�y��X�%���ˎ�4wC�ɴ�D�����I0����:��B�I�du`;S�ڙFq��^0Gq�B��>��*�����v���A��S�'��a�୅�+�4dң ń��
�'�.�JY�?[4�R�& �X�`�'���Krb�bab�2p` z?���1|:�3�"O�nj�В��C�s��ņȓ(Fp�fm�w� -أj�(09�ȓ*�D�[��>oT8�� -	�DH�ȓ2��(0`�&fz��g
ȥrb�ȓ��}P֨�4�����5qwR	�ȓ~2}1� ǐ9)T�����2,���V-�-Q�"�p���Z���,]T��!P��`�M�@����e���`���&yO�u�i�`�%c����P�f�p���$G�2q��Qu�܄�)�<����վ2�vщ�i�H(�e�ȓ-*bd�B*N=l%�]y1F׽
/d5�ȓ[�̓�́*C��$Yc�P�zu`�ȓ���ʡ���x^0�H��];bH�P��s^R0�.	9�������9�>��56�������  %�0�ȓA�`�9s��(d��d�G�'�F�ȓ�ɞV�d'��lʈ�=�g��6����'��aK����He�=`h�ȓ@�TTk "
�E� ��c♼m��2D	%�I�K_#|�'�^\�uOA: H96/Сzs����'FxF�u����4ĝ<u��$����bn����	�>� �l��SPe胊��b����-�$�aM�H�A��'P?�bB-���WM:D�x1���f��5f6OV����e9�ɶL\������IH ��jČ o��ABY-!�d(e�-c�ȁ�3Z�d�F�H?AF��B�{r_����	�/lƔU�ޫ!�(i%��2�FB䉇3��1��*�=��`P�]H�y(�h�3��?�G�S St�heAԷ,����A�BD8� ғ��}}�!�s,�$� �RQ���:�ܘ�y"�G�#��(KPK�J�������OT�a���稟|P�����
S�\ 	WXS"Oh]z����{�4���V*:��r�����գ�{��9O��֎�Gyұ�4�ƥ~!���g"O@�P�+��yR�S�/�A�c<Oƥ�!�P��p>�dV�JK�ur��Y�Y]dR�Zg��҂� k��D��D��ҧ��Jqgi�!�ƖجQ��ʢ[f4jD�Gi&��@P-�/Q?[�ҥ���3R��3 �h�*�c!D���Ø���"��S4	� �"�G�=.:�E�����'���	��G�"q�/�P���B�'В̈U��$c�%#����i=D�D0v��]�bX����*��H��'D��RUN�5O�J᪐�E�H$�,���+D��
�����ɈB�^�xB�s�-D�@0&`�*)�Ȫb�_�2�%�i1D�� �t�1!�~��dg����
"O2����0���{��|���:b"O4���^/*붡a��C��@�s"O$ �EC���:9V��q"O�Ջ�^ {�^E`үF�z!� ��"O�I�vO�
��PZB+Ž}f�ұ��^��P�Hm"�4�%[���:����͊�b���ȓ5��5H1Z-N䱒���Bg��s�(�A��'��x��D���c�X`�$#W-FܙU�'4��׏M�]�v$�����F����{��h�5��"O̆�ɪ@�	atJ	$.�~�	fYi\��	%-�j�Y�NZmX��$�|#Q#Q6g�6����ӕry:C�	 ^Q��y�3$��Ĺbd[�*�O�Ё��]�2)�EE*�d刺(�BQΧp)R�� ZqD���	�T�H<�ȓQ��!�����Z 4Mi����-.�����lAtyҌˊ2b@��DOs����f��]�kPzkG��H�ތ9f��?XvC��/}��I� �������%V�|�L�j�����K��O]����#�xFLh��ʸ.�x%�F1<OB\X!�K�+�l�Nq��Rp�A�$n���C�J�;]���.D�QP��WB���\�\t�D3�,���^r�Xsm̑'�#~R�o�� ��P�L�{���wCFT�<�ᮇ�4+����œ���ɨ��p\h��)}BO����I#��I��E�f�4:���]m�B�	�F�a�Sjޢ
s�ID�J�`$`چ8��!��y2@�8��%�?ɓ���x�h����}� p�3�M\�<�T+��}LUÓ�L�O���<�����=�̈/�����1\��T���M/"� ��ƙ&�a{R�� ;CT����b�j5�I�8��
�P(g�U{D�Ch<�� ���1�&��3��Ħ�y��[}R.0?� ]����:��!��Ʌ�%L��
��Ѧ��l�5��z" �5*��$�'�d�P�O�4�ڸr�EG�H�f`�7
b��{C�*eMR��K��(��	Y��(3` %Rf��c�&���	A БQa�����4D(�lK;H�`���c�L������6���ô�+i>%��I����2+׀;W����@�9I?�I�+�S :S��0P&��D�Y�5���M+4i*�3�,�PA���Px��ì`�t2����6Ԙd�4j���<�Z̀��?ac�	�H���¯`�t��2��Om�"ɝ����B\	7�b|�ד!��;�-?Q'އQ*zHh�@ן@��eN;|�Qxe"F�sd�!Tn�9Q���2�O���M�Cdj�#ak	����J��5~�V�?7_
�����+P�7I�`�R� �f՚!ɷ�:�a��7)�8i��W.|�`��X��>p
��A�Cg�]���R��������,[�D�dA<mt6-ٱC���tb�!m�98f�݊{�&i8�!8.�����тa�����- �2�R��S:7>A�$,z�� m��8�0�NB��w��.�.�
`H�; 66y�Ĕ�x��|���EIH.8^Lx�wCN>%����^u���4o�yB��#π�vT+�,�["\p���o�58�g ��������Ӳj�-x'�u���@N��	F��<��έS޼WX9���#=#��2EM�s��M���ЉE����bO/V�ʧA%�B�Y
�N9s����^w�Us��΢>݆� ��1b^u���4d��$�K<�$+ϻj�P�����$$��2�n�)d��-�ˋKH��1 !�*v괌ֈX�?��Tdۘ���
*�u���.(y���0
'���3F� �P,�g�-���D ��;�|�]T�
 L@ v��gD�}���+D)��2���zM�|���\�C��*@��~�5��{���d9����#��4��JO����:bͲ_;(�1�OF�Z�V(8�~LR�*I4�|ِ���uĬ{v�I*u��x�S�=��C!�L�dR��j����'O>~���*wމ'EXa '�O���s��CY��ߴM��	Ѻy�L(�`��}쒀��O�����Z>�;�� /(<��	=DѤ}��AU?gF�M{�B��~ٚ�kD횦hR�cv��'k\�s.Or��Gdx���g(_>� YR�lF�~H��'��z���+�'P��I�z���	��a"eL�	xEr�G�0 R��H��6͸�T7�ɳ/���?�Ox�E��'1&�z� @N3Q߸��G A�Z3�+��43�-K�{ ��ŧ0"�`7� d��y��~���^E�z��_��@��e�eX�(��W�Iʩ��NKYr�V�5�b�H�l�	Mia�FձHb�K#
V4��đd@5ی�L>!��B�8d��a@��J �0��Nc�K"� � �"�*�D��K�H��1B�mJj#��Y�� \9�Ҵ� A߬܅��aڎ��S[7N(H]Q�N�nh�,8�MH;8$�'i��߮A:��Kt��i4��(��R(.Q:�!`�H�J�<B�	'[�虆���.1ƨ`�I�}��$�h����B�0D�l��<}��� �l�ǖe[��ƏE���K�"O~![�*"]����tH�!�l�얳7��B ��RG9�3����x��c� i~��+�쒯PqO�RV�׉����͋��Ii�Z�m��}>�5zCb£]���F�!�0?1�i#Y��f(�,	�jq�����q��9�M>��!�C����AnY�F�>I��ǩ!�#q�V)��"(Bh<1�"�vЦi���*j.�7e�(+�uYw��?M�����1}Q��>�;���R� ѱ�����(�57<O$���
��8��O^̸�'�W�����f0^6�5�%"O�� Œc�xYYq�T�z�:kW�|R���"!;'+�{�Oed܈bL�/?���!�ћP�\`��'��X� iVd�8�(�K�L�v��S�7�b�'�J�(���>٤D�:z��;��ڬv^�T���lh<A'��9U����YRH����_�P�fT�ȃN_��lZ8V����:O�i�K���'�Z<�t��i$�$�t�C�VM����h ��ԥB�UI�6�Ӌe�����iD�p�� !��%�<x����)�D6M�%�a��6LO&QS���5,r���	�`޺�J�|��I�cٴ�zA!R5��=k���B�t��,(	ys�W7;irQ{r*��U��1x0Z���'��x`��
����$� �jv��� e48s�4�������is���6c��8��_>�a�{���'͒W��Qа%�,|���j@�:D�DH /E�|����v�d-��i�.�Dh��=M�XW��1.��E@ M�/D�~�I�O�	�0��l��f�*y�Q1�(&kP����Y3����u ٬zw.�(Ebwu"A�!o�
^�ٺWGB�W(�!'��Tx�� f�&4ܬ ��!Z9Dl�7"�y��X�BLk�}���2���݂{U<�b�C��0��b�/�Y����!��;6��y��a���ӕE��I�pE�=�'�[�MU9�'則*�Y:���in��7ȟ�94����(�yr"Һqp�UB�*I�8�(���-?% �3w�Y&"����-�"���K?!�1�;�Ҽ#�����
�%Ff~a13{�}b2~*�Z����L�0�>P�G;�1�(_�*Ɇ!s*� l�#�!<O���>U\� �o9��CG鉺8�`2����p�ߴ��{7�^C��Q��dJ��&M5&/�I+�=4�lJ��űHO2�3ү��2(0�Eh�:�h���}L�m�w�O�dj�a��JM0b?�� B�2�qj�E��ӕkB mDC�	=���i�7�b-��D�x��� h����ױ?�N���O�N�a���c!#�,e�$�+�딓jZX�k�)�O��`gl]�x p80�D)*��z���%T(ȁ�҉!H!�$N���m0�,�)wp�hQ�c���`GSj�.0AƠ4�S�	�����̈�,��0ˤ�K�<�~C��>$���{��ρAрT�`�B�0����D�4H��H���)�'s5�	W��)h����QJ )��`�'e��J+���#�g2d�,O�#c�C3�y�� �\ w�^7hO~��Ad¨P�
���	(b���@�<�Lʱ�_ c5
�7�im���8��thg,��4�`��#B�h�F}��̇w�6�E���34���k0 Q4���y�zu*1��H�Y r#���y���,}'���*����1gX-�yr�"Xi�č��0�RA�E��ybDՈվ�h`#d��`F7-+!�ą�F����f:O�@�Y��&!�DW�

�b4�7i��l(5fD!���B� ������x��!�"-,M!�E�\-
8Z�I�brtT�$k�u&!�<k���ւ�M�d�ۢ�Z!!� M6���NѾQ�� I&ݚ.!�!��A�+��2�vq�X�b�!�$�&DҔ��۲h�r���D�!�JT�pS�NL.���2pH�i�!�d��][��ʱ��,Ыq`���' �9��&\�]j�%F�`�N�c�'،%�'�3J�C$��.5B�1`�'���SD�]�\�F��v�Î(TJ��'X��U�^���e��y䎉�	��� ����&d�r(�(M��]�6"OL��g�9t����Ũ](R����"O���`�٤��p���(ɖ=z�"OX�i�oO�_nQ#v�!>Ύ|Q�"O��q0mO�+Y\�1�6��uȇ"O=@�W^9���#� �YC"OZ�YFn�,,mQk����Q�8xe"O��h2�A2rq> h�e�7�fAq�"O��a�,\�G�F"΁e�Djv"O���C���li
���D��i��"O,ܸ0bL?#�LA�Ǐ�0_w��c"O̙8�딾l�q��I��_۶�:p"OTjS䛏/\ i��n�@m�%�@"Of("�M�Y���RM�	F0B�h�"O�k�
M��%�Ϭ�Mر�'�yRM��!�V���j����QR�y򍛪D��X�!!  9b4A�OƉ�y�[ў�����?x��l�f���yR���=Ɋ!Z�E�F ���d�'�y2��9U� x��J�R�)P&��y���'�f�s��M��� 7Iˊ�ybNA�N
aZ���.Q��h9� �y����nl�DΰY�be�A-��y�jY�zoH�+�U�pF��y2N�Y�  R�c�;;���ش�
�y�`U�1;�5C�X>E�0�-�yR�4	���C��@$��c��#�y�b>I���OĠ~�c#���yb4!�1DADۂ����y��$2�@@����t�`�+EmM��y"$
�x����gF9+*�P�
�y���3Hv�Q@�(1��8�䄅�y����z�e�.P�|�q \/�y2i����46�^'���j���y290�	J�Z;	v"m(�O�*�yC"����%�K
B+'�Ħ�y��Y�}26l:������a��K�.�yBnT�BL�yzW�E�Ҁ�����y�-�'g�2���i{FT���Z�y�&�[��܊�,Sx���Ӆ�yr�I
82�PJ��H�S�d��Ao��y�Νu
096a�MưƥϚ�y�B�����
)�!p���2�y��\��)���U`����4�y隮H�q���J�Fu8db��y�Q0NI
H�t)٧��!2�d���*�}�d#� %0��A�]#HhNi��>�\��G͜4*�R��4m
����ȓ<���9���(D�D%�"�Y?��p��W�15�R9M��}yu�,z��ȓ'�TEi������0F�C�tQ��ȓgXH�5��TLp�w�\6�4��ȓD��PP@M�[�PXa2�҈�XP�ȓ$��}��j�b�\����츅�F��d)ho��`��<n�"e�ȓxÔ B�k�$2XY�E,*V�ȓ'M����R%U�(,�$�;y ����6h�����R�8�+M�[V����j5�����?v�q �ج4�:�ȓlH�a"d�Q�w�R����T0.Z<��+�=��	R&4o�i�,X�ȓ)�X���2[W��@ՌH��-��V�by!p��8�R��ʋ	�����������to�Ui�n8h��S�? N�b��P�@F���p.L�=���i�"O|��G^��r�Pb�&W�-R2"O�!�.��cs��C$AX>���A�"O�%2��r����n�(P��$"O^G$T0v�V=�'��'=F!�M�F��ܹs U�!ߎɱF�&?M!��J�l:i[���$5�Vl�(W�!��9Vl�r���]����8aݼC䉎s	F�#D��P~T����8��C䉓,v��btf�p�q���=30.㞌�g���`E���<nq��9�ܸ>쌙����y���S{
�q&�H�ay�m��bD0k<T���PZ��E�b�>�ho@��r��d*z���� ����Ɠ@�|�C����OR�	��]�s.�!Z�ܙ2��`� ���2H���q �4^�*�K��H.����D�5]�>�t�I,���	�<ux�Id�\=Hs��j � �=��B�I=R�	�E�Y޴㄄[�Ŝ�Oڠ�$Z�Ʉ���8�cC���A�C�!���0%mŲ]fZd��f���(�	Ų5����xxDV銎7�Z$�'��-����>�aU�<:������s�ISM�Eh<s�
v[��땣ͬZ*$X0��S�xr�8w�J�X3�غ�
r��sGHZ�/�z��s�A�7����ɣ-�j������
1��ϓ!�.�R/�ov����Ɏrf��ȓAxv�k&�(Q}� ��B~ !'��PC�"Ay=+�'y�O�T��uM������<��y��';��:w��b-��D�0�� 壞,q�L�O���3?�7��:#�>��v�W*� �����^�<	3h��/��y�H��X�d��0�P�r	`�a}�W�1�"�Yd�r�
 � �M��y�/�7unBiІ�v 2�2ՄÇ�yb$�>R?�%�5�W�k��UI����y2#���Ԙ����g��0��h���y�����E�!a�  �pSQ+�y2��/��}��3*x������y�g	���2�O�++�Y"C�	�
�A�t�Q���M��+תa���*�@�lޤw%���J:�Ʉ�&nl��\'�0��_<S����c�v@1��^�8����\3:�n�ȓ� �T�Ӛ!���*�Mp���	 �p�$����6�Q$� �~�`p��
�t]u*R�)
d��IS��p<�ȓ+Z}����t�/Ö
���D⡞<�&��x�!�!Z��QK�x򾥺�޻W�F�EOh�5\�A���FO�|=VI!]�b��@�x֌�O:�(	n����2%����3p�8H��ȶ~n�K�O>%C7�ȶ/躭�0��&"W<H���2uQ�d��ۺ
g�l"b���S�˓o� �I�i�TL�TI�D)Z�I�I��B'��Ɇ�	�M�$H�§ Kޥ�u�(l���huE #CG�i���^�o}PL�����D�x�����1��O�8�"5:�z����!�
(A��>Q�iK�@3Rx��ѓ�N�Æ'���ʧEM�c�DƓ9�<vF�
,|t�*Ԯ�,0C|��a/�O~��D
N�X�δ��	Y��V.e@�ءT��GV�X�Қ��+{,�k�EQ�:�N �'Jhy��J�+1(���V'�v�X
O�YA�
�gK���ө�5��a�>#�xQd�8��Xk�a�![��#*O�D��-��k�bM�O��p���tt}(3�����akq�'6`́5A�?`
��G�m"��a�̣PxQ��*�!L>�"��[/pt�4�'�(���դj���E~�fE���xj�~;NP���/��ɉ�b�����Y�������LJҀp�_>�r�b�
�����35��Qg���<O���a��L5��آ�� }�hT�r �>T��h�!ώ/��G��.T��O��ȊQ�D)k6�Kc��1��Y`Acu`�R�f� �Fd#�%:�	��1R6~�i���4!��(s �X~�'CЩa���9 �� |���P�ߤ��\�$�ͯ2���ҿK~i��	�[c6$��r�|B��/���C��(L��hG�Kg��\�R�z���L>aCE��z��a�TMź����J�	LǾ����5Q��F�d�Ho�? �}�q*ϋLՂ��w&�"��ac�ڴ���t�'O�Rc,�?�F��敨��@����7�&�'�D��O����J^2�N��'�(IC	��?�]��*V�t.I@�'ڪ�;�(�7i���`ƢY������t�&��S ~������I}� ��y0 ߾k_��r���TM�m��_:(�+��¥.�v��p*	m�����B|��T1�J�C��L>�f	�5 ��<�BEM2{�t�xT�[LܓS�Z4��&�K���4lDA�h�ŀV�t��%A�O�H8D�6�O�IPBKA.3t�1��X�E�l;��'��Od@]?u��͘W�V)�O6��$�/k 	(�N�q�$���O�DH�c�L�:!z�i� �F��;(��	�"G�Q�����O1*<�'�:�2��s)�{����;�>���i�x��c�ܙ� d��IB"��1�`@�ȓ: T�����'�J�aSJ[��9&��I#
Z� �%�#�*e��l���1;T�4��d��-�C�I�3�~��愕5Lo�4�pi�<h1D([3�	��I {�v���O��A��HP���c�C��ɃO��q"��"��<���_��S6�$�XP�� ڛ��w���ϓH~qQ"`;�I QQ�wC�1el(�t
`g����	2mx ����M�� 6�`Q�6�@��|ȥ��oz��H󊖕�M�W�� �|}�
�6�&��'��xA$EG$ןH��$�@�K��psoR<z`��g�5qEp��$jЊ5�,�#lT$U��&�S$��F*W���x��7���$!85�~JD��zi��i�,�B�T�G��� �,j*A	�	�|�� ż����?p6��#�+Z.�	ХG�<a�l4n�����T��څd�6\;`f*����`s�A`�,�4 l���S���_c���f�H�U�lx����ɛ]d�4�u��(D窴�c*³3t 2��X��jT�
*:�: [��G!��<Yvɠ)زdvfA0NȴȡReRe�'��|�R�ٚ �2)�rgʗO��u{b(�U�Z0�R#�:�H����ܶE��B�<@�z�3bJ:6j~I��%�J�\˓(�Ԉ���B�{(.[UO.4֐���)�|.e��e�0C2������!�d��Y 9�S�X#�$��,�:-���UB:��1LR�[�\���~bD�d�:蘘����5=��Ș'״����DڇX��a����,�&��#6,×dI�u⤠!��2k�t���S2M��󄓰[��8k�c\�0  �odў��t,ּ.���7`�Ʀ�Z1�B�1��ɲ7昢?�z�Y�C�(��A?=b��Doc\5Y0(�'��bd˸�yFՒ�fQ�0n�o?��63��$��4F 8H~�S���8��)TFJlY!�D�N=���"��hՔ!�@٦?V�˪>!��і��C�e֧A��v�y�ka�@5O*\�b����L����|���Q='�r8Y��D۠��'B��2�XZ�O8��a�����X�׀X�Sx��C!�	�L%k(����P�~
�N���2��Κ�jn�Hiq�Yw�<�p͈$@���Ce��U�l\A���ğ@"�쀾8^��x��>E�$��`�28v�R	ܼ��O�*!�d��/��A;�ț-.0XK�F؂ �"n���X��`
ay2GS�d,	�ʅ�8`B4�C��9�0?)Cb�;;�B-�a@_�X��fϘd�v�ɵ��	��xB�J.F�h���ݓ_a��c�����O��r4�F���~e˧����U�Qd:FgrRd"Ox��ט�V<�5��&V�X0�"O���f쇕7'�B�ˁ{^@�3b"O��QEf�@�b)�p�Ik1��"O�蘶�.I�Q�iG *��!��"OnĊ���N��@���\�=�v	ٴ"O�������qF�֭W��J"O�U[֮��T�<0B��O�%B�,��"O��A�Y2 �,�2UG�=U��`"Obi�r�9;�8(xv��i\v��a"OJ1`��)uH��;~1"}�"O C�I25��tI�%'3l�"O IA�L�k�$<���ݹj
���b"O��A�'ϼ,Nxp�I\$a_�E��"Ovh9��̷(^�Uq���8 X2�HT"O� f� $� �^p�q/��,HX��"O�l �.�	OfUF�G� ��c�"O
�A�!�1S�X2��u'Ь;�"O�ѧ�Y�w���0�˄Jp���"O,�s�E�.)���X"�L6Lp�"O���!�)8Ą��Y�X� ][G"O���2o�-}�Q$OU1I�p#c"O�K�KY�Ui��¥��|�|買"O�\	�.�P)�\�RaC�]n�% "O��vG�,�����i�����"O���3Eڌ!�p�B� 
 B��U�"O褰�AS�c�H���a�4U��c�"O@,ʗ�\�$�̭Jao���U"O8t����HM>EX�Ś?��DI���8��x1Am�$~���$�RW1O�I� ��X��QBc%�"��Ű "O��␉[�w=⸰�S$B�4��0"O,��Y(j �aB"F��w\�[c"O�1���\��2�F�]<���F"O�h�E��&9\ZP0�%�C5���S"OF�!��ˀt��E�(-̝�"O�tU� *`z �q��C}~ ɇ"O����ԁ,��x�J�;���S"O����R�g�~,#WI��W�@�s�"O�h�"n+"��5����b��IPP��Z����t�L��VL/0�,�82F�	1e�mI���:h��㞢굮��mr�I����?$����4^�X��O��3�Ł��0|b�*2g����TH�0k<�`�bEI���6a�zP�F�F
�0|��lX�'&E1��Q��`���J}"	�,�@0��7�哧g*0)1����]�,�rce��#�^�$ӒSZ���u�"���sӈ��P���D���+c����nZ��t��*�����N(]"��EM~]�Є�G]ƀqdA�E��aGC'�F��ȓU�@E�S�p�{%��A�zȄȓ��e�%@��%��j>�rĄ� �r؉#@`&p1�d��p:����$�V��%2�v9��ˑ W�}��X�ʡ���"j�q�D��B��k�'ў�!����/��0��e�S�?�|ɇ�[y�8B�X0N�U��W8L8V���0vPay�Z�~d6���^�+��-�ȓ�q@3&�.?d��d�R0)�X�ȓ+��L��;v��f�1R\��-8�|1.׌v)^}��Ң,o����� �P��͋.ÜД�߹�����;�X�
ա�<q����$�7���ȓ���!�K�2���QH���ȓR � ��-� �c4��!�����*�J�%IŲ�h
 �����0ziS�H5P�	���+7Ш�� �E��ǰ-���T�+0 P�ȓż��fOP�-��C�HH$Ȇ�2A$�Qg�Z2D,�xd�P�#%`a��T�d�a��!�Z	��\?��ȓ�4]jB��.��|;�DҒ*���ȓWUj�X���/.�5k�Ċ�ф�-j�rq�K=>�����:A�>M�ȓ�X ;��S�NV�sDͲ����ȓ#�ז�8�# 	N-[v��ȓ-f�jCB�y4�4���v����P�<�ɢ����AoN2*PB�I�|lj�V*E�
�֩�B�G��6B�>!�H��+��!K��Q�%7�fB�ɷ�,�xf����xA�ĀXW�VB�ɤL�a�v�I�J8V�$ �2�B�)� F�A��@/IX�0ñ�?8���"O�Drԋ׋0$�K�&)��,s"O�5s7�\�T9�x!�Ϙ�e�� H&"O�$C� 	���2@�4��(�"O�%i��X�#v��`C�0~� �W"O���6�Ĝ)��"Tg�]|�Eh�"O� Z�������	El9��g�@�<qC�I3*1Y�O��v��u����t�<%eC�0�\PF�֖jz�)�+v�<��	k�3A-�	v������TZ�<�䕣n͈�C�ZȸL��FS�<)���"\�r����.3�  $��t�<Y!�B!D�t33���FX �Y�<Y���[V� `�6zuXS�<��䗕4�8�i֥�'"�b(�-SO�<�Sğ�n��̫�	P'@��cd`E�<a�ꀂov��;��*4��#�i�<�@�?�L���㜕�:�����d�<ɄR[I�,س�L�,��q�W�J[�<�SÄ:Ծ��nυI�� �/]o�<IueA�(�A2�-̓_��q�vQS�<�ԭ%"[�|��X�oUn Z��h�<a������EV#i��(QAo�B��hg��C�	�7��(�d�_�C��>
�;���	y��c F9SC䉴&]B�����<��鵢�:\��B�	�x����Õ-yxpq��ɥn��B��#߰�����.�%qVo�5#��B�	�G����jF�;����D6?�~C�I�>��e(�Iͬ$	vE�"j/bC��[�KG������+[5v_�C��&�@��G��æ��cnF%�zC�	�`����a:$�<c�FO��BC�I�EG���3	ɡ����W)	�S�<C�I�e��`0d[,}���ډ.�B䉅�, �D�+<���"�L�u�B䉔gj��X���#Ŋ(
���	wxFC�Ƀ�u�nѾd�j�ۧ뙺#�0C�I�%,���d�Q Wt2�����-�C�	�r�@��`͍{� h��g�@wC�I$p�h�D�Ӹ3��`p@N1TO�B�I�71D��UB��u狦PD~C�	,��B���	5�"eA�U�t��B�ɆJ���B��c_ͨS*�B��B�"���B#O�_i����LP�6�<B�I&`w,Dz�%rotݰ���qi0B�	�9Q�ם^nf-ђn�L&B�	�2�T��2燡"�8��k��[�*B�I�4<I��-e; Y+m� yc�B�I�y�@UIQA�/�7*��]��B�.X���B��<GBj�E���B��9I�H+�/+���
�5�(B�I�VY��N�*1h37�	'B�	$u�:��Ȁ��<@P�~��C���P��+	��`ء��)A�C��	1��JnE)E�"a7�(O�C�	�=6z���A�eo�����9:B�	�+�U;C��#E��@�C�Q�!0B�I:*�UPtf�4C�d�J���^C�2{iP��7g�/(t��%��6ʄB�I�]sr,���+;,LXRE'�|B�	Dh�0��ꍋA2���hT�\B�	�E=���,&(0rxp$!�=Q`B�Ʉb�JX��R^R	 SK�4"��S�? �4$g�=3��-�4l�&|����"O>ᚶ��&��}�7,0���W"O��y3o/q��Y*S���o�~8Y�"O�$����C�֩�4�ǿ�r�Z�"O2)�'�϶9V���׊O�<�W"O�X GF�t�&��fʌ���`�"O�|jw��v�q���Rhg��2u"O�lAd�%[�!��͟��e�R"O��7��\���H3/F��f�B6"OD�`��*lI���-�����"O�%��bǤQ��i$M^�j �Ic"On�Zׁ�J�P\��)]�U�YP"O6��#
,=ڦ��h�r^��w"O���a$�"���b�hѠ�"O�U(2��p��:!M�L^,R�"On���n޼|��̲5F��Qp"O��Ig���VȚh����Y@l�rC"O������=gk4���
!u5�Z�"O��C/��#8����R��$���"ONys�bՌF"R��Ӑ��J4"O�!)�C��t�.�S�*� DXp��u"O��s�_]�,�ɖ�5�z�u"O��@�O�4��q�T%+�v<�E"O�\j�MT-&��( @C<Hj^�Ó"O��B'�c���࡮��JHثV"O@|3d�L����"���3*���"O�|@���"&)�p�
n\ kC"O�5j 
�\Ō�f�X�)UT���"O3�ȟ;>8���m�/>z�,�yrd�s��X�R臤h�z��6����yfJ/<ER�XCg��/7��ti��y���Ɩ���d�$2����ME�y��_�v��X���>�<��Q��+�yBC��h\�'Ȅ���+�ƒ,�y��L�*���f��b� �Y@$0�Py�j�'{�&�b�G�k
����D�M�<ᱩ�>C�lm�՗UL�"B�IJ�<��	Y��(�IN�_��0�BmQB�<	���`h�ݻ�כ��(�a�X�<�qk�A��IRI�-�����^�<��*�=M$��G�)Q��CEjN�<a���t�f�r#����z�H�^�<�� K{�P��[⺐��F�\�<9�dܵ%���v��x^ �"�k�\�<qeO�r�t��ʖ4e6~4!��^�<ɗa�'{�|8��bճ|���g*�Y�<�&�̌:�DhӋ\�\��]���]�<	$�Ǘ5��HC�YB=���W�<�C�)F:��$��B��`�[W�<�R���n��B� =w"٘�D_�<�CQ,~]��XR�ų��qaO�Y�<���Z�@(X" &�d�p�Hq�<I/T�1�tu���bZD�-Vq�<Q�`9քd��A�q���s��6T� �)�HYf�f)�,t�����'D�`�Մ�W;�Q1У��g7B�aW�)D������09��Ĉ�mҥ�3c)D�ph3��5=4(��F�D)`�q�E'D�ت�le����Q%�,���o1D���pȏ�p��C�C���a���3D�X�u��0�Xq�ún�M ��2D�49UR�G���TLW�GgJ�r��.D��y�&ځ�&�H2
л��p��+D��h��I�N�\�����;��Kc+(D�� ��ZS'33���#eT�3�r��s"O��s����V��iF��%"QF��4"O�u�EÊCg�[׃�<HKF�!"O
��td�r7�b4��3���C"O&��O�)��HYL�1u�`��"O��*��30�"1��*AqW�ġ�"O.��WKU'@�f�.Y�ܡ��(��y��A=�j� �#���(�2G�4�y�����lS�L��U�]��y�IdY�栉$n�5�$E��y򀐱 ��(�U�#�ZM�䏟
�y"j�&�|5K"!%�#�4�yoʁ��se%Ĕ|8����E��y2�_<Ju�1�A̖2��ujC�=�y�[�_��@%�Y�xX�S���y�i�*z$�QS&EG�rM3���y�´T��|#Tܧs�ny9����y��zE*EBņ�=�DK��@�y� ��nd�K���+MZ{A�P�y2j����Q�F�̘O�	�7����yH�(&x���?K���	'(��y��1�R̓@�9T�eS��C�yF�	)�
�8b�!{��͂�H��y�,�4����v��^����K��y���g~&�h�T���yud ��y@2I~��Ə�VzdB��yB%�W�M���$�Pa��S��y��)RE��C���,��Y��鋨�yr�P�~��ڶ�^�vd)C
���y	TML�]+�J�˼�Ñ����y"��[��M+��Y)4pv|SQ� ,�y��	�,ZLh�䕆?E��W�L��y��ߚ2��@�1��n.
��&��?�y��J�]}����eOPHG��yb-\?�n��0nO�H��Qve-�y��'K�8�ׅײ�E;6�
��y�Ʉ�a�ۄHӮw�j% ���<�y�A�FV8rP�n@��y��*�yMH� jt���
����B��y�%15	Np[p�֎���;ե���y�T#!����.Z�:Ѐ�`� �y2���O��`	���h�6o�#�y�O�w����S�;v����)�yҬ�$ @  �P   �
  �  �  "  g)  �1  8  `>  �D  �J  �R  Y  ]_  �e  �k  %r  hx  �~  K�   `� u�	����Zv)C�'ll\�0"Ez+⟈mZXv�扤���D�R��0AF���p86�
 ��q�"��a��J�ȗ�}��@���{��`��<��A�'+)`D{�'7HT�rU��%%����z*�+U;� ���Ǯd��3q�(���Ie����V���+�eɃ��aJ�H#����J)[��#��I�M�r\qgC�J.�A:�4<=ju2��?����?��4(j���2yu�ݳ��(),t8r���?��H��?�(O���  f�<��?!��&$#�43�� �@� BЭА�?Q���?q����$�OR��w�'��d�OP�X���`[�����ߟh'N�q�n/��O�6G[�@"'�ۧX̨���.�~!�l�'��D�cTl�jDL,ZPh�@�>�`�B/*�2�dLҟ��Iş���ğ�����(��d��4��Pg�H/`�J1:��+f\6�;��'��6m����4>����'׼6M-DǮ�o��8��h��`�4=�b�Y
��	��C8dY~=#���Y9�ȟ���Sʇ�1��HC�Bɷh�X��-?�]�jֶtJxY��i�r5lZ��M��'�BV,�0�v��ҠJ>6Br�C�ׇB��
��k���Ǐth�����Ǖ^Y���L��|���@��Ƭ�r6-���]+�4<ʙcR�$zp�p�#���xQv��9�Lږ�K�M8��,tӤ�n`H&M���۰s���ǋ�4��1��L��@ d�Yz�0JCB����p�$ ��uh�4
k�&�b�H���ܹX�ұ;���6
<�Z���,����&��r��5�	8&l�nt`�DqF�_6i��4��2p��IL����I�ŝ<	��j�U�#vnI[����'��'��葤,nӀ�[��8)��[,Fpp0��Oۍ2����Wy�'6"1�lIP��=����ue�t���8)���r$fޣ1X�%�DC�=9axB	�?!��qKW;�]س�i���(T�P(f�h��+œ�7�@��I֟�b,O�L��
�-�Ze�#���|Hc�'D��'�O1��5eO�̛-#�@6��Gd ��D{�O�7-ɼXf�q�'�[*6��� �R4|���oZp��
�d��B�O�LȈ�J(e��8H�-�du�"O)2r(,�����0t�-��"O��F͇qg�]1�JڬI:�9�"O����%ٻ�t���C:~�� "O���aFH��	s��E�d"O�t�2FN-�����M=<�d9��'��*���Ә�U��M��B�H�F�%�,��D-��B���,R��,a��˥^��	�ȓ9�*��IϔxK��pS���~�����	���K���[�D����ȓ~-p)y�S�> ���A"M\�`�ƓC1��+���L�!{�D�;;�����K�����O,�d�<q(���S���a��r7h��)b�R�o� ��1��ԺE��Q�'\(��M��vex��Υ]�bm#d	�k��X�c�[�Gf$��V
�-t��آ��	>,V�,#TH�yj����F2��E�O�5lZ+�HOn˓��$̹(0h�
={.�,#�:^���'1O���\�g܂衆dR�4��pb�'��7{�nZ��M�(�.���m��]���<q$�.f���E�L��3��П��'\2�'"�铻2��Q)у�7�	
F�'��d��,�P�01�e^�%��q�'��Y�4F�����068}l�jW�� 5�0�C[+�|0�t�ռy<c��X�'^B�	�\��v-e���dM,|���C�	e%��9v���%�˓�?���i�.��p�%$\e4��PăV�E��O��0�'<��H2�0���.F4xL⢭E
=h�6-,��X�z,���=�I�?�+�(��h�$�����!x׊D���ȓ6�"Is�.y�(A/ibBM�sl*D�#�.̪o|��:�H��JD|�"@-D�l[��6} t�Ƥ��K�V��T -D�h@�
^K
�2/�C�$�G D����C�Xk�Ѳ��_% t�k]ͦy$��FB�~�g����y ��y"DɶH���凄�)]ʑ�����&���l�(�n��OC���W�	�j�T���*����aEF�!�ؑu��>�xs��P�
]t<3PJ1�S8<���Oʍ���L�I�����-ɕK̨���'k��%U.�If��4���Ds� N�M3��0c��x��I_x�L2���4%Yt����]���ҀT8����p޴���|��'��@!~�6uK��N� �R��AKB�R�\�B�K����	����oy��J�n�dڔ��#���%I7M6�#g�J(zϚ�Ѩ�38azr�Z�TG�iX�
�6j�r2"^���,�CeсV`<4a����#
7�5B����dĺ:�����F�_�M���L��r���'(l6��<����?���?����I a����Ж?����^�@��{��$]�>���y .�������Z�l��':7��ODʓ%�^�I�i���'ˌ	�W$I�n��HEh�!A��e��'U���T���'�rD, ���C���w�eh�<�� x�OO�[��͓�'��$Պ�yw�';4��H��B��D��wY�7͔�\�R8B�ڮg�`��"K�k~!æ��;�(O����'��,g���z+�p�#6����nѰa(C3_3���?y��O�1O����ѿ@��P��G@�~2��ۇ\���Iޟ`�?�O7n��H�W��8#D(X�R��0���*�Z�������M����?�����dT�?ٶȉ�>d�@E�It�� {���6�?i�\Dd`�����>!b#C�d��ԛe�6,� ����E~B/O6�O>����/U�U��p�~@{�A>?������N>E����L�(��9@���q��E�5��C䉺H�n0��Oʄ\`xA�q
���?A6�S�S�T��S;8x��!�˂Z�Mlҟ������'L	sQ����p�I˟�;M�V���X$�v�z e
��mK6H����-!=ҹ���~���� �`�x�p���
_��#%��f��Г�P}2��	������y���jqt$�CKTP���-�L�vam���DE�T���E��gy"�w鬅r�Gя�Ġ���;q�f	���'�� #����"<��Qè�/�d�VH��������d�<1������dƏT��u	�J�?3��#�&WhD�r%-7K��D�O�D�O�q�;�?�����.��B�\�F�O���VU"�t�&�3�<I�K*1T(m��ʟ�C����F�?vB��+3T$�+�/���0@Ƒ #0x�K���OLą�	���ɖ/_&�战�-6[��B䉝)��9����W*aX��C���OԜog�,�|�!ߴ�?I��V��#�̎�j#\$ b���)��:��?i�"[�?���?1��5)6��a�Ҷ��|��wŶ��f�+)�<���,r��Ó\���C�����qS+Q[>��A�rua"�ʋ?���ȴ��Pp��i9�;��M��1�Mc�V�H��f���7���V�:c�<����=q׈��F���iE*Rh�u�0���?1����(��|�!�'w�(�b߫o�H�CkG�R�	b����$ʰiODil���w�0G���1T��اE\CP��i��?����G2�0A�1�������O�:�"JU�'d����Vl�x�����9֪�=�\Q��S/U3�}�䄄o�:ś�~�Յ��-l(y�!ϔlO�e�'�Q���?؛�j7�I:�ӮbSUL������堂�:�H�O���&<O��%��=�2�R���Wfk��^�'�2�f��nZW�	#I�JA�4a^>1�8a��1d"�<�ܴ�?����?��O��/�������?9��?9�wtd���d[(p ��T$A��$r@�>:�9���J�@�΃���)<�y[�l���
4�p�����%0$c?P�؅�C���9�aʝZ�'o��Ir���$*3M��J��^���*⎅���)O4�B�'����?��y���OT�Y�>~!���E臩���?���0|�7 ��uh���񍕺/a���iv�\�����İ<�(����<���|@�*Q:�09Q��K7X�z9�p�
��?��?���O��$�Od9�ƃK�6�(q�'�$lAD"G��<?�z�P�֓D�~��Ď�s�x	[��ʛC�|2�U,���Hڨ\�L<���l؞L�K�lr�A3V�#4K��*����>hp�]o��'��ם��`�	I�d��0�������v�~��@Q���Dٍ7�ң=��y���6"�8�{ �^���DC��8����O�lZ4�'E���`��$a� p�iմ�6I@�C٣$+�uS���Ot˓�?Q��?Q(ɥ~tPM	�*��U���ۙ'�]��%�KAT("F�S��,�Ó=��;���(`�+栄4U�|��o�r���.�rt<
�c���O����'�7��Od���.8���J�R�
��'���$�O6��O��$?�)3�	9rʁ�5��9b4N,���6|��D{�O|6�DJ�Y4r��f@l��y@�S7cbZ�0�bmJ��MK~�O����'5�ȡ��86�8�N�+�̰H�'+B��;H�=�j V 0����'�TL�2oʝ@b�SZ�+�Ù���'8�!1�
\je(2�&ډ�q��Q9lo��Y���B���(�γl�I�@�n��ݦ�ܴ�?��	�Ku����\�mqb��4r��'��'�ў���hQy���]�H�97M�(@p֣=���>C���o�N�O8�U-K�(��$0[�",���OLYq5�>�i>�<�����Td!��5�ų`�MU�<�U�M�&_�A�r*��2\���'�[�<�tNł]a�1�Ǣ�	Y�j�ڠ�l�<chC�isF��f(����I��^�<�4@�>&�jp�l~[�o�[�<Y��,U�����L�h���'�y�-��p>`�W�]6����cP�x��9s� J|�<� u��Hޞ%s�X�0A�8i(6 �f"O�I��V�
*|QQ�B,qrԨ��"O0�H�	\X�p�{*Q��"O�	���wn�dIF�>L�ލ�'+ p��'è�H^
�b���d4����'�V���fK�^K�epaNYO��EP�'3ڥ2����%�Ȫ���55*B,	�'b�� �b<'�X�#/�2,��X
�'���
��rЂ�GU�5��H
�'���'N3�i���?S��Y�����Q?�@���+��*�[�3
y��$D�d��� �KO����K�"�����#D��P�-M�	� -��.�&�Ifm!D� (3��(T(�U��+dfJ��ҩ>D���f"]�yB�34��2&*!)s�0D�h3uc�1Q[.�%��5�`\�`�O���B�)�M��6B���X��J����S�'0���{R #Ul�.TuR�
�'btm��Rf̌��dN�L�6)j
�'�B( �k��r�٣��E�fL�	�'B�a���6z�˲'��\�	�'� B�K�tHµ�!	;+��xx.O,�� �'�
�9%�Y�>�H����%%�X���'n��E�Q
,Ξ�k�W�$��T��'��t`��>v�q�ǃ�h3xȋ�'c��"�ʑ'	��Lb���4w36��'����0A�#$S�D�W��tL��
���`��4J�-�Bጽ4��c �D3x�`�ȓ���:A��[��8&�ǫ8B��M���Q(%-��ݒSʧXgb��v�>���a�#������"@۸��ȓL�p��Ed��t����@ْ�p8����頒jX;�9����*�hG{�c	���\��0@Oy�B�Ss��1XZ�MR�"O��"���]�:U���&Y�6���"Of�K��O�0c��j��Y?4�X�D"O�J��'��X� ^2T{`��"O
1����66�ţ!��`t���"O�!�˒+[���b���9v�\� �'B�DI���S/���a�嘫$��Mщ[0��X�ȓl�݉�c�2B���Qv��"����nH�&E��t(�E"ˡz����ȓW��1Ā&:���p!c�3��e��Cn4�!Â8j� [	.P���5c�*p-C'0`�d�W��+����'b>}��e�p�@T`
@lQs�lŅ�Y ��gV�F��2���9d̐�ȓF-��̀;U�ޠ����?��U��G �����S'�<H�o��&3
Y��M�\I��c�H�yE��6F��Q��	�9D�	1gJuG���z� ��欖p!�C�ɋ6�Ɯ�3�0�����բ5��C�o�6,�`)G3�ȣ���! �B�	�9@��T4A���K���\YlB�	�.��FG�4�$)�4\:B�I�6Z�83��;ƭ���U�(�=YgKXr�Ob��#�Ϸ��t����e�,Q9�'+TP���V�t��c�-H����'n�y�OI#z�]� ��u�����'�����@7
L�Hc�� �*a��k�@�Z�� ��a`a�u!���%�8:��P�)�p��Uğ��T�1�S�O��A�!A��K�5��@�
䘈�"O��aq��ǆ���5A�����"O� �!z��
Sъ�9�����A�"O�$��+VE(���鐲�H�"O)���%7#Tl�s)Q2(O� Ba"ON0��Y�/	s�O�6�|���T�@��#2�O�h�
E$�4��0�׽j��P�4"O>�:Q!T�J��:���4@�*Uy�"O�Ta��=GX�pjU�Nf�=��t��`�o�?1v|�� �V$
��� 1^�L 
і�xъ������$�'0�$�;�JD����e��E�t��p!�D�	O����K�Ϻy�E��&P�!�DE|:f-��d�0\	t�!��!_�E�AO�9�nQ�� E�v�!���#+h\�ȕ3��EѥD�!�d�2�N�xA_;A��P�dȚ�E�ўءWi3�')[x}�R�\��HH��*�T5��]���`��M��Z1�fա&mL%�ȓ <D3S��>c�.0cb�"-�,��=�|Ac!�2CS���Ȣ=�d��n� �I �ȹo�L�"e��v��ȓR��#�&=E���A'>�"������"<E�T�T�"[r �V�����g*�!�$��f�H2⎽m��$jg
�:U	!�D[$rZL�'D<z�4�ڄ�I�P�!��c��)q�7
8���W<{S!�D˛h�4�;&�
W� ��߂1C!򄊵Z8�Q���:_쬝�ƌ+前E����+Gְ��(�杳Sf��w!�D� o<�k�oV)4O+�Z?:x�ȓ��r#N�-z4�XS�ʅU�0��m�@����ϮF���Q��>�Ұ�ȓ>$� ��A.�,�g���(d��	�q}����r,ܹ�A75�v0��I'8��C�	X�\t��$�;tP4�uM,�C�I�o�L�cJVb{.\���̐	q�C�ɆO�2ժ�� 3� �I54d�C�I�g<���g��p3&u0��T�V�C�r�@�Iŭ��2Hb0�����=�m�T�O��H:�'H�G��H@�4DȻ	�'`\jJ�)�X�"�ɜf���K�'�45�w�_W@���Q�+r�<�
$vw:l�qEՀl�NY:bFj�<qDL��D:H�8�G<�n����c�<��`B�(��-G:"�Dٛp�Lğ8w?�S�O�΍�Ȗ�"S�����\�^PX5ۃ"O�!�F�.C�@M�' s�P��"O ��D	�%@f6�@ )��;�8ڑ"O� q�M�/ �R�zV��7����"Oz�҃�L�kn�[6�@�[�DĘ�"O~�����[H�X�'�8�i�6T��ҕF!�Oz�-��$�C�,��K-�9z "O�Q�[ g�!�q���_���s7"O>�9���8�^
$�5ct�cF"O­�৔$e�N� ���H�PA#"O*=�6�P�I�\�q����zlӖ�'!��(�'G�\�F���nS|�@��	,4F�A�'� h���׋/z��0`	( �Ѩ�'mF��GK��^�(�#�Q5M�
���'��#�̐�C�Ԥ���۰O�@��'i���D+\"Y�n��qNL�F`t��
�'��P�&=����0��t�j�:���G�Q?��l�8z��)+�EBR�fqyA�&D�h`$�	-1"|�3��U\@�ڵ�?D��rR7$fV�"aBM���0D�� H9&��;�t�p�dǚ,�n��"OPl�%蝯\h��Q	��&�%�"O u��a9{�|�لHƂ%>�%�'��lH����%���	?T/fI�� P��(/���c$�@��@��A�X���ȓ^�B9�dH�_1�P�Ѓ:H`���^���c
^�o��h*�]�`�ȓ}LL���G}?ZRm�>SfdU��cx�r�'�Xhä��e�'�b5��]���b�U2�. +� P�~�ȓx �%�C
n�,�h�I(�����r��VN�}ޜ<hBfM�=xd!��7� ڴ��v �5���w~\}��pz6�Zs��=)������dԬ8��	+R�	$)2���4z��a��
{+C��uv���$��dh��i����.��B�ɘ�20��Gːܠ��F�y�B�	�ubXa8�j͎d:��+��A�(�B�I'�D�d�� ���l�ZͶC�	����5�T�W
a�QIW[^�=i0��K�O����!��-�z�C*#VT���'�P�b��/���B�ϘKJj
�'�&�	� ��4�:R"�h�	
�'=�����U/7�@�@☰��'�X�2���L�́ ��8�͊�'��%���H�3��HS���#	 ��� rYFx��I&'L�E�E��	<F:!ZR�E�r�C�IL��d�u��=]x.�YT�A#xC�Iq5�E�5�e�haHؿI�~p�"OT��ꀒM�r8�wD�d0t@�"ORM�@
^m�f�2a�I@�v��ODՑ�+��+H��f'���9ѡL"&E�W8���'vn�R���MS�s���I��9�R�́g�B	q�a�g�R����^͟��"%�ԟ����X�,��<�@�ÃP�R���|�ǹ���0��p��bSoX#>Y5/�nsF]s�V�$7��:a
�m�H��#��y�̴9F�3;ܖ���Į��<A ���|�	�'s�9�&�X�b�cå?L
0h�'Da~��S
@��4q�aߛp��p��h�-���hO�	A]y2�T��P��Lj2,�6ME����5]
��lZ�d`�IA�Di�;V��t�'] QY���&-*�a�kֶd�F}S��'��CQ�-`Ӫ�$�X,��l�|��d�"<`л�׾Z$��4�]�y�f�!|��m�&DX�s���*�\��$��+Ҋ=�А�G%�88i͓|�"��	����?��'>�}&U*z��d�U�Q��s�'��4��Q�U�����,���	R���L�OvRP���ӜxM`-�!���g�=����0#�O����5!������iP��g��7(�B�I�E%xXY a�=��e
'%���B�� rq�����7����B�Ի��B��c�d܈
������G,.!��̞"VXy�D�+!�<`$K!!�^>#}�¤a�@�
��A)BP"���p?)2�O�Fp��B��߆�h<Br@�\�<�v��+t�Z�JC�Қp�,̩Q d�<! n�[w�YzD��iV��R!+T�0��ܭh	vp��?fx��rD1D��z��F�Kݞ	w��$Z�vl*��.|OıYB�>�1@��b �yUM
�W�\����V�<���Z�bά�#"�ƍd���V�<a���0a����0ď�����
O�<97B��lɊH���*b �E!�e�<�w,�21k6�Kcg0<fX���]�<tă+m[�$ B�,sF�}��l�~�p�`�GxJ?1@b����6� P�ds�B>D�t��lF,&g�YJT�66X�ڕ�0D���nN0R�$�[�6<$��s��.D�� ����,����/�_& U[�"O�	p�y���X1�PB!#Q"O�}*�&��J�XD��*aLk'��O��}���L�
�&��R>�P�wH�`"X��C�m��./���Re�Ki0l��H��Rwh�-�M���� �5�ȓ��ӡ$����D�?�I����	��X(a��Db��u��1��ɾo"y�
G�#����b޼�e	$f�cPp<��f֟��IҟPp^wR�'��IZ�<{D�Ц��ҎR7G$���X�dG@f�bKT;OxU��	9��|QC'���0d6�8�����i`��E:7��˓?"��	)"�#NKK�Iw � ����I����?��	\�ln��l�v�ؐ�-IO��C��Q�x���gO);��DA3��BZ���'c��(0�ڴ�?����d�K��3�ߕ%mV4��5�?q2�<�?1��?F����}����V����D�U�>��!���0�8���"�7҈O���g�T�d���HҒ��E�V18ndx�؏5�z%�Ǭ=�|�pJ��(O���q�'9|7��r�S�. �=Ba`3y(���eƙ]�>���O�����O���K�Jѹ��[��b�he�O��hO�ɉt}Rh���(���x�vA�6���t�	������8�	䟼��퟈�'�Ҹ�i�97C�[��֟^��;p�'�ў|��ZM�%녯�#N�4E�g����$�8�w�ɍղ�9P�͔"�xDXD^2=h�	��~�&����|�6l<<��)ߑ�`�������rR��&���~��I�|��Fl�O4�`���F�������-��� #�i��Q?q��9O 0��9$.��; *!����w�\P��V[�A�D�Op�Ou�i�(M�h�竎:#
���<�du�O(��S�93&`�g��;�\����_1�r�ɗx�D�'j��'���J����4=��u�������
;"��'�n8{L�����W�CI|�!��y���@�)�h���>�"1�O�s� (#?AR�ŵo���Δ��R�p`�N?`	X\�(OV8B%c�O �䃘�H�J��w	M�tJ|8����de����'��8� �-��9O���OPP�,�v�<(0S�y'x�e�'�L���	7FP�YkU�ξV�6p����S�B�	Pv=�хI���ݜo3�i�q"~��$�O�˓��Q�D�'.����+b�+� �%oL��f��8���C��L����Z�_@H��E9omx�:0��Y�!�䁐y�RR���$�2(��;�!�DE�#�&����:k�����AJ�N�!�D�&��z0�!Rv����D<�!�d}u�����&-�(8��̃e�!�$ ;<2��2�8�SA�5!򄚃'%��6�;?�T�ᢩE�!��p|^`��t���Y7T!��
p��#p ��[쬔�p[iS!�$�=iF-²J�G�N��@'+sK!�dپ@_` Q�@ٹ�D!�u�2&b�OTL�C��ȟ������	l)�/>D
@�"O�|b2��94��D��Ku=�d��$�:�,�ڂ��3������+H+���L�#��8Av鎇	<9q����ch �c@�(r��(��A�I$��Ƈ_ 0��Q��생%a�0���_�U�é2F��	d�S3k�ĂCc��"���ۥVe��56/�x�ÕP����+Z}6P�0eǹ��E_��3��USGЌ�N�\��ȓ]$� ��L�ny8%�0�͌z��}��k�pMc�B w���"��'�Q���J�  ��H��	�1�--���\���1� _zz��C
���6���x�a�#L�'F��T[ A��
����MР��3���,�}(��Þ?�B�ȓTm�-���'H�h�З���}1�5��X�j�"���h(�J� n:�ЄȓF�m Q��W��`���Y�n$�ȓ!���T�2!�`�3k��TY���e��S�G1+z&���#Ĕ')ⱆ���:��L()`$���`eja��S�? v% c
�;$p��ڼ0��`�"O|�z��#8�6��#j;/֍�"O������V�p=a�G %�$�W"OR9(5�ڂ5����oZ�i���"OZTs�̛e�t9C �)�"OIvj�2:0$Ŋ�O�s6u��"Of؃��AC��R��7��,�6"O:�"p S.RA����-VZ�dR�"OfU�%��TR\�"pK�;t"O<���,�pM9r����$��"O>��m2R��I�i�5w�<U('"O���Ak�D�`�C��\=Oޔ�0�"O2��C��H��� ��)���)�"O8�:f�l�9��Ϡ8��Q�"O@PjN
e>Ze�&��P�"$�a"O hr5F"$Wp�@��
5P`��"O�,�wJ��8�!&h�,
����"O��
0j��&J���a��j��)i�"O%��E�gcb�"�
5<爝J"O�l�6�Z�c9����U=cʹ�U"O�xR���D��a�ǧ��D��"O���0�J	�;�P(rl�R�"O��ڕ��S�(�T Խm���q"O����z��Q��i� g"O*��,�G�$p�/��B�@"O�qq#ْr\>�Ca���o͂�b"Ov9H3�K��0A�v�׉Gj*���"Oh�%䃿ͺ9C�Ɔ8JpV"O��	�tlP+��	�Ԁ�"O&�`, p��iT�8Ur�=��"OD�Ұ���S�~4�@A_�s���ZV"O��5�;j�8�Я#=����"O�3�^�vF��o�
n(�{"O�l�i�m���
ig
���"O�]iB��)	,�Ҕ�00$�A"O𸒳�Te�*q�#��Y��{�"O�@���4ܐ9��߇Ѩ��T"O
xa�F�#Y�X���ġ�\�c�"O�4cӇ��-�
}BH<���*�"O�����Ç[�EQ�̅++�!zp"O�3�T*ND�%#�k�y{vk!"Ox����#b�@��D7R$�"O�T�`���a�<]B0 �i�*a�g"O"���_�f�P�IOYL��}�"O���Ȟ065�`�d��H�%"OL��5��%W/0����	~z"��s"O�x�V��n�T䊒�֓T`�A��"O�,�����9��Ə�O�;�"O,L��d�p�](�$S�%3x)��"O�����t"``1�BG��B�"OJ鑴���Z�v!�7c�4��=
�"O(X��ٰyB��@ǬӖT����"OV�3�I;�V��c���+��)��"O6mvOX��s0�K�YC"O��0&�7V;$Ya��B�-��"F"O&�RG�٢V�Z0��a��E��@�"O*5R4a84��hQp�0���"O�40cS�nȒA �5L�<�Q"O츚q�� ��i3���8�"Oܸui�pu�[n�!n��C�"O�dzs�Y.���ΌAr�Jw"O��R$U����`,o����"O���0���y�Y`E!v\N)�"O�#ьٸCq2dz� \!O��*r"O� t ����i5�y�Ѐ|�6��&"O
t{7��' �dd�p��F��T)R"Ol��%�ؤuQ��0�%�/v�p�"O���"���*ek��d	����"O�(*�	V��j��[�x�"O" �fߚ2=���d�w����R"O�B���3}�)aUa-�p�'"OhP# g�;���@��5d��%S2"O>�������,PP���G��M� "O��Z����)6%`�-�P�F���"OY��`A)dz"Q��Ȟ@ּP��"O.̸@B�㠰��nC'_�L)��"O�a�hA=)�`"$M k"	�"O�\��.�ZD��ÂW0Y*T80�"O���s+��T�{b�f.0��""O�C�ʟ,g(SfgRC�	��"O�t8�@ [3���d4ҌpD"O�p��MǴ3@�A��L���qZ"O.aa�(�P��W�V-e|-(�"O��A�KՄ01�Ο�@_��$"O���K��9�ʹ9��E�E�ш"Oh8��F�-kH�s��*�(�!�$�Ie:]�ť��1�8x�v�P�`�!��i6����L�&���jԶXo!�dO��#��K.�"�yf��P!�$˵UW:YB�ʂ�ƺ<s�	�r-!���'���B���%�f�f
��;F!�D�+&l��ڷm�L�v1���*F!�d�1.�l!��S�/��"�+_9!�dS���� ��P(��2!�#4p�]��}�
 ��`�,tdQ�C +�`����a+��ϓh�iGL�3�"L�ȓB�@+R�
!KԉZ�L �=�*|�ȓ?�8@l�Jz<��#��|X��_^j�2��
4+�q��hחO\~!�ȓs
�%X� -Nz|� ��hJ$ �ȓ{��)R.ԫ/��I�s�zI�3'(D����X
	�T������̐���*O�)�3�کEl� �6j���ʠZ�"O�;� �x���)�/�p�Ca"O�ؐ���,Pڙ�wf72�P-pS"OZ����3}L�ҳ����� "O�B��͚oj��P�-|�D\�A"O���#�âE8i���R��0�#�"O���C�J�T\��Q8em��*e"O��9�UB�T���1l� [E"Oja3Nհ5n���e<S��j�"O^E3%D$~��\���˨O<Tё"O>\ Pf�	3��3tlW� f�{R"O	��k�
G�&!��Մz��"O��4)P6Xr,��6�W>P�U(�"O�IcM.�tB�I�.EF�h "OB���K 4�ap�L�dP���"O����G?�Z��'�N�p�@�"O�si�;y潒q�m�9�"OT|s�GO9+YD̊Se��5Q��b'"O�D�ӭ�[�R�#� VC�iJ�"O�A���o
ı$d�AM�,ؖ"OU�է�-5!ČQ�(�Y7,=92"O���wmG|�l�S�̪���xq"O��x�@!,��9��"ٝWe~	�B"Odɂ��W%l����tLƐ|���b�"O�E��	[�1�め�=WJ�4��"O����ج=��1(U�] /���҇"O� N���,�Ƅ��L˿&gn5z�"O>i�IV�\�Ҥ[�L��Kcܝ�4"Ot�i�>fL>� �AX��Ā��"O��L�Al��C�aP�w�8e��"O� Ƞ��QhV���Рi��ړ"OH��L�=�r���Ԛ4F2���"O DAk�2NxV�S�=v(����"O�EP��D�~F*
��ژ|2� W"O\�'��A��+uO̜jM�%�@"O.�Z�#Q��"�b���*B��Sb"OlM��Ț�����M�I(�yyf"O~P��-�(z7
�5�`'n%y�"O��h�/�8��us�)U#�-��"O���7�n��`C�1Z@t�a"O\�SŏK
 �ϑ����@`"O�)Z�Y</�Z"n�m���P"OB��IFRm^1]� �{V"O��q�f�5Y�F4�6���x �|Ҁ"O��F+=2B���	��|�!"O��sm^�D5��ȑ	VFPXav"O0���R��H �h
��<9�"OVŋw%ǁKc^� UǓ�/�VQ��"O�	�ghA�u|H��:�t5y"OJᣆ��S�:+Pe=��eR�"OV�!#5%�2��^�#�}($"Ol�W�6P.��c�V�u�x|2�"O��2��I�[ܐQB����ܕ�"OI�7��}�@Y�\�[�� �"O��*qjٯT��D�c�[9mŐ�"O�0bFiœ��xs��=��Y"s"Ol�`F�>i�I���=��p��"O�HĮֱ^�z�D�E�3?(0b"OV��o�u�]�����F ��b"Ol�qF�^�C,ȂO�4�q"O�KUi�;�!g�>4�hE[�"On3ҭ�n�:�Q�'�&F:許�"O���I�=�6�h�LM��8P�"O�P��a
 NV((��K�b��,��"O�M⠯���Jt�S��)uWZ$�W"O֕�C�;,�x8p�H)
>���"Ovd�U ��\�40%�^X��+�"O*X�vI��,��`sQ��x���8�"OֱXw�J5�N��2����#�_�<�sN]+ n����"@��]�6�Z�<�veِg��]j�G�!D�p[��a�<�1M��u(�JeK�{,��G%�r�<Y2�ī6zds���6	9�HDZ�<��M��=�a�1DTPQ�GH�X�<	�D6<'�؉�hL�Ia��Z@b�{�<Q6��$sfQ8�]�SN�����x�<9Q�ߍ.*��"���9;��r�<��B�v3iG��-�FT�c-�e�<���[�V�-��.L�����Bg�<I�Fփ&P8J!\������hBK�<Q��D�3�VC�%�q��`8��JJ�<aS	�@K���"�5���z&�`�<��f��T���b��Y��c'`Ds�B�N�2���X5���O�7[�'�D{t
�H�8mi^�6A �3>D���w!�Zâ �$'��#���Hl6D�Pk�`�;HQZ�sF86+���>D�Y�HF�Y�Hp�㉨9�0�C�"D��҆W��x�*�3��Pb4l D��Z��Eƈ!��]�F�k`�)D���Q��"�V�5]�^�h�1R�(D�� h���#_H�1�"�	=M¾Ր"O�uA �hViR�MK�"�xb�"O��g�p68��
��\�2�"O�`�7��C.��1�M��HP"O�\(MU�V���Y)U��Zf"O6x���&M��0�)�'Jt���"O�!!�i#�2m�Q�ȽA��A9"Ox$k�!�s���Y!R��i"O,|#1��18�橂�
�m�n���"O�X���#e�[�a&@�*O��� ��mI�M�"G�y���r	�'"����*�~��!��(Z�z�' D���˴>��90��Oq�R�'\��`�x!bE����?-���'@�I�T��[(�.	-<����'�(l��H�x�����*d	ހ��'ԘP�ˊ�o��P+�H'b8�	�''�+��l��W��:O�41�	�'p��)$������3m�w#<���'_DL��N�."��� ��U�va�
�'�N�#��ƈ-v�Q7g��g�2(
�'�
�Ơ���՛eEd�x�G�?�y�,�M����D�Mr|u���@��yb�ҷ>�:�[�-I�C��x�,��y�냉Zt<�r�șkT�e�G� �y2fe�|ة�U<� 2Em� �yRnY("����Ƣ��&�`�E�y�	�a����g�r"E���%�y�GV���4�2V�$����;�y��G�4�E�W/ޡVm���&�P��yR�^L�P��∖Q�@�p��[ �yB ��,!���Rc�V��ZPHϖ�ybd�9F3���U�J��#G^��yR�X�IJ61y%�:K�����>�y�U#J ���&�G"�pcժ���y��&�n�y�F%U�l�	e���yr��
a}����41���7�R�y�ͷW�����J�/�� �p�]*�yRn�rc���bU����� ��yb��6g*Lz��� ����!�3�y�(t�8S��F�E� #,M�y�A��YV�ra̓$}�4�:��U��y�Kʯ7���U$Δq^5[�cB��y2�`��Ӂ��5�bi���U��yB�K TX�Sd�7�a��I��y�@Y"XY�$(O
��*�y�쏒�"U�W�+p�5��A��yrmѼ�@���!ll5��b\3�yB/U	AD��V�~�H�AR��yH�@؊\A���GO�]�r��/�yr�]�s���Ae�<k�j�"Ӈ	(�y͙{�0uB� KFp�^��y2K��x���G�6w�]3ɔ��y�$�7<���#�.@i�����܋�y��W�+�.�s����s���Y%�y��(�����C9��y��A
�yr�/��e5"��-���n�/�y��T�l���ZMPy�e���y�̆
�)8�N�L$$�;�;�y�G�:u����@�5�.(���^��y�IN�^�Z�+��F�1��y{���yr(T2� ���1^��ɛ��֥�y&L(P��ÍH>`����H���y���/���K��R���p�	��y
� R)WB	�#I`[Q鉟(��x��"O���g������1I~���"O�i�'y�8���"�5&�t�!�"O���X Y&�K�a�)� ��"O�DYP@�S`��a#l���"O�qk��61.x	0G�V�d�Z�@"O^��0��%e^����%��X�r�o�<	�Jl@*���rR�����S�!�X�?��E�q��
��S�ရDu!��Ĝ{z�}Y�EǱV%Z�J$!I�*!�%_�|�����y�$�@�T�o|!�Ɠ�����=~o���,U�!��qf����鎦qX9S�C�8n!�]:'�>�b��U/st���p-S� Q!��=E�����
ۧdP�ssM]2�!�d��-�X�E�5^.d�[W�]��!�� 	 ��F��U^8�7J=�!��.&�+c�E�,�Y�� '!�d\�=]�e��,����m���F�!'!��̸]���VڒU�t���܄E!�ě!T�V}A��[66�آ�*_�3'!���V{j<r���+�Zш��5!��/Cb8��P$\�(�+/*#b!�d%X�P2�@�f�Bt�(A�sE!�$W&�0 ��@
	��U,׿B�!�ڂ9�h�p��_�i~xh���R�!�D��=`�:�#\�>a��Ꞛ?/!��#g�& ō[<pj����c /"�!�$�^�r��QL��,�4i�=p�!�dO��n�H��� eJ�	�$3�!��]�)��]	���>}��0���8�!�DLd-xz*-;�(X�Y&p��'��)Z�'k���)_e`����Vf�Y#�2VH���o�B����.!�U�i�(yF�#�'�Hl�!�J�ZQ��W!Y�2~f%#���Rbɳ֨F42�b>m��F�-�YuI\.z�N틆I%D�|x1*O nШ���	'�[F�O���J=���tJ�<E��GH6?<����/ �[�f-��-�6!�$Y��^H��IJ� A�e����d��{��e�l0t��k�ןў��v`6dh\Q�EMX�]NDCq�*�Ov8e�k��ݭb'����`��Pрk�$���(r�)�O���Â��X8��$�� \u�lPC�ɻM�h$���'M��q �A��A8�'D)\��_��HI�lܺ����N�<	��Ɯ|���Pm����p�*Y�0?h��ïڿNUV8x%�O,)�G��'Kd��������F�Ƴ���q	�'d�x��MɈ{����-Z��I	En��[Z���#I@-o�ؠ�狴�����DV��I�w-P�B�VA� �YG��{f�L �r �T>@��еb�D����$�F�z���2�/�ƨC��'��ի�M#8z<(�a�U�7\�,����f�S�,��yR���J��S�����dك=�6��Ǎ�<��C䉯'�T=��E�e|���-̲d���xF@ųZP�Y���QZ�-I�g*ڧ�y"%�&h�҄��3w��A!�y�8_�����*�Tٗ�M�]H��Ub��Iz,<s�
\�=��E��'��O��	u�K�pc�U	1�C<_�Ac�Nq|r��/$�B\a�c.O��I�A�r��� ����`�0�O���@�B<ah��11`�v��ɮ<"�٣�¥H��Ѫ�k&"@�'Iт�q�fG�0�e��;|�Ȕ�ȓ����t�֑nw��:���5W+J��'4�u����!w��X�O�>����3"�P�N�0x�S��?D�l�Ɍ]����ΨT��܀�˖���B�{#Rl�vB���3���`Jz���Z����F�����$�8�(;@�'URdl;�oM�=P@�g��j�pP	�'�Z�c[�6t!!�GSrE�d��|�'bZ�a_�6u#%�Wt�'R-k��7: 	u)׳TcVȅ�S�? (1�V�	'*�0 ����?:�*f�O8P��	�%�O�>!����#dA�K�8 S�$#�5D�8�)�)ynd��mگ+0�Q0��=�dʏk����dE".������&>�L�s@��q�!�C
��"'*O G�"�
) !�$� g�5��Y�V�4u�G8!�.U�VXBs��7zFUxN��Py������b�I~LI��y�&Sh�%Ȁ��o~D��Ѣ�y"-���:-��G�8&Ƹ��L��y�,	�`6��d�29[���DnP'�yr@�6��1:�Kê3V��T#M��y�$��>��v��1<�\���E�y��;�����U;�f�����y��˺$B��ڽ,+΍(W�Q��y��yI:QK�ϰ*������yBK�"��P��@7GB��C-υ�y�P	L8�Id(2��H6��yR��<�Ly���֕5�L1ւ�y�B��-h�)'�#5�1���y�e�#-tȴ�ξ|��}�,���yr��I�4�6��r&&�r0mL��y���*"���l��@'�M����"�y���(o'�ܢ���mH�����y�*��<ɮ-�1�Tr����oQ+�y�.V)Y����ч�����D�0�y2bD91DdK��
� ,�*êݞ�y"-חOy��)��4���d��y�f\�C�V�ˇ����Fc[�yri� ^�ǂI��E@K��y"�O�n��A�!o��;�&D��.޷�y���/���w�χ#����Ūʉ�y��Mp�X!G)��t\�R�U��y���%v#v@�dn�W�����y� ej���D5t[:��M��y�+�/[ �8I���?c(����/���y¬ǵ"N!Z���<j���c��Z��y����ڤ��.� {fD��ybÀ�,�4f��?M�́�GH��yb#�CdYC�d�
4� $�y��m�e�@e�5�<�#T7�y�A�LƉB!+�04Ϭ�z�$��y�-C�~�|e�Ą��&ܭ�WJG
�y��[`�R���h͚g�f�C]��y2��-T#P"Q�m�jPҥN��ybh��U"^�C *@�`��H�H��yb'�3rW6���$�����ƎC?�yrh�<F��1J�7�T`�i��y�l�|0�u�5k�N�j`�F3�y�JƇ?��MS�@árd�C���yR�]�(�Fq���;��a��y�I�LnӁ
V�r�PI��N�`�<���̃;�p��`�^����$BS�<Y��3V%>Y��JȞr�^Y)��Ll�<���5$��#�O�n?�0��b�<��L
�
�z�9i�"=�V��G�$D����ڪ$���fɡoSL�r��%D�PB���B)�4q��� ��.)D�|�e��<u�*x2sO�'6&@uH�(D���Cg
A��I+�����PQ�6D�(x�萱d8r�[��>D�|�ȄG0�	�x~�d�!L�f�%��2Mv�O����d��͈���Zx�`�"O&%��?���5kK@Q��"OJ�ۥ��0k�B�1vЙ4N±)A"O� jE�g	T52 4A�� Y7��  "Ox1v��}z���3D�'<�:�"O|�GDV�	X�5-:��ȴ"O�5�@H T>�Y���i�B��a"O� �%ܡI�y!҈G�
��V"O��V�e)(���G�f(6�C�"O �RG��K��3�e÷e/ 1�"O���S�E�r$>K�R��"O&�(�G�EW�U����/�Z�0"O�r"ɨZ3n�䀜�΄���*O��5`&v����'nW�l���'{�1��^�7��yI�gϥbZ���	�'�@hSR!�b����Y&�U�'kL�2SdD�#	|<��U�A�'x=XpO̶���Ł��D��'�&��v$ۛ4b�ɀ��E$d5��'C�H"Cd��jYõ�
kU\���'}����)����J��c��)X�'�4��b��F��hSd�`�J�H	�'��`�ӷӢ-�2G6[��1��'�|����.��Q��5N��hX�'u� �C�E�\!X�_2L�hZ�'��`o]1�~�B�ؚ>OR�J�'���� �i�l#u�-/[&��	�'x.�[%�>��-��i҉*�t��'
i������Y����"4r��'�,�rWb�	[��ؑ�/ڦ���'��l�vO��y�XQ�.�*�L��'��`����B$�i�m�!s��)	�'�^����:{��QʄaO�g�ꐉ�'��BIǐ.ʦ�b�W	)�B�9�'TB���
��2ec[8&<���'T���&>�p å�R!�����'����=_�iФaԅZ�e�	�'��D���/f��m�#�O�>�s	�'�t͛ ��q��xS
@�x{�AI	�'X��jd��n�����F�:�L)P	�'�`��&�'--�cuK[]k�@q�'S
���w �ʴIM�S�H���'��1����(S���-�K�����'����	5{�i��"�@��'d�;eiю�����I�X��'!��0F��P�T��_�!"8��'Ƣ���$��D��o�%r�'O��n��a��C��á7��K
�'U�1`Ą�9@��{6E 9�L��'�����Y�KnTl{�	H���'��5����8]�n��n��U� %:�'Y�t�4j��e��L�r.�0Su
���'�c��s���3B]���2	�'Tԙ $�c�F!��y�ʀ��'���[���)�j�K� B�lQ*l��'����� �<�y���P�,�[�'�x\�f�'�@�iP�G~j0��'�FHH�L�K�-��f�'�Xة�'�h�����4l�`D�N�=��'08��K�S@2��D��:�%��'C���Ў�Kaf��UA#HaA�'tT$�'�3����X47q�4;�'Tt�l�/\����F��6�C
�'�����`K�R|��VW#(�$��	�'����b�i�8�iA�1z��x	�'=���&��J�h��*
{�� 	�'�f�wP/dHeA�+* �>����� �У7K�$'�}�ï�/_�V��"O
ix�k٠5�`����Q6a�FyP5"O����㏢2�
ȨvNţ-��P�"O�Q�RNX�$ ��a-��kz�ñ"Oy@��.�&$�1숮_�d1�"OM� ���}:z%�����8��`C�"OI;Wiպ-�֥Ҡ�C9� At"O�1:"��W��I��g��q��`"O����&�)��)u`�"�4]�U"O갚���W�R��U2>���"O�� W����Mے�k�՚0"O�٨���a)Ġ6���1���¶"O�8��/B^Lrdk)H�/�Q�"O�]�B�[1/�Ȅ�RG��U6�!�"Ob0J ��858DHAA�x"���%"O6@���U.H�䰁� Q=+�%��"O��JKh6D�B �6(�P"O0��6��z��c���@> �T"OH5Rs���g��D���;U�Hxi�"OV��d���l�}�ӤN7ⲩ['"On�*$��:�N`Т�j1a"O��˄�@�uv	2�է*o"=A"O&�bs�W3W��T�u��C�`i�q"OV�@GjG&��3͝$(��Uc'"Ov��!��$�� ��q����"O0��d�"z�ԉc�k���"O0%�$ċ���y��ԯj�v$#`"O2�㖴)���Dֹv�F��q"O��i���(`�l1���s�6�S$"OFmZ
��yC*H�b�v���("Ob���#B�E�=i���j����'��|����/z�(Y �1�r���'���s
A�D5@`jR�I60x�P��'�Y� �$4u��D�_u*�H�' eؓl�$���]P-���':��˗��;�DR�H��,1�'����7aݙ"�Z�`@��
2�4��'%jY iJD�@����$~)�1��'D$��a�L���G���z�JAy�'�ph6GRfv��g%�2B��l
�'abٱuA�*N=��jG3m�A�	�'h���D�Թl�Xa�0#қ&�^(�ȓF+�Y�����5 �H v2�фȓSL�ى�ែ?�0��'ߤ`Q(Q��7`0Б$N@%9�ē�@'-Q6 ��d�bEx"gɴ"��(����}�X`�ȓ��S$j]>:�8(��&y���ȓ� PIs�ևe�V�?]�(�Ze"O@�:�%PF����-L|A�̒7"O���c@<���f1	V`8&"O��ާ5�%H��ئc��$��"O&Q2��'[p��-;l�����"O���f꙲>������Om�Y�"O.��l��<rLH�R�����"O�]z�G GF��/�;N&c񞟈D{��	ͼ�P�CG��cѤ[��Y
D�!�\�h(N<:��6q�.�[���X�!�F��`��f�T���B�W�!�$�?'R�d���4 �LY��؉I�!�$\k�9��HA.vpn��#iT!�O�z�F@p��N6kM��t-�d�!�D�7y����39@Xp�D*Q>0�!�#PPT���i���*��Q�!�O�m�⁓��K l��	�Șq�!�� 6!:��آ*�r���Z$w����c"O�d�@>Jv�ɚpG�4� ��"O�5B��	|��E���W�K��0�"O�e��#�<[G̼2��+*��,9u"O8Ii��1��I�$&��y����"O*�`�LK�vD`��"�V�(�P9�$"O4ѓs�#>����f�+K-�4Ђ"Ov,ۃq�����Gtq��#"O2��L��	��J��̾_ol�P"O�r��_&m��L�䚊X��8"O>�xCGV���@z�)UW��x"O6 A$m(`B] q E�<��	b"O^d���	$P���̌$|6F��"O`��ŀ) al�B#�SF <�&"Oy3RbS�b��h�C[�F�x��"Ol"^0 Oh�pL:*�P3g"O��r�L�>��>h<m[�"ONd҄'S'a��,;�*�:k8Y� "O4��a��9�ʠ��KE�6�b1"Oq3�+�d��ey�� �"�bS"Ot�р.,	���	Y���	�'�"e���̳E�@�#��iɜ���'�2�3������H�[�̩	�'ӌI���Eژ�JK�LC���
�'6 ��bژr��y`�&KC��
�'b�ba��0H�Ь�gL)�	�'b9h��֬ [����Pz��	�'i�ȃ5)�y~ �D�H�ltB	�'�]���S�=l��ig9���{�'w&�Q!\�Z�|i��(ѐ8�$��'�88��I�R�	2d`B1ec��Y�'� ��d��[��l
�N5Q�'v��"
�zzP�ل�oX�	�'3���&"B�a���eX��N}!	�'�I���#��103M��\L:�'�D9���1~��IX�o��V2DQ�'���4Ε4�����K����'���jV�ܥ �>�qq��>�N���',V�i���w�VL� �Llj�'X,
3F���N��2��BQ���'��l �Y�rӀ9Y3
M�AXq��'� �c�U?\E�T�1��94Df���'Z����G�e�<���*y��ʓw{<��ӁۼeoNa�V�K+r��m�.���_" !��A���E&ͅ�pjp�FHǹ(TH�1��GE )�ȓe��U�F�=�J�q�K�Zb���ȓd�b����E�_���քVe8��ȓ[�(�0c'�"&�4�@摾����/�qA�n�*9�2$��eM�p�d�ȓF����Jp�Xzԉ$�:���k� �"���O4��s��ܺAvЁ�ȓ:�t5�í]�O����!�F�����T��L��"�#BD��c۱c�P ��[�m8�O�,cζ��uAˢ+�M�\���l �5��ثC��o�VP���>#q'�U�1�oR���|�Vi;���T��Kd-H1Qm�ȓX;������v���#�Oȇ]�ȩ��उPJ�*S˰��ȋP@��ȓ6�(�g�w$�e�6�A Fw���s@D*��i�(I�V�Ͼ_Gh���d^����eL
&��:q��0l9�ȓb@҄��Ȍ"$m&̪�ˌ�E^�u��S�? L����TX)F��,O�r���"O4����֢\x�*t��7ZH�� "OЍ�u(�J�<P�iٕ?N��"OnE{�oʸn�4]���4���;�*O�բB+
�(ꐸ EHx�a)�'��qHp�Z�:g��1�J�a��}@�'lܺ��O�\C�`��a�#(���'�L�k�F��%}� ���@�%֥��'�6���[�-!r���){�= �'��a �W� 2`Q�p��$%�^�S�'"�qQrkC)��@����
##f��'ccŧ��M�D|"CLճD���'W*0����R��y�����=0�'
.I�F��4Rt`;��G���'V�bq��)(c�@Ad�	-��'W�D�Uc�-Q�*�� H�lg�PZ�'��6�n J�*�r`���M	=�yr��2�2�	�B�U3�;W�"�yB�,�z�ٰOE�d� lS��6�y�l�#&���M�~Vѫ5lK/�y�Ҵnr,��lA�oV� á��y��*����WE+�j%q��ڢ�y��W(R�:D(�+�	h�h@�j�y���%�R0�� ��~9D�q,D?�yB`ƶLl�ѣwK�3���ٝ�y�c˴h�H8Se��~0�Xr2-Ύ�y���Z��-�T+u�`�V���y�+"9�h����9j��}��ق�y�!�nj6�ْ�c����� ֣�y����/�������[��ؙd�P�y���kd��:C㝟O
^p�ëL��y�	I�h ����*\��.C���y��_��Y��!�=F�-�`Q��yR�U�b(Vތe��
F�f?�C�I23��+�D{��qA&P�D#�C�Ic<��)4m�91u��'m/\�C�ɗ|�F���G���dB�/�=�\C�I$ v<��K?��0��|��C�J����iE9\(dX"�cQ�RW�C䉣(�YPf~$l���	Xj�C䉤��IA�HǊ�$�S	<MB䉜`�ʭ:E��>3l�dR�lNB�I
غ���bv�ݙ�nN�?��C�	$���J��0����lN(N��B䉓-VX��ՎN$e��h�J����B�*5�U��7ܰX�J�C�I U�%9c�ߐ(0e'ƙM��B�	Gk�<`UF�-?p``��H$U��B�ɇ"jx�)fM�<2��ƽ��B�I�L�k��ύI� D#�M��z�~B䉧A�ƈA��L�$N�i�(H�m��B�	�uT.q��j�l�f���0d�fC�	��r���S�R,����;�B䉆pޮ1���J1+���bB�z�	�'���r��{q��8@(�X;�с�'\r�) 5M�&�&,T'��	�'͆�pa��*Ҋ��!�[��n��'Y���	VH
��~t��'
:�`�KC�~��1���z�e(�'z���ܳ<�x��O��iQ�'=�գ j�Ħ�ǌ�-x�ޑ�	�'�.EP�� %$V�AgK�>v|j0�'�����*^�Zmz)`�i��h�'��Ѡ������2��^g� ���S�? R�AJ���kƃA'l9�"O��a�E&8SlA5T��0#"O�}AvP���� �?I��<ѓ"Of���)�m��U�P��O���g"O�Tå&U47�
D�q�^�$�J��"O� �aH���`	��� �"O>(kEY�k#fmU���oyV��#"O�9 ��0/�t0R��B�P"O0;��Z#$}n�z�T"c�H�(6"Ot`U��[�H���,�%�0 �v"Oص�5'�':4F4���B�g�n�A�"OJ�����_x��k�ϒo�$��*O|l�'dA�YV*�����J�x�'K�d���F.Q�~(Y@��E��'��R�
�E�P�r����+��U�'�R�`�K�<n �Ah���wڰ���'�$�I���D*���$�n� �']p�[�=�!IL/LfD��'��e�a�2o�l ��.ڛ
�Z`�
�'�D�0%b�Rz�{���	�6H��'�f���^�o�jܐ��Em�<J�':��d�H�M(�IЄj�����'0Ĝ#���h��Tb�4�0�'�̀���p�,Iv�R�U����'o 0cG>pW,�l��7)h���''4hhb�ԛ
g2����\�[�zZ�'��@����>��x��޴b�D���'&�SEM) V�22��$���c�'>az���>�H�`�
�1��'4�@B�"�)<���!�-�(��`�'����&'O��H� /�����'\�I�uh��U��I9���|�\���'��8Q�ޢ^~ɠE-׋|h쀓�'Ӯ� �$�wsE85	ϒq|�!��'�T�![.Z��@K�Q�l��1�'T
�:�d[i�� ���^��1
�'�t �7�I>�@ "�*Y��� 
�'W�}㖇�%<�
P�Ti
,W怤�	�'��*�!��B�(D���!:"��'Ò����S��壳�����ȑ�'�̰��ޏ_��"�� s���'L�LKV��$��h`�O,t*\-��'��1Ʉ�D/K�&5S��p)��
�'���p�U���s�[a0zT��'�����p��ۆ� �SJ�9�'0hY��	A�=�1��.��q�(D�P0��#L���Rjݽ	jH�	4�%D�hp��ĴU�:0�fJE(C�?D�P��/̯Y�����J	%> �4!D��@��K�hbĨ"��D�<�Q�$�=D��S`�� �����Ĭ~Z�A��<D�`d�01��x'�ޅ`<�e���8D�����k"�mْd
a���C�5D����<P�֠���� �����0D�D�����c�`|	4�[���Q��-D��CWK��X'�)�*�&*�d�JS/+D��q'�'/&Ƙ�e�ӳh[XLcG�4D��u ϶X��&��3`<t0��.D��J���2g�1A%�C-9��f,D�x��H$ ��˒��*&��;7m<D��ȱ�D>8^9{�j,Ժ��f>D�����ϗ�dI�L_5,�nl�1�=D��U��D�a�A_�)E��R�&8D��УQ�n��d�JA(�y��5D�� ��Y���]r�*�HC�;
.m�"O@���xNV5��G�T��jv"O4U����|�"͒2bȎY��QZ�"O�q� ���a��Ԡ:���Q�"O`l��B�W���~�j���"O�Lq��4"0$�2G�[w��U"O21x��X�t@���Vr��#�"OFɸ"L����D@�LWV�00"O�ܒ��A�V����;����R"OhE���?��`{����f"Of�q��.�J�3䍌�d��5"O�E)�e԰;/4%�5�,z�;w"Oܜq�Β�\e��En��=��aKs"O��d�ڤwX��Bm��=""O$�B���+a���l����`Z�"O�0�V <U<�=����~�"�"�"O)ʲJ��~�q"Ձ�F����"O���	�ZjX�R��&a��в"Oz��EY����!�K����R�"O�p�bţ%4f9��n�)�\�C�"ODZ�f�5�૵K'u��R"OVDҗ��&`�`i�f��/���"O�x��6�D!�ə�")f዁"O��FF�(>@1�2�o	��F�ybÏk� �j��C�-2܉y .\*�y2Ynf�0�	�"u��\[����y�O�ri�EKU�+q�l������y"i�{�@s"�v6U��M:�y"�ǌ
K���'	��;�T�:����y"�e�\��`"ǉ;r��"��#�y򀊱�JdK���	i0v-
�Λ��y�6O
FM��J��2�:p��'�9*�AB+1�&E�3��'��� �'l��2�oJ
6v8z�C��vB���'��y�PF�V���y� VN`+
�'1P@cm��aLpI�^k�IK	�'�(((჌?�"]b��_].j�	�'�p5Qg��-B�s�G�=����'��Y��X�	_��h�Ë�)$֘*�'`��wh˂y�j�s�o]".+��'�N��oWg8��,ΩR]���'n �ST�T�%-\4�$�����ȑ�yB�xh 8A�"?+��#�:�y"�׈z>�u ��Ѧ5���{���-�yb��=��D��J�0O��ڑ��=�y�K�ɬy�"aVj��'T��y" F"i�ح�Ӥ߾]�,���D�y��H�`��6�N�A��p�>�yª[�c����R@(Θ���/�y���pz,�i�
=�\��`'���y��������?,�b�)�h�y�����f���g�B	�y�J�'�����d&���`֘�y�b�J�)0��;rF�,��y�K� }[(ԡ�k����J��O��y�h�8��i؅*Ҷ{�4A���y¢R?p!sB(R�)"8�!�E�y��Q��S��Z�&϶<�E�
��y�
v+��b�C��6���m�("�!�D�����
��`T�q��J�1zp!�ɂ2g���Ņ�Z`�pf		fe!�䄹]�6���2��Q˱��0f!�Dܱ �jY[@��%�����AL�!��>Z&(��aGlv���<�!�� �Yg$J�,��)�+�G��!�"O�r���HJ�x�܌��LJ�'} ��6�E�qt�5�ti�'�NUq	�'|zh����/:0p��GT8�@j	�'�L�C�^����i�Q��z���O8Q��D�M��t**\�VH�G�0%��xs�!L���'v��%d��a���	��!`��6TE�' �tm�V"�A�P��$�P_&|FzBt����(x�f
��8d�)� V&��
��wʶ���gW?�������O�o��MK���)��X�D	�^�Z�����$� \�l�	_y2V�"~�I2w��Su�Ҥn6Q����3���d|���m�����݅|e�Q�.2j�{`�� �!�2��d�I`y�O��6�+�d]�s�0ȋ5/�t�1�kC~c����+N&j��A `F��T�$�D�q�`��w���;��5 ��dCoLR���ڴ^K�H��S�V"�S윣m?d��4�s�i��^|�$�3tf�E�8�&d� ���'gLk���&:J~nZ1+�\3�e�4���Kb�V��ğ���@�hʘo��p#���2CJ�<�D�i�F7-,����]�sb�x��Z�l�5��O?S�Ht+O���������	�+�
�Aa��9Q�4�!A�S*V`�X���� �4=Jv�O�3��-c���JQ�>�	������hi��K��JT� i~�z��aW�]{Z����M���ɱ{�, ��Hb��1h�6�4���;��Y���?YVJ�~�'���'ě&29�\�!�L�rc�)�ꛭpa�C�14Kj�XЌ�ʄ�`�L">��cC�i1�7� �D���<�6���3Cj�u܂�.pir ��[贕�Tǌ/��<a�[�vE �a��p�
� L�ִ�	�:�lY6��8��賂k�CD"?��ƫqD�@�?��5��BZ�(�$�$B�mR�}KCS�XNLa��I �d b� @cThX�/(����B�d�a8��%�ICy��'��	F�'%$ ����"V�$�W�2v�ɅȓJ͖P��H�v�h�铭P����e��bv�$ʓR�L��i 2����5yB:�x���4�ar�`��¸'�"�Q�X&tu����}�p��c��3>zB��'u�tY'L��x�n$B�~�Ez�'��PIT�2CΓ|#��0��\;f?4�S �T	ɦ�-�~�q!a#��"=9�&�џl��43����'J���@=�%j�3},jUZwD@;_5Mq�����O�rZ�������,��&-����t�0�O� n�M�4.b�̉&o�-�,��$B�-�(4�"�i�$�U×�)�I�����?=��hџ������ps�n�����/�
f�4AЖ\�?�(���FN�8$͓�?�+���gy���vyJ萳��	.�J�0�l{)o#B�T9��N��H�j_b����D �bP)I|�1O^xU�!B��{�.�S�ɛ<�H9oZ/J1����Oȱm��`E�ܴI���q�*-���*R��l0���?)����'ֱO���-ЮY/�\9�@�be��H��		�M��i��~�v���N��1H��W@�L��b� �x�)O>��*SH5�  @�?h[��1���s"O�Ԋ��;^&�)&j
[c
�"O��y�a�,z����a*�^�>#!"OܠT+J�z�h��qlN�~��(��"O�Њ�Ꜫvn�L�ТB z#Y�"O�|��i2X�A�aF|X��"O� �l�9�,�1�?Z�Rd�$"O��R�f/6��$kۖa� )Ѡ"O���&���Xѐ�U2!���:W"Oة�#GاG��h"�|���ق"O��)�ޥ ���B���c�Ba�"OdXاό�$�ā�	��*�ԩ�p"O��5-�9�|E(�ƚ
YJ� �c"OB��3T\
 ��$K,h5���%"O����&�9��9��#�9C"8dq�"O2I���Is��s̴P"OԨ鲃������"���x$"O��r��;, H��c�DU�ă"OK�a*Zq�#/n���� ]��y�i�n/�DZ�S7'ڑY��Y �y��:k����k�3ޠH f�P��y2F�f��;	G��H�O���yR�э!�D1�qnQH���P�*��yB�Q(7*`5����=RI��O��y�Ńh��,2�ٞ0��E�`×�yro�5D�&�Ht�ɂ3�n�;��Z��yr��8"��;���,����0A�,�y�e�8zn�P+��$�vQ����yBQ����+��+h4a��!�y���"�$��0-�2 ;����/�y2.�����U�L�Nd8���-�yb�U4pZ�h�e�,2�.06�X#�y��݀`�$% tK���@I�����y��Z'���a"��e1�4CUi,�y�
�p�,!����`��\A��M���p���0?�6H(�(9�
*oҎ�[FX�<٦N�7�B�ՈO,7@�:���[�<)��.D����ǝ[���ɷ��p�<I+�Rv��q�J�
q�3T�^�O���a�L�T�1Oq����b�7E����n+Y�hUS�x2׃[:U�b��|����c�F�
S��3pHrhx0$ʟ41N�-0T�b��~��*W!(r�kAl�'=q���c�{�p�W>�?�W����Y�wj��"���}�j2�'�UpG��)L��ǩV�CzyX�ޟ|"}�D
P�"�t�c���$a_�a
pd�2I��!�mG;�H�Z& FT)�ᓡ}�. Z�ǝY2\q��^�<2���"e~ލ؀��'����3C*��|)�a̞� ��/ߛٲ���n�r��Q.бJ���+����~rK|R" ni�1iŇ1��:���'�- ��Đ��#��s��nځ'�hQ��B���Sf�[�p�BC+�%[c�n}P��4&�����P� -��2�J|"d�+&�v�yp��0W:�P0��K�;a�v(�?�~�u�ؔb�^4���T�T���u�n�<9�.�b�x�(��O*�AvkE�<!�� C(�8��N��� R���<���s@b໗��5+��q�sn�w�<	�,�Y�m�d.X�%�0'��|�<�7׻!}���"���)06n�{�'�ayҥ�&L��qB�".�<�`�F�yR��#v`i��O�����&U��y
� "���o��/xc�O����p"O��2�[�t*��0���"ª�� "O�D2�	;Q
թd���dИ4"O$�/�
�̑��/ζ1�v� �"O|q�g#]0_[�:�]��)"O��!�(F"W���k�Z4��Aw"O0đfI+ؖE�L��-���	�';ܸyb��~m8!g $
�Z0�
�'�d�rp'�=	e4�Q%ƺ5�f=�	�'����ԃ� �pd]0x��	�'��ȪT/�<�D�G'�&E*dy�'M ��!=�.9j@
AVt` �'�P(���=z���,[�;��Y��':�"���2�&߃�f���'�j��A�RX"`��� i��h��'O\ &BY���cv��_ٖ�j�'Ӧ��Ă�F�
�{�+�6']8��'�0�c�gە:���1b/�Hl*�',�C���8�.e3�Q�n��\�
�'���`�  |*���I�gC����'��x+�+n´s�ūe�Ly��'����D4
�$9ҭ�d^����'%�(�)E�fg%h��*R(03�'��q�Q ����12���U��x	�'tl�)e��r\�IZ�焒<�X��'�R���I�=����Td��&XZ]��'��
֣H1���#.�q� �8�'!��
G		�p�2��V,�?p�BU#�'���E��'<�ZR�/˚k���
�'�is�
:$�آl�v�(u�'JDC*۞(��ic�G�=K��I�'R�%���Β)�K��F).F���'�ܝ�r΋�Mb��̅�TRL��'SD .�+_�u��ʘ"���s�'����΅od: \%��� �'mZY��τ�}Ku�ׁVJ��TZ	�'7"��c㓕gK�`�%��1����'#6esW��+�)�(9 j���'����e� �
9�#�A=eRܨ�'*�e�tˀ�
�|سm���s�'�`<Z��8���hАY�l�X�'l4��Fd[��X��cD��>	����'>&�(�eN+G�*܋$��2u��B�'?$��UF�$\�����"̖1��'�BYز������Oθ_����'\&�0��,<��+�(̇c�h���'v��D���I��R�Ckx +�'����bΑ�_���R��<��]��'pl�����K�h9�2�����'A��PEB]:>\�1l��,V��Q�'�ι�Bƾy1�諁E�(��l8�'Ed�2 ���hJ��+1A��!�L��'v.�B���>(>J��&¦���"Oxp���ʦA�IbKA]����"Ot��C�A�1�<�I���u���"O�xђ&�+k�%a&i�g�B��&"O�a3��7���I�!F���;t"OI�ĉ�*�jl9t��:��l "Oځ�B,٦�A���n$>%c�"O܁�%��qn��5I<7��"O�TY&Ꜻ4��d���˂F��y�e"O�xxv���6ێ�k2k�=*��E�#"O��Hv�K6�>\��N�c�,p�"O����P�z~�A5���M��dj�"O� 4�"��[�i�4�&�. l�"OP8hDd�?�9�O�5_��`�"O�Da��8Ը�C��Hw��#"O�I�N@�t����kȐo��y3�"O�E�����H|��*ڠ � �"OV���
��s�,ATI�g�`�S�"O���S�%��h�gѤ{Z>00�"O��y��o�����>@EXk�"O�E�s"]�([��ɡ� "qc*O��s_ W�����"؍����'�0%8���` �H�܋6�i��'a���Eg�4I4z��&�>�a��'y�h�a _DsB-*�_ 0)T�A�'�ν���f�p��*�"3��[�'^F���ɻg�Y�	�(JvH��
�'S�iJV�S�gs���wE;-��	�'^U���k�Ʃf��,���'�V�RD�7>tHh��N%2����'�J���Hh����e�[>��QY�'�yRu�J�U|0ar(�g~�*�'T��B ��7gw���NS���x�	�'��QK �˜��}P��)B���'v�PYgb%R�����P��ZQ+�'>z���-�'Q(�� ���)�$M�'B�3'W�:1�������$@u��'4�Tk`ᒾ;�VD��͑���'iHB�J&&\ִ�qŉ;Zp���'��\	1�J�7.�iP�۷@5|���'�d-k�c�J�|���Ꮑ$�j�	�'@ 1p@Y#Z�tE*2)07�H�'DD��"L3k��c\)�\�#�'2P���L�Y����P�k�H\�'�\\��Haq�pR����O��)1�'�Ra�FK5V�@��U*S&TX4�Z�'C:LB�a�6��8��Ҙth�{
�'�0,2�b[^h���#J9f��@��'V@0��^�w�UIr��>_��x�'8��u
��ʝQ�X;%~P-a�'`F�K�..-<� �JR����'K�!����i%�ɐ��
G \��']�E�M F�)agNs��H�'�&�!b	5��u�.	,.�=h	�'��f�P`R �+��׈��P�'t�غ'4x45��_�t�(��'�*\�qM\7Z.�$���_H@�X�'��bF��t��#��4p�  �'�(�!��yΈ�C3g:1��
�'P�hQ�ES#�$����a�S
�'|����΅�H��c��X��B
�'���x��#3�� K��-S�Xc	�'(4usD��i�hLJr�ʩP���1	�'����$ O�\/�R��K�~�0	�'%ح�uFYY��0��`��q�1	�'�,�C�7ѢX�Ѡ��y� ��'� ��)�#V�<,jBJ���P�'���"�^��N$�� ]� Dy�'�)��&�tuAL�T�"�P�'J�ȉdEؑ4�Zp���Y�PX�(r
�'�ie-���0�I"�D�' ~���a)y�AAR��<Y�t��'b��$��0!f��
�1��P��'��%X'îD�2�b 
<��C�'��m��?0�.Y�4�P1$���'�<�{�U���%E#�p���� ة�)+�hHh�hZR�,���"Ox [��;:���n��#����"Ȏi�	�4rz4�4 P6G�DA'"O��6��>iܙkV/̙{��=�c"O���Ǐ��9I�eYc�]1*����"Oj����_!:������O�8�b�B%"O]�V�04Y�fs�8�h�"O�%!Re��9=x|����B�L��"O��CD͝Mm,*EHn��C�"O��Q�'Y-F�r�#�v��aT"O&�Q�H�'?dJ�Ȑb 0R�A�T"O�l�d�4��S��&T�4hA�"OP=!��̱a�b���/ܒ|���H"O�4�����V�ǉ"w��A"O@���G^�X�ˬ-QT%�S"O�m�	�=��`����?D;r�Q�"O<Y�KQ��sd�a
&a>D�$����%ݚ ʠ@�[��U���<D�HS��
+�؁bÌ�#"\Q*PK0D�ЉC,�5aBP�#K�Q���"��1D��`1Ĝ�;XIJw.Ԣ\�:y���/D�("uAM�rD�JR3b{
qQ�1D�TX��Ю ^E3C��/:M�3��1D��b��/���e+��E��yC�0D�0:��eh���C�W$p��Z��!D�8Ƀ�ȇL�ΈD�V4|����W�,D�0H� q��J��
H���q�&D� A0�d�q�a���:r*&D�q��-?Vձ���?1JX|b2�)D�k�Ê�1^��r�W
F�R�	D�%D���2���p�q�wb�q�bm��1D���v��r)�yp�X�^��ƃ4D���EbP.����l�=FԬ	�=D�L+��/*�ۖ ��`��ɘ�):D��NǦV�Rԃ���7�p=� l8D����Q���P !����1D�4��͝18$�a��):�����-D��"���/b�y�q�KD�ΐz��+D�<��E�u��i�T�Ţ;�I�,D�py�K=Y�� ��ĕ|�l�Sn D�����|�0BO	,ۨ�� )D�|���	tOʌ˷� 1-�`�Xѩ<D��r.��t,����fB��b��s�<D��1������@:��@k��:D�����$:�$�0L�7nd�6�:D�P����,v|^�3u��r+,�K 9D�@��o�)q�����W��4�"�d!D���!mɂ	����'%
$0q� D�4��ݡ`�V	�`�Ӝ}�8%�!D� �2�	�d|Tإ�*��n?D��0�(�1keT,Ҳ`B�>a+=D�����$&���Z�Ϛ@"��H;D��KK9T�Yp�H��pr�!��i;D�����>k?ܘ�˃j��A'/D�$*FD����x5fBNd)�g-D��ZL-����u@U^LV����/D��3�+4u���@cK�j��� �a#D��� ԱS�Fe�GΉG��hp`#D� qc�j���p�J��Ĥ��!D�ԃ!"�R"|��I,윤!��;D�"�O�>5�\�C�H�n�j�9�D?D�TJ�k�T���Z��D�T$�l�J?D� iP
G�+KޭZ��Fk�䨈d=D�2g�ZQ����I27 ���`�<D�� 8�t↵=��4�]=D#��Ї"OpMZg�K3?�<� ߖU8�$�"O�����AQ"�$�Y�|��͘V"O���F(d�f`b"��eZth*�"O2��e@
�VJ��u��0*�Xu"O� �Ï��|�m�v��4ta�"O�L�%	   �*ot��R�Tږ���'�n��-��Y!a9>�T!�G��6U�@�Is�t�b%
 e}��xk�j45.�y7lW!_� �'
6T���}��neV���q�vPp����'�pDHFM�2���ֆU��*�	wLg>�YS���k��X	��7f�����C b�p�	��&n]#V�Ϩx4��D��K��� � R�-� ��K�'�-ꄎ�7 2=�B�o�ԠY��,��'��M�R�h#��-1`X���Ҹ�|�B�36I�à� � 0��*j��`�JP�lWj���7�����e�庆e�:Ҵ9�ъ/a��pJѮi]x��S`̙6��'c氐���վ��!-"ِM��$\O@�/�tE�����m1`�;8�6�S�e�*<�����5���3.B�_�Y��N�-�|3@+��{r��40閁�V���g��AlY���'r�� �����i�LTu��
����T	�+˪����V�r� �#���N�@��aLۍZT~� wM"\OhMK��8�XR0 ��$\ikb��5jz�c ���?�"���H([A$J#hDFł��i��4۷��-���A Zk�Շ�C�I[D�1�i�1�n��	�ɴDV��� �6�E�J[J�UcT�~���vC"�i���T:W�D=;�z}�'.��"�/��M�g�a�$�e����ޤxg(�7Wp�ч@\�\�pKM�v�bEW��c?O-�ߙ2~��ë���h�Of�:V�ы*�%�4��?|�*ѹU��ac���nY�HER��ۓ'q]�0�S	R���s�X�\����		Q���/��_���i�i�0���)�\�p��><����',*��W�ܶ����m��Y�$��y�-M�\�0��"¨{��>���k�d8�pNN�|j�`$D�<�EE� ��a��R�>���Qb��[W�@��1}���E���$A(	;�hA��4� Pq҆ſ6�!� ':��*��	U>�8 2��A��CʭL����;��HCևF�6�*d�%[<C�I�-?�(�CH�+��
C��Br�B��)5TT<B��̋V�Z�a�+֗v��B䉐{&xM���J(Z�>���;0�B�1O��AP.��4��Ԁ�;.�\B�I�ҁ��խ_ 9�p.�#N
hB䉟��Q�e�]�R�����FŞB�ɐ"���sP��+��}�Q'�$.%XB�I>y]�A��"�9uW����޴`�VB�1hՀ��d�� ��Q��<@!B��&����*��v$����!�j��C䉺^f�Q0�	��φ��6_�C䉅�H�3P'�t`R�M�l��C䉰']������#��(: ��4i��B�u�q��P�2���
�̰B�	:,���O����r5`��r�B�ɂ6������X�8�����e��B�I
m�2��p��)A���4e�5)�4C䉞%7�R@H7p��tˢ�ʛo�<C��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   ��   *  �  _  �  �+  �7  �B  eN  �Y  >d  9l  �x  ��  ;�  ��  ��  7�  {�  ��  ��  >�  ��  ��  `�  ��  ��  B�  ��  ��  i�  T�  ��  W	 � �! �- = G �N U J[ B^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�?��+�сg��:�h(+a��Un$��F� U��yz�rMY(P.؁�'2Q�@BۓRLx�b54�n��'�Л�O��@k�b�P4ir��g;D���HB �𸡆㎨5�6���:D�ĉv�%ΤqQ�-׻q�頑�$D����-:*��Yg�к/F�`BR!�II���'\+��0�e�=��d{f��S%��ȓnydP��La�Fe��6E����ȓ�u��
O* ��1��@��Z���z�	�F�^ #���L��"O˭o��x޴��?a0�W}����(Y�J�65	f\�<A��%9Љ(Q�ˋS�X��"�T[�<�/P�	U-zQ��'�>�J�,US��>`Dx��$�ߦr���(�Cu�ځ�yR/�2���"P��9s��i���\�y2�֓zwB#4��4�驴M��y�)��GX�@��9c�}z�2��#�O\������j��<P׊�$Jl k �'4���y�zm��f�"� ����ݼB��	t��JA�Ȋ5be��>[�>��U�"}�'�O�	/?o�*ny G²M#�)����9���D��/r���8zn���	J�2�qO��	8��D/�T?��ӊYʊ<yF�֤f~(�*�K"�dm�H��HAUĘ�^�nQ���Ή.�C��/�f]c`�?4LY�RoH�U=�C�)� ���iP�7�e�diE;٪̰�"O����m�$����>A�<	Y"O$}@'bU�TV�ȅ�ݠ?��m��"O�K�M|��	��P%.�y����f��i��ʍ��.F�:�<Q�����<��`5 ���N����z��:o����ej��4/M�t�4���� ox�<��	c�oPL�QgA&0RdIg�J̇ȓ��i��۵O��(s�\�9D'�r��X�S�'q����g�����dXU��ȓ0���1ed�xZجX�$�f����?	�BJo���I�12u�匔�cDԻq��XZ!�Y�� C�[$�LeH��� lH\����s�����J������ځnw��Z�,D���햨J��	�k���$xP%~� ���>2`$���f_>c�`��QGzB�~r�_.�����q�T� �v�<�NP+$����5��!E�\:%�s�<q�^C;x�ʠ�� }g�z�"�e�<9��]2��<�QDTLz�$ٖ�c?I�:�؈c��@*,���5�Ǣ`�~مȓ3�^��[48E��B'�ꐅȓǫ�b�ɾhE^�X�"ܱ�X��ȓl
Y��)Y��艈AD/y����ȓ>h9bWOQ�W*��n��_�@y���+�S���ٹ_s��AvK_{�D�e�\��y�i�7Ze������ i���U�A<^�Q?i(O?��?51Ȑո2�˷�U3W�����'�p�㣋7on�Y�g� �N=��3�yB',lOޥK�Kʊn��� �n�$��O��>/&1 F�:~�������v�!�$���|DCAj�(yq�4۔#VnџxG�k�O�0J%J,��X�N^��y���!�\�����hXW�T���"�S�O��Q��wp�tB�d�>��]��'��Ȣ	�uL0Q8�e�J���	�'�R����"Kp�% ��u����'����y*�;&.ֵs7�d+듹�󌱃��$S2��3w$4$e�#>���I��*����kGm\��V-X38+!��rH	��H0.l�ы�-5$+!�Ӿn|Ω��0\Q|x�-̝�!����*P�F��U��W��hʉ'gb�Γ[��xr	F�x�1�[%fc��h��,��d'O ��y���fh��D�
T��a:f�>)9n�M؟؃��E#�\�A��T����8�ə�HO��2�7@�r{��f+,r?`цȓ3��Y�«٬/SD���D1�Fz�'�0�Y�M#�骤��~8����'��U��@����P�fO5%���y��?lO��p�≒�TYJ%D.k�h@ "O����nL�>�0�kt��=-^!x�"Ot}Q�N�EYΩq �т'J����S�On�M���R	V$���v�ٷ����'�<�e��*; ��"�}��b�'e�#B���8:��"I�̉�'�
��� ��Bc
ι
p���y"�'`����1�6�bFP�
��	�'�*嚅.�K�b����8%����' L����Do��C�>�$�Q	�'�"!���*p��Y�/УF��ո�'9p���hT 5(���Ԧ�m]�q�	�'�(��(Ǟ��=%�j��0�	�'אYд.� "�Ԅ�kՖZ74 ��}���� ���ʟ-'~��{4эB�MCp�'�'fą� Cb�����&��b��	�'/�ծS-�&Y+R ׫`6) �4�Px�L+*��P�+��_�4�&)���=эyB�T�������mB����H�oDL�<���Od%�%���9�R�U1�2#�"OpXsD�A�41���޶lʑ"O�X�P,�����"ēc��Q�K4}��>%?)�<�_rƖ��4�A���X��''"4��Hլ0.�����}���m��I�O��IM̓ڸ'�,
)]�^l�U��87��3��y%ъk�h�q��� B��(RcK#-�qO^�GzJ|�u���D
V����B��=z'�Y�ȓ0�\5�I�H6 QB����\����'��x"E�Y&���F����X?�y��F���m����*ϴ,7F��yZy��[dԷ_�b �ƿBB�C�����͑�<8,ۆ���8��C�I�#�q�hʝ;�2��`�	>ϤC�I"I�H�ѶGƌD4��z�C�.{�C�/yQl�����s܊e�&jZ�C�Ɇ,�qG��'%XL�����0~C�ɇ��}�L=!���R���C�
1�䤁6+��O����"_45iz�'�ў�?������	M�1��$uTr���H7D���sח9��B��<*5�%1D��8���i��A��&�����)D��y%�����B�+Z�s����;D���Vŝ S)e�7I׆n�~L�a�:D��"�����b��3W�-b.�`:D�dB7� �9�5/�"3g�w�8D�09$䎐_R�w�K�(;C�*D��x�'���4�`�4>o�dR�'D�����6��RHR}-���*D�T���E �mYc�Z�:64L��n(D�����X2EQ8���N��b�ap�%D��;n^�>�s�=v���A��(D�x�E��?�X��E�V�'۸�pFj<D�(�F%�r�H�vē�H�~m�G�<D� {��D!��`�GǅJ(ZU�f�;D�\��+H�G0+�LFN�*�x �$D��q��T"J���E7���!D� Ac��.f���F)¥G��$��O+D�P� °i!���#�3.�<ɡ@*D�|q����
���pE9R�t�`&-D���d���Y���2�E� ����(D�0c��FE4\� A)C�Bs��SE$D��Ҿb�m
�a8QV�ɻh=�yl�Vz���ү�8�$�:��J��y�%Ya�Aq#���J��̍��y� F�ҴBVn��1�4� �nT��yrj҇U84-)��y�����y�Ɯc�l(ʀ�M�7V�=�+Π�yRN
-��qR׃�2�>��7f���y�ḭ{��X���0�t Q����yB��U`�!� zi��'C���ybm��z�����x�BL�3�6؆� �Qk��O���'ZD���ȓ �Z��NA�I%t��*�7�b�ȓEw�$��ڷQ����󃟇8\����n�ƕ���):hЁ��e��.��ȓ+W2����0ބ�d��4�2̄ȓ�����	�%24i''D�(B&���y-�����x��*�;k�Q��S�? ��TdM�+�=�BP�(����"OL�q�O7![��Ƈ�&FB��j�"OT�ؤ��yL����P5IU"O���1��-���C哒0�2��&"Ov)�U;�@��ݏ�J��U�'�B�'(b�'/��'���'`���U�nЬr`͛��шC��Y�K�՟��������ğ��I̟�����	��H�	99�(9�WeUa�`�R��ϟ��	��Iݟ$�I�h�	����T�#מ2=�T:t�X�I�^e�3hJ͟��	����D��������$�Iٟ|����N�r��sIα���Rş����	П��Iޟ��I韘�����W�@�v05$ڊQ�е1u�ܟ���ٟ���ȟ�I����	����֟l 7EA.Qq�@�j
03T fK���X�	Ο��I֟����� �I�l�I��K���-���0"I@E����W����Iџ��	����	����	ן����D��%�&Ex�8c���൓!�
��X��՟|����	�H���H����t	sM=fE6�cƈ��~��3������՟|�I͟P��џ �Iݟ������k��J�(*~ ��P;�:�C�$�����I����I���������˟��I���.8�г@&@=U��� �!��A��������I͟��	���������Iȟ��I�v��u��+U��h��R
�u4�$���0�	џ���㟜��ß ��4�?A�0Y����R�{��0��+�R�|�q�U�l�	ny���O<m���ZD��l��x�@��=�n��a�)?AԴi��O�9O��W����; �3qB���uL��i"��D�O\T���g������l��|�O�>E��hO������-\z�qX�y��'{��c�O!d]�֢ç;���&[I�5�r�u�:!�d�$�ӧ�M�;` �x�OF!}|�`�p(V�� ���?y�'E�)擦%��YoZ�<7@�4UYn K H��(�$�,��<1�'���DN��hO�I�O$����a@(�����lnj�٧;OZ˓��}�F
�'��ѻ��@���
�O֥1x�{��YS}��'��>O��z��H@/�:+��E�ʗ����?��K=<�|����O>i�ol�����ؚ1�0H�l	�Sɘ�.O���?E��'m
� ���*$�⊓F)�'V�7m�&\��.�M���O��С3a�{��8�'gN�I�"��'S"�'gҢF�<қV����'	o�T��n<���'E�_������e_pu$����Ϙ'U<�` ��8)j��q�����Oxmړ�8�'����ȼ<FV�3�/
�g $��&�M� � 	�'�7M
˦��N<�|1��0�������#V; T����}��(�X���D��F^����dQ��O\�g�ɋ�a
��|k`�B�,�����ɖ�M��A���?'`��&�EAы�05�����<�t�i,�O�X�'�6���47�̋b��7g��<X��K]�x���"�Ms�O<u9�)E����M0�i��Dc��	�Q�:��-�09O��OT���O���O��?��� �9Zh�� 9[o�{�/���<�����Jݴc� �ϧ�?Q��i�b\�ĐD>.�0,�m<+�B�Z�G����HR���y��	� �7Mg�<�	Ip9뵆Б'�X���.Pf*����Ի_b2��x�I{y"�'r2�'�RK&��m�Ԉ��6o�(P(�F�r�'���4�M���Z�<���?y,���;�n l��fV?.��I���`�*O(�d�0c��'��!�"O�f��%��:|�(i0G��P ��3��4�TxҰi���&�D[Q�kX���@X>l�z��������Iԟ����b>E�'�h6�	u�v�R���I��	1� :���On�dU٦1�IZy��'����M+�n�9`S�<��l�h��*��F�c�`Tk�Jy�T�Iٟ��P�����gSty��:QU&؁��4"4�s���yBU�t�����	؟0�IʟH�O`����[�|��M�e�ݾe�{`�xӰ๖o�O*�d�OВ�(������]<F���Yï˴�T���C-;��EpܴIi��&����Qnݩ�4O����:ϒ���Λ=(�z?O� 9���?�� ;�D�<���?A���*Y�*���C��^����U��?a���?I����D���ma��������""B�AX�	F���d����S�j��	�oZw�I'g��/eL0<jc�#p؄ꦛ�Lx4�آs�<�5lAG�q�6���?�0� ] XѲ�n�1���#dѽ�?	��?��?����O:9���ٙ=u�0iRKK�o���C'��O8�m�)v�je��ӟ,�۴���y��4[uإ2P�VM�8[��Ų�yR/}Ӫ�n���M��%H>ݦ�'G�pJ�ƅ�?q�E�(#y���@	�\[r���
WX�'Y�	ǟ`�I�������I.f��Ӱ<h!isB�(<��'<�6�45��O��-�9O
:r��7��%GA�ԭ mJ|}�lp�2�lZ~�)�S%RP��'��(NxƠ	�a����"
Z�y�z�'7�;F����M��+?�Ģ<a�K^RȨQ��)*��q�o�*�?����?!��?����DJͦy�Eu��{�K�	��çnlv@Z�����T�ٴ���|jQS�0��48n��'<��$�K @��!�(��L
�XR��޶VD�3O�!;�)I�FH��Y�O�`�d���$��*��� �KA��^�� �� jD�	#:O����O*���O���O��$��.�aμ��'eRJ�p�fM~�����O<��ɦ�
�r�t�I:�M����򄝑_*�G��vH��� k��O�pl���M�*�0�B�4�yr�Q7z���dN';�L����#�v���gϊ{b�Dz�4>��ʓ8zV�+O��$�O����O|��h��h���Wb��+nk#��&NrnDrA��<	��iQ��`t�O�b�'3�T�wF��R 
�;�	#ъ" �H��'�ȼ>Y�i��7�6�4��SH��P�V��[�|�`�K8�:����� %|�@§>���f�}Y��g�l��-O,�:e% ܫ��є�l�d' "M����O����Ol�4�����OH�/��v�I�f1����ݽ~�p�4c�%c�c�'^�l�r�O�)Zy��i�bQ�E:\4qc�u����Tow��d�#E�R7mk������pP�~�IP7S�$��H�'��dڧ�[$r��D��C!�M)O ���O����O����O �'v�ڥ$b�76�͸�#��[��$ҥ�i"<���R�����?�s����3�Mϻr����� (����Ղ_e��)'�'���O����'!��HS�i����<@�� �T/��X!/W\��
 �%�¿i<��'[6��<���?���?P|�S���>��0�u ��?��L5~�B���d�ئ��`k����ɟl�R�`��1��$ɇ7ߪ�⧇d�	ǟ���O�,o��MCH>�D)�0K� ��V#��k�	��#_�<��O5Nerd�*?��(O2Ѭ;Rb��nZ>b��:]`6x5�^(r/�KPET�TO�'��' ����O�n���j�QD��;����"A�)�l�ݦ��r�w� �I��MO>��3�/P�TX�8�@\.c<tĸ7`�\?�ڴ%>���'8��2��i���O��#�ہ;k��S�/~�[�nO�d�.L��!� � ��.O�1n�]y��'j��'W2�'�"��6��0��
ܚ?R0���J�ɾ�M�T!�Y~��'�񟎘a��6s*�Es�&��Uq*�E}��zӒ$nZE�)�:ZΝ����$�3��I>x4��.�=HXЗ'V|��q�8�M��.���< �P"�D����������?!���?Y�t�@�� �������a'�k�U����,�l�
Fҿ}���0#�՟�ڴ���|
�U���ߴj��'8q�ʁ�2�S�A�xE�V�	3��9O �$�� $P���2�`*O������%̐4����`(�j��9Q�h��<��?A��?����?Y��Tc&$��t�P�-z�v�j��C<`6r�'��d���z <�Z���ڦ�'��)�o�/g�b��Z�e��r����ēD2�vluӈ�	��S6�l���	�b��$���E8�5�Cܥ`͈l�BD$:h� ���r�'j��ܟL��ğ��	�_�ĸ�c��S@Z���Z�a����	ܟ̖'c�7��c���O����|:R��<pZ�
 ˏ#3�ۡ�_~rm�<����M��y*���QB,V���*@��ʈ7����L]�F��|*�+��M� �|���1]eP�ɲ�э�C�%���'uR�'����R��
�4(l��bG�}Q�tK�&���P�	 �?�����V�|��'�n�E��� �4"�1b)C&鶹��NT�&��6-��!��Nצϓ�?A�̓�Zh�)���	gm��G��PI �뵅��o���<	���?���?���?�.�>�ӵk5*�I��=Q��5�`(����������I��d&?��M�;?rV0@GU�A)���gA+@	}�e�i��6�J�)�.eB��e�l�G���QS�������uJ�Ir����r�t�IVy�'I�d�*���#�����Dٔ.2�')B�'�I�Mkq 	�?���?)U�G��H}��W�'�R��SIY��䓦?�V]���ܴi���|2�M4]���`�k\H����y��'J��� "�#��!83Z���~�6���?�J�w�L����b�J��S�G,�?���?����?Ɋ���O��ȇ��D>4�r�ݭ��!��J�O�Em��c��TW�6�4�μ���W�_ޤ��3��Q�9O��n��M���n���b�f�F~��O� 40\wMVe���}LXX�jK�=����`V�	vy���$N^XU��νu��Q@W�M��X�P����7��	ǟ���iǪ+��}� ��t� �B��4��I&�MKc�ik�O1��Q� O ?Lq	0��h6r��&	P�.��H�<���$Qf�ć�����D�1XC���s�Ƭ��K$�p�[���?���?���|�*Ot�oZ�)F���ɮ\�h"B � |�H��%��ZI��I��MS�2��>�ǻi,`7��}�u#R%���:��o�굈�	��#�~lZp~B"F3<x��78��O׊P�vM^��ׁ	�F�2�Tj��y��'-��'�2�'|2�i���5Kf�[2y�x�+���b�����O�����q��|y� w�ԓON��5��8~�A��M��	q��Ї�K��M�Q�i���-�,b��6O��U�v�j���l@,~v(�ҥ�JPj-&�:�?���.�Ģ<���?Q���?�Ƌ����֋]���@��R�?����[��k������<�O�0��@U�W���`�D�F���"�O}�'�6��Ʀ%HM<ͧ��'� ,�l�&�����	u9Tx����'��T(O���ڟ�?�S�)�dA�x�n0��F ���m�r��O���O��	�<�b�i̽!�I=QB���Ʀډj�����H$r�2�'�H7�O֒O�T�'��6�H�ZH�cg��Cd�@�.�7�0�o��M��g��M˚'���/z8��)t�)� � ���'/L\���S���9U>Oh˓�?���?	���?a���	�|ה]*��[)]Od#2L0LŬ=n����t�'#R�O��S������"/R�D�Hz$f�	OAԙ��d����.c��%����?��S�X��)oZ�<�r�Éj�%�ѯ�c���+����<�� �2���>����$�O��d��Z��b�%R!��Y�cүG���OH���OT�0r��E:�y��'�rkD���MÖ'��~RTӠ$�,��O8��'�b�im�'��#�
ĈtMf�S�hY�X��!z�O��Е ������ �i�����_ោ����J���X��y���w�Ǒ�?1���?���?Ɍ�9�:Y��"��:㴀�n��c�,�S�O<Do�>nZ��%���4���cF��I�DuI�/D�@ܶP��O��Dk�d�䄟 ���s������(�b�]3��Rj�2撝�'b��hܶ��|2R�`D�%�$@m� F�A֔p�ٚ���F�}Y���@y��'f���3K��>0
���F�:���SƔl}Rjt��o��Ş[�u��m/&]QI��#�x`P�nR/c?v��,O��s�aU;�?��O;�$�<�k�&�Z4kM���$Z)�?Y��?����?�'������xӉt���a�7��\���͊P@Q@�p���4��'��e��F�y�.�$��.͈��G%8O�\
&�{�yC�)��x���9�>d���qݽ����4�w��@J_+xE ���)��q��'�'��'���'�I�p��-iybɓ� ^; ;z�9O����OZ�oZ�-8�3��f�|ҍQ2,� ���)Y�O}�����#C�1O��D��	ÓZf&!咟Xcth��YwZ�f`��L0=�&}�ڬ���v�0�[K>Q/O��D�O����OnM:hs"X�"��$e�)�O���<�ipfdT�'���'v���Okp8���S96�YS@m-t�t���'��>��i�z6-�g�i>��s��c�?� �镋HL�JeR���,A:�p�Yʓ�F��Oz!(J>�Tb
%+=؝Q@��4E{����?I��?���?�|b(O��lZ�:[��DM�2nA�A�ب']�!�VJ�џ �	(�M3����4�2��'i�7�_*C~L�׮�.�dЁkU9y6�n��M���\��M�'�� ��w�re�ӗX��ɰn��"��I<E�ֈ��e��+�N��jy2�'J��'���'U>a�fI	%�Т2(M�M�&Ei�叓�MÇ	M�<A��?�H~ΓCܛ�w�^�P�$����0G�=���Z(�*}ӆ�O1��(��j��~G���,�hu�#h�fm{!N�LU��)xV�@ѼiQ"�'���'���'�
hV�ma�5k�40g>����'���'��U�x�4<�~����?��v�r��%��X��tŎ B�A�����O��'�6-B��m�H<Y�
P�p0 �� t:�Ðe��<q�l�Hp�jZ?UYh�9,O���*�?�1G�OX �J�8|-��rWOFd�(�`E�O0���O���O,�}B�"R
�����X���k��@�Z�$�J�u��B���D�Ȧ��?�;3 t(�c"�zN�`��A�Sr>��.!�F-iӔ�䁃|քб��	YFٙ���H(���E����s���4��`q薰�䓗�D�Ol�$�O�d�O��$�8ٌ����)���Ќ0K6�X}��� f�y���'NR�Oj�$�'r�B�R����T�܍�� X4Z&��M�u�i1O�D�O!#�e�|���"� Vu-�nO1y-��XpǇ"�򤓺=��a���'�ı$�h�')���P�.�}l +5�"!���O����O�d�O�I�<�6�i�jy�'<`9�0͛� �J�X���_��3�'^7�6��7��dIަaJڴ�?I��S$�*�Ñ.�:��*�@�z��5!��Q~���8!�AbXw���&?%�.M�L��H��MS�};t�_�Lr� E�4$�,8��ٺYS��(��G�d��#�K��Qk��{��Z�XZT�ۂ@�ezx�[�A� I�l��F�o�L�fԻ_
l��]/,m.��8t�!Ĭ�
�@��C�� �n!SG@k^Mzt�L �X`W���ȩug֣M�A�Š�l���y`�5KC���P�� ֋	�	��bݵa���Z8h��PΠ�kb�#t��uAҧv�a �J��1��-,nᘥ!%�#�Kd�2��Ƀ�H�	
�(�����x8j 
�E3Bdz޴�?����?ٱ��0̉'���'r��NSr�����E�v���3rEߺ��'�"�'���vA=���O��D�ON�a4�Ȩx`L,yO�1���/�7�O0�S��y�i>e�I韼�'EFEiWI�Jl�%�5�A����ae�.���?�1O~�D�O��d�<��Dƈf�*hZ"�Q�J�I#���c���(��x��'�r�'j��ڟ�I�q�ak�Jږ2���*�&F9GԘ)���<�� ����h�'�`j&�>]wC[M6�8 ��w�XU�@��>����?Q�����O��C ���Ɏ������.��XH6��?y��?I*O�$�ca E�S�# Xq��/�p�� �<^����ش�?����$�O���ԋo1��x���3�P�����I6�U
��S¦���ğ��'\܍�š9�I�O���ư�x4���P���0ዐV��y:ҵi��	ğ��ɛ,ߘb>��I�?7M ꔘ@0���$�b��'8]�P�0����Mc�U?)�	�?I��Of([3��2��\:B�W-7>����ij����S�D���43�ʬ��V�O`�pa
��R�dn�)F�]��4�?	��?y�������d͵���*��D>D}��!0)\�e��7M�%�V��?A���<	�e���;F>lM<��'�ڂA�0��E�i���'��BRnO�I�O��DQl�? �]r��r ��4�˾M,41��_����䟐�3�(�	����ߟ�TI�v��U�MO�L'�]Bs��%�M���>�8�顙x�O<��'���v�&�Q'
3'-@�i���W�1�4�?W�_e̓�?������O�w+Ɉ'���ie���X�̔:7�P�^��ʓ�?	��?A�R�'Q�񰆞?�
DX��P2c�2�)�ҷ�8�OP���O ˓�?�uK����h^�!f��f�)����)	�Mc��?)���'��iZ�q���aشiĘ��%�>~2}pd�-o�Bl�'���'��Iӟ��f���'I� (����#R�����`�����y�V�D(���d�@��}�O������L�#`\G�$��iB"S�<�	�?�X]�Oh�	�?X���B��)���[6L���q(T���'`bG�S��\ �y��vi�R���b����g�03`��7U��I�v�:U����X���4�QyZw�4|��	M�V:zePC.�h��4q�OH���GW>�������~��H��l�l��%-/�6�ۊ)S��'�2�'��$T���֟H�� 0̈́8�sM��)��I�H�&�M��F��P��<E�D�'B�ԩ���T"!MåH�:ѡ��t�����O��$�">���|���?��'u��!�MCR��Yck��;@%��4��=UF�H|���?��' �E��e�8}^��j�aٚ9�jZ޴�?Y�&@���O��D�OT�<:dK�8���/_w�-8�E,[�ɦS���CT�>?����?�.O��Ē�:�q��	�r(Z������ ��<���?!����'����/-c���&&pr��BD�l�2Ԃ�����$�O��$�<��2�.`c�O�؁Aqk����'ڼ(�����MK���?����'���+���شD�yӌӖ�%0E-�7��(�'�b�'_��ȟiңBr��'!�'
Z�n�����,44z�F`ӆ�$"����DC0�LO�"Ej�b�-
�j?�t���i�"^����4%��O���'��D��9X,�#�4b.y���Z���b����
JJ�F� �~�D�E�X>x����X#]N�i�u�b}��'�F�{��'R�':��O��i���7��g�Աa���=\�XlˇD�>i�UN��k0��A�S��s\X9�C�!Q}r�$��0��7-
�$1���Ov���O"���<�'�?����(T�6��D��?O��ʶ္E��ɚ%�"<�|:��H�<�چ(���r�-��=�"��E�i�"�'�2K�3��i>�������R��-��)ҴY�h�`�2d�j����U=���&>��	����#Zv��o�;[� �rj�R .�n�����Z`y��'���'�qO�A�p��(N}*!�ĥ\6%0q7T�Hi�F�Q���?������OR$1WFۜQZ� ���X�S��}���BКZ.O����O��d;��ݟtX��n�t�����=��i��8*�Z���8?���?9.O��DȈS����#Z�t�r�h� a��|�vkA�|.�6��O���ON����E�gi�l��B��j��`;�!JedNc�\�������'XB�׏l��Sɟt!® 8���c�IG
'"�(g��,�M���'��&���asO<Awhȱ&�¨9S	P�j4��'�֦��IUyB�'Ś�2$T>%�'�4�ش{�l�Q��!��l[��U;�db���ɀ5��YhE*9�~J�S���:�ߖG	��'O}��'|�AC@�'EB�'^B�OE�i�aITMN���x�g�Ia*達�>���^L�ꧦ�[�S�k��L�Ɖɕ\-v�ЖkJ�}�F�l��:��Ißh��ʟ���Zy�O"�d� \E
9��E�4^�4���mY,6�ёtCBub1���ݟ�)TBK�1pYav�ݼdNj@) Ɉ��M{���?��t0�/O�I�O�佟9qO\�Qؐ�B�V�7l�(��%�.�'O�m�!�3�i�O���d� �߀'U\�ل`��B��;p8 7��O
 �)�<����?!����'}��3ÂѪD�艒�(f�,���O�ݑ���+;�������Iny��'̐(�V�
;���U�ـ1��X��j��	ןT�	��?I��xɼ��Q��!u�^�C�	K��Кq�_)a*b��'���'��Iڟ8�e��Lڔ&�"i�R�3v���{��4r@&^妡��Ꟑ��\���?�� j�Xn�XX��9��z$���$C,��?)����$�O�E"P��|:�/�hQu��F�k2��s�I�Ѹi���D�Or���H7=��'Τ��!U%eS��(N+�����4�?Q-O���̣dS��'�?����EC"�(�V*-����JƖ[V�O(��ȑ]��r�T?��e*�#u6I�qI߾l�L�pǣ>��M�a���?y-O��I�<��`~�UZV�V�8��ǫ
�@Y�'�R�%Jb��k�y����H�r�l�2�Q�3��e%֦�Ms�,ڍ�?i���?����)O�I�O��#pb)^~�(���O�VZ��#����-�����e�c�"|��c��)�F��l�KC�
�Tq��i�r�'l��A���i>�����+)����tD�jրѣmi"�Je�Ěg�m%>9�I�����2����.C�[����ՉA��8m�џD���Ty2�'N�'BqO|���L��?�0�� H<,�83�Y��G8x���?9�����O�s�kD�o����US�r����I�d��?����?��'�(� � x�'Җ?���� ӄb8�a�d�Th�ܐ�'�"�'��IߟԳP*[fZ֫=oE�x��^�g)"Qr�)U��Q�	؟T�I`��?��4+
hm� :,La:  Uw�ziI#�к��7��OZ���O6���<�a����?����~�ϣU��� ��	x��cH͈�Ms����'�R�̥���O<����
a�h���
����,˦���Oy��'������O��ꟸ��4eC� >n�ɔ�-V�8aC���D��?���ErJ|�<�OLJ	SW�W�Ǵ,�TdE5-V( `�O`����*����O����/O��D�d�����e��|�A���I�Y��I⧯#j��b�b?Ӧ&W�1��@A�M�P�BXs�'{��\� ��O&��<)�'��4����H.K���RfX?\�l}�w��5�0o�����p� �)§�?�7D^�(�P���Wl>��0c4Y��'���'O:܈vR��럸��M?ل!&M_���c�mG�L����/2�1O�X��GP������	g?�v��<WE�P��J֟h�.��,�I}rj�U��	��p�����=	���g�(�� ��"��9Au�F}R�5=����O��$�O���?�&-�`5*g��Urr���d�|�ꉉ.OF���O0�$8�I��s�l��FE�D�r��`��MiBn[�lhՓ��3?����?)-O2�d�\�(���)�� u�Àh��)qm71#�7��O��d�O�㟈�	�1Y�p+P�u�ȝ�JP���%��@D�T�-(�]�|�	���'#��O-d��㟀`��`��+��ݩ��H���	��M+���'$B��iX�=`L<I�
T�|�pؑ�G[�L����Q�Q��[y��'{~aZ>M�I���J��l�Ǽξ���\^g�H�D'��ٟ( ��3Hb��'L��GnZ�[ ؊�Ҍ}�8�l�iy��	pj`6�O^�D�O��I�L}Zw�TDx@A\�O��������X��4�?!�!2͓O��۟��}bG+� U{�|����F ��G�: �G�?=�87-�O����O��i�g}"]���,Xr� �l"YH�Hcᚹ�M�4'��<����D"���� �O�&@@
�����YRd��M���?��c�E�\�@�'G2�Ox���_�Y��a�F/"/�^H��i�"[��3B,k��'�?����?��R�+8�3���}�$�*B֭Wɛ&�'� ��6 �>!-O���<)����d64���I��iG�$YPLn}�ǆ�y��'��'��'o�ɀ#�L2��İDv��"�dVF��a'͚����<Q����Ob�d�O䈠���&cz#AM�.̬��e�)�d�<y��?����Đ�RYv1�'/¹���
sg\�B�[��$mZzy��'�	����	۟��dx��s���dOĄ���R�l�0PI�	��d�O��D�Oz�-�X�]?��I�dN�!���C��������L�9ٴ�?*Oj���OP��Ҏt��D�|nڮ4��b�Ze]�x�҄�?��7M�O���<Y����՟0���?�C��3d����Ìt��hT �����Od�$�O�-a�6O��<)�O.-ل"�s����Aܾ@�����4���8+�n�����ڟ��������Zy���[�0H� �G�0�8�;»i��'���;�'N�	ß�}*��8P+�����@xLh� c���Y�NE��Mc���?����A^�Д'Ođ��*��R�8:�&̪7�d���t�L	�?OڒOX�?��I�|�bE�C�ʁTR�1k��tv����4�?y���?`3*���Ay�'G��T�AN�����S���)Oܡ	��F�'w�I$���)J��?��AN���N�5? )�B�FQJ�R�i�,��e�듯���OR��?�1X5@l&�%)D����@�?=%�'eŨ�'b�'�'�2P����=�
iPd�ƪ0���E"A�r~���O@��?+OB�D�O���:5����.X�̌+�^-���0O����O����Of��<Acm	 Ni�	)$G��+@�E��r���{��6T���Ioy"�'��'�����'G������;G�Rl�C�)K��&�v�����O��d�O�ʓ*����E]?-��>Bo����� v�-#C�*';�}��4�?�*OT���O�$F�Y�1����ʬWj��)&�I5=�N��B坾�MK��?�.O��aek���'$�O�^�!�I�k��L5����7@�>Q���?	���^u�'P�	@RӂǠq���q�/h$H@�\���'DZ-Hc,b�x���O�����|Hԧu�D�p�p�X7�DEˆ
���Ms��?�7���<Q+O���/��a�d�"�_wpt���ؒt�7�8&X�8l�˟����S�����<	� �/p��HceG�A�D�@A_�6S��B��yr�' ��x�'�?��*Fp��@&l�"2���q��@�PG���'��'V��+��(��On���d0�&2����Mو/j�hrqb�ޒOh ���O.��Ok�] h��qҥN$�}�9u"�F�'�^)��L9�$�Op�d;���zs)�][�E)��^)�\�!_��q�a��ʟ��	��'��|@��� �`�O��^u0�&8$��O��D�O$�O��d�OJ�1�#�T�`��$^�2В5�؎]����<����?9���$��&�X�̧�  �.� T|���#V���%�|�	hy�'���'sFI�O�ۥ�=~�� 
��
L�4��5]���I�����oyB M(@	��t�2u.�L�̓AX�db���A��p�IßD��z��	V�� <�0ChV)�r����K)Q-�W�iB��'8�ɨppp8:L|����C舢fx̐�M��M��躢��C��'�b�'t@
�'��'��I-~�6�o�#4�����Y5Gw��_���e�@��MkuW?���?UC�Op,��`(lh=h�̈#����i���'���YC�'Z�'lq��$�><���Sk.{�Q�ǵi�:��'�q�L���O�����0&���I�,��R"��L�^�8�kA�z�@�k�4������Z>��'�HɁ<P5�&2sI6�����,6-�O���OR���EB��?��'��<cVdZ�Ԝ�U���@�(���4�����C���'��'Θ�;�U�Y�%p�"�H�c�&t�j��F�"ϲ�'���I՟ %��/��E� �ð<��U�����.�o�����d�O���O��pV��Ñ�$�h���\��-�u瀕�}��'t�'k��'� DC�"j�6�zBn�pcd�bK�H3�_���I�����y2���VX��S6C�>m��B�@�b�b�c��듆?������?��\t$���D�i �{r��:�H�06G@U:@^� �Iɟ���Ayb��%\��� �D�Ǥ'}޹bsH"?���������E{��'T�\r%�'��i��0"�F"���b%�	|p=o�֟��I]y�,&|��v��kLɹO�W�
�G}���T�?zb�O*���8�b��5�T?9�V D&t��1�@��'uϴ�;��g���O�l����O,�$�OZ��㟌���Okl�uJ����á? 6���	Gn����'���#��3�y��4L��P �!-����NZ�H����4�  �]�ŉ��?A����X��OBB���ޢXSn�@��Ѵ
w�1� m��Q*0+(���?I%��	{@N��$J�{����&�"Iw�9�ߴ�?����?G,�<�?!����)�O��	�J�$,5�Q�D��ݰTM���jwN-�ɯ���H|���?���c^e��Ս>��1u�����ֿi\R!ߝ1��I�����OH�O�����L5��:����/�u�5�Sx}2�OT��ك�O���O��d�<q��T�{tP����z�٤$C<|(���P�������	ǟ��?Y��[�h��<"��W�F�(�!�C��gl8JN>i��?����?a�fo�;�OϪ����B`��^��A(�Ϗ)�M#/O�� �$�O��d�mv�����iT�q+fH�.�j�`�I�"��Z�O���O@˓�?���?Q��?�V��l�2l{��MޒR`��0z��'��'���'(�l�P/�-�ēl#`��0\�֨Y2蓿!��o�ݟ$��Zyb�G%��:����@�F�mD%���;%��#De�R��͟t�	�Xj�"<�O�*����J�观�?a2�;�4���'"�o����	�O��i�p~��dm�� w��DI���ReE�M���?�R��M���OKxHȇ��KΎl�S'�#�v�Pߴ#���T�i���' ��On,ON��E�0,|bR0��!h2S��mx]�#<E�t�'%>���	�&æ)&#I@,ѡe��$�O>�$�;�˓��	�O��I�l����dDˆb�h��W�W���c�L��#'�	�(�I蟘�WV�lO���SA�!M<���!E�2�M��.-&���?y�Y?��	a�	�l1dP(�l�7���T.M�J�S�O��0�ǐ���ʟt�I���'L��ZA�\�L���7-˶W*t��c_;�O����O�D#�	OZ ia*���^����`t��`8�ğ�I۟,�	�l��*�w҂�@�КLZf��1#@�{2-_Ŧ�	ҟ��	l�Iҟܔ'ԕ��4T8�7=a:pA`�#��"B�\�'�R�'aW�`��j��ħ�qS��-�D��O
�5k�1�U�i+|��'*Bf  ��'5���S��
s�\��f�z��(ڴ�?����D�-z<�%>a���?���8.�$9Y�j�$C���C�S����?q�K���Gx��"@�F�S��`�IkwVةd�i��	������4V��Sǟ��S���F�H5�:��9�K�FC�o���'����O��, S�C�lTL��lU� EX@���iH����j� ��O��蟬Q%���I�J����� 03> �E���eb� #�42Ͼ�Ex��	�OZA,��mX"�ķ1c~���;^�n�����	ϟ`{d�ˠ���?����~��B����A>E���a����'1�Y�y��'��'C��y�B=g���`�G%Hp�c��l�8��ͮ$|�$�x��ß�&��X
e�X1���O��P�ޞ?��ST0u�=)�BG��Ja"]p"t��X�$����@yp�I���\t�	��BD�E���KUj����Ϙk	Z�:`�]PQ��tŖ**��6�D-��ňu�
?AC�(��?k�f�k�m��2��u��x� Aӧ샻<�^Y��@�W3���4�)G��H*`k�+�����D�(�q� 
�H�.Qz���%u��!��E�9�t��נ,�,����I��-"ǃ;f���s�MͼG��x�o�KQ�x��!�9�	��\�q<�1����E�t����@����=�r�a����X��4I�1��ɀ�4���7�W�)�&8��3�Q�B��M�Hhx�������9���/����D�#�`s��"G�J�K"��X�Q��5n�Op��!���y	6�sdGA"[lD��q�B�mc��I|����	�%4�P%i$-�����>�OB $�� �z���5͜X����j����=O�QFI`}��'J�;]=6��	ҟH�ɥ&�&H�B_i�h��˒]�`��̎갽�ՍϢ��q��S���'��	  ��(��)�1vK�x�oW+;kN@!MΒ%��*Tb�O?�D k0q��i����X����8����?I������|�cܩl���F��w���F��:�y�� }F�OI�g.|J��$�Ob]Fzʟ�8*��	&ĕbF�ݤ9`\m���O���W'G�8r��O���OZ�d�ĺ{��?�p�Q�
��Zre��[���DfU�; ��28:	æN��x
�U�g�'���"+'0���'\�/��t��OṚ �+Y5�P�ܓ����$�	a�%���'f��c0����ٿG��'�ўԖ'�$����Z�#ꪐ�t�sK���'0V	��6lE��n��qP���*�S��R�d�'n��M���Ŷh�Bژ3~`�rG���?1���?��o�������?9�O,�}�eh�+�L���	C[����J� ���ۀim$4A��'HtA+f�^dȡ���^��d鈀���B$MX .���A��'���
���?Q�eL5w�8�s1�H�|T�&f_��䓆?��������ȃ��8���:iɲ�Z���#�!�$8$Rڽa��)?�fa�!��Y6�Dd}�X���e�Ɔ�M����?9,�35�;mfh!����{?���P��/$���O����=J�����&�� QF*OL��'-��8 ��	���������dѐl(��a�Q��N�q�k^���)�);�p�Bnģ`v�K��
�Q�x����OR���Ot�$�|j���#!�=Bc-߅9��Eyh]��?���9OZ����,F�nq���W�uH��:��'BDO��дl��,����G��#;d}�E4O@U;��[}��'��S� 
���I͟|�ɹS��! ��i�V�`u�ثL4t�+J�r>�X1�툐c�T)S�%ɽ���.����4���^o������Ër�αb��#�:Ո��/)w�a�JзbS�F���V4]`�K�T�`M��%��p�i5 ��?iӼix��S��?�'�|Ar�G� ��h���?�m�
�'�20`��-v<ܸ�$�D�])��H�'�7��O��{1`T�+ީDj�(yP�c���O��UB��"���O,�d�O|����K���?�"�sBY2'�F�a��0gĊ��VhH��D>��b�fOD H����HO`���B�;��m�AkN7n)������$6FJ���ԍ+�8���2m��!ғ:$8��X�"��LR�J/�����c���Ɇ�M� �i�O�OW��$j̵Chjɲc�,V1����' ���×�O�04��zBf#�o&� ��I`y�Y�d�7m��݈YJ�k� ��`�[�H�\���O����O0�JSM�O��p>]y������jA	U�=J���Ǩ�oЭ�CK�R���H��ՕD�tD��Ò���J�$��n��J��ɿxR�l���;�j�@ƶVxX���	>NJ2���¦���[C�J�iŖ�IY|�huJ��M�"�"��<��Ҕ�T�����1�x���QW�<�2�^b�B��3�J?^~<Hx�L�<١S���'�F�#�e���D�O4�'kz��S��joj-�	�?m�xM���C��?����?Qv��)M�����POD����K�u3$x��c��p9�/P�1�Q���KFBUdX�qE��?m��$>)���Bu*nJ4��3l]4Jѡ3ʓ:��I��M+��i��Y>�j�@ #�$��]XH�#�$-�-��L�S��y⎁�r�ڰ	F� ������$6��|���x2�ü0�ܸ9wO9��6�,�yB��'X˶��?�-�������O��d�O6� f�91��DCc�R�P����W`�F��B)Z�E�k��M�Ou1�2L'&S�A �E�� �˅��)+CD�kq�p#�����\O%�1��>T�9���;.�<��K4���:�o�(0R7�ۧ��Cp���o�؟PE���i��t�Gg����Ya$NڨI���̓�?�	�^�2�� Y�,��@U�!,�Dx�k:�-,ҵ��Kc��ڡ!�<"�E�Q�������?�%�ML�Y��?����?�A���$�O0���h@��n%{�G�S*,`i��O�hA�����*�'��I�`�Z'l��S�H@�x���'�(� pbي{gzxϓ.k�M�D�M�V��`CĄ� �n���N�؄��?��S�'��X�pJr(�Y��At�Ո4�hpP�&D��kDn��Vd�xh֮V7�"A� 'F�HO�i�O��(9Ɯ!Ǹi��1�G��V���;MƼu�P�[��'92�'�"&���D�'�󉎤Cҥ!��'����`��u'���dNU>}ʼI�	�v�,���C��d� l�%nT��A��O�3�{�-&�O�8H��'c�+�F�u���/�0`[���E��' �I�D�?�Oe��)7�%b#D�D�;C�@a�'��袀`Q�P�s�g�8瀬3�'������M,,3��mZş��	j�� �#V�Y:^
H��̈�n�c������$�OL��� �h9�`L�lf��S�4��"�J�@ȑ�(�<xJ+�(Ob��	0ߘp����0�P���m��^�q��7 �Q�t���O��$+�	�O�� �@�;~��B�H�!��I���O��"~�Q~8��"蝄:MP��'��H]��񉁶ēB>F�{/ڒ\}�Hb0ڋ7�t�ΓR�dEXŷi
2�'���G�$��ʟ��I�Mre;��0  5� �/ZXFq0�Z�IĒ,	!�������|ZK~Γ�����O�FDjc��>Z������K����	>����B)�4"}���?��&Eπ��RfR�c5�Xb��H�,�i閧
���'�4���)u��:�*L�@�骚'���!ړA9�S�A@�Z��1(�#�.�
Ex2�z�f�lZj�O
����AӮY��ݹ�&�.��#���?CL�F�Bp����?���?�ն���Oh�(LHRX0�c,r�4�b�O�ԛ���Z����`�',O ���	�$R�r(\�V���G�Oఘ�/Z�z�h}�'�>,O�����ڈ����C� \���O��p�'�D6��U������Gy��-v0d��|Hčb�b[!�yr)�3Z�<,z�-�1v]�07�jh|#=�O��I	`nqڴ0�BvbQ��v��b�k�>Xx���?A���?q�����?�������=H��"�X9��l�.>8��*�r�6���	9wP���d�O�H�c!Ά]�L� ���;��aQ�'��l���?	�,ūDlm�ͭ*  ��
��?������O0��'1H��ku)��7��Xc�*>HWb\��^�@֥K� 7T��@U�	R�����	~y��1<F��П���W�d�Q�%:R��U�=R"�hB�Ѕ?V�)[b�'�"�'0����:O��O哵"B��Z�,Y�7�.E�n�T��<٧삮b-s��V�@k"T*0���~셈GA7D�Q�xK$��O�$�O���|���A���3b�v�������?	���9O��;���$?�����#Iߪd!D�'��O�����3[�d�5��}2BX���	Wx�x����1T.�5 GҀ'E.��� %D�d���o10�zBQ)T��x2�=D�,��݌E�p �d,Z �	&F!D� �v)�'f��z�J��2��`%D�����n��0:���*x�)A	"D��k7��m�Dٴ�D�c}(a�?D�|���կ<��u����4W��b:D��yw�57�
��`�k����c9D�*֪Z�{�%��H�Θ�0"�<D�軄��5'xe�p�I�W�p�*��:D�8�A`I&
�L����9*P�h=D�pq�`��#����%E�E�4���.<D��0��������3Lu��;D�h3�)�_��cv`�TU�;�a5D���ti��1�ܷ��(�4$9D�	��ѕHێ�J�\�hZ$�9D����ǽ�j(S3��F�r���(2D��[#�[�PfDP1�+�j3w�"D���N�L|X�׆��W�drdN4D����cL���l΄dw\=P�1D��b��_�w��[�7��y�`�$D����B=t��Y�CJe���j��=D��8�c�C̀��`B[�L1p=`c	 D�t0�[w�0��F.��'�>5��(<D��ȗ界b��T]HE�d�9D��`�Z|�b:�  3���W�6D� ��*\%��xQӣ���"�/D���Gd�a9��"T�ܫ"'�k�I0D��8���va $�!�ƁCL|�I��+D��1�K��P�.Q+|�QV7D�0�@/+] ��EA�fThDB4D�t*&�	�/��U�C�_�Lw0�1��2D��85J˾`�Q��[�O���@$D���Ǎ��+��@���m��¦ D�\Qw��k��E(�*�1W��("&<O����̊4F\�x���>� ���G�8F(��{A�Ą8�S"O�A��D����}C�T����Ց���(�a)��SãSH�Q?e�bb'r�u�D-@�d�vU�#k!D�ʃ.ӢG%� ;�F�
M��mҁ|h2,xP��C��b��'U��%87��ļ�W+���P
�K��q���'V<�S#��2g��+2�˱-R�����$l2Jt&������,�Ju(w�ܟb��&M+�In�Y�6G��ZDl�z���|��Ě�yZ��`�kő-u���'��9F�h�8@�D�����%؄�3���V����@D!��X�_ ,Y�K(�<9Ȓ�'`-ڐ�'��xp-�
HJ�#��%ck�}��'��<� ���!3��uEFx����&v�蔹�]q�<�l�U��JP��%�|"���
I)S�#��D5l�?�'e|`3�����|� c �M�;�\�s��fy�� V��Q�v)�i�'�UơU0��y4�C�9{��1����y���	5��,|�J�B')��<���0���A�T4���y�E���#�>C�:�
��h�'��R���6�0�1����`��x��[����JŠ܎�0�Jf�
���i%�P��	̟����S�6�B�՞SE0���h�$�!q�t�²i��+�l0��肁m�K�8�d� -D�; �*���{
�k1�X8Xb`� ��1��nZ���B&��d��)���	�X��4�J�ls�'��`%t,� *l:�\9�%���y
RJ�����
,��}y'%��Ms&#�=5�,`�D� j�h� �!'���2�4	�`���e���>��~����go���b��V�a�`�'��`��F�!`���/��x��	�D������V S�8Y��+I�/H̒�ݗ�� #��u�'>��6����|�)K(p¸Y�f�$vnUkW�%?9�Պa��!6~@���W�r- �I͟pd�4-6�UjU�5��Ԥ�A���b��]�֎��'Vm�v������9K�"����aHx��Q$!�	~�\ �,_;"a��Ѣ�O!x���l��k��h�(�-4�( �G0��'?�i�O��1��ߏ_��Հ��[�<�Aq�<����&L-���	cY �s��, М�O���2�!Ϝ�U���p�*i0���?�5��&�<\a��6�Og��<HK��C2��9#�e�NB�A�x��4�X~?5%0��-�@C.��D��$X���,h���N��eS��)%��+G������(ѨOt	[2m���.�v��K|�PQF�KV�����7�6����@��D��P`�o'XX��l�*%k#F��"cp|:�ƒ�-�\]�O���D���U=�%V�U:8I�ј�(x b[�`+tq�ԫ��6�UQ0���(��H6B�~B�L^"阇���8�x�H�z��5�c,��Y�܋����q$q�R?�A��F<�<��O��ʷ��X��2D
9s��Rb��<+����	��q�3� �/-��S�D����=R!�2o:wP�	A
�0��'�h3v�p��pd0���I-4R %�Y*��JT(��+D#� TaA�`8����RU�R����8,�ꨣ�ƙ4n8|+V���t	a�\1��C�L(�A��'N��ũ�)סO� ]2��7@��I�J�].�>�r���psV)F�n��a ���iE�D�5.����+�!�����5�/�1ю�Q�OM��1��֎I�"�ŗ�Y�y#��^��)��*I��|��'�`��KP>�"�[w3�,�B�Wx5���>�ȝ7됡[1�B�6���be`T-aO��{�	�U.ekG
�F���dE%G��#�U+	2=���9�0���P&Z� �(Ó\N0x���: ����
K_.TuĈ\�|��	L'[�N���鉇k��z�D#��#)��v�,{�i�j�)���3��'���X�dZ�忣'%I3�ԙ�N�-R�lp��酭����q�~����ԟH���郇W6&IK��W�^^��Q�W3#c�P����-#L#<Ѥm��^=�!ç
�&�����a~��
$V*�`@*v�RQ��#�?��P䦅��V�?�T]�@�ZC�)AfJH�ɔ<�@�h��];b{��!N�3J2�L˗D�v;ܴ!���[b=� �>O8MyR̈����vNʏ���p�ôgU����ݍ,g���5��IX��3�N;{���/�)����oEj�O���g5�Ӻϻ0�� C4)̖ê��dm�5���+; ����@87��"Uc�"��*�HL����R�&#=�;�D�Q
�z^��g���!��ܙ|��I�OZ����t� #N�Gf[�sy����H����'�B!v��7m�x�D��'wo,L��O �k��C2�<�ygi��	!��>�e�ݪ������gh,�ץ�-6ܬ���K?k�Ru���<���̈L���N?�K4�A�Dd�dH�ꏘq�t`��f�c�K@Y�D+���4�j�3��Ȭ �`d�0&�/J�<�e0O��HdWD?q�Q��>�a��C�n	��.�$[�PP0�5l)&1�R�'�$�����)g�`I5�ٵB7�CS�B���rť��Y��r�fZ�g%�	�6jv���'OJU
�镒.��S����MI�Og.IQ'�	��hl��n��|�O���b��"��� ��ij�8cQ���ЛK��|n)j]J0@%��y� �����M���� C��� (����0�	*��i8�		h.�93� B�C֭�@���,m|��b��'�0�8�iͺI��ɈR�+l&�s��O֭�'��H=3� ��M�ș�R�<d�QX֋As���Ѐ�)k��y�wy:h�aaJ6nU��ɓ@��k�r� ���_��$]��M��V�x���,�Ӻ�A\�
R~Pɂ��
{x4p��->i��@�d6OT�����<7|�	�N#��d��	]��l3�,(C.\]���=���D�Ob�p`��7�?٧]�Ql1�$*G&L}��M�� p&�X�Lʄ����ŢxŮ,(U������A��}Ъ�"�T6-��r� N��~Zw��!�p�Ѕ q$���y>,!�	�H\
�O����iI�g�I�1���A�A���x�烸J2�ZC
0��ɡq�>���(RI?��y��ü�w�[?�V�Ul+#\��n4w��qDd�E&�0�m�	OiF`B��4�4�F��f�3�I2|�xm0uCR	�t�	���DB"Iid��uh-~;�%�#��&��)DK�`\�RE�		����g���B峀6���U�fJ�$f�X`a�P�;���%Q�x��?>��i��C~2D>��$���9F'|<� ����^y�7�M;y�bP�ǐ2*Q�|c����*���%Ԣ���h�o}&�k#��?��?%E Բ%3�	�CZeC"���"[��B,Y6�)}R-UV�$�B,)��� Z�`�r%�
�06B�%4]�� 5o�h�B���� #�dX@�M_,s�b>�)�fN
/R[x�	�d��f�5`~]3#��m4��36�9m)��(t7��=ͻ�x��k�X�4�UjW40�H����8=�Љ�E��%vD�S�Y�L=��+@(VҰI�'�	��QNaX��"�P�R">1��!p
�H�&�1B�^�!B�0��ٺ�A�G	��uI��4才�T�s���d`��G�7tF���@I�9���%?�s�A4�$�#���Hݫ�(!D��9�j˾��X��C�(�e�#'��it$�U���xԎC�Q��'K"�t�u������
qb�H�'J2����(Z7[ma~���vVA"c
�I(j`r�T�b��@�!0�a����XDk �+0y\�S�I�'6�*�������p�T�8)~#>I���E��$�q���h�/ԍ@�|P�Z�f�:� 2pXb��Q���h
�����$��T�ds,�[�(����"U ��3PGFgAR��a��ٟ(P�G�t53�$�N8����$'���T��!<9<�Ӕ��2�HO�����U�ʪ̃Q� ���'Y�����@�d�K���"�Zu�A(�/Xqu
�߸ ����EG����5�^���>a��֚
�$q��O� f����k�Ʀ�XW)�nU�H��ȃ3���	�U�����8=`�X���d�yir��$'����w֮A��|2A��bϜl0� *�K�*hR���3%���p"�A�BL��'�l�+,�S�|	 j�2�4�������"t)6x`�I��YO��8����B���<Y�h�q�h�����_�t�vAv��7P����h;�tZf�U��*�s� �>m����I�%V\d)���3@ɓv�,��O�t��E����8V��'6����ԥ4��L�&��Nr�H~�UN��!)�0���/�(!��ed	Y�˘Y�Z�#��|�ho��?�'��1��Ϳu�.�k��T8�*�o�b�<����ą9�֕(�O����t�ك��A7jk�����%̘�c%N/��p���XȨhF�"}����D}? 
s��,%*�����6Q���I�+�d(S������!���_� ��i>m��a��Z�%�ּ8t�ӦΗoN}J�iUS8��KVX؞��e�}`�H���J��m�� \ *�b���	ܣT��0�'�Mԧ�Ob�����|�E��'s�́"*�,JΑC�̛}�'=���l^�y�D$y�M�2��x��'��M���%g�q�bKC�dTyb�'50-�'I�-��E�)����n�lhJ�g}�V4H"�]_
���I��yb�P�db���h���z�9����6��K�C�{B��rCDT����	�T :5y�/�(n�D5C�A�k���d�5�f�(D�ϔ8v(i`��� YQ�`6}��NMy2#UB��eµ�?�zm����4�]�`uJ(ON���	�/ד(#����Ú0~�×��B���b�|���$����f�>Q��>7#_r`>Ib��Eg���Hˌ"�@��	�NW@)8W�̟ �f�jp$�:'��\�T�৮J%D���p�cV�32^�'2�'xrhP���j�'H�1K �-m�&\��S��*M�L�tV	r����Q&�`����"�I�#��QЄAI�g�dI��
�e�"�O�� ��5K�y�`��L�0t��(k�]Pg������V�V,����V1+e�q��?��gy��"Ad��S<_� 8$@Wf�< �~ʒdۓ���\14t�!F� �l�$Y�}����KS'\��	��fħyF�(<)���k��H����4�xN�|�����Hf6�mQ��#�4���ɈO���Ė�m����N�(�!ŕ�
]n��"AĊE�����6O�U�v��5I�VE*6,��F7�n�50���<����$�^�@�:�X��A>g<j�zq�'���L��}Fv�	��>>�1�O��0�M8}�|}g���\s����I+'�K����f�P�5&ƕ������PxR	3��$�4�� ��<˔JF1��2�@_��bޓ)d�O�`�L��]�9~�PJ�������A�?�C�I�D�~H;@�6��#Cg*]N<�P����C�D�':��'X����)(�O�2�;cH�O�`(9�k	���H�`>Ā��؎�$�*q�4�6 I�9�d8(#���LWu�@b=}RN�A�9��'gܤ�(Yǐ����Քj�Z��'��1Y� 
�\�V(�[%x�'�hh&�(� �EC��Qvޡ��'఑yu�ӻr�@���aY�P�8��
��� hm�ъ�_��:�X�+�@ ��"O:�Ѫ�#y�l�Pkҿ7|��Y�"O�b�0�p��C	
xRN r "O&!���9r���pf��C�$"O��4"�/���A����(��ܨ�"O�a��_�T`V}`��~�ָQ�"OB�y��, \���m/2�K�"OP]�ԉ�!�`�P]%I�X\27"O~���[�B�̈́z�	e�V-!���Z�LQ�P�
t���y���%!��WZ1�B�@�T6`}3�M�,�!�F�(�T% � P��r���!��"a�lYQ��<3��z%m ]�!�V�@��p���� ��V `�!�E�����+ >�HڢOJ�R!�I�Z �������\�=��߆x�!�d�!X��c��.���խ�9h�!��AM�$yq W�b��L6�!�$Ռp��2��5��!�wK5�!�J�LQ��"0�^��c�I6k�!�D�y6y�f /"���CQ���!�D�ZbXD tc�=�4B��.t�!�Y
}���r�J&{ʎ�1��<1S!�0^����L�.��\��"��7P!��UNu�������#�"X�
H!�w�2 k�"Y�\��<���ƥa��DH�6����/��g���y"���o�\�0��>4��:�<�y�DQ�~���E 1<�(�A��y�畔Qd�뗆O/wb 
�Ҟ�yc:A_��X��J4&�E� !C��y�n�8J_Xuc�!���hЍG��yK?_載Xv�Ω$��Xxfg$�ybf��1���1Rl��dXU�S��y�g��Uh�5�4����z`	���yB��V����+�.��=��@��yB�P3S� K�m_nf�`�E摿�y���)3�b�z�':ˬ���Bٜ�y!��C%$=�kQ>���a2�[*�y�Q���䠑��8����cM8�y" ����Å� 1���-��y�C�%��1�`L	5����cL$�y���7Xƴ��� �,xff؋�yR�R�02F�����wH>��1�y�@�0h>����M�v�ґp���y2S4a%��%�)8��SUC��y�-�.O�X�%��,o��tγ�yR����<�;���&]��"7����y��T�K@���re�n=�h�����yR*�*�<�ٱ͇�m�p�f�đ�y��ϭLM�q#�Cm� ���/9�y2�Ҩ�n!x��.QjuP��[��yB���!"߻;H�[GGV3�y"! �E��m0H�1�H);g"���y��:V��'�0�!a�ɗ��y"4rM�w�ړ}I.�穕�y�X�k��*wb��#� [���yb��'�
08U&�"n`��!�yE�u��@Y�j؇-�d�;�oҨ�yK޺6k�1��-/�\1q�`��y�i��o%�48��+&K-"��'�y�[pQ����LH[�K:�y�AʢO��5s�b7<��xQ
���y��J"Z�x9��!.��0��ƾ�y
� 
���z`d:q.0B��0"Or�A�&ťMl�cB���$9d}��"O�Ձ�ȁ�!��a餀HG�.6"O����@ʨ�� j��y��*�"O�`�t��.��������t�q�"O��JE��j�=ªY�'] ɢ3"O�@�!�g�t�r�
�j|�@�"O�`J҈�{FМaP��?k�4�"O�a1Ҫ�k`rXq�)D�?K��Rg"O��"���7Z�꩙��	|5|��"O�����I�NXؑ�fH#M��+�"O��d���B$�9�ͮ~�r��""O�����S2l�A�@�O��Hi�"O4��Բ�X|s3OA8	���Bd�I�<Q� �+s��j�%��#��9I��UG�<�F��Z�(+F#�+Dx*qAJGH<acA��2	y������k�Ɛ�(!��2iƄ�d��Y�B0��U�"!�dұsC�ܫBf�j�Z!��(E!�#I�ddb0Ϛ�}bm����`,!�Ȉ�$��Q��3^R�,�P(ѯB%!��X�0�t����-$����	�U!��H�{��
���$`9��Gs !��7r��(�F�D�>���(ʴ!�d�[��� �:*F�(��D��{!��_�s'��Bk�ACHp���*�!� (=p�P�L�M/�С"Y�{x!��A7p��tT)�,)f! �|q!�d�M�V !Ӌ�0l���`!��RX!����>��0EW�	j��2©�<Q!�D�%@�0űA!�V���	�	�,�!�W�d~f,R�L֟-w�)Fִ=!�����@\j^v9+��/z8!�J0P��x�6E7�p$`���!�D��~�ҩU��6B�=aC�	��*�S�Ot�Pc�i��Ӧ�衤
�����' J�Y�Z TԒ�i�<T�����'#�ps��(&��␎�$5��r�'sў"~"7䏿R��� =#�.(�'QF�<9 I�����bO:r��@!�	Nz�<�E^�$d*��'�8pb�ط�^<���R��<�Ԥ�.�FE��d�
x��<q�-\O��Bb�]3Tn<����&.-�s"O�ZD�_��>ũ&$^Y�P�s"O�`�儼zW
 0�āh d"���I�O���K� )u2�!1�]�rj���'Ȫ�NF����p�GlT����'Jr��W牖!;���W�S�1I
�'e�X�R�V ~�bɇ�߼o���}��'��kF�_8Vݦ����';V���'r6�2��5�d��	܆A1��'��ݱ�@ȸlF �b�Xo8�ݲ�Oڢ=E��gN�L���ʕ 
�(pz%91�(�y¬[�}br�D2�t[�oͽ�yG��%@�YB�W	���ˍ�y�N�J�T��!�ƔA,p�$�ؚ�y��SZ�ty��%�0R�4��0�y�cZ'()�F�Z��Pi҃��yB�M��,�W�ɺVtDEP�̆(�yr≍B��3�h�yjш�X	�y� �<�r9���	:��`@啡�yB�Q&.�n!�5���H`��y�e��G Z�ڐD�"���7h�4�M����s�\Q���B���W���r̘"O� Zd3�]�S�8���: �F�q�"OR��L�*J�����΃,�h�"OZՊ��*sˌ|P�螪*D��O^�B�'�=Dl�AMO��2���9D��ș5l�J٫F�=x���E8D�ԑ��Z�9)�i��`��r�Hm��G4D�d��N�/(t�
6P���2s`3D��d(��*��E
g���;�`��9�!�dTRu��3$�X�g�~4	� ��QH!�D'A���A���0֨P����|!��\�$����ײ0�r "��ͅ)!�dD�mr��P�<{��my@`_${��6O��۠���U	Lh6�F1�ر�"O�HTe�F�0�݋��Y)��'2�DС+��QAf�a��Vxt}����v�E�0��a[K��F�^-�)p;�O�O�%$�98��y��C liR��2"Oxp	D˝%�fD�Ǉ�X$I�"O>�)�n�u�ě%L�c���"On��s`�*y���K���q�"Ov%h� G������] �"OE3�lŘVf�@��L�,��"OXI����1U$�,��
����"Op��s�޻DWZ���(Crh؝	e"O�$A�!ڔ&��M�#(�:{���'"O囃�>���Ц6����"O�)Y0/A�P-2L�l݈j�x��f"O���@�`�¹�7��36��`T"O�(����#tlJ��D�grꄡA"OL̰��J�u]��p!DMx���r"O* 1	B*?�0��I#g X�"O��	Q�^�R]�-�����r�"O܈�%c��S$��iD_<���H�"O�u���Z�t@�E��`�9�"O���K�� ����㌫-%�UA�"Oj��� M����W�R�N	ƙ��"OV���/[V��$fT����A"On�s�dеz
�o�S�L�
A��"O�0�v\D�3#�R��H���B�O5��"R.�)h�@P0�%JG>|���'�8���OۥI�T0¨T�)�(��'�rT����5�D���H9)���Y�'��Ճ���b��Y�I8.�J�'�P��#	 �Ի�K�O_zX������G�\A���6�0#a���B�!��+A��a�H�?E�N��Ao�,�!�$Y�xj�,��O��a�#p�!���)(ݪaꟴe�XUi�k��=�!��ه^��9"C�0+z�d�����!��G�|Qg�I��l�uK�}�!��B�=���q��4����d
�*�!�3SE(X���\2f��]�i�!�&I��]����x��b��-V�!�Ău��4�֏Γ ��@�^�F*!��=ּ��֙E�y��k�!��PeTX
f��a 8��!���sJ!�H�}�̉!�j�����Z&#�36!��A�z1{�E$+*2m����_7!��{�&=B�U$2�u���V�!��QƁ�w�J��"�Q�{�!�D���D��dLy�x�RU#A�#�!�d�6"�h �A�u�@p��/�me!�D՗VV�@K4K�?�������0l0!�$ق]���{򂀈EYh�"��B�0�!�� ���Çэh[����K}pT�2"O��0��Fi \h� ^�T\��"O��Hڴ��!	�(��G"O@�#��׸���aƁ΂: �QX4"O� ��*Cb�Hh3�J/e�h�G"O*Iq�D� ��b�kda��"OhS�(�'~�J�i!M�N\Y�6"O2U�ƊR	v���b�2�"O�8Xp���>�(�0�b��;���s`"O��Y���;MX�!*�`G�]��5�"Ox�0�NV8/e�T��n�� ���"O̸(wA�9�D��6�<W��lJ�"O�(&#�:�̚��­c�P��y�W2���K��^)!�fAM�y�EĶU�ܡ�%��>&P��r�N\?�yB쌥5�x 굢R1�"�0�
��yR@!	���Pe�����K�yRc�0�aRs�W��B��j�&�y�ƀH���A�.�V�����C��y'u)���P�G��r	� �L�y���5��}!��.�d��h��yr�؝G� pA%�df� S����yB��,L6X��l�O����#�y2��L^�����F�W���y2�T�f�Z
��@�� ����yr��!����H�, 2�{#�Ԗ�y�CC�S>�Z��!3�aK25���'�z%R�%�<[lU��J�2�*�y�'��U`�<��f����@�
�'�>|9@+�So�1�d(�)
e��'���`秙u�����ߓ�&���'��)���:���zt�2̌,��'����Gݭ~;�)S!���֜H�'�p��e�H�&9Z��`�$K>mj�'�d�H��ن"�5���}F|�q�'���	r��0�����Y6x��d��'���8S	�m  ���̀�:#���'찑M�)h�h���H�I-�,H	�'�Ԩ$��D<FP���
�w���:�'}"�x��Ҳr�E�F�U�m|��'�!�G@_0J���G��m���'xf��%i�~�bA����s�Bx�'�H���@ (fSE|�z��'��@p �>71�p#d�V�`bu�'����F�J�F�#����_܊���'�H��%F�8,�\�B�n�� 8䴪�'j�u����xo�Q:r�δ/V��2	�'�l��!�2���(��2=���'����Ƃ@�U�d�N���'o�D�U�/HS���6!A%v,Y�'ܜu�N =����D�D���:D���#O�&.��@u+�P�7D���u�сqiz%h¨��0ּ5crn3D�󗈔	Q"d9s�Tȼik�-%D��:�.� :H����Z�zĹ�P#D��po	6]�΄`�E(~R�)�!D����j�\h�b�;Th8�@ D�г�����
���g 7L�:�3D����'�&�ѡ�
A
�e�%D���Ge�/�>dsf�H�_�� /D���o36@@��F�q���Ҍ.D�H�!$�-X�xpZD��Z/`k��,D���<�x��m�'#�ăf�+D�l�Շ�g�R�{� m�ّ�'D�� ���񅟑abjM� �+�l�Qg"O�Ya&��z�p�
qF#]}Č+�"O�l1��?2�}k3�ta<Ъe"OX}�v!�2Mi��T�oHR=HC"OT�Hă��W��q�RfɪZ� ́ "O���"��zA鑯ǆ2�J}
�"Oj��4�¥H�<��ڶ<Qx�6"O�@����#ZpV́�&Ѭ?�Dz5"O�P�Avl�8JхŌ(%�8��"O��#���9��R҃v���""O��a��N�o�( Ѷ"ԪL�d�y�"O���"��߸�RQ��X;�AZC"OH�c"�AZR ���pʐ"O�@�F�����@�4&Ҝ< u"O�a�w�51и�T�U�G��U"O�ݫ��G ���(0�D�b�6���"OPx+��3X�D��҅� Hlp�as"OԬ���ߩ��I���v�t8�"O8�@��L��Ik�*C)���T"O�DpwN׵#t\B�	M��iE"Ox���@a�
ѹ�G�%rtT�y "O&��R�Z[E�H�s�]i`���"O��1oc�.�bD�>%I ��"OV�%솼T^�
�c	�a����"OHD3�=5��hā�+i�򨀂"O(�J�`�$]��,�᠌jN(�"OT�*�j�	YrDl#� ܎UA� 
�"O`Q�u#��Z@c�oT�w���2"O:0��J�M�d���8j�ɨC"O�(�!}Y�1GjìU�e�g"O\�q�	�v "��a)T<U>�ْ"O�ɹU,��4M�D�چI7�-B�"O ���*R	mۢ��c�){�]�C"O I ��G�	lHD	�"�:r�@0"O��!��^����� K���u"O���Qh%6Υ�� �䦉�"O�J쀿_��y���]69�"Op��G�n�0#�"����"O�I�b��aT�b�^�xt2�#�"O�G+@UU��p��ɼDs��Kt"O���*��+ ��c�
"U��S�"OE���X�7Oq���0M<�k"O��G�G*Pm2@��)X�0Q��A"O��!Υ<$�}[��­^���X�"O���E�͕��9A",G�<�H2"O�a2��TXؑ #D�}L}�"O�M�ƋP�Y"u�#a��W ��X�"O��	�H��K�擇'����a"O�hs'�ÿ1Y�ȁ�� �$�$l��"O�ݸv��
gr╱v/Ɇ���9A"O>M�䭀? 7�	*Ĥ�J���"O�LH�LQ1�aZ�D����k�"Ot K4fԫ+�VȘ
��! �"O��u���L�1�&{�(�z'"O*�q! !Tw�mi�+�dL���Q"O~���G��h�@�T*wE����"O�LbPc��J�Z�g���Y:U"O(�
���7A�?8\p!#"O&̚#��u,Ȕi�.��W���!"O��(Vn�=}�z���L���U"O�c� ���q�"S�""��P"OE��(����cU>c�qJe"O�5�s�լ�XS����wqV��"OF50PԨWh��0� �\�.e��"O� �Ԋ�	�5YhHA7��^�8Q)0"O�Xxbǽw�iق���u�]�""O�56
�$\B6���wBRp�A"O��H��	ۨ4��M�8[F���"OlHR�Ԑz���cӞY��X��"O��rAg�@���c"�&�9�"O��C�J#��p�fW?Q�Z���"O�P�4�Ų;�$���G���M�"OD�3�PL.�K�-�'Ԃec�"O�h���AE(Q��īV��p""OnM��T�J�N�@���P�@���"O��0&�\K̦P�ak�z!��Ӌ}��2��DSǸ�:��\h!�	3l�D���Ū8�X-bIE+�!��U�E�J�qg�	%�N��/�!�d]8]�<�ċ;q����0��>u�!�䑠k0�׋+g*�����ua!�ړJ�B���
D�C�0e�Wf^�o�!�DLv���K�ʗ	y�������tG!�$	�
QD�ӧ-	9l��x��ňt�!�D�Lg�K׬%h���L��Ds!�\=e� 0���=+2��bfI�'j��b�Cdޕ
���Z#���'�J4AC�<K�q�P"J�!�'����d�2u$pX�K>?H4�j�'Ӹ�I�'�� �P�P0�@�'V���>�a`�R|�L�A�'�bٙ��G?�01 C��T��
�'����&�ƞB�����>�Ty�
�'X8H��e]�F�=�6��*5&��
�'�l�µI�J������Ď2�RYP	�'���iЉPH>�����u���	�'^D䫗-Tu�dz���u�)�	�'��}�&N��3��0�u���s9bTQ	�')8%���J�R=�$��3�,\+	�'b 9���qp\���נ&�����'��@���Inl�󏉯*��EP�'�>�@D/�#ɶE�܍%4y��'�*�	P%#���u��,$4�i��'ZB�8Ҫ��Z�$e3$$ƫ)Xİ���UV�{�zL�hį�%C̪ j!�$w��	�R�O(�����҅Y!�̔*� �;�@]0ZO6�×�T�no!�$�!:
��26,u#�A�EV!�$
��*ɑ'��32�!�fֻ/.!򤋪`֍� G׊R �=�veE
`!�d�2>��1�f�>jo�%Q E�#.�!�Dռ'�v�AueYXv�3��:�!�D$N�����;>#�L#�ĉ��!�d�8~6���!A�t�"U��)�!�I�9��,J���\�2|����w!�dI&
�B�Y$�U�D>FI+!Fק!�!�<W}�p��Z44%�DH�k
�*c!�߂Y���u�8�QajِH!�D�,|��C�TP���)\6XG!�$ٰP����[���d �A�48!�dPB��q�)�N��q��EE�DT!�����6�YֶEp2kG�?�!�d�=��&.�W�0�ɴ�9!�$y� ����3�t�!�.OB!��X,�Qi޷��LI��ݕD�!�D�C:\��Ň�b�J8�B)�
�!��[�X��R�	)Z�j*S��
!��՟T�a��8�ƔI�@7�!�� ҽ����8��yh �	�O�p8W"O|�'[�UpVX����B�����"O(Izu�ҀTI���q $o��-8�"O���*C�'s�%��T�y���"Ox��F�:Aq\��F��
\��:�"O:�" /Z<�TEa�N@#[F�aC�"O�#��R�#{���Ǡ:	�;`"Opl�2���u�,y�#�)��dZ�"Ot���ɮ@P�� ��^0�v��D"O��A��֕FYN�{&�&;f,��"O0 ����� B�@[�
t���"O���r�L &�>�0��Wl	W"O�=x�'������ Ŗ>N�x�q"O
�5���q��|H�
82�9�"OF�{��h60��Cݛv�e;�"O� 1��"n���3��21��xs�"O��2sBZ+|��x�7��r���8F"O2�8�nϻ5Y�D+%�KWS�e�%"O���b�{��/Q 
2d��"OP�H�CM3�Ȁ��oy{�]#2"O��7@�(q�ޠ��+��y�h���"O~�S3!�Rx}S	�$�TLؗ"OP�̶ jιsq���"�N�sp"O Y �I�`4T%+A�[e2B4"O��S�!�,V���K�A�*fS4� �"O:��E��;J���\�$@A"OfP�o>��$ĥI����"O���d.	wOn�p �.��0"ObA�$�Si<�u"MD�lȎ�x�"O����,ٝC����wkR�@�=Q�"O�58��|I�!�	4rC��1�"O*�zH�-\Z�`��G��o?����"O�i����O�:� p��&yH|�"O�Y"�N�"i�@���1��p�"O"�
� ϑ<^�� S/��p""Oj��#��&4�0y�R��1q��ҡ"O �9����A	�l��s����"O�9��ʨ6��<�f��"#z�"OZ�)��uv���h� 0	>(�W"O|!�l�KL��th��|�j�r�"OXY˧AV� �����0Ϥ`;�"O@q�ƪռmt����;~Ä���"Ot��WE�tYr��X���r"O����,�lzU�T��iH�"O"8!`��Q�1���_�ا"O�y3d�n�Vtٳ.ӸSF�0;"OHa�DꌿL�BDpG�ÚUdе3�"O�M�ğ_F298�ɬ��|K"O6� 	�j��D!S�� F��ȕ"O-�1�Ĥx�����Ά5��!"OZU�P�M���1���`q8��"OX�ס�����(f�l�s"O�� �=�Z�	QFU� ]�= �"Ot��t�UY���[Uo��t���z*O�p�!iLq7jx�f��l9z�'F��+��М�HQoW���@	�'�0�BeS�J`�؉@s
$A�'3F�SFF�>��O[�Z���	�'?x�9��
4X*L�4����Q	�'��bg��,�Ȁģ4+F��'�r��h��y�q(Z�#.���E�<�#]�YT�α~��Z姊I�<�R�M8�De:���-7�6���L�<���P �Z��@I�J6�r��LI�<� D�Z�gF�W�"xb����gj�,I�"O��Z��ݹ��hqKY��<���"O>��B��
�(�ɦ���N��@"ORLsCCܺ}���*=�����"O�7�S�a����=s��"Ox�vY��a@��H>cr d�"O<�b��F;i�=���I����E"O(��T�	~,�Y|<�]��"O���1-/�6�!'��?,��{5"On�)�mè+��h�dh�$= l(sV"O:��.W�TАY�T�X�/���"�"O �	r�o�z(����s����"O4�;f�:5�1��'~��"O����g��A8W�]$k_��`"ON��g��̀b͸M��Hk�"O4aDʂ8F7"����	W��8""O�t�6O��,-ٳJN�����R"OVu5I��Ӷi*A�~���"OD�"��
4]\��qkW�bBL� r"O�uk�|�l��Ӏ� O[N9�q"O��2VnK*) �*��f>�1["O U�ƅ"&���Oٷ!'Z�BQ"O��Jchźo�ڌ(Q�W6 !hX"�"O4�r�Ɛ�F���bT���2��!"O� �A<=����G�3�(-��"O�Ţ��<k�e:�ǝ�S�|���"O��򍛻�+���{q���6f�Q�<��j��)��U��$.g�J��N�<�P�C�.~E�e�
���b�N�A�<A��ZQ#�&�/�-BR��H�<��d�5El=��àg�����|�<��f$B��j��x5���WIy�<IV��&X�KGɍ
/=�a�a�s�<�� �)j4���gK�2���H�W�<���¼hG�A�^�Y���2�(D�����_�9(�5
�� �����/,D��R���JH�!�A��J-|�{wo(D�l[�j�$4�B�CJ[:r�R��U*Ohah���3T�Փ��S>R��w"O<MH�PM!�-+0l0Ӥ��"Oh̛VÅ)D��kҐ"�l�Ä"O��k��� 1�B$R�L�W@9h2"Oڽ��kڛs,N�i �@��%�"O�ՙf�+Ɔ��CI��w� mir"O�9��o��l�4�����|Cb�#F"O�� �'È�zM��>)D%�"OΤ����E���XF/�=c,N!��"O<p�s̔	�,4���L+&�q:�"O�E#T`E��D駃��T�ra�""O��h����B&���$#	�t}�8�F"O`!��Δ�H3���gb�=:0�`"O�x��E�m�� ��#��Q�"O�|X	�RՆ�{�N���8�y�H�K�\�c�ɞ!����%�y2!'PN�Ih�U��l�!cA&�y��-W[�L��͠����Cv4C�	�0�~�hE�K�:�"�P��B�	sR�I&I�P�h���B�	�h�ryi��	=��0�QKA��C�	>��PAs.�!a��|�PkR�H�pC䉠+�R1����:pThqvfO�,�C�I�'(N=���2x1zw�K��C�ɳn�f��T�d��K��SR|q�w"O�{��!�7	�*
;����"O� �jQ�E�P�H�HЧD.S%^��"O@%�eMCWĸ�$i�/D�#"OX<5J8oFt����_�Z; ��"O��R��EKN���C�?ޠru"OD�pA���f����C�L�^ib"OF�D��G��z)���$�b"O���W�TRT�j2�N�1:ZT$"O�,�5���9|��ps�$Z�
�"O�T2$�[4@�:y�(Q���"O.����3p��P7G�\P�"Op��W� (m'd���~��%`�"Op��F�x9֍h�N�Y��Rr"O~��qF���/

����"O����g�KB�r�օ^�8��3"Oh�v��(mu�9�����EB�"OzE���n������CM�0�*O8ݹ�;S��2anĕG-�]��'#��rd��9��R��1�'2t�[���"nj��G�*>��ț�'�<T�TGI>ό��c���0�l�H�'�)*��pJ�@F��.���C�'����Ύ��)C�]*vd�q�'@�p1�3�5���8#�l���'�b����r���B�.L��S�'w�i�3�U�0���Z���hL��c�'�R��� lDn]�ACPҶuz�'cd����9Hk"h٠*�;w�|ah
�'�5@�CL8�����rF@�
	�'�� ��W=���O�V�ġ��'%�U(��$�S�#��F�h���'���!��)w�4ͻD��:C0ɘ�'PU�Wg_�Y�&����CH���'X�`@%A�==��S��&�p��'�t�cԆG:6�8���C�
��!�' ���K̸hX��RE�#X�v��'����� �@���Ҳ�(��'��&ʷ�f PA�U'����'����@.ɸ.=>�Y!$F�U��'C�0Pkδ^�ⱂ�܈n���@�'��� ����9HKS��R�2<h�'+@1�t��h�4��%�L`2�p
�'d�!�f�L�B!�1!!in�
��	�'l\\�!�˨<~��j�E0g��$�	�'Ev�#�c�=_��D@�����N8D�xӑ�Ы�R���l]-�^9aǆ3D��:U�-�2�15I p7���1D��k�H�(W2�ШS��J��A�+0D�<��G�t�93�jӘf���H3�ON���<����re��8����k	��<�V�����);H�D���
%�ȓ/����m߈b}���*��/��ȓkp�)R)ϸ[�N����:_����g�6	[ �-h�lk�&�4f�l��+�� ���$CW֑��O�::D�ȓV�б!r�B=>�`UҳM@�S�z%��}v����N9l©	���U�I����Yk���0��2+�2E����H
E	i*��	����	q�Ѕ�ȓCk�щ�g����S�N 6$��Htp��K�P�Τ���Gv^�ȓ7<u�4�d;��3���f��ȅȓ� �զ7gvHH��@�g��m�ȓ. YBJ oרh9��gU��ȓr�Be�e��"��ĠsO�Yü���S�?  ,�'�2� U��D��z��}��"O�L8��f��Y�� ��B�S�"O ���vrd Fe�2;�h��"O�P�4��m��HG�/sm�<
�"Oh�Jҧ�!����)����Xg"O�u����$쉐��>+G����"Oh���+� �ɰ�˺:ĕ�S"OZQ
�['"�ƹC7w���@"OU{��D5s�3�FN!BdbIJ�"OD��o�F{�p8���%���{�"OH=Xc��d�ؘ1T��)K��u�f"OT�F�6*�%�!;S�hLRQ"O�� ��_����U`��(��=�"OT]k� 	�dϤDIt��M���å"O �0��?"�������)7bI7"O"0w-
�V:D��"��4�bt"O֌�� �j(�Ikv+,P�c2"O�9	5'�=w*���)�n���p"O��	tnЃU4�������c6|�u"O����'�1sl��UR8��"OH�Dc�4��5�4�J) J`�""O��
v�B*��uҴl��=O(��"O:M�-1:�t=[�˙h�H�t"O��P�٢8�ie�)Z�p��b"O��j0σ���B�Ƀ�Y��@�g"O �1�
��d�ӈD<o��%!�"O��Iw	V��@]��|�J��G�IG�O�@���MQ�y���zK�/�(Hq�'���*CȘ,U�p@�C #��d��'����%�D�o_�`3&ñw��P
�'񂈫E�'�J�L|^�T 
�'�n�
�A)>*艣
�~ʭH�'��5 ��@�Q�ܼB��V��'�N��E%�@^\�u"��)�<��'&B$�Vg]�9l1�d�"i�y��'��� ��*a�ABt� M���'�(LɢA�׌�g�Ի����'*`9S�͟7r�h�	��U��'[���E�\�tL����,�"yj�J�'�h� b�����
��`�X���'�>�I1[�jA/Q�q�TE����"O~ y��<��!� D��S�,@��"O�A�Vk�X0q�Q�ny��"ObxE�&i'޸��ʂ7_4E�#"Oh	�P�"P7p`*���CL����"O-+�`@)�DT��(�2/�"O�e�9y�R}�0GG_Pvm�!V�0&�ȗ'��k�@�0��+��s�K8D�l����a `#s�� �JZ�G"D�$�!M��4 �̑rLA<xk>�@�n5D�@�]\A��7�fq��{��5D����T�Z��U�A�F7o��y�6 )D����@JT�>8rd�C	cʸ|
�&D��Hwe։�����A�1$`(aW�/���OF��>��N�@����@+ �V��P..�d1�Sܧ<�ŏS+��d�r��l���ȓ
�����Y+Y��,����>�����A��2�Y�h����g�K� ���|%��Nٕ ���M�TO���y�Ҵ"4�2����FN�%[s`ȅƓh��ۃo� �:2h��@��H#���<ړ�y"�.���v'�!x(�2�f���y�K:W�
��]�W����L��yB /P���+�Ώ:YbT8�瘟�y
� �������1,�!�А��9�"O|��׆�2��}�dT�3�6�˃"OZ�P%�
=iɰ����:t�j��5"O8\�'V�G�XxC��!�(�cQQ�4�IW�����U�Ü�"h0QkA)�2���i&�$!ړ��dS�G�!H�Μ�Ĉ�E��q=!��@=~�L�����Ox�х�01�'ha|���k�"P�Ʃ٬,���!@)�&�yU�9_��H�.�v�*���y��(@Q{ �׼�X|�]��y""q�P�2k��f�$�֥���yB��dC ����`�ĕ��J#�hOh�����xu
�HGNƪ=�>,A�hV�W"!�4��� �,��
����!��I��8�F���O
8�H�C!�$ݢU����ᏮAV����'Ɓ�!�� ~��c`��-���Ԇ��!�D�4<��v��e��T"�/� e�!򄀥U���s�G�@X�@� ��'���'���6�U�CA78���4E[=kx*T�ȓUr��8�D�:
�J& �H�,D��E�`��#h̀4�0n֠A�����A#J�,���'��_N�!��M���չ Jei�%�j��Ƥ�RdA�ƖUs �[�}�����0�tm�@ňtdq#�͊%ݖ�'<ў�|BV�F([Sļ�f�-u0= ��[{�<�G��HIR���P� 5��k���n�<����n �X�t��-"i�0�i�<!�\J��"ǖ���t0�Ge�<1�BK*0^��`�\��ݒ3l�b�<AdÑ3��-�0�����
xy�Z��'��F��/G�s2�� ȥ �v��Dl���䓐?�M>���͔/7F	{2K��`�r|r�f�!�D�`�PХ�#�H��M �2�!�� %�1�a�:
�vh���2N'!�D͈a��1���#� vʗ�!���:cd� 8 I�C�V��+ �Py�J2{��)`P��XZp�i�=�yr͕%���8��B����MX��y"��,B��9��Z�������y�L�apP,1#N3�&�#�L� �yb�Z d�&�IQN�&E(�{��Í�y��ߙ�0�˔�K�%^x�kE	�yR�Q5>͜U�P��Q���dnH��yreK�B��a
�MG8�J�qQ��7�y�j5L���e��2� e�'ұ�y"���*Ȭi;�쁗"Bl�3f�N4�y�M��
�p��"�3�B�	��D�y��V��X)J�`T�`
�HR5�۫�y�b�Ne0u�P��Hy��(��y� ^0	$� Ƃ�BV�+���*�y�[2�z$kAhP,~b�`�C��yb�Ĕ@|E�c�Y5& eC͍-�y�g��d��� !����(@��y�猼F��<���#�BH���X��y�oԯ� ��(U�ܮ���c��y�@ڬxx����Ix�>)2F���y",ƺYkfMB#�I6*�����W!�y�Q-G.���c�hH��B��y�
<d3rQ��aƑ~?H����yi����9����y��-)%����y�f�+5�0��C(��z��+�y2�S3f�^ճ4 I5 ɶ�r��<�y
�  7�*��$��*J 1@"O�(%�ӳd��+qBZ$/	��*�"O��Sħ
/�����[�X���۠"O�KU�$)4�C�F!�r�q"O.I��ط/V}����G��y���y��8`&\�B.l1�'�y2� ,>�VhY4�$�����y"ŏ�)z�D�5kv���V�J+�y��EP����g�Thq�H��yb���;\�ʲ��	��X��y� ����.�x�(�7����'f8�Sb��z�R�dC)�|1��'=��J�8�L�+D�0|��'D�(̴D7�@`��([V<(�'(�y*u`�4֤lk���E����'wh��"˺vLdze��0��#�'3❃f�8wT%	 ��9�Q	�'��U��NW����*~��j	�'���4mX�.B��u"�
&���p�'��������%#�	M4��'���BD(��;�zPkTA���l��'��PG�]=-	��ؐ��(=��'F��h%6DȘЀ�Q,y�n!:�'2͡�&߳qh�	Y�nw��x��'�i�喯f�J�h�X�n�B���'��ᷩ)t��(�K�c�9s�'.�����$!x�p��6Wmڨ��'m�r.�>:^�!�s�TJ�d�r�'�z����F sz��aQ0L, �'�����.@H��D&�"\�r�'��	�j��Lz���c�ͽQϠ�J�'�֔2V�Lk�v��g&K����'��r��\�`�씫THÊ+��Q�'��M��kGcK2m�CAz�a�'����'ʝ�H:��& W#_�h��'���P�ļ6�^�iE'�[�����'�"�*f�B����Ͻ���	�'_�Y��R�} ���f��O�a�	�'�̥*�f��^�Ș0ᐨ@����'"�a`�,{��� `E�-N^�)�
�'�T8g�V:S9$�S�@կEUX\�	�'~&0���V-#u)sM��'���
�'s�P�D��.��1�g�)Y�Q�'�xU�0�i��{�GW�� ��	�'���P �
-j�c�):�pQC�'����G/��ꬊ�I��hx�'���s�l�9i�`[����}��tJ�'�0z$�|X�� $>|&�d��'�n�;"���|_p�p�C�oeX��'��{��ɩ,�^��Wfǉ[�l��
�'*,8"��X�84
�
���$���8
�'��DP�ɑ)<բ݉3ΫM��E
�'
��ʐS 20���S�G�t�	�'G
 ��fC�"�K2�D:����	�'�(H����ݫ���:g��y�.�x X� �,#��xS���yb��S0ڹ�bN���>}z2�M��y+�7[�����N��a ��y�!��B7�փ	>����ƒ�y�)�&,�J����!y�J��g�1�yB�цg~������tn�a�7��y�41ER�h�Y``�І@���y2�R	:&�A�sI
e��	V��y2�Բ0��mӱL�Ej�����ߗ�y
� �� ��L�g�.|�`����HHa"O�Q	Q�J;�,ST/΍Bf)#�"O��;c,�v���Z�t/~�1"O�q0U)��)7��K笏}#x�6"O��0ChN=M2�uz�"
9*�"O�Qq2��b�� -��(��QS�"OxUs��ԑ��µ�!�Eф"O`L�$aN'��$��j,LF�<�B"O��3!Dҭ�1�	��B���W"O�,�%Aэ4B(+Q�{ѴeXU"O�p���Ӈf$<�qE�P�7_��""OR(z3+֩D,4E�������y���bE�f��3�����Z�y�EHz��(S��(2z��bF�y�͚2c�����Aq2�DX�g־�y��=F���]$n�ڈ�"b�;�y��6r��;e�
i����ņ�y��ӭW$���K�aՎ�"����yc8��@�5fO�R��4����>a�Oe�g�� qLƭ�5̛�#��Q[!"O��s��vŁ5K]��v�X�"O��Q!�G�P���ߌ+���Q�"O"�P���)q�^ YU���f)s"O,q�ү�W�t�c�Q�a
PT!f"O.i���+���;VO�!,\��!"OxE#"�Z6Kh^|{�Q"YVX��'|���<'���gk�&�fa�d�i!�dQ�4��+��g�0<#�-��Y]!�dʡm!6���ʘ�Ҫ����\!�$�8X��iU���}r�+�Pv!��3F�r�T��:-�~�+Uj��J_!���-?[� *D��=ʦTz�HʢG\!�[(2�>�T�� �0���gO:Y�yr_���'�T�`g��"oP��D�)c��q�	�'� �9��$o��8�K?���	�'�����Q5d(Lm[�㈟P>4u{	�'��`p4g�n8�9��<;%,A;
�'��9�GLC.hx��#��tg9D���e���k<�P *4N�x��$D��5N�J�R�2���&�6u��/.<Ot�D4�I*74>�xc� 2�^���
�V�B�ɕX�2�Rab�d�h໴"M�b�B��8|U�A�@��k*�$����`C��p8UU�٭Y	�A�%�9`�C�I�'b	
Uϙ� �O�lZ^C�I�o� ؀#�D�����L8s[C䉆A���AgɟT5� Ap!���T�F{J?}����`�0H1p�N���.D�ܘS��"el�8!RF�����
(D��E�$i�p`����N�lA�l;D��0�9T�M�Q���	Tn8�@�:D���K �i�:D���?<�&����9D��� �l \Mi���7.�Xi�V�;D�����]���N.(�.�xA$:D�X[ĈS�T��(��(�O�Ꙓc$D�y��O%
O�SV�D��aK�m"D��ٲ�L�<abǬ��u� ��5D� ���),�رʴ�+%��$*��0D��z��ʿr�]��	�6��ѐ�0D���w�1�*�b��]�UZӍ(D�pKA��t��s���b�~��J+D��	Q�Q�7���2��7~YxUD(D��St �!pj�36�^�E�'D��!����:0\j�����t�h�O3D�� ��)�ؖ\m����?D����"O��٣I܏�Wl�_�4�"O�L�Q&H�o�5����$��- �"O>�0A��o�$�q�2"��u��"O ��u�_&�Pqb�GPAP���"O~� �b!�F�C���[�"O��# �L�D~*G�֭k�h8�R"O�ѪcT�[D��{����&NhPx�"O�m����
��E����v� �S"O\��GE�v�!�φw4\��"O^l)t�^ Z`,
��_S�T#�"O�4 D/��&���2� Q:Ұ�"O����'B-9�`��`�ORƸ�d"O �"�/�� ��b�שX��� "O�@q�I>2�8e��	�\av0I`"O^9R�E

p�#�^�ݘ�"Ot(SpŅW��Uc��U*0�� "Ojy���4�A�b��< �9"O���M(h�(IH��Y
H ��ҳ"O	)�їj�0d �X�*�s�"Ofi�-�6$fĥ���C���"O�|��P+3�z��c���N��8�"OX\򦇉�&��k�.ALl�"O�� J�5:�PRB)�O$����"O�� =*;�Y+�
D� B�S`"O<�pK�"���gN***�ݐ"O�ha�!�'5��3���uyh�y�"On4j$�X}MVx�R�؉7b�T33"O���A�;r����فUY��Jg"O0)�'JR�m�8A�Wdlwd`�$"O(�T'�4�x����(RX���R"O2="'oW*Z�FU0����@<K�"O�8�����*�+�%6���C"O\ n��/4�92���?N�E��"O����'ZX���e�|%q�"O��J6F����qç���y��"O��2m
�&%��r�%��@�q+U"O����cPN�!pWjۉe��x��"O"ݪ��zۆ�S�E1?���	"O���'H X_�9�æ˺e�s'"O� ������0��"Z�!F"O���u�K�L�f(	�B�4;8c"O�8�qA�-y��}h �Ã_�B"Od��'���1���e���g�j�C"OLab�k�O�:pj5l΋$�R4�"OX�PR�
 � Υ/���"O���S��T��U��:�V=�"O�-��ު1p�!�7��N���"�"OfM��Ƈ�j��ɒ�m������"O���H�
��� CRu�r@QF"O~l���%WI�a�� �(8r@�j"O�ѳ���$\<�%0 /��ae�"OV���Ò�qJ���+R���S"O4`��"J�2���p��0�G"O�誷��;}q�D�5KL{	f�V"O�<�௅K;(\���~����"O&q8�J�H�p���P�c�R���"OT�cCJ�z�(��xzh�;2"Oʘ���X�l"��T�M$z<��"OMq�Ӷt�����OZjgV�"�"O"-��
��y��"��uyJf"O�ܠ��VX��4 L9Nr$��"O6� "D��8~$-ە@L�: zA�d"ON!��Nj ��X(?��#"O� �h�t�D�
B���s��)��y9�"O���pmߚA��H��(�|k��A`"O�|�b/mqĄa���P-
��w"O�)���Ǆ���jG�_�s"�؀b"O@�Q�o+$�j	�%ə�w�i�"O^!�@ �j�$:T�G�z`~h�e"O�UXPI�'Z~�yv@�b<���"O<���+�]�p�&�ɧA^Yp�"O�H)ed�"��x��CD??�ل"O��#�2ZJ���-4���'"O"Y�GÙ�lH�S��6}��"O$x��=[�}˳�X.3g8�a"O�l��C��g2<�� (S\���"O�lc�O�/V�PL�殒]RR��d"O��24�>�4�yum�TA�e�q"O��:��؆x�Ta!�Z�`0aa1"OlT"v�����@�f؅^7)X"O�ܢ��@�lR`�e��3F*�t��"O�`��(g��d�SFR�zyF���"Or]b�Ĕ zyH���ER�) ���"OR��A�>L�<a'$ל��mr"O��A�Mo��qд�@�|���sV"O�+#b�5>��P
�d�
��P�7"Ov����y3v qe�m}�""O�Cu��N�,*A�F*��P�"Ojhb���J��2�	"]�����"O2��D��~�f�(��T�s�B8"O�a01g�}}U���,R��mX"Ob�3u��"��%��a�~�H�"OD̝�k���� /+����"O(@�&N���H@�O5{����"O8��sM�2�lN��;���s"O��q�(�'��A�MQ�g{�I��"OlawhN�s������YAr75D��{��O��x�P'ï0&f�!#�1D��P@)Y��&���݄q�j�r�&.D�Xx�H�~�l�'�*sr� ��1D����PW�t(A�)C*V�rn.D�2�͔Z<��{�&V�om$EX`�+D�D㤁@�0� 9�������*D�����]~�a��̓��0�[w�'D���B�1�u#�a3^��x��#$D�T ��]awR91 g��Oh� *O���E@�t]���@oQ�!���ɐ"O%��Kع��-'[��� "OrQ
�l
�<m��ĉ ��	1"O��6��+R#n�{���z�"�a�"O�@�L�u���(Q�ɘ]���"O(1sT! ��@� ���Ըw"O�iC��T;�3Qƈ9&y4Ģ�"Of�h�dҩ&�$�e�[aJ(a�"O��R�#ãB���)*j2�� "OR��U��E@`�PN���1W"O�@;�X4E�F��,��|����Q"O
�z���7�tąH6��ݚ�"O��qF���\o�1�$D$M�<i9�"O�͑W�˘p������B�'"O@Ԙŕ�N�HzR�Y*O�4`�"O��A�cFY�,q��w|�F"O.@��
�w�`l@'Dg��	�"O<� b�\=t��ms�I�'vN4b�"O���e%Yi��hA63s6�3Q"O����Ԓ@m��bEN�V�m�S"O ���-O�xB"�	�D>"��d˒"O� ������iPDV�55�3"O�q��+�5|�P��B��R�W"O��� I�"r��5�N�BP��!C"O�0��g�b��zƯR�8f��"O�E�@H�(]�٩�,�i&p]��"O,%;��ٰY�v<[U+q��`�v"O��"%T�jC�@��T�B	ê;%!�D��Ot�!�P!�:Y�&LX���'3>!�WCY����D�9+��"�>3!�H$���0�A� ���0� ϑ9&!�d�f�q Z%o�يA�O�4!��0")�2�ν9�(��#�s�!�dЇo��X��Mњ8�r��v��~�!���bp8(s�"1�>M��*a�!����9f�Ö,�|}!���!��&9�x�����`�U�*+@!���4���⅍�)&L�v��/!��/j�lxx��݅qN�i�e�8!�d
�Yw�Dcb˒�.i��i g�Ud!�ɗdY
��ߡkeZ1����+rZ!�1xD����<|@�"�<T!�>��4Zu��63Į���٬ A!�'x�&q�G�	o,4؁!�
�R�!�U�+�D<�s�\}&��$�A*�!��h�0q��XN%Х(5CJ#G�!�d^�>�R��!g��MR����!��VHe��a^6�,�3�7[�!�Ď�)M&�ڑz���I�"��{!�D<
��ycOX
9�F��g�{!��бo����ƀ��`�3ÂӟD!�d��H
�}a���g����a��?�!��74x������3�	�woE�3�!�X�H�ꨛ�"B,oz��U�Z�2@!���S�P!��$�/3���CV	�jE!��_�Vp�1��vjY��G.5!��h���fnEaB�iCf�XL!�Ě���X2ϝQqv�
����~�!�dC��@3�2h��R�R�@F!���>�����9�ĘsC݀!�D@�,�z5�F�8P�=�p	�^!���s�����>L>�U;s�M`�!�D��R�2���5<7P�� �X9�!�X`�Q{!�$}�l�T�� !�d�9h���N>uz�L���ڛH�!�U��ta,ӂ�
$b���V!�?�N|��25������ՒBY!�dG*F��+��ǯ|?.�	R-W)@!�d
1W��!0�G���t�1�vY!�$J�?=�(���Q�v����n!�ER,�����|H��ڒtg!��^8W�ݩ%-�5b�р0L;]�!� *_��@ǲQ��XǀH!�dӓW� ��O	^�|i�e�7�!�S�
�TZ0��p_r02�O1#�!��͠�$���&K�$Y���c[?by!�DW��D�p���5ڪ�󑌛�e!��K���O?+���k��3N!��3K �d�%X�щ%lY�NZ!�dV2i�p��s�	�lK�xh���\`!�F�Ԩ[qʈ�+��P׈� 7_!�	�0�<�i&�W�z�V�Ȥh��_!�DU�d�+��2�>��*W�JB!���(zLPp��R�F1󆯒c�!�$�%x�
�! E�j�L�ʧ�>B�!�� �,��ݬk�\Ç�6ID�8�"O��h�O�~�%c�E�� c�|��"O��y �?s�&�X��=;t��"OQx�ߙ �ȵ!��ؚ2/"�!q"O�����k����N��U��"O^���M��Pٔ ���>~�fX13"OJ�H��Y1�B`jAi��+)N�X�"O��f�>����e�S$�ј�"O]	�S�w�2�B�g,Km��"O@t�V�G�4�t-h1��1rTNI��"O�5IW�a�Vu��1|��R"O*|;�/��/˒	�e��9�!��"O��Z1�l��{������"OVP[P(��RXQ`1+o�����"O�)I7�!���)��1~.��&"Ob�Ԏ]�7T&�1E��57g� ��"O��҆E�I�qcv(W��.;�"O��i%���T]�Ӧ��"��ts"O	�Ui�b3�4�'��<���"O�0�vG�v�A0�h�Z�P])�"O�@R���ЀhB�Zö$YD"O`�"B�F�li�5)�d�]���"O��9�)��bWd��@ռ/�t�#"Ofp�R�U�|�v���H-b��-K�'��'�剦G�� ��%P��v�(yTB�ɨ��Ͱ$`U�^��q�P�,B�I./��M+��sϲt��u�B�	
�6�{a���������B�	,_�l(�ĝ�+
�;P-M�+�B�	�q�VQ��N�2ij�(���1ۮB�	Q]~ɊR���Zà����J#T~B䉥L+dxҕ@���91��3m�B䉹 �Y ⊔���)�S�ɨ���\aG�)�iW3�Ĵ�@�^l��W$�!�D+u�D���շp�H���!�Dў\]�t�G=U����;N�1O���dQ4f����HL�5�� bA %�ك1�����g̓4���9��E?� �w"��(W�؄�mEH����&+�ā*��ʄ.p���{&��͚4�,Պ�P�&ܾy�ȓ>�����(�DH�kѦ2n �ȓR{Xx��|?d���"��<�l�=QK>���*>��tj!O��{&,:q��%!��^&K��@2�b�+_��R��(�'ha|V/�0P�TI�*	$���T��y��5���0W9[�qѧ-����D.�(O>u"+PJ�q��!��yS�a*D���w�r�ԽA�D5i����!;D���dG�2�hk!�h�i��F8�O0�	r��+b U�1���p���|-0B�I�`�+�O�X8�9�a�/'�nx@5���G{��)2B���J�
�/g�v�K'
�3�ay�(\@��h?p�C�.K�i��!��\Lv��I^�wUp�£)�w5,y�Ea_��	&�X�:�Hc��>I�JP�t�x-��N�D�8<ré.D�k�b�ٳ�����c�5ac���d*}�HB06̐8�=.�m�ClO��(O ���Ɔuxɺ"Jæ,^�,[��ׅ7�!�䓈Z�(b6��LI��)S����!��K�a_�;���C8��Calт
2��E�$�;�0��	N
�I�����y�	ե��Q�2"�/��Ip���� ˄�<��y2c�1J ��R�!Ș,��������>�O�4@M"n�- b�]��A�%�c��B�)� ����X�[!n�#d�q�	�5�'��OH��N�7k'*��@�_�&�x����y"�U�W��Y �j��Q�`��bJ�&��Ӑ��'�Z�)�ӶB����Tc�F�����*pW ��2ړ �.��A���Nո]Z�bQ�@���'��}nB�S&��y� ,�y�2o�_'�h2\�y�JA�1w��k����|%s�@�e¡�[+?����
\,Rja񄒫aġ�ğ*nD�@�A��~k�]�A��y"��[ȼ����l�\��va�8�(Of��dVTY��Ņ!)|࠳O�D!�My�R�Y���3m��0�Y!D�!�dӘ c@�S�[�(�$}	��� m����F{��������(q����ІF+�t1�%C�Ty��'׈�2pf��>N� �!*ϊ,�x��'L����G�l*��kȩ tf�3�'�DaJg���0!����"#�qДxR�7�� �3T�i�䢈�KO�lQ2����|�	���D��TmҼ�Ƣ�� �&)�Qa[4�!���T�YA����Z<Q4Aj�ay��ɾ=�&5�o]-2df����)�DC�wL�(�r�?Y�f����l�*ɉ'�*���aT%Rj
d��n~`-Jd�0�O��D�>�� �(޼a�˥r�<��D#�W�<��� ~Fl ���=�z��AS��?�
�'t$�R7DĘ8����$"�@�ȓ�|!⯘�n#"A�W{;O��0�y���'I0��1L�@
7��J\4�3&�'��r,ٳ%�X�W+\�i�L����A��yb(�$c�`�0@�v1�)k�#ٻ��>��ά<�q��S�Nj��D�9��=q��<�O�|F{J|�PҺv���sa��\Z��a�p�<іe�UF���N ;��q�r�\r�<)��h�UkNDr��拙d��,�'�tP�1A߳-��탴�"^?�ai�'����D}-��p����T�\1ܴ��X�d(�3�\([�*��N��j�`X"%����ȓU����wJ��2��G��o�����djܸ���
Y�J��W(��S~�ȓ_uP��Յ�.�߲^F��ȓ��}k�D4R8hTK�"Ֆ7& ���n����#%�ͩ�#��U=P���+��
�d��K�����8^[��ȓoP�Z�E��
���e��.��Ɏ]P�g\?�dh2Մ2�LK��J���	e���O���[$�W)`��h0%��Ya�8H�'�.�c���p��񷭒1L����'�u�B. �\%Y�@"s����'1��c0��Ng1`��Хk��t �'�l{��4o:��P�ϸ9��RH<��|8���!\=	@T�� ��m�l�ȓZ�(���K��=�Jp�q	J�P�H�IM<�$�ѵM#ܫF���@��6IWl�'S�?����zT�1IL�J��mZ�J2D����囅
VFq1��D���!q�<i���6i��(K7fԍ|���F��,>�B�I�o7<����.O<���	�N��B�>e�Z��\5)�L�����*V&���ċ�?�ѣ_�`��d�d�	0fJ�
BLIѦ��fV葐a�Ϋ����
�q���b��%�<�A�HG�$L!��"5<���"ظN�(}��H1HH!���X�F�@Ϝ.=���
��ӗE���r�H�C/�:p$�;��E�eHY��xX�����j�� �4{����׆�O�=E��� �H���D�ˊt[R�Ǜ.���u"O�:f-^"n�p��~� �մi�ў"~nZ���؃�P�#肰k�'{�fB� "g����K^5_U�2j��j��B�Ɇ�*�J��.<�y�p咽UH���2� mۤ�!��H������\ծB䉆 �0����؉*� H���P^�B�I�t��)�w�A�~�^��a�/c|B�I�lӔ����G�y�$�S�FFJ���7�	84�����bΖy�����m�B䉭m�X<e,�3
�A��D�M���'Jў�?�;S-�&x~��J#�X�5~`i���?O��IB�J��}�jB"j>�J�	�%ZO2 �ȓ6V���;2�:4�%	͝omN��?Y���~:��E�r� �{F`��	 ��y�`�m�<��Ӿ*b1��Y�(RT?�HO��}�8����	�%)$�I��I����ȓL�ݚw�	C��Pr�îI$�q�ȓDf�x0�l�(jP�R)Ln��ȓ,��\R��%a�>�I	��Նȓ�N�	���]A*�K��ehņȓ?���@R+S���'*�"�2���7�
��a�J}Dx�㜅duTi��Y���P�Eз;�aC$�PS�`Ԇ��$Ē���:���ׄ�`���?�bM"�m��*�v����>ͅȓ"�&����	G�@ J@�c�0��;P��D_�# ��0S㚟U�N9�ȓ��!Ɓ�;;�R�2�[���ȓd8\��"���.�b�2���%�ȓmð�#�D�G� �I��鞹��zξ�ځ�߳P�f���Ɛ3n���gpr��� �2-D���_0.�h�ȓ�`a7KK(���d2ʲH��rZ���.7'�U��'W�:�Ԅ�5����]>{�ܹ"�$� \�4��ȓp��lr!fQ�Nm�Egw�`��ȓ�d� B�Z �$Q�Q�%�, �ȓ[St
�(�* Jw�m��-��]��=����!��ԙ�Aږ~(�9��:^Ɯ��U�Mt-� �%sн�ȓqJ�(�d�
83Fr'Fٳ�A�ȓi�2أg8��R��/\�:t�ȓ6(�S��3�b�`n��
��ȓ1�)C�ŧS��!s�MG�,p���dL{S)�0�a��4�&��ȓ~�0A�-Spu25�Ţ�.n����yc4 �)Ű 伀@��� C��Ą�MΡ"!�^.Q/��s(��-���ȓx7����S��e"L
_h�ȓnw�x`0��+L�v�8�a�y!hф�	�Jp��jə(�8��YT��,�ȓP�hPy��F6�]P�O�������0����]j�f�kq��nl�ȓ'a$�էkG�EA0#ٚ��ه�51L(8T�!ƴ�G1��,����9��`̴J��Q�C+V>��̓�p��A3:&������G|��01�J`�P���`g$�k����y"mݮU^Y����6Ad��ǅ(�y�a�b�k���%��)���H��y/�3�*I��"i��,���y������H�CK8`$5x�����y�D�r��T�İa��IS��
�y��ˬLJ@���X:e��!pL�;�y
� �����^6�8��J�"AR��Q"O��x	 �衂�`?HCFE�t"O$����86��!�0\=&�x0"O<ȥ$�&<�DX�'�TAaqV"O@$��o�g}�@p��	�.6<�"OFE;�/���
�0���Y��Q��"Op�;�!V�8ИZ5�΋#�61"O�QeGֳ]���D|�n�""OY(�dӾ}-�p��\�wX��r�"OI�mI�Z�������Ip�("Oz\(���/�T�Z NP<��"OV�p����i`��D�8����$"Od�#�k\W NQp +�ip��c"O�Ա�	�@���!�A1i�H���'� r+�Ǧ3���<ɂ�P�_2x�T�\2��
be@x�<ـ�K�9 �.�?nӦ(RJty�@:Q��A��(��)�0lↁ�v�O����D�j`n1��"K��58�'M�5��h���3
�>�Nt�ߖ�Sp|��hY?"�����O���'��'K�P�3i�R�4���؃>�
��d�<�"�O3	�~y�g�\�&=���J6T� (��W�|���P��^1A���"8�&)���9c�0���Y3pQ� ��R#0�s&�xI�CG@��9�vݙ�LTuPS���jE�m*�"OnyYf�ʗV�DD�!�;*��>O�tIժD�(�A��8L�zQ�a��T�F�?�ke����y��Å[��e㐎;D�<[��I)h��y��Ls��Ғ��0P҈T�"��K䝉�G٩(È�?��3K>ym�!G��0X�:c"m�$�zc�ҍ��L	�N�#3ቨr��ș�J�8��%�7*F;^���r�-�,������f"=	��/\AX��f�H�g�Jq$@%m�<h���"=�w��R�@� ӵd �W�G~CH1#���3EΗ7h�5�P�Ģ,U�GyB�A9"����`��6iq�P��L nlZ���-�$��d>O�ʶ�T#+$��z��9J�dB4䍡lo^�?�Ȃ:�ṕB���]x��] �*�K���+�6L�w���"~��!h��U$}��FI�jm�Y���"x�La�aZ�Ed�\�V j�7�U�|�!YT&Hog���[���Uo����@�� b���I.{o�t�GM�R T �4��
a����e,�\���w!�:;`�e�b$�+r*�%	�~0�����/C�*�'Y�
���aS8>i�}�b��vt6ט�F_e��$B]6[���x`RAy�eQ=N �$��Ʌ�\pv�@-4�Є��#x0u�P�V�(V����,��?�� !,ӗsfͻ2���Z��<��/��"Y��W>.X���?���C�C��|���ZDBl 6�O+C�*(v�p?)20kxN)B��A�F��M3�(]�##4����v�<{�x���a�ǝ�fLR5CA++ψ<�F�]�ap��ǧR<��LH�h�څ�!�G�u'	U���0;ҠZ1�~�'X#9�a�CNfPk��N�Lt���e�ТE>��t�x�kE"C;�l���L�cE�����4�p����;g�j��M^�A.�)��@����[���M��{D�^3\� x���D� -7��h��F5_zh@P�:7�d�`$��`L�e Ƅ ���C�`OC �`�Xxt@@h�:6�L�����jd��� ޤy��Y!�Ҕ�^`A�sN�!�"<1��7(^)ăܚ�Jq�1J��K���
S�lt��-�-S��@ӄ�м��|���r%j�4F��K�aP�2�'��T���Mt��*��N��hK�q��O�PW�b�>-����>��D�95��,K7i@<@n5�5*V`ϊh�v#���`�e Ǹ^�d�!FI�n3�y#���!��*[x�1���l����� �x�DW3T�b��בݴYrA��/��2W�r�5O�QR��+�zU`�吩@Wl=�-��Q���ϖ6]���$��?8���3SWD!�p�M˶���{H.!�J��!ޡ�	P�'��0�s��D���c���Z��p����MsF�X�w�,9:�+Lw-30'%b���Q�̓�W�d�٤��w:]��*s��qHr��!&1vs�GFb�
����OV]��DȰ@Kl�2��F	��6Mӝfj&��C�Uu����%3=>�!fS~9�8yU��U��s��cc�����$՝e)�7��5��O�M �������-3���'$����]^n��C=(��qAb�i�/�	�����E��S�%T7"CKC�iRZ�mڐ�Mc���)mE�����W|��Z"�	p�����$I`��Aq�4:�Щʥ��"3�А'/��t���M(X�9�(�p�*Lrw+38�މ�%�Р0�܌J��C&q��	�M�(
� `���?hp�P:FO$u`b�:@`�.��v�M�f��m
�F(�h����8`QAc�9X��aT ��FW�1���5iؓ�M3� �g˜̂�֠r�:k(� yf�I��5�-�>RP����A��h!�)��⒞'ӈ�{�eZ`c�`�Ʀ]��Pw ʉNr�X;B�u����I?K�������"%�h���	=����t�^�>�)b�)�k4��ӱ�H=N���QC�!$�d��v3��Err!UX���Ɓ��էO�W~R�������^�)�6��J�l��>P]�IjBA�8mf	*�(�U�T��^:I�Q�C�עf��8X�
�l��y�[�,�9��2AR�ҷ��B�,�AZ�M�I.���J���R�5
�6�p"�@�J=&t�t+�< 6�M�p�Ϻ[��S�� ͚���v� 4�pc	&����L�Fo�E���n��!��/̂@h�F�S�tX�ƌ;~�Ȓ��O���lA'����H�6+��+�S�Gl`!bnX=?�`8��>�.�&�����3/��+1�S2Ei@�13��L� ��L�`�c��S*S��uY��ʰ�T�2.@:��%�K�^����,;�P@��V)1�
f�E�i�j�IrG�r�~�2q��+c�R���nF�!}Dp�LV�;�RƮDj�f�	�7�� �d����gP"AA����'��,��>���ǺbG�����԰��Td7���HE��U�P��ǈ�P������L�Rk0�H�ō�?���.����操P�@��q�	�T������l�B �v��C�qB���l�`����n���Q��۶�V�m��d�ߩA�er��Z�i�x��V��k���0𢅙;O��MR�#�ڍQ��]+R���Č�o�0�s2��!���p�b%�T�[s�J(�LQ0� ٗS>)z���7"�@�)�c�e�A%#tZ��SS"-�Rm@&@XV2	2w�	;2(�T�VJ1+�D�A���ecZ�rv�Gk�H�B�t�`P�e�#Z�����ŬZ�@�X�b8UnZ,�u _9I~��'�G,��{�FE [�Ӕ@�/��"I�ScL���8It���'��D*��c %#��M���5V\���2�IGy"��A�Tm����5%DA�ȶyPBi(T�u>Ic�!��0eJApǃN$F���Iާa"��F�Tq2�p�A�\��Ij^J�Ts�J�|,��P��H�*!{Qd	u?I�i߱l�Y�UFv8����p��Ӧ ��7�T�Qt�C;j��aI�	��o �ӏTCz��{�\%�!�P
\��a�CF��0�
Փ�g1���E�4=i.�R����zB�<���T���� uh'�Vq��X#&�X�&EI�U�4�X��ia�2�)��h^�)ƐC��L�l��O��p�R(BQ����lV�{V��e�Z�K�4E ��K8�Q�����V9@��ł[�H�2U��J:����T �}��y�/�VyF��AY,Lsa'��P��Iŧ����ڴ!��{��A�/
PtX���X�H�|u���$� ���!a�¥�O���P��"@=۶.�R������	�
Lb���0i��a0e�,3N6,���7��4�d@����C+}��qC�ȑOH0�L��5C, ��2�� ��I$[�)zW"Æ��FB�a�t�U!�#up�p��Ywo <+�f�$Y�	:�A�
$ʔ�`ϟ"��&�m�4)vJ�0)I��릅�o�Th��	 e��<�2��m_.�EzR)�6l"��q��GVf����T�}�"��c��*�Ra��W�(bJ�7�B�9$
�*�zYSj�>�u�'��P$ �J�N�aT�xa�Q�$�@�swI�>'U�lDzR�1)qJ���ҐU�୓TH�,y(X��jV�D�ႂ:f�SF�'�d����ڭ/��S�1ev]����;M��2h��j�1���&�v٘e��.��i�O�����$�>� G�mp̸�-Q%�d�
�J�	��G _��(2���u�B�����*���Rv�R�[��P���ũ-|���k_)e2��J�7tT��b'�
)����S?_��	�@<�����&X�1`�T�PX�ćO�JI1���L}hP@C4�4�T�%P�)
p+U �@l��^�L%��C�>:�z`��NR$j�,����U�04���5i�6e�V�K�'-n!K�I&"X�D�`Ӱ�@��/s��1���6\L�!F-�u�f�R�@H�#*d�-��i���\ '{�����C*Nو�BW�.WQ��8D` �^.>�F|���I7ʖ�-TH<j��[�B=��[X������3	XU��y����5K�N"&e ��$(��X��i*Q)B��>m��=BЪݐ��̖X�|	�kV�8�n%ٰ���8r`V�!{��
"!·�,���˝�%b7=XL8L��[}\Ź������4Sw*8F���g@��]Y�6-\f�Lu;G�Y���3�˜8αA�w��8 r<���]:�L�K�LE��S�G���đ�a�U9c��T9d
9#u,��`��;�B�#V퍕B��+RGM�f����c���țk<Qa����Z1�DR����+�B�G"�Û	����bZN�$� �_�G�$yـ.,�U���g���R��ۅL���9NP*�C�‰<���0""��n�4��5K� �����a��Փ�
�R�l�6]Q��LØNa��{P�=?��E��%�$|�8���F�?����'Qi�7�BJi��S �ڼ=��]�qeP�?�DQ��L�A}t9%ˈ�?mh��<)kH�;g~��3��r�@Yt'FU���C�W=�H�bh�k�� ,ю!�,���lȑ+�^P���"��X�m�Xǒ0�R�o�$ʈ"��0��A�e�üb�(��?$z��Xc)޶Y"�{F��{}��ǝ�3��I�E��=a���GP="z��(�N�*B�x��">C:Jx�&Ɲ*�j�bD�V�}.��#�'����ģ����i��,[Cb�b�۝J>X���I�p����d��!����4cĝ���)W��/]Ht�q�
�zNpYg��I9f��[�q��I�EDB�Y j@}Q�	`ae�:�L�*_�1,,$��.b�
5�+}#J��T �<��� ����VȚ������I:�KIގq���!�:/�,7�2,�H�[��QE�g�н��HB���I��@�"v�I!�
\�i�&��H�+
�:��AZ�[j����+��PL�?J���5�H��J���+�0����D��@��h���Ґ%��8�؅���!��ϔ�4!���	p�u �i�C��`�YwAx� V�]d`JfGQ v���eo�)��tH�	+�vH+���Q��4���� ��3�K�o�2�	?W-�iK�I3!�� ���"�b�c��Y��� CR�Nn�-J1I�T*��rS��idfƶr�����|<J��$�7�ȃ�jG�/F*�H�f��'�,�Q@N� � ���	Ba�h©���$� �!�x�:�Df�4$� �qp��!��'��B�իa;��r ⁪w������$�v	U,L)R�fpCE@�Q�!!ւT���C�J�#� �f����Tyaf�.;6�� B�	�j��͐�Dc��F~�^ 6�
�X�c�jc'�^�(��Q12@�)]�sv��2p��ɂ�"<�"A�a�nKG��-��iQ�f
%��EB�` t��l�#*e�xr	�O�b�Ⱦ�0=ч$�
j�q�`�e��)3�*K�{C����ិ�b|9&��1T��@��$ˈo+�D3��6o��RW��["?��ɲ�:"2)�榟�G�T)Q��'l�iH�O�w����M5)�A�-ݑA<^�q��8��43��0�1��vz�AGf�¸����"'Ș�q�va��$�8#li�D'[���z�'$\���(�ɴt:T�b�ȍH�0��U��
4�Ls�	�+#s�(p��H�N�	����b�&�*2g�Y�ݘ$ITR)�")ҩ v�$h�%��K�@��'�~԰g�Vdep9֥:M(�녏x>|��f!eW��ca��>[�h�觃WY?�2�]	$�Պw���V�D�4kŗ/e^�$�}ƺP�ʁ�J�Pl�"�,E�0��'��@��Y��֎[&B��t��dj�1)��]� �p���bՈM��ɣy��0��k���LDJ�䘱2ʀ �M h�� gH� ڨ=��c���Ty�Jrs���$���|� ty��0b�u�[�oZ� �35��{Xz��
�6&��51BA�3Wߦ�Ї��H��a{�ې'�![��~Pj$�t �y�HP$��6I��ڤ���OP̙B끬4�n� (�<k�x�ad�D�-��z�� �E뵤݉y�T�� h۸7�`��S`ٷYF؝����	���;3G�= �q��\�|�F���Ț;1�t���'Dn���_�]T��pa��;^�DZW���j7�m�!T��h�C�&pHx��6�^W̓sIp��vG.N�h��2�T�*:����Ufy���(+[�R�:TQI�Gݯ̈Obx�D�E�_��APDdI.g� ����IL��I���y"�ɓ	�tP�� � [��A �D,a� ���ǄHpU
 ���Jv� ,ΣG@�z��$��B�D'O1`bց[�49��ǉN��؞�m����@�8~�$ɤ�ʏ y�4Ȧ�)H�����	�O
�� �O���T@�:zr���DE��f��ȍf��kρ��(O������h�0se��Sd/AkIZ����̵$.���q,�M���2���a	�l3"�����L���6���85�-�3韼T�f���`�f�[}��9Nǰ��XS㊗9�M����>B��Swv��Y�k�2xٲ�k�s<���G[R���g�i
pU`�`�M@�*_&{x�LE��5��d��?��A�7��T|Ex� .�I���ia.���:c��:3��̈$����!�ɋ�1 ��c�)��M��Q�ٝ���*C���0��ܨ�L_�q�Q�/����� �<9)�HsW!�z�L���'(�@cw�;qp(i���[�� �A/� 6����G"�f$�U����R,"ȑ8:w~4Yr�0Y��<�q�ţ3���3G�5��!fL]$IEnUIt�GF����"B:�(`",�so�P��İ ܸ��b���G���J���L�@#�͛-+����jʭN�|٤+D1۶��"�NF���Z�4�B����3N�3g��/=�F4�go/g���Y�C��a�<�nL,]��@��^�02xx�tM�w�*�3�d�)C��4@�F Nߨ�i��'OЌ�*΁1a2)�̟�O��s�ʆ�V�,h2�lH����y��_�U�|p1elåv�q(_6,��c��iO���
튍]N��ҤU�f�N��tAơYۺ� P��,OX��d%d"��t���g�&����ÔZ�d�Ab&B>N�h)��yV.T����oS�R���@�^��~Zc�H���U�Cg�рdCُ[�n��
��v���k�{��Z`f��3r�I����v�.�S9��@Ȍr�*��c�$�T�Y����"}2���:�k��Rj��DMH�'KҔ v���>	�[���M�'��SmJ��� � �&!e�� �qy��\���)G���{�唩PQ��@`�:@���FY�6^L�U��'�C���~���K麻	M���"��bS�d1��	Z��HKp  �O��Q���""F��0��ܥ%EpPAuQ�!�'Ɛ�$9	��JjyB�H�A�'�X!b\W���A�G/zx)��#�Oxp9�C�!�՛���~�(DB�*�9@�^$À��=�x��Z�u�my�lMe�|���A��O��ZpG���.˅S*��5�u�)g�x�Ѷ"OYja�@�"�n1��ǌD�2�b"O^�h���8^`œ$�68���"O$b�� f����L�;J���"O,�90n�=_��X��	2C�H�"O����	�\����^ p�
�"Of�za��c� 	�d��(|2�YE"O�dU���R��H���2gi���U"O܀8��i
D��O>:F"��"O���âX�0��*�!_����s"OL��� FI��!
�d���"O����y� E2��Ҝ$Nn�� "O������mj~P��5%���E"Oڈ �&	2 ��⡒�G���S"Or|�P����亷@N	�M�!"O\�H��\!����˶D�n<�v"O��H�!L�c��Ux�J,�!��"OBw�D�6İXcm�;:N�!3S"OE'�2X�xE��=i!����"O��P��:�	R�L�<��f"O�ū���]:��Q,�1c���"O��ui��%bqf�-9��8"O���V��B�\Ȣ�&�K�>Uʣ"O���H8�AX���1r�
U�"Ox�j�nN<.��C�i�!c�E�"O��&H�"������
��0g"O:��� ���Zu���J�hQ"O�H`v�� PH��P

�^-�c"Opy{�L�+�Vt+n�%�T]�"O`���� 1v��l�o١s`�Z�"Oʌ��@��%�P�e/��rGVU��"O ]�7��,V5p�I�8,DP3q"OV�8V*�3u��TC�&��c��,ȡ"O�H����CL�-�u�ۿy���B�"O� �����J/�A�
�|,ݢ�"Oꠈ�*#fB�A�jL#oF9�"O��b��̏*;�)Ӥ1YTqB�"Ob��t!V9�PY3	O���"O8\���+d<b�B`���4"O�m9�ۍ]T��uc�""�|��C"OX��ԪV�2tT�S�U=u�h���"O@����ґ�7#L��v�H�D^�<�q!�+0)R!T7��a���^�<W���x�qG�W�\�>U�K�Y�<�`�ύ*��u�1��5/�l�T��c�<YB�_z��	�7#ۍ>y�]c�(�\�<	��$aR������1�s��NG�<�1�ۭ#1�PK��D�X��P���C�<��K�昼3�Lx�x���"�[�<��B�
t?�	�@��T�v�L�<IVl�&\ Q3v�	T>�����L�<�F9�ҹ�6�ɢ]E��I�b8�C�fZ�'�r-@����8O�!�T#L$���H��P#mp9�"O �s]3,�pE��]:)P�Y�`���@q(x� ���R��S�Z�d�i�+O-UǨ��`O��94C�(�����A�3 f�����&���2�ܞ/��!"�^)�x�0)0�)$��>`�"١E&P�J�v1ƣ�%q���dɜ:��a��E@%y6i�������'��;\
|h�x�N1PmL�0=	UB0b;JH��%U���� �B�''�ƣ��o) |R�Eۻ218"��
�q4�L*0t�5ZԄ\S}�u�ȓE�y@��1�2E��F=d,ϓd�	���L�r���fA�@�Yx�,P���OZ��FU� �JE��I�W\���'*T�� �qn$�[���}� Q��×T�Pw��9'�y�� �����M$qL�O ���טN�h5`Tϒ�W����>a��%@��#> Ä/L4|�R"�C���� .A��B cs��.(45Q���	�| ��2�HO���e旗��4�I�O�h2e��508{b��#�HO�"�B%
]*�� �	QA��/2K�2��Kv�p('���Є��1ʓq���b!��Ir�x ��$� ��z�E۝H��*e(F��y���-tR��ᄋ�(T�x��Äɓ��b��I�"cR��(3<l�YP&*�d��9����-��Zd����OZ|A3'�����@�I*j�*�Zt!1x�e��(*��ԷU�`��K9àh ��U!E@yK�IV �y,Ӣx�(�� L��&ԥcf� ��~b)�ce|1 .�2 &]ExA�%)�"	��.Z�d�B�) b�> �]� ҇,�i16��)��[2�$a u�bnۗa�V�y�"�<$�]:� ��5fe�W��Y�ω#prYUӽE
�aXui�P�'�(�!��K��p�������R+�,�w"F�r4�q"K!�|͹2�A�y!n�CM�U%� :�(�/������u7D�O8�%7�3T	D�1}�3P����DR��O���s�]�'�8((4gS���D�Z>��hB+@u21�ش@�V�5f'�f���d�|�<����,Sf�X:a���C�����ꦹ�5*�޺[c��$Ў�c�Q�֑7*���p�cΣ�05ڔ% y�Xe��	�u;�<q�x�%R�~�Q�T�E��$J��֨mP�)!��.,G�e�� с@��t���ij��$�)hT��(Ӫ#=�v�Ɉ0&�u����= QD� ���?����܆Nn�k�e��f�i�c+K�e(�E�dA�� VD��ƚ�<���(�Lz�D��C�V�nѧ�O11���%'�I:ў� �GU>XB���L=m�F�I({�Vt�W�;��9J%�J�J�D��G��x�f����ܠP��$�$,�*}�Tt�7K�:��*���N�N��w/�|Kh9�&�l�� ә*p
�'���p�'1Q�
�_�hB��NL &���Q+zF~�U�*#�b��AW,l_�쀰�8U�\�jb�׾-p�&��^��C%nŪ"�hŋ��.iV����O�	���]-y��	��ո1��i�En^ ;�݂W9O\�;�O�_��)�Ac����1ċ�92��E�Ŏ_�1ȸ�`l��*�I���+j��u��͊	���	�hB�0�*��.h�ؠ�P�	�c^RP�g�@�*1�#�0Y�x�e�Hx�('A}�a(vK"̨��υ'�YRT'\`��Vd����i���Yo0܉�kY������eܺ�F�]�'��d�C+3;<\9)F�18˛v��7�3�+�*[*���vC̤Z�R ��@?g�(���"�=k<�P�En0�[F+�*Z&���I%�5� ��k�H��򮄥����H��N�'���32���'<v��-�?Y�S�G�����*O�r��eFA2 ���N[
�L��Ҫ:RbPy�����y�p�'��#5��6
���P���\����aݍ�^�����՗	0R�0�GT-�HěF יJGPi� U�S~L��b��nj��t��
6^�xeǕ�(�DثV �F1ꕱ)B�1<�;��v���c���Z���� >�1g�Z�B7������z`~A�V�J�>KVT���M��Z�`�V6h��X�c���M���F���m�Lx��Ȱ�W}>�І9���ؓC!aJtF�I�hq��9�
	Q�⑤@�jX��}IP9�6���d�	�$ t$��GRƌ�c��!|���̘>W
���͋:�9HB���o�k e �KR�qc's�ͣ�l>Q��wЭ b��m;���vh��}4 8�Or;��Q01 �\8�肸�J``H?�����u(N��C�9kZ�'���f����d��>�������{�ziCF��K�����m@5���ֵb����D�h>���͘$hZ��q7�S�U̪	�7oS�.֖e�&�؛v�<B�L�2{�,ם�c��a�&�"J�J�f�<O�t� �\�֎�-!\��c4J5�n|Y1�K�j�N�ҥ[�G�J@�L��T���ϸ'V,\SW Хg�����ُ]�x�2���9u"fn̼hՂ��e�)F���c@P�a��ثfM�_�|�"� [;
 ��~���E� -S^�Ԡ7h͎3��4�gk�;Uc�"�}�ՙ�X]���_�02�(:�Dޭ!A�0ER����Js�.��*�D@�Y6�Gj�7�4Q�R*��WE�:@E�z������-��b�w}�8��Z�8�����M�<�L�h5��*0�09$�N ��T�~�C��o��`�ֵ�hN]�M;���DϦo��P��=f����	�6J�h�V�lW��#��]�H1��(ӄ��mԛv��"�v�[��X�Q��H�h���9T����]�|��'"�p�s]x����\�`�L�'����</:\�be�F6O̬���i�S]������(S|~@�D��k�
�)��	!8�\�y$D˧�`�h�F��vⷬ�EG�h�`�ֈe�d��@���}�V�i�dJ%�~�8FI.�f0�,@NƼcp�[�HHE劉���6k�Aj9���$�	-&���0�*�$p��M��t	�P�g���B�ы\�u_"iRCVxb�$A�m��U1'�&2I~y��fO�V�)�K\wZ0I��{g�@�P�ÑoF�m�NO7yz�2��<���ӻ?��A��k�^,P�P�[iX<���=���UB�
��a��c��=��lx��<h�A�%��;l�S��F:P�sF��_��I�1��?��p84AC�:e�m�0�����M��0}����,C#�̞��H[�6d��P��00���`��6�&]�!W>�{#�\_��P�ݎ*��\r�N��#��Ue��&/��h*!NT7!�Ƣ<��Y]ưp!��<J�֐h��Zu�R�y3-�x��D�2��� ���6��)&^bV�!��9e���f���8�[��=6�e����n��6� >t�Q��[Gˋ*9<�UJ7���h��F�<p�(�qP��%{��e��12��� �aJ�2\��[p�R�.���\'}���N3?�9rU���\ʔ��L���UFT�N �Ojl����,7�x ��X$y
Q��$_�J�cjƃD$������$f�p!�¹%7����־S@�:F��q�&�S2ک6Ex�S�a�k�\qwC; :��n�}~R�F8���"�ä�[���ay|�ˑh�$k(h�*�3^�Pqafƹ���Q�F�&��v3��xrÀ�*���i��F�2$CG��!=0kq���N���!���uE���3�eeQ�هK�Z�ʃh7y�\�p��
H�A��K�:�lx��G�$�:��O�Z�t�<[�.�<�0	�"/�]x#jƵrq����3Q��t1��K�>�A�c��=Rr��$,�*Oa�$QU�1�|�G���Y��0� h�.P4y�+��v[�0������b�ZU�4�n�w�N�\��ʰh�� aI+j� 5����{v@�D됅D��=� ��0C�$_�8Tr'U�T�P�+�
3.q�Eh�&xLeՉ�;Y]:p�!�l
�`g�k���E��:�����N�~2c1�[9]Z0d��Xi �0S���h���*I��#�d��|ܪv���lf���O>W@Z9ЎG/n�z}��Ɓ�O��s5�D��f̊6,�Ԧ1�
�a���PeQ"�,�$�*I�@pXF��_ �x2H��mMT�F{�
R��}8w�	�����r#I�_� m�	݅v}�D���-0���U�S�'��]`���$��"I��T*�a� �f�Hթ�2�k�T�y���0� �#���$ Cq��:�o�V%طC0��(:0��8Dt��6Ɠ�v�4ӰJ�!n�m���Ɵoe<a�AG�~b�N'3�X{S�?c�yp���#N��Y��ȓ2m1������m��	'g�rdY�o�,�jY!t��zY6mg���5�ۭ*�,�EE EԡvƓ
Ak�k���T1��Ї�M3�iE!5�"S��,-9��@�40�^Bs�>����/��-��(w��$��JΠHN���n���8�L!j��4�qdU�+������t���F�ϠEP�BVF]�$m�T��������V{c��0_�D1�,�~Q!"���9<����K�&[ �J��*A�2EC�!ڛ;�N]�]@=�C�F�6M{��Z�:�JQ�UB�|���D�of�l	�ؾAI2:���om����˄V8� ��T����V�C�VTQbb����1��51�Z�!�H����1B���� �d8�YQ�N���5����!FC�)�`��'[�o8�AT�@��Uؒ��'�F���Azr��q1撲DP	Ya�^���G�=zY(�5O�<��mOVC`��D��%~�1�4k�"��PHE��N>|M�g�I��O����՜�Ԡ�����B�+4K�t��m�>D����Yo"�Rs$N�ט�3�������VB�3E�u0d��x��S�	$x'޽a�G�G^��˗Hݱ�a|��P3Z��!��-{��qӠ�Ӕ\����dsN��'Y��>E�U	��]���A6'�/~��Y�`�Y�
%���Fk����Ɉtfv��3GEL؞I�y�����H$��`��iͥCD���k�
c��s���n��D�p$�x�2�&@<ئt�V	�&NR����
b��[�ʷk��5�3,��!c�O���a�`�$Ϗz�U�%��=��I�E��y�����/�X��������%~�,�C�ɞ3�M��GE�\^t`�'�<���ZvZ@�Ł�'y�"=5�O-w��҂�@LF��A��)P���2P/+s@���;^L�R�l,u�ם�E-Y��R�P=���7"x�0ۣ��bЌ)� �4#�\P҇�3=Ka~�d3b
W�a�1�d��$D��y�ƀ!q>n\y6���WCK�d�6m4jw�e� au�\9��;s�1�|E���ʪOq�Q
�!�+�0>�,��	F]@&C�X"8C�iǎ �rr�m�7#Z�=@�ð�l�P`V"c��d;��^� P2���zb�-n��U���c��"\B:�0/
R����:�B?�A�Q��:C��\jb!�� ���5|��3OA7�E�r�-��$0�%:1��`à�.o�=��L� FS|��I�Enݢ�i�f�Ñ�;x��AB�!֯~� 1��K�?r���gJ�%GdɊ��S��n�ӡGM�|��i:t��=%b� `"��/qn��Ʀ�1(��B����?��F�lm���]�P�K��&S�hz�-Mh�	8q��<kpQBUa�%P�.0�&������@�[�TY��Ե(�y��E�rp��PG�Z�]=�hhflʬ��9�'Ġ�:A@�wy��)U�>�;�E�u����w'�5D�h�vV�$��=�T��pʟ(C�����[�^����
������q�����v�n�#�e��t��l*�z�/�;���稒.����n�7g(�qM���L�:� Đ_tΜ"�&@�լ��1�T�qN�u���2n4�1-Z��@���$?�"�.�*X�@A3(���J*��,1`����C���r�-!�6T��#�,�2�	M�~11e�
�`���[��xy�z@
�:����`������� ����� 4�KG$�,�ɗ��0�L9�!#R<!�f, �l�~R����)D��g��v���J�Ԩ)BԒ�O���]r��U�1��|���A,(��y��2��L�@@/-���bekG�FJ����	),1,�Q`hϯT�r0R��<r>�������ReKǣDM��kgcȪ*>6��hέP����B�٩�'T�@FI��D�k�68)7�I�'��MۃO�*6����C�qSV�&�0&z��H�.8�u�嫄Xl �"�!�N���%Z�L$��C2,h�Ar蕭>�U��'���*
�l��CK�=x[�����Z�����W?9����EY;O���Jm̓L��5!����V/��4C2B$��84� ��k���#ÄR#A��<��!�;��O�$� �A+z q�DL�K}pM��%I�
�haD���y�G�y[���hA�E%` ad�MrrM���	������h��y�0#\�\޶Y��g���M��?O����-
5;�����&��qC�§�h�͙XO�MI�.6�"p�1��Lۊ�ᵄ��'��y�O�X��͘]C�q!��&���k�f��d�ߏ�(O����K�jbp*�/.>�y4KS�|8d�BfɍOԢL1e��<�:���G/M^��Є�˗Q�T�c�x���,���g���,��i���)O�b.������4�6���Mcs��7М K��ܧa׬e��哟2�L,#��0�ER�-P"�m�; t�2G�1c�F� �=2J����*p�+�
6�W�N��<\���*ғd/�]C��C��X�l�=V��Q�B��W'��qD�كw���3��`'�E{�Ξ@��H�LνU��qv��G��Ԓ� A%^�b*A7z�<y�i�/�d	t�'�>q�Iͯ)֦��䝻5�t�{�׭s&p��-{!a�Ό��N�����٢@�V��p����.��Y�؉ �M
�h04���'�,���˵M�v�|I��'�j��eKb��A���Т
ԝp�a����CAH8R�9�P��F�����8`���#ځH��ߊ	���[&�|�c�3��ы��;и�pvB��O�M`�(G8a��÷��t�e�Lu�f�c��S��)�B��_��0�����e�����`M3
���Pq!;�?2�K�-�x	㡠��D'"�R��!ఘ�"�ֳ�����D�l@�hܧ7.!Wգ �<$�iν]a��!�a��_AjZ��B������}�����yOq񡨋;|<]�*� �*y�g$��]���@D���	رL��yN}�qh
9�~Zcٔ���/��MR}ȒnM�1\�8��tib�����i�Vy���@�H�
P�B��ev)3c�:{��$��.�P i�07����H���0�{ܘ\�pf�4(.����<��pt��۔L�P�)�'Lt�a��;l�,����81�u�TW�����V�`���$?��fk��P���dn�M2���
��`��H"U�Z�O��`�����}�%��hb���r���B4�>-���J�7��� ��OS<a����)4:8�m׸d�x�'.J���a�j��)��S�� �B�1�'3���ꅑ
e@����kQN�
	�kSJ��\�@�u`դ�2R�Y�,ĉDT�� �9$�4�b�NWr�a�Ƃ�j��Rv$%�-'��d7�'}n��"���&2F,@W�KNB8�ȓ�H)���p�q+Q�������H���4��^h\�b�\�6�X��!��|P��%I|��@���{�Ҁ�ȓ̆%����K�4]�"A��n�]�ȓ ��4C�/;w�&��uΎ�U|tL�ȓ]1܀��ܐ2p ��ˀ!�Fq��g����✣/o+�Iaѓ`c2D������!��1��![���r��0D��)�ŉkܺQ0�O�!~+��3'B/D��RMj�J�V"�)}���[��6D�@���	M�֌KAL��N�p�Y#2D��sb�T�p�;�P�WdI��C2D�k&!P9SF<�S@�&Lxx71D����c�=#��Xk�nA4T�B�	�}�����Ǘ�r��(�D[�kb�B�I���!�/m�,P��K�h�B�	�u�ЈE�܎  FAA� ӄB�	�# �P�3F��;-<`֕%��C�I:=�Yڵ�^�!+�5B�����C�	l�<C�y��0�THWIQ�y�	
�3��뗋иx�V���Jդ�y2䇳f)�i�vaª`lX�8���yr@&R5�C�B< }�5 �	՜�yr�˞}Sz4K֥ڛ|����Qb�!�y��@"X`��)��h������	��yr�#!'�(3��N�k�N�;��H(�y�ˌ
+$̈�T�Ew7�1T��y����h����kͦY�6(c2@/�y��/Y���*D�)V��� ���y
� j��G �?o��:�D�(�Z�2�3O�\��-$�^X�O�d2t����g5b��Dki���@هvJ��sFF�J�t5xI>���t��V2��ͧPp�]�G.K;X�� �g�nl����{尀��%\�by�t+��X>U���K�a��L�.F�T�mqR* ���D����@�g�$�,Z�(˅f�H�� 싌�	�4���?E��6B��1�f��x�00�JK��M�VHS����ȟڵHB��)���qg_�E~H� �K�'���Ʉ�I� ��	m���Ŏ�;��O&h����O��;��w+<]�.\�q��c6Jěm�bD%�hs�L�7�qO��<d�A��k�N1I��E=k�m�^�X�d�	n.qO�>�礑b8A�6܅L�l#P�tӞ0Z���S)!����Q	`�(uAY�r"�m9��ЋK>�b��9���O��M������ �.T�(������:�@I>�зit*��yJ|*�����JJR+K�oK���G��f.`�)O�)�w�_��1{�"���N~24$�.&:(��&[h�z�Q�N���?i�c`��`�OQ?	�+g��H���؟z5�z�C�/l\5x޴	U�'��u��S�Ha��s*����I �ƿ|����ۈ���*Q���0I �OP�$�!���9�yK�HK"�u�l��S�$h4����2]bJ�`�.h��˓;�v����㞐*  !���ó{f���'JR>E�P'��$��R�*M�{*���'t�Ё�N��D��fW	cāK��x�6��1d�S�I�.��N< �ĹT�W����9SY�a
�l�@�|�Ѯ�<���~nZ@2��-��e�Є����9CׄߜrI�C��&
L��߳tL��!�䐾T�a��JU�
�Ydh��%\\��Ү�	�?Q���E�(R�兎-츙�çw�B쉀I��ERH�HV�ژ6;�ys7��a2ߗ^�z��m��Hc`<��Ȑ!�y�a��sF�@�-�"D0�	L��y�C�c.>)����nT�Ԋ���<�y�iU��q���o��*U/�7�yRXe9�E��g�m�(��`G��yb� YH���12}��NЗ�y�P��xA�T�g��a�y2ƙ9+(����1f�$)%��yrNԛjg�⣭�95�"��"�y��L�$�p�F�A!4�4��ZQ�pB�	�qM�p)��8K�T	Q�+\3gB�I��n0C�L�C$L�#��,�C�	�~�@)�怑�e6�Zt�R�2�B�	6Hsjt���X�u7���p@P�f��B�ə}ް\�ԫ�,1O�)J�
D��B䉉=�!z�!-l�m bʌMhC�	*K0b\�Ə -��"��
� VC�I��!b��9�`�*�	��>C�T]r8IA �yt��k�5�C��>����.)+',�*�	�5V��C�I�o�8�q�ǔsL6q ԉ�<y��C�I�s�^` �AO,E:F肨	s�C�	�ne^��(���ɢÂA (ʮC䉱1�b��T��9��T��S�_�vC�	�c�z`�� E2�@1�)�d��C���PPe�0��<c��͐#a�C�I�qX�H�/ ����"eصRC�	�4?z�e,�I	������pw*C�I�><�H��'���9&�F�, C�ɪ_X5��
ˤt�����IO�lM�B��8�#�D:b]�y��P5�B�I�^}.I�7m�a���8��N�h�C�I�w����ܝ�b�N�zT�C�I�qf°��[7ߦm�)M><�C�I�BG���h��`�n�h	�j�C�I>b/@d"w�^;� 5����(�ZB�	�5�6�ӳ��\ΪЁ��ǋCK�C�I�+_<x8��V�!18�HC�I+)����ħϻP�4�-M"c0C�)� x�j�.�x�0�_<Y�\0�"O<�a+^�rE��(���|�0l��"O&��1��&y.< �B���a"OJ��g����G�G|(`"O���&d9��������ʖ"O�i`w��(6bH��!�ߥV�dA�""O��坭q�
�JSf�N&�yb�ƃG����j��BԬP�taB>�y"�ga�-R�z<pc"	)Wm�9
�'�6$[�'R��.8��m�#= �
�'TeYt T�V���FW�)��i�'b6MX$��M���G�wbi�'�:�����g�xJ�,P��
�'�>�E�����j�Xd\�
�'WV��p	��r�6L9�W	��Dz�'{���	F>���,����p��'��l�
v�� �W� �Y�0���'`�T���l˴�X�L�W	����'�2���>���	q�F!W�j1��'�P9�@�>�p��C�)SG�u�
�'�H��s(ȱ�Ɂr��2 :���
�'�蠉ET�r�Dۄ�į�JI�	�'�N�C�NF1m����ť�
4�D�1
�'ېY�E�Z2�%p5.�%,dPs�'ڨ5���a�&��J߀) ��
�'ľɐ��O
zF��d�L�<�I
�'@d���f�5�\�R#�֬܌�X	�'��USO�=��1��U��i!�'���)���B���s����J�'��]�Eg�:!���iDA	(I`%B�'@��qGK0����@R�5��
�'cP��Q�&�c��\�|p<�CO�<y���3.����	�F[�����N�<�"��.ri�O_�H�sk�H�<Y���h�a"K{"�;�b]�<yA�W��&`��ܔ\�p�{��a�<q�Zf`HhѶ!�����6�\�<i�>vQ��yS�� e��)C�A�<Y,R23� ���]R�$h".h�<acH;#�$����:X���1�d�<��̜�9V�.QѰ�2�*Ĳ(�B��-Ζ��4���WbNE���(cXC�	4Y/���D�P&| �Ec�b�(�2C�	����5B[���jD�M��C�	<��L!R�'|����͋*a{C�I�����t'O��$Jz�B�	u�} re,|-��u�ȌX�B�I� ��U��EF*g�( qkǒB�	;"i�R�đ"+��T�X?4C�I�Yysϝ�5�����bT�9�C�|����QC��E�n�6���B�	�O]N���#���ʃ�˹i�C�ɝ\�ԡ�@ZZ�N�iv/Ƚo�C�#e�fy
���>�L\Z5�.QΎC�	�UG����V�@,�uO��?��C�*����'obԓg��W�rC�	8k��0���`Ll:�%��zC�2�rš�dن.J��W�!B�I�S�:, �L�Z%&Ia!�9��C�{-8$B���7fi�5�0��C�Z��%�7��&vRq� �=O��C�I�~2�:�՗Tz�C �"��C�	�)�Vh#����Oqd����ӴC��8�&�%%ڃ_��e6�P�Lh�C�)� p ��C�Fڴ��U�Ī{mz 
�"ON�JVn	2f�M���+~N����"OH@XD
�#R�BMH@�P(;g��c"O0Q13M�Φ<З�R_�:�B"O�Ma��[��VcY�=�ԛb"O �pacF:;>0p��OB����hE"O茱 J�ttr��V/�X�}��"OvL��c9P&=�n�SAfD�R"O���1��[�h*�F�n�"�� "O"�`�.�4��a�	^���H�"O$��E�I>, ��⎥~����"Ov��eI��8y�
�2p8Q�"OX��G�ƥzr��blii0"O4��N\86I)r�
�5]�$"O��8U`��>���Y,rV:C"O���S�}j�B��X���9#a"O�ș�չ3��|Xѭ�h�����"O�D�4e�1��Ta$b��
�0x��"O2ku��J�L�a���UcReq0"O�(�Q��Ō���.V�,��Ԙ�"Ob�����YB(�&��./	�`�g"O���٦dC���ɢ/�4e��"O> � /o�p�QfS,1��X��"O���@Y���3 eΧ�~�i#"OZٱFe	�n� �;2��z̴h2"O Q2I���<3(�
R�\H��"OAr�S�O����c(���q��"O�a@ɜ0"�d��F
���"O�I��E*+Gt��6e�l̄��"O��:�Ǉ F�l`�!�8C(��"O���e��,��������£"O����iRp���ԪaJ��"O~����#r�(rD��3-�P�"O �� �@+w�D�#ϐ��Eza"O��j�$Ɠ����U��!.	�i�'"Oz��aӕI�I�0#Y^�T��"O�-�C��J�4����	�X���"OT�85��>x���q���FB1[$"O���B%S�X�ŏ̴P;� u"O`���8:zp���OÖr)���c"O�$s
͸/� @� F�n�9B"O�"SO�+f@�İGE%u��a{�"O@���4NU88P�"�+��`��"O,��3p��h�!�p~��c�"O�� '�u��)�ª�/b����"O��+p��6��Ȓ%7Jj4�"O �j#"ݧ$�J��X�Yڠ��"O�=P�G�ڸ�&��&uk���"Ot�!ŋ.I5:�0a�Ak,I!�"O����l(|7���E�e.�dCA"O��s���.�T��P�O�q�B�#V"O� ����=~��2���dM
��"O��P�XH��b��a*`;�"O��)i��LI���,K�E�5"OH�Pe�
����M{~�;�"O�,j��'B�(4���. rqQ�"O���%�,&qr���U88��yA"O�t��}���6 AF-^��"OJ�s�A�2)�9v�X},F��'�bGQFt��c��=<+�'I�$XEB̥%���L�qݤ���'M�tɌ�0������fi���'@�B�/L�/v�z�. t`���'��Az s
��A��
�pt�
��� T���S)r��`@�W���p"OR�h�k��J,r��a-�r��}s"O�e��	��k'�� ���x�"O8TAp)���"&G�"��5h%"OVMje�k��E�G�j��C"O+�۸|��D�Rm��d܌{=!��M{f�Ir�G	�&Hh����7!�D�!J���#��q�lp%��!�$�g�b�q"��b(hyA�k�R�!�$�b��YD.��"d���O�U�!�DخpC��yW+����I�j��P1!�䐧#z�P3$�-0A�.�i"!��Vn؊��
_����� !�1�
�)�Ũ 
�BmN�I	!�Dǃf9��0y�|�F�֞_L!�d���L@"���`�(yCj�;!�@�tC�ᡑ%M�"�l��2'�%�!��#�6!�ć�l8��F��!��ο5��y
�虻\���9rf���Pyb-U \�St+�S|� [��y�E2yJ\%���E,���	�y��(���0��h��k�NЫ�y��]%Lq �ҵ��:�0@�3�ylƈnŴ�f���Q	wM[�y2����(5�N�+� �׿�yr�������6c� �dX7���y�,A��y��S,M4���.�y�Ԏp��eˎ6vV�Q-���y2��ML�l�%%�,m
<$٢��yңF<s�6eq� L�a�n��B&�y�ˇ 0  �