MPQ    4�    h�  h                                                                                 �B=W��IP������M��0d�'�#�,-E�#�V�w3%���BYe���2��76�ä F_�NR.往l$G" c��^8��p����8OD|aB�<Z*s�0R�� j3���C���^��3P�e�˨��T������~B�(��� �ݥUlA��P�@��J�fI#(0���l����y�����<���:p�љL-�֜�嚚�C�u��ֹ᳿�؟}�h;(Cd��w��n�� �m'k�����&��G�WQ�y��']b��Ɔ.����]����W63��;�WJ*�1�H���S����:Dc�=%�xD�=���òɰ.�gc�u�Ӑ,����Z���]���ռ�Jw�',�>ԉ��d���_u%�m��łr|�������_�C��_��o�S�Qr��x���{?�T���GI�O��l2=>��� �5��h� �OЪ^��	��!�5D��FP�:p�EQ#{Xa��T��>ÚC���b���2r(�q�J�{y�s�9��� '����DR������v�m�h��Lߜ'�t�zcֶ�?�e�F\���n� ���?0q,ȴӛ�V/y�ԣq��X��D�f��("��=Q�@���̧R��acz�#��
���n<��S]�v�e�5R�Ɏ�p�=-�-[n�i�����j�����#�s��Q��\Im",k�*>ŞB����)��%�.2n��na������p��_z���_7)5�|��<�S*�ءf����;3��7k�m����d�o�kbK�ה)Cw�!M�"C����l:�z/�'J���W�k9��d���H8?7/����a`�ӯ��y�c>����D�Q|�C�}D���M� �޴T"�#�u��׊�4# �5��8�9�soٯq7wDS�/x�8pФ!�� s���Tm�r��6���p�:E]�����������}M�̐�3��������a��$�O�x���~���t���j%O�o\��$��7|i����c��;�pER��?0_����#��|�-��sn�BwU�>�h�'�d�@���d��A�5��%�kY��u^Z}R$�望'z���c�#���T��� ��ᔸ��T���*7��������.u$u�L��˃�]-���@�$v<)�1��Q��T�C]�fRv"�>2��
a�I� ���6ޙV�,�˨S89��KE�ixm?��Y6b��֞ٸ�M�ܽk�"��ۡx�V`�?d�I8�a�Y$��{i��N��
�29O`W��͏o)�qiqo^���#oE�x͌3E����p:�
Vv�%���C�$�{���@2��C����\[���9��14ZGStL�&��
�ǃ^���bg%I�X@��~ X}'G(���
_����%|��N���Keb�S�q���/Z�Eޓ3ů�T	L.�+��x�Sb�����Q�E7�?�y4!�X=�Hy�0|�c�}�}��z����ؼ�m�,&Ht����'t�+�RǍ�W+�#^k��E�|�R��k���Vd��3Ē!�A��`_,=���@���(��>��8U��͞2lo22l�g���|Ѯ��	n����e�s�x�t+��`������_�����G��jZ��n?7�ؙ��M�~�rd@���i�g�l�?-��ǥJ7�GY�W�i`&ֹ�酻� ��s��F�=���P#u�L�<����I������$��0<��W�B�tyq���ոǘ��kDD<�ڡ��VԧJ=D9�U}�2B�>rs��I�]��{����T0���(/s9$1�^��#qH�i�<,�"�-^[���cI.�琺�Rf�`�mXq��w��0� ��H�U��$�� 6J�AφK��5�GfS�㸋��� C�5����k�4yI�p)A;�c]�H6�1�41J!�`u�w�whIY]�����h
l�W�.��e�-~o���
"�s�^�
"sgH+n�c؈�ŞO��^L�V�cC�n�!��_���;�D�_�ʍt��0�f��Oނi1b�ď�Y@��/��3��J�v�D����F46�A��j�!a��;&I���
��W"��jdr���N�:�ү��U�4����xщ�vo]��'�NE	o�h�7�WH�K#�e�0����W,��R�b��jH��[�|�u�刮AZ����������z�*��=-��ݸzW�˩q(G\>���cჀ�t癭���W�A<=�N��^JW���0���V�r9�^`��؜Mџ�`⢺\K"�}t��Я'��XØ Җ�<�R��I��Tmc���kY��2SL���ȥ�W�%�1v��ݜ�/I䩂Vv��Cd!m��2�iQ�?ؿ%�48�4����l���y�]+���nV��*A��Y-ϴ�q`دU���~q$_`v�`�9�;�P�F��e��{��tZ������E�c|S��]�^zb*����{���Yr�TQb�*sf��F1��w�1�x�ψ=�GH1i����&�(x#L4gY٢���=���q32�vnE}A�.V;���s#>��K��譀�䇹�SK�1ON)�kIKْ�����J��	m�q���8_Aq�A'Es���P�t�?z� 7G�ph��3�
4��FҸ8���4�ZK��ԭ�����V��+�Ą	4�ZO�#T����X��g��.·�7Cۺd��b(�����ou�������⍉�g�������#'xʅ�(��]J͔-�m��	� �������MΝ1�thJ��|W�$�M�񨓲��� �j���eM�N��ȃ�g�����Ġ����IO�������p]�p��'l��`���q��aaq���rb�����2/42�^�7��ɫ\���~g3� `�%����cW?*���Y�CΨG�}�E�R�z�JF	5_��H-0�D�X��"���0��	�߫��J~q�v:�JiLRqsG%�x��J*�4�|�i0��fF@�Ӿ�u��d��|j˾�U� U�.s��L���iK ���� :��%_i��a�˹���lVg��o��A��߹����y�L�~�*�\]w�P����Mɔ�_��BE�o~
y\-!��K�n��h�&�����Xuc�|A$�>9QQ[2��.e#��'�Q� m��oĄ2Q���}�j`W��O
Z���F%H~�����\�V�.y:�#35'[<5H����Р�����y;��9[��3�G.kL����L�Ǣя_��G��)y7��/�8ZC�'h���P��{�����p�PeZ.�2��،I���3�ٕ�(��,PA��xbz���U���\�����x����fɫ�g��+0���/Q��6Le,�����]'�շ�%wlH\��^�Y^��@2���%��=�mk������|�p��c���z/��xx!�J3ʶ���r�z���ӥ?%���q�b�jJ.l����w�W�;85P�í��zO+sM�|���-4䍰�O�[���u�DE�SX\
�Ty��U�š���@���K���J[�y��l���ϻ�\��vD����毱=���9�G�'�z�˶
L3e(ց��FF�CzIun�0 F,#)��OV?y�˳q�g��n�f�RX"<�YQ��x�
���,�|E9��6����/߮�p]�������R����==�`[IE�Hm�����cJ�sQK�QaI�ݘk�F.> %��$�G)��)ǉR�g�vaV��$!�p�h�_������85�H�ח4*z��fܡ�0�m3�W�k��y͞�(�_r�x�K[�)^�!�U�C��d6������'�h�W��)9����\.H�7CፕC��[���vN�4&>���wW�C�:��?B������#mX��E���!ib��s����٪4aw�u/3�zS�D��H� N,�q�m�XY��ľ�]	��=���W"����ˏ�}�4����A��Yt������\џV��S�ƹ�|�	�ƎO6j������:|�|n��<5�v��E�q��:	�_L�鲿n���i?���������A*U�%�h��Ed5:�Ө��\j@����F���NZ���/�'���M4���7T4< �������N�_���7C_���P��߅,u�J��'Ju˾�X-R��@?�<�R��ҫ��ѧ��cܣA��v]�2)b�a�
�{^균�p�q'�,�5�.Зʁ���f1m:��B*%bk{����MO�,kҨH���a[���:_��+a.+)Y��{D�N�;�
B�09J�0�*<Ϗ*�q6,��(��\7o���'r�E���H�t:M��v�l%�C���{�ua���	�>`�9�][>��9��1�<�SO~z&!Q��b����x��	g��SICA�S�>X�YG>�[��SYZ!��W��7PN6�H�ƅD@�^S�v�����*S�Ġ�n3�X/ �	��`+b�����躋@���Z���_W?V�}!���Ç"0W�j�}!����`��n+e�(��&c
�Վ_���+�����y��~��U�N�������}����f��G5_g�g�ۜ����;���л���U��͙g�o���"����(�^DV��{�,O�ef�x�Ft���v��1�չ��۟2㮂�j���i
�76l��&љ�xd�_j�Dz�ϧ�A-;��E��G�!�$a��Ԩ�6�f�����Y,D=OcCPքL��ufә��ɑ>S@��fĆI&B6��q�<����S�ة�2r<C����76��9���}�)P��r.���#U]��{{:��&�@�6(*5�$��ݓ׷�qc^civ�	����^�� �I)v����A���{�V���R��k��tRU���x
J@�.�f/�5�$�S^pO���w�8;� >�H�6UkA�I��A�$c8�6,C�����!�N�����w��Yx�&�j^�h�NOWY4�kn-y(v�X�"ZW&^�e��%�+I��c���9��Y��Ա��C��k!�?q���;{;�ʳ{�(P��^���ʍO�|�1}�*�
4W@��4/O����E�����(�{�6^���)�<,;a��B�x�}<g�P�E-���iӎ�M��Ə��o�w���`ф<bo�x3'k��	���A#�[M��e����#+�1	ҥx}�������6��UuS�p���d�����e�&I�ɥ�g�hھt�z�����G�n��D�L�3Ztb�u���"�R�c=H�i��:�WEE@������ӕ�7�9�����Ml�m`�I�\����8�7��8���;�s\+���kRc�ၔ���D��&6>���~L�(Ȁ�0�`F'�����/�� ���^àm�7��D���z�%� 48�4]��������:!ym낛�Zn��o*��[Y(���̒گFg���$�8ՠ;ws�vg���>eė8<�ZS�A�۳qE8�cW潛�
����]��"�{dn�Y��qQ��sA��FW*�]�1Ĭ�����g�i����]?x�4"g��Mź;�=�5�yOP2�G/n`^53�;rEps^M��椖�J@���@S(>1jԌ)U�aK��%B��X{	h~˧��_�0�AB���q�rP�^�?�@������
��F�Z��\�����K�j�L$��؂���+��]	O���(#/&����˲v�A��])=�7�;g�I`�(���(�u���{C�o�,�Hu��A;͌z��w!#bɊ�`�]�X�攈ĸb^��;��\�����Y��m`�Le����WX[� >���{�)n� wV�.�Mu�N�å\g�	k��Q���¥�����z%��2]�<op��+lgU��N�0�����<�G��b��*���e/���u��Ā\On�YT/�[��%n�e���S?�mJ�'m��,	}��-:Ӆ�85���H(~YDNf���8r�- C��_ݫ��~�~7:YwiGk����3��e�4�ٰD���l�n��u��`a�j��v�pa?UL�spM��#U�S�5 �X�=�����i2 Ra$�Ѓj0ZV�Fu
>A���l�U�=y��q���7Ltw����w�M�|�B �~%��-��~K�L��=�峢����3h�cyw�A?W9̳s[�c.���+����c$�o
lQ'g���`2v�OEEb���4%C$�aX��m�V�@��e2#�[w+]�F|Л��2�;S�iTn*|��3��~�M%%����o��b�G��)�5ؼ �854)'��4���V�v�m����$.���S�F�ho�3-�K��'<�'"��9�Q5�g�p���3��k�P޳�B�Lv�ɦH�g	��	���ِ@����]�{�ղM�wǯ�ʝ��t�����u_m�ǀ�Ș|H��u�ɕ����%{ɶ���r%���ѫ?����,��م�Xl($G�R�"�v_a5�����0O�[��7��H���+�g�6b���E�DXW��T_���!;���(�� ������i�J���y�S��>�vW�
`�DHj��m���쬶��B'M'kz���%x?e������~�00�:�,~���
vSy��Kq������f؛"��Q����e\���B։�GpC���Ե�joU�T�]�lh���R���
+�=#�^[$库T�Q����6��.Zs�Q49�Ic��k���>;����U�)�*���"Ia,���G~p�^>_�>ｕ�`5�4���~�*5ff�O=�W�3���k2g:�9� �Z)���w�K{�)y��!C�Ca�q�;Ұl��a�k)W���9�l����H��7~�}��νV���:l��>�~��:e(2��CХ��L����
1#([��k��*>�D�0��ن٥Gw���/�enڀ�1q )w�eBm/���ri��vڰV�O���U��Ļ��l}��w��SL�I���ADq�x#����.$����ڂ�4(���O��`M��f|_F�k5{���E�.�5*_���z(���Z1�r�A�_���`�U4,Wh��d�S@�c�/�wF��oV�!���B�2Z����F'0���I��c�T��ж�{�W���u����7��v�L�%��7�u@���O��(�-��@zz�<�� �����n���'�ҕv�%2��a����#(�[�f����,���	ח؝�Q��m5hm��b&w�rM�i�k�N��}"���V(>6V���%*aI��YD{;?N���
��g9EFׅ����,�qQu�g(?�dXo�mk���bE�B��FY:$Wv,�2%��pC`R{���v���9]��'_[�")9�-�1*?�S*�X&\�G���:�uy�<�1gwR�IM����X�VGy8�;�_U�����(�INQ�{�A��#S#/еG�O�%�����3;!�;�	B��+=)���Y�&�E�ă����?K!��$�>��02�?�}�����T	�ɞ���6&~���	ٚ�ݥ+A��� ����Μjb���.�t��af�X�>�?��W���e_����ϒ�������(��'UE�͔�Ho�����`������ٞ�˨%�g4�emGx
t��C�ր��LGB�����z���j����d�57�M~�\Y�Ѵ0Gd6P�zC��Ɨ-�N�@��G��߁����ׅ���{�c۔2=�0�PW.L`]�0������g���܆CZIB��kq���hL��3H��@�<�]���8H��U4o�H}�@�>\r�{��4�]��{V����M۲(%�$�=���q~Bi��R��*^��A7tI$#��F3n���n��Z�N���-�u���zU���t��J�汆���5y"�S9��ӊ 9��u�k��I#��A1Y�c+G6g��j�+!�\��-�6w�9DY�E���h�QRW������=-t*ϳ��"[4^��ix+$=cN;���P��Tt�"�Cnl�!Х�y�9;V��(��KN���� OT�]1��ą��@[ܬ/�p-�i-e@4E��ge�6p�63���`�D�k;�=�ݜ_�xA(���'�����j�Ȥ���&E�$���oH�'&��	��&�-r��ڛ�C�e"`��I,&�`����Ͻ`i��A���u�Ո��J�Rş�ix}�A1�� ������X*�z��0��(G�������t��I��}ߍ�=�����6�W����������h��U��OQM'b`�|\O���7��┡�|k�N�T���R�Oс�X�u��2R��:L��.�[����(�翍�6�/��W��e$�yB�mx�����õ�_%(��8C4��r��谁ӤWy蘆��a�n̠*wݟY#���'�������$U1 ����j��|lie�U�f�uZ����6E�{�c2�ӛ#��P�X�wʪ{"�Y��QX��sW�F�C����1� ��>�j����i(	,�7�x�=�g���U��=�+���M-2X�n{_%�W�;M�
s�|�Ձ���4:�=�wS�|Z1��3)�*�K�0%`K�ڀڠ	c3��]KQ_��A]����G�P�h�?����6���Pe�K�
�d�F�����pMKU3�����#���+k�z	jIVP�Y#
��5P��z���h�7��������(w��#�<uX�\��ʞ���$�ī�a	�-�#�:߅�9@�S������VDo��(����P��C��O���M�W���A���%���� Rb��X�,MMž�(gQ���e���9�<�?����1A�*š]DTp��l� ��B�KI7�g�Z�.����bK�0�~e4/��J��7��+��\����4a[ǖ��%	Oȝ҉?�o��t���1 }v������5���H#�D��k��ÑH��Rǫ�^+~�<l:���iB�/)ح��6�����4|�а,�ܸ-�	�nu��xw�jA|���'�U�!0sK��^)�� X �'-�=ɋb��iM�a�T3�E�V�%���A� �o���תy�dt	A�[Yw*�i�7,Ms���B���~@g�-X�K�n�3i�N?	�2��c4�AZ�9GiB[�=	.��]����V��~�o:��QBc��sԚ`��O�Pb�#6%>�1Ǽ��=��V��o�z#�Z[�A潷#(Ж�̍9-;t�o�q�(�3��^�n�nW�:*�>�GlZ�)�S¼{��8E'��`�<��q�U�k�����.�$���ŏ�C+3h푕(FI�"G��� �6��M�+@FM����}���4ɡ�gte��mK$�2���a0��C<�]]phխհw"7E�X$���ܵ6-\Ӧk&�m�>I��F|�� ��r�ɰy�n	�� ��L
r��J���?ی����٠jkl�ǭ�-�]ױ��5�/b��y�O�c������c*����� ���{cE"�LXRR�T��w�˿T��dv�6Z}��L��"��J���y��uJL��1/�%�4D���H�֯'<��lJ�=]�'���z��b�@ĳeU���Ż�����0�O�,�qx�ŵkylq�)��"�fH}�"rIZQ}����;"�����i��a�k鍇�0��]���v�,R>m��%8�=�E)[��ۓ����;X��0 d=s���QO16I޴6ka��>v�;�Z�)�W&�?�zݴaG���Xp�ta_+u�0��5�@��M
�*�\Kf�&�V3���kmC���\�U �..IK��S)�B]!��?C<r���z�K;������
VW?�Q9��R6:H�#x7��a�y Qq[�,GC�5�>���ez�CS4�uk0���ehf#�}�����(���ڪD�&٠�wU�/����?���9 �@Ox7m�-��@��r�k���p�M�i�~(A�r}�A���R��������5�Lѕs�	�E�/�̂E�_��65O�eQW�5 �|�/��FNq���E#��0G_٣�5��lk�����:_�6�U�Rh��9d�g�3>��B������k(�}�
ZN�`���Z'��7ߔb��JT*��Б���4�r=��&7�]c�&��
 u�U�ݳZ�4��-�[�@u�v<:�H�H�B��+��?��A�vӉ�2_�^a� �1	Ʒ����Wl,�Ų�(N�@N�����m0Y>�*�bᒽ�*gME`.k���:�@I��Q���5�z��ad�Y�M+{��N14�
x��9@�������^�qlްⴡ�?t�o���]O�E��q���:��vGa%��iC;){H������4z���`[�jb9�l91�a�SBG&���!�|]���kg2%I9w;�IgX�scG��ֲPg/�����*Nl�v���3�Y8S^�}���� /H�V6E3�	�V�{	��4+�I�(R��K���<�V`?�t�!����0�(z�%}W�d��h/�$2��1&��XՄrP�n�+|�0��:���Z�� �@B.��5���J�3Rd�z�Ò��.�{�_��n�v��>͌1%J���G�(U�[�͏1qoC ��6��T�˃��9�e�qxVit<;�㑫��g�V�Pj�U�-����j+��_ g7���"�ϝ�d�`f���)��A-q��;Y<Gj,A���;�
9��,c��Vtm��XV=��P��L�J���r��FX�4����2��~� Bl	q���7��ɉ[��nF<9O�}Y
���:
}}�w �!�r�]��O5�]�p{1���Dv�P( B$B`|�Mq�q�F%ils����^,w��SI�硟����(��I�Ɉ���f�n$ݪ�;U�%��φJ�iY���}5�?S��C���n�� 4Q��Кk��|I>`�A���c6�	h�a`!��Q���wE��Y��K�`��h�t�W�Y�S�-o�����"�~�^�{��"+�
�c�ħ�o�O8/�geC)�!�+��;1�@�\�^g���[=�w�rO��1�}1� =6@6 �/�z��E;�6�U���4�6N�t�����;��G�x���sfe�X	�a��A��C��|c����&��{��z�on7W'�~x	�������qe�'�y��F��$���ܽ�)[��J-��u�9��s��
��$i��\9�ɛ����=��� �z(6ש��Gm/���vm����tX=*��i�Ȅo=~���R]W�[��M������L��%n�=mM���`��6\\ˮɔ�!����h��)4N�I��R�.��
$t/לOJ���L֠�6����*�G1^�γ^/Zٮ��_���7m���f����%�I�8�94b�@���.6ycf6���|n��*��Y� ��W����đ~�$�I���׏썱��le�3F�V�Z�7&�T�E�SclY�^G����cSŴҒD{���Y�\�Q�N�s��MF�|��9�1�t�ϙ���x�iC?���0�x�fg
F���R=�j��/l�2��n���+��;(�us��i���>��5�S|�Z1��B)K��Kj�'����|>	^󧸿�_r�Ax�K�g"�P��?0�l������M����
e�F#�%�R��K"�KR�0�U�����g�d+&��	���@W#���pˮ��\�	�O��7t]4��9�?�E(R��^Qu�l��]�%�
⾬7�g$͂g��u�#��ǅ��:�NNn�>;/ث��q���Rz��gp��N�ۊEsC���W(�~�������� -�w�\NM���ŹIQg�,�� �N�TR����èM�ew(]��p��lΡۑ���f�]���J��$�4n�b�Wϑy]�/E����F#\*[�����X�%���L�?;�$�����V�}�>ϛ��@��_�50�Hz�DᶳS
x�c �zf�����~":���i=���P2�������4�7԰�YR������`u���҇�j��l���UB�{s&�~����|� �������ih�3aI� �V%@�A	\��ʈ�����y� ��Hn��.we��խ�M�S�p�LBv\�~[y-��Kq��?H�����������c��\Au�9�>�[���.$�������1o�u�Q]������`�zO�{����%9�=��q��vV�K��#�e[�w�R!�БT%��	�;�O����r�3ny���¹� � �p9�G'�)ʑԼ��;8�u�'<A��j��lz�Ƹ7��.�Mv�I%�Q3�D��Ä��&T���������)�+!��)a����Pɜ�Jg��0au�?��~��a��~�]��uը}`w}�������H��ZEӁ\zaF m<������|���딐���N���n��j��?ϚrS�롈-L?6�[��*ٻ*fl� �	��[5!���삐O<���A�~�[�!�������&�E�emXM&�T�Æ~���뙱�����Վ]�eJ,y|/������x��@B D>���#��b�ORׅ8��'Z�zO��[0�e�D{�_�m��HXF�0�,4FZ���y-qq��ܓi��f�B_"�>Qx���;ԧ>���ͫ�f.y�F����>劗�]����ߩR�⺎@e=�[ڄL��y��^��Ba[��s��|QjI�IY�gk<��>�w!���G)|�ǚs�@�ab�)���>pq�_f�����5�lNר��*�s!f-G��3]�Jk�?��o�Y�P�j܉�K���)�$!9��C���ɍ��)>�o�!�W��9�Բ��}�H�Z)7��9�b�L����se�=>"���0j/�[�C�2��0��;����#����d� �.����$�ͪ�ٛ=Gw���/d���Q�b_ ��B���me��.S�n�2�&�]��9�za�|��}���ХU�������P~�2z��:�j%S�������rOG�Sֿ�Pf7|U9��!��'t�E��%�+�_]!����#��hJ��C��q�;Uj�5h�ϽdF�n�ٷ0��^ѩ�7������^�Z�X���~�'���O�R�T��;�l3��ͩQ����\7Tp���F�0�u�������o	�-#�]@pP�<��Ы�ŉ	��"����v\2���a"v��ķ�9���,� ���c5�{����-m+jS[�b���E�cM�v�kc�y�u���Z�L�����5�a�Y�>{�<�Nl�*
~9;<%�;oV�[�^q�g�]aP��So1�����E�H�Y��:~��vb��%x��C -{�\ݬ�l�/���J�b[oҟ9��#1 ��S��E&�X��3�wweO���g��IT�4����X}��G�Ȳ�q��K:��h/Ch%~N��9�7�]�A�S���}4���Oı�@3�8q�	8��+�.�?5�\��5�����?�r!)�,�4s�0������}����q���Y��&�����+2�W+��f�Vƴ��"� �l�������WO�Yֵ�k�����E�_x��)��w��t-[-����U{�c͊�o�CH�S�%���ԭϳW�^���^e7�2x�dt����L�*��k�5��0���3��j��1�Z+T7GBc�����*<d,�����_�X@-tͥ6O�G����U#�%�f���!�1_��
�= ,;P�uL�#��Ɉ��+��F۳[Ƚ���KB��q��vC�Ǆ �׼�<�`Y�X�|�6���`}����W�r__V�jn]�D,{�>�@�H0�(;�$������q�j�i�*��#�^G��P��I���+ǟ>��XAD{A��h�M�E�U��r�*>HJq%����5o}ZS��3�~��	�� /���+}<kr+�IYE`A'J�c�:�6ݜ"�[m!�����Bw ��Yɖ:��xbhv��W
����;�-j��i,�"���^7l_!�+��ec�m_�
���Jv���0C��.!ҕol�;�Q{p[������
����O�)b1�!�{�@D/ Ϛ��Z~6����~��+6ir��V��~�;�e����n��a<�^�7�����kW�G� ��Z���u�o�F'�y|	�X��#}�D���eX��	T�� �֩���V
��� chs�u$�%����p&��y��wa����د���z��u��tGȿ��uD��@tӳ�^Q���S=�M��FWV����:��^�����IpM=.�`��-\����i{i�<�"�vu�������R4-��������W�&��qL�-�\�M��t��PB/��B՝���Omn�(��X��+�O%^�8
��4nwq��m��	ټy�S��g{VnB��*�<PY�<���a�Aّ1�$K������'�$�He�1��Z����,�yE�b�c�^O���u����N��-{^{��Y���QNms�r�F֭.�_1�<���F�3�Zi^�$�J�x��gE��ŋ�=��ߊ�'2��n��)� G;��s;շH��hB��S7�?1���)�i3KEN�9ڶ=T	Y���Tj_-0�A��N�� PZ��?kp;�l)3��ҷq�
 ��F>p��1U&�K�Ub��&��Ҽ�z+�ۀ	�&F� #�����f�G_��Q:7/%ЏB���i(-����uUښ�~0�����y���*����/�P��#}D�1�M�I:ܔ��Z���ጀ�����BPΉB'������Wi��9���8���Cd ����#DMFIRŴ��g��۷��o�i�5��Ã�H��I�]z)�p�a lx�#�L����]Q���(+�oKeb���tu�/����J�ar�\������C�A�%?���/�?��q�Ep����}u'_�����6S�5�eDH(�D_Nb�#��~0?���_�`��~]2:*hli8v���6�d^N��֓4r��էQ�R�k�?�ju�B�-Kj��ݦ��U���s���1%$E �%�N�X��L]i���a�]݃��VSD/��A6��%����@1y��j�����w��S�H�\M�6���B1,�~vՒ-��KLڭ�z}��،����DV�c�'�A�Ȑ9=4�[�g�.QdF�
�L1�t��o�[�Qx}V�i5�`�YO��^�YQ�%4�%�rHZ�_xV3y{e��#�`N[(�T��>hЌ%E�C��;�K��g�_3I�W��T_��R��T�G�G)���q��8���'T�Յr^�g�ڟ!���<�.��N��~��`3޻��^�k�X��J~_fP4��H�z��zl�d�Кs�ɗ�Wg*~���Z�4����ѳ���6J]��գE�wإ���iX��\�,���\Y���m�]t��!�|Yzp�O�d��C��d����zrr��d����?��A�]���
Il�n?��d$�'
�5����:O��	�hpޙ�>�������x�a��EXF�XHDTp���A]t����,-��y~���V�J�L�yw�n i�ϧ�ݱ[�D�We��q������3Qm'^#�z
���v��eTQ�:��/#��4n0��	,�:<�;��yH�Dq�J�DVf�'�"�B�Qs��vZ���������<�!s·���%�G]��s�,*gR�x!�[�G=�#[���u��q����m�.$s=�Q���I��k2�>�}{��^�)w9��S��a}"X�{1pL X_�=�fi5�����*f��fHl�38��k�[��
���K ����KG`�)�3!��C�J"�tҁ8
�Q6�|-�W�6
9���H��H��7/����LG�"��� ��>=�����]�C�o8�������7�#Y#:������Uu�_��zh�ٖ�aw?/z��i椈�� ����m �g�<���~S��`�:���C���Ud�H�}T���~T�Z{��r�/�k��ы��;ƥ�m�{���^�O����NX�k��|�b*���m�b�EY�u�&d_�U^����>㾚��F|�~?U �h�	�d�_VӔ\�Ț|��MJ˲����Z�*��փ�'A�P�
L�� y#T �g�G�S�?���{���/7�ܜ�}{�K�u����� ˪�N-���@k�#<�{�����-���%ң���vI�u2��$a����3"��
���~,x�������	�"��m&�����bW*�`�hM;�`k>  ��a:C G��Gh���y�a�cWY�0~{��N��P
�d]96�זY�"�q���-K���ol��͓��E��z�ZG:9�v}$�%�C�!{�>|�G�}�*쥼d[*Z�9K�1��S��T&F���*�r�$�M�?g�*wIo+��?�pXX|G*����F-��Á0#�N�J����S�IRS��յ�
��3��3l;�T�	�?�+��Z�z$����鵾�Ai?B��!D𼴯00�Z'��}��x���ϗڸG��&Ϣ��z@�n`�+��P��q�
�&�{����y�:��s������(��/ _Ӻ��n�� ���'�|6���U?tͅ{6o����G��2�Jnp�9��>e�Ҍx6�t�z�a���-x��:��F9�n7jaA�Uv�7��5��-��bd���9�ϓx�-�6k�1eG ���>�@I
�"z8�j��E9=�Y�P
�Lq�}�a�"�2-�*-'�6~���M+B�/�q�,�ynf�?�n��*�</���3���qjc@dZ}�E�O��r�ή�Ǖ]�3{�5�{�!���(}$�B��ê�qϮ�ibⷋi�-^�0��c{I���W���<���J��p��hyW����_�U������J,���ץ5��ES�㊋��!�9� *w����k-y)ItJ�A��ec��6P1�;vR!�F��>��w�c+Y��VlhQ�WEmd���{-eL.�Ąq"F&w^'S�_�+�pc�6�ť�E ��L�C��b!!�G��t;�^��Dʔ�����r�-�WO���1�X���E@��/;���:!1�-��[�g�6��������;M�w����iT��@�aZ��/0�9�p2���[�&�����p<*o$v�'W��	�ʰ��2���|9��e�]�O:Z��ґO��dO��
!ۢ��~�u�����&�c���ђ�\ɑ5,넓,�	�z^����G#p��0Ξ�
@�tNJ�9���>��=�:ʵ��KW��B��Qv�U�7��`��'�� v'M��`�%a\}�$M�W�ա���ߋ����R�K���ο*JC���'�=L����h��L��}$���/r]������m�ċ�j��f�%�#8{Z4�����ु$��yYa��B8`n}I<*H��Y.5�8�d��|2�L��$��I��V|�b4��Ml�e�O�w��Z?)��Gt�E�c�q�����!*�Iw����{P��Y�R7Q�\s�0WFCO�ZS1����O����!iy����Sxj�g�.�&��=�H���E2�.�n�"!�;�ԻsJ�p�R�蔲P�N(^S�:1�D�)A9�K ��s�Q�	T�n�_�oA���]7�P5F0?��vj���\P�
�d�FY#b�H��,�K�ȭ�jB���d���+�1j	�:���#�e ��!����Ʋ�R�7��y�3�5�y(x�ԁ�u�g0�w��_��4d��.�x���+�#NNU���x�DFf��1&Ny��N��H}��W��'�{��r*W�t�f��/�q� � �E �	M�Yům�gb����Č��z��Ԑ�^5��;]c�p��l�ƥ��C���B����Ө�A��HTb�ԑo�I/�	�@d�|�e\�����G �GI�%�A��2�?�6�� ��/}�/���٪�qf@5f��H�wD��m��[���c�p��;GE~�7�:�M!i30:���"j��(4�T���៍�����uߦi�.jr��9KU8~�s���fi�� �T�����&�i��5a�$��0V��v�A�/E߀�t�A�Jy.��'��G�w�D���)Mb��&N�B��~��4-�W�K'�e���^�ղ������)ce�KA��I9�I�[y,.��4�.y�ӧ8��M�oka�Q�:����`�u�O12[��#K%/����-�n��VN!��S�#z{�[cD:��|�Їa̞
{;?g���wh��3$�`��R�����&��G��) nq��6t8�7�'�4�rn�bw�|e����. o�?4��?3S]��a�������!���\��RG�A�ޟ�蚸\�ɒ��g�:���u+����%����].X՞-�w3��ʉ<������7v(זqmr��Զ|����
,�Y�������綵5�r���~	]?���ܾ��
lrj�ׯ�b؏5W�����O�<y�#�u޴�)�@���㜧hE�F�XC.�T�R��[z�.�O���z�TGM��:�Jb�)yr�E['��bl�v�oD4<9���W�ة9����.�D'�^zŬ���h�e�������j||vy0�N},�N��4�yc�qw�� Zf�,s"C��Qn��љ���-��%\�����6�V������]������dRo.̎vI=R[���@�-�DY��V�'s�NQ��8IOg�k���>'�I�+Lu)r��P��]a�e��!0p'v+_�C�k�5�$Y�^l�*!�fcH��]�3�tk�FͥG��FE��?�KB�)�-�!/D
C�u�]80�g.~S���ntWp�<95�J��lwHZ(\7j<ƕJuBx@�=,�ۼ�>X{2�&�f��C�إFl�KĴv�D#��2���>�"�P��Wّ�7wf�/ڇ��.C�~ ��7 rm�]��j��$l�ڜ�6UPžc��0����=}�Pp��wO���5�-�ن$��X�����7���"BO�#L�N�R�|K����Xt�|�E����!��_�[�fO��Y_ʝ^S���j���U��th�c�d���O!±�����,�ˍxh�.�LZ։Ѩ~'�n��ś��;��T���"�C�U(����7
��8V��f@�uV'�n��iN-YR�@f�<K���yh��H#/���M��Q�v���20La���By�G�)���,��u9T��p���:Xm!�	Qb�I�{�uM�k&��BL7B��������a�A�Y��{���N�*
I�t91������ѳ�q�فS��Ї�o��B�.�E�J	�L�:��
v��\%n��C�-{�@����%��� �f[�'9*�1��S�Ws&HS��i�mՕ��.�gc]ZI��ܺo�X3�PGe�F����A@\��]ހ�N���-��qWS���)��i��g�W3'�2��	.��+����RW���8�g7�g	�?���!_;U�*��0���+��}(F'��dJ�5���;�&��Y���y�I�C+-=J��f��=q���+9�M���m��+/8��75��8�_.r����;��s8>��u�U���̀P�oT��ɟm����H�HS	�em�~x�/tM�!���=����u`a������j����P�b7��H�H�� �Qd"R[�������8-B�,�>G{����D��[���5;��+ۀ��=V�cP��L�X�A�M�ꑥ3�T߆/ߞB=�qq���Թ���Mn���<�㽸|q���ۇ�}���$r��
��@Z]}]�{¸���*�G-(߇$S�z�~w�q��i�ɱ�D�d^����]�I粤 ���o���:�+����F��{�U��B��J�(��65eX�S���~��?	� %:���lk���I�o,A��c�6S#��ְ!|�꿙�wv\�Y������h,��W�K��$g+-`�����"��^BBU�h+�4
c: ��@�h�@DX�x�WCZ�:!<~!e��;�7y�8u�/z���g����O@=w1���q��@�+�/v�X���,\3�f��"C�6����L'����;��}�I#��d��e������,���斻D��Q��k�"o��'��	]���j.}te�>���i�U�L[ⴽL+6�}@�ީguZ�ֈ��}���-�U��ѭ��+�_n�DCz�Λ���G~@���}�%��t� �=��y��=O�^��fmW~���p봕Tb7��X��;Ms�d`�l�\m(���>_�r�Сl�#úg��g]Rj��{������e��B�qL�<����~���A�	���}/k��'��~mdd싋�á��%�'8 #U4$��qs�?��yԎN��n���*��Y����n����ϑg�<$AS����F�����V�e������Z���b4]E|��c�����:��D���{1MY�|QDWs��F~�
d_1��'ϪQ����Gi�����FxE�g��2���=��+�@�"2DxHn�N�);��s�y���U{����S��1��)�(1K���Lt��� �	OGѧ�܃_��9A�o���qpP�u?�����9�����O<
�O�Fte���n�`�K�a�&B�㏳�x�+W��	�=<R#vE��!���}�0��\.�7��2����u(�"hGu��� ��6�����	���:��E�#�?��gܻ�?r�Oݑ	����<���.������ۊ�5��i�WK%�	�Jʣ��� ��,�D�M|�Ū/�g��ҺQ���>7�+�9M�Nu]���p�[�l.�'��a��E�SVdӃ�h��eWb�E;�j�/V^3����ɗ��\xb�ؠ��ǂql%uM���UH?L�̒��8�J�M}kX�t�Ӭ�5{!H�%D�ٳ���o��`��*.~�u�:`S�i.�}�y���
��l�4h'��� ����u��u�*��1�j-w���2U��gs�)�J�aZ� ��=7�N �i��"a�淃�c.V���_�A�I��4'��)HyI�`�~�~�Nw��~=nM�Fp���B�+"~��^-BK..��G.��p��1d����c =�Aƌ�936[T�.�DW�� 7�"��*(
o&��Q�4�_�`yOl�����%*B��(3L)��Vi�[�#U�[�ړ�#ڈЂ'y��:�;��!ۭ���3�ʁ�3�Ѝ��,���SGX�)��g�R8|Ȝ'����� �]�O����o�..��ݺ����Z�3T
��� ��� ���������Iw�(���G��Sftɍ9�g�7�LT��W�w�����/��]ɂ-ՙ5w����D/��:}�"�	���o�m����T|���ũ����Z���l�w��Er$Zߡy��?GB.���0�+�l����j�ם��5�E@��]�OM�h��wV�ϖ��y��}W��נ�E�g`X>bBT&ͅ÷z$�I}=�"�'�/0��?�J�Cym�X�������D�@Y��yx��l#���)�x'z��B��4�e
�A�����7���0��l,E� ����y~6>q�_?��	�f4R"޻|Qi@��,���oxD�2M�~Ș�|χ� ��[ޱ]}(���R*����=�GM[k��{˶���	��ly�s���Q�Q_I��k��y>b���Y )m��ǫ��ɣ~a�����:p�_�U���5ٰ׹w�*�w|f~�o:3��kY��@+��A��ܚG�K�C�) g)!���C�a���ҷ��yu�2�>W+0S9P�2�>dH5��7��z��.Z=eگ����Ԍ>s����y��C?J���=�����х$#�H�Mm��1I����	રg�ٌf�w��/����h�~�? p.*;Um6X娸��y��W�9p g�970���-e}�����F����V�١�Bс-��u�x��^��.���OX�������|����*��0nE����C�_nR�!��t�$������2�"��U;-�h��rdW���
a��r�y,��hg��i]�Z�-����'�Rj߀��V'JTd���޿~ɗ�����7e�V��PƁ��u��ߓIg� J�-�9E@a��<���4��c`o�yƕ�cA�v�v�2�qKa���������80,nC�Pԋ�,g��X��m][d�@b�A+����M1z�k�k��&D��t�=*��c�f��a�?_Y���{f�-N��
�k�9,�6�L��e�q��W�&%��#�o���ɉ�E���j]�:��v��+%�K�C�t�{4cB�}u� .��[i[��p9E�1�+�SqI�&������h=����g�aI�_�5]X'UG�ߥB�J<s�y���^N�T4����b��SJ?~�NԿ�g���ks3����4	�&�+��,�𠖺-�a�0����r?��!z����~0yvffN}����������yꊺ�&/U�p��$�l+hpA�')� W�1ZE,���Fz����a�f�\�^����b�_�mZx��V/�#`�[�3�UL���{E�o������9ӆ�@CF��V����e	x���t�x��}����:������|j�P��Kl�7X���&J�;�d����fY��	�3-�/�'�LG��d����v�	�*����ۻ1�=��P �CL'_���L�h�֑ Z��IȆj��B��oq��L/%sǵ$�(g�<%U�������\v�~}ۓ��^r�$���f]�'{�����N�ۦ(aW$��:�9dtq��iX����^���!w�Id���M�o:�F��s�t���#C�I1U�Ŕ�;$�J��`�ln5�� S�]ɋ/g/����  *�<�dk�t�I��>A��OcZ½6�K�q�!w�+��|%w1uY�w�L�Eh@�W�I@��,�-[s�z�P"�M8^](9�<C+k�4cu)���^�;���Ӳ[C�!W�#�h�;�0,M������ט��=O��'1����΅@��6/����p9'6������݇?6��'�ǆ^�;��w���_:3�r��������/�芐���v�+.L�f��o�4 '�)a	, ����Eӭ�DMe)������x��k��k�X����u�Cs��˰�`��l��ș�ɇ,�:iv��z��"��eG�0������@otD�$���ߴIx=�+���Wg	��9?��IZ�σ��[�"�v.�M�q`��{\�n�˚P�����Z�ÕcU�5��R驁v���׈�]�L��Ȣ����s��������/Ɗ�s�r� ��m�f��f�6��O%/\�8���4m`�,&S�Z�AyOܮ��n�Y[*~��Y
4Z��`*�rذ���E$��̠]�a��Zw�a�e��-�Z����}�E���cy�ћJ@K�W�,?��>��{Ƅ0Y/��Q�H^sc�F������1�����A�d��i�W���Vfx J(g���\!s=��ߛ%�2��nE��Z;�\Bs�H�ՈK芦����ShF1=�)78�K���N�ڇBf	J��$�_^OeA���S�zP�y�?��=o���	�o�
QZ�F��>�>����K>�/��9���z�����+=		��BF#QE��\�e�'���K�7` P!�ͬ+�](��Jn,u&�C홡�����⪛�$4X�n�C��E#�P3��:�Δ�����7��J��> >�ӳw�:7C��A�����WzAj�J�e��9� �}	�9Moť�g�>[��"���������Q��]K6�p�rl�?��}9׹�H����^Ο� �nbR*:�e}d/��}�{�rɲ@I\�_F�{�	ǽ�%�����?�[ڒv���e+M}�כOiU���<5�5TH
�DpV��?-5�πd�f�.��,�~�A:�xsi)���qE��	.��h4��Z�fQ�����u�Ζ>U�j�
��AU.�cs��c��.��M ~�_�ы	:�i�&Xa[���g�Vb^��!A��?�6�����)ydQ�ۆ\�Y��wQ9Z�+M�K���v*Bb[N~��-~LK݇�+��U.�����Ud�c���Aឳ9��a[/.��d�aɽ{��"}o��[Q�O�ڶ`T��O�hP�*)�%%�ǃXU�q�V��z�
�#0�[ِa��W�}X��T�/;����O^�y3��2�a�%����s��fzG�)6ʮ��]8Wy�'�˅C���X{d�2�m�m��.I2��5�s���m3��^�/���	�!�[�N���eL�a�/��*���pɈ�gg;�MԠ�	5��G�bi�j�]]d�Ք]8w黽��AJ����P����Mg�m�������|jy�G��7��գ��G�W�+&r���te�?��4���'kbl
ل�t����5�d���!O�mآ�+�������X���PE)��X9��T��Y�r�r�d�S��Y �
9��IcJ��$yh�/���I����D*e���-i�N�s��z�$�'o?�z;6u�� e�B\��>n��qp�Y�0ݘ�,���l�"y�qm#�� fo��"y��Qd���xݧ*�Ɖ9�R����1���p���5{]xN�=�R��펬Y�=�[FD1��&��B���ڼ�NOsn0Q��mIE~ek��>�PB�a��)h|������#a�K��Qp���_R��7|J5�\����*��f�<���3�]_k�p���.��<(���!Kxe:)�!%cC�m@�&#�R$t�H��Q�W��M9k%�̹ۼHvO7�@#��8r��dxQZ>������T#7Cz�U�|������,]$#��h(����fk����Kه	w��/P{U��C� K�lv��m�rO�&x�ڦ������Ŵ*���,?h#_}%<����9�k$j����ټ����kf�P���V�5�L�ݱ�
�O�
Mº(鼾�|A��������E*S���_� ���"LǝTܠ��F�]�BU��h�wgd��M��
���K�CvG�ZU_҉�R'RW��;��q�)T��4��Z����,�AN���P7�
䊮k:Ɯu��D�$lb�[J�-�A�@\|*<+q��{�~�w��Ʃ�>Q\v���2f�"a�yd��c}��<d�.�e,��+�3�g}����cm��\�b�����ѧM��k���ae�P��8pzX���!�a�]Y�tE{A�mNX��
L9'�ק��G7Uq��uIS��߅o�&�d��E�;�Ŏ:jp�vΠb%dÛC�۝{o��������qk[[��9`�1�)SL[�&���⟨c�L�^og�"�I�)�ܰj�X��G�i���P�7�&��8yT\uN�	�#Q�=!RS��е�^���I�3�u����	$��+_���+J����ˇ��?s��!�1�� m90T4^��	}^g��Ҭ�����EY�& �x��Qr��:F+��G��4���՛����ҩ�a�m�C�czuQ֡-U�����_���-��q{/�����hi�n�{U�v�vZ�o
U&�?���T
}��]�����3Ke�X+x�uktX��8a���3��k�ۜ$3��lj2��Fb7��.�{>�V��d�P�AZ�DJ�-x>U�"g7G1���A�1֑�e����J0���s=��lP���L������	��vʑ��S��_A��aBBs��q��!����pZ�C5<��Ҹ��&�"��/e}�jE`qlrK�Ϯ֒�]s�{xp��,٣}��(�$	�ړ�pq ;�i������^3�����I��h�z�*��8Ֆ0�F�ON!�ݱ��U�����[\J]׼�#�N5[�S[ʰ�jo�u  b��F�k^"+I�A�vc5��6�)V��!rPH�O
�w쭗Y5���h��W�g\�Zs-V���M�"w_^xc8K�)+F��c�R�vTk�6��.��C�d�!r�M[R=;xIag�_�e�F���>�PO�М1:���g�@}��/�g�5�"0S��2���c6բ��B�9z�;�f�&��Z�ܬ�tJ���&����äs�F���*]�a��o5�b'���	G�#�u ���e��$����k��� �:<ؽB���3 �T`"u�舆�tE����B��A,�����C���z/*���x�G4A��a���[�9t��A�ʨr��ʬ=��ϵѾW�D�����'�J��6H뱺�M���`�Zc\#���U�e��x��b���p_�pv$R�g��qd�;���C���xSLw�1�}]b���N����/!Gd�.4¾��mZ���A`{��!%ʰ�8��4�T���߁u�hy�I���.�n.9*{RY��Is�-6֑��$7���8N̏;��(e�it�I{Zp�����Er��cTj������K:��\�{���YJ� Q:�qs>*F�z����1����`X����i�-����x��g1{����=��3���2�k�n����;oнs�7��#�r�P��_�%S#�1'�)�g�K�	F�H��"�\	Eҧ�_�A�}���FP�C1?W�>�������m�V
�F�I)���7�*�Ky�1�\Q��م��.d-+��	�&2S@#,e���&����������7a�<0w��@2(�xq���u����B6��@x�egU?w���g�D#�� ��m��5*���Ia��xٹ���ԏ�us_�LE����W�W�%�P��߄�u� tI�ﺀdM�C~Š�gs3�Ǫ���&��!/������]�ϋp���l�,�81����I�1�9��[ �b�.ё`�/m��6h0���\n}o�VNV��!%�3����?(�1� ΀�}a	��*�"�"`�57_H D�Cѳ��ޑ�0A�᧡��OP~IR/:��i$�K�J�P-֡"�4^�A�>���ÄuВW���j���-lyU���sm�����n��� y����y��s�i��a��g��V?�GL�A���ߑG,�r��y�[Vf��4Tjw��մ `M�p��7;bB�~~�1K-�v�K��f�	�������;��S�c���A��d9)J9[
;�.=�8��oD�x���<0o�2rQ�12�UwM`/��O�3I��[�% ._�ޝ��bgV��JQ�#�w[g��Y���x��̯�I;pznt��O�3��sC�������׏7AG΢�)Q���]��82J'@�0��l��Sb���X��(s.d��ݰp��e2�3�؝�ʝҨ`����^R�-鐘hV�P,蚉��Ƀeg�/�|�ƨ��m��=;U����]�ˠՏ��wDʺt81/>���Ȍ���mCl����|ŃQ�;g�RX��P�6�"�f?[rZO��oC�?�\��IVA�B��l�<t�O���65(��ӏ�O6ȢT������a�33"�M�E�{X4*�Tܓ��-e�ɑ�S��a)���*J3�vyc*3l""ϓɠ�ǧ3D��}�j*��7OYԿ���'ʈz�����,�e �⃦�ƻ��M�k0�m�,�Kś'�Sy�Xq�����=kf���"��Q_`Z��0��mm�T֔ͩ�����呭�]s������R�e��&�=��[!�2����݋��:"Dss)��Q�dI�93k�>��l����)c}��a�?�La��a���tp��_�����45�(��o�*R��f����43��\k�3�vR�7���PZK3��)69@!���C^�2�Z��o���sW��,9��;�4ÁH�L�7�H3���N1Pd+>���&U/��C��2�� ����TD#E��b���bAI�Kz����ق�#ww'/qB+>
�t' &�����ml��垴'�5���̓k� ��/>���-�}��W��")�ƜD�^>��׵��w���+�rƑs������.LO�[}��פ�|�H��h���N��E����_$�Բ��C�r�����\�)󘻖Uq��h�1�d��Ӏ/K�4�:�o������Q#Z𰄉���'�{���JN��U�T�г4�����&����7Z��i��Ʒ��uwvU����˖j�-*i�@W�O<\�9��YS��:H�o牣�@v5�%2w�a�_�S	\�x��I�,d���jK��������m��-�bC�z��$�M'�Vk�W�����%m3�������Ta�Ywv5{�]N��
�9"_o���)�q��ğ/�a�oX0W����E� �� �:%�lv�%�ZC]bR{��ݳ�s�Ƚ��m[�9{��1��S'�0&�:�:��^m����ig���I���+�dX���G⫥xб29&�/gzN�����$�GS�%w������[�xF�3X���	���+:��f�q�cm��"�x"}?.�[!��N��{�0/��`�}�'��̀b�FF,� �&;;��f�0����+ޘ�]`Ϡ�t���6��B�|\�E5U�W���!���T���_?���h�������Gg��D5U��g�q��oe)^��^��oa��6�L˥Ji��e>��x�ust^W���K��	v���e�wY��Z��j�ߺ�A��7��y�v�q��d�c}�� �%%-�S���G�L7����֬驅(̣x���1�o='P�P�]dL�?�MD���yƑг��J��RrBҳq��[ �+2F�^#�<����	�]�&���}�a4�G:rHX��kX]��J{S�2�g����(�
$d�Z����q;�-iN@(����^n��W
lI^���ɧ��[ہS�����*0`C>K�L�<U�U��1J=�>��5֐�S6Wȋ���8: CV���k�I���A��ic6]�� X!m>A����w��YP�~�Bz$h��W1���-Qp��0&0"2�	^��?ƙ+!~9c뛣�Ő�1p~ԉ�CC�ӛ!���[�;S�]���� �4��U����#Oq��1U���W�@Xw�/'k���{�Jm�w9��Sql6��彥	m;9�H��ҰU��(�V��A�S�%n���f�G��aG�\<�o�s�'C?�	b�H��|�%%te_u���zƄ��}&ZU���L>������u+	5��7���J	���	��}���𾀾��mzʇ���/G�q���2�vLt:�j𥎾�*lu= ���̚zW�G�����e��&�����fMD�3`��\~[^����s�ݓ�K�9��-FR;�l�H�O����ѹ��~L��,�XD��8�)�A�/|#����6<�m�ˬ����R�%e%�8���45\���됁�8yE�s��khni�J*�Z�Y �o�����?��ܯ$�|��6��NS��<e���Z+�6��4�E���c/��������@b5[��a{<��Ye�~Q��sh+F/tm51��[ϻ_���zi�#P�y�)x��Ugl�Œ�=����Q�;2u�n8���;Jd	s6Gpվ���#亍}S�M1B�')-�XK�H��b�ڽ��	@���+_Ԯ�A5X�I�3P�-�?��q�s�8�P���
��jF���4mm�uK�h�����԰���+�ȸ	'�[��#�P��N:�NL{����h�7���W��!��(tcA��Ru\�7�n�G!�� S�Zڢ�d.�뗦�#:�a�8��0���`��:�.�Ǌ�4��Xΰ�/��� ��#W0����� O53���~MM��ś5�gΔ���7���J������ʱF��DW]���p�¿l?8���H{�n���j�2>��}�b�S �[��/g$s��
���\�D�1;��3�%F����~�?] ���KΛդ}ܑ$�y@�]�5�
BH nXD&Q]��~��\{ ����~��:1$�i�O��Ͽq�=>�4����y���F�u�v4��<j^���H�U$d�sH�v��v�+l tP����i
)�a��:�B�Vz�����A�W��� �-x�y�)B�e\�C�wǭ��OM����B��~��-t��K��烡g�<����c�cQ��A#�9�߼[��.x���W��S��;w#oW��Q�n���W``
ubO��`��%ԓ�9�Zs]V��AH#�&�[O]Y�����s��
��;+[,�GT�r3�<E~���[���>V����G���)l����|�8;�'{�I�y �NiB��>	��$.���+}��@��3�e�H��11��N@�H�W���C�ދNК$C��~��g�k>�CF�g���lj-����y]��>ՊMw�jh�u�JLٚ���ӣ)�÷�m�[�����| j����m�W�����9����r��k�jA�?Xb����]KQl �O�*�>�NQ 5�&���XSO^8��� x&��ګѴ�L�E_�,X/��T7����������l6���}��JΦ y^���`��Nӻ���D ��E���Ħ��*]��<'%�Rz�?���XEe{�Ճ�\�VF5�W0�b$,V৛��y�1qc���f偌"��QZ u�=ע��8�oشH�$�h���Bq��,E6]nD9��}�R[E �� =��[�c��,=K�x�,f�}Y�s��QzCI;�k^h	>}��Br)^��Ǽ�&�a���w��p��_�HQ�m5����Y<*��f�@'�c�3
k
ɔ����2aoܫ�RK��)Qҷ!v�C9��I�f҈a0j�!�C��W\��9�\̯ʲH�C7V�P���.쐯�(�� >�w�yg
G�C��#��k��ꏴ�k�# ����^��p���bǪ�֪�}��w�J�/��MF�����L ���~mx�b���a�ڈ���P�Ūqt�R���P}[�ꐲ��!5���j���P��H�����|���9���r2Oiq
8����k|7��C|o�DE`jO�w_�ҲRv���c�J�v�7:���ھU�h~edh���;t��O��������4�|�Z�"���|x'�߱����T��yЎ.��/	���}���s7v�^�$��H�u�k�ڕ��ѪV-Ű�@R�0<�?B�e?o������'6���tvp��2�)Za�e���Κ�3�.�dp�,߅k��dӗ�	%�)�Omp�ub�����M��2k����J��.�o�W���2a!�Y�Q{�A�NΉ�
��9�e�]5���:�q)>�?��<�o��[͚EZE�R��{Q:�� v�%ZC8	�{��Nr���`�l�p[��f9���1ӛSߏ&4�`���pY5t���gOhPI��ܦ�X���GQz�py-�Ὴ��ʷ	N)�7�b�P�S��q��$�� ���c3��u	q�+@0��K����KO��j�?�J!˧���0
��}����tM���u��&V�7��$�l	+]q�����3��B��]������9
S0�-��/R���_�i<����s����_}FU���U���l�o��µ�.������!ˀ��?�be�Q8x�t�v�V�$�I�a6��R�����jh�1�<�Q7i �4��ь�dTv���7Ϻ -��)���G��0����!օ�c�S���l��=�VP���L8����♹�ʑ��X�}��d6B�
�q�h @'���h֩y1<�i��z�����GV�}�x_>�r�	��e=]i�{.�:������(���$����j��qV�iɧҋ�L�^���I�

�՟�3��nSr&ʑ�2�~{���&U��3�L*'J�|�Y:5Q��S���J�  ��Mk�k�݀I�C&A	)c�i�6?�h�B�u!hL��iwb�Yk��vh��.Wl�=�-LI=ϋ`"��8^�9OAx+�+c&�ŬU��,n��'CFb!�V30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�!ڜ4z^��!�֚l�7�\|I�n3����1���D�#J��$q$�֮)軌���tc��G0�G�D#[h��вus�4HҪ��A�>��K0M<�U�"���!�抺��k�=*��r��w*D�˟�Ϋm��`I�X^Ү�B��?���;Jb���ѓLh���ܣb�){�6hFa��N�jr��o���v�yU�!>6-��1ױ���������vh���l�^*ɜ]w
J��W�`DVzRF_ ����$��9�wi��$�f���;l�{t�"W_���d<a�$�� h�9z����>l<���.���.�ݐ�1��C'Î�9A޻~k07���~R?����6��S�g�ظU�9� �.R�b��ؘ�e��$��U.�w r�E���=6�Z��z�C�[����Q��bj���|�^���q�66!ϱ�1�}E���+?�*�h��	B�)[�-��*>��)�l�::5��Wvp�Vh��V���,�W�Y;K��������5��p��Ϣ$�.ߐ6���!WM']���]��s~�x�`l=n� OF4� aG�����ܖ���z�����N�<N��8�?v�W����
��.k�V�,��:*�ìV|�'�v9%,[k)��2}������Y�qv��]�"HRt�����ҝܢ��R[��<���2\b�����4*��������%b���o�@�n2�w��0��lL*���U5�<c;�0�����Z��w�#W|��3Ʌ[y��Q��D���i1))��G�U���%�༷?ߵ�Q��ٖ�a#�����Yp+��Q,����|C��u��9�TL�8���a+��̰w%d}���<_(�Z_F�S8gs�]Q=���T)X�K��n�s��KU����.@�m4֎�ߤ��`#�+��;�������VCS;��������߱*��(e1im�p��S���z�̮��ֳ��'~o��]�PF��:�┹%�\��}�;`�
< ���ݔ�עF0?)+<�IX�?w.ȳ�8�A/�i�0U�FX��d��gHm�{J�gK��v/�M{�2bk�LB��a�}ԨmR��2���?e�>s��G����R��"Q_��m���F�T�Idu���G��Lw���.ص�g!��.��T�Q6��������3㯮�o����!�xfB����?)r����m�څu�S�Q�����?k�xIР@��]�A�+����Mp����������-��4�[J��4j�b��C��տH ���!�̛��鈯�H|0��b������$t3��i%�%ͨݿ�ʯ�P�m5L�	�@�0���J�j��Aa���NbԨ-59��5w��� ��\G[
�ڻz�cr�Td�c��N��̈6(���G3��pעi�Z�c�&��2\:��Lt��B=zx~<�p巾����ja˗Y�r�b���=��-H ��O��jIP��N���:��/�;����|{ZD�$��El�t �R'i��ר�H�"�W%m$gG=�N�޶��v�`��~�ػ�`K?�.T6W^�ÙO�B8��{$=���~�Wc=]D�E+��]h��N��yAp˴٣PQm�=�� ͨ�w���N��D�[���j�(��t�2F5d�:���jBj@w��v��
It =�2�%ꗿA'D���<v��dĭ�CY�+����J�Vq�Z
Y��+"���~�1S���C��1�9�:GY%�Y�G��	��+��a�$�3���4~-��]T�=E�2����@6'���j�3>~��]>�2@�D�NM��N���@ևe��z��ϟ1H�����{�^ ��WҬ;Eߢײ�d���;��h����!��W����4bK������������۩9j��xb��A˓�\�����M��eM�N5����:��
�,�L����j�����Y�NA;3nȓ`���c����I%x���* �́�����!�-u�.���]B�S���˔�:�T�.�=����u�<�:�4�G��Fy9�Oݎ��iǨ�+�g` ��2��Q`M\Ð�}�OZ?6T������շ)?�����\�`��[�q���v���z}�+5)�n�1��班zMa�8�W5V��OH�.�J�]�d�|�oU�C���)�h�L]tU9-�ʨ�G�&N��'5h'��:��h�j`��KP��ri����a����5���u8�� j�Bk����|N:�X��B�O�}�I�Sۯ�͢�	�"�HhS����R!�d�i ��Vi��5���|�N�0�Ko���Hc70)��k�<l`�X�0_aD0���Og��x����2k�ӵ�*�h��WD|�(EEmk���5�x"lȝtM�
d"^iKC����v�P�YE�϶
��i�r�5Cp��Vŋ�C�/7�,%�C됃&($,2SMZr�X�$d��qD�#�8}��J����,<���ĉ���菝x��ǉ3����|>3)��u�J6	6�:V��wz���@�k���H�W��2��3� ��4?��=QXyZq% �b�j�2�X]�:���R�rm� с�:����� ��@r�K:��I~V���a*nu�;:/��<L����8oQ��|U��k��W�j�����y�a�g�"�����+?9��&|>�g�?�UO�beaF2=���3&�R�2;�jh<N$~�.%n�(+ fPV�1�HK�2��;�y9�7a��5HLc��N2V�k�H�`=m�����u�9(��j^���(��k�P"��ǒG�*�����}p�C��X���ʴ~��S�͘�`��ct���w���ЧA[h�)S�ɔ�����:G�����%+můV�Α�[���h~l��q��~����,����VB'�;�l�h�$�Ɨ��Ҷ�Q�&-(fU���(۴��}}�M��� ���9t�B�!�>0�
N^��,}H��B[@�OrBNo�W����.v
VegomL�6����d����ЇW�Y�\��P�I4�I?31�Nq�ꃣdbx?	��&�N>�Փ�f�I�d�31�v*��g8��6��8�K����'����҆�p��ٍ��oQ 媐��]�H��;��b�~&��a k�=(s�)O�	��r�GuS��&�&%��E·�&Ѷ#�k���@p�er�H���P�y�0#Q��O���+ ��k���2��P�V�_X�Z5�Y��^�q6�a^`([=�6&UI͇��~��c��\1	kT���G�s�1jtq��&����t8^��W��1�D!D5�s�T��N��6d���`M��S��рO( �B��q�0��dn{���MSP��IQJHI
'��)�Ne�<G1?ۋR�-j��%4o��U8'\��,�i.y�����9qm�n��eJ4���*X�ჟ����Њ���Ap|�F�}�Cd0R$�������
��s�>�;;��w���߉���2�`�9�-��줩O�}����-�I�z,���!H�B�r�#�"(� �Wz�M�ŐĆ�}̏�_2���BX\��cD�T4���$����|���e�6���Z� K�Qi�X*x�x̥A��W.����(���W��i����B�;��ߺp�JC�g{D�����3����5K'�'PPC��<
�C�Ȓ�D���2T�)���^�]P>3,u�����A��I�;�]���$b���P�܅��]�9��x[\���^t\���9��[����s%��������'�I<F��+�@��M3��e�`�}�c\(�4�u-ʱ^6���U�Ѷ�&��r��"-�n�����^3��C��vpF��z�U�|�Y�Yt�%+0�����e�X�{�K@����ݗ9cJ�>�O��Z��yJ�Wd��VU�&_;����;���w�'R$�F]���{lm6Ѝ�`�_���d�Mα/^�{�95���� Ul�� ��*�M�+4s��߯'9�9��f~��9��5�Y�h�#Uk���l�·��s���Ty /ʫ��l-ǂ��8�e�t|$n܀�m�r.�� �ӗE����x���j�z���[G��/����[\�9�SǬ�H(0�zJ�eߜ���L+�sC�L���ё�!���]#�s��X<8w�f4b9���~a%y\��fG��E���.�͏�׈��G��蚰sa����C{�Ñ|���.
�QS�@�O_�3����9)z�{{��# �a�ͦ���NvU�Q�@��l2� �kr��y�F�ũ��d?�U���b�'��&�r�/�ꓰ6��%7xG�xw��,��:<��Q]��/�-�4TH��6yn�lt�	@(��#�<����0�����x���������	ׄ.N�|�ۀ:�Z_��e��s���[�{S,?����YU���&�n]��Y�Ah�*j5"�u������u��5�[
ݲ��4ᱤJJ)au+5�)�����n<��ώR�C�����>Jq/:��zx\��M� _��[e�Ųm9�$����\��ip(<�q���2~�ˤ]oIH6�Ǯ����_g�ql+���pC�U�~2�K��CL������÷����/�~XEu���zCKKL�з2���l\'�x%Nq_f��UX�m@})�F���I�x���ՓuҔ%A�Z�h�����+�����j�����,5��7���V�c���*�-�؃��i*� pQ96�/s�
9��H��u��c����}�VbfpM��_X��q����?���*k�ĳ-6�d+f�K�NOx�I��O^�,Y�a��ѳ��88FJi�S��:�#b�wP����a���R����.��@H�%����ȆR�EX_�&'^+΁gҹ��Q�X�&^P�,��L�5�Rt*�}�[�@g�9�l��f� u���kA�ǿ��t�~����S�峝��kz_/�$WA�4g��.F/Ғ����"{N}���R��������(gF(�r��� ~�O�D�:m4�P,(���h6�6j`[(���M�G��c	�����cF��+����������?�`�s�JP�w����^�fd4���3����9��W	��p��ԍvu!�n�`����/Gj-5����r�$n́MR$16��+��̮��׳�d.'{^!���!��Nz'�!6K�.��H��g�f�Ka1�瘃�R���o$K�І%]�����E�y8*���i"�`d�kQf���֤�]ɶ�"���/X�.��b7�0������`O�t�$���*O�D�Z�e��7j^�<����ť��L�4~K{V��D����Heh�����b����?�d(U��Y��ݶ��u$�2*+5w͈���hT��j�"K�����0� �̯�(�{����8w�Njw�Q�g-~|� 
���q��匸�BAt����	��SH��A��LRp��ē�gi!RVXi\5�h_+�"q
���Ϭ�$?cf���-�k��l�A>�1��h0
wMO�,rx��~Skɶ���콽��A|q��E�-�GFmxQ�A���j
S��i��Ңl?��]5E�
����>5�_���%Ď��7P�䲫�u�,a��Mi����$3+�q��Ǌ\��	ĺ��M,k�-���ᾩ���G�o�v�7�)L<�H�>���%�/JE��)�I�F���:��k�����r����b�M�����XH�%��D��O�q�����g] �r\!�PǷ:�׆P)j�l��ru,<�~e��P�D�:�ݟ��vL��wÔ�����"�����9?u��L���aF!�"�������9�T&k�6�Q�1&cORI�a���d��3U���a��;��$<z���4�Ӟ-� �K��!Hz�2�D�;|P���̍:�*L���w�V<�KH�n�m짛����9�&����0 �Z}gڟ�O��_�93H��$p�3Ţ9%�q)t��}�S
%��7�r�L������A
5���N����_/��i�k��<֎��cm��XV]K�꡶�ZV��~y��{o��ԣ��D�c��V�;,�hb־�w���Q�l�}�3(5D��5�ٴZ�}�!�^�]�O;@�H@B�q�~J
�ep뀂�}�IaB�݂ON��N~��W�;��ڠ
��o���3�L��__dυ!���ZW���\����Ϋ��z�11���9�d�=P	�LP�= �bG���YV��)1p+�vy����@jv��p��t����P�_~)�������﯃��
�]���3Ԡ�р�&���/m4=p����	��rP��SAP���6�$	���2�ſ��S@?��r@@��Q�U��u�#_U�~��:�W���w���l���PiL���BZ�V��(�AqE�m^O��=���&���k�$��	�ޫ��k��!�V��sow��쾸�t��(Xn��6s7E��`'���00S��aؼ����۸d�&J-�en>N`%�f�Ԏ0���QE\��*r�dͻ-�`�9pw�ӝ+��,5ꐈ����⻳=�#�<c\k<�^�5��&�r'.-YK����N�� �){�wWG�\�*�O5E���an6On��@��f~&�C���}26���7�����nbZ�S�x�y�>����>,oi�]�`�*@{�w?&<̆�6��9���ɔ�$Y����Z:����"�>�Eo��ΌZ�g���f�o�P+�F��">@����4l�Ӿ|�@n�F�>o38At��`��6: ���I���
���|.؁!;���"����a��7��I���k
�9~���#Qx^$X�5�uA�3ͽ��=J�f0ƾ�n�r#b������u:��4�����>�0�6aUf��#PS!)3��onk��D�[�������������g�XErm�	2G�=�%�W��;����z%s��쾫܊�)BQah�M��1rn�/�UnT���v"�U�7�>�X֟�թ����-�H����@���1��t>��9#$oPmo��8��F+9S{���\WHT;ݥl��Lbe�����˘sSt���*}"���F;��=z�UU�e)w@*Y�G7�
6�:?��y��C��D1�W�j�����L��dmn?��D��r�e��}��s`�ڸ�PL��TE�3�����x ���^`GV��Y�j+g��r��4*�����B&�q����� %dϡ�E��qxxVE��%{V�K��Ʉ �uI%&�p�FH�~��Z�I�;��^�f�e�C��������Z�j(���Z������l2?�����\#�V�������X���8~Rh���HBs5j��Z�Y�`F�)%Ĺ���o�y����Y�S����k@[=�#\˖�P�(�T.> O�?�݃h���	l�[�^��52��?l�ė5�fvc?h�=W��J7���Y�6��2Σ&�5�e����>�@��|X�������-'�6���-�s(�	rF=�q�B��}a���%���	ժ��~l�~��{U�� ˍ�	�vol�@W��t�(.�7�K�:T�����Ѳ�v#��[�eш�>ħ����C��q�$y��/�HÅ��d������F.���S�бJ����Ub)������*o�c7$ߝ1"�bh��oИ
nD��w����u*��W�H<�%�ڳ��qU���`�w2�!|�KW�o��YQ��O8�P�S�)�$���p9��ʍ*?	��QJ�D����#����M�+`\,H��f^��E���Y���v~8�|#�Dy�+�6�!��}�_�<�*��FO<8Q=�]{D��B�E){���s�*@��pʢm��WH\ָ'[�E�`�Cg��4{��#ڤB��C�����):����䚶1S��p���H�gzBc�~��:~��V]o�F���A빏x���q�%Rs
=kS����.y~Fy+f6�X�)�w�.|�"0�AY�據3��c�N�����4m����`���w��2̳����_�ۧ��m��2MG?O��>�k�G���k����>_�(�����T�c�u�8kGu��L!Ѯ��O��d�!'��f�Tr�0���?����ݶ3�Ѹ��/�!E��f�����r�|��B>���c��=Kד���$5��"�=��ɩ���Ҁ.rMZޢ
~tՆe�Ds/�RI-�l�Ů���[�b��`C��)�ךgtʧ�'ߦ��9�awN0z�%b�F	�*t}�@�*Ǽ����a߯>��;�j��@&N�S�J�5��a�a��IN̖N-�D�}Vw��j ξ0[�n��!)c܄#dK}�ѝW���C(2z�Gݔp�V�ҋac-}�����աt�&=|��~�:pϵ����T/��auŻ�\�
��Bf=Z������]&�:Ș����$$/��B�{A�$χuE��.x(6~��i�J,��r+� �o�,v$Q#g�x�C��_��
2�~���ߊ)�����6o$ÃuxBb����lŕf�~ԭ cg���������8
}y6�&��'P������J�ť��S����.~���
j�$�{�720�	�L�Tj��w���v�K�t� �:�2���G�DxkV�殙������Nd!��T}E�@N���Yi��飌h�L1}D�������#VG�?"Y�����B+��e�N��3_�Zg�����0��߇%NBĬ���^�t���'q��"�R�}б�V]����q��[%MR�-�_6�^h�-g����~��uV*�m,����2=�t�	����>g�	>lT���=���Z�]A�=��Y�t� l�p���8�0��Έ�-/�0�AD�׆���p���|��s��j���	��Cf��%�(!���(��[#���|mQr�,����	6g�L(gMMOW���g`�.�'cf���ĺ��P�]G,�|+�PbPM$��%��#$[��΅3�����<��_��Mɜ�
P.!�w�`KD���Aj*ψܐ+΁���n�v�M�*v6���]fO�)�g�a+U{�����QN�+��~T�6h[�r%H��g�g��J1���]0h�Ռ�˔���]{r	��@�oo��U"��с��}�3�˓�]&��"���/�5�.�_7b/��X��oO�ad�����' DV+Ze�7G��<1p���7ȫ�`#��D�D��m��#���b�ݞ6�Ϡ������VdP4�J��b������t��+�^��,(�N��ϊ���}��~��M�$p��=8d�����Š����%�5v��I�W�B鮾RǺ3�p��3�ߊ��ח�y����6��r� :,�R�*����CdwQ��T��E&���🰬;�ǟ����0|v�y=l�:�Pl���!Q�xV>.��\���g^��yD�Q��,�K
�2ʹ�S.!�TۣY_���B����B7�a`��4���So���\o��S��d.��-6�!nޏ_`�}�t��`�Q�mf��P
��\-�!��Q=�s���Y�����X?Ժ����.t��0�k� <�b�5*k���~Y�~I��0��n��ɜ!��������r*�J��n�t�φl��yt	&�`0�9�2�9̻ך)��Ren ;SS}��NM���l����i�Z� %@"�ߋ>�&܅�;�֐��ĴU�`�Z�`����">D��(����Zt��g[��f.�4o6���1�"��ڇ��/4����^+|t�a���oӕ�tD���.|/ m֔IH�
4p�|���!��!���w���7P+I������3�b��#�M$�0���)��[����80f)��S#7��It�u�#s4�sM���>��04,�U�!��-	!����!5k56a��s��~Pϲ�*�r1����X壦�������q��Ku;Q��䳯��׌ܨ�*˼)�Vh��u�rk ��CY��zv�<�Uw��>����'/5�4���NЃ�N�_  �z2�����>�+�#��	P��o��x�]\g9�D[�sZ����E���g�e���Ei#�	����5*���(���t�����de��!*��V7z`�6'Dz?I��S5���V�W�����L���[Lc�m�*?���D�x�����d��X-�L�O��9���Ӌܽ��㦨W5����T)^ IL�g��j�P��s�����=���(�$�>���׮]� �9��G���T/&x�v�E!|9����됏H� c��%ƴ̒�s)���Z8�\;&�������슟����Kz����(2�%Z�����2l�K�{"��Hջ�R�O.֬GU���$�8��� 6�BW�����Y. ;FULe%d��$>�o�_ ���7Ƣ)SW�ҧ�[��\k(�����T �̯?9?h�L�	=�[�U��tg�l|Xlh��5��ov�drh"s�r41��Y��P�k8C�Ƣ�5�r2�=&yYd�s\���6�«}�''�f�g��s��K��=8��Yy@~Ha�W��O�7	�=�8u��E�F�����vRd������ .�c	�� �:���ö��q�v�	�[5�e�<�ߧ3K��4�q@.��gm"Hcwh(�=Ԑ�d��;�ޜ��Q@����mbɿ��[�v*_ם���qb'�op.�n��Jw�{�>��*7%Ώ)�<ms��z����'�$J!w�v|$/���o�kQ����`����/)g�&�������j3�?��Q�)�7�O#�q��vR+ sw,�/n��_��L����Xu8�����B�+�%��F�}SE�<)���o|F�8��]�L�◨)�h1�"�4sWd�_f)�B�N�����X10߮�`m5��2Zw���Z��ԀC�E��l߻s��:H|1�u�p����F�z�x�J����.~yv�]�F6�ҧ�%+�/Y��)��Ň�
�TG����JF��+�X'�wx�`��QA�z�:���u���M��1�m����Ϡ +���X2l<�X4�����G�)m\և2��z?��>=57G ���|���@_`�P�,�/M2T`RuM��Gc}L�""�F�,��6!����\��T��_ʑ�<��}�.�q���	!�
f�KY�t�Hry&����$���L�������]���Z.h�}Vv�K�l�Σ�M�C�����&���t��s-��ܚe�A�~-�b��C�ӕ�ɿ{��V�4��|J�5p02by�ǨئtH2l����݉�/��sL��L�

@�ډ�;�JG��Iw2a��yNl�w-\���w�HZ�
���^��[�$�څ��c|"�d���q#�����(��rG}�Epa��r�0cͺn�|q>�u��t���=�~���po�5�`v��haW���_ܫx�p=�³�t$.-yV�S����ĉ�/aX��1"{�B�$o�|E6�F�fi=P�P,5�ܰ����$����tѶ�ƕ���~8?��*��_�6��Z�#�vB$�˅���!x�~t�c���O�U��d����y�w�˾�mP�~#axY��X�����昉���38��
7j����0%2�Y���ԥ�~�j��fwu2v�U -� �,2�4 ��!Dy��pn����R�o�y�������ad�Y��lKp�0�1�Cx{�hP`�Ã@G#YYY����S�+#�I���3��"4Ȑ��� ��皻�<�B�@�(�᪝I3 ʨ�)k�����D��W-Ng�@��1eiRb���r1�XA��B{i���j�����,�,�.'8�E3h��������!v���Kٕ�=w\߻��ڮ��:�d9���x�g<�K����0��ꙑ�:� DVe���N�U���j��3*v�h���MKot��~؜޸�N�K338"�`���LWg�g(I�=��� (����V���u�+��������;Ӕgz�B7f^p� ����H�Ud��'�,[&�6/�߰D���4YGs0x�7eD���F<j�]��$/9��4b���e��ف	�?��1�<�ˠ����F�˭�޽���O�l�R	%
�Nɫ4�NK�Z�������y��k#V��\q^��i�8�����ѷ��:�g)�	�|�H���R�\��>k9i0_V�Y5�f�V_O��C�����Z\c!���k[27l��%2�y�0�_�O3�xf�{C�k4��� k��_�|�+�E��r��g�x�Э��M`
�%0i屪��׳j�E��.
&HCst�x��d��-�c97�#^����Mw,,7Mt
%��$�/$qVp�R������E�,�����¾�1a��y]�
�j��>�B��JP�qӔA���V�ej\k☢��[F��8������U�X�%�3䄃1�\8���C������r�
��8�:�a]���W�|rPS��~p/釻C��:	���3L���p�k����;���*&������&�?va1X"@���]��9C&�ˤ��\�O�)�a��:��͎3 �.�l�y;>��<�V���|�)i
 ��&!JH%ld�M�;�zo��4W�e�L}v�bl�V�U�H�})m��Q�@1I9�-�Da���E�������D���a/p��#�d���u5��[�SU�k�:<�} ��9���z�A5�ǀC|-��*���� �i������m_�7V�v�u���E��Pk��v����W$Z�.�V	�;��-hM备`c����yQ%���( ^��`DH���}�gq������+��S�B*9���2
(�h���}�ΥB��WO�$N��XW��A؛*�
0�4o4��%�G��dzl���X�W��A\a�v���cD�1���7�d<��	������x�-���#��~�1[��v�i�Ȁ����7��k��$	��&�J��
��t.�	fZ�ݐ�Ɖ]�����弬�&<� �?`= �`���9	_��r{��S̅"�o���o�m��5�=�l�/0�@
�Irkk���5����#���)���E����&ķd�"�P�7\��\�Z�P�����qPy^���=l��&/�,��+ʙ�!;����k.@U�assڌ�t�F&��B���8�r*W%����!^�s;j���ŧ
,�4#M�_�>�c�)Y1닉=����~b&e1�����+Q���ϳ}���<Z� ĨF��8e4)]H�V)��Ȓ�~�sK�+����6&c�k��LU��"%g`a&T��i�{���V��C�����ȿuD��/J�.�1g�Zp��'�\7�z����_���V~��]sF��W�Ջ_��}|���9�\
єe�-U��W�F.�+�		X�o�wl7t�6K�A���c��6��b-�%��m�I����t�S���2ෘ�L�%����;LmЖ�2��E?c��>1��G������=�'_T��<t«#ІT��6uA�G�q L��&����s��!*���P�MT� 1�S�M�.��q9��(~�B!Y�f�6��,�rm�E�V���:ʮQ�<�����8s߶�9ΫE�q���G���Mn[Z��՚we���9�-x� �٪��rڌbO�C����=�������&��y�uGq0��b�k ǜF&t�@�&'Ӽ#2�}�ܯR����a�~�@�A�g�0J;�L���ax�N�-P�n��w���~h��RՓ[���y;�c�Мd�K?�>T��x�(F�)Gq��p�a]f�cA�|�p����t�Ȼ=��
~zNsp��T�CKa	<1�p�.�l�=���K�J�Js�̘��T�8A/U���V��{�5�$��E*HF��:��i�;ȨD�E�u̲�tc$e~������ ����~�^����,-6��×��B�����4�-�~�Fdc�����[��sJ�Loy�Y�2�P����B�������L+�BU���Z�j���M2D��0�h�^j�14w釀v~Y��� {��2�#�}�.D���z��1w�F�e50G��%�T7�U��Y2�`*�|��1���b��\���7��G�.Y�-�Gy�+��Z��)3s�54�}��[�3�۔���V�6[@4N��q�3�]���0��D�Pmˋ�Nb�@�e]ښ�eL�1������{]r &5:��6yߠ:f�"c����h����W��F�1^�K��@��86ӫ�N���.��9hP�x�1����i��G���X��Og��fe�zN3呯����o�j�œ�C?�/�\������N?I3,Tc` �@։��ĚI���e�� �F������u��/
�Q�{͉��:�@�l��;�|�}UuS|5:�c�G�PF70�O[]bЧe����g&yGd���[\�ů}�ڰOث�T���&\���V)��Dl\�k�jH2�|A�)�涞�X�)t/n�z�� �z��Y�Y큶���^E��b�纒S"��wl��&��s�U70�F���=fdS67,5&t��H���Yj^�kKd���\��X�_���`�l�<8���j�\ϖR�|�˱�a�@xZ�;ݱ�����0	�ZH&���*�R_8%�b��i���V�B�58t�z!A��m���N��N"c5U2�G��k�"lOL�VM U"03O��x��}�_@kX�w�h�i���n|���E�t׆6o�x �ǝ2ι
⺹i��f���>sE�v
ʳ�gSJ��
�P3��˥�A��7����0׃d3,0�lMS;-�$�1�qB�s���Z�.���K\,:@т�1�8[,���-�œ��Xi����>q�#��NeJ��Ӹf�Ե�p��h�k�֔������A&�1�āPb�y��X�ؤ%��(�>����x"5���[�r���ѿɠ:�'����{jyr���H~l�����p:-;����<L'ߢ�v�t���ݵdܟ��ƌ�?��[�7�jaU��"�F�����9�G{&�d���l��O��a�g�S��3$�s�'[;b/�<�xd�,�̓� �#��t�HI4��T|;�*�u�~��/L!����V+�H�)Zm����dvU9fz�h*��_� i�Fڎ!��y$��)�@�0pA/J������%��v�S�*��^�c!��]�P��_AYg��&��*�N��8jɡ[�+ �m��V�@^��.�i�0��:�òS��?�{��҅YV@��;N�dhq�ʇ���.Q�,��=J(�;���֗��{}��Mϸ�0�����BN��|t%
L*����}�]B�s�O�N-��WQt�?�
TOoؖ�B�'��t�d�8u�M�$WJ�\ꆩQ*�G�1@N	�(s;d`O�	p�w���0��:��G��"�]19vh	U�\���˽eM�b��*z�>��nzﮰ1��=���~���B�]�b݊�௼&�[���=�xӪ��	��r��Sp�哝k��׷�u���x�S	O@��8r�v׀,2���=#Np�MI��,r�@A��[�C0��P��O��Zs�!���q�^�jv=��&S#Ç��/��Xޚ�gkR,$��s��t���&��2�ϊ8��W��}�/Y!܆s_Ӎ�P�@��L����M66��YրMͥ gq�q��|�b�K�M�6`�m_T��'S?��2�:��?������ ��4m��U�C�'�9i,"҈y�<i������-��4��}��v1�_z&���k���`���F=3U�A��R�o�g�=�E
���fsoj8����S������Ƹ,۰H�`ϻ�-\��b���E��TbM�$%��z�~��_(NB�Z�#A
�~��zXV��GL��K�&΃��BVb�!
�T�t�b�����ѽr����U�X���~� 	,�ih�*X�Ȝv�AM�.Q����(��;W�ji_�׮O+�;����.yCA�oDLn��5\ۯP��'N�PNr)��`Cr��Ƚ�\��x�T�g�1J^7¢P<�&u����S��A6<�9���Q������"������(��x�Ά��������[G5�O�%_�F�\�G���5I:��鹔�U��$N^:>�!����m�uk�^,Y����4���:�p�8"��ū��[��o�^1�C`"NpĔ؏�a�_WY��K����0�7��B��#w�ց`Ɖy�����UZ�Jmˉ�|9M�0�ѩU�)[6J]�Wb�V��_�����LG�\\w�U�$-,��7�Llks���=*_Fl�dRC��s�9�`9��U���l���f�����g�i������'�"�9z�!~�Y�`?�K�DԠ�����ef��+��a��(
 -a%����E�A��Vte�Z�$,�����.L3 눿 Ӯ\�P.i��Kp'�Z\�
�t����N�kk��T�r�5\"!��p��Y�7�����+��{�	���.���a�����)n��2ϸU���1&k^Z�+Rl2ll�Iмc��n�|aS�x����~�au���G�i̞�r�@�:Ѻ��X鐕�:��B�ȶ�� WZL9��=7"0E7H(��\Z&a�gM�_f`
�o�|�nZ"иӇ�/C4$Qo�J�|f���\moEVDt�{�� !} ��I�sP
�Gg|��{!Ӑ���#�Z���	e7Q�I�������Ӥ��!�#cz/$�#'�7�n�U��%0X���@�n#t�o���eu�>�4����"��>elZ0&p�U��9�56:!T���"�kg���me7�0pϤ�pΤ��y�X�L5��V
��M�i��;Q�䥗,E���������)�� h������r������ ��9v4;"U)v�>�a��Y�8��r��$Ƀ�ڳ�
����`=�>�`�#�ΌP��oF+��O�x9%a���������7����ˠee���b��9}���*��y��&�f���'��e;�W*�fH7lb6Y��?�5��J���W����y�e�.LU��m�i;?(�D3P��+�O���[�
��L���kT�Ev��g_�����,(�^��8�Yj�Ɔ���5����~�V;����#�`1 ��O�yWH�ƽ~x��NEo��%S�]��pW Uq%�N��XT��гZZ*T�;X6z�xx쒕�s�����}& �l�(�GZ�ZS���lD(^8��tҏ��}������g����8Pw���/B�r,��B�Y`�F�"K%P%y�o��\�!�'�T�SI�����d[O��\_!�x�&S� a�X?�~�h��	>1)[�z�&0ͭ^[9l���5#5vl6�h{%��:����:Y7<�]�ģ�qj5&(���aK�X���4T�2#� s'Yq�����sz�mh=j�W��{0��a����S���������ā\��಍4̄vy�����/6.g}���PJ:&:
�(�'�#�$v��[g�}���������VRqr����ӂH��UQ����X��NS;�C4����b;x��T^*��	��Cq�b���ob��nUmw���>�*)�-�Qv�<�f��,Є#��V��wDb�|�b�)i�Q��]�T%��\�)�V_P��'��\Fk?�n�Q\����IF#x�բ�0+rs�,�>����g�Q�k�7Pp�8��k��+i�s�}E��<[Y��TF�g�8��j]M���T<5)T�R�,|s�
��v���M��O�֊!�� yg`�^�$�i�����T�uCO��r���n�-�0��@1�p���ZxUz���<jԑ�Z~�b]�F(�0�I��ܔ���(���
{��+����BF���+8ߜX���w*TR���rA+Sۓ�/qB�����E�c�ym4��c�����I2�2ޡ��
����C�y��m�O�2���?᠌>o��G��>Ƚ�#���_�҆:K'�ᆆTR�-u�G���Ls��8�Bر�!(���T�TM��J��,�f�/���c�*�R�!W!Bf>�~�f�r����T�{�����͉����6���t�HL?���)��ǔ��&M�ү� ՘�����r@-��B��H^�08�b�dC�Ro�;%���)"�H�-��DT�s�0��bk���i�t��P�༡t�ݻeϯP��i{���@��_�eE.J�N��;�a���N��-��� w�� �|/l�|�[�$ ڷ�zc��d�!�c���ȵ�(D��G/�pS~f��>c?�>�.V�gBt�c�=��~8�paO����OA�a�͘�����=�D� ������rJ(ʶ�i/���T�@{VT�$a�Eh�R�� �i/AѨ�;o��,�Sq�$���J���{C�\�(~*�\�A���6S����qB4�"��zJ��6�~f�c9��_"�Y,����?y�C�0��PMϣS����ե�_�J�X��à�ޘ�j۪��|2��Go�f��j>��wg�.v��v��+ 9��2r?����nD��8�<��۰����3r���<�����ߘY0��[��5i1OR���X����2�GU��Y(1��N+�� f3qP4z���١��:����c��M@����܅$3����'���I�D�S����N�,"@�=�e�L��c#1D����{�ӣ$�IҨ�y��{�`3q��mh��.���5�STެ/oK���/�K���L����Yx9�IxO���W��X���+��ۙ��z�eI��N��j��c���R)(L��L�}�Q�Z^��O'N��<3j-�`����	�"I!���c� ����y!��%	u���-���\���S_:��*+�������uQ��:�@�GFw�Fu4�OY���eq�9fg\!Ek
�M��\?�X}=|O�U/T�m�iH&�*e)�����\y��c�D���H��1��u)r�Xn��i�cOnzI��?F��m�*l�����x�����������K�H��U��Ʊ���I"�s�5dN �FA��>Nj�4�KL-{��M��h��ݨ!���̷j�58��jD�f��y1|��&�xľ>O�ys?��YY���|	]0�Hd}�(C�R����i�x�V�c5�oQ��Uސ��#Nּ�
c�W0�"�k}��l&'�^7[�0�TOc_[xr��TkV��&�*�`�F|ޙ�E��X��Հx�ǝpܠ
���iG�J�o�p�L;�E�&
����/�� C�Dy�R?�ҿ�7����҃"@�,�jeMV9?�$`��q��4������L.,�X#��̆�6�&�t�m�C��疀���
X>/�Q�rOJ2��Ӷ�,�s�ˆ.lk�K����������C�����wXuXu�%|y��f}\�~P��6��-����r��}�+:s)t���y�cr���\�,~R8�ݼq�:��1��eL%V��4��������ه�@�f�Mٓ��u�aS�["�{֔�f�9���&�H�c<0���O�+�a���� 3�� �N�;`1(<J�6�z9�-a ��L�eaH�<d�2�;	���3�]�G�L_�=���V��QH-иm�2��b��9$d��߼��9ag��L�(�C��&[��>�7p�
=��	�>����S����ܒ�_K�[.���VYA�XJ�%H�sJ�2����򡙞H�)�"m�q�V*�/�W22�g��d��A�<��L�y�����ZV���;�ٚho1���3��NҔQy7�
R(b�����Ƕ�}����������5;�BLȷ�:�&
ʓ���i}��BWTaO�RNk�Wa����
�V�o�O@w��3ld�ȅ��Wxx\�����@�E��1>K_��Qdރ�	�\g��Տ�����`4�1}7Cv&��Q/����T��G�Ax�|�q�lGv�l	�F],��b�|7�� ��]n*��L����&�?|��=W3��]d	��er��S��������b"��C��Q��@l��r�_׾WS��u�#	���P��'ǒ�>#����7P���ۼHZ1�h�uҪq2~�^�js=ΚV&� �������Xa�kв��C��s�/�tm�Y&5����8��iW����}A!@�ys]��X��I����]hM4AJ��Ě����>&�o�q�v���s9��LpM�_���I��FD�'�̨J�nڸk?�|��>����4뷨U4�'���,�'�yAJs��fR�gu���*4}v��&�u�].�|�k�LĻ���<�y�F��ӿ�R HC�er��َ�(s��"��E�Kk�Ӫ��ۮ8�`���-�C�젊f����芚��H.z������B�Y#?��|��zӾ�A\_�ظ��$����uBԅT�_��T�oW� :��z��������7O�D@� G�if�*֙�� A�k�.O�AD�7��W_�i]���B�;��l��C?6�D
[\�k3���q�w'��P����85�CpS��{�PfT�r�/�B^���P��u_��QfgA�ʪ�����]��y�ජ�X���ܸ,����xW��_�BXY�����[��Uz��%����Z�����[I����'� �S����x�>��_wv���u)��^�?�ᎋ�2�(��=��]�")𵫈J���^��~C�Ip/�v*�����Y��0���y0�P��{�¼a���Ԩ��G ��Y��ݓJkA��:Cv���G��'��J8W�k�VQ�A_�lO��`E[�w�P�$+����H�l鍩����_D�d�C �����wL!9�!���Il3���f���a��'fI�^QL'��9x��~���.�f�Uq�B��gg��b�0���B��R[�P�; �U���g�Cݭ���ae^d$j�e����.
C\ iE�����N�P�zN��[ ���$����T���r�5c*�(�LH$R�z��ߘ#����+�3����7�ŀ9ǝ��Y�/���X8�~Ҭb5O���jyXپf�*`E�W�.�p��ಡ-p:��Ҁs�Ua���{k�|�t�.���OQ�@���_��S�B��)vF{T�� �s��"r���*Uo�Z�<���� ���0�{	yή�A�^�`�=U��(�NA'?Q1&�M�/
%Ѱ2#�� �G�q��e�:��5<H]R/g$�4P������h��	�����<2�V�|o �t���t��E=2��B�	S�N����ٚZ��k�Կ䃱YD{O�Ǩ�)��U1$�I���j(��լ�h��5�]���哽d��������!�ٹ��W��Z�J���+1�o�тj�����N�[���s8J�`r��۶\+uX���ܤ��PŮ�w�����������(	�qi �2z�Ĥ�P�Iɣ6�����`W�_c��q�#�����C����z)|K�L��������H�(/�¯X�8~�έMK��.г���+\#�%��lf�wX7�k}%���0<�I��#�x�l�q_%���d���]���l��#(���4����� ��`?5c��R"�-˿��I0����Q��p�4�ن�ԚD�x������'o*}�(�f�^��[����;����e*g8}��k��`9Pf�܂K���xfv�������a�v��(¡8Bd�����C����{J٪���]�/�. l��?+�]:�k=\��G�� �����xX��
�as3bx<�ԝBy[�f&�BEY�.����ED�D��'#�s�����R�{���|�.�.�u�҇L@p��_ފ���6)y {�L, �@��E|<�e�AUR,S���������Q�yڭ5�d������Uul�#X�'₹&��_/mK,�����K�Gd!.�Ht����<<�1�]�[/���4��ռ���+N	����b ,<գ��{H���7!V�hn��]�	6N�ޠ۟�ZMU�g��F��<��{��}b%ǘ�G���m���8��hX�5�t��MᠽG1��!��zdܾނ��|�p��J�`�+�֊�R$��.�����Qs�����~��˷Ԫ�����3���ZM`��Lȹ��H�������qcp���i��a�M�	�h�Wƙ��'/�&��m�䣽?�}j�FT���� 4	�U���'�,���ymQ���S�����4�3���Ɖ�|�(���x7W�l�F$hBF�ɇ��$GR̖�ۑ��ܯ�����sY� ���������h`���u���\`9A�-��|�L;��%�����#趛��o�zԈ ��w�B@�l#+����.z�J�m������Pb�E	�B ���&�T�j�̝!��}+�\����@�W�p� �i��G*�%O� U_A7VB.{CSG�1�c�8WſSi�/���}�;K[K��,Ck�D��Z����ۙJ�1��'��P�����&C�k1�'<W�|�Tu�[@�^��SP�3�u�s�}�A�n���;���@�⌶K��S���tx�����j���y[�)�8%IiC��	��h�UI�Έ���|+�\i�<�굖�Q9u�a�^��ۿ�w\�^�<I��"�N㫴O#�,��^�uCJ�p���"����D�Y�7x�͟�0�����훼w�� T��츅���??�J�M,���+��|���S�AJǉvW�V��@_��2�1ޗ��wl�$W=�á��lwI����_p�d��ǃW�#ѽ9�N�f�l_��Pa����-�ӻYƊ\g'�J[9��~.��Zx+�Xn~��)ƎB��j���E����M ׂ���:To�T�eCA�$>&�'�.�fQ ���E<�ز R��j�zz��[�л�P]a�qd�����q�T�hH�W�z�ȥ�DDW�<�+4/:��;V�q&��|�s���X����tb�f��&��y\}f��EB5E.�n�
�Y~�搦�s	���T�{�_|i>I.����5%@��_GgK�nv�)"�e{�<E �)��N�P����U�؀��H���X���l��y�o�m����UU�Q8��:'k�]&6��/6�U�ް��C�G�V���ߓ6�G<D]�+�/��4����ޭ��>M	�&���`8<^�o�(zfΠ��� n�qX�����	��Ncx��(��Z���0���/�E��{�EG��+��y1�u�6���#hA�5�P{�v>[��3���������e�����Y��J�5+�L@��_u���B����F����]��J,�E�\W�����F�v��Z����u1�b�X�?0(���q��B2&���>�I�[�6���oh���>_�&qB'���C�<��&��K:�RLf���H���k�DJ/,�X��*�z�K�!�_�M��L�\Ϸ.%���f�3_Xcq}�G��\h�I`H���z��,�%�&��ad�����.��H��K�Ͳ�!�n��ČCc��3+C-w��u4�9 9Q�M#���ٲ4��j�@ر��؞S߲}-��f���*����X����*?x��GV��'f�sFKLHx1x|��R���сaOiĳT
}8��ė����e��|��2w�卺nR�2��[������1��G�R{�_A�^ӫ�gzL�8� ��k,2)���#et��ߕ��g��'l���y��E�fA@�+��t��6�vU6�[�����/p�A�+M�z��'p�oI����#�oΟ鐳�z����;��Z0(,�ɓ�U&�4���m�LM,мl�}�6|2(ru�M��T�_���^x��\Zc�L���a��U��hJ���k��PPxOZ�����ƾ�G�]3�K���������V��5v�!Lc`6���=��j��ܛ�q�զnƞGM�K�6�H~שt����B{Rf�;g���tI��p�6���]��H\*�gKJR��q1HU��gu[�����x��]ƽ�t�s�!��V:I"��6���9��~�e]qK"� �/ [0.l��7-����e�ꦓ�O�e���<��Ҫ�Da+�el�b7��<\x��?��ȖƄ�����tD�!�nS֧�y��&�Z	������:xV�w�U9<bx89�m6쟂��Mȃ�aʰ����5���*��l0��sp9��=Â����e����G"3�@��c��"���ٲRR4�3s�~�Z�:��V�`����� eOR"�]�o@d�t�uᨬP6��H]
�{}�����0g�4y���:zX[����Q3&>�#��w	��gI��y�@,����K��$]�S�'YT���{��-V�GB�7�_�`�w�z�U
��o�S 
�
3��8+{�6���/M2�,Pt!#|�`��ɩԘ�jL6��#�Q�nݼM�,C6V�~��xe�@�n:{]eN�r吃����X6����H�"lg�Uf�J41��~��Rny��^m�/�]]]G��e;�x�ӵ�F?"�>�
�+��~�5e]\4":�/W��.��7D]���b��}/�O>|��c*�IK�D��e���7)��<S|��-��M�BT-�f9�DZ���f־�	�����1s��G6�avlV���㬶-b�`Z�֜|얔���V�D�"�0�BϬ����`�����/�p0΀=��`�G��łQ��ޒ��-�=X�9&���^R)S36�3p���n�^s������L� \BVR�J�&�dYL��H��O4��Ɵ�HƤ鷇�y�D0Vy)�:���1_�Qj��>�~��}bag �y&f�����Kl���[/+SAgT��W�6{��k���7�%`)Ƴ8�4SQf��~����c�dЮ|-��n �`'F�h�B�Q��,ut��w-�����Z��8w��'��M/�za!��ya�̾��k���*�5���l8���YM'�^���l�����y���⫦�\�l�/n8_��(���[�&������:2x���F���z�ndL�S�5P����N6�@O�i<�����@=L�A����6��ֲ6��&�,�f�Z�L(����"��t�����Z�>g���f��/o �`J"@���G=�4�cӀs:|�	_���Ho�I�tf݉���� �wI*�@
V�\|0�$!CF�5�ʩ�c	7���Ibk�-��;��G�#�ML$e��wֻu˞�`>F�0�-_ѰCM#�0!�k�?u<�41����&B>�U�0���U_�N¥��!��b��q�k�����Py ɛ�$��{���;Xޣ�K�4����2;s����Ι�n��L�)Dh/Ժ�W��r0�c�We�Wm�v�>�U��>� ֟�}�������ǃJ����\�C���>�oZ#f̠P��o�D���9��M�U�+
H�ݧoo�	9�ex��g�(�u�q�+\�*�z�J�0�֋"ӗc|e�M4*`�7܉H6ə�?+���u{��Fa�W(�_��"���L�Y�mQ��?�PmD���g��п<��@�z�hL������޵(��$��
�B!�m^"���~�jm,��U�'��G,������������ 'k���,��6AEx��E��dR3l����j�� �^H%h�L��G��@�Z��;ȳ���#�~��ef��ۨ���(T��Z�Yy�@��l������	��]���1��i����58�pk���B5쭴��YЅlF7f�%���X<o*�ρ���ılS���I�`[��V\��4R	��� ���?[ؐh�	�	���[��k�����l
I�5���v���h�r�� ��IY�=���M�h��5��5�_���UK��+�7~���M��+'����I�]sꛓt?�=ڊ�;]j�a�a��@�0��<f�_)6n�&�4���(�Ս�vq�]ׂc%��J�.���F:��|Ø��ēh�v%��[ד��5�U�Z�E~�q�^�I�^H��)��+�2�Ȇ�޾�*г˭�0�_b���}��*q�9y�{���b*�Mo���n�Jw��B�`P�*��8���K<OB�ۜ`Ąs�&��Ew�uv|F�=�qش��QmCS�ĄUDq)	,��ӝ�2���eg?K|\Q�|�Ys�#���Rv�+�f�,
���h�Ç�������	�8�g"ن�w+{̛��}���<�F`nF?Fq08S
j]������)��W���)s�heA�=�dD��Y������ߐ��`��������)�r��/�C��$�⺚#t�ߝot�\��1U�pa���c%z:���L�M��~[4]1��F�@���o�8��K���'��
`4�������qF�+���X	��w���$glA���3b���P����n�m�o1�Ӽg�bΊŹ��2NB�z���)#�馐m>��2��?Q��>��G�(�-FJ����_@��f5�QXT�@0u�@G��L�ؙ����!��!�=K�~M�TttP�`W朆	ş.���(�,�!�yf���֎�r>%��'��F}�?�K�8����r���)�;���-k���-�M\BL2���@�ⷆ-&V�G\����b��CJ�իp��)�秸n��3n��0<� b�>D�Jw�t��T;��̝�+�_������܉l��@R@u��p�Ji�i��l�a&_NNj�-~���4wD�ԉ�ʝ΀�O[�[�'�Gc^�dc��;+�8�(���G���p�%%;�c�E���!�t41=�}�~���p�f�����a7���^����=����Mv�*�PA5�A���|�&h?/�$��0�{��$��YE����@�i�pg��X���ê�$Sz�ɺ!�o���A�~�����1���6ÏBÅ�ZB�S&�g���C�~֗{c���1���Eb�:%�yx)�ˠϞP� q�^[܌=�c���lQ�0{��N>�j�. �=�{22��[%e��G5j���w׻pv,���� ��P2➖�+�bD���Wz� s���/�������B����Y�cE�4��j=l1�G�f;����%r�G�*Y���uѐ+�&q���3�c[4�<��IQˉ�e���d�:@"�e�L[%3<��K|�i�DUa�9��N=V)@ �e�j����1�X�uE/{Q ��U�yߎ�@�����')�h�Ϛ����A�����K��Q���X��z�f�\��9V-x�� �-c��%���U�3q��he�R�N!Ж�-1y��������c���ʺ/� q/N-I3�jb`|�unP��y��I�p���[ J���������u~J��/�_�?T��79�:��:��,)���+�u��:�y�G�ތF剞O��E������g̦"��=��Qh\��H}}gOF�rTOġ�W�s')+<��r�\�c�>��s'�W꼶�[0*D)���n*{���z���$�b�T���\���I��I������A$�E	P�|��(
U%f6�7�3����X5��$��t��ߩjL�K��D�^��=B��M�+�i��ځ�8�j���D��|:���Q��.����� �?mg�9rM	���Hԭs����R����PilN�VUBF5fa�h��N�ő7ߤ�,#9c#�#��gk��l}�,D����0���O��xx9ijŘk����r�И�|N�EY��d�3xC۝�<
Pd�i��D��?����#El'�
�q�U׳^��\������/��7-���/o���)�,�ZM�"���B$Ф�q0e���ߖ�u�H��p,(��0Bž��3��W��z��.���e)>��N����J�m��&H���w]kki�4�g�-8��dR��D���[�X�5%����
ŭ�<�f�����]c�rY���t�:�8�-���nZr"����{~�Ap�M�N�+:Z�����L�q��xD�}����臂�#�ֆ�����\�a��"u�o�!9e�K&h��m �nNO/y�a2���9�3����f�;�d�<�[9�J��{� R`��>�H7Du�(&;y�����w�L�)M��VY%�H�GRmI������9��ۢV�$�׾�/�ڼ�c糥��0e�i�po��v"N�Z�j]rS'�3�L�ϐK��!��L�AG肀��Uɀ��|ˀ�&�š	Tt����m1C�V������׏������XK�Σ邃� =�V.T�;�6�h�<��2����yhQw��zT�(�@P�r��7�d}i1˾{�9���ե@)B�{���|
:���]�p}4
�Bǭ�O��N�.W����mq]
B7o�;�����d��e���&W�1\3�J��%l赹f1��VI�dN�	�)�:&��w_�5�$���1�rv�-����G�sB���꾱t���������"�����[�����pչ]ީ����N"&��a�=r�(��	1�Zr�ԅS�H����A���I���X5����@��r}8��.�|�eq�� JI\F#��C��r8 /*�96�I>s��-��QB�����?�KR�����ZrJ������R�q�_��8^�X�gl������r���w�,$�)��tD�镵1g�	�l��y�:�r���:A2�j]��t�蹫G�博�΅�/"�6A�;:��z�D��!��V�U�^��Z�N����j�{;(���E��R���mN\�,��/�1�6D��(��LMl�Q
�YÂ�c�ܤ���k��=����ƙ�'�>�P�\��i����Z�9~3ҡ��S����
W(�g�+!�hd`�Tg�/(j{3�S΁��n�qyM,}6�H�����f���>d�{x���5���Є۳�6e�}�*HN�Jg}��e��1���Y���*Չ�K�*�2]�]g��q[����-�"{�|�EX��0���0��]c��"�Й/r�.R7�j�����3RO9����u�m�D�3�e�7�<������H�����!�UDu!>� ��֙w�:?[��L��BC��"_VA�;���|b*s���S��1ܞ(㍃?�B��s]�g�������x�
�pkv?=5j��B����S�y,���2�� �����R�m:31���p`̊��P�yc0������� � �R��G�!:1d���i��*a��ߎ�mV��$�Y��O0#�yz�y:����L%�Q�+�>�ξ����g��Ty����K�^=��_S�T8��\�Q���9�7��#`Dbr��S,u�عw:�P�Od��-s��n�~�`B�ʅ���K}QB�������m-�N������v�s��ň�a��<z\��Hk�)�"��5G�GH�+��Y��Y�_��<+��2���,�.Ŧ�1����n�<��#4l�/&��ܳ�32����s���n��PS�[�V�������[mqi�u�����@xx�ܭ���=o�x-�m��A�%�}��Z������";�����>ZQw�g؇�fKW�o�fa�C��"�a��B�Z4�h��;[|��D�d�o�[bt�*��+�1 
�I�&6
T|KM�!�S��������h�7��I\4����V�T��b#���$U�+�Jлp����=����0��"�+�#�CM���u�Sw4,����.�>�i�0�)U��C��!�kM��kҲ��8���[hF�/��Ώ����l�XBb���!}�z��4I;.DU�0��0SZ�I0�܇��)ߍgh*ϱ�	�r뜲�r�1��<`v�-Uԁc>�⩟Ē�qb���q�e�X|��7`?��3>���#a��P�^�oqe��#�9���0��E���B'ќ�keӊ��"B����˽�D*�ǋ���z�q��Ӓ�!e��*�@�7��6D��?dn��AC����W#(��R����L�<m�5o?sf�Dޑ���>кH�P���5�+L
���V�^ސ���'��I�=ێ���^�UE��7�j���0L*�     i  �  �  [*  �5  A  WL  X  c  �n  �y  =�  M�  ߖ  0�  y�  ĩ  �  J�  ��  ��  B�  ��  �  w�  ��  G�  ��  ��  8�  � �	 J � t  �' ?. 
7 �> �F �L 7S 2V  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�=A!L&�S�ӰS�����<l༛L��5_�C�I
/y$Ցr�C	ʔ3d�O��"<yϓ|���q"��L��aрFF�1����`�^h�Q��hPN�}�d�ȓ!��x!D�<Tt
iz��ޭL�e��~��TbԀ�.͒��G+/���ȓr�]2)��ԭ��
�Vلȓz�<���!�P��fͬ3���(�����w���t,\�H���K�D��`���58�Y"���)A��=�����v}��B"���sΝ���l�{��ı;X�C���zC:T��'�J�x5��+s(T���	ف����ȓE��G���V󨤢�.�=x�i�ȓ�P��dC)'�l1�c��
Ѱ����`��C�
iv�@1
N ��Xpz��)k�<Bd
�>r���ȓ��
�h��l�R�ѻ�����)�J�0���Rn
顂�T/��A��L���S�)	�T\J�c��>�r��ȓ|6`IV�5^���Y4��E�P�ȓ�b�෠�3%�`��/@�J���NQ
\K�HJ'�]	��Fp/��� ���b�BA�;�:��L��K��@��}vMc��O'�=���4��9�ȓX,,����W�Δ[���L�&���T���'-JH
��ZT��,Z
�'	�p3Bl�v�`CRCς\Z�'��$B���q�(����"M����'���Z�Cq��%��K	=d���'�~�:�K
�gM+t"ݚ8�4����� �����H	��hT	�&`M�jY��HO?���<���K��ˉ�a�ʇ�<�!�.
��9����"�!�D��?�!�$ݨR)Ҙ��F�3\}� �)�i�!�d�%�����d�	�� ���/!�,��e�J���H�G��Y!�D��� 	҇��Q��U�Ɓ��B�!�
Xۄ0��݁�L5b��ՙ%�!��!��)�wI��'��L	"'_�z!�X�`�┥�6>��pQ#DG�!��͉să��w�e��ˤJ�!���6L\I*��n�����'JB!�ۂ�|�b�RS9��JC�s8Q��D�t���I��D�&�S EN	��n��ybh6S���HO#<����gR��~"�)ڧ
�~m��%��>��%�\\m��!�L��Yq����6ō��R��ȓ2�|�0s��+vS򹫑!<6J��ȓx�<y��'C9Y�D�3`Ν0{$�ȓs��MXIE=)�����*oHd��]�hX�Se�;�̵qEg��l��C�����8��1�e�^�F�dQ�ȓIȐ���C�k� 1ӱ�2(����u����呼	vzQ�jTl���ȓ>ܒ���!}[� �0�V�fxh4�ȓiw�0����)��0�%*D�|��ȓ*������J����\k<��ȓ1JX��i�,*����C�Ϩ���<2��(��6Q�6|�Gl,^�hx�ȓ�z�yqC�i�Eˡ��+���ȓ"�qy&��k������Q����[g(�(c�\�j�a��_6�M��A�Z���/t"@�A� 
�%�ȓN=�)�����jF.��+<@�ȓmTY�D)@)X�HARd��e��X�ȓ��u��%J�=��eb�K�N��Ćȓ������Ƅm�`�V� �Ƹ����i���Bvu`"Ԧ͖��X���ޱ0��:)VE�RR,HЅȓN��ra���R��hg�-n`(��F�D F�'`�,����G$�]��|�J�:���(��	>� �� ��"���*k56�MC��G{r�'��A��� W��9��J|HYY
�'F�z�*�*`Q9�%ARC6������x�,8/�V���L� W���c#%Ư�p=a5 9扡{�*`l�q��Ff�4��B�I�q�|���	,}�x�NU�b�E{J|juG�7`��H�G_�N(p�VL�<)Clə	d��)H�hlT�#��^�<���9)�����j4R��;֬v�<�ǒ���@R	��5�(�Cd�L�<�G���;��@��"ƪx�Z ��AF�<�0�X�%jFL��r��	p��B�<9�˙9[�$8dOH'��X!����<���)4���� �;j�ny�g�x�<���\0(}�1K�-�<�*�LWq�'@axb�H��H�2$�k��\�j�<�y"�.m��A6. ]�P�s"���y�N�61��#c�V�AB��y�Ά5xr�A��W�Trt����y����0h�J��R�P�^�21�ʂ�y��ۨ1*��I�I����ע�y�n��P9,]P��4Bfh��ɣ�y���� ؍��C�W�rAWF,|��Q
��'ԉ'W���\;����R��7x�Z�Q�'V����y�e�"�J=��
�{2��L����$��f����`�ѰZ���"O|�P���9Ct���
'� D����O�㟐&�L�,�GG��#�kA/(Ѭ�*7g)4���`��.f�Q�&)V/\=��h]n%!�$P~�i��M3LWF��4�Y0w-�y��I 
��A���`)�ep�!P�mښC�ɛ9(R(ɰ��S!~��M
�dC�ɏ"��Y�h��:�(兌!K��C�	�}!H�K�G���&���L�L�*B�0g2H5����h�6h{$B�&c�B�	�:X����3V��=�a̳.�DB䉜_��V�pU^@�vE�1�.B��(8�U �"��21\���N��r���d*�Ĺ�
�-�������SVν	bi:\Odc�@���*�`��7O�v��"�%D�����
囗b�4�M��N�40Q��>��ŌÊ)j�G�4.:%o%D���D�R����+�e��6���)s�!D���N�1:����}]��D�%D�p�ǡ��Ez�����]�1D�H�Ç���L���'o�����k"D���CĘN�p�kD�%~�Ci?D�t -��H�t��"��]U��aE�)D�|�Ѓ�.�qIW��TeU�2D��Ņ_���1�M�-�)�Af/D���4eտ;���r�g�Si(�K4�:D��s��/a��I��zl��m9D���榇�2͒�
1�P�C��<D�l��d�f h�hN�FI,m�Q*O:,P3�>0���(��'��x"O�倎+@ܨ�pE�9Hz�c"OD��,ܲ?�:� �$Q�o�1`!"O �����*mL��m�=M#w"O�����ӽCE�����/$쭙�"O�+�DN)ܦ����1Չ�"O`H��/ZF�� hb��2��u�3"O8�A�7q !fe�
pt�0IQ"O�����+A��:	�Y��"O���� L�Q����cT6�i"O��'�Y2!����߼GN��{�"O�H9�74�X
3kT�#N�Q"O.��ckN-E�|��WI�'?��9"O2��K��z��!)R�v�|@�"O��A�lM�/��������B�X�
 "O"Ԉ��?EE�`��.;� �8�"O�}�J,Զ�avj�#w�� �"O>�[WLPj���A)��v��� "O�1� ��b|f9�?�JM#%"OZQA�C�'8x�p"��a��`:"O h��P+x�lJ��,*���a4"O\���],|�>�I��Y=f��0�"O�G �(rޙ#��Ʋk�	�Q"O �RvfB�v�,�zF�:)�^�+!"Oĝ�@��pH|�P6�[h�*�"O@�G,�(v{&A�����^ѸG"O�8�r.V�p�
w'���r�"O8r��V�NeaElU$u�ڢ"O��ƑR]*=��k�*W�0}A�"O��p���DE��+�/d�|"OZtk3�S	�D�KS/i�u��"O��!�%z�^�9K�3s�*u0�"O� �- R����W�D�<оy��"O���ǙR.±r�
��L!�"O�E�a��4+�ֱ�B� >6	2��1"O��f *~��;d�Ԓ@�j�ȗ"O���f!�`�J�*�^�>��xs��'|�'�2�'��'E��'#�'�I+�A^$ܴ��P��E[6�{��'�B�'���'+�'_2�'Qb�'�{`�˾RO��A���'|�x JT�'���'~��'���'<��'���'�R'�X*J��l1� 84���'���'�R�'���'F2�'�'�P�._�Bi4q���H@�h��'FB�'�R�'j�'r�'}��'W��s&�y��E#uÏ�#���(&�'M��',��'Z��'���'��'oh�Ȕ�F�O�͛r��|��l���'m"�'o��'��'L�'���'���8�͙\E
%���D�4�v��@�'���']2�']��'=�'���'���p�� -��)���1`�'O2�'���'s��'��'��'�V8Ir�ߘH�2%B%*Y�`��=�G�'��'���'�R�'���'�2�'�b�fҲC�`�ZU%����q9�'B�'�2�'v��'��'���'��3C��xz�A3���k�e��',r�'x��'��'lR�'a"�'"8@�"$N�I�mY�	��N��g�'=��'�B�'A��'lr"`Ӣ���O��ac"�>1T����
y��*Q�Xy�'
�)�3?y�i�8p�aa��0f�'`�~4́���$�ڦ��?��<��4>عR�Q�gjH��'
�(*�K��?i��ʡ�Mk�O��S��
H?	P��ǡ`ʄ�����%�>Q���4�T�'��>���f�-$��(�6n�U�Τ�Іܹ�M;���Z���OV6=��|K爎�A<N-��K��6���L�Oh�Dv�`ק�O[�ysr�i"�� <�0ň��'f�z�����'6��r�tj�{+̢=�'�?���$C�`X��8�� �G�<9,O��O�qoږqwRc�xX6B�"�&��ݹ{�6�a��G��="�������<�ON���b+�N��Z��s������U^̡�3)�+U_"�韬��$Q�}�<쑦a��?�$YŌ�Zy�W� �)��<�j
:zⰅ���£G�6mY�$V�<��i+�9q�O��n�n��|�RN�%1�
�'Kغhi��AC�<��?!�na@���4��y>m����(���CB���E��*i�0�2�$�<�'�?����?���?��l�Z������ܰoon����O!��Ď����0/�]y��'2�����̇�ln$���.��ݹ��I_}"Iu�<�m�9��Ş��,�.\0A�u����,��,G�n�	2�u]҉�pMУ�j4�^w��O��'� �ppj�=�شΆ L[hĻ��'���'�����X�"�4|�@Y��_oB�O�b`}2�9'g�d̓�&�Q}b$j����'+`��ރ ��8���]\^X��߿X���>O�pC�˫4B�J��\?J���]�2��`Z��܏�":	Y��I�D����`�	����Y��5����$��4�A���p��{+O�������%|>}�I��M�K>QSOA gNT��D7T(���k�4�'�$6�R��v��$n�L~⦞�@�>�CPh�0~����e+��=B�����w�|�_���?G�Y�1����)ҳy�&<���	L�'06mN>s�����O���|�n�:}0��"��9���hT�U`~B��>i@�iz�7_L�)b��.�ڸ�C�dB,�7�%4�p��@#H1^<,O��H��?Q�9���u0��1A׺����� b���D�O(���O���<���i�v��NZ�b8xR%��"{�M�D������'��6�/�4�>�'��/T��Ф��&9��d�	�9r�'����i1�i������?M�]�T���������w~}s�}�Ȕ'Ur�'>��'���'����X���Ҁ��@c��5Y���j�4�zX�(O��$��.���OB�d��6��*��L�_ ��ꔖH9�pi��M;Ǜ|�'�r�'p{���4�y�$ŗhh�qcq�A}��P���-�y�:x0�IE��Iڟ��'���'A��c���%��iR�?~��'���'��U�kܴB4@,O����;���h�69�lm�&�>ƪ�Oz���y}��'S�|b��AKP}�R
Ի���0��Y����Z'��K���ɼ����s���.�DX)sxq���6:�Ի�G��3�!�DD�J2�!�B���,�w�U�uv^��ަ�	!�Qڟ��I'�Mی�wT��`�'㨘x�) �0P�8�'��6mDզqشHafߴ�� <a��9��[D̓�@NԴ#"d�,5a�i�'d-�ĥ<Q��?��?)��?�m�=��*���P$L��Nġ��dU���0Ilyr�'��O�R&��Hd��'D�%���x�aAR�l��?���S�'%DJ<{Pቓ%e�1	gAύ]�-pToM'i��(Orq�� �=�?yJ)�D�<Iw��A���n�cg.t�6i���?Q��?���?�'��Wզa�hP��L�bş�b�:t��O'E|��×A֟L��4���|Q\�p@ܴ>�����q�V��P�ɲ@�2[����_ ��qog~RD^�~���S�9&�O� �p@
J��y���4t!�!8OB��O����O\���O��?E���'#�ȕ($mǕ)>ӗMUy��'�6-C3&i��O*inZF�	�:�����e�]a�d(1 wX�h&���	͟�S0�nZm~Zw��P�#W�+6��#�.[�$���A�:7£�m�	Pyr�'�2�'[2'~69h�(�+ )��@�rZ"�'���M6$F?�?)��?9*���!�
E<.
�sc���Ұ������O��d/�)�K?]I@��udL1N����I!��+!.^pG̨�.O�8�?��3�D�S����+_�z������@6 ��D�O����O^��<�&�i��{3j
�'����d�¨
��Y{#@�+7���'r66�I3��D�O��S�-!b>Yc#�6	�p�4�<1j���ic����EGL%ji��&�Oy���K�R�Iԧ�������y^����ݟ(�I��p���(�O� �E
��2���h�3y��Y��m�r�3O���O���d����)f�t����/9��4c@l��5�f��	���&��ן�I�6�l�<�7G�Qz�V#"���6K��<�g/x4.�Iw�I}yʟ�A�ц�=T�(��+lp���'��6T�[o����O��բ,�����ȴ-9h�*FGI���RϨ>���?�M>� AD�@��`$��c�AJ~�*�>T��(R�Vc��OE����c��/Li�j��B�I-�I)�E�4g���'�r�'q��S��|&o�&������l��yā����۴F�PC��?��i<�O�N�5I��)) ���i���>:d�d�O��$�O�=	�l���ӺC����´@�@l��##̓�'�ŢALD9d�O��?���?I��?)� /�r��({�ܸ�1i�iv���(Op�oU4X��ğ��}�ğJ3�*��5a���0��%^����O�$/��I�`��b��"4`��j�$>憱
��A/cN�˓@�L�����O�9�M>�.O���AAW�D�x���%�"!8�m�O����O����O�i�<�a�i�b�ʖ�'H��iWA9N�8E*a�`��cKr�u�D�`��OL���O����%V�H "F�M��5�>`�h�S��b���ޟ���	ԊM��D�nyB�O:��C�GYb$���O*2�P�4"�#�y��'��'��'v��)z���`2��W�X�s���C�����O������� �Rvy2�a�P���<Q��O�B #��N `0���V����?I���?�҈ȫ�M��'5��.kK�шUʔ����pf���QZ�9���OX�K>.O��d�O����OY�IЀd_NP���E1E�d�c�O^�d�<���i��´�'g�'U��*b�5�eX�P)x�e숯!�J�}���ߟ���S�i>M�	�h�,t娂�W����gT�����¼=���{5�@oy��O��4�I"��'U�2���qaA⴪ʧ}� 0��'���'�"���O����M��&@�-�XŪ㒇@�0�{t�>cݠ����?���i��O�'f"�ِ2ԞD�R��_��8'G��	���'�����i�D�O�=9�����qN�<�Œ�Xiʄ���D�6�U+&G�<�-O�$�O����O����O�ʧ`9��9�uy˵M�
,-pE�vmۣ�M[�-$�?A��?QN~�Ǜ�w� �� 폠:t�l �&�GR�ؖ�'2�O���O���D�.��6�f����N9k9
q[S�Z1N����Ix������4"�b�uy��'Z���& ^(���KD>@�!�S�U2�'��'(�I��M�Ca�%�?q��?1V D�d��pʴ�"#���@4��>��'7�ꓤ?ɈB�C(W9�� O��!����)����$�R'��;wIX�g�ؒ����e�J�D��_�)�3��15��HV� ���O���O�$5�'�?��'��S�� ��	��X#AH^��?��ihB�2��'%�`l����ݲ1MD`:��[z2��E��i��	ޟt�'���HW�i����^�8�V�OHD�j�`�3Chʉ���P�L��z��Vy���X�Laq`�M�(]z���0�,�c�v@�r:f��O��?Y����d���kJ4m�0ت4�R:���CΦ���4Z����O�fa����q?� ��g��j�i`aύ�xapW�����<>��O�	ByҨ��Q��x+e/��,җ���0>at�i�Zd���'J��B�\ x��Hk��k��:��'��7�4����$�榽Yܴ%ϛ�j��-H#��.ܤj&������Q�i����7Pv̂�OR�%?��� V�d���M?,	�.��`3O����Od�$�O�d�O��?Iȱ���[)(� �?vtrC�ş���ϟ��شL�8ļ�?i��ir�'9��� Z�1�na��>;t�᷃)�G֦m���|�r�˃�M��Oz4i2��NR^��C�*���"��*W@��8��O��?1��?���r�M�D-̅� ����$�u����?)OPo�n���'m2T>���U�͆x����&TO4�q�%?	%R����4)Z�6'�?ɩ�]�I�EI��p7�H"�蘝z):�I�#�\�JȖ��TG�̟P*��|�o�BKqCQ�=\�dX�3^�"�'�B�'&���P�Ȋ�4&B�KT@��z�ܤJQ�K�5�5KA���d��y�	m�	������8jWl{W*J�O[�I>�������ٴm0��4�y��'mr�����?HrU�� �@rk\�b
D�r7A�i���=O�˓�?����?a��?A����0Jtt�F��<'TIA`疟.DIm�f���	���	y�s� ���c���/N:!�4��!��i��	�?1����Ş� <Hܴ�y�P
�w�H.0���!�b���yR� 4qp�������4���dH �̩
��� v#��9a� ����O��$�O��A�����<��?ac� ~Bvđ�y����$k�O$!�'\"�'��'H�j���vVՒ���	��O ��&/�8~?�7M?�S�q���O�K4O
�n�A����(�Zp"O޹�a����.ś2�ډc��huB�O|�m�.x�I����@��4���yW(ڲ4�@ �-+��t�U�y2@dӸ	o���M�c
��M3�O��k$(�+�r�揃t���3��,NZd&�עs�l�OPʓ�?���?����?!�I�tUض�3=F��b��	zm��*-Oh�m��L��I�X��]�s�,� JU4}�a*Q�M�5m8����OR��!����<�&��3�K��l� �L�@���>L,ʓ3MJ�5b�O�0�J>�-O�����D�s��re	%/dN�Pw��O���O����O�)�<Qa�io �e�'h���gH�g�3(���iR�'6� �4�dq�'v�7���1pشr�p�r���>��D���%U=�(�@�E2�M��O\���d_��ڲ�(�)���d�&�Y	�<��la��>O����O��d�OL���O��?5( `A�)��Y��MܑJY�<�	8?����vl���$M�%$���Df\/LqX� ��[�@U�2@h�����i>��1,�����'�"	7��d�
)�t@ӓp+z�	NT*B^Y�����4�6�D�O`��5������O�̱��I����$�O>˓ۛ��ȗB�����0�O���S�[�B��!���!B��p��'.�>1���?aI>�OM��yFE��S�*�p �U9j�2t���
�g�E95���p��i>�"d�'<��&��ڲ,��%%�9�!$���J"l�� �	֟��	��b>�'��6�Ϙ-�*��$ɞ,D�a�ؤjhq�(�O���٦1�?y�W��I�e�m�"a���P�%����I����'� ɦy�u�d�����%by2l�c�z���O�u��X��H^��yBX��I�����@�I�ЖO������,PHǍ<FaC#�k��9*��<�����?�Ż�yW�A�'���S���!#f� !�/UR�4��$�O^� 4�a�b��xƖ��7'ÌW�hl�T�L>"�D�I?}E2�h�'P��&��'�r4�p��\�k��݃6��1HVihp�'�2�'�W���޴n^Eϓ�?q���t��!�Af@O� $
h���k�>���?YJ>y�K�^�9�dd����� ��<�dFJq��Ϟ�M��O��)?�~��'�(D��\��}�ׇߔ��� �'4��'(��'��>�]�M�h�+���µ��B�%tJ���I-�M x~�p�d��]��\1h �?*z�Qc�	hr�	۟���ʟ�Pv�����?i������?mxj��t`B�.�r��ҁ�:KlD�'�������'���'���'b`���$X�J�:
vb j7�h6U��zٴw�jT����?����<�R��*u��T��G��2�����)s��	ǟ��Ie�)擡kn�9 ��#��k�"��cf�y�����8�'���p������s�|�V�8Y�l.9L�q��"�$��U�T�ן��	� �I��jy�`ӂ���G�OT��� ��`d�<h׶�S�&�O��m�C�i>��O �d�OP��Ӎ[�T=��!Pbȉ�G�/_ށ��oӾ�I
|QT��0��J~���UPT
 EQ5^� ���0 ��L���?91�ǌ'���weO3
���4�ܗ�?a���?�r�i\�͟� m�V�	!6Rd��T�P�"\Ȑ���w�v�I<���i��7=�*�,}���@<����]+T�b4�o�n{F 2N,����F3�䓮�$�O��$�O��G!��� ���;ĝ�p/�BN ���O�ʓc�F��PR��'��X>�[5�˝`h����K^���z3l=?�`P����ڟ�%���Z h"�**P�p0o�;ľq��� K2�ѧB�4��4� e��T��ObLtЀ9���xPm��2��(����O���O��$�O��
?FK�<��iO||#�
�]/��YVi�U���v���B��I2�M�J>a�O���ݟ���7��������U�8A1h���I:USlDn�<a��oT	�թ񟠜1(O������I���s�0��W;O�˓�?9��?)���?�����V�cv�s��v�B��fk
�F��m�F�RI�	�`���?A���ş��ɞ�Mϻ4��r�a��P&��r�
&<^(�H�����T�'��o(��=O `'��x{,�@ʟ�p5��h3O��8�'��?!W�4���<!��?Q'I_�����VH� �Rg���?A���?�����Ĝ˦C�������C�#܏;��9�V�̹2ǲ��Èx��ea���8�Iy�#=�dR��5 Ą��JՔg��j�������~�<ВN~� �O(���p0-5c���X��%i!�i����?���?I���h�V��D�dV���+�5uv�2�%p�K��'��6��"t�	&�M���w����gGa4	��(�gn}қ'�r�'�rlށߛv1O���P/1����π ̙*�dún\(������B�<�d�<ͧ�?����?9��?	�_@_�Q%� �ݓb�U����5e͞՟��I㟼&?��S�N�[U)Y"�)*Ş��5B-�>�`�i��7l�)��G#8�p C�w�y����2����A�5z�'�����i�ş��1�|�Y��;`��S���S�*L�S�`� �o��l���(������IyB��O&����' �\����
U3[�M��D�'47�8�ɢ��d�O:�k�(<@d��3���dH�7P{�Ea ��M�'��nO�(ܜE��g@��?U����$)�F 2|��!�d��[ˠ�	ҟp�I���֟p�Ia��}C6�kbǉ51*e�3�ƪ5+.�/O��F���3��h>��,�M�I>���P�~���ʀC+2꒸��
z��'D�7��ަ�S�*=o�P~"ѓ����K	u�a����d�
1������0��|�[�������������5CI��(`Ȓ)nta ̟ϟ���By��gӼ�<O�d�O��'KMX�����	U�82�N�+Y�R8�'���?������|
�`�<�u��r�G�+]��;�c�LlA�4������'��'�9�pD�0>Tz�Z���d����'{��'hR���OS�ɓ�M#���1�%+�G��1|^�KZ',x��'��6�,�����O`�C'�lh���� ?�U����O���W�W�66�e��I8�д{��~�*���H'eŠm� 9CQ+Q������$�Oj��O����Oz���|�Q���u0$9Q�	�F��<x���9ߴN=q.O���&���Oмoz�A�ŌX��`�j�c_��4���H��V�)�S�ve��o�<�v�$4�e��;c��4ۓ�<�1 I�W����J3����d�O����$v���u�ƌt��2L�o����O���O��[��HT��y��'MY'Vt��v��p)	5���|��Ox��'�r�'��'�ŀ���/kl����'�m�����O��!t��/a�x7�>�S_����O$�`"h��|��{�h��C':y �O���O<���O�}��DW�t�Hf�a��!�Ca8��%ӛFj˶,�R�'7�6�)�i�E�E��KQ��1���<6%��h����wy��A)6o�����c#�Ѱ[��̌#J�E�#��Kׂ�zt��<\+'���'�2�'�R�'�B�'��`�B-�$���d�L�p���Z��R�4u����,O���?�)�O���f�ɚ-�@&/ �P���+c��n}B�'��O�)�O��e<~}�"�ϗ=y����'ؠ��Eؗ.Mjʓk�`�"��O�4�K>�*O�t8��J�'��qx�c�9T�����O��d�O���O�)�<�P�i ��C��'fr|8W�	�Q������
R��Zp�'�6m?������O���de��B8~�=�S�S#qi�!��	�M{�Oƥa��ų���6����~�k��3�E�d�N��s�0O���O����O�D�O��?͂���5C
�%�r�P�>�P��H�my"�'��6�G4l��O�m��I"&�8b��B�Q���/�6�c��	Qybg#"ԛf��0 ��$!dL�	��K��������~l�'���%�d�'nb�'�r�'�X�	C��=�r%	�G3QH���'��[�h�ش8�H�q��?�����iC�t�F�('��4��y�i�=n%�	���d�O6���ʟ���\��슆d��DRސ��,�=@���`�O�hM�y�'���Eџ �v�|�o�dB���0b�	�c<�b�'���'���Y�ȊشrR�$�U�÷|�& #�ᓦ5*�5��b~"�`���4٨O��D6 *�ɰ�Er�2a�I��o����O���Oc���Ni�lr C<Cf���a�]��r�D+��V���|yb�'U�'�"�'U�Q>1tNշ��p�-T6[��:,�0�M�$��?���?A����9O�lzމ4��
R��j���6g���!ʜ��,�?ͧ�?i��S��۴�y�o�.+!��KF��!Z��{��ѣ�yB��d�H�I�'�'��	ş���e�]X�%H�DG"�!uf%\���	��D��ܟ`�'Jr6- 	6���?�u�4WFT%��l�=e"��Ȧ����?ISZ��#ڴ̛6l$��0&����� ����9�+�:\Q�	1#���W�6u�|�$?���'�|��	>���w'�+{�!S�QV���IƟ��	����	S�x���'+НÓhՉ���0����@�T���'�27���2'���O��o�q��李���Ӵ�T�\�n��'I�K��	ޟ4�I�,��(�IΓ�?yu���6����U�J&\��K#���XԂɟ2%�(�N>I,O���OZ���O��D�Od���ڞdUfM��"[;��d��Ƞ<��i��y��'��'��OK��.�� �O��Z��Pr�"Z�>j��?���O�r�'f��2��# ��Y��5 �4� -��AT<(ze\�@�ǂ����c�	vy�&B�[NXmٲ�؎{���7��ct�'�2�'u�OU�I��M˥e�1�?	�ć�-���7��&i����2�?y_����?��Z���	Fy�F#Rf�P�!Բ@�|��� �'d��TK��i�����A�O.�M%?���LN�+$o�
`ɘ1_%~X�����	����ܟ���B��	�x��G����ZM�lKΌf~B�'�6-X���$�M�H>��ʝ ]��NbQ:�������?a��?�d"��M�'�%F��� D �a��Xo24Se$G�r�@��~��|P��S����IƟ(�5M_>S��x���j� ��w �ڟ$��Gyr�xӼ�X�?O<�d�O�ʧ|�ޔC�26�����=�F��'�4��?�����S���Z$Ms����@ڝVs���'R�
���Dk�5u��&����$-��D.���Uq���S(C�^�p,A�k ����O�$�OP��<��i���
 �ӥO�H�2͚2c=3��:���L��?�f]�8��&	��в�C	/�ll#@+ɛH h������`Ԧ��'�,aQ��`ܧ>+�z����zP����Jg�e̓��d�O ���O>���O����|"�j@�)���;A����\(`�F���m�&�y�'���'�26=��P��څ^Hn�)U��-̀R���Oh��'��i��o�7�v��:�#Ҿfi�5��.e�0!)D-k����f/X��$)�$�<�Oڲm1�VC.5`��E�D�Q
Ó��&�fT��'���%P����M�Y��x"4���\�OX��'��'��'���IA�I�x�(��(G�����O�Qx�	�jk@S=�)��?!�Oz	����L��l�iA�i�h�rR"O��R�G(���.vHe�F/�O��m3�q���L[ߴ���y�M�/C�Qa�r|f�b@��y�'��'-�1饱ii�i��c FI�?�2�B��&���b)�9<�ʁB�j�ma�'��	X�'޸!����.^�ĂS�Ǫg_bl��O �mZ5H��m�I����V�'J�f9x!�G�J�8B���X?�Za_�T0�4��6�'��ɗYz�$ �n��u�T<�dF���͙�U�b��c�nd�G�O��I>�,Oz��*T�tIЄ+�@��2S*�O���O<��O�<���i\.M!��'��ի&�W���pґb<�vp�1�'�@7�3�ɓ��$�O"�$�Od a Ɓ45{6�aa�)z@��D�H?<7�r�,��yٚ�P��O`�L�'t�t�w�:LQ���-AKx�`@���#�Լ��'I2�'���'��'�2��ƏM�n� ����؂p{7��O����O&alZr�d�S۟���4��N�в���C�R���M�w�Dp�L>����?��?{���ش�y�ԟD�O�#@�P) �]���FT?9����䓻��OP���O���ˑ�0=I������J��=y����O��uśf��P���'C�Z>������_��A�b�J�@�̝��O<?y#T����`$��\����r�C���R�ٸD��|���+i\y��/��4��H��%h��O��RD%�46�t(�^,/>t����O��D�O,���O1���	���ˁw�J��&���)���0aF�[��p�[�48۴��'��ʓ�M��G<h�J��T'g�z�NZ�q��&�r���f�n�"�k���ad�p�K.O��d��?2�@�1Gē)sEz�#0O^ʓ�?Q���?����?A���I�:r�^L�A�_C�m�ࡕ
�x`o�~i`%����	\���H����{��@>Rz@ ��^��lug*��G��j�Ĩ$�b> ��զ�͓<]���1%ɒt�,�&DV�qK�ϓS-����On�SM>�/OV�d�OR���:AK1DZ:8������O��D�O���<��i�����'Y��'P>��F�2����Կms��`��'i�'����?���6Z�@Kr/	�a� X��y��'��x�dZ(dD0u�X���Ӑh��a\�Q1���Nq��)�M� u�y�4�Dܟ��	ڟ������E���'P�a@�)-;���4.��g��8��'**6�0V�����O��o�K�ӼC��	(a` ���%80��(�<����d�(�<79?�c�E�/�h�iщ_Xp9�dI؜G2��b$E�L���O>�*O����O~�$�O���Ol%�ta�@��$!c	P�Pk�4��<���i�~�S#�'���'T�0x�]	%�����)ǛXXM�E�D}��'��O�	�O4�D@"�	[��H:U���"T)�KJ�s�E�0��jt,a�n�O�;J>y-OL<RGm^'o���I��8L����'06�̰yD�DJ4�X����V�y��H�ʶb��ăȦ��?	�S����4{ڛ6d�V ��ŗKP����P�e�j9 �t=�7�7?��U����I��䧔���l���U�*ޗY&t(Ee�<��?y���?Q��?�O~f�I�c�la#�b �\����N� ������?���or��-��s���M�N>�$�?��eԦ7�n�%�Ox̓�?����?Y��&�M��'"D�%+��`��}�=�����|X�,�&����|R� �?YS)�	\tq��k�7+:�Tb�u�'�:6mv,�D�O���|Z�2����5���u>*����q~R��>	�i�D7��)��N�H�|���N�d �\�%��!�6J&B��h,O�)��?��9�$�j~��h��ڰ�KY.y9*��O����O���i�<yV�irzTz��"Y:��]�F��e!� (g���'��7�8�ɐ��D�O"�RE&׷jf�y	u�R|�u�� �Ov��H�6m2?��Gf�q1�'W||˓
j\E��N o2��{Wc�"Ex������O^�d�O��O��Ĩ|�����
=���ʤq$�T�#T�]]�V��
uR�Iޟ��OV�'�d6=����D��l\�r�̈W�5Z�L�O�������I�ҘDm��<� Zp�a��(� 3���I*�r�;O��1s`���?���'��<����?��`��a ��@`eЫ oD�c ���?Y��?I����Ħ)���U˟�����X��!��_���
�L�
�"�L@g����"�M��i)O�EE��1�� f� 4P�	唟dA��T�SN�|
C*TL�1RG*ޟD���h�&��!&fytSDm������ڟT���pE��wR{�D �BŞ��#�T���h���'`6��8'x��d�O�EnZA�i>��;,�h����Qu��6ʽ�6�I�M��i��7��($t6m+?i�m�t>���-O�`�Y�ሃk�(@*���4Bf��N>1.O��d�O����O����O�My�&�x����mC�͘���<9��i_L���'�B�'d�O��a�)6�Aj� :V�p�T�Z����f�`�Ɯ&�b>5w�y8lԚ��o��r�e�0_+����#[yR�]��z��	�l��'�剰]�	��׌D����3D�'l�D�IΟ���؟D�i>ݕ'-�6-H�M����!_g�,�V�ҥb;|e��` �D����զU&��S�����k�4w���"��N�0�g��h�"�!�G��fQ�1�e�i����P��O7��&?����l~�hb
؇W�p����Ѥn���l����\�I�|�	S�'x��؉�-�$�����Yr�����?)��S��l���d�'��7�?��V*Lb��0��/w�Š���(7}j�Op���O���]5�63?�;abHc�O��(P��A!8mH��e��?�q�+��<����L�j����Z�<�(S�X3�O��oZ�x2!�	��I`���T[6� �Od�.ܙ��@����X}��`�ޑn���S� R�9����A.�>ٜ%c�b1"��c(�[�y�Y���&qz�ev�	9��[F��3�ؔ���O�09�����	���)�by��eӞ}ٲ A�4��U
�:{p܁a<8
�q?�F��H}�K~Ӑy �_1#�h���c�Bڧצ�#�4U��M��4��D1v#���,�<�ӥ��,z1�O5{>��do��<�*O����O\�d�O$���O�˧"������PVǬ񚒫��4pXоi�F��'V"�'L�OU�q��.�}zP!9��U�0�eH�?ݲIo
�M���x��d�[v�&3O��If�C�ca�A`��n��<O64x��҆�?10�?�D�<�/OXiP���+'<�r"��],t�A�'{�7�ȣ=�����OB�R�vt�S2
��<����UW�"�(�P�O4��O��O�"m��^��X�$0a��a����CeI�(�x�c�j�ӕ)��\�����K��b�x�/͑]G� Ӳ������؟L�	���'?E"�kt>��I:(�>Ȁ�k�y��L�:E�a+!�'}�7̀1n��R�Ɨ|b��y�!�5"V �(E`�:�"��_'�yb�'���'@�c�i���O��EFJ?��FD-g��tjQ� L�ꥠe��cf�O���?���?���?���2S4P���-7�Q6��
'����*O*l�*i�T�I՟h��V�s����O���S�À�D�cҨJ%���O<��>���I1m���R�&	2!��	�R��	{,\�bD~��;���a��� %�Ԕ'Ɍ�{�B8q��Ve=�<ɐ��'>��'v2����P���ݴI���y�∘��/;����F�_Lل4̓2#�6�DO}��'��'HZU)�`F.tl:��e�V�*��!�iȤ��v���#���VSQ>5�ݲ+	&�q�K�R����.D���Iݟ��	���I����IV����D-S+y�ޥ�#*K������?��<�fM������'MR7M/�D��K�s�\�-�ĉ��̌m���O����O�	Or��6�/?��f�&�B�
=�`�XԨAqb�C5G@��?��)/��<���?Y��?�I[)VK�x�JU�+ 98��^��?I����$��},j����O��D�|:#�0%�1�C��n����jG~�l�>����?�I>�OtptH�\��j`MT-$*�Q���G�0�+���"q��i>1"')�	�4���G�Ue��G�
2�K4�g4�9�Iȶ-��H�@Z�^��������;�L��u���Kl$�PrOŬ�,��bG��,"�9�kՈ�j��fB�8+s��9��p���
u�zAaB�9"P	�iQ��:=��g�� ��>Ŕ�Q�-��%�@骷���C����8Ê��p?�	a@��4�$��(��	ؐI�4�<�B��Ȑ�C�f�
Q"�I
��1gȰDWy��营
���u"�g�|�����W����Ӥ�f`��S���� w/��:�>$�%(:�f� b��r� ��C��'��|�P��KҊ�?vL���G��P8 �#���b���Iϟ4��ny�ɓ�8��~���n�O�X���J�[ .��?	�����d��c���u��az���95��xqP�ՉE2��?����?!*O2�{�&�[�S�e��,{T��,U����&�J��Qܴ�?�L>�+Oj� ��d�0@���A�C)�����C&>N�f�'rP�,��)W��ħ�?��� @�(
�[������F T����a�x�Y�(( ?�S�T�V�_�Y�/�*�"m1�.0�M�,O�)	P٦�3����������'�p�R�ĭf܈PB�����Hٴ��䄱��b?]�#O�'�����+w��e��duӞ!��#٦=����,���?8�}�NX�u]V�Ѥ®W����Td�+h7��'��"|��5�X�[��W"�h�J\3`="�"a�i���'��ַQ�
c���	���� 6�����,8U�2,ρz����@�1O��D�O�����5!`DRgC�?Kbu�J�j���m�̟�CI�ē�?������s���5��l��F�EJ �A -�W}�,���'��'��h{t�Uo
��!��4@��1I��`V̨%�����%���';^�pg ˟@�$l��jƼh�f���յ�'���'12Z�@��+@,���d��f��ԛTJ� VP��f�����?�O>�/Ob�]��SF�{Dy�T�js#囫��$�O@���O^˓]kM귖�tF��#�ʸ� �]]��"�gK&s��6��O��On˓�l��>�5�Ѵ5�)����;�ư0�)�ߦ��I��ܗ'*n�C:�	�O����4u����M�м@ǁ�{.i&����t�X�g*�1YNLpe-Ջ�7ͱ<�WD�(��&�'�r�'��s��X�!���&hP8�촁�딎"p�6��O��K��f��!�$8��"vN�����;�I��I?&�7�^$M�<o�ҟl��ɟ���1��ĳ<�#�~����"5����#��(}�+P���On�?��	�B�:�`��5gjY��d�7' ʉ�۴�?����?���9Uq��uyb�'���ya@D!d)N"J�;��E5Yg��|��U�2_��������i���4
�O[R�*$�ۿS	D0T�n���d�B��x�'����d%���/���e��AwP�òh��J���H4�?�$�O��D�O˓Hg�ə�m�ni@Q[Fi�
n@��`2�ٜ���sy��'8���t�	����B4D�8�:A�M��SG/L��\'�X�I�$��oy�b��U6�S�rł�3P	C�&V��#ɕ4�.7�<������?��v�vs�'+�*�:A���˾M�t�O����O��D�<3�̿h����*���[\�C�'�*k�b�R ���M;����?1��Eΐ�b�{�K��>�j��e�TZ����ˊ�M����?+O&)�4C�_�d�'��O��P�A&~���Ŧ�&V�,A{�M,��O��dѷ+�:�t�'E|� �"S�]����"04LAm�^y��ô���'��'���X��X1[bF08�%D$$���c̄ p%B7m�O�����4A��b?�"ǣ� ����f�3N�u�CGp��C�@�A�����	�?=3�Ol˓���R%�B�SʤXǄ^�#�T�ƶi�8��`�$5�S���ӎ�n����Yz��xc��y���o�ğ���ݟ@s֊�����|���?��킀.�*(ha��b;���ĬJ�sϛ�',r\�${��X�'��i fm�g.���H���,�'e�F�h�O4�)Ub�<�)O��h�פ�:>"B� �Ο�~���0
��ē���<�����$�O�P8f���|�@	bM�Ff�(ia$��?1���'�2�O�|p� ��}���+�����i��8�y2�'���ߟ\;�or�#$�T����H���S��������D�?����dY�ěgQ
D|�s��!9N���o
���?1*OP��PA��'�?������[���t�B��T&\Hڛ6�$�O�ʓA�m%�(����K/>=y!�X#~��;$v���O&��rA�Z4�ħ�?����#�+5�����*}kTl�G+�h�Ky��'/����u7��$/�h���M_V�B�)	�����O�S�
�O���O�����Ӻ�ԚC].�jt�Ɋ-� %�U��̦���Ey��N�O�O��e���PZ	��m_�h��H��4�&9��?���?!�'��?����e��|(�86mX�����MS��Jp�|@�<E��g�/�Y[#ڊ'���Ԫ[�Ur��'+�'mj1Q5W��'��$*"$K�!��n����2���$9��Y�y�+ԩ
�P�d���O��d��a
^���o�Z}���	 y�(5lZ˟lۤ��&���|������O\�z�cWT�P��0b�5l�xMC��D|}�'1;�Y����ʟ��	dy2�S)(	qul؊XݒE@�s���;��2��OD���O�˓�?��E����`[<EF�
SI6J��Y�"���?9M>)��?1-O��u�W�|"2�G�X?�ȃ��=��B��a}r�'���'T�៼�I+X������
x�].4��bg�ߝD�tl�$�ۑ��$�O��$�O�ʓ9l������T)1?������D�D?���M�%z�7m�OԒO��P��}����S yW���1��9A�h���ДZ�V6-�O���<���ۼ_��O\���5&�E>90��3�&��=��J�%��ē��$ί���8���?�����\57D�%��+e���E���h��i�R�'�?��2	��(>7D��"�=l�����#<6ͦ<	W�X��?A�����ܴDg�B6��;`qީ�f��"L�2 lZ j������0�I����{yʟ �$�H��Px�O�"�lh*U�צ	(Gx	�����rL1�����h	-|xy#����M���?���ǁ�'���|����~�̿ta���x=<-�-Z�0�BP�H�6�]���9O����O���_�8��]�#f
M����0Z��m���lBE�	����|�����Ӻ�gϜ"�!��L��3�� ��X}R��hv�U��������	Vy2k��(p�G���(p���oďu��i��"�$�Od�-��<�� ��ҀC̣M{�,(q�ݟM(���d�2�?�-O4�D�O��$�<��H�
N󩟡K���剓9P^6<a��[m�I��K�	nybhU���+7n��DD�h�,b�� �ꓼ?����?�,O����P��'�iʥ����H���p��\B�Fy��d�<a��?Q��#��<Γ�?A�'y�9�G�Qyz�G9�l�۴�?�����ě">�L��O��'����^(S������f� ���N�!���?I���?Y� �<�M>��O�B` �%�!a����+z�۴��$Ļ��Qm��D��ោ��������(V5/v�C��
Ct<m1�i���'�L}x�'��'�q���:e�,�d���N��}+��i>� k��rӊ���O����"X�'���'[U�<I�O��>�ry��0J��u!�4[������Odb!I�y(=S�E*c�j,Ҩ=��6��O��$�Oxi�G@R}�U���ID?顭I$�ek�ȇ�A��d��æ9%�T�Rhn��?q��?aI��u��%�G��\��������'S|1�Ģ>Q)Od�D�<Y���.��y�P�c�(��%�ԄSLUT}����y��'���'i��'h�I�S�<�ˆ �ZnZPR@�	d` ��r�����<������ON���O��鄭�G��)��G8;��Z�c���$�O|���Ov���O�˓~yJ�X�3��@ 䢔�^� �(���5)PH�Y�i��	���'���'���ɴ�y��ŵОɚLF�i 
�g���{{�7-�O���O��D�<	�o�4d��ܟ�X�p-�1bSl�6���D�3UL�6��O�˓�?i���?�Ed
�<a+�f���@t�����9\��,���ͦY����'_�yK�N�~���?��'^��!k �Y䄩0��(fp�(i�R���	ş4��-3c\�'��Ĺ?��QF��3߸|�gD2k�tbc��ʓo]�]K�i>��'���O��Ӻ�&���z���jb��ECrͨ�/ئ���ӟH��m����yy��ɐ�G�Pc��rl��� z�f�D�j��7��O����O���y}r_��RwhփDu����)Il@� ��>�M�&��<�O>a��$�'BI�J͌ڌ|	�팜GF��t��j�D�O���'����'�����p��I�f �y0�my"��%�@!o����'w��r���I�O����O�k1�dct��g��VP����U��0�N��O�˓�?�.O����-������d���MxtQ�d\�Ry�ȗ'J��'�2_�L3R��Z*H�X$�Υ�z�a��G����O>��?�.O<�$�O
�DC Z	��҄
��֑��)Soj��0O�ʓ�?!��?�*O"Aڶ�M�|���ɠ���Jڃ[a��������'�B\��	�������I�AT����<:��Rd��-�V��Oj���ON��<a1LQ����'�4-�I'hd��q���M�����O����Ol��$:Oh�'[N$u�D�S�����&gOrR�i���'��	6=��ѹ��f���O0���u���i!�) ��}���[+O^�'���'�����y�^>�	k�k'B��c���s�`:�h�⦉�'߾5�Shs���D�O�����`֧uMXyμ��O9y*<i"ҏ�M#���?)�"��<�W?��yܧ1BT���;��Yc1��T��em.-��:޴�?���?��'"��	my���+dP�3EO�,H��#¦�\(B6퉜Fh�����2D`b�D�gr��$���Q��iYr�'���
�*�D����O��	&(��u�D(F?u:��Q�jV�IB 6��O�>@V��S�4�'YB�'��E�T�ߙ w�eS#+�-F�B��s�a���䖆{k���'����d�'�Zc���W��,�Z�;P�M9r����4�?��JI�<a/O����O����<���T�0 ���6��R�U6F�y��Z�d�'�2T�`��֟����?��@5�? Mpk0��W��R�y���I��x�I�X�I}y�B��+^�擾(	���b�> ��-ѤA��6M�<����d�O@���O�a @=O�i��E7ʝ�U�A$ r>��qGЦ���ן��Iʟ̖'��Q�tN�~����E.�9{v�(hǢ؝C&ԱB6I�̦���]y��'��'*()��'��I�s�R�>���w`^"7��H{ٴ�?a����d	���$�O���'���JYj��S��	8����J Lf>��?)���?����u~BP���'P���:��y���;�%�1�<Yش��$�:�8�mZ����ioZ�?��O����T�1�ݜ3�TY�D埡!��'9�
��y��'*��'dq�� '��u��Z�Ɏ_-J��$�iz�+rӼ���O2�D���M�'���6	� �w�ܤ[�*X[gZ�EGD͋�4^�JM��?�)O�?)���z|p�r�#�x��j��β,2���4�?!��?Y`I&��	Cy��'���`Ί-9T� 2c���	'�F#<�V�'��	8�2�)����?i�`��ѽA��rA��?��@#0h���M��4��uZ�W���'	�[���i�����8�>Q�8B� �1:(�d��YΓ�?����?����?A(O@�XR$E�@:�`���Z����AE�2D�Y�'���ҟ�'�r�'JB�A+
�V���zb ����%1^X(�'���'&r�'��s��fI6��D���҈s�ߴb5Hf/]��M{*Od�ģ<q���?��a�\Y�$"H��B�g=�m�!��(",< �\���	��D�IQy�F>-�Bꧦ?��"NAX�`��ns|�h3�ȣ_͛6�'���ɟ������:�j���	�
� �Aj�!�j�����^���ixB�'��I)�"�⨟����O����H����cMW�5�|m�����G����'���'�B-Y.�y��'���T�P(
�`��0#��9x�i��cĦA�'.����#s���d�O���蟌i֧u!\p�\�Fh;~�����޼�MC��?�0A�<���?�����O؈H e%T#�n ���*�-�ߴ_�0��W�iO��'�r�O�O���)�6�I����\L��O'j�oڭ`�*�	K�F�'�?�G�b��D�3$'�r���%Q�pқf�'r��'�j��!:���O����|�Ʈ�:W�(��c'�

=^I���w�ГO0k�aUo��ܟ�	⟴+d̉1�8��[�
��%��n�؟ܪ�â��'���|Zc��AC����(�pq�TKR?P��ڬOް���O�ʓ�?�����'<��
Uc�g�(�[GI�	V:�b�٨,6�'��'H�'��'�
�R�E4#�l̘���>@��@���yr^���蟐��yy����F擳az 
�#�+0���1��R��O�D8�$�O�D�Y���A�5В�zs�W�"Θ���زK4���'�r�'�V�\ �����'d��"�jS�hԸ\�@.H��<�y�ie�|��'d�����>aAʋ�,����� J��yk6˂ߦ���ܟ�'�&�)e+5��O��ɉ�.�b۴ė=w�z�)��2C�8}%���	�0�DL̟�&�t��j9���U��Z����L�-g�qm�wyBI�f�h7mW���'���6?9P
C1D��a��eY)��Ś�֦e����`*�e���&�(�}�R�܀	$Z�0@�-r[i�eM֦Aa�Ė�M����?I��%�$� ����`��0^ü���	T*1��o+S��	v�s�'�?�G
�N걑�����%��3қ��'��'H5��):�	؟8�)�8��S*��XH����B(oF�IBb�)R��?	���
�q�e�:z���ک(O4�ӻio�.:2GDc�<��U�i����$�&y �)�(��@�JJe	�>)��έ�?.O��d�O*���	�'L��}���B��\�� ���ǐQ�dd&����ן�$����ן�
Ц��{0�=;�#�`��!����Isy��'X2�'��	;@X !��O�6�3D�m�0����&m����O����O�O����Oz�/�y�ΈT� @ �獯d�tř�$�_	,��?Y���?A(OVt���Gn��4 C��F�L��6���,�d�F���4�?aJ>���?�o��?iK�t�1�J��>��A�9�T}������D�Oʓ<����e��d�'I�4���#����fB�A^�=w����O����O0�� �OܒOz��n�eQR�<����5 ҭH� 7�<A�jL,P��6�~
�������	�xєY4 ��#����%a�<��O���FG�O��O�>�f聽M��桓6h,TH[�!~� A{��^����I˟`�	�?uH<ͧX�����MO�)��וn�ms�X� �If�S�'�?9H��4��4��P�%���E�<;�6�'^��'��D��<�4��'T*�HnG���/��aѲJ��MS�2$8�)�O�D�On$��fр�@���+��N2df��Ԧ)�	4(pE	J<ͧ�(O�hQ&oա9.�Da�$]u��xE�x��'��I���I���'�E8 �Sy�`�sa ��֢�P�KS�8O����O���<����?S��L��a��̐h|����/r��U�<����?�.O|��O�}���$�V�4;C��t1�q7I�H�>�m�۟����`%� ��Ay.��M3J�r��Ju��:ޤ�&K_}r�'w��'X剼h��5�I|�Č��6�Hmt	P(H�i7#D�N���'��'����=. >��coä~�Ryi����F��7m�Oz���<��mUt�O���O>,�m�`R���g �<[|d)%<���O ��'[T�L�'~�Q�R"7�l�A�*�l|o�|y�#U�u�6-�w��'k�Ԉ*?�@�%C�:G윒,��P`�ަ��	����:��O@�DQ䓵_���S2�
�j����4	(x���?y*Od�)�<�OS��b!�;e���Õ䒖3LDܓ���>Q��Q���O��#ۇK 0n��#9�[�06K�O,���ONh�Ɵ@��ß��{?qeU�+�`s𩅡�d�(0	�y؞@�Iǟ����&��9
� Ƹ0#P���a��D2�4�?�5CJ&�'�"�'-ɧ5�̝�D�|��`�;L)&�ÂE���F�G�1OF���Oh�$�<qU�ęF�=���72���E��a���x��'�b�|��'�2��4�j��O��I��l�AG'wb�ۊy��'02�'��	�h�|��O��sK�I:11l%J�j�K�4���O˓�?���?���^T}�.
�Z4��dn.�4��C畇���O@���O>ʓS�	�U?]�I�Z�l
�-���ܙb�
2�F���4�?�)O����O��D��z�$�|2$-3Q�UcEiεX��ؠ͘�����'�[� B�#��	�O4���D�T���]!"���N�h�}�Y�(���|��qo���P��' �IU+��р�舕|�V� �%�4K��vU�,�����Ms��?������U���5^x��T5e�� p�mI�'�&7��O �dM�Q���d��'�q�� ��"���B�l�W�A�= ]�C�i"a�A"|�\���O��������'�	//�N�����-P	�$�sN+Q��K�4� �'��I�'F7>yo� q��!�c�||���"���p`pB�I�>(��W'eӜ4i�A��D*^��Dފjxx��oV��Q �,"vu�0�����`��@�c,z�`c�P�_tl�qm
J#���#�8
&չ��ʝ*�N  �
� ���0F&1f�[v��:�X���MuH
��w�Z�{2�b���D��%C:O*��'�C�-���PrFCK"����'IT�=x�% l��'nB�'��� �'b�0�f�w(}���$F�W�r��*�&� �y���J	�|b�~_��P����������J�F�V4��DQ�r�'��k�h�:h�����f����@�|��'�b��?��C�)�� "��(v*��+gk D��i��ٴt���kQ#2��p02h`����4�?�-O��˅e���'I哙'eB�ˡ�ӝsU�"�ʏm��[�)�����Iݟ��# �%"�%����D`m��S���E�h�UBK�0jL2�X1�G�(O��`CȲxj�rP��(j"��x`�&Q���˘$NT8�Q�I6���Ol�?i�dN�X �lYFB!@��uj��q�(���+m8�`��8NwHc0*����e�	"H.qA ��!S1(yԦ��8t:�Ie|V2�OX���|���� �?��?�HT�.����;	��ы⢗)ښ��,߲vJ��CP�I*�c>�dC0L똝�)I��,��r�6D���{�LLɰiN����)���(�x�|�Â�Z%Ĩ(5&/x�R �I���'��(?�<��4{�BH3%�H�l���ȓHn��6C���1�'�2�~\Fx2�*�S���9&��c��D����E�K��'���fа]W��'Y��'� ��֟�ɚ��j腱1���3���y����pHj�����]!@��Ơ۳����99�B�U�ָ��I�R&��:DA��<(�[�	٩j��	!R����OD�O����OH˓\It8@��>;Kʝ��$�	�� ��-bS��[�N/�8�4 K��+��)R�ʮ�<8id
����A	3�y�XD�ĉ*�iN3��<�$��y2j�w�"���ي�H����y2�I�f[4����fPf�j�c]�y��2$��tyRÐ/XZke,��yB��*p��iK�A(M�d%��y�Ǝ�F_�Yc�m�-�x9!�ґ�y��G
�8ZG���Z�ha*��y���q}`�s�]0^M^��U�G��yb��U=� �șOr�� �'�3�y��TTc\�J��ËE��t0TgO��y�#V�~��1��Í6���-�yR��y�TT�3�.0L�*�ŝ�yR�T�G���6�����i8�fA"�y�	��XgT-�%��O�����[��y2��:94���D�%wfrx+����y�-F
.ߨy(v�G�q��AG��y�k�4T��Q���e�֝�qo׵�y��0d�H��O�R) ���"�y�%�4B�5�s!���k���y�-��>&(�[w옳d�Ѱ��y"��U�q����,Y��P�����y��"�����N-K3�y�h��4�`���ńKf�R��+�y��xx�J琴�j�)A!�:�Py�,f}R��OܹU�h!�U&�[�<AF&�)� �{QfF2):��3%c�T�<A)UFv��7O�4���UR�<��S�%��y��֫P_&�ɦ`�F��(ڦiخ�N}�@fB^�5�Щ"@�4��gH<ɴ�< g�H�I<-��АM.�k��tΘ$1ј�>]�F�[����Ī�ݠ�x�O?D��	"�M.s�Xi+��+T�@�S�M�`���0���v0�H�F�i���G�,OT�Q�8v��	p�*� [d�P&"O��ćdbIЁޟ4�8� �(K����B"��D���Kw��)�p<� ����&:(���&�Y:AG�݀ �'�LY�$��cXnA���7v��T�n�+N䮅�,�6�y�A\e(<����	����Ap����J̓������i���r�I ,�
�>��o�zM����MG�p�X$�5�"D�� n"Gz�=j4�;kI|`i�,`�!p��̓�h����1?�|������.%f�69`,M-5�"��$��b�<��i����#p%	lѮ��c'�@��ZRX�\K��^�A�>��N3?��OB4CJ�o�u IH"TD��'��E�@P%UD9
�Y("�^MK"N�3�j��K�04 &�Ŕdb�2ס��=�Rj�%V�x`	�J�i�VHƪ�H�'�FQ+1�����z�m�+ %a��?��gH�l��(a3I�:E��"e#D���eE��G�:Ⱥ���Pƨq��}ӬI���N'�>���n�<�!�(�k,��,ܙp�pWZ@��U�F�!�؈ ��%1�ע2o��cu��s���
��N�,(��W��:�W?�p��d��"�Q �f1E���K�C��1�a}�D�2[��l��K5'�r�J��,An��nF%i��Qq�"G�D��0��A��L���+/j���3��?E��ҭ;ғ.]&�
P�7u�p�����b�������%!]�|�}r�Ñ1(����p"Ot9kgr��QVCS*�h<#�i��m��J<|JjiH+�'���p�S��5��Wm(E�� �`�j�奋)�yb Șx���mn�j!a��^�����0�R�26�P8��Q?�s����g�D���̡_,*��R��+Ea}��?
ѳ���GU�Xbb,EFh|��o>7�]sP��fFRec`��W���3	�9i��bK��6%cw*ғs��� ꌔERN	��␟�����)S,7/��d��DW��HRw"O֕c��0�nţ�d��2�ű���_�/aV=��@mS\$eM��S�I�2	���*W����Ԉ��תo��C�	  "$��c:��,�E![/;�^�(R(�&�qš�����%§���	�B�� ���.���j�,�BB䉵l*:I �� �؄"U�\9����@2�	pŀ]ΔA�鍕,�Q�8ʑ"K)i��;£ٍHR���E�-LO����Vi��ݠ��A�T��h���P$�Qҡ�{6���N�Fx��2��<�
���p���@V��<q��� �V��W��!_�09X������O�����[@�t9��<O�� 
�'��qR���KXJ����;l���8g��8���D�j<�����ة��'��ѐS�I$\�i������'R(� CU�t�l ˵�ߐ�|�[�L�TtI������×��R)D}�L2U���d�6��Ht�_��0=1S��"[Qn%����l���@�Ğ�Z�09�dT>��d�7�M)��8�A#�O��c�	�v'�1i`�i�Nēq��7)XNőu�M�xv��is��FfJ?�1w �6d �EՆ$e�屡�.D��{�*@�.�������A^�D#��-U�V�(xZ��m�O�"|�BF���2G��C0mJ�҂Db�ii@=D��a���uҲ��q�NR�FD�1x��)���:C�B���a@Lc�'�p-�B%H�s��1V���J�����'K�!�U�Q�P_�lb"@�� � d�%D��I%,�~$�"�G�V�tqs�M;6�`��D��x-�<�N>a��4*3�s��MqU:XA1��c�<	� ����}Hu�ߋ'����e�ɟW��9���鍟]=��c��2U=�dsb$�"q���3�|�N�&�&���r�Y�.	U:�8���!�	��ұ�M@��*D)��tk�Ze�R��dE7:��͓Q.��p�%O#uFFT���i�*��}#��bME�mW��!4H�U��%ԎN`VT��DȄT�:x@wA�)Wdp�*���: t��W���(����5�h)��BO'Oh.�sa����1�|J��1j� �P'�C�N��A�#\�� �O�"�i��B	CL�u�s�
4fԢL��d�/묵3��G}w�AaB%�]��I�4�#��>�jأm�dQ$�ѻN�yR�he�'�@-;4�Z�(�T:�����#�ʨ�4�U�^�~䢠K�+���8��(������_J:��P����Ԍ��)N,��0a��-{6��
�r��D"���S��.�=s�ܱa/��w�T�)A�_�g����H(xĮ���üRd�D���13*��s�<'vࢢd�1��\Q��+�Mc��X\�r MŬK��U!�� �^͂�E�g��ͻ	��c(@�Ԅ`O�s����ɻ]YmP5�	.�(!��J��0.����^*�aƁ)e4�I��P1{��K�
,�8!�TJ����Y��0��<\Đ
ْD���"�)�$Y����R[2�I0WX�3� �P&+��<%4�Jp`�(X��D�p�r��UNK�dǖ��#�X�O7��?�gNM�\s��J�9�$ �<����7SҸ�P�L
�!��?Q��#�bY�% �ÌX>�i1�G�Q�<�{ЇT>{�v�k�kA�V����Q���$�@Ǚ{4�EO<w�՘ ki��x��$D4$<&�<�ϰ$C�z��$��&��NG:� �0��`��	!�N̯3�a~��֛]2��y���<Z��"�E7r�v��� 3"���c�"�Pu!Ca� -q�1%��>����D��S衐�S=}�Z�`Df[)<!�D�Φ�2�j��c�*yZ����1��}Y5j�O��8 ���%�x��ɷ#���$ýߖ�3ɋ����sP"�Dџ|YRn�Ħ������V�.Ib�O�+�bx�g�;�8��	ގl�hCF"��?��" �-,0���.X�=�1kˇ����/}Xt��퉮�.у�� �+uHT�V���`\!�HL���:�z�k���y�Ǟ�"3p�B�Î)m��D 7Y����j��p������Kv[���L|2��εHd�!�'�����A�}0�����F)z֦�����(��X�W�2%Ćb�Ū�fL.̞zu��PMj�O�>��� D�Hb�'��\S�L�&����Ɇf�������$������YE65�`$w�	S�\�p�CE���~��<;&Ŏ�5}ܕ�@�'$H�J�$	nu�b�c̞%"�'�8!Kt�TS�$9R$~$������x����BV)s�<�`Q)�� Y!��vk,�@�*�2���h7bZ�oS�W�����fԔ&_�f�[�V��?���M�UԔȢs���Q
��CX؞Г6B>6V u
'i��L�V��&�4X������9z��}p�fޟL��!_�{2�X%�hP!�ȺYH@B����'�HA@��#U�4Sv�5R����<�$U_��8a�ݵ�x��cA�g�B��4>�&��شa�L`�� C�D@L�`���L"��2�H(O��Mk:���u%8S���TDĊ�O�yYuE�{��b�)	7r��E�����Y�d\�B��џ�@��>�O8�r�� CC�Q���` *5�'ÎP���7 �!(1�C;
}�$'��,C���6�F�xԚ����?�6��+.�l��AȚ��΀,g�(��x]1O�)��
,8� P���Nay��gy��*L����P�'l�q�LE-W�����[�^�{�>:��DI�A��L�q啝����S�qϔ�O1�Л�w����I׭8[��`5˥/�����g�>�اh�~�ٲ+�M^K�`�*LreX �>!�$Ѭ
�ȴ�/�v�����˟�$�Ȑ���Pa�P�E94���9w�:}r�݉v`���<�r�ͩ6ఠkw��Y�\|���ˤP��MrU�O+<i9�d��3	��M��E����4'�qGz⍚1��m�
"y����c��9�j���RU̓y4j���B�l!� ��	,l�湦OB7��c�8��H�� ���"�x@;���|��D��^
�@R��ב]�hhK�N��N��u� �z�ᄖ���	H?�'4��λ�t�	S��3N��T�ï�p�,��.ԎQ2U���@^�0�"�G"�>Q�#�H�d��+�$	�[ ��c�MįbĄ|�rO6}�JFE��!bZ��`QĖ��ɶ VE��}�%�Ѡ��j[>��)�ԍÛ ��<�OåxЦ���ڔ]8�V�ٳ(p4]�eJ���#=iqlK�*��IjG�
e�r!G_�[AD�!�,�ɍ`"��SN"���4��A��%�2�����ƶ	����:�XZ����0NN�E�����gs�m4 	�^:��s
_7&�~9y2�	�-%��''�ta�w�x4AU@G�b���u � z3�1"�'2*�P��&�)�'�p:��]�x�`yc棂=|X�O�����W%W�z7m�a�mi�&.��O�)�'~����ʰD
�>I���1D�O���pA%���:6Xf���D�\�	ۄA�k���ی"P\�ʐCa0ibs�.�2_��G0C�(9��_>U�IK%�\��㞤T&U�	��'��H%���祅�&�YG��1��`�t���5�k�����"§�	�����sV�0���6������ɩk�l��O�p��#�D-	W��p"��w��|"��O����Q�����I��th.���:o&@����0���� 	�͸G�޻I�D��>	`l��������'%�9��"�4u9

 ��J�h��K�4h� ],���hǧ�0�ا�ɛ�2'r���@�*���Iǉ�)�	k�"*����,,O�],y���+g'ā�U%D�8�T�{�L�13���I�}���/θ'���ff� ~�l��kY;F?Tػ�'E������U@��f�8�b�'�>�B�`��4KP��?�}���34$�s��2(� �%fq8�,H����~r���qp�(��m(��&��'�Ҥ#��'��W(��G;BeC5hA|7� ���d���F��/Y &��@*�-
nY��D\u��% �O� L�b7d@�E@\ՂQ�M�X?�x�S�i�,�4)��~2�G_���YS%?D���T`F�h�ȓ'F}��M�,�u(�(�Ext�ȓ9&Aҧ�Y&)d<Ї���tt ���*����y��q���?\|a��,�l��i�nS��Y�`=�P��P{�e�rn�5���dER�3�`�� �!�bF�.�q21n�O
���-��l��kK��l:���N�6��ȓ.��ݫ �wu~���ԏz،d��x:�)�$ܨ_����5E�GT�1�ȓ6nz4��d�3+�<yU��%@�X��43и�G$�	9�*uKBo TTn]�ȓ)$�J�P���b��$S�&���?��P�Ѩ��$��83C�EAm��B$�}a�/��/D|h'�[�ұ�ȓs�(��T�a'�XK�5ɖ5��.w|�ڂ�: .4@��HZ4�pm��d���CU/� `r���SB��z%�ȓ<� T���b���k�AƾC ����a��Z% (Qk-�j�(Q��F^�8s�ʾs B[���N!���ȓ�(��%^�;���B����7�Z���~e<�V���;�n�J�%�:X�ȓV���'�ȵr��)2���4,��ȓL�0��Y<	A6�B`ElE2�2D����.�LK�iS��<G�ѷ�;D���Q���C�ڀ�eE�W�ơ��+<D�����3;��5�&B�)�eؤ7D�xI��W��-Q��]�Zw6��G�4D�(ʳn�D^Vlk����-*���,8D��"��xj��a�ܣvm�Ѩ��0D�,��nL�?�:A��[�<J��)D�TR7G<n��`c��]�
)���;D���eʗ.6�>��@��hŪ`1�O9D�ȳ���	a:*�[ �C�'~H���j8D����
Ц��#w�,-XD��"D��&X,Z�����'.�0tP �2D����Vc�j����M�O�*xؔC2D���#��L��	w�ߒbT2[./D�2�ձ<Bxa��^�&4ԙ�f8D����!f��P��o��h��*D�H�!��,W�Y�w�B�k�A�*D���𧚾�p	s�`��><ƙ�4 'D�I1	T>�f��GȎ�d�����1D�L�Əۇ]���.i\�lz��߅~�!��Ү<d<�wf̛fD���D�4�Py�`M ,�!� �iV����j��yrb%xQ�&���b�B)r!/߽�y2��<x�F�!pJ�"��F��y�J�,>���l�pBʽ8�)��y�L�7)&����,ٽ���y� ��y_�)h�x��'�%�����$¨�yB��tUt��Gڪ
�R=Z�_��y�"Q#�������Ţ�C�yr�(�n�X&��)R�J�I�3�y2��)M����-��"j��BV��yb��:���8)#M������'�������+�OӸ;H�X�'ר���E�,%��-v�:t�N�<Y�"��=!Rpk�m��,�8JGiH�<)�o�Dݸ(��K�}���a���D�<�w	��
� ��dF�缵���E�<YVǜ�%y����m��i�
<A�Z~�<� &�(U�ۦ7 *���훅?W�T�S"O�<����8;�
�R��	NI8aK"Ò�P͞�KCBu���L@�UA�"O,����e�����ǀ@-<9���(|O^}�b��q��a��dP�oFT��"O�1����+|Z0��-��2g���Q"O@=����
���p+N�~lNU8G"OVI��*%�����  /�@8iv"OZ!s��	ƕ�s�D�]Dx��8Oz�=E����/M�L� ��|'L����	�yr��m���$�Z/t��l���W��y��Ʃ.m�y3F�oh�L*���y�I§Y�*��1Kb��x����Pyr&�G vp��G�$�y+2�<Q�].�! �1e�Ts6��`�<a�����B�#��0����E*S[�<	�FF=`��0�ЮЪ���1hT�<�cWf����q ��<�F�{�*�G�<����$h�TH���nU\�0���D�<���(F�h̛b��L�ν됪�G�<�rLN�=��и�CB]NmR�D�<�����f(3�bU����'k	D�<)qh�9���`�A�k�4�� �B�<A @�s/:�x� ]�>�����{�<�i�U�bM8cb���NT���w�<���X�mV u�
0Vh�=ɷƓp�<�毝�[�^P`���s���h#�Ul�<1��_}�4��� jźN�g�<��&v�
i;T�6P\����m�H�<ɲ�
R�􁙤l�4>���Ȓh�A�<�bmS8�(	�I�O������B�<Y*ٳ
�&�!SA޽'� � ��@�<yTB�, ��\�W��7QA�肱!w�<�V�ʨ�ȴ��.'����&��\�<�T쏓)�,�h$�B���HVdY�<1�aW�}r����b2~e����W�<��OC
~�`xiDڛkX�髣dGR�<1�I�	v&��oF�*����ëTv�<!�K��~Ȅ�#q���D �ђ5`K�<qGa>h��D#�f�H$��%\J�<��c�$fh.9�� ��"r��L�<��LT�r�>��t���^L�<&ߦ^�<@�F�Îj�T���K�<��#�1���A�y��Az��]�<�щڞ	]Č��-�By1��@�<yr&H�&z@9S�ǅK���p�UX�<	��U�#sʑZ�lHWo�(��Q@�<�]"3��2p$�7�NȠ��@�<�Ro�<lDÔ+��c�84Zp�[V�<y�aB���� �,�ҭr��T�<���_�z��h��
�i�v�$�L�<�v�[�qixy{p.�}�j9�A�c�<qc�T�`Gt��"&�#i~ A�z�<Ѧj<FX����`��`~��H%�Y[�<y7�\���T�MP�\����Eb�<�+�:$@�!f���iT:| !��t�<��tT�qdHa�L�S��U�<q�ě�5��D׌84]����jW!��qKh`���w�H����	�!�J�B�C�Gє�8D�-b�!�Đ������G�"B'R-Pb�17�!����p�7���	���� �0U|!�ĈT�\�P�͚A
ęx�� [F!�DY/JV��S�V1��6�P�e�2B�)� FE҅�А{�.���F|Ur`�r"Ori��� �\�
���8�^�;e"O�;g��<u��� ��U��Q�"O�� sG�&Da���piS���-Q�"OpLs�5D��m��gT?b�1Z�"O��D�+����DF�x4�4��"O>�p���4�r�Y��[%-�6n7D�<y�Ax�۵ �dd[h7D��@�!C6��(�׭}9>[I#D�\i�%>����N*� �#%?D�� �(	�-A�(�oљm.�c��On�=E��d��H�Rr'�xP�����?z!�d��@D�4���gQ:�!��L�$#���I�D��兜'�!�ڵc��8�K��`��{�N7uZ!򄛐O�r���ω�e�2�{�mOxg!�$^?<�֐��*P��a+T���*�!�D]$<��DI@���,�z�y�(�=�!���߰}��)R�.���aHŰQ!�$^�-����f[�@�D�����
Z@!��O��X�BJ	+-�Vu���Ȋ8!�$�"�D�bjG�N�R��B3�!�D�-\��@f�ƥ1�xL(���?f!��
Q�Dl��Ȁ�0P(5A*Me!�Md�)Ӂ��Q��b޶+G!�^12��%�&o��@���+]N+!��-��q�!��c�n0s����~'!�DQ�gT�A��p�)q�	
�2!��ի7L�eb��͘oY�(��ƒ�b!��V2��l�񥉏g&֭[��ƟSM!�N�H&\l���@u �8Q���d6!�$Z�Vc���a��G�e85$�p!�B^� �� ۷7�����!�D1J�P�� %a�����k�!��Z /���D�:1�P��d�:�!��:YMεe菋��ڇIQ��!�y�R�'nP�Nؼx@�E�LL!�U5Gw�U�ƅ��3�����'+!� "A��5	�ဴ_6���	$�!��]Ƣ���CY-mO^"" ��!�$�p��m��@n��Xp7i�!�D�/��q¡��$%Xv��o�?{�!�d�
?q�P�%�XE,�y���`�!��Zi��	w��;3�LPN��e�!�DFx�<mB6蟇<<��R�0,M!�$�<$��6#[5	�@�E�/!���W\���D1� �rs$]#!��\�X~�P�1��4��"��!�dJ2�Ze3�E�k��͋�"?~�!�DˉN�0��S�M�:Ҿ\p���q!�D�v���@b˙o������2o!�D��k�B�3mI"�8��ǄWj!�d&�\�9q��^pp�c�	 j]!�D�#�t�ǣ�7dc�+/�K!�䙧1T"�GITQTY�T�V;a"�O|�)� �f� fA�X��Yu"O��A	6m�����|����"O�,JN\_o�d��o��|�,�W"O��X��kS"�z��ӆ4{�%�D"O��R.�e���brU�g�Z�6"OƘ�e4"]��"-צc8�PG"O�)R�ʘ�{gY;�l�0w���g"OJ 薭��NY�\�P�M�!�(���"O� ����	��܋@�١�&Q:E"O� ��K&KУ=�8�H�N�tL3�"O���"�6 7ִ��G��p�p;�"O�(Kp�#<���(�_Z`Ÿ�"O��	X�e���R+��g#�iH`"O>�a�#���0���Jt('"O<�b!QL�D�&�k�`T@"Ov�sj!Uj��Y��"��7"On�iD�ُd�X};v�H�=~�5q�"O6�Bp�dB
,��!Y0Pĸ\�s"O���CxbЀA2^�� �q"O��@	Ǽǘ�pmO�F��Z�"O�8�'O�nZ��a�ˋ�w4����"O�Xj��U�|L����w��k�"O�5�	HNf���#T D)��"Op�@g	S�B)Y������	1"O,<Z�UB?칑p��< ���E"OB`H���1�p��
L���"O�a���9W�P0�Ɛq���Ir"Op��$�15t�QT����"O�p{��b��a7�σ)0�8Qu"O����JL��hH:�� ��"O��#�˶'m���Ƿf���V"O,�z��_�\���'�d���"O�%kX=��z�&�
�p=��"O.Q���_ $�D����ۂͨH�$"O�Mڒ�"H\r�x�C��D��5�1"O<�����8�!`#["jP��"O8$KCN�9g���L��y�"O��K�W�-D ����� ���2"O~�
��ʶy� �+�h��X5���@"OHD��A"=^�0@v���(�"O�%�6=��ٲtϊ#h*�B�"OT���.��c\�9�7���A��y�"*O6]��	?v]���H�|���3	�'�P�A�_�6MX�\�+N����'iE�j�U9�l�n���D�J�'6XtUE�fZt�2G�"/���
�'�$���A�7�ᘁ
�������'�Ȃ��B6\c��;DG� ����'v�f���t��t�I�r4��	�'/��"��N�L]��Ԩg]F��'v���$ek*5"��R;�D�'^���mߤ<
��@7����'J�� Q{RT�����0x��' �0��n�)Q�p���ɸH�����'P�`ғ�Еvռ�1)[��B�'���I��Ĉ-��5�qj�]:��	�'a�}AUBf�QF	�iW
H�	�'�.�Q@"\]T�����ȈP��d
�'�lc��_�`*�#V# ��	�'�
���C׆
f�2TR;j����'�E�rb��XUDKc�Z�i��e�'&�����
-?m*h��>]�0��'���*vXyy3�Y�0Ȏ�¥��<)�����Y��fk�H��'[A�<A%���7K�e �K�EÀ�c��<�e`u뚔9P䕐n`|�7�SD�<AbH�v^:�A7�&{."�h�}�<�'D� �8 (1E��{A���/C�<�G��d����ጟit�1��z�<�
Xd�ؤ� M��}a�ՈeXz�<y�K�T�WH޿)��D	��Kv�<A� F��d�
�:��� �.o�<�T����9�3	�(�ʵp�h�<� �݊���<7��YR�?���"O^�;u�5<�A��A�C-Z9�"O2�������^�`�"O��#u׏l�bݱdΔ��|�e"O�`�Ø$%��p��31�P
�"O&��'�ٮ:�����;q<��à"OV`��ȃ�����G��!"OX�f�Q���9�6��_��"Odi۶�Ƶц��t�֝f�Pq"O0�( ��!p*��iP6?~���B"O�����R�����	�eF���"O����l�:�y�FG�OO:`��"OBL�G��kG�`��Gޗ)9(RU"OJ�Xw�N'fB�9�L�4
v���"O���A�ɀ/a,@����9�2<6"O��uI_�9�0�2e%C��Hta3"O���C��_  T�Gk��`�2���"O& � *D/G&)rB�qJ��s�&D��a�ʧe����!B��aOB1�7E(D���ً��tSov6�ǯ$D�,�`��il���ϙ X]+�c/D�x-)ty��/�4Y}�����wI!�$ʒ`��!;�Ȁkv���h�4p�!�D��r���Έ��ͱ0�M�
�!��}�����"C�
�X�Z�C�-�!��8~�z���aܑ��|�F֙�!�dD#,h�p!�V�Q�V]�����!�9msx�k�Zc���T� !�DW0�����c�F���O�S�!򤛎7�����f�6Mn�q5�K�i[!���EϺ�#�e�1uW�B�U�(!�d�+Y����JNB*� f�(!�Di���TG@�h�&N�&�!�V:uT|�Za�W
%��"��!�EyM��o�{���R�Ď.W�!�$��)�
|�Ձ8�2T�DL�u�!�$�<�&�P��b��R�BB.�!�DS7+��c�*��%�E�Z�2�!�$�2�1JT�͹v�$����9!�d6y����9!��r��K!�M6�mq"T�s�,q��0.!���?.��ik̈́W�@�)��޶S@!��/m(�$�M�@I޸���:f!�d��/��B���A<�1����!��e�L�	�OTFJU�[�@�!�$H/i�6�s�L�X7|�	1NݍQ@!�>U�̺V�;>=(����*6!�ؒ��]�dk�]9�e�a�&!�$�+)�i
1�Z���V�V!�Y&i'0�hV#G%
n�5�4$׉=!��M%��H���{Zb��$ʀ}�!�$P�B �Ci��%Ex�Q��-	[!�dQ�y <yI�R#w1\if`O !���,-�� �s@�-#,&�"��	:�!�d��x9�ER).P[�/T1�!�]-7T(;�j��9^����/i�!��<����C�w*fL����&yp!��kv T����wv(�ԍݩsW!�J�<>�;%�T�,�媴�VGZ!��ef�2AG+�P��ỉE@!�d��<8b)� j�6Q���b6!��6��cO�^�r���,��v�!�dɡRD�9���%�v]�􈀸[�!���.1&D�� حR�pmb��܇=�!�� X���H�S��P'.;p�<x�"O�2'G�Qo�cs嚞D[�{p"O���Y��F@hS^�*�"O�����E�(��=8F���<�"OT�� U��)C�#�{唨pV"O����\�+���Bh�+=��}��"O��0.�N���JD����)�$"O�,�"H8+�	��	I2%���#"O��@��D�b z8�r)�7&*��S�"O��P�O7DY���qB\��0�C0"O�!Sk`����a�7��0��"Of�b#��.��8� S�'�=z�"OH8���H����n1h�1�"Ox�3�D� �:`g΢hV��"OY�އ+�歑��II�1�7"Ort���ޢk5��;��Ў3~0p�"O��֢U�=X�ȓ��� �y؆"O�L��N�=��#�����C"O�hy�)��%���G��$B(��"O�	gG�qf&�C`-��B�����"O�pS B�)h�U���X�3���G"Ov��$J�Eg�$��'}l�+�"OF�)�%ȞQ���2 ����g"OF�
�R�E��L�Џ�1l�D|��"O� 	E�y�Eʳ�$(�.��a"O��j֭Q�Ey�U���G9J��p[�"O�BD(M8s?�5�U�Ȼ.J��W"O>1�	�5��y)�(�
HS���"OL���6/Op�J@(ӍAr��"OƔs���p؎8�Sg�#�jUw"O��9e��]�$)r�4y�$��"O\=H�g�%BT&i�0oY�J��'"O ٷc�?Nsv�Pm߷3ȼ� "O�!��73�v�x5G�Y��"O��B�62�H��#�BGHIH�'�hܡ`��b`��-Q�Cv)
�'�|qP��Ĕ:+�D00�Їq�2�`�'�zE�C#˛J�E��+Gq�]c�'��1�C�*hH;q���|�[�'�v�J���N���Z�NĤ`;���'�X�u�M�N�P�A���f�b)�'�)M.B�00 c��<c�'ƠT����~sPk�Ѽ�~e��'O�d*U�u<�c-�$T(r�R�'�F,����;z+6��ɚu��]I�'(�$�a�Ũ1h�+�H�=i���k�'B��p�l� p$��(��iexջ�'�ư�v.���Ȭ��Øh�A	�'D�x���?jd���O�	�<��'w:48���+D����U��u��'A}Y(� �����H����0�'h� �m�9��4h�!�
�'Tf 8#�U�-���X���-����
�'JTd:V �9R$�Z� W�W�,K
�'�zP��#Ԯ���*�R��	�'Se ��E�,�!�c�:B2�!�'Yd�{���I��W*_55^p���'F������6"��@���#�=�	�'$-+T�N$4Z�颶�ձk`4��'��e�2K�b�� �\d�t�+�'�$���N�2���%�`2��'�6�P0�U:}7T�q'
;&��*�'dp���'�u��C� Y!�*��'�� �f�w������b��� �m��C]
�ic��n0L"OlЈ䮋�P�PH��A��8��p"O��¦��+����L�	��5 �"Oz�z���p��]z#�C�\���"ONT�&�<c4�]��C]�z"�!�D�=���1�եX�\(���!�Ċ�4��������!Ԧ�s�!�d�7=��%Qt&�d�1�D�2�!� %�>�K�\Q�.X�)˲j�!���Ua�JG(@X�5ɇc]S,!�B�\t�u���?B&a�C��Uq!���S���թ�� �mb�7iu!�䛄e��p+�>opɖ�ʊs!�$�@	�tHT�	�U�b�@��@]!���|��xY��=g `�j&�F>!!�䂵y�� �G�a��tqV�	&!�dڸr�LՆ]-~�ňD�x!�D�$0bF&C5L�:1{�iQ�!��4
f���GnՒ ���&�ʯb!�ė�zf�`7��q鲩J�J�V�!��I\�[���0W�R�*��Ƹ�!�$��L�� �7n `���:CS!�$��qDS ��,�fX���D	k5!�$X�:N4a�/I� �����Ɛ)3!�Ńh0lE�'�
E�*��f%M2@1!�$�;G�Q�:��LKd��<A!!���?L]���)�Ȝ�F�Q!�ċ>Km2��e��e�����N	~!򄂄i�^�p6J#.��dq�g߸ ��t��(�:\P�F���e	�*a���!"O�H�A�Wh��ДE�W@�т"O���A,ʝ���Y`��E
(�"Oj��oҋD��(�
TS)l��V"OQ����_��b�KI�	r"O�$��Tb���>Q��ڃ"O$�]�=�&�� �v�"`͂ b�)�'b$P�!@l�L���ǉ� I�$�'P�!戄:N�����).#@���'���/���b�I �����'��T3b�?YHn�)����,Z
�'`<��7c��t�`�P�/��Z�'Rz��g�����'B��4�I�'	��%�V�`�9+��$x�@B�'�:��C5+X�83�Ë{+�A�'�^���A6, ##�@�f3�]{�'�T p�AW�E�4�s2]����D4O>���٣f#t�	��I��"O�x�hI�O������E7
�"O<���cN�a�cе�`#�M!�dӓ @J��g��2P6���k�%�!�$sڠ1 �@�FN���+g�bO�X���Ld���S!߄a�:���"O��0������	k�J��^�dX��"O�(�%!f�$ԩ��l;�P�%"O��S��-�(`��`���"OL�� 0Nz�LSZ�8���<�y˘�iE��3T P��8�(�e^���d:�S�Ou(E2�:'�\d���A4V�)���xR��
;9�E�e玣x"�!KF6�yeZ���Ɋ�Hm�Te#���y��K@0	a�>e�6��w,���yB��A4ęw���l��j�ݻ�yR�ҖJ�YK!���vzͳ`Ǒ��yRڏ���� �c�(P�Ε����?Ɋ��� v�!�Q�r[�ԅ(,��%I4"O��@pE�N�,��&�R	i(�{F*O��2��2zr|���Q�߬���''������.[�1�SH�<��,z+O>���ǵo�X�Q�o��G�4� �Dٛ)�!��J�ɳ���uz�9����!�$�
r�=�TLX8cލ�F���3�R�'��O?ɡ��¾T�m����E
`���h�]�<!���s�(A:� �6h���m�2�yR�%/^d��q���.M"�'�"��O4"~�B��5̲���O�F1lm�uK�<�f���ubx�oH e`*�3q���y2�Y�ocV�3��o�4}A �y�c��;Lڬ"Ԫ0o5p�0Ņ��?���,ړ;������C�~Y�����\�j
�'�����D�u�B%�����
�'��0���
9$Z��[p͛�- ���'��Y�W&�"A�`*@'�z�\���'{���b<�98��M�H�a�'�$��sK։<��Y���$j~>��
�'ۂ����R9c�v}�u�+^���
�'��mF�Z�nJ�2I	�1��!�"O�L��`W&�ĠV
V:ieVx
�"ON�D�ҜI`��Ǘ�L<-��"O`tC���k�Ziൄ O-�M)"O���e�٧���z6�+g)�lB�"O�
��|�4�2�Z�8�Q"O����r ,����d�<�Q�"O~m�4KX���``��}�x	!�"O�[��5yF��7K-v��!�"O���Uǚx�)ٴ�D�(Ϻ�0a"O���`���9DH�UN�
W� �6"O�Y���'{h���D�<R��"O���dҫYd]z� �>@�Z"Oj�!�^�[l��-�f,؄36"O0x#�/�1cd���=j%ޡK�"O��Y��� ��2FdݍL����"O�@h#!R9"��-Hq�K�eQ�"O4�@A͠*P��S	H�����"Oz��Z�c8�m����-c����"O�y���b�v1� #v]�:$"O4,(2��	Y�����֬X�T��"O�1��)T�vpp��/�(D����"O��g挀#`U��Z�|8�D�"O �)G�_ Ev�]�K ����"O�*�M�x�b��j#`X:g"O�a��$&=�ȃT�Yg��̨�"O�P���Yg��,T�E�>q��"O�
�닒1?L�)�BC�̀P"O��%Gئ:�:Y�5c]�T0w"O�h����&^x�-��BU
AJ"OB�
GKT�;�d�%�� f/�G�<ѵ"V�X�� S�N�V�&I��+�~�<I�ɛ�b�^��a�A`��,b�
e�<��Y�:f��F�R/|>8�a��k�<i��$M\����O�p)����Q�<A�J/�@�`�<|'�i�/BO�<��'&D�|	tb�>>Q.%���U�<�$��K����%b04��a�Tl�<!`�������[�G���C3a_�<���B1
C����&�v(iR�^Y�<��c?B�q��F�0$�Y�<����@�4�b-Տ
�b��T��N�<!@�Q5[Zhɠ�N"	F`�v�U�<� �U�B�3B�z̩P��j)��{�"O��sJن|��EX5M��`$D�@�"O��a�/#~
D��]N�ʷ"ON�rvL�
Xpx6j� �"O�I�B�F�g�*(�'LN�"��"O���
!zyd��3�z\����V>m�sIߪ��H0��;iBr1A��2D�Ĺ��@�;���)6� ?5r���M1D��X��"��I�i��)�х-D���(4:��Z�#Y-��,�6J&D��Э�-���`�+D�l:�����#D�����@//!��oŨ:_4����"D�Ȉ�j.o|D�T�A,�d�%�.ړ�?��dV�B����&ک�<rF�	�(JB�I�!ؤ9a�J�w�.��̅�CV�C�ɌTPZ�{fFU�e0|��ߪ;�tC�(FЈ v@�!{��Y����t�
C�	��FEq�O�3Z̹���U��B�I�_����CCO���%�xSrB�I��|�ّ�)*�TMC5�;:Y^�?!����*(D%�e�Z�?�2�0,Se�!�$�'i��|HfZ{PT�B�ȸ=v!�$I��~hs�؎_^���G�!f!�Ā�X�	h���=U�١�]���e��(��ܠ"�Ʊr��E0eõ�t(�"O��B���o:I �$!��l��"O��Rnʯ�U';E��؀��'���4��Y��4�d͍*7�4��P�/D��H@b�&,�� A���T���#/D�p	��*"�xȐi�.w&}�,D� [��Ӫ@Xt���4�
%*G�>D�l�R�5��l��Y�v��؂�n7D�� �A�r�| �AY3R�8(f4D���Q���x"9�d�&MU� ���3D�(rb\�;)���S8K�D,�v�3D�`�P�J�06��O�0'>���/D����%̉8�`�;C���M#2pJe�.D��8#	
�#����4��L��� �,D�1�����[��^%z����)D�t���U�#�.��S��^�bY�B"'D�d���*#��0���9yT��'#D��HƊJ�#ʾ�HfPΒ�Ӷ@5D�,١�������-˯�.H
 d0D�@!0�*,.�� ��~d��Z�/D�ԣ�'��x�׬ܟ!���ע/T���'$=X�lB���R~�(�"O�U�@/F�pvj%� �=8N�(�"O0��E�,V$Pr�	�9U,�Uw"O�����M��f����C�_2�a"Ob=�n��9�"i@�	�;�TYg"Ob�M��?m�d
��;#� "O��4�-J��;W	T�g��� �"O�[�i��('�%�e�]7��"Oұ uGٌ+^�K#H[�3Ҫ�S�"O2��O�-1�x��c̣L��p"�|"�'�F��a���*LfPk��ÃP8ja���x�B�##� %(k��\�r�L�y��	��9+S��4��<0��ƾ�y��į@RE��O|O�+���y��4Y����%1p�ʉ��ޟ�y"R�`�����:d<:b0��'�y"�A�	b)AB�\14�@L��B=�y�Vze�X��8 2��-���!���'n�b$� ��	(Ā�i�1#��� $��R�]q�Hiu ''��"OA�'� 7�������(:�V\��"O�X�d͇"ӆ0�������|!�"O:��L-I��0��Et���"�"O&����M(Z���â�Tq�m��"O��b6ADZ����A�8Y��0��'f�ILi,)�B�V�Vg@պ���{fB�ɼ�\(e��:yT�@�Ġ-5PC�ɛ>�V|�J@%&f<��D�þS~DC�M+�-�W�:��#p��'@�B�0nAhmzfb_�,<�uR3�)�B�I�x2�a�1�W�|���PС�{˨��0?�a�O��N��ߪu���S��T�<�ć��.0� :GK�%K��R@�M�<�ÂB�~��0)W/^�XH��qU�I�<�2+�A	�O��Ct�i��H�<yEFF�x���sf�ŇJ<���b�G�<IwM���"�U?b��C�G�< )��>��`Z'ZD�nd�"�l�G�`����7�hIwA���p-y�'D��{�F�4i�`�$��I�l-2�%�D!�O���B̒&k��!��#�R30"O��ZvbPW�(�"���^�6��"ON�r3�F�e8���W"éE�����"O�y�Pf������9P䞑C�"Or�	DX�yb0�R�ȹM;
�*��|B�'_Lɠ6 �/�V��CX� �ݰ�'�r�Y�p�q�C���<���'g�l�Pe�=��a-�7���
�'fH��H�9`��(tj�.���X�'N
t��e�9t\|������
�'�B��Ʈ^Ț��)��6�+
�'ݬ�h��ɹ:��I�,�C�h�a(Of�=E���sZ��%�τ	�`���\��y�%K&C�(�y�L� 4�����<�y2�Ҏ#'��%��JX0O�5�B�.a������+(�ؤ�TĐ�N�@C䉌t��iq!�B"��C��l�LC䉠F=c���^��KʈF�C�)'`^`Q������G�EF�D�O �O��g�':p8��&�$|<�!l	)C2Ѩ�'r�R���qK����� �q��l��'s�Uk��$t�yt�zR4p{�'G�K��;G,Xt���T�'���'wR5�����1!���U&�i�'�f��PbȆQ=�\8�͊%�M�'s&!2����Y�^�۱L�-'x1����d�OF�S��{"Ђ)�dU�$,><(�� @�;�yB��f'F0?L�פˀ�y����jH��EM�)/}�y�v��=�y"�N9$َl�G�Y��	�n��y��w�R�(E*`���L͉�y�����҂��c����Ⱥ�y�i�:�J9��@Ǝ=�Zq�f���'�b�'���A��)��I�3cP�
�ɢ�'���u�X�.�4��gֲ7R�8��'�$՚��H�b!��E�'�v]�E�M������0�Z�'�zm)�M #S�[�%Q84� ��'Ŷ$� !R����B6���']�,yt�E�J����sl��7an���'i�\�TNľFzE�S��5�ft	/O���,Z���)wI�,T_����k��C�ɨ9�	���+h9�\���˓EҦB�)� �8P`�;;=���
�tHF+"Ob���Q�&�sdc�K*��J�"O,�8�=Xꅫ�"K`(>bq"OĕH1M�VDy㢠�,2#��^��D{��)��t|l���� �`ʢ�N�K�ў�������5,V:\�\�`�U��dC䉽�l$Iu�A���4� ��-�`C�	l��E�]��&�A,Q-�tB䉃[�:0٢IC�gD ���D;;�C䉪J�zeõ�
3k(�L�3;ҲC�I ��U ��T"�Wl
t0�C�I9S��I ��(E�0�ĜW:����q�P�'c.�8aGƲp�聁w�A!L���	*љ�" 4���a �uY�9�ȓW�Z��iՋmZ���@��(�ZQ��>e>�DhP=9��	b�(��9��n�2H2�C�A$���G�p�-�ȓJ��nI*3� `a��D-s&h��	@iJEۆ>P�Bē�|
���2�ɠ*�ƀ��MZ�2Q����zJ�B�I�9���!AQ/a��́��Xb��C�IC�N���$wp����O+�C�	�Zm � ��V�c>���$�߄\rB�I0� U
D/@!B}�i��Iû| NB�ɞkpNP3ɕk�J!�Q˅�*b�=I	�'d;޴CS+ַqDFp���#34�!�ȓ*�A�I��T�@�)��%Q&<��ȓs��]��S�K�֠�V�ݠGaH	��D#�Ar�
](�zd��V�q�TلȓD�TѸ�-��K%�%�&�	/\V���ȓk�x�C�K��˰�Y�� ��Q��l��I���պn�b���5o��5��NA��I��V�vڒm��E�<�jy�ȓaC.��G�s.Q�!F�#g(�ȓ}��i�bcJ�p� IG�Dm��U��xm�sa�-tٓ-�,9Ҝ��0��ܒ��:ܼy0���e��ȓM��j�C��lG~X�A�G!S<��}����'r��1�@��'S,X�ȓ��	�+Civ����#[3Fޒ���I͟��<����930�!*��`��b�<AV�S�T&����)�%g�D�c,�V�<�E]&��AA� �n������i�<��(�
*�Ԕpd��W�z�2�c�<م�����s�ʊV+d �roUF�<�'U=�4	�/�+�Z�����C�<	��_#:��K
_)	�v�z��B�<1H��0�{�O�E�Ԍ���c�<��T/iwx��3�]'GpȰB��\_�<Yw� PPN��׃W	^�Ґz��Q�<�pH�d$r�J�k���`��I�<Q�
?�&Qb1�S�W�Fm҇�k�<�A���LA��:=Z��B��m�<y��V8����2$7���3͛l�<����?����ɷ#�H,b��d�<Y�9�44��F�6����"l�b�<���1Z�Rb��*%��	�Ãd�<�A��E�`��I�(x���x�<�㡏�I^2���/j0�h���Z�<��-�r8��u�W$5� aF�Q�<i�F��Q�¨�6���S:T �6	�d�<Q4-�G��aia��/;��k�	H�<��S  TAa�#��XR
�3TK�}�<	�
F�{���=L~���D^�<� Ā�3��. h� w�Ѩc�Ұ[P"O�5�q��X���R�T����7"O|�7ES<NU \��ٱ۠�ss"O����

'\Ē�
G�) ��1"OH��-|�l�Z�(G�,-�1�"O���a�N�E�W�ג}��s�"Ov���D�uv i�@Π8.%"O��&ʢQF�!����t�d�P"O�tlֱb��u��YpK��y�,�.d�S��Z��������y���1j�$�`q�ͳ&��q ��
��yRa�0cL�I������P��ۈ�y�'�?o�@����վٰ�Z �y2�/`� �1akK�|4"�ؒf��y�m��r�v�!%'��m"�AJ�'�
�y�I'4&a�A]>SeZB�iT9�y�"�4��;S��BTv�y����y�ɜ?*�R�!���BeX�k����yf���� �ǝ:'��`��yү�B�QP���|�)��C�y�J��d��DÙs��9%���y2��I���0�҄i���2%�Q��y�+NB�d̢p9K�1
�S �y���+��l@�"�?ɂ0�QdǇ�y�aE�[�@X#��e����P���yҧI�M$e��ꂰXQ$�)��=�y¥�{Є��F�#Uk|B�'�*�y2��+
:�1���J)"�B���yÒ�<��}k�'K�G/��q��E��y��� ��ES C�\���\�y���%\�d0�@n��?v��be-�=�y��H\�ԯ�;��	V"�y��E1r�Ҍk'85^M��a���y�����f.�)�`�{3���yR��`�hi(ǧJ(x�l�.��y���q�x�#i~���"H��Y!��![wv����٧L�LEb5��#-!��;���+�FX/%��@2D��1:!�䉸�NPp�V�q�@��ܮr#!��ަ�N�"Ug�����jp�_�:!�d��.�ɠ0�b���tMO!�dQ<>8�IG��Gˊ�a��R!���f怄�sN��r���V�i�!�$�12�$pר�'9w��T�L�n�!��O7������;˴Y��ɪ(p!��1l�Z#Í<7U�����M�;m��џ��?E�aZ�'�b͘%bS�$�D�D%۬�yrEI#C�0肅�,Ed�"��œ�yߢ#p4� 4\8
�Y¤�5�yB��R�<��K�+�+b��O1�C�I98�ŒC��%r��#��]-g|�C�Ut�l� !�bq���޾��C�� �l�f$ �)RQ�\+b�C�I2�L-D�ܷ-��HI G�(	j�C��}����nC+A���t��O4*C�I�����Ώ�d��B��)8u\B�I�Z�ڸcv�
�Dmҷ#�^	6B�I�n�@�@7�#s8m�t#?��C䉞aFUX!	�i�L]���N�"��d�O��&�O�苦��VpB�眸m"a��"O�J���]�X�6�;}iƀ�"O�<;���L+ ��$+	HX�8��"O��rdl`W��	rM��Tɮ݅ȓl�d(b���-�ƨ!
v��T��S�? &ܩ�FS�G�T����?��ȡ"O��ct �F�S��L�f�g�'t�	C����L�H ��x�# �vM�H˰2D�|�怐j3��K�ΞD�h%2�O��NM�p:�o&8\a�-H�I���ȓc���#B/S� ���� Y�H=X��ȓ g2лt�ʥz�R�X�Ҏ_\��y��k@�X�
��t�g�G�%!6l��b�f���蕅M#d�1F���dz
��'���'��M�f�܅b4W�}>x���'}4)S��^W� ���(s�$�*	�'�ơ���;$,�Y�R1h1(�8�'�ztˬ84�G�C#f�t�'���ᓯT�'K���,Wl<��p�' ��%%ߟu ,l�&�Q�6�	�'�.A˵I�-3�h��Ȇ2�و�'�1��/O�8 ��T�ɑ%&��Q���?Olq2�8Ut%�R�-I��Z�"O6dѦm�� ���@�3i�S"O@����N���T��uT�`"O��iÔa��U�u�ߺG#R ��"Od�A��S�*pAE�rĂ�"O$hsE�1a{^�w��78��4
�"O�9�e�1J9y���e���x��'Jў"~�O�~�|���
�l��L?�y���-7��:�'2vq*+���y���A])�S.� @vܘ��M�&�y��o�Ε�D��n������yr-�*	�e����a�`!i�f�yR	�"��ђᄒ:n>�p�.I7�yRcN��p���iZ��r�N���)�S�O_МB\*r�j�㵬CLc܌c�'���(WML�#�� H6�ۇ=���'���Bc�^0b���f�~�Z���'�n]��y��<X��%�J�Q�'9�d��M��S |��4"�%�n0��'1�dcbZHq���ސx0��'����̘�)R\E�	�(	^|����?���i�60I$,�"LB&;��B̃�f�C��$9A�������-��\�i<j�C�	�s%4����pk�|�� JjC�	+X�bY��L�<U�����W�&9@C�I�{(�)� P��\ңL��4�C��w`�v`�'iv�PQqE�[4�=��'@��hADٝ��n�O�N��IU��Py��� %�@|م�'7T����0u��B�I.5C�+�7V����Y�s3z�O�����ZHr���!{���"O�=!!�Dп}�*	 p'� ��ȵ�B�H!�$X�� ��n�L����*Z!��HX������FPx�ƶK!�D�N���4l�'D��v�[�4��'&�f��~h�cCh�� �a��0b����Of#~��@�/A��I�G�ɋz�.�se�{�<�����'�"l�bھe%�Ы�y�<����\4`kA.�<���y���~�<�'�p�JPzf��'��\��-H|�<��`��i��B'8"�erF �b�<�e�s_*�M�9����`�<�mٰu�xpr�֑\�}��F�<�wi�3\Z��X�Ɗrr@��'J�I�<���>&٠���Kщ���b-Q�'ha����D�!��N�:��  �]��y"a�t$Z�ƌC�8�,԰�i��y
� ���2@U�	�hD����>c,Af"O�}h��
3 �L���eK<(U����"O�A+����O4��
�"WOJLi&��v�	O��A5*����M�/��Ih1�F�y�@)2�S�]~Tq���&�y��B:C��!�K�<�*F���y���'�� ��µ�R:��;�y��1���S L�|^�!�c���yR�[+0�$LcU#��c���5�y��,����lA*X����Q(�y�̝�l��U�шQ�9\r-Qq����y2k�'A���vfې5+&���g�y2�K��Yq��*�t����,�y�f\,
*k�'�
���%ؔ�y"�;k��!VK�o�b��G�ÿ�yR����	3�b��oq:At�]>��=A��?ɚ'�&�`W_i[���v���5Cܨ�'uP�C&.�I�H�犋&1;0�h�'��'cAK����F(.�.�
�'Pz�$�Űj�`�3��P�����'��D�f�/3�~�1�ۖD����'�lɛ����
��5%3D�r��
�'v��j�kT1ss*�ŮVH�ƕ`	����v�����
'�琴h�*�� �8D���T�O�k|�	�F���`��f`6D�ģ��M� Z���ױ`v�4L)D���f���] ϙ�|�n����%D�HP�b�ƕham���b�X`�-D���ď-9ʲ!3��9�R\k�6D������#)��P�%� a����WD:�In�'%�4O&H�ǟ/g�p�"3Y5��"O&�y���(ks��2F�
s:H���|B�)��"J�H�`C[1V��LХ�S<C�	j�F��RȈ�m�쬩�K:~1JB�	1
��\�����!�
�z���x�B䉫$�U(g� �[��U�r$��'� B��+�N 
3c�Y���)D�46��C�ɓL��]#�k�7p���4�
�=�ԓO��=�}�țk�<��f������Ɓ�s�<a�dY�%��сB�Y��ĚcZW�<� ,��t4 )��R�T��DRS�<��$�/v� �U̒wǶ�A獗M�<�Ł10��Pt��B��	�J�L�<���J:.8~��5@PW�h��`L�<����
�ڭr���'!^,QP��Ky�)ʧ3k�xSN�DY���}�h��00"EkR��,��Q�ċ�9R1�ȓ*�2<!0�Н1VP5)��B�-QE��6w�:�Ő�b���x �� �K4D�ۣ����+�#pV2��c�<D����߰x�J��7C�4u8��6D��5�d��c)Q.�EÃ�6D� ����:J�<�R�
�a������9D�L��=bM�@�'[�N\�4D����m_�-�$����,I��N.D�@���Rܤ��cC�V�(X��1D��P�o�%�5q��?*��u�0D��
4��1?.�&ٍG�p���&:D��i�i�cD�����N�J@"��;D��PQl�'xL�Gl[T�:����+D�H� D�?�,�k��ۑ5���T�*D��Q%�	.E��Q�W��;��ղ�A#D�Б�$H&v>� !��W��+EI,D��Ñ� ;Hxf�zR�� �t�"G�(D�� j@뵡߼~g$��!��$ 2��b"O\�Gɖ޼�sP��9�0�$"OC"�'b��K��T	���g"O�L�T	ĔBE�H`+��|"<�2"O�m����63,d(r)�n�,H� "O�ps ��G^J�hP��; t9��"O^��g%͸ ͤ���h�8cSV�)�"O����Z�R0ȣ���$��`ag"O`m���) �P�&�E${\x6"O��"f�� ��!3X>Ax��"O�I�4m��3�ӌD�ڔ�"O��� ��J2D�2)IE�<��"O�U�4�	����۱�Hـ7"OT��en�>=�N�;F_�Z�<�Y�"O���Ń&ZFn]���q�6���"O8�Ƀ��e��#a��[����"O.m1����g;�]C����|�{C"O�K��H�����S-O���Pr"O���)�:m��Ms�`�\�����"O&Q�/�8��@Y⮚�B�Z�YS"OZ�����g�q#�6z����"Ol0s��[S�8��,>'�|L`�"O��{gH66n��4�:\�(�A�"O~`rq�'!�̨Z��S�]�U�r"Oh�a싊HJpA�"�Dn�L��"O�+��K3MOPhQG�g��"O���A�q����f@XМ�v"O��SO�/|ސ�4��\�l%��"O�YUa�2g�Z� #K��&U��"OHL RB���R����g���q"O���T�)g���2�)�_��)�"O|%1 �3�L�h���~�����"O��yb۔B�>��lN��|aV"O4���Φ�|�x�j�j簔�G"O�h��J�g�<�����|��"O��P�o��[�8��H [�A"O��3�'J%?��8�5��1f]�Xqa"O���&ժ'�p@�C�/z~p�'"OzI�`�MZ�Y3P�@�#z�]�
�'�6pq7%� Bt�l����;���'�2��kT?��
WK۟;Q��'�����'�	~�6:��Z�A��� �'�43pd��d��<��-�N�Mi�'�੢�C�6>HXQ�ȷo�t@�
�'��,)�@1L'��PE��:g4*�P�'��uh�U#!iB0����z��'�!ץ����@c⁥a*����'� l��(H6{Ӽ��"m�7%�|���'l��@"#P4A��,B��jD�UZ�'i��T�ҝo�`���*��N,еi�':D�z4��H�C�W��5;�'>��P3b
o�L�AgO>^�%(
�'�)�p#�_�"��PfzE �V)(D����ٓTR�����f}c��&D�\�HH���p����6@� �p�%1D����GN�L$���p�Y�ڙQ0D���QiA4}�@�� _p�ٛ�l:D����K�&r~�hPr��.
���k-D����jݗ��Iq��{4�A���+D�H����dC2��ԋ(+�BІ?D��)(b�����R�
����"=D�`�	_73��yG9c������9D�d)�%�&0 B�"k�z�d���9D��إE�;�p��p�W#g�6�H��7D�� ������� �H��i��S�x5Y�"O�QG/ȸj��g(F���@W"OJ�r�ǔ �8L(J'c갺E"O��qCKD)��8!���Ia2��"O��R���[���$��#cT@hb"O�(���yD�ѡU(R��R"OR�7k��C���s��Ī\�)!"O"1�tE���"$�E�f&��!"O&<�¬�->���$H=[���"O����%!>b�(��v(���'w숈 ��	h~��7��E���'�nm"�	iy��:���(3<�)z�'������_�B*��h�lUY�M���yrb�+#D>ɢ��.
(��B�C��yǇ �z ��A�~bz���^4�yB ��U��	A��>Z D�dX �y��Jb�I��hŌm�ƙ9�O�<�yE�ߪ��@�ݠuz. �K� �y2�������	�Y�ͣbl��y�3�J�㔧��H��ay3Aˈ�y����4�����@L1� ��y�] R|8�F�65ƤH��M��y�oʻv�V� �d�<)D S� ɫ�y���RW������'��Ҵ�7�yR���M޾���*�������y�n)R,�ݱ��M$m���m��y�*��m�"��?	�2���ɛ�y��J,� z�$�)rb�j�"�y�/�^
��@�шh�n(r@@��ybn(�`��R�	�ru� ���yr+ҪJ�<�;i�&~�*�r�M���yR���3���qf�y2 uei#�y���,�0��g�	�z'���Q�y��8)��!�#!|�j�ߕ�y�E2����A��\qr֬���yrϜ�MOF]ɦ*Ƞ��6��y�_�%�<�E���*, ȕ�!�y��ڢqv S���}�
`t���y��=3a,q��O�D��Y3o�:�y�茝f�~� @�=JHx�d��yr� s�2��ԏI�	�(�wE��yңQ
	��st��
2�K��3�y"�8װи!��6i�/�y�ՄXP�ǅ�8wA04�D�2�y��/�F{��ֿt p!��-���y��r��\�Eဨ:e i`�4�y"l�%PBڙ"&!�';BSӊ��yRC�.� %�@%�0.� ��L��y��	% i�1�Q��F�y��I�ک�Ǣˋ&JHyR�y��Q�i_�A%F�u�4��l�y"�7~�l�Q���1�`�K-�y��2j���@�:r���w͏�y��?;�*�ʰɂ2r(lBkH�y���|����\=b��*��^�y2'�v�!�E�go�t�3#S�yb�����I�F�n�	����y��\���u�׫j� q�����yB�F�M�|�(N5jV�p���y��A�'�,�i���1T"je<C�I�/<x#E�]�=j��߸E��B�n�q�3O  6PSwS�B�	�@��A�Ď�6	��p��#[#B�I)lC���ŝO�M�振C\B�)� 4�;C�G�O �ySA�1l.�d�q"O��+��F�/=�Ț��.E<%"Ox�#�ܻWK�%CPĀ�c�	��"O����ʀ[�~dHd�����y
"O�i� �{止� �2s����"O�	둆ʖ�{%jμP��"O�谳j�<Y��)A)����"On�"!b�\����ƈ9��])�"O^R	.�HS �ŀ{5���f"OԜ��D��bP�Ϗ	w����"O�xp�]:@�͐�o!G:qj�"O�S����P�^��h�>x�\���"O�B3��H�xg��pYb��D"OT�@P���)nv$zT&� .J��7"O$0�1aQ�X�e�q=� ��"O �W��G�r12WgɹT��q"O�=�s�Q3���P&�*/� �"ODA�^�@������:�5�+B��y��\ V@��B����$柤�y2�D5f�zb��^����W�a�!��gG��6��xv�y�lR�E�!�D�+>�j���"GF�D�^7�!��Fz��wC�8b/����ʹ0!�$��(�I{U%e�q���T�?s!��t�0�PF�l\�{�hL�mq!�$��\E���Th���PeH�(!���yۨ�@tI����1�){!�Dˀtz����_�D�N01�m֮<h!򤝋0�Hy����9~c���U+Q/99!�D�3l ��2�R4D�i��M�u!��$&3z1��ǺT��R��3�!�$
�@.�x ��c\������!�d�n��Y1�K�xl�p��GO�!�C8d�(�[6�	&UW
հΔ��!�$\��� �CF8r"��i�K]z�!�["��qʃ��"(A�+����'F|;Iֈ:x� �^'a�6͙�'A��p���l�`P�DOͽ['�!��'�&��Q�o��d)���[H���'B�
�"��\'�lb�hٖS�j��'QNhqfW><�D8@�LSF�:=�M��m�W���0���z�;��
y��<�vc5�OP�n��1'ꅛ��x!#ςC��)r��d?�>��	ڂmx��cH�:e�J���d�b �O��N=?)c׍޵0p��%☄�`$x����4�=����O�20��6E��0�Qur� q�"�S��yr���6�7��rlh����y�aGw�"lsp�ԍ �r�k҄�	�y��ԛw=|(��$�mSh��iR��y�aI
�3$e�c4��#��D�y�
N�V4����Mړg,����՘޸'�ў��`k�	�,M����!k�S���:�"OD�� ���l���vI:V�&Ty�"OP�!�-$1�O�1-@���1�S��y��,_i�1�͵Ea���S��y�k�0�����.��)xg��y�@F���+�-9�yr��y��?](pu�7���'?`��E.Z-�HO<�=�O��y+vď�8h>�����7=Wv��	�'W�Y
'.
�BM"� :@�d]�	�'�����*�Y8��ӾdƬ�	�'<x�p���.;G�h�Al	ZP�Q�	��~��/3�I�vDJ?�P��$���y�`آ'kx	�ጟu9u���ך���hOq�� �)-ןԸ,AǊ� k��p"O��bG)�+( �hp���
@~� ��"O5sv�S/ad��qŐ|F`j��|B�'1�t:���<�4z�/�ʞ|I��$,OL0Ƌ�Id]��kO]4PY"Op%q�E�}�d}#���3�~��"OD�Re�	���s�iI0�B�x3R�tn�q���O�~��6ˊ$�������Y�j�'>4�V�s<��H�)UZ* �'�a�&w�:-��c�,W�ѩc)ݚ�y�,�+:]�dܿ"��&��y���l�B.X6����P-�y��"�����e�$���K�����yr��1~m ��m/����)J�M{M<鄧�>%?�O�Lcƿy�Ȕ��.�<��쀳
OT7���p��ubƥ�"1���Ɔ�i�qO�=%?	쏱!�p��DŘ-��02@/"�?�j"}���aV��4���Hu�R�Qz�<Qu���m��0H��DX4��3��y�I�A�Q���yҬ�1'����˺k�A+g����?yp���x�j��J&��г ғ:��!ʅ	>��M?�O>i+O��Bq��sd	�CI\09��#?с�0�u���o ��Dk�am*��&���M��'b�	a!�!��)E �hV<����O�b����$"�*��NqP�-Y��"ĤO����Q�a7Ѐ���,9��8r�����!�Řp�T��e��?v���bT�$�!��Vv��%�a$�{��HV���џ�F���͡�.i1��X�<d��1E����<aM>E���>P��1�B��A���C!C8�y��S5[om�"�reh� �B����-��Z~r-\�T�[җd/yM������8z�'-a|�n��Z[h)�7�S���1 �K��HO��=�Oޖ��w� .ol���i�oY4uh�'{Z�3���@ �� ��(I���7�S���)�x@H�Mv!���yb�&�|`i/�p^�P�1M�>ˡ��:j��&̇`&��13��2z�$)ғAU�&�D�=x�L��o�UL*���B-�'a|��J8�ra��?��ڐ甆��	Z���O�$yZ�+ǠA� !C!	!=�ĩ����'H�<b��pg�ɂ@�5<*���'�@�o؊�F��7��8�9�
�'8M���<�4L�P���
��y�� }�@���� �5��o6ў"~�%T6Dz# 
�^~�g˓&�t���H�-��kV`�ț�.�$�~e̓��?Q�ix��Q���HWz�7O�YB�I��Th�(U(e��X0���&k�BB�ɱv������]p+�	Wd��{��'�S�t�����O?�Z@�f&�	p�C�I�vl.�C�)Щ }���A�0ܠ#=�Ǔi�h}i�đ+_X� +Ҽt�ؘ �'�*Р��1�4�Bsi��j�Q�'�h�2Ǉ�,w��t�'NRq\Xb�'�NE���[V���'�!gG���	�'AШ`��D�Qj�7�}�a�(O�=E���1/�pؔ#F$e�p*T��y�ɺy�����ӇRmp%ɰ����'7ў�O��=��Tb⠨�n�v��8���yB�*�� rK�����DD��y���"��xBg�?b��C�Q���O��~j��՜����&��z^%p�Ok�<94.�(}�	��O=$����jy��)�g�? ���,�^�8�8�k]r6��s"Oؼ0�b��rr�J��uꤓ�"OV%�eOJ�Vd;��:@�(2�:,OE��X,{ʒe㇀&���5�q���'�<сm��<��R0��­ِ�'m�>@���m�: T�{����@���Ӏ��'N&���N9eʐ����@�����D'��>��݉ *C/8��0�a.��6��$�',b�)��	�l�2(@���l┬˝^X��� �	�W$fyk	����x�W��%�P����'x�A�.�&%����+C�D!)�'r�5�v�ͨ!����. c��D�ɦC��D����å���E��Y���~��OT� k��5��ɒ��osp�9�/�$t�5� �'�'m��*BF�=`�HY�&���-�8YT�b�@m�3z��OԒO)�� � :b��3��=��"OT�Y�E\�dPT�&ͯ�Y��74�P�3G^73����� ��R�M)��TӦ�ow?�*O?�I5}�a�/n��!�7#��	d�B�	fX�\caL�ꐋ���8I���~r�)�3����wœ>)
��U/�G�`��$�>���K
38���ҤG)YG�r�� �1�O���$��vb�2%��%�e�$�"w�!�7�(#`ϕ?ʹ;$�Ŵh�!��i�<۲�T�j�g�7!�D�
Zzu�BG�,ѼP!p(U8!��	�P9��Ƈ�(yc��6e�!�$�&G,�w��<y��x��� 7�!�E��D�r���`M�i����(|�!���$1y,�Z4EJ�T�O�]�!��(U�hz��� #�2Y)AoN1!��M�_L��`�CM1)���!�d��	��UZ��׺5Q��O��J�!�$��B0�1�$&1��B¨��$�!��0�HM�'C͐o����e�/�!�$�)I�d��,��u��M�E瀽!�dQ���2#h �b���	e�R�w�!���h'�L��;!�6!I�%čGI!���<H�݉��W�`�J�k�iȏ3C!�0>ND�8.:U;�i��<U!�B�'�$`+�n[�d��fնp.!�j��Q�g��]�s2�V!}1!�S�(y�e���46�xM��d��%$!�$
65�b {T#��	z����j�:7�!�J/C�B�y�$��3e e!ƮI� E!�$�!$݁C Î^L�X��Iq!��&"� ��C��$����	E�!���	а
��s�BT0b$O�!�$�4J���I2��!&�@ �Q=S�!�\fy�D1�ۊ,���"��!0!�D�Vx1Zp�31(|ܚw-�!�ޑ*�L�@DdC/)���!�ސU�<}��Y�����L%;�!����,���)���رfEk>!�DH�
QDaA֊Q�n,��gB�h7!�dN0k:��d��n<ɘR�^:C�!�D��f�8l���a`�������gja~2��2m*3���[5F1-m�V�h��4^pU���e�A�<���X2	Z����z,�%�r��) t��H_{�)��s�>����ҡ�"5�CϘj�E��dQ:Њ����R!ADo�,�8̆ȓ9�*���l�%1 =ᄊ�_��C��L���=[�Z��o�?��a��S�? @���dхp>^1��,�8V���T"O�+�KK�K4t�h@j��x�P�q"Oʨ�qN�$TwR���KϚr���9�"O�A��C�9N4�J�+��5�v"Opqʠ*ԛ5D�q ����.A�"Ot���,������9��@c�"O��1 �Θ�eȂ�w����G"O4�2&��) zL��h�w��bA"OX�HF\�E�Qza%Ž\y�pZ�"O�f��}׎I��$�	q�$)t"O��`�@N�#�0Jb$�4]���"O����. ��E1�d۶l<�p��"O8��g�!�N��pE�52�di�'�v��!ẻ&2cC�nv���'���ش@�&��0���%-�h�S
�'�r�R����##_�?pH��'V
]��ß�7Į�rI�8,��a1�'�H��L�ULzM6�Kq\��	�'�<QH%Q.�4@�@r��*�'{��Z�,@%B���	�Ӆx��b�'C�P�+\#'^���ݔp�u��'.N�{eS��᧩	 %����'��hw�F'h쬳eh���a�'�|�sFK��	�$A�+g�\��'/�a��`KT�����!�[c� k�'���s���?.mʀ�\�H�n���'�ْV,Ϩ&�� �4��(M%HU�'W4Es��]�|t4q�d�<X@M�'d|=�mM:{�(�J�H�$ժ���'�8��ʗel�������.�!��'�PS'�P���K��9Lt��'��P�ï��dR 0�0���j�ش��'��I���kaZ��Gʀ�\�L)�
�'ތd�K������I�6H�N���'��i�A��Ih)����C���C�'nR���A^S;��wR�G���:
�'����$'��������ܸ	�'?�ՓfB�3M~�b����:j��	�'���JGfU%_��ŻS�:G���
�'�pR�_,@_`��C���l��	�'*������6I|�Y�j�C��I�'��!!΃F��ay�җv�]�'��]��k��%��j oTb*$��'X�YUl*�v��_�ԞB�'�䩂N�u���{%-�'
����'�*���A�q2��T�%��``�'{e"�|��#�Q,
�h�!�'H��ů��lϼ���A�3�n��'�8I��c�MY�!�g$�'7v��H
�'��q���i�}#.�{���y2��F�0�@o����(5��y�.˙1�����P=��Y��A֚�y�L_i<��PǦ�	�D@�uk�yB��\�\D@�̟p�i��#��yB��gAyqB�6"7���7���y�@ͧ��u�`�#-��xD$ʔ�y҂ʂ\:X Fj͐��1r�أ�y���oTp�1�aR�?��a@��ξ�y��-	���lB�X�t��ԥ� �yB#O#���EI)Ur��4f��y�K��
���=H8��a����yG��0�65@d�6H�4 K��!�yD��RB� ޗH���$��y�<0��kA��0ހ���
=�y
� �0s )E�z��T ��G�l�BdK��'�P`�w(
EX�`��Ŗ.	�Ja��u�X)˧�/��[� :�-�<�{�l��?�%�Oa�*D���=��:�� 3��� �'��e&	Ε7e��2D)/����O��	�Fְj"Lu!u�O�A� ���1i`�N~��Nd�tx��M�P�l��C�W�<�$��L�(�.�|�@�]*O'$����Op��@�RA�	�б��ҕ����	3{�F	�d̝S�@�0f�>=����O8s��mJe�Ca0�:�ka���F/�)m�0�!&��-P�:�QP��n������	8	�t� 2�ێs#�y���E7���X��1q��X��I��JԳ@+� iv#[�c7���l�/�=�࢚�n�" h�#>��?� -�@��X���^&�h��Ɋ�� kL�8A�U��i,K�����N�B��L�$'���$e�탲OP:Rq�rH��n Ѱ��9D��6@E�7���[�N!sN�8in
H�s�'�0��'P�T���>4���sA`�#yV�t��V��84 ��Ɗ�Q�l��'����B%�0�Jq
�)����R (ā�p(���
	M��eɈ� �Z,`0*��[\���ϓ�:\���H+i�Ty��È�P�v��'D\Yۅ�i>�X����0H҂$��j�@U�ɂV�b�p/%f<@Њ�GM=~� SGFSM�q�C��	ya�	
.k���؄K}��'�S#d����FJˎL�*����H�{."
Vi�,o�����'��'���yw	��1�C2AΙq��IG@ٓ�p?I��'y�HBa ,������)I��¯���x��N�.n��2�$ڑ-�>IR1�*����V�@�M��b�s��pv��6��$h��H�jAY�0�e��Q���@;N����D��&8
�X6>6��!�$��ڸ��P,^
���� \M
չ0�J .$ ��B�?2��#>�E��%V0e�vFR�`֔e �@r?��i�6���������
	L�(�<a���2m�*�0 �'���k�O�EߎX*q"��&J(��W�p�,8a��(�O��r��D�~]����n��GZ�E�D|���ևN���ဠ�L��"t�ŗ
�je�D�?Y��wW�I�eb ���A�%��s����Y����T�VC�U$I���S`͑�8��ކG܎��!�<��ٱ�OB�]��
����M��󄊝\b���!�Vq�$Zj�,y�qO�(�6�iݍ�U��-zfA8�:*	� "aÙp�t*�`[F��2@� w(�Yg�Φ&�ԕA���{�'G�i&,1-ռ���@9΄q�fܓb̬�3g-�Y�&�ݎO $�I�FM�&�>�6,=9ߎ�Г�I~�)�l��lČ̣���J���`��&�ܴQ �A8a�1�P��U�c��� �
�#��"`D�ɑ2&�ؤypKA9`�!��hVHɰ@�,�󕈎(Q�jH��I!n��r�>��c��*��u�U2X�.��j� [9�L��_Z'T=��I��wP>��%��[�"���Z��3�)Y(N�r���#�~�;�!�	��h���4���� �8LV}R���!۠m��V���A�ŕ&G:�����'<�&h�c�P�%�Z1���2�!$/@�6L5��d;�*.X֎�����OZ AQ
��5V/١���੝�C��K���y����J��򣊣1�r����#����tn<�O��Yc�'A�Q3��!M`r�k�"O1bwk�7_��`�֟9���P"O�`��.�7t���t��iu�E#&"O�=��a�� ��8p�g�$|er���"O"�ZpDߙ+��|�4��\RM�"O~܈�Nۤ 48]���J#co0�3"Or0jD�Z���x`� (:!�W"O$��Dm9e�X�W�b����v"O�4�B���p��yD�;A�|A�0"O��qWbS�*n�9���c��2P"On9[��̡^^��aUG�;|���;d"O�:�V7I3"�aE��5�p1"OB�Ռ�[}l�[�ş�F�0"O���rBGt�����Y�?�0��e"O�x ��5^5�@%����,�H"O��� ��eӶ,��j�1_'��2�"O�5�#�2��\�"�[�$ =𓑟ԩ�R�H�z�е��A��[�Mb��
�eT3��>���)UC��ֈ9 T:E��HA����� ��y��B)@x���.E?W0F�B
��HO*��AT�#�D�[���@K�>�θ���]On�������y�	�%L�xё,�:F�6�0��K�M��i*0�b��>}���iofى4�E�<��y�c��^��4��'�F���,xT�9�͙������O�ԛ�LHjĂ�@ϓC`�e�Ս��t�Е��P�$
f$��I!dN �0�H�9�� T��G�LF���2���#Jμl�"
54�DI6�G3]�9�C��QY8%s4�4ғp��{#,H���?5���H*8ؙ�j�	sHH0R�'D�1gb�	b&:4HtmƬzDd�xe,e�H���Ņ��݈M��}:G"�O��R6��)B�uc��n��P��n;�|�sh��g`4���X;6��3 ��>	��ϖ[�ԩ���<9ԬL'<^f	[O>V�ѳG�l�HBc��"���W�qx��K�c9�1eV�xRv�[҇M�DVh�`�ChyB.	5�E�5K��)Jԛ*T�<���ha(�:J�">)�I�{�B�|*�j��␉��d|�&�՟��j�4��O���gܓ�P2!�
z�hb�݊)X@1����h'��"�JH#��"�z��慌p~�b�'m��z���X��Y[��yir�����1�QՀڂ|�����@�y�S�]!sC�
�!��xqg�+A#DB��&f� �"HN�@?�S��V,dB��R�/���1T��?c`�1�"�g?٤���0��8��/��A� գq.G�<�5 O�`;fmB3�N	&����	B=Z�,!փ�7��@�5�0̯{�'� �Sb��v�X�j�!ȋ?�H�X)8$)Q����M1���
�ڽ����7�C�@7i�@@�[؟�� ң:� �b���8Ӡ@1��-�I�*W���S�J��+�+J��OC��L�]{I���*8as�'�5+�<�x0�F�"8~��g.Z0%'D��S�W Rh� �۴0��>�zF�-q�ѫ/�8��L�7�\؇�_�L1��G]�(��=B� ڙI�|o�Dꘋ�E�0EJ�{�{�\�Th];#�(���J���=y'd\ _�p�e�OXd�J�����d��^3���"Ob�(e�I�wO�Y��"ɡ�dCt晰���h��I22��<Be��'���:H��"OƘ(�ȅ�Q�]0���B/&I�'�0�Vx%�|������%ZȪ�e�פJ0:�n,D�xK��J3e�>i����q�څ��y�0C���O�|�^�(��l6&��`��Ǟ(�yD�7����܅؀mr�Ȓ�yr��(�
���δ��i򤟉�y�^Ux�Y�ԢN�����@�E��y��M�������~8�J�'�3�y�����w��P8�7ț(�y2)Гl�q��7�����c2�y"�D9HD�Ҷj��0��t�S��y�!S�<�H E�Bv�*̂#�y�o�i䖱�����4�*��R��y��\:2�0P�@!�SC�͈�ybMO?��4+�A'X�{�i��y�
Z��>��K�4(90q��e�y�'\��y1�/��'���҃�:�y��ή�f�ӵ���V�@�Ŗ��yH�D�L����F��Ω�AgȌ�y ��"��Xc 
_P푃�N��y��hR�� ��4$ b���yr�X�Q2�
��J��l߇�y�hC$�+�m��K��0��yBHTsf ���Eب�d���y�3I���g	Y�Ƞ�Z�U��y����u�:� �kĦ	$��(�m��y2�� tڡpqʆ���T��yB��~��[�,J�)=�=X� ƻ�yr�
O+`}S�A��]�p4��G)�yBoK�a��r&n
�W:^�f%�yb��@��(��լO�ʠ"���yrL��Qk�EǪS�z�y���y��*+��z$MăkN��e���y�\ ���+��Q4�
�1���y���"p�:�����}%���F�Ȱ�y���E�tU�$N4iqĂ�b�1�y
� "Ax֦"K�85���W	z�T��"Ol�Q�C�P�hB��6$2�S"O�)�f�̕������țzN�T"O��ĮN:NЭʢnی��[�"O���	�7MH��1*�6��d�"O��)��ޗMIRH�	
$>�Z�R"O���F�t�ĨvG��"2���"O���/E��l�G g�L��"OV�x3���Q��u'�Lc8|��"OD�H2ə0d��H7�PA�Lx�'�8�k�g MJXx@@����	
�'�hqP�Nǅ@	��"l_��4��	�'D�!2�"���"X3$3
���'1�5k�o�V�ܸ��L֬Kv4)�'��]4@��2@Lp�'�(:����'a�H[d� ��Lȃ�;�
L��'����'Z/�!2K���PK�'RX��/�3_�U����#��9�	�'�����F҅&��i�C�+g�Ւ�'N�<
!��Ѐ�&�� ����'Y��!󨖥N/Pi�&��^����'��xU�Vy�h�F�ra����y®�>���҆�+e���b�gϗ�y��߹��0��%���`���2�ybI_�
,��)@�DU�fx���*�y¨��'�&��p�@O�|��ab��y� �(� �D̳1Qv]��IU�y��.?|�]s����6���9EO��y�%ާYe\Y��O�{��� �f���y� 5��@�㨃q2�@���)�y"�8p.X2%�i�z��5�#�y�A��2� �pHP���֫��y� �Wc��R�p����ŷ�yr`�_��T;�/�i٨l��FJ�Py��J
qצI��*u�'"OV�<�Ӯ�:82�
�,߄"��4va�S�<��Cר�J����)+�Z�pďDK�<AƮ��|�"�"�[�!�� �U/�D�<�gŉ>!X|��A��*jw�A�#o@�<!`���� jI�dJ0 Ðl[�<)d&kI6�f�Yz�gc�_�<qE���/�<M[���D;y��&�W�<�#�	;^�a��)�0e� ��1�P�<��ɏD��yWeZ�:�IT�H�<YU-Y�4��a랭@��4����G�<)'�+l1��)�FA�v��5a�LC�<)"��e!	[U�?x��-@�C�<�tJ<�l9�F�C�MdB��D+t�<�F ����$J�@��<�3Kt�<�@�:_��@��-k|�I�e�Mz�<��Ϟ8�FIB� [�I�]m�<G*E�)���0�ιG�8b��@�<� � '�` .�#Y�켘�T�<���_�P���UHL��h�i�<��L�^4������� MQb�h�<�@
�W�X�;�cT=C�|a��Jh�<��JǯO�����h�60+�yu��g�<ْJT��Re�vײz�>tГ��c�<�q@#d��iC!,{#ܸmPwj!�DX�:�{�R-�^X��ݥRv!�N�Vm*=kq� �v�b}!�4l!���vV�xS1eX9�$z�ǒ@[!��ȅ(��#c"M�@�,YӐ��:D!�$X~�B�0wJ��H��%c�60#!�� ���s�@�f�([Q8��"O�x1�dE<J���Æ�?W�8y��"O��RQ*&cԹKR-P#<��XK�"O��r�P�}pf�����4_��e�T"O,K*�x�� f�M� �є"Ov��#u{lQs&��8���(w��Q��U���h^���)2y�]��NE/L�!���8\?��#�&*j�+wJ�z�I7�Dy��y�)�'��i���>8yѵЎV��ȓ[���u#=�����	�rL�OZi�Ý���ÓJ�z�Ʌk�F\n$Y�`D�;w� ��I$�:����m�-����54��(��a�#� ��O�0('T�$�h�@��"r��d �CLQq �ΪdEZ��ю;�S�i
���&��,m�q��+mt�C��)w3�d{@ԇ �J��2A
3���ZgcH�VJUh)U�+&6M�_��������@��O����m�h�!�$���ɤ��= <�a`��7%ɒ�H��O��+��p#Ll{��'1��跈�	�<�g�����2�N��9� A5y�@��^�C]$�`�?a)��*W���Vz.�
�2�x(�i�\���5h�8*�P�v$A��l�Â�Nnb�����@:�Y!���uR��*:�1"ŏ�7N�͊G'N�3*���c8�O�p���K�L
� wkJC�Mh��M����Ks���9��&x�x��'����" �w>����e�;
����r����z(9�'S��z���
3�<�j�
}�>qsS�X�'��pа#	""�L��g75S��B"�9�(
�*D
|�:y[�'�e9g	�-D A�L�s�T��IԊC⥝7�C�E� �����2/f�(Z��T.�.<�@�^E* �2���tDŒa�á��#>�`m� ]f�	v�*=)��A~��J�P�߄iU
�BP��1p�^�)Q�m?�R`D�fܙ���	���k��c�Rd
v�\({�a~RG@/j|�ѣ�M8I#X|�Cۚ8q����8p̤Ô��-0�����-bp���;O)Vh�Zwj��]�a�2���@4<+:��
�	��B�I�v�!!��W��&G�
Ya<
�U�`� �P9ot��������)1��������	_k
�ɤ[Ȋ�������JA�,ۄ��/ќq�%,�.�Dcu�S*Nv0���M*�j�"��T3S�.��䆑OԴ���-�J#>�(';	*`PW��<"��!1 �L�'0�ZIO�̥8ROC	%j\<(�#�!"�|Mqt'�#�@9�%�h�*Q1%�Dp�(��'�����,�;b�h��/��iBD͹���>�s���$�f��f䔝����q��:c�b�0�o�Z��#��@�!�_�� ��FOƊ !�^�Er�8c��G4�¥��Nͩn��Ht�M�5�pa�]�ބڶP>����+snp�kZ���(�3�����E�^��IQUC(�O���q��G\l�	FA�6z��2$��6m��)�d�b�i�g�I�A�d��g�cu��-4y�L���D}2Y:WL����ǟ�� .Jf��N�8nkXaI��ӄg����C�&�!�dV?.1�te�"�"�Ǐ�2P�!�ě/V��m9 �ǳ�H�۴���!�[��DY���<�N��'�4!�D_K�f� ���i�Ak&���!!�D�t���	R�\j�l�G�ԁg-!�dР
��d���1QH�
���3!�$�8G�R,�t�Ɠ�V�9G�M�;!�d��kA��XE��ce��2t	!�d�>n$��MM�sH�s�
:"�!�$����C��o��X����Q�!�$�6��Ȉ7C��,�Z�iC�O�y	!��:)Ӕ�f�����)�!�,!�V�5� 'X�9<�h��J&!�䙼%�
�h5J؍9F��7��<�!��J�t���!���%�����-&!�ě�$���Z�` ��QfG�.a�!��4o�iߴk����e���!��i����gM�#vE�EW�m#���kE䚖�'�y�CNJ;D�B����ˇ,�\�X	�,�T�pQK�86pĻ�@O�l	j����+a�X�	�'-�9�1��N	�� Vk̍U�i ��d�	ʒȠ� �'��O��6*�&��`�ef�q�Q��� �HR�%/e���C�%D���iȸܠl��d| Q�O?7M�T�e�C/Իc��೦^4�!�䝫��9�㫛/nZEQ�O �����]ڈHjK �y�dX�lX��MC��Ƽy��J���>i��	�^�$��M��~( |xBfF�QBje�g�um�B�I1(&n�H�{#N<y��ϋvߢ"=�FE���$:t�/��ED\�ۑ	-��2���2��C�	�!N���Gb�+/��p���v~6�	7�\�(eE��)�'!L�I�R�d��2�O
p��5@�<"C�	�ˢ̹�,��W����ea�;#[|�d����$L�	i��9���r�
���"�;�УK����y龈��Ix��	��)�y�d�@�8� �"�Т�*y�'����tk�-@���OQ>-+�VR��!��X�)U�2�e�F�c
 ʧW\���'W���SC�(:�,�Q�>��g��T~�iL~�=��'�6��ŚSgB7+Qd����g��t��gՂ����Ѽc@��H%`V*_>���ɮ�a��� y�a��ˎ.���1�C�O|�Ё!��A�5�4'vڐ<�)B�gR�x����	��c�X�$k!�$
�ԊL��Ϣ��M�a��u�� �ȵyB�0��N�7A�[����e��B��X�gg[�'�J�hI2D����&��^ԠA��Fy���yc��R:�,��kڵw� ˓��2�*��{�'&��`dٹ����u��1��ۓ]�b�3�f¡}�>X���eN&�!�\
<���Ӵsx��`�$�I؟xP6
�9J��I�%�C�V+�����/�I�!;d͉#�2�,�*v��1��Oȶ���)U�c��j�8B�'�vm2BCّ0�q�b���L��r*֥$8�q ��.�L9cٴsW�>��"ݘ�%B!5�:���oK�F�5��C��ç�D�h�$;q�+W,Ilx��Hҍ�f%�{RhO+,��@����nረ�/�.��=���P���%��O�U��!_$ѭq���	lV�"O���0n�P�
�Ǖ�	y�m�U�D�x�d�;��B8�h�����i�)��#4�ԳJ`ʄ9"OP��r��>lH�ʙ�	a�<qwD�.��Ӗ|b�����2�vL�FF#%�Y�)D�l��"U6z�渹!HJ0C��Y��g�`�)���|B�Z�b��!��ש*�B\�0"\��y"@o��t��
!�
x�`���yrj�l�dr�O8�BQ���ߛ�y���2���)%Mܟ�bIA���1�y����;��9�ĤJ��PTEK��y2�D."e�A�x  �@"����y���ERD�"s,�x��d"R�9�y�K�E��X��Áx�,%��*�%�y��ԃ+`JH��F�(K��O7�y�I!y�|C��+n��4aΚ�y��"~��C� #$����ĕ#�yB�M=(#^�yũW�jm*Ջ��y�[%yQ�C4�L>'J�R�N)�y�fR�8=��3��;*� {�D���y��C&�lY`C(%4�5��L)�y�̞.8I*�H�&���c�K��y�#� �X|�Tf�L��pV�И�yU 1N�TS��7j���.t�D�
�'F¡�\���6��01u�X
�'��)��㑪6�5C1�)=H>���'�t��Ae-t��P�gnB�0t(���'{4��AEӞ*Fp�	���(.缝 �'P�U�Q�²v�n1B-S)�U;�'-�x�7U(02�vLA "�}��'[�0RE��*(�#v���^̊�'"���G�އ=�^0Xfg��V�I�'�p�Z�!�9U� Ui$k:�
�'
�����.�HE���T4��'H��X2�N�f�a�/ڲ\��2��� ��zc#Zy���SaJ^��H�q��'+�Q�irE�0��FJ5��H�z�(�7}�JN�w� ��A�O:f(R��^}נ���7;�XI;*O�Y��J�P��tj5���Q?�W�޳*e".��R�ʠ)�l�O�9�BF��r�� �LBɆ��)�
P��%�U�VLa�dZLI��#C
�����
)m�)�6���If�A>x�A��ж#/T�`�kd��'H�<YU�OZ8��d'�C����F��e�ذ�S:Jw�42΀�M���B�a�4n��5��{�H�X+�\`%��
�4mPCi�1��Հ.*B��)�kj0 � A�$���*_�U���V�@�$#�+|�T1��SaoN�Z��4V��<�!�UCj�i���qc�+:��4��*e8����Fb���m^�gN�	 qzUa4&��q��O���L�l	�@M�8����F�' �@�� ��T�}��S�O[�$�ތml*��V�=Șd+f
ĖC����&`�I-a��a�$H{ؠI5���<��Y��K���H&�T�`�׈oa���E��U`�O�%y�Q���B���ɲHJ�T�T-G��S��,cdd2V�V�}��|��"��oL�]�"f�c�l�w鎇L,�S�OK��ic]Ȗ�p�� 7.ERq���]f1��ٕL�H}��]�'E�u!*�j���c�;�  ���C��`p�,�~ I�-Ʀҧ'� �0|B�-��:O�ٓ���b]��;��П���$ڽ)�Z!���=S�� ��S�n}�@���w8� -�c�b@���я)��s�K�q��ulL>ɫே.]$�,��)�64��m�7��<
�x��U"�X��lK㋚�rH��	�F��rt@S�Sx$z5M��z�4`��[�G61�7�"W�ֽ����$՟�O��P+��cT��Xh�:�%�O5"nR%:a�P2�>��)1ʧ2��2�J�51������-.���!�'��]�'�n��r-M������O
��Շ"M�p2q�H�D�zU	B"OT��̏ If쨘�i�/9���p"O(YI��Y6yMtj�U�!�zQ!�"O�!wK��~�����O�o5���"Oܰ�(� ,����&0���"O��"��[��Y"CJ�RzE""O�`K���:��P!]�cd.8{0"O���� D20a��� -:Vڄ	D"O*x˳o܄)ݮ��aZ�"n9("Oځ�mp�1Xe��1��E	u�<���]s�-�#�fG���r�<i j_)'�&1J��W�`��@���]l�<iT��Ka���cP(T�<J6�]k�<I7n��~�
	�K<H����ng�<y0�9�*	���4tzݚ5��e�<�c/x�x�QpH�v���g�e�<��B�C��!�-�%G�\2��Mf�<�	P�h8�!����C�@����b�<�AɃVPt�p���,P�nG�<�υ��c� 5ݐ�I�Áj�<�K͋~f�� �ea�}yrJEf�<i�j̦K6�Y���lD�m�dJ�f�<�GoG=��(qdG;
�����\�<��`ǧr>晐F��qz\c�iL\�<���2{�*s�͛��tY7b�[�<i�aثs4��@M��y���4�T�<aWFc����jى(>���dWQ�<i�(�4a(�h�C��=����'K�<m�!^��s�@ʾxk��4���y���� C�!��5�� E�*� B��3f�X]��"Ub�LKr�:u�B䉩l��p)��U��ᅍ�ѺB䉝�*�h�b��4M�]���@�P�B䉏A��'M�&�N�+�-B�6s2C�	4g� ,�⣉5(e҅q�%A�%f$C��)3�|t(h�LՀ�[��2W�,B�	�H�x�{��*]�(�(g$ѩ3X�B�	�mRV��b��,X���gS�B�(6��LN�>�"pZ�&�+>�~B�I��r���nȁ^�բc��4bB�)� �MB�%w���L���d��"O(���`�/�|(ړ+�t�4��"O���C	V�p�0��A�Ə qN,�"O�3	�a5�8q��5Y��b"OV\Y!#[;9���Uś�vGvl0"O����;]�IR�M��r"��Ȅ"O�A���^{��sLI(�Ru8�"O���śU�~9Ise���N��p"O��#��.G�$-�oW� z��@"O�����_:h��*b�BX�B{"Oy�(D�R4H���#G�=�"O�hRV�ð~E��X�AD���"O�<6@�:l�� "�@BY��"OH`k�i��B
��1ԻC/��Kg"Of����� ="��yC3Y* ���"O@�0�>'&}���7E���U"O]R��C2+6`���.�|EY"O��%O+z�N�p��(Æ��S"O��2�JU������TF�[#"O�P��$�*~�8����z�g"O�|���Q�6��#���r��+�"On��v������AT�b�4YQ`"O�d�R@�9��`��b>t�`"O&��F��#|���h�.�UMJ���"O�H��� +G�<0��	;1I���"O��)S��.Znl�ĺI���:�?D���Ȗ�3&�Dh�BFj�9��#D�x0C%>�꼚�"�l�I�D�"D�(�����ZԘ�P�TG�0إ.>D��B����j1�B-N%;^��S->D��jB��/��h��Q�p
�ȇ�:D��F�[q���P�8ơ�v*OI�R)o޽Y�e��P "O6�),��\@���P��-k�"O8����<1����7@H˲�R�"O���AA�f�� 5ŀ�z (��"O
���+t1��C��Ve�pA&"Oh���Q��8�,3+����"O*<@��S }Ak�G)V�+�"O�$P���iZd��� KW���"O��A��� 
��` ����r'"O�ݫ��� PJb6���!����`"O�tv�&�Y�6- �m�"O�\d��A+q������ 05"O>u3���F��<;�A���2Ѫe"OfU����$r]F��j+l��-z�"O��aBL�'��Px�	�d�~tSb"O D�$"ն3I�q E��;>h&|�"OŉFAE�>�������w�bI��"O�q��eܳUJ֙QaHG"VHt��"Ob'd��-`�7�����J"O�HA�^<`hH� ŋsAڬ�"O��1ǩݽv/hP+�AI5t<^�XQ"Oܴ(�W3qV��q7gQZ�1�"OT�k�*Ң,�TQi���)E�	�G"O�]Ң,���^A�YH�Z�D�h�!�X� -�%M"�R�\�x!��U%x2ҔI�j�62@#��Ɓ1!�$];�%�A��d+�!@�X�v�!�$���%�� W�	��`���D�!�d�'4���Hv P�sܥJ��,m7!�Dښn���6C>�ȑja�6E�!��̈r�n�qc�>^�E�زP�!򄆊L;���+C�/W�q�%N�4�!�� � 
'
�_�i� eP�<�Je�"O2� JSO(�Ly�-�r�!�6"O�HcA�J�"����':�A�"O�)���!(,�����X����"Ol���$L	vd��hW�M��uI"O�y �ěrF����
6[���d"O2�BR(M0��Z�)�S�Z�C7"OD �r��[�����ȧ"�z�sb"O�l�Ǩ��c���I�l X��"O���DS
 �0q���QXVi:�"OD-1��"p�Jy�i�5V�IҒ"O�V�?T��0@(׮ut���D"O��Z����48tX#�fOZr`82"O���p��0�y���	U:\�d"O�=+��Q�b���JO�ڶ"O���E�Ek���"w���\�<HU"O 	ig��#U@���T���jU2�ʖ"O�Y�	I�Y&�h��G[�#^�Q)"O����(\P���b�$,ڱa�"Oll{��b���C:7j�"O���e�ͼ{����'=�p y"O�t`�EA:Nh��@Ʈ �J)��"O, ���
�'><ȓ�T$E���f"O� u��I��e�;Q/h��"O&�� ��ܜ����$�}2�"O¥X���z?�̢j͞
�B�"O(4#q�8d���	��P` �1"O��Oυ?Eм"g�s�:���"O~qs&��n"���&�{��ds�"O�ubU{ìys���:!����"Or��#M�J�(ʦ�إt��f"O�0�mN�nQt5p�l�K�֡�"Ou�u�Ι3�*��RIQm����Q"O�mI!�L�Q�䉃w��1��S"O��CFA�"P�QW��<Ӣ%#�"O��j�j��1*́D����P�C�"O�8;�h��z���f�І
{��7"O(X��g
:�,���.��y[8�;�"O<��B��~�h���,��3�N0��"Oh��[&rR.�Q�ʏ�N�x���"O�Ё�L�0<���G�M��	e"O�����9#@�ˤ��E����P"O�����%�����D�@��T��"O~T)r��f	X��C�=yn�8��"OBU`�C�Hz�� !>Z�I��"O48�7���|}�" �O�Oj,���"Oq�3A6
�rM�eO�3A�Ę"OB�qŭݯ#�H��]����sd"O��"���#B�� ���� ~�*0 "O��s�Αq �Uqc�_�Q�;0"O�� 0g�1]�@uiBl�+��9�"OM92g�:���`�d[�E���"O  8��"1����P)V4l2w"O������� ����3.��A"O��0jߺ=�ġ���+N0p��v"ONiq��J���P'�.b0Zٙ�"O�Q�pEQe芰�v�Y)aw ���"O�
b�]E�Lӄ�ϳF]"���"Oʌ�p"��3(��{E�:f["O|$@gk�SH��P���#U	ʴ�yҌ�k�ء�1�T4`��s����ybO��Zh����W$,�|y�I��y��@�VB����6�!�d��ye�2ލK�Ô��4#0&�8�y
� ��*�-�WS�4���>�P��e"O�$�"�1����D�f���"�"O�Y�R.D8n��ɣa�7e��u�"OR�*�	�
��e��3�t�"O���c�G�V��X��/l���"O��s�o��zĸ��;<o�Q�"O�Q�V��'�T�0�	i�iD"OJ�$��]?��� �4M[ڔ��"O�-hP�@�%L���-Ld�C�"O`�
�E�N���c�]�M/~� �"O��s��1F��f^�'���w"O��8���IƜm���4H�z�"O�p;��|.8|����
��e"O6���M�<��{�X�;�dE(�"O~�kE�?�Jt��`҄:�Q�"O���WcD���3�A.+V�2"O�	lʵ� BG�/: ��"O�4�7oC�n~��gG�[2�Rc"O�eӄ�H�@UX$h�G��5R�-�"O��K�cU 52�!��:u�"O��#�
�8<���Q�_�P�ٵ"O��9�g�R@��"�[��F��P"Op`��*������
kD ��"Oh���]	-PH�%@�:X 2��"Ob���`�2�����D�@%��"OP�C E�HY�j"��s�	��"O.D��N��L,�볇�%����"Of�bv�R�O���qD���b~�`�"OT����6�j�2ƇQ�"%��"Oꤳ ��g��嬓�^�^E�"O<��f   ��     G  �  �  �)   5  f@  �K  dV  b  =m  {x  ��  P�  �  �  Z�  �  .�  ��  ��  :�  ~�  ��  V�  ��  /�  ��  ��  B�  ��   b � D + �% �, '7 > �D 2N gU =\ �b �h �j  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>���f* 2���y�#W�@ݳ�i[)�d)�OЉn�g��|��?�u�)[�^�(p�
��`O��?��sY���ٴ���u>������\�a*���Dl"�i�T� b�h�Ioy�퓚[)r��,�6d�B�10�mIܴr��<Y���g��O�>"��	$oZ�a��Hb�ϣDp��O��M}��� V�P�&=O0=b�DݔI ��g! =���p3O����?� ��|��+�KW�՚�;����VxP	����0�'B�'�.6-ʫ1O�y��K�zM�ii#/17�t�ӄ�;�� ����O��}�ʧ)t����Ȏ��;��A�eG,��'=��-�\X����K�XX!�'�0L��]2h�ΤȃDO���e�%_�,�'���9OP�T�P�i��2�&@�5�5�d9Olmn�j�����v�4�f�a�`MkU��`+ J�7OV�d�O�dK9,C6M3?�O�P��eE�m!�m�:�����(tL��YN>�*O�)�O����OF���O�Y�����~�0��(P����<q��iP�C�'��'���y��  j&!{�it�Te('�C!<8j��?i���S�'H�
d�bnK�q�Z��&*S�ܕ��M�6���'5�*%F�͟l�'�|V�T�4��9R܈��٨m���(G�����	ߟ���ߟ�~y¨|�N)����O@%��������l@Kj,�L�O�Il�f��ПX���@C��К7tR�b%�7!D����BՖ$͂em�o~"/�U��5��_ܧ� �� Kx,��u��P����F-�<����?����?���?y����MS���pq���C�:�:��$|��'��nt����?}sش��?���bR�@�_
4@v��^h⤸K>A���?�'qɴ	bܴ���O�-��(Qb�@	EE�Vj��,_����ɒ�~�|�T��S��������*g�œ��L�W�t �����	fy��}����"�O<�$�O�'-MT�p�e2rR�ْ��V'
��'�$ꓶ?����S�4@R�'Y`��s���r�@@a�	$�x��.��q��T��ӚbGbeNA�5מD+gQ5� 1�
��Ԑ������I����)��|y2�j�x\��I ,�,��O>Y���H���-Q����O��o�[��;��	̟�����Rkf%b�kS�Rd��{�
՟(�I��nP~��T�Y���}���>r�<Lzc�R�G�z�:REE�</O���O��d�O����O��'Z�f9���C�0>t��-�2K�v%)d�i#e�3�'���'���y�z��.D ��	�j�@��i�%QB�$�O��O1�:��}ӎ�	�M2���%�<?�mBR�M�.�J�;�xã�'��0&�`�����'�m�5C��;��Ѷc�<aK�DC�'&��'.BP�\��4{'lS���?��0�Dh3G�<� P#�98���>i����'��Z4��4)6(��IM�"��DA�OPl���Z�Z�ɡ��0�)�#�?����Ol1�%�KbT�$�7�(W��ON�d�O����O�}���vil��!����`�@��X�T��O �oZ�{2`��џT[۴���yDM�/���/8���ÈM��y��'��'C� ���i��I�w��j�ߟ`�S�(S	J�t��DU eQ�X$-&�d�<�'�?Q��?1���?I��4�Rl_������S�������hd�Gǟ���˟X��"Ĵ_���q�o����E��"��۟x��o�)�S�|s
њ�mAG�|���d�N\��áE�u�+OFp���N�~��|W��Z%�Z?5�j5铄��U@.ui�a���D�	��x�	ş�Svy�r�8#k�Oʨa����L-P؊A4}��1&:OX nZK�
�������'��ɚ5��n�hQ�FR�jxZ�P�Kͅfٛ����i�@իx��d�[m����� h�R���bɪMq'�&�*��:OH���O����O^���O��?u��(V�9�P�k��>�~����Q֟��	ϟl�4��<�'�?y��i��'��T놯שO�JA)��3S��Ē�y��'y�d� }n�D~��ϸn��U{@��-�⣉G[l�}Y������@�|�_�������I� ��J'��X�vNN�,�xc"��ş0��@y�Nn�θx���O�$�O��'`N$d�Vg^���Qf��~��'�d��?���S�MחgӲ����Ǵ
A�|��ߞ[�t=x�W�~d�O��F��?�6(�DU�ʹ�"F�Dz�`[��]8E,���O�D�O���	�<���i6a���z��D��͂
3S��҈!���d�O�Ql�V��h����p(�n�r`j%���,cw����ߟ���d<nZv~R��Z�p�S_��Y!qf00�2'�V�qP���m��D�<����?i���?	���?/��#�n�M
h�X�m1��1S"���-�l�My��'}�O��a��ͅEb ���O�f�bg]4ZX�$�O�O1��̺&�z��I	����ӥ���҈*X���j:uB��'��&�`�����'�PT��t�x�P�T�Gy���6�'��'/"U����4.��\`���?�� ���갡M�,��q��FD(y�:�A��,�>����?�M>1Gf��A��@���l�eJC}~�(��5s8԰d�ib1��t��'�b"?a���24A%���g>%8B�'��'g��ȟ��o7�#�+�+h�:4����4�4-G�!X��?A�iI�O�9S��U��f/	�ш�@��$�Ofʓ6��p��4����30����Q��e�f�[�4p�������m`F1��<Y���?9��?��?�����<a�EZ
�LA�bD]����٦iQG,
ן���ɟ�&?����:��"U�B	�<�I�J�IcV���O��D�OD�O1�xa�5EO�8z�٫�ODN��P��B�v���δ<I$cK-��$������X�V3��Ss�TȠ�#��wy����O����O"�4��˓#��+*<�R
�B �t�/�@ԋ`F��yBci���0H�O2���OB���aTL�#�4�B2D2HJq�7m����� �����>���.�V�!2#��6@�c�A�"ǲ�	ݟh�I�|��ǟh�Ij��L�=r�"�?Z�um�<t���+���?���{�E������'��7M>���1I�h̩��B|�*/Q H�1O<�$�<A񊋻�M��OH#eMl�RX�7�фn�;<�x���'�N�Op��?���?���q��	�c�کcG�&kN�X+��R��L��yrn{�
��$�O����O�˧abAЀD
!`��4�����%�i�'�6듕?i���S��Z(�jp�0,X+@A�G��;0"���i�)$��M �O�	�4�?� �#�d��" B\�Q�@ *K< ���F8`^J��O��$�ON��ɩ<Ƹi}�k��A�(h(��.�u�`R� ��	��M��B.�>)��ZR��W+C!tlU�$�Y-!�(x���?tB���M�O��J�J��2N?a�B��mA�`� S�f+����Ho�@�'���'���'dR�'!�S;ˍ��N�Ezh8Q�/=�����iy�8@��'"B�'��O#r�g��n�'}\��GB%p�n��pe�
 v��1�)擼a�tm��<���N'&��X�TƵ,��0�lF�<i���J7j���������O����F����D߁���#b	�?�����OV�$�O6�nQ�6��\t��'�����&�HCWlėUl�d�Hŧu�Or��'ZR�'n�'ҥqČ�"(C��s4D��D(\�r�O��Q��c��6�U�s��'2S�UҮ`�wF\�],��t%Ee��'\��'l������͟'�U襨� ��(PD�؟�۴X������?�B�iK�O�.ԉ��z��W���&HE�
u��O����O02�&}���Ӻ$��(�J�D���q�b���My��4weڒO���?���?��?Y�j��@�!��#,��6O`SK2X��Q�4sBJ����?������?���$��j��)�P�P�J�5fb�I����`�)�)��*J95��a $�7]�Z��r'Z��'�t�k��
]?!O>A+O��#�)�� 9���(�2A0Ђ�O����O����O�)�<Y"�il�a��'K��Q��6X���bMH�EL��؝'�7;�	�����O����O�X{G�</x}�&�U�w�$0r�~Jj7-7?���'���I.�S���#��(v��)��A'��	avba���I��D�Iޟ��	�x��NG�H�D!{��K�'船�a�W>�?���?�c�ik�çS��A�4���Ҥ��`sF���D >Y��<����DZn7->?��K�7����p ̺#6�i�iN>.��83�*�OʬcK>)+O��D�O��D�O0�;�8\�W��`���H�.�OD�D�<)��'�H<9���?����i��L�lx'EH5$%��u�Xt��������O��!��?�b��rBAIV��*��1�EW)���,Ǧ-�)O�	U�~b�|"�͗u�����AHf|�'
^^�"�'r�'����P���ڴvPT�^�m�4��V�$��E	��?y�R�����D}��'7B��Ξ?z�.���-i�n��t�'�˶h��F���)z�*���/i��)� n�ië/*Mvm�����]���d3O(ʓ�?y���?!���?�����I9q����	-+t<���N���V�mZ�/BV,�	Ɵ��D�s��B���#C�)?Ӣ:'Ε [�>y�j��?�����Ş[�Mb�4�y2���7�.CF�=l�nY��L�y2�B'dn��	�h��'���I�8C!�,Zd����Sg�fi���	ß,�	�<�'=t7m�j�L�D�O��䎠x~���l�h4���Z�T��⟸ۭO��O`�OV�1F�]g�m3�����*s����f/9:x41��&2擼:}R&�Ꟁ�l֡ ��l����8�aqB���0�	���ҟ�F�T�'����'@�>0�	�tn��G�����'D~6��L�����O��oS�Ӽ��S�/�PXSq�c���I l��<���?y�r/��޴���)<u��'J�6�)��X�O}r���	!oXu��E3�$�<ͧ�?a���?�Ѧ���:n�,pTh��
TJU�p�a���'�V�$F�P2��'Q���������B��h�N�j����'wB�' ɧ�O/���S]�&؈�D��tq@�C�P$��k�V���e�4F��I�	uyrn 0�ŀ*�>t����@��08���'���'#�O|�ɪ�M;�mW��?�N�DV�d�'�:^���+�*�?�E�ig�OY�'\R^��* Dޒ$} iY�i\�wZ4]�͟_��el�E~bi6��@�O�w"d��䀕Ó:{��r�'Ȇ�y��'"�'A�'�����8)�|���%h"-�NH@����O �dU����u-YyB�r�@�O2���&�1#w�B��0x2�#���O��4�z�`#�uӂ�D^�Y0�Uj�����;VM�B*����D��䓏�4���d�OP���Q�����<� Qѫ	�(+����Of�>2�V���9�'H�T>��-%1����0Ax2�-xV���	��?�OQ�"ׅ�\��$?θ
�Q r82���� �i>�ذ�'F L%�"�A�?��ɓ��ߣ@�qC,��8����m����i�<���i���6�e
e����y��kV)Tk'�	�M��ƭ>���43X��[H�)�����}Θ(�D&�O��dC��6+?�;H�!���x�ʓS_�b��� 	��d�6D� ��͓���O��d�O����O����|�W�ݰ[�6���-I+��2�Γfk�6aX�r�'��T�'��7=�y�@�z.�˔)��$����`F�O ��"����"7~���������h^f�FX0�j�������hS�IKy��'��@�0w4���ɏ8'�v��'��$=�'�B�'��	�M+ $ԓ�?���?�#��=d�q�'L���q3�iՄ��'�4��?�����8:��ʒ�e�@�I��R?u���'���SM�;`��v'���(�~�'G�A����6N�(�E	S��q��'�'kb�'r�>	��01�^y�0�M� ����qMQ�>� ��:�MK/��?���}`���4��%Q��4J)�s�ܧ(��x��9OH���O��d�N�P7;?i��O�8_��� �6�jA���ӜE�6J��Kpy%�\����'�b�'���'� D:�ѣu������I�P��^���ٴW�H����?Y�����<�Q_�]?ո�,�D�0R�c������ �?�|�����,�q�F�~"(h`��f"9àH��򄁙c��� �p�O�l9��
A$A*?��+���s)����?9���?���|r(OtPl+	u��(%���'�G��{u�Ԏ)�4Y�	��M����>����?���{��Rg �<(;��SiЬ6�^H"�c�3�M+�O�<z#iܲ�����D�w���1
OH0�V�� �DT(�'��'��'���'���1�Y#"�p+!G�
`%��ia�O��D�OZTl��$"��8�޴��Do
4�c�0Ou��Z@�9��SL>Y��?ͧ16D�*�4��$ћ"M6U*�Q}A�y릈K.5�%�Q+��~|�X����ٟ@�Iퟘ8�N�sn�T�u˙L�髣��ޟx��Ry�li���4L�O��$�O�˧		"e��Ƕ^/����6q�z��'�Z��?��ʟ�)�`��w#>�F#��@�
}S�)�it9� bX�c����|����O��H>!T�~Ι�BoC�+��|��$�?1��?����?�|
(O"pmڎ������Ȉ�
A�	^�&ZMB�,�KyBdӾ�p�Of��N5�v��&�	u��	��ָ0Ԩ���O�`�s�p���h ɡ���V�O��հS�O UY��P@K�f^���'��Iퟔ�	�����ß8�IB�T�]=f�ܙge�FY6��5�N��7�ƥ��D�O��$&�i�O��mz�� ��ǂ�\,IXv��U��d9�)�S�<��o��<9@kR�sF�*#�0~�ڭ:���ybΈ�Um ��	�U�'o��ß���>[�bl΂����vCߤv���	�|��ԟ�'�$6�ܮvL����OF�Dg�r5����J2�Db��T��tӭO����OȒO@\�1�\)$c���@b�?��<�D��p�g�?s�}xI$�S�s�IDȟ�Y#틥UԤ�a����;	��k�NB՟,��֟����E��wo���"	E�������!VOR��@�'�,6��/��ʓ+Л6�4���'�#M���P������0O��D�<	S+M��M#�O�0�����'� h���gS�zM��Y��8ԡ?���<����?���?���?�!��1�� i��\�`�Y������`�L�ßD��ɟ�$?M�	�.�hQ�A�/�.1��-$�@A�O���)�)�@@�k%/�"�c�����I��*����<��l�a�|�D�/����$ހL�ʔZ��B�Y'V8:�n_;tz�D�O����OP�4�X�+��)ڪ	��KO�h ���II�:���XGc��yB�m�6㟰h�O����O~�8z%��їp�����l���.��$�{���Q>��#��?'?��� �5��I*���A3��	ßt�I����	Ɵ���y�'(�Aj�j"�'l�J���ԟ�����<1�4@���'�?a�iJ�'�,	���H;'����NX�a���r�|��'��O4�y!c�i)��3KltDb��O%"dA�Ī�1H��5LܧV��$2�ĳ<ͧ�?a���?�`��L�<��@@�� 0� �2L��?A���Mǟ��s��O����O��'kfz	�b�)2�,b���+n ��'\���?�����S�����[��Y$bT9	Y��AA�L0��L=YFF�#Q���7�R�V�	��4#�J
�k �R%��6T��I������`�)��by�a�x|�%S.y�<Q��H@�^>���R	>Z:˓g�&��AY}�'%bY��8n�	l���L��V�'#�).q�����֝8j����剸r��9��*ӲS��#��f��	Ry2�'"�'��'��W>U���>q�6Pϐ?0�l��*��M ��?���?�L~���u��w¨A�ʙ��,��sbɕ����p�'(�O1�����q��I�v9�F)*�x��E^�S�
��X�`���'[�1%���'M"�'>�1��
]��a�c��{ibmc�'�b�'�W�X3�4+H������?i��\��%�R	dR !�O�>��MÍR�>���?aM>1B[����W��\w>��G%�H~�  zF\�S�ʞژOqDL�I�ZG�*ڑ
z����+(Z%q����b�r�'�B�'�B�s�i���8l|<��*�xK�@wO�埐xڴC#�!�)ODmn�H�Ӽ�L��NyJ4ol����<y���?A��/d��ٴ��D�s�@q��'7	θ:�	Q{�EMG�lDa���,��<ͧ�?����?A��?aI9j$��˘t�j�����D�Ǧe ��M� ��ƟL&?)�	*��Ś���>4J��b`�$d��@��O��d�O6�O1���0��S��J6�Ղ�>�A�׬wJ��`Ր�x2�-,Y�b��Q�Ilyr�X1:�y�A(�P��l�vJ�#e��'�b�'��On��=�M��N���?9�1l2���q �z�hBG&�?i�i2�O���'�"�'DbKM�Pd � �'��f̊���΍2E�B]��i��I:7��Bc�O?��$?��ݚZbL�@Ў^�dQ{�B'%H��Iɟ����h�	ɟ���I��gt0�� A}`mrA��U6c���?q����V������'��6�#�D�F~;b$5h�$l��f��f�t�O��d�O��A�
�搟�؃�í:8TXy�%C�(Ĕ:`�I���?�6�4��<ͧ�?���?�fK�>-0h��'Q�`vj����ߟ�?�����=h�G�ğ��I�H�OK�,�3 	55ߔ�[�mL���O�!�':��'ɧ���-����rN�d۸Z�H�;>9P@hZ)l8�֔��S04W��IW�I�[e|ِㄞ&(o��x��o2��������͟ �)�@y.q� Q��kV�0�}�"��=AVJ5q�
ǭ�n�$�O��oZk�:��	��jݑB�� 3S��dU��۔CFwy���S��Ɲ�)J�02@�EImyBcKm8�"��=f:88�`IM��yrP���������џ���ޟt�Ot����#W1
8�����_�t)UDlӤm�u��OZ���O��?�������!x-�p!1E�d��31DB��?������"XH�63O ��V$M�N#��]�q��鳑9O��1�jU��?1go2���<����?�BM���\�"�.]D����i�	�?y���?i�����립�gW����ܟ�1ĩ�"Q ޹R�@��Mv�HU*�Z����ʟ8�?���H���ʶd��MԲL�W��f~�mI%75��(D�VZ�O;���	@a�x�zQ��6*T��p
A+%�'���'���S��Ȑb���0����IJ"%]�E�sK�ϟ���!٦,�'
�6�.�i�] ��P�*�2��BKG�$><��Sls����֟���DHm�D~�*�O�� �S�B&�<9��؈@�����)�B$ֱ�s�|�Y��ҟ�������Iٟ��%�M�}-��wG�.AŽ� �{y"�{��`�p&�<I����O�E���tS�_}ᐽ�bh�>q���?)O>�|b��#*0E[4��8O�j���/�i��e*!@�Q~҇_|�b9�	�#��'���*�jQ��f�<��5�b�O@���O��d�O�)�<q��ic�i��'���6,C��A��|����'�F6m9�ɳ����O����OPɀ&�I�V���
� غ��ub$�U+U/z6-"?9׉�<^3���4��߉.ԬÑU$D��R�P�<��������� �I�l��`��w�L�wF
�3��p)M� ���j��?Y��)[��ɗ�M�H>�"��0-tVm裣R�2Ĕ���?���|22��	�M��O��95� p�A���@�F�&0+�xz�チ�?q�)�d�<ͧ�?	��?S,��!���Y"f-x$" �p�!�?Q����dEڟx��O����O0�'o%Ne´ �:=yBpw��="-��'B���?����S���H�c>Li�3tCvl᧏�%(������������O����?y�G(����B��s5���/Q�Dp�PoG��$�O����Oh��I�<�·i)1 ;��aW����H"bD�����M���į>1�i�Y:��W�j��So� :
ɐ+O�9;�`���#Y� u��|�A*O�i�"PV�dT��f�%,�TC1O��?y���?���?Y����)̟H��4��o��\h��,�)a	�m�	;p��I�t�	X�㟤)���� �3��}��&SkS��e��?9����ŞS��13�4�y	�YC M1$��$�Ht	�F���y"�T`����䓫��O��DQ�>�eyڠg�@0�5�� C<������	񟐔'��6��A!�˓�?)eC����*DK��Tp��
ˠ��'GR��?)���)߰dSAE�i�2��p��=6�J��'��eiC��5I�n#�i���~"�'K�@��P��`�b��9�-
f�'���'z��'�>5���n5�D�ͷd�r\��,R�|�dy��:�M{Uo�?1�5ߛ�4�0P�C�ì\eQ�/�l$�;O��d�O��ѻ��6M(?YT�C#Ht��;����aɖ6R�F p��N�s�R�%�4�'j��'�2�'�B�'=f8�FkR�F�0a���-E�B �5W����4� -j���?�����O�n��K���n胗M(&ELXI���>I���?iJ>�|b��V�A��*��/0���� �m��4��D�;B@��'�'"�� L� �!AY	V�`�Jjn�5��ԟ��	����i>�'��7�ȜX� �D֫M3���O8��T{A�z`�����?if\�������I>�^�Q���B�>9:�h�b��r������'bX٣��?	�}��;Lh��h�24_��ȑEĄ$4,��?���?����?�����O���I�&+�\�@�� 4��R@�'�r�'�P�������'�X7�0�䏈E$P�°+�"A�����H�$��O|��O�I�%
��7�$?�#b	a��y���^����d�Y?Hk���
���'�X�'�"�'��'��X�J
�g��[p��o���yF�'��\�XZ�4>���Z��?����i]/P��VD&D��Px ��;�������O�.��?!��;4h���-�>����O���ԸhF�+�~��|�a��O��rK>y���uF+Ѭ��X��Hq���?)��?���?�|z-O|�mڕe�z� �O>3����������͟��I6�M�ξ>9��[�D��a�ytd�GEA$�u����?ylI��M��Oh`8�_�I?Q��j��Wc6�PvbT��y�V���ڟ8��ȟ���ӟ��O�@DN�IN�B�,>��p�"�i����'D�'k��yB$x��.�9h����*zd�a�r�1o����O\�O1�@�z���Ʌ\Ҵ���
��s��+�b�%m_��/�p�(g�'&�x'�Ȕ'���'&@	�S�(�������q<&5�A�'���'�Q��3�#vU��ǟ �	h���9�%�;����W͞�J��?�R����䟸%�Tr�N�pr��0�
X=Qf�hS0?�a.��j�#��E�'�`����?�qA��/�`�( D� KQ����(L��?���?���?���)�O>����KI:���/]�U��!j�O
�lZ������ӟ�X�4���y��Q�q;�ab�'��oPJ�I�d-�y��'�"�'*쪤�iu�ɔ(tQ ۟����2-��33O�b�<肥6��<����?y���?����?�%��0�\tÈ]�}߾X�&O��$���yC ���	ğ�%?��	*�0:��	&*�a*"jZ?x8pa�OH��O�O1�������lZ-��ې4�٥��"h�Ҙ�&��(p�H��E��Mk�NyrH�D�vY��g�
'�F�N�X��?Q���?���|�-O��o�a�T�	�G*4�j�ɢ2���8�L�'�D扠�MS����>����?���j03P&/Hm��/ع�Jlȓ&�-�Ms�O~���AG:�����w�d��"K�Xj�4`���p��y˘'/��'cR�'���'Q�"Y30EP2%iP@�ѕ�huX��O���Ov�mS��S����4��0'�qЁ&	 h������B
ʲA�'O��'���'�F�b6�i&��O���Ɓ�"Q�~4XX������NU�	14!:�W��O<��?����?���7dh\�eG�i�B`C�6I � ���?�/OF�l�_s,��I��<��g�d��l��P� �#F�d��6���J}�'V��|ʟP�f	C�^��hV�
�0��� A�v00
^�c��i>�*0�'�Y%��H���a���ς�f2��Fʟ�	ӟ��I�b>i�'.6���, n	��m�1t�*�� Ϝ6���`�O���Ц��?�T���I�z��f�٧2o��r���5)������D��=�&����g�Π�2��I�X��[��]=>��!���Z"�zyr�'r�'�r�'�Q>����@'g+��b@�K�n8h�B@�M�΢�?���?a��d�}��.�D�̺$gK1`�a��K�2���O��O1�n���e��� �9Z(x7⑻w�H��ܨ�7Op`!v�_��?�q�-�Ŀ<�O��}(��[(q���s��r��4��M��$�����O �Jbm���E�k���� �#�	���d�O&�-���-�6mC̃I�*�۵G��	|����Ηk��x$?ѐ��'��\�	�|y�� Q��44M,��Si�#t4C䉹e&$�� �75���$�*|FB���#�M��R"�?I�oɛ��4Ｍ�T#�4qVb,����\��a8O��$�O:�d:K��6m4?᠄�2�z�S�-���8WeĎF�UD$��&M��$�X�'!џ��wF	hw@%��N�=�.����7?�7�iU�̳ �'f��'��� ��:�v���A
YB���k�O}��'�2�|����E�ȥ����?���� �#��$aT�i�Lʓ �������%�P�'�Ĝ��� G�z82g��1�t���k��ə��?��L��R���d���,�h�;�*��<� �i��O\H�'�r�'V2��*�xP�QHȰz�xI�&a�.��R�i��	�}�8�8��Ob4'?��]I�u{& �)I���4�}7�	w����&� }�^����1����V�۟�	ܟ,��4M����ODB7�1���M&�`�!Q�YĖA��E�\���O�D�O�I5D86M*?�&B�	djdQk3O�La̩��.ߓi���ƶ�@'�p�'��OX�؃$K��<��ڧ3�T�����Mc G�?����?a)�̹�G&O�;��x1���a��������O@���O��O��#�U#��w�i���2W�hh0b� lB$l���4�(d3�'b�'vP��	�8hR8��bCآYt>�A��'���'+"���O	���M"��
*�0��p�I�'ˌ삓ⅶ!�H�����?ٓ�ir�O�,�'#�,�$>�r���&H�M����4�\Y���'�0�;Ųi
�ɶ���ԟ˓\ʶ�4�ށ}V�b )E�2��Γ���O����OX���O`�d�|ʀ�I:
���Q�V�EI�qz��E"֛��V�:<��'������'�>7=����&���˄���;a�iwg�O��� ��IY�[�6-|���+K�I�buKt�њ$�Y�!l����+�2DS��;�$�<���?I�`s!��,B����M�[�Iq���?Y��?�,O,mڮ<�V��	䟈���$�*�O�D(���<�f�PE�5�ɢ����O���*��۰r@F|�4�MG��2r%�+��	��ٙE��ߦ9�L~
#��p�I7T�δPaK�%�NQE��P�8����L��ڟ���}�O�B�@",�!Đ>��=��d��8"�e�lu ���O��������?ͻ��} "ni���9enP�H�E��?����?��G���MK�OH�֦����c�G�С��|����nG�>x�'��Iޟ��I̟�����I�1��Ⴣ�xP��R&@]�-��,�'[�7͐� �����O��d-���O�x�DC+O�aB� [A�jH�uo�K}��'�r�|��t.΢��	ÅQ9������R7
��S�i�(�<�X�Aȿ�t%���'��|�Rٽ0(��#�-L�N(Hr�'OB�'4����4V��۴l� !��f=�P�-�(f�N��g�
o`��K��jٛ����v}R�'^��'�\�I��0 ����.@��&���"Yڛf����Z�Wj�i9������R��?h���X.�r�B�ya6O����O"�d�O����O��?%yq)P=��r��"8� ���,	ӟ�����rڴo!�'�?�źi��'�8���H�9~�ڱY1�W�7E��!�|2�'%�O��i��i���0N~�	����6NZ���UwB�	s�&�������O����O�$�9R(8��sტvn��r�P@���OV���i۹��'��Q>�Qb���@p���1�J�x6�:?!g]�p��ßt$��'�)��Y�����$<���Q�ё6���ݴt>�i>�1U�O�OH0S�"�F��z�́q)�0P O*�o��B%]8��ʕL
�j8@���$	K0e�I�p��4��'$���?�a�O�c��m���5ILPN£�?)��,�-:ش���2^�Z���OK�I)f�R5�ab�%&�l����v� �	Cy��'� j�J�6a�2X)��ߪ��;cM�O(��]�x��z��G��w)�Dӱ� d���I�0����'d��|��d:��:O�MaIE�0�6dK3Ɲ�r̐-!�1OPd�q��6�?y�,0��<,O
 BbL]�I�ܛ�D�� (�A{��'��7M
3(M����O�����0�a�舘 (@58,�=��D��O����OD�Ot!����*�Z�33��4�&E�����8gb��jJzlZ&��
Ԝ���4�K��$uI&�¡H������0D��
�j��$��I�1	�1Q%S��49{�X���?I4�io�O�Wg��82�O	t�JҌ�l���Ox��O��2édӄ�\�4�W��?������;�N�Yɾ���^�Ly��'��'~��'5bf� ����"D�IA�YF-OA\�	��M����2�?���?AI~Γ�^%I��߂cW
����M�y�@X����|&�b>Qr��(� &|qC�)4f�9�T�l�Б�SH�2b���d���+��'nĴ&��'
8��ގQ�,��h�-���@��'�r�'�����[��+��w=�I�RmR��>O�l*5f�f*��ɛ�MӋre�>���?1��$�R4a���Z���e"C�JI��i�(��Mk�O(%a�����ğ���w��QS&�N�I�������-�����'3��'P2�'�B�'��D���!X7��ĐBJA�w������O���Ob�mڛ&=��'.3���|B�L?��9�fgE�y���rt��2H��'r���鏔L�V��*�ˇ9T44+�Ë�Xv�ɡ௑�{E��O>�O���?���?���w�Q���Hvx�Ie�Bm�y���?�.OjM�I1d\˓�?A,��U�L88���0$p�ٛ򒟐r�On���OĒO�2B��L�f��D��SkK�8��%#�J0M�N�n����4��m:�'��'l����-(��Ѱxd0ӗ�'!��'�R�O��I��MKB�Jj �2�F��D�Bů��8L���?�%�i��O
��'q�/K�{T�<��b
A�eƟk�b�'�&���i���,Ϻ��"֟ ʓ$0>�XVM��-���:���|f�̓����O����O���O�D�|r��TPM��a	" kL�E�­Oś&��;)�2�'���'��6=��<�6'"�0ŶhaA6,�; �'�ɧ�O��PJԵi��8�hEX2hu�\h3��
zX��V��Ty��3S|�O��|j���]��kC��p�[�^���+��?��?/OƖ�@X��;�'���'m�u+ж n@��1,>�C���BG}r�'�R�|"�L+\HP� ��@�J��D����dA"3�J	{�jW/!�1�nS�$�F���C�b��+bP\�W�A������O�$�OJ��$ڧ�?��ňkVZ%#c&��Q��h��E(�?��i0s�',rk�����1nA*(i%��\X�4[C���_�H�򟌖'�~�)w�i��	�5BJ0�5�OD*0A�N��x<۴.�Zp��qdSA�RyB�'�R�'or�'!�@:c����N�� �PDCV�	4�M�b���?����?1O~���YZfe�1��"'Zx��m�?^�~�Y�U� ��l�S�'�dУR`�1k�<\�6���j�(j�k��z�E�,O�1��(D.�?Y�:��<�p@R!�4��"BOԞ�da��?����?����?ͧ��D���%�7��ğ���٧/�>(J��� ��(�7,w����4��'����?Q/O����IYL�.qPU�[�:FP�q�$K��6M+?A-��{f8�������s��5LN����:u��0f��<����?����?���?i�����MQP��\?|�Ka�M�\b�'��dv�d%
��<!'�iM�'� 	s�(ϊ3hraN[�͸Hb�yb�'m�	�8@nn~R=sz����
�u	t#�$w������韔�P�|�W���ğ8�Iן\i��L�'<��a��a[t9�Bh��	Xy�m�Ľ�b��<���	M�Jq��	Q��`&�9���F~�	(����O���߀�)Rm�)3��isF	�L$��Q��.3R�����4��<��,4L4r��qe���jAa	[z уu�]�|_P��F�S98<`Pd�0B��5�6�bP�cbOR��B��V�P� ���^#T����#�'�@䑠�20x� ��T�YM��ʐ� ғ�Dp'�Y�p�"�j�.�N)hf�S:�D��W� �>	�UϮ
j�\��kq*R�
�Y��̩ ~���'E�,��uIS�*j Lk#��ug�}q�l��<ł�gڛU.�"�E�m��l��JV'2h��)�d�/O��)�2ހ]��!V��E���E��w>����G�.!?8B K��xsg�>�)O��:���O�dDNu�r�3`)"��_�ڵ��B4���O��d�O,�J���*�2��M�R��#Daԅ�4F�:"�Ԛ��iQ��ğX%�$��ğ����Qt?�ԡ��67z���DV0���m�D}��'�B�'*�I�|��h�\����?����@��@E	`S�,l��$���I��\Y�LB�T�hUS�cU�?�\����RP��`m�����kyB�?|\���?����Tm<��y���x�liC�x"�'�dN)3�O��Y.܉��������Gh6�<��N�f�'\��'��Tż>��OQ�\���i����� y�Mm�۟�IJ�"��?��D, 7I�a20��0Lzq���&�M�e�:1�6�'X��'l��ʠ>�*O�I"�a��qj���w.؁Ȧ�1��a���O��Gǘ
l�7�I(w*T��Ť@
f�7�O��d�O8E����~}"_�t�Ic?�5���w�2!YA+ޞQ�b<�q����$���&QF�I����͟��>.����aL�P�"I֦q��7�O��[Y}2Z����~�i�1��ɻ@���z�*>S�29�Rλ>I�����?I,O<���O���<��N�~G*���.ٴ��)�&�.12D �AT��'�b�|B�'����j�����A�%������`�2 Z��|��'�R�'��	�v��ИO^&	Ka�;d���ĈS5Q����ߴ��$�O�O��O8�x���O8�[���=_�	�p��5 �r�K�d}��'�R�'S�I.El�髟����=w�Y3u�¶G����@L?`yl��$�,��l��H<�	���P�M����a�I6��O��D�<١�8U�O���5��	��!S@B9�	�&`�9�����O���<�9O�� d���e�	R���f��i"�� ��i>剸&�6�	�4n����H�� ��ğ�P�4�h<�!�7m��P����Ο�[O|2I~nZ�~�S3D����Q��a�7�Qk��l�ퟄ�	��8�����|r�#�=x���dY�8�J���,��`�6�'���'�ɧ�9O����h=2��� �d����ĸ2�do��	�P Vf�/���|����~� PI�vY��8W�P��'�M�����Y��3?���~��Ӥf��Q��0��-���ǭ�M��EQ�)OZ�O��O$5��E�?P����a�.�e
�	�[�	�!��b���	iy�'r\�i $�ﴑ�!��-8|�U�V	A�	ҟT�	q��?)�'�����.�?Q�Y�f۴X���4A*�<A����O��
�d�?�!�K��l5�٘3�L�<���p�H���OD⟐��Hy����M+$�ەΰ�#@Ț�G<���WH}��'��'��	
lP
�hJ|�v�ң-�𘸣�G�F�t��"�N"����'t�'�i>��I_��O�e�j��`� �R�qF�{����'LRS�Z��ۈ�ħ�?���S!%�,j�N|�qk��[��T��.�[�vy��'������u�
�7;6M�#�a�����Q+��D�O~M�6��O>���O4���l�ӺK���"sQ9N��Z$
��ʦe��by�����O�O�r1a��ͰS� tR��cШ��۴+�IC�i�R�'/��O�NO�	I��P
��>L���&cߌDm����	͟&���<9�\`�$� �	� 2ʵ0RdF�X�0�гi"�'G⏁f�|O�)�O��Iz�L�� ֹ&W|�k�꒧GX�6M�O�O�\��yR�'���'�L�)a�E1(�������#����R�s�H�D�v���$����%��r�8[�� C+W�J*09q�cE<�ē�?K>������O�����/t\9�')=|��Ѥ�G�%�ʓ�?����'W��Ob���&�(R���j��C�N5�i�.���O���O���<��n�%��	�!&dHbǒ���͛��Ò9q�	ҟl�	l�IRy�O_����4�$�����H'���3�O\�ħ<a�=���,��Ā5��I���Pq�eI����
��,od���?�,O8��d�xr��,q�x9 F.t��MN��M3����Ozp��m�|���?)��c2M؏l�N�4*���@U�A|�	�� �'=��������6Jƿl����b�>^����X�`�	�X
��	��h������`yZwiN�ZT&A;<����bK==Ml�@۴�?a/O���)�)N� �@��C	g)P�:�gY	m|�6c�BI�6�O���O�)T^�i>�ņ7.�|)6�X� ^��ȃ�M����?�����S��'��z��A5`�!tT
���*�6��O���O`���@W�i>��Ip?��#� �d����z٩F`KЦ��I]�ɝ��9Od���OB�<_�,�@H�U�~5i
�����lZӟ(������|R���'K���"�1	����&�n�A���x��'���՟��	���'&B��(���fc��f]��#���!�O��D�OD�O��Ӻ3T�D�B��/�*��8����!��jy��'���'��	%>x�!�O/���ՙ�Kf�H$�۴���O���?1���?�b�_�<�3ȃ&b*H<  �|����SnfR�I؟`��ɟ4�'��=��~*��b*)A��6:H�g��YtxT�b�iI�W����ן �I�V@�nyRa�.(g>h
 ��$o'�X&�8�6��O*�Ĥ<��O\�G��˟��	�?�� JL-D���3#H�)��dc#�;����O���O$h�a��t�'��i8K�e��tN��1��>��vY����$�3�Ms��?������T��ݰ:���*�1J�y��@�F�67��OX�� �wq���f��'�q�l��w�F",��ui%�F�F�<d��i0J�At�~����O>�����'��I�K�����V>�����%>��a۴a|������OxB��%
>ݪ�A���T�2��4_��6M�O,���O�}Y�K�W}�Q�8�I\?�eT�\�ݢ!I�->U�Ta��S����Iby2%���yʟP�d�Ot�DT}�� ��L�-ۢ�b��V2��n�ԟ���F[�����<Y����Ok�Q�Q��c�,��{pBL3��	�;�`�Cy��'�җ�d���:�^ŉOg�Y����3/â����>a+OD�D�<i���?��f(P@�ucېC� 1r:(����K�<q���?���?�����ď�k�P��'+,*�A�J2V��"Y�%�^�n�Ay��'�����8�����s�x� X���%&(�sc�Zڴ�ckD����OJ�D�O���e!`[?�I�%6��q��-nc6( ���7�Pb�4�?)-O^�d�O����	��|nZ+6� �����^��MbTl��6�O2���<Y��^�v]�����?U�bjT.��h���A��b�z%����d�O��D�O�Lc>O�˧�?��O�*:��D�{�|E��%��L�j52�4��C��in��0�	џ ��������e�E\S!ϓ��Jǽi���'�v�1�'��')q���)B"��`��T�XP�lp%�i�,eH��p�L�$�O^���B�'��I�*�+uJN�cD/�0r�H�޴\��������O�ҭ4� �<YF+I�]�:0�G昆p��bԲi�2�'�U
Xt\����O���%�^��L���аP�O^~�7-1��'s��?�������i�<��Gg1X��� ��G	Jo��,H叐��ē�?Q�������gH�
T�kb�W<]2��fk}"OҌ�yRX��	�&?�culM)g4̴�cnJv}�]���0V��tiN<����?aJ>���?��$��E߂T�1g�=��d+�)O4�N�P�����OJ���O`ʓ&�n@�78�Lm#�nļ -����&�t�0�x�']�'@�'Z%��'��Ȁ��]�`��G�uT
��q��>���?����F�8l'>�aD떷O5j����Ѳp�x�Vh��M������?��<V�S�{�J�ޘ��t!'g���&�U+�M��?�,O ��FZH��� ��
w�)�O߿R��5��F�i|.�N<a��?	 .F��?�O>��Ok$�+�l�/-ë�F��Qȸ�@ش���I�#Ѐn�����O�	�h~���iU�H��Y�w�\E��.J�M���?!���<�I>����������kD�'�԰	a円�M+��^;p��6�'m��'��!?�	�5D�8�mC�r���R$��{ҐY��4*z�Y�����OS��=r`t	���ϰ�x��Q!H�t7m�OZ�$�Ol�[�Gn�	ß\�	K?I���.r�r	)�NDSL"���$�(b/?�ħ�?���?)��C!V]�!��Vk��F��J����'�~ �T-�I�%��X�!���&�� 6|ВW��.=u,��=������O �� �	C�\e�.�/6/V]���	}���Vʊv��?9J>���?��@�?�2}aՠ��x�|��#ri�l�����Oj�d�O^˓uZ<b�6��<�"�Ϯ�:���ܥ=6���R�������%������(�"L��d@��q�	�S�����	��S����'I2�'��W�|�5�P�ħ_�yi񍏸&�&D����$�`ks�iL�U���	۟4������K���4���(
]���|LTH��4�?9����"8" �&>e�	�?�Qņ٪��X:"I V)�1�� �ē�?i�=��Γ�䓞���$(R�*�k׈��u��_��M�,O�)��l����:��^���V��'�|�!� �K!��+���!�&x�ٴ�?���|!��b�"�I2��0�ơ'*j��Ջ��L�d6m�O��d�O�	\L�͟�AU�`Hth���\�nz�k�CŊ�MX.\d�?�����'^����a�X�h*eM�hks�r��$�O��$�m>U&��Z���	)�T(᧞<�H�!qs�����}��Ο���L���/ap��Mf���g�5�M���k�^�b7�x�O�Q������@MMda�os6HO��d�<q���?����4���s�@�dI:�X�EȺk�Y��ҟ��I��'J��'��d�p�x;�z2oE�k�j�(�m͑��'���'��S�09Ї����N
%�@9AŃ�|V�Lɀ�M)O6��<���?���<Ix�'^�z�J�.3��.�;`�P�O0�$�O���<��nM��̟�z���/�0��m�C�@�
"f,�Ms����$�Ob���Oj��s>Ob˧3^�\���A����	C�D.�8�ir�'��I#&e��ۨ�0��O:�	�{"j]Y�d��u/��pW�L ��A�'*��'f��\��y"R�<�I|:�H�cAָ�[,6܌=a$a����'�膃iӎ���O����=էu���?th�h����'��ݺ`� �M����?駣��<\?��	C�'9��\u��6[��������IlZ�����޴�?���?	�'H���uy�R-u�Ґ�m��Jy�&H*E
6�ʻ
���O�ʓ��O!�*��C<ah�o��3�̌���O�f�6��O��d�Oҁx@}�_� ��S?��ᐭA��w-P@%�,Q���צ=�	��	!|J�)���?Q�C� ��e6H$��GD�B���K�iZ���pT��'a�P� �i�� ��/Zy���ܺxrpH8�O�>�aNZ�<�+O���O����<AR$
Y�q�m�8DJɒ򌙵6�R�P�Q�x�'�U�|��ԟ4��+I^��%�16����X�bR����/g��'�2�'�2�'8�.��p:��X#b��zF�X 6��PdK�WF��'���'��'��P�DɅCn�6��e�1��k	�<Mvl0�S�p����8��qy��Q�}���FlycOU�2�c�h�9e����h�˦)���h�?y�+�g�'	����D.bЪɨ�_`�n�ҟx�	��P�Ip��O�r�'-����8aH�隬n�`��c�r��O�$�<Q1�U��u��4	��%⠏M3b{th��Z��M���?�iP��?1��������׃Ei&�M{%S�A����w������	sy�� �O�OX�⡯w��&d>�@�ݴC����Ծi��'���Oo�O��;yT �6�KL�~�2�e��L�~�nڙ?\�p�?I�g��?	��p1L��#Y�l���!'����'z�'��p!��'��W>��	S?�q"ߎw: ;�G�'$�����f���M|���?��|;��7Ò�����߈R���肸i����8c��b�h��d�i�1�@�yF��r��Ⱦ#����Ac�>���z̓�?����?�/O�y� �� Q�����BW�~�&u��lOn&�O���9���O����i���0��$-�����^*F�E�@���O���O<ʓ3V=#9�NġRb�7^���O��X����x2�'(�'�"�'g��O��������4`Q�V��P�U�����������I�^�DP�O�"c�&}G
�*�gR�h���#�L�0֪7��OڒO���<Q�g�IY\�K�ѿk�t���5m�7-�O��ļ<�"��,Zl�O�"�OL�T;���"in4�u�_&��t��w���lK��$§�n�� �!�נQJ�-���H�z�Z7-�O�dG�Y���$�O�D�O��i�O�����m �D�!YT���Y%YF�ȳ�iA2[�4�U�!�S��<J\���J,O�QSRDԴ$R�7��/8��\mZş�Iԟ��sy'�L�I�\2� F�\�
�6S�H� �ٴG#��Gx��	�O6(I�}Ӕ�S��Ŭdrd���Z�M����I�A��0�}�'<��?��M;��� �d
�d߱Oz����D�O6�D�O��rǺ#��U�S��> ��1��������'\���}��'Vɧ5�mU�G_欛�D;rubL�` � ����Os1Oj���O`�D�<iP
mn��+���/'�2���1w�������Ob�O|���O���t� �=��2�)ԜH>
� M%~?qO��j�]�#r�88v/ڝv�:��J�\�e�bF��$=����f�����H�J��t�
O�T@$�X��&��q䇢_�c$���.s�%��C D��@XĩT�*,<AHr&~5HIP�=A�f��$�˷/5t��$��=f7�`�D�T-B�[�ո{~"h�5d+u��%���ƭM�=���#R_~�����3H���Z�J�m�06� �#+Lo���̚CX��DJ$x�.�1UGGn|6<+s�R<\� ��!"����^vܛ3�Jo�Z\�	����A�'=�|���=��⡂�?�	�|��σe<Hv!��$�� �!�W]��3G $Q 3�Z'�tx�g���<���X�1�Ô��rр�Ja���a*�'����?���I�O�@I4�|�``h #l3���aB0D�48aX cv���Po�S�ؽJr�/O��Dz��-.��82��!_F��6j�+	�<ꓨ?�|�&�� %�?����?A�Ӽ�qJ�j��`8a�@"�$ɂVHɧ+�$8���@�$q����\�H��L>��	��<)Xa��̎��иY��	�����X����Q�D��}&����Ɲ�pw��G��
�
8�p��� �'p��|�����^����I O`���%@��W�!��F*:x� ����U3��QD��@��ɏ�HO�Sky�"6�hADR.�D��s:>�f� ��ߴTB�'}B�'#6�]џ��I�|wF�hz���� ̰|� �M�v����E��'x)X����'���J��!U�l	s�G��$d��(p_�*F�ң���<SbV�����!�B1#��8�HT�'�R��D�� iX�P���6�`�m_|�ȓ<~V�[r슟��y0� �7<A�<��U���'jVᒲ�{�����On�R�+s	����a��*�����O�特U���O:�ӜDeݴ��V�4*W��>����CϬ ϊ-�㉈;�2� �p׃� �H�E�?aH���V%<O,@ �'��'m�D#�
W���]R�L��K���'��8�l�36J`��&3w0T@�'E|7-T"rn=�2��7�h��Ōt;�1OJٙ��TϦ����t�O;��[�Y�� �+�|���ҭ�2	�4����?AW̐��?��y*��I�F� �ЂCP�c@6�rvB�%%d�'�^�s���I��z��CF��kw`�0l@�7%�Y��,��C�S�'f�&��V2<�\��l��I����΂8k�M�	 ݠa�Qd�z)�`��$�HO��a熻�`�C�k�*g+9�,�����	� ��>x�Rm+w�Nϟ���П���� O�׸�h�jȤ"��!�c�`��XI��I&<�|pE>?6�1��Z�/����+-<Ojl��ր��P�AE<�ĭ���'�>�����|��9SA�4���Y�4e4 �����y�I��o��"�dY�1�^�1���$M����0�tɓ�h8��"��NA���)�8�ᇦ�O�d�O�������?Y�O�x�2���uix����TH0��A���x�G#\�B6�W�ND�)���tO�x�'T��c�U�@
�(S4l��7�T�JD)��?Y�:b8l�(���, +����tS��H��R;,��՚����
�D(�	+��'��:�tӐ���O�A:F�M�8U�Q�@�Z$���8��O���t�����O�� 9R��;���;�b�y�bP���$��;F�xА��'�����D�j���6���v�Ǔ=>��Iy�)� �:��k���iT튕 ��4 W"Ot|�d��P���GG�o�*Mz�O��lZ�-d�:c��_��I�˅�3xdc��S�#  �M���?	ɟ�=���'�6���C\�X=�52e�:��'Knh���T>�+�< �E�)Apb��.I�6i�O�����)�^}̠#7M�;f� !�<G�.�'��9�����O-�@k ��7�{�T�U��݉�'"1��k[- M���E	R=|���ɲ�HO�m3��8"�8�^��ȹ��im�ҟ�I���9.q"(��ן,�	�<�]�������'
��a��+�� �<Y�%yx��a��J��M6�+4���
��(�ɋb������I&(�:U�΂B�q@C�� %c�l`Cd�Oq��'Ġ���z�6�yAH[6&2�r�'�e�UjJ�d=1��'(l�$��O�4Ez��ӫg��TkC�I��Y(w�1S�@��f��4-0����OB�v�P�;�?1����$*��u��9(���#�D]
�k� l�t�{�'��A҄�k$p-��2򄺑D>�x��2cnh�NQ�3	.����8+����?�5��F|]�q��'==�X;ub�w�<Q�����ݛE�I�r<z8Kt�Ar�ñO��	��Ц	�	ן�06`�j@�U��B*^=ʱ�Sޟ�̓k/��I�d�'I/F���^�ɋ�t�Q���X*��1�9��L�O�$«Qs�d)���ʠ3v$��'6�����Fv� ��8G^���D5T��ȓ"ؙ5�Ɣ1��X[f9��]蛶�/l��9�/�`�HB����'�
��3bp���D�O��B�ք�	���H��Jj�^(q�NF"(E�H��ٟ�Dh�˟ �<���d� nZP<���X�(�=�&� %e��\��Fx�����mζdh�$�T{����%���3���d*�)��p��h�/��P��p�vB�"�C�I��6����s�քq@Ks����w�'T��8�U '2��ȓ��//*�Yf��>1���?Q���(Za����?���?�;p�@�q`ړR
t�E��%Us�MrԨ�%%k~��2c_D����լ���n��l�u��4_�v�`�Bϐؖݚe�H'gKɛw��&x*�`r��e�g�	8+I��0�\2dob�*���_���	o~"����SK�'� E� N��ad�,�(�;���H�'�J I��(`P��bFhG1����O^�Dzʟ��~i��G�J�,�[��\�a8�}C��mx� ���?y���y��>���O��ӝ>D"�BC�Yb�-%�ɗ�F��,�X[!�1��h�1�� 5�F�G
ă�VC��3�r|�B��p 6��2j��Ȭ���O���]a�Nu	 b�yR]��MP!�!��R��K�i��lc&�)!��Q�1O��>��Ƈ7�F�'�R�G���i���4X�%�o�98�:O��E�'��5�4|��'�'fT�;ӏ��-� |�mɏz�P;
ǓenH�?�E���x���a�� B���Y Q8�H��O�O���G��Q�XM����ae��b"O(]���	�Z�h+f�Ȝ+2!уO֠mZ�Jǈm�U�eĠ�Qԏ��>c�8Ycm>�M���?Y˟��4�' =�
�PdņO�H0@�'��g2�T>���tbBF�,Y�g����O<pjv�)��(Zא}Z3F�yI��'ɩF��'�����ט��Oa�i��o�q m��RD��C
�'��C�� � ����:_XX
Ó1Q��L�$�,j��h��@�8x/p���I��M���?q�eA,�T���?����?ў��%V6�8�kā�Tt ����'���*ϓ��	xU�?]��z�h[<)����=yF��Mx�����M�'g<���ҒpZD
c
�[�tZT�)�3�$�5B�`����,���Ȳi�B�e����FW8vH�2r��c~����"|ҥ&��+�Vy�(������"��d�d���?q��?ɞ'��OH�Ds>��F R��۷�M�[�B�	��� ,,C�ɑeX�	����Z�FW.\ht�"-�xI�#vj���C�	j���R�9#��'�O� >0�g
'q��p%�5(	V"Oxt�v2���c�I&)�J�rV�$�Y�s���u�i���'0�'�����
�k��Z؂t��'��ɗ �"�' �iӟ.��|B$X�LJ犈7��R�狱�p<A¯�r��D0�	 ����sA'����I1b�~��.��7NuY�c-����膶�!�$�� �|�g��6!�H��!��]Ȧ�0 i�.�������oR(( �M;�ɧZ�� (�4�?1���im!��i���c��*���*�Aԇ0���'F\��'1O�3?)� /L����ߧN���NY�ͤyi��?-i e�	,+J�P7e'b��c�.*}����?Q�y��t�@���	5w5��rr[&�y".J�. �$+ 	B�M`ْ�K�0<�W�	3s��A�V�؀�:�+��K�}J�9;۴�?���?�W*�$faJ�����?���y�;g\��!؛f&���A�g�*�y�(L���<y����Q��%�R?E�吲b�Zܓt�؄�	��Ѣ��j�� ��ȋ�x�<9���ʟ�>�O�I�6�:T�L��2�,�m�A"O"���蓽fOZ�ꗄ��4zUˣ��Hy���ӘP��H ���V��DJ#`�h3 �|��I֟t���<)\w)2�'��)��.\�	Fau��8����7�R�"dO�ah5	ʚg>< ܃*��5A��K�!��ʛ��,+A�	�\%�*�� ��'����^�"�F��ІI�h�.T�F���y���T��t��Y�y�梊��'�`b��,��M+��?c�N�ZG���Sf�P��Ǥ	�?)�'L�$8��?��O �����i�����4�DeC� �H~����:B���n\�~�-h�"Tk���{G
0O�	{��'<�'mjp��A�,	hxma�dT�oF����'-�i�t�ХC�`����%e̠}3�'�b6��&�pe	4Ɔ�o���:�꒸Ov1O���U��ئQ���d�Oe�ة��uv�QAp�G�0�а��%C�0K��	��?�#�  �?�y*���� d�P�Y9<?҉c֦� ���'?�2�����{VH���L�z�hDB/U�
{�6����	k�S��x
8# ����s˅#D�u�ȓ4j$4����.�uɄ �$���I�HOx���_�bi+%�T�.�Jy���G������P��1�8��GeI���	�����iBB�$h�ڹ���N�J��Si \̓mђ ��	=�R�j4BMp���!�V GO���i��,<ORd��(��G�n����/y,]1��%�I.{, ���|B��9��σ,NZ\��eH��y2�\/��:�INJ�trՄ����dLc���.��F/YU��b�I�;@���T����m�W��O|�d�O��	�c��?�O���
�3��8����F8z!
3���xb�" �
d
d�R&����h��1t� 	�'�d�7��*f� ��_���:����	q����G'��@f��w��r�X�a�/?D��H2`I!_�Ā�n-%2�r@'�ɽ��'BXpiU�d�D���O<��%� \6:xç&�s,�Q&��O��I�j����O\�ӱkZ��d;�䆔��ᑷ U*<Y�Ԁ��x��-��'��l@�M�B�ʕ뱁.3�L�rǓ^0
��	D�&䂉	T�=�l��,X&�fC�3*S$!��`�$(��m`q7�B�I��M;&��.
7��H��]S̓W"]X��i���'���M���_�g��5���H�Zւ!��A��'<��D�O�HѦ��Ofb��g~R��H p("
A`n`5ò����"<���EZV?�d���7HL¶��`��^0o����,A�D�R�ݍ2>N�C�`/U!���E̔����j��"�9haxR�)ғqH��I���c����ĝ��	��i�2�'�"BБ1�/l���O��Df��.�WG�504O������K�xD c����$'<O�Ep`S�+Eb�S5�P$!^\���ړ&K�y���1r,+�E[��h�A-�!D�1O�x����������:A(�8"����L��S�? r��#�-d�����!��d�8՞�ؠ���"Ra����(Ӫ�f��"ۛz��1�Å��\2��	럀�	�<�Yw�b�'@���Ӫs�i<L�Z�{a��d'&4BvO$�1���J�6lՁb�q��$^�Z�!�D���-�������F�*3�~����'!���8��ʥ��m/YI���y��"d�i�<њ%�(����<a����%x؜0lZȟP���K���2��&�������>��$��꟰`T��ʟt�I�|�j�r$%��ㄠ�(3�t��$H̜{��3��,O@H���ߺ�'����R�у<� RCY�+�<�j
�Gz������蟬Y'돇S�������Y>�p��'9���SJN�[&��,;^���&C7^>B����MC�O�6DxK&�ZZ��ER"��<�(O��Q�����	ݟ��OT�q �'�Nh�.�� �L={2,T�j�J���'��/����T>�a}��DKw�1yƤ�6'�O����)��Y=�A�v���E��t"�O1P��'��������O\�1��%"2�y�qEJ�5zXh�'� (����b
��`��X�L�Ó{�����j�G4��Y�aVZ��6D�l�ֈƳ=�h����'61qC5D���!� 6������_���q��>D��t�_��r �a�˻w���#3( D��0#͒UÔ�@{8��g-�)�!���5wF4����*�t(��,ǇQ!�DA� �`�z�L݋B�f�VJU=�!��JnN�Ag��/��ӓ��<�!�dJ��TlJ�B�9�8�"O"�:S�<�,@s�Ω/�\��"O��hg�]/�\����;"�|��q"Opy3Ň�����c(?P@��3"ON4*�D�K@���p,��gL���"O�tpc��>2���ؕ�+�z͊g"O΄��l^Sx�C7�F?g�-)�"O��J1�\��)zE�ݼVH>��G"O$hh,�b08�q7��_th�"O�q	�D�CD�\#7��l�Zm��"Oj��t� 6ŘqH� ��l
��w"O�Qy��?:I6pbD��[���e"Od�*&k
Q�Q�׀��B�"O�m�5eƳ<Jj(\�}Y�=�q"O��@
�H
.�����$ES\$�%"O�x��7@,Xre��O9fH�"O@@c��mf�9�D*I���`"OR51�JۻjI��R��Ѯg �ŢG"OdIw�?��e2� �jh`�q"O�KE✽�Š�Oh����"OH���,,����&:=h�m D�,��ނw�̍�6�؈n�~�c@�$D��Z&m��3}:��0H�V�l01sN8D��C�-I&==7/['^�*����Gs�<A�ϝ� ������(:�t5�wLy�<��j@��Dtr�L^-H�4}�!&�@�<�
�~ABx�a��$\�U����|�<qS.�y�(Kǡ/��Ͳ%��x�<�g�?0��tm�m���Gs�<���ش�x�i��bVipLl�<�J�<sZh��䝹9Lq�rlHg�<�E�U�����F������Ec�<�p�>x�rG肳& B��v�<YǬ�gw���шC� ����h�<��"�#/
d�HQdѫK���&�g�<�b���-��l�R�L6Ak�<	��S�r�n��'� =צ�y�l�a�<ٗBݮ'e��T���zu���]�<� �d"w����F�(�,�?Z�u�c"O���5�?lc��h��\��(S�"O��CBN=�PO	
	����g"Ox��u��:}r�����t�m�a"O�B���(4�q,G�J���D"O�i��i؏=�-ca�G�B��M�"OX+� ^����b$c�Z�l`qe"O֐bN 1lM���4GeH�U"O�Ґ��
 �2!T8(a4	��"Ob�j�%�$r
v�rq��:%D2�r"Ox%�6�:�d�;�b+C;�<��"O����N�t�|lSa�_�3T΁k�"O��y2�
��MQ�"�Z:���"O
ӃB�<gĸ����J�m7V���"O�q넃L�.�tY���Χ3S��0"O��9�֍o�ňd��K>��"O1�g0 ���(S�H
=p��"Od���݆cq����x��qw"OT�6E�Z�d�#��.���Y�"ODY*����v���+��4�f5{��'�v;BH��F�����kՔ�B9F)����!ӥg-4��j��
�H�4d�.R�D��&+ړ(�����,�/	Qbb?{3��>K� �0�A�O�%��-*D�(  ��
a4�2f��R�m�`b�O�@�F.g��P�H�"~��o���|i+&bͨe��!�U�ԏ�y��\�R�e�P[�^����������FU|�:Aӹ��<�1$��&"���BL�*(�� (��K�9(�}���E	��غl�܁"T$��y�6�0�!�8���ē�����-��5b�/:����I�o�� �R�x2���?�'nC~Y�DnYV�85R��^�H&Pm��I!T���R���C� p����P�V��ъp�y�(A���[�S�O�P��`�ղ`�(4�Hf�����B\���#~B%�$4p��5D
�@Um���K�Z��H@���ä�J����N���	�+@�·`*n��U�n���tP�D@-��'�dp�'<�����Nz`�8�EE5o�� E�8�z4;��ݛzz r�'rѴB�	sn$��b���q^����#�<���pgFC�+�xX��9>�R�E�/3�$����Oq��+����8�P�"V+��p��at�'���
!"]+�򤔖]唠P��<:�Ċw��2Jh�QF
@�|ɧ�'�Ȱ(�iY���	zFi����>N��&A�n{�DӠ��9�0�}�D�Ј<q�[E��@�&r�����l���ѝ�
�`R g�xI*��6O*Ȃ�+��K �v��4|�m���.l��c�LY=�����/� IKǯϴ5�*ɀ��>�f 0`GR�*H;U�J%m7P���'r͒�H�
M�Р�	��/X�	 g�=T��-z����0A��D�(�?%?����'��t���F#؝��P���=!��܋%��ɀ\�f����R�$/�h@A�,-����cj?y5�'fh�ߟ���&y݉jD�>A��ثlϪA�E�-N^} w��x���~|[��ًOdn]����7J`1����~2V���"ˊ9Hl��I_ )�#k~�������&�0<��aYsgN�jWEn౫�#^�	��qO>��+N�M���3s���P.���'p��[�� �D�B�́u$�$��\�%��	No���#hg��H��=�CU.'&�9�򎛨 v>X2��A4%2qaU���b�T�'E�	�C���@�.��d��S�D1g�zXhg@/�O��W�Cy}rI�N�~D�q�S,|��d�g��8VWtq�.Op�ʑ���#���B�[�r����\Y�IK��%�G��,yE��B�
m"���IH����"((+Nv$;��
F����Ƽr�$��v�N�3J:�cB�ѳJ�~�)�B�	-�9�O�u�tk.�B��M���=AG��ghݿR��⟬�S��2unИp��B	��Ȋe���������Q����D-_U�f��D�Im}���'n�az2�O���kq�Z+n��J M���sT���VG.���`אd�߻I��Ɂ+-�ʧ[�$1�ES0A�]:T���a(�x��M�Py.�� ����U��$����@ ݳ'H9+�^DX����G�_tIn�Ѓ�m>-�3�i���;,�J0) ����#�*q"��*TO0�(G�p���{�hC�G�d�p@i�/L��1�T�3E�%y�DF(G���ش](����)�f0�c�:3�*�9�B�j��<��/x�F�Z���vNQ���-s��$�g��N��1�B�}��ya�X�?��,*<���$�J�P���ޝ}W��犛%a����[;>E���+��P�
Wڢ�ͧ�LQ�w>� NpZ@+H���5q"Ō?��"O ��2#٨(�bH[���/p6�H�H�H����&���N��k
�$9�Ȳ�?�	� 1󮌔gm�t�S N�XM��`�!𤔤����7�כ%O\���Ϙ*�ju�ӈC�t������'+~,��j�c�'�\y5��3��Փ�)�Ě��Óy0��c��,19#� ?�?	����Y�A�\�P�|HCCYc?������dv���.g�H@լG/+\��OD��6�A�>����5����S���0u7�$! '�!�0��V�~N]�"O��;��T�6��y
�)�f`
��ѣЉS��ThW�� ï^�wo�b>7�^�����\��@��=_lZ�B$'x�<!HL 7A���p���2(��S1b@Dq��i���d��$��9Ҭ�E�c���>
az����fMt����?�����U��x��] ��A�F�<�r�Ty(��I�
�pɤ�A̓o�Hqʢ�1�������c��ݛglɕQ?�e��"O�q�҄p���0�ՃK��*�7m�(�O��)��3?�����
m�tZ�@�/s_�e��
�C�<i��E	n��a���	Rh	�&iܕ���&�O� XV��
�@QP��YIdԸ��'���<�6��;g/�B� (�B�j���O�<aɚ�p.xhc�����"P�M�<���U��,h��cL<tʣ+�G�<��v�-�2�
�P����#�\�<e+8F�������<�#�ZX�<��OU�m�G:
�\�#c�x�<	��T-@��"�˭#~��7�Bx�<�����oz���>?������NK�<A�\�*4@�+G$� T��Ļ��k�<�`�K�z���ѩ�2RF�LS�i�<�R.�,��t��T��8{0p�<Q��Q&f���"��h�h�d��m�<񢥃�G���h���UޡӂgN�<QY��jeSk&F�@�G��o�<�`�B�[vh*�/M�oc�4Kd��v�<�G)E�J�"h�@�,�0����n�<�Λ� ������V�O	p�"��Yh�<��w��Q�K.����c�<��,��D��h�i~B=��R{�<y��̑
wҩ�g��R�։p�&��<�ueM�z�([K���i� �y�<As�ا|�r��c�j� �	��Z�<�W�����"珂p(��T�M�<�'�#L�{7Qw"�Č�I�<��`M�G�$�n�*�)`w��B�'��U`,�'@��%бB]�1i5"�l�6Y$bH��FD�#���T��sM6I"T@c�d�8v�p��=E��Jhb��W�Ko6�Q��J.ia��?��-M�V&,�D�$́�k4T{w�ޥ?����4�~"�۹/�>݅�	
e&y�GLW3;��Ƞ��ȌL$���B�~�d�O��>q��dG$�����ċ��N�MBr��F �M�!�U.ܩ���z1$Q�u��?c�R���Ly���S�8kG*��ا�I����R�(�[92��".��x��{#(�"���=O�큇� Ya��"��[� ģu"O���C�F�t �꒩ �,�PP�D�'����'�'��Q3�)����C��Ԅ�C��ۃ� �e[���d�-���Q���9� &��E��'����fD/1��ᤑ7N��4��'զ}���x
�a醅'Xi؛'F<����Q�0>ɅM?5)�8���O�x־���c�<Y���V �iэU�9���e�<���~jB���[�A!p� W�<��%EQ�h���	y�b��Nx�<9�˱$��+�?��rfD�<��	�p}<5��� [�\��&B~�<� dU���K�3��{gg^�IА"O��0�G�Z%&1���J�L.�h�s"O���i9b3��'H-=r��K�"O��p j�g��!�FH8|�:C"O�`��� �!��1 �E�<sk�Ia�"Ov$#d/۸p:��O�V,��"O���@�h��T;��'�H1�c"O�ysր)m����5V+ �̩��"O����^4���Z����f�>7�:D���{�L�(��ya ����9D��J)�y�\=xGꙮ1�⌀�	6D��;�G>������D ����h5D��	�A;@���Qn�;����d�2D�(���Ȣ6t@�c�U����0W!-T�L�kL
��C��U6"O ����-a�2 Hw�[�1"O�1sd�ײkۖŢw�Z�.X�I�"O���U ΍�N H g{kd�t�U"Or|)���H ���U��,�"OT�ؓ�̾=;h����?;~EY�"Ou��[��i�l%a��;�"O,�Y�jF.4�����j��i˔��"Od59��ڹ6�h�#H�&��"OP�y���E|��;H� ��"O���QgÜ0ybmy�	��h��"O��	'̒T��z2��y����E"O�xƕ�f��(GFHl�03�"O���@U�v���[�kܒ?]���"OP���Jv�$D	�Ɉ�uY ��"O^��ôb�[�n��$�RI��"O�`��:�6���29�B`"OPf��6����A抰 l݈�"O�����9,������%�%�q"O�X24�@�vLl�ʧ"ݴB�����"Op���Hк���S�	E�0�"O|;�!T0A�ϗD)�ə3"O� �Q��HDnX;/���K�"O�Բr�X�e�|(0�΀Qf!!"O��腨޳0[蠩 �+=�Ѹ�"O��*\c�RYa/Y�B80�B�"O��*�Kڞq�� Ch-!G����"O\�ʶ�V(6
]j���C`��3"OU��J�'d�2��ĉ�::~i`�"O(���ER6>� �e�э(8�i�"O���EK�=��i˅(_y#���Q"O��S��^ J�x��G��{����"O`&LH�H�B� ��e�5 �"OD�rV�F�C�H'��0N� Qv"O�������f��2BH N�u�w"O�e�$ň).&^I���86�01"OR,�v.B-$�<;�)hc %8�"OHY�Њ;8��,H!�<\X��E"O�LS��Q��<����c��|k�"Ozl�oI<�J]��)܇S�<�c�"O�=��lڐH�4���G�	M� Dz'"O4H��l�9,F|P�7	��F��� E"O��H�iJǮH�����lsu"O���a�/IE$����('�p�"O�d�D��'^l�"�.P�t��G"O�8�܅9&`sQH�6wR�#a"O��Y@��"=�|S�'�'Ze���"OH]�JK:HrX 5c�A�"O"��w�/`��bFD�@P ��E"O���2'�6WW�`sW+�*tc��$"O� b,��h��[�l%�@��
"yŐ�"O���s��ZX*�u�X�8B��"Oz�9"M\�3$���K�A
���4"Ov`X��5��تp'�(u��z�"O����O�[�9�`�߂[^�Z��Ik���IA�&�ΰ��A�JVAP"d ��!�$�w��U8@&A6666!K)��C��x���]��I��J�(�FC��S�V$:�)�	e���Έ�RF&C䉡9����N�P�,�fD�,d�C�	n�����%8�p���}��C�I�x�H��F�>v^U
��85��B䉀[��v�XeL^EzA�\�C�ɽ$��T��� �86G4j3N(D���'�VN�����%l�f��pj:D���J	,����S�@�tA:D��b�PIV�!6/A���C7D�,��b��=w��!�)ԴҔ�[�e(D�D��Ӆ�Hth�E�;�p\�F!1D��F�\�L�y��U�<Ik0D�|�K�F�qƄ��ZN`8� o*D���BJ�
h� (+���~$���"D���W%1�^�xQƗ�o�V����?D��`���6t�����S� �K8D�pS��
8�$܁�`�6e1��4D�@����4�B� R���j�6�<D��ؐ�H=w2�2����(�M<D�����4.�\�rG��w9��"%�8D� *Cw5,�pA��}f��ha�)D�$�RAǳl����)�5X~�H��,D��IvjK!T&¬�Q�d��F�)D�˗��?�ȴc���u�,i1%"D�Р�+��x���@��v����a�HbD�5�Obٲ���j��Y�Vn%LR$���'�(��O<]� �E��v,��k�$Z3�BU"O\�sB��m?�00�Ƕ(#lZ�	q������? �>�SG�?9���q��6�!��u��u����#QI�p�Յ[�qV�Ҍ��*�g}r�V�p���N�:���&��yҭ�8y�Ҵ�����4T[����?�d�'C��P�I��|���0�U>��	�	�9���`��#��Ą :0��%��'�ИF�N�L(!��n�m�0BŜ�X;�g�#qO~���IH�S�=F�v0��,A�L�J1�O<t.0B�	��L��S5-�+��w�-J��LS�'c�"}�'�6����
�<s�Tـ�FJ� �'m0� S�6�^�����|��H�'0ģ媑�<�Τ�4��=�ޅ�
�'�Ƅ��Ώ:]�:M��DF,6�@�
�'��b�I����)p�E�4S��
�'Cf=P��ְ6v�;�%D�(~΁I
�' hk��Y�,�h�-� &��p��'*�`b���_�V����.���*�'8��㬅�|-`�Ē���!�'i�@7�=��*C��Ů��'�z�J#��!�AP�	�(H��h��'�`�����;��A���Q �h�'���x6���(a�e�HG�'C�c�'%�lKwA<��U�"d��+]$���'�v�Q�MQ;"=C�H;��M�	�'�nT�ei�����)��8��I	�'��D���7܂`�-��Xx2�b�'���@2�ڂMd�=�Ţ�)I@.�H�'׺�PM��}B����E ������ �@a#�/f����`@_�6D��"O�a��^�R�R����an~�S�'��䁾s����%-��6 ���w�!�$+"z��(����n�C�Ŵ:�!�j��0{��J-B��fN�[!�䘆f�H��#�%c���@�7�!�Ĝ<]@�isȔ�F�(@ׇn�!��K�І� ��W�8���Ӈ�@�!��_fgp�k�a�T0�L�!��Q�tm�q{��$�P�B�@��^^!�O�&���㤊8��V@�iN!�$ջi&d����	l 8M��.։.�!���X:����U."��ݳ!#��!�$��!
r���cY�>������j�<	��]�ņQ��`D�B,h�i�]�<yP+�J�B-+bl]U��Ej�b�P�<�&�ީR`	����'��Tha��u�<i�ȝ�>w`p��ȝ�k�4�b�^f�<�a��CK"�s�%�>b���c�KZ�<�"�Ь;�p�2�mW�y�����j�<��Èe�05�/rD���m�<�d���B����ũ���x`$^�<Y��(w�D���kؚ#:���D VQ�<����8��p�v��s���*"%�s�<i���-iORlY��Y�X�Z�hr�<�q�C
uz�p雿>�Hh��m�<w�׃/'^=�_829�Q8G�p�<����;t4��R1�ڱaN��!%Ph�<1vMCzUȉ�㆑�p�ɳcBy�<1���@ѪaR6oR�ʐR��-S�!򄚟W���;�/K"΁��ŽR�!�$	̸�$��[W��B��@�q�!򤄹�đh���c�}�SL�9�!��$�l1(K'��œ3���97!�U�~,�"g
'��A��Ś�!�$B�b�V-3E	
�Ap&%6!����&��"͗�ܨʢχ0�!�$ֺt����E��(
��X�1�!�YL������R5ذ(V=|!�d< >�C��U�V#l���酟/!�$'5� ����!6@��B�,=s!��Bw�D]B�fΒC~��s�\*S!��'j�ι��!P����0u���1�!���5hb�B`�"If,Wޅ^�!�D�;fA�X4�L:jt�B�1�!�ԭl��H
�kېo��ƄW� �!�/C���poŀ5��,h���(K�!�DZ�(E�b�|ƨ�CШĐ'�!��%���7��1m�l%���1�!�D/.X�{��ޙ#��	:d�L�8�!�C����0� -�j͂�� 
"�!�dGB7Lp	�Z`T|�"�f�!�Y!l��c��\3s�@�����yB�[� - 2O�+|��Y�8C5�3D�,I�HI®� ��)m`�2#2D��ՉW#��te�I�O����*D�����
}����ԭ'$\u�P�+D�����%��H��k�N�*�rf�(D�\s#Ο<7�h`Ğ)	���d�3D�@c:V:�k aR,`9�(���&D��I#b�ZG�9�7j
�^�4�4F%D�$�@ԾD X�' I�/�ES�#D��2�慐OXf�;�Ǟ;k�\s�n?D��� �Lʜ���E&B
�L���<D�� <hzGD�>d�Ɖ{��$^jň "O�U�rF!�b��V���Q��D"OX
A��r&�|;��\�c���1"O��/A%�*���۸J5r�p"O����`U-W���x J�F�ȕ"Oe���H��`˱c�6i Ā�v"Ot������H��U�����yGJ��f�)M��aբOhC�	�)����GƃV��4A"$��8C�I�Fn��hPJ*�� �����4C�	B`�C�
=��"� ��B䉐nb���� i�y����B�ɟd��CqC�8s���/]5c]�C�I��8��G��e����&5k�C�`&�%�"N����゜� :XB�yӑ�Q��x(�sb+Y4rB䉌n�xKrl�~X 1�W膐N�NB�I�{�f�k`��9Y9܌ʅj��?^BB�I����.���"R��Y\�B�IK�"�0H�]Vb�s��X�_q�C�	U/�8�լ*��*riV1g�bC�JYFr1�B6FegI \J(C�	�I���[D�c�N�5�U)|C�1�)Xw.2q�v�Qr�F�B�I�D��ͳ�!	~x�4$BSB�B�0D$d�D��lϢ=���A�X��C�	�N*bP��M֭zw�9�5	Z"	�C�	�	��pƆ�q����Df�%w��C�/
�NH�6e��DrΠ�P`�-AafC��t�&�� ��U�,�J)�C�I3�`�:u��#�TY�Ȉ�2+�B��!Pb�S	��,K�DF�j6(C�K� ����W�:#ĩg��B�I�f+��-ֆ��=p#DجB�5#��Ph�EU�˪P� +8cn�B�I�"6��`IȨ?h�\#e".B�I7)0����0�N���+(B䉒[)hB�ۉ"u�X�@�,��C�I>wsְ����7�0�J��_�22�B�ɯJ[�p��!��e��h�M�pC�I$R���V��0#C�u0���:%�xB�ɯ�D�2 �Gd� ��=~)�C�I�j��E�%Z'v�N
ԌB��C�I	���a�� LDU�5@Ԋ(�HC�?mm��)��66���&MR?�B��u��ĐT��@����R��1\�B�I.Z�hpC�oU�(�	caE+Q�B�	MF>�#�BAB R�(�ȅ�z��B�ɚ!�<�Í�c4|�Q
3q��B�Ɇn[�)WH�~xN� ��^�7�vB�	�,4��k�Q�S�D��X�h�lB�"
za��� >mn���4B�6B��.�	h��t;X�S���?C B�.C�^qb��>1�	�A`�C�I9��Z6/��Y�B�+��x�C�ɩRRJ���C�u�Xp��ܵI �򄎥]z�d�!�tL�F�<�!���7�I"`j�&,��@�C;�!�����*�A��0!;��Y�y�!�U�g�MѢ��`����3i\�!�)o��c�H������蟣$�!�d�8Dp���(�"�� 3e�(P�!�D��+��UQ0�F~� 5���[:MM!���V�Y��	:v %)��zl!�� "hb�:E'��(��)-r�2�"O�9��O�9t��1��>u��yv"OB����Ы@�"�!ŀ�wE`�!S"OPD#��
�����`9����"O2�z��N�$:�r�(*� ��"Oܻ��=U <��W���i�"O~��i�0+�
��2l�+HP5P�"O��2���L&�A�J<9N ��"O�4{�O[`�:��P��76�>�{U"O"@�E4}^z���C�t`��6"O>�8�o\\)�5mњhQ&pz�"O��y¬�0vo���@�(�H��"O0�`��V�L`�;��=��(1�"O���"��sd0	P�V�4�؇"O\���OG�m��a�a	�i�ł�"OP���)�-f��0�ڂ
ND���"O��Ģ��lPܛD O
}�p���"O�I"v��56�x5*e:4�$ �A"O$\9%�ڊj�50F2CS���a"O �1D��=� ��s���҅"Oм��!,SvQ+`�+����5"O�Q�l3c��Iz7�X;��+�"O:<s��,��)��n׏n.�Ж"OT��1m�	p��x҇m �X�)JR"O��x���)'�,��,۴ql�A"O��2�2[��Xk�l؏&lvq�"O���v�L�GpŘ�j��]N�G"O��j�%�9.H	V�,�
�"O:Jp�̐����I�4����B"O�#a�VQ��JH�_��H�"Oj|+�"�9I���x�iֈغ��"O���S��k a� 4����"O��Y�AC�F�<�{��K�U�Z](�"O�0���֣0�]�$ψiu���"O�0�T�O<:8vp�s&V���"O��ݩ4U��Ѡ�� i�µ��"O�0�M0Vu�"Ȱ`Ǧ	k"O��i��1_�|�6��0��Y�g"O����k�	/.t"D Ǯm�.��"OԸS��ӽec,��/^)&I>ܘ"OL�� �?4͊�� ΄,I�P�A�"O����	�%t�k�G &^Ժu"O�Q�cR��Ȃv��u8��"OrTa�+����W0�x*�"O�A��&��_D~P�$�
�X�XK�"Ol��B��HK p���U����"O@�4�Dք��C� :��j�"O�]�G��t�l4���E0,-�"O!��鑴c�T+�'% ���t"Oh�:����f�h������""O���t�Q�ώp	�����Y"O��P��6��b�� V�ؕ �"O���RD#M3�l�p��
R��7"O�ɛE"D�c:Nq�"�ܶ=_<��w"O9ه�N���r
��d��H�"O��� �F.S6E�3�[�F ��"O��zF+���v)�E��LN���"O@�a�ɔ>=��h��ù0�kW"O���0od>��S�Ȋ3�v�S"Oܰ�1�)n9�RB-՛0z��30"OH��1$�����̕c�is�"O�IKf+X�M�����,L�N�l4��"O��`��Z�^������^X[�"O�@q�*�?X�]���
�n��"O� ���@N�A-�&�H-�ms"O
���`� �������&"O�j��,if�c��;��"O�Dď�8' �Qpa�`uyg"O8��� $j4Ԡ�/sެ��"Ot�!��Ko�" �,\�¶$�T"O���䍔)��t�Q�^/O���5"O��t��~��H��/�.���"O<���V�F��iW)l��"OD��q(΅v��[aH
�t��aT"O�a�5����0!���%tQjq�"O�Y۷ֱ:����'�w���7"O&ub�Q3o�`���گ=����b"O���VM����BAԓ>���A"O��������Q�"���l�v"O��D��gR����>����"O��HG�`�D��b�X8/�HeH�"O�Z���k8ԍ2࠙���e`�"O�I��mɌ���oQ%T�(�j�"O�ݱ��?t*���S�U��t#"O�Y�� �_���NF���<3%"On���T�p��� 6�H"O���/֏(.���]�1�K���x�O|9��ᔅm}�XԈN�~U�q�
�'��0d�O�C�%h�&t����'�L{0G��V�I�l"p\�ِ�'�	��M'(H��ڿR���b	�'�8)�̅.��lx��^�D˖xB�'+`�[�	٤?���]��2�*J��y��c����+��M�%c�����y��a��b�d�"�I� :��C䉄`�Ε���X�Ά��B�I�_�2'	�+i����;Y�&C�� 5��T�r͌IV���EҮ`SC�ɰ]v��5�ϋ/�Y  �'����<�J>�ϸ'P�!c�	��Oeܔ{�S,��0	�'D1󣄊h��:�nX�dd��'����C��P�-	�>	�Q�<1A@!�]�ԣ�9/ֹ�SK�<�`���g0TۧJ7+�is@�]o�<��F5_�v}�`m[4f�����_�<��O�"+U"�[��\�{n�2�J�U�'uџP�F��~���3��?*��)Fa�W�	u�Ă2�*s`�	�e�z��|�q�?D�<��IQ�4�ӖT�g�<D�XB�M�6^�����Mծr��u[�?D�4�e���?��={�AYFX��p��=D���4�N��jP�k�M0t�A�
:|Ob��y!��|3�xwDOb��s�6�	h�����:��a�gٗ� �H�+M^P8��E{J?Q�ԉ�{ô� �+���rXR��0��3�O�<��ɘ�UI��ŞS�f���"O�h��\ʮ��ժ�M�,��"O���̈I�L�$H��l���ǋ�y2�A�F>�( u((jt8�d���xRI�\��!��G��R%�7�۲s!�d۝g� �BjJ >������%�!�䁛1�Ɯ0�K	�"D�}�f�Ϟ2��OJ���D�B������y.���%�^�,A!���Nt�Z0m��$� g�ݿ�!�[x@ũ&� bV��84 @"_�!���2x��g�9J-P��(4�!��-l;D�(Ԇ
�C˘�C�ț��D$��|ڎy�
G��bG�X�n���3��S��y
� ���F�]����g�2kA�S��G{��)�~��5�"��?��=�#��3'!򤓻U��y9&���L�d���F�K !��j��R;k����F�c�!���x�T؀��
_a�#��V�!��.g����A
u4��ؤ"�4I�!�W�F%4��t*��?d�e���x�!�d.aㆉ#2'u�xJd�W�ux!�Dhf�����%��JYQ!�^MLq�1�9h�n�ʂ�Q�kG!�$�4�\�bT L�L��
`j�#%�!�D�:��a��U��+��n!��Į'�XеbŽpN�⢉ 'm!��
m��tk]
�:p)F�5�!�V3�H�Xt�18���(�2K!�>G<0��蟛n��]��f��_-!�86��S���q���a�Z�	!���7+.|�L�8���K ��[!򄌛v���xU�.vLİ���9a!�D�$T]�@Z7��B]ڔ� ٬x+!�\]�� �ݮ?�x�a��R�V!�I�C4�m!��W3�✨B�_�BvbO:�Qfo��'���ᱥ��r��T"O�1���3@	��9H�c"O��;f#ǖef���s��4�]y�"O4�@J޹��1K�̼f��|0A�'��I����pG�a�B�3TŇ�[^C�	�8 (�Q6h�'p^g�Є��� �@y�ʝ�`r�s ��:�9��<A���SRv.�DɂF�HT@Q$_3Q�B�I
;/dԋJɔ�Dt)�]�[��B�ɏ|�lxȑ@B��
�S�c�֒B�	�F�&m� ,K��i�V��(k�4B�I=���H���:`n��U<��B��	:��Ly �ؑ�:��E��4\��B�I(��HS���J��*�7�B䉑}5�Y#Dd��a��ҲKٳp�C�I�R�09�JX�'�p�ː��4J�C��rʲMK,n*")�tM�Z;�C�Is����T�G���#`��E�n�=çm+�di�IP 9M��;Ӫ�.m	�A'�4G{��TФ@�}���Ӷdy|��"@�8�ybLF1a:�Ÿ#�`���SAX�y��J+��XA6A~4s>�yr�Ԍ5�ȩaޒ0x"�U�y"��Q�B��T��p�8��_��y�(".,<�t��(aTH�x�����x���1:EK��ƨe�|D���FO!����F<2J����=��,�HK!�ޓ���×C�~0��Ū�l�!�d��a7�m�0l�Beny{0�1("!�Ĕ�~��E_�)-"MY7(O8[!�K)�r�/9����^!LJ��'��EC�di�0-8g�����X�	�'�<4B��Y�eqꬳՀG%�"���'�� �J�`	�J�)O�P��T�'K�i�)� ���+�/��e �E�A����'���A��{Xi[JuI`Q�'�.�P�e�Z��Hɦj(gϴ��'���� )A�FC�<b7���`�zm��'wґT�ڤq�"��v���@����'W���@��Z��{�hR68HD��'�5J���0�PF�� �`� �'=Ҙ���j��K��Dv�]�K>ُ��� ���M_�R����L	�3u�[�"O�@��$�6��x�+�{�V�	�"O�]	a�C3u���d��!.k�\`�"O !X��\+�59�k�WlV�0A"O�D+�O�4]�&��#ܛ_bt� A�'���!�`N5��Es��4g�83E$�O�J�>k'����l�ց�(i����+�h �
kI\AP�o� x�����p�	�q��z%��C3-&q���ȓ,%J��.}żA�To�#&���ȓ,.�y�F� 
<t�R��7 $m��t�$��D�X?a�Zy�6��Q����Is�I�
 f�@���=j�7��!�����	�<��$ЯI���I&ESch�)����}�<	�M��L�*�e�ypRt� ^�<a���X�Z�cs�ɒ/t����<����O2T�I��Yy���Tk�c�<��%�s<���`�82j*aq�*ZJ�<�d̱!�:�A"LQ28&�C��FE�'�?�J��!mt��1��-�x@Q�,"�OH�	1���G޴ �@5����B�	�D�P�1uf$?NeI�L��`�<C�	�=N���U��1�\16�EI �B�Ʌ�l�ec9_�q��X�I�|B�I�]r��	4HI�&�
/L�JVB�%{�zI����X���p�G+C�FB�	�m�|8���V	��У�-�(|d�C�	@jN�c@����T:��5IRB�$$=��(�(ĺ��U��HOB� JJ���@:�ā�s˅��C�	#;S�h��(�l�R�d�& �C�I�Uh����HѪ'�Z�Zp����C�I:�4h`�,|����'�M"�\�ȓm�``iq���;�Sj�2q��	D�'���YD�qkRB���?��p��'M��R��6�n�r�l
�:-��'�z\k��K9��X���6��ܢ�'�ͨ���j��aՋ�#(X�'&��a�7,����揫!���
�'�T�`���_�dU��k�$��	�'v8�0��Ґ.�@�S&=p[V�h�R� ��	�A\�@Ȇ��^�𰊥lK�Y�B䉫Mm� ��L44¬iS�	�_�C�#$=��
��k�l��DG�3~�C�	�`wR�X'#]F���A�F�-�~B�ɒls0ui��
�}&����|C�	�DI��%��nf8�����u�J���/�I1Sc�-	`e�L2ՇM�_x��)扪,�T%Z��@�4TBT������(��I
��XD/2k����J;E�C�I�Bx�, %0�.9��@G�8��B�IE����ҏ��6�Jd���E@��B�ɠTڸ���_/0L�&,�4�xB��;]@j�r�1��ó#U�4��+$D����ӧ7"V�§� 	w߬�8��/D�t�1"X�^����fߝ*�9��1D����	#~�`q(��X�<ud5QF�$D����AQ�8\���"�.8g\��E>D������,/[�y�W��b�(뢊/D��Z%����#t�A'��	�.D��@�@�$�u��P��%��,D�d�rDJ o+2]� ܄F��š�'-D��t(	)6L��t�� 4)���'��n���P#��:�U�Q�$
����'+D�� b�w��X b|b���4���W"Ob4h���EI����
��|��)�5S���bQ(�^+�ݻ"�D/+":C�I7
�,(�W*I�vS����Hçg�XC�� HE:"���r)��W�_�,XC�IC����'�2Mİ�]�4�C�	8+U���A�>h���G)ٰ'5hC�ɶ_o>XB�J�9<,A�D��8C$�C�	=
�x0���d�(mAI[!o���1�o2�iD�?^�z�k�6L�]�ȓ1�Q��U�8!و��@��D��i�Vɸf�1z��H􏕘8ɰ��+�:;�LO�*,��.��@�ȓW���I_�Wr|q��DW�<H�ȓ�,�QNB!$7.=����go���ȓ;n�\��a\0>�h�+���V`f�G��7J��if�ڵ�EZX��C�I�d�ԡ*��wn�A�,�0^�C�I3����1��'F��� ��W�8^�C�	�%Ϩw��.����AJx�LC䉳��9E�\k.���f;Ek�B�I�8�O�*}��,ƺj`�B�ɰr�̒�ϓ���I�D�>$߶B�ɂ&��$bg6G�" U�-����$�S�Oc���S����Q�`@�$�q��"O��1���?����@��?�쉣�"O�P�ce�/���1w��D"OnTI�fN�nB���CQ��`�%"O�Q2�ӎMp�ɒ��"l��(e"OP�s��v� \��~�D��U"O"��`'ٮ[�
5��#�N��D"O��2:M�'���Q��"O
�Rْa�z�rǍ�`�H���'�����h�"*�s��z�O���!�D���d힔ʄ�XЅ�3o�!�9,x~�9�EQ�H��L���ΦW�!���_$�u��>v1�u��p�!�$� Ul� P눗~U��@�
y!��ӆ<f� �4,�k�r�ȷ�ҥ!��(8�=�VGU-�>�pgI�ўP���([]>p�R+<o����A�
B�	{` ���:pi�2&�P�w[C�	 f��ٱ�*L%m6Q҅f��%�,B�	%,Ƽz��ߥr\�Sd⍻e�"ʓ�hOQ>��Q���Z6M��I�~��ag.ړ�0|2¡ 2�� ! 
e��Hóc�~�<�j�`�}��a�~�6H��Á�<qI��QB���!�<&�B�C�/�c���0=!H�x��)�bf�>���DD�\�<��C��:}�ɕ�F� n΁)@�[�<IB��&2���iSM�7l�� �e��G{��iӞ@��#�kV8S���s Ю=EBC�!PJ8F�v���ȆI�tC�	�k>F(�VM��� f*��Se&�=�	�'#����X�i�z\{�.}8ՇȓW�����AX�E�p�*Q+�r�B��ȓ�ּB@	��8�6(J!��7 ��O�ٗ舤4U<����N��؄�Y搲G
F�O������эWn�݅�I[~r� �5�\�c7!U�%�@]�p�Z9�y�^��>J�⊍}&�$,Z��?�'��$H�(�d�.�(�Eڋn-fi��'JZU����?Ҽ\����B~��'���)s�_�y\ ��C���Q��� 04u��=I������	\̬9�"O&<�+J.9�pC�b.xܑ!"O��˧%BaI�%���KA��
4"O�1�� X�P0�Q2P��3)��IP"O$�kS�?h��ȱM^�;(����"O�TɆ��Y�}R�	nX�8�"O,�1�Ō15�����;\D�Xu"O�u��k[� S��+A��\X|�"Oz�Y	��I��(B �K�B>���|��)�S�
WN�+𤆍i�
�ӥ�M
C�	-��X���4�w�1c �B�ɯi�
����P"|y6x�$�dM�B�I�"��頏�6Q��$H,�8N~B��3a[r0# �2;������M���C䉟��Ӵ�� ^T�� E�C�Ɏ;||�"B;7�H͒�c����O��$I�#��Db��OWr��S'k��.�!��ȗ.	��%'c4D��,VV�y"�I�6�^�J!4<�J��ƥ%B�2 y��������a-S�2oB�I�=��҆���xJ�h��H{�B�c���8t�,6�$�bV+qL�B��+X��T��#�Ȅ2���5T�fB�'[�D�#�A��|Q��5�DB䉢�|���!�z��i�7w�B�ɡ�n�Ӵ�@�BJX��� �.C�	�1Y��#��u�N�k҇V%%<�B�	6-�l:�f[*3�>�h���=g�C�I,���d���d�2S�L�)�0C�	�mE������".�D�4��?D� C�I7axe;�
\�0�E�$!�6c>C䉓|	�Y�>)�t� �*C�	�%�R�����6~C�@�%�J_��C�I
Pe�����6#��9a�7��C��#u����
V�zZJ��Di�x�xC�ɆL5�S��5:4p,ʲĆ.1lC�%jb4�
���������;^�B�	���Jߠ5`�Ń7-E�x�B�I�1�����엑ڮ�(r(ִw�C��3|��9�-V�*���ֆ��FC䉪D��p7�U�v�9��O.M�B��8�@
d#�-:fqjq�M�x�C�	�;U��jQ��55���c̣/���D{J?5��m��0�fep7nY�E���<D����aȸSYt}�B]o.�l�  D�l��G�e��9��h�O^BM��+)D���G�.x����>�4)�G
�O^C�Iu���8c���Z���c��� B䉼��<{�a�$ ܐ�G �f�C�ɀ����"��[Mh<Y���C�	i��#*	$�D(���mIC� �A�K�phδ5��1OBC�	6"ޢ��CT�r�:�I&i��B�	�7�:��W�[�n��p��y�B�Ƀ+��)��%ҙ )�X3r�O�,̪B��;"��hk�+��E�͊1I�B�B�T��2��:��5� �˘-ŸC��&3���F*_p��aqV�:~����5x��4��B48�h�S�`�3����ȓ�TÖ�� 
N�CE�R
6c��G{b�O�Xࣗ	��8��FMχ"\ �'yđ$�I�yZ��X�ʙ,F�N;�'����O�`b�8�h�hxx���'�4�R�c�5�<��e�M[v�E#���)�� �Y��N�r�t4��$ɜj�z�*O� #d�x'��"��B�_:����'�vp�F�?L���ǦPH ��OT�2��)QT�:�#t��ss"O.=��K0�����Β��-��"O�u���P�J��Б�0Ԋ�"O<ݰS"ȏm���C�sN(��"O��a�B�ܴCE`�kCf���y��U'y�᫶��$& :\�oX�yR�� ����5*L=�H=�+Q��yˑ	� �ůJ<jv�ۣ+���y�h۾,��Z�S��t����.�B�I�R�V@{sKU�=B�@DN8�JC�ɞb{�Q�I���QI�� �bC�ɖIkf]�a[�@3�E��Ě���C��O��q�"W��*��rTVC�I�7��h�GP,6�։	�h�+�fC�	;b��$�gN޿
��p��XC�I�D̕1f�[�]�y�r�YH�B��=6��U�&L��t����˥CC�ɿ^�.1H����ѵL6_��B��-S"<�iKn�ƕ� ���B�	:s�v����O�r �(� �LB�	���%2�(T����%B�I5n��-Ha_#����6&TJB�Ɏ�z�jb���k����:�(B�	�$(k�!Σt���#7̏&�B�I��
�����7W]� ���	��C�*����D;yz��H� �B�	6a�4�h!˼),L�����C��~�"�Q��4t=���d(V 4O���$8?�U�6-��!8�GQ:,)�X:a�t�<ib�ü���X�X���(��[[�<��ì� �)ŧ�
)|1�Y�<17I�2ҡ��.�(��`EY�<1�'@�[
x��D�0B�2� mL�<�1�>y��hr)�,(U𸓷oKK�<a����(���Y�]D�%�f�J�'[a�B'/��Sa� �J|�w�Z�y��S�p sՆF?�F�QF���yr(�,���o+0���h�	���yb`ӀDG�R�3y^�hr)��yrK\?䬥�ׅխ~d>��i��y�G��P�a���\5�( p�g���y��L�"`�M[d��q�����y�Ǔ�l�X0��a��ڜ�y���KH(\��I
)�yQ�̭�y�"��*�b��G~e#r�_��y��G(g�:���N��I�����V��yr�A: ���6:lz9 ����yҎ!Qȹ2.3L�9u��yҀR4�tx{a���Nj���i��yҍW*	$T���$&B`D�1�݋�y�#V����Y��N�SY|9�g��:�yB흯`���[צMM�=�F"�y2J֏#�¡�4��A�%�dH�#�y�"ߧ*��q�gǍ�3�V�S4&�/�ylB�U4iذ���V�FPj3DǄ�y�.��f�:T�B��U���Hd�5�yb�B�b� "�%�-7�A�	�'�^(ɥ ��r��-�-�����'�黧j��m�5+Ĕ^�a��'ټ���S��0���Bd��'�.��&�=61@�0;c�x���x
� T��b#�X�&�;R\:�k�"Ol4cr��	ru��3@���\W�e��"O
 څ�K4��m@�@:&`""O�4i� 	�Q6�Ko
-�*�zp"O���'i���2��C�Sn��S"O,rSX�Vr�*ݝUl���W��E{��)I$��c6Ȓ����Sʐ5�!��s�JP�#>F�tG*Q�ad!�d��F�����Ǔ�0�(�(�ɕ"�!� &Y��xt��3�2�:�ԙ�!�DC~���CGBњ	����ֲ&!�D��Tz�٪+��Dk7'@�g�!�E�bw���$I�,hŠh���0{�!򤆁�^��jƽ4��lC�@�;0}!�dɞ3l*��uB�;�t��t�B,!!���6:�N��@g['{��<�� ϸB�!��ۃ��A6�Q%�}X�  m�!�d�w�U�eێO�� �����!��W�x�`�5�Z7(���ct�P�!��ѮoC>��E9r���h2��t!�DIV��5��aĶ<���+־�!�D�����0��n�LJ��M��!�Lv��RĀ3oȺ�$�(�!��+wm�ԃu���
@ �,W�!򄐯}�N)�"�ּ�<�`&	�}!�d��laL��Ј
A�:� �%	�_u!��{%��q��+a�{���8jc!��w��c�ˏ�`S"�h�hۈ��OV���NXŖ �".�+,#�D�[�P��'�Fy0��_tDD
TEl�%8�'�n����\�@|�g�;��	�'9B)	2c�o���&e\?n!�e��'H��9%��?<����a�bL �'�L��K��{���r0aI�ke�`��'�
�Bp	��&�Z��Z1���kO>�)OR��	H<�eB �0hL��Gǀ���IM�����P�&t�� ��-c�����<D�����Ɓ7�0�X5�T_���x$:D�\�0.H+T��̪�H�)��`+9D�X	���-=^��Fk�&u��2��5D��W��6�Iq�J�X�����-��<!�' ���a��9}B@9�懞�Z���$� ��	60�H���@8#�x�s��'�T��0?��#��$���d7�l���A_�'?axR+ۖ ���1��z�޼���2�yr�p�4����t �c+�y��f�~M�@��f��	����yh4a�v�#��
��Dh��yr,	}���
�I�Y���8�䓏0>��b�o��-H��`�3F*���"O�<�5�ơ��:���}���"O`�e�@#)���+��B��kF"ON@K!C��.<���E�kJ�"�"O�"D��,
��#�H�]E���"Olx��ήv?�1���+W:�H�"O���D�vaS`�0[�jxq�Y "�!��Y$]^��Rh��$)�!���,�!��$V��(x��\�#�����de!���p>��⋌�'� ���,�@M!�D�s}614��=U�HU�֊��I(!��շ*G0H	RÁ:]k<	ʴk�2+�!�d9`�z��c�BhB�,̨_�!��Q")/.գ�R��`�v�M��!�d�?��,��1}��y�F��'0a|
� a҉�0
܌���ó���2��'�ў"~���V1sX�4*�銎c�ހ"�+!�y-x��x5͕4Tm�șR�
��y�d�Y��:�lC&A[��E��y��.�d]��!ݪ$��Hk���y�eW)�L�Cg��Tr< f/�&�yrT�$F��:B1�1�%����?I�b�S�5�FI��T͒�	�cۦ���	A�'9�1� �ݔ⒮X�@.np��'�(`B''�#H"����́;�T���'����&g�(�.�2"��5`�'��I
��A`Z�!�f����TJ-O��=E�t&ҭO�H�t��y(�:6�Ǿ��'�az"'��`zD)��of`��ZH$@�'zYHe�B#�bl 6�[(%d�4 	�'k"�p  �4��d{��Ў�����'�	�A�T� 銄(ډ^T��C	�'�pS(�:��R���R"(@	�'Qd|AC�ƱB�l�C$��+DS ���'�����C�Ol����C_��1�'P����2n��iǐ6���
���y∅�H�*���
"M��e�W�ٻ�y�� ?`|l�b���f�Y�W��ybI�q[��Z�^��ar@���yҠ��n�Ȍx��Y�$� 4��A,�y�@�v9<�F��&�z�M�*�yNV'w�1�Ff����E�P [��yB�H<�Rlb�Z<p��X &�&�y2�%t���߼7�`Y�,�y��V2^�,��e�ѷ3+�
&���y��r^-EL�b�H���D9�yR�<	2$� ��R9�XH⯔��yB肦1�H{@��CI���	�/�yҤ�,w�Du�gcJ$A��!����!�yR���<M�'�D7B}�����y"�W�?~�Rw�ٔKQfɱ�-�'����'�>	�)a)t峲��y�@M��h�O�C��C �;�<1l�\�!.Q�>|C�	�-�)C�*�X��!!Q�r@.C�I�W�ً�瞞Ӫ������C��3~>���	��K|б�&N@�B䉲i�VS��ӝJ�n�ڂ�V�O����0?�,x-����Q�!*p���DNx���'/�pǁ����P��L� UP
�'�hU���(D�|��e�J\x��	�'j���@�&�ɥ�W���+	�'��p�Ĥ�0��3��
 u;�lP�'��$0"��4�� y@Ѣe3Xh��'��q��oU$u�VY�ᅎ5:�
ϓ�Ol���]�J��M���G�a���)@"O8��O^ul,hI�R!�ީ��"Oڹ����"C �J�-E����v"O�ҧ�S ��y�F�]�(�Դp`"O�$J昡U_�i@���cq"O�TH�Ղ�`���-OpH���"O�j7,�	 ,�M��B�&v�IZ�"O.���+�mC�d;C�RUX:�jF"O6�2 H��u�D����ON���"ORm;�h~������L=D�����D�,�^�Kd�C�6�z"�8D�|0&�@�U��h! ��^�.Hxe�6D���@�F�
�Hc����P4�bb5D���������D0sj�$W�w��{Ҕ|ª́kU\�9�BȾ[T�䘡��Z�ў���3� ����˙l�����֏-4B@��"O��Q�%0p���D� �8@Z�"O����$T1�
��P9=~�[�"O����Z;M=�!�/Y�@�\�P�"O��A�#00���Bo�c�@i
�"O�]�R�Z����O� G�83��'ў"~B���6BLDS�$2Pࠋ�P��yb�гQ�l����62�>I!�N�y�ɔ�%���Fo�.�f�P�W��y2	�T�p�:�޽��M��y�H�13�nQ��ŒM��9��'���yBd��$����(�+>�� #"ƈ���=A�y�틳9x�б�J�L֍����yRŒ p�� �I�[��wIA�2�O��~�p�i\�#�v�!'
'[>��ȓo�:�XP�Էd���Ҩ���ȓ>�بq�R��*��N�o�v�ȓI���`���xl��A/I�d�Ć�J(d[h˦�F��Ă��_�YF{2�O#����1Y��`;����':Q��"�X3@���ϖ.���Y�'� ����<c���[�!43���R�'q��
�G� ��-���T?E�%[�'@�)�Lso~��C��Xt}[�'��Eψ5��D`�Y?2���'������Z1�!P��.��њM>������*��, ���k�$m��ˬ��IS��Xk7��3]�P���ݧ+�n4�=D�,#k���lQ�
�*6��T�>D�`sE=4����C�<�(�D"D����)�C��qD �3�e�t*:D�xZ��Nb���K_p�l	5D�,��]
��ly���6 v�˃�3D�� ����_jm���D�_G:���i1��#�O4\k�15��81p�ɂ�=C�"O<���u��@Wk8��R"Oȼ	ǃW�XMpI2�U�\j�[ "O��0�H=7��Q�
�p"O�����j����ԍ
 DYH5"O@�oR�<�(д*�l�FiA�S���	��H�?�}��N�a��0SCqNl����f�Q����yR��0��2t��1���f&ɇ�yR�]=~h�E
vmJAlԋ����y�"�{�e�aӢj��Yڵ �*�y�`P8%jR�f�Å]�ny�E��y�!=vD�t��J^�l�ldb�
�t�<QT�O�-��X�������o�N�<��g�:���U&� &bP�C�Us�<��%[���l��E����ЧFm�<Q�._�p��IwG�{I�X�U�DT�<�RݡD���C�C��I,�X!�J�U�<х�I�f}c� z��=)&��T�<���@���L�l@��CJ�u;!�D� ���7�̌��U;&��1!!򄏴e��m!�U�v��,��O���!���e P�c��6c�ᱶ�;�!�]� �x��G$�1���xY�gx!�ۀ@sR墐�_o�>XӠ�N%k!� �������"Vc8$�C+�Z]!��Q�(�	*R�Q�!4� cu�ӞY;!�D֗.��\�͙�@]��Ɣ)!�$\�P�����kY�_����0ƌ>p�!�d3".HJR7_��t�sk��,�!�-K�ZT�5+_�8	Z�$_!�� ܉ZC��*���	��P�ļ�4"OFM�&���"9{r�̄,��]��"OX��f)�oK~� �E�P��u"O���4hщ �
��S�N�F�^ȲW"OVY�T�]%�pTZb��3Z���"O������#���&)�D!*-�"O��c�.�7��p�2��P��@"O�=K򋃪fp��QƦمW-�h�"Ol�0(���ً�E7E�.!�%"O��cPL�{��"d��D�����"O��dOA"/���p���\~Ɛڰ"OL0��#�~��s��gs֥	�"O��Do5$ni�X�>ț"O ij���s�1�4�_�c��q"O�R��]�{�u!� ��T����G"Oh����ܢl���#0��?<����2"O�$���x]��y�f����ȗ"O&��w�Þ(���Z�$׎K�"X�"O����Ah��B�Rm㚴# "ON�҄�b���G�ZE�"�:p"O��а˴GL�Qs���6;r��3"O*A�f���j���G�H�t�"O6�R[	ߤH���>b(�K��M�<����hT����"���%f]u�<I"�"yE2q+d�	�j�����Jq�<���<H��T��EC�<떥�j�<��.�):�	j�$�2J����{�<�a
G�e���)#F�.&r�UKAĞx�<��oبh�$QD��U�h��6�[�<ɶO:' ̃'d	��ڽb  �`�<Y��ز!)(lk�]F6�qu�H[�<!�!T*J�T� cH�2nf�)�TY�<�wf�"W~�}sp�*�J<��i�X�<�T��k���I5DT36��P@�R�<�P� m�ш��O�8]�v��i�<q��K):7�B��-X�p|��Gz�<�6�=	2�� ���J�K���t�<qЎU����V�Tf��7� I�<)g�4@��B�u�vDC���G�<)G"�bͬ�FϬPb�*P�C�<i�$ݔe�B�8���BC䫑C�<��Ψ=���gl�1?�XT
0�H�<9G�q]0�A��)R&T����F�<	Q��!9nܨPe^w����� Rl�<isY?gO2�j��	����`G�r�<�⁁�=@��)�-w=J�%`�v�<! G�.Ⱦ�Pp��&m� ̹��n�<Y�H�6��P�_�<]����f�<qA�B��eYԮ�&�\����\�<����550���g6�p��]�<� ��?�$�p�<z��EY�<�2���F��Y��m9/f�˕eU�<�j�At�E���݋^�e3fkQ�<9���[i����� 4�� �ČSL�<�1�ʚo�2|�@��$}Ot��$��s�<��O�p�쌳c,�!6�R�2��Ir�<A�jأx���M �l�so�o�<����{��1rRLў}�Ľ(��G�<�A(i�N-
��nM¹��C@�<鲁U �օBD�N��X�Q��1D�xrUď�r&*
�K�e:�
�//D���e� ���m��ɵ}��JV�1D�8QFF�j����$i��r�3D�H��CG�Tb���C��H��а�6D�� ���@9E�h�B����ss"O� �KΙP�9��Ƃ]��`Y�"O�}r�	�[<)�@�FX��!:�"O
i��k��IPU���
�h�"O�<z�h�x�z���b�LY�#"O^,���8���EDT�&@�#�"Ot�f� p~�$�KK���D"Ol�*T��/���"ӈP�6DͰ�"O���7ʺ'(����f@t*"O�!����>-��F��Dy"O�=fJ7lR��FET�Lat��d"O����yq��Z"�Q�]��R�"OЬ�v�#��R�BŵdV2�R�"OF�'჆Q�l1sĂ�xL� ��"O<ّ�[:W�>��@��bD� 7"O�LR(�m���i`L7:9d� 6"O��2!�9ܸ���ˋ�8	h|z�"O8�٦jP�A���kE�F5(�H!�"O:�F�<9�� �1I��(��B�"O�P�@L ˖�"��>!����"O*�@�_#f*��ݷ�̫�"O���㓳pj\�����6@LL�#G"O�u#s�١v�4B�^�C�F�xT"O���w�V�$%�eW��4q��"OԱ�吢z���CD�pf5��"O4����n�j�y�Q�G$�5�@"O����,�9rD�V ]����F��n�<����>2n�i����V�Y�E�c�<�`�L\Cb-��/M�n�7i�]�<��M�,!b� ����97H�V�<!���%�\I$o�3E�R�+T T�<����~-z1x��*3-��!�EHu�<ђ� ��ݢP�	(Kst��!I�<)D#�"%W��qHڞ|��D�E�<��MG�u�pE���!f��D�^j�<�"��F����F��9J"%��ƍO�<	�Ӎ6Nl�(�o"Ep"��H�<) �ʭef΍��O�N6lV�n�<!��70p�jH�%��|s5d�j�<�l�I�x�i��?nT�u�qύd�<���Û*k���bƘ*��ч.�F�<Iƛ.otv\p���s6�e�te�<	��{=��!���
������P�<����@��XB4��!$Ɇ� ��t�<i�˒;\�8�Q��6�H�ԨTl�<��
D���Sn�!O��a��k�<��w���y��\�,ze2�A]d�<	7&�T:���^+\�Z�-Pb�<�e'�,}�ԁ�
�)x��ih�^�<�Q�?�}qѥR ,�}�`�PV�<�&�H�i�	rON;Ur�(���Vx�<9!�ť9T�)�3��M�ŏ�i�<����dV'��dcȡ"t��y�<q@�C�D�d'�v��Q�@Ox�<�� �.>�6�8�!�q�D���)2�$�W�V=F������b�&q��ne�}S���$
�F�`Y�ȓa��k$ޙ\�Z ����6v9�Q�ȓU���c�/�M�|�,S2^�Fن�/�pM3UO��	�y�С]0B!@�ȓa� ,+�تl1�-!A%԰B��!��^Ax;w��Q��A��%��N�6X�ȓ p0xC�Y.1���QMׇY���ȓKkt\zT�U=g�Ns0��^����S�? ����nCԆ��$%E��0DS"O�����*x`Q�U"[\b��@U"O,��Ԅ
�R����L?;E(s"ONA�ej�� �I��O�=8LJ�"O���⨌�,Dx�s�M�!$�%�"O=�0�\�Fy�Hr0G���T�R�"O�DUAZ�`�x)���ƹ.ɎPX"Op2�I?S0�:c�k��:�"OfIk��L�ƌ�*Z�T#��P�"O�M2��J%Ľ�ų=(�bs"O��c�U�� ��Cf�hhԍ!X��G{��)�-z��J孁�1���1�r!�$��^���V�vͬ��V��7e!򤞹J0n���O��)���͝/gT!�$2v����CK���@&����v�2}J|�'���"A<����c�Va1�ѻ�'Kҽ����n69ʡh�%L	�ٴ���}����P��K]�2��
U�q!5�>D���F��5(������'��@�.D�p�@6�}�F����G.'D��S�U��.�q��R����e*D�H�P�V��J�mM�'�f����<�	��`5t��8�~1!�˝�f���D��(�X��(�7L��X`� Sk�(B��0>��2����\����1hD������ӧ.W��{�M��l8��t&\+IO�C�	�8m X��Ş�}]�!�&ك�C� 
O:ћ��]�=[�����l��C�c�D	�!K�}h�|�wj�M,x���dq���>%?y��dP*��L�'�-n�:�O��'BZ����@��Jd�E�e��K�'������)7�@�F�IKv�8��$8�2�v\�s.2M����"̈́]zr��ȓS��加i�><�Ycq+رn�� ��=a��I��1U��L�pC����ȓ��aC�mN�%����-�,w������A���@�J��q�ƅ:����U��B�/ґ��%[�+C0ʎ�� ,O�QA�oҘU�*�k��wg����"O,�J�)�3&zh��+��VX4@��"O`����<	�b�B/I0i�W�K>%�$�G�G�x03oP�l�0c7D��07)@x�����Z�UubT9梟��Ӹ'�L�"h�b}d�9�Ν�X�ݘ2*O ���Ʉ3�<m��@^�Z�
�c���
�J4� P�[�
�hS��B+�����g�d�<���̧1:&H������1����<a��*mܬ1��)N�Z`���w�'��?���i��V-�q��"U�0��đ�&4D���VH�<]~��D�����У0D�@���.?[L��)Q%z���A#D���qέ4eZ� ���$K�*�&D��q�NN.[M����сB6ECf&D����۽"դy!�ї
�l X�/D���7��#�Da�	N4e�dZG�-D���I�4H���.�?0�+�A0D�,cs!���:����ib�R#��>э���4���#QFv�����^�C�ɕ@�P��(	�F�	�!�O�㞘�� V�Rz��I�I����[>4_�C�I��MQh˭|4����7^dL��f�$D�<��8yq$3p�(��SB%8D��0�`]:����BŘp��@A�5,Ov�<A�D�(��t@``��R`R|Y0��i}b�'l�|
� @Y�v� (������lG�(X�?OD�Ic�S�O�$I �˚�1�.��2�Ǽ2\\2
�'0���oP��`B��%�,)Of�5�Q�b>��vD�3|_F��$ �;t4���?�O�p �'�&����0@�����9)4���g|yr�'*���$+Q���=�^Q%C���'���&6?����Ξ6�H��A��]�āZD/���y2�|��d���VdPlRA/;�������OD����	.�,��a�H9D��0"OjQ`��|i�0cE�
6ec"�'U�$�.}mL�6�[5�d��b]�!\!�D\�U_�d�)C�t��AI	XO�O������~��/>
�w�W�O<���'�H)l���{
�'7�b�E1$G0qqD�Z>��s/O�ʓ��S�L��IA�:}xL�ؐI�7^[Tl��/��"�a0l�4̱�^k��C6�çF	�'��|�$כ?D� �Y��@H�X��p<�N>a�O�p �>hw�*rΛY=��P"O"���Ǥ�F�9J����I�W#�?�z�)��5 h��UD-N��3D��I4�S4����T�1���6D��m�ȹ��`���b4D�\�� �=R$%��<Kb-�A�>!	�Ic�X�T,nq~(��)\��Q��	ty"��Sa�a4��D���e O�y�ȩ4ȸ�h��W�=�8 {d����HOD�=�O�|sSc�Z �lC0Ì�Bϖ��}��)��$x&��sI	8	h=ʕ��2��d�[�'dўh���T�N
����Ѧ�5��	��HO����0>U8��6��| ���ٟD�!��ܭe��ѩB��e�(l2��Y����F���e����G�>b�t�p㞮�y��4�&	1���3����1�F��yb��;Pu�5`Ӽ3���;q燦�y�fP2BԀ�!/?f�r���&���8�O�`@�����u$ˬ��cp"O����͢.�X\����+��t��"O��	uK���ݢ�kO7*��I��"O���D�!XXiH�� ?L�-���'��O��Q$K��S��|J"��{���h�"O�����\�|%bQ�f�
��0��6"O���b���.u
s�ZJv���2"O�i�P�]�>��LJ��ڧ}�̉!"O6X�Њɋ5�f��5����ܚ�"O�(�%�I>$�r�{֮G�r�f�q�	^���i96�"ɛ�A��^�R�����!�d܊�Zq�e�׭��� �
/b�!�ڼW��7K��a�<1�D��9kca}R�>)5��2<R�
�鞖�����\��?�(O����TMIx��ݮ�̬"ע	L!�d� -b�ٕB�����Ƚ~?!�DY��)q��D�~�����`D'Q�H���'ux�S@Z�%�,��c��'gxB�d6�c�[${�&���D7��C䉧wa�+P�
��-�1DZ�HpB㉢%1zı%�U� [d�se�T*c���ȓ$�ze9�@�%2����`�"I���[�'h����X�	�A��ܱA�ux�'6�`�ú$Ǯ)@�/\':۪0�
�'=@e���iO �RWgց&���:�'m��O��<�8pi�m�=���(�i\�	��?��}�e=�S�8 $"R��4*@�q`$�S�HzL���1��-7��AK��Y3A��m��OY�
���]��朢 '��A�GN�(5��=����� >Lې���l\��&ɼE��mkR"O>���و6�4I��l@���h�'���9H��{�a]�(-�T01O�74[2B�?T�6-ۇ�����@V#
7&�B�	'8m6:탪1�x��-&�C�'t�p�s��R@/(4��	מC�	KFe���eF@��۷�d#<��A9�S��<.x�Ĉ���8&��3�y� �W^�	�`B�tw����Dܩ�yR�)�'h�L��g�=>��Ɗ�b ��G��TID�ՑF� %�D��{��͓Q�
��䇫C��p�"�.!gJ�ZE"��Ha~�X����Ȅ�21��
 ��\)�K(D�|ʑ'��vi8��G"�P�`'��b���'*fbu��@S�z��$HZh�݄ȓ;�J�sD
*OSH\����	�j���`8�8$�5y�0ܐ!kK%=V\���H�P�RHldp�h����R�ȓ(��:b�GR'��8�ʎH�͇�>;���P�(0�(�S�R<|��ȓ,����+ԁ��z�
7���ȓ.��xR4��4�U���j�>m�ȓ�I'�ߙB!j�y�o]�V�F��ȓZ�(���J8�D��.h��+�"O&(�ckӨc0����fA%2�L4J%"OjeZk�-c޴�R���"O�	#3�'�r�0� Jv�)%"O��1"�H?sF`;f ��L����"O��١�՛Y�HQ`C?p��"O����ڨ3�
�:R�E�&��"O�L⁧W�6���0���R�"O�djqI�]
ai ��&RPЍ� "OB�81i�g1jI!�c�97?b�Y�"O�x��&�%;��w�@
?ʔP "O�Fhȱgf��S�n.Z���"OH�)B$���Qd��H�: D"O�q)��++�����	&h̥A�"O`��HG&bk��W�(�0c"O��ڠɛ�Xz8Ԙg��J��	"OJa�ƾ<2���p�K�#+���"O�0b��wC�tYc�S1�Pb�"O�j!l�+=�pɳ`�q�j("O	��@b� ����D "����"O`���ǖh�N��EƐ!�r��"Op�B�\�p���D�>+�,Z�"O�c5u�z9رcT�|�䍳�"O #gD�0y7�yZ�Aη9�̄	4��uI
4뇣Z$b�@�S�'���5��/=����0�ߙIi2��
�'�x��e��2�6I:��R�@�Uz
�'���)s��D��YǪ�A���'$H����q�Щ�v[�>+��!�'7z���Ȓ�1��x���-E���
�'d�M�W�۠}��mc�_��|5i�'�2`w-��k�ƈi7$�9��Y�'3v��2 �������Ԯ���'p����`��d}n�X�d�21$����'�����_�i��fnګZϚ!Q�'�xl�v���,كe�@�J��C�'�rՉE/§|{l$�B%U-G)D��'X�"���"�T�{r�aU����'FTX[���+�֤!!k�v�
I��'������7]��:�g�m���'�.]BBg�/���bgUm���2�'�N��W�_�P[j�����MÀ-�
��� ��+���8�0��	�!!p���R"O��z&i˞{�K��Cb�I�"OP�(��]7S�1#��xdv ˱"O �jV
_�3J�H�!D
�1vޤ�f"OZ�Z�� �\��uc��xh����"O:��5G��,i�ĸ�ca��NӐ�yRmB�ז�X%�ى�>�����1�y�l�w��$�GޢP��I�y2���e�x�A�O+�-E���y§�+��U��/*�\	�i���yr�Q�E����hF�p�`͙�A��yb��E0K�	�M���ڴ!Mu�ȓ*'|Q��A >�t�Q#�_6Q����ȓ?�����	N��I����1�@�ȓS���+��T]uty1F%:`�m��f�{���)`]�Y���. A�$�ȓrߨ����,����%\���������c��	4`,k�/ۈoW�T�ȓ~v`I"7��9:zvb�M\����B�b�a��>�������!�ȓi��1�!~��J���*�^9��-�f���޵Ik��Y�|�*�ȓ~Zh<�C�;����B��:J�ȓb�JA��G4T;pF�53���V�������|��R��5�ĉ��N�&���Λ|���#�+�0|lF���Oa�Ċ��ڦS|�I��	�zt��R���%��1'�\i�Z8!8�x�ȓR8��XvoGCurI�F��A�\�ȓ��)��[������Ɖ�zЇ�&�mY��S8qhKBށr�����)�T
�O�=$��`�&��ȓ"k�� 2��=rz<�% �H�ц�Gm��2u���K4�*R ̥8���F�����<d`\�pD�Q�	����uO�ف���9\JN��7�ڋ$~݄ȓh��lңKB�[oQ��CZCq�<�ȓw�.e��&��o�.�ң�;^=�ȓTŒ�2(��,^B��s�Ը�����Q�HQ#��+C��P�ď��P3v���O�.��ѷ'$�Z@��aklȄȓB�.A�3��8i~
� u�@%Q�E�ȓ_Ӝ(
��V֐PHE��:%�&݆ȓp/>Sl��!�z�)D��7�h��9z� ����#�n�����J�̘�ȓ��ѹ�(W7/��ٲ���]V����6h�`f�`U
p�eQ�xU�ȓT�L�H$��lP�UY�!V ���2�7HR�T)�kyE�J"Onm ���~�ܭR�咋.L�
�"O�s3�Ҵ.Y��#ɋkl�jq"O8��H�����(5�	�4��p��	:�:³�S�_k0�၊�.,J
eJQ���C�	�8ð��*\1.��أ�5s�H7M�6r]J��?��s�����d�H(NI�PG��X���"OH���ڮ (�1ç�`Ƞ�OtigM�=ʀ��=T�C��ɂZ[�#�
�1]Z����+�dA�D��"! ��K���}���Єj�4`��"Ol�*� �S�jd������[�����i+��Vy��U3^�RX�Mn��S�T���PяB��F)Z�lTP�<	`Dx�	y�m��](d������ D���7�ڒp݆���b�>1���wڎ��fl&�>w�򜻣�/�F0j#
�
����"� �2�HM�GQ&p`�o�+<3@����	;��z��G��Ys�'�2T��m� 8m��09�<:U�K�OT����GÆN(�"��̫�#�	�xR��C��x�'��;�� ،�$�V< n<�c�DHN����3"O8h���-&P�|���(4��$�$�҂ ����e�O�ޝr���K`4P�H�,'Q��O�P*�w
���HCr����+m��J��E-�s)��'b���kAv���K��/���R���
� �ܿ��D4��u@&�0*�u��FҚsS������~�?�FOg�e
-1.r<��l�=`H�[U��/s��qxЭ��<���(O�={���O[�zBh��4�!ި4��0F%�-b�1u�(���ٔ|��M`�p�OU��
�!�/Hh�9k��ބ�ڙ���pDXj�"O�88��D1,:�z��K�N0(��a�M`�@(�bS�v��X��#� lZ�g\p����dFȼ;D������M�m�y3bI�R��$$癎4HF�����J�����ǘ�t	<#$�� &�Uڴ)ڈ;�˓U�����)Ҥk'�O�soY#V,x����4]�� 4���d�T��U��>�(|)��PG��nC�df|�#c��@�B��V.�I�<��`"�A� ��y�GǞT�-����dbȊ���DY�Q���p��AU`��K|B����$����V|��#��!)̠(	L)AmĺBO>�h�� ��	 �/4�sE�W����	��~!�"��O0�5�\����� 푚wf`Mo�*r��RhӲ���	��{sʉ�U��fl6m���זQ���xD�=��em�&Mۮբ�J�y�G��/��t�m�.,��<qq�F:n����
\1(8#�[s�'/�� ���7��qa��Fe�Dx�'���4N�6����m�.Z��
�M� 	83h��_�(���@Z�P#d T�U���\�h�0�CH�!���T����HBY��']��吲.X7sK(���V*�����وJ�hy;U�z��I�Ɠ~AY1�l�X��
K�}����� ^q��$?��� �'�0yM E*Q՗�yR*�v�9�;e�=񔍓�t�$��P��`�:���I2a�0�F`dBL�5���#�����^�<(��4*�,|�4��$ކ&�д�rKCbB�	��y��9qx(=s��:�\�S"J˒�hO���2�O�� 0R����i>)#�ž)e`#�-\`8ٚ&��0�T̻1Q0X����'��M�C�(sB�
���8�:I��a:,��g��f���c���A�O v;' ^q�06-�E��*M�~�J�-���"F9D�ؒs�:5u\a1M�]��4���W/<޸sc�vޔ���M�m�|��ӱih��'�� �FOv�)�Ɔ"H�� ��ƌ�;���:�3�O���O��5ez@J �&�P��K-8vx��%.MA���4�|�'kj�HяHT8�>�qL�[&���͞�v����¯�Q�'G~� VM�2M뇃�(t3��;s4��}�V�pF�#� {@��T�'�d�)p���9'���,�;G/G	_�T,�&�K�D��I0r�x��umD�oX�$�'���-�'e׬h!����:7$ϦlmZ$���R�j"<T �e�R�<ٳ�B�v]���ư8��P��$>� �r�ܹY:j�3��q��dʓ��|�O���;}��I�� ��db��-����,��ɢ8���BF		'��@�*7�:���G�
��H��L%\����I2�hL��G'��(���b�6�>)��$�t��![�P�H#���0yT�H�4��!���V�JS"O��Ԥ]�y��1j���F���]���V;%
e��h��?��,W$Zuzm����1b�F�H�/D�|�G/
T�D��Lߐs�(X���Q�~����a��+��	)��B�ic>c�<+��B�0j�!���`�*9� �8;�*�yF �����L��}��f�|�'��OD\M��&#e~��	�p�z&��8^Z��DNr=̣?ɱK��vPe�;��w"ƿx1ըFF�:Y�i��M��	k�7$��:׌��X.�$�ǁ��__�$����<a��W�j]�3,�-��s�d�	$M�c?U�����Qʉp��S�+���rgJ)D�|�`��D/
-� i�ZƴåL�
,.,sT"�1�y���M8Z����m�M<ye	E�_��$ 	�
E �� ��T��@QID6bAC�d
�Vu��)�CT��8�c�sF��A%gKE1��h�'���p���n��h�r�ΐ�4ݰ����up�!�M�"<IxH��C�)h*T��)�-	��c�
8Ug2вGE��x��f�Z��ب�z���˄+��$�a�6��V-���$���o� 8���܏m��$��q	x���c�"�y��2Gi�t�E�[D��K��1k9"8[�f�Z3�m�AO?)��N~�a$/񤇾y��:�[D���7@� (�!���{����!!Y�Hq��;V��)`��ၨ�I;ҤCE�)<OL�DEP �.!#��T��$��',����R�z$p��8*U�0�Y��t�[���9�m���q�<1G��
Y��yc��wŌ�iqo�r�<	r �1bKH�	Ү��
�����l�<� B�����/fp\y�$=r2��X%"O��*�)k]*����C:���c�'�<� �)��I0E�Cn���*���.�~%�B�əV�u`�ǃ~	@=!G�+=��c�81V�֪?�ҍy��S�6
փY�rP@8��K,1C��$(��I�+C
�!ö��6�P�(�`�Ѐ��L�T�&!�&��FМ$��MUh<ٵ�0[��1w
�(�l�Q�	�/��P�vo��
�N�<yq5���e��e���[LG����	g��U�g!ZI@���:S�e��αy~�hY�A��>V�%�ȓJs>��`� �elʄ��+CK`~�&����kB�Ll`��DG{�O����L�/�`uu#ý O��J�'5H0�1(Y.��(hՍϯ.�>��0��Q�*O����#.�3}�.�"�2��Hɕ|*�t�Q�Ў��xbDρ+zX 3t,��!F��S$f?��Ǆ2F͒;B�'wR��3�F�{�����LV��څ��{��������Ѝ��'�b��4	 �i�| �F${�F9��'�Z*q�X,C�Lx��
L�Y9�y�O�N�M���a�O��p��&U!�q�!I�R���'�H�ԢYI�;`P�A������K/��O���Y�L���ܼ=�2ҵ-]�X����L=D��ᑥ��^UDIˑ
M�YޕpPg<D�;�$�m|]��MPs�m���;D����,!e�X�u.U2gDf��d�7D�``� X�����D�o�T���J!D��K�΂�p/�a��́[�� ?D��[5�_�|Q��ٖ�\�w��m=D�@زn�Y�4 Y��k��B��8D�`�$��'LBm[EH�;9^���ׯ;D��hS�W9\Qd�K��F�NVnP�7D�,�v	�r�m��K��}�|��"�7D� �"@�(>��R�AP�"<a��7D�4�sO��&~h���o��0�fI��3D��ڐ�G1(z�a1�KզK�B�1V$.D�Sn��>���ƍ��+����Vb.D����f�8��!k4��7`�a�� ,D�s@��)v>0���a�
=8z���g+D�d
�AW tvtp'�bNI���2D����dD*�`骆IF,y�L�`ì/D���r���5
cI��v>�T�+D�P�Q�	B��e�&�Ėy\VP��b=D��#R�����ǉ֑|\|X��/D�����.a�*��uN�dRdjN9D�|�wm��j�,l��H#C  Чn6D��H��J�=jB8��!�LS�aE�2D���э�>Y�ݰ��	� C�-�E�&D�@�F��K��1+օ7�]҅D+D�0�	�2a
$�6�^�Z-�ld�2D��3�eѺ(2������Z� ��N-D�ti�i	��%8@��XCZ�s".D���@L� *��@oڷGȐ���)D���+M.-(�9��J��Y����E%D��P�σ7}(a����W` �p�#D�qv��C���"�A�.zF�CeL;D�4��A)�"#!�]�h��D�4D��r�� |庴x�b[>
 ��)1D�d�f��I���I�4��``o.D�� R
�<XL��g��&� �&>D� �Y,O�-�� O]ֵ���>D����p��Egʧ{��4�pb<D��b��3`�}#��T� y&�!D�@{���!}��S�;'���8�:D�D�6��!
��ŢJ�x��3�'D��ZcD p�:�A���0�"`7K"D�� @��F�1eM�ZeO
�pg$DZ"O���*F�b�� � m� V�� $"Ot%9P�
=:@��_�@�h[�"O:���	�PXЦOi\8��"O��;g�_�;���VMH�*T�=[S"O����^g��@���35� �v"OL�a�E̚7�('W9.�� s"O8 p0���b�so��viPP�&"OX��T]���9���)�>���"Od�����y;F�0FP�3KZ���"Ovy�#�����@F��`#�0s"O�Q;����?{ l���]�n,`hYG"O���0H��&k�A"O(���J��2�KU���	1"O���x�6��C���,3�"Otv��%F��I�<��|�'"O��R@a��X�D	2'�b��C�"O�I# -8qU�d{�G�$����"O�����@�Jq�,���ƤVy�ͳ�"O���ԭ�Z�~��R��+�"O|��%�ڣ$*j8i��X$��9��"O�Q)C��=B�\��Qě�&yt 3�"O����	�4T���CcV�DP�4�"O�H֧�� k��%B�5�RU��"O�Y����/��3A��%�xp��"O���!H�����3���(���"OjQ�Ѥ�W`֐@�ǚ +��t��"Oa��L�T���ʰ>����"OZ����=D���{1&^1�Pt�d"OL�S6�38�D�Ae���Jkt=Ф"Oh�㤍�ffڱ;��	�^�*�"OR�P#͌�R�IT*K� ;��k�"O\�Ð���S ��)q�Ös<�tb�"O:� $� *#�Z��#r�Śc"O.%�eG,v*��a�z�.���"O�ѕ%��DҜ1� ��t��"O�q��*�&rFvT���7MJ�)'"O����
��RS����DH#���1"O�����E�H���Qʪ�m##"Op����H.93�D�@���s"Oj�O	�W��Qa�Eh��h�S"O`uP4bX	+���)��\4��"OF�I.����M�2�Ё�L�"O(Q"�g��Q���τa��"O�̐ҩ��5/,h�!K�^�.� "O,�j�	�;?��a�!��$ݴ4qu"O�pR􊆶:?ݻ����l�z"O��+�=@�F	�C�� ��-"O�m�U�P�3L�y� �4P��C��8����R�@���j����B�	�^��u`�̏lM�L�#!_6+�rC䉮z����1��5�ڈF+�B䉜9>���ԇ�7v��t+�_�\��B䉵3F�$���F�~�P<��Y���C�I�HFȉ�Z�f�헿J��C�	�$3���s�mn��Y��ɺ�P�=IajIq��"}��#�B�vU���'������<!�����^	���I�m��������Bp�����9%�"~n�)l��C�ԅkD�4*Ƅ�f5�C�	�o�T����+c�Dr�.+O�~�I<fR� ���2w�az�߫*�xR��	�0ҒY�eNߵ�p>Y&-�;x��ڷ�
:�D[*�����L�x��F"O%�rO�EZ�Y���S��I��%Ѳ.���Yp�Yy%��@Ŧ�3��Q�S׼c��ނ9><���C�/��3whL�<� @x[�L\3t6b`q��ƭ(e"��r�g����'�fԂ�O�)KfY�5�,Y�y"�tEf�΂J���#���p<��K�9	 !�b��iP�"]>4n�-�a�õb6��RB0KV�ɍ	�%ӱo�`azb��+�hTC稖�j�9
3�W.����-wЮRtf��Yr<���囌h��)�<ţʻA�@���ĭF�h��G�� ��B�� qS`����� ZNR1�a��<�$p��w�<=�f-Q���$4@��S��[����'�~B߼۳hK�f�4�#L��;�#bP�"�O�)҈� S0�l���0ԫ	�%cХ�х�zǚh� ���ŏ,��d#%���s�#?[���A� BB<�?��/N���D�s�BS�9����!k�lU`��Y��݈�R��bL�/Od�Vc�,KP�z��b�-��Z;gTʈ�a�-��D�"h�mI���
���RUĂn�D�'$6��ǋT�,n8�@��9J�$a���30��'(Fqۑh@,��y�X�v��J��6���bH�v9�
w( /6-J7�QZ�]{}��m�!��K�}8��1�آ��l��*�O�0�5t�j���T�JeN�:�H�w�x�pV��d�ԯ��ɿ�~�	�Q��'���	�H�u���3f]�4�lM����O�qtO�t+ֈ��J��u�f�0��Ձ'�`��t�2�/���N�Z��0ӅG����<�@��I�wI�{�`��R�J����R�
Q%���?�2!��C�5��HM9ȉ?��٢V(��z��'���.�uA��e�ˡT�x�a�{�P�d;���e��v�ָ�'�V5��m>��D�&>�&mx��t��PF/)D���񏕀0n�;�m̧d � �D��V��׿F��tΓr�@�|�'��h��?G�^�
�I¹U�Ԕ��'���H�kIЉ����U#F�p/��O� p�6D�Z3��x�'�4ظ �0bP�%o�]���q�d�;���>4w�� c2-I�l�mLF�;�JW�nr�)�Ɠ��HC�Cvh��$�)���=�KxY��O�ZC�ߺ/��و�L*'���q�n�<�JQ;�>hh�-V/i��EJ��D.����BT�f���'#|�|�'������}��*��MTɰ�'H2��Ҧ�&x>�h���9.�i �d�.e�BgRu��E��I�dό��D�7̲�Ҥ�� ����3n�:A
��ªAp�7m͠C��Mz��@%�����,l�!��+T�h��CP;��s��]7u�O^)[�L�M�D7�,�'Y����f�T� H<�����,ꞈ�ȓ��pH�ț6���zR��,]��H�+��e���IL��~B�.#�Hy K�5!�,p��S��y���?*��遤��'Kx�����?��OOPR��7lO�x`�HI�V�~��&��.� �p��'܄eYT���l�d�[+*�B#��ZGLA��FC�y�)��ɒqӄ��xnu�c�W��(Ox�۳i.����L��i�St�!bN�"X q��"O��!�V�GM�T(��9::��!"O�l�Go��	^x���ӥ3����"O����5�����L�j�����"O�mP1e�td���Q�:(�"O���̝|5��!�˃�!�Q�G"Od}C'k�u�m�c��D�NL�bV7u���
p�Y�9�he[�D�,Dq��'�B�cN�E��d�`CY�#8�!S	�'�F���(0������{!
u2Q��]�*�+��_j@�GP&��yR���,Ɇ�RdY�w_�= eI +��O�,3R�f�aI����B�����$��Å˭%-�#�ş�qH��c	�'A��#-�'
$,S##�!L�p�+O�8�0�f��B�N�.M�`[����O8T����6dH��
Y�����'��ReBZ$a[6�BJS�0�[ԩ��V#�mrv�«&�>�������'%�:O��Si�=���� �D�]ъ��%�'Ж��ɍ��������R�[3L��%�ȹ!݂md]��Δ�0Ď���w�iiU�VwJāh�`�$�&�?��Eկ\Q�q�"�Va�����CiVԼ���N�uf���eQ$u~8�5-$�dyv�W��\�۸Fh�ѡa�<�2�Dj�����W�^]�=�u�ļ)�Fb?��㬚 y��A �F�'3�Z(4D����&G�{��0�Ԋc;�����S�}nx���i	�`fD���(I0��N�N<�C�r}���7�Ǧ��B c<��+�	�|@+J�9M?��9�o��DM��NG5`�����ÎQ�~4�	�S�? ʈ��`-xV��@��D��6\ �'��Q��B�?���`AР3 �4f�� ic�#��]B��
��Pv�<��%� �0���k+.��c/�p�<���I��z��H,��jd�r�<)��<� L!�_$����r�Pm�<Q@�=N�f�1����q:��x�`���s�#�$"���'��9*W�һy�V�ҁ�ȹ��'R�T�&%�'z����1��8��a�y"���	��Ib�e�O�$��e�]�(�T�s6�\�Xn �
�'����&�E���5)E<T�M�'���|gH�Q,ORyT�?�3}R�Q�6hyK�圹f�TUJ��˛��x���-\�uУd7�����I�9`����bE�8@F�Q3�'�*4����t�rÐ58��Kϓ	�z��C�6>��[�'蚨�h_�$'��� �#$��li�'�f�9 D &8��ȗ�^�q�!�L>��cޱ~��t��������葢�J��`�!M\;�\�2"Oޘ�h��2hպ�L�+B�[�b��n��e�V�� �.\I�g�UFP(����x����"��y�񄈛K�����7�N�[�%K�1̨��/Ѩ}��I�4�OФCӪٸ�4�U��2A�|�r�'� �%C�41F�h�b<O�A��CG�
V��5PPm1�"O��#!؂`�����͋��ppc�$M���dX3�M.���:u	"��~V@�I�m ����&"O��3���>e�V�!>��2�Y=B��d$� ��<y�hY�? U@d��.uµ���w�<!�B�F9��L�/0��اcF�<�GQ�4���FJҭ/��1�ĦKh�<Q�O	N6��A�$ !:���ef�<��䝄N��ÀP�Q��^]�<)beE"ȴm��ҿUH�t�g
�s�<s�L*? ����߮?��q�u��j�<Y�"�u�\�[�ʨ����KI�<�@[�]�Q�E�/�  �m�@�<�ǔ8PXp�/��-@�gl_U�<!t�V<�x8�ᄸ69��k�F�S�<٠J�<!t^�[�/,H`b3+�M�<��!ŏi��ò��	b��Y�g�J�<��!�4)�]{e�Yw�M�E��M�<ٴ�%}����lB��ʆ��M�<�&mۮ@�Ǧ�%;����mVf�<��i/"̩�eu��Y6
\�<Y��V-\E��FM�&Q9��G�<%'�2м9YWG�		�Ա4�Fi�<A�a�S���&�;ʺ�yF
�e�<I��O #ˀ���Æ�Y��i4�i�<�Gʊ"g@| � cN�	Dy�BAe�<�v-Ѧ#��Cgg@��=�fF�e�<��T�{�,�qr욯/���V��b�<�H� ���j@/G��I�U/Oa�<1�I�R�<Uѣ��'N��)�M�]�<� �=;��C�E!Ri�!%�X�<�eꇵK���HD�I�VO�aj7��_�<�g�C(3��iL=]����E,D��qD�D�M-�
�)�U4Ph0� D��1�V"D�@#��T�a�����I�$6~:Gͷe�Pia&(<LO��k�
th0�'�o��"O�)��� P�S�U�h�r�"OhU�w �3��x���P���A"O����s�� )�(8� ,y�"O�! ���6{�\j�Hڌ<��ib�"Obؘ � w�12$�����j�"O�qqe��+9.�dD���
��Ղ"O��!� ��'��H�&�];�p��?Or�'�t���ܞ"�Ή 5���u�ЍR�A���9�$ _�.;�l�*��'A~�� ̐r��S�g�? ,X��ƨOߔ�B%��;�YB��E?�V�Qo��w�R�0|jDK�b�)r�"�#I�����Ʀm�BL�E/X y4	 }��)�'����:|{�)Ӆ��	I{ta6\�W[^�˧gܲ]I(���gW榅#��O|�Q�NM&-���C�ވXx�#�ǘ�5��`��B�ئ�@y��Ocq�f��"�>���s��ʉt|��7H�9 �u�'&x��
�`>����L2d���ࠋ�u����e��j~���c�&-+�$��I��"��L�d�uU�A`����D�	���r�,�)ʧj��[D ϐ8��x�j�]BlL�	=E��}���^�4$	�&ȎI��I���@&9&��`l#�@B�b�'p�����<�J�o=D�D�Q";n��
��W��$���g8D�hȧi�#dŬy�U���E�<�S!9D�4���7k�J@�ň�^&$�{2c4D��S��M&�r(`�A�`�Y��=D��@�Ӧj��TC�G1kd����:D�`�h[892��E�mV
��1A7D�L�sN
���sJ����%�ǡ'D�����W[���H �U��I3��$D���g�ӗЭy�&��"�����7D��Cqǘ5d(\�E��(&�)�t�9D��"�i�)3��Ɋ��W�'�N�(U%4D�\*�DB$PQ1�
j$J�	a�2D�|�w�J4n�ГDR9��`��1D�la6k&�x=�3cR%6�+�C1D�8�gO�z+8���J9"ވ�c�3D�l��n�L���#��;g�`2i$D�x9e�ض�.3��G,wôԘ�,$D�����Ơ6���WM�$ex��#�!D�ܫ�.��N��|�B!�"(�a%D���i�2h7,� �W�xV�@e�#D����	��g�e
��#};�pq �!D���lA!_m�|����"D��� #D�Ty��9� ���"�&%4����"D�l����zڑ�5�C2a�4�E� D��'IЧ1O�p����)�h��f,$D��[�Պ*�0���Ț?A��R��"D������i��hֆ�)i@4��� D��;��K6n9��@�BHyl���:D����F_���M�o[�~�<���9D�<+�F�",��� bX0����Ħ9D�t���H:&]�,J��&o@�)�Ј"D����+'S)�Ed��;��� Q�$D�hqǋ����D$�/~Nt���k6D������Y@���i�3R�4A���4D����c�ZfV0�$g��H
p�4D��k��Bp]��)����&���k1D�h�:�4h_6Ch;��2D�H D��s���z�Ǜ�H�Q��$D���CcN7J�Y#��,�z�H4�$D��pr�9k�p(і�5΢�B5D�$�dFP�\�$��� )@b�p�E'D�����+N�DN�"N�xP6�"D���@-�k���hD�I���Sa%T�xR�&Zsv�Q�ˉV5���4"O�����0OT-��C��֔cT"OB�s�mLhY�����O4Hy��"O,}��I^Bf�X"�ڬ1S�!�v"O���7�Z����T鄑=<J�@w"Oh������ 8�k$�'	/��z"O`%�WELz���
��ƴHK�"O�-��K�1�<4�0)Yx�jp�B"O�� 
�54�p���E7Ux 	7"O>i����r��}���N+����"O�i�#��,~�y�"جC�"O� 0uH�n�-Y��8e.�#�(ݹ�"O<�b�W�S�.�[��އzjz���"O�-����<$��\[�9��"Opx3���H0,ps�oP�M�B�V"O�}{Rĝ� �j�9ro �5��x�"OH�S � %�&�9�CS�g͚���"O�]TᖥL;}��Q�Q��)��"O
�h�G�5 ��+�׶�(� �"Odm	�Xw�����Y#�v�kG"O��+ޞF�`���언y�X�y!"O�ŊtFʝK�	a�k@N��y��"O@��(d!�@��
t~:Ar"O���pdX�{H���ϗt�}��"O�j����Ih�Ң��8��Ã"O��@�Id���S>]ީ�Q"Ox\{EǯL@�W^�fRx�r"O�t�ӥVm����T�5zA|��"O�Lx��.X��%�5@�I5"Or�u�176`�XÀ�YH�÷"O$����O�P��N�&X�R�"O��㍘-,��Z�ٴ&��$"OLp0�
MR����q���"O�y���B8dq���6
�Vi�"O�z7���K4v(  ���n�z�"O�����RR�ƀ#Q�G22� q�3"OVMFHD��s�T)Y�����"O�=�`�,}ܨp�������"O��+w�2
X������$h�"OlI
1G�P�*�� .Q��/D!��ۿ�"<���8Cf6XЌ�8k�!��1pR�L�D*�(J�Hv��G!��<W��2l28�����q,!�č�NW��C`C9�\1�M�3!�Q�D��6���]��[�"X&(�!�ć;u-�E���iI�mq���t�!�O�xx��E��c<Ό����/iq!����\����>_*v�[&gɇbW!�dW- �|x1s�G�@b�"�N!��ڑ~�`F�Z�X{ejC�3!�ڹR��,z҃�gL��(c!��5M��@���h���#N!�,vL\���n 蠡c�[(!�%e�I3�o��8�1�*��!򤍸jt����W��EA�o�K�!�$Z�tP�g��3�p��wlM�6w!�$��m�\��� Ŗ����!�$�"Bd�\q��G0b�4����&$R!�D+dI>�3wK˰|�L��JH!�$ή)����� ��������ȩd*!�D�̈́���
)5�>��j�. !���o֮]�W�H}q����ִD�!���=?�&�#m]��ڨ1�(R�|!�ݴ2Dp��eU/O��9��'�%{!�c�����dޛT��ʧeJ�h�!�8*t�)��)چ$D24��Y�B�!��$~"��Y��U$)�:�He��]�!��^.-h����/^�=�����N�E�!�S2�܂��)yP��X��d�!�d֨c����`JC9O�0�`,!@!�D�.��! P�F�)�(�#&��!�D�?J6��A��d��X1�V�r�!��.LJ>���Aj�q�����!�D�r��(��Z�uȸ$�"lY�7$!�$O�(G%��`�&�0�<!�� `��*q>B,��a�&"X�q"O9��@{��#y|�S"ON��p��)R��A�J;]�)#�"O�<����S�����֑p,�G"OPX��fDK>TTխ(Н�A"O���ȫf@��I�X�Z��M�7"O�mSP�h�d$��`���8�"Ol�1cl!?
�C�J:8u佲�"O���c�x� Y�hK�� y"O�zB�%ȦMS�HS#ch�xz�"OV0�cJQ	���bUHƂee"O��z7HI�)�zЫ�Â	3K�E�"OV4�� hq�'�Ł?D�A "O��l��:����%M\	~�:�y�"Oj���N
IA(�ZuF��Q�tԨ�"O�,�4@!(l���A/�ΐ��"O�x�朑4��@�Dؿ;��S"O���P��/c��a�#��K�L��"O� v�ٝ߼w��o2l#�"O|`	b�ߩV'%;�F�~���"O̴�v	KT�6�g�=n4@�S"O�EH����Ps��ב�d��e"O&�B�cF �r��͘w���K�"O�x
f ��oX��юV�}	�ݠ#"O� q$�t�x��-A&x�$�
"O���"�ӯ^<�� ,ˆo��\y"O}qtd܍?0���sKؚz�v��U"O,	cOS+&��غa��2V�03�"Op�A1E}i8Qr��oQ`�ҵ"O�d�u�$q$���gX6 ���k"O���bn�XVx�0�N|�P��"Ox���%=����ŗ�L~lu�A"Od��a,�����䞮p��Pp�"O��9@��]h]�Ff5�j���"O6��q �C���2��
��T�"O>e�T�L)�<�1��I���$"O����"��=��!�pዊ��=*�"O�E �Y��PCOK�xv�c3"O­�B��. n�yq��b`��"O*Q9wB��!C��p��OGO��zE"OP���HR�s̲��"ь+�R��U"O� ��
lؔ1��k�r9��"O�ts누2&��SB̨l%Hu��"O�L�Pq�d�B��fÖ�37"O�]�$�ŚU���I-�@��h@"O ԪgĞ,H��3�FM�Z�"�z�"Oʼ������bF����#"Ol��2o�y4������?n�0��""O����z@�٦��e�����"O���Q�
S
,���\��}�A"Of�k�H
6�a8�!A�$�@"O�X����e|T�a� [����"OV�����+Z��)"�hS�NM(S�"O.�'[.R2n-Bǈ2jE�d"ONXj��I X���� ��4\�dq�"O�{@�̙~>���ĉ%q]�C�"O�LC���>ys��x�-\t��t"O� �:*F:e��Ֆ<r���"O�ț�$���ԉ�D�H=a7"O~D�C���v}�mC�HD�b�
�
d"O�� V%cBt����*�V"O��f�&u�����b���0�"O�!��8���
9����"O�K�̆fp�#��T9c����"O� 
�H�gɢ)�ȣG�v�̘S"O��ઋY�<�x�	���a�T"O���b Ϣ��q@Cfr�(��G"O|�����j2ѐ���!s���w"O,��F �T�����:l��r"O��{��J�QtD�Vc��D8Z-X�"O
9�S�3C`��3��U��ԣC"O��`�� �yY��WLiU"Ox+m��Dzڍ��/'4��"Oʼ5�*�*,!7��*d
��@"O`���d�x�(��D�&Èx�"O4��r�3��҅F��~�l�`7"O�4ɆE�n@h�'%��R}X&"O�9���:�^,��X��	 "O�3��2}�xQ�����"Oh�ѦHم;d� 	�eg$���"O>���}E�8 1FTRB"ODq:�__�X��1�0hi<�17"O�y���p���Q'r\b5��"O.�Ӆ�*5����&�:���)�"O�I��   ��   �  �  �    �*  �5  A  ML  dW  �b  Fn  �y  ,�  G�  ��  Z�  ϧ  �  w�  ��  ��  >�  ��  S�  ��   �  P�  ��  1�  ��  �  ( i $  k! + �4 �; �C M �T �[ �a h �i  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C�d �S�)U=w*����R�|cC��<H!�D�0@3�qJbʌ�h��K��I+ 7!�$O}_�%��h��F�h��d�S�0!�d��K�X�a�R9����Z��	A��H�d�ɀ�XfΪ܉�T�θ��"O8 ��)}�!pk\�'6.q�f�|R�,|O�Xѷ�������fE/��0��x2���&?-yN~J�ݩzGd�bp� E ��Q�
U\�<�������Q�ae�&
�� ��_ߦ��Ol �C������禡��b�3\����퐀h�މa�".D�$#!EL��8�0�R(n����>!�S�ԛ���3K�tI:�-�n;�q��>L��H��S{�@q�̴zn@`��JQ3m�v��ȓ	f
H�@��?%��q��V-L�V�ȓ��ґ�=�ޝv(^)���ȓ=\���wnX5o������&:��D��h�JQ���C:n�cn [���ȓ-�<s$��x����b$�F��O�7�*|Of����46`u#��
�����' �ɴXBDx���<WW�={V���KنB䉻���%13q��B���h�>i��	ڪ'�n��)\դ�B�d�/!���R��:1*  �#T�8��K��h����)Z n��1��ăQRD��"O�p@�� �K]�-)������<k�"O� �m� }�X܋�-�)c�T7"O^�!vB΋�����>#���Q"O� ��=tiztk��-g���"O�0��eLx��p(�G�~S&ȫ�"O���Am�N�d�R� i�`�"O$@�Jǀ\0Y�`�� =Y�� �"Op��#	8��Xc�e�䰸"O��x$��3��|�уSP�L��"OJe�����I|�0�4�3>��-;$"O�`�F)t�b5+'b�?��DjF"O8���������c�#C��`��"O�qB)�3"�f�9R����8a�"O�X�)7��0�g ��q�< :"O�YZ�׋i��zɎ5Yq��§"O�-�� �y"nta��be��5"O
]�ŉ�#x�R!Fa:�{�"O� �饊\2^�����J�cH��4"O��p@HH�s,�E�1B�!i�"O�ݫ2�� l�pi�!��~*DM�"O��;�U%�l�+n�1�6��"O��%�S�6����LN�o��{�"O���'�09k�8Xp�nF���"O�4�Ty�T�� 6x5Х�C"O��S��D���]� 3d��"On�H%�F�L�j�z�.߈w"��J`"O�Y�gJ"���E�U��Q��"Od���G�1�f�3��]%� ��$"O ,� )��zGLy�ѩW x���w"O�E�É�I���p���x�yv"O\���a\�Zn��!�.�-9�"Ohc�@�VLR��5h.2�9�*O
���<�8��t�[&��\�	�'�2� �S�0ȓ��˄r�L�
�' x�J�|�xԦ3~	��'Wl�9��I��h�����i�V�z�'�D/�3<���GT9*��hQ�'��p�ƍ'�^x�����(�t�q�'��� ��*7F��AI֮'(���'x����`Y�K�p��
P����'*t,x�.G�V�RljsC����Y	�'�f(A�0��8p��S<tdz��	�'%Tl;a��>$s��Gj�8s�����'�x3d$�*%~�	Rŏ�5�j}�
�'r�1���ty2-����)����	�'9|ɥ��GnZ5�`JA=	|�	�'馴xwl��)t&��W �7$��2�'��@��I��Y3~h��h�	�R��
�'�̘�4�E@�����/��1�	�'�P��ӬZ*%���E��#wLY{�'��bkZ�}�|D�#�@!@A!�'��84	�̸���%������'�T ��*�d�0/X/��2
�':������Z���y�/ҍG <�	�'7B�f�;A���h�m��D��	�'�N���N݋Ei����h,C �U�'Ɇd�VӼ5yX�B�D�H|��'�Y���?�<@�I�;�ZA�	�'��l���Δ�z�Mۤ�R��	�'Mޅ��F� N�(�R���[pE��'ڽa7CG3���ϓeF:�	�'��(�`	 d�T �C%5҂�K�'���G�7N��3C��&x�X���'9x�b��9[����S/?u��� �'�j��� X:V�Hè-t�0 ��'�,��"	�Q�X�����!����'���H'B��a� ���0��'���0��� GJ����I4e���'�@X��_-U�h�"��5AX����'܈���@��.���\!@j*}��',��#&�? ���"d�41��R�'"���u �)N:�˔(���B
�'?�H�$;�Xad�����	�'���1�!�5Sδݐ�Ɯ��Bh)�'�e§��5��8BtmI�����'�hp�O��C�vȁ������
�'xT�DR:p�����x�!�
�')5����J�k���p�^��
�'nP�#5f��%�� �"ɘ`��	�'z�|7�ϛ@/�(�A�9W�8�H
�'A���H�0h�p�`�#R>�,;��� N�)uj�+�ļ�㍙��*�0F"O�YY�GKh��Hq�_�1�r�9�"OdE��Swb�Tհwf�8�"O���j@�fj"��:g#�"O���KG�N表��49P@��%�'?"�']R�'���'I�'Z��'1h5x3��Z^��B�	bW��r�'�r�'�"�'���'L"�']��'s�)M���Q����6Ċ����'���'���'Y�'���'fB�'�xxK�� {��pO��
D���'�R�'�B�'��'���'^2�'��$�!������am��"�'�R�'���'���'nr�'g��'r��+Êd�([��Z�&��xS�'�B�'>�'���'"�'���'{@-�%�J\���l^E����'�r�'��'���'|��'O��'S����K�!����"�W�q��3V�'J��'�B�'R�'�B�'�b�'F�e��AK�g�zD�0NG�`�`��0�'�"�'���'("�'�2�'+��'<h����Ky�-�c�&<�Q�'��'�B�'$��'[��'���'��$c�V�L�3��"u��Z��'��' r�'���'���'"�'4�8�m���e��Y�L8��KP�'�2�'*��'R�'�r�'2��'����# �#c1dypd�)O�d���'}��'�Z.���'x��'i:6��O�����%�ΑW�Bha���@��S�%�<�����P۴&0P��F� '>
d7H˂�fm��&���M����y��'�aJ ���sN9ys�	x�.���'�����E4?I�O����+���?��@H�1,6E�&�K�'-2^��F�i��gǒ�"��V�/n�)�t.�5 �^7�L�~�1O"�?�@������͎0y�!3`�`fh�����?	���yBV�b>�$��̦U�h| �"a���hH^ql�y��y���O����4���d?Z+��r� ���F�tT�$�<�O>�Ծi�ę�y¯��s���K�kX�|)	�+�#��O��'���'<�D�>pm�>bx���t��8�%��"@~r�'������O���I)⎏�/�f�:��=n�X�G�*��by�����	�a�TA(��Q
�|��KO�qN��Ϧ�(:?!��i��O�	Q�Yz���E)�*�����
ߧx���O�$�Od�	x�P���	��d���(J����آ联Ee,Ez�C�����4�V�d�OR���O|���{>���#�^��9U%�>&��j<��,;*zR�'O��t�'6�T�w�6&���s��9}*�{���>yg�i��6�.��G�s�-����i� ɑP�!7A<d���XI}���e�r ��f���]��� ��"oz�q�b⛛Wt5/P8a�. ���Iȟ������S^yb*p�^A( �O�!CE	�3�U��ka6�K����̦}�?�6R�`�I��`�I+3�l���Ņ�4�J<�B`C�˓�c��7�/?	c�RQg��I*�D�pݥ�ݹj�x\Cb۰s��irq`�OJ������	��,�I���Ic�'U|�T!a�1A�H ˓,)J"5K��?q��囦��7f���M�I>G�!k"r�;�'M._$��	�N���%�d��ɘ��6m=?G���2�U�lѡA��)���>l��I0��O,O��o�Ay�O��'/ҩ��On\dᶎT;"�Wd]%�r�'��I��M�4��'�?1��?y*�����
�7t�XC���渂E����Of�nڬ�M�N>�Ow8��Rf�$Y������&�$�a�Å+��qQA=��dNǺC���O��.O�n�#���@�a`�N�L�&�D�O���Ox��ɥ<�3�iȈg��i���1���g���� K]p5��8�M#��>��O�,���k����O/*4�}���?�u�^�M{�OyZ&����K?U���ǋ
\m����N���EW4�M[)O��d�O:�$�O.���O��'/�Xi�)�HO��P后6I�����iMn�r1�'��'X��y
k��nW�D���`"�[<&S�I�+.�ao��M�L>�|��N/�M�'݌ a�
�BI
�pa���{���9�'��0+$�Pɟл�[�ܪ�4��4����O41?PA�@�*7r�8$ F�O�`�D�O���O��g<��� �9&��'<�"��E5��v��e�Z4�&ʚ "�O��'�r�'��'Rr%�d�'JR�ܪ�ʓl�@��O�8T��; �r��U��XyZw���	�BS�/$����=)�9;�iҴ7(��'Fr�'�����P�PB������O�2jje#u�֟0
�4Q�j@.O0)lZc�Ӽ����4#2��ra*�9F��W[����O����O���תa��B��MSA���M��+]0?�NՉ��N�mv���FS���Ҧ}���d�'�r�'7��'̴��O�=#)�ͪkX VhHH�1U����4,m��Z���?�����<i�Ұ)	B��12�.���X� A������	M�)��i��qy��˫W��]�Q"�$�"m���D�'2�!I�E�$��Op<p-O� mey2�CT� �1Pk��~����Sa��h��'���'�O��	��M����?I��Y;9~�a�Ϝ-�2�6��?��iH�OX��'� 7-Cݦ��O�l�@������$X~�p�`�����<�R ���='�����L�Ov�}�=� �xAQ�ɜ~�F�(�n�q�4!#�8O��$�O���O����O`�?��F߬]C���E� �f]A��ɟ�����,aشS�V�'�?1�iO�'�$�K�̆^a��4H*Pen��ę|2�'��O/�b'�i���%	�ҍ
Ag�,!�9�v�մc�
�����,p��<!Ǳi������	��4��F�Fq���Y��R� ���+�t�����0�'l�6͔������Of�d�|*��L3s���s�S$7[���#�@R~�˪>����?iO>�OY���'��H���r8���ޞ;�(���i��*��N@�~X���&x���AQ*o�}
�!�$QR��	ğL�	쟴�)�iyr�{ӪL@�N�\R�y�m�J9����e�~�d�OflmZ_��J�Iݟ�1�b w�*A!��؁`MN�kb����\�ɋ�XImZ]~b�]�JDJ�������]��)�A��f��Q��	C�Z-mzy"�'s��'���'��U>qH���uDh*N@
`*������M��M҈�?���?����h���͔/k�����/	ﶼ(p�Y�M+\���Oz�O1�N�hs���I�yQ�!����1��a\�o���	�b�}IP�OPʓ0ě�U�������s�E6�hȊ���*�p0c�N��\�	���Cy�h�HS���O�$�O���֣٫�M��e�OҲ@��]�n���dl�L�	$�&�z2lK?��A7���"��0�#ȋ8�M�T� �Xwdi���?!�Fڻd�Z�9҇Q�3����!���?���?����?���)�O.9�%΋�dU��ati��"2^���o�O6�l�#,9�I�l��4���yn��g�9��ԔJ��Jqo� �yr�'�2�'�(���iq���F�R��gП�`�pƛ�8K��x�H�$@s�HhBh�<�"�i�Ο��	џ���ܟ�	��J��r�L<��@� GM�J���'�P6�	xk��?�O~����:8�����!��Q0g?8�w\� �IΦ�<%?I�ɂۢUa�BL�6��<H�ٱ��lڠ��d �hϬYh�'T剃�M�.O� rElE�A~�l�2
ЪN�l<����O���Or��O�I�<�w�iH|�J�'��T"�M�/'#Tk�O�\h���'f7!��4��D�O^6��O��3����:��� h�3�8m����r�n7�4?�%�.����hyIk�)���P��SBD+t�@�į�"Hq��I�����x�	��P��z�'D9<h4����ܹd��CWJ�R��?��o�v�:_���6�M�N>D ��W�l�!^gB�!��,@�'<�6��Ŧ�ӵJ���m��<�B�,C��R��S>�=�	��S�R��僘�&�f�#�����	�<N�Iڟ�����h�	���G��(J����OV$���䟐�')��D+'��I����O�؀o�3<V�Ѱw��X�x���O4Y�'kR�'�pO���7z�����SX�BX��R7��P{���d�h>?�����E��Ӽ[���F�̼�fI�g����@��?Q��?���?�|�.ONLl�(���Ύ]���h�h�+��#s��iy��g�Z㟐h)O�6͟/�d ��L�4!v)ZU%â:C��n��MS�	�M;�Od,C��T�
M?%��k�3&�\��c/N$.��tC5��'�Mk.O �$�O��$�Oj���O4˧'����R�-7(9�7�+�0���i��e��'���'���y�Iz��N�@�(���z}R��"�/ĔoZ(�M#s�x���)Ȩ/�V5O q���mB�)��7#�?OtZ���?A1��<���i��i>Q�I�p;���ч^���[�@t��q��۟h�I��t�'#�6M1Rl����O �D�	r����� eRp\�ΝR��㟈x�O��l��M�A�x�.�3#��\�uB=�3dH�����R:z���+�",d�I��u�j^��H!��'8������9�8=24A6@R����'Z�'V�'}�>���	L�����HP�E��&��j��I�M�����D�����?�;d�@{�e��xhR�	��õ4[͓�?���AX����8��&�����Z-��� �̼YB�Ve�&E�uŒW�H�'�7M�<ͧ�?1��?q���?�%�ĤdPa�b)�K*ްǨ�>����=�"�U����I�P%?�	�l�Tp�C)�T���ϕ�0C�O��D�O��$�b>y�+B�l�i��I0 v�Ԫ%g�'��0�f�;?	EK�0DN�������V�-�'�
i�e�51���J�/M'�,HW�'�B�'�2���$]��*ڴ}����W�i��'�]���ҨBD�}�.n����_}ҁqӐ�oZ��M�SM̐+�Jk2�S�Ҥ���"�5[ȥ�ٴ���S�Lr�P;����S"�u��w�2,zG�,Y����: 	y�'p��'_��'�r�'�]2��yV(��݅w�@��n�Oz���OJ�l�8�E�'g$64��M�?��%Z�H�R	�0���ʞd��($�$k�4jz��OfT���i[���/ށ�E�E���!��^5]hεJ��_�_Q�oZby�e���S��O�]ȗ�T�J�HLz6@�2<)V�*v�ɹ�Mk	����OD�'
-ᤏ�!`��`�А��X�'x듫?Q���S���5D6m�c)�#L:�rI9?��0B�h]�X�R6T�擧t��H�B�ɐfN����b�y��p!"���c�C�Ƀ�M�GA�9�\����ܫu��X4FˬA��+Ȏm�`�u����8��ۢ[|�H�p���B�{娙ß$�	<L�m�\~Zw&�� �O�B���� x|jO8�`�"�z\�C9O�ʓ�?��?���?������T�%葠�MBd?���!	���UlQ��Y�'�B��T�',�6=�%2wGQ9=U(��Eh�+#���T��O���"��I�23�.6�p�p���p�2L�3�L�~0��x�@
�+��:�b��ay��'ҏ¨Jy���%��-[�e��Ё-��'L"�',�	�M�7#���?A��?q@I�9E�[Q�E�(�v�c-	9��'��듉?Y����E�hu�K�E� z��X�Q ^|�'�\@�D�Ně�l8�I�8�~��'��� ��-c�Ȅ����N8X��'1B�'�2�'�>�]�^ꄺ!Ȃ4.�ڱ�e�9.`5�I��M�Ն��?���f>���4�"�@("���V����e18O����O^�Ė���67?q�&�'~X���_�Ѕ�HT!��.O�\�$�4�'��'Jr�'��'�n�"�@|��e�6"�� c]�T��4?�����?!�����?q`�L�0�pE� 	�v��h"���a'��ԟ���Q�)�%E��d�0��"obR���l�r�*W�̦].O�`3�k��~��|�[�@q��_��>q&��4�,��%\ҟ���֟,�	��\yraӀ�� N�OdDr���'8�����[!r@�HX�?O�<n\�L��Iǟd��͟�cǡO�D}p)��J�/�䉴�7P�|l�z~�'�&l��e��]�'���t�LMS��e"�]��@bƌ�<���?��?9������q���7�N�/,I�V�O<��O����ۦ�[%� Gy�vӴ�ON�B�"��0,��Ta@� q�n4�d�O��4���Y��gӎ�R���aAϴEΰЙ�	�у2��4��D
�䓕�4�l���On�����̣������BN��nD�D�O,�_қ&BЦ{Gr�'�2_>�aI Bf��l�x���fd(?Y'[�<�	؟&��'��#B���8�4A���./A����1? ���4*�i>�Q@�OƒOfx�b&I��!�F/� ��U���O����O>���O1�˓?��voQ�N��u!�K�m�@��S-�5Wt����'��!vӺ�\�On��S�<��hJP��(!g�U�g��~��d�On�U�w�T�=��T�7ʨ?͔'�V��1�<U�B�\F���@�'F�I͟��I��p�	П��Im�d��z�f���O�qXC������6W Qv����O(��?���O�Tlzޡ1����HhJ��[�#�<�s�e��Ia�)�Ӱ1�*TnZ�<�*P�[��\y���;z��M���F�<���ƕLI���G��fy��'�b�ɻ.�R���%~�b��جU��'O�'9�I��M;���?����?��J��K��<��@Un�j4�iK��'v �[��&aӨ�&��+F���Vl9eK�[�|ᓯ*?�rJ�4a�����A̧9e��$߁�?9��T�^N8��\b�ut�� �?I��?A��?���)�O�`auA �(��0�.F�?p\�w�O�@l�	3��ɔ'��6�)�i�قvK��B_��#�kܽ[��d*�e��:ܴ.F���v��D���x� �}� ���FI�D�\�&Cc��5tN0y�䀐����4����Or���O�䌨RՀ̀tǢ6���)֏
N�:�������O`�?�ҥ�:-���..�\�q�*��z����'v��'�ɧ�O�R�	���A�,Q�׊D�L�����2$�����O��!�=�?9m5�ĵ<��lX$�3gfR7�D4�%����?Q���?����?�'��$�妝C�Ɵ����F����s�=	��h���f���4��'H��?���?Q�k�r�zlxƃG�a4�`��� y � �ܴ��D g�<������O�W�H=d0�� ���92jȡ�y�'[b�'�B�'B�����	�	I9Lhd	��V�h�0��)Oh���؟�R�?��ڴ��Bn�͡�ָC�"!��F[9}�`	L>���?�'b0��4���Rs�u��j�*Z=�Mqc�G�.��R�D�?��C?��<ͧ�?9��?�Ҭ6��rFgP�;L� �̉�?)���������/	ȟl��ޟ4�O;���7�ݜn���"��	q�l��'�"̴>����?�O>�OG$<!$fܼL9�a��'�-F��#���k���,�<ͧD���	N�	&30����a���a�op��A��� ��̟ �)��IyB�a�@ę��n��s�ܧ$-a�	����$�O�8n�f����OP�D c���,O��d����S�&ܤ���O��耎|��.?=kC��?]��e�7*m�� 5��w���<�*O���� <@��\��G[(R�R�diJk��po	��|�	�|��B��O,��w��c���1v"}a�ܲFK.�I��'AB�|��TɖH���?O|ԣ0mU�+���i� !�8y�8OT������~b�|�Q��'ZruiQNԣuanq
N�"<�ÓT���!F'���՟ �KV����=  ��HR�b��I��\��U��'z k�D�pb�v���-���Y=T�x�B@&3[R��N~����OF����gG�e�&W� ��D@���� ����?����?Q��h����W�6������5�Z�AĂ�E�d�dHԦQ�D��Ky"�qӎ��]7[$R�ËP!'!"f�z����T�	����Ϧ��'��PYD�^�?�H	� Je�DOL�G �Q�ҸZ�$�{�4��<ͧ�?����?���?��A�1F��[��ͼ,����
E=���Hզ%���������۟ $?��I4����"�I�̎H�YIt��O����OڒO1�F�sc�P��])"�
48���W��O@AQe��tA�܉��Zr��Hyb'��`p� K�	���i�'L��'�O��ɩ�M3ǐ��?�ac< "�qBŅ�<zdc�@>�?6�iJ�O��'E��'6R�� �A��Qgj�÷��3~�e+r�H�M��O��Y�Mŵ�z��4�wp�a#����\	Q���S's)�(Ә'���'���'%��'\�,�pl�9 Δ%a�-�4*y�:@�O.���O��o���$�'�6�9����dM�ic�Fz
��'޻��,$��I̟�7��PlJ~rG��&*ZD���T�C�l���JC�������(9D�|�S��S�����ß<��e��V��xBC�$Y�d۟��Ay��i�h)�&Ǹ<A����I�P���,����֭*�I�����O��D)��?�	w�әx�X�Kq��q�p'<-�b���I
*O�I��~��|RNY��x�;��XD��3�S�~��'�b�'c��t_��2�408T�Ʌ,�=/��G$�
-x�Õ E�?���U����Q}��'I����|����s'���h��'��9
�֕���<>n�i�<���E�xZ�t9B���b/(�a�M
�<�/O��$�O����O.�$�O8˧n�����cal{� ��Nh��#�i����"�'�'5�O%o���@g�<qcHS�j���JӅ?
���d�O0�O1��,[�CsӺ��=V�U�s��(aH,���ɵ!�.��A�'��'���'��'��<id�Jq��d�s�̬(]x��2�'�"�'��P�0��4�����?q��l�zN�"T-�X	&
,fyq����>y��?M>1a)�]�عh`�֪�r]�$�c~���U@�Y:NX;on�OU�E��9o'�g�Qi��*��!GJ�
A�$aX��'���'���ޟ��V��U�Π"T���0<Q2�۟�;�4hy���?i�i��O�Ԙ)wtQRT�d��-�c*O-��D�O<���O���d�J�Ӻ#a�ͭ��r�S�Thp#���+�6�5��(Ю�O<��?���?����?���8����J	��P4�%H,��H(O��l�81b,U�	x�Ig������DI�G��1`��Cn�,E饦1����O�d*����`&d5iB��3�x#�fL3L|�41��m���'b�a�ӆ�h?�O>y+O&��� tX(���	7_�M����Od�D�O���O�<9��i���x�'�(�CDNY�D� �h��9*J�I�'$�7m8�	:����Ŧ�i�4G��V'ID�U�����4�b��A
� E�� �4�i��I(\7�ir�O�q����.7�Xı�J�yq���VB��E���O����O8�$�O��S�'~
�(��Q�I�D\y�"ȭlR<:���?���" �b�G$�ɗ�MJ>���[@s$��F̊�3k�a��ћ?��'hұ����|7�Ɵ��a�&�"�t�x�g�;K�{Z|�C@e�?q[~�'f�i>e��������L��ə/ȸY^Tr�G�+1�ܭ��۟ؖ'�6m�*8��ʓ�?)-������^�<��G�P�DK��0��H#�O8���O��O��7,b��u��z���E�~�4y�&Vl�Ĭn���4�(d��'��'R(eY���D�1��p<����'3��'`"�O1��Mc��s�H�J��L�qm̫�@ h�����?��iS�O޵�'��&�Fq�$�pC��u|�zr�8K.2�'ʊ�ꗿi���?I(��%ԟ^˓|i�EB�&�o~9��^�$�͓����OJ�D�O`���O���|J�S�dZlB@M�31��uBꄚ曖CM�'LR���'�j7=�$I�v(��n̹�a[�tip���E�O���<��)�TF|7a�Ԩ'�T�p�$��HX�Q�Qg���L:��	QC�Ey�P��S��T�sZ܅��%���*OR-oZ�Y�b�'��D���j��`#��H%�u0��ӈ%B�O�<�'{b�''�'޺eҐ*ԅJ��c7�֦p��y�O�5Y�N��f�~���2�I�?����OVr�����)����5m� A3��O��D�Oj��O�}r�IG���f�$h^�Yc�b�0-s�����hD�/�k���'^�6�;�i�mp�dI�9��8�Fװ0e��@�q�$�I�,���W	�MnZF~�,L+?R8�S�%[�Т���,<n�I�5OĬ ���餕|r_���������4��ߟ�K�L�)o�4;ǠԡHܶ�)Smyhy�n���E�Oh��O���l��	EKn��=n?�Z��Ǫ-����'���'7ɧ�O�l��!�J�-Z�I�ae��fY�G&K!F[��H�OP��O��?I�`+�d�<�0�qN*0k�jϝF�@Ā��?y���?���?�'��D�ڦYX���ǟ�2Bb *g���i��d�Bt� n����4��'�X��?����?��gZWJ�t)�ږ@����b�l���!۴��DG� �N��' ]Z��j��M�FKdYS�M�>/�-�&��=S�d�O����O����O��D,�S�l	�ԅP�~���W����	Пl�I��Mk1�ӻ��d증$�𱖧�T�E���8@݄rի����&6-���S�v��im�[~��ڈ�� ���v�<�I��������LB�?'�3��<ͧ�?1��?a�o�0(Dd��3���Y��02a���?����D�Φ�in�ş����O-z� RM�$#q�RN>S|ys�OzA�'��'�ɧ����i�(�a�ǲ9��#'&ԥ_��8��l�"G�d7��ey�O2)����F�4Z�-��).��Gls��	���Iğ��	؟b>ݖ'��6̀�$$	�׹rP���Z��ZV��Or�]��u�?!�_���	`a@����	P���DA�������������'���p7#�or)O���t%ժ �x ��p�Z !3?OX��?a��?i��?����.N^d��/R�7J�L����)�RYn�>hb�Q�I۟���x��۟����{�)��;�r��3�߃M�U��M˜�?����S�'p��q�ڴ�y��E�@R���1�|}�����y24Lh��䓦���O��ąb¢��Pl�42bN���F@`�$�Oh���O,ʓZ\��J�1�'2Ŋ3&�Y�3J£)nt
U��^�Ort�'�2�'�'���a��6ո����ɢZxD3�O�q���Ǉ~)���F�<�)E�?�F��OĈQcO�s,()��ޛ0|�ë�O��d�O��D�O��}"��Db��<=�V��7�M�DQ#�Z���	���B�'E�66�i�*Q���v�8��F�	�p�P�l����L��+(8Tl�S~Zw� � �O�:���Ԁ�åkĈ2Ȱ �5%c��Iy��'n��'5�'���`ā 
�p�P�"��y4�;�MÔM���?���?1M~�-�6� �/�'a�[���h�Ա�Y�<��ʟ`'�b>i��e��)*t�p�,?���"�� Nn�=?9���A��D������d����0��&�ɲ��!|���$�Oz�d�O�4��ʓS��FƖA���Z;24�(�2�	j�����m�?8B�k�h��p�O����O2�d˔D�:C��[��6�C(%�`ٔ�s�L��x"��?%?y�����<��a³7�TP�#B�5m��ß<��͟4�	��8�I{�'d�T#���6>Z�u�D�B7
�xk��?��l��	���4�'��6�;�Ēw�ԑ�D]�}Q�YCA낢D�(�OH���O�iջXY�6m ?�$�պg��QD ��E�*H���,?nLmo�S?N>)(O����O����O������4�p�IwO��0��O��$�<�p�if����'}b�'W�Әc��H� ��}J e�%�5��R��	՟��	d�)��
�>�Ҽ[��
'`�`$a5!����1��Z��Ms�X��,?��$8��[�g�Y���ZR��{Gd��l��D�O��D�O���I�<���i?n��5&]v@p��a��h%�p���C�X`剝�M{����>yűi��5�RȞ;e��q1�\�7�Hcs�y��o��`�XoZO~���e���SG���{�~��a�62)*ḤŘ�2�d�<����?��?����?Y,���A�E�M�vݙ�`NV����Ԧi�E�������%?�Ɂ�M�;;Ѯ�憓ME���Ӎ]�;��ų���?�L>�|BE�ɨ�M�'�HP:���=a�x7'P\I�ă�'�.�٣&A͟���|�V��S�����i�t^�5@G� �<�a�h�����	П���LyR�x� �c��O`�D�O"4+u�̗-�����/L�1��8�&G"�������O��$-�$Q�	� �ZȐ�"��]�I N��-A��+b>I��'��I72���A�=�n���HC ������	�����r�O�b,D/e,B(��\K���4~��d��|y���OR�D̦��?�;fF��&�۶���,V�|>͓�?���?���	�M��O�n]�v< �)1������/I���ʁ�U��FI�J>�)O��?Y�`�Tj�(U$�+EF�P�
�q~�.mӘ�	���O����OR�?%���8�`��萱( P+�K����O���:�󉌖3Z�  ��p � �ׇE�Ъ1$oӠ$�'�>,cw�VL?L>�*O2E���ş/|X<��&ܿi���u@�OT�D�O����O�i�<14�i��3��'��Q��1r���*����X؉�'�27�4�	���զar�4F��6�L51�2d�f��S�R�YA�@�{S�}j��i��I!���Oq���N�,��4�#�
�L�bh�3!�}��D�O����O����O��D"�S�b�^����߄����$_q���'үw�2Q!�?}C�4�� �e�&��l��Q���7@��A�x��'��O��2�i+��p�2�Is�3�4t�ť�)("\��5`2LG�	_y�O�r�':b�×TL@a�`�(]���PIٜV���'N�I6�M�T��?Y���?�,�4�2'�1d�.u:��̠!$x�%��la,O���w�B'��''~�㖊�,I�H���BCT��pZ�G���QkVz~�O>���	�t]�'o4ɪ�-Q�n�!�Θ?VɅ�'���'�r���O����M�&�4S�i��]�l��1� ϔ�eK�8Y���?�`�i�O���'��6-W;rx���.R�Z�4���=q�o��MS����MK�O�*�Q��J?u�$IG:z�>��G���j˷���y�^�H�I�$��蟐�	Ɵ<�O"h&��,����r7����dӴ���@�O��D�ON����D���]z�x�2D*ٜ��!ǟO���Iܟ�%�b>�ZUA�馡�S�? j��`�#q�b$[�g�W	B�=OB<���2�?!�`9���<Q.OP�6�$l�<��ӫW�X���'Qx7�\�;�r��?�� I*v�T��QA��djQQm���'���?�����wn�gD�`��t�Á��+�XE�'�����H�^�r����������'�H�u���N���Y�"�I�Z<�
�'�P�C��@�R�J��B�m
g�'� 6m�H����O��l�Ӽ�s�W�e.�+w�YCFБ����<Y���?Q�TP��	ݴ��d��1t�h�O;�x�TF�� �4��[��ݻ&�|bY��ER�̩K�p�򎚾=�(T�u$ܤ��d���*qɗП�ͦ!��x��E*��z'���L��Q%�[4mŮ9�S������`'�b>�C�� q�(��n��,K�(�#]��o��@�>�Щ��'K�'��I�����E3J I�-�,9��h���T�Iߟ��i>)�'1�6mO`���L �hf�ƧGh�HH��3YB���ʦ��?a�S���	����	(:��i��f�
y8r�QPK�pA�+����'d@-0B��OBI~
�;�Ay����D=�e`�7/Z����?����?���?�����E��_4��9�h�F��p���0�?���?A&�i
���O��bsӂ�O(����T&~��2'
�B��"��O�4�:���s���Ӻ��CԮK�t�NY�A��b��0:�j��^��Ol��?����?Y�r����X��VI��G�ؐK��?�)O�anZK�q��Οl�	c�T$���k")}��I�����X}�'�b�|ʟ�P�Aڵ�d�ˎ;�`�p0�^
!N|r�'I;K��i>���'��u%����'�h�8��'�Zv "1"2�����I؟(���b>y�'�x6�Yk�M.&�jC"�7S;��1����Uͦ��?	CR��	�IǄ,��Y�t�c2Mׇ<�����:�LҦ��'��A8e��?e�����`�Y�:��80����1�(#:O���?y���?����?�����I߰T#�p�d���I�ɒ�l�o��R������h��|�s�h�����#�'~>�Ǐ,)>ĝuި�?y���Ş'X��8ش�y2J� ^r�$ �%�̔�˯�y�%׌QP ��ɫX��'U�)2HU*�vD�EJ$��BTTr�P!�4i���h���?Q��c;�0�A�d?�-�BD��:�
q[���>1��?�J>9���)��Y�`�1O�=�5�e~������iƞ��6�	�'�"�^[՚a4CZ".ռ�(�,V�R�'*R�'X"�S쟄b��F�E2�o���j࢐�R۟�1ٴ�b�C)OZIm�X�Ӽ���ˈ2x�d���Th��G��<)��?!��]��l�ߴ���D(=��9�'*#2`�W��@f�ҩ �VYA#�Į<ͧ�?���?Q���?`e�S�`I�%؟n�N\(�����ܦ� ������I��$?牬[B��T)��p���E*��1�O
���O�O1���0@�K�InDY��ν
d�t�������ē���T��?'2�GB�	Ny�`��y�cV3 �\�jV�XV��'}��'��O��I��M�	��?)���	н邬��X�0���
�<釱iV�Ob$�'�"�'A���\�D�""�-o|U��o�M[�O��V���b���w'>p�`7A6��&ݽe���'gB�':r�'sR�'R���B�#Ƭn���
��Ĺ>3�����Oj���O�,o�+|���͟4��4��XZR|�	H=5}`�`⧋#P_��M>a��?ͧjn"P�4�����|���˧Cm(-3u$��P(�IE��'����Ӳ�䓓���O�D�O��׏���0��ȩ%�!�֦�&Hc����O&ʓl��� �XXB�'�"Y>�)Q?G�R��]4��۲'*?9�U��	�'��'q�f�R�N )*�rrm�,W�ag,��4b�d�7��<��4���a��J�OJ��� �:��VH�4Y����O����O����O1�4ʓ4F��GR?N��`��L�2qp� @O%3T*��4X��J�4��'|p��?a�/��J��d0��;��c����?���\d��ܴ����:d�����#*O��
f��fJ^	��đ�J����5O˓�?a��?���?������b%����+@%<-��"�Y�[�m��H8x�	���IG�S������!��ex��h�dC�X(�����?Y����S�'Mp��ܴ�y���
���U�2V.�4C4j��y��ةY�29�����d�O.��V&*ո�A�mͧ3��m)�%��1�(�D�O����O��_@���U9c�B�'��g�<�laOW��'/�Up�O| �'�b�'�'�؜bԀB�Y��uQ !

a�D���Ol-��K&�46��x��L$�D�Od<�&d��4�h���=:"�$�C��O����O����O&�}����Y(���7��Ҏ�9	���$���� �z^2�'��7-)�iޕ3��ҋ@�bq��c['=�r%��$t�<�	��|�I�PA�Um�q~�I�\��%��b�I8�ݹJh��
�ԥJu�%bL>!,O�D�On�$�On��O���&C��3�`y�h�1	�=i�m�<ჶi��AR$�'Nb�'9�OLbM�
7�2�*���,��p ��K
g��?q����S�'ij��� �㠇��kp�p ��	ˤ�ѥ��Pp�'0MYVl�o?�N>1.O:�Qb��b��Xڱ`R?K�t`I+�O���O�d�O�ɭ<Y�i�B����'�qt	���x�ϖW���Q�'WB6-#��&���O��d�O�Q���q���H�(J� ��	B�w�6-??�,ا~U�)=���QcuBV6Q�v�;�kڮ
�X���`����h��ȟ����D�
�-[1k��U�`�:�pH�Fٵ�?����?���i9,�\�<�ش��^�%K�!ߑW2 �⧁D�@��M>���?�'$[ґp�4���W�k�laQ!�8$~�[�#�63x��2+T6�?1A�7�D�<ͧ�?��?�$��&1`�_7���@�3�?����$�ɦY�A�E�����؟X�OA8d� $ߘ,��MR!�2Y.��OB��'��'Dɧ��Y����֎H-�|l�ڏjJ�U8���.f��ղ����]���O�	02f�3�V�Tp��Sg�Ex�U�I؟�������)�Shy�i���� ��*�|��܂��; �`��`�O���]ئ�?W��	�#�2pI2.G*>�C�'�&�H��	՟���˦-�'U�\�a���?ͥ�4Maΰ�M��IA,I��-k�cx�ؕ'�2�'���'���'��Ӕ%�2)y�Ax� ����h}8�4^:�����?�����?I���y�/��T�Y3�ܾv��x[��_�zy�'�ɧ�OL�G�i��ʭ[��G׺ 7n�i�둵V���)^�+�'��'����|��^u��p��;Wct-�o��I��0�	ݟ��IП�'8\6
1�����O��Y�t:�W삣=A@�
���j��OV�d�L}��'���|��\Ŋ#�hհL0"��ҿ���ѪL!�A�s�F�z7�I���7|�d�i�N��V�ʕ�Д1�ER�����O����Ob��7�'�?���^�~�`i@d�Z�b��-��	��?���iȰh�c\��J۴���y�m쨋U��'��<ȑ�Լ�y2�'��'W��i��	�>;r�3u�OE�]�E�Qq�d ���,7�Ft����U�Imy�OQ2�'�r�'p�:-Pt8U�C,']�;���F��I�M�e����?���?!I~Γ��QSB�U�zcf�F�q�����g}R�'!r�5��	D��Ri�O�N� ��I�:�d�BAR��I�Z/�8��'-R%���'�P�`�
�3y,�Q'#F�w����'�"�'R���X�d�شFe�����|� *k_�12ƣ p/����B���$Il}b�gӀ�lڼ�Mcp�Q0d�PQF�pB�Y�o�j��a��4��I�T0�A����O
��A�
�����/%8~�R���y��'"�'R�'�B�I@�hK}Zf�@4�c$�X(T}���O�����uˀ��@y�fӐ�Ob`3��O�@��vA�_q E&Gv�ҟ��i>�#��M+�Od`�ͅ��1R��֛�ܫ2�5:Rx����R�n�Ot��|j���?)�s�2�P ��wRF)x���\|����?�-O��l��)�BX���	E������I��d��1�a�d����d�N}�'��	>�?�*�ȈV�Y��� e�����խ"Ќȉ!�]�5uZ��|3��O��H>�E&1�u���Z:�h���?����?����?�|j+O�!mZ�N4X�Q��ݵRDv�෡2X�*t*A�UZy¯}Ӝ���Oz��H�B�֡#*N�{`ʀ�,��$E�-3Ʀ��'*Bi����?��������zʸ{�N�w��<�R?O�˓�?A��?���?Y����	Ĩ3H�8©�;��1K$+��<nL:���ßP��H�SßP���oΉ0r����ն�2�� d��'�O1���AC`�4�	�;���P�fQ�(�nH2�/Ю�h�		4-��'��&�$���d�'�0Ⱥ�a� A�d5AP�^�>U�\�$�' R�'_"P��y޴4$����?��qx�Q�Ѫ��Q+%B �p�9��>Q־i�:7�H�I>%��I�9���fOr�H�q"��E�Q����|b��O��A�"���e �2k����B�K���q��?����?����h��NI!�,��bͪPR�����J�Ҍ���ɦ�4bJԟt��=�MsJ>��Ӽ�*�#j�|��_1��T`����<���?��[�.��ܴ��$̶pl��OAސ�4�	b�n�cgJȤy�f� ��|rZ�$��������i�Q
tñ^�h�B� ��C��QE�S`y��p�\0�O �D�O`�����.!Dr��Us��e	�`��'�2�'Jɧ�O�N��s`�06���T�ޒB�Ȱu��y�f$�QZ�p��Ɩ�P2�{��dy��J�榥y�.�:�0m&f\e��'���'|�O��I!�M#%��2�?9v\��`���+X#&�ʤI�?9��i��OV��'���'�r@��_C8�	�FIb�;�	���@$c�i3�I'NbLX�ԟ.���NT
ha8�qGɋ>z H:r��?��O����O���OJ��*��43��Uƌ¼�U$i��\��ݟ��I��M� ��|��U-�6�|P�BA�8�P"�A)R��8 �|"�'��O��9bs�i�I?Be`�Z�,�K��e�w�E���%L-5��:��<����?����?Y��]�)l|Y#a�J�E ƙ�?Q�����ʦ�iƆ�۟��	���OT��a�C�|A�5H�80.��Or��'�B�'#ɧ�� ty��X���������8 �3�A�g������w�R����ΝM?iN>�RF��}l<
�h��/�J���&�#�?���?���?�|*O,$mZLX��{�J(�rGdχ�R4Q�m��|�	��MÈ�ʽ>i�c��t�"�xtbc�!q��0��?"n���M��O�C�����P�d���LD��PP�H��H�,c�4�'!��'@�'.��'��8��t��쑻(���
���H4f��ش@�8Z���?����'�?���y�ˎ��1@&��<\x�Õk�Q���'�ɧ�O)�H���i���v�vX
Vh��T�HYD����D��@�,��'��'���t�	�^n����*��%�q���	۟��	���' �7-��3@��$�O��$ExH}��'�&>m��$�1%�X⟴��O�$�O6�O�E�B �W*x��%��!5<�������NP+6td�K&�ӯ6�K����ܷ*�p|�$�+YT����Dϟp�Iҟ,�	���E���'M���P�3#�طǈ=4��'j�6m"�0���O9mZZ�Ӽ[q�؃=�P��%�?�M3�Dw?���M��i:�*5�i]���&�	0�O��j� M^yD�aRf�!+�&��#NB�-|8Hq�@Z��ꐮ6�t{��q$����cW4?�v9ʢLG�1DH+�dze,)i�ē	�����K�,0�A�� &�ɰp
Z���(zS`�Y �%x��[����a�d7+��˳��1&�@�]� Ch1;-�6�l�¯���i��9�J�2��;2�B��a�Z�ɞm�Ҏ�R�+0��8�~T�Sk�� q`�����d0hiD�5�NP�
<��ik���,�.�8�hѕ]n1X�k�h�
Zb��6*A$�`�")Đ�hŮ��'baoȟ�I���S����X�ڴh��6�n�ae)�G��o۟��I�(���?�����)�ʁD�6�0�bE��?�ԧ��M���?����S�4�'/���Y����"J*<�t��G�x�$�bU��O�'�?	� C��e�P�b@��:�����v�'�B�'�6J��>�-Ol�Ľ�9���$g�r8q��Ǻf!N��'�	��^Q$���	쟰�ISv`K�")�� ʐK�&,Z��ܴ�?af� �	Zy��'cɧ5KD�"��I$���B�ʅ#��D�5,�O��OH��5?�Х� �r�B IN'=}�P��H�	�))�O0��?IK>����?��%N
{�Բ��H�Abl)�fԬ6��<���?y������=Y���.i�4��*�>m��r�b�2u%�6ͽ<������?���3&Np#�'B�b!G���!�;!Sv0�wf�M}��'�R�'��		.��O���_	zP
"�%���,c�}��i��|�'��&�.�qOF��.2h��:�N�&C��R�i��'��I�{����O�r�'����]-&оxa%�Z�\��2�,^P)�O���O��R3�:��JBV��1���"p	/#�"t�U�����'($���io��'q�O����p�<L�x��O�*E� A3�+�榙����XԮ�a���Ocr#c��^�����O��W�X���x�T��4�?Q��?������cyb�L�l������&��3�S�e��6-�^�����<�D�0�ç� 	AC�i��'�B+�!�N듂��O�I�L���He��7-(@�d�Ck0c� �$F�[�	Ɵp��ȟx���
,~ـ��I/�����A��M���
i���P� �'�r�|ZcfqF��<0�V���-��	�O�\"D%���O��$�O��-¸����!i�����J$ 1Af�˞����<i����?a���1s���+��I�b&98T���O��䓹?���?�*O�"A���|�p�/�iC!O��LT�t�q}��'*R�|�^��蟰b�n^���Źr��p,>�#��A���d�O��$�O�˓`�BP@!��4�F5J���&��E ��a�j�<7m�OؒOf��|r����8��і-ц5��e��敞PVd7-�O����<9��،�Oor��5V� "�p �1��c�ƕ�To������Ox�d,�9O��,��M[Pd��"%��R��΁6���U���d唭�MC2Z?)�	�?y��O�a���$l��MKB��O-��B�i2����� ��'��禩�$�ɚz�xೇB�t�6t� �iӀ�kB�Ϧ9�	�@�	�?��I<�'8MH����c�&i��ȯ3 �=z��i���',b�|ʟ��OJE3�N�	�$�K����|��P�g����a��䟼��'v�N�H<�'�?��'_����f�0S)�4*�f�to�Ecߴ�?N>��^?��i�����(�~HK᠂�}ux���4�?٤�����v���D�$Y����2鐣�v�#w�N<0�$'��)���Е'VR͇..|> ��`M�m�d*%ȉ�
����W���	�0�?����~�%K�!Dh��	3"����U;�M��kW}̓�?*O���A.����&���B��4p�Q�'Q�O�R7M�O��+�	؟d�'�$��4,�PтM7�Y[E�K�3��$�\�I[y��'��U�X>E��*B\u���?T��K���)��f�i��O����<1`��P�	�M��+��@�%-2�a�"I���6M�O�ʓ�?!�����Ot����k숭|�<��T-�Q�ޕ�!�ȃ(M�'��S��.(�Ӻ�td�IвL��kQ�+�$��N}��'#����'|��'Q��O��i�� Py�����h��Տ&�H3�i��P��"ׯ9�S�S2Z�r5r�iC�2�0�a��aZ�7-�{Ϯ�D�O���OB�ɺ<�O�r��ÆFn8���E_YP| p��>�4�r���Oeb�C��RX��c�f��aۆb9K�>7��Ot���O��v�g�i>a�IY?��/��'R͉�.��7\Ȑ�G�ᦱ�	j�	���9O@���O��5`��03�%+R����Ӡ4ڸ�l�ҟ�0�FE����|����Ӻ�1�D2@�@����q���� k��꟠�''�'��R�X��و@��J�MG�
,���L,ט-L<Y��?A.O`��<�;	"��ҭ�?�(t+�e�*}LmZϟ��'���'u�Z�L�%�����z��Y3S��/�H���,о����O���,���<ͧ�?)R�5
����@Z',�Ԁ7���S��'
"Z�T��,w�8�O�2�Ԥ2Z^����.�Q��ϪA,7m#�I˟h�'��%�L<���݃�Ā�6%�,Œ�!&H�ܦ=�I̟��'3��@w�!�	�O�����0QΊ)�h黴�06f,(0��xbY���i�M�K~�Ӻ�P�4~$�HB���<�Tm���XԦ��'��|IGk�$E�O�R�O���_�$�y�F�*@�|mZ3 �EY��l�Dy��'r�&�7��i�jr���G�%�t�W�-]ĥ��4����Ÿi��'�"�O^O�I��<�^-�D!~��z�$�*�L�l��^�B��	П �'���y��'�� ��\��I`u��:c� �qmc�����Ol�d�4^`�'��Ɵ���[c�a*���P�F`y��V�%�~l����	�L�5�s��'�?9��?ᇹ^4t�T�ûW_��p֮�$p��o�Ɵ�3f�K���d�<q���D�Okl fȈ�5�T�4���Iݿě��'>�4�'���ǟ��	ǟ̖'���9���mQʽ��ϋbR(�{�3f����D�O�ʓ�?����?�tC�_��lF�>�䈈�({���ϓ�?����?���?�+O��Ń�|��\2M2���P �"�|\��L�����'A�R���	�� ��
@|�	�'S�E��ǐs��@犇�(�l6-�O��D�O6��<�g
�9x�����@)�e�"�H(��3X��lQ"��7�MS����D�O��d�O�]#�=O��禩(�%J�q<h� O�?�Tlh$Nb���$�O�˓%;搻%U?��	���sIp��ǃf'\�9�/�" �!XƠ�K}��'"�'����'��	֟���W�t�E���O&��tϕ5�°lZXy��	3{�7��O����O���u}Zw	l�y��
����'g��Ua��4�?���^6�̓���Oz�>�c�"��U]��p���<fЎ����v� a���Q��)�	��|�	�?��O�˓�"-�e��X��X$�����`qкi.|x�'��'��n����*�H
�"�7jR<�U%�*T���l�̟d�IdO#��$�<����~2��8��y�E/n4�4r�T��M������P^��?��쟬��b謙�K�6`p�!���!�"0B�4�?Y�.��@��	ay��'��I���?��yyb- <XI����xbX7Mg��
0O��d�O�D�O�d�<1��ɔ"�TMP"���� �j���(H�]��'A�Z���	ӟ ��

V�)te�#��$`T�Ղq���i���	��I���_ybA٣B��(i��`��q�"|)#ɗ�c֊6-�<1�����O���O�y�S8O� ����6q9���F�/p���oRѦ���������H�'Z�(Ђ;~���/���&�����C^�}m���'"�'��L��y��'���Iw��z��
�k/L��"�@���'Ub]�\JC������O�����=���Q�1q��Ǯ	���bĤTE}��'=�'!��'��S����,��,!�/��[���9��yn�Zyb�`7��O���O\�ic}Zw=`Z��m���s%�(:yaܴ�?I�7"4q�����O �R��/ ʐ�I��9=��ش���ĵi�"�'���Oj����đ2ɮ�Z��W>8��f��>o*)l:b�����*�러A���2i��c��P��+��M����?y�x}��v_���'���O�X�C&ٞ~��b0��O
F��t�iw�_�xI��a��?	���?�CF�!	� �i�!�+#y|���oɛ6�'}d�s�K�>�.O8���<�����L	$u[pBB+�&�L����q}2̏��yBZ��������Iiy�-׵v:�c��@ �*a��ǒ�4� 9b7ϳ>�-O��<����?A�,0�,#�!�A����5(��)����de�<)��?Q���?Y���d*A-�T�'D�z���1N��ad��g�nZMy"�'o�	͟���̟�"!g���>Ĝx�U2˸����	�O�r��?����?�/O���c�W�4�'��ɍ	O��I2��Q��(��a�����<����?��V�6̓�?��'R�P�#Ƀ\a\Q�F$= b�4�?�����o���O]��'��D(�P����B�ԘQ��F���?����?�!��<�N>�OXZ�� ��9@�(�"5pM��4��;��l�؟���ß��������BTJ�[T,�7�!A�YѾi�b�'�x�k�'+��'&r���`����j�X�hi1�؛6��r[Z7m�OF�d�O��i�k�`�Ɋ�.Q�%�����\�����i�uК'�'��4�dQ:i%\�r���Y�*����a&� oߟ���ݟ� 섢���?!���~
� �)7퉯G�6AC�'Ai����$ϻ1��OZ���O���ܴ:P�a3��u��Qq)|X&1m�� s������?	�����S2�S8�j!B�!L(8�#�C}BD��y�P�d�I�����ByBbO
R֩BA�	�#8��ҧ�e��(�=��O���=�$�O��D�.�H�#�0�������6��{P=O���?���?�.Oʠc���|�#�� �n�h�I�AB��Y%��u}"�'k�|2�'j��+F��K�	-���@�ۂ1��I�^��V��?����?�,Ol�R #[U�� �t|��l�Y�I1�NYe��dJ�4�?�J>����?y�ʑ���'O�8����
���(K0RH!ٴ�?�����'o��&>e���?y��K������<$7by��-dA�OD�D�O>�D�s)�$$�d�?�e��)r��	�Q|0��C�tӮ��䌢��i�H�'�?��'����/`]�`��O��E���ς�\7��O����2�D2�S_U��y H��I�Y���(('\7&<�$l�џ���ɟ��.��'Q���jN�b�%JRc">@�!��xӐ@�w��O`�OZ�?Y���9�^`jqK}{�؄8$"��4�?!��?�V��'���'�)fZ�rd�R�.DEh�,����|��P�_[f�D�d�O�����p	K�J��K��2�eL�b�.Hm����ރ�ē�?������	߆&rF�����A�^��B�O}R��F��Z������h��jy�_G5�����:�z��@�H4J'*dx�,;��џp'����џ�J�!�@Vx��h�]��82�X�r�����wy��'�ґ��a�
cY�瓱v�,x�c�4yW��sh g��듟?�����?��0�����8o�Y���Q��U���02�͸PY���Iʟ���Ey2�Q$j�d���i5�5Fw�\b��+.<
�����%��Q�Iǟ �ɸW&H��a�d�jtҸI�a��t���!�bo���'��^�Ha -C���'�?��bt�R4ɂ_"�ԁǨ��ݨ@r�x�'˔���O���?DE�`�P���;��a�l؆��6��<a�%F3���˪~:���6��P�̙�-(��� �yؤ��Bi�>a����;����S�'}���萾@SЀ��
�f��mZ4�ߴ�?���?���U�������/R	�2�G���@�u&��?���d�'���E�4E�.�i��"A�q|Ӓ���O��$�6��)�	�O��	�.>�-�R�	�n�~�� �A`�\�yBHхJ�h�����O���m p�!��G�ptb�j] ol
@l�@L0�ē�?������ò�/�đ��I�"�����(W}}�HJ���'�B�'="U�ؘ �E2xX��(v	T�s#��l�Xd:K<���?QL>��?i䠑4a�Tl(ĭ Ժ(�Vf�#,�*�(��ӟ��'=�蒌���P(y;¸ђ
�&���k�
<B�'X"�']�'Y�	x�4퉰�k�`���		]����E�[�s��@]������h��ğH���s���	Ɵ\�	Li\��`A�i�܅�Cz�~pp޴�?�L>�����S�'l2�%�L�>f�f��w�m�ܴ�?q���ˀX�&>a�	�?Q��C��u�S'�4V��y�vGҕ�MÊ�9�����i�\I0*�(X��s%O�Z��y�ش�?���M�ȱ��?�*O����O:��ƴ0RFU	Z->-��C��F�E)�iCR�'��K!�ט��O���BgȞE�e#VB��7f>h��4-7t���i���'�"�O/Rb���R�ܙH�����U8a6�	ҁĦ�M�p�C�'d��DD�*�RB�ǡpF������h/$�m����	ȟ��Ʌ����?)��~��>�Z��ׂ5R:��lM���'�n�ӋyR�'�2�'�xȩӡ�~f}�J�܀����u�0��Źrf����ӟ�&�ph0��)T}�(Z��@i����%����ć"l�����d�I˟���ly�!G�|T��K��Z��3��
��0`q�'��O����O>�8S�,,;�+��l!c�Ʀ2[,b�$�	������	>,7`d�'2Hy�T��/\j�T�S>l��l�`yB�'��']R�'��YCwۦ�M�[	̤�b�H�#�i8��)Y$�	��x�q%�'EЂei0�)�'my�2�M�YиI��iȑ��T�ȓ7O���%ݍ�fԛ�J�3-�rY��j��dc�R��E!E�/p�b�/�C*ޡ�u	ZD��1Y3���.��X9��V�Y.���BB3�ܙIbi��e���8���U���`N���~���Y�mFFQ[DO
�l���l��KH,غӡ�0Xl
�c�`͠��� .��d�՗������w�j����8(DXw/�O����Odȹ&�@={�i�z-
E��H�\��hB�e�0����Dd��J��t��O�1�GJ��:�`��̟C2l%��-�?Q�4��鋴�0�qv�Z9/����֬�:��dے��wc&��񮋓}@L��Æ	䈸"1����"�'�)��'�dCO��Ux�ܥ`�|bD`��> !��N*%��+�Z�,o04�O�6u��� ���?�8@�7(���KDء^����ϐƟ��	}���N�̟��	� �I��u'�'>���=FHV9�B��'"&	r
��D�d_�C�d{Ӥ�8�b ���hOT`	�D��oԎ\���ʖ���1E��ϟ���MZt�;y�$(k��hO� ���!��04P�B�%�.��@	E�O�e���'R�Uy���8tB���K=�8d(#���y(A�7|�PbJQ���mHu%E"~�#=�O��ɇ.�VB�4@PȣB��#:�Iȴ��0vP,
��?q���y���"�?����H�+D�b�"-R�q��Ύ�KiN�s�gD1t��)��(/�0̆�	&��J���D��xXE�ãm��0{���-᜕� 	��cd����'���S���?�q��.f���m�6�z�{rJ�_�<�wD%L}^@��n�P�*�Ӓe	u�<"˞�4�H�b�?,3���D�<����d9(��'"^>]J�ݗt���G6�0t8gLՃ@�9��ʟ��I�[�����G�L)ɄQ�ʧ6����!�`&Ts�A�r�$`Fy��;�:�Ѳ'IPH��>-�7 ]}?��TDn%h��&1ʓ-m���ɟ��� (%ZS"(�t�ܭIa&���Ņ�<���5AP=[u �xQ�i��nW7h�bą񉙉�B]��ѮP%������\<0ÐAϓ�ܐ�Q����p��Ɋ!RF��'��/\�1Y�`�5!��	T��b)���ad��S�(t�^�T>-�|�	-:tJ�P�;e�z�q�K�9xZ�"�!��Hb��΁'��$��S��?�ӡS�8��|�P�pk(���ß0��r~J~�O>��b�+x�%�kֆ<���00�W�<�K��C��E�v�ѭ#�n��m�'�L#=�O�T<��ج	����0D�2#4�Bb�'�T�Gx�!�'��'|�dwݥ�	�H��D-9����S���I�#����0Հ+�O��q�d�/je�(��ȑ�]vDdY��O��J��'k�k�M�(q��I#�院3����'L������=�Ud�(���)ԁ�3��@�<�t�Z��"��QJ�`�D�Բ3��"|��6Nv���~�����"�� 'ܼS���<4��'ir�'�|-@��'��0�x8j�'��F>>0t��#����Ă��_��p>A�{y���T�@|��Ч��`��/��p>����ߟ0���|H�)*¡W��إP7��<: �'���Iğ��?�O놴+Q�6�r��h! ��'`���;]���s�,�tP��'�D��򄓮��lZ��H�Iu���#\\�AI��}�b�'fR�O�4ၑ�'�2�'r�ɚW�'1O��"`Di� ��|�բc۰*�>�<��nz�O�Ո#/'uz$]���R������d�;B�S�M��X�� �Yr�͗!;B䉃f�z<����-v䲜���S?m����j�IU������$�\�'���W���	��iH�4�?)�����;+��'��5�4�7ł?��!ʡl�3'���"��'R1O�3� ����rl�bMz�#iʥ�F��O?�D���(ٗ�A�E�\3�n�(?�t`�w��Ob�"~�I,f�� ��7�ܓ�ʍ)H��C��h��H"$o[}���MW�g�#<��)��KT/P3���d���Oٸ�Hɚ�?I��-��=��mՁ�?���?Y�'X���O����u�M�`��d�.��sA�.M���-�}B�^�7p)tM
�x�b� ��׹�~�E���>�Wn]d�����0O�v�h���L?q���՟$��I	c�6m�al�[BN��կ@B�<B�	�'�b���a�pg<�S�.T�����ᓾ`��Pp޴-�
��.?��tR嫘�4J�����?���y�H���?i�����O���?��l��䋇@<(R��ʏ8�N���ɳS*�d�~�	��ؠl���	��דn�a��3\O��D�O^�"�@rf�3&�4L�!@g"O�T�Ķ�|p�*[ X!���y�<K����[8hģ@���yB�.�ɕ{,��ߴ�?����IDu��à�V9	V�I��4{�Dx렡�Oz�d�On]�d��O�b��'����rgt���)��hGyZP�r��		�"1��`
T�
=��_�b�Q�f��O2�}�&�+WBN�WF۶j�|r +�h�<� P�*ؐ|0s��6{Ĭ�ŁKg�$�I<1��ѴV��dF�``���<��YK���'4�?�����O���Oެy��*
�����" `s`��4�@��>�|FxRDܙ�������b��2NPEJ!(R�)���ƃ� ,�!��ĩwؐ�E���bk<��	g�S��?� (0�(�+^���Be�%"X���"O�ع�$�9��%�_:CK�Bቢ�HO���8 �kf�X�d\�(��E�	��s���~�i��؟@�I��P�^w�w��h�ɒ=c�&m#�ӫDN�x�'���g/� U�ڙ��G,Oj,��f��n����FO�/��}��O̡�� ��i�p���v8��s%SJʼ,�D�?Q�h�8�ʟ@���K۟�ݴ3�����D�O��|jx}���3�DD�F�C,8�r4��[˒�BOM�`	� ��&�p4KB鉨ej���<yf@=Z��n�aJ���g��I��s�F�����O����O��أ��O���`>ũ@��O��D p7��ʃ�L�Xc*�sȢ4���:D[!��&�QB�x��"�nA<YSs ��:%��C��A�;D�z��N	�?)��/E|`�f�Qb�� ӣk�J�8x����?a.O ��6�)����;e�D�r�G܄b�B1�U�{��G{�LZ'��@i�� �h�8S♅�y� �>qI>� �����2$ޜbb^@��I�dy�B��T
��r�☶NdD�&�JxԼB�ɧzn���F�؆;zF�!�c�5N
�B�	�&%Р�C�si.}S�L���c��l)���mQ���MΑa8��g2 ��ZmF��/A�̅��+�ZT�&�˺_ Lp�휼Ts����J=����I�NT��)�U!$B�	�3o��i"F	�ZE��ͣ
B��4�^!cK��_9V��Fɉ�B74B��&J��+'b�d����d��-"��C䉛b'����'J�`Y2r
� d@0C�I)NRɨS���B���=M�C䉉d�D�1Ɓ͔<g�Y(aF�:b�C�5.O�l�3C�p���	G��bC�-�B�@�&�V�zФ�/C�I%@�RA@@L��� ȉ�Á74C�ɒ+��8J1N�ܡ���ʮ0�.C��/J^l�3��Tм)+���*o��C�	�ZJL��((��53���C�2H����½,�9Je�>K�C�I�T|�(��G%cؠl��J�7
|C䉟Wr��ĬG$u�n��o9;>C䉝'@r�A�bZ�9%D�@l�-�B�	>���t�M�+~`(`��4$�B䉙!�u�V!ێ.	��(`& �/�`C�IY����O�}�ȉr���	c�$C��5`S�=��	�^��a�I�GRC�əOк-	�`
e�FhP'�"O�(C�#qVT��g�2�)�pbL�(X����'��p ���_��h0oQQ8=a	�'�L� �h�Yo�ݡ'&��D��|"
�'ʬ��$HX����a
ψ:c1	�'t<@��0&�����ޯaG����'d�P�I��plƔ#V�\�p�pPLG	a���K��& ��f��P�: �� �*L�|܆牵T�* � �h~"��,?��,b�'��:��yI��y�-�{ӞԒ�G�b��
qAȧ��f��%J�Aɥ�0|��C�x���"���v�ޅ1B��<�5�F
I�Jh[oD�9#J0��Z�x�$�Q�@�g��ѪK�N� m�'���sʙ�@����qe�YJ��%�����eQ!�R�Y�Ɲ� Yj��$���f��B�AWX����0Q��yB�E_H��0����ϛ�$�8�έo�*L>D��Pi��]ib��残�:����Ц=����>����P�<�N�ІdZ�U���P�A�EO!��"OBy�́OZ��Ya�M(F]v};s*�J��'Uf]{���>�fi_�{�l4�� πa���2��Ch<	H�'��	q"�[<|c�}h��D1��X0-��0?��,�*�=Ga��r6�px�0A�*�?Ci��槀 ��	T��u�ؽ�U��
x�C"O�P�� l2ى�˙�p�pa�Ę�`�0��O���xB��/�֠�आ^hzա�'-�8BƊ�t� ��(�.\b.��	�'}��Ə�0o��2���;	��a	�'�Z�q�#)m���1��͌0�-��'�DK�ht���W�JV���'��xSņ�Z*�q���U�1rĭ��'r�1`q��."�Ek�̗ +Q����'n�s�N�!K<. y�n�)q�y9�'��\����VH���DԒ�j���'�VtXE%�3�L�Ģ��^��SL>�D���V�y҉��� S��@�B�������?�V���r�y�p(�I��uq3�k�0�ä'>$��J�
�%o�<��!*����>�,膜�r,!�)�"]8�m��;�4<Y�H�\B�I�8�D\�r� a\�R �W�� �Z�1!J �)�S�/"h 1�f�^��mP��_%kN@R1"OFt���hr7d	�Fl�0�d�N|��'�@5�"�<��5���b@��	�����uEC�(E>��ybQ� GRL	���s~��^���ؖ��{�S�O�t�+-P谼��ڻy����'#f�R�E�J���Q���w��@��y���:s	�a�
Óy���KU�0�r��(E�zφ����9� ��s�BA�0������{c��r���>a$��%�OR��ak|<�@�(.QX����'cR���g
��'����n� �J��  #��nR�D��,��jy�8!�+�}붠�`�1���ΫS2*�p����.�Z}B�#*��SW*+-O꼘5��$H*�١C�9X�>�q��|�<��a�&j�������S5�#V�V�X��ll�;:�ߴO�u�W"��<��<1Q��"�n�ϻ��2�kU�:�� ������I 	�`�ڤLL��L�w�L!i�!�dM	�x�L��!ö^�N��j¦)ϓiפE�P�ȹR�lA���R̓U���Aՠ=��Ac���>>F|Gx��ר/+�0P�#���6��� U�?��x3�x�@j��OdD��G�L�<A�1ϓhd&��BJܱx�DY�鉚&�E���<�g�Վe>��kV�I�`���U��#8�\�Z�k*?yկZ�g0,�ٷ��U������d\�k�j�<���B�,��yB�]-2� e���ƌt9�%�	XD�� �O�ʣ)�o�J�!���?YGkV�\Z��� ����Z�\st�١E�1�P�)��]R��"��]�nn�Q�@%�p:PiqqJI�<y.iK��Q�D�] ��7�����Y��KR-�50�PhsuBY����y����4��A��H��2��-^��O��IUi)3�T؇ѱ$��d��[��HE	�<0>T�vSd�xmA�B�.
T@0��[����C���6�0=I��V�*�XP��J&��*�cћtm��h���Eu.1�`ꍍ2���'U�-�q�Is/���O���U�� +��h���#F޹1�"O`q�ć��<@0EK�I [����
���`n6H��\}C�$p�M
�n@��u�2�HsHȳ	�B%@V��;9a|"�:ܐ�Uh�ML���Z�G�(��cJ�������`�t~�τ��,9��٢	پY�� %��'��`�t�C�'9 �h^�7��q!�� nd����@��{�����=?����U�:I wC�>4�Di7`P>*��a[���$2�D!�G�'�\��$���}t��Ǜ�*Ӯ���Ո���sHG!X��h�6�<��Ok��
R��4���E<	�5a܏�!��2�4���rgbP񇪚%:��+g��8U5��9��U,�;�w	 ��I�fpE�f�ŞC�8�s��]�/ԹD��A��=�����d�Rq�%�J�$�kH���[U�(�вO�]��O�q#,O�|�0��eO7yr.�����%7�8<B�NH�y�`�'h۾.r��xb.�As	�B�r�i@�Ţ/��X�#�:t���* "����=Q�h�+c�`�k��T��pb�$uF�6��0��H��*g�@D|�w��j�%ЮMc|t)��ڗ��ܪ�'��p�FG�D��0�&=\��5�����O��
��@<f��堃C�f`��L����6'ͫC}�pjdڣw�a|��C+P�1Q�I=3�-J�ʑV�I����>�p�OtѲVG�@t�����Y~�[��ɚX�D�4K��t;��H���">��"<Q���u1��a��iv����Eɟ�S>�čj'�� <^��!�ϣO����SÄ6�n�
�'a�A �ߵM�F`8uBB�"NLy��0D�\� b��$�+�����3?�缻��C!��!T ��p}�@m�O�<�  i{��y��2`cV�`�Zq����^r��C�f�ɬ���ŗ\}-�\�i��x��ǐo��Ѕ %�4��L��m9Ԭo��z�C��y*�+ �Sn�*Rg�G�����
ߙBR���$1f6+ `�i�t�޲$6�$p���ֹD.�ab�� �N�67�,I޴��1#�#� i��)	��/yPP�s�Q�X��C�ɽb���@i�1'���A�UM��)��JFq���.X�XTҰ�~�5aԁ�*���C5�ڥ?��H�������ٔ��U���ف����dL0}��T��(J;+�dy��g��ѓ�iy
d+���@���m>髒�A�6־�$� GΊ R�i�,y��A��-�I�5�`��xCN�|��j� O>y���6�)������?��d0�g��)���u�>+%���'��۔�<l���R1��<�t �I�xO
�{�"4��O�]��P&���)�:I�v(�C�,<�a���

bbC㉉k�$陵j�
h��r�ɁR�����B��#&��OP�*���i�đ��4M|H$J�g'v��%0�K�/C�l�
�������J��/1i�dA�����I7=��h�T-�,ߦ��Or�r�[v�	�X�8��)�}���c�
����+\�|( ��j��4B�+�"�S���Toj��s?$����Tk(��k��G 9!a!YGN�hV�|� "��*��Ȱi�0���P!�o�<!���=9�8�r딲C��̒T�.	��ї�n7Nҧ�����Wvb���7>#l���k��:�!�ʸq�x���'p�q��_���0Q�((;�/7�p=I���&��z�>j��!��My�P��@0�ڤ�t�i�Xdrd�z`]�и' ��ȓ#BN�X�J��K���iW.+k�"ExbeA�eϔ�����d�O��<�w�/�R�����O���h	�'�8��$�
�T)t�;J��A�ЇC�U�ҍ��]u��s���n�YĦћG�8$ԩ	�g D��s��q͚��G�.^�%9��h�8Ӥ��:��@��'�������t����d�];,8	�g�����hѩ
pdӂR�){f#2���~�VxBk�j�<��قƘ#Ȑ�C�BŃS��i��8���91�ߓE�<�3��i�U8���L��fOa13�=o8!�O?�:�h�"P56�˧+ Q�zA�����
�, Qk���0��Y��A��;K3��H�S�����>�\�<%D�F�G���5W�6�
�c�/waāy@	�)M1�QqcӉ`���������:�L�Xb�[�*��	�7er#<�S�N1�,x��/h���,�
���F��cA�DL21O��ƽF֖��L�	>�����MQ�'.������`�i`eـ-O���������L˗�� �$$��.�*��������0���|*D�ô�����x��)�:�ãJ���S��yb��#7X$��V�rD��BC�>��O�� ��0����#��X �F-y�B�	�&� �a�:K��DAK/-R˓[F�Ex��I�6g��))�H	�LS��w"�L�!�d��*�A:���N�����A�=�1O���V�'�$p,Y�l3x �ʙoM��@�'֎ةB��(�����μ^}���'�h�sT�z���g&ڼcj"I�' Xy
�̀�0��aW@O�V��Ar	�'¢�!� Q�P��HÆ��V�L�r�'���u3�MF�>-�|k�'�<9�����<'�H��oε2���Z�'�^���FB�P��3�&(�,�y	�'��q!G��7/&��Y�k8&���;	�'�>ٺ�V�w� ٺ�m�M(�a�'���s4�P=C@���IX��dZ�'Nȝ3p���;K�܀$�y_�1�'ct�;�nJ�ʬ�'*�!
dTc�'�ٹ׃]�`*�҇ɔ=����'�qbq&ӥ{���E#�w���#�'x�)ȐJ��t�x-�5�+q�� 9�'l��
�)�;�dIslʌr_��
�'����i˼,|RȻR/�*]�F�:
��� �1C#�� u�>)�����K�*�	�"O��t��.W�T�xq����I�U"O�9`�g�,:p�&�V�wʔ�"O��R	�>պE[Q�H�5�H�"O��)1jиI�Fp:Q�3hԜ�"O���R̈\�V�ӣe\	8B����"O��(ĭT�O6 �b��O�S=B!6"O���!&H�͐e�[ �1H�"O��bkG�[�����ҌA�<H�"Oj�8�����r��L`(ذ�W"OF��N�L�JÌ��Y%��3�"O�|Q�G=0��H�I�/m�Q"OztK![�TL,JTJF.<Ƭd�r"OP��V�'U�B]s�Iͩ
���A�"O���th��J�1q�Һo��<��"OX��۟~>\ض�;yp�eX�"Oh���<2�q���Y�%��T{d"O�u�E�ƽ19���0�W�z;����"O� 晋�P)P#�@3LI�q@�"O�5�@ᖴjo^�����v8P4�""O��6�ZDR��Z�%?�AI�"O��B�Ք-�����T  �qD"O8�X�C#��� �/I@��"O��b�������r`�լ
�R�"O" ��D;��8�CB�u� + "O,-C��vl�"�%L I0rI;d"O����f"@�Qp���#�PB"O,@1�k��&�k�䐍(�8�"O�c@ᆎ\oC��i��"O���L�����	=6晚�"O��ږ��:�ũF"Wb�!7"O|�ps��|Ff���
\�a�A"O�!%�{]�$��wg��"O��s�-B.�"���~��C�"O�����1,>%�B��s���s"O&A	���� �9SW�Ũ:��@I�"O�):@��9�|"��6�&��'"O�(��H�#*X�J2C���a��"Ot�;v��?Y��a�5d��B�f a�"O�з��ټ̳S"ĕ?��hr�"O��"�J�%?��;bƇz�4	�"O�`I"JH!P���q�4����"O��Z��\/l�� 8u�-J�����"O����D�Oa��ѭM:*Q�0"O�Qi@L�d��/Ձ��@ "O��B�ȣ~��Հ"/ҭt�|=P"O���c�ޠTZP3�͝V���9�"O�m�&�W�'� �Fm�5-�XܚR"O%�f�])c��p�l�9���"O4y���{}��T���u���"O� �N)K�X�&�(^����"O������?B� �R&[�u̕q�"Olp�s��h<:�8��ђQ�8	��"O��wEB<�Fm�$@ ��\��"OJ�I��ц="�msw��}�`\`r"O���%��%*=^ѢDI�;A<��"O��ǌ *wkh��T,���c"O��	r��!

���2ߊa���"O(d��!$(@�%e��7cL�)�"O�<B0AP"+�|��<4E��C0"OL���x�D�ч&�+#ڪU@f"O(�X�
�g���@4�^�RAx�"O:@�ũUWw�M;.� �v�2"O����d	
,!sM�s�|%��"O� �q�gK�S�:�He�V%�@�w"O
d��3�6hPĢރk�Z��g"OF�@7�3!f�ْ�A�6��A)"O��Wf��
��m�V���3wP���"O��P����1r2hB�s�b"O�ā�t}`��F�6b�h"O,���/��XY�2	�w�x�"O� 0cK�5}�h��Z��%I"O�QPD$�o3��FBS�KzlhW"Oޅ�P!	�M�|ƪ ���2"O���S G��Q�+W��)�d"OR�B�?,��I�J._ ��s"OA�ƫRG/V�zŌ�2�t���IK�$ �O9&� ��z�����#D�"��7?����ٓ
��@���!D�0��'�0�am�U�>��WM>D����M"Wq<���U�WQ(P`�k)D��{�ˇ�h�0�;�'YDj����%D�P�%B��?y|�b�ܨQtj�rƉ%D������y�ޜ3C)�;a��{��?D�������< ^$5�&rp�Aa�0D��c�EM��|�Q�I�)yj�-D��0��� � �W�F�%zbʔ�+O�<�ѫ0�ɍ&�[�ԧ����!¬B��� �`tg̳/���e�����'+�#=�P��3~�v�ҕ*� ������p�<�$�̂<�h���S3\Qq��_X�%�F��d�+xp K�kљ 	�*4�.I!򤖗+��Њ���jcHM��UU3!�$�9!�jiB7Ϙ;'y�%�G?q!��:\��$G�0s.�ش ��!�dO�=\HR��X�l��1bF悷*�!�
C}��k���-|�|(��8T!��/!���wG�D:!����h!�dxpIL�#(J-�ǂ99�!��<;ltyQ�D��,���E�e}!�d;^���. �9���x���Ky!��	�Fq�M�OS�N��ث!���!��� �1Q��8j�)z�JU1O����ʍ]�K"�@�Dj�8���%!��Cj���dO;T_(0Tk_ "�!��� M�����)�'q�@������!��;�����E>~�!%O�!�ρP"��#c��<6Bda���y!�$N	�LHw�_16uR6�\"m!�dM5�
�(ʠ\���pI�m!�$�H	�L�N��Y��X�"�Bp!��^fp�0様{�V�ɠ�q�!���
-7����]r�Xpȍ.u!�d�!ATA�!ɞ�f\��f)��+!�d�FDz@�'C�~h�h���4&�!�$?w?:�Qn�!j�tDi6U>f!�df�H�(�e� U�
�yT�gў�ᓄP��[p�?t���ª�5��C�	�@�2�v� �N��q���ˮB��'v�b8!e���X�#(�'J�C�	 A�4��cB����Ζ?v��IZ؟�� ��-g}�y���ݶL�R壡�;D��[��\�~��Tn��"���*O���ř$i�̰��)`�*�(�
O�7MM�#�$���I�MXEY�h݃th!�8�l�R)I�+��yC�!�D�r���W��`�h3�^m�!�3l�J�	����� �f�.�!�� |��c/OZ�Rh�c��	{,�z"OAx�c�4i��e�_y�Ԉ%"O^��ԥ��YT�M֡0jJ$�p"O���!b���1���,WX3�"O��@�*�S���Еi�+(��4C�"O,��G�&#����C�!|��C"O8�aE�S�7q�4�3��&VN!�"O
�)�2g7��+SL�u�x���"O���R@�e�l-+�לMȔ)�"O����R�d� X ��#�� ��"OJ�׉��YSzj����=��"O��Ql�#)�Шӏ��J���"O��d(�;���@
� �`�Z&"O���ǈ\�V���"oWO/z ���R8�(��Vy�X=y���H�8�JFE5D���2)4a��8�޶y*�)E�3D����N4��H�ǖ?�^=R�1D�|��$�z1k�@���)Z�##D�� P�W��ڱAT�H)n�5`�E?D���4耐'���JT��%+�N�3b=D��(�BZ��\aRɸ2
�P�!�D��'"�(1�#�����C�d�!�Ă�&Qd���T�)����ue�2
�!�$_0�J��ы9���J�v�!�DBx+*P��,~�yh%o��/�!�d�,a����]D��)�O�l�!��4xN�!S�2+�έ@��6�!��Ūo>�,���A�ui�u��Ǟy�!�F�OJ]C"'�m/�H��.J6�!�$�0$HbD81��A"8a�5N�"�!��_	{����!U	`1���U��h�!�E����Z�p���K�{!�� $J���K��� 4���4�!�$ӨxB�J��Cw�M�!��|�!� �d�(�a/ׅ!�>�[��	��!�߲ p����&�&+դL)���R�!�(��0��N)=��y�bO��!�d	Wx"ڶ.�wdF�z���!�U,����h�#G�@���h�!��$Os�e9��V�5)��Q"fӊ!�+���ӌɹ!�NT�GF�J!�$F(�@EQSN�8��3�ř5e�!��Y��s �/A�D`÷�юh�!�ғL�$@����4��e`R˄a!�d)Wؒ��"W�����!�d±]t��u�K�*�ҸĂ�!�!�Nmb$���%�4��A�_8'!��?"�$���B&z1��6L�!��M0�l����op��Q�,�!��+5�Ԝ:P��	E~.���"LD!�$E�.A�q�5EMR���@#!�J)P���%� �b�r�H!�@1(йz�GTW�b�1�%!�D� ~W��@/"B�T��!��!�DԊ�"W
534��'�2�!�$B3��a��O�Lِ�:�D�)p !�dIc͆�#���
��<ԃמP�!�d�C�0�Wr������[��'�&�j�C��8���*8�<	�'�z�$� ��,��fX�*�(�{�'�z|�*�6E߈� ���"-��8��'���+�m^����9G����6�'��%1B�T�#E�TʖA����R�'Jt��r'Y3��@���������� �`�����g�8gkILH�C"O��@	��z�09�	�K� ��"O��YEKO��y��gŅ�.���"O��%�&4���ၼ[w�k
�'Ț�i���"���'�J
.9����'Ofq�U��
8�X+'��pT��;�'*���s��@��炰4����B
m�<�����(缥(e��<.h��C�_�<��@6;Y� Eƀ^pT�tƖq�<����0ւ4���˿Af��E�ZH�<)R(6��M�"�C<B
�V�D�<�a'C?B�ɠ�̶4r�{&M@�<�m��Q��'Яw��Ip
Ny�<A�a�
l,���I.4�� �I�N�<�f)�rP���!	�9v̽�s��M�<1�J��D���'�ȣD���T�<y���W"��ʔ�\"gD��)�P�<���<�\`���*�J�[�/�H�<�I�2���:n��<����%
}�<1TP��J���(H=m��5�͆|�<)��WƱ!��;�6�1u�x�<ɡB�8R�,+�����֍Lj�<�d�I�4�W���k�V��G�Je�<�֯D�,�zP�LW	��I��@d�<��·6�5�����6��y↜�w=���s�ʈ:�t�J�.�&�yR挗A�p\�q��.ۺ��GbW��y��¼^��MBf�'�Py�&ӗ�y2������z���)�\*�#A��yr(��M�0R���	Ř4Z�����y�i�	�O4���Ehи�y""ԆV��cA"�8��(:5g:�y"#�.E<�q�B֚+XPi�� "�y�i��A��S��;n<�s��Q"�y�-B�8�P�6�Lf�,��!��y�g�q��qc�EH��;%���y2DP�#�l��c" 6<`�(�4�yrжv�z5�"�V+���H.�y��_k��ItB�� !@�qU�G��yb�W�w�^�i�E�Qz������yre���n�x<eֈ�5�y�K/@���BIC��(��.�y�LĬT[�
F�[�u�Z���g��y�!ۧC�xQDL+���J@�q��k���&�ȶ3��l�7�۱�RЄȓ{*�!���K�* 3@.���X	��7�\���ʘ9>��I(ƨ¨�����.�i����21+�h)b��$=z��ȓ'PPu�C�!�0��Z67�6P��OP̰�vK�=o���ʔ�;�4`�ȓ|.�!�Q��	
N�m�nA�E�ȓ�3u�S?D����iŜh�j��j��e��mʹ�QB$ːpA`0��iI�R��Rc@ sn��u���&A�V
31�C%�WW���8"Od�F��5䤜R�71p��"O�� SF �^��ĨO�A�0��"O����
�<��8��璑@�̉�"Opq�Fݩ_V�E���܊@�p�``"O�h���:yZ���Dd��]#�"On$sWi��(%�����"O��$�=8�� ��*ÛJ�4j�"O�W �9¤��8��E(���J!� �j�$Q�N�2~��LgM��,�!�� �y���گ	�R�3(�:䐤�"O8����^$9�Ԭ�P琪P*Z��"O����-�*(��� �9��%"O��pǊح.3��GOD1f$G"O��Q��R"����\�="����"O���撈=��99s%�&~Vѐt"O�Q5�E?�"<B��* ���"O���Aj���pgÍ/LH�(�"O�a2�2z�2`�hN}(ơ:"Op���йW#��c�ֿV�׃f�<	��1J��a�a��D�8�+%�
I�<�%�~�$Ty#ɓ�4�vds�!�A�<�3�P�,���q"�t.��!v@_u�<�"�3�T� `-��8��ܘF%M�<�!T9hX(v˝=HO�H�mWH�<�U�<g��@1
��	�Dip`�O�<�w�E�g����C�N�H�@�#�N�<	��m5�����H��mac�U�<���a�I�L̒Qg�N�<	S�۬e��s`o���)�H�<�u#@�<\:�B�iB�QFH�<�W)ֳ�z�C�(E-
��RA�<����o-�u��.��W�t)١��~�<��A�B�a2�j�lx�3��8D�����։MXޔ
�-�C3J8iR8D�x�ϕ8k�X!�f�[�'�ju�:D������{Y(L��e��4 U�f+#D�Ĉ�o=�����O� uh!#D�\�t�Q��X$��Z?Ǵ�y�4D��@���+6��E@�i�%�/D��z6H_7EE*=�ekVkr�ڕ�/D���%Ŏ_�FH�B�Pr6��w�-D��J��K�H<0��f�/g�&�4
!D�����W-*��]ɤ����:��>D�@sՌ��z�n$�Ћv�$�� (D���5@B'C�r( �@5;t�a�'D���Bn��1xn9�P����I�A%D�� Ú.!�ڠH����o��e��&D��JT��
�T5��aĢ6&�-��j$D���V�,'m������T�� �� D��@v�)2fr����5L�Y�`K+D�PY�)�N�l�9	^'��-Aa@%D�X{�&X�bYV�c�	^��E��#D��0�(Ϛ,����JR��S��"D�Щt�T�T*�0Rc�I=.�5�1�?D��y�+M'#���g[/#.�"��=D�@�4JR5u���
D�����` �=D���V&��u��a�#)%���")D� ٓ�2;v\Y����2�ĥ���2D���J0�}�rl�;�i{w�0D���@&��	�LШ67|�<J��0D���0�ŋ�\(r�#�%Vː��j;D��+��"�]��I�vTh�@��3D��3��HY ��&���N�Շ%D��9uL��IT��KR��PB|���&D��r�Ŝ|�~�F�_+$r7*O��i�kرq�ڐ�#�ۈl��y�"OB�`�ǦE\�2t�L�����s"O��&�U8.Q�XӔ픿4�*�P"O�L���M(k�����^�5s`5x5"ON�"bx��c��{f�!��"O�P�'��(N��Z�g�.cG�I�'"O���B��*_b�yiw�#b-FX��"OB	{�E�>��ȁ�є""��S�"O� ��Ɇd���Ш"lݢf��E�"O��*���!y��7�\!�ȣ�"Or�;D��#�C��)2��"O����H(�X���&	�2�
���"OZ���H3��LP�.BS�,��"O�Rրˮ$}0���[2^���Q4"OU1ulT�-o�!G� �h�h�"O�1/��g8�QA�O2��Y��"O�SGFQ�C$�m��ϒ�^�J��"O&���,��Q�Nʛ%�V��2"O�A��߾]4�$iG�{ h�B"Oh�B�dP�_-�)r�kA�U	�"O�-ڤ�]�X�|ɄK�k�*QP�"O���Tn����Ц��d�dт�"O8� ��U�7���@�
I�(�0ʑ��O���$�"�@!ړ)��e��L8���>%!�$��:����*| �u����;B��'ў�>I�qa��3x�ā�a�X��9���<D��+�!�u��� (�g)���*O8�0�ŋ<�P�B�J�/��i�F"O��!�Ő�N$���/.��HqU"O���Ř8E@��
 ���It�\�x�f�(�҉�cQs ~���,D��R�CמM��(�o�koVh���Oh�=E��+��S�Ҩ�'OL�Q2iF� �!�D*g&��p��EN�4"Ԡ�Y�!��'f8j�c��4��uHd �nq!�$�|����%@s0���^!��ۿb����a���CW�<����!�D��(�r �C� r��Ǥ<!���*`��A$i�Yo�eB��ʘ?5ў��aBxY@��8��h"Qd�
Hm�B�ɭ9k%����B2�PR%R�FB䉈NP��l*4e�T���%D�C�;�>��ꛡ5���Y��#9�B�-jlLٗ���DO��ۣ�(����hOQ>)��hSnI+D��o{����?D�T�BQ�s$,᪓	�Y� �w��O8㟴G��'��ɻ�%��p�ӴЃ��M1M>A��?�	�$Ezza�q�ڀ�7�-h�-�ȓBX�}���1��E�b�  �Ʃ��|+z�:ڰI["��F�j�V����rďd��[ j�@fX�	{��?)���ΏeVL(Q��&H����� �[!���-qHF �<%eV<�@�W��2��?�g}�d�k�P�R�E�1
@�`�@�TyB�'��D���F�h�4M��I�1f��'���53H��m�ãދeh���'�V�Spf� ��3�b��%��'�:�`ӌL�|���3��O	��'��ɓ#y漡����J<����'�������;�.݂��A������?���L��+���Y��������a i�#�%�D�O0��6O\���K��.��a�G�Ǭ �)@e"O���W)
%�x���$+��T��"O�rp�6�5R"���[�"Ot(���� ��]�A��'D�@��'~r�'Dɧ��8���-��#�d驑H��O����$4D��㵆�6B�T�ZF-�=�a R�0ړ�0|B6�B'� HQ��	}���w��\�<I1��)<��i��C6����	X�<Dh�:�z����.�n�H���m�<�B���"&Z8�vb�-}��rAM�h�<�.�\6�����Z���պ� cy��)�g�? >l������@%kҨ�@�͢�"O"x�'T�<��H���@<z�F�2�"O�1��lɭI��uq�m	(Pk1��"OĴ���X�!��b�*Ưbat�a"O8 q!����`JH�elQ�"OB��s�	rx��
�3oc��T"OQ@�O:,Gx�J�D/�����|��)�-a�Ĉ�΀FN�|ae	�-bj�=Y�' �<P���WJ��!wٮ����m���Нk�h� _o�1��+���K��B"J\�;6.�Q%�E�ȓ<�!c��S�
2�9#�,��[��4�ȓ� ؛���[n����N�=�B�ȓr�m�u�ѤS�P����
�<ړ�0<	C�4���� uI��e�q�<�m{�R c¬��k�
��7�Im�<�SFƿI�r�Z��M�
�Z���j�<aG�ڸi|ap�l��O���ϐ@�<I�(oz���
A/h�T 3 #T��ᝢEA� �C��9H�(��b8D����9g�8��T��;�զ6��K��<�b+XI��c����a[�o4D���qO��U��*�K�V:�3`2D���F�]=P0bQ Q�:�!��<D�l���
8x�i1��		7f�xt�?D�Db�h�s��aӌ֥g�:!�Ҥ=D��!wA��\��D�pkF@�ai:D�8ct@<?� es��/	�<|²O=��0|b�JݬD�
e�� n���pk�t�<ɒ�k��9(4��30#�����x���<���r �QW
N�"��gs�<a'�̝,H�܈��YZ� Q�2��U�<��N�
6�h ���Ƃ��E�q��P�<�p�J_G~m��IA�X@��)�u�<!V.Z�V�d�C�S�@e�X�7��t�<���@�ho)�g�Wd��Z�˄r�<�&�-W���B,��`��
���T�IK���$??)S��PPp	��޿)h6�w�@Q�<��D߬�v�@��pӸ)��DKF�<u�ː]��R�̍78*(��"�D�<�eoج�F�re#
�!��9S���|�<� �^�6�SFe2���Щ�@�<)��T�fT�7ˮ2�%I��c�<��NY�x�hT5Sp$˖�_���$��I2�|�œ3%����ʎ�B䉧	�ĩ'��1.��Sed��r1B�I�Hb.�hV@�1RCX�dd�r̚C�#�|��jC��J��Ο�9j>B�	�U���Nچg$�J�]8x,HC䉒kF��c/P�5y�8moG �C�	�F2��sI�?c���@��)�B��d���K��<E�XMӶG�C�����z"'�"g'XE	��N�Gq�B��!a" ����i�ꔳLf߂B�ɓ1�p�Ehґ9�hBȊ������<�'��!�i[��)�-T�p��\���n��҅Ȗ@�*�XP$ͷԥ�ȓք��g^�r���FY�<-��i�|�"�<[��Z4
�.O�Շȓpk��I_*
y�J��֍q�ȓG"p ��.T�x�eY}T-�ȓ�� v��oR�G���}P��I؟�͓P��ثT���S	 d��b�<b�H,��_cԨ�ŦS�?Nd��F��[ǈ�'���IT�S�g�? \ ���``%Z��K$,HE���'B�t
�g��D��Y�j��.���&)%D�x:tƃ<5D��Q� ^�b���#D�|csN�h��)`(ۚzŪA�.D�h�3͈"C�$�z�@XyJ��(/&D�d	WF\�0&�D00)��R"�`�):D� �AᄭG8�
�<w@��q�3��'�Sܧ"��� !*�4)�1�r�Ɂf*�EF��
�fĉ��C7�M�* � C�Ʌ,�}Q�#��z��Ц�*B>�B�	K;
��댍5�N���iΎ��B�	�d#��&뇔�6�1�+�(hB�	$R�rds�"�#K�4$jc]�q�츄�%0!a�Nr�9U(��3]lUD�'[>����iG�� �p]�=X��!ړ�0|r��"%���@уԂYְL�%L
T�<I�ǻ7�вE�ݼd�੺v
Z�<eo^�"��th���#?8z�1SJ�j�<�W�H�.�xܨG�Z�j&xD�5�p�<��%MĐ�0�6Sw���ŭWk�<w���g�Liӊ�&��!�S�<)��	*3�	A��_�X�"��N�<Y%T�|�F��!	��=z,�p�H�<��ڦG�r�Pc�ܴ{�xr� z�<����Kk����ʶj(� aUs�<a���
|]�A�28;jѱtʊn�<�I�:�\�s"���'/���,Vc�<y�훊I�ֵ��W**�,	A�G�u�<�Bv�¤�c�-��	PI�n�<�2L��|b��T�Q. =�xr�l�<i@ݰjYJ)� �+p-`-bi�j�<�bꀟmر��¤P��"�e�<��A]l )�@I�"�c�j�]�<Q�f=e�@!:�ےs�&�a�fq�<�H��[^�(r��ߑ/R���Oo�<	%�O2/�Ҍ��F�7/��T)*MT�<aGo<T��P��Z=f	��P�<Q�GH�?�N�����w��X7�w�<��"
�"��C��>6D����W�<�O
,x����H5��d�\�<%)Ǟ�p�['K�m�,�{'�WW�<�c�LKD~���g�[SN@N�IE���u��S�ҕ#Ѡ'av%��%D���g�pg��L�8{1BI��5D�X��װ���AfN��	��(D��pUO��`Q4�T*���XA`&D���tΒ4�l4$o=r� #��#D�[%�ǶJx����*J<� �a<D�DɄ���J-I�%��\l�f��<I�JZz��O@�B�M��B^�49��tD�3�X�wgT���K�4dŅȓ:6��"��v+ɂr�F�Qv��ȓY����F�d����1�Y�p�-�ȓ1����� �/�4P�R'�2��ȓ75����ݜz;��a�@Y�|�@��ȓi�PY@�,��^�9��+j�nh�ȓ�5K��,$��QA��3Lg�A�ȓy*��!Ǫ�oM��
%��/TYD���e�dZ��Ǚ#ˆ���¬-��ȓ.��<b��E)Q�pb�P�C9j���q�>�#����j�A�� N����ȓwNxE�0�_�������� �☆ȓ(Az�a�B�e�>���D�"V�1�ȓT�&�p%f
�N�hr���@.Y��S�? ��k��`�́pc��.l��g"O��!U)�a!������b"O&]2�'�.��E�!���a�+g"On�C1,�:b#��B�$K|��b"O�Y����-�B�����N����"O�,��ȳD�|x��O��s}��Z�"O��2$ϓ[	�AC�M# z��[�"O�Y�T���&���ȋVx�A35"O�D���cՐ�1֣�S�b�"O:�A�
�(��1,�= ��"Oteq���\��hw�	(#����"O��2B���q����끐2���se"O��c������L��P�T"OJ�J��Ÿ�|��o�%�΁1�"O�Qs��:�p�P#�RsꮡX"O��r蒒5O�T𗠛�����"O�YQˀ'|o�A�/@]�p��s"O���0��-zo:�yG��%�(�C"O05�v/�24��Ё׌G/#n�5"OݙӉD%M�4���@01�j�z "Od�� E
�1�.l����[��V"O�y@艈-��m���4�$���"O֔����A�(�k��=3�z��"O����_�����d]�Zg��7"OBH��ۥ5D��Hb#*N�\{�"OjX�Xh@�`������*L��F!��6Z�,��3`��r
RdK[9&��)�'|����v�M�.k��C�WFd1�'X��@G+�*
�2����N��Uj�'y�xq��@ 8��RFL�@�a�'x���@mYA���QM�:�H�'5dP��K^+����͇�@0R���'��I�O'`�`�ǌ�^���'�yB �E�z= \�ϸ ��hs�' ���&��)pB�	��[#r�ȹ)�'��A��BO#
��y����u�T@
�'"LA`�D�j�p+�^j�<��'�#NX�V�. ���9A@�'��H�C�y�
xq�h�	(ܜ8
�'��d�#H˕M͢��OV r�H
�'����2D��;,Tj!f,��OE��y���7���ԍ�9��l�Q����yB�\1+ �+T��dq���A�yb�ہT���9r����ҵ�N:�y�dX#� '#�\��k��y��;sN(��r�
��U�B��yr�A�[l^	��(܎`�&��%�Q5���hOq��l�C 5h��6��8�d�R�"O�E�uǈ��8�S�/��)�#"O����;��2�AƌJ��)�"O$�a��Jrɞ��s�[��i�"O��h�	�Wp�k7��q���B�"Oډ8��Ĕh�J���E�{�ZH:�"O>��Q��E��� ��ܭ8�
l��"O��¢�Ⱦm���X���Z�2��A"OV�l��S��'k�1��n!�$ֻ{*���&�;RF�(� I��!�$	�5)t��R��!F�<�g��9G�!�dF�ncn��t$�f�𰴏ǯ{�!�$�I�r��hE;{2	9��2s��5O!/t��CT�Yr����J�&	!�d�6z�,��e�]�[��A.H=Pb!�'�>d��k�=��t��#[�$!��*.ې��Bƭ�L(B�L�J!�� �p2���T'���$��lP��8P"O�#�=Vd`�kGD��5H�d80"O�a�1ND��b&-�l4�'�	�3�6ȓ"Z�1�Y���ç��B�ɜzP���U��k��6UXVB�I�VG�Y���N�v-��0+��
*.B�I��.Q��JG�V����%-�=GnB�	�/��Ղ ���� �1�ZB�	�~����C/�p�c��Ku�|B䉠~�|y�"EU>nx�E蓊�5�pB䉺�������3D�bE!��Ϝ!+8B�	�aL2�C�̈́JH�Ypȃ4P*B��|�򡸒�U*<8fd�f�B�ɂUIl�Pp�S=>k @�Scˬ��C��60��j�'ݿUK��a4 K��C䉨Vٰ�O�F���p�ܩ{��C�I<;(j r��9f.�sQ�3|C�I�S�T�J�����D��C�a�vC�I?4�vh����/�lLѕ�(E'8C�I
&�HA;`���A�}�����aJ2D�$��G˃3��C#�#,b����,D����@�0|�R-�5Ĝ�8��	��)D�,h��,)AV��v.Y9j��]���%D���m��:��;DH��>��q�vo0D��r�a %o�~ȉv�_4����.D�X�����Q��o�r��A��+D��(�ၫ�"�j� ٠]1 ���&D��%_�	�0m�@'V2���A&D���b��|0h6�	�2�6m�q�(D�Dф�2�X9�KF���P�.&D�Ha�fI.6����D$k��D wO9D�@Ҵ�@}4>4��)�cļ��4D����gL,I���`����vT��3D�X	F� �~�p�E
�I��4D�$��UND��`�fP��<D� K�/J�o���P�]�T�<�a:D������4!*����$�-	zT`F7D�8P��8���ՉKQ`zAS`�2D��� \�#���qSkJ�{�v1�51D���w��rd}x��
�E �+��$D���E�">��p9�DJ /-�B�.B�ɡxԦ@�A�Q�g���z�T�>nB��$	���@���8t nl-�#fuC�V�~l����G�<<��$�S�C�I�T���3	i�\�˒�ς) �B�I�NY(b�]9�HTA�M�?�bC䉾L�jaS�HPS..<�q�U�74�D�O���d�&��s����3�)�'|e!�Ě�F���hc͍�2�0=sg�8&V!����`��Н+�x��eRM9��U���ɧ�Ϥk+
�Xg��,�����%D�0Q��F7 ����/S>�n�8� .D�$3U�Q%0y�pRP瑃e׊���-D��A��N�*)L�y�C�aE��z'@�<�
�S��c��V6p5�����q��ȓ4x6rB��=�����֫(8��ȓNm�W*�Yr��)pR���ȓ�^4 S�p�|� ��#D��a����Dـ�P}�:����X�~��ȓ���u��0/	�ۢ��_X<�ȓ��)B��U�o�ʀ#���k>D��ȓ'�<H��)�@�n'A;<ńȓ��)�D	��X�P�RUɝ!{l
Ն�2EH�U�L��2QG@ZH���S�? �e����La�!"#K�+4�!!V"Oܡ�eM�*T���*H !�m��"OR�ň�/F���ҨB ���"O^<0��4$�dCF�H�c��e�b"Od̘W�ѣ/D@Hc��qg�pȅ"O�4c�,T�]�$�*����cc\��P"O�1��NY~ $�"��J��@�"Oȑ�0H�dv�\��Oͥ9U��"O��;���u��K.N�(	��"OT	?/ļ��RFޭS^Q�""Op=���.Ԅ�Ce� CoZ� �"O:���HU�)�D�iJ����"O؝���ٶI������?V�u"OT�BHȴ$�L<#C��=hZ��{�"O��#(ϧW,@2��Ͱ>�B8C�"OZ�Q��^2<d�@ �K���"O��j�ix呷OE��Tp"�"O\ �r&F��f��,C-Z�fAv"O�M���( `�\�ԩ��1z(�*b"O.��p���p�!FƐ/>޴��"O {"�K�D�V"�/R�&���"O�c��i�r���Kȕe{nQHt"O䠩6��=yS5X� ��r	Ȅ"O>d�ׯ��+jj�j�N��uN #��D.LO,�9&��1 ?<�!�Ne�� ��y���-��x%�¶_z�({"�Ա�yD�>\���j�SA���9�+���=y�y�Yu(1�G���N����v���'�azB�H�{�vX�U�6?o�L�1�S"�y�!�-�|�#%�6����D ��y�֫��%�5���R���hO��D)�*���8 �¡F�S:p!���*k��5J@A�.���j[*ug!����޵�iNᬑ �	�e�{��'^���<ZF��f+�3lt����!�!_��D.�D�a"K����Q؂-KP�j��>D��p3:^8B-ZٔT�@q�cM:D��BPԈ6�kRFՉn\��X�@7��a���Isk�JM���v���~�� �3!1D�X"$υ��b�Lќ�f��-D���Q�R
j���V,Ta�<qKĮ*D�4�u�֕Y�B�S��4r5.�j�l-D��)R �jD̻���h�J��(D��x��ӜothY2J�4o� Q�e�+D��I�#Y0%>x�E�=wn2=���O�B���A��xH�,B!����4/'�C�I�R
�CS�V�/STI�҅+_�C�I�~�1��MP�����&͆C����+% ت/��8�)ɻ#ZC�ɿ/r��AGoŏHe�	Q&͓})�C�		7X�,�v"��V��9Ko��f��C�4]�z�ˢ�
��x�i�B�2q�'Oa~B$R�h���qh�=`d%WG.�y2�N�?,<�Y�lS����,�y^�P-��n�v>�������?9���0?��[�CB_i��xZ�ƃ;H[!��A�	'M�я�I���3�ܬI�!�ۋB�Qav��9��B�Uj��'^�a��@!Ԧ��E׉$o�����'�ў�E|RgD0��0a߹0=	�)R �yb*Tx�#�.�� ��9��	���y��5\���'A�}�HH ӡZ��y��N�W��(��_�s�ܕ���i�!�$E� V8�0��M��|؅F���!�� D���n�-Z�����
it�B�',�O�Y�0ǈ�X�`,�5fB�)R�'o�'��3�i>U��F���ܘ���:x��Tj�<)Eg�pnh&bK�y��(aDdh<ɲ���}JD�a؜9�����%�+�?��'#��d�ǩD�h��ϓ�t�*���'@�-!Ч
fs,M3a}b���
�'��Z���8K\=Xë��vШ�{��?��'�0��i$6���j��*q���1�'�����qM��ӗ�F�t��@�'o�E!p���1���&��>t��z�'�����_�~eXȃF�4n��d��'�:�Yf'		����UA׷e#n��'o�����J�N��eM�/k7�hX�'n 0�'!�_V(dCGa��QNj�c�'�M��Z�
�iSf��E\$��'�<C�,]�l��J3��{��'��x����8<��'D�y�ZD��'�(�xB�\���*��lm�]��'V��HӃ�&����@�/�>��'��IB�M�������� S-��'���� o^�."�y�D�ͺ�0��'��1µE[4^�^���;l����'r�z�P�v4`Q�AO�2bYX�'3z�p5nA<��)�a�+#.�]��'O��D�x%t#�lQ�  �	�'�!"�'�^�t�n�"���Z�'$V��@F̣+?���w���8��	�'1�T��_�"uN�s� ��%$X�'�8��ˑSn�ͣ�X�1Fn���'�`��H�����ɑ�0��eS�'�����z�,4yā^'�zH��'���Y�J�!h>^�2��B>)�0z�'��{uON/Zd4��N&qĥx�'G��p��-/�a��#�J���'�8p���Q�D���cE,�Ll&m��'�<�0jـW�í_p�X�
�'��؀fkM�%@P�p4�G�|:�̘	�'��QHӣB>~ ���Ưn�q�	�'L�5�"ˮ[�.Ш'O;[S�)	�'N���O1N~���6o��P���'�:�R��!��D��K�{E�T8�'4� byN4	����e���q�'R�	��h΂)�����E¼���'���؄�Q�G��s@�Z�_�f�
M>9(OV����y( �ᰏ��>���(�jшs�!�DE8(Oz���1�x	*3鄳.�!�d�1G����
��Bz����6!�D�  Qb�5&��[_�M �FŒ^!�dC"Fy�EG[�HH��i��	M�!�d� N ����3ILA��I]/?J!�$�41��lڦI�-P��Y����+:r�'���'"�'���@�!%ֱ�� �
7�Y��'6�RrJ�+WD�i�d�xv8��'�zH� J���N���X�r�Y0�'�v�[U�ѯp����h� }P�'�"��a�F+�6K�K�Yun��'�j1��n�%�i3����L�����'�q`��(z�P��ԘM�XM>i���0=Qaݹ0��	ڴ�X�b3��
�m�d�<9�O.?�`��S̅ ������W�<	S/\*H�z��̇/z-����S�<��'I/<F� Aċ�����O�<����"�Us�j�
n�=rŋO�<� \८U/v*pPcg�F�4�!"O�D��hCa��s��:p�`��Y�P��ɀ0A��5^�Ti�oN�`$�B�I�|�1�B�O5�$i��Ϳ�B�ɨ}de�E��+n蜨���'L�B�<!��ə�!b��X'
�K�nB�	J3��y!�S����R���C]:B�	�к (4��,Rی8�͵FOB�əd�X1+�Ʌ��$��+���Ir<�@a�-V�z�p�MDx�X�# d�<QAƌ�v�.��KK>�}S!��h�<s.Z6&��ƍk�
(�3˔[�<	��[�L
�$��(K��z� �T�<I3�0}_>� Dbْ1�,j$cA[�<�Vj2?�tk��ގcx��� �m��^���O��d��ضR��UX �Whn�y��'�!��C�K���A�B�`�����%ƛ#^!��	/a� �!���pK<���AR!�d8R����W3:$%f�W'C!�$�8�TLJC��`Q���AO� !��F�ޝ����\*}��ڦM
!��#��x1P��q�V$Ӕ��:f��'�ў�>]AdNL5S��\�����`APQ�?D��F#�O�,4a&�Ã}�~y��#D�� u�T�@�`a��B�����h!D�̺��.Ξ"eΞ�%TB��;D�\�MD�Z
d����;�B��"I7D�谁�#���3�8q�`�!j(D����cEsW�0�pKT�s�p�V�3��^�'h��'o~�㗆@-�h§Fk�l�s�"Oxh!�o��5�i�`g�I��y��"O�m��)�8#3��hUf�
�$ �!"OJ�с��&3�^ ����HY:9�"O��;��t}aY��<�dG"O~�IP+HtO�QG΋�u�h�8�"Oz����8[���3�DpNi%�r�	���O��1�lCs*L �釴y��a��'��`�4dWe����rN�j�L���d7O�eZ'K�'�.�b��,���B"Or�Ї(�.�X��v�0zJ�m�S"O&�ɰ���r:Ѹ��͋D88xH""O�)��ˊuc���v �4�Z��WOI6EЯ@�j��ׄ]<qI����*��0|J�"���x��ҏ!��ĉT�Nf�<�A�޸H%�l�4��9�!p�K`�<qGF�,2v�w�"	f �$X�<aUȚs��Bu�Q!H�R�3�m�R�<���-�N���,�R�<�2m� <X��L	+���'�K�<�0A��k�[�l�$]Z�WHG�<� BS)�n��p������Dͦ�y��̍B�Ș
tn d)�����2�y�GQ�wD��$$s�T�+�
���yR	!�Ƶӵ ݙc0�y��-I/�y�a<
��Ux��ڻ_���iΆ�yr�
CQ�A�g�Ԕ\�(�`R���yba�
-���ֵ
1\�s����>��O4�h!��X�����g��T!�"OD�ggX�l�R����9�<R�"O�l��/�!Y���d퀞N��}	c"O��x�B��,��8H�Ru�
M��"O�i�D�ժ~�B|8v��?�R-[G"O�\���+ �܊���)\��!aq"O�P�a�ȲE=���Fn��c��pa"O� �I�d�S U��M��U�����"O�Ѥ���p9Z��ƍƙ@�J��""O�1�åީu���Vj�����c"O^���/T�R�d�T�E(0rd�Aq"O��8�+Y�QEx�RB��!e����"O���`Q:U�h�1!/�1iH6�J"O0U��������#�[1B3�*�"O��	�B߀?fE�o��"Ơ�"OL�����:��ճգL�Y�m�V"OV �R�����%��%}�4�{�"O�(z����nY"�2*���Q"O�dJGHф��:ĆQ*�Y�"O�=ʆ@MGrNui5%�<� "ON�HԠ�	s�����H�/Je� "O���Ua�7@��9i��ș��`;"O�@�UMR�r �<��.Ҥ\9�"O ���S0���r�N�"[�G"O�1ۗhS�C� �����Z؂��'����cĂ�\v��e!�'Y�L�'���U ݍ.�����S! |@U��'��P���!j�����ʠ}��`�'�X��Q���Sb� �iw�\(��'T.`���"T,��FDѲt����'��}B���C�r��J�x{(mJ�'FE��X/+�m��J[�s��	�
�'+��"b�	}jDJ2c)ZψL�@"O���ǭ��|�e�2@�J��"O�̙"-�s���P6�ӊ@�����"O�8�w!W=Z� |��,۪�H5�"O�X�#7����2&�=����w"OE���]�`x5�@
�Z���@�"Ozh[ь�:-�J�m�:� �f"O(�B�.vxi�snZ��jp��"Oj��PE' �����-b��d"O:聖M��|���$l�$+�T���"OX	ʄ�G+R��Ԩe<@��JU"O�t�Q恀��?�p�k��]X!�ޑF���O*,@�Q�b��W!��v"3a)��A�Eb߂V�!򄘭[I�X�+��,��-ˣ�� �!�Q���Ѐ��V��	�*ӗ(�!�D�=>z�B�	��Z�L�[��>�!�d
�Hdԥ�2BǽY��eb��Y�O�!�D�'W�`(σ(r$�Ȥe�"�!�D*)#�*��V�P�9�eNz!�V* ���w��=��H�Dn-q!�$Q�o��-��Fq�)�^�wm!��N�9��(y`|6��*s`!�˾Ur�(��b*�"Ė�O�!�d�2iL8(�E��J�rQ˅�N(Z�!��0����`�,m���5��d-!�Lq�X��1�P	h�k*ԃ�!�$�<K�zp'�"�����.�!�ʹMx���K�rt��(�$��!�$�m���SjA2otl<9�A�P�!�$M�P� �bϩ@g|�i���
s�!�)I��\����`(\!Ɖο+�!򤌳U]rf�?J������P"w�!�䅘2�����|�Bg
r!��U�9f�j	B����Ʀm!�$ɪDWؙ�BRsȤ
�`C\�!�ۙ̰
���R��Po�	|�!��S�,��v�TL��eba� p�!�T+c��t��jp?�ЃW� �!�� T1��ַ��+0��1@��yh@"O����\�nR��Hv�ܳd�b��"OA��-^� �.�;C@���"O�����_'A��E��C�NyL�A"O�m�F �>I� E�ua�qi��"Or=�I̊IL⩀��C�/Y@ՠ&"Ob��WA=s�>4 "�L&*�ʤ"OL����y/���g䙕U�%٥"OlX�J��|ܦ��"DK�H�Nź�"O���;�T�𶂒wH&�b�"O��Ћ�OF����B���"O�E�֤�!%�R!q`�Ǽ\���i�"OQ�$�-9?��u�3�z�s"O������[prͨ�D�T���y�F�-
���J-(��Q�V��yB[7T�TS�]�%_���jM�y�	TV�t�c�^�4P�x�����y�,�)϶yx�m�7/a�s�E ��y���,W��"P	�&Ƹ30$�,�y	ֆjˆ�� ��*5Εzr)�&�y���_��P�ԯ��9ٰ��'�y�ɗ=7""���JΔ��!@0G�y�$V ���'��C�=��̓�y�̀Cq!���P?�Ӷi\��y�k�r^�PF�T�: �8BV፡�y��/#b�h��X"*y�u�Ł�yR"�6%�|�a .\'KO�q4l��yb@[�M:}�pN��,�R����yb��nFn
 �Z�/��c�"U�ybE�2;���w"�;|�m2bU/�y�+GG=du�Q��5KU*q)q�T��y���n�Q�_-��l��yRf_��PQqA���p��d/@=�y������h7����0x�bnِ�y�U)	v�i���� ;�0AR�۱�y/Df倘HwoH.m�&��qcG��y�Cļ2�(����
Q'�h9��ӳ�yh�'W��b�؎yb���ቆ��yR�
L��Aa��t��9I @C!�y�k��F�y��Ǖ�>Ƅ��N��y�.�V%�i*��Y�g����W��y��D�e�n�f�_A��1�g̙�y��\�vrjX{!��a���C�)�y2 �+W=x����t��K�ʍ2�y�؂;�x9Ҥ.� ��g���y��$^V��� �J(b��u���yb�K#!͎�`�E*q���ek?�yRخ~���F�f�~�	&�M��y�dK�EP�b��4H�����cO�y��޻/ ����@��>��\�o�)�y��Ԓs�y5O��2�\������yRmX�:�ڈ����%-�����y��ɾi>�-Iƣʢ(� Y/��y���j�jR��%^�<c�K׭�yR(��n�"6 E���{a���y@�չ���C��:A&B�y2�Q?0�6�77vi2!"��y�����za�_ }�D3SB���y�HJ*(��WnW�l�,:b��y�@΄��8���f1����$�y"��A��i:SB@)ޒXx��S��yn�0q*���C�� Q(����y��}�6���c��������y�HK%�"���X�|�Z��F`ΰ�y
� |(Z�(MM|���N�v��\sF"O4�R��w4�T��
�U�0�c"O�+��=]:J�"�ƞ?fn-��"Ox�Yp!�!0�xRƆ��V��"O��Յ��"��sC�d�N�("O��#��!�9�HO�R��=y6"O���5��r��Hᒩ3�H@Y%"O^�i���d\� ��Ŗ(N}�-KG"O�,�E�\�*���;V͛ʔyk"O�-ҁ��(�&܁�gED�༚	�'���j���t����cJ�UCn��	�'���Q����0�R憩^ �y�'k�&�(K2Ĺ�M)@Up}z�'���F����2��$��>$V��	�'��\�q�
� łѸ)ϼ��@k	�'��DE�Ʉ�9G�͒��N�<��%͞�(t�="U��AdCE�<�Ϭ^�L�� � W��(�u�<�p��l�lp@�J25����G�u�<$NK�}���yBB�*q?(UbǮ�e�<�pVS��0�f&|!&�f'�{�<�%_+�r�1�%K�!��cV{�<!,R%+[f��Ġ�}�b��s&Pr�<	R*�13��t���>XI��DF�<A�fӮ������}��"��_�<1Q�P[(�!6�
��� �V�<!���6�x�ZL����DG�<Q5(�;�n,� 'U�=E���qeKB�<ӭ�v�ĽRwa\�<e� Q�ˀ}�<y�#@�j�閆
�`�*��BD�n�<��膑M2V���׭%-6r���+j��E-q4��Z�A�2o�*Ɇȓ\�0b���V-ȱ&.{Д��7�Q:$φb��}����=���� P@b"A�l8
�(�K#f�fP�ȓt��mib┰
�^I� S�r(��&(�Ѡcd<E�<��� �܆ȓ+����#I.Z�*c�	�u�a�ȓh8�`t�ŤH~4����f���\�\`R�#J��AV�X]�L�����H¶��J�Dx��P- f�ȓrL�B+;'���IP�h
���ȓ�<aCg�u���s&ʝ;8l@���J���p�gަ-�e���;@���ȓ HBiJO�-�XD���!��ȓ �Q �?YD��dQ�z�Jx��FH�X"c����a� �v�ȓxȨ��vI\44��Y֍�>;*<�ȓ]�$� �1:���@R�x�8p�ȓv�N�i�-Yt��Qiش^����ȓ{ hxBC
9Sj���w	��T�e�ȓlr�1����Z�؄�WI pL�I�ȓZۊ��G�P�ڈ�7d�!@q���j1h�J��,)ذ�ł�hm�ȓ ��Vj{WP(bD��M�@�����T�e��36�y�$WK����ȓ@�
S�x<�С����@�ȓf�d��u	�-}ԜQDg��@6>q�ȓv�@m��&X7	�,{�	�.�N-�ȓd�uHV)S�@�cVHs�e��e[08S��T�x��%�1	�u�ԡ�ȓ>,rk�![Tjl� �$7�L%�ȓYdm��p
(T*a䇟M"���J�v����j��QH~t���S�? ��B���6Z�4���=&r(�AW"O�B���k���ɘG$��q"OF�{�&��}kR��qd�4;��y�S"OН![	{�� Q�_�8���+R"OȈ��*Y&��%cS�c\�Z�"O��r�1�9�V��?�N�8"O0��E�8c��AwF�{ϸ$[G"O2�C���p'���p�X4�� �'����[3U���\4n��T��t��'h2A�(a�N��S'����'�ƭcf�91��$�sj��F���'�f9�Vd۸:vj]i�IR�JYV�9�	i���'����_�7 �1a�۝ 6l-��%��i0W�*��2����ow25��;��`��E��/4��� �A~�>��ē���4�<����q�ժJ�p�$�eH<@E�k�|�LF�b�4���K�<�+ \(�����?V���cd�D�<�R��)b�h�i<�pԋW�x�<��A��g����b�L@�x�t��q��D�?�����pq����4I����$G����k�0�p��s	k炇:e0��<���?�S���1�KP�G�Va��ـ"�C�I/˨t �h`� $A
1r�B�IKH���%�2�,2��'e�����)�I�o�� a@�=X����z索=1ÓMlP�z���yP���/��E�<a���0�WM��&V̠r��ؽu"O�D��4��� -��	l��F"O����d�+_���* lO�N^t�b"OrI�dc)p� ��&!ǶeơI��	]�Od��j�h��Mᆜ���\�9���'�d�+A��z90M:�	Ğ-E��s�'n�P�����x�9�Ј�K>���	]�]4��"	
#0Q4F_![��'a|Rō/	�ΠQb- �Zu�yz���O8�=�O�����ȚMz�i��	�8/�13�'����
�VT���gB�%�����=D��	��K+VX��T$^�1�h[E;D�4�"$\>&_D%c��� s�B�,�|���I��J!}�2a���(X��zǄ(D�x��I���Z� ѣ68���a��Ɛx2%^=b�Dl�"�[84K�xR'���y�n�.%N(l��k\�b�u�#^:�y �3*����V��Y�`:6j���yҨ5����g�N��q;u`Y��y�D(i�乢eۺGg@�D���y2�!b<�!���0Fd�17NG���x�j�=O�b��V�Ƃ[���s#���$�!�$U9+�s��N��8Q#bJ�"�!�	�_�<T�!h��x��IKG���!�$K�:�~ap��W+&����B␰s���x��d�gD�6�J�ǅ�R9H���
>D��P���$p|HC'C;aB֥3֭1D�����V^؀�� )���v�/D� ���>�6�C�mY(r�r�a�gL�<����S�`��# �!{�P@SѤ��o	��$�>ьy��	��I�Щ�K�2_q�l*S37�T�'�p��D	��с��G>l���c!���?��O��GV1&�x�fZ�2~`�#�^'�$�IP����C��	��̀%�C$a��]��,ړ��۸Oc4�K@�ϥ,1�) n^���tR
�'��kq�ϗba�!2��̇"�,8q��M��X���'-���S09n�kC���z��5�өXj���hO�OH0�S�? Խ��J�7�2�(3��
�"�#�"O��c/ݚK[���Т#�>AS����t���O�X����14�~š�h�?p����'*�����Q�3�p��(�4�VX�.O��'r��O�����/@�2m��%�x`�U `�9D���U���	��V>#n`u�Uyӆ��?Ɉ����'M�0�A���T� 5�#È��0<���$!���H�遈 �ƀ[�DO�K21O|���I�T�P$%߸yT*�]�v���hO�O8��3nJ���n�*\,�L(����D0B�	53�R��'A+p�4���Lܹ�ؓO����2�8	f��<W:��j�,�:}���:O�H����uY�0�3mŬB����<�S��y�/!"�{�%I(U� ��O "~��Cϊ��%2���P��}�<�GOr�<�6 �Y\�ہ'L}y��)�璇�٨)H��dm��n��Y�w�<D�̣��(65����qú�R�K����O$ҧ�i0�I�^B�[�ȫK���F����C�	����f�����"s�2'�DԨ'ͷ>�!F~<a�kU)�VM��ρ�@��ȓp��EQ2_�^�P�CP�+Pj)�'��~��Fc����MB gL,�+�	���%?����hO�i��͠��S� $����*�!���O�T�Gl� �E�i�U���p"O`�
�g�wN@��m�[V )0�'2ў؁v�ʌ5�h@z�Y�N���'D�t�!kY�:ψ�0�n�n서D	$�� h�$l�ɕ˒=\��)Q ��i�|B�I�0Dpu`��H�Mʨk'��,��ʓ�0?�Vܪ,��m��CUA,��c��Z�<q���K��K�>����k�U~b.��O>��b�vjt %�`�Ed�*D��HB$	���p,��<.�<�&<D� b��-��`��Ł�j�Ӧ9��hO�Χ�L���CI��5'�R�LA��`5D��2�g!WJ^�"g&�o�Aja'�<a�J(����&�d�R@��� 7ĜH�ȓb𘧭Uz�T�X�&��:��!�ȓp�6m1 ���H�,�qoƲn/*q��K�,��wM@*� �Hc��5Af-��N��j�˖�j�~\�椖;.��a����s����&>N�b(Dc\�|����E-D�����H�B�(!�1o�s��`a�m�Ї�I>	��A�ЁN�,�P�kǥJ%�dC�	�y��с֭��<�@d0��g2|C��?L��h�3�T�Y�����[�"<����?�Sbj����`��0
�<%�7h'D��С!{��,Z���m�$u)��#D��V�R?@܌�PG�HY�p%�#D����a�w�&�he�M�s�ФSF�=��hO��.*{�"������`UؑN=D�,���A�.Έ�Y�,�) :y�ǆ�HO��?yI�T����$�N�N\5��c���':��xy�L��<� ��k[��$�+����y�D57�FMBgR�	L�᫶i�4�y��)�3��@�n��/@��0���
�e�ȓY��n��o��ec� ��(�' ў�|�aY�/]
аnT�[�85 ��_e�<9G�g����ʕu��<���{�IH�̪3��6��}�GB ?u�Y6��<���0g� �gR�`\"�`�.Y�D��C�<O��I�R�$,�v8Q#��6?�ʓO.b��Gy2��2x�Yp��������X��?鞧�  uȷ#2мA�!�5ek���"O�4fKϹE��E��O�A�><C�'�Q�,��b?+Ŕŀr�^�wZ=ɅK8D�$���%3�2���I��K#�#D�le�*`n�IS��'WZP8�# D���t��3g!�y[��L�S�D � �<D�Avd� J��+��P�[b9D�x�!b�3��h�JN�j"��Ap�3D�8a¬V�B�((;F�J.Z�"ݠ2�-D����U_�А vM	u���!*)D���V!�+.�șV L)����!D�P�cM�N�u�I�)�>D��S��^<C{�-`Fk�<]@�!b D� :�)[� �|з#�-Q'tI�)+D���%^WᱤM1(R -'D��C��8��T,��*�\]�$%D�����v6 T��ܑ"1�Y3�(D�0	a�"p틣?W�fA��,"D�$�&��	SI�t,@�qR!D����ȏ-��u�D�ņY�J����=D�T�����(���Dȅ�UO���1D�Xr�S�t������v�� �s�0D�$C��7F�)
�H|����(D��"b���� �U).��ȉB*2D����̕YyL"�(T�r�B(4D��zA���u/��4��[��l"20D� H�N�v����"I��b,�y�L-D�����$��z&��{a�mɖ,D���,�'x��"��8"b��k(D��b2���lv5P���1�J�à�)D�\cA��v�.EA��5;Fjx"`�%D��9b#�"z@h Q���.��#�0D�d�b'��7�q��Ρ�4U�t�,D��	��^�	�H%��H24��r�$D��b`��P���#��UKF�I@.D��C����D�"$D2#��A��6D��鑻�hC�*�U Pa#u�޹W!�D�,7d�Bg��s�,q	CG�w!�D^59Y"LA!90�P��"��6�!�L7�H�x
-9� ��N"�!�$H%{Ϣ���J��F�y$�RT!�˭4u���˷Z��TQ��n?�\��B%	��I���]-E��#f���A���t���7ǝ�<n�݀�&)D���'�ݫ9a�7	ض�<8@�L;D�(�IX�iK<��EY�&����4�*D���E-&����K�LQ�w�*D�i$���\S�-bn�M<�e(D���4h��[H� �qf^(�&1@��-D��sFo��&805�B?�4%*g/(D�p�Bƀ�K
��E!�
��X���2D�l#�l�>�%՝3H���.T�Da(�
6�X)�c6}.���"O���H:U�@;�ĭ}�����"O� Z3�۬w�R$�V�"��"OnXQ���Lt���
_% .�b�"O T��@�^������n�)�"OVT� ���@|Qê	{K���"O����B���t
�;U�A��"O�T@�D�cB|PR��" �䈊�"Oʙ�1(O-$�@I�k��o��IY�"O�)7+��N�d(���N���s"O>e� 
�')�t�x /\�:��&"O��g#Q�q(�Mb1oЍ����g"OYJ7ψ�&�b�Q2��>
F��"O� T�WiA)����G� *�0�"O�@��7;nIr��D�(.ZI�4"O���nМB������T�Ab���"OLdCҮ�ϐ��1Ý
~ió"O���D�޶���Qc�f��{��'�r�@��x���-Q�h��m�t`k�KX�y �z���A�B�Y�@�BK-��'�J�zb��my��#b�&?�	q��8�V�!��f�L���")D�Hr�9JTIb�"'�&,P�I�"��	
�-IwA�K�>!h�Ox)'�G�& ����lH�J���"O����NJ�.Z��c0�M,]�� �I=^�(��'o.t��ǉ;I��F}��&}���z4;\�<y�!H��<i苹Y� 0�v�<�;�L�[�|��Q�lw��B��U��`@���.�OHT�7m�;;´�y�b�I���x�`�Y�|�0�O2����ڙ$�ŊL?�FŊ�u*I)���*]�s�%D�`�1��NXX"V�)4�����֖���P0�P��$L��s���$!ks�����M��Q�q�"	�`P*l�B�;$�P��I_�K�������\R��K�c�����Z�tX% (��]�'�	fV`k&dA��Z�jg� 'K�l��$�r�P-O� ��`>{H|��f<�u�� P�Q5����@��p?鰉�8�pQ*�큸~f��S6�CW�I�s���\����K�(n��#C�~ʦ��`׍J����CĂN�<�4�ɼH������8�X�ಣ�]��$]t���Ň5��O1���'4�i���:'�DɤL��
Q����'x^�K&l�0�v)��b�)8ؽ���D
����~&�$�&h���(��Z��(��lk�C�:e,�s�� G.bb m��9t�C�Im%�k�oL�-�n�����((]�C��&�4����ڑWؒ��力�|��C�	�5�@�i`m�B ��WŘB~nC��7 ��E)���7�&���5I�|C�ɠ1�l�j[4��u�1O
>B�	](�E�	Y܄c�bN3I":�Oތs�"γɰ<��R�q�Hp��W*��	�%~؟��g��$&U�-�A
(��	p� F��Q3E�r(<�!��56�'	�#��i���L�'��m`���bt�t�|
"� �p��N=*x�0k�L�<Q��[�e�dD��h�~p�q��c?���'&p(eK��+}��i̭@(ֈj�cQ1ws  ��jǪ-����D��(��	>nq���*�.4���8Wh�w�
�'j���.�q��D�Ď ���L�@@Є�Z�=�D�`���@���?�P�h�@]�`���9��Ȍ9�6��b��) V�I3ٌ��ѣ��c@ny �;O)�ab�G�YzQ���Ѣq:�	�!rX��P$71�*�#X0(]��L��g��A@����Ǚ�[������AsG<G����)`|���� .�\���D�~"�
�X9�v��0�H0\�v�ra��Z�2��]9�MD22�����gi�a[�1�1O����\�gG4	�c�M�B	�t�>a2FG�4���:��:ړk��l+#�Ҡd*��c�O�[`|<����^ -
&�ؘ2P�Ģ%�'O���P�1�f5�	A"h*��dj�'9z���M6��*5x�'Z�Xi���S9��7��}���[��6Cږh(V�?���
�kvnc?E��C�64���
2T=~aې �>���Э~S���a+�� ��ЀAÛ��)Տ^�2, �O�4���H3e��	{�(�5K�l��'�0�n	�E��;��ٗ����d��d�\dH�;Q~�}���M�a!F�	�D���+��GY�Mr7�X>{@|��_10��?	i]�a��������M�al�"/�h4Bd�^([� ��@�H49��#�!C��ҕIQ�	q�H��n�0�|"��)Qq^����غ>� �H����8-��b���R�c�k��vJ���r�,G=N]�A&��m�N�Q�$ɧ_�B\���G'9�ڤ��ҽ^M�l�Չ�$~��}���a��1��H�#�Ќ�G Ѣ$��Y2�o_(���`"�L�x5*��%c��-���N�!�мɧ�P �y���I��F70D��Ş,C�Z��I�7\jy���π6H�;u+M�.�bV�ɓ)��p��ذU��p�"�@�g՘��N�3B�U��,�,*��Ȑ/�&�N� �2�Xg(ƗA�t����I"��O �$✢U���F·'������ �X���T�U�K����aKM�/�jp�%�P-IN���O����L��,$\�����D�%/��ѳ%�GM�����J�$��I��!7��,��<{@��$qD�t�P�p�*�����3 ��t�c�G#U�Ҹ�ŏG
D�����8ql*EhL�Y��x� ;T�� ���ua|0;�_CҮuX���>�ԁ���l�"~3e�fa�:G���+��\�Z��C��j±ϻB}D�E��'0��ܙ&�횴Gz�� =%���"�Ǆ�p�謊Em�.'��jSk�2l�XsW��)_�>�B)�"2����6p�����m/%�뎍�Ϻջ��@��� uo���ϡ�"�B��vӸ$K�����Z�&��x�� BЌB��M+��K3^�>�a mB�EȐi�����@�R��%�C��*py�l�7,�;��,\�2�YP�	�:7p�B<g���5��!p�O�%[�)k�������y��2t}ℒ6�J?\��BGF�g��1�Ā
�]��[7[eT�Z����f@�Ǔo�x���O�����#�e����SN\��,�+��:.Ha Q�K�n�&XS���mZ)'�qa�w�Y���=^8�m�� #�0	J��3qϢ����ԪU��!рT*%(\eȕ�o�@�z���X�.�y�
�6�����ah��)��3L�* �%�.X�`�۝ �Z�"~�挋61�V8XӢ�	�(c�aB̲p+Ê6'���P.�3�0=���Ł#��&�^�#�J��px��F�߃&�Z�Ag�3Y�P�UC	/p�� �K >[3�=SS[�<iсK*�����nS�E�:�(�[��7B�ZhR��d�B�j�O��}C�+ԍM����$��Us
�'-p�`��_LO���g��
o���$��e��m�t$-�?��
����	
V1���n�����m�/ro8C�I�I��kd��i�]�5˘'\r�d�޸@�T���_��}��I�!^iK2l
M�`)�q�GK�T��$N�t��-G�I�^�	���+�Ce�
��Dh�eB�#�(B�I�&G���R�"JJ��p jk�OH���ޡimyR$�=�H�0����6(�$5��l��� �"O�)$%�;�ԁ�R��,�hٺ���@P��I(*|������g�\P6�b�E�����{��_�F����/D�����IT�e䴙��Ù�t`�yE�ԕ)�%Hf)i:������@<.tb$T"83r��@)Χ�ў֜�C; hZT�#921�������e�4�W2qT�\a�"O�C�1 T
�˖7O���'m�0Q�@çe�|AQ�T�"~zc�Ӊ ���B�dُb�X�I����y!Z����Cc�ϰe&��T����D�<Ɏ����ѯ����Ă���m��׆�D#�eH�@��'�T;���#���`L63|8B���%E���*��^��EbCacX���f�D6d|h'�ϝF���05C��V�͂C鉜5*��4gO ]{V��|�SB�$Epl#")'g{�0��\�'q(R ��Q�'QوX*򈕸'J�֥�32���	� �H�+����h[2�����,� ub�_6�}{�������G�>����3_l�"}�G�?��yK �_��,���i�ny�mA�|�l��"��P�ax�ɂ�d猸��LLh��s �N,��'�� ˗ <�pvj��4a3y�`la��,�0*'��1�`��.&�Od�Ά6:�ͻT�S�	�V�)�	�/,�D�q��d�x��y��>���Z��P�5�<!���
�K�4!��?qsI4���l�rl��$�>�h2�� ��"O�,�Ŋw�B�#Bf���,�
�"O��P�Z���!�%/͞H6( �"O|��I���$W'.8|p�"O��pr�R�U.��E��h�l-��O�@��}�$���*���G
OV݌Cቺ@t���2���w��e ]B�@��ċ)q%��2�O�	n�?5���P�N�!YV�哥��]�D��
t���r�'�����1	��yz�l	z갢O�4�TnX��剞��S�D �u���^�?���,Z��t�1'��� �����C?D�ؠ��<�Su�nȔ�+��)l��	�f�Nظ2��Q�1��s��s�ĝi�mz>�˅��LzD��AY�Xͨa��;����ğ
#��HɦaBQ�LY�P�=��HB

�h.�u-Tg?�UD���ϻZ)�t���'��l�c	H�m���iwkŘo��a��D�<���|�)§�4���`�#N�X�p���O�=x��?��%��.l�h�C�%�	���/[�BL�ɍ7=�Lx�Q0S�n�h|��S�~���o�,k,��&�H;��V�^*>�SO�Kb!�$ʖI��l &
PE �j��e�I1P��4:`Hf�JH��J�K@26��Z?qV_>�$c.���[r-\�UPBAh>�O���PD�>E�h�ɒ�ˇq�j��E�U>F"jq���Ԕ/_�THǫ*^���r���O*x:@D��`)�X9��B9�*�cS�X(-@b �1X��A�G�sx��j�K�'j֊ �6�'�~�����e��y��)� P0�O
,Z��S�� to�ѣ�i$�U�@�ʹy^Q�O�O��SC-,v�B�Q�V4�Ǡߟ�Zq����yr�VE��"�#H�<�eCŉ���U�KzE���[+O�\�qkHJ�S��!�(a�~�%n��X�`x�o���>�f�_g�$�#u��u6���i[�y>l�H��B�I�T���B��(V�]�E�Z�!��#=Y���(Qєx�/��9�z�9Đ�W^��3'��X�C�	8/�Fd����z$���ʭ��7�ԉ_�ԯ�%��)�禥���u� ��f��:1�db�4D�:�\4���rHT�
��I��>�q�@�\M�`�/<O�#�C,4���7��D���G�'����\0cO�!@rN_�twFm)����]�0"O`���,��t��@u+އL�F���I^ݞ����qأvf07��I��w�<B�I(B�x��S�P�"B�}��f�Q�@B�x\^,&i��&��A�Q�x��B�	(B$�l�)��mS��T8���m�>��rh�|[Tx;5��;:�`�ȓ����C�e�.4�
:t���ȓ(����S9:�����)G����v��a����f^-�D��).2h��
�H-�RA�4�@��&@?�L���=�
���1P�.YA�n�M�����V�J!SK�Z�صc�q�J@�ȓ7/���L�U���u�����{��Y3d��+�r�`cO	5	i�ȓwc$��b���6����aK�~p�ȓy���� �Kzp��)M�Vd��<�xSK�"0
��V�B�/d��ȓQG.����;D�]�&h�܄�ȓh"J3�N4(�� �e�)�!#�'�PcDܕ6�i��� �4���p�'�B��3OXX䎉 eE7"~6E+�'k�l�B�0m|��mU,�Z�#
�'���07`E5X�Х�čtu>I
�'<&M�4텨�x��e��vr<�`	�'Y8%�c�O	\Ѫ��N�':pf�x	�'������5]��:�&]�34 ��'g4���䄌i�{F+` 
�'v4t�WE�L�҂�A�ƾ��	�'=��"�)��J|��(�����yj	�'c��jAb�a�]z��TT����'����e�>Nف�H�=lhţ�' ��j�JAR)f��*�����'N�T�"kML9�+h]����	�'��I� .�(���3�-Ā���z	�'��Y�ȓ�nQ���X�|�t�B�'��`�؞^A6���. }x5R�'�VM�PeǏ\Glm�#Z��YB�'���:�-�'� 2�J�Ķ���'Xf�a!�1涑SA*��Q~�)K�'tj�K�f˳m�^QJ�
L0�X�
�'A�A���s�"��w嗯R��2
�'RD$�	�&s��sT΁��H���'��!�e���I�A��(�����'�>9�a�X�H����bkˁ!�`!��'	��	��|:��s��m�̈p�'.usb��/�v����m:)��'���釮�+�fE�Q��h!�'�,@�� `R�|�e@��A�T�x�' J +�H� ,VJ(��BgBT��'�:�� ߧU���끋H	4��'�Ԕi@"�	B7(�S�gú1��Q�'�~��Mڇm~xu怹sc�E*��� �\�fdM�Ya�L;d��3J�L�'"O@Q����[�L)����Q"Z)0"O����[�~	>E����F<sE"OZ0�%���Kh\iZt|�"!�S"O`���0:g�Ч�A�"��R"O.�r�m�:g��zt�K1��,�!"Oڙ�W��;���)���	a�S"O��3c��Wl���$T�	�,�P�"O,�+�B��_�vY����*l�:�"O���#
�)M~|�`�
=\�%2"O���%nct)H��ߚ@�V){��'���B��_�	4
��a��֝J�ށq�B��|�C�	%9�JL�,��V �x�g���L�'�D,��oLw ɧ�O��A�-�FIP�Z.6hL���'q*�p#���R#�(���@�J�d�V&�R��D�5g��.
!GzuHc��b!��4d�65�e�V�.%Є�'"�y�P���/ҁZd��
�"�d���Jsm�m�F_�  � ���Q��.B�2��a(eS	�Z����Q>����q�xq��Ӱym@)��������'�МҩV�
%\%�O>���$?�$���w[��tJ3D���Q�+As~<tkW�E­���K;'�_��;���U�gܓZt����-�(M�@���$_#�B���Xr������=� �^9Z���!ZH�bA��j����BL�fzH �@� �y����..O\8�#��!�œL�����9pSJA��rqk,D����xh�� �^7Y���d�/}�=l��Q��|��d�Y�K��!: ��	 @4i�E��y�d8h,��G�h���iA�/MqO�<��@_W�g��� s�ٷ4�1`����dB�I�.�a��E�,�-�'��YwzB�ɒO�(�������Q�T�c<!�	B��ĉ��$$����/%�!�đ�`�"�*4h�X ��ڭM�!���$1�����Vm���ŋ !��-�<�rڌ%�J��!!@�R�!��؎V�R	UIMzu>���",��'t:���bMlX�xA���E���B�D�Tݙ��9�O�<�Ҏ �0�X9�˞��-���ŤN�rU+S�%��a��@������7fR����$���H�T�i��c>%��g��74��O� ݰPA"D�\��
#�FPQ�ɚCg1 �����T��/E�S�>E�4n�"]���ׄG�. i��[ �y��ع{J@�H��C�4�ʁHq�����Jn@�cQ���{�ax2aғ6�貤� .	��A"���p?Qw�\�O@�h0��6R�Vi��`�٘�!�$�P/C�I�� �vi��	H<ܠB�w�l�>iq!��k�>�Є#��JM�RjQ�1��#%��P*B�B�xiaL�5�R��o�
?����a����7�I�}q�S�O�Tx0�K�y����/a�����'���G߼v�I��'�C� 
I�� I��`0�'�\j�.Ҍ^��ãdE?�$��D,5l�b
�{��x�A0ǬȽ
�&8�
O:��� ζv� <2/CItyb�ɂ9��Y��	��<��Pwګl����ä��%qO��qr�]�0<�BE�(@�R�g�;�b� �+�D<�bł�hǌ���6s�!@����=蜠&L���?�BFѵ`��T�'V<}Jp�
��H�'ֆ-j"M�[��!�Q�?Uɢ�}>����[/Yql�Ң��վ)l����o�`͡ejgU� ���d$>7��󴉎?�y@�,��^�I&8�DD2�r,���s���f�0�U�P�<2���a(9U��q���Z�4��X��x�s%�9�O҅ d��<����F�־z�
�VÝ	A�n���K����h��@�5ϟP�hi�dk_�H�i��wκ �\3/��ӎALƶT�	��˴%xP�ƌ_
����(�]´�L��`ĘE��=p��Y�b��'H��z�G�Z ��3GϹ?i� �V]:�� J͸��(V�a�c���������2E_�h�F��X�Z��R��É�/ �
U�S��*�>`�s�>4��r�H$; D��"o�$?=��#c	�,�HO���Ǝ�>uLƅ����I�Nx*�^�89wF�6\2�B!�]�}���93�*�ђ	�N��ы%\�
�@M�c��u�8E/?h�x\���J;��K�wo����	� D2w�z�l�7���#x�DR�R#���g�׺6SL ��A�H8�s5��z<r��6)Q �����Xr~�p�gE&�jB��6(U
�'m\�7��$�V%Ŝu�t3!w�ލ:cJ�k_F�i���4Bx�1�-ݩ2��4��O��P�C��(��uO֤HF�@�����p<��I���փ���~��R	0u�M�@���P�M"� s�[5�t)q��V꼤���3r�QGzb ���(�Qc��zFr@b7���'GvPJg$��%��A�ݑ`"`�D�e�������`O$	Z����:�
؅�	�"��=QR���J̬��bY�w��h9�.<}�iD�E�:�"�ݹ$O�9�F���F(K��SѼ�`�]�O�z�{��Lz���H�<��)K�v< �$�����r@ 2<���+gCAN��ϓ(5G��O�Q�d���PLBsʊ|uX1�#O�h�1W3ctHA�ӌ&����� ��~I	S���$�PB�/LO��bS��7{z����B*)����'yr��$��(-�=�c��4�N��B�0#��Uj�
�B�	*"O�L�!�c&aK#i�7�B��#�|� 2�Z�SE�Iv<Fᓯ3��1�^�S�V�A�?9�B�I!S5`�[���*C^:���*]��)R��F� ������OF��E�:�3}��Y��(���RPJ�J@�G���x�A�*�LE�%M�7�|�A�`����OU�Z�xMC�
�5azRk�:�P��!BO�6�������<���BJ�"���I��c�B�î٬rMDDba��S������"�y�dB(j�6��I��eʩsń����e��K�dIK"��fJ#ҧ	�4��A�8d���Џ�`�&E��j���H!��vԈx��T�k���,��yR�Hͩ֫�@���?d�R���ݪS�ӓp�a~ҩI9B��5K݁%��A�� �͘��� B��H�/���0?�J޳e>��!�?M�0LXT�^�'y�����Yl|\Q���Pznb���@,4���ؕ`!�dW�@��tZ%�(ԘP���� ��ͦQ����⍈��)�'qt����2SX�0��*?n��1�'��(�&�ٖOC��0�l]"O��H*O:�C��s�$u�c)O�R0bD9����$J(+�,�7�'�&����/�����;a�,8Z3B՜md~LX�F��y!��ġ+�СZ��"������ў�
�K!r�\2��l�'0��eʥb9��zq�^3��(��6�<b�d���2�ˏ%E���I#dFnP-&�p)���<E��hVaN�K#�~i����l�!�C������ARe0U�]��IiUA�!� t8`���ɗU�h<�gօP:�t��F�1=r����
<�����	_	ȴ�̚�2Xn`B���4t���'��L�e�$j�1k�J+)�����I]dT�Q�&;��9?$��"6K��
�X,��J�C�I�_��$�W��	$f���+I�׀C�I�y�h)�D@��� 4��c�I�bC�	8 >BD�f��]������0JNRC�I�I&R,�g�ĭQ�	+�i��nC�ɕ<�z�Rp�E�8p�'��I�HC�I�N@��J�#�L rU�<v&�B�L�z�k[!vC^��j 
hbC��#�(1�r#N�?�<4�sa�/x�*�I�s����'�~p��=1�M3�>y�x-(�^b��{�����?��LK�,�����b�{B�c�<qG�\�O{^|i���a��P`f�D���4��n8B��"}�$�,��0���*u�`ph�O�<��
�胭J�t1BA�
��M���� �<���h���؜tP(d�@�5�l� �
B����
d�Q>%Z��]
H��(J�DQ�ߊ\0��Oڱ�t���rE!�ۓ0��xpԢQ.�1���uQ���J92��B_�)�3��1-��B�~�VA�G@��i��Y��=FQ�)W"O�T�� ��\��G�\^N�ӕY��$ҹ}8&��2��J� ���,}�Ť|� l��5�ڥV���dCt+��1�'�^xy�n/����ъM���7-ǰR�>���Q�����d�=�􉢾H���Y n��F�̂q�&�"���e��� �l�Z��s�) '
�4܊i��8�~5�Ί�7�r��k��Ļ#�s؞h���̔"Ҩ���!>!�8��t�6����۶s2�O���(1̀����DA&�� ��φ,p�=����5K�!�dP'
]05�����`J�>q��I3�M�HɁQ@����������,H*�y&l�!b)U�h�a}bd��A�8�(�Q5k� š�F��]��T�!".]�Ɠ} �£�=� e#�ʓ3cܖTDz���Lс�a^�'U^@�TF�����F�8�f���[2�-��ܿ)q��b��(+���nڹg[����%ϾUN�S��Md��"Y����'��u�b@:'��B�<1�&�7y��p�Z-h��!B�e}��P�d];�G�Hx�
F䒮=� )T��T<�9JF�*�O�1j
�bF,1�C��*4ph �dէp�����*D� zT�8��P�o�&-����n+�D��H	�4�'�:���"ZWn(��D�bў�ȓ`�AJ��C�VF��gL7u9t͇ȓA�"�bҘ�+u	2j5��ȓO�4m��Fū$6����4e��5��*?�
��D�<�[�I�ST=�����DC�DZ��T�\+:�����^���ǯ6��[1�Š_?�x��WbR`�`Kٶ%�ܩ����jP�ȓG�H�#T���>�������2��Єȓ���#�L���*u�d��ȓ1/$���l�}Cb(��W��H���M
��h��x���w#&S����-*@a���0iH�a�����c1��G�yJ�)�_�}{�f>t�`U�ȓ2~�HQ�ĩD���NUT�z��ȓ�j�SɁg�r$襎�'4�$H�ȓ�j�H��V .��u �4Q�ȓ#�ک�R�ۈ06@�����'�Y�ȓhx���G�ڶC ��LI�@�JH�ȓg���&� 
vp���%F��ȓR�Τ�"�e�D�	
*v�*������<XO\@H�J\5��Z/���.u��HԎ��t�v������&`P�1��5���»\_ `�ȓt��!cD�
f�B�y���2M�|�ȓ6�"��s�&>u��X�)��h"-��_V	�p�ޔ�珎�`v�ȓ{��xsJW%BH�HuBr��M��\�� �4�ɏ���#�C\!J�$��%q��YMx
i�d�ZX�Jهȓ+	���&��mf��ϝ�Ln@͆�� �5Ҡ���K�s�N�ȓm��DYua�$�T����#���G|B-�/�0�crd���-�DT�y���hOk��&,��%@�lC�I0y��i�KU$�,Y�hȤ!q�C�I<p���P#n"�b��ڒ*6�C�	�0��[@�����R�X�^�C�	���6oZ��x�r��<!W�C�	�{�h���$��6�Hݱ3C�C�I9u�[f_9��������0��6jf���\�c$�A��A��DYz=�'��+)O��z��i�=H�Q�e_��*U;&M Mk"�xƣԛ[�1�Q�i�&��IĦ���B;��@t �/Z��U��m].���I@�D ��Ek���С�+�"%�C���6AV�j�	�*b�����8
-`D�즥ZU��x���i�u�8 �!K<\e��7ʊ*9d�Q��æa����#�D]Y� �?=D��¸("D�CJW0.����4��6`�2bԼ1�v�,[)J��h�'����%`��B�T�2D�?( �h�k���"4h�CUh��m�p#}b�π \	HǤڛ%V��Ĕ�O�8Є�� tM��Q�A�JN��D�˃M9a�4ϐ5\�q�-��P�l}��߹�Y�Х�����'���31���?�Z��!����)(�6���°�� �̀�JE9�a,?E�d�ԝ_�����B�A�(-�1oN�HJ��5��()*���"~"]wĜY �oL�2�.x9��]I��Q�م��b����ē����0�0�I�U1Ad���n133b���U쌌�0|Rd�\&dJ�S1�P���-6-F	�O���M�
۸��O >�y@nZ�LX�I�OD }G����'�Q�ѤEd�1O�>E: 	�) ��BM�O��Ղg�&%�s %�)��5��7/�����$ �ܠIP1D���7N�z*f1�B��j.��8�&:D�xKw���MQQz��DBلT� �:D�X�r��?u�t�L�AI��7D��RpE�05���K��P�h�i1b(D����
ڜz�nغDB-Z22n&D�(�4��/��؉aOɛQ�PI�/D��b�gH�$�yaG�)D�:ŀ�0D��Q�̔/�X��d�9�l0Bҧ-D�(�蔁]�N�Ypǌ$0@�l	E� D� ��Jъz;~5�&G��=��*�=D�4 �G�/�<�1&ŔW(�y�b�;D�d贄&+���B���7*<�p��9D�l�Ī3D��5��I�]9.P��A9D�Z�-�1h��9A��n��j�,D�|H���-y��)tǐ
Y�x�*eJ(D�\��iK�t7|PyV��:Q��k1D�T�q�J7X�����Z9cCHu��+.D���o¸U��0@Ģՠji��2D���lP�o��h2R��L_
M �"$D�0����y���k���P��tRgN"D�d(d��!Z�Y�q@X&/��1W�>D�D�Bʋ&:�=����\z���U�=D�0S�'@�N� CFh�?5���*8D�<{�h�jZR��)7��]���3D�t��I�R�f�G*6�ݹ�M.D��sc���~�`�Y� �ziC�E,D���2)@'��	+�	�8$~6d+�6D��	0�͸?.����/�:]Z@�#��4D�@j4�Ǩiq�1��!�-�&X�I?D�P�u�3pv�Ӱ����e�0D�8�R�L�&���1J�i��2D�T���M�y����L4T��8gO<D��r �Ê=2(��k�v�֬K�j:D� ����4d92̻WD��/q�\�V�8D�����G�~�h���+��U�h7D���½2S�|Xf"�LA�ecel7D��[bnI�+'��h���,Z�؋6�3D���o	n"�ĺ7-�-cn�K��$D�@X�*�a�c��U�^��$D�p���O�h����u��}7B"D�d�K� Zrc�K��A�|��%!D� Ӥ��?��C��"Tܰⵁ?D��hc�Z+S,����)3����J>D�d��'[�4��A�&�(�^hy�J;D�4c��%���G �6[\ E�5�4D��Sҏ�
G�bĒB��7>��I+3D�(�C��ZD�����܅1֌�I��&D�  �̐l�L���Y�)<tӨ0D��
0iH�lPSGI�4*�h�m-D����HN;-jDd* �*.�i�Q@-D�416���R�b9c�T�o\4���,D�@i��(@@̺�m�(o�.�ѣ,D�Xt.A�S�P��T�5n[:]I�-D�4c�S�ۤ�;t'�Alx��4(-D�� ��U�s�R�P��S=<�±"O~D0���Y�@=SӨ�F	�,Q"O��&��?~�ApÇe�0m�"O�!7��?����N?M�H�"O��)�^4)���Պ��zD�dz"O<���-߹i���*�G�`12E��"Ox�S(b�D��FI+�l�f"O0ٹ7,��6�tI���'Ă19�"O����۠q��i�j��P�~|�"O&!C��E�<��x��4{Mz��u"O��A&'�>G�tX{�m
&�ԳS"OF܃�&S�}Q-T�@,X�"O�y�E\�B�)e�օd`^���"O���w�\�;]:�h�P6�X�"O�I	6S�
9Ria���":�[g"O�<;�'~И�(͕��:�"O�0�,�>y~|�0E�'�h�"O
 ���S3�8e_-��8�"O� #�ٿqYv�Zs�2+���{�"O��#�f�s�����W�`ʙ�"O���Wh^�K�8�8��0@Z�]V"Of��જ5A�.d��
ݻ2A4���"Ot����DP���I�?C�B���"Or�J��Ё��mr�i�KO|5��"O�AS�@�4$~��!i�<���Q�"O���2�F��$(*�(� �Zԩ�"O����M�J)\e��.[h�X�S�"Ot��eJK���Ed�>E�@@��"OJ�2�Ӻz������imZ ��"O0���̤B�i0�h�7Yh:�"O���u �$so�ar�C+'OV] �"OJ@�ā�3� ��Q�UM���"ObL@t��"/���i#o�/d6!@v"OB0���@�iT1Ĉ�l�0�3�"O�$R��q,:5*�IH�d���"O  �1IZ�a�9�E�ʌA�F���"O$��Ҥ/�N���,�#3����"O����"A��8C�,@):DHȉR"O��ґH���l5���G	=:�A҇"O�� "��m<i$C�'J1zD"O��1��ƾ��}�C��=KlT���"O��3gDQ4a�P�Pc��N[��1"O��x�/	�BB�I1MQ�RLdQ+F"Or�2�M	B�h��K���@�:u"O>Lx@�H]��`�K."8�!h "O��80�N+_��y�ȞL�H�xf"O��8���)
�`W'_)mʶ�"O���"�͗�,���'�HɲU��"O��K'j��\FPyA'��Ag"��R"OB���*/��y`���rQZذ!"O���mR�*8<���.7J�HA"O����Z�e�R!����>e��a2"O��+1��;W�PP1�i��]/��4"O �j��rJ�
�nŇG#6�g"O��R��ڔyLT92-ً��HR"O��C� @:U7���ʊВ�2�y�H�+���Ip��'N
B��y�L�C0 ��%��7���XW��,�yb�^�l�����Fq�/>ڭ��>���8��Y�b���y� �Y�̐�ȓ�`�pE�+��)0G�4d�>1��Z$��{��Mj6p���7X(l��ȓdg���.ԗz����
vQ�ȓH�T�#�T)I����B�jV���S�? ���T�OMa 901�D`����4"O<�IC��:�"�*K�8�r��"O�\BP
��2
P�ЌlY����"O�8�7�):�:��?w� ��"O�qK7�P5�La�`�ƻh����"O "A�)B�r���L؜VBY��"O�`�!e��p}��Z�/Ut�P4"Ol�:ծ��H�������U;�@SC"O���`d�7���he惉+W.\`T"O��¶�P< �h�TeE�-D����"O��(3 ӵ%=@�c���E�ظ��"O^ � ��-�I�kXc�
���"O&`�$� =����[(�����"Oؒca͉�܈�FD�YN`(�"O��1ڑ3�zĘv�ϘmS�`��"O���R�F2\P�z+�5J���D"O�QC���|�F����G,��)�"Of,������n��_&�(�s"O�9��8'��d�ÂF�7w���"Oz��U�1�tف� �nv�pr"O6p8 �F.�6(�u�����3�"Ot@`P��&� �����6��g"O�$��S.
}0��؈`���b"O�=+�m�]z2�!���.��4Jw"O�Y�*�.P��Y "kJ�g����r"O$�Q3M�--�hQ�$*_���t�%"O05��'^�.}��h���� !"OjA��)ݑ^b�ɂ&�\�[g���U"Ol�x ��<�L ���V3*U�6"O��"q��7�~Q���ςL�r"Oby2S��*<���qf:+	FE�2"O�����b�2�A�θ�I�e"O\U#��� ��<��$/i��ˢ"O� ��E�W��ɺ�b^6��9�s"O0��eT&up:�1�bλ����3"O�m��Aӛ!Wmj����zԆ,��"O4\���ͼ:�Hhb�/�4�b�"OR�"H%R"��u!S��0'"Oy����CQ�|b��"[��Z4"O�=��L��w4D���$�B�"O��6�@��e`7�a�T�"Oĩ�,�5f�������"�d�(3"OF����*E�<�R �Q�i���1"O��ˆ�۳_�R�y[Ȕ�B,Σ*�!���
hء9f��%�՚1���s,!�d^4R�2S!��X)��*�u+!��2r�H�Qt���w^����=�!��V�Vv��J����2g���*Ō<�!�N7����h�@8���ΐ�!�D_�%<�̡u&���C�ޕ!�!�ȸN��|�WK�<FiX(��-�s!�ě �p���� Y�Xb�"��u!�D�4C�(��E�l04e;����tE!�^1A@��#�N�v*F=�!�ǹ9N!�$ҲU�Z�ss+ɋ) x�K�F"K!�W 3R��$�� l�*^��!�dxkz�+���.C@)i�aWN�!�dQ	Z8��R�F5�p���Ϥ!�;h�d���g(��K0���!�d� 2�����ļ,hukb�P3_~!�9*Y��ڑ�M�f�|2l��oj!��<��@;&���p�%�!8!��C��mT15�d��$U�u�HB�YQ ����P3izl����DB�)� Z�!O��¥#�<�0\X0"O��V�"㣁'��8ɦ"Oj|�#�ߍT{ � t��L�t"O�t ���*S?r��sJ�(bӎ��"O���d�[¬�[@�>����7"O���̼|gdؤD�X�>�"O�1��b�4*!"-F�!&�l؊"O��3�g?��x'ϒ�I6�lB�"OTU2jٕU�h�W�@e�����"O��`H�5M��a�#�*U���2"O&�q�EI<rY��)eˑb�6"O�Ya��Q8�$1��^�ԅ"O�U3�$��(������.�ą8�"O�ڕ���&�CP�<@�t͒�"OƱIp!��B�p�)3��"g���c"O�d�� 
  ��     G  �  �  �)  (5  v@  �K  zV  %b  Wm  �x  ��  m�  �  �  |�  -�  m�  �  7�  z�  ��  ,�  ��  ��  m�  ��  �  ��  ��  a � � � j �% �, {7 c> �D �N �U �\ �b !i !k  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>���f$�2���y�#W�@ݳ�i[)�d)�O2�n�g��|��?Y��MwPf=Cp#�_.6�;c$���?��uYf�;ߴ���~>р�'��S�
�9Kb�|$$�UO��e<c���Qy��S<�-P��>f��#���.���0ٴ%�4��<!��$�g����:PO�a9d5[�8$5>��$�Ol�IO}���m׫E&��4Ox�"�.��/�ʑK'���0��G3O��I9�?��+#��|��D�b`p#�]2�� Q�ժB;$Dϓ��$��Ϧ�٣J$�I~l��!���.����Bb�!C�d��?qRX�������Γ��䎔�����۾֕���@v�	��\�(���b>]��'���ɡ0O0��%
�b�����% �'Q�Iڟ"~��H�j���=����R8�ra�'�6M�%r`�ɻ�M��OÄ%"D더�JPzR���hYۘ'���'�R�ډ��V���Χ[����P�7x x�!�\ZI���C�7^��'�X���4�'~��':��'��U�̬^���it"ܖQ 6_�D+ڴ#�4�
���?�����'�?�$J��._�y�3甧O���j�C��(��I�|�IB�)�S�6����-ûi�R�kr����z�£oU����T;�����O��qO>-O�,� ��|�by���:�t�p��OJ�D�O��$�O�<9S�i�Zm���'�,]!��Q�)�3��)\huȐ�'+X7�<�����d�O��$�O��$ ��r\�C0'Q�g�N�z� �D�6m ?1a�~d:��'���	��Jz/�#͋!-Q�1ۗ~���	�L����\��ƟX���� Q�M��݂�7`���+O*�Ć���a�&���i?�'>:h����b�`)��J�H��`�|��'��OQ�@j³i��ɏ�2�p��B�sYa�/X.=�����B�O2�Oj��|���?��=�����>p��2�/�l͆1���?�(O��o�f����Iş,�	w�T�ծ�H��H*��U�b������P}b�'�2�|ʟ:x���_([��hpB��[Lq�5�6|�Y3�"���|zF-�O��kN>!�#C`�����6���c���?)��?����?�|�*O*xl*�X	�oA�]h���mB�2�^�K0�H՟p�	��M#�RB�>!��Vt�)�J�� ��2�D���k���?IF��0�M��Oش"&GD��O�҈0�b XB��$aD�tʆ��'-��ğ$������Iן@�Iu��H��$b��1L�H0'%�0Y+�7�d-4���O��$#���O6	nz�Q8W��
J��9RяL�Q�4�埨�	^�)�*�l�<�9<�pU��I�9��T(���<�c]q�.�K����4����Z->�Jc�O��XZ�0i�/�!�<��O"�$�O|ʓ ���S�-M��'�"��U��,S��t)�u�p��<��O<��'h��D#B`�Y�d�2�~�6�@
9���,0S�Փ����w�%?���'r��I�&~ָ*���S�D`+���?��	��8��矰��D�OQ��C'5��u�t�*y��A���*96��z��x4/�<�ױi��O�.��%z�ݣ��H��D9�!ύ>IV��O��D�OBy;�E��UN&��/�?m�� ��4	RKa�X�����m�F��Gy�O�r�' �'�lH$�:��3`=�`Ⅺ|�剌�MN[��?���?!����ʀ4 5�sKҹ LD��$G�-FӮꓛ?a���Ş3��D1&�0FG.�J�� _�.��ԪR9�M�E\��tŅ V���1���<ٷ'Z�TE���E@��� �?��?I���?�'�����5��C���4�����w��-(L0���0`ٴ��'�^ꓻ?�+O��A�-Y�@��U�jW\z��իɺ6�X7m3?��Q/-p����:��'��� &9�ģC^�f S�x8���;O8�D�O����O���OP�?�sa����m�.G�,g����Uyy�'U�6��D��)�O�QmT�P�V@ː	�;_Lp���K�Lc�p��hy���'��v���i���1$7P�Ό��!L�ZP�1�'F�U&�@�'���'7��'�
��FM8���� �UxA�'P�]����4j�|�����?!�����A¨(�EZ�[��%8����q�I����Oj�*��?�Pϙ7)8��i�Ks�(!�LD ���{F������|��,�O8)iL>��'���HA�Z'>�iI���?����?I��?�|�+O�m� �%���R54�ЦA��BL�95@ƋLQNʓOY���ĊV}"�'_��4�^�h��3�ڇG��"��'+"��{�敟��Wa��'�T�~��k�<s���eȞ�C�	�<q)O���O8���O��O�ʧZ� �$�9J��%���{�m!T�i|&�+w�'5��'��O4�y��Qn9P)%
��nXz��0�Q�sG���O�O1��q�t�|�l�Ɍp��x�k:(�z�R�h�+(z扁w�v��"�'���&�������'ȴ|Qk�o�P�@��(0Lt�`�'��'^�Q�8+۴V�l����?i�w���'�;'H ��o�LE��r�>���?�K>�!ƍ1� � �G�=p۴p��@�]~�{K�ɚ�i1��`��'!�!]� �~���5{�������� �'�B�''b�ǟ�0D�2�H:�,ѫP,L�C�iȟ���4=%�!Z���?W�i��O󮄄������q
�q���0z��O�˓<f|ep�4���Pl���'}�ތ�DG��W��a�F"k��Q���$���<9���?����?	��?�5b��r<��@��y0X!b@�����Y̦�	 ���ß�'?���3)
���=�n��N�3C7��O ���O��O1�:8:�Wg��Ȋ�.� #|�1��`yYA-�s*�	�0�P��'�΍%�@�'�xP�%+\%}~��p�ډ:�ށJF�'���'Eb���DZ��Y�4?��!#�
VV�!3fE�bH�JC�G�2��H���P`�F��X}��'��'6�{F��:_�����ܤ�Z}�e�݉F������j���������hdJ��^BA9��$Q҂��7O���O����O��D�O��?yR�!�.7�" zu�[�:�ñb�������X�4�6�ͧ�?	ºi�'�X<Y�b�W`m�#�I�w�%�y"�'H前_���lZC~B�E�U�����,ncX�:�J�)}�V���%����⦒|�U���	� �	ݟH���Dyr��	C�a΀���*����	Ty�y��PR��O��$�OD�'[��+ab&4P��L
Kz���'���?�����S�4B�I{b�y��4i�V��.ԯ-!T=���ڧ9��a�O�	�5�?�6J<��Ǯq���	�a��]�~N��d�OL��O����<aP�iX�͚�o�!|U���x�*d���<Y��'��6-6�	����O���p�i$�L#S�2�ү�OD�D�$��7�4?�CC����5��,������7�Ǌa�t�y/�#�yRZ���I�x�	���������O��`���o!���ə�E��T��}�ܼ���O0���Oꓟ4��ܦ�]��dH+��ծ�xe�EdP�5�jt��\�S�'N�||"�4�yBf�:Tw�9��ԺOԖ��s�[��yb�>nH���.:��' ���x��0mK� R��J���(��.H��ΟT�Iޟx�'
�6��(x����O<���P�a��C	3�X��Eg�x㟌��O:���O\�Oh�Ӣ\)j�@9�+@�=Z
�h���r�׉{���mZ<��'��Iퟸ1F�\BQ�<JF	>~�hH�W�H՟<�	�h�I��0E���'t\�8��R�\�j�zQ�(`"��'�P7��//����Oz�n�~�Ӽ�Ta=���/%��٦�U�O��ߟ4��؟P�冓���u�U�N���ސ�F�P�/G�kJ`Az�G�W��)$�T�'�'z"�'���'n����N��	�t���u�T�� ޴/ 1(���?���'�?)TO��)�ҼJ���DhV�!��&��Iҟ$�IJ�)�,clXJ�"�S20Ihe�٦W�n�1O�����'�^!��,|?	O>a.O"��&�P�Ti�'��=C8�| ���O��$�O��$�O�<	��i���I5�'q���`�P�T� �%jb��'�7m#�������O����Oj�b���n�\�QF#>!\�4I���078?ApE٤�R��:����=�`�ԟ8�< �0Z���kd����Ο��	�l�IџP����U2�
VDݐG�$F��?��?�ſiFn�+�Oc��h�|�O�XH�U0(h*�ȋ�X�I*&���O���۴��$����U��(�W�TpA� MD����%�?YEj,��<���?Y��?����	%�\Q�5��A�8�bT3�?)���ĖŦY�q�@y��'��?~3�&n\�ep�lۦ��	WX�6���ҟ��Ip�)���DT_4�2F+U@���8�C)��$8�T��M�\��0��$0��ܥ rt��w��f;�P�A���H���O����O���ɢ<���i�00�g�D�
��C�>X���5�<SzR�'�N6m0�I��d�O�%&Ŵ�4��Q��$t� 岔��OT�D-�H7�9?��"����'q���S�? � �D�;(�С��n��B���BP:O���?a���?���?����)�.�py�qB[��td#����n�7�Nx�Iϟ��IS�ϟ�{���KS�ù7/�h���A�rc <�1a���?y���S�'r��ڴ�y�֒E�\}��%ȵ-T��R',Ǜ�yR�ULM�@��*u��'I��@�Ɂt.f�a��Mww�0����v�D�I͟������'d6m/t�d�O:�$�$aR��+�bY�J�v b�+�hSn����O��d�O~�Oy�ЋX�3�n��A'�?�T�S��Ԁ��N6t>ZAy*�ӳt;�J�i��cC<��p�K&3�D�#��D՟���ߟH����4D�4�'=d��qC��kk|`��BDʬ��'6m�A�����O��l�A�ӼK����Rh*"�i[�N�V���E�<)��?��� ���4�����z��[����8\}��I�d%W1<!��Ѵ��.�䓼�4���O����O��D\�Dh�H���#j�<h�g��.��g��f��187B�'B��i�,]���Ԭݕ7�8,��T|t,�'���'�ɧ�OXF 1
C���z��U&����͞�ɹ_��X�-B�6|��n��Ry"�P	f,P�A	6T��)@�I�F-r�'?��'Y�OS�I/�Mk�,#�?��ڒH|Dj��|��@���?�B�ik�O4�'��_�X���WA�.��1"��F9:}AF�0N1m�y~��0@������K"�O�g+�f��0��L��d�\7�y��'��'N�'�����'��	�b؁��=���[�G�(�D�O��$^��]���x>����M�O>1B�K&56<d��iM�v����S���䓖?���|�fO��M�O�Pk�i�j�0��`l�RT�P��׏8��ŀ��ēO���|����?���6�li��%il�I��F[mZe���?q,OMm8���	����l�T*���dI+��C5f��A����d�G}B�'�O��Y����i�u�pJƔtS0Ma�H��L���FVuy�O8�IY��'�v�q�+�4+b�R¡�2�D��'���'=����O(剮�M+ �."t9��(]�O����K^�~]b���?iǴi;�OH<�']2C�1=�x�J��X�C�VذaNՒ���'�(��G�iG�iݡKӥ��?��Z�w7x��C�B�R���aa���'��'��'.��'��/&cL�u�A*U���s�ĆH�4�۴�R=h���?����'�?�&��y�̓	��JP	�Hw"4���چt]��'�ɧ�O �����i��� 8*�bisÐ�V|�L����h��d�7"QR�?�B�O$��?��:�tY��&�}�s�O8��a#���?���?Q(O, l�E����	ß �I��!�d#�j��#��a���?�\� �	ɟ�$�<S�͏�d�4]�A���\��f'?�0�V?	�\M��4%��OZ���?�	�D2r0��@ڽ>�|�y���&�?���?A���?�����OL�$�̱0�Xk��Z[P��O��oڮE*���'o�7�*�i��c��	e����
�xLHEIi���ɟ����}[b�o�y~"B4P]�'8�,8��n�*aT�}+7OL� ,���K>/O�i�O4�D�O2�$�O������[��4I�ކF�X,`Ă�<�2�i2�Z��'B�'h�O�@0?3�X� ̄�W F��#��b1��?���t ��@�c�K�C[j�q2l�RQ�����^�剰A�Ja)0�'�z�&�l�'��]�����`i�lƫi4�5�'���'�����T^�@k�4m���B�-����en<P1#�+w�U��\(���$�J}��'6�w������6�H0�r#
|����Ā=-�6����J\+h!��1�I���<1�`]+BP�a���;�(�3O��d�OT�D�O��$�Ol�?ͣ�Ƭ$Z���ϗ�,�B}��j�����	�t:۴sԉ̧�?��i��'{`H �@̚?����M�< ��|��'9�O��p�i���R��+�O�}��� t%N��IA3��8B��$/���<����?y��?A���k�&0s��3 C�|k�mM��?a���O���K�F��H��ҟ�O햐� �%	���c�(��O�(�'���?�4��'\��d#��e�k�	A�ؙ�D �2�������bS������|���'����'�1��D�!�'��'R��W���ڴ�,��g�՘+~@��s-� pL(e�)�?���\ԛ���u}2�'��A*Ϋ*�ȠS@.:I��'�r���������J�G,���~����]ְR���N�h������<y)O:�d�O����Oz���O�ʧZ��1��,YXp` �T�S�!��i���#B[���	l�؟������G�|l�p@���?B!�(�,�?ɉ������$ԛ2O�qC�٦y�֤Vn��H�ɔ=O�m*�h�:�?�9�$�<I���?ɏ,o�lH�� �a �ʵ�;�?	���?�����JԦ�i�%\Ɵ��	���
�[  ���	wk�FLD�	c�n�Sb�iM7��O�O���&j!�j. ?��;��m���,\t~Ę#�P�c>�c�'�y�I+Yx����2\���55��x����L�I����	l��y��h*��pg֥_l���(.�"ao���8�b�O���N٦m�?�;P��!��zP�D��l��/-x��?�*O�yee��8�:���"����� ReYI��B��+�Da D,�D�<	���?���?	���?�0��(O`N��V�ՄG�� �����ڦˑc����I�|'?��	��\�ʤ.����v�ɣA3*d0�O���4�)�Ӏ��԰!�S�-_z̳���)$��@���A.�ڵ�'���r�F�kG�|�Q��C��Z�u-��4E_c�l�� ��H��Ο���̟�ayB�f��/�OnIq�Q8@�xY�p�8-�(����O��o�o�A���ӟ0�	�|RT�K�1�14��!���{���\[$ lj~��Y7g_��'��'��`�&p��CE�F�_�b]f�<	���?����?i��?9���xz�5�^=�`D.�pc��'8�aӸ�Y>���D���]'�h�P.�=\?�:bn\4x�>!�&�d�I� �i>�R��ʦI�'�&,q�=��i�� vB
�ҡi,������4�����O��䈿9���iԫ�g�`�cj�$['���O$�%��/Z#A��'I�W>-@����܍i�N��;�Tq��-?Q�T�p���p&��3�����,T�`����
(qpX1�:8�:1I����4��lB����O��P3)�8ky|X#���	� 9�B�Oz��O����O1�ʓ&��0h��9p��I�@0�E��R%�����'[cd�:���O��ǉJ�z�å�O�Pw����@�{�����Oĭ�CA}Ӕ�Ӻ� ��Z���<�pEϓ\]�mJ�o�^�hmJ�	��<�-Oz���O@��O��D�O�ʧ}�����+4!��U(k(�S6�izz���'���'��O��`��NT�Y��BtCVZ�~�A�YGЉ�I|�S�'?�H�ٴ�y�6[c�wM��!Uh�&o��ɱ5 �I`��'�vd%�@�'X��'�"hק��|(���a +߬��'Fr�'�r\�����x��	�4�I(�
 {3gѰK�xt�#Ո_��9�?Q�[�����T'�(`r��@6�+Q ��/S��0�7?�W"F�6D��!�s�'
>�dڳ�?�O� �P���Ǉ=�(��d]��?���?1���?��9��"
ˢ�
$�Ŭ�n0G�#���}Ӵ����O������?�;h:^`���!$�P����v���?���?1�,^��MK�O
Ԫd$C.�*�)B�{SP���Hڐ0�D	�"�{ �O@��|Z��?���?��7&��E��<=���
G"~� )O��ɸ1�����Oh�D.���O�mxFZ��� ��?nr��/F}2�'u�|���eE��S�mK*	
ΉI6�oP�
7Ͽ��DL¤��z���O�ʓ}�
�:�bN&G:�]�0&<�>IK��?���?���|�(O�tmZ�����O�!��&C<y�ʐ���1OR�a��O��oX�
�������i�E�� [B�t�(�fК5��4-���o�R~bkV�B�&9�S8t�O���@Vj���"d7�$y \7����ڟ�	�$������IC�'W�����:��ո���%�Y럐�	ޟ���4[Ӕ1s-OzMo�y�IP�bfa��j�:83��^0j�u$�8�I��� ��7�-?�����o�h�ɐ�c�Qx�NG�o��&�Oy1N>�.O��O��D�O�� ��D8�����:��٘��OJ�d�<���i&d�w�'/��'��ӓT�V<@����Y�����6ujR����ޟ���B�)Rsh�&q�N�"0� �4�Ҍ[��G<4�&i�c(�I#���4�˟聖|Z�R鈑U�^+��v!U�jvD+���?���?9�S�'��$�Ϧ�9D�I9ON%2���|�0�i��t�����4��'0@��?�"H�$���w�
�a�4���[6��$-la�6�>?A2
�zզ��!��Ā�3�@i� ����U����o���<���?i���?����?�*���X�(O�(+�|��k�/XG��kd-X¦�YF�۟���ڟ��B%��yG)٩_�0f�ʵFV��_`t���I�1�06-v�8Ғ��P,B}���&��(Vb���!�|�2�_�IEy��'��kԀd���Fm�1�^5;��
	�R�'���'��	-�M����?I��?���fK� ����;^ʀp���'����?����ڌD$�� -ؘ_4tY��)���$Z�*�4��@'c���(���%c4���I\�A���Q����b�4
E����O��d�O*��"�'�?���ٛN��rDŌ�
CN��BoP��?I��i~
��t�'P�I{�X��.P�,�ۦ`�)4Bx��ao��I�L��Ɵ��!N�Ȧ��'��$d��?��$�ӺI����r�ǔ
�H�Ph���'��i>��	ퟬ����D��>i����B��#>^ҥ�2�̀*? ��'��6-�l��Ob��0��3J�X�h!EK2RoΑ0������OR���O��O1���� � "�p=9��H(��u꒏"d�H	p2����� �D�BdZn�	Jy"�0�j����;����Y�eS�'3r�'��O�創�Mӡ	�2�?Q��;%�%��(�'��I4����?�e�i��O���'���'���{04@[�Iѵ��h���*5��S׺i��I;��(W�O�q�h���N(���`�F(���7C֧dF�D�O���O���O��d,�ӒP�I1y�+VN��X$�Iٟ �ɶ�M��EX�|"����|mM9-�,`H%��/���Gѭ��'v����d(�J,����L[SK+� 6Eid��$S�.M1%ͤ7���R`�?a��2��<�'�?���?��P9EjH	�M�)J�s�8�?���������s�\py��'��S	�L�6eL%?Y�D�#G�x�hI������	K�)"���'V\x�#�ϼ_ʭS�e4c8�|�bp����Å����|2-ԁsP$���jΧ=�2����Œ\�B�'�r�'���Z����4i.B<"�/L���zb���eS%�Ug���'��6M:�	��D�O&[A�T�(�%+��J'�B��k�<�'螳�M��OJE;���2�Z�(�<I�(^�d���_�G�����*��<�)O��O����O����Oʧ&�t�K�/vH���=��$���i#.`���'�"�'D�O�r�t��.�:���h m�2U~H�0o�/Q����O��O1���0�Ol�@�ɒ)RhLS�@U1ڼ�F�Y�z](�4%NTI+��O��O�˓�?��B��q��$���v���R�r��?i���?	)O�mZ�_.|q��ȟ���7&px�&��?Yd����:=U�M�?	�W����˟�'�h��"�iQȜ��-�8��	�u�9?1�S(.i}�4^��OK����?!q'�r����ئ-�^�rfŧ�?���?���?���I�O(\�P!�%X�H�y㢘� �Hx(f�O|�nm-^ �	ȟt��4���y'�ƫg���qhu@�3���y��'�r�'j�T��i����c�ԟ~�:�H�&$�X��/.4Wh�U�>���<���?��?����?����c�p�s	��,yn(��fN���dH��*a	�`�	Ο���A��8�DŎi\tCrC	(����L�	P�)��6���r���&@B5XU䃯b�N4B� ����'��1:(�O?YH>,O����F2R�Xѣ�/Ks� ����O����O����O�i�<�#�i�!��'B��"�EP*K&�j��\B�5�6�'�7�)�	���ON�d�Ov��g��.@ĸ��E�]�0����GW�MS�O����8������w�m�w%�}���{6��e�P8�'V"�'���'�B�'��$!+�C�P�4i[ve��{�X*��<���}ț&cǉ����'S�7M>��	BŒ<!�Ƽ@Jz� C# ��O���O�iQ&7-&?	b�X1[���2c���x* ŀ�Ǎ ~�|l U뺟�&���'�r�'�R�''v�C3��=Pn�ZQ���y�t�y �'V��"�4%�L�9��?����	��>\KW(�n�c0A�lA^xr�OP��'!�'�ɧ����J��2��.	�J����ʎP����C�Yٮ��0���S@�"ai�I�E2|�^��Xc�X�qk��	ϟ �	؟0�)�OyB�v��A�a�+i�t�1LJ�hEQ�Ș$0�6˓K���Kp}b�'�`{gC�@�ݫ�������'>ˍ~�����&��m���~�	�?nh��a(I��8	2*�<�.O&���O�$�OX���O��'Z�hM)�h�*Z�,��&��zj�*4�i%t�Y�'���'��O��Cb��n��V'����ݙD��C@F:6l�m��џ�'�b>�{�/ЦaΓ'�F��`�D �S���p����f��A��O�@M>�)OR���O��Y��I�MXh5�,ކk�5�"��O����O��D�<)2�if�s�\���ɉM�ʽSJ�;k��e�S,��9�"��?YW����۟t&��2��à/��)���ۙ�{�.?A2ǷX��a��XA�'S����Y��?��9�p������H�9p�N��?����?���?���i�O��#�	�+8-QЎ8����'�O$En3c��	П0hߴ���y׏�O�Y�dĩ[\n�s5�7�y��'���'��@�b�i@�ɗ�\�ʲݟ����J�]þEӖ	Q<O����##�D�<����?����?���?�*ß9� !q��ƥtec�����WզU����6�i����'�:�[�R��j���C%n˒PZų>����?N>�|�M��KyNPB���Iy@��u��>��}ۑ�Ey~��\0^vje�ɉr��'r�	X������2[���G׼#����I��L������i>ٖ'ʜ7�S^�D��g�8kU��B\2�ٵ��1�<��W���?��\���	�h�	�3�>��o�'F�z�ha�`L3�L�)�'M�h ���?��}�;N�ĸ��!��͐��΢RQ���?����?���?�����O(�!�ů��~�D����:}���R���ɓ�MK����|���:���|�H�X��bK7��)cJ��ۘ'���'4���@�v7O���A�E���$gg�)�O/ba��SV��?YF�8���<1���?)���?p
�@�
MyC��<m��ْR���?)���d�Ʀݪ�D������h�O�����/�}'fu�Ճ�{����O���'Y��'�ɧ�iZ��m!�g�rX�p��/��5�r���/&� ���據q��lN�ɽ|�ꈢv��� u ��+}F������	̟X�)�Cyb�x�T�Q�Cnڨѡ�?t�
g`�a����O��o�u�]���ҟ��Ō��H�zQ$DL5|��P/�����uG��n�S~Zw�H�j!�O?|��'N)C�T4��yJeiߎ��I�'���埴�	ߟ��	����}�ThŁ ��})�f^�Q��KQn\�~�*6�*���$�O���0��MϻS�.$��d͔G�ђs�3D��;��?9L>�|�p@G��MӜ�� ��9�*�v���'�D�_�r��$?O������?�E'���<�O9(L�"��(RB�H���vD�-pÓ����ѱ�R�'4�-��yM���P���R�a�p��O���'���'��'���en��A"���P���+Gn��O@�;��'j����5�	]��?���O
����U�r�0�X3 P�Wl���"O.9"@hG�\�`xCv�'1Q�Y�`�Oo9������xi�4���y��;����F͋�98��1�yR�'�2�'���־i��<kN�b'ܟƑ@��ۛl��0�S�e2.�QdF5���<Y��Ď�K(T�%��:	ʨ+��D�(P��3�Mk`��?���?���G� f���� A.�HRb�W6����?a���S�'BpP�˒��?�t����Ҷ)T���cNV��MbS�H����s���/���<	���|�`��5%���)��_��޴~���)��V��{��0t�$tS1�",������u���D�~}��'���'9\Q��H#vI�&�75VaI���_ٛ����X% EVS�tȃO������Z�e&�����U��|��n�P��I��D����/���6K	�c�`�I� ���M���[�Ԅk��O|Pa��洴H�Êf=6�`�'��O��4�f���}�P�T؄�B�s,D���敓C��H�S[H(��n�Imy���~F��TD41$ܡ����s=�p��4l ~0��?�����[�j��e	����}��*W�H��	�����Ox�d8��?m�������m� g��J��u������0�ŉ��	P)O�i�/�~2�|�1v~\�B��ݻ,���S���FZ��'@R�'���t_�@��4j�3�nFv���0��M&�}���N��?A����F�DYo}"�'ʢ�b#�X �q�0mC(BvY��'rhWk�V��D8��q��ɧ<a#�O$I��0��N/����<Y*O����O����O��D�O
�'1C�!��<�>@G	�s�X�ҷi�n��'�"�'i��yrn���ˡ��|�P��&lf��a� 6�|�$�O�O1�ؼ���bӔ�I�:U�D# ��&�1i%C&v���	4�1��O��O��?��E)��8�ӽ<	v£�����h���?���?�(O�n��R�
��Ɵ��	x!p�ClQ�nq�lIЧ�?�Fl�?�QQ���Iɟd%�dcĠM)��`/�/J%f0�ը9?�Vg�����4^��O�(��?y�ȋ_Q:XD �2��q�m�,�?����?q���?)��	�O�maG˷X�
H�0���:h���O��oZ�?Xd��IƟ��ڴ���yW"��/��	Bؓa�ܠ���y"�'�"�'`�Mh�i.�� 7��UxCԟd�Aɞ�#�"Uje���!��k?��<����?���?����?�ɏ��(����$Ui8��d��+��$B��� ��矬�Iğ�$?��	�C�D 0�C�}T��2�@�`V �O�D�O�O1��m��Ą�;r�G�¥8O�I҇/�	n47�O\y�L�.|�N������ٳY���1d/&ۄ=�%	�Kk����O����O��4��˓rq�F�55���Cʞ�Y��K%^��� ��y�i��{�O:���O��$(:ҞI�Ĩ`��a)VF�`j$��Jn���] ��
�?�%?���&6-��eG�#�s�#��0��I��<�I��������I[��q�*qꃢ��,r�J��j(�a3��?q�L��V�������'�7�3���%~��󁈎`xdq#�{n�O����O����7-!?�qI� F\���W�[!r�r�	�k�.͹rD���'�P�'��'�R�'x@�2���	d�X&Ƅ�Ô5���'iU�ȣߴd�a���?q���)Axi��Z�2�v�	�B�
A����D�O��D8��?�� B	�Q�ɺ���FT|"פb����Xæ*O�i�6�~��|r��1B�:`�eJmf��x�H��xbDdӜ-�*�4^�i�̌:�ԓ���	~���d�OF5l�_�5��������&Pf�9�W	v�,�1b/Bџ`�	~�.n�y~�	��x��E�'���Xhx0�6�� �*�q�Q�X�$�<���<��K[�Sw�Ԋg��@�u���i (�(3�'p��'񟐄ozޥS&⎠5�H|�'҃}������]ڟ�Iw�)�1&��lZ�<9C�L�IB`A&IUo�3���<�$D��o�:�$]�����ĥ<��~��d��k���ʁ뚈r�|��æI�n�럘�I̟��C�]�Ҩڐ(�[��][֧Vk���I�	R�$(\HK��P�JS ���ݹ7���d�& PTM@��M�`��ԉ�A?���VEH�i�xD��k�MZ�L���ȓG%�a�2+�68z���e�v��2��V��r��'FL6�,�i��ܖD�>rƋC�U!8���(C�yB�'�2�'�D�Z�i���N}�h��П"\��*&Ȑ��ۚ.=ҤӦ
+�d�<����?Q���?����?ɧ��<���i�8�f B/Ƚ����)I%'AП�Iݟ|&?�IC]�@K	����;�߲cx�*�O���O��O1�j<��� �ya띔Z}� ��>w�0e3��C��I�}��=�6�'���'�0�'�������f���bR�w3�i��'���'3����X�p�4 h���}�}Ç���{͂�1f��'�<��������B}b�'/�wW����'�;�[�ѐ^��4�`����@c�Ґ7���+������舜~��@�e���� �8O����O>��Oj�$�O��?����'o'���������z�M�`�I�DI�4n#���O.7�*�$�j�>��s�F�!CGʔBkƒOF�D�O󩁹/��7�4?��!{��r�\�$0$�:��҃U��]i�ǰ� $�8�'��'�r�'�r�x�K�3`�ȰHnN|Q�p���'��]���۴k��8���?a���	Iwr�t�O��P��?7���-����O�$*��?���@�
a�����Ӏf��y v��XNd�"dy��%�Ry�O�
I���SO�e���ϋu�<=��o�J�|��?q��?��S�'���Rܦ��Bl��-0���D��A���ƕV�(��'y7-#�	�����O�]z��U��t�Hg�+e�j���'�2&�i��ɏ꤭�ݟ2ʓ)M��2Q��):9x���M��������O����O����O���|:��WY8P��X?!^��d�R���fA�*>��'�Ғ���'_
6=��1*��o�R��7e�
74��
r��OR��5���?Qu$6�b����)K$�`g�z�`pڳ l� ��A�9s
Fg�xy�O>�K�t���!Ѱ��7q�2�'���'��8�M�v)���?I��?�rg��0��w�%_41��#ײ��'�z��?����=�n�pVc:�0�9uB*=��'�!����z�����-�̟����'�2!T�M�2�U��&�����"�'���'4r�'��>}��>[�8��D�@�?��b�ʞ�R����I��M�`ꁐ�?�������4�.\;'�ΜO�J�˦b�:�p1��=O����<I��X&�M��O�M�#�'$B�q!(Ѩ����*RE�˘�K°�O^˓�?����?Q��?��#4썓T�#P_�����@��|�(O"�m�(y�j��ǟd�	j�ǟ�p���!!�=��:^�������O��b>Y�hѭH%DU�%H�?sp2�b��Ԇ���bZWy���/RJ��I�i�'�	�]u�W��K12�@�$t`z\�I������ �i>�'�|6�(<`���Q	V�#F���J�Ɯ�b�G 5+:�$���-�?_��Igy�G��^�Ȳ%�کv�� ��R�Y
8��i���J�f�A��O�li%?��  fM�4����vy[��[��:O��$�O�D�O��$�O��?�kG�N�j}�� 'gܖ�q'������	򟼂ߴum�T�'�?Q��i��'.��St��.p�&h�gi:az~Ń�yb�'��ɟ^��elZ`~�B
6EKJd��NM�E�	!go��R`V��r����XD�|T�������Iٟ`�[~
picaO-%�(ͻE�T�����qy",q�:�-�O����O��'OD��x�O0f\��CiW5$���'���?�ʟ��n�c����R��y��#�fQ��d���Կ/T��|�U��(o�F�����!Z��x(w	��R�1�S�3�6�AnO#B\�$��#!��Q����d��N�F���P�����J�hB9v4�	W
���ͨ�)�-��f.h,����HOzL�$�Ƌ\� �V3��hu�58,����ʰB�p�sT�/.=��c!��g)��K���?MAH��?,ZyU���n�2��5UFA��&�����[��ҌI!��1��8dry���	�/Zv}����y���a�����@䊡`��fGdh $H��ݫD��(�YH����Nx�éR�;���L�>�/O �$=���O"���	ib��&��8p�PH��OVE<٩B�&���Ob���O��o���S7��T�v�F1|���ڇ�nR$���i��ޟ�$����ޟ(�#�O?�� ����ڒH� B��iitK]}��'�2�'Y剳:)I �����p�ry�b���ָ�R�S�Ί\mΟ�&��IΟ���VZܓ
����p�O�!�(�ٱ*X=I���l�̟��Ieyr�ޙh�b��?����"+ݸm����v�ƙ!N�!����'BR�'J}���ĥ?i`0l���Ѯ�$l���o� ʓ>W�$�W�i B�'���O6l������r�м�$��T��l��Q�Iڟ���DPk���Og��aH�c���`�*�h���4)��-�T�i���'<"�OP����d�]�|Y`�9C����A
,]luo+*�4��?��d�'���3��P� �J�:����G�e���D�O@�dT�&����'��ȟ��tϦ0x���  z�Y1�T�N�,o�T���M&����؟��i��ۅ!K�u�eib�9��A
�Lz�2��ǆL\��'���4$���5�Իu�n�V(�W7������+����Oj�$�O��V�80�R1 d13�G�d��t�e�M5���hyB�'I�'�R�'�f��wK�^��U
5�� �}x#&+r��'0��'��^����ƍ"����d~�"���	7��x'�[��M(ON��!���OL��L��D2,y�����R8�Ё�M:P����'���'W_�X�f-Ǩ����O�+ N�wu@X�aXG�t��ɦ-��`�ϟ(�� k$b�t��M2nX�4C�J����p�,�$�Od�AfHJƖ���'*�\ck�(*�HK�*�ZQa��̅L ��J<�*OP���O8����� H@�Q��+��"A�C17�9���i1�3ql�ٴ5H���ӌ��d��bJt�+G�� 6Z��B�!\�F\���ܟ��J|J~nڵS���V*5	4p@�C:{��7-�1v�Ho�͟��I����S����|
5�6�fey�$�j&r��� �+D͛��'���'�ɧ�9O��J���Sb`��;�� ���Y���n�˟����|�č�$���|���~�a`1��2�	�@0��h��M����� ��3?���~R$�-inPp�'�>,�и� �r�X��P/0��M��Sq�[���J3�Y#a6�" �!u��y��x��ݏ��'�\�8�I.�$d;��N�D]"������Kpivy��'Ur���OL�	1-�l+��l`�	8a��0w�86��/1O����<	�{Ƚ��O!���A'_n�刲J"zVe:ٴ�?����'��W����b��Ӆ�ݫa��XG(�<���Z���䟄�	Dy��ьc��v�8���=��)��k�P2���]Цq�	x��{y�OB�~"�'R]'X���\.S�������Ħ��ǟ��'4.)��"�I�O8����U���@�w�6ٱ�P<L�$�x�S�����'?�i�1Y4`Z�B�L�Es�����*�>�Eu>����?���?��'����(���v�z�qE�&��D� �i�^�ˡ�%�S�S:�(��"L���hA��I��6�	�W�Dn�蟔��쟔� ���|*EAG;V8\s�W�r9F��V/�+uM�V�'b��'�ɧ�9O��䇕N���o��J@�0����m�֟h�I؟P��&�&���|���~rCƭ%�<5S���!��c5�+�M����@.�s���I�����%x ` ��U�gYf��kGTJ����4�?ɱ��R�$��Sޟ�&�d S�xŸݠ�B�&�H�卅�ē�?�H>�������OZ��5�XuV���;s��p��K�OB<��?�����'���OjL#q�֋6���s�ԣg�0��жi�(��O��D�O8���<9A�)~n�I���p�c�(��"5j�H���ݟ@��i��]y�O����5!�d��0F8�J��p�Q�#��O�d�<���Y���-��$��V�����A�b$��o� �o�r��?Q.O��KQ�x�#T�=H����X�s�  ���Mk���$�O8� 
�|z��?a���Cϙ�7��Q���*L�z9��OUp�	��'1"A������ak�
��i��OZxk~��\�T���y�X4������I����syZwؾ���Z�e����e�&����ش�?�*O����)�)Q#\����W+ϗ{�T`��ߌ$�&%��X9l7-�O�$�O��)Zm�i>�W�X�,UP�xU��Q�����߄�M3��?1���S��'B,˽L�j4Y���L>��m	
�6M�O����O���2A\�i>��Ix?��J�q�(uQ�d�H�Т�`	ڦE�Ie����9O���Ob�d=l�T�GB��)�d�{,$HT�mH��#�6���|�����U,���c��)~�U�ª~`��`�x��'������	��d�'r��5��8�e��J�'}l��ٷ��X�xO��d�O�O��ӺK�d�NYv�W��>轩քF��	Dy��'+��'�		��p3�O&j�q�P�����Җ[����4���O�ʓ�?����?id��<	�&�4\)���(R`�5��J3n��	���Iٟt�'��d�~�������уi���%K\�j��İi�\�����������Ily�N�qŰ���L�WnPu!G��{d�7��O4��<i�Ȑ����ٟ��I�?U�F�A�w��1�� ��0M��U�����OR�D�O.�������'j�	BM��F"�X `��TF�˛�Y����O^�Mk��?���jUV��]�A�$�a�
Хt�b���H�+\Fp7M�OP�CgV�dn��'�q����` �\l�����U*O9�;��iw�d	a�m�,���O����ܱ�'�剩 ��lPv�'_ �Jժ�4D��4ID�����OAEك��=�Ej��Z0$�� |47�OX�d�O�i��Pf}BZ�H��e?���z.�	�&��'J��}����O��Ŀ<!�� ��'�?a���?�Ǜ�� �`�ّd�6�)��^4)ʛ&�'æ2C�>�*OD�D�<����
\"\�c�`�HR��p}B.��y�P�h�I�%?�)^$# �9��̊�{`��#�_�b��)�O��?�+O��O���]V������LL���7���r;On���O����O��Ķ<��D�S��	Ŕu�l� �,Bj(��f��5
~�^����sy�'B�',�͸�'�����aJ�1��Yb1ʔ�M�>����?�����D�%K�H-�O��tH�C�jA	M��Y[w�]z�T6M�O~��?i���?qԧ��<))��&n�|��`��kz$p;'.���MK���?)+O.(����O���'�r�O�zx��HC�m[ށ�2-�-'�ҩx�m�>���?��R�L����O����{v�UP��e	��Zf<�6�<Q�k  $כ��'B�'����>��[�4�2ʏ�f�F�
���4-��lZ���2�T��v�	hܧ�&`
;I�E"�	�1Y�Yl��};��Z�4�?����?Q��+�	dy�&@��  V:|J$$���2�b7-��k:��)��$��� 	� ��C B�ve����͟6m� 2��i<B�'v���@t����O�IBb�*�KvL��I�p�:7m,��G*s��?������?�Ma���?&5D���,�7w*�l���\�a��6���?�������d�<o7����Ή�1,$���M}b���yrQ��	ȟP%?񋱣M��<��b�x�e@R=Q؄I<���?�K>����?9�K�6��Y���)f���3�f�r\������O��D�O˓ "je!!8�^�h`f�4�\��G� 4���趜x�'�'-�'�	���'	��ޭ2�j�ІX�z�h)A��>����?�����=4
'>U�G��U���k��U2/�V�;�ʊ;�M+����?!��sXLC�{B�E�Z��P���Ҍ(�x�c�b� �M���?�)O~4��"�m�S����S�Z����o�0k�P� \0�p�I<����?)�A_��?)I>��O�r̋��\�BQ��DG�B$�t��4��$�=;�n����I�Ob�iFa~�ߗG~isP�˞!&����M����?�UK��<�H>ы��͂.sP�5x�Mܕ@@�$�"��%�M;tB��hl���'�b�'����-��/sR}�U�OL�0`6���#���K�4vĢ�͓����O��+WS� ����<����#�Y:�7M�O����OĀ K|�	����t?�r-��zOؐ�dIy��;�	�$�0�$�\"��'�?����?���8Yָ��#+<�����)�?I��E�V���D�O�Ok�����x!��D�~UL2'f�E�	�O�N���yy��'6���E�Me������[��\C�)�]�BL���1�I�0&�p�	���G��z�4w�/�f�b���.���cy"�'c��'��	/F�h�O⌭����M?8(򍚹.�S�O��O�O�$�O.@(�B�O�HXoIlTV�p�ǒ	���K�$�{}��'���'0�ɜ~H��iI|R� ��@�$ͻō��-��v�<	��'��	���I��@���l��OЭô$�m|������|�x�I'�i���'8�ɍd���AJ|����B�D�b2�
��_��",X�l++ډ'>��'tl�'f�'W�)V:U6�1����Xy40��\7hě6P��Ն��M�D\?����?�P�O�Z�i�}O�]	��O7aH��»i���'kz]���,��%��HP��&	��,a$�ֺ��6M?n	�1lZ���Iៈ�ӌ���?4��{Ŋ��ՑXO����i�;\���R2�O��?�	���p���]q��(�q�	[~�1�4�?A��?�aK�/Ae���t�>	�E�
�V膋i�2��N�����?�'��$�';"�'� i�gϱr��) �ˏ*�n��~����E��%��Sz�'۾�	��<M��a� $5.|�#�c�Iԟ�' �'wRT�̑�M��7p<�q���}ْ�ِ��<�֘`K<���?�����$�Ot��P��%��o	�`��2��RhH���Ob���O4�~���a&<�.�'�oY4�pgގ^V(���i���ӟ��'���'N����0�����9_���g�ǒO��Iʟl���x�'��5;G��~���0��*�K5�R�D�/|��u��i�rR����ן�Ɉ��I|��JW�UB��N�� ��Ϗ�(� 6��O��D�<S���~"�S����	�?1鉞�)�4G�qy� �/L��d�O0���O �*2O��?q�Os�����P��e�&��Xݢ��ٴ���.u,�n�����	Ο ��������YY��@#ay�d�q�Է?qv�Ӈ�iJ2�'�F���'�0��?���됣%�ԍ8&�V�[���!3k�M;�B�:ně�'yR�'��D�>�+Ol-iQ*
2�D�چ.�1?�� AbM�ͦ�rU�p���IZy"�	�O����iD�� h�\�xmJ���ͦY����I��R���O ��?��'�RxАGN*����p�"�8:�4�?!��?I���<�O���'��AC3B��e��aW+#�8�)')ږkOz7��O^a�w��g}rT�8�	]yb��5��G; ���i���@�΍�e�4��d�
gG�<���?i�����Y*��f
�'����6�+f������k}�]���y��'�'���z��,�M���0)�h���lL��y"^����ៜ������	�W|=�	�S�����N�00 P�z���ǩk�D���O���.���O�ʓ1�2l3D;^��BK�%V��=�ʟ?+X��?���?�(O�$b�jB{��Wa�ā�Κv2�Bg�4yuBP�ٴ�?�����'|rݠ���
�$���ѫwb��钒�M����?q��?���$�?A���?)���bU��&�VTTD��g랹D��*D5�'�2X���CM=�Ӻ��-G�XR�� ��ٍ6
��pG�ʦ���ٟ|�IA��IOy��O�2��5�/G�`U�U0�J9���Q����M����P+���*\y��X�)�pm�D�ĕ�*qK��i��p�Ot�F��OZ���&��V���j��,a�2$�$����r�4z�����Ϙ'D"���ԭӼ#h�H5��`.�z��o�����Ol����&<����O���/���D֠4�.ѐWR�cou��^��៌�I럐��dN:Y��H"ℜ9J��}X#Fʎ�MC�	!0��p�d�O�Ok,E0�6�
pg#��A�3���C���G	b���Iğ���^y1� ��;C��*��x"Gԕ;Ep�t���O��O���1���O���K<Jj��Q�MK�}(��򀈉u�>��R��O���O��RCzٻ�:�$�A�,H�}[j�� `�7��s��x��'}�'���'2�� �O��+f�G<O�`����2? TY�R�|��ܟ���ҟ��3��U��ߟ<��1kaD%2CÙ�m��c�%M���Go���D/���O��3FY&�\r�c�7 &ȍ�P�28��3i�6���O��j��=����4�'L��bS�&Hb�9WG��^��΋)�6-)��|A�"|���50E%
\s�!��A$3��@��@bӪ�D�O�1cf�O���O����b��CW�O�0{����π�u84}��������	_yR
�O�O�����$֏9Ѧ�1���.A��4#4���i,R�'�b�O�O"���%txa�vA���-2|@���l��V�)�'�?���0Xd��:�"V��p�diX	tN���'�r�'�U"�)�	ݟ�5�t$��+���: �$a�>��>y��z��?I��?ّ�҆�5b4��Z����*�6E��'̍9��2�I۟|%�֘.(��|�Z�
 ­SPo"i��'O^P�<A���?����MV��p�n���N�#��(j��Ӈ��O��?9O>����?���_��*��GC%O�8R釶4��=y'��>�N�"#���s�]�}Vd�	�/�[ŲM�7�?Sr)V"�D�qG*S(<!�틱X��d���L�Z!zs��tܓE�����Ya�˟�k� ]i�(.Ox��H��lDPT(�jO"3���.8*mBX���G���T��BI��0���(P��iBlB83[L4�r)&����J�,�2A���@!4Y�d�0IP�Q�Ͳ ��Ñ D)$�ql�����(Ds\����^+.Ί����'�.�P��l���D��}�Xĺ��'E���0%:��OI$M��`� BY�>u�����)շV��q�޿Zd��˖dŰ$[�W� ��t+�Ri, ��Ɗ#	��p����*N�J<�O/�u���u�0�*�Tⴽ K�dy���O���#ڧ�?��a]	A��(����= ����T�<��.K4��em�>V^̒��
O��Y����6�Zr@�E��\H jP4(�l�' "�'��Lrr��7v=��'?���yG@�6�n��v�$%�jљT��)
j؉!1͚�X�N��܆s�� �Q�|�
Y.A�l ��Y�2d�Թ���9�\�@b��DwV�$��!�$���L>���٢5��Ef���c���
 ��x~�F7�?�'�hO� �2�.wE��"�*~���0�"O�:2B�)2��+B�P��� V���i���?�'{���ӭ�O;��S��0	z5q�f�4 u���'_2�'­a����ӟLͧ����bt�Fi�+%4��1@ÛY,|�bB�K�K��8�퉻m8�H�EG�%Rv��aKM(L�@"U*B?mT
���AK���=ї�
�$�eB[6ibE�+�t�^M�	���G{��dP<� $�WFIY�P`����!�d�6\<�I�V��^�z�bU$T�	}1O�=�'*�I,%��s�4�?1�I���%����7�{ ������y����?�������?�O>1w�M�Z��h:O�&m=\s�ʄO8��`o8�I�3z�	ë�Rq ��Pb]/�l����:Z��|bj�>W��xC��B�� �
̯�yBW�G�LaR�_�L��]�1�Ó�x��h���v��|Bޝ*#�I �Xb���&�\l�ٟh�Iq�a[8�?�S T�� �0R���Xbʀ;L-����O�ȋCa�Ob��g~�坌s�ƥ�ɉ,.=�\�����I�n0�"<�ztm+W�vl ���4�b�X~���%l�����%��x	�A��X`]@�2N�!�D	�Vb�!NYb�9�	P�axB�/ғTԘ��	�?v�@!I�c7�ZU�i5��'�+��i���A�'t��'���w��]+�@��œ�0$ms��$[�z�y�A^)�~aR�bN�d9.�ؤJ��̸'Ђ�s�d��+0�Q�RV-:5<j�,�yB�<�?�}&��@��~�<L����K�^v!�DELO��q窃8(P��J�����HO>%�c�؆u���%"I7Z2���N��>eh�g����	ʟ���u�'M�4�֬��� A��dc� ��f��C�R���'�ظ�*
�x?�9Ce�K�B�M.�xr�
�D �l8Uǝ6�����+j����?цlU40$sB�O Y>�����}�<� �����˕�F�gN��1 U`���O�P�sD̦��	D{�ctGL�x���Z_���iM� �D�0��ڟ�ϧW(��IC�$mU�9u�>�Zl��I\9 ~���I��O��6���H��a��ʎ4h��4�'�*a����S�? H�30��H.p����4�xq��"O6qAO],^��䱵�X�R
�	�OȌn�%x����	���P��@Zb�c�x�!Ő�M[��?QɟfT��'�@����).8��nT�~�v�'�b`[I���T>�12v�� �U+u�6�K��ǴW?z0�O�����)��EO�sv�K�9��L�=(��'���S������OA���l%*lR���0�h�'yz� ��Z0^�qx󥗎#�CÓX(����%m�(5.�}AөM�t��1 H���MK��?9��5�ecW�� �?����?)�����ǿ}�t|�k��Kb��B���+��'%Xc�3M*4P��J�p��9`�±!����=	�g�Ix��A �	6S�J!� LH�~6u�&M^�z6e�)�3��O��ZQ�#A�~��M�hF�s!���<TU�	C׭�9^g��4&V
k���HO>a�mEXdJ�`��_������L�q�� 柴�I���͓�u7�'gR9���Rr�'����H-���:�^�~�!�D��������
ett� �$^!iV�7O��N*`vE��n^�yf�3֥Υjy��'�|��.��)�@��30�R���'m��s��]�	D�����-2 �;�y;���EJI�ڴ�?��o>~��,�4j�Ҭ�e�Y�<�B����y��Ӫ�?��������/�?�M>a��ֽD�8I ����10���Bd�O8���0�I�=�:� s��
�U�䏑�a���̌z�|�'�~08XӁl�*=4�9ZsA-�y���,]C�a;��B�8��2&�
��xrbp�f�@�	�|Tv� �Ƃ�W��9��DϽ��o��E�D�?YQ͒�ncx�Aaؘ\ش�a���?���SX=������V� v�R�C^<0�j���С��I-O\#<�z -I�U1�	�Q��l�6�
���T�D\ 9����ɝZZd#WnT$��Pŉ�)�!�D�nJ|���l�%)	����axD3ғ8�MBtg2��$hDG�f���X���������K$&a�	ȟ�����&�L�&	,���%�H�G0�رc���]^�$�A�Ӛy�b�HF�g�<d2�ai�ob�9j�OJ��0tr%�W�@��5(�&��N�LP��	'�3���!6���+J���r�꟎*���*?q��O��8ړ,��$ �ВT�:��#��*����ȓ��i�#mQ��#�L��ǀ6?i��)�/O�Z�&�PC�al͵gLa�#F 3"�y�2�O��D�OB�Iֺ[��?Q�O�8Abș���o�$�����1KL!����.���ưp�.Q�d�^r<v��O ��4�N
0T�3E�
�k|�������'OE*�j
���u�ǔ�BXZ�'�긹5�ׅ2p<!P��d��8�y"6�	��f�ٴ�?���N-���*5(z�(�~�����y"k\!�?1����f���?)I>����U_�Q�Mh�P�&v8�`8��+�	P@�٢&Et�\�����m����d�-�|� �Czȭ�C$�9P�gJ��yRm2 p # 6}��=P����x��t�d���8z�t���M9���W�C���mZΟ��Ie�4A)�?���"#�
0��э����u�<�?1�k��m��ݘ�򙟄���12A��OG�[�(�7}�)���O�`��֓yΊ��0�$$r��>	C�ğh�<�*W&�7I��qc��8��ђp�HH�<�2�ǒi��BP'Gyt���O������9t��1�$ �3$L�aҨ�;7ܙm������0c�$;0�}��؟�	�<��x�L��\B�Z��D���<9�I
Vx��EjO�/$����?�h�u) �	E>|���vuq�R�p�P!B�>:D�c�,+���L>��(@�v�;��� 
-���5JMx�<�aI�!SRb���lʾ$6کa%o\t~®&�S�O�FI2�/۬N����!}��{VL�*���d�'&2�'��k�5�	˟Lͧ�r�
��θ^C��Y�G:l�8���r<14j�v�EWB�ft��l��s��ل��u�ipB���yh��E*92��B�e�ǟ��)� ~�1��J,@��q/���-I�"Oҁ�'�d�L�����0ʐ,�P�dMY����JC�iC��'Zd�ZO��3Z�us�O[3\����'��d�
w���'j�[�>R�|��^�b祙�K��B��p<�%�N�'-�hb����D��\h`D# ǮՄ�	����<��کV��u��5�d�VVn!��W�q�<2u舌����U!�52!�$��ytאl:кv���3�He��;�I�l�m��4�?�����޽oe�ě_i��)FAR:x�����V2J��'����'{1O�3?����2{��p��H 9�Q�K�䏊4$��?M����/k�������]0��-}a_;�?��y���O�6kO�-25���k��0�H��y��?AtX<��	� h�L��K��0<Y4�ɱ֖ɨЎÙo�h��Y�cӒ�ݴ�?����?Q�	�c�B,����?��y�;;���[F~��"�[4N�x���yRbV/��<i�QY������	�?R��
�A�<Ɣ��I�!����F�"Y���	�|�*��<��	��>�O��裊�t���S,���L�H�"O©���W'	�ԈH���	,�����T���S?i��3p!�8N� t�u�&$���? ಍�I�$�	�<9\w���'��I�b��Q��.p����ʜn��đ�O�50"K�(Uz �ʢ�սcF@iv"
$*�!�)Uj�e��#%�L�t�оX�n���'����,)h� 9#�����QDH�yb�K�I�ֽ���'!�����dD�<!2��� 9�n�\�I�:�PhP�gה)�*I��BL�VT���<���R柜�I�|j"��͟`&�l�Y:�<�)kQ�ReXh�+$O��3�� !�l����zx�Uy�B�O�x+�?�O>�D�QI���Ԅ�71
���ft�<�E@s�$]��׻#���R��W<a��i�|4b��+q��t8�f*?��#�yr(�6M�O���<����Ȫr
ɪ(6�<�,g�2,Pr	�,��'z����B�S��O�m�0�P!b<��ȃ̜�?�Z)��>�c��`���O��Y��J���^D�%��(ʽI������O,b��?e� D�4ft��OBYX$�c�a5D�����n&P�jJ�p��4�0O~�Dz�ɑ�P�Z�`T�pl8$�#M�7��O0���Ob�C��3XJ���O��$d��.Q�a�
\C����Jxa�`4Uc�dp�#<O��	����#|q��KM*/3�x�&��]�/0�y� �4%�qa���P)�Y���ͼ"1O�I����A����� ��,|ȓ"W��`�+�=��	���Z��'�v"=E��L	B#L�1��<-'~\c�[*y�DYzĒ��'�R;ON�]��I�|*�od?������-T��	5� ����GPJ��F�b�dEQ�C5�� qʌg<�AF�#P�$��B�ۥ���z|�-�	i��x#$��v=~�0��)E��I�C<D����{V�{���E8z����9��"��'�&��~���d�O�yIf�ĴKvH@rC++��Oh�Ʌ`&���O��%|��D"���a}�0�5�U�dD�=[��[�Ls�x��ۣ��'9*WA7\ȕ9��Z*
���ѭ?O�`!�'��'���fՔA�����I( ��(�'r^e���P"|	؉��J�&,X�U1�'��6M�Hu��BW)@��p�b��1O�ᠶ �����I�,�O�aB����$��J�Z�JG*7+�j��?�����?y�y*��	81Q�Mxq)	�/V�ZT!S�f��'L�S�����.�")y�0Y����H��c����P�S�'P#Z�PVY�,��r.:O�`��ȓ/��1#Q ��r\��7��OWQ���6�HO�}���;;��D�ϛ � ��v.�Ǧ���ܟ8��#7o�-ÀH������ǟx��߽�%�ޣ;^1#�%^�errmB�)�K�F����ɟ
�0��Aտ-�pT���U(3���@3�8<O�!����N}�L�E`A!_��<�af?� ]�����|�β���O�>uAhYuj	2�y
� l�!��R���0�KD�j�l������ ����7$���
�S,N티�߆�6�����([@��I��P���<�^w*��'4���ň���87�P���M�_8� 8�Ory�AҏU@�镏@#B�YKE'�vt!�ҎUUƘb䜬ͨp��"L����'M��o���
rgɮ8K���1c��y��M�6��gа�Fp��c�͘'6�c�<�����M����?�r�*���,�=�%�j2����?	F�Γ�?����d�Q�>��N>��-r�~�Q��řs��1) g\f8��f!�"�O��3fꞪ:�αi0,0a.|y��'�������?!���?f��&2ʸ@���T�%0>��oM%��D�O��"|��E;y� ���$g!�,��FGe<1�i���Þ��H	8�. +}����'J剁T�"E*�4�?����iҀow��$]"��R #�2F@��Oց.bF��O��P���Ofc��g~�F�883�	��Ƶ#�o�:��� ^�#<����%<R|8!,O����7�MK��X�2���N�Q���+"�: �Q@G@Ϫ?!�dΧs��#��F�x���RdQ�$ax2 !ғg��́'i��g���ꀧD�K�p�ȓ6�����A�=�D<iҥ�4(�6`�ȓ=�l:P@P(xZ�XS��E1*2��ȓ=_�qX�$΍&������z%���Y/,9�m�;Eҷ'�%0|���ȓU�����ȟ�Q*%��צ<E��Q?l���-d5��a���!dj��ȓ/��p��K�@�r!�`��/$�y����9�UL�����h++&�ȓ#���"+��x��5I���y�<���z�@���E2Gnʑ�Sn�JdTąȓ,��Xw^^	x7��K�B`����UÅ �ʨc��XB����j-s���e���kumƸG�����8��w��gd�H�'o���>)Av� Q���n��m�P|�ȓ5R4:��Ǳ?�0�����V�R�ȓuBj��s�S%���0Dk	��#'D�t	�k��P!�$�)&*J�{�3D���A�&zlYA�3k�dH�/D�,�VV��Tsv)J�gn8Za�.D�<�2���>����Ʌ:X���C0D��PdF�d���\��H|�do"D�|�'�w��) )�%kV�)rT�!D��!����}xP��A[�H#���2�=D�L+F�M�0OZ�KRhY�|�1�&D�3�/A�g;։8�&S&8""	��2D�Db�Ռf�.|�iݵ !�L�$I0D����ftHLГP��4�@��I#D��#l��P� ����Ӡw�0(5K-D��öG�-)�����B�4��-D�l)��*p�Z��9칛�b)D�0����|��e�
;n���$D�����``h��!$U�NnZ�g�%D�p
ؕ<�19�i �:9�5�?D��* ꊋn)Uҡ�ʡ2F����<D�p��U��	¥��l�$�j�9D��)��e�V�y�	Q �q��3D� �Ό�Fi�������(�)<D�X��	��o�@����
[�p���%D�<bI�> �A�l^����#D�|�AǤ��ᄭʚ��� V D��ٶ��a�Q��)F�K؎�t/*D�X(��7�m�O�<����b!.D�`�Q��^��I�Ȉ��ư)G�0T����ˀ�B�����!( �{"O� R@zƎ2U
���rt6p$�"O�-��Ñ8�:}sn�-!�ՙ�"O��Z��hv�͚Aˌ='�غ�"O�!Q���a�͙��9A��S�"OR8롨b�����,��,�7"O\y�B�W�5��\�'r�|��"O�U��冔_7p�j��,dR�}��"O��4��#4�K��*d�}��"OjѫD����%q�!�,w����"O��_eG�}����.�>l�T/z�<����	rq�̆)-�!���[�<�WJ�B�l�$��D1�`�W�<ن!J,�=�pMR<F�u�caCZ�<��� X�b��'o5~�H(���VU�<���\6WQ4�ز�Ŧ)"�L�g �g�<�G��F�X�)���?Dfׅ�Z�<y�I{i@q��|p��bT�X�<�ea��~���s���51$��+�j�<���3��dZ���0B�4 �bq�<9AI� �!�wHӫE:@���
ix���c���qI��G�0"���%.�Q�����x2�̛t��Y(_>=�(|@��	��hO�as&\�3I� ����aH�b��K&";~��k5��+�y��p,��:��� ���_4�?AGB��W�(-PP`.}��	�[i�"�@Ʃ<0pJ4�<�4C�	�:7��K&h�)[Xj�a��4m�ʓo�L9ੈ�
���D��G`Ah�Gz�av@�����;��0�	a�OR����y�C�*B�H���]�,�wOt�E��@�`��TKC�4r�f�'��II�J�I�j���4������1|�(%�
V�vM;V�'��` �i�v}r�� ���jC��E�fъ�MI��y��܎9�O?�P*�JM�� To��D��F6�I���肋��R�L�b���_�|� ·^k�xU)[ ���I܅I��}�!,O�����G52���Í��$�ٖi�	dhb�4�9�xU!�!ہx\iJE
Y�-����!L$���.ʹs����@P�t���'�8�r�('=%dD���[� #l��Ԏ/c�"P��JV4<���
4��e8�p� �?�}Z�O�l��Q�! 8bD�D+P]��XH���U�4˓lz~,�$g�4�r���ʻQ�Iˢ��2�I��#�ݟ�IM�Ţ ��'�~B4�ݏ6� A���.q���{�V�<�l�����Ï0T�D}�$��.��wԴ0b�S5	����CBZn�8{CE�p<a`�=h�}8Q�ʛ~�9�! ����Îy� ��|��hȧSը��䯊3Z��hbd��Tl~��c��s*���eֈQ��K��'���!"�WͲ�ʄ��ABj�����"h3U,ڊ�J� �FI�����E�����"�>�x����� hIw��2.;�����p�:	�'�z���G�3f��㦀��z��A��,/���ן�����nR�D�9�u���w���9I�V���M�oŮ]x�*�&��OJ�C$Y̓K�Z�Y�,	�3�0�&�[�2�`Ǎ3
�B������A#��v��4��i$~���Ľ4<f�b���5�&K��ƙ:R\�Cc7��ֹz�L�I�k�F)HX�`�d���aL
h� T�IC��@ʯY|:�¬���~2��p=�c���<'��y��U�P9�F�x�jɉ��Ω��D"GM�3�Թ�'玴r�M2��K}?�Y7���e�T- 2hJ�E�:���E[BrUQ��d+S-'�D�BtQ��s�#*v��1PE�D����Ø���	Ed~�!�z#��3g�ʓq�F��Ō�<��{2d��I˕%�'��0)L�\�Vu*r�ځ5��!J ��R�ʣ`L�f��Z���D�j�k�;�yr+Ϩb�6�2�T�3�z�I�����'�B���F��l�cf��^���(q?)�L``@�qK[*/ǈ���f�DQ�Q� ^�XyƬE��|ہ%��W01
�b���pWGۗ]�29yK�`��9��<�4|؇�Ob�[>I�6J��+�l�)`4�T�WgZ�^/�M�ȓp�vԲ��1~�2|q���>&�nh�e_+{��C#�7'Kl�`�柄t�f��4��|r��v���Әw���	�"�5t7b\�+�,���'l4�J�	�[x�8���]* ����@C�{R ��K��n/\D�(Y�[�4�o"{~p�rR� 8����7g�t�έ�0&��y�r��䗍Y���b]�QqD�`�G�>N�@�c@ҹk��4R�Ȃ�<�0�j�*ğ��v�I!!�a|BAUz�4�v'N'6� �6
А���^�.�� ��`�Ak����F�fR��9�V!Z2:�� ��K�怿l�5%ӡA�Ɛ��"O2<Qb������)��a�<5 #�#E�@��&F�b8`�J3�"�?�I1���I6z<:X�1�1�2��!�;�!��Q��M��kK�yp���q��	u�^�pE�;}&u؁�yWZ�RC�O�������OДڇ�L%������'+x����'לa)�\�O���[Ǐ���J��nǁrʘ����w���0GԄ�~��7l����u�`�8(��Q�g�@��'��4� ��c@�0��[�A���'}�`=@�p>9��G&t@U�+i4�h$�0D�@ ¡E.+ں��elJ���Sq�4@��層��?��$��gv0 �P�i���%VΡ���,���;��7t�B䉁e�*I�@mH�+�5C6��fZ0��mU��HS��x�@�Р���㴣 2O��4	g�.LO�p�W������W?Oz�%��@s^$�Չy�,��"OB����,:��P�5]^�	t��h�ޱ
r)�����X�b�݅.c������dK(P�"OdYH�,��gbd`��n�86��xEJ��$I��%� 	��,�g~Rប,��9 ��<h�P�L;�y" I+�f�����;Z��Ii%LM�	���gdFo��}B �	^j��s1��# 0�с7��0=s� U��'�vi@j_ z��i��Kq[2�	�'o�и�
+�p*ӣ��a���1�yҫ���O1��:уV@���"��S�l�b"O���;C��(�5	�L>��ҧ"ORU` �<g&�uvH�aC��"OR�p�KK�\�LM�&��_���!"O^(y3.I���M2�%C�X}�ӂ"O�$:3��6R� 7��\m����"O�} �ME3�Tԛ��ՋK^<�ӑ"O�ģ g҄{2L4s�O�]9"M�""O��ң�:o՞� V(�5�H:U"O��"1
�m�N$5��x�ޜ*�"O$:���9�f{�KB~�6y��"O�H�M��2&���A�V�2��9;�"O<q�ை;\�2��Ფ嚅,�5�y�f� ���9"	���_��y�+bf��0O�h��!fM��y�Β$�Xs��	)_��	G.��y2�2e�XxP!�����k��y��F�o�PѠݐZN��c"Ĕ3!��9:�$�8cOA�+C�Z��2'^!�D߯mI����d&(R�����p-!�$�6@��q����.p=�� XK!�DI�RY�}Ѓ�.YҲ�q�G�w�!��g���"'MI�҄Z�I��Q��:��㨟p��M� hBd�T�F$9ƌ�+"O���r?^]���ҳh�t��`�J�+��УU���O`�+C,�?l �I�!�>5x�q��d �6�f����ӷ-Nl�`�BH�ze�]�Ǌ�Z�H�	�J�k��'�l�[q �;y�D�`����Y�����W���O>����Cƍ(�\��&�Aa#ݪv�H`�r���q/����ġa�S�T�����5R��H�I�,�	�Nh}�D� q�b��d�Z�Q�  K���)��\�r��̆�	����j����<�6��D
1e(��oJ�TPu��N�<��b?`���šU�f�R�3 �A��x1c�C�>����,��fA�>ti�NR
K�Bձ�"O�U��A;f��$!��
�cF�aR�^'e�
�#��|��Qgc�����q�j��*�ॠ��9D� ��
\T�d6�V<yS��#�Ce���A$d�|��DЍL�����GD��y��t'!�
���$�ޣ[-�4�"I��3{!���Jه�C0<=��#��c����ȓR���І�W�^t"�nÁ~�\t��|��K�Ԋ)l�b�F"����	��ͫK�VKt`�&�ž!m�,��S�? �˲Θ����ߓ���@"O"��S�ٳ��i�bE(F"T¶"ON����L�4uH�����9h�1"O���]�m����1�${"\u"O8m�. !eR	�C�R�c@��XA"Oh�iG�Ī�0��0���a9��I�"O�d�T#T�v�	�#LS#�=pb"O(AJ�GZ& %*��P�0�E�A"O�8Зo͂c	f�r!E?Qʜ0g"Ox��m�(�x����_�Nm�'�`z7�ЊJ��]����m�:=��'����F6��x����F`��'˦=��^-��x����\�
�'���c�C6$�j��Û0 q�	�'0�aBR�K-�(4B�g�|�ܨ��'x(U��C%gwJ��@���Ƥ��'�As��Ġcm��* ����l��'V������R���0W銂μm��'br���BD�k�����'	<�|��'�:]�W!�-;�\�A�U�]��'��U��ț4zb$�B�d�L��'.F����
րY�	�V{$��'���0Rc�3M�-AkO�6]��'��M�S@�rnQ)�G�U9��s�'����@��h%�e�N�J���	�'�n}jU�;5�v��e�	�Iz\89�'rmx���vnC�ďy�A�'x���M�'o�X3�ʢq�8X;	�'�@(�M�I�1�w͒X~	��'��u�(HyC�Sgā�~�TY�'k$�r�DޜH%s��]�l���'����&M�b� �2�ĉb�\�'N<(�1ck*� 0"�%W."�'�����HT����D�-�
�'�
!s�K6��Yآ.C�6��
�'VEBT'�,IG��yq��Qw�r	�'�$�صmơ?� ���c��E����'E�L�@G޸@����Ɖw�$%��'V��
�(�R��9"��ij �`	�'�ڨp�����uPA�ޅ_-�Q�'��l���m(E�!.)P�H	�'�X5�s)s���j�m��Is�C	�'����lB�r*(3����@�6 ��'y�\�D��a42�Q�L�N�x�'9P��qj��V�~hR�ȗ�hA��'Od���H��C{�d/�%N�H��'�h�0�$ڑh��DY@7Fl 9Q�'g6,pV�1!��s �<>4�h�'}�(w'�'mvq�3. 2H���
�'�(Y�cT�j!�\���=m%ƽ�
�'���!&l
&M�Q
aK�Yp�	�'Q,�����#�l0�	�	�y�K�WU�$Qv�O�^G(i���M#�yR�G�\*PZT@P�Ywp��お�yb#�=z��go�JHX�R����y��ZK�V�;���-_v%�"�G��y��M��p��П'XM�&LS8�y�"o6���ָ?���EI��y�o�1j�B�iDi
�o��Ӹ�!�D&B���O��|	flr�ě�U!��@@E�G&[��(�⛭=!��� P�"D�d�t��GDc!�Hd��@4��&�`�� -I�!���>�ܘ�f �2~ܮ ��S��!�� ư�ÁC�XH�a�̒:r&��" "O�ˑ�E� `�|PA,W-&8ԩ"O
d�,�@�8A
̖J>�KQ"OH�R&��&�v�i�
����X)v"O�	�kD���xf#�p�q�Q�Ig����@!T����c����P���"�!�>i�.�@�I��
P��$�Â?[!�I$|���bi�hK�"��9"K!��M8"X| 3�ϧ5/L``��كf�!��/}ژ
UNG&`�$a�;x�!��G��y�g  D�㊛e�!�d�"1$5�[��z�/�*��
r"O�QK��F+o�j
3*����W"O@�{4L�,bQR��
Vw��sC"O����[?C��a'K�u�vA)�"Ojy"��9��t�$�^�o�r�"O�P:���*-�
�����w �8��"O���BˉUr�T�4)^<��m��"Ot�@$��(cOz�j��&MvX�"OD�@�1��:��L�� ��"OB��j�W�!r�'Q�xi��"OȈ)����]��h�E�]+��y�$�>a�D�*#`��+i�MQ®0�yB/�- �z��e�����`Re���y�GǠ���x��O*~�f�@���y�IC8"��up�䕙% ���q@�3�yr��\H+���	-5zġQ���y�	#> HT C���N5`�/&�y��dPj4�C�D�ݘ�x@����ybmC�G�4aׇ��T+7�"�yb��FL
0�6�E�8�4��K���y�K ����L�f��|�#�ߪ�yR.3l��kv�\ܤ"���y���$�0?��S�(��I�D�-j����a��P��>ɖ��81��:gn
w���q���V�<q��R�c�X`��d/r@\tq��}�'� A ç|��D���t�a(�..Ṅ�W줒"�׽�Z=
�a�F��� �I��H����5f�B$��B��T�3��?��B�I�:�����)~�%yv�U.C-��dG���;�F��oC@�H�"U<T ��m,\O2�6)��}D��}=jiJU��5.ʐx�P!e�P��o�����%K[��1�fG�,Zp�=!�0J�O�O�ZL�f�D̸i�d��bvt��	�'�>���� rh�,̉`j��3�n?�K&�>�'X� ���j��a��]�r�݆�6���-��o��Py�/�6;��i��aL�1�	C9:�iZ0�ֺb��ȓE�� ��`��	�8�q2���3�T��U�����G�so|���c��m�ȓTS�-BcO�,(����\����`N�@'@�6MX��bExApl�ʓV���F#�/!�����Q8h�B䉼D`mƏ�4��Ԩr���WڴC��c��<�Pb��3P���%ڒC䉐8-������
� +��=q�*C�I�"&��9�.[�|��P�\�f�JB��y��KG�ӑ%�����٤'�@B䉥�p|%C��&➜A�(��mP:B�I�-������Y1@chL�cJ�5�B�I�6oJ���@���\��7�W�`�>C�ɃR�P=��N�f�l� e�ԣ ��B�	"t����C&a�<�`��^Fu�C�Ƀ,�Tqފ<�,H��[:C�)� ��q����dʦ�E�|�@`C0"O����&���H���Ae �I��'���
�a`�O��CF=qL�5�!�?��#�
�9"�!�'M0&|!�D�'� ��oʀV�	Ѣ�GA�!�$�z,����%d�F-��KX��!�$[�����^�Z�\�;V�+�!�d�ʐ�9�(��!�|b`̾*�!��+N<��k޺r�R[7τ:!�dY�O��a�@+��P�<�ab;
!��e4Z���(׺T�T��,A�!�$E�#e� ����4X���eZ�z�!�D��D�4�vÒ�3� �C��*rJ!�M"��X5�͸?��Aì�
?!�D͗vT�8���P��2���`N��!�$�4T��B5+G���(pP⛛z�!�č6��1d;]�`���K��y�!��%h{�����R��YԤK;�!���D����΅�>�:�����M�!�$	A�P�E�@�0!i�g�!򄐛2��%����:�����Q� �!�D� t��)a�C	����VdȦ�!�D\.�Եq�E��y��`����{��Ш;j�h�E�C����qGW�y���`���h�"p�vT�@%�
�y2��V���k�	�4�-��yRN�3g�h��Lǔ"JX���H�yBF�IN̼�3(M�!6�y��#��y
�^`9�'�3#t��h���y�-�	�4X �X��@����yk�!�l�q0d
whԻF�H��y�g�
[��*��W�s���s��J��yb)�+R`�� ��suB	���W�yJ�.��M�D�M��>�3%I��y�X�j�F8˵%D;�� ۗ��yҭ�96�~�+G+߻����f�_$�y�I�pȬ �!����`)�d���y�$�kML%��� :0ׁJ��y2���|�:��s���G���W�Y9�y�2 f� �-��9X�Ӵ�yr��U����7b��5p�%��o���y�1M�� �ꆆ&�pXІmA�y�+W<~Zi;qV7]��S��'�y2��'f2̝� jY�}�BD�Å�y⩖!+5R��ť�t@,� R��y�*�1@`q��8m-��±��9�y�"i܌��PAúal�d�!�	�yrϙ)��5�ǦZ	�ԭ�a
�+�yr<"5JMb3�U�s<T�a��y
ԞNenh%��c�0,��H3�yr��	9���Ǆ)�� 1L���y����n|�C$I�(�ΰ�����y�oߍFN�R��HP�8|�'f���<���D��8Ͳ��5�rxC��T�!�d�8 �
���n"}�⩈��9!�.�
�Iud�*8&��s�šv�!�Dĉ+��P���ڴ*����f}!��.3#*��!k�	>���`c+�u�!�;���w����A‪��Py�Jw����t�H>;nR�qs���y�$��?ʹ��2i�>7����Q��y��' iұ�^�c����s"Л�y2i��`���V�(+�kvF�+�y2���,u��!��[%p��D@��
��y
� Z�뢊�2P��{C�F��$��f"O
%���P�2�:ӌ�8��@�"OT�)B�> 1���W�n�$��"O�!�פ*u��r�K�;t�"�{U"O���B�_�&W ��#"OL�Cwo�e��C�U�~�j$I�"O��0p�R
0H��k�>E��t�U"O����H]>	D����.���d"O� y�ٚdL2�p� I%wxY""O�r�9>�<@���`�m�G"O֕ uE�� �X�w��;�,d#g"O�4���O�	(r��W;-��)1"O�D�noN+X�c$2M�"O��P/Ǻr|��)0�΂C
��"OF\Y���&_���3oܔb#����"O���q$��-k��0u(J3�[e"O�����OV�^��5G�7q��x��"OX�����axy�e	%�<4�"Od��'�҉2&C�#� �i�"O��hɿM|t8�v!E�#�tܠp"O���.�����[�u�T��q"O�Y*4�E;T�N���
�ǖ �@"O�U0S/��<p���!�`�g"O~=�B�J-��H���a��)b�"O�Th3m�X�&��4�٫�0<�p"O� *����y&����F���5@�'9&����Q1��K�%E�?*�"�'*\LGH��u�Z,J�K��>�-#�'}���(A	��Q�� }
��
�'�T��MKȜ)�cG3	 i�	�'w�5�����r�|c,U�{���'X�p:��[���UjM<t�&�:�'{���DͲ$d� �L !ٙ�'�n��Ӧn����?#��%�	�'�<u2�B� c��`h��&(����'ih�j0c	بH���U- b*�1�'attaCꚱ ���	:i7@�(�'q�I�!�� 3hMz�`ФɊ�'o���ō�v|�C�R醝��'m��O
$vB���p���x)@�3	�'=Z�q�� p�rgDr�^M��'.����:����@S����'<����J�?�Y6�׏7�fY�'_ {�Y:�V431H�G�d��'f�uA�bѻhWbū�����d��	�'^nذ�[�{2�h���%���'ޘ��i6��a��N���p��'h~i2�h��iR`�U�w�t���'AH�Cdלw��d@�^p���
�'����֮�L��0�"헜x՘�
�'�]�-�6E2����K�e#�QC�'`*�0vJϭP+�Ա�`Y�Y����'4!3Aڲ6�)�.�E��0�'� 
��©5����O�O��3�'�����a��7Q�`��F��A
�'��4`��AϾ���u�p��'V��G��=�,S���i�k�'pzxpE�:m�x��ɧ�V��'M�[����[_dX2��7�2L��'_��D�*K�%bY�\����'�"m�1m��;ŊB1IQ?;d�Z�'�.����1k��J���1>����',V�Q�^�*<�U0��J�3��
�'|�AC6m�[0�����*'zH���� mk�O���@���6Av�SS"O��K�	TTR�F��E<�|8"O�Y
�*�,(�j�q �EX-y�"O�c�3K�^1��!VF��"O�В���N㜄�p�PӪ1)4"O�H��"ݣn�2ĹQ��~+:��`"Ob�#W �}��Q�c���!(�{�"O�5�S��5�fl�S�%fHW"O��XO�b��$Ir�0}��k"Ox	�Vjk.T�+9�x�"�"Oh3���Y��l E���i�"O�ppD�Y�P�Z�CF)�X�P"O~��0ɑ�h��s���7�*<��"O�H�Я�:a�v`LY�er�"O�+e�;/�T��dJ։k�D��"O��QN�'�A@V����`�G"O<�H ��=Ҙxs�g��`'"OT`�Q�f�Y�& �^<kr!���"~G,K� �0Oԋ7R;1>!��.W�!S�nsa�i@D"L�r�!��:5[�h�7�N�+.x\"����!��A/f�j�O7*��PaP�Ru!�Dbc4�a��D�+�0Q��Z�!���A��_�!tɈ�b٧*!�dë)�ĺ�L� ��A�%A�+j�!���(C6�t�� �]�c�Q�!�� �6Y��it$R{n�㡃ħR�!�$���xtB��%]��QB�)~!�d�c�� sn�t�ԭ�p`֯z!�d�V訝F/Yl�2l��Ɵnv!�"k*$�r�bאv�0��D�W!�dE#�l����XT4�h�ؔN�!� �>H�k)��5B$i�s$D�a�!�dQ�2���;ҋܝ?�\P��!�Y�^�M�f�?�$ݸBl[�1�!�d���Y��,��T[���_�!��%K�M�& �[4<���9o!�X�{���A�M?tv���	�o�!��F*�B:s'+It��7 �)!򄉙>R����'k�+@��K!���h-����l1�D�X�ɦP!�D0����A	{"p���W!!��?��ɛ򯚤if@�ZU�5T!�d�G�rt�ԋ�.<\�	p�؎p�!�d�R_���fo
�0vQ�A���!��
"���5OڭK ����L1=�!��<\7<LC!Y-bK�س�DˋQp!�_�`K��s�䤉�,�?:�!��˿b�`D��B�4�y���.0\!�d�2=��X��&]�
�7�
�YK!�:뫤ǱM�
9�b�$~_BȄȓD�>l�%��6e!~� ��L6A�j���t��q���>m>�Z�/V�� ��oj�� 'ǐawn���""t̲��ȓ�
}QKʍfV\}����Ή�����#�(��o�bj�yG�<�ȓ}U�P� �"B���#J�&��xr�1�@�$4h�"��<;�����jgJ���	�c�p�zv(�h�`�ȓ9�e�E)VD��Ì��L��ȓy�p1�q�R��2n�O8���ot��� ���tc�!��&��T�ȓ\
�	�!�N#�u�~@���?a�؁DD �Dq^�C�������S�? ����+ ��R$�cRpA3"O>�j"�<!��8���`��*"O q�]�԰pPȅ�#�p�!"O0�E#��Y��V'F=9$"O�m�GF<ҒD�C䔄;���4"O�eH�
�L��d�`B�0n�|���"O~=
E��&ZO�$q����J�Px�e"O���b�~�h���ǽW�`�p"O^DR��m����$�_�ܝ�3"O����
��Z�I�a��YZw"O��P$l(4�>��A�@�C����4"O� ��F��sM��i#Dތp)�1�"O:u�a.�t x��D�I�`�"O��@�BM')p�a�#D:�d@��"OȲ��M*��E�	Z�j.����"O�yQ�_� 㪭�DB-"�N�"O��"�BD��*Q;=s`��"O&�pU�R*i��6hCT"O�|�,�1��<�'�/�^8�"OL��ȫ�r�Y�@�̘��"O��Qvċ	������t�����"O���A�,�B5b�-�h�DJG"O�e9�C�?	��̹K1B���1�II�OL\I�N��Q,�ie�:c;Ʊ��'Ԟ� 	8=pD�e�i� A��'�XUoҘ�^,#
�1��Q��'�� �#L�6%�4K�2"nd�'��̣��X�F�Tk�DR�)e�q��'T�a�w+C	3�L)�Q��r!�M��'�`jd���|v`SqE�k�'����M�A�hҷOřN	�yI�'Uz����3R4`�GJ�*;�贺�'�X� ��k�
M8'
ɟJ�^��'�D���C��D9�F�B�L;"�Y�'���Ӕ�����q!��t���9�����#��?��(��(C<-�fE�%Fі5�u@9D����AP ,�iJ3*�x�"�A:D�ܸlQr���#E�F#=*ԑg�:D�����I�|�D���@����y�1�7D��Ȓ��v�j�+v�Ń�t@��4D��:ՉK�k����$�(<VY'&D� �M����C�_�f�:Q;T:���O*����5x4p��NO=C�b����>�*�O.��C)B���d��,ϰ|0�"O�TC�n�?�9٠(h���I�"O���Q��:vh��J�q�4�hu"O@����(.��x�d�?�p���"O%J�� e�ߊkp��'m1Op���EB^�z�#L2J5)���#�S��
3t�\�s�� Z�*d	}�OP�=��l@ ��/%���g�JA*�`ؓ�|��'�إ�-]K�J�)�-� Z8��
�'͚��BC����T��Նr<8p�'	�m��/E<��)R���+y���'�{�С��E)f
�(�t��'׆-�ec�\}�k3aG,DE.Dx�"O��!��s%����`P�=R�a&"O�L���Y&d=RS
Ӹxs\�`��*LOpI�s�Oy�JE$G'kL �!�"OD����V��7��!=,}�"O����Gԭf=��b�:�t"O�8�BK(Q��]��7�Fذ"O���mƨv?�a2�KJ�\�&�[&P��E{�O�1O��E���<��e��
��`y'"O� ʥA�i��"
�-+�ƐE�p�Y�\��D{��I*��Kԇ�nyb,�6��V�!�Ȟ6��R�Y�yLp@��:I�!��@�	0��0��Uf�y"虪K�!��# �fBp��5o��yǡ��o�!��2?�:y��5@,I�qjA�!�D���t������0+�n�=S�!�X��8��Q�	�f���ǇY^�!�&R�B��"�YDv������"�!�N4��s�B;ce���ϖW�!���T��RKT"d4|�Q��6�!��+s���a�d�>]�C� (�!�d̠iD0��O0ĸ�/.�!��(e2T9hWC�)Gs����J�!򤟽Z��Z� 
��>�Sw,O�U�!��|��qpc��F�y;tb�5Z�!��4"X��%MG�Y5�y�~�4݇ȓ+�d��.7�
����ܕ2��ȓBT�Q��04X�u(Fh�>1��ȓ3�Z�h��Cy.`]����;�`1��_!z��q�H:6켅:1�V6�H�ȓ+6�0���\.^��iV�]N���w<�E�8'�13҉�]:�@��q�<Y@i�N���c�_k�Hx�Oq�<�p�$.� ��qY%jC��S0��b�<�AW�?<ڠ��O�63А���%�^x���'�j4oO�F)Jm2��Z�mX���'B�����j�8���+ sQ����x��άW0�Ԋ�CO0/�h�U�X��(�S�OO�����î}�@!��H�P�����'��5�CD>* �P��'^���ь �?F����T�)�bU�
�'��a�e��.ވm{ A��p|���' �\�n�?i��R�d	�Q�~��	�'�pp��iD�IAX|�W�^6O�=�	�'����seS��`'hݜT�����'ڐ�vC�:�Zm �$�/Tꨴa�'�ި��n�*!���ꛚF����'`��a���4�d�3Wi!
&�m��'���4�/Z�H��f�ڏ PI��9��h�rN�hd�:6���jP���`�|r�)�S�,d�#g��<��Ѐi��r�lC䉹2�v�+gV�RhM�cL݀�2C�I�^U.���E>(|qS�
��c�"C�I)	�:Dف
�5I���S��m�C䉸<v��]o��2�J�+#C�I!x�Ѷ��J�����juC�ɸFI��	5�����j�E-��d�ȓl~� ��	(�zar�C(w��d��;o���a*�85J��N0,3�Q�ȓSr��0��$4���G�x0ф�$�P�����`����Ao	���؅�V �\(n��q�ʉ.�D̅ȓ!���'�a-�&�0���	6�y�"�$&�!Wl�g�I�C����x2�p��Av�P'?��8vɖ_��S�$$�"~��_RV�2&���G_��g��yrh�	Sw��cmFn�:���`P��y��
l�85{4i�`!0 3d(F	�yRL��1���Y�bJ�-Uz̲��y��A?IӤ=�a�F#���3�K,�y��eu*eSp�Ö�=:V��yҪ�<�q2�U�?�Q3��[�y+׸B�L;���`䔡3�)	���hOq�� �0���l���`��e1FE�"O� �a/��V<���!J��"O
1��CO&���S���"O�����l���{5l�%�)W"O���p��0�.�ԛ.�r�bE�'���I���"ʶ��h�?^e�I)�O����ehAN\�f��uؒ)6dߴT�ȓ���9VP�'��PX���5*ub��ȓ���#��_3�R�Cć0l �͇�2�F��1��	Ae�	D���t�<��ȓeL��X)�/���@� (9�z��ȓ<}(�P�̍#q�2bjF�(8P���	y���.�QAo��pp�2�.�h��(����<�V��Q�����Zʈp��f��<q�!]�m� p��GRE����V�<)A�d����K�,�^H�qF�\�<!"d4�%���"þ�U,Ho�<F�**�5��`�?Yx�ZB�	m�<y&e��i�fP���o�lsw��N�'?��,�"$:0X5��։;�%�O:��!�6}��MO�S�:|��m�8�DB䉻-z����P,Y�{���'l�8B䉺#�6�K���	k�i�W�P���C��5Sd5�"h�_��ɠa.ЊD��C䉱M5��r�XhE�u˦��
L�C�	":�I�g"ˡ[��%� ��x�C�?wP�x��J$��x���("��C�	XvE
�f�� �0qP7�G���C�	}s��BͦRq��C�C�P|�B�ɖeA Ш��Q�%iʔ��`��+G�B�VV�����]��ĚG��?3�C�	�a[��v$�&H�^ �-���C�	3w��XAF���46�C�2i�Q���?qqBH�����D!T��Ђ�A7i��,�d è �.��ȓo��$q��M�b��a!զw踄ȓɜE��Ƕz^v��'�R���Q�ȓGCȰ�SA�=L�eƥ;l"j͇ȓ�l�E�
O�����}*F��ȓvX�0�����d{�M���� �Ɠ*Ӑla�
P�,J��{�	�+s�ͨ(Ov���*s�j��6�Ā7 1�֟2c!���W$J�+d�9����&�8l�B�ɀ	d�T�*ٴ")t�i����B�Ɍe�H�e�#K�Z��X�#b�C�I�o'N�ɰc���XC�i�f��B�=�������?8��{&!U�M����"�'��F��Q"%x�kӺf#v��D;�	�r�ȝ�
�+|�RPI oք%K��T��ɩu�#��26�ġы òB��<~4]R�`��M��0'm��MժB�	��t��^�9�VE��f
?j�B䉺n'�m�N:N�L�1�G�kp�B�	g���B�o�$�p��#b�:@C䉏D䒤�'h�"I�	?d?�B�S�m2�̥�8��AE�)��B䉀Y�dir6�Revb��!%�xC�	�A�$�!2��+\��tĀ+<C�����cDN氁&kGyHB�9)q.\Gɂ�F�x�Q.U
X�(B䉖W���%F47�P��O�-�B�I�h�`ܲ��?���S��$ �B�I¨�tL� gz�r F�wj:�h��Ip5d���9�yxт2d�C�)� �1@��$W5L���?<�i	"O<�CԦǈK��e3�+r3H���/��;�SܧHOD�
��мNY�!c ���T�Z�&��=�i(`�� ��ȓ ��l)�E�

�	�+��
Z����Pizt�$��4%��86eJC�pl�ȓHW,9� i�'8�XEk�PI*T�� ��(���>+Ԑ�J�'WE��%�ȓ!*�7聰*�vd�	�rP���i�'�h�s3�T�\7ht�c���"�\\��'�|�T�.u=�(3���TN;�'c�� �#��|J�kȩW���'�j�*���?v��Ȓ�B���s�'�-�S��	L8���!
��;1��Y
�'��j�_�Qł��'�~��C
�'����ĆNp����}P��B���0� �
W��.^�2Ə˿�앓�"O�p83
J��dtS�鎘qeؽ�"OY���J�ӆ�[&
���C�"O^5��Y�T��m�b�mѤ���"O(єH,#�	�@��o�$�k�"OB!Y��.X�dc6H�9;�"Ov�b�	�)Zb1ض'�<c	��"O����>w���&V	16�'�ў"~�&�v��A �G9"��]�`
�y�o;O@���k�d�H�7	��yBT� 9v���,��~��R�y�`N�bX�$B3Ν0�0��o,�y�(��D��t��G�1~�pR�o��ygJ�64I�E$v� #% 	��yB���@� 5��E��Z4�=������yrc�+Bn
<@�E�'C@8a���yB��.?��% A���0ؒ�	���?a�'���Q/��j�3@MԬ�:���'��@!�I��,j���G��	h����'�I���3lWS�r�Ll��'aNu*Z-��u���l5��'srdI��?R��m��,�-[X9��'�@]�!	�䬻K���ZQR�'dU�p��7j��p -�6aNt\���<��Eʳ��^���'Ǖ{�����"O~�h�ww��c�Pv�)�"Oؚ��H�Z=�(0U��KM����"O�q�b�Z�d^t1;�gW(N;��V��D{��iWZ��a&eM�OU����EK`ў����=�x��$ c�x�fI�|ɬB��5Fe�3�Jh��}a����.W�B�j�fH����&c>��͋�8�⟐��I�W�$ �D�"GTd��5C�B䉜gƲ��s�nJp07	Ǽ$B�	�u D�6?�P,���""��D)�S�O"�m#��k�>�Se�Ø|t|0Q�"O����R�H<���J%cJeI7"O��T��=�����̊I�`\C��@>�*�̈	fS�����[�-8����/D��z���>N➔h�nݓYH�{��9D���N��K����\���uN2T��Q�o�<u(&�*l 94K�"O\�`M$e�AX���	��g�'G�	/}�D��!��G7D���+�jC�ɗi���k'D�6zEz���Ŗ�7�����q� Bo��	��
e��9KJ�ъ*D�a&C�u�F��4K���a$�*D��y��rE
	�B瀦<#V�4D�� &Y��hY�`9n ����M_�E�6"O�m��.
�:D�A*,@���"O�L��a��iU̅hC�,P��yV"O�9�4�؀��
ŉ=\Q�h@"O��c���d=n ���+gDr`s�"ON��4�ܬa�܌��%�CA��ҧ"O�TzU �<}�`ѱ[�3���"OMل�.
�&���D!-��C�"O�8��ۢ^$�bO֠��q��|��)6H6�׈M�<��u+���0*B�(g�z ГN�)J���iCa] >�C��J�4��Q7I~����Z�s6�C��&� �Ss%.\���pvK��$��C�����#����r9�E��RN�C�	�5�2�rg��{��9)�B6xC䉚���B+��		DN+�T�O���dG>J❫�L;��h�o
<+�!�H�� ��#
�W�p2U.��Ai�y�	�H�ɩd�A*�biyaΈ]��B�I�N�Z@i��)R.� RO	Os\B䉪!������ȍd�N 9��i�B�[�k�!Y�yx8DH5Ç	V�C䉷-� �(R.N#2�h��Ŷ%OB䉣C��`q�cR*����]�C�Ij�:�CN	QF��#m�4r��C䉒A d�zP�$� @K j	�X �B�c
����dƒ>�8���FF2f�B�Ɍ^Mn����T��`��,�W�0B�1}5n!�"U���qǯqB�I	/��a���ga��j8�C� 9{tM��	0b�r`���(��C�ɔM2��X񮇾v]`<�ᦈ�w�B�ɔ.��)����8��h�&�zLlC��5���)UY=n
�dr�&��B�I%M����+�o�z�A���I<�C��8�D�c�(�hHp@���C�	<\a��%��Y��(C�FP'^C�?$0��H�s����L���B䉾�	2$�_�C��D��D�1pR�C�	����	vH�Nd�4�5l�*J�nC�Ʌ�6b�$�,i ��U��{�B䉄P�&賁@��@�Je���@�:C�8*�*Q	��8;�2���Me:�8F{J?9�%�6m�ha���eDT�٢�=D�D� Q�P���!� !$ P��:D�� ����! �4K�ꆟZj��':D�d !C<-P��5�'Y�,��f��O�C�	;Rx�	���*(R���E;H�VC�ɩ@9Da��j�6 9��8R�P�t�C��>,9Q�h��L9x8[�`Q�c"OV1��].�TE�䀓�RԡV"O���۬M�գǏ�0xy"OΜ��/��t�&��ő�:�H��"Oܨ�����4�0L�
���s�"O��F[e~  ���H���<#T"OJHZ�]�j`BI�c�L��"O���#�9D�Y�d^�Y"���r"O��J4��tH&��C�G	�tQq�'�4E�\ .L����M��H0."D�8r׀��7�Y�fҍF�H�Y5* ړ�0|��fӔh����LE��۠B�e�<��o�o%詛��0�h)q�@�]�<�g�<a���QPi_vLH<xtQ�<��$�FV\= �� �x�W�L��hO�g�? fx���#��̂A'�Z4xd "O��S��3E��R��?3Z��1"O��yF�#T�L����y�h{D�'��T� ��*nŚ�MY�Uб�?D����������;B��+� �,9D���@�V%�5 ���l��e��6D��Z$�&��K��fGz�Sf�4D�l���ۿm]��V�7o|M�3D��T�I*�.����͆%�vy��+/D��{c�X�""L�$�K�/>B��S�+D�<��B�H��	�*@er�g$D��x�Ǣ<�` ��KB�y�fH�� D�XP4��W&|8���?���@ D���'CZ%�=`.D�T&8D���D���n���+ro��J�&:F5D����AL�pH8 �!΀~k�y��)2D�Xj�ܻdf��:�*�*,j"�[ǉ"D��f):	f�aQÐ>�塶	 D���ga��f�`��C��FLa1�+<D���\+W똠K6F�{3J��1�9D�L#Q薉�N S7+�-E�29 ��<D���bCсZ��x6L���#)-D�P����r�1�� &��v6D�h��L�`��!*P�an��뀮'D�� �BSR��؇&N�A����#D�@B�'>|�س�b$6�y�"� D�P"҈�������b�&���*� D�< �	T�8�"Ά�H�qS�>D��r��C�C�~�h�32Azh
e�&D����� r<<R6�F����$�$D��4��pP�(�3Ue�Ъ&�O"�v5hP����V�����*�7J�ȓd�l��Cb̆xb6}�uaX�{Ȑ�ȓeJL��E�+.��l�eϬ�܅ȓ~"`Jh��f�iz�h��`�'��*a��#f�t�Ke��~zD��'��H��B� �, ���x���B�'�Ą���+��4 ���Czf����%��$9&��-��eD�!v��"OV "S��1:eBFV� M|�k�"O�9����C^=�"�B��JT"Oz|HG�չg⠀�&��+K�1a�"O���7)�N=b"��P�8$pD"O2����D-��#���~e�"O�غ���U��`�wh�,a����"O�!q#_s�{�ݻ5�J���"O�QqΙ$�p�;�NŇE�@�٦"O���N6Z�	j��
>�Nu��"O���ro
$P�|X���]�y����"OfP`�� ����Ԍ� x
l�d"O°s���O���f�
a�yX�"O�Y��� � �ㅅ̏CV��B2"O�3d����B4$T�Q=��"O(��2�ږr��Z��a�
��q"OZ8a竇�
㆕���M���Ё"O08�Aњ1�;q�W"*�Z���"O� 3�
"t�����R�)��e��"O���I���ӮDWި��"O�-qC�N�l��Y��'8��#"O� H*۟T�0p��Pt��x�"O^ȩU�ՁV!@$`'ٹ�k "O I�" <�:G��"D�ȵ�"O�9YJ����-��@�[�H� "O.d�Qb����d�_�*ǌ�J��'s!�� �����$��V�ɓk���j7"O2ѡP�7.yF��ФܞV�L�g"O>���(xp��ȸn��{�"O,�Js�^	B�}��E9Y""O.YyRO�g�4ЁM�q��-��"O,��艰\d`bL��g�@	��V�D{��	WgE�QJ��T�(�$��U&\�e!�$ފ b	s
�9e�S��R�P�!���x�΅���QU"�"#�58�!��ҒzF�as� �'K�TA��Y�=�!��!E|��q��`���$��!�D�;H�X�����*��#\�!�$��5E`�HWeV�,r�r��ө Y!�dЎ+P��&'ڹJf�8���8-$!�$�0h[�!�B��0@aXt�J_�!��'N� DW8\d���֫�!��{�x���I�rKp��$�K�V�!��\!}�X��V�5LS��Ak;P+!�dM'W�Zг&/Z2�rԁQӼ~�!��K�M��H��$?�
8!�K��!�L+a"�0��&�|�y��ޒ5�!�d�t�h��͖(lӒH�$�=P�!�䅆N��@��ٺv���%J��!�D
�^��f��o#R�I ��'xx!��	�0w��� αrd��v��&)!��p7�U��JUl��0�l�t�!���{�8�8���3�~���N��o�!�DÊ� ��⍛I���5��ў ��a��ܹ��'m����u愕<��B䉖a|m@և�'�24�ЉA��C�����VCZ�J�\�z��^+vC��4�~���� � �����B䉐 ��d�K=m�e1�(%p�C�&y~�0��hN6g� i���Z�C�	�k�~����m�m�B���O���O�˓�0|zC���	��J�懚F�P�X�N�ly��'V�ո%g�H�4Y���A��!�'hP5��oі��z"ͽ@�J��
�'���d��y$��ɛ�*����'�&p/��XBU�ʤN	JpYנ|�<�A���5Z��Z��Dy��q�IBy��O�� "3L�X�����940b,xJ>��:QF��F�)Ex� #cBD�s����'�a~2�W1� 7,� S	 T���0�hO���>|�D�T*˚j����	l�!�D�Gb��Q� ��>����#�n�!�?-��e�R�>��HkA_�@�!��E\�i��������#T�!�$�$�f �����sꞒc��'�a|뒼P�b)U͙.]uЩ�T�V!�yB�3o��<�T'��Kbf�$4�y��R՜�@��Q0 f=A׭��y"���
h��&�"~ �K�e���y"�Z gL,�G��6�Xع`¶�yfW;	 �=��8���ׅƤ�y�B�hz��p��3~�)ҶM��y" T�K��|���Q���Ȗ� ��y��$48���?{�����,	��y"� �j�X���	mN����@�3�y�E:|�FT�D���S&Bq���y��O�T`p���0R4�(��3�y��)'
D����	op���yRmH�;O(�ub�DL\XDT�y�@���]��
[�)˶��B�9���0>� |��3�&,��
�.�!
\H%06�'�ў"~����0]��
�0<jPHJ�e��y�kĿN��LRd�I;���#��M�y��k$}��
�C��#&Eۉ�y"˂	y��)2$"Ѵ;� q)�I���y"EZ {hs�a�f� ��*G��y"�ʂܑa钩F��H��(�	�?���al��� ɻvl�Y[���37*V��	t�'2.���f?F��R�X�P�����'� �z2�N�O�^McmK�J i�'�&�3���A&�ir�@�H���B�'��B1�@�M�Xx� ֡PI���'ў�|Z�S:co>��b׿t��Ti�Y��0=y��֭Gjڔ"�]2�$���%�R�<q�o�-	V�J��]�j���X�<A��*G5��N?t�h�)����<Q��W��ܺv�� aFxQǅe�<iE���UK\�QpJ�
x}C���^�<��+Bv���I��Ns֤��"O�q1"��(7)�PP���?AH�T"O�	xCa	
e',)��)&Z��a��'���=��t0Ū̘l�F	�`�Щ'\!�q�(tp�n��c�j9!c�3oP!��i�0�k�$X��l{���[E!�d�_;Vݹ5�֕}�N��5i_f8!��V��m�t�I�mpdI ��ډ$!򤅕.'�<rG	�`Y� Qƭ�"�!�D*'J��A�
�XP~E��-�)?e!�D�� ���W�6����XE!�D��,���0*V�F7�`��� �!���trT�ӌγa%���bL�
B�!��r%y�)�X�D��U�K�܍��/���!�]�V[ƴ;L�vh ��>z�0��70���3�,
%l�`�����1�)4z��r�hn"��tʐ�Am����qD�$���$���?���i�BWYJF*g�`d'�H"O4�!cc�f�r��`C�9k�`�d"O���gڔU�J�sO݉L��"Oia�H���:cc��!3�\��"Op��#.�83��t��¬)�f"O�AئnM�C��b7�����'=����Es$"Y# �u$��B��d&?A�i�:�m���	-��҅!�H�<1Q���z��0��bV-0�!D��R��F,39�1h��n�Aլ:D��#� ��Q@j�j?F�����+7D�ܹ��(C���@��Y��9� #D����Ӻy�\8QkR� ����L"<O"<�T,�&Gw�T�� �X��L�mD�<�Ė�.���(qJإZ��b��|�<b�Z1%"���u�b���`�e�{�<����>	�)i�K�s������t�<1qOE-{��蛄j\�5Iҝ(��Os�<+H#iF��"��H<��](%lXw�<�$DC�N��z�,���0��
j�<��j�G^"9r,�(b�`y/�b�<Y�-àA; �B��>R����\�<��*^m�*h�.B�T΢�%�]�<QS'�X~��2�$	V[�x��Y�<��D�S����X/[��k� @R�<i ̞j��4{4�L�z{2��E�N�<YP��o�>A�!��g��=�V�]I���$�0��΍N�Z��Aw�q��K��hO���� �U���0|/��B2��4KBuÒ"O�`鵩@�7��Y��)��H�"O�	aR)q�*lJ�IЏ,�~�L1D����\�(s���E��8d�Qu/2D��JУς7�j�n^<<` �V�-D�L�ƱH��CX%wo�2Rn�O:�=E�#��y_����2Қ<{F�iP!�D��-�H�t�^
R�|�S��N;{0!��
�KcJt�@DN�6h�	��:J
!�D��Hy��Y�j_r����M<[!�� �R��hh҉ܸU�z�o�5B<!��;X�`@��/:��)��{��O�o 2�k��ԆzG$l� J/!��B�מl��� .l Zգ֦#�}┟p�c��7܍��Ō/�D��S� D��؅B�b}1��ϸ�
hy�O2D���#h�5�r�;� ��||�	{�6D�X�Ԇ#P[B��덺a��1xqM5D�h�I�
m�Ъ�L�d��	���8ړ�0|���H�<6�\Q��I=j�s�a�m�<�R��%�!kF�I����PK�D�<�A@@�
�r��5
�΄;��[y�<��������1i�x��J\�<A�iӰ7��{��Qn$pG�_�<Qp��C���J4�ʔ;�`����u�<��,��x�acF�u8,H��f��x���O¾)#���28��@"	�|��Z-OP���k��Dy�̈́�?©���A�!��\%t�,u	�dH@Za����~l!�D>b5���^6.X8��%S!�䗧=Ib�q�D�rV�ٚ�`
"fL!�$�4�<��t٢
��(P6�51b!�$���P�d�&�����OW?!��Z��
�F)
�������r��'�a|����9F�p���0=s�ݙ��[7�y�!̺H��iIT��?
�����EO3�y�a�� O���EL�|�@�cS��y2"'Q��`"�IRr����(�yR�V�B��j3���>�$|�!m��y�♨#�8�ؕ�		t��"��X���D�O���7�)��b�"Ƞ��S)} ����W�8ڒO��&�t͓>��x[�%�3[&� C��z�H��Ug��Y&M�p���KЃS=5�JU��x�%jrz�L�GCA54 ��ȓ2ZP9cS�u `df�F��A�ȓ;"���F���F�
�� �l��ȓ%<c��D��	��S91H��ȓsk"���Cw����H�o�`��ȓ3��!ڵ��9�x��Gb�Lx֐��4���6�İl��Z���,2��ȓ���pr(�P�N��v#��f���u���h��N9'VU���Ã\�E��r�v4�&-��g���ABC��K��ń�WfΔ���Qw�P	g�=bRy�ȓ"�L�e*��Y���Iէ�.]xd��-���PWcO4cz\�S��9=e�U��������*l��%�H�X��Ն�	��qOFc9�hS�A�� \��?��q��N=Z�~	��^ ��x��E���D�B�����ǘ#��ЄȓH�tl�6��/��=)�
ư��9�ȓE�M�v):b���t��*&kن�2^i[�D)��AA�RW����uU���bgB�7���Y���E��S�? �4�TN��%� �"���s�\ɹR"OR����j�X�F�#P�ތ�5"O"�J��u�I�g��{`2���"OpD��E���I���yY��"Ozq�qMM�!�LQ����_B��:�"O��,M�`WP�C���78��i"O�|�H@2^����^�p2v��"O��`�!��0��0��M��p[�"O�$J�I
x���c�'����"OAՂ�1Nbl�b�:i�>Eku"O�"-��v�T�'�(q��� "OJi ��O4s�X�"�V ��@��"O2�S��v~�j�蘜aՌ�YD"O^))�
'G*�0���5�Py��"OJ	��N_5�|��f�E�PCH�'"O�$���<o�&�i�̆�&>�Hpe"O��i��t�r塛�V@N�b&"O,#���l�2�{��R7Q*bٲ"OTݪ�n�T��h+� �(��""O�԰��Q�aC����LЩ:��Q�"O�����ը7����
,�n���"OZx"�[5�fejE��P\l�0"O�؛b+[�|I�A�(]j"P��"O��i5�®Kz�(�)-�Ks"O�!`�A��qX��(� ���x	�'�*��!CҚ#�9�4�/�@�`�'���JB�O?>��40�S�y�'����SK)K\	
���p(���'T���I�N�$�;��;h���
�'_L�2�łx-BM1�*?u�*�
�'X���!�| �LK��k�"���'�6�p�ݡ}��i��*{�D�i�'W��x�d
���������J�'��	3I�[_z�1�A� �T��'ΰ��βc�4�v��7|�r��	�'e�����ۿ-߈<�u��L�]I	�'&h���h�h������f�8	�'o�0#  Q?��ٓ����6��'o }����}��3
W��H���'��#1��x^� ��5����'(�i���1���K��fl��'� D��f\=!B$��i�CZy��'�hPK�d�2Y���BK�8� �3
�'�ֹj%ݵ7y�kb-�cR2�)�'�♒��18]L4��RV����'�l���3tix����%��'�l[qhB8oQB��C���n�	�'�X�d�|�a�.���0AK�'���[�.ۃp�4E�J�5:�i��'ut���ID���ⷃ1;��D8�'�-Е���-u�8jgh?���R�'�����Dne2�
��O~^R���'#b`��
DT�QL�t�Z=��'��br-J�����`��8 >m��'el\0s��?��aH��͉%m�d�'�������x 6�r͏�#�B$��'v<�'����u8ҢK?����'B�۔�zL*�(i��(�r�'�,�y���(FR�zOW��)H�'��Qq7�_��]�C`W]�����'����C��\��̘��j�(e��'�R ��Q�*�K�iX�^�L�'�niJ�j &b����T�8llS�'A�5���P	 M���J�줳��� ��)�Ꚏ[r�q�ũ��d��Z�"O�,��Fw9r!�����+�h�4"OʬӅ돠G����m��u���{$"Oڰ�Ԉ��_Bd`G�i��e��"Ol	�FQ�~-�u��J!U`9�"Ob��1L��݈����S��4�2"O�80��c��P�U�߉-x����"O�yb��G6l9-#��}r>��""O�x �+AZ(�ba%�O�5#a"O���D�J�tк�i�V	>��"OZ��l��q�x����Y��"O�h����4m>���e�؂Y�b�Q"Op:C��4�p��U�ُ.�tPA"O<�2`� v(���B+C��p�"O�̢Ģ֤&x��u�܎>�̱qV"O��xՅ��&���C�EC.�j�"O����Eͮ%V\�A!���be"O�B��¹8͎�#rdß@v�s"O�૔�� Yz$@��
�6q(�"O�� k�	^D�g��;[p���6"O©2�iR��0�p[y�B�"Oܵ;E�֧Z��݈�3x�l�"O�rDɝ&�1Q�(-k~y2q"O�L�E��.-� A۲�2S�Qe"OL�נ�R�P�8��I�"O�{e
��$�m���!?�2�5"O&%�K̸}i����P'v��hr�"Ot��/eP��x�[�HƄ��"OƤ�t�H�(Č@�,�,ա�"Ox��@�E�S��up��Q.d�0!��"O�,�`�� a����A!��g"OH@v���R�iV�B��@:�"O�s'F��]�p�  ҰP�v52S"OV�+�L�9N贩$ �e����C"O�q�r+�"_�^�����9G f���"O,�इ�aX��bt��	{ r"�"O2M��Yb��"7� �w"O(#� T�0ذ5qק̙ �B1��"OZ���"[m*t Q��E���""OX��%_�t��e)v�� m�d�F"O��6�y�Vʴ�����"�"Od��Ìدj�iy�LS
.�>�c""OĘ�ELt�;d�L�s�v=��"O���Щ
�k�hy1!��{���	3"O�< �B
�npk[1#��!��"O������Ip���Mk�"O�xև@�b�T�X5ㇻ�``9"O2�	��\�I7 ���B�0E���"O�Q�A��^h�ъc�˿U�=�"Op����2����&�Lɋ#"O�A�&�ݎ8���U/؀��"OZQ	�g�%��2 @�M^6\�!��D
R�.���)��u��yY1f��`$!��K�O�|���3��,���F�I!�T!0�Tq��܀S�v�Q�
44	!�$ �:�I��Q3yw �����!��C���dMԕA[F�ӧi�G!�$0K�8��Ϙr<�)c'�L�J�!�DQl�S6@4ܘH�� ;�!򤎁T��A��ñf�:��O-�!�9�~�`F�u��MǍR��!�ߡZҐ	��`�Ϙ`�$*òX�!�d�r#�CS附+��lSE��.I�!��6�*țrl��<�r�[�j�c�!�� 4�g��>�Ȅ�1FΤZ"O�Dд��<ɺ���ȳ&�di�"Oz���%�,�>�8ׄ�w�z	��"O��`�iW$+�|�)s�ؽ~L~4��"O(9���Z=L�j,��#�� i�a"O�ȑH��i�n 2��;wZXx��"O��#)L�~�q)��72K���5"Ol((��	�&�1CA-�>'8t%��"O��ӕ*�%Ò�c���4n1�A"O:�S�j*�B�.-6$���bH�p�<�Ԯ",0��j��)f5��/�ny��)�'=�~u�*E=j�	o�w08��ȓ�hd�kص2n�$��*�y��N�p�:��֭*��� ��Ȕrv���{�^�sS͐6 �(��B�'�d�'����)�Y������c��A'��/��ЫCm<D����ߵD%��� E [L���R�'l���=� �ns�顆ɘ
4�0y�k�o�<Y�B�&�@�'� 6��yc�R�<�5��ژ�ش��Od�5;�i�L�<�b` �<�)εt	��##�T�<Q��@�B�%���O�*��;A,Rwy��'7x��ak�� q�|����r���@��6�':ш�R��߾t��l0�
X?�NŇ�v>��H��d�s!K? ~�]�'-�'��)�'n�4��7��x�E���X�$�݆ȓv��y�m�9W��mcGV�m��h�ȓo�©Y#�!	�F� �Ý=[�bD�ȓw�h��Ҧ�.q�� 3O���'��	�<��}J~"��A\Qrܠ��t��j�BX���O\m	G��>~f�Ӂʅ5C��:0"O�tt�կ[�J�ya
��y%��[���t�O�ZA�'�R�xWz�����&�4|��',���C��u��EBԪ�6]z-��'N�ySJ@00��T�3��3Vy ���'X�ȧ� Dk*���T:LDX[�'����L��<�`�Q�T������'��Pr�͖k�:���G�l��"�I|X�{נ�gJ��uF�>q�����?D������}�ݍ'�h��@�3D���Q��:
ގ�KƊ�x,��1ړ�0|�Q��o��$�5��L�,��c�<���A�Wa�A���@�+�ACz?��'qO�"=�af��{GB@��DZ\�9,�Z�<iB�͸U��d�ۼ|�:�c�X~�.1�OL�d� �MCÄց�y���'@���$ƽ�4I뀩!VOx��kÊW�!��u�ndy�ŏ�Od��tI�2%�Q��F�%^�L�W��/L�\I����y����wM����n8'� �B�5�y����G�Nh�0JU(HO��yů5�y��	=�QJϣGC� �bA=�yb��N��W.G.@�B#E"�yRf�����Bg"B�/sP�:�)X��yrh`�����c�$*�pQ3n���y�b��Ӱ�\
9�hd@�$�y�*]�=��b�U�0ĸ$C�H���!�S�O�X|��T�HN^L��oL�P1��hB��r,S
?
�1���|����=aۓ;��z�o��>�X�(A�н(�����M�����H��Đ�ϛ�
6�u�b�VE�<�˛�*����� 39���:6��G�<���	r2Ek�,N�L�����|X�tDy"a��gv�`A޲>��@��������OH��� ��K�
\:@\z�'!2'��B3O���d�S�O���c��Д~������I>��p��'W@�`��P7�^Ex1��K���(O��7B2Q�b>5��A�d�����n��(��h?�O�ŋ�'�dCݒyu���`¾'Ue��
`y"�'���3I��(��$0@�+?h�;���i�����O�Z�EK<�� �B�s�E��'����#�A�J��M���>n�������(O?�ĕ'<�⁺�e&T"�-�(L�!�'R"�sE痐-�e:��|���:O 9 #jհZ�F�Xs�D���"O�e�nO��x5@�)��E�$�O��w�g?A�P?�8��#�ؠ*�	�,�y�EZ;���3�gȲ����'�����d�<iH>���m�����`�UV@�3��R�'SFQ�-F���9j�'O�5�=�7��g��D8���VC�VR Y3��]�%:ĉ���1O��O�����eɂ>��p#�o�`����L�e�@�'b�e�E���B�
Z�'c��D��Õq���K蘽`%����y��X�2�$Q�G`�A�e�$@���y"�ϹK�����ޓ3 ��#EΠ�y�CZ
C���BC�^�0�� 7���3�O�ӧ�#q�sa,O0
����'��I�4�4KT���Y�z��\� u�B�	QT��e�_: z���.�"=y��T?�ce#b�}�ɟ�b%X�3��)�	h���'s���`Ë����#D�O�N=��g��DD{��?͆B�mX.p�$��Nݏ�HO���$D��]9�LҺ7�Lt*6-�u3!�䛚*R�EZB�)�Bݸ���hF��YT!�� �@|Ptt%ī�y"m�;[\�s���C2�[Ci �yR$޷7��}h�*�4i�Q��J0�y��u� ᆥ�>����S���� �O���Re	Ap� �E�i�tLʁ"O�H�!�+<��j�D�+_��0"O~�Z��lJ�����J/+U�|�"OF�Նٴ}-օ��el��g�'��O`<�@�ΩP�t;�+|3ł�"Ot!���E�t��ȈP&6�a�"O"�E��	*aJS�VvU�"O�1�����~ތ!�WFG��1누�y��لuJ�	���&Y<�)�Ñ��y
ی�L1��� �G�W��Oޢ=�O����S럮;�x�h��J�e����'J��!�]�$h��揖�bz]��'�ҹä���(��@6���*�䁅��~���K}d\�TC�7��21�FXt��<a�2P9Ө[>��\pvˇ7M3�ȓW��-��ňJ4�SM��8���F�W��X��7=��}��N`�'�ay�V�OFqB���7t�윋����yb��"�H�A2MY@�0�#��y�g«qS4hi�-4;@�dk�3��x"f�)>�� ��R6X;r%�Wą#9!��]=h�����2�l� ��(1.�y�I�3�̣ҫ��W#n1�6J�cŘB�	i��m*B�Ϲ@k~��#a0�ZB䉥5���a!���y�5��{XB�	z+�8�ÃԈWF�Ix>��m�F}�L�OTb�Q����ͼN㼅/�E�|$p��B%�0=q�r�V*2Z�U�� W�̸�����q�<��DÀF��L RLܱ1-���&WaqO4�=%?� 4)�f�q+�� ��'?Pp���"O��P	H�f�ڍ�O��jid���H�'B�	���zǜ�5�z��f��M� B䉶u>�ti4٫}�x�� ���B�ɠ^�6`:`G��W`������f0B�I,A���X� ������1��C�I	Q�6�j���?I�M17�ż9�
#<��e>�S�d��k��$�&!�k�vx�+��ybė�y"�$��0�64� MR��y��)�?��@r�L��}{b�#
��f�"���P2xQ@0�D5���U�5AY����$R�;��i��>�pQcR`4H&a~�\�h����=P������ΦnK���`�.D�h��웭!��2AJo �9K�E8�	X���'gT��̔��<ѱLѲYC~C�ɻQ}N@�j�R>~��Isa"O8�`@fӢ&�����@? ���w"O~�{ǋ������#��:�F��"O,�B`�ɩ@��k1m �4垍+"O�����Qe���BiW1rĸ�;�9D�D�#��;E�,ى�(T:G����i4D�8
�jE;l]����и,��-Ӣ�6D�0�l�5*a"��c$Zw�╰ӥ6D��k`�=\B��"_�\�����yB��-���6J�:FE�x��	��yB��0��iСJAA`�q�CF��yb!�3���"҄ݖ5m�[��%�y�(�,F�,�C�5'�A3�I���y�'Q�K$Ⱚb�P�p�ГD��yF��\ֹ��D�
�.���ʜ��y��Y438,IS@9}�@S�K��yR�V,5�fl�&�M�%��-SR���yr��<IZH�C�G�i���"�y�� -�X��u��
VN��3nŶ�y�D
Y�V��P/( `0H�^��y��-Lu� G�� '�pd���yb"�	\����E!�ku�� %Eį�y2@G=n�b���(� N���D��y�$Qsi�s��G�.�BC��y��4�B�ctrL��������y�
��R^�8�HW)j�1��ㅝ�yB+E &�f�t�S`��A��S�y҇ ?m���s�֪:f��B��S��y�(\$.v�cņȀ.�n]���� �y��ٿR:I�Q�.LL�sG���y���{I���I� <�m�����y2�Z;
�&�r���������$|������ G������0=�s����t!�O�&5P�
J�<�#���H�����䃓��l�<)��$X�@�#P�+��4q6�n�<1�C����,�pK�Ti��0%oKe�<A6o	
o*�d�Rg�&/����fɓX�<��n�m`H� POU!`S�RT"[�<� �Y*y��LAT�~0��)|�<��㘶}7~� ���&�R�x�eOa�<���ǒ3�v���<z����\�<�����.��!�Bo��� S��Y�ȓc�������j1e��>ȆȓL� ��ξH���y(� 4��(��Z3��C�!�q*�	"�<K�|!��x��&�O�$�޵iР�>>��?f���� @�����;2]�Յ�L� ���$"1 
ā��>Z��ȓR#�\���N�?�2�GK	�5!5��S�? �ȸ��I0C�,�#f��BްI�"O�(��ȦgL 5�CG/rO*<B"Op+��%b�m�E#g ��sD"OV���ԗ;W��w A_IV��c"O����J^R�MK`O�E�䩖"O$�H$Ӥk����m�$��"Ob�C� X�E���T�;r�Jq"O����lQ'*M�%��r�l�"Oz0���B�W����܊�V�G"O܄��a��9Ui���Ի/҂$��"O~����sbD�����@� �	�"O汫�g���x �E�0,�(���"O��cJ�!���e��̵a"O���E�|�VU�w�Βu�jh  "O�T&
@t����Q�kx@� "OR�B��X59�hcB�d���"O}�6��"zȠl!���)j�<H""O<�cUk���]�O�?p���Q"O���$L�୩7�(OwZ��"O��3�^�(CF 	��ú80���"O\=2H��|�ԅ�*2�pU!`"O�M��]��� �!��1>�8��D"O^j���x���!��̼�ެ:�"OB	���0
��MC'�z<C�"Oj����M�@�%T��(W�4�"O��"CG��!M�ءbkׁ	[r�H�"O 4�������{F�(��q�"OB<;S�Q�PbB��%����}��"O$�s�ƉS� 5y�*�֐��"O��_�z 렡���b��3�y�+�T��7�M��:������y��W�[��⡈����$K���y�G�$�DyW�4|�,�#�O�/�yZz�����ԬD��Q%�3�y�MςE�:%�͕+k� �dn���y򢀘-s�A@V�\/w�p1��̐�yb�ЍM��\HTU><�ȝ��3�y2#�
n��P��+¾�R¨׉�y�?E�N���F-	֑����yB�M�k�$퀧���1kG�yRI̧%� ����
}�H!�H_��y��7+j���K5y�(��3L��y$�3p^���X����F���hOT A�,ܗ�H�T���痔LT�������"O���ꘚY�>�`���M;�A��� K����5�C�S��?�`�%�eFH�<�P�!�C�o�<���uȅ���~�	��eͫ�!�$P0&�.�:4�>�5�Ί*+�!�$Y�Uj8]pB'�-?n���d�L�!�d�Hؾ�;�j]� �Qp5�Ƣ	!��ZA��ܱ��67�=!�b	�8�!�$�*g��q	gf�#v`� !�S�ўۇ���o]�>���iI"K����F
�37,Laa�*D��!/�[���f�
�B�,ŁFhh���A%+԰Î�O?7��_�0��EeXO~~X�Q*�i�!���j�p	��Đ/��h�B)¾ �dX%��d�t�˔�0=��A�	��aXE$ӟt���y8��Ԣ��b��t��%ʥ	��9��@�rndp��jÀQ�!��ظ'�ĭ
��)59&�P��aT��k�\�N\��'�Ia�n t�H8%?U�;��bU�.=O�����9S�^���wef���j�DUA�o�w��qw�֐^3���M�v��2����!o�k��b�TZ���L���m
�hL��))O>  ��7+j(�Q)&'����댕nH��:"#���)r�4�~-(�X(��M�Q��� f@��	F���A�C�t�a����Ս»�t����� v��?1�'&�� BH�W��>7{<I���AKh��"O��(6���G�de[R	�<l��Y�ɏd��7'�����F�W+��FG��F��D�Oʴr�w�vkVH��6] hB���j�I���z8;�hLP�@��6�V~İ��mA$��@)U)E*hv���[��$ʩH,XUːK/�I�E���ǁ����S��J���?y��<.n|J�ΜP�2Y2�Ѥ7�HtBS�[6`S���9Q�&��)Olѐu]��z��ک 5΀�T��v��]qu�ߨ��d�LQ��+�%�z�~\��jI�0�6˧W����MZ) 7*EI�F��(y�'�xz�=��'�t�p��
4��(i�c��q؆P!���� �x�g:x�yG�ɗ@�6@�jp��s}�epޝ9�� �u*�g������+�O��	v���o�J�)&��=q_ҙp�,�(n��`�V�dv�{�V��ɡQz�]�!�v"�'�r��QL�%G*D)vg�#V|"=��$Ǳc��(ŬX�|�\��� �2�u�K�% ��(�c�L�1�������C�X-��R���<u��$�$���ת\6�xPg�E}� Y'T�\a��i;�,�&>���%�na`��%�¨Z�� !ވe�2q X�s	�'��L#�>@t�xz��ۻ( 9���13��'v)��Ð�'��|c�c�Bv�D���y�;]��5K�1343`�(�Ve��I*T�|���/�5;Dʁ!d$U��*�:`@U&< 6��7�������<��"�hq��+H�*��Y�tB6O��F�
v��1-�8���*#�N���!�#�
\���%:�^�Ӓ+��2� �DA1��E0HC�-�P,VW�� 5_R��Ɂ8|����\ a|�	�A�8Τ�!\J�*F�*&�K��� 9~��<�L�`� b���ӧ �D�*Y���4/�A�A^�1gB�	�D�>�
����l$,�.C0*�X�
D)C)AD���u�( ��Mծ�ީC
@͓t�&(��t�!�����b+6E�U	��#��8r��/�O�4R�B��P�ǥ��H����/�/N#�ݘ�'�Ԧi�C	צ��'���R�%f4�l�1�@̓V�J�:�Ι86D������ �&F{R��8��+�.��8� y���=��)�>h��Bk
�@D��0S����G�,��@Q���p=9���S�Ƅ�BoE�IJDȆ֟�!ˌ	?*R��'A�|t��\]
�6!�<Bĳ饃�H�]g@�b�����ǏpD�B�	�Th0kOۋ�~T�"���HL�`F�$�X�G�*XV�����R��$�v}�%��P�G�`X�u�lz��'$5P*���5R/ 9hG�S��0@v�˒
D�e�Ŧp=&jeK��MS2A�Hy��*_`{��ID�*n���&�+Rg�1'��"��D{"�Ju�$�V��v�ҩ��Am2�I���I`�䟸5(T�*nԖD'�	�eK�k�Ul؞ط�J�}m�Ep1�8�b<ЕNa�����݅k�)ѳǁ^�l>�DN9
~�C0�Om9��F�1̔���B�:�,t@
�'�b��`гuQ4����U��蠒��<�9[��$���/�f�˘���\���95h��3GZ�x���2W�M�~�$�i����舭�4�4
)�WJ�/��Y���'�X2�)�+X%n��� C>� hK��
�B�:��B�?m:��#-�~r���eD��͑2J1�ap��r�<�Ŧǘ��cVg��6� A�\s}Ҡ�3;p��QD�ʕ!��F�ԏI��{3c��r.�S",���y ϴR88K!��Ot-����/
�D!��`�H��W")�:���y��QXz�5L�i'�����x��9S��i!�ƌ��t��cR��:���ɝ�k�8G�b<,��!�'1,ܹ�e�~4��>	P|	a��Ă/��	��T�[�.H�Ed��q$p��ȗ������N��e?����h����x"̈́k�JXc`�)&�&��VÅ�����Z��l�`���>�x��[�ޔ����J�'���iT�//��	Ռ��yB����|���7����]5
XR�à�Iw��iQ#Aݎ��}�H~js=��}\:�� /+#�&h9����{n��&٧xP���I�=���bV�>�Re�Kɂi��`�#Y�/�~Ż��fX�|��T� ��mA�h��0���5�	6\�Ch��=ړ�ڥQ�l��@�Ī8��8�`�Q7���в�[�B�HB�ɒv��%!@��i{r�J�'H�?���6�͙k��%����d]"pC�B� :�ӆ?��� ���ݛp��;�"��I��'��""
9��G�g���T!ު@�Rb����d��$?=�x�DS?�����M��ZR�x�+��x�S�=�}����Y���P��)�J�A�X��q�5iK� �����'p��C,'�5u(6�r�xǓ��ts�lT5�ڄ���p�����=,��J2M�T�X�h:D���K���DQ����x���G�9D�DQ�ꙗ>�L,{Qn�t[�i�6�7D�� ����\�o�Ti֣O'0�|��"O��h!b��G���1��G�`t\�R��'ge�qf���I�]�<��l�H��i6�McpB�� ���D���op�q�+̶v� b��a���7t�
�Q�e�|-��7��3iӶ����'0@
���z�R�I��T�q�)xt�%#Ѐ�/O\�9� 1�3}���3����6����%	��xR�ֲ=u�P(���(�j��Vgʩ	7d5��'��wP((���'W�i�Ӕ"��ARU��z,a�ϓ#��i2�$�|"u��'u"�A��3mtp�t��rcj��'ND![� �'�p�sA��i  �K>a`o/%�C�T����\i!��p߄����Ƀ[����"O�Q)D�<b�̹�vM�s�^�#��dM��F_��R�΍E�g�� �U�zQL�jg|�s��76<���J9n��I���TJO�P_����&�6x�XU���*�O�X�Dˁ�M�ص�r��4��E�'�ܡ�C�17����U6OH�т+[t� l�P�ԖW�*��"O����I	�&`�ʱJ��4
��$J�H�� "��	񨟨d+���ZM� 〷R��P�s"Oj�q�"��DB�!�ʗc�,��t��V)<'���T�<���K5��p&m+h��H��O�F�<y�M�og4��$���C���:��o�<Y	��&���`]� c@��	NO�<q���≮u� �32����^K�<�ĝ>q�d�v'ƨ4Z"�S�!Sh�<�G������c��
+_�}b���e�<	a��>�x�Ѥ�M�a�ʡ�1[~�<�q�a��E�q�'TT���i�P�<1��N:#ܠ9t#,�~�c�@�<���MR}B��0=�EH��Nx�<�+� �ԠuA�eE8��c$�L�<q&L�a�b� 3�̓TS^DDi�I�<���1s�U�shL�ij�`1��VK�<����'�"��QE� \���w�SF�<y��;`����v%?SP ��F�k�<�#(G& (T�gK@ ���m�m�<���Iܑ0�B�)��)5��k�<�piY0t� �
��^�)�h
b�<Y1Ş�	��M�M�������_�<y��h�!�gٮ��y�c� |�<yq��>J�Z�HcM�7@ T;�`�~�<��K�tz{�K��u@pdA��^�<U�1��]�6AA���0Ԋ�Q�<a%�}�v�
9'T!�B�c�P�ȓ(S� bF��+wŶ�tC�n`��I��x#cI�)�ެaGJ�7�H\�ȓ0�Ӕ�ڧ]�H���]�$3����?��҄̄����"�]xE,��G�@vD�#{KΑje�*�؄�3j8�&K�"T�xZ�d�b-p��[`\�%���a���a���j]���ȓT��%
�H
�*��	u�[TQ��ȓ&�P�B�
Ki�-1�k�x��(TA`5g��l:��H�b<|���s\:'� 2z� �̱>lņ�tW��c&I��$ģ���5Z1�ȓi�Ѻ�	�� ґS�f�_%�4�ȓ:dH���a�%*Е�#�zV�y�ȓ���0�뗡���B�����[
��1�ܷ:�
�9���B��x�ȓ/���V!܍j�T� 7�8ik3�(D��z���5ִ��+r����p�(D���� '	j���A�yb��&D���C��,�"���'�b����3D��  �JG%��#a�$p�G1���"O����B�
H�6�����3l|�j�"O��ɭD�,����D�j��-k4"OAr@X(j��q���Ѻ,�te��"O���ԋ��tg�?�zň"O�m`��};h�7L֠H����y��6���� J�@X@�K�#\��y��0�X�al��A���@�� �y�<��T!�#E�j�HQ��y��6Q*IkD���49H(˥�ő�y�D�"Pm �`��wz� ��Ԁ�yR��$b�:$����X��"i��yb�	W� ��ՅF���D��y2�L�0g����>�h�0����y�o�B~X���C1$�i��-H��yB�ҩ*����w�߅3�0}!�+W�yr&Z9(��9�n�.�@��KH��y�J��L�b��d9$���ף�y���}$}y�FÅ&^�����0�yB�ѫz�Zq�ai�'#.X�	���yj^k��j�GO�(@��CmG:�y�k���� qN�C��H��y"/�r,��(h���@0kP.�y�[�b&�m�Ņݼ&��qD)�y���:^�v��f�@ ��Y��/�y�k�+M4�`�c�W��B-8���!�y��A�`��*������
X�y�bJ���Qr0�H�\�±��(�y©��'��Y�iMOA�%(aV��y@D)"���N=N� �N(�yrC]�_�
�I`�)D�Jݙ%)�2�y���?�\�[���:��̃���y�%V,[�jy���6��1���yr� (����B�4vFL�����y"��E�p䊤�̹E� �+D��y�҈%@�y�1�7<��%	�a/�yR
U }l�y��ٴ#���4�J3�yr��wJ�t[���3��%(t$��yrfn�HK�ˏ�B�ڡ�y"��W�0�ɥ�C��@$��	�y2`*$)��́#���� �%�yRB��b��!�.0*�G�[�y��[��Vޔ%@��!RE���y��̯5T�a�Ѓ��(��D�!A�5�y2D����HP"R�*�N%F�yR�<��yy� ��q�ar� �,�y��Pq��+j*@	e���y��Dk7��d�l^.l ��yb�ǉ{r��8�D5\d��	��y"�==8�<�sf��S��۴
� �y&5~�j�P�J"9��6jG/�y�W�N�(����(��t��+ņ�y�%L�9`��Q�D���¼h����y��A'���K��I7	�l���i��y�
D悰�0Q�z[�% ���y��U�)�2xc$l�;if�|*�O�hOF`ju#J �H��� A�
\����͖�Z���X"O$ي4��(B|$bmB���!#%�i��	�D刎%Bɧ�����ǹ2��ըQ�ޤi�"ő�hO�y2�Ϝ|(C��/h�����Á�~�hX�7zv]�4-�h��,C�8��5R�o�>1�8mf�.�O���4M?Ü�����H�\,�eF7m��P�'Ú�y∀	==nD� �Q? 9��튭x�����
˓*��B���T(���� F���ÈCL�d��J�,> B�)� Ll1�	2 0� �fK�'A|�4�C�Dq�S�c��k��p�O��c��Y�I
H��{R�A
�u1K�+!�ڭAg��B8�,��D,8��4R��]�!�@y���+"�P��U��$"�(Z��$��7��H(��Q0�0=����(��\�S�#Y��I�a�x~B��E�ͣb�u��4
��ߒ��4X�p� C>��T��S�q����b��#5!�W������4v�6��!�%�du @{�<UK')�5�p�ɗ����O����y'�^�ynrHɁ� ��"���@���?9dF^�|�µ�CfϊR�0�c�U�[li�l�>j�`���;PV^a��OJ�qs�D�v�㞨ɱ,X�TqdZ�,��TT �鰏5��a4\�)P�0TJaa`'�=P`|8�Ik�ђ��)c<H��D���d�7I���0�'��I@��3ϚT�׎F�n��EY)O�(S�8ߴ�*�%D;zX��A��|�j��A	�EYM�6�+�g���Z�Fa��y2�]�� ��8v��s���uҹ���Q(d�{GK�3a���3a}�:�a�eݹ�'�H�58%��d�MCd���H̀gXR��d�4;- �P2˚��Dup�Q�t�i6dC ���A�Մ1�2h
�_��&�S�ꀙ|��F	M���� ���!� ��O6�!��ƳYB
�K2��] 8$�Yw>
01�Y
-�i0�ʸ����OV|	P̂�v]�I��|� �	�d��4�X i4O����'hb�h�Ȟ1QɧJ�(�R:5zG�օ:]2��)�-m,�PGS�O�Xd��O<���v����D�u�%qE���:Ŝ��A!���E�OZ�	��U�|�e-��~?��Y���;Sx(��fC}�<)e�
s�>%�Ϣ �ڲeT�Q���k�!f��8�'ZB�D�,O�2p��29�ժ����94f"OT��S��,v��]����x	�dp�HU�>��2��X7:pq�Ǡ,<O��'�
9�W\�M�$��a]]��܂�.R<O�zA��ϊ~6@x˷ѓ9U0�2P��I����G$4��5�	�Q>X
�h^E�e�F*�/ �&t[�E��HF����2��[��yq��":?v]C���/�jC�	'& =��р�~Y�`J��\��Ӡ�x�η��`��<�K.l�bPpsJM, e�Gßk�<q��\ }xU��A݉rք��gGJ��@r�V�)�� Gm8\O �(����Wܶ���a޺Y8�!���'��q��.�i��`(`�i�f9��&A�b1b���`D�D�����'��I�4�ʫj~��z-_�n��j�}��~�Ӈ����H�F���fA	/�`4��Oq�L�Q"O�����K2?�pI���Q��	�B�>q���d��&�g?��OH�\�0�B�Q���D�RN�<�U,��dRP�2Y%M-��dk��l��Ť.$�A���'ƀ���̍�G�"�IA�ʝ����
�ZU��դE��?)�#�|�IA�3J�.WmM�<��'��Ҥ��Jn&�(!DJ�'C0���gXy�O�v Y��x2��AV*�@��'B�lk6�C@�t�cE�G=u8��'�2�p�̂(:��5d��
�l��'g��Ag#�u:>���f\4BV!x�'l����D%_��<����w��yx�'���Ya���NY����g�Y.�5��'�:8jg� h���t���T�8����#v����X�L�*�Y%��;����b”� ?Z;�}�2������b���U:;j��r��ƞ
��8�s�<MT�����*Nj������>��yb-[�e�d�(R���Bj&��'��O�i�EC�4d:d�3%�h��D�v�Y�X�� ���ӄ :'�<T���'�p1�DA�I~ X�̑��Eb)O E� �0B$��I%_:y "�R���O�=#��͵��!Y5����H������hTְ� �O&^�
��[�x��6%��p��A9��%?mʵ�x"��pOTTk�cBr� I�F�І��?�s��v��]���Ŵ5v=A�"I#j��J�jYO�Dd �W2 ����;,O�� /��U��A�s��쓄�	<
�B��N.pع:���� �eQ㢓�1SJ�%gхS��R�?$��P���HҔ-�V�ԝ=&��
�<A��[V}�x�`�(#��c�6fO�c?�"��=zy�tjG=d�.�bk$D�$@O£9���X-<�π�7�.4R��!*Vv���"�>R���|��M<�q(L�W�fQ����	=����T<�Q�O70�c�̏#=J�w�ĿC(��$���T��0��#Tz"F�3�S�? ��G���2@;��F7+��u���'OFl� ��2ߨ$��)��9A�1�޲V��đ��[0sq�9�5@�c�<�e�?�TI�p�ͰDƌ��EcIR�<	4�D@����,A�������SI�<���J,1�Dj�/�?	�R��EA�<է���p��e
к]x � �|����n�>%�'��$ҐbA�&D��%ИvW�d��'��rS�_(;��K�bZ�^�i�y�"Z \�}#i�O&m�q�'t�N��Ĥ�����'<�5&M+<��q/\�*��� �Zeؼ�(OH�p��3�3}oB?c\ 2�n�_NV��B�	S��Q�Y,>d 0��~��!�_ +��sA�F� ��h�'M���$��4k�Rq���4<O����7m�JY�Юt� ���	�M���{�@��QA�\Ӓ�!D���m�&v=q��z� ��>��×�b�@w'ߣ�""~�eMV3W���p�$Q��Iv�<I� Q����1"���L�y"���2
�k�_Zy�GI�'���=rm���Y!%��L�H��u�Ɠly�@0��E�9����Cᏼx~�a��	&�H\ȣʞ9�0>)B�\
Ib�I���v�� &_x��Y��/u��3PfL�<�`��$0>��r��O
ͺ�bG��Y�<��)@����qyN��ÍZ̓yF��-H�� �~�3LG�~�8D%�l� BP��P�<��ÜN�:�"S�j�J�q'��9<�q�T�|2�WS���d�HBE0�A	�;��P�n!�DF�/x ��eI	.�ͪFU�F�!��L�?�Jh���d�|\��eע�!�\�C�4�x3�ȇ)���؀�Hx!��W���G&�=F(��:��QXj!�dM5�L8�Ŧ�b(Q@B�:~!�$�s<�낭�n��9��B�]!��	�R��L���K|~�����2T!��7Hf������$Wе��M�_!�D��;U0������^J��J!�$8WkTA!R�'JީH��̧UO!�х@�pd@�N�Hb��G�$ !��@�J�a(�d�pa�옐g�!�)�е�b �4�}[�k�#kB!�d�#t�j(��	>K�*�� �%;!�D��yt��8A�^�F����!'!���䡒��J�*���Kw��!��u��dh��$f�$]i�GC =!�IJY;i�4p��`FӃ�!�č��2.�7BjR��q���6!��¤x���R�Ť	D�hc���&!�!�dΖ;�N�� ,��ŅV&a�Yw"O��*���$U�Z��EI��d��LS�"O�e:E���J犀
V+V�V���H#"ONEё�ڬ8�<x6�� )��v"O�Y5)Q�E�R<����K$���"O�|��aҵ:b(�0�ӆ^HK�"O�lǫ-u:T�1gQ#" �U"O>��H�I�v%��F	�!��z"O�]2BU{!�Q�V%ȁ8F�9:�"O����kŦTHh��/$+z�DbϞx�HP2udG)L?^�:B�'mq�� %�B�k���R�#�'��@�U�D��
���.I�J�����'kH�ic��_�� �(L;3߄���'5�@�!M�q�X9�t�\�+d��X�'H����#I'
�qd ��(�����'[���s�N'/� d���$� m��'oFX��V-?r0�FDd���'9� ���E%�����13)�1	�'_��O�5�N��u�F���O�������]:���J9WH��	����IQz�+�^%�R,�i �3� ��K�M�Ɉ�`��H���R�DYz?AFlG�gGѸ�(ղ�0|C�t5��a�h+A*�F	Ҧuk���07�	j5h �B�*�)§��DoRz�Y���U��!D�M��$ѩ��ۥ)�LX�o�Ц�A��OC�o�08�ݨe�ݝ@?���'��8��� �#�ͦ���G�{��O6q�P��V��Z vɐ��P0Kq�d��$o�z5�'�.�!�!�R>�3"�ݝM������N�=�GS~~¡I���	r�^f�����2� ,������թ�ҏV{�DI�n�AhD����S�L�L�a� �-b�: f�J���,�O�r�V)�������UF�j5r�r5N�?��+%��Xd���?�{���d��T�bT
ǥUx ��:�
�yb�\5cE��r
�<H�� �����yɒ/1��]�v�˫6��(�%��y"�Y'��s�Ë=w8������y�B�=M� ��� <�����ɐ�yR#�EvY�
4j��A�_��y"+\�e���V������`��yrMʪw	�"�@�b�A�s�Չ�yR)�3f�D�0��40or �Ѷ�'�n%˷KWq��ȱ��͊�(���'
��@M)5j�D��K��]�'��U���:|�T����&P��'�M����f/z�;��H{�,�1�'�@|is�2�z��P%��t����'��B�Ǐ�!�$���svz��	�'VJEJd쑇.�����	Ӱ\�@8	�'6�X�'aH�h�r�򐥒�M�����'�����#ޜa(��BJ����'�ʤ�u�^4I���
G�z��'Ej�p�EV�Ci�ǈ�ׄ9D��0ₚ88#}J��$8�D<0��7D���g	�0.����� Y#&� �,0D��z'eȨj��=[��؟Mв�`�e1D��s�^=pJ�����W���Z��.D�,��^]T��J4!Ӵa)v��h:D���uA�q�JX�S7�Vpp�6D�t@��>=L�i�̳]K2����'D��4N�Iʠ�{#�T�&X+�i&D�������9t�x* 50ʩ���#D���VAު����/]�x���y�&#D������:L����?@g��0�+D���7��,��u�s�8`!R�-D���v�Z1`����ق&�2�)�( D�𡳦��)�lm�v.֙����+D�$8'�k�l�K��)To��$�-D�<��B v�y���ܛ��4��* D�Tqd.I�EX�I '$T(l��k:D�xI�m�y��L�Fė�"�@�ul4D��1p�5�h �áս6�8��E�2D���rk�	�L4�/Ԝ�"M�a'$D���w(]"7������1,��h*c�?D�HK�h� �>H� ��,}��C�9D��(��]*f�p��k�6�.�5D�X��
px=jr��J ��S6�1D�ԡa5iv��&(��E��Ur$%,D�$���	��I�i�6c��/D���)>sVZ�c����%,l�!��ы�&433H��m����c��"_!�dM�q-!���6Rd�g�S�M!�$
�.4��� |��mI�-B�J!��Q&	$�9;7d�2�}�Q�ɛ6!�ڈ[��&ߨ8����<��dɎf��CaI�[����%,�y�BXB\�)�D��R�2Q��g�<�y�"�{��-K1�L�9D���J��y
� 
K� ]9�8��7@P�	{f"OȚ�lC?	)pdH�XޞP` "O�t���' TyA�ۡ ����"O
�2q���v�͉�%�:J�ɢ3"O����ʝm��T�j�87��[�"O���!K6I�֥�b	�"�:�K�"O ��C
�n��$��8`�u�$"O���B�F�\R�ta�*TO��!�"ODȨ�NY�7t �)�%9�|�"OڬI��-jI^	���K�JڄS"O( �W&��<�4��IԈT�0!�"OBR�`R�-��p`�H�'����r"O@��Gޘ8L�°(p7��"O�h���FV�ũ�n��%&p-�@"O:=;�Ϗ+5w�˃.Ö\��"O��hB�W�s�����H� ls$"O��(�.D�~Fi�3.�)�ʑ� "O��G���m�bE���@��U��"On1:�K�9�&�XB@^	7�q�1"O
�ڰb�@��ԛ���?LL8��"O�̢��W�PFh|X�/	!\�lV"O8YP�`�� ��-[9���ZP"O��)���:�$@��ߍKx&Mp"O��{��N#\��ዷ�L�	k�0b"OD: ���4�\�)׭Xc����"O6���H�Q����ge�uZ��b5"O���1��.QxZ,#Ge5����"O�\k���y0�3��K�!JH`h�"O*U�w'0�1s"Q�9*|x�"O�	r3�L�Y41K�	��
�2"O�0�O���=�uB.)�8�8"O�M@�M\g��Dj�jשp�t�9u"O�9]�R�q� ��T��R"O��Lڈz)���U�Ŏ2%���%"O�3%�	�VQ����
t���%"O>pd�_�+����c�5�X�7"O����aիq �4 W�<-!"O0��A[�{�DR�HHd��K"O�$aW�=�j�2>{T�!5"O |����~8��3f)���^��"O�`��`F"/�.X���� ��2�"O�\���-#�a�E��1f�7"O�U�����T0��T�(
$5h�"O@x:���>� �ЂA�a� <ے"O�KTIɰE�I���ގM����"O�Ey�,Ǳ��܃���ۜ��t"O
�0i˾@�Q�X����"O��Jx�:��������V"Ot����[�L���г���D`{D"O\@��J̒T�YF@,sF�"W"O�����	�&�걪�8ru��B�"O�Ъv*UA1���ޥil�)�P"OF����ЭFB�i������!����  ��bE�sh]S�H��&p!�D�8l�8�v�ř�1����dn!�Ă�hId�Z$�E|պ�� P�_X!�$�%;��Ha��ɻD���'<!�¸4М�f��K��	���ߪ6!�ēJ n��s�F�^������ե !�d�9��]y��]�H��b�f��A!!���n�:,R ���N�����T�y!�䐝BV�l8�kΒV�Q�%F�E�!��t5� h@+óc����%��"!�Ą/��T9���y�`	�mذ$]!�� �@�!�X�i��SÎ?T4T K%"O`�X`\.~�<�c�:%�*Аc"Od1K�g^�<��p.M�����s"O���u�2����\�C�����"Om���H�9s�l��Ed�q�"O��	WJò	��S�7kz��7"O`���ՄAS^T�����@S.옆"OPm�e
Dg��ă��=�6"O�]S���X�P���WLTH�"O�z��eh��zt���
9T�R�"Od��$�@/W�\��F=�=�0"Od"��	���E�`-"u"�"O��RU&�{�a�c�%+���"O�в�lN�K+$ͫ#��R"O�� JQ@D�;U	U|ؚ"O��bU��g��L��![xy�6"O����B�pI�1��؍6ļx�"O�h����j{]AV��
���+�"O� Pρ9�e�`Mmo��2�"O�Q[PLS3%(�%�竁	#i<�Y"O��5$J�Vi
쩴 �Vjp��"OT�Ǉ�%؀`�uo�*kVbpQ�"Or����5G~�Q��NOb�d"O`�W'�-Dˆ�9���Q��� "OPy�W�V�~��(C��ݮ�A"OZ\�`DN:Q@����1�6q��"O���Qk1]����2e^,W��(�R"O�Kf_�_��L�#��=J���q"O�X�'��va�-c���,�M��'�ja�"�,	ء�6g� ���	�'��2��Cl�5�S(N**p5��'j�8:w��hԶ����&����'ȼ�9�s����G�/t��(�'���w��.@�lP�c�(�0P��'2�d�G�7�(A�v!�QO�̈�'�<a���� >��A��$�=~a�'q���7N������%�HĽ��'m4D�
;�(�����E�͋
�'h���p�\�L���Ѷ���E����'�.}3��k���Fg@��k�'�4��o��S�N�b-��9
�'�(�.�G��)��S�rFJ��	�'k�����=qt�S�߁X 1{	�'�ҽ��Eϧ ˊ,b�b\RXT 	�'���'�
Z�Y�acAH����':�4Aц��~��	�B����'����A��h����뜄q.�h
�'e��(C�4lgXٱ�FI�e_���	�'���� R8�D�	3G8(?�)�	�'�%��#XK&y���V�'g�y�	�'�x�h��A��U G�#j4i)�',:�׊S�#m&����*�P��'O�Y��QGǄ�y���7z���'X�9�4�5m���%I��:��@�'V ���� 	�`���4m����'���R�3R	����=i�
���'Bx��a��z!M�8eȲh��'U���[1s?�yCq��.ؽ"�'���*@�LMt�!����~H ���'�`�! �;2�
i��#I0�'A�
��Y�0�j`8WLj
�'Â��0'0_8�|R7��P���'��#3�G�r�pQdC�.u�\�S�'eN��Ccǀ[�t$*��:]B�5���� ���'�5ir���@�G�:,cS"O�t�d!�p0�]x2E�G"O�=��"�4�$%R�N�V�<I��9K����dq�lI�I�N�<��DU0jAv�r�\�t2���I�<Q�h��Kpb��ǨX���D�<�&d�_�`�[�萌q&HxE�V�<���i��q{�&�*Z����O�<�r�L�fe2�n�g�~�ZA�B�<yp�����TL��;w�����i�<i��=ZН��.�;FI�toTb�<�c�Ety:-���J�x�<��r�<Y#~�2����ȋz訐!���i�<��C�*��a"E�}���2�]e�<9ԩK�p�8���4\�8��b/�^�<�����}(�d�G�$0���ys��Y�<!����?����R
_!7��z��@�<p��i:HT�� M=j�ZT�y�<����߅F���G��(N�h���������
�7����d�I)W��х�K��   @�?�   �  �  �    �*  �5  (A  nL  �W   c  �n  z  j�  ]�  ?�  ��  @�  ��  ޲  !�  b�  ��  g�  ��  �  j�  ��  C�  ��  	�  K�  � 
  � y! , �3 ; �D 2L �S �Y ;` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C�d �S�)U=w*����R�|cC��<H!�D�0@3�qJbʌ�h��K��I+ 7!�$O}_�%��h��F�h��d�S�0!�d��K�X�a�R9����Z��	A��H�d�ɀ�XfΪ܉�T�θ��"O8 ��)}�!pk\�'6.q�f�|R�,|O�Xѷ�������fE/��0��x2���&?-yN~J�ݩzGd�bp� E ��Q�
U\�<�������Q�ae�&
�� ��_ߦ��Ol �C������禡��b�3\����퐀h�މa�".D�$#!EL��8�0�R(n����>!�S�ԛ���3K�tI:�-�n;�q��>L��H��S{�@q�̴zn@`��JQ3m�v��ȓ	f
H�@��?%��q��V-L�V�ȓ��ґ�=�ޝv(^)���ȓ=\���wnX5o������&:��D��h�JQ���C:n�cn [���ȓ-�<s$��x����b$�F��O�7�*|Of����46`u#��
�����' �ɴXBDx���<WW�={V���KنB䉻���%13q��B���h�>i��	ڪ'�n��)\դ�B�d�/!���R��:1*  �#T�8��K��h����)Z n��1��ăQRD��"O�p@�� �K]�-)������<k�"O� �m� }�X܋�-�)c�T7"O^�!vB΋�����>#���Q"O� ��=tiztk��-g���"O�0��eLx��p(�G�~S&ȫ�"O���Am�N�d�R� i�`�"O$@�Jǀ\0Y�`�� =Y�� �"Op��#	8��Xc�e�䰸"O��x$��3��|�уSP�L��"OJe�����I|�0�4�3>��-;$"O�`�F)t�b5+'b�?��DjF"O8���������c�#C��`��"O�qB)�3"�f�9R����8a�"O�X�)7��0�g ��q�< :"O�YZ�׋i��zɎ5Yq��§"O�-�� �y"nta��be��5"O
]�ŉ�#x�R!Fa:�{�"O� �饊\2^�����J�cH��4"O��p@HH�s,�E�1B�!i�"O�ݫ2�� l�pi�!��~*DM�"O��;�U%�l�+n�1�6��"O��%�S�6����LN�o��{�"O���'�09k�8Xp�nF���"O�4�Ty�T�� 6x5Х�C"O��S��D���]� 3d��"On�H%�F�L�j�z�.߈w"��J`"O�Y�gJ"���E�U��Q��"Od���G�1�f�3��]%� ��$"O ,� )��zGLy�ѩW x���w"O�E�É�I���p���x�yv"O\���a\�Zn��!�.�-9�"Ohc�@�VLR��5h.2�9�*O
���<�8��t�[&��\�	�'�2� �S�0ȓ��˄r�L�
�' x�J�|�xԦ3~	��'Wl�9��I��h�����i�V�z�'�D/�3<���GT9*��hQ�'��p�ƍ'�^x�����(�t�q�'��� ��*7F��AI֮'(���'x����`Y�K�p��
P����'*t,x�.G�V�RljsC����Y	�'�f(A�0��8p��S<tdz��	�'%Tl;a��>$s��Gj�8s�����'�x3d$�*%~�	Rŏ�5�j}�
�'r�1���ty2-����)����	�'9|ɥ��GnZ5�`JA=	|�	�'馴xwl��)t&��W �7$��2�'��@��I��Y3~h��h�	�R��
�'�̘�4�E@�����/��1�	�'�P��ӬZ*%���E��#wLY{�'��bkZ�}�|D�#�@!@A!�'��84	�̸���%������'�T ��*�d�0/X/��2
�':������Z���y�/ҍG <�	�'7B�f�;A���h�m��D��	�'�N���N݋Ei����h,C �U�'Ɇd�VӼ5yX�B�D�H|��'�Y���?�<@�I�;�ZA�	�'��l���Δ�z�Mۤ�R��	�'Mޅ��F� N�(�R���[pE��'ڽa7CG3���ϓeF:�	�'��(�`	 d�T �C%5҂�K�'���G�7N��3C��&x�X���'9x�b��9[����S/?u��� �'�j��� X:V�Hè-t�0 ��'�,��"	�Q�X�����!����'���H'B��a� ���0��'���0��� GJ����I4e���'�@X��_-U�h�"��5AX����'܈���@��.���\!@j*}��',��#&�? ���"d�41��R�'"���u �)N:�˔(���B
�'?�H�$;�Xad�����	�'���1�!�5Sδݐ�Ɯ��Bh)�'�e§��5��8BtmI�����'�hp�O��C�vȁ������
�'xT�DR:p�����x�!�
�')5����J�k���p�^��
�'nP�#5f��%�� �"ɘ`��	�'z�|7�ϛ@/�(�A�9W�8�H
�'A���H�0h�p�`�#R>�,;��� N�)uj�+�ļ�㍙��*�0F"O�YY�GKh��Hq�_�1�r�9�"OdE��Swb�Tհwf�8�"O���j@�fj"��:g#�"O���KG�F表��49P@��%�'?"�']R�'���'I�'Z��'1L��$�FP��-1r��H�,УG�'M��'���'#��'��'���'C��m��/Kl)�WFېt0���'�b�'�B�'>2�'}R�'�2�'薔�ȕ�5�xX���#
�Ԑ���''��'���'�r�'�R�'ER�'7�����[*@=����W�p�h�%�'�2�'b�'5R�'���'	��'~�Se�*gG��b��.`ː�'���'���'��'���'�R�'7��+ᦄ�78�s���U�����'���'W�'+B�'��'_b�'_� ;�	��}R��2pG�?�*����'h��'l��'Mr�'D�'���'d^��#*
%�X-A�e� p�ni��']�'v�'@��'���''�'�� QêG�KȔ� �NC�g{l�AG�'�2�'��'E��'���'��'���Bé�kj>�!dOݾ\-�]���' ��'f��'�R�'���'��'��'�D�#z tb3�M�H�䋁�'r�'(��'���'lR�'B"�'ΰ�fOS�	�t�����7l�T�'���'��'���'R�uӈ���O���f��)`�"�0s2V�R�i�MyR�'��)�3?�S�i+�m��o�$+Z����fݗ����2�N�������?��<�|#���M[�g����F�J����?�%X��Mk�O��S��I?-�C�
9r���k���#h�YC��-�ٟ\�'��>����!�8����R�ZE��#�̘�M�.\g���O��6=���R���9p��a�G��P�zb��O���x��է�OEm�v�i�󤜑b�@��� F�P8���+��da��i��P�X�=�'�?�FAnt��"�O���R�D�<a,O<�O��m�?GOBc�H�ȟ�o�ʅ��!P N&zXF��t�����֟��	�<ɮO���-T��i[�i������ӛ�L��:d�$�RW�#擺d�B���$#�n�7M�dq�1�Ҋ,�m2�ry�Y�h�)��<�Fm��
���� �� -�%�#�<���i�B��O�1oZV��|R"J�>��%���Й��m��<a���?!�-=�`��4��e>u���M����ǋ��!����	�y�R�{֠9�$�<�'�?!���?���?YS�0G>�H�I�z��i��	��\��`h�������&?��/`�-�Q��.�ΨA��R�ZT�a®O�hm��MH>�|��,��� "�@?��!�IG���[Zx��?����B���kZw���' ��'���3'K�T���s�( ��6�'���'�B���t]��+�4N`�p;�;�lc�L�fƄMˆ��|��]���sЛ��r}��'y��'A�e�>i���C���y�(�� ��
�&��8�t̃l]�$�~ZV�������h #&	ޘ?��%"&�ڽHa��O��$�O��$�O:��7��%1j쬑�@۬(��h��RT�	۟��	>�M��	�|j�JI�&�|�N7Q~���gD�ݨ�S�	��'�7-��S�u�$lJ~�N:̨�K�@��M�D�N�3��cs�
��p�TP��"ڴ��4�����O��$�`Ψ�c\Gq�4�"�	YRx���O^˓&
�����0M�ן4�O�h�y��9��Z�� �`�H�O<x�'�b6-\��$��'^���h� F:yN���f�ٮT�ei��eBn<:�d�V~��r�2�'a�Ė�y�&S��<I �ݼ"�H�(7��C��'��'���Z���ݴf+��6KA�Od8\���S7�~l�pD?�?��z����d�b}R�'���h�*��GMV,0�o�4i*�-��'�2��+��&���
f����~j)��b�|D�v*�	(?���˒$��\�D��՟����|��ޟ��O9 �0'���8
����76�S�u��A �a�<�����'�?�"��y'fP�~���	��2`ʴy���
-"7�Xߦ�%�b>EC i	��ϓ%���1�Q���hI�̛jR�Γ1�r�@)�OԼ�.O�@n�Gy�OaRC�1�
�z�*K/�VA�dL#txR�'�B�'�I��M{T�_����O&h(q���D��B��W�L@9�L"�I ����Op��6��
� �@�`^.gj��,;j����O��ҧ&ٓzi$�������]w���?-��c s�N�J�M��VVbM��ȕ�-��'���'�b��ϟ��Ec#�y��M��N��uI��K�?1�i�����'h��u�J��]�T\�2�G�>lWJD�gA�7�x��۟��IƟ����զ9�'�u��?}p�'�#{�pt����!�$�p�VV��'�6Ͱ<ͧ�?���?���?a��T��ą2��������aO���DEɦ�	� � �I͟�%?�	�G
�m�����x� �g����O��O��O1�
�bo� �9 dۯd�n���&̢[���n��\I�Bybct�N�5���d�ƃiA.����E��,����?	��?���|�-OP]o�$�Լ�	�wu��F�F1�v��am�G �,�I��M����>A�i�7�OFbgk�
�R,�u��!F��U��@6mn�,���4j�4�V�u�~�u���� ��A��qR,��,��)��+s:O�d�O���O����Ot�?Q� �P�`���M%7|E�ŪMğ����tSٴ\��ͧ�?	Ըi��'�6�"�[v"RQ�Rb�?��ط�|R�'M�OfM��i��I�M턼IdM�D3�@į�Q�:UňD��d�<Ad�i{�ڟ��	����T�.�@pap��ĩߊ:3�9�I����'g�6��[� ���O��ĥ|�W'	S�^Ae�k��Y�7SD~b��>���?iM>�Or���霆d]Bp+�쌿<��6ǋ-`Î<S�i
˓?_�N���~�\��](=<攳W �+��T�N
,#�m�	��h��۟��)��^y��jӢ]ڰ��R(�I
3��*���r�&Y0:d�7ԛ��$	s}��'C��ڲ���3����"ܲQ2�x2�'@b]T�6��a'�L/�)�<�HӉ+�r	i�.M�X�N�6��F��&U������`�Iڟ�����O�"��䏞'2$��%��
��T�W�g�<�(W��O"�$�O��?I������J|�@@2�.�p��P�G8�?�����ŞNn
�۴�y�JB3 _ X�fhA5B�U�Rg߲�y2%�o������ĦI�'=b�'��U�$.�,Y"@+�1���'r��'x�\��h޴#X~(����?�P�d�x�C8 [0�x�'�G�)	��j�<���M#L>1�N�1X���W*��VDm���l~�T��<��i\�y��n���~r�'��S�J�/�4)Q���"���'���'%��'��>��"R����F��	2��*��E�Wپ����M�-	��?���V���4��l0�3�� 	#�X��:O.���O$��ܥY��7m,?�D" ~��:�n�(g�1��}��)�	*�l�'�r6M�<���?����?����?!gC�>���ZU��(�b-�W�����\Ʀ%Y�L�����Iܟ�&?��	�A�F�K � �6Y˃�A�:@��,O �o�Dc�����X�GM���I0J��,��
e��o+�7�`y�W8v�h�����X�͕'l���C>7�r<� =E��\�P�'��'�b����^����4;��dH�SM��9`ػq���a�Z�v3��;�6���d	@yr�'2���'Jq� �"yt�d*�����ej�̗�&�� ���RX���<a$���.P�*�&!aDD�:OV�2���V��D�On���O����O��,�� �a*ׄZ1A�F]�ag�|�t����$�I��M����|��q����|b�ԙH��=��EՈ3��@��ȉ\JO|oZ�M�'o�f0�޴�y�@Ȋ\L�DԩPU^%��g ;(8b��ejT�F�
ee׀mn�:��˓�?a��?��$2B1�u��w�Р���\i�lr���?I-O�m�s����	���Im�䩞�6���/~�ĠP�I#k�JD�'>���?��H㉧��ʍh�m�FN��Y.8=�.Ȓ1���Ȃ�f�Y�嘟 �YwH>$��,G��i�]�R*ĺ@����ぽ#y¡hԉ���ꟈ��۟b>��'��6��:<bV��T%M+�労g�4Nx��01&�O��d^�=�?��[��lJ�0�q�V�;��| q�͐8��!��4'3�@���֜�0�q�V;��Ԙ~�F�	�6ը�jT�N!8Y�N�.cu�Q�p����	����	⟰�O~��4�Zrl�;�fx8%�}�t�E�O���O�����d�ʦ睜fJh�'M�F���*�EC�HA�`�4"̛v�1����i$7�d�<��J��}���h��ҿ
�Dk&�l�����&����'`�7�<ͧ�?a���9�6����")��CtjɊ�?9��?1���dE��q)MQyR�'��u;�bRk�$Pj��L�k�^)����m}�Jr�zLl���kb,iBD	4od��%����'��Ժ�T�Vw��{�O�������ރ�?�#�Z�0�M��C��sݢ���\?�?!���?���?щ���O���?Fh%+��]�Rp�p���O�m)[R���؟��ش���y��)9r<Hh5�ñ}�����y"�'S�!zӖ� `�vӤ�Ѭ�A�K�X�h$IFaQ�
�� )����/���	�����'9B�'R�'ar��gH>�<���ܛl��KR���4%2b�p���?����'�?3A�5�m9r�O�C7L�v��("����	5��S�'k��<�� �t��* ���=	�'a	�	�'o`0n����^��i�4��$�6�^Y���M 	�EZ:c�,���O@���O(�4�vʓ-j�F�&F�lR����'T�=�rEF<,���z��$p�O(�oڅ�M[�i�x��`c��T\�`3�oTbmj�NF?9�����8�����^~���~� ���������5:Ҹ}rv@ҧ0C��On��O
���O���,�SO�j��v)u������ #\�J|������I��Mc���|����6�|2��?=�؂��&$1��ఇD�q�ObUoھ�MϧQ���)�4��$Zش��.W7D���`�`^�Q� ȵ/�?�/�<I��ix�)�'\��C�M�(�0����z�B�:���R㦑�F���	�P�On9v�M60�Mc7e��D�� 
�OVT�'��'ɧ�)����!��bX%�2�"3HB.m��H8�*Ph$ '�<ͧ::��DI��Hf���F�|���ѐ�J�<Ԅ��nJ��B�����T���_� �1V��
)	tl���'�2a�r�P��O��X(W�n����K�s���M�4?����O|d�u�r� �ӺK�
���ˤ<� ��J'�\�"Y�`Z������2O���?���?���?I���I�J
��H{^� �R<,�l��DMb�	˟�	W�S˟�y�����n�1�XY{6�`
��E�� �?����S�'(kJ��ٴ�yA�����萁Ƚ^�Nx���
*�y��I����	A�'�	П �I 	�浊Wkz<���iX#�"@�	����ٟh�'��7-Ɏ6����O8���1 f-y�o/�(��}���c�O��d�O�Oh��`�`�2%� o�b�x���`J2މ=^X�nZ��'z��I͟��֬8�V�)7�
8ur-s�'ȟ��Iݟ��I���D��w�ܽS��Y�CE�Y�#�O)@I����'��7�Ԅvr��[��F�4���E#�Z���C�l&��4O����O<����4*7�!?�&Ӈ���Ӎs���j¡A:��|���NL
��%�h�'�'��'R�'#jH��Z�VPD=�¦��5��ܻfS�pp�4�R�����?9���䧘?)�aǴvA�Y1�	�P���#��(A�I؟���X�)�5T�b��QIУX�H��A�e��P��`SΦ�8.O�-�vf���~�|T�t8��BR��ꀧJ+n�f�����0�	���	��SDy�~� ����O�����"LnP��Z���Uk�O�mZl��xX�	ןd����
&�/ui�����d��]P��W�F5��l�v~RA͇_����Xܧ���7-�5�F�A�O�hh�\��o	�<Q���?Y���?1����.���A+C<K����H:aD�D�O*��������h>m����MsM>�"n~_<ߊ=�ա�2q��K3�*���O6�4�ri��-j�z�)�FIxu��(�N�;' ɞ)�jE�q�_&����9����4���d�ON�Ğ�cW��SAO.x�5٣M� ���d�O��sV��/+���'��Z>U��ĳ����s�QY��>?�T���I�4'��:X$H%94��J������%H�I�9ߴvq�i>	b��Op�O��>|�nd�f��%��Ӈ"�Oz���Of�$�O1�N�#*���� z*�hP�E#���� �D(�`���'��h�r⟜�O����OxMqC�S4,7����AV2xQ~�D�O��yUz�z�ES\�K��?�'h`���D#
�41Hqj  `a�'H����IߟH�I����IM��蕾|�%j⊌�Z�H �a�9�7�yLV���O&��0���Op�nz���!��*q��kB��K�F5�����,���)擽Y�Pin�<�����{�6D�ࣖ3�0T�����<��mK�?b��V��Cy��'k�cޮ�|=����qS��ZԯڜZ��'?r�'���!�M;��8�?y���?9B�/HOHۆ�1BH�
�B���'�b�XM��Oc�)%�T��e����t)I-)<��a�+?�'iD�[9�� C
�'V=��?�?ѡn؋F0����BʢW��\	�IR��?����?���?q����O�c���As���G��e80���O�m;m��IƟL�ߴ���yE.E#~�"�A���p�Fݾ�y2�g�D<l��M�䋙��MS�Or�A���b�h��d�ʰ*�" +6����Y�ؔ�O��|����?���?���}� <���-B,���堝�A�5�-O�l5m�&������I`��U��9"�]7��ah5�V�e¬�b^���I۟<'�b>1�$���<胦��"X��RF�֯JTbQxA�7?����-T���ĕ�����D\/[_��Z�*��a`Ġ	J� �b���O��$�O��4�T˓>D�6-͗N�b�����ʷ�8-D�Y���w�h���X�Od���O���c���{N֠k0���)��Ђ��b���g�� �t�>U�]K�(�H�m``�!�ކ\G\����I֟$�	ӟd��M��tl�#%3���(�Ƈ�x���Z���?Q��1@��)���)�즥%� �sk݂l;��Ea�D���g�a��ןT�i>� 4)��M�'��[��	gڔ;5h`���YC&ô	8L��ɻS��'=�i>1�	ܟ��ɭKV��s��0Mw������"�.����\�'o�6m���L���O��$�|���ӯG�
7.^���������<!��|��Iԟd��a�)*�F�'\Sf�	����K�&� F�Rit}"�jp��.O󩂪�~b�|�[�eBƤ"��<(-�����B#b�'ZB�'���V����4CI�0��1]נ0���A�1C�F��?��
'�֓|��'~��?1���5�49 �M�7S������?I����ڴ���(m`u��O��>]��R$j��� Tz��Ny��'rJ�HW�5#hLh�W�^B��1X�#aӪ(zu��O��D�O��?�����W��wS&A��̍6B���q�5�?q����S�'R��4�yR���x���[q�ͯ]j�S����y��̮��������<��oK1n��a�q�Sv� !@��n�@��4c(�T@���?��gL	��d���,��N#1�Y��!�>���?�K>	��B�L�
PZ�C%I��ksm5}�L�J�E���Z(QI�O�Y��*Q "��4]�ȉPh�3�(A��C���'���'�r�S��d�Ҧ�' 5ԥ)A垩*���5jM��Tc۴L�,�+���?�'�i��O�ΐ2x5�`0�o37��A�g��o��d�OV�d�O�M��O�2x����!��К��O�j� ����A�/ 4� ��;wL��ª*��<�'�?1���?���?�P��5W�̴��'�ґ�%�����զ�ʰ����h���&?�	/=\��C��S�78���NO�0?,m�Oj���O�O1�J�*$�&
�X8�ȃ)���6��:�ve�������n�PqB��X�	Xy�Cɢxͼ�X���4~��q�Վĕa"B�'�r�'��O��ɺ�M����0�?�G�&}��ez�
��	
�TR�A��<���ih�O�	�'S��'����`��(;���e�ʍ�ӧˏ!Jzm 	�����O�CJt��'�O,w-F�\7"�s!iG�h��b`���yb�'�2�'"�'#r�IހG�8����'��t����lF��$�Ox�$G̦Y0��h>a�ɥ�M�I>�&`�B�H�����9 �m�'�����D��I�����O�	ȣ����񳇒�Yd������:T�~����8{*�Ot��|*��?Y�;�0 � N��;0	��#�������?Q(O�nZ+c���	ß,�IP�a]�Wڂ��%�۟d��I´!6�I�����O��;��?��T��?n`��G �b�		L�H���Lߦ��(O�iH��~��|r' �&����!GIoh�#��C�mG�'B��'����U��h�4WE,ez4aUK��z�Sc4�=�&�?��Y�&�dDP}��'c��Ꮖz~ز�P��ah5�'���%;'�������������<�bƂ�w\�y���'��@���<q/O����O�d�O>�D�O��'6Ry[r�Xv�U�wiM-�4@��i;��[R�'�r�'��y�gx��N��7ގ� �F?\.�R�A	�3tD���O0�O1�`uC��}Ө�	�O�m�'C�]��\�"A�<��I~�0`�%�' @'�d�'�"�'<L��
'N��XҬĈg b� ��'���'�U�#�4l��-y/O��d��jX��w훔K������Ɛ4 f�@تO����O�O��u�ʙJ�Z!��+�S��%�t���BT��1�Z�I��Fr�S�0�R����q�H��[�4�:s/ &D�3Eԟ���������D��'��*���8Jb0g䞕\wT�D�'�"7� �����O|�mZs�Ӽ��G�4p��pG7g���A���<I��?a���u�ܴ����
�hal�h$��� �s�f�r�]��@pa.ŷ�䓕���O\���O���O����4��y�0͐�Z��:�/�r�ev��)'|,��'��$�'V�yԡ�%?JE�2�*p��g`�>����?�H>�|"D�ܸO0��GO��:-A��B�8�tS��$�J|<��'��'��3U�`I�&�$C��� ��̦q�6)�I�P��۟t�i>Y�'"�7�*=����J�U�k��C�N+R�رe�%�����m�?AB\�$�ٴY����}����UA)����]B\�򬈖*�HQ���$�R�Y� z�d�����m#��9@9=���~(��5OZ�$�O��D�Or�d�<�|zwM��=���٦ ��&�6T����O����O�hlڄ,���؟���4��j儤����h ��/:��0�v�|��'���O%�9S����$Z9{��+�D�C��-wE�.��-P`�_��?��?�D�<ͧ�?q���?邊юD��� �׎fQM�#l��?�������13sOG�P�I��OM��F��$EС���C!H.�%��OR��'n��'ɧ��]�n
��PЊ�Y��횀��u�څ��\I��7�ly�O��X����H�� �$P�/�D��vG�X��eh��?��?�Ş���ipG���}���܋tĔH"���$��=����ߴ��'#���?1�Ǟ*( Bi�&aT6i�Nd��� .�?���m�<�۴��d
�pڜM8�Ov�+b����@G*J��ǯ�S��d�<!��?	��?����?�,��}7�#fsjq⇢%v������ܦ�%cN쟰���h'?��	8�M�;{�.M� -,4A���� 8KF@q���?QK>�|:�$���M�'��d�ӧ3~.XӰ�E�dب��'48;��B��,H�|�V�@�'ü��H%���Y]�,ؖ�!�0<!Ķi8�Z5�'J��'hXy W��7@TY���2i�~=�G���i}R�'���|�GQ�:IJ1���F��=�G�˅��$h��Q�v�ۗP���Y�����d��hqҜpF�^�x�䡃Է&�@3��?����?a��h�L��Yh/�8�#��6m�T�q�GԐ=�����ئ���ITJy�.l�>��]����׉ׇWN�`��@]�-�L�͓�?y���?�1���M��O� �֏J%�*�!E�<81	�p3� Qm�. Ġ�O���|����?	��?���(P�`�s�Ҽ�J�8ՎG4l�9
(O��o�- ~�u������IM�s�<X�'��,IW���N�ʢ-���d�O��D4��ɛc��9�サ �ףD��JP��CN�V��	�N9����'�>Y$���'���b�[$��k� ޺f�1�2�'���'[����4\�\��4N��L��c� h��E�,,>%�¢��{�t�)��Q���DR}��'�r�'ry[UeS.�v*¢Աn�M���	�o��Ɵ������F���K|���A�k_�6�1uOF3��p��b���IɟT�	ן�	Ο����,Ϋ%��SL ]� �k��Є�?A���?�G�iu2]��OIB�{��O��OH����#a%R�	�H��g�K�I,�M#�����
ƈSD�f��j��?� ������I��C�.	P�􃠮���?�*/��<ͧ�?����?�u�P>��0ط�݊enX؆���?���������H�nyr�'��S�F!Ќ���@2u��i2�"a#��|�	���Ih�)"1�G�2b� %����� r���D���Ms6W���w��D'����wU��aԮ�/�L�K)�.,����O���Oz��)�<I"�i ��H��#S��ے�:4��,��M�4�"�'B�60�I����O�!ʢ$ݷm�����X`�%���O��$�k<�78?Q�m�> � ��fy��%A�	ڡ �9�P�b�Q�ybP�\��ɟ@��џ\��՟�O&�$���#v��T�w�8(-�,���mӚd��n�<	��䧱?Q���y��?q���a}�B�xl����'ɧ�O��0a�i��dTB�Li�M.F���P�L���䔶~���'-�'|�	˟,�	�/�L���P�kQ�,�vg�.�]�I۟8���Е'!47M��WLN��O4����G� ��h��G���@���!�O��d�O��O���b/�ui�����ݎ�.�����tk�FU�5_�� ��KN��4X"�ܟ��en�*Z�,B]�J	Cn�|��d�OX���O���8ڧ�?����h9X��I�7M�����b��?�T�i�\����'q�	{�:��+�(i�>q�&��U�>��7O4���O���.z7�&?�;x��9��L�`�0e���S��4ӕ�j.����&/���<���?���?���?A�I .*%�plڭpz�Zc���d������ڟ��	ԟD$?��I�o���'�D"*��@*�4,h8�O���OƒO1���2�B'nȩ�'�ޒ 1��2-�Pq���� A"i_�e^�mWy�	jy"@D�Q����ħP>f���Ţ�=��'_r�'�O���"�M{����?����"�0���-i��d���<1@�i��OB��'��'��W�!az����\u��3B��Zl}�i��I�~6h��ҟ쒟(���@��e�Va����b��	�:O��d�O8���O�D�OB�?I�'өs�Ԛ��D/uN4������I��ٴR���.O$-nZ|�I3��R4���:����"GL�"<'���I˟�0|8ny~œ(�^��͟n�191e�^�F�*@�Eo?J>	-O��D�O���O6���!��bH�5�%Lɚ�b�(eO�O0���<��iB|���'�b�'7�Ӿ/���S�\�z뮽�v��vl��K���������)
F�W9������2(�m+1�`�������M[�Q��Ӻ��$*�$ɖ:f�i��׹ f
(k��5Sn>�D�O��D�O
��I�<)p�i�(E3��|h�ψ(��rB��"R��'�6�5�	����Ѧ����P�m�s�E)����CF��MC!�i�%��i��IQ	���O��'$��4U��1(.�E���|<������O0���O���O2�D�|�B_m�>�p�#��٨���J���D��I�d'?���$�M�;��U3� T7+�"��F#0Ia�����?�J>�|R�l���MS�'|b谗E�7!hRJT��b�'X4�yÁß�zp�|�Q��֟���l��D�q���43�
� �A���0�Iğ���]y�t�b����O����O,H�V��V��pJ&C$��)S�"�	?����O��D1�W������J��8�A�|���?d7����M޳P��b>����'�̤���|�fA`��(.p@���2*�6�iV��'B�'��>q��8�,}k�m� =��+�(WSX�����M�#a���?��b�6�4ﰬ�&&[?lg�ٰ��R����9O����O����(�27M8?�;����'nb��AehZ7klZy1D*�hw��h��"���<���̡�2�0���M��p��tL�I �MCc����?���?a��D�D�0��y!$]r�r�:�$��"~��?	���S�'m�d��(S�I	sm�<%�8����M[�Q�,qč��4��$*��<��l�B��؄v�-�&ض9b�'6��'N�O/剠�M���
��?�`��y�������:`[�8걧^$�?���i�O���' �6�_ަa�ܴEE��1�тQ�
�I��E<�XA/V��M[�OzQCR������w�R��`�� ��=a��;�''R�'UB�'�"�'d�l�/���s�&^#�~� ��Ej�$�O��Ǧ�j��"�V�i��'��-�����b���-m���
@�?�D�OR�4���vBhӘ���T�u/K�igV��%�ޚ3W����lӸR�����+����4�B��O��d�!��y��ʯvL�x�%-<�n���O"ʓV��v̳@�R�'b2^>iZ��=U��9a,�6n4��h��7?��S���	ڦq�K>�Ol��)� �
NoP����F�C��z�Ɵ�B���w&���4��q��5��O^%�%#�h|�D�䢑�!,��O���O�D�O1��˓q��v*��/�.��p��)�H�Bã�.Z��H�[���ݴ��'�H�gX�&O6<�qF�s���U�#`��6-�֦mr�%+x�6�Z�9�Dc����O���:��S�pqs���O�D�[�'��Iʟd�����	�����q�t
L� O0tB�gR�|��r��A�u�6�֍1h�ʓ�?qM~��+��w�\�8s*�_� {�&§*�@����'g�|��%%�B����� <pkM�o��	�e�L�A�d12O�-!ԩ �?I��!���<i(O- B��hR"Y�s��
\�(��'֜7-M>C7���O���
Ky����jئ0�l��Z�n����+�Of�d�O��O���f^r�$ ��eb��Pӗ�4H��O�Owڄ���m��Np�����l�!U�4���F!�ܰ�?D����ov՚p�D��?E/� Y�*�ʟ� �4>P>U����? �i4�O�ы!�41ۂ�'
ZfhK�.Ľ4 �D�O��$�O���an�:�ڒ��a��?���IC/���6��# �Ir��PZ�Ipy���8K��a� �Z�ع��.��#v��:���@F$<k�'x��������l���d�{2�֗q6a�'�"�'�ɧ�O ���D�"�TٛQo����b.��V�<�Цޖ*���k�	Ny�g@�qD��c�J&c������ɆRV"�'�R�'��Oo�I��M�0)�?A�DT�B��M�#��-Z�xi)�h���?q��iv�O��'4R�'Kr���8�T�!�EP Z�9�E��K`X�µi�	YJ��#ݟ*��l��Ӄ��TkC�A
h�n 8&K ��O`���O����O���#��0���1/MDG2��A�\(iJ$���ޟ��	
�M+4����D
䦕$�<��됌Hvb����[�	�|l� Kc�Işl�i>I�������uw�,i�f����0=ڎ���(Q�*yܜ���'�,&���'�b�'���'H@��2!AnPp��W�oP�l��'�W�p�۴ou�pa��?����	�n�T%�3������U z}�3�O��'���'�ɧ���9c�
b��.j�(T�6Ⱥg�\)1��T���ƕ��2-�B�KE�ɼ\�J��"
5?9�x���ؓL����	� �I��`�)�Spy�r�
�s����go>���nV��AT�x.|���O@l�P��I��|�3`�;/"B9�6jĳ`�Ik�e���b�l�T~�΋�P����S]��Z
:�(-�*�> 8%O�-���<���?��?1���?�.�$�C���	�~X�1��b�p�x�ǋ����ǄYϟ��	͟\$?��ɇ�M�;6g6�jq̂�j��t�����a���?9H>�|B���MÞ'׀sI��T��7Ĕ*�p��'�D8H�k��d�r�|�[��~4����-/˶�L�zr�`���M�%��1�?����?!@�L��|�a�CC�3�lta��'k�듽?a����6�����[�T2 58 k��uY���'�d@k�F��p���$��� �~��'��2��Js{j�����c+�@7�'K"�'�"�'��>e�	 h��,s��^;Y� \뵅V
Kz1�� �M�wfU��?A��Sțv�4���� �̯X=���ܠOu ��15O��O��D�>+b6.?7�YB-v��4$)
th��f?��#go
!k� �HJ>9/O���O���O.�D�Ofy���O�3#`���S� Ykþ<�w�i���$�'�2�'��O�"$Z�c���E�0�f-p�a҈$e���?�����Ş|\�I"!@�!�4�U!6�hia���'@l�Т�D�(!�|�S��BF�p������K�<_d ��,�柤����`��ҟ��[yB�j���%�O>�h�K܇P��h3�J0U�ʽ����O�l�w�	͟��Ɵ�Swh�'*�r&	>H���mp=o�J~aB�;��	�Hܧ���m �Q��0i����X*p�J�<���?����?Y��?ɍ����7^+ !
���Ah��BϾ!���'Wr s�,)0D�<�C�i�'B��#hQ�u�č'�ěqC�� �|"�'#�O���Q�iB�i����J���EibE�q�pu�V�H�����ɖvi�'��	ڟ���ɟh�ɇ6���4��a��Z�ʚ�E\L0�I��H�'N7�6����Ot���|��Bȫ	4.u���A�YLH;�kF~��>9���?�H>�O#(M�ъ��찻t��O����R���\9������i>MJ�'�n'�l���E/� (�N�+nHV�F�Ο���ȟ`���b>=�'W�7GHS&%�щ�4YT]ZSIKH(�p3��O~����?9uY���I��(ZE��oa�p�Q	X$�	⟤�GI��u���nf���Q[y��9#�Xp@�1�����ؑ�ybR���	ߟ �	̟������O�\U� �D9 !Rݳe �7K:O �$�O��D;�I�O�dlz�A ���4]�|[DOZ�b[2�{�l
ԟL�Iw�)擴%��l��<yłׯP�pi��^G���$���<��R���	v�	hy��'��K�>t?a�A�`����"\�?��'=��'�I�M�E�0�?Q���?���Ԯ1g���G�� Y&4bo����'d���?����\�u{ �5ь�y��^
���'j�:3 N�웦i-�IB��~"�'�@0�J:*_��(�G[�րP��'�"�']��'"�>�	?3�ʨ{��I8,�@mH�¬D����	��Ma�R(�?���m~�f�4�0q�ֈ�	��X�j�?y
b,AS=O��D�O��$2��6�%?�O��J��S|�\DQq��1Q(�)�o�u���$���'1��'���'L��'b�M����^��̢���({%�!�uT�lb�48S����?����'�?���]7t��x&�ՙ��8����Kw����d��M�)��K��� v�6"�4��ʟ~�l��#zӮ@�'�|�Z�V?�H>)O�$b�E[��Z�Y�E�!�P�"��O����Ox�$�O�I�<���ia�4!�'R�(`ÂPa�Dy`.�Zhb}�0�'87M �	����O����O�k�D�!�ZE:���T� )��� F27�%?�� �N�P�))���Q	�n ��%�\.-�bՑ n�d�	��`��ٟ���x��Ci��)=h�#�3j$
�"��_?�?���?���i����OURE�0�O���0J��!��>.GlZ�o(���OV�4�:"Dz�$�"F� �`��<1���m��B����$�ԣ ���ȡ����4�"�$�O,��ǦB�R���l�>KoTL{��@�8���O��`_����6j���'&BX>u{���
H��ʗDP�*t�� d9?�^��Iן�$��'W�ƴ�ա^G@��%!W.I�0�b�kFIA�U�wD�B~�O����	��'� �QsOӸ7NFH!w�(�b8b��'���'a���OB��)�MC`��< X]Km�Qb�a�.)0�|��+O�ma��Wb�	��,H�N��Np:T2�!�Y^���$ ����ɼI:]���>?�ӉHM�<��*��M�$6e6�8l@��u���	Z���	XyZ�M{��?A���?�����	�M&R�CO%M�j�@�~{�Pnڼ'Qv���͟8��F�ϟhA������"pnyp���'wB �떰�?���S�'1h�� ���<�fNM���a�b�:S�_	��D�.}��ՠ�'��'��	�l�ɲTd�Q���U�_��[!+�5Xnlu����,�	� �'�&7m�	d��?�@�4��`S�]CJ�DC@��,���?��_������<&��2��_б9P��q�($?qs�ۃcr�1�P���kp���Q �?�d�ՊE���(U�Ȩ@^�QWe���?���?����?y��)�O�|p���Cg��j��B� ���zq,�O`9l�< �XP�����9�4���yG(� �ą���ۿc�byU?�y��'<��'�B��T�i��ɳX�@i���Oq �6!Z�]���e��
m6���'J�	@y�O
B�''��'��Ԏ�2�����4���R6%���	�M[ ��%�?��?AK~��2�` �� �L͈h�ae��E�N��Z���I��BO<�|j�b�+W�X�3�;N�F��T�xl�`��]~�� �� ��;}�'��	4&�T��T\�Ӗt���g��u��O��D�Ot���O�)�<�C�i�:��2�'��,��W�Z� �&
����k�'N7�;�����DP즩z޴lf��.��6�(�	�(�`]J�h�(߬0\����i��	�|�b��Orq�����
X�zI1�� �<��Dg�P,��OB���O
���O4��'�S �҈C�*zkj4)�|^�I����Ɂ�Mä���|"��G��|R�No��A0܉_��	&���B��O��D�O�iE�vJ7�#?�Ug����В���&	˴�J�Ԫt�P���k�O�m�H>�(O���Oz��Ol����?�L�BUɛ�}N	�CD�O`�ľ<Y�i*|0�4�'�"�'���fjq�um@�8$P�M����I������	��S�Gʍ����\:Rdr�p�΍nr��ip.���ʙ#�O���?IG�,��Wr�8sԁ\���}��E�D�$�O���O���i�<��i��}hW�Q6H�r�s�+|��� d��v�R�'�`7�2�I3����O��j��E�`�J���ݰ`N�%��OL`nڢ g&)lZi~R�&p�Ra��s�i�-Z` ��"�D�� ����Ħ<��?��?i���?i-�n���%`�l�{ M$8-��nOڦ��I\�d����$?�I)�Mϻ0_N�[� �3�QQ1딍)��}���?ys�x���/
2���7O��i1dƦ\|f4bJ^�h �	�7O`lǧĳ�?��' ��<ͧ�?A���M��!��ƀ>��Mȇ��3�?���?�g�;������h��?��	��`��Q�gt�9��K�,l�4�A�ş@�'�rB�>�ռi��6M�v�I>k��YS��4� k�`�!U�r���TA�Rbd��Q%+3?�������T&�?����"i��݀w-��/�A�����?9��?Q���?��9�$� N��a�
��F!e�F@�W��OxoZ9S�|��ʟ(*�4���?ͻ�P2�(���K��f���?���?���~���'�ri���aR��#^�% F뛺<<��e������D�O��$�O`���O�.BD�U`фѠ��4�T���Z�x�`���Iܙr����&?��Ɍz�!��9:��MXr�\iEެةO��d�O�O1���(��H�2p��uʞ�(��(9U��{f�Љ!	�<1��_	:��d���䓀�Z,)L!���D�����\�d����O����O��4�8�8���ꖬ�rxxXy�2�Z
}{
�!v	Y��y2�vӬ��a�O����O��$��H�Xa"��5�Ή��j�m^�P�@H|��}R4y����?y%?��.� U#�Ʉ>��H�!��b���	����ßp�I韰��y�'Ǡ����J�#u�H9f��R�|�{��?Y��C*��e@1��t�'`�6m1�D�vF�uZ��ަb>}��G�X�p�O��D�O�Ɂ5=46�3?����z<�2�Y*k��pT�̝ P�G��|&�l�'�r�'?"�'�z���D��	\h�؀eȸ1�h ��'srT�@A�43�y���?����)
]����k
�
�I��G�*�	��D�O2��*��?� �]��˹gRx5��U�kozi�f�x�Ƥ�$j������$�~?yM>Yd�ξL�"���ڰbg6�a2�X��?	��?	��?�|�.O�)nZ�R�t4��M�"E�fyC�Up�0�[�hby��n�p�0y�OZ�$�"iE�!O�21��ɑ����q|r���O���vbӲ�s����̬?�'y;��q�C��z�X�Ҧj��yR[�X��ퟀ�	�4���̖O{n��4͐(<ܼ�'���N�0(Spcs�v%i%�OL��O�J�d����Z�r�� 9A|���PG*^���	ȟ�'�b>H�d�Ѧ�͓O����U�ӗd6��p�'��h���I�ݾx��O0�O�˓�?��ww8�ӂ�$I�T���B�q�(�����?���?�.O�mڞ�N�����H���>@1�+��@yZ4�^*OK��?qdX����ɟ$'����� m���b��qa�e��.*?��/Β0?L�KCA\|̧9>F�]<�?y���wƊ|�'�S�
�ҜC�K��?a���?���?a��	�O��pw�L�OP8�5�תȪT��O�O\�l6���'�r6%�iޅ�eMH#���� ��&;Ơ�����IƦM��4x�8���4��ҝ#cx����lBj���J��:D�	�!�Z͈�'�4a1�lF	t�@�@a,׉Fb�9�����>$��
�
m�e%�>}0v�QՏ�R�����-V��aLG(k�p���/�<��z"�
�d
w�q� �1�+2h�'C̸�Ƅe��0I�8gp)��M�lA��AgR���س���5{^�ĩ���@NEڰK�2O ��&�J�p"ur"��:��a�!OdTQ6��v�t
� C�E��R�Ck ��Wς�V'X���l1I�G�VP�e`V?Pt��dI��\}�iK�e�f3�-�H3p�蘀D([�M���?a����X�(S��6+\�@D�U�� "���1�M����?�'h���'�q�x<�d�+H� 94�Nm-0�i �i��h� hiӬ���O���� �'��I�$��i�B��$���#�щy�
��4�@Dx��)�ONdq��T���0�I��v�B��NΦe�Iޟ8�� B�4�ҩO���?��'m����%����)�3&���	�}�$Iu�'^��'MB�� �̛�A�4*ŀ'�J�}��6-�OR�`�e}R\����w�i���
���6u`ӦĜ[CxБ��>��\����?1���?*O(�G�Ŋ!�=�7��|#�q��d�-Dʡ�'��ԟ'�L��ԟ�#�Q2y<9'_�W߂4z��%�c���	͟8�IPyR�عo���Ӂu�t�(�#�9b	F1��JݝK<�6��<A�����?I��r4���'h�U��/\?Vld��ҵp���B�O��$�O��$�<)R���xB�S�P�a�]֚I`��ֹI��5öM��M������?���=9 ��{�F[#=x4	w/ɺL$@��%O��M���?Q/O�P���]Q���'w��O%�P:���;ݢ�p�R,9XB��C@9���O���ݩ%�t���"*<��pk��l��"��,6o�gy⃊*�67M�O6�D�O��f}Zc�hC7���i��"��JJd`|�ܴ�?�zO� ����i�7�<��)@ʩ���0盦�ՙu�<7�O���Od�IGg}2^��(�2s�NS�(`�'h���Mq͖���'o�t����MTٺ��g�t��(e��n���$���0J4�������<i���~r��	/�`���Q�"!�!�RI� ��'	��rd�|�'��'�&���cț8� -Q�*�	���f�p�Q.9#���'x�I8'��؞_�p�	P�a�Pd��&&�"�w���M>y��?i�����\�Sq�����*gֽ{q��o�dy��P}�^���IK�����I=L��$��F�����ڙD��ѓI�`�ٟ��I�l�'�h�bT(o>��5�Ľl��P�G!؞)��ZK�>I��?�H>A-O��O�X&�H�C�6hC8�z�0�c�J}��'��'Z�ɺs�@�[J|2R��3��9��E�?j.f�[��Ƭk��f�'��'��i>���Q�	وA�[���*%ܠ�a��Bd���'hRP��ɂOĚ�ħ�?)���j��Qqb!!!A�Y,0'��k��dy��'������uW����0� o^�z�x��c�M�*O�!���L��������	�'4bl��:�J� �� tJ�a�4���OX��c�H�s��]��犁?^l8J��>�^�b��i���9�kӞ���O��⟌x%�擕?Q���Z:$�p`�!T�f�
۴�?9���?1L>��y��'��}(��<	��Pɦ�L4sLCal����O��d،Qc��%�������wK�0%`A;`m)`��X:²�ڴ�?a����dV��^>E��M�&k��(�,!��K�e~�P8&/
ݦ����c�~��'K�ꧣ�'�\�x�Ի]j�Ea[
u�Jģt�+�d	k1O��d�<1��w�Y���43���נ YĠ�S"�5����Ov�d'���������1�d��VOր�ЋI�/��lگA9lc����cy��'�,�)eߟ�aJǖ3N��=Zׇ��������㟨�?y������g�6��!e�h��'e$^��rL���?�,O��V�:�"�'�?񤌕�/�Ve) ����}*pEJ
uH���d�O>�}T��%��უΐ&� �0ӫ���q
5�g���$�<���!2���)�N���O�����1��!�&���
@;Ej���x��'��Iq.�#<�;�� )ឞpވ�3DB;K&��'��U!A��'t�'/�T��=� <����Q�$ ��戒�G�|���i��T���@,�S�S�]�]S��ì){8a�P�?L�6��2x���$�O���O:��<�O\�)��%G�bH�͑�7�z,�A�>�-�G���O"$ǚS�n���N�r4���Ń7Q�6-�O����O؍p7�AW�i>��IC?���f��`���ߤK���U�TԦ-��]�I���9O��D�O����2(��;��N�.K��;CKOf�lZ��c�F�-���|2����Ӻ��oؘx���ЧF
�����gI�ߟX�'���'9r]���B�6�4�3c�-#�.Ub��-�"̨H<����?�)On��<��>&�qHe�=zF�@������ioZ��\�'�2�'�bU��X�����4��$=2��S��w
�l�t����d�O~�+�D�<�'�?��g(_�ΰ��ͨ
��@K��V�pˉ'%�Y���	�"JDQ�O���U�1��� �	ˌq��K�~�6�>�	şԗ'4r�
N<)��#U�v�[�OI.J,${�J[馝�	��,�'+0Ux��1�)�O6���f���L��Nc��h��H;|�~�X@�x�^� ��͟�&?�i�ICk�*ehVx���#Ҥ=�cp�j�]ha�im맴?Q�'r��	�:q4�A��7\ ԫ�&��6�<����?6��$���4t��,)�돊e\,՛�+OR�m+;uxJٴ�?���?���4*����eɕ���!��
g�䅨G�]�%��6͚#S|�d�O�����<���Ax���T/|�p$.:ǰ�cR�i�B�'����/t�lꓯ�d�ON��3#�RccnL�Yb�R'D�7�On�d�O4�+a>O�Sݟ8��ϟ�KՈV<  ̝��[�_������M���3Nd��[�P�'�^�T�i���M���l�O�`��e��w�����ya�<���?a����$�3t��yg�0^X��h��׊]$d��Q}�\����Ay��'�B�'�,YIf��S|�2��<vc02��'�yR�'�2�'��'t剂\��O"6�Ӌ\\� �p����4���O^ʓ�?���?IA/�<a�MXo��I�2"�'���PV������L�I���'U����~R��`-ʐZ�I�
)uj� ��دFxLl�t�i*T�0�I柬�	�jP�	b��4Y0�x!�HũL��iHq���61�-n֟|��py�B�����'�?������E�?p�Q�eÉ8i�)sG- p�I�L�������Bn���'eRџ�]b��.�BP��1��a$�i��ɮ?�BȪ�4�?)���?��'%��i݉ʳ`�Df6����Fg���� j����O~��?O��?ٌ�t�X�?����D/@�h�f��M�bꎿ(���'��'�����>�,Ojآ�įc�,����T?�q˂�Vͦպ��y��&���j��������0�(]2��l�6�r�i���'���_6$듰��OJ�	
u�D�؂��(`ĺ���1N�7M�Or˓[Ƅ�S���'���'�D!zÕ�BmH�P-\
�4��'n�b��]!6�P��'q�	��'pZc�z�3���k%�M��f  68��Y�4�y2�<I���?)���?q����@��y���y���2_�>L��Bv�Fw}�_����Iy��'���'�P�RТ:� 1:���;1��/��xc�'���'�r�'"\�p	&����t�T� {H����!Oy���%��-�M�)O��d�<����?9��e^������e�P����Θ V��̢a�i���'r�'5���}c��z���B�E�\�h�<�Y$�Ѣ#xzP`�i�"\���D�	,&���IП$��8�R��U(��HK�$�#n�$hm��P��Vy�lߐ�'�?A���bw����%��K�%]
��HڿA�I�,��ϟ��F�e���IRyҟ�ɻB'�%�$@�̾e<њ��iV�	"L�a3�4�?���?��'e�i�[tNY:�0*蓚M��- ��r���d�O&t;�8OԒO�>i!6�"ecty�4���C��шƮqӴ5 ��V���韴���?5ѭO\˓�ܥh�*̜;T!��e�4y�����ir����O����OF�U-p�PU�Sə�fIr�2 �v�6m�O:��OĜ��n�R}RY��	~?��Q&;u`�@��,�������1��Ly�'�yʟ:��O��Q�O��(��M�o�@�%+\`� �mZܟ�Cv�6���<i����$�Ok�I�S >P����q?�0#.ǓA��I�i�P�IXy��'��'`�ɑPG�\�1d˹j�`AD*��e�}����+���<����$�O&���Op
e",)+� B kZ�7~6��1�k=��O��D�O����O�ʓ=�� �9����f�209�DWY���ˣ�i��韄�'���'��g�yZc��E�B�і)��4�q艝@y�q��O����O����<�!��R6�S��@�b�ܢu�b�#NO#a@z��R�H��MS����$�O��d�O�$3O��D����˽}�e���7 ��褉|��$�Ob���y��U?��I�� �0/��HB����o�L�*� 	����*�O.���O��d_6E�2�D�?�If�C-e���t?K�l;$gc�n�G�h]�Q�iB��'d��O�l�Ӻk����Os`�4��C��@��6��Ob��V�&���On�$�O��>���e���FܘBхoE ��t�}�D��G�Ȧ]�	џ����?��}�eޭg�����%!��1�Č�l�7�P�0X�4��"���4���5t���$��*���1�K��M+���?!�1e���%�x�'��O� (���֟&�8��J�>�����ăy�6�OD��OH�D޳?��us��@;2	@Ǉ�AR��n���*�MG8�ē�?�����fh]:'7�I �� OZ"8邊�h}R��yBQ���	՟P�IEy2IM4vR��B@T�B�sv"M�\=j�J �D�O��d7�d�O���$o��s�	�Tk(� �"�3���I�5O���?A���?�*OP�!��|Rw�ʝ���B�D[�
� �A%�]}��'���|��'�Rk�R�η"Ȱ�Ǥ��x<(P�r�\h�들?����?I+Oh���E�3,���R�iA��e�Ѕ�~�*$ߴ�?iI>A��?��H8��'�j(;@@8ya���N�H�ā:ٴ�?q�����b4D�$>�I�?i;񠅎[�Z��%D�-,n��V
с����O��$�O�q��3OޒO���OU؁K��)����W1^��7��<��%K���F+�~r���כ��(�l� �>�YU�ڽ]�}�'�xӒ�d�O��V<O��Oh�>��Fm�;/�D��t�X�q���j{�Ra��EF��������I�?)�}m�9|�I�Lr�`ѢK�#�>7�[�R+���1�'�S���M�"�uR1� %�4��t�U��MK��?1��A��x2�'�B�OZ�R-B�n�^	��`�,Hnb4�7�i@�'��\�o&���O@���O�T�6MN�:�Xq�E���vViA���Ȧ��	����O<����?yO>��H_���rϑ��)e�^���'x
d{��'�	֟��ٟ@�'��Xʤi�;4j�ڃJ�U͠ xSCM6Lb�c�P��\�	�T��$Z�<�0�QzG(��P�5RI q��ʋß �'���',�O��D�k>uʐ�\����%���Ph�>���?�M>����?)ZeT���H`Z a�[ x�B(6a�$��'��'72Q��*�����'HJ0�"䋳LݔD�U3$�NH��i:��|��';¢|���>1CH���s��-H���@���u�I��'H��+�i,��O��I}��8�Q���\6�%cN�$<%�4��ܟ����Y����d�]$lꂬx�/\ z��X��o�<�M�,O��b�%D��y3��R�����Y�'����#B�@���r@
$u���خO0�$XD��#�����<���ɐ�Iz D� ���qܛƢ�8��6m�O
�D�O��FZ�i>5!$e^1K0�%*���/qS䨳Lͻ��d�O��b>��	#KI�%r���e*�E��`^�MXz�P�4�?����?�dH ���?��IO?9�/��d26M$Q�X6p8b���N���ħ�?1���?�D���.��阣�Ψh������7���'�B���2��OD�D'���(��M��'�b��4IXu�Ő�R�����>�Iߟ��	����'���`�e3# ��%#ۋ"�@����6��O��Oh�O�$�Ofz�(��	 �)6uR�/ƨ��'�r�'��	���3Ͽ~�!�7w7 �惕�Y�l���F�̦���0��a�by�m^�5���=��p���N?�����T5f�F��?���?���?a����	��8;� � ���c��Z�H@��
e���>���O�ʓGJ-%��K���.cA�YZ���Ȃ�fo���D�Ot�;�v��Ɩ���'6��⍑%�YSCE2}��@Z�^
��6�5�ɚ2Zv"|����	�㙒DfF�ؤOK�a�tuAMn�|���Ov�'��O.�d�O��d�����H/bD,4Z�M�*"%
�ɂ����şb��;~�b�b?u3��tfY�h�J*�F�M�gQl����'sB�'�b6��b�F1�⣘�V����u@؂7� 0�ش?n�aFx����O�p97k�,oYft�A�0��� 4���9��̟,���C�p�O<I���?a�'�^�:�ŋe�Fz�ܹS�\{�}b�T��'�R�'��D t�"�8Rg�<�d�*h~��J�~�`���?�+O���?��S� ���J K	'(l�*���;}A�h�'�*	I�d�����O����O�ʓ`U���՚Ɏ,�f�*U�4ܹ$�ڟ'}�'�r�'\B���������q���b�@ɲ=�h�b�d�ON���O���O�����O
�%�*i�0�tꑰ|F"xp	Φe��Ɵ��I@�Ɵ��I�8��}�f�ZdJ
� {b�0īɰbPK�Q�`�_3��P�sJa�ȣ~*�@A�Im�I��ǔ�"��Ё�Wk�<�eW�-t����QN�ȡ��~?!P�X�i�������u��0�%�QG.:v�P�,[:�8��&ӡ	0���=S��ے�P~M����4@9����]�`&!ܿ5l���	�L؁Cр8/�3QW+@jm�uFZ���Ã^IPH�Ae
�t�:�BEOn�Y��_�&*����\��E�'���'��l�9�� �0!�u�N��E
w���"8(v��X�c�N���ƘϿ��C�'�V-�e���J�j�t�B�@�40ѯ�:k`�Y�')[�v�.t��gN�������;b]��q��X��
@��6)ȩ ��/�?������$�|�KN�uzRp�O�&U3Z�ӭ�y�痆(���ƅJ�H^m����OB�Fzʟ�d�AY.�JF�$c(�\�)��?���9[�X�c��?���?�b��.�O���49���i��Q�sI���R+����1ΙH��	NI�1�֟ў\Y���:�:cM�bּ�`�G�?yu/0���`#d��<:��3�S�? 6M���ʯ(G�|�qk�0y�L!���OpI9�'�r�	ey� ��6�n���gS�O�2uCr��y��Yn�3`�S,�z�a��d"=�O��1
�(a�4,6�T1�䉟|�(��!���/H�����?	���?y��W�?�������-ɜi@a��Jg��*�NF
]:���(��	��w� lO�#tF
����O�����n
r�T*K�*i�P��IJŮ��ߦA��bȩ
�����oԆ]焅��M+����OL��'-��-�d/�>E0�ɠ`J-�$����R`�$����� �
��hΓ]���Ieyb(D-.��ꧥ?�(�2�ґ�S?�r�[U�����)��c��$�O���Y,7�0UI�I�/��\R�O�:.����E�5�T IW�Ԣ�Т<yS�Ù-Tn˵!��q�(d�Q��~����Tz0�x���I�,^f���O��?}h�MW�X4}�rJ�5���h�{����	/Me��"��H!b�_1���3�'h^O`�c�N�<@0�����|�(��1O�ȒGy}��'v�U��A��џ@�	�dx�h�J:B�5(�/ڰ)���ʲ ��ଐ �R�p���S�D��'S�-:%G]'�0ۖ��1p䠫6��i
�psf�I|��J���O?��[�j���?���!��߉�����O�$9?%?�'�|/xR(�Qg���RU�c#�m=*C��0�6�J4�-3�$�����<�2"<)b�)�
Y��>�b�	%�֨:¸8h��ǟt3�,h�T9��ʟ�I� ]wBr�'�X��!%��8H��Tޢ:�\		�'$�Hh	�xѲ��M	>p|�p���)l���K+6��c�6ӤY�3e Ol�quaL��L���@��* zA��O֐3���O����O�Y�d�Iy�`=q�Bc�K��"�R�
��xb�'V�xq%�5h���AF�2��<y��0���ɤ<ɔ$�?)��&/Gq��*���"}4iba-�i���'���'ntКV�'D�8���[��'��,�l���H#{$�#�/���p>vh�cy�L��A����߆�ʠqC̸�p>1�"��<���i+�AR7*X7�<�QV�j��'�$������?�O�ڭR���`��p�@#ƉN����'Д���ƭ53�,Q�&�~=��'q���hO1�x���n�GP�!�V.bA*i��"OD����"/�����vQE�s"O��1����<1E �>B�h*0"O� � *>w��ү\=O)
l�D"O6T�۟�xqiwD�&"�8�b"O
��@O8]P�"��4I�v"Ot|�F�PaV�`���7|q��"O±94+C�Ux�ً�n�\*응A"O� У
:.d�k��@<`��"Oz��H�{=�3m�����)�"O�D��gՠx٦H�w�8,�2�E"O`m���tRd����!/ڀ�c�"O��r KK$����L��� 4"OP��0b�57laТ�Z/v���"O�}�W�ѸdQD	�w-�O/��["O�ȶe���2��1���k!�Xy"OrTz��N-^����u ̩f"Or���͗;"�D�TK�K��(h"O�t������%C�JCU��1��"O���h���z0�u ;;�:�@Q"O�!1Ǝnq���>D��qZS"ON�
�
-	f`��T
�
����"O��V���$�����vdVh�"O����$P3��`��0��!��"O��(��Vw�>�*��	�3=\�)�"O֐��
��H�xr��')���v"O� ;'��!�@�vn�|#��ځ"O��bF�ٟpF�)� �� 0��`"OBev�Z�/�����Q�fL��"O��4�3m��U0�%B=��<�7"O�I3�*�؈��͆E�Pa�"Oj�hqEƋI�����d�
Z�(��g"O�  ���#�5k�I�7b&HϾ�6"O�d�@�"��|�#���`XWOx��IM("�X]J�J�)�
+�ĤbB�'���!V)%��(+��$�P��	!��k2�f~Rˀ8{0�&jH��0���Y��y2�	_$��wCУ��]B�OD���
��}3OE��0|BE$JBl�83��N+\B�-��`��c�y�*U􂍲sI��&�qv��e�	��6���O�q0�!�@�(�'7����OV�ďOg�f����|x4,)��N��T1�o'�Or��ŉ_ SvRV�����'~B9K֥��	5�|3�ɏ4%����t��`�^B�I�B``Q�AO	k����k�*�:�O�,�k�.�*��I�v����kF8/Z��稍� !�C|UR����βq�ڱ.�*�ו|2.����,5se�_-bN�+��1 �Ƒ�Ɠb�~!6��,?!��6T�(�)��f{Z}�
�B���!!f�><���!��|����	�:4����]~2��#�Hȓj�[\�bӋ���y�= �r �l�To<��b�����'g,��⯁��0|���R-M�\0��+��IH��{�a�l�<���)g$zu��#��٨l���}�<Q����3����]��iU|�<��ɕ�Q�`!�g��mH� ӷiG{�<g�nX�� �ÇT^04�t��!��'u뚉�%L�&��0�y�!�DM
ڊA�dƐ�df��bB'_�!�ԍ@^�L�R�2]R��A ���!��G�EAv�)��H^�h$ۧ�ƻJ�!򤕘2(L�( E�M�<�IU
fz�'�,�	�-<O�T�ɼk��ň��wb�LA��'��Y��1_F\�qH��H���ܝk�8���x[L�`�`�ZSC���GbmD2{�a�~�P	�	_��ۦ �|��c��|�<���J2`k��JrƘ�.����wy�+�g��(�=�~RC-ɛ&>�p
E�G�7�)z����Fބ�k�'8�]@��yK洊6Ø1�`���y�Ù3�p�5����$�	���/-�t�k�k�f�x�"O*@��*
�+B�әI��K���bҌK�w�c�"|B���14����K/d�d�Bc�Qq�<a��X'"��aP�E(\0���]r�� �#�Lp��s�`�&9�eä	"u&��5��1ehB�~���ώM�(��4HK�����O<�I|���G}"*U�<����<N��+�����0<!�Ǡ<���<'�� M��FP4��!��Fצ���`�����×>�Z�b����c��J���/�:}�Ǣ�
F�x��3�ɉDIN�(�	����zy�� j8|x�A8kX���1-�|B��+/�BT`ݬ~�T�#7AXs��ͳ�*�O���GuӶ(���ߢY��d}��!3IH636��/)o>$�Ї�{0}b��	�����;X�N�zp���w�H٩�� �'�D�d��l@@�+S��肬ۧ]�6Mk��c��	{�t��GکRI�c����$��"C漲@/�gc�A�c7r(r� �OY*5ņ�{a�NeN�9��?��щ:d8�`g����E�-;y]ȡ@���:v���ۆ,LO�𰆨�\�`0��I�d�L��/+���qaڜ5�E��x�	<�49j2���)~p���4yV����

w�ո�"Q.U���E<�-�/X'00:���#���R���r}��١v��7��~&��	�S��f���Z�݈h��)��[:�-��HU�/����d	�*z}�oT�Y�ᱠ�|��6�Xp�1d� >K:��e+�Oa��z��㵨�-<v ���?j���c��M�:����Q!�O�!(���3?Th���C��^[7\�����بF2h���I y�i	1FH�&^��f(��h|�S����0=a����J,���+G�AjШ�v�N�ԥԢ{PΡ�v,�F*��'�݂p
եC!�4kR�O��@��W�>�y��۞rpP��"O�} 2@ڜ2�j)3��*���A��'`��	z=s���K}"��CZ ѨF䁛]�Nj��B���G���0䙋A�'}4�%�L,B*hQa$d�V�d�� G�&�f\����fV)�'̺͢a��Q�b�>�`�*�{
� �	a+ѾPZ��g�ǂmSh���	��d2�F�=!2� ��ȯE[��e5�ň��w�T��1Ɠ'8�MS2�A�H�x�AE�]sa{�)3B�5���N0��R��db03G(�>���� 뎹ou��C����fy;��P''����L�dc�5:Q"O�qk�(>*�s�	�$n'�ѳ6���XR� ���$p9�����y����]�D)���;NP��p�+�	�0>�ϗ�LQR�E�C�����п������U	�O`3����]*"` FV1� �����(|�%1ÅiǶ�!���S��p�u�x�(Hf�NR�lG(+?���&@q:d�W���Da�!J�`i ���F*=z	ߓOQ<�AA��Z��q�/� �����9T�����#P=W{R�bY{ħy7�$��7Ě>$ʂ�ˇjɘ�y�m\9L��$�[��X�2�:w]�䒏�$�)��eC�8+ߦ�C�6�L<pE�8!z��D��	0��Y��'�N��"h޺_���㣍}����A!'��=2������EO�
8/.��a&o��v�����D�2�,�@fiU�z�"�B�:>�(QCʗ�%��X�,u�@��O�)�@�=��
�( ��&#ҋi�2��ʓ:.Љ����+G���$��*�L��
.�%��1~%&�yû��I��R%W�����?��|�;L�I��)�%=J��3,�B����3nqŭ	������?��0��ǟ��U�۹�~��u>���\�xx���o}B Ǘy�i�Ũ� j�|��פ�p>���"��m�0�E����`j@2WG�*C)'iI4�i
��� �';�,0䩟23���Exb.��|���Y7���[d�C�M;��=cuxqđ�f$��/S���'�04�ذ��L,z���s`I]�$A�<���-��Š���G��J�3
=�7퉛\��q1O~λNKn��VΕ lG@��F�Ζ7☌��I;i��L9+Oܺ�ȿ�Ӳ��bن*�	э[���R6&�ftF$��8�S�?�:E#�mGE�	�F̪d�%�X18� x�c�e��L[!̙��'����2J�A�0�f����N���/U�i�a��f"y��ɻE��)yR��f�4Og�y*��-J�qZ�M�6�N�2g�j�"	�"�?�$�]@dP�MY�:�����曮��
��>N�����Ȁ2`[C�<4�t�G]n�Q$�X�v9�I���K��T�a� ="�$k����(;�u�O���MS5�N�p ΐ��ܻY�8�ء���p?!�O�X�gQ-]M�Hy"�P8@A���S��hL�1U� ��PO���g��%�h;!�3y���^?Ğؠ2�'�O�yf��0^ZNI����&�p�g,�;r�a#l��OF!���J�}�n�� MLG��9c�ɖ笍@���X{Q>�A�&V�|�G�kn �c�=D� �Ys�jH�ǫ�v��pa�,Ѐdså�$:<�S��y�%~v|dJ1jBK�/3��	���V��7`E1Y���E�lu�9�V5�1 �a�h����vT�4�K�X>��oL?T<a|���;�ꀠEg��b��4����xq!s��j�'ve[�ªs��(���iŜ����Vw��2,���(�\�:��e.�p ����Yk�"O��y6(}|	� NK�(��'̼'�P��cɇ ��)��<��#J�lD�KBn��{� ��P�<!�(,ƨ�s�דn��S���<�j�:{gx<�i:\O��;4�ƻT���v� �-�����'��m[s���O���&�er�_Rld{'���y��7C8��P��\R���r�&Ę��'#��5�83_�
�K5�'S��8v�ň5��t`D���,��_�����M�}��{�-�\��a�X<^_t��!�'^@Тƕ_���D�=�*��Ql�1a�d�*��[�n`џX�Ԋ&ʧ�xܳ͌t,0I���+;��ԅ�+Q�IB��T�����^�$��;!N @	��'����H�<A�%�I��u�T�Nu�寁��b��G�]a���L�*
?>͂���$?ބ���/d�0ʆ��41��dC�"�$L$��R�K�Pi$M�FN�,�lM���E>��O;xT�7��=}2J�ˤ�A	�d+��3ht�WJQKf� *5m�)L�j�@@�ݗB%��`n�Sv� ���D��'���{�f�%�HA�g�y���S����Q�Q>�ƌ�E%�0ˣ�(z[�A:�,(D��7�ɪZ98�)DX�qf1���<���{��(�����FK�(V�5�A@̈T�2x�"O���U��%)��ш2r�t�H`�0v�az
� N���L�R�;��<I�H�"O\�b�n`^�Z����7����"ON�æ�L��Dq"B�Z���P�"O\�J�dB�LT8�d�"���"O.!s�(
2p�� ��T3�:�I�"O�iP3��*�Py�bR��V��""O���K<ā�pB�G�j�H�"O��A�H�&�m8����-�H�Hv"ODI�¤�>>�� (#��=T�`hX"O�[�C=_e�TZ�ŉC���'�Z��m��fK
Ę%J���`�
�'1P�;�
�`���������	�'�)��8 �Lݩ�FT�u����'��ѹ���U��G�A_�e��'wqC�οd�T91腩5����'�����I�<��%;u���#蘘�'J��U�" C�	�7-�.h���'$$����'���Zr���?B����' ��9c̝[���
Q�8{����'�b��U �4�1�a�ʋF�<�
�'�R	 �jč([�P��f��Q� ���'�p(�J+9�QQ� Kb }:	�'wN�R�f
<_T�nL$H��Q	�'-�)����ܩۦC�W>��[�'k��ZU����t�F.�#@C>��'�r%ӥ�-7Խe+�58	�0��'Dn������`������5;@x�(�'Dt���AL42�|]$�ۡ
�t�0�'�$ݠ�C�6���cffZ8oҸ��'�2���ꆹ ��z�(Ře� �'�B�`��B��LX��fE����'�q�(�:HP���N ����'i���@ V��l�I�(݁o'����'H�- 4�G(0ΐ�f׃� �x�'+`�+qK��Ѻ�zv�Z0��ia�'}$0���̨�F��r8�'V��� <Pv��ʑ���R�'���G��\i�P�#My�v���'�$)�  ֈ4���j7�	3�'�&���H��`�7�^�&�b�'o�� �3�h��`�X���';��Ѧ��'�`@�DP���'2�ds¤E�*j�䂤[�Mi��*�'m~�D�H4~�L�ićB���y�'��H�ᬈM�-l����)��'AnH�1Z!X����m�)q2�'�n\���D9O�dh�U�%W�Q	�':҄)�ǘrA��"��o�F��'�`��!¶���)V�^H�E�'�e���+m�j�*�
=P$��
�'I*��b��L���)��G��53	�'��E¶�+W�\��%PjB�H�	�'����E�H�%�T�\��`	�'����K��剕m�2!4 4��'Z� !�<:x�25�օ& H�'ov� V!�*m���3������'H�Q*ؒ	k�MHC�C0||~1r�'�&�*�'�hu�(�%�q L���'��qA�BefJe,��	�'o��i�I�Sh��hĦ�2,4�(Y�'���� ���4]$+_�d�'"^К௜�*X�]!��Z)��'��P¥�(��!k$i�|F,|P�'_*p�T��+A����jʕw*�J
��� ��:�OZ�z�T�%��P�����"O��)ݔ8�
a�b��MT���"O�9���X�Iob��3B�*L�h�"O��z�
�B&�h3Р^1=K6H�p"O�¥��=,Ґ���
Q-�IJ�"O�)�6◽Z\���6�ۤ2G���2"O2Yx�$Ԗp/�E��H�%@*�q`D"O�\�CcY���t
��2ݠ6"Ox�X�@� 5���EH's����"O�@��G�C� }R��I�.R��R"O��kQd-�(u�pC*bv��"OhDh�� a~�#�ǁ7h	
4�4"Oxš%	8W��c��"�� ��"O��kH�h�8X*F	2=��}�C"O��g��`���s���%7p�!"O(�y���.L��z���eѼp1T"O��آѡ�D4�%�+��(�a"O,��ǆ�Y��L��Z"O~|A�B[�Xh"�����0V"O���v0�)��.(� s�"OZ�c��T*}�#����� �"OʰX�%ֻ=��]A�Ί�3{��K�"O&� ��� b�;F0�ԍQ�"O2@�d䂒s:��z�Y�L��� "O�(�6�AtQ0p%Z��EH�"OJ����\CM6� �m.}n����"O4U(DL$���
�	���"Oj0A�Ɍ و�C`�%����"O��2d�xF������i.T�"O��)*�5�fe�eKW*���s"O.�	��U'ZL��B���-{ҍa��I_���CeB7}����%i��H�z�+9D���O/;�69H*$<��i�l8D�(��sb�H�V�[D��d �m D��
1��-y	XQ����VJd�#@:D�Ȁ�
������&�7Yh��c��9D�X�,>�6yb`��!���+D���Р�[[Q�a L@
�@�B�<D�D�$NE�h!  Ó/N��m�`8D��i����Xe2!�`���b�0�Ԫ7D� hP ��o�XD�VI�;fn�I���5OJ#=�&ơBtJ|��̘J�m��\L�<��
�X���XP�n���8bE�<ѕiB+E��P@�1*;��DB�C�<''��n�uJc-�umիb@�T�<��C={�!�Zir����P�<9MҾ�0��i8Q M���I�<Id��"[PEHv��2h�����F�<�f,�D�h�4�أ-���j���B�<)�l�4ːL�m�]�x!��@��<���?<�dRD.����(!��~�<EC̯O�*���	������|�<��"�$��9ĎTжDBL�<�A.�8I-����`�7s�]�ML^�<a�Ȅ�"x���ٯRG�\��gM`�<1�������7�ت>N����m^[�<Y��{c@���ì<E��áJM^���=��Ð9��a3�C%rcDP�hb�<	0l%_@��u'Y!�<�I5"�_�<�E�Bv��x �m �(\9�)r�<����jȆ��b(4 ,��Dn�<�d��e�$�1l|�̠��j�<!��� 	���2IQ�B-��Z�E\�<��ԯ7�B����8��!"TF�^�<� ��i���r����' ��(�"�yC"Oꔀ���-�dx2�P85���#S"OD�)��6M��yr��tv����"O�5�&"ɕmFH%�bI�3t�z�IW"O���CE����J�F&p�B"O�#w��9E(����S(�3"O��H�/ڷ�q����(�Y �K>���X2��� �Q|c8eG�-D�t����i�v�xE-�-H֩cu�)D�HZ,R�3�F"HT����1f5D���0ǯjZ�<�`F�-yV�M	O������4��d�k����+0�fB�I�"��DPGǫ��T�99-B�I�b�����)\�RO��Ci�0�C�	`rǓW�8�{��Z�R����:D��!䈟�aa��9s�٧t���<D�ث��;�`h��ևXo��*��&D��0Ce��g��ҥ��Zzt��`c!D�A`㕃o�6�����b�k��?D���C�G��%�BL��#����*D���`E���E�5�*\Ѭqp�'D�x
c��<w6й�OD�t17�%D�ph7ɚKr|�������r�e8D�d�ۇTd,��@�:�^��֡4D�D9����i������Rk*���o2D��V��0F�<��T�n���y@�;D�\�o�)�ظ�Ȗ+Y�����%D����rDm��͔�3�����%D��+���M��A����l[�F!D�
$$�#�=� )��T�Y��=D�ġ���O@�m	��QVv%ځ:D�@ #IB�l�\ ��d�5N��8��7��p<������l�m3`��j1���<�bD�˘!�h^4.KdM�y�<	Pǁ\�8���hq��Sj�<1�Ҕ;^�Z!"q��"�Ai�<���/&�ek`
ދ;����db�<�Gm�cH����J�L���hH�<�4&�=}�^h����<���y���G�<	��B:��2�� �,� ����~�<!EdR����q����T�z�<1ᡖ0t`��DZk�PD"��A�<�A���k���bFdeA�1z� B�<ɴE:9���K2�	([�4)��l�B�<Q��S�;6|Lڅ"ΪG��a�FS�<q��(����F�Ü?����b�U�<�Aˌ�b1���ƕ�x9f�E�<�g�߯X%��p��G4y�
L�<A��] ��ǌʈV�p�ѥ�J�<�6��'��L@#��'� ]�VEQ�<�ul˧'|fX�!L�0r�`���TA�<a��Q�y�lQZ��R�N@�<�];4�U�e���qH�~�<A��_�?�8;���t�ڔQ�Sz�<9�OX�3�v�(���JI����x�<��nы �8��1��S��I���z�<����H���r�Aĳp��u��BO�<)"�k��QӇǟ�t�(�+ƀO�<�`ĩfsZ��b�����]����P�<9e᜽}�P����M&d��E˧*M�<	�T�*2vH�:]�dԂ���Q�<�G�+������#q40w�JP�<�QM^�Q�jP��X!nx#�F�K�<��왏%��s���_Q�	{2l[�<� J����!ӜŻ�Ѯ:�؉�"O��`"�)�d}�w��$hb���U"Ol��Q��9*�bl҅�G6i�-Qa"O��i  ��m<F���|�AH�"OnP*��.K�}�%lG�T�*8�"O���E�
V/,��_�&|�֏R��yR�´�^�%#�lz%@���y�A.!	7o)�(��ͣ�y���:rI���04�2��'�y"�>
��dM{��=sd4�y@Z� ��`��*tQ�d#��@8�y�d� ��L;�� �X}>�r�D��y�"� [�\d��
ǸSV��Pɇ:�y����HI������?�F!�Y��y�����2rc��1$@�3֤ƪ�y�D�%0�$������.>��Ŋ4�y�Yq�R� ��(2�t��+ �y���o�NL dc;,g�0�c���y��ÝXg�	��>w���Z�n�+�y2O��:��`;�gԷs6R9YDeǧ�y�\w�<��H�xi���c����yb [�|`�yBuJԉ%a�t�bO�3�yBo�{Z��9�Dd)�C��y��#D�T �B��a&���y�kѾM2l��ȇ�hD�y��_��yr��5B����A�K#ST0u�@E��yR≵hQ\((�D�*G�x��c���yȖ)T#L=WߣY̋�O��y2�9u��qya�¤~F���I��y"�C�`��L�f(��K�<�y�k��9�и�A!oN@���y�DL�(4�H?H3��K��[�yr��Sl�� d��6@+z8���[��y�,�6r\�(���U7iXA!@��yR�(2�(�͒;6V@�@�G��y�ܥ`����n�6��ѣ�F��yBiQ�-�����O�Y��(7�D�y2R4(}L�+�)�Uz��ӑO���y�E_�������2M��m��K��yR���h�X!T�U	1D��PV/�:�y���/O����D��-u����m�5�y�Y",Π�g�֧Z��9��DJ��yB�܏	��ك�,�!LU��ܚ�y��t۶A�Eh\ cb��P��y��
ذ���e�X���(S��?�y��J�.Q�e�7�	<@<X`/\��y�A dN�r�-'@�> (5��y���nI�m�GF(=n�uj���yB*�%w��Yq�#��6tph�ܪ�y�b���9�`NmHu���0�y��Y�	if����֟Pqȱ��mt�C�I��^݈�B| �tr�K�|!�C��]�L�b��w�D�u�I?%��C�	�G;���O�`���	)�OTC� S�e�Aܦ]w���pKF�o͐B��+L<FM�q��W:��Iu�D�F�JC�<*���E�OM`�D��d� X�C�I�^UT����*C�d����?�C�	�c"r@����#Ȗ ��۷P��C䉍\:��@H	u((|��!�7��C䉭l�|A�l��.���a�VF��C��-?�����7,z�j��G(��C�I�N�j���� �,��hẗ́�~��C�In�b�)BJ0;��QHA���C�)� $qcb(W����KR̒�<�V�+C"Ol�(8g�xęc�]�P����"O,d��E���X)2C��Q��ś�"OH����7,��s��Ϋ�
�8�"O^)ďӹ`�p�8C�����c"O0T���]z�$�j��Ѣ'D�<�ލ.ujU�V�35�,8e�/D�Ē�-:��p�#�2�|hr�c1D��B��O�|�u	�Y,uef0D�l���%wٺy��#vs>0��--D����N��ži�����u��� �=D�\	�"�-��pB	���=���:D���H� X����#d�)\<Ċ�N=D��y�h��a@H�m�8L�C:D�,!�ƕ<w��͓����@4�1a6D�@��{�(-�#��\���BM2D�Tb��J
,��h�v��-{p���+D�|i@�aŢ�`&'I�@��a��=D�����6WV�(f�F�s�����9D���M���ܛ$��ZT�9��9D��h��,<�F�A���;���S6
=D����	2"� 1�#Hr=��:D�X��	&\�$,;bÞ�F�X3�7D��귣MxTLɓů�2`�a��:D�`X���_��`P���4ۦ !Q/#D� ���#�j�"�!l"Jp:�?D���r/өC�ޔ:t+��_@АǦ D����h�w8L��t$��06l��*D����$%�HJ��A#��ن�&D� �gK�mF�˂����҅�&D�0{҄A�qd���T�����a��#D�``@ T!���a�eK�g�,�@6D��y4�FZ�����E�I#�Mz�5D��#"N�,>DfL�
@/�dٹ�>D��yG%��;���M_	Jl$T�c2D����-.�������)uI�8���0D����-]�mQ�_�(6��{�f.D��۰�ʈ?� ]�"���رt�-D�$�����x0�A%h��٣S�)D��X��J e�Τ��B�J>���(&D�41���	���!��,P��T��$D���W�
�Qb�Pe�΃!
�X��� D�aU�\Bm�hꕀ��C��ś�K?D����K<�T�Ӫx��)C�*O�ʅK�U\Ne#��5��E�"Ov��M"Q����6��v�|D�"Ou+P��->�����Ӵtd�#�"OT������V�d|R�!?X�@C�"O0xq���~�>�aEehd@�""O�%�`���SCH=���W�e8�"O6][3kY� �������"oժ���"O8()�D�`�F�� k�;����"O�IR��x��2�Û�9FT�2'"OP����^���"�M3VmC#"O2 �K�2-O�a�tb�:V����F"O@"/q�d����=�"L�w"OPp�p��c��DS��SM��yr"O��n�:^�y���	�E~f��"Oԑ�G��z5�yT�ց9�\�"O�}r�lv&�:�B!7����"O�I4 ��]�Piك陚��)Yp"OX��U�P�f>����I8��E� "O�1,��{��[�m��|�ҍ3c"O�	AF�m����I�z��|a1"O�  pJ\BpC�A���"U"OJU p�I\d9�ҍ�ۺ�X�"O~�
Y&��fc7Z튵�n�<�֩BH�àD�]�x�"�.m�<�0�&�h u��)l�Z�&�S�<)Q�B�T���Y�
q[2�m�h�<yqdJ:a�Ջ6n� *��`jMa�<��Hб\J�q�5�A�H����_>C䉎����3h	'��25��	ORC��1n~��H�ét���e�[=v�&C�6 a�L9E�8N������(3�C�IB��EE��*u��c����C�I�4��犳Jd�e*�NY�/4�C�IXL��1J )u�|yړ+��@�C�I�'lv���OE(\�
������vC�ɷ\o�x!Єݘ[[ՙ���5�XC�I�obj�`�!ͫV	Ԡr�φ5[.�B�I�Ӓ� �B����F�9���"O�H!F�>�(�,*��Q{"Oi��݇y�*���@�.K��Ɋ�"O����f��f�Z\pTiԡA�(��"O���Q�rQ�$[`ށdxVHJ�"O"Q�7���z�˄-^9EcX�@"O�&Ú;?X
(��-JT:�bE"OX�d��Sb`���	V?b��"O�¦h�t\���B//L��C"O\���oV�,�p@��7(���T"O]ڀ �^=��P=eT"tH�"O^l2�?PƸu*��4Gl=
0"O�����W�#�����͎T"�}�"O& ;�AO�|��x�T��8-w>�B�"Ox�VA�(�Q��]�Rq�	��"O�YS��{1�Y��,��
l�g���OD��@S��[�V���@Ɂ-�
!��?(��[�(�Z�4����PR�'�ў�>q2S��2 �����NP�e?D���E�'u�L����0��"D�`���x���i�� �.����E>D�H*��E�p*��ȃl�ۀ(>D�$a�-Z� V�P�S��F��6�8ړ�0<���	�@�&b�Ib@j��u�\\�<���!-�lQ�g(E���A�ڟ$F{���P:w�r�*��S�x��:�xB�* ���XZ�b4��F�M�@B�']�	kS-9}�~D�t��D�<B�IW���ɛ�m�j�a�g��	��C�'P�^�u���h�P�(A�>��C�	�v&��!A6�$)��잍.@�C�( ���ji*8�Do���X�=�.%������K�v�!1	O�w��@�ȓh��� }̤�Q�n̓xR�}��'��3 O�<~D]��<M���ȓ	����B�XA⍀�kR�B��G�<Y�Tu�p8�,Y'�ʙC�NFyB�)ʧ/G|�I�*L� x�;W��30%�ȓE�VMڒ�Y*��YC��گ�Pi��a��h���Y�'0y��.^IW��oC�'�b�'�ax��SD��}+�)ΰi`ld�M�yR��(��Y��:f��=�S���yF*_�~��'�Te��t���y��J�8�*����X[�𲡄͘�?����'��A􇙏�(�3 �Ի���Y��:D��ɤ-�<b~����9[;��$l�O&��F��'�,ӃK�.&C�������2��E�N>,O���� �8�IR* ܎��u�Rh�K"O�A⬑)*����dԗWMl)T"O�����Μ;� �z'��?���"O*�X5"��^ȭ@
�>.�PH8�"OXM`�ÄO�Թb�j��%�6C�"OZ]��2+��ds�j]��Tl�7�'��'���>Q��F�5 `f�І>1�ٰ��V�	㟸�Ip����K�D�2ԡ���$�.)�b�6D�8�5G�&! �r��Z�A��z�k/D��SD��3�ftQB��F���l.D��ٴ�V�A�^����_G�1�"f�O����OL�O?�RP�FGqV��M�<K>@��\@�<q'JC�)!�J�(2��5s��v�'�a��WL�Q�'�S�p�%�P�yBbA$ �B�[%cCH�ȨZ�#W�y��\�Yn�	W�"Jq�e$�׳�y�� 5�,��N4F2��ٳ��u�ȓ~͎��Ə8H0���|��'aў�|�����8��ݔ|�dx	,Hz�<�ti�(�<e�⇃�Gv2����P�<I�.M�xXd;4t�6���H�<a�G7���37�5c��7�M�<q4JK�e�� ��cH/���0Kb�<pmԙgʕju�ϭ��iڬ�yB��x���ء�$[/�hH�������hOq���Э�r��}8��М=�0���Iq>�9c�V���	�ǩ [[¸A�N0D�4��K�yP,hQ	�PED,0�/D��R�_�9�2���_2��J'�-D���
[*��E�faȍ�P�-D�@95NV�L��`��	JK��[�,D�d{E�)7��4Y&�U&P�~u8` ړ�0<�Sɉ fs�рe螟t�0@��E�<�dN����yW�����M1P��U�<AP��5}����E��]F��*�P�<�	Ʀ_&�*���4���B%!WK�<Y&�
<}�h�F:��Q�DJ]�<�S�9|�Yc�iڬib���SH\]�<y�dA�s�^�����@2�Iq4�d��0=91$�:;T�iX�k��z�0�� �w�<Y�F�:yf��e��2�<:3ll�<�af͐-j貓�
vLr6̈M�<�c�݁jT�Y�BE &p���̎Q�<� �I <�>���/ʾ%�`1�KK�<�cL���4�tb�|<�b�\G�<� ���.��m�D0Ҕ�m�'�a�����P�1��M�$I3��b��S8�y�G>y.����'?��`��!1��=��y�!Y�"dUp�$�=�(��(���yR���1d�#4$��k��D���˛�y2*҅5�p���ӓ[i&��Ŕ�y��M��`y��ƩX���9���y��^:}#���K`��g
V0�y�F�};�@4艉a����#�y2!��6�d�)�c�<�t��-��䓃�'��	^~b�C�K��e�Q̀�t���1�V
�yb6	�&�`��Їv��Y!��ѕ�y��SbW�y6��lyĭ�Dʟ��y2�P�Wج=X7�қV0�JS�
*�y���P1����A�G1����7�y��Z\.��seFB��(x`O˟�y�,Œ<jʹ����x���͟%���?�*0�]�N�O�y4�D(�@H�ȓe��9"��ʞn t�ѣ���(��S�? h+2��,x�@�����#�m@�"O�1�S.�I��!4KA�j�rl��"Oܽ9d	G�I�6�$A�O�RUP�"OUB�	H={��C׃� @?t5q�"O�e���3,�LQueƙS�Țb"ObX�u���j�0�5d��A� �"O����d�*�H������!�"OX���*��d�p�K���k�"O,�`�搒h�D�v.Z6?�.�`6�'����<IQLEEk�D2�-,�z���y�<YG�G�y��i`�F�?宩Q��@�<�PD�F�p�W�N�	���!'g�Q�<qs,ܯ:�b�s�F��m�La�h�r�<A�n�mJܕx�$�?L�x�Xp�<�H�F��q�OG�e���!�Vr�<�"ܐ2��+�-�1+���6�Yjx�$���<	�)��W��=bQ,H�n�:aI��h�<���Êb�)Uf@0JQy6E�c�I���?�}rs��2<���o�*T��xcx��Ex��ЁU��������KQ��>�y2�_�zn���4+ՃwYƵ �,C �y��t�T�b� >�0�Ad��yB�����IL<�r$ M�b���
�'����s�_�p�p�M�[�z���'��	�([�i~�m��i�.�H>y���)_# Eu���~��y���[�NZџ(D��kAx��]��pR��W��y���)
�,;*HUa��7����y2
L)rˌ��&��$��ʥ��y�{��i[����+�=�%^���x��R}���jЅN�1K�1Cg!�t@F�hD-Ć	���#��8�џ��	{�O�y��^
 ���Hע���j�9��$=�Zh�ƈ;���Jc��3µ"O@�Xa+�p�8;(��=����"O��aF�\�&!s���\����"OF�c��E6'h��"�#x��Q "O
�S�!^,_G��h�d��}��"O�����B�ېD!�UQ""O��W�߃���3��M�j�r�*O��ȧ�K��W ��&�@�'>$Q�AD�?Tf�����O��^��
�'�p���7R���/�z�2
�'����l�Q�!��F,La�y��'t:P0���	�ɐ/�WVu��'��C���`9�)�6��R�r���'&���[�uNF��B��@	�'��(Cwn�)��!&��K�#�' �ʢ�12���bu�U�L����'��p�e�3Crt�TI��G����	�'K�pp2��6U� !*�˛)V		�'|���.J�7ILu�C�A��ĘA�'oĕ�B��A@�H�CeB��Z���'WV]9���"4���!$�e$R��'�x�Elٴ�BPєj�>N>���'w>�B�9Ew��$LE�j��3�'e�᷁'<����3	�d��'�p!���>g6,0�A��)o&$a�'��1 S�N�	Pbu�p��"L<�:
�'���p��\8v�P��H�
�؉�I>��L�r��ף2(���}�z��ȓ7Wʠ1��H�`=b�	Ib���Q�L�@É܏;AD����M��H��Hjxաו:��Ѱ�B18Շ�S�? $,I"K=w�:�0%D�I&�lQ`"O~J3MP2�PG��"Oؕ���*e���F���*���%R�(��I=	��0z2ɨ{>�|�&g��zuxB�ɬc��ɱ��ZT�̝����LZFB�ɼ�E�@#�1�ƮL�	�pC�	:`\������ ؤ����	o�B�	�'��F�K�Vw�91d��f�B�I�Ṯ �m�X}����	';=�B��7Z���0<�D�1Ae��0�B�3��p�3>E:�B'��hC^C�	5=:8A��\ޥs��RRC�ɒ�b�Y`��D��"W�ҭM�C�1bʌ(C���H�8���$G98B�� t�f<ڗ郈Y��+�)��#�PB�	|�h1AD5>Du�"��7�B�I��I���:D�1q$��">B䉶wzJ�`��14���#k�
�VC�	�M�$���H�_\�	JR�E4}C�ɬ �|���Í4d��N�+3fJC��70MčXD L�EUDтB�Ι	V.C�I�_�|iH�$�#�!��_jjC�I%I�6�R I<*E#�"A�&0&C�	�}�|��f �	����l�8C�I�$�����̓A�p��	߽��B�ɧ>Sn%X0.Y5ue�˃��iX�B䉨GNh�af!�'"w�@S���>��C�	X�ƙ��(?YCB��אS�C��.��$�B˞�4h����1RB�	C��`�Ă0�xE�HY�w{�B䉹:f:�hу�88=�6�W#�\B�I &�jȱak >�i:�`�=�<B�	�_�,��R3z	�-{#����B�I7Y��!6 �@4�1���=kF�C��#���`@�`�F�BJ��U��C�	24�2iR�Bڇ(aZ�@��M�N5�B�	0iS&š���$�y��I�RY�B䉴X.4I(v�L@�#*
B�	�ݖD�W"޲ah
��� 		NB�@Mv����+aj<H���o��C�	#k��<�Ň�rB4 9���3B%dC��;vYR̠�π��&�²Rp^\C�	�s~z-�q�ڑ3$�ٶ�ҐHC�I�sJ��*c�H�et&�0���0D�,C�Iz����	��K0<XS��,7�$:�S�O�L�0�`E����IӤ͸;>��#�"O�=�t�'MTrH[0��<0,�"O�Y��K���E��AԄ����F"O:�*c�ՏH��Ր2A�6;��8� "O��KUDk��[� ���v���"O��+�!F���o��K�����"Ox5Xw��8Q`y�pA�:n�P{#"O
�0v�''
�i�/N�$,��ZP"O0Q2u�ߖZ�� p�Vn����"O���_�'w��p�Cg����"O8Iy��D���d�ۛ�ĥ�"O��I��ȉ]Y�|�DII4��8x`"O~�B���xT0Kb�Ȯ k����"Oh��EmH�!����"會xL��"O���aF�B�Eъ-:Eqt"Ov��tD�&E���tN�Y3���@"O�b#J�>��C�,ϑz2����"O���i��yk$�HC揌r�И'"OH)H���5S���r��@9�9p"O� T�2��յx;�Y۰��>@2��|��)��8a�]�t]����rO��ZC��$!���b�H�*Z8�Ukv��.C�
�b�C�CJ$0�p�C� A�*;0C�ɗJ&(�oL�n=��;,C�Ʌe��$���n�R��K�s�&C䉈4�B�P�_�}�^�8�,��?dC�ɝm��Pu#��M�(`�e�X=��B�I�A�0�s/�{\�ջ���'�nB�I�^�,��uG^�;��=�V�C�,�8B�I3T�r�(b���e'��y�J@�nM�C�Ʉ*��h`��V��8�n�KU�C�	�|�V9�F�Z��Ц\�h�C�ɲg��TyR41�܄S�a,0���D}��)���u�\q��A%70�C�
8D��!5���\Yְ:!HJ8���6D��;��RE<AӐh]�"�`��*9D� �E�-Č�2�
H&N��j3D���y!
�+�EM�w�(�F?D���g�#,cH��̷x"��9#n>D����ʜ7Ӽ����I34X��UN8�O��P��!�cG��B�0��@Ú�.b�u�ȓb��e�0��l��t��C۸�ȓ?����^	N�r�G˚-V�8��|u�$�F�X7D$+⌈��e��P�Ȩ4$��p�֙�U��3I�6��*�8B���)6�HP���̄ȓL��q���3\���ؘ9dd��'���J�i+S�DC�%��v�x1y�'�H�!�)C�Q����+_�qHt�q�'_z���B�cؚ#�y����'� ��P�3W�p����
pL��A�'�$H`p�
0.��-��ĺk�x�J
�'�q�d�6�p�S#��$6ظ��	�'��!bu�[$@�
CIK%5p��	�'�(B��d@]����*0�4�:�'�r�Rc�,N���,�:'�DA��'=H$Y��*x��t�.,��9��'w���Рq260�#�R`y�1L6D��@�ڂ�����+mf]u/9D�h	Ӯ	6A4�)��
R�昃��7D��s��;s��� ��9�$��H;D�A3�ڈo��r�b*Lnɘa 4D��*���~}Á������2D�L*��u$�RDk� 'x�B�-D�8;�"�DUdT��J� c��2Ei+D��P"�I+��0CH�j�޸�WE(D��XAB^,E��a@����0�e%D�<b�-	/_��5%�2L��ҩ#D��IGK^�k!<y����_y�xx�e#D�p�r
ҚYNt�4K�M���ǅ=D�X�6�C�MP��{���v@Ev�<�ӮC�	]0%pӡ�A���JHu�<i#�߿H:q ����b	+��m�<�a,�s�J$�$.T=y��s��T�<��OQ�y�ͰH�)B���A�B�S�<��Bѡ<�Z���K�JC-�T��K�<) -,a,K���"RLxF)�S�<qPj]��p�HU��*zsrыv�TR�<��@3k�ظ��D$SK|�H�`Pi�<	E�)WJ*�ؒ
���5� �a�<��&?�Us���+�"���M`�<��F�?��p3o]2O���7fZ�<�"J�C�$!�rc�,t�l��g�S�<� ~��Ԫ*ʸ����Pɰ	(��'���'h
%��m�+4�鱆�0Z�fE�	�'�bq�� ,��� ���N�T�s�'�H�90.� 7���U�uSX(O����c'�qs�A͂	��A��)�!�D�h�~�q�mP!y��U#An��!�d�8��)�r��7-��e~!�$� ���5�ޜ�(�����W�IM��L����e)�1��T�O!�����!D���Q*��8��XT#�S)�Q���#D�|HVg����TR��Rzbq��/"D����
$r8�8��$#8���K D�T@5�r�B<c���v2��[E-#D�X0`26y���͐+&�A��>D��"��B-<  ��L�.-�L�ţ:D���3!�/C���?OՒ�3D�h1��"��_"vv�=	ԧ3D� (�O]2r�yP��ہ$t-�,D�$��	C�Y�����(ܩ�N�ɕj>D��[��̇9���+|�X20�:D�8�F��%Wl�"#��a������:D���vɁ���b�1BdpD4D��┋T�. �`bI5݄ �$D����=D'�a!�8UB���%N"D�\���Zu�5X��7d����f�+D� �JӔ)R��ۡ^u ��m+D���gk�;el~Q�w�?f��S��4D�DpqHƢc����C*��b�v,���1D�4b���A�����h 2e��HGe1D�L��m0P֌yI0.��$.�!cÉ"D�������J� b3��y2n�?D��B��чY�P��6 Q�_����0D�����S�lp�a�b�?L�<E2փ2D��C��DN�<h���6$"�B��-D�B���x,h�[�	�`��(8D�V۵��Y�L�	��m�f��/�y�Bp� RN�{�rQ�D���y����;D������3���yB,0���Q0N]LY �o���yB��$V�9S��sp��R��ݧ�y�ŀ�o&H�+%��ii��Q���yR���J8(���#b^6@�b���'8azB�N	BX8'�� ^�
��B�ʸ�yB)�p��Ȳ�A�B.�I��ᅉ�y�
�q�@�B�̚=��# 	<��=��y"�Y�ɴ��K¹2i֨�p����'[az�L�\r��
�l"y"������y��C�=nQz��U�{�0e;�O�'�y�Ꮖmh�A�^!l���������hO(��$ ?P0���&[^-ĥ���s!�م>����,�F"�5�q��=+�!�W--2�2�O�D��)B�l��{b�'��I8iU�	RkK�׀	҇��:'�x��0�\+�)9~b9�DKiAJpa6D��P��,X\.y���sh�M�!�dG� <���d� 0!g1&�O ���Z���X�+ߓ!f 銄��!�L�>�����oel!��C�>!��6�b�ȇDB�m\�����.!�D��2���ñLT3�VP�e#ΙQ�!�d��j��#Pi�$X����6�(�!�J�t<�hHK� tTZ�F�!L!��p����e��6��3��?CRO,���ʕ��	h�$E�H�@C"O� ���A�8������!G�PP2"O&I�7�H6_�f���bí�x��A"O�L�2/-ˈ�w!H�W�ra"OP�)�Ό6�E�/[�@�؀(d"O�Ç�V'L�
� ��F�8EOz�����/g'�y��$[�B3bDu��<y����'��h�x=�"l�2mr�ȓU�ޤ��� �<#�)�E�(u�久� zPY$�.\n��+�(L�N� ���󟐄�������eA�Eٳ��+D�DC�	-�j�A���J^��:%\�Q&C䉄3�-#���?Hf��M4 �D��$�O̍j�A@�v,�DZ���VU�, ��O �=���$S�r�y�ρil�p$ā::!�$C�*4�V#A(yЕ��F!�d�)�f�0k��r���� �;.�!��U�M�JͰ���6�F� �!򤏘zÄ �����=����:�!��ɧ|ngc�ix��Zq ��W����'y��s��@;��p��K*"�Ț�'���|P>c���\���hּ��ȳA�.7�N��ȓK���I�K�� T1��aa��_Jh<YG�I B�BvGn��xs5h��?��'��X�O��VF�Q�I�%4$J�'<r�A�N�=b�>�(1��2�ܔ��'�\h;�X�"��x "ؙ'�֑���?	�'��)�F3P�j��7O��pI�'�|��Ԡ��¦?�*DX�'ޠ�2uꆰ:k�ȳ�Is�I��'b��D��v22�#�JL%v*���'%��;0iH�6���`�U*̾8H�'G����M:��ak6P#4�b�'Y�+R��"eG�m�fS�'�][�'��"����M�p��g�8���'e*��� "Z
婄JV�b��ŉ�'�F�F	�0HC��$�8U��d��'�N��*I44�s閭W�`���'�`<�B�m���*�ϷK�� �	�'����a	-4�z�	��ۡp�PIY
�'f�e���Xr��JU�S)V���'��1QbV����N�:N @)*�'8�8�K�\CqMγ>v�9�'��C�L�+6>}����*�>Xj�'�jTˣ��h:�x���(Ep-��'��
� *a��s$+¬ �y9�'��e�tFٶy�����+͋yL���'lĹ����Խ20$���E1�'���8�N�^6)9���vH �'�tuh�9<���s+H��u�	�';�$��&�$�څD6�y�'4�U�ƩǗN0�U��'ȉ}�R���'����#()P6�A�1ʄ4{vz<��'k��P�(Ŗ��R��6x�|���'=�A��GC�8�JL'h�0�
�'�t�s@5A8�8�uO	�\̈́��	�'��v� �&\ ���L���	�'L���&DҊ`�E���{�|	�'�~,� 珖O~����\�rZ�q�'D�HH�nȃ1�"$X�v>�p�'��Aٷ��.5|�ZF�.tB�'��4j�덢yp�����@��		�'8.ȂnQ$T�ّ��#�L�	�'��zB�9[��%0��6!%��yI>y*OJ��Ջ*{|(��hȄ�d���2A!�� \����A*iZ>��tL�:6ˢ���"O���v`΍Q���1bfғ8���"O m{䠐'LX�-"����[5"O����FM=}����ģY ?��8b#"O�� � ��m8 �#�:W��*�"O8x"K�9\�%���Ň9z� *0�'a��'6"�'�ax��R�zZ0�Q �W�j�Sn� �y2m��P�p0�L����"`��=�yB�J�)�̼ۦЬ	:�O��ybK�~r8m�L̾YĀH�J��y2/W�"Z��B�F�6�)H��
��yJT�P�T8�լ�jx��1GOT��yR��=y��T���U�2��vft%���	w��ԃ�OQ���OC�PP�7D��Wi�,��QG�E���2�'D�`�BK�=M����C zʠ���'D���fCH�f�����*�i�L����9D�0���Քf�b��%��u[J5��!D��	"nėA���CB;p���ac:D� �1�
.`sd�Y� ^�X���O�<��i�8��P��"+�R����đSm�8��AblU��%�D��ҵ���M�ȓV�DV��Bgדk�`|p�q�<�fk���8!�b}w�Yy J�n�<�o�pX�� Đ%�\��$�l�<I�"\��"b7$PD| �h��gh<�c�v' �+g�б�Dl��EC��?I�'؈�Xv�,c#̸�-׶-bJ����'��4�vJA�u"��{1�Ϛit�K�'�h�b��1fZ!�a���_���'8��AD�E�DaE��]���'8�}�f�=p�����`!J��K�'���!���l��b �<߾IO>a����@�
�nY�c� J��!���j���1�X�d!ׇW�$��&��
ώ@!B 4D���4��<#Hə�L��{�Z�y�,4T���aK�-�8�d��lt��"O>���vڝp �)���ٱ"O���t�
�G3VAף:���#"O��`��͉&ˠ|��`]�I�2e���|��)��
*�3���-n>�A"�>�TB�$�\I��LB�W"0���$@��<B� ���d��%
������l�,B�	s2�]
R+{9ԝᔡ��/r4B�I���kc-������&G!5`C�?2�Q��KǺmf�Eq4��[�&C�I@¶ᚢ�NK��`���kB��tE{��'9�r(�����xȆ�g�׳
�!��N8�%3��Z�E��U�g�ѧDy!��/w��q(1lǝ{��U�W�٭l!�dŜ!��A�C�� !�F�G�Lb!�ě�@`QSG�����LՃ�!��T�u��N`:>�A�*̼mQ!��!H棛 3�ak��E�D�ў�&�P��x�Tl�v\0���H�>����e�%�y���:?�t	1��B}�LC�
��y���Jg��1��n�,,��-��yr�Ԟo�&!�ք�����2EG���yH�|��ARfM��z�z�C_4�y���2L��k�gگ|-�-cD�ָ��xr��0��G5l�\)�WHĈ"ўl��
Y�2��OI;����e�M�z"B��jD �hքU����6YB�?_�4HL7O�� ��nT��8B�)� R�a���@Eځ�#��t+��;B"O��"�d��J��������  "O�+�(Ft!��7+��
�"O�E�E���;
h;�%ӎ)$��[r"O��2҇�/�h�$��m|>�"Of5�C���?4:�����7�f�3!"O̡���@ir8ac]0h[�<p�"O�|ˤA�<GUtݐD�D����"O��ӷ�}L����a�$y�d"O^�0��	�tHp��栖	7� ��T"O�L����r
l$`Ҝ�-���'���u�v�S'�4�.4w%@�S�C�IRU�E�%b��~'�Ҥ��NB�Ɏt�r�z�m�3r��1	P�\�Im6B�	i� ��VDP������=,�bB��F�&k�b��b$���T�� _�jC��%P��%�޶�yI��}(B�I:	����ЌAz,HP7� 1Q��C䉵U�ܵ�����kB`jW
�2b`�C�@K�A�%�	�u,P�a�K.l�C�I(Ss2�Ѕi�!��)�l��3E�C�I ����ΰ"�p�J�B��C�	6P�U�5`��.����/&C�ɐ-ЉV�D˴�HbR�]?$C�ɦMÌ��C"r����S%��C��o�~I�%�P�@ɒ��HB�I	q\%�tNF�tܒ��t
��\eB�	!F�ސӆM,�r�x�dڽ>�C�	���S ��h�BH��Y���C�	�\��1�����Tkw��>��C�I�T���ՏA�z���1@�Mj�B�	9K�.a���	��A:v��8�B䉆�̜����	9��!��됊��B䉡_έ�R��G��Y2ƭ��&�B�	&�lt��MD�:V�n�@C�	
c	�%I�L�4Uf��7�[�D�>C�I�rĶA"҂F6=�6�X�	��C�IFI:��k�MS)°ȕ�@'\B�ɉZ�QQ���.�8ɚG� _E8B�ɭ=�0�
Pk�?(�\a�0��ZB�	�56���S�*B-+�!��=�&B�ɻ@�`�q#ۥp*=!���&-�B��7�l5�G^�i#��	�`B�ɝ �V�eΡ2N��u���C��e�$�РlR&F:����&M�B䉑c,0\���bcy��D�g��C�	�}
�$�䮐�K�L�!Û �C�	� C�`C�!2s�LR���o��B�	�*�`���"R?qچ�&�T�W�lB�	�rӊԳ�c�+7�0A�KS�t�B�	&� �Vgv�eF-�JffB�I�J*͐D�2h"�!$�9prB�ɘc�xlq��z��,��G��T
�B��")� �!N7�(�a ��BLB�ɳUQ�i)���%q��X�ș�X�jC�ɦ�����[�4XH!��VbhC��g�Y��S�*��g��
ŠB�%
c�к5AԱoP%�G*֔I�vB��&2����8N
���<m�B�A��)�JƘT'�𓁦W4C�IO��\ʦf_�~�x��G��4__C�IY�tj��ԞJy���r�ü@oBC�I.?���`��-##�L��*JqXC�I&@��X�խG??�h4q�h�rC�)� h�F�W("��Y	Q��UІ	"O���Ĭ�odf�S�F'9
q"O��;�!��o�	X�Jp*��R�"O^��diK0]h�%ˡ�E�a�"O�}2� ��i)Nl��� s3d��"ON�z3�p$�`�#G�O���{t"O��!�%Xn��DR0$d�`3"O�yK�c�z���F�_+4Td(�
�'��i�ԎU: KA�(K���'w��H�^?er�9�D�Un��'*� �A�uR	�ƙ�U�
�!
�'��y����&
L�1ǈ,N��	�'|�J��x"f��nבL�x���'�ܴ22̯ ��mi񠍫�HlR
�'f�
�b�'2Ϥ�Z�j�6T��@�'d�|�T�'~l�R�,�?���'ļ�u�֊�x�J`řw���'���BS�B��OD�W�����"O���&�ô_���j��J����P"O4 ��l�30P���lY4P��5"Od��̀�t�]�/=���w"O-1g쒣
NDY1��Ф-؍��"OxI���S@N ��#�k#@	�"Ofu c�,}���"�T"9 H<k"O x�̶v�YzK��Wv�	['"O��{�X�/0$!��C�/����4"O>�[u�P1s��`��DDiX�"O��2t^�6V�+S��c0�p8�"O�����	q���9�JK4��ɘ�"O�("6'��V�\|�'͛
�$�I�"Od���[�R�D�	�Y�"�^q��"O��(S恭���	�_�����"OK#��f��%'� �j8J�"O�La�ۼBxza��/Nx��C3"Ol]�$W1CCx�Ar�!�"O����a�����T�[�J�;�"O��@a�`Q�,�%�T�F��"Oh\�t���5J\�"RI�>|��r�"O>L �EP5>��3Sj�g\\���"O�Y�m�8?ZH@
Q�J��[�"Oţ`9!&��	l��=K�"O�p	�L���6`)NѴ$o�9d"O��%kΝ3��D[�Ζ�S�� W"Olti�D�9&2B)�SM���hi��"O|t��J��a��,�䌓6r�"U�P"Or�@�e��(rD�QL�*+�n1[�"O��Ab��Z�B0��K_�j��h�"O�8���T Z%zdꌝ`�.��"O��P�Ds��U�r���H�<A�0"O��7"�!lBP���C<Y"O4���ç{m����\�X�ȅ3�"Oq�O��~���M�l��p"O�M� ��=OH1���Q��"Oniȱ!�mf�I�f�J�ᙣ"O�� �h�.,D��� ��4��"O�5"b����q��_�ڔ��"O��)W�āT���R欑�5�&�I#"O^S6���+�{$��o#!7"O6���L�20F97���5"O]���I�iu��	Q*�ޥ	�"OАk3��=��z�)�o2(� �"O�xp ��/KoDH���f2�lRQ"O.��fk�w�||s�j��R&�-p"O�*�,��Q# ]�F���ss�*�"O� �E��Z/Rw�M%�Q�7�8�q"O�������p�v`1_��<6"O���䄋#�����Z![~�|�	�'dd܊��^�Mpy����	!1�h
�'	|��꜇qw���X��t5h
�'�8crMV#q��x"�+y� �9
�'�@��C퀯s<�m��~���'4�!8 JR.�YB"��,�*��'��"���Nh�x"ã�&�xX��'�d}Y�	�;d/t-)B+W�XȦ�h�'nzݛ3F��"�L�k�!��@��A!�'n�؄l��>�H9	Dd΍a0�`�'����$�*&��acR�V���
�'�,$������YPSH��W�q��'h���犌6�ʅӂ� W���'B�e��f�,I��1$U�P��Y�'m BFқ#�4 2�?oJ!��'P�%3�3�|�*q�	l����'`�t�-La2ڀ_�g`0�:�'���A���1�0@��ˍO�6���'��:VHS�a�`����/E�0���'S&���N���Շ��I<zlz�'˼��gQ7s3�0ave\�EEb���'D�p�ͽ.�<
&ͅD�䵺�'��0s�
+M����ŀ��9N��i�'Ţ@`�ER<Vp�b��Q*��E��'t�Y"v ��4�"�1�J������'��!�di؝'�|0U.�B�	�'ô��%	ӑh<Xt	�jN��p��	�'��ܢ�S-R�>��B\�m�d<�ȓv��p�Ti�;�(s�'	=o|��K̽X�^&�pt�O�*��y��{�&|�$dT�4W ��&�o9� ���Re��Is���fDW�,��q�ȓ&F0�B��/��}+�"I�/ܢ��ȓ��8a1�?'?dlS�J@4H#��ȓ
<�h�5�L2U'�\�Y9�NIٖ"O���Uc�|�/_5Hy"Oh��Cg�5f����OnS�䈄"O�U6�Q�4����n�FMR��3"Ot,�C�U�RJ���9?+��@"O��'PsB�zc��a*�h�"O�R獇�'��`1@QXXűv"O:�`6�U#7�8	kf�5�t(�"O ����f��|�tM�A(J��"O6��`�~�ʃ�(ԭF"O�#4�S�ļz���?B����"O>��6�G�̠��܏,j� "O���%��;D����"2%�,pӰ"O�
��I�����Ӑ)���"O��AlA��f�B���>��x�"OL	Lf�P��o�8yݸ���"O�Y���)~.�P�3��1"��{t"O�H��ic��C���%um��hҎg�<a�%�c0%裇��w��Ux��Qi�<a&�, ��Q�܄3o��A��P�<�f��wF �1փ��L�6,��N�<!.&�}��D"z+�t!ѯ c�<��J˄[}6���O!|�`�C�<A�JD2w2���aAE�l�0�ǆj�<�T ��m���0�(�>S�� 4m
a�<��fXJ`�ӬU9v���k&	\�<����i����v���1���Ir��[�<y�X,1!҅��l0$��@�Y�<� .!�!G4 M�ɀE�J�\���"Of��#�2&(�L��F�M��YQ"O>`���2g� �:��+/��[�"OL���)���q�e�r�p�"O�5b"ܯyI�J��z&��U"OT}�pBN�w��-�d��M&���"O�!��^�����Ri�0 d%�r"O����,QUn�i#Ѝ�Ɲ�"Or�x�l���d)Z�M��X��h[V"O���"�%�j@�6�"z��E�7"O�d�4M.e�l��m�v�Q�q"O<i^m���A�t�[��H�<)��U0&d�w$�&?H��Ъ�I�<ywW�cÜ��Ab�������F�<����@�i�8	��2��D�<	��H�r���f_�L\�M��
[}�<��K��9�m0f0�	���y�<��ׁ-��aaG�(S�c�NFt�<Y��="��Y��̞#<��"�f�<�AAU��fK�m�jT�s�@_�<��-�'+G`�2��)�dBcbZS�<���s#pp �
M=n$|`��`U{�<�W莮OPtxW%ƱJ����3ƋA�<��V�s.�1Ë�)���b��\I�<�ëE�2�Y��ĤM.4�ڴ�n�<1v�W�j�+��l����Mg����'�����*A:@��H�DA��<�TK8$���G_�n&�AX�ő0�Ҽ�E�0D�d����>�D�� �D��3`C2D�xc��Z�[lŀfA��#�q�0�4�I\���!����A`�6bȲ��6�B�ل�5���@� X	 hP�_���)֠���C[�%�A/xG>܆��f�r7�>^��E�f암-�H��jdH<1�M �{p=r���s�R��@�O�<����Һ({�d�#pSl�X�B�T�<�g/�2z����!Iֈ&+��X#(BF�<eo	�6BrH�UKO��*e�ci[E����?IF�T��l� �_�l�������8�Z�yg��&_�)bC� �4�<��?�^["���<_��"4-��zG�B�=�VP�cG�/�� �6f��B�ɚ'�.m�Um�*jی�b�&T]�����%�	�E��dQe��lRA�1KТ=�
�<l�� g�Z67��u�EB�iyX�<Q���I�p��4����&mH}���4|!���7V�j<�c��	oc����,Gp!��Wx�h�CO�'f�$a� �M<!�ƶ��IA ��.X��4�s� �&џPG�T�+�J1s��իQ��a	��y���� D�rs�L
F����-�y�%�C+|��gV4S|�������hOq�<��1����Q���KHPuؗg�z�IK���q�Ò
a,�Z�֢P�x� �(�hO��'�0��q�p	(F�ܔ|ܲC�ɏ:�
iJt߱`ȂH����o�~D��'z��8!E2H�j�@�h�9n�M�'�J��A.��b�Dg��T�΍�yB�'[,�`���* ��4�V�I:�]��'Evܘ��AzHK1dGH�J��U�*$����.
����A@>PԍP�?D�Ԩ���a��+�o��*
�=��:D���o�J(h0��!N7xĞ��=D�Xȡ�K�f�c� �/g2�9ہ�9D�� ����%��]�S��B���b"O�j�L��R��W�\^\��ON�"�ϐ�J&�QFH��4���K�4D�t��'���*Pz�%W\��3D��k&�(k{0�Z��4 �0phu�%D����h]��B;*'#��ڴ��<��Fh�x��f��
P�S�B=��p��{���se�)-�����ȼGq`��ȓMV0��R���1k��"`g�mZ�`��C+*X��n� sV�Jd��
a6��X�'�ў�}�a^ f;ʩ:����-���P�i� �'N1O?�d���~ j�i�)--n�xS��o�$|8���q��1�6Ĳ���(�D����?���' ���O�}{�f�I��]��O�?[�l<P��V�<���&��آ�Hj6�c��C�f,G{��x��i�&\x�D�X 
�H���n�#Y!�d��,�j;2o\�U����LH��iz���?�~���e�ā��Z��"�	E��y��)�)�ty�]��Di��
=����@���yR�D�`�sj��a�ly;�ET?�'��#=�|"W-:j�Y�(^.v�P��,^r�<1E�>Z7��cr��-.��(�|˓��	��ϸ'��A�J�_�����Q�+����
�'_���+ӥTR�*��SN$��4����Ov�b?w�ϡ��I�E�*�(C��)O�=9Ѣ��]~�&De�������t̓K�a{b�͍T.M���3"��R#'���d$�S��yrm'W:´[u�	�Y���� �y��Zl�����j������
=�䓭0>�K6��$j0	�;{�t��l�y���Γ,���ç@p��X�1���s�l15gÅL����R�x(8�#������`:��_&jp�)V蝁9#�I"OvQP!�1]�F8�dƑ�7f�B�_��G{��	F�S�@��sa��D��D�ċ�S�!��V=/Xy�5`U���H�3�?~؛��>1H��'��'�PP���h�����d�� *�'��
� k�(��0,V�8�3檜���d0�OJ.0bu���ڟ<Xp�a쇞B8!��
p@����][�tӳ덧I/�IL���&�ӒD���-
XdP��<)�O0�$?��|�IQ��X�S�b�n��ԋ�'RY<)��YZʅ`�����F�8qM��b��ȓd@ ��b�G����U��	 Jb����[�'�a�z/$��wk��(� �'w�q���Q�wlz��@�P�s�����'E����/�XU>�����t��T���
�y*\	L��9aK�- _����C@���$(�OXdA�ȓ?����cN@�I%d�*D"O*��F��+$����n����t9��Mr�S�O��1�f�*�l�-t80�.S��y"l�p�`���(N0'��b���yª9r�8��'&F� �qq댾�O�=�;�~�ڄp�6/�$.tG
��y��ӨrG��!u�W���F>_:nM�'�a~rIV�D��I�'֠i�����y2,��Bb��6iw��
5�I�yB*�uyZ|�b͕�V���"W@���yB��;T�8A���# �ԩ�F��y��V#m�̋��\'@Op2t+�R�ў"~Γ)�T� �!��a��l��ȓsm%��b�P�N`Iq��fϐ���?ш�&�j�B�K�960Qp��g�<�%m)m7�$�s�2i�2}���He�<� ���sK*k7�#d������[�	q���非.o$�qe�׎tR�[6�"�!�T�c-"e��Y�K!3��P#�!�dBP�ީ�p=7��X�� ,�!�Ni����a�U��\��}�G{ʟ:��!,R:��h�	ɢ-�0IA"O�� �)D8.c�JGԎ�>m+�oEh�'Tџ��%#T)�0��Ɓ�xID�R��(�	y���)�<��j��Ӑ`0�/w�����L�<�#�� ����-wKJH�e�<	����HK�(s����֊XU�#  �B�I*R��	B"�a2T�A�����hOQ>-"��I/�D��7e^�=��$�g&D���j�~<�8�HP���!�E?��>�O| `3��0k���ǌ�<�R��\�xF{���B�.蓴gE'3Z���#�!��O��h�T"�38Q��E�c��'�O�<��]0Q,�8�P��J�Ąq%m�w����(����rD�	ǎe��H/a֘��ȓvmґ�޷aW���g���������j�'Yl�� �J�&���T@p�'`Ȩ�A��&�x)v/�,t��� 
�'�Pa����
��g�k{�g�<Yq��1�d��1��!��kNN�<�cc�vޚ�xf�֩u!`�q��p�<y��,F$�]
=���ђ��l�<��Ɓ5 e2)�t'� G��HѬ�f�<��N�~I����Hp�ؐ �_�<Q�Ꝃe�!��	=yf�(�(f�<A��>D^X���J�s@C^�<Ԃ�R��XC�oO�V$8Kw�B�<A�C	a�5��KT�M�,��z�<)`/͙8����ۿ �ڈ·JJ�<!*أ�,���H̸���D��H�<�siޥ/��W�?$&m-ԒTJB"Or�,%�����n��K���{�-^)�y�cu�^<��mV�U�� ��y"ŉ�L�1w�
3<��-� ^��y�b��h~��[�-��
��y��+P10t+��*#Sh�/� ��'����6mR�}@�5�!�^K,�ha�'w���p�]>��0�aAM)I���a�'��!q��!Z����o�:]DQ��'�I`1J� Xz�I�	�7tP(��',��)7�l���۰��)I,�k�'�x�`KA�B��eXЁ܇*u\��'�td���:֐�"�SN$�l2�'�M�G*ߑ<bF�BB��G� ]�'��H��F^:���B�#�kR2݂�'���q�쁱X�՘@͘_2�x�'*pE��+�� ��y2�L��[a^٣�'Rn�収�h��p��!:��'��#1e�y��H���bԈ�'Y4�IC�r�z��7�\
*�^@�
�'��)`F�O+t�R8ig��P 0\��'�re+�ܐm2�[pWw�h��'�n�HrkO:Y��g`@6&^�i��'�\X��	E�u�>��V�O��@�'TzkS�����U&Q D�Uq
�'�v�#��nF��ӄ4p���$y���0�+>��]�@�A�$ؖ<h�HI!�V!T���`� � 0!�D�8i\t�𦖨<���M*�!�D:_��zr'զ#��)��^,Sw!�$�N�d���DGz��c��&`!�� b0�t��/�B�����9c�4Ke"Oz8¤�KL�3��Yd�!E"O�Mq�eV]�*�P���$5�Tp�"OR��&)��M^�����=J4fMʲ"O� 5�ɸy����@w,Ur�"O�#%�݂j��+��-f�b�"O��'���E�D¸9�"OPWHAȎ�������컂"O�hH�]%r4p�&$K�pػG"O\���![	f��|��dU�8��1�"O�Q��I�
&�E E(��)�(J�"Ob ��L
4]d�<�"��Z2�"O�Ek�HY�S=ReCAF(zOtkC"O �#⭁�^!t�"�LYfO���1"Of��b�&f�ݢ�l�x8���"O"Dk0��d��0����n��Q"O�Ah5��x�P�,ǀT��"O�P�fIՄ|v�1$D�"ns3�"O���P��+c�c�$�4M�Z�bb"OX��"^�l�q��Ms\�#p"O=�Q-X�(n���=oS�!�V"OX�k@�ʖr�v��S#IW��"O�w��OW�ai�l��1B����'Z\5C��x���:�L\���[�Y�\��&U{�< �R�9
����������v̓����B�<��^:����%(uaѧ x6�RA��?�Y�"O���Fmʅ@�E���t���$
���$-Hl�P�/��r��'`�i������$��Sp�y�	�'���P6!D�8h�ԁP�'!TX4)��bL���8%1�"�!K�~�>!�A5X����;t��cʄFx��a�N>s���9���3҆�c� p�e��q����$]:&g�pf�'Ԉ�" H�;�q���%1ԒN<����Ie�1!�' ��kqC�BX��d@�j�f�6�ˑ�9YV�U�r"OΕ�-��1��HX�!F,y鐀��i}r��=|�#_����~��N�:�~��YP������a36��̐x�IC�_Z$ȳ��'Fƥy4"Ԓ01e�5��}y�F�UG��@�	VT�'Yp=CɎߜdڦ�A�O1��˓���-�<��+�E�\`�ي5�b���ȿ"�����uO���$h�*Xs�HՒ����wOQ���'pe!'ObyB��D��8ص%}�iš �T����}��	c,�=w�!�D	�
-ơc��I���,�9��2�:��a�q��?=S�R�x�T�������Œ RS�8���;D�xRg�6�b�y�JNZ1j�bk@�7H����x�B߿L���9����Ac+N��y"��%E%c?xZ&�����
�y����mI��D��	|�Z��s.���y⣎�Y��J�Y�i-^���jA��y2@E2��a��U�bƒq��Bڵ�y(/`��`He�ʎ\�j�H��=�y҅��AK�*6�ݷL��h��yB':ϼ��]�A���"��^��A���2��>,Oʩ�\�x'���ŉ� ��%�'�@�{e�(W��աՊp�8�(�J'k N�b5
O��r�[�k
�@���J�]�dE�a��,VE�	�֠L%n1�01�s�$�b4��?��!�"O:���ϖq��܀t�����|���O��D���~�8�M��}z�hG�,/pH��G��*��6B�#G�t��=��1�gyBŉ"F��s�B_)nc��˵HR+��	>P�Ҡ�W+P%T�џ42um� �20ui�7I=�H��:R�P��KSR��y"�;W�N5�3��1/V�u+�1G��p�Ě�<��G}r���Q�Sdn��&M���X�3�S T�lBWm�
]��F}2�?</&5��Jf̧O��Y[�� �JJUJ��x1���'��
ԍ_�hC�i;j*�>A���-�M�5D�g�,q�.��`a�h[�$�4 [E�>E�D�'/0`Ѣ�*ot�{5��9s�h��b�, ׽U������y
� � ��U� �8�i�ˮ]-��Q7�>A�f�^�T|�N,ړ1���%��R\����Fp u�q��05X��0 /ė-��q$'0O���2lƀj�f]'��|�-��+�95̊M6�*�l%��o�� �f!�Sg�[Ҧ��~j���#"��9�@�<It�?�S�ߺ��b?q1sE�8t�a��;8�8 2��>��#L�<����V!ɒ%���r)���)�5B��Oy���⦇�$�Y���7|���'x����a��6ఙ��H�j��怇^t�)�8i�B��v!N�t`T�����7���%�I/
���"W�@v�A��I	�?�7�	_��a&)N3�M�@ Ŗ����e��>)K^I�欌!$ L0��*�	YZR����o��R"�D#+������I�2[d� �,Ja	3*w�&˓r� $eͪy���Ĩ���\z����CW޼a�\?K��x�LA6_:�-��,O�?l�Qґԫ�t���ޓ}��}�K�!=�L�ӯ�1�b�����*$8򃍄9���H���;
�Hp�aK�#;�P���3�b�����yGMP�P�R%S��xIP���M�����[�B{Z���i_'|�l��ƫ^�!|<�����^��y�WΆi���"���N��U)�%y�`����^=#z,ȩ*��MS����g�` y��9"��p��l�'��e��dH�V�Њ�!�8�l@��#L�� ��
�`�����=&�����E}�d��K/m��3�@�/T�E{2C7H�l#��1CC�H�T��ly���%��S/�^���m� ݆X�,ѓ<Z*͈Rį����d�vJ��j� l��"�ݮ?@ ��x8���F�
�<q@n�&n�f��Rb�:;�)X����Bu�fo�>/&>��c���`��p�:Y������i�MA"LD��$Y� ��7�]=L+�eD���,"=�4�R�BF�?I�e��7�&`"�K��U�D�FG�E�p��&ξA��OL�� tD�7�2HA�,�uG)/>=!��c���$G�+�z<җ���j�<x��i�� ��E�O��?���"~�4����æ�	�)$��\��a��>��Y�jʗl��-Q����+��#��&��d����&��@���0~�Ҡv�Ͽ	q�)��DZ�:��I1 u�a��%&����6O�`g�9�PRbml���t�;�8p� E`�iꡨ�5a�j��-6@�x�I O݊A�Ɉe)� ��"<��p�S�	�P���H��<��i��&;F�V��' �8�(���M;�(Y��N�_�Z4㆖�BW����^7�����U�L�[/�>�؃�8/������J Zt�J��T?|ġ�bI̞ɪ扨5B#|�'���ƃG����HT?:K��3�n?p�Y����[������-F���(����3��]0P��o���$��	Qj���ϵְ�92��?�fU1g��Cd�y>�r}q���Dh�@�@-Ƅ[؈�Ӯ�⠩�Q_!��CCR2	jFE�m��!D�4<;�'��=C���79<(4Q�eR!db>9hV�6w:V���Q�[b��xwl"D� �`+9, �;!n"}D��y��ׁ������P����DT�f�?�'��58�̇3���y�$�Lh}
�'Ť5X��P?J��a�P8{u�찳 ���$1��G�'��3��'p�t��q$�!x���q�x���d�"|����:c�a��A����0PK��ot���'�LT�s"D��x��	׈`␀@O>���W	c垘h7��:%@"}�tZ�X���[�o��h����*�w�<y��߄���@=K]�}��\	%uBY��'Pأ��Y7.Ɓ���Or1�E띱_���sW�ͭraD����'���A�+٬XAf��W�]�T?�=	�	X�,��U$�}'�}@��������gO
����%Q*D{R D�x:�1ZR+��C�1�}b�As�b����/��8E"O��!�o�$�r%1ÇKk�0���'��p �m�6v�|�VX�"~�׏ǣu�\[�O�`�m۳h̜�yD�9�T�V	O/ ��RG��$л[/$�`�ʟ2Qx��d��C'V ����?]���c"� 3��'���C�	
�<�a	�
0��{��Y�hh��/ �t����q�xX�4��ƴr�BѢ�e��(<x"��`���0E�|a��CL4�|2�ְ<8]�uk�2�z�����t�'��ͩ`	n��3+��Z3҉:~΄��-� gmN!�ɪ750��C�͊Jي����RA�4��y��jA�N�$Z�Z�¸>��했?p��"}R���2��pp�n�-B�]� �Uyҁ��b{���Ñ#Uax�J&�D�c�֨<D�+dC����P~��K'�&�H�P�Q�ӏr�D�w��,[&ș�C_��	�l4�O�1ǌTx����D 0e������a:fܐ��$�6� !�,�S,u0�I��@�;5n�$IQ88a �?q���!Bv� #V\(k%/M��԰"O�QC�f�Mh<u nI6L^<!�"OfdA�ߏJޤHQ�L:K|�r"OZ0��I�P� �ץ��R�9e"O� @ �`�ZJ~8xS�	lD�	O.�I��R��;�$�$"4���6,tC�	!�8�j��@0[2�	�L7F�\���]��b�@�O�m�":��9�"�(h�h2s��2]u���k@I+��'6Z��$O�a���0Wo�qr�\�K�,���_�*��	�{u��V��A3���?1�K��O(
5�d�$��I'I-D�H�E�X:�<��g�,X~p%be�<�T�Oh�EH�6~	�.�|n�,C�b��'b�@�Z�o�<ٔ�����r�:���M'z�i�N�t�5�b�Q�&����E A�P�t_��T��H�Q?YP�����D��+�fT	`��Xh�O�*
�,�S�S�+"�a �<IРn�	a�`�<xx�A�G�Ɩ+�أT��Oٻ'��{�dxY�d:Y� ��=O��� ӡ����l�Ʌd6��DZ0n�
���0~9���f8kL�"5*�����9ZM���g�B�Y�!�K_)�Q@4�.P��4��yw�I�xz��&gYv��C%-�,6M�o?qgP>)�qiͩ
"8tKe��s~|	Sp�.�O��"&�� 9"�i�н)�l�(��
`�����C�u��ˢ�W� r�O�>�	�n�:����̈r�԰��/�=
�"=A�g�5}���{&$��n-����aҬV�AF��s�d:x(Ѳ �
��=��nҵa��H(��V9�"$��jB��E�F���i��B�>%>͡W��-U�I�	++
�KR��7!6�ZA�=��C�ɳ�vqkPCAI�P�2%^�0��/� *�*�V��0�ُM�qO�S
���#��r�H�#@�<�B���5z�J�A�?+85�5f�7�jQѢ��2R�	�
�'��P�`�@70�;� ֋d$\<����	�A@�#�n���O�b
g#�/e�8ariM]���[�'�P]s���Y 4{`ΏG�܀�ߴj�4 �K��e+ҧ����o�4jMz��s��7f���i9�y��^��`��	&/�f˗����O~>e�� ����<����ZVd�,������6S 8���D6Q2�k����x O�-e��EpA�W$��B䉍e�*��vF� u��av�
7��">��l��̢|"�MҰx�8�w��%%`��A��Q�<!`�&�%9���WG�%e�t�<	�D�|�$�z��:;��D9C�Nd�<��k�x���k�ҷ�2�lDf�<�C"�+p���x�f����B��FZ�<a��W�2y����K��plr5��^�<y�k��j�T`k$fO Q+�y�"�_�<酬��It8ZE�X#=.%�G�X�<��U�?D�)�"�9�($�J�T�<1��!WA(�	��W��ȑ$�R�<Y��ğ���v�P���iB�w�<������ЀĽf�*aAf�<	@m��o���q���4Cse遥�a�<�f,�\�����0}i�ذ��c�<qB��*������*of�H���p�<!�&��<K!���2�x�KG[i�<��%$ ���_�2�����O�<���!|�p��L�5o9T�Е�\K�<�  ؇!��3�l�+#[0pX��_z�<)B��`D�Q��e�g����k�I�<)�@ٔ#z��A�A�TLӣ!�E�<��$�+���wO��n�^�we�<a��صP$h�� �3E�6�(eB�\�<q��OZ�"�`'C2�@��SJNX�<��#��, �F?� �q��Q�<��/Q�D�x���A!��@�B�S�<)Wi������3��yI�iSa�<�B	hl����$W�8l�k\X�<a�$״/l���`�\+'�d�w�	U�<��y��ZU��?K�c�"V�<WP1���8��5��M�捁i�<yF&1��[�׿}o��� ��B�<P�J%Ő��s�	�3� h �Z�<� �PJ�:�� �C�>*�Nh�"O�Q�2,��S4T�6e��Z��*Oz�`�0W�&yyA�� $��'/�hrBhƕ!��u��k�#QB�2�'��Ÿ��U.c��l��өb5+
�'Ȧix��c�b���(��\���!
�'��8%��Z4��-�\x��ʓN�P1�WfMȡ�0X��zE��9W�:���&3�#�L�����qH8�c!ݖ��a(��Ts��ȓ��t[���08�.��r+^1*4�ȓo-��bǪ�	�:EAA��j���i�Uqn�/��Ig���p�ȓv�l��gM�$X=�$d%����ȓ`��]C"J	5NF���	�*l�E�ȓ%�f���_e(���,4̤��i�Jq�q#Ւ/Ю��E�G�%�~�ȓ	�W K�v~&Ukg'�V� �������#H��~�᧎���͇ȓL�9P�ȥ����щ�����ȓ{���a�ٔS�A����������Ւ�@W�pF�"W'݆��<�ȓ[0���T�P�V�Q��+p�����8���L
aɰ%㒦*,��ȓ16^�;�B�>XJ��j�*%r�� ��:�0�Շ
z�|3�˛6X��q4 Ү�,6`��)W��czRQ��"XnH�������BN�)HXa�ȓ�B���R4f
�������I�i�8�Q�|�e�
���	��Γ`h��'B��y��WӘ4�g#Ҕf]�"gό/��	�(ɰ0Z��Y�)�,..u��E�9�LY�Qa�t��B�I	yJ A�@���+�W,4�q�'xK�!�b(�v�Q�g�Zy�a;�O�y�ޝ[�獤#6¤��[}�A��ޢ:�|H��	G[z�K@LI}[��S�'�O�E��+ 9B�{�!�.|Z@�E�'�
E��
�0
�~ѤO��!7�S	Wz�8pe�	C
�q%"O����]�u��P�GO�ZK��"������g�!���e�>E�4&����Pg�۴:=Xs�J��yҋ01f�Kd�E(T���g�(b�2�O�d�#νW�1�1O�t��Oƃi (""d@)8`5O�d�L�d�6�&?�m��ҵY�$X�tA��p?I�甭2HVQ ����n��=��U`��Q�J©&�0`�5�>9a�H�2d|z��4Z�<h�f@�<ٖnָ�|8�4Ɠ�>�jd06�BA�D'5x|��@L$����Q�����I� )�}�&B^
^�!��*;�mZ��ّC.�9�6!�%=��H�0������8]�ı�xa�p��Q�`�ȓG�\�,��[0��CŌ�(6J ��\�㇍Жw&�8�1(
}~��ȓH<�A��T2=(�5���4O�L�ȓ#$T!k`A�1*B��&@�����D+dt�G�S�9���Е(�� ���%��]Kr	M7u�2�k�흮
�P�ȓj�>���Ǒ9gC�Y{���#;=%'�\k��\#:<ay��b �6�S9��(�S�Vٰ?��
D���.E�J��A�i_�x}�tc'���Px2��6^ծ9j���5�f�ʥM(��O�d�5Z"iFU�����%\���w*��^Q�f���yb H�����CP�
J��v��~MM4��|¦w���E
*���ݳH9��'���X\B�I�Z�n����f�Q[�]1�'?���v��g!44��	�DTɪP��-L���vX?�����xf
mY�C� �f��D�c���
eA�E3J<� ��8V$	�16��=yPC��	aB��[�#ҁz�1����ڍ9���yei��- �Qf"O�!���J� ��'��	�`x��O2@z�a-8�ȕXH��}J�%�r���2R�~8���t* Q�<���>��K0p	@c	�M��"f�*�f���0<���ϗT���*��U�D���,WO؟���Y-��,Q!O
$0Ĩ��-gOڹy�i�R(<��d�<�>�:�$U$�4�U�}�'5���4� S���3B @RR���8���=�#D�]���D�~o�t!M"ZVz 	Y��xr�D|�n]��E�	H�¤�/�8p]�АNִ>X�"dRkʩ�DϏ������:��OJ���Ӽ<�0#$:J�G����$�n��oD�Zp������4,�j�/ļXt�D|b�ձn3`���x�Z.���$G;�=膨9��]�Oݨ@�d�Ԫ'm�0lIP�a����k�*�Y�V�"�D՝ʉс�'��}i�Je.R$�g��F�L��_4���	�Tn�p狷r���at�J3,٣a�F!q�l�;P�B��˒�1�FŒ��.1����R�4����xG���`�<�bM���G��D 9| ���#+��@l��@�}M���П�Hx�����M��擃 p�S$jƲg#�A�P�'h��ϐ�ǆ��&��p}�3�ͨ2C]Ij`��A���mV8{�kP)6�A��ǝ>T�F�1�#=I,_;p������%T�fa)��vy"��!:�D%�EEa���'T��t�Y�/ �4�6���pp��棊�aV����% ��Z���#m1��#6�/�OB�ʂ�^�J�"`)E��>L���U�)����C*<l����x�Vq��Y�F��J4��$R���w�\`yө;�4�a�K�n݉�'�XpQ�M@�~���)MI�'V:~�D� ���Rx�D��qz����@�t�0ڰi�?�s+�=n���J�29�I�C\�l���$�p<��`D�; m9�-���~R�P|{���!N�Q���1�/,�����J�#��@%O)Ԍ��"�|��Dz�	�a�
��Z��0������'�4���A���I<j\��D�5Lt��Uz�����<^�*\R�@�',@�\f0-�5�'A��X�L�Z�V�@���~%�(@0Ĉ��ɉ:�N Q��Ȑ0��s뙊*P��ӯ�
�ՖVP6 s�-�5(���3̧2�!�G��tѪ�-ܑBD�ȫQ���G3p +K����	d4O�aZd�3?���<Zc<�%�J
�BRKh<�w��VX���@c��y�&�*5�F�YE�R���>�	�7�®�0=Ii����-��Ǉ:6�l�%-�\x�$���83�p��͖�A���Sd�D�cyLd��̘�I�6ݩ�	�X�<y��+�0i�A!�7Rt�	�U�	�Px`�i׫ؔr��2q�v�O8H` �D5�4��C'(bq#
�':(�(��I4Qn�ċ#+��?��CR�QE�lCe�O��?��k�3����>�Ah��+F���⃍-x`�B�I�p�kuE����R���`pp'�P[ �hAωb�,��鉅	 ��(�w�@�m�����<=��f@+o��I� ��N�PSe� H�	�D�K�ld�C�I8b�:٠�M^�S�&\bRo�;`�O$TJ2�G�8j�3����H����b��q�
yB�@$)$�u�%"O�9:���@V��hA���'���#ݢQ�~�	��̀hR+̐#9�g�t�v(��ʒ?�@��*dݔ%��I�oΘ����A��XꦇHh��+'^4�a���ox����ݵ@�R�,�&�Ȕu�О+ў`'�/�p{�Ij�';dri#%j"�\����?5 |�����Ǩ�Nh��PL��>��I}�j�G�-�I�������1����A�AU6P��*:D�
d+QW�|	4#9!�!��<���P�B�4��f��0<qA��n�xu�fIѝt�% �$�ix�,�d��d�>�ء@�-qv(m�r��$�
4�!��9Q�h�Ƀ���<�/�"�ўT� U�4��I�PK�i�'@�l ba�
�0��1�o��~�޼�ȓ.�QRA(Nf�d��C�,8�L���%��|0��#;8�Ŗ���( Rd
CܐI��4}�3��'D�����;6@�	��S�~/�쪱f�<�d��LV����F�0<�-K6@�����H��a�@����� �j\��1��j�4�P�F�"��|�]1z���7��l�TJ $�����G}bc<p�r9X��	/߼!�%dU�JH��f��4I<!�� t��Z�6r1I��U,.�<V"O���AO�+yV$��5[�����"O�8�V��fvpp�G�� DVT�"Ojx�R�	1�2Q���ox���"O4�W�ٯ!w����]?u���"O�$�V- )spʬ��fA�$f<4C"O\��%P()��+�/��Sd"O
)��a �6�p(d�*�f|	G�O�����á�0>A��(lb�b��_~��0��j����#TC2R%�	}|����hX� {��k��պ	�.C�I�Tm<�U���<��>W���$ҷ*\G��l*`��*RH��4�כ\��O�p��B�o��B�M�.�5��Ͼeܙ����(aר��I��G��'����Q+=���3�߮6:`+��Dݿ29n�ȋ�Q���D#�؛+eVU ՠ�#���5'��"��E؞D�tJ�Q�@�iL1x�Q
���O�A�M�c�ĒO�S`�=���0J��V�׿%F(����Y*`j�@��y�	Ԏ S�R��"p��YP�ف���`���΂X�T��*�+���哕!��		G˂v)���ܣZ����D��D�B����;_���`c��H�,�%n��?�<�E��
<�`�d�>i�鳟p���	+y�ލ��խ7�ɹ3#5ғ���*!�G�B�?}s�O5/�)(u��$�8X�.�O��x�B^Q�"E:ۓk�*t�GI9m�p�ve�fQn�L�Qg�ݏ<��S⓴*��i�Ȓ��ܳD���%���2ů�/a�͛�E5D���/Cs꡸'��9g���
䇡>��E?k�;�L >���C�T>��!`ݿdUpQAg�5�rxg�=�O�:PN�81
��� ��NӶ���l��m?��p%�M��8�P<S L��%���B3.�GzR��h$�@��f�'_T9�� ��2��i��G��l�ȓ&��؅���Al�RcX��oZ� }���,>Q�S��M��)��G������	���v��q�<�w�޽(�UA"��.�v]�4�l}��JZl���dx������H<ʐ��#P�T|���0�Ot��gP	8n��Ň�.;ڍ�0)C�	ԉ�E/D��	&��<l�&P��OJ�I,�E�v
&�>��5���;�'Y�nBg��c.���2g�~E��#�,<�2�P�Y�����G�$v̜�ȓz��)y�̚���$[4C��&�\a��Uڬ��KH�CoH�Ae�D�-�Q�ȓ2&tx��
�����Ӈb1�j<�ȓU��{d@�1rъ��Un4)-���ȓ���bJ�$Ҏ���e�2T��$N�ի���t2���l$�ȓl>��ǬЖh�%:���=|^�ȓf#*�t����d ��O�$�~)��8������ U~Dѷ��0Ͱ�"ObH�� �Y�D	9m�$��"O�H�h�����`B\l�4�С"O8���IC�G���U@�z�����"Oܘ����02avY����-�6"O4��&HHiX�YK�c@(�T"O"3a�F%[�")�C��:��t�1"O�482�5i��IKBb	j�pT!4"O�I:P)��}����^�w���i"OE���֙?�\ ��)P�q"O��ђoC��& Y
diz��"O��-�;�4=� e�;*oV�H�"O����=d�}ZĪ��aNJ�W"O��1D��$�Թ*�B�R �er7"O@��a�ͩ?P����A)�A"O,d�0��hU�x�D�Z��TBg"ON�"C&:�|��@������"OL���)Q`��B[�g�2���"O�,;�nr!Va5Ǩf�l�R�"O� ��t�-.�X}kV�_�j�t�"O��� ��;n����툒2����"O�P�6�PNL����ק)���"Ob��O�3~��{7��!.�,���V;�6O��v�x�C4�Z�'[F�ɡ-W�<��60��A�ODS�:B�ICl����V+��<�!�13J$B�	&���c�I�rV�i��cFl��C�I�z��Ct��L�p�0d�d5�C�52���`�W�
�*92W��2B䉏.�*MI��)Y@i��E�[�C�	�Y��!����� e@N#e����DC=��'�Q����Y�&/�$+T��ʮO
�h�_� ����
âA�Dƭj-[�Ŝ�n>\иaZLubآ�b��e\�]���Eͦ��I��dT�穂/J�)�"ܢQ!Fl@�a� �(<�����S$
$���oDGk��#P�(p0��P��)Q�D0x��ͦ�%NU��I�6	,ܠ����3C���Ľ9�Vh���M���svH�@���''�?�G�4dY ��M���I�S׶���VbB�ʚ_^��3eMK�1�hq(����� �.��i=@@02�Z|�L|z3m��r� ͓�#D�#�����dӤ#}r�O중
�j��u�̰�e �8]� ���nZ)p���QG�L�]���u)�0|�@�VMw��g�/""�T�ջ�p�`�&;�z�;A�W�t(��]�t��Og�4�Vկ`R�	 �N�	���'�|�bm@(t[4LH�O�>	�u��0���M�%�K���^��+������]姈�zם�F)p��4v�aX�Gߘb���@Ԃ��'	`�3�/��	��a�>�`V��!j��!���"��'I�1���0�N]�r�#�����9��0�>i%ǋ's/���?M(�g��R&� VT2$h͝�E�Ē�<�NjUB�)�'x��C"˸<��2#�gG�ȃw��:<%��s�y���'ֱ�҆�7e���CS���]�'B�௉�7URC���j4��	�'�0�`1�ƪR��R����:%��J�P��o�`n�aifN�l'`�ȓ9���B@AJ�S���ѧK�*{�l]��N��FE�,�6�P7��=�����W��h��6R"�����NR��ȓ �U��� n�q�`TP���b���s*S/7ޝ�VBT�e�ؼ�ȓi~�|��
[��)�BV�p *��X砄ʆ�*s6�a[bاxD�����$�B��bA[�jۇ!��Ɇ�N���b	 ~<#Lx.�p�ȓZ���L�%αKa-�(����=����ϙ;&ྍ��/��t@���& H�I�&04n����g�Ν��z��+`j�V������.�h��ȓ w�8�A��@�9Ѧ՞>�Hl�ȓ>�T<�@ ��k�J�'k֘G���ȓ�z<x���A����FJC�`D�ȓw�� mWM2:��U�D�T��E��B���QC��x��G�C_>��ȓa���"�F������1J���#��|�f��z`�i��nH�:���ȓF��0�΍�vUL(�b
�joƠ��SPj�wn�#RN�󃦊�a�ȓ>
�.܎q�aB�99��5��U}�<�q��4�^�j���e�����JR�<yՋ��MMNqQ�����5xZL�<9�� �ܵ���I��AC�}�<a�!\���i� _�($��!\d�<�s�J?
��z`m�R�)S`�<ɲ�̱_z��K�-ґm�-�E�]�<I��L�d��@�E�'���&�D�<q�Z�Ֆx��"B�:�Q# )�V�<��A(tGdtSfA!����v-
P�<�#M��S��4R�Dw��4���O�<� 4�wh[�l�&�1r.��hn���"O4�!�cc"A�����Lgx��p"O+r ��A!x��F�ͻXW�i��"O���"М7�r�bf�ƪ@L͹v"O<�i��΋H���x�,�X��H"OP�+�눴s):c�Ӭ��1"O2M�� �h��4[���m��-Q�"O����S3o,�C��-HA�R�"OT�"J�A��q��6x)�"O���1O�j���ƎtYr"Oj�vK[�A�\�@Ùr�f�xG"O���1d,�=��/Y�$��h�"O2��d�Z�2eX��P=Z�n$!7"O|}I��S�8��I��+$�X���"O�����8?0u6�Y*%�jH��"OJ`�!�?!�\���'�,}��T��"O*Yt�B9s�Q�W@�9��y�F"O��	��Joݴ��D�D9(p�ABd"O����Ô+��Oެ*l�x"Ol�#e��)f�v���n֕ki�$p@"Ol�q4L�*[�e�����-��x�"O@U�w $�X0��B��(�5"O�UQP�\4,�(�gA��K"O>l��ʙ29ve@C��>��3�"O&��0�
�)T��'_��q�q"O�$�b��c�Vͻ%����p�G"O��"�ٵQ�  ���A�z�PC"O�x2�ݞ���$��D��� �"Ot1���������<��t"O6���m5R8�
<���"O��%'5��]pE4xH��5"OH�w��!�`��'��}�B"O�x"IJv��p�W�B"B�e��"O�\�sK!�Z%����n���G"Ot�@Fm;.
=RVc�b���`"O|��T���Q�ʔ2�*\��"O�*$�&AZ��B�ɋ�Õ"O�噵�T�n�1�tH*e�r�)"Ol�r扎1[��q���L�٪1"O-�C@x�!@nL�i�����"O��p�ӝ��a��O{�ʍa2"O����þ`�� �� �h�$"OpE
q~��qk���9��� c"O�IB�p�xl�c�AhѰ!�"Or�jt`W�bֶ-�6���]�٣�"O�Hc��@6��6���+�&8�q"Oᐵ�V��,���'	�ΰ{"OF�T��-D�60�3CVI�蹚"O0�
1n<���Ũ�|�R�&"O��4�C���@W��z��"O�ts��,)�X��a�])i���(�"O�ѣvi�Cʰ ���ӽe� �"O�@�_�`
�aB5/p�C"OR���kI馠ㆁ�8���
"O�q� <���!+
��k�"O>%�D
OG e���ߴm���@�"Ox���G�^�p7B��Ƅ-��"O��#�S	^a����aK��2ie"O����j�%�X�����j�RŒ�"O��i�#��P�����].g�HE��"O^q�5��3g~h���E)I��!s"O�����z&l�����9�2E��"O���D �.J��b�"3"hX�"OP�Y�(U�©�b�SYNɉ�"O� @��G�edI+�e>�U�"O�����^� ���ߤA�ޅ��"OP|����=}�L ��ؽI8j���"O�U��%L!o�>���T��}r"O��Į$�R��1$�b��2"O|e��K^0@�R$Q�"�+X�^yr"Of<����@�� i&�L�b�<E��"O���B�ѤmI�\b��"ONqY �9�f� �O�����*C"Ov1�V��;�i��F�D�"O�y2��nB�����T���"Ot$�����w��Z7HXH% ���"O��Ç!�0�a�H8e�R�PA"Olm�����6� �[=b���"O�9r(+�4����5W��`��"O`�1�� �5F��M�1"OHu��k��Q�CΗ�W$z`��"O��a�ע/�bE��=q��x�"O���"�{�,���KұZg�=K�"O�#��8�N3�ݽjI(m��"OX �UH#�d�M�
BL���"O�l�W�4`$Z�nʁk6@���"O���,݈8���i�.$*��"O����e��X|�w��}t��"OB�(׶���AT�_�F Y�"O���K���QI��1�@�"O0}8NJs��!�LUm��X�"O��5d��n���z���X"$�"Ob��ѯ�W��hkA`�.[N�D��"O`P�vhGF�`T[�nM�����"O�A2��^�g�jd@f�](B�B!��"Oȱ�4X���,U�"�C�"O2q���]Z�J�,֞@GM�e"O���g�ϴP�SB�	59�1�c"O���IP�.qiS��=�����"O�Y�c"Ōi���G�jI��"OFib�^ )M��iD�۩xC$%� "O�9�����d�g�CE���E"O�y0&G(Ř��v���Y|L��"O2���^s��]prE�/<��"O��Ag�	I\|�y�c�2
�ԉ�"O��eV�&�*}��B�k&4���"O����ܼ@��i�ҨR;l�}S�"O��9�ĝ.bo�A��g%j��Ag"Oސ�W%H3<�&�X⥃�N8��"OB�+��W* �@ے�K�N�x�"O���� !>|T��[�a"�"O�"��M�Z���+U��6|C5(B"Oʔ��l(�@4+Ffчa��ҕ"O����Ιy��xa���`c���"Ol0+��	y���d-M�>��I��"O�XRą
�乂4�d�`U�T"O]P����r;��D�фp�T�"O�\;�Y
Kߞ���(D:��9V"O��Q�f]\5Pw��b�`�"O�X t�O�%a(�p�G�_8FԊ�"O>�і��.[�� �A�>��S"O2��ы��6pt�ۧdQ�!�����"O����DZ2L����b��vr��p"Ow&F���B��;�%`�e�J7!��P=L�����83� �ɊB!��LD�u��M&�x1a��&,!�̑D�Q�wj��x(p�$&�8!򄆊���.t��飏_�'N�0"�"O� R�J� ),������s%P$��"O`d�3�Կ!�E���z -��"O��r�jւLDЄ�(j��"O��@�"��N��#�kƖeҬ	"OD�� �È$@�kV!�
E���"Oh��� ~�R<���.?��X�"OR1j�/P	y�йc-��U,��qu"O@E���,}�]��F߲<z0�"O�LY�I��8����
']	�0�3"O<��4�5=z�#�&�i�l�1!"O�U�b.�u�bH��ň�j) �x"O�u+���@�^��W6[�к�"OV�`�H޶VD��d��`W�Py�"O(mH��	��r�c�3>�B�"Oް�+K1M88���	�T��'"O�h���;+��<�aOU�y�,�{�"O�� ��t�����.����P��"O�u���M��3����T�"O�Xtn��7,=�p,ր	��@(�"Oԉ+����t����$����2g"O<���n��^a��)A#���� �"O�`��XY3�U�w����&�+�"Oj%�AY�/�1�m�	��肃"O�A����-���*TF�ָ;w"O��;��N'^g��4��b`Z��"OXh��mXF���aC�J�=J� pB"O�UQf���&�X �I= R�	"O��[��ʥ/�d1�ꖝw��  "O�E�bC�?h�蚤.�n��"O�L�MǙ_�zL�R&�}��uɔ"On�p�:ɠ�IŎC�]~�c"O0�R�'�w���Y���Sj �0q"Ot(�A$]���Q�藄jV()�2"OLM� 
  ���M�2v�F�
�'g�Y#׈ִ6�8B�	��v)�ؒ�'�
�iD��9`�xbK�2Fu �#�'�� �X�ش�Qb�ލJ �Z�'I�0�O@=�<0�`F�uR���'J�����%��T`1�o��@��'�H�Д�ڀ:�� �p*��}�Ɖ��'�HM�7 ��%� iڲ-4,x x�'�\�h���3p����"e��%oZ���'8���������Jy�Qh�'CA�T�*;]��ӥ���g�eY�'�X���%�(����i.���'i  ����22>9���4{9*�
�'>�y!!lA�)`d�6%�9g��C
�'��	S�+G� za�S��gy�X	�'�*�!��Δ`��v�LLZ�$9	�'�@�Jjm�M�-+�hJ6�@_�<9f�&	}����O�	�Y���F�<���h�V�Q���v �b�Z�<�q��r�&�gǪx����s�JN�<�����p��D�D%k��(�B@�<1e�?LI��Hϵtt�[��A@�<�˭
~ �Y1�ƭ"vأ�	�F�<��J3�J|��"ȫD�D��v�D�<���яU��9R"W%�MC��T�<�P�͋U{�TZ��� T(Vȫ��L�<��ˋ��|������Lm+��L�<�G�̳:�ҹz�ЀX�-�F�<1��A�2fθ��[���l�n�<�a��H#$9�V�?_���K5��k�<�wG�I=
uٕ��>q֊����i�<���'�i�`K�#Wbm�G@g�<���1k�ޑd嚀+]�M��H�\�<���]�t��y��|�j�J�j�X�<�#��,yȡc��N3kI����K�<q�Aj*8� ��<Z�	� WD�<�kN��,��@-sf�'eDC�<A���T ���+�J̘Um�A�<9&��b�,tȃDK�C*���GOF�<q��l�ب�ʣZ�L��R��@�<R�U%,0��׀�Nq��[�a�X�<q�NV6���a$�T>)3E��G�X�<	F�	e��	�`(�0P��U)�,�m�<qg�[�o)��.�3n��4Zm�<R��VӞ�A����^gN}`���^�<���j�X����I걓���\�<Y��	gX�c��n���%��c�<YeN�� �J)@/���1�R#_f�<�''�>8tAZ�	,W�j�!��F�<9��!`aN�k����}�F!�f#�<�`�Ґ6�^�8Bc��U2�PS�
F�<� �(B�g�>,�^=[�%��j� l�"O�[��AW��V�B,l��MKd"Oĸ+V�T"J~��CM� ���+�"O��0�NV	t�	Y��`�"O�e��Aĕ8�$uQ3D .V�ʈ�"O���K�"6Rس�w�r�Y�"O��MδTH|�A��Tծ�x�"On���h"f�C�j�t�Le8a"O:A*�o�d��[� ��j$ȃt"OPl0nA/\_��25���]J�s "Od-���z�IC4��{4���"O�����Jy��a�!�ĠG"OX	pmSFƅx��I�-�VqY�"O�Y�d��,䭢���8@���"O�D;T�I0{9\��C��%&�r���"O�)�5 
  �F^�n�Ld�M�6c6�'���'Rv�1��'��'����/z�45q&�9!+���K)k�V_�H�!���M���?y����\��X�N:L�:��&6Icr�[#Ua6m�O��d�5F�(�}B���*��dK�.݇�f�ben������@�!�M3���?��z�]�Ȕ'�\a����B�<�(U��0qt�#�y�n�!���O��Ox�?��	��ĩ;CG�b��%s��$�����4�?a��?����[��IJyR�'����brp�YR�_FM~����h��O�E!:���OH�$�O��)�d-Jz: �ǥ\	F�:v�צI�I�L���0�O���?qH>�1Q�"f猆|�B܂�ć�]���' ��y�'*r�'?�I�K"D�Y�$<����@N;C8ݓ�g�/��$�<�����?��U������	��|�����X�dN���䓁?���?a)O�P��O�|����{��؋��G�I)6h�@I���'���|��'����m�$#�$l
E-�?��5�VӞ+��I�L����X�'��-�`I�~����p��c�YFm0i�5(�|���iY�D��؟x�	�a?����dH[�+��\�*�T���ϟG����'BU�*!����'�?q��c��!<�Li�B�Kj��2���ͦy�'���'L2�'J��yZcŸ��ȋr}L����@p ٴ��D='�}l�����O��iG~2	I�8)�ⅻ8DJ��)�M+���?a���?Q$_?5�'��s���2/O�v(@�T�8<-K�i�R� ��'5��'c��O,�)�2���T��A���>H�����@�>d��	b"<E��I��X���o��|"�'��Y��7��O��E����,O��r�$�<N��=K���=�� ӑ��6(1Dx2�:�ݟ��j��Ub<Ҫ�S�)�k��umZ؟�R�euy���~�RGȨ4h2Q�u�C/PKD�x�޽JvOhu�$�O��?5,��DF<\a�B�W�,���H�:�@,Oj���O��t�	t?	�G�!o��I��n,W��`pA�ܦ5�B*���'�2K��:���O4b�Hd3b'^R��(� �����'ER���O�˓y�l�= ��a��Q�p*��#R v�O����<a��s���+���dP9;���v
s�ڀ�Ǻ@�Pao�r���?Q.O��!w�xbD��ZNYCCL'k{��a�0oZӟX�Igy�%ȑU�D�����k��(� ��,ǩn��#lz�'�������	G�s���
8��m���M�ᒶ%�)HT6��?i���4�?����?i���*+O�O"O�T|*�\.��Q`(�-����'$�I�<Ɛ"<%>!`�AЦ+o���Vv��i`�t�,<�d��ᦝ��ş����?� L<�'���cI�wc��i%�%k^Bq��is2�'�r�|ʟ�$�O�����"�n�c�ۧ`=���G/Pߦ}���t�I����K<ͧ�?Q�'��,y�MW	4�P%{����4�?�H>yU?��͟t����(y���Sd�� ���������o����I��7���|B����z�� ,*&L��Z�!"��oN|s��x��'������Ο̗'͞�v-Ÿ&RM�B,�NOH�$d];`?TO��D�Ox�O��Ӻ �?+����Ǆrh���������I[�����'=�̗�T���E
+�([�o\�}��}ðO���&�';��D�Ov˓r�Yo d���e��{�G�cV���?Q��?�*O�A��,�b�ӱ��h0�MƖ �V�x�]81)�4�?�J>i*O�i�O��Ox��#�×06A`Sᑝ�a��4�?�����$N���Or�'���;~L��ʚ(Zz�;��R)����?����?�"`��<aM>��O�L)ś�ZRB�Z���E�F��ߴ��D=n�T!nZ�$������������a��ς�Hܜ�4�1g�h2�i��'"89�'K2[�l�}��ðZ�X�0d,!6�,��d�ʦ�0$l��6���I�H���?�#�O,�Âi6�
 U&lht�N Jp[E�ii�[�'�T����L���Cӣ�^P�%��J�6����u�i]B�'��� sF�����O��	�< 1ȴ쉏D��z���X��6��O�˓L��S���'YbޟN�0HA�NwxMzdf&� �KӸi�O�2Iw�����O�ʓ�?�11����
�r��LI�����'�!�'I��'2B�'�T�l�'l��O���PE�\6b�Y���h�d(�O�ʓ�?�,O���O�dS.hV�1�ElD�7m� ��)�j�xQ�5OV��?���?Q)Ob�t�U�|
���8�4Hpƛ�F�:	3�!HҦU�'��X�P�����ɁX��	�+�~�{T�-'~��p�[�) �ۮO���OX���<1��/'�S���{��V���؞�%p2g�%�M[����O.�D�Oȭj�;O��Y�1�,mX�����$+$I�E�d���$�O�ʓ.z��X�]?���ʟ���4ly��Yw%��{�lM��`��?�p���O6�D�O���A�4��D�|�����4O�FDB����3~'����㗡�M�,O�傂�ܦ������I�?Y��O�΅F&(�$N!Il�`�o�I��^�F�'cX�Ø'� ��<���4�߿"^�X���G�yݜ�͐&�M��A�m�V�'w��'��$b�>�+O�1�HO
���E��_�X�@C�Ӧ%s��t�$��Py��i�O����b�x��p5�X5tH��a�Uͦy�	��I�;h�U��O��?1�'߂�����5�h1����8J� @�4�?���?QB,��<�O���'6,/���-�?��i�׬�RN$6��OZ�Q�GBy}bT�0�I@yr��5�"[���D���2~��������M���6	���?A���?����?�+O
��#M��4�נO�Z�ͫ#Y�g1"��'v�I��'w��'��ک%�ViX��W#��NH<`�P��'E"�'���'�BT���P*���ĨU9Q��ڲ޼9�p��@�2�Mk*O$��<a��?���x�O�H8�6J	}���g�׎��ayݴ�?��?A�����/Ky���ORZci�1��*�=t~đ* �<nm�ܴ�?)/O��D�O������	v?��n�!`��	�GF,U|�C���������̔'���z7��~����?���U������8��S�Ν�G��d�vX������8�	C`@�g~2ݟ��{�ʡ;P�(<DL�i��Ib&��ٴ�?)��?���<�i�q�g�)�(�H���O�$�p�fr�n���Ox5�;O�L��y���K�o9���Sp�m�j�4|ӛfό�`Ԛ7-�Ox�$�O���s}B[���A$׽��e��,A�b�.9���2�M��.Q�<����>�S�����Q�#;��"TA�)�0B���M����?���{`P��[�Ԗ'�r�O$8���ВWǴӧ�]�FGj�r�i��Z�\��+i���?9��?�����|�ĆФM����C�Q�
,�F�'�^u�4�:�	���%��(Xz�����V�)Tk��5`<�iD�̓����O��D$�I�$).�ՙu蘪���6�7#eȰ[�b�]쓂?H>���?��N�U��u�H��WX��B� ;d�\5����O���?�	ƫ,�@��'<���;�cK��L��y�0��O��O����O��b=O��S5�i�ql������H}R�'"�'��	 x�-�I|ZGd�P�<�P�%R�wt0zAi���'��'�'P���')�Y
�{�h��I��h���C��oǟ��ITy"�������D��*̣�'��5R�H7oրx..}��Ty��X�I�v*�k��iJ5�M>��m�MшR(��t!�𦱕',�0K��Ӕ�O���OR���<\��J�	ՄAȆF2閝n�ǟ���}�`�Is��pܧ�`0ŝ"o�l�C�(B�{�8n��&e��H�4�?���?Q�'o��OݘC��ns2��ü1�"��f��Q�Ս�`$������"dy� �_�q#1.��4�x�!%�i*��' �JP�4\�OJ��O��I��
�Zb���������f7-;��A�'��&>M�Iϟ���BSpI�QE�+R �=��-�k���ܴ�?�t��[Q�O���4�����7��2�Aq�4��Ѱ�W��c@�ʟh�'�r�'n�Q��s��0�h�R���f6�Z�][�K<��?�N>���?��AU�@�`�H�D�i�
�*��p�p̓����OR�$�O�˓J�H ;�(+���k{$��ҒN�:��Q�x��'��'���'Y��9��'��� �Ui�H�##͊<����!آ���T���ǟ���gyb�Og��ҷt,R�$�42倔-��r���ʦ��I\��˟����<�0�W�D��o�F\�Cc��GP��j@� ��&�'Q�X��11cߍ�ħ�?���C���\�A����!�3d�a����O.��?a��P�I Z�A�R��)�@��?ɀ�F�?A����$��$�?��T!S7�"|`Ή�U"z�� �d�(���<�&�y��ħYf4��򩘿q�:���#�A24lZ�m=<��ߴ�?���?���d��'I�m��Lj�Y�7���E�9���$�Oh�y`�T`ԩ�W��j[�`R��T�������4�	�|I�x�N<y���?q�'�����]2;gP��o�r�&���?)��?i� 7-,,���'���Z=����'=�{r�#�d�O���4����@�@�D�Gp��@�T˼�RT�$�6�?�˟P��ş��'�~J�dG�
�fP�A���z�)χ(4�pO.��O@�O,�$�O�l�'��.�x�B���9 H>e8@!XM/1O��d�O����O>��-1����.&��@�5Sg��ya�C�|L@LlZYyR�'�'4B[�|c7Kb�%!e��q:9��}]%�2l{}��'��'"�.K���I|e���x�4`rC+��q4,W��9��'}"�����*�ѓ��M&:LR�L��Y�����i>�'"�'�����'��P�@������I`��b!�\e�r����M<�������4���]�\����o<ɢ"�\M�>7��<�V�Rv��~�����`��xy��5vJ�$�VLM.pJ��։wӘ�d�Oh��q�'m�����%V�? Ry���-��n�$P�l��4�?����?���q�'��aG;m/��Z�@ߒ\(�5z1���$r87�Zp�"|���5�D�Ĩ�)=0$��*�":*�S�i���'��*��Y�lc�0��b?�A�U�8����]�e�ܽ�Əf�]�d��<y��?���WA�i���ˏ$N�!2�)ߧ�,�#�i����D>8c� �IK�i��9Bo\	Q��j��L�𬂄Ȣ>Q�]̓�?����$�Oh����G*m��C��P!S&��I4�҃)�Xʓ�?���?�I>����~BĜ�d����L?�m0s��<�M�eKD~b�'���'��ɒ�i؞O�&�@��mjT���݉(�:m�Ob�D�On�O`�d9�� aH�h��^�e"8|�wۏL�H��?���?�,O��ѤL�G��$���ȓ���]�w�;j�z��ݴ�?�J>9��?i�!�|�kf��雝t�D9J��T�Z�oZ�(��hy�!M�3<V��������BGl�2�����I��Ir-v�	�����'�"<Q�O��,��.,���1�*P�5��	 �y��\C�F�F�����'(.xA�OdiY�cA�t��3�e,jz�"O,�j� M�6����rI\���*0�⣩O=g����W%�0@�b�bI-$��$���faJ�c���$,9��:C���vU�͋S���(y�PQ��G�	0���ҹ2�R)hR�	?�V����ˇZZm���Ϻ��FJ��V �Q�B�*���h��4^�Uzt��,45��u4������G��?1��?��4����O���0�`ͬ�@i��P��-[�L�l�`���Q�"���hc��넝9@�9����&��2{�ȳΖ�xȣȍ�j;�hc���������XD��$�d��0	Z��@eR���>;�`�	�a�^���O��=I.O�hV*Ϛf����a�&m0�Qp�"OV���@��h��z��T&\�� �ZV���ɿ<AF�@�4'��d;
��`T�M2xX���'[8C��'F��'1�U���'�b�'YX ��<NB��9�f�)��� >X�D;w#�+�p>!�+��D�N����y2��R� ��X�!���Xń�I������O^ ��ɝ+p�� e�Y� 2�a�+�$�O>��)�$:��Ͷ!rpt�A!��6�yթ$_�!�N`��Ĉ!k
�)�H�VI� U��d���IXyb��KR�ꓽ?�)�Q8�:1od��/��X���*a�G_a��D�O����:%��x�d�#!'�)���G��';��$���H�l_��Q��@4Y�&HGyҊ���t����L^>&e ���-L(��x�I7�z=:�k��(Ou�'2��[v�9؀j��]\�#л�Q��'��
�5Q�m��ѭ�P���0>ɠ�x2E���v΀�4'2)�C���_�*��}��qCsZ���	_��er�'3B���Q̔a��JD�6�@r��n4�4�V��Xǈ�H��R}*�Pc>�ħc���0�3�����B��( @<C������RQ�������On)j�ᄝmf^=p��.x����V#w ���O��S�^��

D>�ەN�T�ν3��
6 B�I�R�v9X�c�[e���3�z&�"<���)�d�R��uk��ĳ�.�3լ��<�p<@z6�M��?i���?1��i��O�ʿb>-J�+��;d�TI�+>$����h��}"��)�Ѫ7��<O�����#�~Bl[���>� �4��m�-L��3$Ɲ�[�����O`q���'��{@T�4CI٥IH0/��}�����y���"R 9Y�� (�f�h\�4�#=E�TeC)2�
7-��J�@�ʗ�<��1$�
.'�$�O���O�*ub�O���}>�b��O�d�H��St!Y5L�j�r�+�|r�ǖ���20"bc�,/��]+�O^(��|-X?�?i�t۶��RB�9Ay2�E

53F2\��X�<���%$ܠ�A�@.� �ȓP]�4 �u���!�!R54㤼̓_ұO��{c��Ԧ��	���O:���	K -�!�' Fd}�a�'�J
�r�'b�fҽK���T>�3�Ƅg���S%h'\p����;ʓ{&`�D��gR�c���!D���а(�T�C��8d{b�>#��XQ�K��<�5���V~C��O_֜AG�A7��݈�C��df���k�	/o����$\&Ez��@��к73X���tmZش�?����)�AOd�$�O���3U�,l���3<f ��K�>-*&N�O>c��g�'1���w��V���q�E�*2��c�K��"~��m�rE"�C��\��1��g'j%�i��,W�T�<E���x��f-לz��c��' d��G Q @�0����/�N"5Fx"?�S����5{�X4ct�Ł57�lJ�f�A�"�'�X�:Ӭ��dh"�'���'5���؟��2Tp�a؂k� bT�·,{��	�,����d[�;8`1��I�QrU�q �2kn�d�*�}RG+w� X�c`���(�wEB�~r@�?iߓ[���D�ڥ �g��E�4��ȓ1׀�q�(B�R"�d��3�����)§���	c�i\��jW�>�H�x�,��O���'�2�'�rk�xVR�'���C�%�r�'��Y����6:�A�"� #
�	�w��'��q"`2m���&i>zxv��	�J����I�X�qD̏xzTҀ��=,��c%D�`��mاl69i&a�?NY�-�!(%D���uχX���3���Aт��m����}��©$�6��O*��|
7�Q�P��7��+��xVa�iraA��?���oR�����Ԙ��)�.UF�s��Q�H@I��	Q�L("�4��A�B�����*�c�7|vDy����?����'G�vxr�lҪC�X���Ӳn�!��5J܈����2fiJ	I�a|��/�D�;���%J@;Z���3�,20�$�*m� ��'s�R>7���?���?i�)
HL~�ڱ��Pr�L1����|��7"�*����a¬7Ҧ�)�tb>��L/R�b�+��<��m)5�J=N?̴[&i�:1�́ɒk׍d�6P����O��x̒F���`��;�l�c(��~�'��)�I"��-J��d��h��J���cp�!�G%l�*���f��*s-^"�8���?�#�b=0T
*�J]�r���1��J쟔��2���qG`ݟ��	���!�u��'�"o�"��R�N��#� Բ%N4�~�*����>aE�@s�j���o��D5�l��H?��Dx���W��h�0,�7NȊk1�8!sF��\ۄ��OZ���Q+&��%�&H$-�5�vo�l�!��C���pw��S,n��ŝ�z�©Fz��i�>�8PoZt�����E�D�嬌'oj�0�I럼�I����2i�������|�*����	�s餘�F��e���E��<~����d�"���[�����f�
�;��PV���b��'�~��MԦ7�TCw�,<�*)�
�'�fU�B,ܸX)��i�U�P	�'�~aBQ
@<a2l�#���N�n�x�'Z�c��16o�M����?-����%#;g�	RFo<E)r �3'�!2z���O�$E�
��'�|j�펆F��5� ��Y� -��L\�'PH@��I�2mY��2�Ë�Y���ʔ*SQ��Z1%�Or���O�ĵ|z��L�KԚG�%k DY�����K�S��y2�m����ߥS��1&���0>aq�x�Mv��R׬M�=o�����y⡈�j��7��O��ı|*q��?����?yB�Õ����U�f�|1��E�/����������ɇ[-�瘚P'����H��f}pC��{����2��{2d��5���.�X1̟<S�x�g�'n1O?�� �u���#Dk������jAq�"O&$9@뀈��0��f���@�"�HO�:g	`�Zq�Afg�qQG�V<v�������v���p�nQ����p�	ޟxY[w�wf��$N!g�����VG�PQ�'7ԉR�qL���j��l��b&c ���t��m����2�p-�K^�
�<xɧ�Q�i���Z��+|O�Y��`��Dy8M��J�_�n��7"O.=ʶ͊�J�6}�t�Ǳ6���{u\����T�椒æE��)�:���0�ғC��Z�ğ���ş|�	�g�m������'`�ʁ��Ɵ�ؕ��-(��(E*Tx�kf�!�On�)�X�	7��	kA�ĩcj*@ =j��2�On���'N�� sV�۔C���5+�Y��y�g$D�P��2��-yRT��`D/�y .Y�.�a�˄�lDfP��&��yR-��a �Hߴ�?)���)^���`R�?Ҁ���k�+��y�%�O2��Ov��!��O�c�ʧjA&x򤭏�O����$�S�|&��GyFT���|�Dh�
Gđ:�'
n�����I NH��=ڧ`hݺ@���=�`��1�̌�ȓ4 �6����9r��N�����I�ē��z����{�|<aׂ��fE0��8����i���'&��/#Ȟ��	���I�TF �cB�9n���iA蜭S�e�U��O� �<�O��Oj�؀㏘l�8�AQ啦;}��!1��=T8(��K>�)��X�GI*��y3!��─�`�%y�\���IȟxF������Ǆ�)��Ըp�\�	J~!ϓ�?9
�\��Sd!�:�ֈ��O�LV�Gxb&5ғ��G � ��(��^��d�D,�2N����O(��o@�5���d�O����O�`���?q�W;�șFd�(��M��B1u��'�
-�)���9MF{��+	�@12J߂U(L�j��R�u�D\.�,�Ɇ�R�5��hO`�� �fm�mcl\"�ֽ�$�O<8k��'�R�|��'�R^���%�M������9,�IF�?D��ـ*W�KJn��]N�||b,@'�HO��qy��#c46���*�� @��R:���aX���d�O��$�Ov� ��O��$v>�r#��O��d�+�F��e@�+�$Dz� KK��|b����?� \
��ڠ����R�:��|R���?��&���Jf-\C�^d�uGрkS&ԇ� ���0��]�*�����I��Ն��ȓ$��=vFA�r�̀����=fK4����O�	���G榹�	��d�O���g˿:�V�κJ�${�gN>,{��'A���q��T>��F
4݂"&~�BAPj1�#��yD���ǝI�j���k�	"������<�(OF�#��'��>�Z���XSFBTq(��I3D��0��)��P9���J�6,3�6�O6�%��K!�;a�:�2�薟c�<Tk%s���V%O��M����?�/�XȨsk�O����O��#3����9�
E�j�3��X.����*�|Fx�D²���3���<Y���W$��RN����)�矔�u.�?/V�0ץNQ�e;1mF9\�"���ϟ`�	���G���$�0�
��Y� �4��#k�Γ�?��19s�)'V�ȠFS��	Dx2�&�S�d�޵0����MO:(�	8R��9r���ʦ\ 1VN�N���M]��!�SV`
�\�a��)_�U!�D[6e�T���#�t�`��rN!�D��a	DЪ��ӌs@��ز�0E!�,��lɤN�?6h����k!��$���k Ҝ 0�$�'��w[!��,
=<����%�IF&J�u!�D�3@�I��H"���F!�D�j��Y׌Y{Ҙ*u�,4!�� 9h�K�K\�&	��@H G�!�d�':N��Βj0akt�٠+�!��;��DR!�=�(=ɢ
OBP!�D��~t!�f8�$�R�H���!�$X#+L�u��+sƘ��甦V�!�$�;[�F��Wm�3S��t���	vy!�� N�z�#3�]��j�=SzB�E"O,���'�b���U ��z��%��"O��V�A�z l�S�\S�yz"O̘PQ��?����ƿ�f��"O�8�1���;FD@7��;� ���"O��H�#8��j�'D*^��"O��h'�#'2u�R�ƩP�Ju�"O�}��b[�>�V�0R�p抭"P"O��#G��"���ǅ_�A�����"O�����X�09���L���$"O�}`���$�q
�G�F���"O���A�1:���MK+��su"Oд�c�ڴ)�:����ޕzQ#��>�������O꼄�r�-kڒ�����!����'β0���Ȳ%(�UcB����yB��Ns�̈́�	9|�6XEΰ���řk�nB�	<6��#�!�+�Ў#�T�S�� ��}b�@��>A'��1�pY�C�N'�����)�I�В���<R����5	����H�<�s���P5L�iv'�Zo!�$�hJb��@8X��ت+;�I�0������fe�E(�����(�&^���C��:8X���p<�x �h�8m����P)
�Cx�CC˙%T6��K�q;p��]�g̓s�qdc�>�ȥ�#��5�hɅ��3��p�҅ۦI0T�X6�1���:7�[jݸL؀Kԯ!��<��I3<Z�*�f(a�tͨTȖ�HT����@w#@)"cW�>4e��5Ot����B-=4:�r��F�f�l�v"O�P
Ee^)���d�%����᝟�1�����l�|YA�!W�O�Tp�i����%�14K2���'#a�0Ώ����蓎vӼ� �� Hk���'
>�j3�-�Ϙ'�V�JRĀ+x�J�H�ܘ/��y�'?V�H��'J�XÅ#Md��{��-��|�c�������
Ğg*����Åw�nm��	=��=Q�G��>���cr�,��o���b��b����G3D��zǋ�b�<·�X,
��a��#�<�� �&"1(E��S�P$��F����n��RqJŲU��
 K��yRD���Iz�c�_����S�Y�j��`������M3�#��*0�W���}C	%h2L�Um� ���	�*��?A!,�2
Pv��ď�=�H��I��(*��(�cG�|牄?���	�k��H��Q;6.��'B�=`�"?�rN¬ڀ�u�x��W�(gzI t�I�V�Qz�O6U4�zG"ObH�$D$g�n�)� NSDk[�8p�\�D���&�'�$m�*b�>J��܊RI�l���Mn�@Sf�>D�hA�LM
���9F�̓!됙1�B���Ģ�&���?��9S����{L>bA�'6��zCD�9��� MDn���f Q #�A��ES>jn�y�m����Q6
�|�4�Q�7\���U�'�P�7o��}ƐA[G�K�`k���
Ó9�d�1����Yw�5( �A�G�Lb|��+8侈�Yt��B�	�w?�5���O�')6I3R�$�ʓ���� %�-��QF��/;�~q�S�'{�F����	�L���ǧ;���V�D Ub\��p�Bw��  Up�b�FY$�Ɣ��S� ��'�	�4G��'ORq�O �R�4��	��q	�b�����W�S=N JF
Z��IӁ(�)�z9���4ᤠ����]r���'�2I�mIQ�z��1,}f��J��Dڐ.ˢ���#E�yh`�1'�G�)�d�.p�)�Ǚ�;�X���Y�����'t��* ���s���s��n[���O�������t٦ŀzj`�X���vȋfݜLB��At-�|��xB�"O0)B��8fw]�u�)?:r��4��b��ar��e}��ǆ�ħ�,�𧛟��d�J/i1��`"�Y<���;�O���`��)\̎����ÍD \��$�F,,a������
i�<�J ȕz|���Ą�M��.z��(���y��\x��R6fS\e �$LO.�PF!�i.2j�W]N�b�AƷ���R�M'=� �k�,@
��'�ԕ[ 	��'�	˵i0i33���B�K"��c�1OB�I*��#�]�	�s�x�]��>E�Tk��=���Q盜1첸�׌P�&�^�����CN��"<pK�JMV��Aj]�KF,��@7$P��l8[$քx�l4�?6#Ҝ[|�7Ms�� �u�`фC�-��	�1�l���X�T�7�_e�ؚ�!ڱ!l<�x�� �i$l���*�D�X���1��I{��D92���Z���3��/Su�1S�<����P &�� ��GϪkZ4 ��	3� `�o�m���R�iM��X1��KP�;�<H �eTD{��9�t�'Ó�aB:�S@�X�G X0���I
T\����U�@QPV)޷�h�(���!4BQ��b� -�� �����%7a�T{�Dӑ^��m��<6��jP�7�����_jn�aw(<,O��rQ���v�Xm�N)���h}k̎�z �qB�}&@`���/~�F��#���Q C�ٟ�*W���j�hB�Q<XG�MVMĚ?� �>��;��_;n֨�7��t_��h˘cY|4/M+��B��Ll�
��'~ٯ;Uy�3��#�y�B��F�
b"��@��[��0?I�N�����Ul6x��2�JM��رiZ|�fa`)O�4 Aoߖ	�p���]%^��͡�\#��I3Q���Q1|�M����)X��#>i�+Z�>!�4�&�_�i1v�9����"5#Ul?l�X�%�E1`@�2���Ū�5!��`�4�J4C�d��ቂfa��x��̎Rɮ��v��,e�I�w���*��
�-W���Vn��&�6mS�}e\ ��"}F	�2��HHF��J!��ᔱ(�'?zEV!�	I�pm�q��/1z�Y�G4 ���'�*����@5�b�r�>�	��ʿ*nx���
s�XI���',$��'@����%r��ˎ7Òq�G�=�𤌁�ԸI�B��]�$� ʟ�m��I�J7��{�e!zv`E:!k�X:�">)R�V�5/�m @���dL�CW�<��Ѽ,}���Ď�	E���@�:����o�l(�R�� �1�����پd�� E���)�]jG�PCy�����v���6�3��ɞ$C�4:(�n^0\*���$̴��r�M�c �����wF\��ã
�Cj
����'A��	zc�U8���PWh�7F8`�w��a�i١p<`4wn\�(\c�`�"P�¶4c��
_���X5���i��	��'�$j�	���(}k&G�#Ul�J<TC�I��KaD��f�1�mWd�'�� ��F���ʘ8��}a�O�9h���5X	��h�"Сe�<:�.��6�Z\��h_�v�X�#<O��K��U�Zh0�*5iM=�*(C�FH�4HZd��È������$�ax����.I�K��n���AG�̠�y��ɵX�Υ���u
Ra3M]6rϞ]���:
��(J�%�5Y��]�bB���'iO `?�H�ħ��e������2��pV��� �r��SEC�x��z7���)�fq�,O☩c��4>n�����Ä��U���	Q��xg�� ;��sd�M*y�#=�W��h�^���l�=&�8��.�j}�d)N���A�=1Ó��	>�֑�p%P�[Ԁ���	�0�fEc�爯ls�����-W��"<���9Z�J̈�`�1Y�EI%�]�����!��2D�S�]|10uF�(7(�B�ɉF�bbHQ
gn����2z�|��UhTf��u�(+h� �s��i��?y�D�6J���#�̥ ��Ť�r�<)�G�"�*F����)K���q�<Y7�K�x-���S��!��cE��w�<�6�u�K��(Vx� B���B�I5�e��M?+�8q�T��~7�B�_4��ᨍ�
]�̳! �� �.C�	�#�z�H��["վ|�H�z�lB��V!P�D�د<j�����%i�B�I�Y�r<3Q	�76�p�ULE�	�C䉙&t�j'�\�/rP�2Mΰb�C�ɎV�еb�cMpm�΍5\1�C䉚cF��a�WN�рG�&5�`C��<.v-rR�Y@G�� ����@d⣢L5~إ 7�#A R|��+� ⦪�t@��S�"oP��ȓ&wp���L�%iиxG䞵S����do�	��y�S�OҢ���@O�	ꈉ�ѬK_�Ձ�' �d?��m#aDɟn�$0�N�����;�^i��"�z�1�ٕt^����S@�����1:�x�u�A,c��db�x�R �FcY�.O
B�	�`�HԘ��2"���'��[@�>Iv�E���É�$�[s�v�p�Ԯl���Æh��y�( ZO��s@_<]�l�$��~�lޞ���Zu�|�����I��"3�@m5j_�a!�Ĝ�6��@�l� �t�!)�36�&	�DCS���<���=E���E�$EX�9R�]��@�$�p�l%�!��u$?�S�d��K�� %H?R��=@th�5U�.�����t� z�Ǌ��5��Xt�&{s|�����t�hsA�A��S��{�'Tn��b0�G&P3��yG+�T�F���P퀷�@X���;���C�&e鶑��%6B��"�O&	7��'���h��aZ��G5��U��E�I1^\xUZ�4����6�8��T�{�ƙG��@�B���+��-X������I�YS��W�'��%hwL[�D�&�)mE�y�d)so]�rϤ����F��NA���gy���,��"�H�� c6B�>�氋��'@��Bb�8N����BkV�X�A/�"LG���ēJI�0SE����&�Y�1���EBL�3\��~�D��(��	;1���q\�Y�bQ�<I� ��Gʜ���N�9d~9sG�
fy҂9=���=E�$	�!2��Z��jj�h C�O��yr �-�dP��ᑜh����̦ޘ'��Q2�-,O"���c��A�m��P�}���ku"O�}�$W�6et|��b�8W���B"OhXP�NK��(s� �6}�Lc"O���D��&�|�� ҟlw���E"OjD;c���n�$��$Gt<��"O���G�4tY�i��5N���%"O��!�	4G�PW�@�P��Ѷ"On�:��[^��Xxހ�Vœ�*O�͠�D�0/9d�fË�w����'84iz҄M&}��`k�Πq�'�=�f#�<�^t��b.��
�'Ϝ��E.��_9X��n�c�8$�	�'uM,9EN 2A�L�D8�rf��p�<�#/%E'���r�O(+�&T�p��l�<�@NB�ke� %)�R5�ta�t�<��J�Z�x�ǧK�}4-
Ҧ�n�<y7-�)!\�P�g��"H�ţ�O�<��R*)��,36��~~e���P�<�v
ӓ{p�������� �E�<!��@:�(��3$e"�Y�'�L�<	W���`�-(�t Yg�R�<QT�T�K�" ��ʨb��b�Qu�<15
����}	�EB�}�ll��+�l�<���_�eO���'IB,b����&�h�<	Ɔ�2Q
��r6 �)(_��:���<�[hq��̍�#����'��\�T ����$aˉ=6��{P!���ȓrҤb5H�\@$܁�̉�Z�¬��yR|�s��߶G��й��V,�����g��� RC�f�����_>C�*]�ȓw��J�i5wb2���O�:8<�ȓJ���S	ك!�2�� ���R����"�dM{��Ղ]�r 1��oZ ȅȓ*�V��T���b���g�O�Fs0(�ȓ	�*��F�3
��JF��->g�i�ȓB 8r�AD�sɦ�A�c\+k�`��M#�qC���D�B5��(dن�w9"]�����l*����1l,E�ȓJ=�=oאM�HMU�$���1D�X����
+��(��Z0:*^��n"D�<w���s?�Mk͕J�*����>D�$z6�:U�r����<X��S�<D� ��H�����+ ��M	�;D��bb��Zn8�a5����s�7D�T�Wf�/\F�a���M3Cڪ�s��?D�h��)�rR24{ƌT5����+<D� ��+!_���4"��ss����E:D�8(�I�*#x<�#薱�X� ��2D���6d�3t��l8����($;6%D��1��6%W|E�5đ���u�#D���B��9P4�xh!��Tv
 D�� b`V ��R�h�C����3T$���"O9����P"ԧ~�T|��"O�zp���`R�=�T
�"O��\�>�2T�@�H&Ar�Pv"O��[�e�Z,��ɼ8Tʼɓ"O��iQ�GOV`s6��ZR�I��"O@�Z�F*?\Yp��)^Q����"OLk3� �\�b"E*���"O����*�i^���\#�Du��"ORA�oŅ,�С�a˽��M)�"O:uJ�)M�p��P�0M{+��y��*tfA���.7��c�D��y����C����+p��	�a��3�y¢Z�X9�pr��R�g�v%��Mߎ�yR+ϒ!z�X�oY�c[0jA�F�y�D�S��b�/�;l�ȃ�H��y��"_��
����hd�x�g	�>�y҇IT�.Qy�EExTy�J��yRiB���� q�Z5�L�hP���y2i'o�tٙ0�ٵ�(�gͪ�y��S��c&N�r��%8�#ͤ�y�D ���GꉮbBTS�+��y�qۮl[�ȿL B�c�E���y�}-�h �GA>Fw��Ї
��yR,2I��qO�C���� �y�Mpꀻ����A��(0���hO�����J�y Ȑ�i��$s�
�� d!�d�>�t(�l�]�d��)@�j�!�h�!c���S뺼A㎸_�a|��|�"X,&GNd��嗐iƠ�� ��)�y�)2p��U#s�4O�Q�!⅀�y"�̜r�t����H%�����M��y"h64����B�N<�X����{�<I@C�!dH� Bb��>��ȩa�<qv�-f�Zh��% 	n�� o[[�<�VhIv�B�2�S�N	�4��S�<W�ڀ
$fI�T#�"���&j�u�<�`�է:8�V�\�.)��Q}�<i�ᘱ?c (��C�%I���!l�a�<�ϛ>{.6��E�O$"�x<A/�]�<9M&�4�k��:[�\��ӋX�<�b�U!ͮ����ƸQ�<�q�MW�<�g�>P��ϼ�V%����]�<�w�1;D�ԣC@�=O7�A�ǧW�<�'
	]���yp#��f���-�U�<Q�e����=)l"�V�KO�<���EZh�2K� N@��Y�)�K�<�f�E��}Y���pR�i�J�C�<ɷ&�4'�.d9���>q7�|����B�<� �Pp�$G�_�^ma)T��Q�T�d!�Y}���/8D���`'�3x������tD�B)�hO�S�2�t	 ���>| ����3dlB�	�LЬ&��Jl�@�@B�ɖ{
�=�N�n]�+�;A�zB�	� �T��t@�*�	���	3B��#$�ɐ���H��B�׃��B�%;��d$\n�$���E�Z\�C䉎;"�0S�mЯL$���-B�b	*�;S&*"�<D��C�C䉴�E�����Xyp��-��B�	>}��b���;)�-�:�B��"$@�[��L)�Xa���3��C�d�xr\b��<�3`���C�)� .̛�đ3\�LHs��%<�&U�"O.|1�$�#���)pC�m�q"S"O&%��E�w%x8SFb �8�Zu"Ox��L�,C8U7!E Yҩ��"O �iFk��&	4�rр�,<�Q��"O�m
0��?M�zi�� 
)<X�l!�"O�T
#X%P�(-��A�
sF���'��O�usf��% �DN������'�'�=P��&,( Jwn�-S}�����2�H�nh���7x�&!0�P�O#�4�ȓ{�^�G�AjX���'�fф�'[��BS���ZLz���E�"?"��k�p�0��Ãk咰��������Z��"'�
P��bҭTg��ȓf4�B�)i��	R��+�̭�ȓQVnHS$'˩oz��%%&?�a�ȓ)UZ��7-�P�r��Ǒ9z�昄ȓy�x�G7;��I��Y��J݄ȓi��ӷÝ�W	hM�l2 �~��ȓtR>�q��9���	�$9�2�ȓH� =J��ܚR�Jm�!H',��ԄƓq~t�8���&.���1e�?��1R
�'ZM(F.��j�(
�]OȄ3	�'Iu�j��8|���L�4Z� L��'p
 �#I�A��칆���e�x� �'2�hq# S�)b�IAk�`$�r�'�~e��Z k�$IH`�2B��ab�'_z!���,[�d$�`F6	�B�j�'e^Ș�L��a�ɛ���)qQ
���'�N�����冈iaG�:g&�xp�'�����)X� n�e��'�<4 '۟sg~x�e�R!h#�'�B�Sjӥ��%!��D<�)�y6��Q@�Q� 2��@�y��\�H'tpڅ�Ez��x3�
�y�B^�8�
т�s���Q���y��S>,�F���bn(�쀠��%�yB���eS2͊򉈢_�F��B'0�yB��@$�$$J�T�4 �c��yB��8��|(��>BzHRP'�y2m&E� a�a��
8�mD(�y�#ư=�,�ҕ�� Қ,
�@�yB��d�H��A(�u^��Ud�>�y����Ej��Ć��a������	��y��N�BIabY�S8u����y2(�z��a8"E%8�V�Ѵ�����>�K��8��D^7V9Y�Ę�z%�q�AJ2D�D1��# �1�	�ɖ���/T�HS�'�(^R=��
�7�$pYs"OLH�@l�4k	z��`�_�*�ZēB"O
�UNN����B��)�,���y2DW�Jv����i� 1�6A���B�yH?%�h�j�m�7�J@�Ҋ�5�y"��
��T��/���r%l]%�y�M�$�p��1C
;����#��U�<qb�O<r��E��x"��K�G~�<i�cF� ϼl��ڗeԔ��	�{�<�E����S,	s.�����m�<�$Z�t *�xƉTrȈ@8YA�<YT�-i��i�>Wn�P�Bg�<�U�� ����gΊl���X�<	eՔNT�;���yY|	�&�SR�<١�At@�@"R*�v$�U$Ms�<� ��RI�5#q({�6ء$�v�<� ���RjS��L4;��C'a�%��"O���&�|j�5���[���E"O x��kNnUf���c׭>>ޡ�P�mӐ%�<��t����|�!qR�ͫ3f�Eړp`!���Fm �Xd��C�f�3�)DF���/�����X<L��)㇪ :,�l3%�**C�z�	K�#�杈S\������HS0�)4�Ók�$X�!�&?A���.�p�ɷ��{vHa�^?U�xB��0T'Dd�4oQ3~�.��0���.˘B��M�z�#b�Ѥz��5�$K?\�<B�	�Tv��r⊖{���D57��C�	}6Ri9��d�LȓTL�/T�XB��mAR��d��
i�K�%@RB�!��a�J�r��]I��ʼxjC�IA B�[�'ڣ? ��@caǗDtB�I�6��Q�rHW�a�P]"��;N5jB�I}g���''X<�6!�V�B�e=*B�I=	��h��m�tF> �r߁[��B�!b�*	Rg��+6zIa_�\e�B�	�+t&�kW%�cl�r���5O�nB�I6�z�ࠅ��(T����%a="C��5� ��i��F�r�+)BB�I-QB�t�s而
s��z��9�B���n�!�R��U2�ߜ8��B�IrѬ�0v� ?��s�*�
(��B�J�L�q��á��Hp�Z��B��vi�E:k�$D+7h^�b/�B䉓"��h�4+��4'��B�J�B�I�3��	��ņE����*U!�B�9h���8�H|�T1@�Ŝ,�fB�I$C�v�cgC�K�ꡢ����<|B�ɾ?�8�����p�De���&B�	(O�Ԭ� �TGP,@��ݎg�C�ɝM�Y�F^�k�X ����"}��C䉱JX��F�8-��J�.��i�C�	7g3������2򽒣""{�B䉄d��i��IE�ڝJ�"A�*{�C��8{~��+�傍C��}8dO�<3LC�	B��QX���a���[20C��F�R���+_���T�G�I5�B䉩Z�Z)��H��vN���t�	�3jB�	�X��(��J��M#�t{�I22TB�	4l\�CHvӺDb�+�t�ȓ}�,ѡ��Be�95duxS�OU�<1P��4�n@jFM�,7���FPL�<Y�M�C'��w�^.`����˞�<�f��	HjS�R��xj �~�<� V3|1v<�D�T �$)�-Vt�<9-�I�v�1�O�g��ms1�s�<!v��?l|d��k�9j�H����S�<���9>Ƕ����5� �a�N�P�<V�:Q�U.;���uN+�~B�ɲp�`51�·���	r�؊ xB䉘]>z�v�^	�~a	��<ZB�	�:���t�-`���偏:	�B�	" �.��T�X ��H�o��D�B�ɗG�@�Yp P�OO����� iB��w�`��6J�!-(��S��(��B�	=C���#a�0��0�i�2E�B�	�h����$�7[nH�"J����C䉆LP��KІ�>*�rUQ�$1��ȓ�.9)T�	�#�`<�&��i���ȓ!<r5b�Z?#+�8HE�?v�t���bQ�zbCI�>@�&�� Z(�L��S�? ~�kp��,q�]�w��6zl�"O�a�l��!m���f �uZ�IQ"OVM��oՕr[�%���3S�=q�"ǑV�����t"�z��%"O�48��!LaQ�!$��d�F"Oh�B��\�:@��į�QE��!"O�F�$;"J�+a�"O>�1EG5d)5�]%ުQS�"O�9:UAǱ\M�$@��S���"O�\�����n�a�M#����"O��G���`p��] 10E�b"Ox}�7�+<�p(�l� bR�KF"O|��d�E"Ⰲ#�-V0Є��"OX,��26���V�'����"O`�:���Ge��1�F1y�3�!��^8��Z�铯:���j4��0n!���|���b�Z�"�VA;�/[�/h!�D�M��� e�J�o��)�T�	n!�A$е�Â�),�p!"��[� �!���B�|�-	��.m��LV�v�!��"޶�U\�5����d�B K�!�D'Z��fEZ�њ`	ꁀT,!��	%�  �"B>hʀ�5��!�!���
L���=;'J�e'� 8U!�,��i��	�g#�|b�F�,R%!�$Ìj�4��Azv@�q`�K>X!�$���,�R�ƓSdf`)t�V�l`!�$���Ĭ3�l�1CG�q���5/\!�ď�4�yZ��a;��KrB�N�!�D֧3��0��Lj2��(��
3^{!򤟲y�P+�Mr+t!	���MC!�$�H
 �PnL�Š���)�!��Dg���h���#k�h�V+ڊ	S!��#<����7|�.��&��!��L?q����R(��q�����)�!�$@V��)v�V�zu`p-��mk!�d<Lͨ�AҎ�m�>@��)�f!�d�@r��a��5yA�ɱJۡ!S!�� nЄ;#�Y�z%��Q./!�d_��v��1,	�����$f�s(!���8r��x�����D�"!�ҷ-a�Ib1j]�lZ�ɰ,>^!�d�F�4�H�cA�D�^��5K[�z�!���0t�3���=�m�J�
V�!��d��;рQSPd�z�
'3"!�dԨnyE��*
�NA�zd,�67!�dр2�� F��09����z?!� Fp
0&�ԼAȽ�C�ʁJ?!��,���K��U�A���C��4HE!�
}f�]b���
������4:!�DÈlj���J{a���VwZQ"OL�C��,|��0Kr,�b�.���"O��FhJ�]�
P�L�R"O�Y"$f�*_�I�,ĂDx (˦"O���W���D�Z���xo�0��"O�X��fL�:̹QcILD����"O��j��%�J��󈂚��]A7"O���t�ݨyvl(@6����� ��"O P�؜d�.���]��p؀"OdE{DDBŤHSe!�/�Ҕz�"Op��H�n��H���	�^��C"O�݃`lM�@�Б�C3En�A��"O�ҖAJ0-|WH�L_�EI""OJp�Q΃���	��Z!bV�M�B"O� (L�3hQ�!PJ������yM���"O��A  �u� �!a�ߦ	�n��V"O6���Ҟ�N@��Gk����"O��b�
�ga����C:=��S�"O��hP���pH���{��S�"O�����3V؅�`�Ww�P��"Or��F�kP$
�'��Lն7+!��'�b1�JJ�fq80��KH)`�!�D���u�D���<2���6�P/R�!�$��!$��g�� öI۲�Ĭk�!�Ğ6y��� �ȃ�>���CB�o!��[|��a��)tH"��r�ֵJ!�Y�BOH��+�B&�h��ҩ`�!��¿<?LYʱ��V�!���D�0�!��\4
�$d����1*����D�I��!��V8���Lu.A���\�p�!�d�#iv<9G��8Z �3�ڄn�!��C�.��јVnկ��4�˕�2�!��55ǐ%.5�Љ�7I�Z��1K
�'��0��g�,�('�$f�H�	�'�Q���\�J�_T����'�zi��Ĩ���ڗ_yD���'�t�	�5	(����!6h��
�'뤥�s�=.r�|b4�Q	��qH
�'纀p��-/*|�Qug��	�<�	�'��Q*S�]�XpMs���˘��'���[#��;o�T�s�G�F[����'�.�aWb5`�ha�2I�Ѳ���' z�a(ѯ{�R���[�z ��[�'7�`2���H[BA3aE���8M��' ���7:b^��UR��'��z�bI�
���OD�=P�<��'�(�;aPW�t�'�Ă���'� t�eǎ,��s"� �z���'d(�
W�Vch68�3�ѮB�T=��':8`� �2t<��TB_6礀1�':�Ļg^�� A9'i:�����':.`rr��!�� h�OW0�65��'Ц9�a��=0�Ѫ�� �����'3fppq#�#<iXU� Sf�|ܐ
�'S�¦�8��Ԩ�O/��j�'�X4"� ^�<�s�_(�2�x�'\�5�P"�b�������8�'9ƕ�1�P-':��I��1��'�@���X6[z��7d"on!��'�b8�(�%�hf��~�D�a�'��lX��� ��$:eH�#�}��' p���cX-;t��J���$O��']��(��֔?z��0JҦ! 0h�'�v��aY�.;�Uٷh�A����'Ȏ}�$	�.f�6A�6��`di�'� %�7�Q�#�%�%�ÅV� �'�Ri9��$R0��t$�=a�0��'��A��`X-^������
p��Ms�'���.2�!�ClP�`�'�})d�6h6���-��iŶ�"�'N��S����>Ju�'O�#_`,	��'��Q`�30``��3*�va��'�ڱa��2v�Ve�DÞ.T`��'3 =�4%ҸH���Bd��' �>1��'Eb�IE�L�B�A��ʚ�G�:�S�'>� �w�"p?(��@�L5=�&	��'���a�d��gvJeP��?g�L���'?�I����XM�����u���� ʡ��/�5F�zY��N����`D"O`�1BE2K{�m�AQ���"O�C�Ǖ�$�L@��=-&���"O�A�DU2N��B��L&� 8�"O�t{$��e�t�들�03�ؼSE"ONyP�@�x8�g��!lu��"O 1�#��q�ި"�e`n&��U"O��@T<����޼Lc8�I�"OYw�Kq� ���Ȁ�m�8�S"O�=h�Ĕ�[�X�2b�V�:D�"O�����'$��B#��|4]I�"OXaqC�69�2�:BΘ�q����"OR�s�NP�8X𩙔���E@D"Oh�kԥ͗Դ�P��Ms�p��"O�y:�0|k.h{��I�^ꎜ�"O�aUgA����� '�z�.P�q"O4�i0��e��"��!]� ��6"O��C�HW�������f�"O"�	�n�o�|�a�{Ebm`�"OT4�����`S��Ե�S"Oġ�A)�����N��B���@U"OXI��'/�Z�bE���s8n��D"O,h�'!�@BCG��	bR"O��Zei�
x�� ���L�pBc"O
-��)�/(>ʼʖ�R�n�4�е"OH�8�j�<]�p"�gI�5�8�P"O&X �ܘF����ť�75Y��P�"O�8�F�f`Xa9�A;	M��Ӕ"OȰ�4��[~pJD#I�PC�"O$lp�@u�P`��\!�18'"OD��"l��Eu��@#��i�zͻ�"O�� �._�Q@�'�(:�f8��"OT�[P�/�.����U;�)��"O�͓�Ň�#��!��E$[/�	T"O��;�G�'hS ��2Α%Z�#�"O�]�  ��6�\�8��3\]�a"O0X����dgĠ��ۜM����"O܉*�'W�g��\����C�*�R@"Ot�"�D�#0��E������2�'8�M�t�֗G2L���ۧX����'��9b�� �#M,�E
�<Q�9��'�t�f�T�q���qk��H�L�
�'^�)��;�^PApb˵?)��*
�'���T�Đ5��p#G.�7���X
�'�b�;��ބL��P�eM�cGf���'���6���H9���$�M�V�� �'Dj\0�ݶ�p����EV�0�'
��UB%����C��88zbų�'��k���X�K		�`L��'0�QA�φFǖ��+��:�'���2A/U&�4xBIָwH��'�p���ľư�	Ҍ_ N�謪
�'��8�،(� h�G8N��5��'tb!� j�NZ����xb�-r�'��9�B��F}����딐&t����'���ʤO*x*��t�� .P�'{��"(Y�j#"a1�d��L��`��'�f͸6�Q���QD��q��'�H�����
	pQj�9F&V��'�)��P.td�P�F�Cج, �'��c�ٟL�\��Ȏ5����'6(�R�,���]SFn 5d+�D�'��4�L�7^���EJ�������'��t�]!
��X��8G�1J��� \:�ͦL��ACAO+V�I�"Oj�p���8�� �-M� +�"O���V�� ��0�c�1b�����"OU8 ���\@ڕ�g��W��%�"Ofћ��?�n���iO
�M��"O����óY��c7�q���2"OBL8e�ހ���:�dٛczإW"Oh�ʢD�1}*����k�eF"O8	@F>v�P���≣7Z�2�"Oĉ3B�Z��̉DP<_G�	�"O�Xj6�γ�Ba�VNk*F��"O޵[��^"G\���d�ǮTY��'R��� N�'��+7d�*!�X�@��6D���*
%B�,�[⭛�o䵉�� D�T@̑,&O*x���/:��q ��4D��/}Lb<��!�;]7��*�����!�S�n�!R�[�`F4�RD��+�!��<��h�a� ̶�����67T!��X���)�&��!�+S,>�!���3PgT�p�_�_
�x�E^��!�~�¨Q��"d�j��'e�:�!�D��Y@f䃵��
|>p#�L�n0!�ZU4Z��2$g]0E9�eG�/$!���/4���Z�̊OM�u U�$�!�DX=4R9x��<��� �Y�C�!���X��1,�8'�LZ0'Ϯ<�!���4c��!���&c!��Q��KD�!�č��������M"n�3#�� �!�Ф~� � ��4J{Ir���%S!��	q�VF�<,z��x�σJ!�^VX���?p^�-c5�X�}/!�Dj�Rx�􋟗"�x��� l !���$ �X��GR�w�\�w'�0Mg!�B"�6��b�C+3c��vF	�W�!��!!n��T�Wč)$��!��(+Y�u��+$C��Qq디�!�� 	c��@V��(�YHT�=�!��F�{���#+ڱ�� ��!��H
16JlyCDłdk� ��)�>�!��B�-R"��f���D闅v�!�X";��	r*
hk�5a�3t�!�d�qbR�ʓ�ƿS��z&���A�!�$��SI�$APM�
xl$
G ;w�!���o���+��(\�<��m#b6!��4�y	q��>�H��T��>!�^+�^A�`�_ �p��p� -!�N�.�Tw�[chy����F!��S�H�1 e��X�ܰc(ź+�I]��(�&�+Y�e��AbSI�m\|�"Ot@@sF�fH�]Ca�K�:%�c"O���#d�4I@l�����#���+p"O
���ꁹJ��DҒ�Q�3g�m�f"O�) � ̋U�X������QP�"OfL���5)�بF!	y�!1�"O
����XE��X���ߠ-��"O �[�R0��ZF	��G+��"O����+�WR��b���+q>-B�"O� �@��fҸ���FL�O_���g"O�ԪC{@̔a�d�w5(m��"O�=(�ΚH�B�Z�$=##̴�D"Ofqq7�_M ���]K���:�"O9�pi��*f4Ⱨ5l��� �"O�d`ã�!&� ���!C��e��"O|l�dO_�ril�����5|���a"O� �1��M+l=k���+8�<[2"OHx��i�8�����(q@��"O��zG�N��N���ID�T̘�"O���ҋ{�ġ(��ܦH���7"O�Uۑ�L�c2���@	¨.��(�@"O��C�L�R�d�#�B;��<�"OH]�f��+[��P��Nؖt��"O�(���B5k��LY��������"O�qAGMқ-�]2��U&s���s*Ov�{F��h�zݨ���_Җ�Y
�'�:�͜8�(<!lRU3\I1
���d7W��d��ME7Z$�A'JÄQ"!�D �G 9v M�7P��� �؆	t!�ć I��)��P����i���!�d3��D�F舖 ��%㧉P�!�!�J�����u�C�B��+pOZ$�!��&30��RtOH��d����!�DK�U0 ���/�|8�Jњ��}B��/}G����_�r�H���!�$Q�k����g̷K3"�bbI&j�!�DђBU�H��c�:����!B�!�F�.�%z�KE�~.P�ǻR�!�F��iie#�Wc��s�ʕe,!�O�Y=h)���A�3aʭhP�Ģ1m!�dU�����#@�c��hP�
�w�!��҄	�"� �	�4/��O��=���٥�D<�iy�*W�L�� �P"OJ-8�������Z�J�������"O�(�e� ��@iߤ���"O�-h�BGC��E	 n�'��9A�"O��cd���5�lZ�B>\�F"O�I�u��Iڄ�R��Q$�rG"O��Zc�P
X��(� J+{օ+�"On�§���&aH�!ц�-�(�W"O�Q*�(ȊVxx�t+�?�d4��"Od�7B���'��)o$h�"O�9e%W�=xTQ����hh�i;C"O�U�f�/+ɖ5��U�P]�-��"Ob8��-Ñ1���CcX?PR.�KF"OP�A�a�.G�u�6�
iY�1
6"Ofy�4D�93ICpƖH(4��"O�iYn_�KԪ��C��);8���"Oz�IFڎ	2��1��]�{�T�P"O��pVHZ[����^����s"O�K��صE"N�i��_�^��@�"O|���~w�p��ޮ\�ձ�"O20���H��$�p�i�3$ժ��U"O$��E邖GD޼�q����x��"O&h���ۖy��iP[�<�d�y���m��1%G�|� ��NN�y�
���5��M"$��4�����y�㚊�ȉF�T}��#J��y�M�F;\C,��H��M3ӊF!�yR��=��pAa!�;E�ike,X��y�?7?�d�#+�9Ҽ��uō�y�NϒI,p����.@l��N���y2Y7e��-9soSm�>@ ��yR%���F���C�%c�����n��y�h���vL�ԥ\_h>�k��V0�y�Q.M���I�h'O�媄�Y;�yB@�2x&�Xb�e!�*�-;�N�a�'1J�ءK�H����
�3d�A��'����ԉ�1^`�$��/�P��'���Y�-\�:�-c�B5%	Υ���� �`$��-���&�+tհD��"O)�ҏ�(5J��eĉ5ѴU�"O�yk�Ʉ4�*3p���`(A"OP +�@�^�D�AF6N���X�d2LO�	�l��@�8(qB�U�V�\i�"O���ŭ��@���!����S"O*h��Jw ���w��$6�D�"O��dD6C�������u��Lc"OT$x�g�0G���AJ�>��dR"O�D`���2%��RFiS���9f"O.����<x��@��DV���"OЈ��_�'s���%,VI"w"O�9����5T������&8��С"OV��>i��)V㝚m���q""O��!\�VH(��*��(�!"O��V��D�"�2t�\:���c"O�q;��޲m���Ca�H�%FE�D"O�єH�:���KgA���1ۑ�II�O�ܕ�TD8:��RH�{��h �'�$p�V�X�4� ��ӊڅ	�6�a�'�$DYg�J1b��#Z~~�]��'�ְ�w�_6E��� ���w��l@�'��y��%m�j�F�inN�P	�'��dqp��={Fx�ڀZ�,�`i	�'�Թ�a ��H.��ceß+�JU;	�T� ��'��iH�
�<	�b)��U1=�ɢ�'J�8��)_/��Q ��@'�����'��hţE"kx��'F�2V��r�'S��q�L�9�т�h҂˜�@�'�p������eY�
�*5�2���'��9�TI0=����	 	4���'�F�S�_P�B�Y���9	�u���r�<C��Ы4��L��j=2r���ȓ/>�8yg�ؖr��0ׯ؍G��لȓs�M��ڔV�8,�g�U��`�ȓA�����	8=U�y�W螞+\f��ȓB�8M
(Dђa�"�$4Z؅ȓ7sD��&!���������K�����	�����O/y������R�F��ȓ�����L�&����PN�1����-�r��ӡ/t�D8�a�7��q��J��}��釁Q�����L��j۴\�ȓ��y�@��R�L22�/X��d�ȓ ָ��V蝔p'��"gݩ)��݅ȓf4���3
�3Oޙ�VkB�`~�Q�ȓiJL���. 9��R��2�j��� �����M5V�*&�F9�e�ȓ
d.��t"��1��	��
��ȓ!F��p��H�\d��cI�w�j���}l��SFL	���+��V�KrL܇�>���vf�56Ԣ|��I������U"�����),-�s2$z���ȓk�ܭ�T�)txD��d�	8q�l��Lg́U�J-�S���d1�ȓt�0!�@�(pՎD����VẌ́ȓE}V�ۅ�B�s��%һz�����P�#���=g��q�l�8,K�L��C(|0���;]��iEn�3��0��{uJ��H	!s�t�b�0"�M�ȓ���h%�5�)�э�~Bp��ȓ#4x�G�G����'���� ����`Ÿ#�v4��P�j@<�ȓ&H�Z%
q3���؁X|�$���i�� �n��e�ϗz�Շ�S�? �5+�Y�f3.a��&0Zsx���"O*%QW.��JL;�B�;eN��"O�e�&l��ă�rP��s"OЬ��l^T�F]'T�D��"O�����i"��R$�%(�h�"t"O��R�.ؼCڀBe)�VB�3�"O�� �Վw�ԭ(wF]���h4"Or��I~3�i�v怮X�4()�"O|�!�f�X�|�/U��U�%Ξ�y�MZg�(���PM@��I��y���	���b�+���ԡ5F���?�'	Z)p�JOj؉�EP���	�'4�݋F@H�I�fP�0���I�X ��'���9��fJVQi%�M3:�J(A�'HyA#�3�����CB/�,���'��(y��,�U�4S�Nn���'�n �qᏺT�A��e�*@��+�'�ܵ� ��;�S�l�$I��'������cq�@�`�9j�h��'S��ڴ�E1r�t�!�	��lPE���'�$	��ꩀe�7l���'!��� ��2�Є�N�N���
�'�h�a�A7s�r�#�hU-8r����'�t�E�3O��)B3�;X�u�"O����9w�	��D� ZG��	"OʝY�ՙЅ�V
^#u?�t�"OT!:E�C=T�!XQ��q���c"O��0�˼w�Z���.d�~��"Ox�귭�/���R�	�P��%�A"O��c���#,FPs�G5g�&�Å"O�M�v�@/S��A�E�"O͓2�xy��[�k?/T(+�"OZA��4���
�@�:JdD�K�"OPȹ�

Z����ga�,n3�J�Of�9���F @�A/<�� D�PZ���]�DY@��u��R�k3D�40�s[��Ǘ�7��)`�D3D�����4(��#עF��)p��.D��!��Vԑ��Ӷ`�=��+D���W#ηZ�*Ȉ�D�
c~�����=����$		��%;0(�7��D±K	��!�C�ar�dj���x�b��.'�!��T� �Wꗰf��Ȫ�����!��0C<�cЧ�'��	����`��}����ǐs���%jI1Z����7�0D�T0��ͤ?-丸0��>LƁ"!�.�O��<�d��Fb�-~%x�@V Z�K��ąȓ�䳲mE.= �����D�ȓs�0Q��CQ�`erq%ƺ1���]��4��b�
b��jr/3p�ܝ�ȓ7ш���l�h�Rā���,V�ȓT����E�չG^�p�M�1,i�4�'�a~rLJ%~\��G)��)4hD�ƉG��y��[����Cc	�c�uYei҉�ybC_=E� 	�d�(nX��,Q �y�.e�-��
����*���5�y�@KR�F��`9�`������yB
"OՀ���6):q��!��yB.Y4T�ᆥ�<'6������y�Jϓ�3Nb`ee�&I	2���"O6�ӗ-���θ$RLpp7&V]�!�d�i����rm�*#N$�EW�d�!���f鈔뗢@�t�I�E��
^�!�ί#|���/t@8⣋�K�!�� �5�ף��d� ��B&�LKc"O����1�*���$q�,u��"O؁5N�7n໗I��L��"O�m�Fe^�0$����q�R�1���5LO�PHN��{�*#'�M�E��"O�H00%�$��I�6e�6~��a"O���Kq�¹S�H�0s��c�"O:Q�-�s�.�bC[0S�4"O�,s媇�2<Ys"�y��qz""O�a��g�R���Z�B�*R�ԅ�"O�m�ӢN43�TTx�L�x@�u"O:L�w�'j�I�bX�a�9ـ"O�[�
����qdA.��%yB"OJ�)Dϒ�c9X��
��"O���dƺ|�y��P�3�bIQ�"OBy�ߋ��� @L�ղQ1"O�𒳮�w-�������hA�"O��1�ԩM��81�@�p�5"Ovlg�юP���Z�/ͮh��1�%"Ol���+?� �xGN�7xpX@�"O���@�J��c�mW�9u��s�"O0A�W�U09U�E�ď�^�Yz��'��?O0=ӆU#D���.�  "�E*a�'	�	�`4NYydX�y,�Փ`�,a��m�ȓL#��цn¸��)s����Ѕȓid>$�Ø�?�>�R�%2T��,E{��'���'eԢ+������^�"�)�'4u���Bm8@ʖ�c
���'��
҂�Q׈P��@W�*����hO?��l^�*Ԩ��Lݬ;��P2�(
B�<1���
vF��uJ��|)�@�Q~���ΓE焨���-���uF��D�����S��!�ۼC|][�>����(I���<T�4;�� �Y�ȓX蒌"A[���`�[eR\�ȓa����ĤiȌ��l׉$�����^�]�B�D�=�$�ꎋn����ȓR�Nٰ�eكMXՉ���8��'ў�|�aOhx�"ҬȖb�$���,�_�<1f���D�&Q�a�C/��p$f`�<q�HD�#׈�ڢ�w��ݰ�́s�<Q���	J��4��m�z�p��O�U�<�1iP�H�
��*.���V�<�aLSo~~Aa�Dn̚�I��NԟD��[����ɻ+��lPp��p�@�ȓ
�xl(E��"�8tz�/�~C�8�ȓA2�3ƠC]�v�#@"�kKXȄȓTjx�`r
&X��seJ>�&1�����q��	�$�→�@Q���:d~XXP�ˬr�W�(Ժ��1D�`���c���,�L��#D���dS�'4���-��c�����!��O���4O�0��gAy�� ��
��Q�"O�h{�&X+JÜ����4�^���"O���!��}����	G��d"O�4���k��ث�"���s�"O�y�D��\��!��k۲i6֥�f�'p�'/�)�'2���j�L�&o��6��*/ZU0	�'���9���lE��#�jѸ^nYو���O4"~��U�`b�;ХL�c&P�(%OQN�<���
(M
��5C '�}��fJ�<ip���|��Ȳ�F]��U��M�}�<a�'��^���*���UU���1�ZD�<�� F�&} ����rw�����v��hO�|�� �W����㓠� ZP���� �S����]vb-i�� ����]�D�!�DMr����g�6��1HWI�%|!�DW�\,����W��p�i��'i!�Z?�|H��U�"�{�"L�h�!�DV�S�M�p�¡^]�Ca��K�!�D
�"�p��$����T �ў��'��y~�l�4P�fؐ��W�~<j[�.F��y`��hሹ���J�cNP!e�"�hO���)��A6B<�HN2d�$s�IK�N��g������U�uut`HS��..imB�J'D�����@�.$0� (�!B�0@�&D�(�G/	?�L�Q�.���ء��#D�,z���-F�\P��)�IZ�mʓ!�O��>ڙdb�)l��l� ��6�h��YM�L�B˘Lc�ˍ
f���ȓ`$đ��D*6+�݊��/���'�a~r"X� n�)st��f���1P��y��6^��Q�sc�0/�d�h���y���2��c�I��'��-�&
���y�A�=��qzpk� �0E�v��6��>��O��!ECTc�p����]�EӐ"O��y��G�/`�d����.�M��"O> ���ٱi	�pF��G*N���"O��at��+�����s>(��"O�"��CU�,��l%y�b�U�<�iL���8�����u}�𓵣ON�<	��=�|!�BV*6�XtH�J�'a�4�J�f��:@iԸF��\�����yb�3l�Q��"89��9Y��Y��y"�H80^�m��E1��f��=��)�O>�أbCY*ѓ�Ř� �n�Xc"OJX:�F�2_��=PB��
8�����"O*�1 ��+W�����@����!"O d[C�M<%�,�1,�`s杲�"O$�`%��X�⠊+�d�(�ɗ"O*8h���rh�1H�V��ꕋל|��D%§-�lQBsg��U��5�F`
8J6a�'B�	S���IAM�N�8b�L&""& k��0D�8!��
pp|����͒��q��l0D��x@~0�0�Ɍ&Q�5!�!-D��Ã�-�L�fn���&����/D��hE��@eSb.��K�<|��,D��##��>V�t�u��/^��f"*D��	ЅU12�BF�W��t��b(D�\Y$�݉,�z,����$�\R��&D��@�	G.>F�=@���
q�	/.B䉸J�V �Ҋ�@F�A9��Z��B�	v���*F�["68i6MK#4{����&?!��N�!�Lt�m��t��H��
v����D%ړ�����*����W�@�Mm`�����ğ��P�!,� ���h�\�!�C�}`��t�� j�P��\�X�!�٥
�$�"�hQ
kwnd*�'�0�!�0h��X���ө)jT�� 7~�!�dHF�N�͌'<e��b�!�nl�	��?E��˕�{d�c��ֿ>�2][`��)�yB`�`�q5hR�FL��q��ޗ�y��[?@��T�60qZ4��M2�y��3h�����&"&:����Q��yQ*���+q$R�cҍ���y��e>!3���8� U��y��
o�ШfD_�}�8 t�Q���D�<AO>E�T�۾;  $�W�0l6�S鑯�y
� |�)d��v���RPK�]R�P"O��ei6G���I�)\/pB�eiv"OB(
�H4d��}����2�8�j "O�{�J�4��\�fZ7.�:U""O�J�FW#f�J�E_�ZL�"OF����W+�����O2�b^�����%��|�����:قQJ�ܲ`Ϡ��So�r�<�αd��yR�)_��#�KW�<��O[�PQǭ#AAF�:U�Tm�<Y"J�T�cOOH�R���A�k�<��V��q��MR-<њ`I��<Y�
����J&�Q(O��!F�{�<9��	�Pq45�Q�(�R�ɤ�y�<��"G����B`�L�c*����z��hO�>���V�T)l�b���JE�|�����:D���0͖&�-��C�;]$��j�Zv	��mӼdAA#Z�t�ȓ2�����3G��7OA*;���H<�}�4)� ���V��vxX��ȓ7����g���|��I��Q�؆ȓQ���l�j=�FꋆZ����?a���~�&�K�In�8 pb؏&��q�Fbk�<q�F��;&IZ|�V�1��h�<9�j�u�$ܡ�&�Qޖ�D�[[�<��Ȍ4_��U8g�_:}�����V�<��ʑ)`����T�ʊb�"���K�<94��<�&�%ʞ�Bin5Ё�N�<�j��_�Hu�ч�$E�哆��J�'a��CO3�6Eѕ/�,zD=æ�ƥ�yrKXH��IB𩟛6�<;KR��y�H{��D�e뗄/.�� V5�y�׺�n�`�,�//0ݳҦ���yb�M__p��q@I':(2�����y�g�<	f�1r�hs��2A@�(�yBmA+��!�C�Z�pxPh>�yR��3qV-V���a��.�y�M ��y��$�#JI�ēg$F/�y�kW�V�b�@T�[2;k�" L���y��Z�1!��k
�1ؤ��N��y� ٣;�0����(��L����y2Z�<��l��FL�o����L��y��](%�Ӣ���<�� �9�y�/~��\3�0\�~�tM� �y�%� ҄ô��( F�e@�(�y�� �!h0�2�O%%��t�CL���y�Գg�� Ѥ,		&� �h# O��y�J�,qiH��.24\���BS��yo�>|ґxq�ŧ-�8��$�3�y�LP��ɩ3a͙"/2$�Dg<�y�A�17ό1��j�UZDO���y2j
�)�ث2�ޡ
z��V�ݏ�y"�?h ^��CoÏUg��a�H���y2�&P�DX#	y"�2c��y�Q�G��� ��+_�h�[!�Z��y��˜Y �Q�ǎ�PԆ���y����l���u��F�&I;1E�7�y�H���i���9ʨd�`�"�y�H�I������P-�>]c����y�M��?��#@�6�30���y�%]1>��ٺ��G�3��R �:�y"���B]��dD�|��)�D�ybDM�UT� V:|�la��P=�y��ƧC�2,y�
�u�<hZ����yҢ� v�͘�B�n����d%�y
� ���uX�[�����?[��Y�"O�������(��잉`���"O������<�a��^3e����"O���&��j�mSaC�����"O>���M�-�j����!]��5��"O�t����CH�����7y�v���"O���@�����G�ft��!"O��h�OHp-�%���ӿ/k|�S�"O m�ХF�}�࠲�_;��"Oj���kўEѶ���� �$���"O�dK�J�b�3A-�%$��be"O��"��fL���m�E:m:�"OT��F�Y \3����L��/��(��"O��ĥ �Oְ�H���N����4"Ox\�2Nѡ#/j]�ɓ��
� "OXC�\�<stuc6ʆ6�,Q��"O:��6%N;��C�T�ܴ��"OƄ�t���E�(���	*U���b"O��0 R4B��Mb���7"6�A3�"O6d��JU�T_(��F�LC�"O*A�P匽W�����!8�Y�E"O�\	�fV� ���1��� p"O�|�#��wh5�)�<�� a�"O�٠C�HzƲ�8��I&Hsh�#"O���u-7K���E��^(�`�"O�P4��7C��DP��6]>*uA�"O�uxT��`�2j�i����S�"O�X ���'Z�=�PI�!�pe�"O�dZA�G� 	(כ-Ѵ8��"O l�ō6�B�t��6w�zt��"O��"S ��(@���H�BT�7"O�<�"% H(���Ϛ<����s"O) �Q<�x��h]�+���#�"OڵY�J��`$�)
���$�"O� ��iX�T����V:�z �"O�āt
:}� ��F�
�a��"O���@î��q�
)5��w"Or����d����)ȫV��̰7"OVE�C�b���	V�R�"Or,�v�M����(Ob6��xb"O�4R�� � ����r�@�S"O֩�V*�N�J��7���g,�P�"O���7��_��yC ΁�m2�P"O�ڵ-��伻�Q&�@�"O���Z�o[�O�fbL�"OLK��,1R�A=VI�Y&"O�H�욈A&����C� B���"O�	c���?�Xpy��Ƌo���"O���e��ʝ��`�L4]�"OR|�p��,Jf",S��yښ�
G"O�pH��'��@�#�G�Ò!��"OxQ��[%Le�V"̔?��}K�"OR蹶蓖2;&�h����ܳ"O�@"����6� |r�aO�<�&ah$"O���W��;���J���e�
�!��]%I��[dNҨA0�%�(X!��,x{���l4TțF�=c�!�d�B�{�c��N8ۆ�A�c�!�dG^V)���X"U�\BWcS&f�!��S�;���0&���M��� I�!���8V�CҤ�.���R��14m!�d#U�&��� ��~�� �I�VM!�DS�G}2YI�a�]v��FLU�S/!��ԍ-_0���kH =��*�ۥp�!�� @���dE�Nj��q�◶J�pC�"O�u�Ȓ�D��cAʞ����"O���w.��Dj�L�T��s��Æ"O�����T�B�DS� Az�"O��	��$D �m�"jH5�!��"Ȏ�!�E�,-�P$�R�㺄2a"Of��wb$���׋�t��"O0���͒Co�p� ��*�^��"O�	��C��Bx�Qɴ�r�J"O^ݡ�F�@`v���՞e��)R"O�m��d�5G����� .�x��0"Oډ��*4�Z�%N�%��Y!�"O�H��#��dh�4��$�	��H�"O^p�M�|��j�A�]4h�"O�} �L;G:fݲ���+n$I�"O�U�A�>�	�B�F�c�Q�"O���^��)��`�M�Na�"Oʐ
�
�b��5�����(R"O�%Rw���y�\ih��O��]�"Or1�I��,{vEڔV�& ��"O,���^����<%h݋�"OnQ���)�>|����P;|�a$"O��b��E=p!���c��>pQ��"O��h4�ɲB)|�Y⍃�4T|�Ã"O`E�u��)X��eLQm'��{"OhX�,�r�����ߍ�nZt"OBM
�Lȴ�)�'ɒ3���#�"O���r���k�)P���E�N��D"O���
�7���d��-e���"O������s��Y�j�SF���"O�кq�M��V�ŏ6=�}����yP���TC�4��B��y$֓n��P�L]�$����&.���y��߲/����s�< Fq�栌��y���4`�8����
Xaq)���y���i]-�F�X?��Y����yR�A+;��"7�����i@��y�.кXv�C �N#��DJe��yb��%q��
%"��	�����yb�ސv
�U"��c�IP1�@ �y2ᙀ�v��M�]q�E!���yB
k�4��� (�홗��y2	ݖ
�(lX��6f1x�+�!�y�d�Y�(��o�-#��z7k ��y�G3�l�
�*,<�&%lO_2�yR@T^��{���'j�q�+Օ�y�b�%v�;���B�M+�yҠ_�8k��{�����@���y�d�YX����
�,��R���y2h�Fp�( s(�/���
��yb�A>��@�K K)��1$��?�y2ʔ�R6d3c	�IV�%�Z1�yB�?`xX���9J8�)�я_��y�]Ud���Q�F���ځL��y2��'��T	��ʐ'z��i@�՗�Py"A�R����@Όn{�8��@t�<y���>����#�J�<�I��ʟK�<1b��9?���z@$�008�qy��Mb�<��^!^��iK�J&<qtcT�<9��3BΎ�8�j�%n�؀+�`�u�<�c�
'Ғ� C-^�_���I2�Fo�<�mK�r�� ��9�~yQ��C�<)��7.\$���PT@@�%KAB�<1$Lj>�h�΍�\�\]p�.�u�<� d�ڦ�	W��,!N�GkR��"O���d�!H]��O �0M���"OLl(v���b�ĉ���3�"O2i�������gC�gV��"O�t�g��)Y�X�k#�l�.<JW"O��q0#M�A�$���GG�,��H��"O�9��-?��|�&��)7` Q�"O��u�J�"ě��# 3,-�"OԽ��YT��q�����7+Ό� "O����Ȏ�c X�AR�N:q<��ٷ"O0H��d��I|́��>"Nn9�r"O2�Q��[:!i��U=i.�	!�"ON����+�L���\���Ѕ"O*���X%���*���F���0"O=��l^�X�A �A��H�� �"O��r���#2���'�d䒀�A"OZip�Ə\T|��E��>@��s4"Ot���A�z��	��°ư�)u"OH ibݧer���V�ŋL���"O qp���/gt$�Dō(<��"O��c&G����1�X�T	jlئ"ON�z ��D< t� �
��R�"O0с�!{˨��� �	�~���"O�l�p�Ӽ}JXS�@�1�Y�"OZ]S1���6��4"/��b1"O�` �*�F�LkV��:�`�@�"O�a(�/�7��̒ܳ��H�"O��CHG�lt�#���"���H�"OФ��웑IO$�c�*�����"OR�	�
�g���9�
�)t��!�C"O�2� Jexڀ�c�Hc��y��"OBqz��ƄAC���Q��/���"O ���@
�uB���_��h(S�"O� ��P�K���`��h��4"O�$gB1��i���` �<��"O� ӌ���Ɇ�M>|�Z`se"O*���K�e$\���NE
E�p�y0"OZ;��H%UxMڵу:АXc�"O�-jՌ�%G�P ��@8<�8���"O\��1ϑaYM�@.X�R�H"Ot��g���Hyx�x���1>*��R"O�e�D�b�LM*m\�-��[��'q�'KdYh��W����R�(�*"�(�j�'8�0�1�Ζ'�4�z��fDBM��� �S�$��r��a���f�F�x�l�yR���Y����	^�Ơ��Ƣ=E���x�{��E)w���8�ZV)��g-ؽ����D|Y83� :w����?	�!�O?:�(��ʿs@�գ��s؞�l�_�ɒI�D���d�<qg���[���C�D��� ��<���兘�P�HC�8Y�N���>_�`�w�B�1gH�1����R��U�6T��B�I�l�4���
�B!"��2��	�fB�I�iP�03�&̈?A�C�"�8P$B�	/#�dQ96��|!�u��&+� B� <^<�̑�EP���.��C�I
+6�����\�D��a�;6��C䉤ue�d�,
A�l� �d�� ��B�	bM�
�����#e��dtB�	nb�[��C�4��,����~B�ɜ��h1&�2�8��G9(�:C�	���݂�D��<�Z��U7�B�I�h6�� �3&�1z�|��B�)� tEy�* �pK*hxMQdۘAkS"O<�Y���L͂�"DAg:I�"O\mS�'ɱ0U��ip��K|1�"O �A�Q�;^�ɠ�O WfT%a"O��1DHW�l�h�7���w��l93CH<�pɆ$<�(
S�J#}J���Mi�<I�%Y�����!z5�	���n�<Q0�ǔe��P-�P�Pao��FyB9O�L���iи)��\�Rj�7 �	�D!��!򄊪2x�q	�`�"�[Q��+��I�HO�>	�CM��@��׋4�P�k)D��:��	p:b��$�X�[����'D�b��
i��S��W�Q��`+e�1D����+)g V�C�c[�G���ySA/D���Ā8l��peL97nZ`��-D�\��g�_�e"w����я*D�$�"��%.�Hz���
~����,D��I���I���"T��	$ra��+D���!��%�l�D&E$����)D�p@���=븨)Q��4���
2D�8�C�H�/�L��$$�* �����,D��0���N��@�d 9`��� )�OO�aK3Đ�@�ft�p��pp����"O�`V^�P��N�?hT;"OZP�t�S�uE$�RR�>I0�\r"O�|@˚�=�d�k�PXâ"Ov�Y��)VT�k��Ԋ#��O��5��_ԄZ�ÑP(:$�b�&�|���㴔�s���]	N�K~���t~B�OV��6ǂI�*|{rܝj����w�⦙�'����<��'�.��G�	�S)�JcmH�{��ɚ�'��t�a�K52T�ۧ�4���7E%4��֋�-���j�[CS�-Ӵ�+D��X�A�`����ė�y���;1O�����'6ފA�Ȕ:`,b �Eo�-qX*�OF�I覥Fx��|Ή#)S�x��d�9K� @���ʿ��<)I�ȕ'fZ��s�D42�p�̞3t)�]*OVʓ�hO�Dnj�
����̝#��#4>Y�>�E���E����B����D5 �mp� �	�HO�܇��s�<uRi��"��1�)��d��	ӟ\��L<����#��e�Ҩ�A;� D�8	�ua�X��(X�0�Z��W�N���t�<Iߓ3$bC.ٖ)����
\L��R≽Z�^�{����rk�y��� EXB"<)ϓ=�Q���J64����T�_�isDyb�|b5I��X���+QN�*;Oa�r��y}"�'���E(��^a^P�C�g�Z�����c���q��(/j�Yb�/ٺ?F@B�	�Y_LxFM�;����eZ�w(�O���DJM������� ���͖T��`D��.ٝ),�]����8Rl���O���;�S�Oܘ��b�t%����I�ǌ5���D1,O*�)jZ/$�L8(�g!'n���|R�'��R�޺X���C�t�>�"�O�=E���	=�@(3$?�@@M7�yr̔r�\]B'�E.3i�'���D.��O�I3SI�]o�0�A<P��`V�If>��U���`Qb���c3��z��:�$%�S�'^�y�A9}AP�D��jF����/*ܪ���& x�D��*Y���J��"��*����8~a�ȓ y��]�d�b�ڲ��R�<��Ș:qh
d�V�������ȓ~^�q���Zi�BQ�c)v�h���S�? ��y���!���X�HNG�hY��"Oz1h����
�i�%P�a���qǒx��)��DB,�k��U�0yĄ�@��I��C�I�	�yrD���<J�y	��*;��C�I?ز�@�d���e�7��(��C�	�6i��  �Av�\��B�+�C�	�u48&��,�ܤ��,�f����d�<��4��Q��ߘuu��lGu�<�A⁲M�dx��k8T����u�'O�?q�N׎,�v���0�°�<D������F�.]�&���8��9D��:2��?MP&�k�@�z� L�w	+�Ov�'IR���,��A�a542H\�O%����S�)� X���&)p�Q�Tʆ �(#=	��T?��C�4�����%id���>�*O���$��egl`�I5u���ɚi�a~"bM�j��ǜ�)�R� &eąi������Р�y��8P��u�è�	lNn-� �O,�'%Q>���a!"dz��W!h�Pi���=�O���Kylq�6=��X���)MNv5D{��9OZii����C��p�`ٸC�.ӗ|�>����a{��1e�/I��"��x�	�<a	�nj<*���p`HI�p+G�7A�=�k�D QQ�N�V�2髆ꞗ8�p��
@�0�7��4Gu@P0N_�A?�iD"O,MP��ɂy�N��c�
�AZ5�@�'<������S�#.\�y�l	�"�*�+D� (� P*mZ�l���U�}���)D�P󢥄��! ��M���%D����(@�
m�ٛb�A4���$�N}"�i>�"֣��p�@ �7l�)`����#D��HU�E9`���#�*�e��H D�0`p��_��-	Y3|�@�2"O 9v+		�|#%d\�qBQ��5Oz��$;(*�$��
�' ���GUx�!򤘞��-1�#p���R��Z?bD!�䑃Z���cp��,�Z����!���M�L��%�tQ��Q�j".�!�DUdUx�7�_���t�Щ]*�!� 0J~� 󦉥F�Nh�a��M�!��OK���7�DX�I۠I	0�!�d�|��88r��@,hYT(� �!�ĝ�XwZ��e�I$+�����@�!���.3���,r���ȃ�O�!�@�2,�p7��{��T�q�
�!�3~G�䑐c��!A�F��.C�I�+M����R��A:iW��C�ID"��3,��jdMt�)�B��a�`� .6� C αk��C�ɇ.��iZa�Ù!���uP�.�C�	<	8q�N��kHܴKs�̢*R�C�ɥ:�@�J�P���Rf�I(w��B�	E���t�O"t�`A eDE�L/�B䉕1�e��C�\Z6�h�f��&��B䉮^�A5A����D��("RB�ɸ2д���(�&p�����^�]�<B�I�J�t�#�� ���i�G ��:B�ɍ Ԏ�a�E�!4��%�s bfC�I-k�*#J�7f��!y*Ʊr�PC�I�k�����-�_��Y���A-=�C�I�%s�̰�l��4F$`r��@<�LC�ɓ/���aW'V�F���
�� �!<C�	�F[<���H�,p
ԮӤg�C��;b����ԀÎ/�"p�R!ҞwM.B�)� �1됬[�I�����4�jPȂ"Oz�����? ��f�6t�f��u"O����/��T��8�&6J�cs"O8�)��ؑ
��H�"l��4���"OF�I�bW��Z���KI�$d��B"O�;�CC<etT���&�h���"OvX:��I�g�U�8�f"O�u*P�ǊAŲ�F0j�ɚw"O���j�)����G��k�"O$2R.���5f�7��	H�"OTt��L�Kݾ=�E"������p"Opy���G�45�a΀a{����"OY�L�*��0<P���$P�yǺ�8@�'�,y �a@)���K�%,f���	�'i�q��-@�c8 I��)%�z0Q
�'��5B]�R�0�����8��	�'I�lc�
��u���I@�B�'�0yałR�K'2D�!-8)�~I��'�� ��oY4�R8y�W� �j��'����⊤M��a�2#.��
�'�Č��hȥY�f|P�@������	�'�tjU	�U���2��p���'2����	&F|$˂�κXA�Ԙ�'����.�*�@U�V#�d���'������2ڶQ2e,4H\��'���4h��l$�PXp�6g�(��	�'�0{a̅
7a3�쟣UE ���'�Jp� ��Z�Hu���P�_�\�*�'[,�yA�Զ<�ڗ��Je��h�'���1�N�!�2@ 7�B����0�'Ř��~��x�bB�;8-n�1���O�<�4��#O�Z�q !ʳB�TS��AA�<�"�T	/��8�R�J�b���E�d�<�.ÿUD\hφ�E&f���O�\�<�4�<lxz)[��PI�x����a�<avd�x��U�@�8�ٰR�X�<yt�X�+�ʁ�v"�:qkH�Ȗ#�X�<!'�]�AŨE���ȣB!���l�<��k̀`������R�Vs m�g�<1��(P14,�F'��U.�i��#�v�<��Ž+,,���c��[�x�p��8�	5)Xu1�Sv"�hTֈ+��<�h�=o߾B�'5��� ���h�4���-�,��mz�!�������|�'iBp ��w��Z��F�C$p=��'��u@r�� ;hp�&gőf���'�����Fw8� y�" ���a�.�n�i{��>LO�x��2ָ���'(l@��c�#n�����	g�$T��'�$ɺ�g;�>��aD�S��IȎy����V��y�6�l�O@콉���=�HP�#�^�=���Z�'�Q0PB�. } �!Ղ*r6���"���O�x$�3?���L+;nD,�SJњ!�ʬ�b�~�<i�!/Nx��ʈv�$�"\�Wd�9�"�y����$T+(r�y��lN�|oq���,Raz���3�����ʖi?�a�:^�"�ʐʕ�<<u�S�D�<���٘mm����Y�g�zع7i^�g�p��G��K{��~�������̕�p�u2/LT�<��ˢ��b3'I~z��0ab�}l�<:��|r"I���$G�!\��p�
,'�Q��;%!�ܾ%��P{��?��t�M69����k����I%^�n�kS�Q3ye^���M�<C�	�k�
�a"'�2N>5���	��B�I��,�� #�	3R��xDF�6\�B�	�'5Xu��́���؃���#�B�I=��HP�����?�\�j��y
� :afL�=N2��ғ"W�?zn�p�"O�1�W�_�i�TA	"*[�]l��J1"O�a���!e��ų�$��F���"OXY�#NOhn��`hY�R�����"O:�Q���lM�§�l���r"O ip�3wג��� vf��"O�����Y�ڙ�Ƣ�-�.���"O�XRlN}�zqITa�0z����U"O|��d�J�F<
��Ӡ�4?�u�d�|ʹ>�q�=�}"�%�?P���{uA�'\����D�	R�<)�/^� ��Ơ�b�HS� �fU�Oj��OP&����E D���)+�PADF�{ m����E&H��U�Ϡp�Ci��W�*l�B�&J8X���l��=�a}�8�N��%=�	#	���O��FBЎ�t<�!��	Ir~�S��֘ �莬K\V A� ��B�ɽu�@uZ�錎�ƅbK6��Ld| W�T�\f���d�Ǩ���4�I�ڬq̃:F:
��"OY�w��>{�Fk�F"�I�#cQ�~����g��m�ΕZT�::�g��lx9�B͇	��Y�L�
aԅ�� qB0�aŗ 0>��2��e�z����B*Xfn!RCc���B�A&�'!�����!a��c��2y�(�����VT�z�LV~�}V/Z�2@�I�&55
QǪFs2Nba��_T!�̺x��;Sg�6)�pba��(rP�$K�1p
I�1�	$Jx�j�E��{��}
�T h����ě!�)���~�<9�.�R	p��4�tp��8B�������;L d�q��N�${��(�.�S
��Op,�-f��r�K3d� R�'rYt��+&�O���CX,]4t��cU�X��8�g��.�pts�BW4Fy�u�́~\���Ƿ�?i`��&_����AU�,�r��>1'���T	T����J�O�������r��x�c���g��0���F�A�'�:d��4١NG����)�;n�$b�ϺEÒ�O�L��˶ሣu��SÓ1�$*��L&:j[�;0K�9�ɠ ��!�W3�v�[���2�("�O8b���94M� YӠ� \tPQ㥮��
�2�g�;	ހ=�%��u<���C�t��ňwe�wx���$�
�,`Si�~[�-+g瘫F\,��j6s��ŸǅX�rt����D���}��
U��5����^����iX=D��{rK�U���ī�S	���4B�kaz�8�HB�l����FI�M%2�Fֈ�0�vNO=l��訔b1hgp� �؟�I�J��,4�����;����d�����ȴ`߈ih@j��t�]�,o> �%'�D��&I?x'03�� 3�byZ���v��=~+D�;O�蛇��]�B��(	�.�}�X�@�Z�Y*��wO�b��䓯�*�2��	=}�[�^>I��ja͉�o��H1��
-b��t�E�Ϊ�x�c˶>
D�Z�<��5@ݦV9�|�������� H��P�ez��K6=	D��.�>��"U��'Կ���ٺo*0�qEc�%xL���DW0��=���H�h-��j�;mI� �S�4�,jJ�O"
I��L"8ŢqAs�3r�����M�0�lZ5��g}r�C	H��8�#�]�T���ʾ��'��A�c̈́�\aQb��o���V�?����\�^��Ԃ�zq4��W��O�}��߈I-��7����<1�)_�4+��B䆐?Z��v"@?Q���-Fl����@�m&�G��'\ �S6$t�1ḼcU�� �CϺ�yR�/��:7`�M��tJF$���?���	)pب�ī-lO~Pi��٨��cU�W�Q>�K��'��� �]%>rb�@�P�	���)e�P��G���y�aےd���C�4Zd��茅�(O�P��![�e��#}����L8�R�.H�i#�
�i�<�S�X�`���x�Z(K |����T�K�\'�"~n� _���D��R">��B���B�I�]:��qc���C�
]�5���i�����%(��PazM�w��8:qkEq��8Xua��p>���Շ0�`c"�ݓ6��ܘbLs}��b����]�FB�->�~D�1	�Hy����X_;��<��/8�fl�aI9§2�6���"5�(R�Ϟ&c� q��X�8 Vl�sM��9� �? `E���Ke��9a�OX���OfI��L�W����7�r�X��E"O�!£��Y��&ꉍ��e�"�O�)���4WEb�ӓ�T��Ӯ�S��T
�l�;Ӵ���_�`d�B�:���U�I�@^A6�//p|@�s"O�y��)�L���BA��,3��2��e�ga_(�>� �C�.�t�QL�}�l!Z�F>D�� @E��a�!J�.e#��.j�4�׸iX>|�ڤm�ɧ����m�r߰���瀛/��+��K=�y�)�+ޜ%'!��PDd3R
����D�i�vH	ۓ~�T!P�5�!IЇ�E*)��J�d�Cפә*���уM�KF�`��I~�r��ǅXz�'	�j�0�ȓ8���dC�1z:�*�@�$�,Շ��ޠ���8z�,q���<r1E{��6�`�i0�DuXh��3�>ls��&ÊC䉡�$)�B��+�����Q�BZa�3*����!A�}}�!@.L�J��23E_�H�͉E�>D�aE�M[m�%Z�aZ4+d�0�z�걉0M�G�2P�ō:ay�&ܞ(�z�����lj����N��p=qc�f$���3��us����dM �x��Z�f����S-��xbl��PqKv���S�8EF�� �'��c� �;f��HHDʚ31��V����>OΑ�0���b[BEc�"OR 񢥖����qD��M���]��b����!4g�������<��
J;c:A��O�d�^-Jc��T�<�l3I�1��*JH�X��.//�\-���09=���DdM��ay�F�5	�M�!nɭWE�����5�p=I"Փkbx���(�,x��G��rm��:ABҿq�^�ru(���0?1�S%?p��gG׸Z�<�A�)Y,q�	��.��,s�Y0�ϐzqz����\�db�:��;+%�QUW��DAF}Rf(Q�T��B��6yY`[4��*\�f�閥��}rJP�W�7G�r��5Hv�@�W�<�Ec� �8�9�D��&�fm�"�I�<0*S J�BbO6}��)0kv�4�4-={�̲.â���K O�����K,Z�azr�����S"b�5X5|xᆊS��ķh�~РB���ēn�~����OjX�	�v�C�\�qty��O�%[�2����,J���SO���Vd�U�F�v��IAT*�F�
-(I<��hT�5jb8�D(��C�(�����h�h`�!E|���0~�`�cőUܧ5��:D��-h�=b��X6B�h�h��_�@�ݦO٪��Y���!(Q�%�ܭ c꛾fCRNb��p҈�	6���#��>E���Uc��hq�&� ]�5�����M�@ޖ/+Ь�o?h�)W�N�+�>`���|����'U�e�T��8�f��<�t�8�d�{�����H�R�+�1����V��%�#���$�����P)�d��@�ޙT�xZ�
O*�{V�A�A�܍�!�|�Vx��	�fA00D��x�'E�@e���x��D2�O'�@��ȓ��S�ׅ~}���6F�R"���'�*�����w�S�O�{ �8Ĭл�"t�t��'��l3!ė=�	Q%C�&�����'LD���^pH4D�)�D��'RY	�@J�W�>�Y�&M�%yb1��'d�W�=b��*�>�p�)��4D�,���L�Kh��(s	�%J:�� 2D��#'*˲P�
���ψ�D`ԙk$M0D�pҵ�H�F�d�7��gsNu�C�+D��EkT�2�(:�-�(�$�-D�<�G%��1�{Ў�0dP��閎+D�0)C$�]ݴ1H��@�?��df�"D��	�),ra,=
�j�qܨ�n#D�Hا�O�t�hQ��%_(��i��� D� �斚"duzM�8��0{��-D�0����q�4�pe�)|�f��I!�Z?*$\����N�0�%��?#!���y�F��eL�x 0xJ3Ƒ��Py�c�{V4��3�ӻ�Ą��Z��y�@K����@�-X�e�(�6�ybD�as8�0� Ӧ)�l�X5�P��y2�G*:���b�])�PȚ�o
�y�E�)�T)Q�V",�H�����y�mA�`tr�JA6#3f�3����y�G��]xQ�Wò��K��y�i�'.p�)�`زR\��Ӣh�=�y
� �)Ag� 56��V��4#\Q"O��D$J/	|������W$�""O�%��8)<�DB��X�{�"O��a*�e�DD���Y�!�d"Ot3�$U!k\A�`�#�6U�"O�-����?&I��O��s�-C�"O2$��"�����c��DN\��W"O���b��|_����_� t�ȓgb�؂B��-OX�۶����<���0� >6z�A���&of8�ȓ(�j����ٞ�iJ�L􆰅ȓF.�81�A7&NL�y���#�^0�ȓFW\�3
� )�'įt�"8�ȓ(�[�f«s�Is�Ì?|6����FYh��_,�r{WKБ?�ȓF��`�Fe Sd2��ҫӥ��1�ȓ7LL�%�j@:V�]fu�!�ȓ)�4j��ɕP��!f�S�oE��Fo�(;�JD8�]IëG:RBe�ȓm�"�����5�ƕ��MQ�r����ȓ98��"L�+qV���.���^=��q�\i���N����V"�؅ȓp�-3���E�Ryu`�\�D�ȓ{��r��5-�a� �l��݇ȓV	�-#�V�WJ:��Ca�x/���"ޖ�����R�z�+4e
�x'px�ȓkZ����&Q/��'CQ�x�`!��iBuaS��U�&y;��"o%TԆ�=΄�(Z�3$+���5I�`��Gd��ؒ%��e���1r�j���fW�3�k�);��� y�������.H��IA��ʇ :�ȓN$r��# )P�^��w�Q}Nĝ�ȓs��Œ�B�*����L'vu�ȓe�t#����$	��gB�s�Z��ȓ�=j�CX F�}�w��e(`܄ȓ!�$��&�D�X?̩@�X5��E��27&��Mq��I�BP2uB8�ȓE�rL�W�S�r�B�J�6�"u�ȓv�$��D�
�Nz�N�<����h�%�\�h1u ��Z�L��ȓb����փXG��P-F�����>�X2�ʔ�����䔍� ��y��UZv-,l�ܴ u�� n�C�	?v`X��"
J�"@��G�sg�O� sT�̥��F;�d�Q�P���OP'lE�"O�4{6�'��Js�G�%����2egt%%����<!��8m�>��GI�?����T�<�@�L?�AJ@������ِ�p��c�%V���dݟLK�ᗅ}h�� Ώ�$�az�KB?>�h@���R?��K� m����M�<��a��n�<�K�Ex8�,|��d�7j����<�W�5l�����D+�'j�|� ��!o�����J(X�0T�ȓ*9���1��%ej��5�S����b�,&��'�:�я𙟘AUf�S0��BaY' d�1�)D��J�
͍B�, �+��c�b	�V�+���8��	�r��|�*��+G�0g��3����i��0=� %��x�t ��J3hS%��0
a��'ՒXAD>D�,�$�@_`<D�Qb(g�����?�I(f����I�#I�Q?}@���6\��1�G��Dt$xqf:D��b ���FS
��U�N�D�;�aث��bL>1��8�gy�/�1W�@�ғ�R�J���)����y"!	�����R�ިL~�I�$�-�M�`=XXH��ןx������E�4 �ʞ+r�!�� BpZ�a�7i�� 7f@��ֈY�"O,T:%���rmtLpP�[�$?�AJ�"O���0`O�D���Ä�,,�(4Y�"O�� ���tX��3��tĶ�k�"O�ty�
ǬW��pSa�r���T"Ov0�w�O/�bAQ$���x����"Od<p�X<���� ?fRH�t"O���[N�f��Q�U� N����"O���Zcu���Q�Z:?RP�Q"O"Ē&��MX�yf��jLx#P"O@�{7H��{�.T�0�GP&�-�"O�4*R-�z���g��
Dp	3"O&<��G.I���5Fo<���"O��Ql݌o�V\�AŖ�@��"O��,X��^��*� $̄�"O��"�9w; |QwjB�= �Qq"O����$ص6�v�q��F�mpt"O<����%bb��iG��	qF"O> Q�	JBѴ����C1\
�!rt"O�-(RLG�_ЦEa�CMQ�j�C�"O�!�f��	A���h&z�X 7"O�\�A���k���Hvr���k�<���%M�	�kI�Y��I�Wy�<	�M�3~�0c�=����v�<)�*�5q+Z!��B���@\H�<a�� :��s%�	n�P�[��RE�<9�W�m�B�z#�� %�t$Ii�<	V@��*�G�vo��K���d�<��e�1k��+�ǂ[�`�9�x?A��ؙ>�'�����Ӳ�5���'|���O�P%�i1����n�1�����w�l�AED,c���`s茝
��gdB�8J>4j��*6��̉P�ϱzC, ����O\�BS�,��>Q�Z�y�ؘ�ڸCp���G�
k��W��MY� �4B��	WH�4�O؎%8e`�/h�D�(���\�NM����Q ��V�T
`����IT�0<y�CE�<D S�T3Q� �ŅڝE.����4ZS��ԥ�.�Z��[ e��@�shA�5��x��aK�R$}�`��f4�aR���x�"�H>�f����@�f���?�����i���h0+Oi��DX@�J1�����p��O����ޠn48�j�i���E�ɭ��=�f�_��G�h^���5f"Yb �a1�
P �
���Yi�5���Y&��@@*sT�����,O8���σ�&w
1`"���Y3�$��=a�A2QGA�<
2n ��#lڴp'#�s�1�u�\�d�!�F�	q>�U�ag��^{��56O��
��b���q��4E�ջV�S��8����m��OJ�O1F)���I�~���j�x�4Hr�z9|�i�'ȵD2��7��A<i�C��c��@� ��4,���V�
�N$���K�3P¸�[� b��l۰���(3UlK�|zVe܋%�
L��D0��������a����SŜ
q]p�Gfi���ED��6,�����:rfd9�����YFF���/s_r�?�=K�l���14��u ԁ1H���?1����Yv� �M�bj<c?A�C��'�T��%3[R9��OZua���_�R8�u`��<At���8L"�P:*:�GʘFъ�ۃ��!p"��h��dV��[DW�!��e�� !��Q�Э�E.��tw����0]��A�;^���y''�A؞����C-0�����K�FI�f"�OU�gꂑ7���X�.ĈCg�����Ȩ�`׼/�!���z��Ğ?T&`9�K52�������?K��j��$ҧ�0�`RC=P@���R蔙itvфȓ	��q����#BA��@lڞ1'a����u�)���q��G#Tq����/MvKq  D�4 $%M5:�r� �#�y�4س㣟����$���'m���slI�4�&x��O.j ���@��!�_�2���`
U A)� �� �@˗1D�D��o��. B�pP�]3X
$��o/�A��l��+-%F#|�Rʗ�2��AS󈇷����A/S�<qB��عٴ�\�9~�qÓJ 'v�%��i��H���O?�$VV�őf�K�����l!��G�-�ΐQ�NJ�)�0w�:	���̫tX�| e���0=� p(#oT!نyx��>d�Εz��'��]z��<����臰e�f�ks�J�3�~�	�.Hc�<�ÂO7T����((zP% ���Z�'mڹ��b�6W���E�dj�
P��C#F�"��#G��-�yb��_"X��.^�&k��¦h��M����i2���K>E�ܴl�zh&Տq��p ]�<���ȓv��jB�$~vBE0�S�ZL�@�'���5� S؞@P � �z��򤝗K�A�e4D��ٰ��9�6 �o["f蚕��5D��1[e��C�G3?�@m��0D�X�-J'�>,+Vl�6�*%Z�*2D�$�� @��W��Fa1iԇ6ړZKj8� @Ю���CC��<rw��3g�ۜb�: �"O���"	ئ2� �sv ]=B�|A��	,��yc��:e�듟h���K�B���v G�����^*�!��3�uٱ��4�,5Bѥo�v�A?,>����F[$EN�9��J�f$�s��	:��\"�D�4�х�	�/�(iE���F~<1��l˭{���G��'u(���B�iz�Ԇ�T1@%� @[o:�Y�f�Hl��=Is�Q�<ވ����TlÉ�T���)�L�ٱ�.e�&�� N��yB��!u��q!Cͽ�DPP"Ɣ%2-2ǌܔ=��Ca�OfXa��Y�|q�F�7�zq!eF,uM����3D�@Y$�8M�h�7gſMA����l�D72i�#D$|N̻�d��<���	!�F �'��V�L�2�X_������2H��bv�c!�e!���s6p5I0H�i�D���F�V���h.��f���@�G�H`f��R�B<pׄ1�r�B=sߐ��f	�Sv<�$F6��;]��a�j�z�s���i�b�>��n�+�������P�e���1� ��H���UOR����X&je$��o�<�ċ&�gy�G�Q'��D�Byz�z ���yb� L�`����j��S�z���2��4����a�0Ÿ�HN�,�`y�KQ

4���(m�v���B˿pz��[i�X �	�}�䬱S�3��'���	���C`n	�t��� �L
7$^x�Y��)Hnx��	�&0(�S4�{�6�)�@��fPF�x�.��M��xҠ����Jݖz�2#~R�)I�(M�\��dM 1<v��Dx�'(>9��Eȝ.��}.u��AK�Ά(P
�|��F3|�εIcΞ5&�n�'�.�G�,O�)��\T#B�W	Ѣ.���Q�3O��y���w�9�J�"~�Bf�ekֽ�PȀ)/�B�g
ʦ�!�̍;��I2�49Ó�)a�M�6b�,}l>�R�><�V-�<Z��b�8�vmE<[��	�~��qy��5���[ �«9G����U�"0L_�y�PIj�Ň	"�):�h�1E�YI`J�d(<A�kP=Q�uaS�E:@.<�#1b�|�'�U�C�]7��^��@	�80�F�iRÊ*rF��f"Oz�� � ��hؗ��*B]�1�uZ� �C�EqO�>��$ƛ ����X{v��d3D�,��
'bT:���Xl�R�Y�3D���ë�S�61Y�g�+@�8�0D�� R�w\f���ۗ�D\{V�,D�4a O�31r����-b�^9�g9D�h�ӅK,o�R��^�Zx�B`8D�Dr4,�%60�_�3-7�*D�l:W�;;4��i��\�u������5D���$�Uv���.I>
��)1D�T"���*7��h�I�vؑ��.D������$#B
�p���;��¥� D��Y݃Kzn�@IјF��}#v-*D�P�f��4��A�w�O�l��1���6D�RX�SN`��`��2�#2D�dq�a���AR�I�2��H��0D�PЅ�E�:8pC�$=�i�( D��֧Z�1MdPɐ�5\�|P��d?D������ʽQ�ĕ_�FH;
;D���I^!w���b��QV�9 �;D�H�'�Ð6��q+Y�z� �"7D�$�犼l~iq�V�nr(��"'D�� �j��çLZ:�DjUm�\�d"OH���M�@DIEV��$��"O��"b�l�X#�h
�gk`�Ґ"Olh+F���;����C�Ms�@1�"O��(�
�[�ex�/K�ph���"OdI����	Yg���qH�c��዁"O�M�e�O;`�Vm���19�8S�"O�\ڃ�G� ��Q�f*�w/��i"O��TM�:=��"�	L�2j�cW"O^�҅���J3��đQ��P�1"Oj0c7�[l�X�0�Ȝ?{"�Ъp"Odq�ԧs�8x�&K�\	�H�u"O\S�/P�7m4LACE�*��]b"O�8���5k�(�
ㄝ!@���"O�y��N�W��$��T�uB���"O�����S�����nJ37
,M�'"O��`t+��uܴ#vmn�vh��"O���g# �x�4tѷG�%N�V�S�"O�Bǀ|G����GQ/XrVݸ�"O���	�F�����C�'tB=��"O �s	R/0p1�Vi��ykK�1:�>�z��A��n����w�)���+���e��]��R&^� ��8,��\�΂H�)ڧ��Md&ӫK6����38�po�Ag0�ҡ�|��i٥U��5s�D�$_�@���,$��YR��s≫YI<�����<�íW3�����fy�Z�%�4��ˍ��xםK�>��Qx�F�rW���NWjy�L�4�Y�+\�ݨ��7m�?+�1f.	m��y�G����c砕�FAN�rק���DW�͸N��J�*�6�>Y�r�q$ވC��)t� l[览��^w�t��tdĦ@�pٓ䃞Z�<�Cdj��IFDhT(׽I?���O��"}��O��x�)ݐ	��8��U�P?��T�G��	��/[/\����H���O*H��e\%�P�1�١I[H�2���l_�!X�Auy��0�ɇ<g�$�S	$��P��?�,�X��	��1�`�d>��a��ʦ��"!��0|�eE'H��Ր�M�S�ʩ*◢\W�u���ͦ��a��U�@�Zç��5++�#!��7�D�j%�b ��O�9�`�y�J�F��a���iGv����;Ъ�A�ޔ/RX;tD�+K�8�k���D�I�r�O�>�ӵ[p�e��7U�Ȩ�ψ�&rJY�G�X<|[��y�a2�4��<��-�ƁړEW~���@�N)��8�M\(=Xvq���'�����K*
2��j�[�HB���'�Ԥ����.��\�RnW�A����	�'ĔY� !�@�΀HR"�:2��S�'S�J2�ܴG� �,��"�|��'Yl$������m���Z�4V���'�r0�WDӬAxD�KB[�L��'���g��&��)��$�!�.�C�'�6a懙�(t( ьB�'@ܻ�'�"8`3�6��3�n�b���h�'��ؠ�k^*v�K'�,[L\���'�d��gW	Ԓ�8��Z�Op�� �'C������P�zЙť\�EP4A��'u�m��$�#NRjp"�N�A+�D�'�����\�i����ģ=�
 "�'z�K�X	��}��#�m(��h�'[XP��l�'m^���s���aX����'*��Go�Q�3�܇Z�|���'
��	c�!u�ԭh��E���'Q�P��Ё&(ֈ�a�Mcb���'��:6o�"$F5�#�Tw��DX	�'ix`A���Ё�3@�vܢ|��'<���o�2J��Tr#�،\<$��'�t�hQ-F�$#H$�b�[:���'�x찃G��X�8�'a��
��':f��E��1�$1&e�>�rt��'��|���Ιu��ɫ5I��#����'�p���Hn\8��٥,;\x��� ��o�B�؄ 7�l>�-V"O�QQ����h��e����I=�|�"O�틀L��q�P��1��1#D}��"Ov|�EG�>�di��
p' ��"O�,q��PV��,��hE�$��"O���I%{E* &! p	���f"O>-��jV�u�́Pf�˯�Di�"OJ�p#�m*��¦%p򞉚�"O�y�S��P�x�K��1�ʉ��"O.�B�� {�AC�F:�ءRc"O!aa�2�6U��lYe�R%bu"O�p%�9�p�Kí�5��|H�"O4�h��κU]d�;�l���b�#"O�MY��K�&��u�^���ܺ1"O2	gg�,Ю]J�K�c� Ur�"O��$��< ��A���t��	�'W^�ӰJ��q��5�&��q#���'�,�3�Ё_6^��拎�8e&ٹ	�'ް��M��vb,ͰE�E;)`ب!�'�ЕZ7��M�th��(
.m �'��I�2�ͭ�y�C52x�`�	�'�~��0?3�8��&��\�Aj�'=vt+��*O�L���ߌf*֤i�'*�t a,ظa�
Pp�oZM�Y!�'��!��K�h�~P�4���>�89�'�E�g
�VY�	c���#|eD���'�v��foE#"�D�����
9:D#�'�R� E̗�y�9IѠ��f٨
�'�,��s���c��У��|�[�'�F�k1�I1f�B���"յ��${	�'���(Bۃt���j�A��e�,���'�E�dm֖���Ç�enB�`�'�`���$�	_�iu���y���4:u�)	p���o����ʂ�y�D�D�� c���{����d���y�F/Q~ e;����k���/H�yB�E i���	��I\�^E[Dɖ�y�/�}T�t*���k���Z��y`�*&$�]�d�˧�R� r�͝�yr*	�)��hC-&a<�9�����y�ŋ�nvH���/����j�"Ƃ�y��E�I ��f�*~0�3�Y2�ybKT`S�᷍S�C$�m9��7�y�	G�pp� ��2sSt��dW*�y�,���x2��e�Π�WiĀ�y2��{H�#��0�6�����'h��sk��%��!���KΨe��'�\� ᎑=2}LARc�I�Eę��'��ӱ��+yx8T"͜E�^��	�'?�E)0�05�̸��\�:����'K��8k�Y�P�_�����'�� 3F �4E��"�[W@���'_
!i!�>f���>�����'��� �Y�&��`�nP�8���S�'��'H�q���~��,8	�'�>I���a�a �ۘ}(�l��'�����L�46!�!�	��@M����'�,�!`�'^��m�&זk{�`��'�d�0c�*����6��c��s�''� �@J�**&Y�$�M<a��Mi�'��0P*��W�(�	#��#����'��}bD䥬�-vY��NV�<����K�@�"�D 
�Z�x�(�|�<10��"m�h8R��X
?���#Z|�<� H}!��"_@�� ����� "O`|���
Dm!!\��<��
�'���`���;#b=P�mʴ	<��'�������1Trf\�"(3	˖�Q
�'7"�#�j���xYd�.rXP�y�'���[��*O���^�{$���'��|3��C$_��a�ėfdT��'Ɔ,0��EP���`G4Ű���'��I�6oMg>���+�>�e!�'k��P�V�I�zt��K�
���
�'`����)Bp�)Z��xH6"O�(���f�80`�(Y�~
�"OB�hF��A����X>H�Рw"O���N$����$n�:j�X�f"Oj��$d5NiN���-M4aox�(�"O�V��~Ta��, �d��&"O����)�p��4�*v}�9"O��D��U���	$MK�_c~�+�"Od<��l��ܲ�I϶t#,�"O*��B�BU������R	�8�"O蔂��Q��h�SE��9��r@"OnM��ۖx/*XK�d��~W�0�"Oġ;7g��'�pD�tM��X I5"Ot裄'*��K��ϯ;L�S"O��1����̋���K�(`��"On��pD�H�������!?�����"O�a�"�S�D��O�A�D"O�h���(Z�}���h��s"O&%�#� yP&���Ƿ,����v"OB	q��h��`:'����0�"O@�ʀ�_
_�� �AKȩ,t�a%"O@�B%eӽdԐ<�DI��Et
��B"O�9��<�Ȥ��&�:wτi/!��N�A�<�i�CT!RN�Y��-_�!��B&[,A�t��N["���[�s�!�D�;	 �rc��Dƙ!�A�!��ԋ[����i�=f�.uX4�V�7!��<zrc��J,"A�>�!򄒭s�����k�DhE&��	t!�I�ODj�*�9fތ`{�c7W[!�Ĝ:z5���q	��+��D��lޖtE!�DZ�E��,k��خ��$�A,E �Py�L�+����'�
�Gfv���@��yr�ޚ����/W�9Q��ӕ�y���L�N��D�f��F���y�/ݱ5�j ��b��,,m3e�^�y�+�k�����*
Ai��O'�yr�$��9)� �������)���yB���v:~�r@u�I��.��y2猢5Lz��(�;U��B��\�y�л,h����G�}Ir4��K��yb�El7ȅ�����kvb�s�n��yR��g���W�H?A�%�U� �y�F\�<���nҕ	��)�,���yB��.x;�4��nT�8����sS4�y���7WN�J�F@/2	�4h�)s�!�>d�t,�Q��k�� ���.?!�d�.Z��=��h;43P�IU�
=!��A�$L	���8CD���6'��	8!���pu�}��(��gB��S���N�!�$O�.�p�x���U��!�/_��!�$(J^\,C��0ۼ|���0qO!��5Ƥ�A#K%]�t�:ը�-!�d�.}ڵG��+%����%�9A!�� �4�3�B@��]�򃁝X�-J'"O�-S��=_Ж�A�̈́�k���o0D�p�G���P�wY�m�<��Wi;D�XIQGO�U���jg`�L
va�V-D��r�ᜌL0� A!��:3�d骑m,D�pb�b�T`�رQJK3u29�,D�H��	S�(�4���!��U�hɐq�*D�PcqI��(d���|�T��Q4D��z�ɐ/;	$�Yt��#qDx�X6F0D���&���1HsC
94*p2��/D��C���M@��zr���: � �+D�����iڔ��v)Њz4�q�&O,D�4H��P�2��rGDJ�x��)D����MK>6��	�g�;r�ڑ���2D��0mS�|�3����nܔ���/D�@��H�NU���.9�q��g;D���C��zP�V�Ԟ@�*l�;D�L��̂\UdىbaN. �5(Q#<D�4x�j�)���b�:z�ِ�l;D�$��؈H �d+�`�lՂ��cC:D�|#Ƃ[f���̛�B�U-;D�<(��G=bz�Q��'r�B�*�:D�����6 ���0�/�s��Ѱc,D�t#W���](\��dV�,��[�$>D�����S0:�,}�� �;��ԛ�0D���e,�9 Z&�XwEB�)�t�V�.D�#Gt>��P�]�l�a�/D��Xb���gu� �寜;"�(��."D�0�'��8g>��u@5P���I��>D���)N��#�)#����3�'D�p)@MQ%�RĨ��"j�$qTF#D�P�qEҴGj*��k��o��ś�J D����gI�v�:��5��+����A4D�x���--�:Qkf3a��@��1D�ȸS��*VÌu���»<s~����;D�\q���S��P��tv")0��8D�4��J7>u���	�be
ţ�8D�x���w�u@�mJ�9���7D�D�g�W!xUh����|��9�Ĝi�<��*(����L+	a&Ă���\�<Y�'�:έ`�ͤZ��tZ�#�X�<��L:��ň���$�Y���S�<����0(h�H�E�1��bU�<�K��.����OS�Fh��R�<���,E�XQ��ǈ�p���pI�f�<9�H	C��e��0�BJ�Id�<y�H÷v��	iƋ��I k�]�<��և&�Q`q�Q�*�:�hD��t�<Q��až���k��x`aڱ�Dl�<i�gZ�s�逡���m�4�!���h�<17�Q   �P   �	  �    �  �&  q.  �4  �:  NA  �G  �M  ,T  nZ  �`  �f  <m  �s  �y  ��   `� u�	����Zv)C�'ll\�0Kz+⟈mڄc� 特m`�DB�6%p� �f�q�䐻"�m�|Mi+��.�c`e�	��IuJ܅b�"I�;0�4���'Y8��J��}��1c��)U����	��l%ʡ�bC� b�Ԛ�@�����B&� 9� ���X`�-��H���9���=vr�,��$�3b��4�WEXB�b5���1���G��z�*�4yir���?A��?A�⌽�g�X���`�r)X�������?��й0��F[�(�I)es2���O���؊\����6&���� T(�����O�ʓ����O���'	���O����tI���R�~��AY�8�O�牐�>�+�&�)������۴0�(��y��,���I<Y�D���ⓤ9>i�1ӑe��D������I���������q��?�P�wB���Q� �$/��5R��'~�6O��m��4כ��'=�6�	�y�޴`����'��3�
��K���{#��<���*�� �G�?}� �Ϊ'�0�W���LF�IX0�����@��m-m}[��i��6��1����u�?���lY�Ik^��5�<"�J�A��;:Ȕ7mP�K�V�i@DN�Y6��PA�,�D�tk>E�mn��MG�i���Y���` �="�5�j����B �ŷ!��7���ec�4v� ˃G�)�j��!ǔ(���@�֏�V�K� AO��Y�*M
g@x��pB��\��	�´i#^7͎Цu��\�Q�qR�,� zR����G(3~M"��ڵ��p���_|�,�I=^5��u	�"s��31��
d<|���U��sA6y��N�i����9=�6][U����2��'���'	���O����K s�I��'xD@�P �-nY�T��N��]�R�:Q"O�mA"�\�VƁ!�Ə�7��eB�"O����96��3R��-��%��"O���#ȁ1�И�F)��D��S"O��Jq΁�.?�	�R�7/��,	A"Of���Aif��Aj���j!;F��fU��~Z���<�n-�4i��	��y�5��c�<!v�@�U��y���G�]t�Ѣ�v�<�f�3Y4��*ʢK�H�!ʞt�<I�͝�3Ft(��͠q|�02�I|�<g"A�������ic�c�t�<	�mS�f�(�n�>�h�AR�����3�S�O��lٱG�;C"�,�B�:.�ʧ"O���a�ލ+�D*4��:�F��q"O(�#�>�:��R�� ���6"O0|�D�K�%���*�M&��"O�峕�O?CMh4�LZO_��z"O�ep'��8j�XaP4+�.2T��X�<�r�.�O(�LN �0�"A�C�(��"O&	���Rvސ�AaJ�M��%�V"Op8��K�3s��
0��[�Lpu"O����MD�ufp��Å0����4"OB�a�m�d�x��з��G��<y��X�!��������J�x�2O
$��3#A�O�ʓ�?����t��$0�npʂM+s��!C ���2㟿e�X��B�6�t�)��I�F�J:c�M=���� :B�rL�%�z�:e"��C,!s�,�z/�� T�ɏ@�F���O�4oZϟ@K2�žM`�V;dI�Y�3GSy"�'��	S�OO�Ɣ;� �S0	�K.Y; #��1!�$e�����.\����G*s� `P�f�Ox�D
ߦMr���ß���sy���y�2O�T 􎐁CJ���Ba�>�XQ��R�ϳ>qO>�ف� �3ܑ�&�^�K��i)��;?1*Ƨn���"|R�O�F����N�9�H@�ľ����q�j�D�O�c>��N'bhR�Z�o�J<�r$4���O^�����j�
tV�na
3���a�џ�Q���L�WMJ,{Şb��c���$2K(S�O���	k�,@@Y�~ni�%�Ҩ";<B�)M�Х+0��\�>��"��:-�B�I,}c��zu"��c��|`V�P��C�I�=��d�h^�+J�]��I!�C�	��lE�$�"V���#���
��C�	����0�˟.I�Z�ASKT(��KeJ}�Ć�d����P��*O&6�8׍v�p7�?����	<kD��"�[;����W�c��C��=
kN=xw�=T$*�j2�Y;s%\��Ӣ�O�̇�I	|%P�8�@
02��M�r'];��Ǳ*5��h��'eI��a�h�vr�'�`6-1�D�=o�`�$?�a#A�B���z���o¤�Q���OV��?���?���>׆$�'�%^��s!��� ����ۖ4���艟rb��*s�4�G8�l9��O�^b50��1eڽ�Tgۢ �8��0��	f��1.����Ox���'�򚟘�� �Ca(�!��7	rte��A%�d�Oz����T���A֫M1�89��+]2�O�O��(�Ȏ}��S�B�_������'��	$O��2ڴ�?�����iI4��Dд2O4�
���(_�0RR?���D�O\��c��Sb�z����(�T>E�Ow�(�`�f��s�k��+�\�X�OaRT�Lw�-r�Î֨��tô�F�v�t����2 L����O��lک�H���)�7<��ѳah�"X�r#���XB�ɖ$1��X"h��("Mh��[=?�N�?1��ӆ!�B%'��q�Hd��E~��8lZ���'��D�a�X�$�O��$�<	�����	���RV*Y�������8.:���\5T�N�(���)BS�	8�䜁�*4:AF�2i%~��0j���	 |�� i]�!�1��ORP1-�4_N�a���U���C�'k�6��O 0�*�O c>��?9�%Q�+� �	� X&xC�j����d0�S�O)X�V��>o �b�d]?���I.O��m��M�I>�O��	=vp	��K�d:Jx ���}�z�*L��M����?9���|2�O�B�pE��f�% ��Hb�ٽM��]����Vm�ق��N�џ�\c	J3�$Ul����J��!�X��0�F�jm��s���iږ����%5s��Gy"'�u�+��
F�d�I���0����?�b�i��R�@�	Qy��?��TI���V9`��Y��*��6�OJ��"��7<�	1��	�(/���'�6��OUm�ҟ��|�	�LF�H�v����d�B<��Xj�J׏� I�ȓ�T]��n���GC�^���䊵� ��9��=;�F�"p�ȓt��gC+7��� �[�Qoj��ȓ~�^%��(�,(��S5PB���o��P*S)��Hf�
!�XR�F{�'D�̨��9��^ }Ŝ��A*��wR���"O�ܛ���O²`��7m4��c"Oȡ�r2-lI#�oÎ+���R "O>$���B��0q��Z�`�� :"O�T�0`�Q?�=�Fni�X��"O�Ճ�i3L����-�>��d���'a��8���7$� �#CҬJ�R�8&`F�n&���Exybe+I4%���u����o>~,�B�͇~onA����P�4��8�BL+e)�1 �UY`��� ��ȓ$^p@{�;w;΅`������ȓK�^�A�S(M)0p�ە9�n9�'^�X;�)%I�de��8�$�7g_�-��A6�Y�3H�	8T�zj�
 �Ą�`�	(���:+L�" �!�D��ȓb�ڶ@�p�-Ąe4:���c�R@#rG�.��сD�ԥd�Ņ�	5��	4��Ȁ�@�Rs�� �U?�B�	8"<R��3\_�1�6�Wt��B�I	P|��VI�C�8����U�TB�B�I&�<��%o���G���a�nB��0JJ�$8�"	(�[�O�2x �B�3%"�s�����ѵ&]ZȞ�=��}�O�:ܸ��j�&�Xs��=>&�B�'r���B��J_4E3���0�&;�'�
�����p���pKԺ ����'� ���ΰs{�e��l�;i~��'14�X�+��g��C@�-��c
�'��)y�$�m�(�C�R㖝��X�||Fx���I/\��,�Aj��5�u�U�8�C�I�\�Xb��ω(�^5Ps�S�J[�C�	Pl�I�튦a�Hkmѯ}�&B�	4>�`�1v`چ/��D�P�mPdC�IjwvM۴�ʈ�&Q����&C�j�*��5N57g�{"LY n6˓R+"a�����(c�*K�*�"��C�)� ��ZĮ	�&4S�n�*4���@"O�9Z���24ҵ@$��*+�P�0"O"0kA�&?74�Kc��.t��"OP�� a5^�[��H�]Ӗ����',hP�'j�d�s��%^L��u+��4��'�hr4EY<E� Eo�bO��3�'�H��I�l#�'�^A~���'�FpE��7�|��D!#?���'8�U�ax��U�cF?��T��'����C��am��2��Q�v>����d��Q?�h�����(���L��aZ�!.D���d!��U{��sd�L�fy��K�9D��y�����t�4��"6��1cS%6D���e@�#"�U*�HM�6�~���6D��B��!�heHV"�a�
YR��'D�a�L�_�& �flG;-1�D�P��Oz-��)�'!L(��_<F��)6`�',ҖDZ�'���DրE$�"�D��:�a�'��|�P���_��,He([�<�2�[=|%�DR�e*��k��TW�<���d�]��f��ea�T�<�T�Y"8�
U�e׶O�\5x���Ry��+�p>1 -C���ʆ�ʵ��)f]N�<��+���D�χj��i�2�DH�<��اs��12EoT!,q�3��G�<)�e�,t�j�m��aB���&X�<�5�A	/���:��8AU6��⪉Wx�H`E��8��_�6�Z#\?��;A�4D��	q��$��)'��FƆ��e3D��c%�8K�Ƚ�g��,�z�"1D���v��U����C
';Uh4�� 0D���D���1�l���Ʈt�*p�Ec D����.	-gNb��P�)��SEG*ړVK�@D�$/�F��4w
�}���G���y���;>��a#�W	n�s����yr� �Fd)�R�/Pت�j6 I0�y��P�v� 
���O��e����yB�Д6��p n4L��1["�P�y�� b��q4-E�/�xҪ���?��F�h�����Ո�π20 �o�@���"�g%D�`�ƥ�� ��r�mK�F��o$D���*Q�PR���$��MJ@�J3�"D�(
��##t0�kG*�B��>D�����Do6��7�@�?jr(�A<D� ��+ʸ	��7��d���<���C8��A��ݍC(� Z'�� aB�\"�(8D�$X �M\C��Q�̡U��SrG"D� ��K4�R\�sb��{ي0A%�!D��z���n����
l�p�>D��C�!��erz}���_�B���R��:�O$-� �O� RF%���>��0.�9;v
(�#"O������A���P��a�s�"OP��d�_8J��d"�E k��K�"O����!O�/Lxsu��t���`�"O|D��%R
)pDE�$�
lO��	`"O�A�� H�m���F֌6�ځ21�	�o��~��F�I�(M@�2_�LҒ��B�<Q������0���^��� ���v�<�p��>e@ܨ�B�� :�*]�ȓ|0�y+D��~���4H��n���>	�Z$�+{�t�X���
|$�ȓ.`>�gb� � �R*Ɖ3�9�Ʌ٘#<E��N�1��lPj��r�$q�S�	�!�$\,E�ʱ�d&�����!T�
�!�� ��)��!<Bp⇭��-�>�y�"O.���cǚ2>e��͉�cw@��"O�hQ�G?+!���E�*`�S6"OVm+���6Ծ�3��"�yQ��  '�O�)��Mê2~<��E���M�"O�͑WG�d���u�I�a��9��"O����V�M8M�D�4/�@��"O�]13(�)$���AE	H,2���"O6�@a�"y�biI�N��Щ��'�.T�'~�<��U���{�e�-u�\�y�'f�mz5咽O�~D�fH�0��T��'3�m�S䖰W+��*�.!�&�s�'�t!�@%�z�ąkENCJ�
�';~� bɇ(+���ڙ����
�'Ǣ���gslr�˴'N�ڪ�+��DW�Q?�#�,ȋEg&�2�:yq k(D�|T��q���b����{	*D�$�F�(I�y*G ��:~�(b�+D�LZ���#�"t��E �)Lp)��H*D���dI�l�lE��\(W��8*�"+D� �ٝ{���4�A6�Y���Of F�)�'f^��q¢]>n�j��s�RU�����'c�mK��[���#�M�TD�x�'����'U�Y|E�@zkt8��'��3��Qp��07�P(h4u��'�.4�R��J��C+X%xdB���'�L,yk x�8-�d
e�l+O�C�'�h�����13�}��Aèl�#
�'⁓D�G�H.�� $nzǮ<�	�'�su�1Y����y���	�'@���T�O!P��52�]�v�\Hx�'�j�%���%��!�R�&eff})�������Aք�=���s��{���ȓc��A����3��`{Q��!���ȓ&c�Yk0 ��~B0��Wc��,@�ȓ[?��b	*Mو��c��SU@���cm���IB%��{`c�\T&q�ȓp��ㄭԃ^�@u{�"K?=��mD{B������8tI[�P�jy���^��"�rE"O�Xs7�[6&�i���'ͺxK"O�L��`��NÚ���P�j�"Oa�tm¾$��Ac��A{G���"O<��-�F�D̊�&ۜ��ɛf"O4P@#�$�UI��V���e���'�Dݻ���@CX���m_�� sA"/�B�ȓN0��+��J��8� M���Մ�$��r� F6T(t��,9
q��fۘ���ԈCm��HO�x�@�ȓsLLр�kW�$�Ƹ� W$?�n��ȓ�h��OY�U(�=Y�/�[��ї'�\S�I��	V�?f1ir�� ʡ��	#(�S�V)H=�1�d�^��܅ȓx�x(BC�CY Vjb��a�A��m���#��>E��4qvO٦El�Ɇ�I�:,��H@�Bu�-�s@]�k�����h:��*Yx�!CS!28}R�M �C�I Y;��H��͹K5��!E 9
�C��0l���g�.�n�PsF,	�vC䉞rD<1�j�2T�Ҵ!�&6B�ɡ	e�m�VIR=�:ܲp�K�C䉪y���於��P�ǐ�_)�H���0�z$���;
����rb�D�ȓ~�"h�"¿?�8( 'řg���ȓd���� !#y�4m�� L+�@���S�? ��R���M����FBWY����"O*\���A�p)��^��L�q"O,<�W-P�w_
m����t�2�$�'*������S5k����FR8����%(s�8�ȓxo@���_�3�H���i��B��Q�ȓY��:P�T	Et�[Wk�� ��ȓ<	�IS���<�����r�P��ȓ?�� �e��]��,�g M�!2N���9`iy�͜	�6�i�C�76h,�'�ڹ �g��E`c�!&��y�g����5�ȓ>��=����/5�TŘ���m�2��ȓr09� ����X�Ɗ�3�\ȅ�%�\5��D�-'�:!�l��ȓ]=�@P���xJF�[�N�?2���I�M��ɹ_ܦ9PV�j~�5�vHɖBwB��* ,SN�k~��e��/C#B䉦a�by�Ff�C�Iس��')��C�ɤ;�u���N=���s�� �C�	�z=ҙA�˗<Z|j��F,�6chC�ɩM����D%�16V)���9A���=a���S�O�`Ʉ)34���6�( ��'�H㗩ֳf@<�h4�
|�L�
�'n�5���T�'��l�@�^$yT�p�'TT�a̙6A�[Ã�;k+�� �'^rQ��h�lHZ ��a����	�'����HT����R��L�K�x���#v�Dx��	$5'4̹!��
*�`p�C�U8B�	r��A�
X&��]�+,,\
B��M���ޑj��=�Ph@>P��B�	
}�2	��{g����C
63ĪB�Ɂs�vL�g��,2��v�y�B�I�8��|B���2E�T�̒xc>��=1H���b�J?9H�x�w��06�CqN%%Z6<a��	Uy��'���'DN�ӣj�����o�9Ai�Qb󟮝K2H ?p���d(D!Z�t����!D=Ե��^-r��I׭\7cd��r�C�� �&mE�H�]&�����-T�2����I�f���O�b>I�����.^0D��΍�>5�xKSξ<��wu�aҏ�
aE�LCc�}�j���	����ѩe�H=���jP�5���W	9���!|�^E��ҟ���d����Z��'�j�R��C4���G!Q6����'E<j���P��R7�DO���T>��|b�N�md:]8�L� svJ��2���<Q� �D��d��߸�Z��I�>q\��A��h!1�X2 M�d;!R�'��)�	:?A!ˈ�!�z�D��:	Z�����H�<��FL�JI$�*Q�	 �e�P�B�'��"7K^�!��+PB_9���䥎��?)���?�3hÔ#?�r��?)���?�����d�%�����B��rp�_K��������Ò41�)�4�<Fx����Y/����< B����d����':z��8N��i͟��DK�%(d�����I�`��)5?Q!X������?ٜOp�Ԩ���,w��u�5	[:@=�U��'�f����2A�i�NO):^Ȝ��0A���Sٟh�'a��@�鈶2�2����A%*-@1&�9
�L�(��'�b�'s��h�������'q��Pa��;\��rM�^]���B��%)P4�ǅ��X�F�'�h� ����=y#��q\z�@�y��V쟁�� cs�*,O��+�'oy��/� � E����]��@�P�'����3ڧO=
���	�;��ZD&͚K��	�'��X����x²uZ� �!HD�I,O��)�Ir�:�~䥟�p7H�	j���s'��L_>��@"O��`�$&��Ex��T�bkz�Iu"O�SPo��8�<0��F�=}6nYX�"OTX�dI�:g����8º���"Ov�҂L����+�dĪ�۳$"O�hr��/~T���.f��t���D�+q���O6z�:�ٯ[&]���V�E�\9b�''$H)����a`ˍ�6�b\�	�'�P$p c5\�J����6qd=`	��� ��5Ђb��Qx��PY�EV"OЬ�ѭ�$}��5�2�.{�6�!4"O����)j�0u�!@A�28\P�@�΢�O��}�A�f��D�I�Jȶ�C���ZF��>��kB `�|5+@W�Z؂8��	��5�&���A<Х�gf΢44t��(��5�wL��MC���#�(u��ńȓR-��b�'@ a�;��>)�h��ȓXX�����V7q��EM�W��<�I2Q@���d
�E�R��/'T2P�lZ!��9v�䃵L� N������%�!���~���K�w�ʤ+_�!�$97vbPKa�� �8�	�m�!�K��q�����%2A��џ,hf���M��?�O�� *�[�@�$��ӏY�]��K��^�H�Q���?���\�B�˦	Ir�d���ITY�6=�2���L�O�Ș#W�ޗ3������7a]v�I�+� c�"L�1aU����!��127���4�b�LK%x��##��O�#|���Վq���CS�ӔAI��c�\�<�� ��M�EM�JZZx���.OZ��=XB8�9'CE
��D�#V���Οؖ'�O���.�P�0���rT�Y"�Q�Pׄ��:�|%��C�-Y�,yx#��[Rn��?�4�ēA�8b>A���Ԏ.�hdq�6z�y��(?��O��q#�>��y2DJ�@��{4E�41��Z��ֻ�65[㓟p�I���.}Rk/���ck�8hUƆ�n��t�!-^�C�ti�I��a�'��>�	KG0�C"�$dߔ$�ƀ̋aHx�dD>}�"}�`	��I�����pE�-3сv\��s��A'Ę���I2�N�*R���F���cb���6�N��놫�?Q�(@��v�$ɷr��V���.��B}ތ����)�$����)��$��c��sQ�?����?A^HQp�2Ad�x0��{��I�/�ҧ�9OhT���*�&�5H^�ʶ��`�T�⮃�to"T�'*�mJ�O��x��)�r��cR*D�;1��AIɸy��@C?��MN~ʟ�dSq��$@+V�9!ꈁ}�i��8N�2�_؟x�uD�<u2�)���A�R>��2D�.D��)ai��q]��h�
(��lm��4$��٪���O��4E���x��E V��k��^�Jh�&T��$�tG{��	{���g�H(�C�0P�d���"O�%�P#�\�d��SD����
E"O�#��JV�-�d�3{f-a�"O��k�#�/���"ʆ~eP���"On9�W�M����!/�5\v�4"O4A*I-+n��b���"O���៫(�h�3-:c���(�"O�L�d�9Ȁ�5+K�6"O\Б���<k�0���+ި���0s"O4�	�Y.Yt��kC��#R�0�"O^�JtM��`@ ��d͎�	�"OXh�i�>P98��ad�/\T��"O���Z�I������,{��D�dZe)«^���=�FN��<X�v!V�,��}�gꍋ	"y�QL�sͺ%"�֬k���8�C���<��*V	&��쀑=J�ٙ�K�O�J����۶_�&\
�� E���1�0I�|1���îF<�Y��J�P˷l�(�$���t�6h ��j�>i�dqQ�%�=[O�m�tc�7x��B�	X�lL{�	�<��@�K�G�hB䉍:G�H #�Fֈ���l�2�C�ɼV�
�%����9�L�Xp�C�	/M�0�AB�F�݈U:�+$-�B�;R�L���-����"��+vB�	� 	���h�1B�����x��C��qc�� �B�m'P�J��^,;ΚC�ɫTl�IQ#b�.f_��#���bC�����yPe�~ �0+g(X$�ZC�Iu���h�P7(����ɿt�B�	.7Ťd�!�ǖ������E�I?�B�I�x�Ɲ��"#A���ڱe�8{!B�)� xys�w@�����
��#"O\�z��?i��	vLQ�|�~���"O���'ď$���K�7A�:��`"O���`J%z��S��;]|�x"Ob��Q�K�y��H���7�<��""O���`bB/Q2�)BW��7�H�2"O�P�*�T|���ӮH��Ss"Oh��q�W��p�u��bD 2�"O�y�ai�4��"	�7C�}Z"O ���˒+-�ry*RF�#8��%"O8M��y��\ �ZEs"O����;O̘a�K�$5�U�"O�vH �����	��q�� S	!�F�"�Tepօ�!�&�yQ!�q�!�D�6@^)a2�ܻh�"�)��NL�!�d�F��ѱ�I�)�N�P W h�!��/�la� [�XЬE���0q�!��
t���&�lDR�b�2�!�$V�(G�pC疿u-�}�5O�}�!�d�h�ˤh� L�x8�߄�!�d�!UfV��C�^�&���)����!���*l¤��2|���h[�8�!�V�S��(7!ގES�@��gOi!�ݽr��)$�XC��ArM̞Z�!�d7D%P&�E� ���P��ս-�!�d�Jl���K�C�,��3Gو�!�<q�,أ�~�<P�fV9Uk!�D\#Z��hfA� +����μ^g!�߾J	X�AчH|�� @*[��!�$[�z���E��dj��xц�t�!�ΪU�\��&!��ze�4�ckB?�!��	T"��p�䕑:�v�jBj���!�d��d5��hM�'�q8�+^*�!�	�}�d�0���N����7��}�!�d�@2@���ڷ���D��&�!��\��H��
�J�f��	�%�!��=~F<<q�ʕjmde�I�6�!��&2���h��7&V/'q���"O�!-%�Дӵđ�c>Q�
�'��ժU�է_�� �fU7����'T�8Pe��`2�tI �)b�p��'����G�3J��Y���R��<��'�4���#�	GT!@�(��X��'���H� \9Q��ǡ��mR���'���`�Q �B�ҡ,�h2(tc�'��<�$�X3Fm�l �È0�R5��'���(F��r�NN�QV�@�	�'G�At̏/o�0���-xC��H�'(���`啪*U��PR��*#��A	�'$dɱN�"T�4PP��H-j- ���'����/7��<j�ɂ�`H*x�'v�����Ύd$����)c���'��]H�BP�@>���й`8樒
�'Y�HX���C����)X�h��'�L�����T�A��}:�I��'�)Z�	_���Q[�ɍ�|��|+�'^d��'�1_FE��Oc,d��
�'��1��Ї�x�S挐'!�
�'�$�CBDR G�PE�0h�
�d$z�'�ƥ���]���E�;m�~ػ	�'X�ܓ�k�:i'���`���;N�1��';�J5'D;k���p��.��h��'�^��Rh�3#��ʑ��,��
�'o��'ˣd��P�Q^4<�s	��� ���K�Gft|2�K���"O���a�����bg¢ ؈�"Or`9W"�5�z����>��r'"OB ��Ԑh3̨*2���T�)"O�I9f$��
��qri�+��`"O�!�(S3
�r�����T�8�Ys"O<���g��X�0�`�*�*OXH��`�\��:�g6@��P
�'Vr�fk�/=e��ҕ�?�z
�'��Xq2$V�zش2rD�=�<̺�'.p����9}���4L��.��9!�'�=@fI��yAoܘ&�ތs�'����B%��0�=4�|<��'��D��� 2�u�� (�fE��'�XU��b	����Y��B�ꈡ��'B@d�G��;JF���ĉ�j���'��Y�Fl@-��QP � ~��<��'��<�u���4@�)ҥg�h�h�'�,�sB�U0��$��g;�A�'�ju��B��BPY3ˀJ�.���'�����H;?	H5��BH�>7(h��'��u+�J�K�=F[(:��y�'0�$�LZ�`ܚ,X�X;
�'r6��L�L ��)!�S0[.�q�ʓy�xą��,���B�!������3��I�<�X���f��&i�ȓ] d@��������j�*C�ćȓ	*^�b��F�;
 ����ц�� ��I�T�%�d��MÚ����LU��հ0@�|�0��5j����N��H� �4܀l���'^�6y�ȓh����,į;^V�����\��fe�����I���G�	�3Q]�ȓ0(f��q�9,���:�냭D�"	���}c	A�E*����lH�l� ���pXe����~U�Iz`#��>�ȓH�F�`ҿ���I��׭q��ԅ����j��ѝn� S�.N#�Z�ȓM* �ЫVÜ�&Ό������gm�4���`ü%F�݄f���ȓC��ʀi�"ڠ��	Z=	�e��tڤ1��c�N��)sΚ>&��	�ȓ^m��h�0t�����>~����|�h������Y���̷GNP���:8�h�\�p�6���5r��ȓwĠx��kN�S�9�B�'x�"Q��D�Q�#�*ihuu�[�JH�ȓn���yB�VF���DL�v0��ȓ@��L��:/*���� ��E�� H%�b��4r�H�Q�1#q��ȓN�X�s�>�0a)&�FLj]��Z-�xi�\�Q�v�*Ba_�L����ȓy����>X^�j�疳>� ��*��r)�.�Yt��M�x��v��(��dݏ9:=@�=h/�a����`�uꉘo�0ĠF���q�ȓ.6Vv�7]6p��t&�A'�܄�K�B}�"L*%��SEHN�E^�Ʉ�M�\m@��2�h�&��S8΄��}m�!���"��L��G�7̴��#
���!+}��m;g�^2��ȓ?Y =÷ ��#�
\�ၙT�Z!��y�dيG��/]����_�R5x �ȓdF�ծ��r͘#kQ[�j���S�? �P�,��JEN����(\Ș0f"O2�:c�IYB(�e�q��٫Q"O�A�f�?	�B�Y�bNd�"�;P"O.X+�d�(�vDrrˈ?+��U��"O�z���<~͂ܨ� �>����"O��B��B��\�4NZ�~�V�qd"Oݚcn�X��5	b�>޾�2f"O��L�"/Ў�r�j�2����"O��``F48��BQ�W�^,�6"O ��&�ր+ D%�"���x��mP"O�y��F?q�\Հ	]�()"O��&�^ 8��m#'ϑ�Z��"O��k3+؅n�*u�EG.2��1�"O�(�k���O��1�zR�"O ����΋h�<K��m�Aq�"Oz)���)T��I+��=p<l��"O�9 ˀ+���b`i�%��"O�=IG��H�������W.Yr�"O
iQ��ÈyD�suA�RQZ�e"Of��Q-��a�(�Z�/�?k��$��"O���
�;��a�`Q�=�����"Ob�d,� b�tq�J�G|xU��"Obq���юd�$Dqīyu���"O�	�'Bۡ*�4ܻ/
 r�̊�"O��R�߷$�����o��qzن"OT��"^'HlH���Ƭm��ca"OV$� �"H`���"�_�f:�"u"O�9�6�.B�Z �eKGd-�"Oh�2����T����<;E�Xq"O�+��զ\�Υ��H�o�L��"O<�AVGq0�5���W�|b5��"OH<���#�X+dgYx8P��"O6 ��J��n�&`��[?��#�"O���o_��Q���{/�)��"O�4z ��Z���ҧ�����AC�"O�� S�=� 䂲�D2�j��"O�1�"��O6�(�bϟr�N$�7"Om���0����_� p`�S"O� p�O
Fr���U(�1Z`�x�'"O�����"R��xg� ]"���"O�p�@N�X�*-�pe�~o�Ty�"O��Q`��^rr�i!D�0fz��7"O�U�1���l%��آ��eZH<��"ONdB��ҜnojU@�W7F�L��"O��ؤ�G咐� �zͩȎ�y�Ɔ�S\ �##N@;��`h�A �y�� B"Ver�ڶfۄAJ@"��yB �%F�h��PŖe��X�K��y���E�Pԙ���,� j��
��y�H�q �ؗ.X� 0q3#���yBNθ7��H�%��`��x�U��y��� N����͙4by|���%F(�yr�(K`�}�6ȃZj��H���yBh�0�M���5T�V�P�L�6�y�M
�dnБsC�M��U۱���y�>_�D��t�@��P�ƫݙ�y�g��>}8�!ɞ5<5|�21+V���'~��Ȁ������!h�,�K>)�!
�}:d-��B>��rmd�<� ��>M�I*A��K=_�,��'�~		F�Ր7tQ�c�
;\x� ��'���l�+N�<PZ���%g��'l���$�T�IP#�gѶ��
�'\YT&�$c�T���Pv��`
�'9�Q�/��r��4 �ȣ=�<�
��� &Dq�hףdz�2�!��+ژH@�"On	&�M�-h�u!�4��,�"Ovɣ2M�1��;�g��m���B"Or��B�ڣP~��ކv�P��"O��"
�>�`�O	�vfҨ�"O � q_�3'�4��-�r��9Qw"Od�D�PF�d���앻
wLi�""O��m�m'�$�0# ^��x�"O�U��4E84�c cɐ- ��8�"O�1�1��C���Z!�ݜ@�\�q"O��ǬśX�V����9u���v"O���P�T�] \����6�:��"OP�q"+�-lf���g6��4��"O��Xd�3[�Ȝqvb�p�q�"Oм�oR�X��I���*|hx�"O~A�*�@��D�.�."��""O�u�mί����UǍ	"��c"O���2�D�K��yӰ��].D�g"OԨa6ȁ�K8����c�B�4"O*в+\�C%xqs�dǸ�""O>T�Ҍ	)ܼ���]�N_j���"O
�#���n$�9���1��X0"O����V�Wh6D�@�T�#"O�����E�`l��C�� �/!�	V�Q���7��1#�!��XC!��0+�̰��`!��b����!��_&q�Fف���uk:I�g�Z;4G!�$͕=�$��ĄnV"\QԦ�$e�!򄝺3�FDy�m�"HK*,i �V�!�$� -��V�^�eWJI[$��#�!�DZ�fƎ��-� T� 4�W�޼/!��4l�MK�E�$�b!���I�@�!�d��eh�q�5~>(��E���!�^�)����D�2V>�P��M�%�!��a�����D�x���7�!���a��,L�!ihI�n�c!��ÏE�Pt`�HвL�h��j�#v)!��d��@5L�^[���`Wc�!�$ˉW8��p����nEt5���Y`�!�D�~�ԱQ,ڰp�m@7����!���	_� v�+wOH�q��Ѧ&�!�O>�Z8k���B�)zaKF�$�!��(ꅬ�(<P-)��Ȑ�' �%��>�𼛓`V�p��h��'�\1�@U�<^U���ѳY�l@��'i��R�?8�UA M�q��'ɠ�UǘYq��HVAͭ[t���'�p�xe.S�d��x����Rj�x	�'.V�H�(�(0�i�¯C�]��'K"�A��0Y��!�bD2u��%��'�� �V��!Jޒ��4�CAV��#�'l�C�O�"��T�a��-��4�
�'���1Td^T
��c�Q� ���	�'j� �w*Н c�N���%n�}�<���jdL���J��i�͋R�<�A ̀=��!#��[�`R1���m�<9p%Ԁ���������H�e�Zu�<9B�!����6��wi��&čO�<9�/�{#Pa �Q$�wJ�<�g�E1M�`���$U�ЉF�IG�<v-3��А �P��%:Q�VC�<�(��fuR9�wF�9zD�Q���M]�<����F@0�a�@�2Y �I�C��X�<�� ��v��"#�)-%̨�LF�<� @�Pq��7D� p7��Fv�1�"O���'h
^<{0� i�t��"O8�"�"	(k?�Y ���6$�!�"O���ϐ9~�� �ַ2�^��"O����Q4 �8��Ņϸ���0"O�x0G�̹}���%��Q� ��U"O���lQ&8�F��@���t��"O$$��IK�7�,���@�NY�"O�Y�V�[6~�Se�^����k�"O �Uh(������@,F�<-�u"OU3$j��W���Ĥ�=s1P"O2}ZƆѥfGָ��O#bh��A"O@Hz�+P�p��-[�͆5W�aju"O~��f�����	G"�f�@�b"O��[�#�!L،8��2r�`a`�"O�����Jt����HŁ��4"OΈ���Wv��[�
 &��Җ"OD�sJ��%���T���dX\K"Oj��%Z�9�V�Ď^B=("O��؇���(�;�MT�kG�h"O�� ޘ+V�����C�D� x	�"O �x��9U��`Ze	3�8X�"O$s3O"Р5�4k2'�H�"Ot�:୊�O�����i����(�"OL(�2۝]������W��()�"O�͓E`��?�fL�7cܑi���j�"O�����>���85�m�"O�H�
1{�N0y#�P�*��5"Ob�S��>hO���C�p<Q�"O���PÙ0f�m
�J
9�4r�"O��k�C�%&�����/�t�ñ"O�,cv-݆�H��'EMV��AIw"O�#�)�6�&��s)�==�;�"Ol�#n�&"�z�k�h0O�Z�*�"O���6��5�L0I2�I�.�XHV"O�	��B��Q�(��3-��|�u#�"Od�z)�t�5y5#�9�`���"O�p��*�,4#1�
1z�� Z�"Ort��V�&�*��/��t�"O20��׎57�x;t�¯ij�e��"O��Ĥ��mƲ��4�	g����"Ore���+%y@8#@��;\���"O�H�-@�F���oҠj���G"O����$[R���ΜR}����"O:D%��{XD �3�S�Vξ\J"O�P��O<1M��#��2G(�(i�"O�M��� H�V�z�eG7	^�X�"O0�S�'�y+���W�
nL�b"O.̋W(�7o �#�*�,EQ~���"O� �)�n�}��#� i�X�#�"O�arGM'�����,�h���)�"O����*�8�����8f�P"OP��T ��j����a(��2���2�"O�(���]��谛��E�8�t�c"OB5�P�Z"!�^i��'�]�x���"O���5��k��,�v	�g�.4��"O8 �KBM�(��"�S%I���5"O.����M�n1"	ۑ ��$Y0"O��@sM;��<���L:$��"O�Ԙ���]�@��Cd,��"O��ˢ��
%;D���G ���:�"O����Y-'����g�-j�DM�"O��y��[:�.u��޴j�"O|9�[�f�*�srJT�"�[�"O� �`c��A& }��������C"O\��3g�3e�\([��X7Vh��j&"O�K��Rx%45��acT hv"O6e��̛(
� ÈU��"O��j�Ë�\z�`'H�m��Y�e"O51�I�4N�%�l9M��1�""ODT2�#����Ӡ=j�(4�S*O9��ʇ+�T[�FpM2�'HI;���J�t�1eŔ4���'�0\�6B:6��T�!fa�B��?DjZ]+�'�*��=	fJ�$y�`B䉾3���B�,�2anE��S�|��B�ɰ2p��W�
�M���QCаT��B��5>pj�⡯���d0G�"��B�ɺo�|2�G �@'6X�B�	�Ni���'V�.������A2ԚB��62�>� �R��P��#F.pPB�I�)I�\2�-�0�4����=J�\C�	/E<m�-�]]J�P��?k�B�I���}23��P��y���ʒ&pC�ɑD�VaM�Ll�������P� B�	�_�p1��F8�x�apmQ�z�BC�I�C��@��
�0h,nAGL�&C�I	CNMX�@�\|�p戕j�C�	�[��	IEBޯ6� ,@
W _:�B�	0k�
�gl�#!O�MT
�~��B�ɧmd��cH�?f��i��װ}֜C�	�<(8��앎c��쩓���RB�:h:+�='QV$��ՋQ{��P�'k,�c�H"`	F���O�4�̼y�'��	4$�:��H������ޒ�y�`͡[���Q�	{hp�X�B��y��A=v����ٹteĨ�uI��yB��M|�05�]Ѧ������y�M�Rw��� ��%��[�GP��ȓ-@���B(�l�8�0��g�rh��V��Թ �p�)��ȉ]ӌ��ȓd�D���\:�B�3fo�)�ȓl�v�HcIW�WvQ	U [�qr��P}dU�'��4X�zy2�I*����'�,�k��
lt%��_v�����!�h���PU���ŇU�VM��,P,Ms�W&�&������i��.���gg�duI�Ro�t� ��ȓt�KǢ�4"J:(�0��e���ȓ]]v���h��t��@�t�n���D�4L���0��Y�2��D��W�r(1��?��9�j�\Q�Ą� �@�[T(��)̰�B͝�b�fY��nB�����-U�@��OC5$H���Bې$�c(Ӗd�����
3K`m��'�"TP��^l���Z�-	l3�m��v'�#�n �VM��N�1K�,�ȓw�i3��ME�.�2�K
u?J�ȓl�.���@R�C�d�8�K�K�
Q�ȓ??H�)2��t�*��bD���,��ȓq�@B&D9��p(�L��6<Շȓ-? �{V� ^�Ni��'//�F%�����`��S�ipv�!�ì��%��ih`<Z�N�6`�r�G�V4|l����X���������FC;&��5�=�#�w���%��5X�$���f�	�-�,	����FȰ&��5qC�I�}d$T���H�.Z\|��76�$C�I'X�֔�l5#(�E�!Y�C�)� �ZQ�<��a�v��%*p!�"O8T"B��q�� :�.A�~!Vp�"O^���ɖ[>�+��R�;9(LrQ"O��S�̓�T1��t,
_+xd��"Ot���	� ܢ�%;.6��"O�0x`��"��A!a��M��52E"Oƽ"�ߴ#���a��)�����"O.Ԫ��ݵK�p9Vb�z�]�W"OfqX&ʣP�bL����WbA��"O�D�w*�%P:���O�Z,Q�"O@��� )O�mH��pF�S�"O�M�AdX��I3�P�H_���6"O0D1Ɠ�}J���g�>hOV���"O����14�XY�2�T�*6|���"O`��ꁻ{D��X Y�:#��H�"O&�I�uԬD12h�<�)A1"O��B\?,����W�I2"OEر"�12�j!��>#��V"Oq�L˹@Z�뵯��:L<A�"O:Ta�G��39j|�c B���ʈd*!�D�q|�+�$���J�.�+�!�?N~a��V��%�����!�d��5y��1AI�(M2ɓ�|~!�d�4��䧓�$��AzW�*�!�d����aXtc�x�hp��CP1!�$L�&�����^29^9ӧ�լ>1!���	-��H㮔y.���wh�%!���
d�(D0�/S)� Y��8R�!�Ѷ>�}z1��
Y�( V�)r�!�,�.�je'J�f�¼��DVV�!�DO&^h��s�O�jP�h31m^6xZ!��1L@��N�I<�x���C�x!�Ď'za�#�N�#CXP��!J!m!��/�J=�Gb��N���#��Ο]l!���|,����;�D�82jɐ@l!�d,�ݩ[!"� d�U7H�|���'wB��*�ޕ��A�8ʥ�'C(0�!��c���#��4��(��'�~X��zL���L#.rpy�'-xxr�2e��A(�o'\�F|�
�'�P@�#�̂q�JDi�)	d"O 1�ˑ�v�J��\��
��"O���nO���a2���s	�q�"O�����_֒eA�� g$*�Xb"Oܠ�
X�c������E~���`"O a1�ڋ0F8q�e]�>d©b"O�-��
�,9���%EU;G^�)G"O �cS�*P��e��M�%�T�"O��S��f;I[c��hm���"O�<�"�Z��U��FA�pÆ�r�"O�l˷+26:Yw+O�\\f5p�"O|u��^�gN\�9�꓉wʵ�%"O:�CD��#������$Ev���e"Ot�Caڀ2>�usq�1);����"O�)E@��JC����p��8�"O08J È��pPU���R�5T"O�M:IG�b?2�:a�]�f����"O�1s���W,��U�
-�H��3"O.LP��%XC�\y�IY� �M�"O6@�g%�Y�jܨ�����D��"OdyZDe� |����/�xI:,P�"O�$�����
���Α#���X�"Oz��@��î���2V�2 �&"O�	�#� Z6"ǋ��I~|�ѓ"O� N��>'�=`Ԭ�Yz��z�"O��b�mF I����TA>~u�@95"O�`�WCW���xtIĊ���"Ol+w�ˤA4}�Gԟ]�~���"O�ꖩ~i��#Bgkq8�0�"O�Y9���H�V���P�@`
P�U"O����J�_ � X�Ꞙ2T���c"O�8�(�NZج��,̽��pu"O���,)z�.�@��X9:� A��"O�ܨQ`њ+0x)�r�[�D��exA"Ot��`N�T69���2*�"Obp"�oH @�AiCmC�h���[�"Op�h��'YW.�k�k���Q"Oz\1cM��f�V��1@�?���7"O�����|�`4��!�8�"O���D僧#��mi�/B+ֺHҒ"O��9�(�q��M�/�6I+~M!�"Op�(B$٣����Aώ��z��"Ol q6��9<tMb%o�!r&��"O��1i��$X�I�YYh��"O�p	T�\�t���&ʴ\eV���"O�OGZ=�h	��4THP��"O�7 G�b��IKw�X#<hM� "O$A����#,@�xa璯^8<p(�"O0�4��9|d|E
�"M��35"O^��Q��x)Ԧ�	����"Oܱ�!�G����rfͨm�T��!"O�I9�'�2��R%�#.���p"O���6kL�R���p*he��"O�<KaD�S3��ꄠ��m���:�"O��C#�A�ne��ؖ�$�{�"O�T�!�7r�>��/۷j���"O���S�Z�&KBE�B`P�!"OJ���G�^lX��ڹ��a��"Oz�Ca�׷�DA��q�@�g"O��UDS=�ju�F�o�"�d"OԴ�W퇤6�N|Hҍ./����"Oz����Z;[F� �q�����"OΡ"f��$� �96���&|5"O�$�eA+Q�J��B��ٲ�"OҜ��EE�m@��mJ���)HB"OP��"!�5:��M�Uk��%���"On�&�%���s��3/`lEh�"Oh�
�Ry!��JY�zD�Y S"O��I!g��B�0�	G$���� "OT��o��$���iP��[#0���"O�ɋ��?+nNTʄ�
�	1f"O��0�0/X��z�E�{�Dkf"O3E�ۅ �4ӧ�Y�%�x���"O��0����R ����.�v"O�1�fӐ|���U��L8XJ�"Oz�	�U0i�e[�İ_ї"O�!؅���lM�pA�� 2}�B"Ol�Y�M4M��Pf�1]L!#Q"O.|��K*n��`[�6"�\��"OB]PO��R�n5#��,w���"O�(	��X��p���F��5�$���"O �:��V�l�9:wkJ.h�.�8c"Otu�q�Q60{Z��#�7vrH�""OL[eO�x�2������]h8m�u"Olh1�&]$��t��L�q\b���"On-� ���� �A�K�5f�I�"O̐*�-��dp:Q��?\�@��'?�DG7Dv]bUM�R���C���%R!�� ��f�B�^��rm�?TE��"2"O��Ԁ�	U��ƍ�*o9�I��"O��!c�F��dx�+Z�����"O� ���8� �t��j�R\�t"O���i8T4�aÏ�l֚��"O%8�&h�H�
T@4��4p�"Ov(@�kG� ��Mkq�>V����V"O���V�T�XD�B��˟a����"O�pKrJ��k���(D����y���;��"��T�B�L�� ��y�6Z�Eqs��=֮�B#f\'�y�-W��]����DlQR�U��y��X�j1>�[V��4.�Qq`:�y�C��Đ,R�#��{������y�P�Ix�(�"�R���B�yN5��ʓ�M�|ָ(	Sj�y��Q:R���u���s��A�b�L��y"ғ`��x���V�W�4d�&	Ƙ�yr �� �6�:i�"O�$��ˌ�ybn�Nv�� � �K���ZuC�?�yB��*`��=�vi� G��ɨq��yRi�6F%��
�ǅ�B��L����yR�ۀ)XL*�L�A��1Y�iѩ�y2 ��(���	T1Ì�q�N��yb�+��- �Iw��8��һ�y�C�[��ɳE�Hk/\,�v��y�l?nNĺw(*^�9�RD�-�y��)Ť\�'MGD�`���^4�y�bV�Vv\h�����D���k_1�yR.��[��,�B	D�\r�T��yrf�7`G�q��`;
x&HH��I��yB��$���i3���*��������yr+���ˆ*+^�s7�P��y� �[䡓t̗���m���B��y�膮�0���J�C<v�Ӑ�_��y��?>~��GA.5;>�@��y��T*�N�(�fЧ43,iY`���y��r�Uh�!�DL)e<�y�AI!s!\ jrE�|�L[Q��/�y���\Q̘`O��AH�� ̖�y��6O�h��⭅�Mp@-�"JR��yJ�(x%�ys�J6V/H��(ҕ�yҠ�=]��)�@*�;}ݨ���E֯�y��[�$+����x��h�϶�y��>�������6#p�q�W�T��yR�ƫ+c����^�{��#��G��y����z'4�� bK�U���qL�y"`�N��RA�J\h@�Q=�y�����(���^����_�y���_�L�w��"��"��y≔�3���Q��M8��	��y2�ќ>������5j�m��#�y�#��;D����W�=X��)�9�y�MS�1���,�/�a�n���y�J[�l�f�砏?)'�MY�`���y��G�� �$ا(rV�ӥ�׊�yb���&m�$ZA�\� �Iه���y��X�ع� U6!�c���y�L�� �˂�,�u�N��y���#�\����eGlX����:�y2A��Nꓨ�d:Z�Z��@��y2�[�}��%��*�0]����eڹ�y���<-��2fnZ�Ud>Ei�����y����p�ک+&�N�xTXQ �-'�y
� ���%��	B��
#.�q{1�7"O��#a 
F��bb�'6z�x[G"O��2�Ϣ%�`��a�h~H��"O�0s��M�b@+� %"}�<�"O�X@!.U>Du���f��b�b�"O.8q�E�h&@�$ωzY6�%"O�L#���\v\��� L�T��"O�I���Ѹ=�x�*��[e@Q�a"O X秇 hd�$�&���0`�}Â"O�H��D�5"~�IB������"O�ڢ,�ms聱2�L�u���3"O��s`n�N(V�j���-j\�w"O}X��moj��D�O�Kp�"O�@r���
'mĔ+P��v=H�� "O�Uxr����٥�D}D��*r"O�d���ŻB�NM(j�h�"OƘ� d�>c�bx[�T$���'"O��(U�
<WYHDx�M�  �8W"O�3J���8`�i�y.Pp"O��Icd�k��	Pf��(T�|飥"O~��핃K�p=�Q
�&,�B�t"OV �V�Þ}J��IP�N���U"O*���\ Y���#e��y��J�"O2�9���#Va�}�I1s��"O~�(1M�*U:0�5�$�
�E"O�2���"s�R�:�j��܉(�"O��A$](Fx�T��c�k�����"O���t�@
j��
dɇ1b�Yh�"O\!`��R/J���)�.�"m����"O��T��p��1m
 ����2"O��I��B�ᶽ�lC��Ecf"O�xC-Os�fêD�4�Qˆ"OR)Q�gM��HQ:��\z~Ř�"O<���+`<^�	2�G�A� �"O�yeH����٩D��v��j "O)hdB[2�J=P$����6�JV"O�A��[-*f�@��9.� Ʌ"OZ�D�;t��\[���$�B���"O�(YuaЦ;�p�ȏ�g�zMڤ"O@���շ]]:m�R烂Q����"O��sF�g��0KF]-�ͺw"O�,����T1'�	��"O�qJRaPoc`4��΄��D��"OL�8u��]���C�	�}��\P�"O4�#b�5Y�lp�Ē�Z�t��3"O*9� c[)>0�ãM	|���"O�Mq �:e��WMK,z_� ��"O�8���	�=2&�I\�
T"�"O�9���J�7�P��AkD-P3���"OƐ�e��'O�4Q�H�?G1 �g"Ol�g��!`T�1�C\�@�'"Ox��C�*.��s'R�1�8(�"O�{Ќ٦LpB�[� ʬ��T�u"O�A�QM��hP"�-X����"O�=3`/X�m�^X����"�A�"O ������aEG�1��E�"O�0�v��d?.̉sg
�=x�X�"O�[��
�"e�&�s�(�"O�iyG'0\J�]���A"Ox��C�&nS�K6�#up���"O�����j���s���b|�x�"O���D��-[�Hh�˚�pH���"O4乢H��O{0�T��F:��"Oz`�b�	6aYP��Ӯ8�Ep�"O� �����n�x��+^�x�`"O�}���ws�m�F��+g`XM�P"O��(w�������S!*R}J�"O֌z6��'3>��k�/�7F�$a7"O�M)EI�\�j`�vDF�Iނ���"OBL���t���x�<�f$� "O*�i689[�(�!q����p"O�Y�%o\쌲5���;��1{ "O
#��K����K�i�ܕ��"O�ڄ��3�q��f�?D#�90#"O�y��'i�$@a�c[�o�5��"O.M�Я 	Jj���p"�
�*D�w"Ov���ӛ'��$�� VQ���2"O�Z��[�R�l�Q�7s�i�R"O*�Y/��̝S�8��qD"O�]20O&9�DM�uc�-R��k�"O���B�E$�H����/?�1�b"O�Q��RIBH;"�B�5�ճ�"O���+��2a� ���Գ9��ܑ�"O<�;�����s�\��F��"O��)AHǕ1r`�8�M�'Px mB�"O��J#E�][թ�-�'m���%"O��ҁع >�����kN")��"O~���j�>\�㫄�<Ne�7"OLHZ�Cy��@��GkC.��Q"O����G)4t�a��B-`�"O4�@�Qau&�@g�^���ʢ"O�d�FnȲ!G`S��B���a�"O��"�g�hHF���B�.(p�"O2X���)S��pq��Ԇ|��D��"Ol�3q�k�d�.N#U��h��"Od@���3{z<�sa�I,<�Vl�%"O:���M�x����W+Ιi�p�yS"Op�;V�P=*�<T6K�#BK���"O��a#��:e�,b���+����q"O�E�� �Gz��ҵP+���U"OP5�+ֲw��3!ݣX��m�"O�aIA���f���(�E^�:tP"O�Ts��Q�"Dv�u�&+~��a"Od�i�bɺ��ҷ���Π:"O�8*aJ�:}ڈ��n74<���0"O�a�bɌ9o/M���kW�=2U"O`1 ��!A���S��$� ��"O�a5�̒9�*p��'P�m3�!�C"O���̛�vM)��_�x+���"OH���,2C.�{G;����b"OHd� Ȳ&������Z�у�"O��k@G"��i��� ����"O���$���� ��GI�\�rmZ�"O�!
��A�d���q��[�"O�Mst�;s�TP��D��,���"O��S%C^/24���^�z1��"O�dbU�P-���j0G��af"O���!�[?T��2�(C�T�x��"Oz����6_��"AF�N���C�"O�Hi�O�A�c��
PM�d�a"O�Yp�
����(��[L?��a�"O�d��ᔙ��5"�m��_�-��"O���c%5��Y6��*e(�	"OJ(@&��(����1�Ŵk����"OH(+�k��ʐ�	���}��qH�"O��s�a��J�)2K��@2��p'"O� f/	�9����J�	:.rm	2"O�� 7�C
oKHЈ�A����"O� ��2���"*�ȉtM�!g�@��w"O�dȂl��f��ӟ^���Ae"O�mX���.��Uk�e\�Ht�P�"Ozթ�i��"�$� 
�Ҥ`�"O���(��k�r�b�早[؜=Y�*O4��4�I-+j*�S�RD��*�'�E����E�EjӃ�+�<��'�*Ƭ����B�KrސT��'��ҕ�^,.����OҲdU��'~�]�s瞉9D���ٶTB=��'�n��팬l�����f�&�>���'f=��s�,�p�戄=!j���'�����W-0�e�"g�^ɎQ�'�rs��!�V���׌W(�1
�'jrm{��S'�*��Y�N�Y�'�52�L��X�p���*Y��}��'6�}3�mJ�V/�Y�U�O@���'��-@)��5�V����J�&���'��U�q��!�|=�CfMpT�+�'��Q�E�D4���MY�X�D��
�'N)��G��j�����S�~�Y
�'y�]:4(��N��)�6���Qφ�
�'�dʲ�Z9*�]J��9��	�'���E	�X�~��!��-+NH�'��wf�U���rCD�V�`]��'1`A�B"��n�<�{&�UeJ���'kTղ0i+�މ�����[�p�x�'7��3���u <X"g��!I��
�'����+��Ed�,��l�:��YJ�'�Zt��N*DP�[7�A�	nn��	�'�&ă�%�g��m�`��0ș�'�����@�a�f���~Ѥ��'����d�4�z�q��N�s��b�'����u�0	�|�@� h��`�'{ DZF	�N{x�7iF	����	�'���W�L�r&ӆ�5cDe��'z��1�l��qʰ��DH..����'��-�&o2C*�U����*��Hi�'Fh�m�
x�\hd�Ϫ���0�"O�X��&b�\ �ȑ=:�v�s"O���F+"���1jT�$V�:"O�ic�JQ�k�Z��q��;��L�"O6,�����<�f ��g͌K��`��'3yi�
�_L� 33 �,`��'�*�3��3w��y V'S�k���'V�;4�ۃIF{�*ưcD<�B�'�n���ٔ#0R�"PJ�'M�$�:�'`�8#!�Ո.�d��̯-z@��'��<2ЮA.���bD��*���h�'2�H��,+*@�{e���ԉ�' ���>nD���ɵAF�
�'c��+��K5��
%<���
�'/����K�ޑC�����1�'�pܻ�_�!Č�)AD�`v��
�'-��� ��7I�rDK�J���'����҂F%�0̚!=yʡK�'7���&n��Y0����Ϲ%tjD��'�ȤZ�`	�iY����p70 �'㞐@��,B���ޔv�D�#�'�D��f�=15��X��3S���'�(�1� =4���G%D:|@��'�*� S�D:B��)i\�.�`�'�h� �+dED��s��4S~���'�RI��CI�.�V��Ɖ����x��� ��0�M&�� �
�'��"O�<��EW�qq�qqc�G� ��Y9C"O�k�*H�I��+A�6�Ae"O	�r�ě*�,���3	� H�s"O��s H#��2���{�½H����,AS�LN��iũzl>��%�M"�dJ�GA#g�qO0����SL�A����8�F�s2�=~ȅB�O<�+�������bpO�.7�������̴9�]ڢ�x.��$h��g��p���P1&˼�)�(�+q\i���.-�H�r@J��b�`<�"a�<)����t����MS���)Ǻg,p��%}HcǤ!Ȱ�ʱ�'L�O£}���$ΆP�eE�pHƝHP�T����Ğ٦�(�4�Me���)8�q�LT;%����$#�w?�*W:g��f�'C�)�L<��/�"m7�]S�
C�iV��2��G.,�4�Sݴ]���	�i��f��e�Ţ��O�����b��w"����Ȟ�i�n lZ�z��,��'X�[¾ �2��;6xȜ`�d�,�>��%L�kl��j*�h`坘F8��:�ቯ �MC��?i����O,>7��?+x�2�ᖈ
Ұ�$�W#
����㟴$��G~R�U��ʨr���_: ��L��(O¨l����j�4�P�$�48�
q��]B��]�pr4�:�M#�|���x�g_	N��f�J_�d��NE�����4`�RĨb�Դ4��I.�OxQ�A��=x�X%R͌�\E4���"ۍ/t�}����|�%�],�ݐ��Y���*b�n6ܕ��4��j�<`�LE��(�!-:�`�DQ��g*�O��Oe�r�$W�p"�*ؐX�nA�2�")sjS����hO?�ĉ�wܒ��Eӓ"g�U�Á�(S�����4K��Ɣ|�O���W�x��	�sܬ@3'f�w�Q &H�L
���Fʊtx�T���lr.6��^�����/�3��5��'C�<�R�p�	�l�:$H�(]�o�"?i���
{ހ�ׁ]/ ��xE��𐪥 -��{AB�1Q#RO�h�伱/Q'#EXt9(O�����'_����5���ɵ���{0LH�H?�7-�Onʓ�?�(Oxb?u+ ��r���އxN$�ӥ:D�TK�4t��@�!N���zRa����ٴ9�6T���׻�M����ħA�5Z�j�MDD cGS;����=��X�����(ܲb�P�A1�O�ڱ�vKz>Ţ3a�4�0�;Q@ߦR���k4ғy¤E���R�b�M)�ɟ1Qr($��,V�;3>$6�5,��a
"��Uè��R����5�+4U�H�.��t�	ܟljٴ�?����yBj��:����N�e���f(_ҟ�?�|�K<�F����ఁހZ�pm�4��g8�	ݴ=C�6�i
xu
wĔ�I2��R���P�@j�'�R�ۢ�v���<�'�zL<���uz�u
V�M�Sg~�ڴ��;��)�!_�pZ�y'�3yd�x 2�Z�'���8����F�9= ���s�^�$6͑�f����I�A��b4fE� 3S��"��åU*����hi�E�3�d˂,@1u9���7�i'x����Z���<%?q��M�&�;E"yXW�L�i�
�-s�<�GU->$�MR��^�)��ӓ.�y?1I>�p�i�T#}*[w���� �ց`�a+D��>�~5���(��9lO��9`�  �   ;   Ĵ���	��ZP�viė:&���3��H��R�
O�ظ2�x�I[#�x3۴|f�v�J=|L��gJ�'��l� j'�6-�轢ٴ.q�$0��\�I�F�p�� I@��4��X����f$?�!�r#<) �d��&�R�~��� p�<
'��`�^�xQ��A�Μ��'?����6}6-L}�D��$�A����36�̣ln*�c�CN^y�C�ODcs�ʎ��9O4�y 
�/��cEI�6\��L���X����b�8��D�`�葰1����'H$�n��$iq��%F��P���q�'�dS�	�lu�'�����K �R�	�7
�j�h�'B,FxBDH�'I���vjƓ4�T����ܥ/I���O5Ku"<)pI�>C䆚�J�PMV�M���/�H��OT�R������'s<!��m:����)�*rY�8i۴;WH"<	s5�Fa�*�Ɏ(75Z� +|�;qh�Z�>��#<1� ?� �B����P�¦.x2�Kc��Yy2��~�'���?I��ؗ	h���'��MY|[Sj�?t"<�e8�2����н)����B�R�]v���s�C1O<� ��$����~B���p�� 7|��ukƐ���lT"#<�m5�k(:�R�^6V��-AfՈs��x��o��X�K���i��mGDq�����|y�@�3z���*��$�B�<a��"T��P�<�2k�3Uo�O�2��>R��#%
�f�>I�s\�l���I�-C��Qe�:2z���P�:Y�I�"7D���'K
   �a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  '  �  
'  �.  B5  �;  �A  H  aN  �T  �Z  >a  �g  �m  t  Iz  �   `� u�	����Zv)C�'ll\�0Dz+⟈mDԤ�57���DB�������$)�9�R��<5G D�Eg�  !Xm�@�߶>���VƐ=-�I��~)�U2�'Wꊠ���(I��A��{�>��`��H�t)�#GJ��x�R�<2�¶^5���Q���������,���0c�Ш�aA�H���EbN�R]e�pJ�8Q���5 ���"J�9pX�q�4gn�<����?!���?a�K����_#>�xؐw)M;9
�����?�1�i�*7��<���hܘ�'�?��v���aD��[2�%��_c��X����?S��Ɉ*48!�	�fl�l�p��A7�̠$�.r�F� A(�,q(@����<� d��1q������℅�F�g}4O�㟬���R*-��'��8�Q�B�s%���Pl@hܼ����?9��?���?i��?�)�,�ݾ �j�[4?S0���%C�=m� �d��a �4(���i�����nZ��M���i��fg֌
f	�E��+ZŌ#=!v��s�O������9Ahd "%.��#0�,���[Q���EG�u��� �i��7��ԦY�Ӯ�RdK:*��X@f�z�Px�E�I�lQ\{r�t����P�[�.�s����h���I�Dk�7���޴�z욁�X�E΄��r�ZRːH�𢅮)���5C�����GyӸ�lڶ ��9s��%{Ӳ���D�<(tM�gힲE>�Lˣ.�:yע	=��i+pcϰ{�I�ߴ��/o�L�X�g���Y���� cvO���`�ϒ�d��CĪO3d�܈�iZ�dz��N�`xv�a���AR���'�O��aNIa�+r��R�
���g[��� �f
����شj����O�4�;Ć ���@+"��l$����ވF��i� D��'!�D�h��p1�`�V�#�25�!�O�W� U@�G�0�H�֯��!�$I%Yn\�PJ%M$v�&�O ,m!��JנxXҁZ�,��cl�:=!�$�0@V
�bağ^���yeL24ў r��/�NothP��'u�(y���%���"�X ��-���#�Z $~�ȓY\��CHĨ}�x1� �M�r����=�u�8l�]cco�b,��ȓo�$�D�;��\��?l��d��@���:�遌|w�!g��72��	b�#<E���שrm$<��%�"l�Lp��ږQ�!�$ۢh�n�iUÍG��\��NLA�!���#�QN+���5�F#�!�V�=��M"`�A�\ 8�,��!�d�3H"�B(�_�P�	�`R'�!�dBn&�C�Kg�PR�	C�)`�ɑ2˺��ĉ�s�(ib����0R�y�B	��js!��(&��x�Ņ4���x�悚 !�D� V�����=B�&�CE�	!�$ݘW����I�j��8C��܇/!��.q7��i0痍i���A�����yB��>d��6��O��N��B�y����j�c5��$�O�H���OL���OF�p0��O�˓�y��Z�uÑG͙t����A��0<�BnU��h�	6mz�		��M+���N���В�W���D)}�2�'x6��O���IB�L��xd6R$1X�%�<�4;��O�d�ɉ-��̣#�OhQj��ܓOcZ�QSD�2yx8�qd��*��|J��'�L�	<:�dRQ�I 1x�������!�����O�˓�Γ�y��7���6��(e�M������$�`g�
�{��	S/m�>�2��ڝA��q�q$�K�	%� =ʗ��S.P����%BU6 ���
 6`��K�� ��ٟ�%?a�|����O�����Ul�-� ��k�����	�q����ʣj1��ň^EF�?)���A(|��@пD�hEz@��>X�H�� ���3ʓW�����/�(*f�$�<0���/� �)y�bܲӈ� <��z�\j�̢~m�Y#sL�3�����yZ؋q��cr�$Ӓ�ŌBv����&0���Gݝ.�	��^:E�H�Ɠh,`�#q�&Xk�Qņ�.;-n��G���<��q���]Z�L�p�T>]EZ��D��z<��#p��)��wL$i�ā�}�ֽ���'p�@�"˲Lۀ�	b�"����B����� �ز�R����e˹v⁇ȓ���+0�ʉGR䢑\ ;�,�%�Y�4���� ����N�;Bt�
&�O�l�L��w�@��?�,O���O�����,�\���e�.�.�P��!D��� Y��&����(1���ټA'f<�}5�l�ab ����J��Fd\1pq��!XO(�"��N�/�3�BN ��On1�`�'��u�"}?8����m��2!*�D�O��(h�)���'u��1�D(z�����O�yH�f�aI�!��xq�T�'p��O.���4�?I����9H�b������Ԉ�7n�d`JF	��.g��'���r���t��ɣ�@Ը2���T>U�O�|,�@*�5�m��K@H�O�JWO�(�\�h�֖\w��}J4�U��!��F�R��h�F�e~�鍢�?���h� ���0��88�kR�N�>C�<-�iʷ ��g���,*Pq�����h��d�Ԧ�St��&���4�g#j����<�wS*P��'"�'��I�H&\ӣ��	MӼ Z�a�z�>�d���b=���P~���d
�K�d�O���O��s���0�@1I4@�
$c(,��_$7Vx+�L��1��܊rL�~�UFI���F��,$��p2��$�?�´i��Dp��Y���	�N��8����;*a�����.ٔ'�ў�Gx�)�>R'���U^��`J���$cӞ���Ozqn��(��ꟸ�O��%#�)�-9�6�kF�ܰ6#4�b�ሄ*�6�O*�d�Oʓ��Id>���_���1yÊ��&���'�;���"�Ͱu�Co�@�FrJe�5��+�.8iꁣ�"`#lR-�=r��ˇ����_�+W� ����(O�E�D�E�$�1U�~ĉ�B!j�b�'�6M�O�ʓ�?i,O��'[N�]#iL��Pe9�,G$R�%�l����}R@& 9����ނC��������M�����?YC���y�5F�F��׍ _���� B��y�kҙ���$��5mzy9׈ ��y	�T�P�Aci�!�4��Ù)�yb��~���2�
�;�L�����yR�\�k��ѴǏ��(Qk�I"�yr��(Et��� �={�(0����hO������&!�,PmV�\���Kp ]�8�C�I�
���cAL�v�j��v�گ&�C�I)ee��K��0@`~-Z�� o��B�ɣ>��рh#���7-E�B䉆CVZy�'덡m�,�`�ҵ:�B��;,v20��\9~U�aQ/us���ܬ�"~� �G��t�ڳ���:ǔ��d��yj��
��c�� 2 �c�� �y�b��c/���A� �}�i�A@ۥ�y2G	�&�����jM�
Q�U3��B�yr�ТiF����YkP��#D��0�yR�I�^���XP�_�c&*4������
�|R̀*��B	1Ea��flW��y�%Q���Q���&��0��bF�yb�_��b2���Q�.��e��ybKq�,x�5>�`ti��V��y��Η,D`Cf�$n�n-�%f����>1҉Nm?Q�%�\u��e�)]�ڡ: O�_�<��(�,"�6*�I��X�6ِ&(�C�<��R�#E*a� !�䀐�<y$)�CO�� �K�� �2�+�ov�<)A��;,4�U�Ӝ+B8<c ��r�<�1ǉ� 4E ��A�"�0�Vr�'6�1����>jT���Pe����J�P!����a��F{��rn���!����!*��X:4Xzx�,Λ"�!��t����K��>���t*^�!�$�o#��6��=܊,c��D~�!�ą/.�X�ѥ⏬-�Na0CF��&2dZ��O?�J�"x_$�jĤ�)Wԥ  ��T�<)�m�E��ҖL�Kl���k�M�<	4�VH�8�2��jT�1H�H�G�<���&6Y^Lk�� ly���� �]�<	7�S�|���pEWc�h� �\�<�F͗�%dH��B	}�̸�Uy2l���p>	��p�9����&�^����6!�� ��B�HƲh�:=�-��N$�9""O`1@cH��'K��D�E	�B��1"O�y{gǁ�3�܀��+����(�"O<�c��ҡ<Tu!@M�='��"�'� ��';ƘpP���f�{V�T�}�
�'vt�ڐ��:c�v(���S��)�'a$���G6� �vK�-I?+�%D�z@�Z>�ȍ#%n��O����g1D�T�EC#��I��E؇eq��"6f$D��;�ۻDx8c�	\�����.�D�AG��gZ��T����s�M��ݝ�y���?L&�m��[�'��)I��y�	��V��-���K��B�"�ybMŶQ�YĄ���}؆$��yRV)��ǈJ"y�Y�����y���GG���`��0�~��TeǑ�?��W�����Kr/�0d�"���a�h��o���y�"Z�I%���dC�
 R�)q% ��yb�
�t̠�)��u/��p!���y���
3J2h	�)��v��o�4�y�-Ղg�e2���^���헣�yR����l�O��[K��"�����D؃*��|B��%�:��d�CH,�[ƥ�y�HE1��J�2D���v�ʷ�yb�Xb���qdű7��M��&3�y2�/t�0-�q��4�tm�����yҧ�n�0��B�[� ��H�������>	sdWu?���0`�i��;vtҀOB}�<Iw�F�F�81ƍ�?P��h��z�<�TO�G�ޡ�2�Ć6��E��s�<�cD  ���h��
�T����j�<�r��5����LǔVT�Al�<��h�>P���@�i�n�1��L�'��š���L2R�D�Q㘜A�0�[�o'!�)Nנ��u�W�`Z,"�cҥr!�Ow�d�F�*&xǌ�9$!�$T=Sz�+�8-�����(_:!�D#�������8���zTA��R/!�J"2����� ޲�ˑ�Ͻ�R��'�O?i �PSK��3�h��q���@�H�g�<�nW:DL�	��:3�R�x I�b�<	�ǩe'��G!�8>f~+0�Z�<�VI̸n�������5K����ΌR�<�5 Ҕ!��3AW�8�bl�vʟP�<!T�Sd;p��%FhqRĪ�Qy2N�(�p>�!� �c�:��e%R�>v>�a2ɎQ�<Q'���P��'��s~�ę���L�<���� �§	kn$����L�<��*�Hݰ�� w��R�%$D�X��ł>+D��*��%-|�uB,�O�E��O�9��-Z�Vİ�ȖM��Y=�y�"O�]&�Է|��Hp@4�!c"OV�����A��ʕ�k��؀�"OB�ʢ�<M�A�O01�hPs"O
,�P�X�.�NUCb�z4���D"O�mqe#Y]�d� ��@�iE�DB��	����~27@X0e�ؠ��A�O�\���g�C�<�ǃD�2$IWS/�<Q�"l�g�<A��ןo|92򍐑K��8���}�<���ϦQ=��Q�
$����+�a�<���9̢�iˆ+V!2e$�`�<��oR!Q���'�Ļ>��Y�fEß���j&�S�OI4��Rep�,ЧO�Bc�M�4"OX`�,B�B��<+& (�)u"O� �XG��$��x3n@:a�.q:�"O��`2���ex�J=G|��"Op�rW�L>S�����;4�Р�4"O�hr�n�Q�΍(q*�� x��V�d��M;�Obu 2�ͳ
h~Y��IB��c�"O.pr�Io�z�#���%����Q"O����&	)Wb���&H�H�q�"O� �X�0�썒��[��Y�"O�UM���+͊(��T���Nx��e��"�n
���ZR/ĿW����3H!D�)�%-b%bC���dp��`�#D����⑓��C0�IU��wA>D�q�O�yz��CE�WmB� �?D��{r�6bL��$� �3�F�M=D����Ϛ ]�.,� .�
o��E=ړ
�D����`>�T! 9?Z(Бp���yG+V�I;'#��9�M�l��yBÚ5�|4�E��(]�`��DT��yR �*JB����[3"��Nޒ�y�"g��裌��H g����y�R�d2� jE%�^`r�ܑ�?��l�]������&��"bi��Bu�ޭ?۠�:��'D�l!m;/K<-�bG'[�L���'(D���HO��
ࣧ������*D�p�#��'h���D�BF�1@6�3D���-�d��ɳ.T8*��]��`0D��X�G�$E�(8c�7/r>d���<Y�Sb8���ч9I���ф9 ~���)D�(���-��Qr�9�Z���(D�(�.E.8�2��mQ�xeN��4D�$�2.W�I�,9����H)3o4D�4��j���`H���5Ԅq�g3�Oz�p��O��rԤ56�����JQ�N`x�A"Od�0�����M���_{��ɀ"Od	yV/�NH�a�M���W"O����>1���"`���""O����(!f�Y,1�Q�w
̎�y��Ξq18e(B�����d�&�hO�CD���:�h$�E�{�V���W /��B�	�\>xܪvdN�l&K̅b�V��1"O�����b�*0�0`ȶ&�8Di"O��Q��_���$�P��t"O(P�7EΤ"$9(���L�9�"O��	��0g�$8��5h@�d�'�0������Vk��P���
�2��� h<��x�]�ޅ&�1��C@���ȓ^f�P8e�bD��R�Go	.���QH�)k��L�'<�è$f|��ȓSX��� �X4X�B�x��ZC"��gt��4��4�l�q$dԜ	)J��'�.I�e��@@��68��X��W&���ȓt�Jp`G�:zG�YCc�@�oʝ�ȓP%������+'9����-�P�
E�ȓ=��,�!*F5��4�U�G8m�=��X.�8q�^�%�Z�2�"N	c�<	����}��	8
X��OR>�bJ�5��C� ,0��5l۬ļu�� ?w�*C�	�+XZ����:(�H�'�1Xt�B�	#Plj�j��G�Q0H�B`�ж|�B䉩�D�:�G_�&}ZQ��a�a�hB�cU�E1F��2P:��BV�=�)�j�OD�[Ƃ�4� ��tB��;�@I��'ۂqj2�ӬL�h�B�1�v�(�'�Hl"1�%I�@{���}�J�x��� �Ð�V�f�賓�*Yܪໂ"O� ���6j�F�� F�@L�t"ODL2w���z��p!N�C��%i��'x�R���ӡ��\C�ȇ6~�$L�I�+C�|��<E�	:�I�Aߢ�L�4�^̆ȓYҘy��!�#��؃�R�dԅȓVi��ע�$m�|K���;�&I�ȓ��zC�G�
A&�q��O�q�*��ȓK���΃6���KL,��'�$��W��*r�b���Qe��\��ȓ������S������ۥ�꜄�dC�y	���+��l
3��%򪑄�O\Ea�i`OV�26���i�ȓ�Ф���R�<��Z�+��p���	�m~��ɶR���H;7�Y��@�7M:C�	 v^�� %P"���b���<C�	*+��m�F�פ�����B�\�|B�		�;�T	.p�Ѐw
xdB剷=ex��w���%W��2��V�@�!�$[��=���XT�2`��_�ўаt/)�5�~�xR�e�px[5$W?v�L�ȓ]�PP��{lB�!�M\�uT1��9?Sq�j�E�Fg�
>ε���Nl!�����	�$��&���ȓ�2��%B&��m(�չ\5N-��!�4R#)��C��ř���3=8|T���Jm�"<E��CL8�S3�ZMc&f�rh2"O� Iwb�bT�A���s�!Sb"O���⏿E�u�r��7���E"O�s��4 _��)֋��E�4�t"O�Y�B�%������D�OPp�F�ޠU�����/<�z@!�f���'{��n�,��'z��z���B������� 8#� ѻ,O`���OL�䐠G����;=�2��	'@������!B�D`���L��I�]W��">���F?�TI��+U$ �j2�j�U*ld�eb�rj�%T1r�S��à�(���jD�$�Oc>��pj� �s������V,�<!�hp[�e8;�[�8�H���0��D�j�@%�#�"4��#%兪T�剟8	&\��ԟ0�'c��П4�I�!�<�Մ�4���: �g����ɷu"0\9 �~q `ī`�"�	!��u�O��� DCO=9�(��D�Ν�`�'d*�@L�!|���P�(L,؈ )�eB���x�}�`=&�(����%*p����<Y�����	M~J~*�O�sTAM8 �dQ���jޠ�E"O&E��Ǆ�T5"0Q�*�i��]!����ȟ�`�d�}،�ʹ-�lK��OL���OF��C��(<��d�OL�d�O`�)�O&{`B�k`�C�Ş������Q�1Oem9fiZ|j@F\�*;���O�b���G�Kf��R�D��VQ�5`�[$G萰� ��H].c��&Yt�'x�x�)6,i~��G�.��]zGLZ)-"|e��D��dX�Rz2�'�ў�� sщ��T��)�+c�)�� %���fM�'A;�A��]�S>��I��HO���O�ʓV�8"�8OȲh�� �媀����7y�ڀs���?����?Q���?9�����F�����')��DU�	�N�-���8Aa��*�haGC�
6��&#�H�'D8i�酞A��]!�l�1g=tE ga�A�Qiۇ0����E�@x��q���O��Ñ�'S h�wd�����F�	fE�yzD�'vў�E|�����[�:FJ'oH�o<R�ȓKyL��dJԒV�����Q�T2Bx�'��6M�O2�\�9��N��i���4�\JЊ����_&��B�_-�?a@���?q��?1Q�2ۦ0��U�gH8��|�Cn^�w$T����G�x��1G�[H�')bH���Rf����Y�C��8�*tH�	YoS�M8 �	�7�4���ORc>��F��d��ط�̝US�(�b&�<�[��!a�ϔ}yx����l&q��I��d�-c�F�C��1xI��	�H9[��O�4ِ�9���?�	�K��v=R-��YvJ�$�C��&��c�p�uy#�;�PC�I?I�8��p��l`�E$	�S��B�)� (������huRb
�z0��B"OȌB���B��юV�0���
�"O���m��T�A-�)�LtR �Q�O^�}��W��p�b
n�13��+�䑆ȓHg�%�F�X�-6N���7�
@�ȓc�n�A!�N�1D�Yۡ��N�F��ȓ`y��P�LyI6i`ceٱeT��ȓ!��kPck�X���/)Ϫ��ȓo.R���:p��+%l�6.p���&>����$ۊe��	I��3ΰmƦ��C��G�=��*��L�x0��1|�fC�	<�q���ɻ4��ك�6YbC��'e�L�ȀGH&3Ȫ�(���u�VC�I�7�ȳ�A�A�0��g����	Z�P�'N28�N�
f�@�n@�r��U��i�'n�d��'w��'��h�u���~?�iK ���a��7-��uw�E:G��pW-_�8�����m��O����fekA��-�p��)I0��*���E����0���(6��  ���On�d-擔6��[Hsj�󷥍�PI��0?�p�-���R	��
.ȵ�V�U@x�H)O��J  ��m�-��N�?a����^���I�����|�'������� ������JMm��	U�'�ў����ʄn��z��X�?�l�!�
:�Ɍ>�Oxb?�1��6��	{c�@4xЊ7M;?��OԂǒ>��y�M�x�0T�T�ؔY��$�$��Lk��8�O���@�,}�� 񩄒N583-�I���g�ER�B(K���'��>牎^D@��6��?Rɒ�[$DT,����U�+}�h+}�������i�h�@
�m��\1^�a�F:Dh�aK$��ɍr�Т� c֤j��q���J҇�]�?Q!��S��@��r3�_��,���L�%���p	TⓂ��:$��`��?5�"���CV��r`����XSv����~�$	���|�fL�Z���?��n?'�)S��JV�͑�a�7M�d�'��H��O��B��i�8�z���պX�r�yrc�_�mV[?t�MS~ʟ��T������8팯[c�1�ԡ�>k2ie؟�أ���]�������,P��5D�4��>`����Ĉ)���e�4ғ��'�"�'�Paɳg�~�ap��X)/�	��Ʊ>�K>1��T?��\M/�4Ys��/ZHX�
�M�y"b"F(�(Q��|{��Yw����y��Q��Ь1b�������V�yR��0
����!���Zgm^��y����X�v�֕��`6�U��y��?dZxU�0JM��Ys0���y�O�!ҹ�w�>J��5�FN��y�Bߙ�J�[fF0,�,bvl��y2�� �FAqf��?W&^�yBM9�y��fL ��g�RI��P�fA��y�n�r`���XEN���!�U��yB!��$�����-g����f؝�y�-�:��0�&��2	�6iy�����'n�}¦l�-q:����m�!r���"b֎��7a����̀>њ��͎�X��@�
��%�4��Q,�?�48��b*�8��Qˍ$,�jH�0ʁ�!0N12L�!?���b�L>`���h"�7gp����
'*���fiɓ϶���6$^lq�1�'T�j�O��&Ď��*p�c£
�ؘa�IBx�X� Ϥn��Y`�ƥC�Ĉ�'.D����a��L����FR�ZLK��*D��8�ˌgY��2A��(�l���&D�0HrKM,>� �����Ufh�A:D���-�=NZ���Al8}"�6D��A6���zV��x��A5D�X�a�'7#��;Gb 6���HT�1D�T��,˕1�VP�H�U�r��u�-D��{���Q"��J��c.Bգwb*D�`XDA�)i@�r�CU�HWڰЫ&D�8�#-�,qF,���2 c��d�#D�P���ѮVxz��Q.(d�v��+#D�� �d���K�?�r��O�9���"O�1*�c��z�����i���e"O�0q�/��Haܵ�W"z,Y�"O���ōT|�����v,�1{#"OV�K��.ঔ�vA�;����"O`HЊP�\���h@o�!o�&��"O��i�˲8�EKȗ'���g"OT����>Q�M���M8p�d�y'"O �P1��� *���.,-:x1C"O����D�n�x @��Q"O�(��$�1}-N0DŒ�N�aQ"OL�`b�Q�q���S:Z-���U"O�(��\"��� GŮ/ (�"Ox(P��I�2�QO�&2�T� "OЌ�E,R+ e�M�;�*�"O��з=l�3�^�v�Y1�"O:� ���0��V�]-O�0�h�"O,�)�j]�s>a��	33�"O��Ħ�ck"M�'X�c͎h�s"O>�S0-N|>����׆�b�"Ov�h5��0s�����0�J��A"O��9�b"+UJa�����a"O~����&��!���A����"O���3!}Luk�	̀��]C�"OHa�@Í�%]�պ��\�m7T��"O�Y�if~�u�'�V��"O.AS
��O+(� f╖��ڑ"O�E�*讁(C�W$+O�"O���P�ӧh����HQ�(�c"O4͘�JW>�<�k��/�x�"O�Q���k�8hKed�lG���U"O��B���NV �A�BJ�J��ܑ�"Op��`c�$����ʠS���*a"O`s�V�p�T���W?{����S"O`���# ���h"�t���"O2��U�R���0c�� D����4"O�ѱ��8&^`�"��>m"�ݨ�"Oz��cOC�*�$ɣR�V�IT+w"O�=�@CY8@��O
�)���a"O�l ���[�(Ĺa㛃V�z�#"On}�A�C�R��$A�4�T"OX�VF��)6��86bׁ_p�yC"O����%�GY{��X�eD`M�5"OzH1�ㅅ��A�" P�q�-Q"Op(s��2;j4��W,��G��K�"O]rRo� ^j��&��CӾy�"O�Pq�b�&E��@
!'}
"Opa����{��8�&k��^4� 8�"O�y2Vㄺ���E�?��J�"O�ev�_�d[49:���dĳ0"OV���D	)C���eش&�x��"O"�3� T�/V�C�ot ��"Od@c�I'C�	LY`��"O�D�$@B��y�e�D�ȫ�"OO�դH� ն��gA��y�Hʐ%������C���Lkf$��y2F̛X5�)1g۲|��ı�$�y�!�*n�0�Q�b�+�|�a.�+�y$��H�~YA��n\��sH��y��/}Π�Hs��b=�t"$ۚ�yrl�.�dD�QIюU5lK�+A��yR�7
�h�b���L�,��'%��y�Ws�~��&L����7����ybH�W�N�2��_B������y
� ��P2 �Yk�%���ƈt�~���"Oލ���'Y�Bq�2�¡Q#���"ON��	ڵ7��Q��Fdaː"O|�3l˰A��PS�ζ:i�)"OVѪ5��%,iR%q�nT�tc���u"O���Z!(�� p�+�%��)�"ON�R�e��jg�X�
��V�`l{�"Oxq�J�g�@���5��Eڐ"O�$��>���ףĭ$�b�H7"O��* MF�G�u�5h�o����C"O���#�P~ ,�(4�ͮ�HT�"O�T����-��,�t��O��mE"OZ����ւU1D嫒cU�t�$�s"O^����1$��y��A~�U�"O���g�A���{��
�{F��"O�������H3a��"CV000"O�U2�^�>�B�Ceꑑ\2�x#"O����P?lq:5��O6��"O,�����(�J�RL�5Z/�X��"O�hR󀑴C\~,�jߪk���@"O�չ�f� Bh`��)��7�LԘf"OvK��&-v�:���9�B�8�"O��'��OU\��ՏFK�483�"OpL"��)+$T�z��:@��z%"O:���$B1eAZ��6*�p�<�[�"O�T�t��|t`4I1�Ƚqˮۂ"O�\Z�\9CA�YHUO,Wa
%3�"O����ރXb �@.�(#�(�"O����GZ�v�X�C�Q-Ӛ )a"O��O1�>Pr���W��)"O&ؚ�ƋZ������3|�p���"Ol�A�k՜W��G�)*��â"O�a���rWT@T�&�v%�v"Ov,���a��D�o4!A"O�Ɂ����Qj�
wރ>C�-��"O8�)g��*\%�
@]:���"O���"NF�gj88��Z�k�ȩ�"O��BC���a��8@��* ���f"O����n�n��'��Z����"O��!��h�T1�G��W�д �"O�l���B�Y�<-zD;��	C�"Ovy�B�X6&	�5��#�P���"Ot�#��U��� x�̯F�-�v"O�`���G�.!0@��8'~�k�"O��n'��tcl�)s��q!c"O�h������R��ǻBB*��3"O�D��Eՙ;L�X{egՉ)4x��"O���'��Z�2�[�^�=��Cb"O�$qC->A�5�C�(F��p�"O�����2*H��$�K6u�t�K�"O�M��EQ�q�5�2ۜl(�*O��'邉=C����b�W\+
�'Dv�r�E���gI�!xF��'�vu�q�ջ�.�" !�����'�F=j�M�-W�Q���ދh��j�'�����=u=�q�ʼft���'��% EQ�ڍ��mޛV��Y�'�����@�_�fe	��P3TZ�-��'˖C�
�O,���V��B��C
�'uR�ӂ��'&��aN'�r����01펩Z���h�Ϝ[
�'!^�ze*�.
\�BqnZ�\n�@
�'��t� t��|����&o�Y	�'HD��V��?fLm9S��F���� @�`�])^2�e�d�c�"O�ȑ%�3�L��PТy�F��"O�<�t�L�a�pdM�|-:H�"Oz$�bO���C���<��B"O��p&�=��RTEʓy�T�q"Of<�b↑4�"���M]���	S�"O(-1��3$Xm���q˂��"O�d�-���3�ǴJT>Hh�"O������3*��b�l�wD:�`�"O���4Hú0��I!�K7�[�"O܌#0�Ӓ�(P�@j݊=�p4:�"O� �b��`>T�J-8@���"O��9e��5�Af/N�W*0q��"Ol!�CM�d�1�/	�D��s"O�1���V�AmF,���()�x���"OnU��)���i�(��M�"��"OH�C)�-Q�N�'R�<I�"O�%�W�� 0H��r�&�\�"ODIٔK�m0��Ci�<Y�v��"O��V���	�vD�3�ˢ9���p"O�t ���+}�R�S�~�,��a"O8�Q�˥@�2a٦�FH�\���"O�8
��$*{2s!�^1d�h�H�"O��y$��
3��*���/{`]p"O�+�
SUt��m�T"O�!v)V�T��y�3�[0-_* �f"Od��7���P6>0��Ù�;��)A�"O��Q�X�(ȅ��	YΜ�:�"O8x�bW [����@-��,�C"O�m�u`�+t�@�MN�fL"ZR"Od�wM�-ilts���X7J�"O�p����n��ِ5mT��H�A"O\�j�BU5��yUꎗ8�h�"O��Xu`�7 �|R��4m�ѩ"O�@{V�U�"��"Ā���Ѷ"O�!6mַ��Q��%�<��"OP(��_g8�(��b:�d�C"OBm���R=w%���1BE*z2:TS�"Op�aC&P�>�"�hG���x�+�"O���0��2"(��2W���.pPI�Q"O��R�� W��q�S���h_d��"O�p"w
,{�6	��ϯ,Zp�:d"OT4*���Z�ֱ0�%�}Qp=��"Od�(�+�M_ �q$F�>���c"O8ݩ� �%q(W-I���q����yr̦V�U�Lď.���k�G�h�<��P��j=R�.�C4�x��.�i�<y�	Ȓ�\9ȥG��AP�Hq�<	u��*rK��p�`ƪӒxy�-�o�<��R����'�V�h(��ۂ��n�<y1`�g@-�B�<�L ���h�<ё���3U�@��J+���t�f�<	�H(p����X�<� �1&��y�<�'�2
L `�ڢTa)���a�<��JX�����ݜ*I�"�_�<�J�li��pbAN��QdI_�<�#.sZ�a�⠘���XQ�Q[ܓy�Ԭ�ЬE8�����'�,�%��i�삌i�P1%��6x0��:$'/D�@�b�:2j�ܑ�ئZ�Z}Q�!D��`�o�Tx�a�G����*O�l�F�O�{�YPB�� �x}��"O.�q `�0ā�,@���2"O����G��С% مq��`""O���t+�v������| �*���y
� 0�@fH� Le1�Ŝt�B��t"Op��%�d�"���%֭tߠ:"O��X�ǔ��h����#!�I��"O��pB�� E�ڔcD������E"OX=��M��/ڶ���*�	J�q2"O0-(u���R"��8
��2���Q�"O8���M�g�.��ЃZ��) s"O�p�'���?���b�CP7la�I�!"O�}C���+,I��HJ�xE<}��"O����c��|;�Ua�����"O*@��oX�L��\�.�&l�ԍ9"O�y� iƘpQ\�"� 2T��=+�"O�yzF!�	G�t$�W�� ����"O�iچ��|�\�Y�BJ�r��Ȱ"O ٗ �%m#�8�@C/5l�L�X�<1��R*u�豃޸^>N���c�\�<2LR�G4���
�9�4M�t��`�<צ�!?�\i�"� �<�qS�
G�<iǠ�_6�5,���2���c� B�	�%X�eҷ��;_� bu�E?B�d�p ���4.�b�X<'0PB�ɸT�
@:r�˦q�L���,.gA�C�	�o%HX��}�p(@�tŘr�'*l�0glI:Y�1Rc��OުT�'G��#UL°ilf ��JNL!X�'�<�K��aϖ)�5�ȸG��9[	�'G0���&zdd��M;L4�a�'VF��Deڴvqx���H,B�T4��'�"�)uG�� ���cW0>!8�'�-c�/�k.e룁�"����'\���Ǉ�5c7�@�F֞XR�*�'��8z��X[tU�h�1:���'�@�G�?9(�W�ܜ7�!	�'>���V���r�6qj���1���8�'�X�aR般Q�Z��рNP萫�'�\��E;ޖr'�9ox�0��'{<y�e&��T Y�HW�d�ʼ 	�'�N�cc�m����sǎ�nV�Y�'���a`��J�����Yz���'rT]��&X<����	�O$��	�'�z���L�}},��-_ L�Q��'���%��z��a����B)�|��'��K�E�l�`5�`%)�B���'G^xU`;�l3&^2w���q�'E�D�"�$CH���,m��'^.-h$cW�^�~)��d�4A�0��'Z��D�4�� }r���
�'A�8��h��J��f��o�Ȩb
�'��r�N^�)�`X�AB{�(��'B�Y��'�-u�8	��쇷p�^���'��t(�hI�65
�������
�'֪�r^� j��S�l�����'(��;��D���]x��1^��}y�'��t�d,��A��AcF�\�����'ͦ}��
Ì���!c�=Pzyc�'O8��ߛaU~��E犢is��'�|1SM+-K���䣊�DA���ȓv��z���1yǰ��`�B<h�lЇ�� dkTY3p�`L1N�Af����a;Q�БTH1�u�͊s�D��s�9�6I��Ĳr@�-C�6���W�����À-;�j)*�X&'�T ��E�re�p, 5'a��I�#j@���^+l�3`Q��-a�.��{��͆�S�? �D����SH��Г�T'A�|��"ODt�m����h����\���b"O�QQ�aוe�ư�˞&~��s�"O�h�1�No�p,X�#�
#�tX�"O.���h@^L5xc�.=���*`"O�IBFb�4DL�yv���tY�5"O�ly��/��Ԩ��4��"O���W.9b�2��L�=�D��b"O i��b�#' �1.@�e��-�"Oހ�@��J|z�K'l�gN����"OZ!q�.V4;�<�"cbTa�F���"O��ѱ@�8$��,�GE�X��m�g"O m�6jI<I��1۰aF!EW�bP"O���dc�v�� ��02��1"O����6 �������$*�2"O��ց�M�ʁ	�̓(#w�p�"O4a��GU!e[��c텦D�|0�"Oܽ�b]�yC61�`e�
a���W"O�!�M�y�(�if�D�J4��"O҄�3b	��D4@b��Q )c"O�C4욃f�4���I�J��"O��2��ɹ{�ZM���*jR�# "O��#s�^�tRRX;DK%bj4I"OB��1BU��Pacr��IM�@e"Oj9�*ީ'za���q��Xr"O�<)Æ �,��	��]6E_�p��"O^X�'�P4+�YABL|���"O
X�t�%3�-qUA�Eʴ�P0"O�Ը�m^76�L��'V���8�"O�$Ƒ�2�z��� �K>��3"OP�;(XXH4[�E�
pj��"O.�s5��	��)���T��1#�"O�I�H�U="9���/ߴ�s�"Od�#Bd/�:]��0<���b"O��0G!��LE�|�ŇϥP0h�kt"Ol�� �ȍ��(��d�!	7X��U"O�US��_V켹V�MR����"O8Q+l��:xX��"�$��v"O���7ꂚ��1�D�P�J}�8p�"O@�W�S�<����%6�4��"Ot�H�	 V�d�H ��9bf"O �B��⺵�眃�J��3"O�P0��t�U�U%�2!�֘��"O��)ňr,$+��7P�H�7"O>9c�dw�~-qAj?Q"ୢ�"Oh�r��؆h�tE+�(I�pau"Oez��7N�#T�Y��`�3"O,�i4��1.JQA�M+I�b�� "O"����Y��@K��	�e�na�3"O�xJ�2R�ah5�
!k
�E�g"O�t�AdKj�t��왕t(X��"O �2	B�~*�)I"E��]b��pU"O�C�F]&9�j욲ˋ�d=���"O�0�AC-pcr�� ��{|=�%"O�8��)M<0s�i�@�r��1�"O�)Jp��1f�*7g�.Y�D���"O���%K�{D��@�E#��j"O:ؠE�)R,�p�O��Y6�(�"OlQ�`��{?�l�Ä�y%�t�"O$=��^7��!󇢊�M@���"O� (Q�&wH2�1&��2L�@�"Ot�����~Ā�v�"B|}�"O��Z���Z���X�`X����"Oj0:M�	If1��cU$,_hI�f"O� xl�@�f$�E��Q�TB��""O�͋B�]ۘ�X@��f�YH6"O�-�����怙�S(�&}��"O��9p��3`�@X`��2;V�"Odm�4��(BY��^=+mH�!�"OJ���D�h_� h�N)T9T�u"O0X��'�%V���4-]�<34��"OTA��X�E��@�F,1TŐ�"Oܘj�)A2{�D�hV�T�2P�ȓblܱ��!V��P�%`ڿF��|������щ6���y�eć.���ȓ2H����.r�$Tw��n���!Ӑ���Ѐoa���vh=8�`�ȓD�H�!�)m��8a��A,	\���ȓ7��BR4�tY�SI�*Q↩�ȓ{l�;�հ�ĵ! M�R��(�ȓ�T�����;��Ȃ5C� �ȓvǖ���f	qx�q��|9��}����$�/q�*컷mҚ(6h}�ȓo(d(�KĢ#��[ ���@�ȓh�����*r�2�AC<�ȓZV|�[DE@>L*�jd�@�j��m�ȓCx~���d�*re��H�� {T	��04�Rp'�����S�/����+����U�N6]|��dO�0ʐi���"��U�V�s����TeL�T��-�ȓ(j��h�M�n�&�üi�*х�7v9p��S��1���K�$�ȓ]�2�tp؂H�i�c�`�ȓU�V�cCJ�1m.����Ԓ/K�e�ȓq�Q�!��~#�M��A�Bh��V�( #`bN'G����1�Ss���ȓڂHRĬA�T�HP��Ї��i��Z�$���(�+��Y����4l|���5<T�D��`�A��!ɚ���1�R�3#.��کP�A]-�Ɲ�ȓb=��$���ȳA��'��m�ȓPQ���gA+TR0xs�Y+E)��Lx,�FTq�(� _t�ԅ�K��֌��d��s��
L/8���P�8��(� ���"CTB��ȓ_�`���/*w|��񃀟1i�d��,�. Pv郅E�H���K��*g����;�Tt��'%%�`��B_�-�Z��ȓb���Y�A�0-���A6#����d��i�F:(Z,J�,� p*����Yr*`Q�&�y�V*�m�m�������giԧ_� ���x��5�ȓw#��s��m�`�R�� )�Ň�n<$�'��5H���C����ẍ́ȓ1X)�P`Q�y[\Kfƃ�v�*u��@2,iz%O	, �6���f�8�d�ȓK|���¥�~����A��`���{X���-��d~���!�T�0�ȓ*� �SkU,�0�"�A1Dh�ȓ�֕3f�Ɠq��Yp��96���l�N))�g��03��h\+`���XΤw�3vX�@@�̞=�p͇�q�έ!(5	�Jq���`[.�ȓW#�� 5�3��XPwB��,uL��jy�Xe�X �ə!�ׇ2���=���K� �Q��j�:�b @�I�\�	�g��A����?9J(x[�K`�C�I�F^ȸy�A2pQ�Z�I����C�ɐx�7�H���}��,9i��C�)� n�@1'ZG1<	�1Ĉ2v����"O�zG��gj�Sc�]AFL�G"O
��K�FIl�ۂaS�*<��G"O��@��	6��lx �-����"O�I���:|�� �E��J$���3"O4���ɕ 2D�PnHP66��"Ov�
 �1C����mp'V��"O��� 6N{��r�e�BL�!���+~�٢�d�nc�T���T�!�d����s�-�(-]+J˚$���ȓ<Fj��q��:#�P�j�犑{�*@�ȓcl�{��oT}
v�]�v=�����!��Np&e�$�@�2�d���!�p���~t�t������a���ڥ�wf3.Uj�	1j�:>w���gF�Z�	�(j�z�*�K��J[a"O�7�^��@L��`�o�̅ "O��B�*!�Ip�����s"O�U
4��^(��7Ξ�E*]!"O�Er(���a�'k�)d'�<K�"Oċ����V��j }d`�d"O��	��
g�P��D�ñ?=*�q�"OL�zS���G���(�=;���"O�q�F�]6�u�#R�B/�%�S"O`��֮�k�yCU��Ы"O�{�ʘ/Q��7��<_�٘"O�E����4�L�G�	�kSV���"O� � X����#��8:�t#�"O�����*{,�P�ac�?p̕�"OJp����$�d"`�1
�$�&"O2�#��$]����vR�}�h�`�"O8ȓ�d�#�UaQ������	7"O
I��B�I%Jy�`�C�A}x���"Oz�e�?ÞM���L�e��"OB�O�	�5cHXԖ(�"O��	\�t@{�j�
L�ʉ��@� �y�#ֱDŲ�;',�*@����y��7�X�� �f[ ��f�՗�y&�*�T9*S($/?d�a�́�yr����N{��-)��A �,�y�I�'u���S!�H�6�B��y|�@�\(�J�KF�nK|�a��5D��!�lL�f��(��mD�qz��ZHB�	�7�2H��%C||`�ch�5}2�C�Ɏx!�͙�gV�g&L`��&"��C��;qu��� ��F6dq�k˛��C�	_��b��~'�@3�Ŋ�RlC�Ip�b�*�C%s�p�!�J `C�i�� V�@?���W!��U�m��'rz�S툼n�()7ŏ4���'4x�1�g�<�8<�'�A!u�,A�'l��`�F�?� !�J�|�����'x#�!uA��K�o�Lb	{�'�B���1S�L��ECT'�m�'�\x��Q$״̳�
��Wu*-��'�z����%:h�B�ՖR��|��'9����C�c�Z� �d�;%�Ex�'����Diو@���4e�n �
�'l��b�-D�oݶ����оeB<��	�'�jw&�;h>���
Y l�X�'a�M3�Iscԅ�&�Ĺ�
�'l��悍?���`��t��);	�'�b���ŢU��K�
;t����'>̭���7v(�B�F�x8���� D�C�՞>؎\"�B��$���['"O��"D�6L��� ��*Mʠ��$"O���P�����b��_�ڡ�A"O������0Z�	K�E��I� "O��,���1�??Fz�#"O�@��nF�T��T�@l�㬽��"O���R�M�B-hƭO�����"O~- '�#A�~l�"M��?&���"O�� +��3��@��[��Ÿ�'�t�PCn�1'��;�I�2V���'ܔ)�͗�)�F-S���<YF�h�'��bA�4XKvA_:Xv����'�.�LO6Y�$�Vc�8J�8��'��X�mɉ�}�����LQC&C�I8�d�+�� �TEy��ǜo?�B�əY.E���D�3+B�$d��6��B�Ʉ_d3�Ĕ�D�R�U*l4�B�I=$��0�&HI��9
�	�>�dC�	A����B�8^?�ո �$o�DC�	�M����dl\\jP�0�f��y�h�,� �A��Q�"-G�4�y� �
؈$i�D�
O�����7�y���+�D�h���^/�M�s���y��߁xQ�鱇*P6[8����)H��y� � PyD��!\*<���D�yR�¤n���S`"�=�� ��
O�yBHR)H[°r�Ț�5i��A3��,�yr�4D�l�#B**2Xɓe
��yLF\tA�1���zjxГN��y2�S�*�x�*6(�8lDIᢄ���y�͑��
��ƫչLu�d�� ��yR�қ/o�M�ե�;@hIs� 
�yb�^�Lz���!�L:D������y��sQ��4IN�`��ҡ����yB�=
�D�8�gS(eb0�t��3�y��ʡ���C���$%ҹb����yBT�S��]��'�3�phB���yr�'�r��eUI��@#��-�y��ԣ]�N<���:.~ET�ھ�yRj�"[l��チۃ@�:H��HD��y&�=v�^���,2A��ra��y��U;(|u���M-�Ȍpc�Ґ�yBD޶*L�$@3f)�f������y2cB�2\0��!�S�P�J���y��,Q���Cʸ�$a:3�J��y�*F6�|M3Vʍ=[MJ�K���y�-�wc�a�j��r$�2�u��jb6��E�$��eG4�.mE{��'e�<�EA��b��"�.D������'��������<|��Ɠ�K� 3
�'͠T�g J$#���8���F��ِ�'v��K��uH���@�˭;�^|(�'r~0�!�Is�\�0ē1�䔚�'ƴu F��0SCE˗JŻ;����'�L���d�&e_� ����/߂a�'4��"�柼<U"u+���j����'b�!��ȏ ����#:�L��'v�DA_�C*�� ��^�7��
�'(nsVB_�3PNtc2H^� !��'��)*��۔+`F�c!hz1lX�	�'�@=R���lD	Q��E����'n��4�Z�y�R�c��R�Iu�Tr�'~����4�����˼,�\���'�ʴ��kF$x���2#b�9vIZ��� ����2(~�}3�E�%F}�Q"Op͒4fV|
��z%�O-Nu��"O@��T��[jDMѥoSO��(`C"O�b��0I��m�����b#"O�T��'I�����=�Rq�V"OΑ��F;O F�lǘ:���w"O��؃IĤ}J\@�X6ry���"OBqc��A�#C�끊L�,��9"�"Ob5y��w�j9����O�d	XT"OzBB�̜����3�Ƞn�ԵH�"Of����n�AƩ��k��E��"O�!�a��)�B!BFW�n�.T0�"O��h�,Z7v����V�*��yE"O.D��Ϝ1V�b����9y�j9XW"O��Z�@qS|��R2A� ���"O��J��t#�#��ԅ.�j�@'"O�F��L������3�f��d"O���b-�X2h�"j�$|�X�J�"O.����yY�݀�		U�r�R�"O\4��P�V���P3*I*F���@�"O( 2'����j�O΄Jä�Ȳ"O.�I��Ӷzܜct���K�0Y[E"O���ܲD#l��B����`�q"O6=��I8RxC�+ʹ�`	2"O�����͜̡ 'k(d�|t� "O8�;� XE
�a���\(���"O�h�!�O#Uy�pbŗ}�(�e"O$D�kQ/sT"�"
+� �R�"O�U�e���Fo�����!�"O���P�7�`��E�}��@y�"O���ukA� �>zP�ƦTR"O���?PJޝ1��NM�y��"O�tB�� 
a��d�U�I(�R�"O`�{S���12��3aX� �8"Oh��F*l�.��D#a��a"O�hk�&IY�D��/�/Y���"O��i�-
�c��@� _�t�r"O
�$%@�J�d���P�(�ޤ�$"O�Hr�S�Ah�X�c�:����"OL@�B��Gr1�r�D$�<1��"O���S��^����GO]$`����!"O�%�pe1��0�X�u����'��,1�рO$��+��E�:zT���'��=���˯q�4e�th@,
pdh�'�>q����`E�����$�9�'�L@�Аt\ĉ��͜	E�d��'�^�D���r�|#0�֒v*��'� �X�oX�9���<YL���'�e@�#�5� z��S�3�*x�'�t!�E�-?��x�`��%S�Ё�'�Z�
�jW���H��"ـX0�'��P�)8����F��d���'"D�GiT���Z�+HJ���'��U�h��'�fx9%�����'�\��H��0����̘�2k>���'�$\R���.�f�+���.?X(�	�'�Z,"`��?Ш���D�M�($��'h�e"!CU����r�[�K�Uk�'�T%�i�-1��K�K�P�Z0y
�'b:�@�-��"Ud�W�Id�y	�'�2 `�'�x; �ޟLA�'�,�g������7���z�/6D��b��P#�,X�D�:i*��2D��I3h]�upt2�BK$i#���+D�� <�2���!%P`�%�@;q[�m��"OV|�в2ǢYB�B%l��"O�$�#ШJ�v��BX�i��Y1b"O�h"�
��'��y5�I���!�c"Od\���0�L��D"�C� �J�"O V�#tR�`�b�C��x"�gLj�<a`Ş�\�b�	�1]�1
"ʝf�<ө�	&��d@�g��h�V�kł�L�<9��_9/ (Q��׼*$D���D~�<ّ�U�lϤ5����5u�jt�6Oo�<9gJO==��8y�-������R�<�7�
�#@���� Z�<�a �%. @�fnՉ(�ȝ	�N[M�<ဢ��@)Ze�e�Ӌ{Zl,��Qq�<�,S��IZ�`�/q�A�J�i�<	�� �&P�R��ۄ	�F� ���]�<ц�*Y� i�6<��T�G�[�<I�ݾ'�ݒ׈��%�r�`�T�<A'��yF`鴪��lŶ �g�[�<�g�'Q΍��A����"�Z�<a�	���ji:�lL�B"����BR�<��,�kZd�FNH�5�[GI�<q�h�
f}K'�7.����ƊB�<�]�C�� 0�kݱh9f]څ'YF�<)�x?<,k"�P�5��Q�!�}�<�2�H�'��)��Z1x�����_�<�cEċTBQ�lR-fu5�@�_\�<y���?f�N��ɚ�;
�!��T�<�gH	�4�^8;���"=+�X)V��R�<�P@G5;c�I�E
�%~���Qb��h�<���N� �� �Ŋ!h�,1�o�<a���?����%�G�a'�Hp Sm�<�ÅFG�,�#��D�CnTՊ�,�f�<y���B����eL@�JH����G�<�E sx<��5A�	4����D�O�<!�/,-$���
�#H<=��lGW�<	P�O%8�9Ο�#��R"M�Q�<���0ftq32,�?>�I#�JN�<��b�uׄ(pV��@��U��j�H�<1e/�_gp�E�hi�#�E�<��#�������^��ഈ�}�<a1��Q����{+d����M{�<I6�ȤW�\�x��O5���c�s�<�s
��v��1���2*Ѱ��I�<��b��K��:���+	a���"
[E�<��j�+:�Ma�.βW~줚�g�<��KܤE?<y0V�L�_��T
GIZ�<�&F���5-^=��8�L�A�<)o
�q���eOe)"P�N�k�C�	Hc(��"�#2q�p�ңr��C�I�Hz!SF���@�u�7�P�GۢC�	����5�� d�)��B�4E�iS���M�ָ3!�0��B�ɘq>��M$Q��;��[�u�lB�ɪ@�����aHQ�U1aO�k�.B��%FyP�F��`�v�Sv�L�>��C�I:lKpU� $]3+J���-׳-u�C�I	V!�1�*��l�(��3��n��C�	�Mdq���2{����b���B�I�]18��7`^9�d��Ə}��C�ɀ#�,��J�vo� ��L��7h�C�Ɏ4^�@�WJ̝X�fL�c_!nC�I=��0�q�E9iTi��۠@A�B�I�`[F%����o'��*p�B�)� ,Qs��$[�X[0E�(h�Yi"O��rˊ1�{^͸Q���¼�ȓYZ��/�� ǲ�0vNA?�J��ȓi��H��'g�& ��ٻ�D�ȓA����яĘt �U�Uc�:Z$����:T�а��޾?Ղ+���6W��TZ���C!PS4iR�^�����ȓVad Ⳮ�	%���5�˾Cc���ȓz�F��`��
\�oǠงȓ!���0k׷b������݁eB��ȓ�d@է�VĜ���λN�Pq�ȓ)5�s��*j�Tېƚ:jD�t��C�IA�0zf��rU�L�rZ�|�ȓXy��!�;B2j��S%�?Tie��&RTQ�fKn��Qg�7O_}��%�>�C(Z(�XuL�
v{ZX�ȓK�|� ��1n�0�iC�LV��ȓz�;���pϖ��D�a�ȓ?��y�s�"q>"�yv�KZ,9��@т=!�@�������q็ȓZ?�!�uǀJ��X��&^p3�ȓ5�}�� a�Ń�Ij0��MR6��%ČSlH�� j��i��|Y@,Eft-�aQ6�>}�ȓmɤ���c�'��=�q<�<�ȓ�9[�(�+� 2�	1
d����83慈E��7B�m�d�22�����5ΰ� ��A�P#
O7� ���$��<Z�Wk�b�@0�Y�6k�܄�F�P�
~:�I##�(Yq���ȓm����f��m�Ht��ƌ�@�2������g�ַ!p���ǥP�:�(-��BRj��$\�7��9�MY�LK,��v�d�SwmH�s0Ґ�v��aR$��N�"�a'm��7-Z`�A��?DzB�ɤTy��I���->��y�lA�/n�B�I�nK���G��:U�La���]<C�	�{N���K�?#(<)�萧w9�B�ɑ9 X���Ǝ0��a���Bj�B�	�d�F�@�o�l��%`b��B�I�a:r�c�k�+��-(P,�f8�B䉼=�����x#���fԶW��B�	7L`�M���W+T�xᨳ+�j��B�ɹ`��$�U�ۓH�)6!G+f�ZB䉽g2lY���"�"Q��㊈3�HB�I#L�hP�#��2�ElH:T�NB�$mERI��-	j2�����Ĺ<�LB�ɗ�~��`(Z���0N�6��`�'�L��G
��t���u��tX�'ހP��H�[����@��h�lm�'���wÉQ�i��?_���[�'-Ly����n�|0��@��5
	�'e�5�R0P�T��"�25�2��'�l
�_<#���n91��l��'���&�
<F��V+=�8,{�' �|*t���S��-s��� fƴ���'�N��6��l�a�&m�3t�jl�
�'}<)T��;a��{�Z�Z�pI��'�,��m���V���e�j�'`�x�  �$��a���
[�.��'�Vu���I�b�H�BQ�_	Z*a��'<���t�Z�A��2!
����'�(�cثp�"xPcS��Ԑ��'�v4#C+禙ز�AK�A��� Bm��@�=��ةV�P�Z�����"O&�"���a�|<�@ͷA����"ONA��NH>�y$c�p3F��f"O��'��!�B�����wD�z#"O� �@U,
>�33�O���0"O��j���H�ް�a`F(y���"O�����@�p�*	���>��т"O��ۇH58t��@3w����"O�+%�п4o���2O�0�\�Z�"ON�zwG��w����-�.H�쨋�"O6	���
k��5���Z$QB��"ON�#��	2K׌ ���L��|���"Ou���B'{ƪ �M<3��R"Oz�K��
l��a�G�K�"O�����]�^�)��#'��q"O��q�͛�Px#PG��Y]"�G"O,�Q�N�'je���.1��g"O��8�p:��ڲLt�チϸs!���@E��e�?-JB�f'o�!�$��k�!8ݩd��Z�\�!�D�-XO,5r���Y0�y�@�l�!򤞹k25���Х`ݐm9��"B�!��4+�8h�&^�*�0f���!�J(H����Ą�G��M!F9U�!�dW�i��,�7mB�Z➽��-�9�!�D��h���E�N�8Φ���ݙ#�!�$��"��9���'V�ʴ�޹v�!�d�%>�r�P5cB�J8���u!���~�8�6¬r���� �� e!�d�q#��� �B�W3rh�7�>M!�Ϗ��P�!�'6mf`U tK!��F�j���uC�����	5S,!�(,V2q��_
>���_!򤌸)��ݪ���]^�p���a�!�䎚:����\P\�vlb�!��/Dh$�mߗCx��Ta�4�!�K4��-xp�L�0(�|qQ��)e�!�ӆ��PD�߽�{W��	H�!�D�3'L�́��ɝ
K��De�!��ոMXdmi  � 0���@�L �j�!���zݔ��#�ʻB�xX5,��7_!�$_ |Ʈ]��J�;�N� ɍ�!�Dt������z��!'m�3�!�䂆G� �������#�%�9X�!�$w���Qnͤ�6���%�&�!��dp�1��!�&x��F8,�!�$�c�.��V݀v���&��V5!�W�e�.1H`h�	���Є̃I !�$ޗKR�`�J��w�N�K'!�l!򤜷5��ꤋ� �j%���C�D"!��@K�@p��VL�A���I�,!�$Ҫ�f��
�g?j�h�7�!��C˼����B�m����\�E�!��� pV��x3k��"U��^.$�!�Ĝ�V�)5o�\E:�C�Ѻ�!�$Q)��5{A#y2��
�S5!�$=] �	��-K!�	���!�Or����	�I��%B�`#|�!�ă�k*:L�"J�`�x��`�c�!�$V�r͢���)^"�Bm��Y��!�Dʔ���x4I�SR�\���ēy�!�d��9�q��Ą�t2�-���U�P�!�D�,6��Ұ흽6u�2Ύ�h�!�ET�T+@�� �*�LN u!�� �(��F� r�`�\��-��"O��!�@��$���Yؚa86"O>8�b�6D0� /���@p"O��9�(�m��8���M�!����"O�m���ӻs,�5�5�y��3�	���+%��<u�)�&�$���)pDj� @�7qO ��9Jb4�և�X�.���4u` �O�t���1Yf�K4�	wY�����ĦpR�Y4B�8��Hɡ��@*$��_:�9q��/uf���)�M��-���I2%����O�nZ�(�O�P��+J 5N|hPBj����E�a	�O����V�{}��hj@���d��ۤ��p>�w�i��6�f�8૱	� 9��ѫWb�4N�$�a�
�M�fV�p��	qy�O��4�x����D��d�#�9t�7L=�¬/{=,<���)z��ڂ#ܨ��O��;-�`�����9��� ۓw]P�lZ�FM�5h��=A��ncC\��I�<"k�t�|��sj��S�׮r>Yk�J�d>�o:}h����ٴ�?����il� AwJ�%����-�.���'tBT�t��	<rL�Wb��DSD�3=�#=9�4Hq�֟|�U?���I��I�eA��N:H�Q�������'{04�lZJX��@��ƂLy����-սs�����b�&����$P��A����/��H�'L1#<�Æԯ-�8�e���t�Rt�!�ܷL�Q���I(e��E*5N=)����O!�fO�d��'B>�q�3�a�&��kâq"��OJY�0��O4dlڰ'N��<�����d-+�T0�� ���HQTBѴQ�Q�P���6@��m���xiv��,uq�M�t�i�7 �����X�����$�����Q��G3��1���ox���	��P�ȱ�ٷ)ab���oMƨۗݙ+�`X�h�2n�
Š'�� J瑟@����+T�V�Ru�5+�"���a��2����LX��c�'�+��h�ūN�)'`�h��Iڦ���E�E%��5��j�jy��oӪO����O�O���h�(��k��h��آ={"	��OF��d�9^^�X��/�1T�\X���y9���	��M���?�C�i�BL�q%l�z�d�<��89_f8�a�]|��MҖ�oRT�l�ɷ Gy�1�ђI�tBG�ܯC�x��A4��a�צ`��B�AF?���i��	�C��A��]*~z܅�c��7O��;XjV���̇]��DR��?%��@��cJ�OrHi`�'-��nӐ���~B1�ֆj��h�eJ�O̬TZCN:���4�"=)1$-,%n�r��93f\�v+	z8�d�شM��i��2,ߨ[F�u/��(\���'aLĚ�jy�N�D�<�O �']�aJ&LQ>��,R H���L�.Р�ru���es|PJrCϹD`KY3�q����w����t�I!0�MV�;� ���4z�6���(9�hI:`aW=cOl��6�	:'���|��5�Bp��J�澔ˁ킒��`mZ	�����O }��r��i�ZU�eIܛv�0-���ĀME@�'�b�'��P�z��N�XLX�H����~�Q�ߴJ(���|2�OD�N"<�ik�OR;;�A��!��9�$�&����	K� ��   ?   Ĵ���	��Z�:ti�-���3��H��R�
O�ظ2�x�I[#��y�4g�Բ �I�n-s�E�_�]	p7m�䦕��4E�� ��q�	x8�Ļ��My�֠�B��H(�Qy��7U�#<Q�
~ӨP(&m�r��xp@DB4F��r5X�T�$�����1?�E���/��7�f}2*,�1��l�?)��0��0L־�iP��uy�`�OvԚ6F� ��9O��@qJ��0~
�rt�
[bZ���(��L�@���'�,��$�ȄyQ#��!Ӹ'=�TΓ�|�YՌQ�����fn��hJ�$�<�ቭ!�'���#1���{�L:�I�h$�'�Ex��|�'�!�f�N	^PH�$$��}��-��&#<���>��I˟R��X�H>C���w�Y�D���O(��{��]�Jr؉[�B��K1�=S�,�MSV�1���"<���	��pˀ�8���(��[�HI�>q�	)?n��B�9Bw��2b^�H�����<�fȕ'5��Fx"��N��|� �%�L��t��'	��F'|�1 �?�@�"<	(�O�e(����.��L8��Ev�����$Z��O�D�O<q�	�W�؜1�O�"
�j$�wL]?y�3(o&�O����*�1	�D���N`!GK5F���l~.��>(��4w��	�/^5� �O�h�q�סe�8��F.[e�0�X����M b�\c�0�'�ǁG�'�b�S�������$�C�2��ۨO�����d[3�OL���LR&����f��0��:F"OL�y��  �~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  -  �  '  %/  i5  �;  B  IH  �N  �T  '[  ma  �g  �m  3t  uz  �   `� u�	����Zv)C�'ll\�0"Kz+⟈mZ�p|�57���DB���H1�ѯ&q�5��7�$�b�ی>��+�FRH XY�f��%e$���;F�FiB�'>Հ,y�'mx�a snQ�)�8=s���(-��(:0Lݧ||<Z���I<���@�'�A����4���蟺�d	�
`
�c땘,�z���0�	Z�DΐzRf��	��<��@*��ߴ+��9���?1��?a�n�>Pc�(�[\>�j��¢;����?�
�;���q*O��ğ*K�����O\�ě�a�n�AU��8C�"��%S��v�D�O��'�b,	!���C�?ٚ'9�t-K1Nz�Q�m0\�����ؗ/��2OP�Z'i��P�2���UI֥��Q��̓��'�P�2�#L�	?� �[$��)��}���/� ��O\��O���O���O�˧�y��ېj@�@SS��/m:�A�c��?���i�R6MSȟ�n�˟X�ڴpr��md�lo�Lce'������3�U1�X���J۾�HO���k6�'x S�����0�&/���v��o��@ؖ˞�x`���ڴfۛ�{��I���CwM�
P0����W�k��f`H ̂ �fyK�4c$z���� '�YP���,S�h7�5��aP�d��4l���M�V�N�0�rw�<8��1��!z]�}`pA��G^~��u�i��6��צZ���A:���v%�	Xh���M-�4�@�D����G�#`���pKJ�H����ώ�M#&�i�>6-^�q%��φD����fo��XJУӂYO\(�g�A&H"qo�����1ʉ/m���d�c5�m9U�ٟ��?�C�. �R��$�¾eu�`a'ǁ*Su���$�
����n�8�m�?���� W$�2�8�	0|�8xC#Z|���K'�5�ؽ��t2:9��(٫A�#f
�T�ȓ&�� 눓��#!�ӣMB$B剄�t��+�Xy�p@ѯ
sVB�	���'��Cf��yүY�3:B�	 
�,"
(�J0q
2"h�=Y�g]T�O�d��q�KiP����\�"2�R�'��jT"J"{Ȯ!rP�X2�X���'��:�� �ĥ�WH���
i��']�0+qo� Ub�@�7�������'ق����[z�+B	Z�wA.l�
�'5<%���hS�I���8l'4��#R��Gx��)W&��4@�T�9�%H�K�{�C��05��e%�� �\�%Iרz48B�I�c(@�ȋ~��Pi�㔣p� B��o�^��f���b�+��b��C��,9ej�j��+_%"BR�1p�C�3Z�ֈ9��0m��:�H3M��˓/=J̇��-O�����)e-ь�)"C�%��I0�F�%��̙cm��C�Il��ӷ��2���	v� *o,*B��������Q���h�fѴZB�%"�ޘ�R.#�bro͏�����9H8�n�۟\�	�)p�E���9�nek$�V�T��I������V��`�I��Lj���ƟP�'��N�zΠ� '�
1Ϝ�2�F7�ax2!Z�ː��X�CQp���~�pgN�P��rF	V3{ f����;8s<��O:�o���ء�+��s�$\�Sp��U`Sy2�i�R��)�=,�J�h������L19&JE����'MP�Q�m5��a���D�O���B R5$��"�&V�J�ã�'��I�L��u��ӟ�'��'K�$F�L*���]3�*M1Q�z0�	+.�A���;�l��9���p���M��)�@��.�)§m�ȵ��.�
J���U��j�I�'�����?K~j���h^�Q>6%(%	�9@�bI�K����?�	ӓ*�\Ĺ�Hϵ6�N�Q U-��D�9ڧHՎ��wȾ�p�C��>f�	����?��g�'P��F!�����B���<Y�'�(+�&k�|�ǃ�^KؔC�'&��@��Y�D����DK��MLM��'�T2@��9�V�kW�����@�'�,d21-�3< I��#~�r�'H\��H__t�R7қG��ܛ4�Ĳ�yB�'aH%Bg/��q�6����T/���A���x˚�Cw ����!o�`�2q���Mp�m��'p(���(c��Ш��~�q� �?�@�'��AB�'�(Dô�D<��0��'@�s&�1
W�49�A�7˔�N>�U�i	�'1���<�I�;q�6�c.�d��y��@R���\������	6$ $j�ݳ^� �)�-��f�,�� �I(�산 4^l��)W'.*���*0�"�flr��o�����?w`�*��-�FYJ�f�'M��, �����O:�u�'V2��XY�@%�JH"qO?��M���%���O���D�ilĺp�
>e�����۳�xR��O�u"���Y�.D�G�<ɼ�A�'��I6fך0�ڴ�?�����2��R,)�7�����(��kρ1��'#�Dh�:�p�%B�k��T>��O��̓�*K�.Q3T�ߍZ�����O��3�.��ڴy��A�@���}�El��aqЕz�b	NPx���M~�.Œ�?	��h�@�Ĝ�i����r��!��"J,B�	6b1,��4�ȡ	_����!r��?I���1D��`�@V�bc�z�j�-ZC�$l�ڟ��'Y6��pa�����Ox��<Ycl �����e��|y�"݌�F��"	�;�"QX5��&D q�*�>�I�o�	�$L@@h������9���E*H�2�a@sc,�6p�)��>�u���q�O�L�v��p��
�T�(L�bR�'{66��O�����O~b>˓�?�EG�*D�40fe�:d"�ec����8ړ�O̸)"o� p��x��3���{В�$oZ͟��I��M��������)��#�T@ce6ţs
7\�X=�4�	Ŧ���� �Ioyb^>�ϧ�^���%B�?i��c�,(]�0��A(�5������R�쁪V�����O���t�iY7��"B��<��D�W���D�RN��#���;R'l�6N��Ipޣ<��ݍY�
��b�("y�h;��O�UL9�I��	�4�?I,O��D�<A̟$�AU�͗��Rr��;qM�K!�|R�'� 2��̍1�4!���&{Z�����'��6M�O�b>���>){0�	/�(X�g���5'@��cb]�P�C�	�u��%f׎Xp���e���C�I-���ac�Yr�8����B�Y�&l�p��j��:0E�[R�B�I8
�Xy��U�;�z��'.�"�nB��;g�<T�ʹ�~a�f
�<�,�=I!U�O:Ԍ�P.��z�O��n���''�9��ҚE��@�EP�X���
�'��ty���	OS���f���M�
�'T�e@���G��!K�����4�
�'~D,J(/L�V+#a/\TX
�'v�H@`��`PE��?R�^�{�{��Dx��)�.���c'C�b�YҰ�ƓSTjC��%N�VH�3Μ�-�*�#�MD��.C�I�x|��`�U���E��>]�B�I�$n��ӷ�ˈe����`� >$B䉜3p�l�'+�%.�ΰj�@�� B�Ɏ,<�'�jh�őp�P&F>�o�T\��I&<�~��"�ŷ���%+�F�hB�*D}Иd���} �!�'jȖi�,B��v�ي��Y�X>~qK��E(�0C�ɲ��X��N�&n@ kH<,,C��
U�N�p��c�,������$�d
�$�6���`�K�(���*R�Ūe!򄇉v@ة�	M�o��I�V�M�{�!�����ʴ�[�ER�P�%[�ZB!�)pL}z5AQ�.�k�e�%!��RT/˗'����%_1E,!�� ;��K��C��Պ�$8�ў�P�/1�'i�PR3�����B��Vd����N��h#�c��M�le�q��\A��h�42�ԯ?�����jР�ȓu�Z�?PvN����479��@��x��8h!j��&`<QOẍ́�t���D��`����'*H�	 ^վ#<E���N��9�S@W�t�bEkuᕯ**!��+V�p�o�6�P�
ӡ��M	!��ؚ/j,�8 ��Z��XQ�V��Py�&�S�\@ё'��X�JiFؾ�ybI��S>)X�O�6I&��y�ə�]�����+�\UP݋������o��|"葬�"U��ŷ�eҤ����y
� ����,�nM��ʟ�v~h �"Oܝ�눢��£��t_:
�"O� ���4h,jO�DZ4|S"O�Cg�4�V�����cS�p2��'����'��AR��
�~Yj�a�L����'�4kr��q�Z�;�l�6Z�5@	�'���1I�'H�`�6m�T���B�'X$�$l�b�Y�#�Jr��#�'NF�ph~m��5+X]~�X
�'�`��엣G�}�ŅM=���ʉ��؉~gQ?=Hb,�d�J��"�A&d�,|xB)#D�ԣ+Y�rBi��!=3���@��!D�� u�V��@��2�da�W;D���W�6x۾���O�a��0+5D�xA5�ǄU���Bb���t��2D�܃�n�gl���ȑ�vU�0D��O���a�)����B�Ɓt��ѳ ��V��	�'=r�1�n�Вqy[v��#�F�<T�� H"�sw�H�mg�$�qO�A�<� �ep�T� 	Ѵ"�ZQ����{�<I5eН=�*���K�3���AK�z�<ٶ��
d�xh"e����"��OyR�W+�p>���WC�����^�l��z
d�<�!m�;Z~舡�Q�\,�"�^�<�v�0vo���f&[V΄�,O�<ɵ�;'�	)�
ƊV��h2S	�N�<��
�吠c� ��>d�B�Bx��Q筺����^�b��Ȓ�)^� ��!D�tr����O*4H	���m�Iæ� D�D�fl|_�Yk��� ��XR� =D��Q��4Pn���I��r�`ມ�/D��Ӫ֡@f���8�Z(���?D�L C�j��-�`gD=m0��k;��>mG��Y
�T��q[5Mj�zGHߖ�y��H4p�N�~<��c���y�@�O�n}2�B�,q��M�W�G�y��$"� �5"ޚ{U�1�B�(�yRĝ�6x��;U�G�x�>�@S	D��y�m\�}�B���_w���i�%ΐ�?! ��c��������Ŭi:6�� �Z�+�U��;D�\ÃF\G��<HD�9�؜�5�:D��B��^�r����KW*m@n�H"�7D�Ęu-Я����
Z/+�`A�g�4D���Ԯ o���i7�W�'�B��)4D�x���ۍnp��.
��"e�v�<9ƍE8���u��+
� 9k1�
*f�H��dg,D��6-�'Dv�4C΃�)"��C�.D�lZ�J 0�Q��_6F�L�PD-D���d�+N>d��蒱V�ȸ�N+D��@VgW�}]��9tH�\�l��F-)�O�3��OX	ad�8`�>�k�d��?����"O�j��.��!��c�/<r��"O��Q��4Bk��J�f�B�"O:����Σn��,�'I� �<%�r"O�,"�i��s"b!a@A�Rh�"O#p��A�r��r�2.^�xT�8<��~�$+T;J. ���)�~3܀���e�<��.қC�� ˳&����/�b�<����3���:��+G���[�$Rc�<�Ђ�2r,���4��le�W�<	T���&��6�W ]Ö��|�<Rl���P@�ϋ�@�P����@��*�S�Oʪl��oٜ$� ɜ�X[�4��"O�x��!�����)uX�SW����"O� ,I�d���Hsjȉt��8�"O�����ȇo�8�Qa��#6�ɑ"Oxh�e΅�a���	􊕙`��5"O8�X�"L-�����e��=��X����(�O"A��ÃN�0y�T�S�~l}��"O����U�;\A%�F<m��4Q�"O�9�`A�z���ǩG�D��"O�$Ȕ��K�RHh��z~D��"O�Y�ԫHW�|xU��΀�a��'1~��'�i��6^w�H8&�ֶ)��i!�'	�p#�E22V>�8�k'�����'��QG��O����ⅉ-��h)�' �<�nI�	a:YR`A6!X�j�'�N�1��r��ԯ����
�'�lL�t�B�k�^��ceF�"�҉��X�d�Q?�
rO�(�Q���α'����D$D��PB�&hL�zG�A9�>�2P� D�l�a���%��ISID@�B��?D� Jգ�9L�-i��)Ya�b8D���M��]���In��3��4D�L��%�>��z0O����O@��)�x^���^��X��荃�^U"�'�l��O�IYڐ{T�+Qެ�
�'Be��$��l�xȁ���?:�ܵ8	�'������N�BM<�X
�/���	�'����bN����h��H	<�}��'�y���ՂW�$ŘdD�6`|,H/O�$i��'���窎�"��k'��%,�}X�'?lt�B�'[G>�KbjT'�`��'c��)DNO�{N6AB���	�-��'�A	�˂�8�l��E���}!T�p�'�ܬ�W΃'�I����p ���������HE��
5�@�K�1h��ȓ��})��ѫ �B�h��L-q�����h��iծ"�X����E��y�ȓkߪ���#aB�Y�.^K�t��_�Y��D/[��H5��3;�E��DA���`H��Y��#-(�&�D{�쎯Ш��0B��M���X{���	�ňa"O��Ru��"�n�����,�>t�1"O��(��6=�(��Î���h�g"O\�w-ӱ-��{�b�"u���{�"O�͸u�2NhjUX��T�5��%�A"O�Y�%� V&"5K��߄$���'�'��������>��J��Z(,x(�S�f�4���ȓ=A���p�ʩN��T#�D	�i�ȓL쎁�2#�3.<�����YG���ȓ7�͋���ҨQ�NZ?588܅ȓ	i8�hg�S�&r�8A3��/b�D�ȓ��U��*X�#�X��#��S�`�'�p�
�>���+�뉂/������X5zd}��J>d�tϜ�S��H��R�U��4}h��`���0����Gʘv��T��rnd����U �p�q��0옅ȓn�����&��k:���eI#ȭ����r�6�ɲ(��Ɉ!��|�f ��R\���מX�̼��@�)=`�;��L�G@!���
��ٲê7�hPdeX�B7!�$�fJd���$8�:�i�c/f�!�_��E��j&;�aF�L�!�DK(I����̅�+>�BЁS�:ў+�%>�'W
��#B�B4 2�h#�ʆ?r�̈́ȓyun�* N^�)���rw"�ԄȓZmb���")��h�6!������S�? ��o�-6�%Z�͔+�X��"O$���F.©�FK�7&ۊmY$"O �aS��G�႖�{Ǝ�t�'��p���S�q��)t�O�a̜�y��Z��z���P����
 8(�y���ͩ���ȓ#ҒR!Ҟ1��i�@�nS�t��q) 5�ል�*��D���E��H�ȓ+�D4���'�8��Rk�-d�v���g�����3�T1HR���V��'1`�
�8�r����@e�bICS��"k��Q�ȓ��Aq6E�q`pQ��[.����i/�Y� �<l���R�י
|�ȓ;-2���'�k����Hx������j������4a[N�a��QAx�h�&��XqW*�G��m+b�ԡP����Ў=D�Ԉ7˄!09x�Ȥe�*|J�31�:D�$����	���C �A}*X1�e9D�$���/;|�Qү�k��d���2D�<*�{��a�9M� ;��5D��AnǴ����Gf�3a�2�4��yD��+����7��E��)I�y�k��P����tcʚ)ZlA*�.$�y�h
8�� �A/|ک�&E��yDY<l؂�kς!��t�&N��yҫ�}2��j�f-/2<�c�=�yѐj�(8a�S�Թ�J�?Qb������R!�Z�)�����"4�|r:D�أ��W3I���26	ɓ�|���4D���!Zd���,��>d>@ �3D� � J(�4�P�*�8o  �6L;D�ph!mu�6@� ��th<���/Mp���)L��C��yR�����O� �Ϩ����O��`��ԮF����ʊ5+l@ັ��<����?�cujFm\�;�qKG�n�y��O�2�I'F��mI�IBL*��@���}Ԁ�1Z/�ik�ꀐ��$����j"8z��0X|�!���R�&Gy�R��?����On �1����o1h�8��\pz �,O���d��d��") y4Tmr1Q�2q�}��<1�B�.Ǣ��D��5�D�[��\y/� #��'j�I{���'k�BͲK�U< ��	� PV�-��.(�XP��J��K��x�j�}���!^�
`��D�Cd�X����<a�)N9"�4 G�Ƽ	52Ё�E9h���c"8�JH�!�<W0օ��(��dF�I���$�O��S�V~�gO)"�� ��p��y0�`�>�y"R'5
� ���kji`����hO��F���э�tz�+�+ִ���ܱ_��'�R�+�����'���'5��O^��Y�H*-h�L 0W���$�Яs=\��G�}�J�&��j�Z���
+���D�4+G���`*�׺u��E	������A-;�ΥH M�@X��#�?%�Ɨ�ysh�6��I�i �qP�av�8�R��'������?����r��:���-d�$H�7KH���FL2D��	�鋊H���+Iغ�#�O@UGz�O�Q�|�ՈY�k���wa�u�\$WD��mY�;3	J�踤����H���?1�IΟLΧE6�\`S �8&��,��"�:���ĦG�k�PR1,�+D�I��4H�"?9��O�"�2���:��\j��`!a6)�h�N=j�A>���� 	f�ʽEx��_��?�%%Eq�P�0ð1*Z��� �?���:�hx��k�v@���>E�ȓCOHA��+N����c��U��'�7��O�ʓd�Չ��h��1�����&��(u#��� �i��	�?IńO�?����?Æ,`#$��@➆=����|����?`ܝ�d��Py�SPE�~�'gŹ�3$�L8�#�iK":y�钮�Ow�d��k����pQD��O���(��1]��㲨�/��D�c*ɪ!�˓�0?a�	�~{:��5D����elSx�<�*O��1ŋ
J���t��7B
^����4J���,����� !V.��9��`��P1�Ix%�-D���%V�E�d0H�ڕ�ne��$)D��9�JB�J�4Mrb հuI��<D�� >�xf�:���1%o��rl�M�"ORYR�»B}���-& ���"O�萱(�*Bt��#��r�����Q��O<�}����Bs,C��3ӡ�6�(ąȓp=���.��8�a�1
Ե}�Y�� ��!�ł�:XRL�īƭ;��0�ȓJo2(2�������$�#g����ȓ^���5��;_UB$`A�V���s����GQl���D�r���Ƀ3>p����&L����ō�:`����Ɣ26!�$�����c� +l� �c��?%!�Ď�*�M�D@[3����C뚈R!��?5)~P觌�K��%J3
�n!�D��'B��J&�p18 r�[џ�����M�I>"��=�|�[7`�{�p����X[~b�'�"�'R���aؕM���!I�����j#�����J5�=4�<؀�sz>�X��I�fƚ1��0i��x HK:.��M�ڀ�a��ŋ�Ѝ
��˃A�x��2�I-���d�O���Oh�S5���;�T�۾	a�A�r�P�D�Oh˓���	>?q���L��"� ���,3 ��c��|l���d�u싮Qo�E�f�[7�ʴb"�꟨�4�?Y���?�.O&�d�OX�5L�Չ�iMt�r(��)�(@���'+Q��F{� G
W����e�5d�V����D'��'���K<�g-�O:�'	���qE��i=��2�OW���d�'�z�	"�ӧ�9O�@����$I
Y�'p����t Pb��Op�,�&��OV,$?�H�E�<U�܈��ꅣ:v���5M���Ɋ�~��s�L��M�M�V�K�a(�`ABM�rn&�'t�';:q�J���>�B�`��!�8df_�mt�,�?Q�@�x���U��?9pK�$wҁB�M�bxr�q4gV��r�"}b�3}R*����ə�Mcs��#\�b|)t�Y��`���ĝcyR��9���ȟ�PA�v���f��* �����z?a5(I�T>�I4�����֟���'B�|��i`�:eo؍� �\{�u�޼�'���D�T
�B�B��GL	{O�1�p"��?9�L�����!?��y2��~��?J�(�a"D\��䙈Gヹ�?��m �O���f�J�pt �Ie)ʿ�Tcw"O� G��9_�Y;�A�31�x��xRP�0$��Sٟ,��9S>h��o��n�I���#��X�O��O8�=�OR�Aqo��CΨ��Ȁ�P�؍}�)�	��~l[ЄW�z.�z�_+!��ش���*�3����7�+\u!�Dc��� IX��h$��*�=!���yAb�1k��� Bgk�!�D9;\���(ʇU���goi�!��0�����B�ks��`&X�!��3n��p�P�R7Xtp� �i
!�$Q�'Ʋe
��K�9�:pz�
ʔ�!��/l)X5#�O�:m�=Є�ūE�!�$K
A2�V2I~�x{�"M$Vs!�dO�������@S
����O`!��Ao,U )Œ&A�pQr�
 %d�O,Q�$�J����	"]��y�E�KR�P� ,F�h1�1�!/���7DU6�W�Ly�a��C�t���"�M�DY24p$;��4(4)x=椨ԤA��o�D�NhUÀ�o���BD�O�& ^y��o�X!$������s���AG�u���Q��F�	 .���C/ �D��&��'Y�#<Yϓ 0�d3S �"O. �"��!�ȓJ�d�A�ʃqk�}��J� %�Q��Y�Q�rI�dn����B�\��@��<���a�N��S�.�����M#���ȓ �&�0k֦���C3���0�����_@Y���	�2܊$�	>j����	��sXn�
���d1��b���6�[�r��b��;�de�ȓ+��31�����6�t]$p��rX5S��|�$B#��*ʢ,�ȓ	leX*��f"u��S�"����@�2i]�=ҵ�4�ʹRFp��S�? R�)�D�."~��RfƘ�N@�D"O�0p���wK<3GG\Q�b� 6"Op �#Q�=��L8U�D�{��|��"Oܬ��V�4����Cx%`"Op���*zX>��B�%<ʼA�f"OQP���@��<;#���z���hD"OV]�C��$3���ϖ'�<ɪ�"O8x	%�Ւ9��T�%��P�v"O@���Ub��En�2X
��"O���a)V�C\����j�>CR]��"O������9���)�<\*�"O���wE��U���R�G�' ���"OhU��.J7?�F��򋝟uR"O���(�}�H���F�Np)JB"O��)gf�0L�yp���%�Z��@"OdY�t���+�)x��\	"O�m��D��l`|�k#h�.�Va T"O�@Ѝ�{e�0R"hؑI2�̀�"O�$���C�V�)�MP�2�R*6"O�ݲ.[��t��
>7�
�s�"O~��mX�r���WO��D��"O��QV�{� u��JعWmz�5"Op��^2s�J��J�RUjl�"O�!��� �"��sc˄Y����"Ov��%�C��||z�D޼;B 1X!"O��0X����# O<�A6"O��%�:x�!��eΐ\1�"O���R�B3�� fA0�E��"O�h����>���B�
��*����"O��#M�9,ԕ��)G'}� ��"O�лэU�gj���A	���"S"O2��ݧh�V #� �2o��Q"O�)�TK�]�$�O�-/�>�Xc"O���O08���z - �Iߠ)�"O!��0Y����Nk�B�r�"O�M*��Ӫ�jPY�#¤��E"O�t�mշ �r�8��+"����P"O�L��F�{%�=lc*��Q"O�%�.@z�����1{v]RT"O��!��0�b�ģ�,Z��"O�S���RԠA�FÃ�S4��8�"O������36
���"�<mмI�"O�	kUă.Q��TCS�Í��"O� "�F->�����/.g�~�iF"O�D���Q�a*v���ӛav��"O�ä���y�,
��?U��"O��.\�,���-@T kRkɅ�y����U�ܨ����h����y�DŁ HK��+jJ\Ј]��y�d�2��	xԇ�&�\0" �2�y�χ�k�`@��"R�'rN�@�9�y2GƫJ��ĉI����O���yrb�I�f���ӊ�v�	%C��ygE�td&\[BB��}�����y��}��E��*� � �bE���y�5Ѻ��ī|6���Q�yR��-��b�mtԞ��Ѭ��yb�A�\���D��r}�+� C�y�e�5�J)ЖAęc��yK��N+�y�� <XЅ�«U�DQʷ%��y�#��;\�ьȋGdm�G,���y2�W"<ـ��@�7L�p`�Z��y� R�"�I�'
=6��)�#��yb�$o��8�����3�Z�hf�4�y
� ���a�E!��#BE�2N˘�2"Or}��(V��^��ġ�'(��x0�"O��x�o�2��
�J��>�c�"O�ɡ�	��\Q�*� 	Ϛ��"O���N̈́`t^��lѰK�`�	""O��@V��hچ��b�F

 �v"O�̀��ݍ'�	��
m����"O֜hG�ЙT1P�1�B�?��Ȃ "Ov�cэF#A�j��t�K;\�Np�#"O�yqt��0F�2��_�K�����"O~4��+�i��u�0����H��"O�ȷ�T]I���q��l�]XG"O�(�#��|q>\{������"O��(Gg�cTt-a%N޴N�^ْ�"O̐:$O�P%��m�Uh&�b"O�`�T`�s���U�X){b8Y�"O(��E�W+(��L� PThQE"O��qB�I�>}j�˶�j;j���"O��A�(�w�Z�X��	R2��`�"Ov<����!X��=KGL��p0&`b"O��r*E#d/�����G,P�Yj�"OK#m�����C�?�^�"O>�$�H?аt���&�1
�"O�H&���t!(�b��S0%-;S"O����&��Q�ɣ#4���"OLApщ�����6��� �P"O�+��=JWF�1�e�	>Feڧ"O�4�4���?KP���?$郖"On�YUm���l�$b��d+6�s"O��3��Uv!y��H5�5(�"O�=4K�h�����!R�W����"O����#�3j��b��0j	;e"O Z4���D51��ƕ^cfm�"OZ2sn�pFD�:�O�CEJp�"O��{�n
�\��܊�gܭ]).��"O,�3�+�q��Arc��	u��A "O�4	 A)����!jņX����!"OjS$h�6A��K$i�6l�"}��"O m�nB:=�8h�P�h��$r�"OȘ�Ƨ��sy��P�փ>�L<s�"O�>;���bn(=�b�A�"O��`�CK�oH8�(c��k����*O����`ؿL��r E�T�[�'ֲYѐ���2l˂g�PڒQ�'�FQJ�)��䀡a���3/X��
�'fZqh��h�"�!�
(b�<�I
�'nd�Z�f�"�����ϰMK>͚	�'V�p��\(�t�ǌ³?VD�A�'�E!�֓X:
�@7�W7��`[
�'Ω��.U�u��Y��z��
�'���Q��/=�@���^�b�t���'W$� �dI�;�l8R!�0O���3�'w��eG!T�e�򍊗PFν�
�'f���f� AD��ѫ�H�F��'������\�%���H&ԁ�
�'�R0�L"FwV� ���r����'Ȗ�A�܂8�����lа���'ȶ�y"/�wġ2eˎ/4Z��'��[ATU�"�i%F�0��}
�'ܔi[a	E3+�"K��(�z��'� �j7`]�,�N �đ��z�;
�'���b���&��@0�� �$���'�8E E��l���J5D�	{���p�'��tf�K�3MF����lf}���� ����	���@q���3�(l2�"O(QIըW$r��8�D�	f��
`"O��A�іxI��� �<�\h��"O00Q�70A�}+�$N/(`Y�"O+d@�e�V!,��\q ��.�y2+@=b��!���""�
�b��yɜ8;��0��!������Z��yB`�뎤��E�K
�R(�0�y�l��Mo8Q["�D����a��yB@�#�D@��7x̠�搕�y�h6��$Z"�^�y���A�ņ3�yR@�(-p���Q�n�xqi'X�y�ؾ+��h�����3(N)�y�ܝBpf�j '�H�u����y��+Y�J�@��6"��b�Ά�y"ƌ�!&����9to�������yr`�D�ȓ4� �g#&�{A�G��y�I�_`݁�GAg,,<BBj�$�y� �#gY��I���X�"@wa�y釻J8T���%#��P���y2�ћf�.�*scM#<id@���y�� k�
��$\ANlz.��yb,O�.���D��UP2(�OC��y��
�p����� A3Q�����Ͷ�yB��n�T���!��5h�8b�]��y�$v}�s�� ����a��;�yr�^?*��55g^?����0�[��y��R�t?���d� �RXd �y�d߭K�T�g)9_��J6����y��6>#��b�G"u)��;����y¯\&G��	��)��$�U�Ǩ�>�y�D�5)��cҧ��r5ƌ�� �yC��dN�a��S�oN	���y"l7'&a� B��hh:�.��yr�N�@>�r��
&@�s$�F��y���9��,;�"H� ƨ�+� �y��@�OI�4�������u����y��:7�n�V�	┽�A�(�y���
��L���L��d	��y��Y@�qQi_�J�>`����y�F	:��c/�%U������8�y��ǆY%$����µO����%�y©��66x�k�D��������y��M:*/H�q� �F�����f	��yR�~*A���9�R`:��3�y�
W��H8�LΏ!p\v����yBF���h���z3T=�%�[�y"�Dh��𢠉q�0�T'��y�G�[�1H�V�d�"XCi+�y]5_�渑�	�f&L9ٔ#t!�$�q�x�WD��e��eqq�ڊBq!��j$��A��7ux8Ԉ�
��6f!�d/v�������,rR=R� F�'f!��G�$M���፹t�����ԜML!�_�w��z��Y ��94�z9!�'G7�Ո�*�F?hѤ.I8/!�6T��B�02'�]2�F2& qO�P'0T�������6J�8��|"�ֈQv9{'�A),�mh��yr���Ko*�y�� r�B����W��y��M�O���l�":o��U$B��yB$��>Qԑ:�E�&*T2x�Ȕ��y�h]�orhQ����R�\���!��y�
U�	�"L�B��T�*\��yb��- ��8خ
�fI��/��y
� ���6�I�)���c��ϙ}0RDJr"O�)�	�;��!��D^p��"Ol��瓣<� ua̵�J �"O�XQ�g@�hl
����y�L%��"O���b%�9qw$L��+�>� "O�����؇q���{��:8��"O����W�M��I�bG,d��K�"O�U[a�*6an����D8DP"�"O~��E*؄+>0��[Ve��!�"O���jV?x�՛���+
� ��"Oƙ3���E�>H�Ħ�<ǐ�!s"O����F
N�ԳC���1��s�"O�e8�jG�.|1�w+��n��$�4"O�Ջ5��=��ɞH�@d@Q"Oh8R�/ż`���7��.Z2��q"O��[E#L�@
ژ��_2��h��"O�h_b�8{���i9�"Ozܨň�)C��5�Ġ_�m	�hs�"O�D��/]�a��Qs�I%R�0}��"O���@��$�RF���@["O*	�,s4�����èi�½��"OL�"���,�p��0E[���+�"O��q�AP"����Q��,E�"OFˣjT��}c��Q�97e��"O�e�`��m�v�BT�̡(+$�kP"O꩘T��,y�PȔ8��5�"O� ��`��F�YC�׷q�t� "O�|�-�8���H��E� �:Mx�"Or<"Q(R�^�RmA��̄s8 ��"O�����ɑ�예 ��O��"O�d���7[�t[d	�:HA�1P""OrM�J�)V���$h����(˴"O̬g'�D � ���[s*��E"O��
e.lDj���ݒ[b� Br"Od����PԀ�����, E@�w"O���'� �u��胀
*����"O@�$D	-]"�B��A��.�"OTx9v,�:O�L���+G��"O��B��6Fl�P#�O��,���"Ox�ю�P�XՉ� �!P�yc�"O"�
����%-ӖH��T����	�y��N���Y6
X@�
=��̉�PyRHT� -<�3Sn�O��!p��e�<R��*a�=RC�ڙ?�Ʃ�b�J�<�w���.�T�����.�>�&&�D�<�$��T���qjP���Sg�I�<�k	J�����?�Ҭ��o�<i����LДcɾ�[�'�n�<�$���,�$	;�Y�'�S�<�flL�T\���� M�n��-To�<�E��d���×#ZԐB���l�<�r�%pPF��g-O��~����Us�<�S K&{�>��$ѓ;��ۢ�M�<������"�I����#�e�E�<�cN<
Kʽ�e��/B��D`�B�<����h�n�Ze-G� hT���y�<�kM�@�&�J3	�-�֦Np�<9��7w�n������ZW�ɑχc�<����,0�a0���hRpԲ�Kh�<�� O
��Pum ",���S���b�<I�%�"SX%���=a�����h�<��ԗ� 1�kŵ� �N�E�!��%95��j�(X�N]�����$�!���8%��A�dÕaun��t���!�� ��A��*8����J�U�"O�,H����r!L�ل{�s�"O0D3r��:�"�ó�E'���zc"O@�"��B�T�8e�'�ł���'"Oh �3*P�=Sl �bj��X�����"O����N�.�ts&�
<�H!"O�݂U���F��M2�(u0�T��"O:]���B	\��.ѨB�0�D"OƩ�1g�(ֈ��n��}��!z�"On�S�`_�q8��r '\�'����"O��S�s�"m��/�8�>8��"O��¢�H�}~��s��^R}��"Ox�p��M<&p�ؠ��ٕoB��Zd"OԹ�$iNJ�"Ҫ���E[�"O�J�J۔P0n��ǬY�T����$"O��x"
 � ĸҥIA�.�a1w"O�E�G�*u��XpH�7����"OX�H3h�nвI�O� �"f"O��h�K� E0�L�ٴTP�"O08��Z0��	r�@4Y�ܔ��"Ox�s/�B�.�!j�|�J� �"O�aP�Z$Hf	Aȋ�v�Kt"O|� ����M�`=�q�֝ ʆ��"ORq���ɭ0�F�ѓE�e$�TPv"O5B��!���fD8p�� �"ON0� O�N���.ǽ&4T� �"O��5@��~�X�
�D.�#�"Ol�P���6,3և�(,���C�"O`,����9G�sG�h����"O��`F��s�
���e�-���"O. Y� X;�����R,#�"O����3w���X��F�Y�xK"O��0"��[QN0;f�^
U��]�"O�)$��~x���D�ޚS$�T��'p��+7��W(�Q�H+6�^���'!(\"�a�V���㍴.$nU��'����D�
+R�� �g����y2�'��$j NT�����QA]m���[�'O�X
�KR�4b�9ڰS�69��@�'L��L[<"F�K���=f.��!�'Y�`:C�K�\��H�@W!Q�� �'�|����1�N�����FԈ1a�'Z��r�F�9��10g�U=58
�i�'���y�oO=)�.q���\�*���x�'�m���s��LP���*RBI�
�'�~C��4tJ}0�ܾ$��Y
�'�8�r�L�3$�T����>�D��'�np�[Yf:�"#��H\�R�'���b���:tĉ���B�8�>y�	�'m�2mR"s�(���bZ 2Ƙ��'�D!0+\�ځ����+��P�'��� i�?$�|����Y�� �	�'�\(
�O[���CʳW���z�':��u�#X`��3�� �	�'}��`g�00�����)�\l��'����e�O�7X(��/��&�<�K�'@#�$ѦZ$D�&�����p�<�PE�$h�|�@�ȚzZ&�5��H�<�ul@�_�Ƙ����*6l�R��G�<AAM<E�q�D&�$J�3�CW�<q�b[z.!B�uqd�˅h�<�iH����sA�;��h��˃l�<�A_�U窜Q�CFhJn�P�/�B�<�d�?q��=�&�P*&�^U�RhQ^�<� �,���'E%<P�FK�2�=1�"O1@��R�c���s��@ψ��&"Oj��e)T�QV*�2iȷN1�!�"Ot���h�^���
I�"#.��ST"Oh���O\!yD�! �"}��m�V"OLi��
�bF��!�:[��D��"O��(q�X'h�hl��l�2o�&��"O�Dh�ꕢ�0l8��"�.�p�"O@�:G�ڌ^gtq{G��aϺ�s"O���TƑgX<�J��V�_3n��g"O\�"v�A0k�f�����.���"O"�A�りTE���+	z´�2"ON�!�H\;l���B� ր���3w"O�1�bF��e�<�yQ瀣9����"O�p:`Έ%�pS�]���*�"OvA�F��L�r@��(��	8�"O4Y�ʖ�O�xѓ`0;���1"O�� ԍA��D�d<J�Nx�"Oz(�E��Z�P����J�r"O��墈�
��B��06��ڡ"O�(�մ�H�yF����,�"O����1��L� n��r}�8��"O�qx��[%���Y��(JA�=D��¡o�7�I�+B�Eh�<�#�0D�HZ懊.���Ǖ
=$��l=D�(y%�E�x��lU�F��U��?D�� @*��W��y!�$_�t�cN;D��z��6��h�����H�a�:D���!�0PQ�`O�Q�:��Ć4D�СP� �|]��)�k�B��%3D���E��@O��{��G�"��X��2D� k8tز1$đH��@�1D������)M���m',kڌ0��3D�|q�n�?!�蠢ҴD��2�'0D�T1&"K�'��\{��%\����1D���A�_*u�a�.O��m	��#D�@�E�~Bz�X�O�=��xѣ4D�X�����H1.f,�5n\�=蚌���Z����;V�f�R��=:�
D�ȓAX�|{�T�a]t��`(��4F���ȓm��9ɕ}0mj���F$B��ȓtAn|�e��v���SQ�U�¸�ȓ@��XQČD73�xHk��7I�Xl�ȓX4r�;�e	e���@1f.���v�,(W�ю&Y�x&o�05��ȓ��8zbH f�lD����(3�I�ȓl��h�MH!ft����*VF��ȓ\d��#D�y��ӓ+Z%�:(�ȓ}�t�D����}�a#�5/�A��3���9��9�: o)�4$�汄ȓv��؆jʖ"�����a���ȓay�Y�
_�{G�A@6�	)kf��ȓV "aԉW$��'�6�v��ȓb7�P�吹�� 蓪��]R�Ȅ�NV�� +E=���i�C�'q��q��d�e�K�]`��ې�ˠD��ć�_GLգ��
\��|��S�/���z֪e�`(�lhx�f/Ɨ&*��ȓW�^	j��2Z$��g�J�V81��P �A��aȏ;�� ���$��ȓs�la#��714�q�!
��d�=qԍ�v���a`1m>��S�I�v��,M
|6ܝ�rC��;��C䉡@�h�Srb� .U��W�N�s��C䉠{^��`���~>qH��MtU�C�)� D�A���&j<����H2E��"O�Y(�l�!�B4#U:m:�	s"OFHu'�X�zM pk�<0��@�"O�\��E�.tY*Yq��<[��Pc"O0e�l��|i�!�Ĉ�0=*�h�"O�"����셄�g��H��=^�!�d�r��ے���;�&U��&�s�!��Z>|
e�`.H�5�J�0�凩!�œ.0��쉺]�be�b$�fY!�d˾R�2��ӎ8?�V����>,o!�$
�)��T���U��-���	$ZU!��\
yi�M DQȥ���\�!��@�C�����MY�,!e�
��!��0�����l�F��#���{�!�ϪI$(d� mD�x�`q��K� �!�ĉ*�}B��>W\Y����0,�!�D��Hwň��%BZ\�d�i�!�?#@p��G��(Ḷ�#Z!�d_K��9d�E
^�lI��E8-�!���% �����L�fE)˽
�!�$� ���
w/o���[�x�!��05�2Ap�E1+�̂�Ոw!�DW�.��t���S�6ǲ���>a!�$��Ԩ�IueX(��U�
շd�!�$�z*��V��
�k�?GY�� �'���v
V�w|l1�&Csc��{�'A^<�4��x,1s���_EB@��'���ӭ��y ����: ����
�'4p��%$�5J� �UoN�t�8]k
�'��9��� ����+B��N 2�'��!!�Ð�慨�᎐y�``��'���L�60���C����'w�PC�M�,���eiU����'����G�^'1z@���N��*�'0F�QvEE�Op�9vF��-W�(��'�0T�6�G�"��E�ΦTr^��'!$�A�O��r�#àFƂ�y�'c:X*Q�%<���ɒ�˷@
�<��'���rO�{�V���kC4;��	�'�����ŋ�6��r�K�[�z��	�'�K�(+�Zyq��	�x�,�gQ�<aԀ�7	��$[��yG�PO�<1����	�� �;4z4���Mv�<�O.i���re*O�?N<�`�n�<)��G:
D5&=��9�Pl�<	W�̌_�d$����5�^�q�g�<qu't���!�	�O� l�f�	=�!�ZP]>�sA!Q(~20�c��!�$>x.�;�I�|h�=�s��cA!���3n��ʠ�MM 9iDT�j	!�$I/T���t'�a=XK ��!�D��1Q��R�mF�P� 9aQǜ}�!�$ٽx��������r�+��b�!���2d�D�&R��� �Z�!�$��@�e����w�a3�MT�d�!�31C��3�h�,�I��,�!�Ďy���pQ��;���t�Ѩ�!�Ą?B�h +b*T�X��D��!�Ě�j�<�����#�|��\	�!�	>X�(0j�	�*��q�`�=#c!�D� д1;������C.l7!�D=I�Rђ�׫I�[�CP�MT!��Ϩ/v�P�F�5if�y�f;!�D�/����R7��Q�NG�Z�!�� �1!W�0��j��߮`�~L�f"O��'IX4}��M(Ǧ���̡"O���r�Zy�h�҅��`�$(;�"O���&#5/�\���e6$E�#"O�`�t/��F��s�ɐO�~�H0"O��{��ٶN%@vd��К "O�T��	ɔw�X�"�B@��l��"Ov��0)�((~q��!So4AJ"OvP��)O�ಯ��8�X"O蠪�HS �����m�6t�����"O��6�Ӧ0�dm�VL�fvD"4"OVP�t�ƷN5�	���΍aO�x��"O�E�'g@
f�P�D	!	4b���"O���ƃ��n���B���7a` "O�X�mM`���iG�y
���"O00���/����b���/�1i#"O�ࠧaHPH*Pʆ#7����$"OT����<2����\3F�00"O��NK�7a��1H[���͹�"O�Q	�(P�WT D��[7>|��"OH�P�e\�n�*l��a^6h�pY�c"OP�`���VQ�<P�'{*�s�"ORI��(����R�e��Ȅ �"O�-xa���]!6�`�E�d�zl��"O�V̙"<D��$�w�4䲥"O��9%O�7���`J�"'�X�@"O��b��E+�nH	gh�ZaXf"O�֭�*,��#���`���0�"OJ(	R"�iL��SE˪6vq�$"O:�yf���H�)!���#DEbs"O�p"cWX_�$:�C��ޘ�"OJ�c� ԧc�����- �4-["Or8%��E\r-��	U����w"O^<�bX�^���
��E��"O�Й0�(�Kԍ$�v9�&��yr���j�r1�׀I�"`	&���y���6w9�6�@wN��	0�ybgל?#�xaCjV+l�D	���y�F�i(���	8g	DD���<�y�ɳ}�RI���u�������y��
	�Pl�w�B\&BɊ�	ܬ�yª
UR��E�S�
���$��y��̓(t�=��ā4�d�D�ޱ�y� �E`:�jT�('܌��O��y�Z�4��IB�l��H2C�N��y+݄]��� Ym�ک���Q���!�S�O
���o����K 'Մ͚�'��l��lM�0������h��m��'����ߵ��P�"C@�~�<i��ïS
t�x��E����~�<�烅$;����ŗ�U��2wo�E�<A1,#q�RE�e�؁t�شJ�MN~�<�5�G�en@;q+�>	9X!�m}�<�C��(i�qWo�7u�u�R	Vz�<q�o�1L:����˵H���A�t�<YQ�۳e7��D	_1{yF �@ m�<��!�"#6Q�G׈(��M�ao�i�<�l�t�.ɠo߆d�(`�d�Nz�<���
��&��Kn�跉�}�<��/TOnQ"T�q��BBR#�!�$�@K�ak�˓�]�ȱ�@̰T�!��2_9^ ;a�F<h[LЉ���'>�"��L�+ɲ1��囱a��p)�'E��y2�D�.2�(���Q%3�P���� 4��H��}��{R!>��l�V"O�-�P�D�[u��C1b*���{�"O�1�M�v� т�g�+;�� �V"O$	 ��aڂ����=Ђ B�"O�Ģ�
".�8m+����)�b\��"O@�Ԧ���E�+ݭzD�@�"O�ݡ5K�<E�P����2:qa7"O�`�u+�(����u	X�f�Ա�"O�A�ՄU@��(]���S�"O���S�D�F�9b�'��Z�*E"O��)���&~��bB�� �T�#2"O̴�j��241Jq恷<�0И"O�)�@@�>��@����@�\)c�"O�� �O�{�p���c�z��j4"O���&�4LmӆB�*8j�i��"Or����݃"�P����gĨ@!"O^����o�0�e�Yv�����"O�e`��-fWb%1G/�7_��"T"Ot��%*��qS�9�#�Id� R�"OR��H�8�8�a���M�f���"O�	��)#��\���|�|"d"O���B�,a�x��؁,��u�"Oa:wL�Ȑ����Ĵ�.�y���d�T�oH��#�y��\~D����*b�:ĭ#�y��E�z5v@��MW���WkA �y�	Φ�؉yQo��}�$�foS=�y�]�&E���� �@s$����y���u���"��}��I�)���y玄H0�Zv�Y-�|�3�yrc�'j781xEI׺b���H N�y��X�9+4�欝.a<
d��٣�y�����l1!�T�] B٩��[��y���kB�x�1��!`,��L���yR�c  �cT苠����y�G�25��s�I� ���4�H��y�(��<���{�Gճ���0b����y�_�}_ح�q�� ��L�К�y,�6|�Xz��R�x �����J��y�۲J;��[��]�^�Q�i��y�o�O��D�S�C7u;L�0�y��U�������;qBx��Ś*�y2+N��u��n��I�Ԁ�PybG ���Ɛ+'���5&�\�<���
O��
� ��7Z�lH�JU�<q2o�?9�`�" "5�d�Q��N�<)�&	�)랔���ܹ:�a�`Ht�<飡�/4����6jI%��n�<1�C~|���1tn�Q)Td�<�!�T nE��!ѻP��t��T�<Q�F�t�8������d�5�f�<)7�B��&FazR ���v�<��E�A�����=F�4h���x�<�u�d0�g���-^'^�C�I����f@;$D�M��b�>C�I�qy����H%�m���Oz��C�I���@�G?�����xC�ɶt��di��[�c�P�Z2oã �ZC�ɐ{�QÊӚ5b����B�@[rC�I���h����t��3�A+U^,C�	(-V�[P�6��͡�d��VVC�I�l\:���E=5�����1.G2C�I?V���Ɓ~D>�0�E�X�C�	�j۬|x#aN�M\2!��o	,� C�)� ��s�a=Dh��H3W�(�"O�T"Ĉ$�21j�<H;V�r�"O���c/�<�l��"i�48��"OPQ W+�%xSHY�⊋<A��� "OnȐ�(O2FL���cڋC����u"O hC��OGZ�=B���p��)"O��I�L3h���P��Y�[�{E"Ox�;p�ѣ
��4&,��&N�b"O�(c@��*2:Q)��ƿ|�qɇ"Ot��/[ }_~"�)�3=��qZ"O��K��)�([�Mq����"O�D���$38�`�'6�j��S"O���5�Q'H�h��5�]�5h>-K"O�Hc��>nZ��ʳ�X�g"�3"OLP��)WII��,[�,[{"O~L���_�,u�A��]B��s"O�%�fFD�J��h��a�'K��@A"O�1���jzhM�����T��"O��G�Mo|�ya�*C�J��i�"OB�{�LX���:4�����[�"O ����L/$tE���t���(�"O�@r�D�.��І͌�;k�I�""O���W
��!~)[�[<RS���"O���K#W�, ��	�a5�pj"O-����>T���t)�$\"����"O8����˩V,* Ѝ�yA$� �"O���i@-{��D��+	�8D�Pzv"O��Ɗ�c������]3t@xK"O,Zrn�\���$� z?H�Z�"O�ۣ�ː"���$�G53�2 B%"O�}�v�D/h�+��ߠ3.;!"O�R��MlP�f�!>�m�e"O8� q��)���8p��(Q�؈q�"O�����.3GP0���`����"O�a!�	:5ܰ�PᑻZ�t"OB�)t�vbƜ�B@Ѥ���j2"O�� "�1�H�e��Z{�i�"OԀ2���m���y���"O�Z�NA�2�$�x��Ͼ=&d �"Oh9Bc��m.؈�'Gu@|!p3"O�(�Iw�Hi���a*p(��A6D�kC�Ժd6�#�Ή	^��Ł�'D�4�Gk�'����B�<���2D��q��׌uv� �'ϔ.�M�3D���2 �[��������
1D�C�%�,ZP{�E�z!�`Q�,D�ԪP�O�2��3AL�!�X9��+D���˗�W�`!���H�B��@�+D�$	�/ơa�аRug�'�t�Q(D����>/�� ��`xh�l0D� �G@Lg�� r^�x��1Ao1D�����Y���Z�!lr��p�/D���R#J�?*|dHv
� C2� �B/D�D��E�7�P �e�4j��u:�+/D���S�K5W�4�ZR�� ���6�(D�Q���f_n�e/~F%��h&D����ޣmz�5 ��� �Ҙq1I:D���i[�)y��$E_�K��X
!<D��8 �L>�~�3V Hf�|��#'D���æ��:v�[�!ƄswD�6%T�:�#ܔO�E9Ң���� �"Oʤ��%��&jXpR'P*�8IKc"O<=��/Z�B8�H���S�&uB ӧ"O�8��%k��)&$D�xX4Q0"O� � څ"�\�����ᆺٞ0s�"O���b��(��w�0f�e��"OtIBf�RVH�P&��OO��"O6!9�ObIF@[���B⦁�y�Ⱥ��Xid��>H��0�A�]��y���T�����
�n�6|�� ��yr��!3W��j��Z�]����yb鋮uX��j�BZ�g6!�P��+�y�K�Yu�5QU�A�s���0 
��y��I�.|���E�D4c��A�E2�y2��41x����̸\�z�S�'�y�怭0�~��g���AHN�1����y"��7i��ITlڅ:�`��3$���yr,�n�l{�&�4ڪa����y�Ā
(��9ya�P�0�9�u�'�y�ۗ:��;F�V�3 (P�+E:�y�Y���RnY�*fl����y�V?')
A���@�D\Q��I���yR -b�X��K;�JUX K�y�+�MO��jr���$�/��y��;g��8���J�MP��F*�yҧ�RۄAY�G-H����+�/�yB���:=���q��8�Ń��y�耀>�1�'LǠpe��hX�y�$@|�sFh��ѓA��yg�`���ZKJ]O�����y�i�4D*:u��)�"M�v�j���7�y�E�)<�TmbNܵ.ɾ4���5�yr 5Π�q�nJ�#��Q�Py"a3�N�i�#�mn� ��J�<GI�* 5�y��F�p�����C�<1�U�����'�H�aʕw�<�e���}M�����A$Pʑ��Cq�<Q��ץ^�L5�'a�<���l�<Ѵ�G�K���Z��N�s�2�cgc�<I�G�p�d���.=N�#��t�<)t�	?PL ���(�<`�D�Es�<Y�E@�x�^	�UKҌ�`�B��E�<�S�J	B��Cg�
6��	����B�<1��P���"d+nt2a�]|�<��I���؈�Oۦ:���A�|�<�� W\���#Ǌסg����E��v�<aÁT�0z�� P
q�81Ӥq�<1�dF
|p��p*Ŕq�n,Y�a�w�<Q�)��(t�WeO�jw�)�g�\�<�t,�
p|҉���D�4Z�U��Z�<��C
�tl���ě9	`���QW�<9�&%Qm��Xn�x���S�<)�)�6j&�*���zP����N�<	��R� H��ӫpA�uXeęS�<���4a�ebE%	���ˆ�Q�<�#��*) �k�g^&=����.�F�<u� �Qp���c� S�:���C@�<���ru�yY�Ƒ�@�K�&u�C�	 6�k�L����i�C�O�C䉔q���!�Fͭa7�,�OދHC�I�uV���˲hd��
H<>�,C�
|�A��Tpb��Eż�@C���!�G�>q f�(�p�jB�	�R�`dBC�	�O�nX��.�v˜C�<�n)*S.3-���	@��^?PB�I3=uR���E��hn:����S��C䉨$��Y�4@X�� z�"G2B�|�.%�C�C&l���Z��N���C�)� �䢓EQ?���26gM�HH�� "O���dƆ|_�y�Te
;_1n|!q"O�WK/q��Ǝp�l QJr�<)��:t�c��L�.�D$�DD�<�Ս�;	�~,R�Ɲ	k��K�g�[�<q�Oٲ3�$HI�!BD;����<7$�)*��-��Y�+�<�2�KA�<!��Z$*�k�>l�b�9P,R@�<�MA�~n;s�f|B�C�IWx�<!�G)+a������1AѶU�K�t�<����z�Le� .)qU^�2��Cu�<�a˓ 
j���`m����_{�<�c�27�P�����0s���BI�q�<�Q���J[,��aŝ�uΖ�[��l�<�6�L��,m0w��X�VYyF�~�<9$KAO jPhPoЦ��Dq�P�<9ݼ1��c�� Y<�ts�#C�<9�hӹF�����&HN�)&��u�<�3k�R#���ߟv��M{#B@g�<��O�eB����]&aYT�RU��f�<���(}F�r��C&	�8`���z�<IS��08&tb�e�EM��ɧCN`�<q�m��Yk��z��@}��8JU�_�<�+��6r��"�T�����]�<q���#�'��3�<�T�HW�<Qf�R�@}X���nF�@൐�`MU�<��I�;G�� �J3a��P��H�f�<	��=1]LԠpׯU�,p罞!�䕫P��hC(ٜ%��ɰ��)�!�D�W=��R�@_�QT��XU�)�!�dG��¦������Q�	�!�_�|P\�BD�C���@�)ʲ)�!��^8�i!@ f΁"¥	c!�$
�� �A�ŏlX�Yp��,#!���0=`���&͝;S.m�Dd��I!�� k���kP�"�r����>.�!�$V
ž��dn0>\���!�)V�!�D�,)�hHT�Ϧd@��jbY R�!�t�~H�c+��2v�jf��}�!��A�T��)U�B�*��9H�����!��Y"Kt�ר�+u����ϙ�yn��$��<s���=DpZӆ-]:�y2��^8�u��W?%���q�]��y�
-��r���"v*$h��ɛ�y2Ň�|�RL $����� Y��yBm��8p襑sl��h�����I�y�g[<���Sk�>deh��B��y2OH�X�: �U��%[���(�y�Ʌ��t�۲)�*Z��0;�#Ʊ�y��O1I �IơFM1� ��߯�yB��<����$�Da����y�T=��y{�Ǘ�D�BF��y"�5 ����� 	t��83�I��yb�� �N�.��	����"�ڳ�y��+����c�$q>~z��X9�y#N�]zQB*jC$��'
7�y'O.
�#�
�c�=��	7�y�2�t����X��wg���y"���	,@uR���N�HL�qE]!�y"��~v�� f�R�oh(	�h�$�y�o�u��H'
2� �	�'�0�y�@�o���K��0yb��(B%ަ�y��X4J��d픤({�!1�K�y" K�dy��seҞU�n-ÓO!�y
� lQ��݊�ʨ�v�֠@��m�"O������'�P%�%DD�o!����"O�Ź�8MG�$��"V;<@�"Of�r�䒫�l�e��G;0ɑ"O~Pj�%iwP��@��(� ��I��P]����i����AsV�Ұ.�<`y1�[>������O�h[����S�huiŤG@`˳� >���JJ"���0g-JFײ!:sD��HOdk&�X�L>$�'9Y��9H����T:��G��G���*W�3X�4A�%AޤK��̓ti�O��$������F�oN�i�Z����b���4+0A���!�i>�$���'���xV�Q�0�zN��I8�@�Û&/fӠ6�	�U�|��-Y�t�d ��FS�P`ݴ'���"3R�ܖ'���O�'�'���z21iC�\>EB�ʁ�ɑGC�ć�&VM�3�X6,�J�i���Ͽ{��Ko���$�L�;����l�ʦ�E� C�����x������w~A�t@�4{�1�k�L�dK�(ɢ̈*%� 1 �	s��L	��?A��in6��O�#~n�-
G�eQ�������#��| ��ß��'ayb����ȴ��[?�	�%E�HO�7���'�(�O.�rhQ�F2��*E�ʘ]�HQr'A�<�Co�7(k�v�'̈�{C���@�*S��@K� �D �(0	P����X�F�2k̊��ψ�O ti�i������;,ޖt��N_�� 0P�+KLV��q�D�!���ڦ���g�ɽg������7a~���T>s��k�(+
!H�aݛfI�t�,O��ķ>1g��v���To���%��A�h�<!�  2DÔ�^�~�Ǡ�,#�� ��a���oZ_�	�����<A�����0Q)��?��BcωG#���E�_���<I�GpDX�� �h�)J<1�|��CÛ#�  `pN�C�H: ꋝ[R�"?�%&��Aʖ�#D �d�Xxap��;M�m�c��3r�~�A�,I<gd��ѦF�Fx�!�?�۴Px0�#�����Y�T�X8�jPlD��͟\�	[�IF�S1�~��P�I�A����$G���IE؟Ԓ,A�.T��[Æ�*,a��r�A��?�Ҵi���'B7-B��mZ�t���[b�Q
i�t�5���q��a��B�B��?y���
�L���:c>�Tb�)�#%�擩X:����,R7H<��EOr!�#=hX�{�
�FR2/JV��s����u�'��-�U��.-Ԁ�b�se��	!l]p�d�O���	E�����T��V%S�	�d�7�H�eά�D6�i>�Fzr�8��Q�ʕ_ �8W����p>y��i��7�wӆH�ьW�O��6�F�D�����Oi�7����	Qyʟ�O%Q�&��M���4d>�5aTk4 ��caH9j�����P
q���x����W蔻Mv6y@�E�o� ��k���M3�O�=�tH�c��OC��{S���@��̻��e�����X�Uƌ@��H	�f��x��˦;���ON��_y�����V��?�8�I��+Md8����~"�'�azR�O`{�䎖%Wj'<):Ф�M�Q�4*�4(���|��O���ʿYP�t��Z3vJ�(�LT� ��4'��퉏e~p   �   9   Ĵ���	��Z�:tID:,���3��H��R�
O�ظ2�x�I[#��C�4e��B��.�=H�n�,��x�$�#f?V6͂���H�4;p�1��\�I�$U
E9�`[*P��2A
��l�tD�UE/�7�T#<)�&i�Z%��MX�J���$[���DX���'e �jm�,6?i��K) ��6Mp}"��t�Lc��&q�N�3�jAg� ��
ry�.�OB�6d����9On��$J�)Q����Qa�dL"D�#
(6 ̋v�H���D�==�������'���D$�q��Ȫ�`����H(��%����3##�'(����Ð�> ub$��T�M��'��Exr`X^�'��E.��!���Y�P����(N.#<���>ѧ*�4e@>a����Ty�F.r��)�O�ڊ{@�Y�V-;��ΠZ�<K��F�Ms3�-}n�"<��/�G�ld"sf�|e�Z0�E9Z�p�>�Vn)�n�4�t�xEY�(۵#H��U%��0�� �'(��Fxbn��nfR�� 7{x��K��Y�0վ�a�:$"2#<���Ox�$��q�E���6[�ٱ���OB�8I<Yf�;t5���Q�I^��p��ZS?Q8�\�OR�I0K��p�"�Q�Љ�ޢ4�.���h~r��97�]��4*��ɏ1qࡉ��OT�qakHn��SӨ��
,MɁ���H��܄N�Q�����>%f߷&.T���	 ���3ǄI}R��j�'ѪGxr�H�s�NS;2F�� �%�y�n�J�  �O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!6�D�O���&�i�O��nz����j
0mb �(�Vy�W��%�McS�'���t�O���iWBW�V:O�И�F>���Q�l�
/wh�y&>OnD0bh�?�r�?�$�<����?�pD�1|�%8�#�/�0��gC+�?����?�����Цm�1�̟ ����"�;pp]SW��*����w�m��$���	�M���i�Oz��3�U�&&��2ª
{�U*��D�%������.�S��RϟL���oˠt��d����e��GM�����T���� G�D�'��@�2��=&���cD�N�v[�ٱ1�'��6-�V���PE���4�n�+sG8Z�-Yp!�u�8�w�O6�i��m�l٨�m�M~��\�Z��S�;�*��Q�=Ю�@���/,�n1��|�Q��Sٟ���ӟ�������X��Ʀ�v���Myy��}�\�{���O���OH����ܸ:��vƈ]}<�w�C�����'�D6�ӦU�H<�|���o���bCY_(Й��ԋp�܌�Ѐ_~bߏ�&���>s�'��I�9�*a�q!F�fEz���$�:���ʟ\�I��i>!�'�f6M��w�L�Ю+�����+I(v �jV&V�8�����=�?��^���ݴ(���(w�X�!$�8m¥iqEضv0�:%��(}6�%?�Њ��`��'����1  ��<m��3��[�L(��r1o|�����L�	��x�Iޟ��bT�U %��5z�I˛q��(�h�1�?y��?A��i�x�:�ONAs�T�O©9��݈g���Co�E,��]��Ovo���?���Y�B�lZm~2NM�'�NŹR$�A�g� �>��4��ޟh��|Z���I˟8����Z5���r�� �㭛�Pa2,p��\�����fy"Dr�Rt��$�<����Iׂi�s�ɱ~� �U����ɜ����Ǧ)k����S�A�
�0�7/��hZ6ܲ����o�� H:A<���$Q��Ӣ0�b
�V�	�!R��)�$Z!�����1o�y�	������<�)�ay��`Ә0���Pz1��l��I$5���	-e�V���O~Qn�`�@��I��W�0i���VxrQF���?	�4g4\�!ߴ��DK�)rde��'<�8�H���-�m��YV�T�B��IΓ��D�O~�$�O��d�O����|r�扳Z'�| A�Ěiʮ4hch�#T�V��%�'a��'R7=�D=)e�3L��EÝd��i�F�O���4��	Z��66�e�������|����&x$�p�l���l�(	��.�d�<���?9$�SѢ�1'�ىb��%:7Q��?I��?Q����T����r˄���	̟��7�� 1PJ*l�%�3,�x�[��ş�Iv≐h���"`Id�U�n_�o��4���+Ĺ1�PH~r�k�O�)~�P��c�o	B8�5-Q���?q���?Y��h���d�$oDX=Ѓ��6Jz&M�%��.���̦���k�埀�		�M+��w��c	�A��)m�	9�r�J`<O,���Ot������6M$?�uB���S�y�vL�.	�  �'v�P$��'��'U�'�r�'�����J/�Nmi�F0K�v�Z����4��]/O��4�I�O
|�W8;mX�r��E�tTc�KGg}��'���|��to��i��I���#�b�a� �(Ԙ��ihfʓYp� P!���%��'SL��A �)�@Ekf ?���C�'m��'U�����T�p�ڴZL����wDm�oG4+�~���dxL�8k���$G|}��i�`9mZ9�M���\^�P��BP=vlƼ�禋9R��c۴����t�r���'��O"��֪��Ta���t��t�r�8�y��'�b�'���'����W0D*q�կ�4آ,s�!R�p�x���O��D����k�K�oy�z�0�OL��*R|���7�B�L�k���z≽�M3����T��C^�&���Hg T�t݄0���Nč��
� �fyjw�'8�$�p���t�'���'�n�r��[,)�B v���d�'��P���4O7P����?a����	D9sN`�kR�'��x5LD�Td�	���d�O�7�A�|��ʛd�`u1�-��$
pY���;0����ɋ�x�
���l՟D���|B/JB4������L��+؈i�B�'J��'����X��j�450J�"���th2�Ї:Ĵ,S�� �?���j+���D]J}��'���@+/%�֌q���=����e�'�-)K������OI)5g�ɽ<��)�=Q��lS���KB��<9-O���O���O����O��'��-��/O�7s�}��?���M+�
�?����?	H~�� ���wB�Y-�f|����˻(����$�'���|��$��%T��=O� d0�f�	d�����5LjL2v8O��@4M�8�~|rQ���	���V��]���y�,:t���5�����	ϟ��Oy��p��U+�Oz���O l��� �jF@�����")��P�O �	����O���?�$J�9�L貢�;%�~,\��A�O�S�.cض6-AF�\���O�����H�9�K����A���O����O��Oң}��.|2Tab�I |"53b��9H_`Ձ�� ����2fE"�'c�6� �i�ݪrj�y������o�p��q�8�ߴh#���{Ӏ��F�m������xe���f����7;�*���ͮK$��#ʛ��䓏�4�^�D�O����O2�Dک,ײ]	��'c�>����C�!+��>��v/:��'�����'p���n�dh���3�EWb�$���>Aa�i�\6MU�)�s1g>�&T
�oY�h�(��3�߬�r��J*?��^?T�������$�f� :�k[�c�P�)�Iu�����O��$�O��4���@�F.	�Y
RS��� �0�@��	�y�h`���
�O�hl�?�Mk'�iY��+s�E�]�xH��+�}(�Fٻj�曟�����k����i��(0�!IӼǒ�a�CĆL�dy��:O6���O����O����O �?����^-�7�PC��k�O������T�ݴj�J�'�?��i�'�Zz���'2�9k�H�,�،��5�	��Mp��|2U	���Mc�O����#P.�����o����&��#?� R�5.*�O���|���?A��(���AbĜ/�F�zJ۸/�L�0��?q(O,4n�O����	��	W�4i�d�\pB$��[KLİa����Q}MӦ�m�?��S��ȹUi8}ґ���:8xñ��e���Y�+�:tʀ`�O�)�2�?Q�d'��B�1\��q-�*->���F��>=����O|�D�O���)�<���i'h�ɖM�.t���H��^�"u��l���'��6�:�	 ����O������aI�c�*�G�,��Ģ�O���I��B7M6?!GjPL����wyB�T_ժ,��k�Nv�h�����y]������4�	���؟X�O�V��f,ܛyz!��Q�"D�i��rӔ���A�Ov�d�O�������]_��<`�)E��pcĭڢ
���ݴG���%��iK
M��6�h��y��6&�f���� sV=*��}�xcba�I��`�c�	My�Oib ��<,J	��L])t�
-��DwQ��'��'��ɜ�M�6�Z:�?y��?� }�T��f�:X��r挹��'e��S|�v�m��<$���gF�ri�xI�"(74Yp�3?�l��bަx��
Nv�'lݨ�DO6�?IWƌ��� �'呴C����'�R2�?A��?����?��9��Y�fߠ2�ƥH���4�u�v��Ol�n�{t�'��6M6�i�I��Β@������>�J�Cc�g����4s�F�oӺXh�$v�j�@2���&䟔�閤�Mx�9�`�^9>��� i|q'�������'��'���'w<���#T5���X��N*0x��V���4Gl�qJ��?������<� ����Вl�2~ �[�g��0��l���S�S>(A0$�jZ�2נ�qǠ0����Q�^�$�b.88;���OTI�O>-Op�9GgF)S�0ڔ)����P�&�O��D�O����O�)�<���i�X�p��'S�T�%]2g���b�

�6���'l�7�9�ɔ���զu�ش,c��
��Eb����^�PK�<�A'&z�� �i���q����O�q�P�.޹��e������h{垾B8�d�O��D�OJ�D�OR�d'����@�d�0>[�8� ��4�|�I�$�	!�M����ߦ&��*�M�!C�
$M�t�@a����h���Gy���Xn�D6�"?U�R���\��b�7$p��y�#?1իE*�?	�-)�ļ<�'�?Q���?��W
a��1g�)�уԅ��?����$[ئ�������I֟D�O������]<yp�aG��좹c�O��'��i�ؓO�S�1Xq�K�	_��H��^hx�۠ʁ	m�fSPe!?ͧ�$��˂��W��("��m(�P��)���y���?����?	�Ş�����Rw�ĲS|�BTC��zt(R��/y�L ����j�4��'���fJ�T�)���	~ n���V!�6�����`2a����'�E�q���?�&>���V27t�yB4G4���2Oh˓�?���?����?���;>ժ������4�/.�HoZ(�������	A�s�<����+�鑤a���p��1
�bek����B�2�iFܓO�O:G�i���!�����͕}\��H�æ��O]��P���A�2�O���|��j�<a�$@Hp|饏�
�0�����?Q��?�)O$��	< ^���O��`��|pw��.D����@ܛq)�tk�O|��}��$��3f�	t�<���#�&�9��??a#�@�yr��#3B�/��'}q�����?�R�N	t!\)6Ҿ! du��(���?Y���?���?ы�ik>=h���p^��s�� ��,jB�O@1oZ:l���	ܟ�kش���y�@V�l
m�dɻtܼkĂ��yp�,%��ۦ�
�%_����'}�Tkd��?m
ч	%cD�0	G!�;����s��e4�'��I͟d�	ϟx��˟����<�i�f��+B4
�k�J�V�`�'�p7홞,T��d�O���5�I�O&�S�\ ����Y]��Rp�EO}��v� �Io�)�xl�� ��E��&׾x2�@G:!v�MI6�U�]e�����1e�Ob�!I>/OJ	��
�X8 ����K���:3��OV���O�$�O�<i"�i	PUa�'�]�PA�>����]�B[ ���'!P7�7����$����
�4Ǜ���cV��b
AtZ���HU�
���i���"U�F@ZR�O�q���Xt�����lj�XI )܊ry��O����OB��O��D6���T�����T�t��fl�5{�D�	؟��Ɋ�M{�#A]��du�B�O&�0.��e'>dz�$ VE��i�M�����lz>Y{4'J��-�'ht
'�E<h*PbvK�
mF�+���3\���'f��Q�앧���'���'dJ,�Z?9:qh��=����',rP��i�4=�x���?Y�����10|��h�4\��U*raY2v��	���d���ڴ ]�����bAD yS&*G��R��
#_�2����;@)a�b����v�R(�;P�'���e�9O)� j�D��C	B�2�'2�'D����D�'�Bݑ5P�ȫ�4H�tH�	�I}P��dG�\��@F�
�?���?�M>�������%�2��,&��ڣ�E�YÜ|	`�0�M��ic�1 �i�$�O�l��g�P-�̺攟4�&D�IF �M�/x̃CMo���'��'Eb�'	2�'��ӽL%��H�"
�l������7��*ݴ,�@���?���䧶?aѶ�yGG���,a��Ҭ�'FA�t��$l�|�&�����(�nr���ɺ}Y�����E*LӀE+ӣ=A*�I�:@\��D�'7��'�����$�'�0�Z�)�.c��s�Z�]Q2D�'�B�'wbQ����4~�=���?��7��+5��I0٪��_�]i���>)�ib�6��H≥P������Ty���T$xK(�#p�J�W�1��T�|�5�O�T���`��=b���#z$�3�N+2]����?���?��h����M�8�r!AY��@	Q�G���$���Ѕ���I��M���w�l�K�>/X��X��t�'P�6��æ�#�4?b����4���193�-���5V�
A��hP���B�	˸�*�B%�d�<ͧ�?A��?���?1�%�1y@��ir�Ӯ4��y���H�������������I��(%?�I�-I�}�!�u�`	+���^�ɪO<�o��Mc��x����k�"��EŘ0m�B�5��V�9U$�)����3N�:��V���OD˓gfx5	r@��,Q���rʃ2~����ɇ�M�v�+�?��G�FfKJ6>�^���*�;-:��/�M��Ȭ>i���?����*��W$_�hp��@�Y*,��U$�3�M��Od���
ĩ��d���w���3��@��'\�]Bl��'��R�R &��Q�
p,�r͋9n0�I�q޴7��u�O�6�,�$�'ws��R�DÉP�r-K�bU�|�6�Or�d�O�)�32�7-0?���՜S~����j��$�6,�@��6	&����� $�̖'�O^�*�K�6�^�c�F �*w�Ɂ�M� �����O��'�����,
$)q��b���d����'m�ꓤ?1���S����*BHK������\%,
�\��!��%�<�'t�	~�I�d�2ȉ�bY{�T�@��G�BC�	��M{0�B�*5Tő�!�2�N ^X\��o��Ċ�1�?IZ�\���و�BA��V��,���Y�qC�)���`+�����9�'�P����bJ-O�*`-�'mʍ8Rd��$��9q?O����=���x�L�:��Ì�@
���UP�����[b�Iß����yG)��m1@p��c^0e�($��"5_��'?ɧ�O��}�R�i��d܄���U/Z�@�h�r��Xp��*�'a�'��	؟���6Z@�0�`E�f��/�Ow~���ǟ��	Ɵ��'W�6M�~�6���O��$�/:V ȃ��J18��Yp�KL#G���ty,O���xӆQ$�\�f-N���`�D�Ό4.�:��"?�t	
-�|�r�U�')��$�?)DgJx� � )L].|"��ŏ�?!���?q��?���9� ��m|~��
�9�y�ׂ�O��mZ�
�`��	����4���|λoY���"�27T6`�e[��ϓ�?q���?���*�M��O�س�����f��V�
�*�kZZ>h����l$�';�Iɟ��	⟰�	ڟ��I�R�T��ŋ?B!$	e��x���'�p7-E=���?�O~�]X��K�a�/����T[�Q�U��Iȟ�&�b>eP��Zke��O��o.ҍP�Y��|4o����D��2�1��'X�'��I�60�9q���h����%'�N��	џ�������i>��'K�7m�9l&��D�&�Շ#
' ^��a��.r�p��*:�V�|�Odp��?���?a'��Q�� ��+JV�A�c�WOZt��4��$�5n�i�Ol�O&'�*U�$q3��8N0{d:�y��'�"�'Yr�'���)P�B^qX%f��=0�����?�5�i�����O��r�p�O���'�}��q ͂K�4Ey�8��O4�4��Dswӌ�c�&�鐺��Ql�8&���� ZO1@��OT�Oʓ�?��?��!j����Z&���i�h�`Y����?q)O0�o�Z�1�'�B]>�1��ЎED�i�0�ڤ-�0`�G,b��������O&�D&��?� ��H��Ϧi�9��F5(�8��a�
�4F�!U�cӞᕧ�$h?�I>iUB,�F(��&�2 (B|��]&�?!��?	��?�|�*O�elZ�=��(2��T�X����U�W�u�ƫ���I�M#M>ͧ8��Iן�Hg�I'8��xC`�ݻk4\��.�ٟ|�I�J�@��F�=?���e	��cy"[!�YP���x�P��@\��yQ���IğX�I��I؟��O_�H�W�\4
�������+^1�3_�Mk�_����O���.�$����2�N؃���!j�<3aBېY	�-���('�b>]S3��Y	�	�HG^)���,G��aU/�/*W��ɢK�`�2�O�O���?i�D1D���F �A������]�p�������?����?�.O�LmT8d��	�����1�0c�Ȃ�G�����&��?)�Q��s�4=��f#8񤇟hvŁ���<.e��+��/�Ɍy��dy����x3�b>	YW�''����V� c��²L�-�\�I��,��ɟ���O�O��C11M��C�S�BHP��'���wӂuxgJ�O���TǦq�?ͻM�@��
SZ���4gQ�<����+��F�|�6�m�C? `z�8?��G:0��������4:g)�j���E�L|	�H>�-O���O����Of���O�x0gCN�zA\��ۦo�8�ŭ<9��i66b �'o��'��Om2�G�zj&II3���Np" �GI�5*�~���eb�8�&�b>�p���=7�ԭ#B /�&;7�'85*�{sm5?v��Ct~�d�*����D�G����@^�B�Y q�T�i4���O��D�O"�4�D˓A*��'Y"92�Wrt<آ��$� �����y"gӐ�V�<Q��M���i�
���!U�|��܈`țsh؈`�ؤEP%��O���[ ���d�w4�qBtb��I%jmB�G'�N�Y�'&��'NR�'��'�<�D�H�� �3�	�8[Q
�O���O�`lZ�gqH��P�4��{�VuK`��;˺�@��5!�����x�h`Ӝ�lz>�ta�e]��y�>t�f���re1�ډ(�-�P�a���U�����4�����O���]-���� �c�\̊��4����O"�2���PM"�'"�U>yv�J�#G�y�C� WM�( �8?	�Y� �I��(J>�O�>A3+�p�H� q����|鱖�c�N�$�Ĉ��4��x��a,�O�d����'�����ٍb2~(�d�O0���O����O1���e�F*��v� BpgJ�Z� �#H�$��aa�Q�Xz�4��'�Z�"���8$2��eM_��@D�n�6MGæ�r��rr��l�+�f����O����d&�;�J��SC�?q��Þ'd�	͟������	����Ib��(<&�P5�Ȩ<�L�6e�#Ɗ6��$6� ���O���1���Oؤoz��*�Ɏ%{�,:�߾RNrɨ����M�C�i��O1��|15lt��$@�0�s�>b� L��Ɍ�*��� �fw��s��S�ΒO���|Z������-^��`9:�I	���Z���?)��?q)O��oZ-e���	ʟ���f� �uH�@z��c���1W���?��Z������sK<��LʒJ�nY�dc�y��㴥�k~R��1��AqeIK��O��i�Iw�ܑ%`�Y�#K� ��D
�@Cr��'���'R�s���!��Y!���n�����O�0��4 �qi���?q�iO�O�Ή�r���j�dX�H���d���-�ٴD5����NE^��O���|��S�a��X�Ӄ�-�5�T��%��EQ��|rV��ȟ��	ޟ��I���`p�@�g'��d�"m���h�IFy�d�vh����<����'�?y!�N�Ҋ��Ԃ�f�R�)��  �˟�oZ3��S�81���B�C�|��h�/K8���A(+/<��]�U9���OPLiL>-On�B�e�[�BE� ���t�8�,�Op���O��$�O�i�<��i9�[&�'��<�$̔�9�'.+�Y�'�Al�⟸ �O��d�O���Z�l�tiR�Iؒ3��U���H�UM>��`��&��I�n���ݟ����R��u�b��$j��U駡��n3���O��d�O����O��$9�S�F��P��a�'��)˔�8�a�'��t���8�.�$Ʀ&�T�uNº?���A��]>59nd����e�I���i>�Pf-ٝt/X�J�NI�W@O><rU����m��D���هw���G�zy��'���'�ҏ�?n$`g,�?n� 5�L�.�"�'��I"�M�Lډ�?mf��$�|*�]�J`٤ D3Xr��#@b~B
�>����?�L>���M�sL�6��Z%cǍB���D)�:$�ؒ�*uz�i>���Of�O���$O��v0	T�̯>�i���O[m�Ɵ��	�b>�'6�6�Z)DǼ���^�p;�і{�< el�O��d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q6Q,��M��w�8���D|f�04ʖd�2�'�b�'�r�ča�:���O�Aِl&���@�T�����T�3������R��'����$�	Ɵ��IƟL�I�j���Xp* ��Q�K�(
�P��'��6�	I�N���O`�$4���O� s��~Hѳ(�
��aI�r}��'�r�|��T!�)�>)�%f(&v���ƞmK@�cɓ�x*�	<;�iq@�OƒO�ʓ��a�F�W35 ��d�~!�M��?!���?���|b.O��mډEȤ��Ɏ)���yCi��g!���rm.���	��MC���>���?�;�B��dG+R���+ʬ�Z!L�:Hv��'V�YЅ�RIbO~����F��@
\"������(>�ϓ��?Ї���Y�$1baL&�����O
umڎd56�'*I�֘|�ë8�����Z�M��2� � O�'�������77G����O�`x��37��	�M����mk�͗M�.9S�'��'��h��9E� ���I!j���td�7�Fx�eaӖ�c�<����i��h>��W
N1>VV��$��$cE�ɓ����O���3��~��B�?��H�KA6+�({��'^nD�۲fE~��D����O�[?�N>����jl�(��ގ}�H��ՄR��?���?����?�|�.O�oZ2
/� Ӧ/WsM~�!��_�g�V��5�J��	�M+����>���2v�] d-G�x�8�AŞ=S��@*��?)��1U���'���	V�Br/OƔ�� )�$l�5*�^�B��5O���?)��?����?����I��d�u ҃e���� :����Ld�p�B�#�Or�$�O���D�ئ�]<�n�0��,$�0��:H$�	ޟ�&�b>�1N<:���2rL��HĊu��PC@���F] 牬~�D�Pg�O��O~��?��d5�a�LF�/xP�舚��(���?����?�*O���	�y"���O�( �by9aU`�z13��:��$P�O�}m�:�?iN<!�G@�6!Z�C��E�:�d5�M�x~�f��&}�a��&Q,�Ot�I��$Qer��z���'mΤK|�h�Ê�I��'�b�'��ퟬ0�!��a���2���0YN~��0�ȟx�ߴlqƑ:��?�@�i��O�ʤB���R͆2�~U��!��l�DP���Y��M�e.��%�
��'�(��0�Z�?=��!VG�ҁ(�=m��J �ܜ/V�'n��՟@���L��֟���%�tY�!3o���4�A ^VL@�'ʹ6��}�l�*���O��󄜞RP��o+��eHsO i����'3d6mƟ�$�b>�Q&ˤ{a��[�����`�]�#x=����iy"��w���I�F��'�ɷAF|k�e�.T�.)(#����ڌ�����i�n����~y�'k�,���f�O@kP��<���*')-7�J���#�O0�m�W��Sh�I��M+��'��L�1e �u �F_Y��QC��@�����X������i���F����.�.��]�'�[ ��%�V�A��$�O����O����O��$2�S�^�5ѵjR,��)1��V�EhR$�	ҟ��	�M������Ǧ$�X��@N'�t��Р .�K��%�ēa ���O�4�P�Y���O(]�!Ǟ�%n��ڝob�5P��՛P&�E��2�O���?����?	������GD�=�H!vk��H:���?a+O�������D�O���|GOI����J�$��`uZc~�n�>a���yR�xʟn��@��w��5�p�ϐG޵ 4�F4���#��fn��|�&C�O6��K>	�e��B�j���+k[�h����?Q��?9���?�|r/OЌm��H^<I��_�C5xxa5��#�6)Ia��ҟh���M��R��>Q��i���QI�D�3Q�&P4���D��O&6M?S�\���H��*�G��$	_y�J\�E�	ct�}��!�i-�yRQ���	��	П8�Iʟ@�O�~��񃀉kq*���A�;.�i�np��p�bM�<i�����?�Q��y�X:{�r�!�/��~��n��%.�o��M�7�x��D��(*��,y�'�J	�%EL�5l���N�R5|	A�'W�X����)E�|RW�����JR'gOr��VAN$iࠆ���� ��Cy�H~��	;3g�O�$�O�J�S�%\�2d��N�@<�a�0�ɇ����צ9�ݴq��'�L1�ɝqK�ఀ���F'X��O��ea�1�
�x!��Q��?)!��O�B��CJ�U{%��-#���5��O����O:�d�O��}"��v������;�v��vAE�&N8��j0��Q~���'4�6m:�iލ�#��.�%�[*X�(X��������OT7�¦�pC �?��,�`� ��0P�l�7tjHY�ŋ�T�z���a����4�|���O����O��d�'E��D�3'��Z�H��w*�j��\�F�F S���'q2���'�xd��:l�9j����S��PB0j�>Aa�i��6-X_�)�S* �,��!��q��$�,N'��4 b�1HJ�L8
�p$�O��hJ>�(O�h�1K��*u�!$�95Nq�(�O>�$�O�d�O�i�<	2�i3��
��'#�d�U"E��p�� �D���)�'V6�6�����������۴g�� ؀�IWr�s�����=rA)�>Q!��� {T�R�1���	��ʔ"���0AxT\`���%�2$��5O^���O ���OP�D�O��?�d�7?�Z�8�ՐZ�)�T���d��ϟ �4�Nͧ�?YP�i
�'n؊g�ĩQ �"en�)�djb!��L�i���|�φ�;�F��'k���M�64@yh�)=�H=��؁�q�	�v��'��i>I��؟d�	�lt��Dk%t6TP��^�#�P����d�'�6-�3��˓�?�*���{�GM
i"R��s�U�v��5��X
�O6�lZ�M��xʟ
�*�J�'!H�T��!x�mB&@/?�f�	4��DD�i>��c�'��T'���e.��Vh�1$�O�V�kcO�֟��Iҟ����b>��'(7-��A���9,�-����%�Q3.��̬<a&�i��O���'I6�D�N�DU�B��WI��y�O;�Mn���Msw��m}ޥ�'�.4#AL�?���&m�󦓅PiSB: j��57O2˓�?q��?��?���3G�ʡ2���:i6)�,S'�u��i�bQ�5�'���'���y��d���\�[��1�a��P۬q���lU��n��M[D�x��$���m�`��'W8U �F��Xl�G�н*�ϓb1Z�pi�O݃H>1(O���OX��$#E�,�hjE:M;�i��O*��O�Ī<ᒴil2}+��'W2�'��8��Y9tn�zE�Zt[�d�K}y�(�l#��NV�%Zd'�kxhMڕ�[�'�L�'�𼘤j�e�5���tSٟ���'�|�C�@�0(<�JT$��Ģ)	f�'X�'��'��>��I
4\�l����bOS!J��I5�M�S����?9�j�&�4�t4��'�<^褠���b9
��=O��o�<�M�D�i"���ٷ��$�/98�3��jxB<���Д+�L	�`f��m`f����J�VK�0�.�9
�yF�<W�����%[��a8⃖�yH6�t�M�Js�9`0J�<>�DQ���m�vp�ϔ8�,B��LϊQD��$��e��2]�H���@�[�恚���4OD��A+�+B~�T�ݣP'���H��Z��C��U�5㚛/�����N��Dn֨d�=X�e�7Q$���eJ6��
όp���8Y	D����=W���M
���s���Q�l�0�&����Q�2M14�pd�s���F�,~,}�)�)dZ�8�T��v�4s�̙7-���'���'��$	3?ٳi��H*� ɛ|�[6��I�'kP�������={���"�BT@Y�b"דp���	&?F6m�O��D�O���H�	@����,�<���t0Ȁ��:�M�fku�����$�
y\�hKDH%FW��3'�)&, �nҟ��џ`�@��ē�?���~�#�)T>�]r!��uĄ�@�F���'���y��'+��'�P���!�,X�t���~Y��k�2��݆y�>&�p��۟�$��؁E-T���B��蛡{v�Z ���<)��?	���H�@�0	�M�WH e�1�N�wv(���
P�ܟP�	\��\yrC_X�2ĉ�$ĕA -�j�|��1�y��'���'J�	?��Aa�OE�����#�dI3���Z��M<���������;��	�"�6�s�슘�f��V�H�|�H��?����?y.O��a!l⓸�XY�֍�Mm�NB�-D�eP�4�?������<	�O�L��O2���/�\t��m��DU$ɘֶi���'��	h��)�I|R����G�I3��RT�W$1ٔ��%f�)S�'c剒��#<�O�H�B�k��d`2���l �<p��ٴ��#J��m���i�O���T^~�	�Gx��Wg�e�%������M�/O>�;��)���*>x�G�	 ��e���{G�7튵s�H%o������џ|���'x�귫F�X�"<{��S�\�h02�zӀa�6�)§�?qT#ޭ^8V�X"���<��,�-��V�'J�'N��5I7�D�O�d��@���(_F����ł}�83#�2���R�&b���Iʟl�	�"���y��܍	@Jl*`��8Dw]��4�?���)�'r��'sɧ5��Wk�����m �6"`� �ʠ���əsY1Od��O��$�O�*6�r|�m�DFP����A�m�,���䟰�I˟$��N�	˟ ��A��*Ï4h��cW��F��Qo�.���?����?�����<�?9����El]ҥ��5��a��*�,5��'�R�'%�'�BU�T�!�}��A荓'Z��ˤ��9��P�`���\�Iݟ��'�ց�Op�&P*�F�1H
E���c�	��H��7M�O"�O��d�<bb�d��]�}z���zʠ9!��D�Z��7��O(�d�O����"{��d�O����O���#),<I���¯)�ٲ�+��%�<�$�O0ʓ0���GxZw�$�ȡMV�04е�����1"tP޴���1lZן��	Ɵt�������`JP)K�;A�Ar��6a��=���ib�'��b��'��'�q�FђWgӼ��P�I�_^�dB��i��T���a���d�O��D蟆8�'��ɰ:c\TX��@	5�NX�DF��4B��ٴޘ �b���OR,����$�� ҉̎|3>����¦��ܟ��ɛ3W��@�O���?Y�'`r9S#g�q��8�$�j�����}�cG���'b�'5�L��|��sv��]�F0�cؿ%��7��OQ�+
H}]���\�i�͘�+�
����B��.@`q+0�>��L!�?�)O���O��<i�Ѓ閡q�'(t�F�`V	�#fm�9�^���'M�|��'L§9� 
�ǯ]�V6԰��͛�T��P�3�� ���?��?a-O�1
Q	�|�!'ԍE�)p�˗3��y.�ܦ��'�2�|�'����O�����$�|ИU� B�P8PtL�)��������쟴�'�H,�æ�~J�$�����[�Kմ�����&$6P�&�ibB�|r�'c��ݾNPqO�)��@�]�D��a"8�Sǵi��'<剪.��Q��p�d�O��IV�(��^��`
y&��$�P�����z��8���4�.o�����C64�L9S�@��M�-O2��vJL��]�I�I�?�R�OkLəG�T�#��S^~D���.=���'b���sx�OJ�>�1r�צsY�QQ�ԬG���@�"d���f.����꟨���?%y�O\�{�f�Ab-�9P2ii�	A�������iN<�d)��ӟ��@��i<��枂@6�%�7���M����?Y��|�ZYb_��'x��O�}�𫊾DPz)!���:`�lzQ�M>����?������Ծa�tՈ���
���ռic2�=9����D�O4�Ok�����j$Dh�Hj��U(f_�		�b�d��֟��	ky��Բj�3�EG�9�!iFjՁ��!j�>�)O��$0���O��d�7Ry���H�\=R���K #b����5���O����O���^���3�Fa���{���DlT�?��4�CU���I���%�ؗ'0~TaR�'X���Z��(���L�)��:�@�>��Ӗ�6�'�>l*9K|�gM];I�ָ�ڝoRp��"K�@��&�'��'��I�����_��{�<�A��9b���i�ad<6��OPʓ�?�V����i�O���k,��D�5��x�	AS�ǵt�'���'�����lW*�����E�4B��IP#b�$�x@��'��	ϟ�w/�̟���ܟ��	�?͔�uWaP#̴BU`%=��t*�5�M��?y �1����<�~bЎ�(	&�5�� ��8�$�b�ئ�Cv���t�	џH�	�?�����ȨFQn�����d5�S��\%�6xm��9~FͣgC9�)�D������C��(�QM��B� P��i���'"��� ��)�I�l�dm�8O��,=T��)������'�
��.8��O��d�O��uk
�Jy�e3tI.D����E��I͓u�,��M<ͧ�?�I>�;��	�m��'a��*u��ts��'(R�*C�'7�	����	��ؔ'������=W��qb� ,��O����O6��?�*O�͏!Y�1����"��cԁM�Š�D�<q��?�����䉶r9Χ��m���D&2]�0�d�] ��L�'&��'��''削F�Q���m�v��iG"H8	SO9+�굱�O6���O@���<�b'DSb�O�=
��5�`g�2q̉�E�m����&���<!"B�:�?�J?M��֘|�F9{!��f�����y��d�<��i��� *����OT���\�#��9�P�*�fF98�\��xB�'q��)"�i�y���%H�5�F�����q�f4p�i��.}�����4O�S�<�S����ݦt|���H���)c�*?7F��^����#��1J|I~n�o4X�N���X�)#ig��"bӜ���%F��e��䟼��?e�N<�'@�2��	"r�ǈ^?u^��i��(���'��^�'?��pz�H2t�R�z�Ċ�6�m�a��M3��?��'�H�מx�O��O��tkC�%p0����3��AZ��i��T�d��T1��9O��$�O�ЭP�*ݸǯ��7r�������q��l�<�e`N����|*���Ӻ{#��.ta�]Rp�hq� O�z����P�����O�d�O����h�NA�u���3�-O�ص���Ƕ�'��'>�'��	�$�h{g�Ԉt���q��9\�)�QG��� �'�"�'��P��RT�����I��+�N���e� 2��\���9��D�O���2�d�<q�jʸ�?�t�Q9z�Ѝj��2D(�5�ŘG�'#R_���	&eVV��O�"��y��=���N܆�0
��4��78�	����>Eb��e-?��C<cU:$Z��S�7��J���ʛv�'��V��Bw�����O��꟬UY3D@�e��ySg�F+dP��P�-�k}b�'4��'N�,�'�b�'	"ӟ�iS�w�r�ę��n�$�M[+O޹�t	�ᦡ��؟<���?�+�O뎔&Z�b��
s5���L]fڛ��'CjV��y�L�~Γ�Oqpрd �#a)z��".M ��޴q8"�A�i�"�'���OĎ���D�pUحJ7�վm{���'�!G�!o��b���	W��{���?��-A�� s�2LtM8�1M��v�'hR�'�z�)&&�>+O��$���j�C�c���0R.�A@ĩ2��>1/O���g��������֟�P�(�#d�x��ܕ&��쁐��Mk�f͎�{�T�h�'��[�l�i���BMy6��0Ç+*��>��NA��?y��?Y)Oj!9���\p�A�fN 8�b�2%�9o�8�'{�Iӟ<�'z�'LlHO�Xu��qΑ���,^�ؼ�O��$�O����O��h\��Z�6���S��ä<P�`��Dd6����i��Iӟh�'���'L���?���������D��Z$KV�S53����';��'�rV�hj�ɋ:����Ok�gt�pa�Q�<�j�!S�ſrp���'0�Iٟ����0�pe����y?� :�I6�[�$]{�j�? A4�#1�i���'��I�H�脀����$�O��)۴_lb�1��j�T���ڌu�v�'���'�B�Ν�y��')�	nz���x\��)�]�� R��̦e�'����2ed��D�Oz�d�V�ԧu���!� ё3�I���;�L��M����?�&n��<1����� �ө1��� F*�F�ط GW6m
�Ho�֟���՟��Ӽ��d�<Ѵ]X-�!��(-tu�7��).���d"�y��'�B�'����JT�1�a���� �-*G(�m��	؟�Rt����d�<����~ҁ�#nS�� O -Y����M3,O����f��?��	��x��#n�n��D��&0�@�A��0�Iaڴ�?Q�&�t7��Vy��'���֟�ز|��܉��	H�.q�uJPA���Eϓ����O�$�OH�3`�M@�� ~�Z5�*����!���4}w��jyR�'�����	��h�c�'�b����I۲���Y���pyR�'K��'��	-}�"a��Od��3���@[H A�iƦ�@�4��d�O`ʓ�?i��?��+U�<�gh�
/������
-�52�+J�?������	̟��':��XaΥ~���/���02�X)�t���a�ʄ获�M;����d�O����Of���?OR�'���c�X4L��I	�d�9K�F��۴�?!����@�\w���O[b�'��$���i�
�X'.����ڇ(i�꓀?���?Yǯ��<!���D�?)�灨�"� 0�F�'嚭��g���Mh9��i�|�'�?��'Q��	�r�m[�O�V�`�S��˕5R6m�O���I#Y��$&�$0�ӱ;9��c�-Բ,JR���l�= 7�G�L��nZǟ8��şp�����'=�@�M��}#&4�q�	)���djӂA��<O��O��?)��;a�L ��ի|`^y�rڅߴ�?q���?af�L�'@��'��Ċ;�I#0�֗ ���� ć&I�&�|B�?r����D�O����EQbFB�9=�8�"jɊCpo������G���'�|Zc���+�D[഼{��	}���Oт�5O@��?9��?	ɟx
`əa��Y���P�jQ�� �͌; n�O����O��O����OJ�/	�r�b-�R�&8u�$��e��+���D�<a���?I����	ƾ-{��A&z�@��] `!��F�J�O��d7�$�O��$-W��dG$�E1&s.� ��_y�'���'��X��{��E��ħaQ0��0J
���v�Y)��ʀ�ix��|��'y�	�y"�>�E���O��ݳ$�ݼu�@i������I󟸗'��5�b*�)�O����&RlM��GU�I ���\?AH'�4�	�����ퟬ&����L�����F�~���!'�ݦ*4�n�^ymϥq307mWo�t�'���l3?Q�7A��[&�U�j�l��#Ҧ��	���"�&�͟�&���}z��� 3�T�z��N�K���ɱY��	xP!���M����?a����x��'L�f��̪@(Wh]K�d=�+���w��O�O��?���7wԔ@���]� b����+X�;GZ�i�4�?��?����E�'B�'�����N���4LR>&��D+�2+���|�X��yʟ���O�ā�1�Р	�jE���
�⑩?��`mZڟ�������'"2�|Zc&��##  ��X����S`a(�O�h2��O���?���?q*Ofi�$�1:�@Z��S�(H��D
K"d$����̟ $����̟X�p@�꽱 ��c"�4�7�6a#n�IZy��'���'h�IdX���O[ �G�Kz �x����q�ɉM<������?���.Ȉ��u�]���<X�P�W����R]��������zy�j�J��� �V�J�R���ǉ1T@������	n�������4*��=y��,H�8�qw�
'o����]��a�I�P�':���!6�i�O�	�,d PqsU�� a*ʙ����{TX�'���I��yb�a��$���'A����EԞOk��%��u�4oyyB�ǲx6�p��'����'?��F�r���B!/�vd��/	B}b]���I]�S�S�-����1��CP�%�`���q�6M��w6l���O����O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J 3��b�h6��Op�d�O�����D�O���rG^i��	�C� 9��;��LN�'sb�'	���b��ʘ���ͣS��Ԛ�lT��!0$ &#�f�'��g�/=��'�r�'���'yZcn�93p��+7����Š
I�dߴ�?��4����Vj�S�g�? �HD�P2զ�)�,X�3��a�i.Jls�zӴ�D�ON�����T'��/z��e"��
8�>��b�3d��(�4'$)[���Ϙ'pb��Q�
�#�ݏFmʉ#F�N-Za�6M�O����Oh%`Bk�<�.���d�����`R�hM27�۠a~8���2��'�حb�	.�i�Ov��OLR)F��`�J�4{����ئ����S�R)�N<����?�N>��~�Z��M�z������Q�c��\�'"���y��'��'��I�����OI-r��(�Tnν]XX+��ē�?	����?��*<>�IT.Y^�h�T�P��Ȑ����I̓�?a���?�-O�yRB��|�e��9��x�g�J�{]\��du�I͟�$�`�	͟�hp �>Q0��6�����P�=x(@��b�r}��'�B�'z��|�b��L|�s%�1c*�ɉgvNAPէW՛v�'u�'b�'".�s�}B�>�!Qr�N( X�$@V�A��M����?-O2훐aYM����(��3aMǋUTn�����D�)J<���?	��S�'e�i��a��)��K�C�*pCfEZ�d˛&\�| !���MC�\?E���?��OQ� Ą�?���ۥ
}��ib�'F ���I�E�������ø��q�<Q��&��0"�6��O~�d�OT�I�[�e�
�AO!-��Dk�*��(þi�Q��d$�Sɟ����(&EpKG`اI��Y3��N��M���?��7���&���O�����p�I)5����t��W��c���BK?��������r��ҳM��Ha��M�)@�ՃqDE��Ms�]o�� U���'�bP���i���G�-l�����h��/H��Ia�����t�Ġ<��?�����$^*1�L���"[�Pɰ�m��9�0 B�_}2Z���ISy"�'�R�'�� �H"a�@�B��^=�uȅJ?���?9���?����V���l�'z�6���N�4�^�У��$V�&5ldy��'��I����ӟ�B�v�d���`*�b���l�Y;�*¥����O����O,�Gw^=xER?y�I���	�
�.�*� \譢�M��M����D�O��D�O�$Q�?O^�D��x�dM��2��
�&,'�5�lt���$�O��=��a�P?����H��1W6 ;MJT)v��>+�p"�Ox���O*��ʃFD��'��?�"��T0t����3��yh��S)g�2�1��+�i��'���O]�Ӻ3�#h$L:�I��δ�!�ɦ���ğ��u�q� ��Zy�I�381 �th�J�~t M�.`�m� ]7��O�$�OR���a}2P� �!���h��*��C%U��u�ڑ�M��<�����$-�Sߟ(���H�!dȟ�P�x�hʙ�M{���?��f�=�wP�ؕ'�R�O�I��*�55��2�*�%�@�i4P�P0&n��'�?����?��
#)
ܕ�����JܝH�6�'�hBo�>�,O���<����Q���Tx�gE�r�AI�x}�E��y_���	ߟ�%?�B��>UKpS��K�:�JH@�ꐃ^��	H�O�˓�?�(O��d�O���K�>m9	¿��p!�R3p��z�<O&�D�O2�D�O��D"��a���x�®B�3�$�(&�7rQ�J�e��M���?���䓕?�-O-���iL��P����o8�!
�4��L
�O���O4�D�<�aiF�C����Ps��T1��2���7�V0X'���M#��?q���';qO��(!�&��]��U)�ZLX��i�2�'|r�'ª��q\>�'��T-�7
���D��#㤕 5�P�.O��D�<!��Ko��u�+��A�5#b�ܰ*Vnύ�M����?Ap����?��?������?��/F����^UZ�q��(.#�o����I�"U�#<q��4k3pUqF!L_��H��S��?����,��s���0=	�2�Fm3��V�"���[�<��`�5?���ԭ
�.3Y��[�0k�	S� L
Aɂ�J���.I�թre�?+9�t�U��2t�2Q^�$C�����U01�`)��DV=��՘&�>LpU�����ZLuq��X�2P@�P:%�0��a'Q!ܠ5X�� *d �#���[4:��g���Px6�Ĕnv��k�
�?���?i��Z��.�O��D|>��A(V�S[��	ďRI��\���N�8C�	I���P��͘�-A�k>����D���N�� �D�e0�� ��ph�/T�.NH@���Φ�#��9-$!4�E���@J<y6hFW�¨넅R0��[2�G7J�(H�	��TE{2���M��A�14Ԕ���bM/'!�֟pt�-;���<<���Ȅ�p1O4!�'��	D=�aB�O �]�2mb�0��+l�$1�V5^`�$�O( qi�OH�z>�I���9'�ڝ03�خ�~��'�2�Ѣ�"o^ � "O�p<I&��}��� ��K��Ӆ!/�k׃�}�����a5H �x��]��?�����d�am l��/�;M��&T�	�1O���DR�
n��0��F/�r���9�!���!۲�
Q Р�0k��~a"��̔'�~����>�����	��U����Q�KG�-�샞q�ƼP d��X<���O�`��)d�AI��ͅ0�?�O*�S�4mj��#��#�!��o��G��'�
7	Ҋ8�i��  7A�>)����'`�n���՟5H��d�)}b���?���h���� ���R �\x��נJ�<(�G"O�9rǃ(l%�1�դ�,��P�'�#=i��Ɉ!�Ȁb��x�0/��W�����@�I<M��T*aŎ����	韄�i��F�c�N=b-���@E�_t$�A�^�L���@�b>�O6�@��*2�$�E�a��e��tc�+�O6��Ɇ�и��a�H)���D�A�,Igɣr�������$ʒG��O�ў8���?np�⠅�l�ZCe=D�7e��(�jm#D$�.��kpM??!��)
/O&! #�ǰT��<�1�D�9.8��K\>����	�Oh��O��D�к���?��Oz�Iᇏہ;Zd���̆�]�D� ����x�k�&ɠ�x�E�)8������*F��@	�'Ψ��vC�3H��Dާ���@��!�?��o1t}B�N^M8��r��	o��)�ȓc��TKQ��p��(���X�dS�`�<I@�DP��l��t�I2Y=L)z�J֓x`>�kƪ	#"z`���<�`����	�|Bq�����'����^��YK�O��1��$O��� �Ĉ3m���0e*T~�1���Y:�x�C���?�N>��X�C��t�!��?D�����J�<���O'	���
�o�\�z\@b*�_<y�i�x<YӣI�_X8!B�P�"�,[�yB��&�듓?A+�������O�����0-q��;1�[I�=1�	�O,�d�*$W"����S
#�:\:�f��$UJ�O���*���Ɉ}�.��v��;F,�'����+[@x����٘*�>�PBI?�/2�X  ���U ,�LG�<kD�'�F0p���?1����OJy8$�D)7��$�p���F}����"O$�ڷfܫy��E�D䄽d2	S��'�"=��ɝ"i�)S����>\�V�M�.���'��'�H��)N�'K���y��N���8�cd�+ag �*�C7.1O�%K��'�(d`d&�/&�v!�eGZ�xM�{�� ���<����;&�p��)�="6�P� �.��'1�P��S�g�nM6T+&ܠD�!�kֵhC�I�9r@���F7w�Q:�+L���ߑ�"|"u�T�Rr*�c�I��u��c���72�+@��5�I��p�	ݟ��_w�r�'��	:*��:V&�#����1Ό@!����Onu[�/�B�6�{t�~���e�NM���'~$�G�֨E����#��Q�� �r�@�?1�Z΍�wE�C
z�3��D��ȓ`ߤ���v�9��ZB
"�I���'t�ŋ�m���O�<��	�5�L�5�F�3E(�%��O���� �|���O������'�W�+JXy:���2'�4�A�/��x�E���'[jE�w�ϭ���� #L����<�Z�	D�ɷM�x�It�˵{��HK!\�M�~B�I�( 8Z5�V�3YPc�x%�B���M3��A��0�⦭4 xٓ3��P̓UZ�h�#�iM��'��,s��0�ɯ,�|��6dI7N?V`Sb�w�^��	ן4���<���D�!+�@���*u,��P�o�a:2�Ex��A��uIJ!�ߎ{|�Id���ɾ��<�)��&.#x�[��� _,Ż��Z�;a�C�I	
��ȡ�����2U0!M������r�'�Ѱ�+U�4}�<�u듾w��J��i�B�'��n�[Hؠ��'d�'��w��!!3��:��Ų���E�<Q��i� OP-�P���_M�S=*�1��'Yl��RP�?���U)�I&�����B��	��ȇ�j�T��DU�����X�,)	ׁ�?�`y����'��"�i���'^��C��d�'_��'"��'t�T ��|@$"��F䰔btO� �4ƍ�EFe����r(�8T��p1��d^}rX���	@�t�CΙ^��q;5!̐\I�D0��şD����L�I��u��'\r�'B֙(�0f�pxD�63e��cT�z!�DD+W�,H�t`�]e,+㎗�(�4��F�y'�ؖ��h؞��5� "l���5�ٯnx�X�Q$L�R���d�O&�&���Iɟ,�?��_�K�
M��&�Hwh�`�$�]�'?H����0I"r��#�pd�%Q�c�6wfx�O|\m�Ɵ�'��*�ê>��[Q�5B��D��l�@���Z�,�i��?��b��?������n� ;B��#��h���#V�6g2��S+<�,��K�<����9%������)?� ��D��:�p�	�D�6z���b�1�@x��'�0����Uś�>)�N��$��Y��҇w6�=�� r̓�?1�S�? ���CƘ*
�D��jͩ4�Y3FOulڮXq&��$߮6D��RE,E3A���IG̓�MG�,O������v"N<A �D%�$�P"O�e�ņ(yL�����15���"OZ�r�$��a8�b���x���1"O^��s��PH���	��dF��2t"O،���^e\4\@R�ѩT1�t�"Oԙ˵B)s"&c6-��':H@�"OV`��S�eX h�Ǭ\Cx$z!"O�<b�E��3��\4��$�@"O�s'/�b|	��j՘||ȕB"OT�"�ч�$z	Ɯz�)c�"O�T�G.�k'd`Sw�;<�v�t"O�Rrc+C=P��Wf�)��u"O�a�'j ������I�6��"O�أ��, ���)]ְ�a�"O0X�H�)�(0"�b��X�.�+1"O* �H�.0�%�Uo�"P֬��"O�,�S		 d��W�ϮX�"O���0$�7/`�}r���"� �a"O�]��C�$<�1��D f�2��T"O4�$f ;S���9��o͊�"O�Qu@�)W�$�̟\M��T"O6(��mE5Q�d@���_�7O��!c"Op�m�%K�(P��W(B�y�w"Op�ǁO:䒼�"�B�����"O����ȏ,v(1��O+/�nXk"O���d�V4V����wLJ�#�Lec�"O�`���%P�� IE���X�"O�5ۂH�.m&A�e��4+�8Yɦ"O]�&���u:�ad�V�z��Qv"OhIg΍�M�:a��]'f�D�D"Od��+�K���%��
K��2"O�� v�
+/Jؘ���٢g���0b"O�p�/A��MJ􉍢~��̱�"O��Rg��
�p�@E��#'�n�$"O���� ��Xh������+y�]��"O��#�D�'��S�PE�x�a��8XD;B���t�/�g~��ԗ�tqr���6G��v@W�yB[�&4�&c��ID2�9�. �wL�e��aCn:f���)�����^�*�@Ra�L{bͅ�	b�J 鰈\�9���ɣO��]R�E�d�zi���)K��C��/�(ؤ��G���",o�zc��ӄ".k�j� �#�'TޖHB��)��M��Q�S2���a¢�ys�Plpeh��A�`g��R�,ۚ3�q�'��@3��0�^�Z�<�7�*$�j2D���[�3��+0��YN:!��͹zr�x� ��;�����$Z9򜃗�/vȉCr�4:=az�Ȅ?���s��y��C7L� �K�^P i����y�&N`�p}	�jL�fr�-!��'�v%2%-#Ed��A��IK�N@�1%,�.����C��x!��˨[D��EI2޺ЊD��<�����D\��'zq�#|�'��9Qe��c�J�����y �i�'j���ŝrb�����Ml8s#�"�N�i�F�0>I�!I�}�4�E�8x��D�T��И"l�	됩�Ek��p�i˝hٮP��`H�M8]:�(D�����&�R�Ӂ��	�LXj�*��
�\x*e�˃.#~�Ă	>R���j��c���X�o_P�<A�b�74�� !0�U�/
����J�<iF ��V=� R��$!}�t#Ch[�<��NѨN�كa���5��h�L�<!�,�0?�`(��D!cT\y!��GR�<)#� <�j��D��Y�a��L�<�tE�>,�5�A��!�di�'ɌK�<� \=K�?l��ّ�X�����"O�aХ�N�Sp�%�I"p���Ƀ"O8aևI�[~��#��>���q�"O�]�g
^�����w��A�Q"O��{dj�:��P��>�j�C�"O�pf�-|!�,�3�_�����"O=�p�^8M�R��f	�	�|�R"O(ě���m^���V��4 �����"O�M�2�	q��Y�b'�"ai��� "Ozܚ���8�0��֏�!gNr"OdT�Ջ6ɞ�Z��!6(:|zW"O|8����"��;p4�U"O`5!��S%`�@Han�Ct��0"Ob�Z�GX���1G(z����{�!��%A�����#cK���n��%q!�Y$��X9Ff��:8�����\W!��ƞ:��1��ȝS(n��P'� ':!�ğ�#>2����ǜ#
���f��O)!�D�-0�fH�Dʅ�;Vnd��,!�_(���q���>eCr@	ep!�d�M��ˡkI��D����� ��<����'pB$��!O�P�2�b���8CF�
�FL��I�=ƪ��aًD'����Ҝn�z����&0��' ̪����z�)����w�ъ���^���J��I���p0!�I5x��q��2Vt�O��2�4�)�.�ꎾ R @T�])��'�=@!�)�'v��CQBʀ8��TQ�Q�7\T�!�C�T��'�D�G�,O\��go�7���BEQ�Ig�D�C�O��A�O�צ����M&�p<���ԤJ���a�M+�ʄq�(�y+^l�p��=Q��#?��&�B���qbB%<~,}�ʂ<�l�UN�.,$t�c�3�D�l�$u�g��`,,��C��m�ԟtȠ���?�@9�Y�!��y�D剥Ld��3��;�`y4�� fe ء Kc �-����#ȎbR�]��e3
�|O\��S��cH��S	il�)b	S,X y�̉6[D<����G��M��	$g��)��@�`�ɽ{骰ZS*-Č8��I^����u%�� EĘ�[�`֝5fw�EyR�]yh���A�&�2�5�B"����ƈ��pq(�(��\>�`J<�T�A96}�Ŭ
�\z�)�#Ư^Kv�:�����	����|�pݨ1l�s�#<��.!F)bAS@��d�!&�\�Ed�Ȱ)�c^�+��f��O$��Sd�+pL��i����V�6d@�D�I?��O�>��-υN�����W�:��,)p+G�T�X�u��?jq>T���iP�>E;bA��U�+6!J�eF�Q�'��0�%H�M�Bs��q��ϻS�MЗ@њE۬ԱF���Q{�!�y�4�Ko���10�w���S�v���ω1A��lq�G
U+ 4���'z��d�6Wop�R1��"٫&d�?c�@��'�3>�t8qNў,.�#`)�|tr���A��͉b�_9�RO���t�7Jz9l̘��jM�L@�O
����֬)�:���L�$Ty�#<�*�6.+�����][����-�|P>���!
Ypu�� 
��O����QTܨ��ڇ�:�"@Y�擛>��P(�	̒E�7Óc��p$��Df��RTjA�4��D���I1��DnV�s�-��_2y�L���Ѡ.dft;s�"A���)�S�yW%<����A�T���e����5�*B�}���	���a�X��;��99���d>yf�т��Оs���_w��D{���1�Ä@[;Q�e�M��t����'�z��/ڲjB������	F�9	���.y�x@*��#�z�\�)�p���r1�Ys�X�����*}=S)�f瘸r5-���1�R��1A�b�	��%����ZF�R�3�\��J?����6 ��`�bS5q����u�#�ts�MCҀ�2"&uS'h:���45��KSi%k⎐�R�5N�PM W��TUP� �oe�PD��O�Ă`&N�"(�a�2N��VІ}���OZ4�ʔuJ<�¶��%�0|!L����1V�k$&q !Ц�Y�#ɅX���f��� ���I,R��x���SQ�!r��^1��b�(�������K�¨�ם~r��3Wx�R��C2E�I �h�\z��Gn\!� 4��ǋd��p�cEBæ(y�M�3
��5pw�ÜZ��Db��C����^����*Ҹp���� 7d�d���2qhNt���S	c��E4������Rg��*���(�NŊ&�^+2	UV]� �D���R+ԭkt��Q?�V�>����m�fś�������#��w�<Q��/+��X�㜘�>�xd�ͦ���m�{���5��U��y���T��&M��3U� ��=1��	!8&j��D�g($@;@��KT�R2C���Ԙ�F24�� ��Z������W��8Hz�Ѓ��_�X��@c� �Q>=I��Ҹ$����*"��J�+0D��� , �U��ev1��a ��>���'�Ȑ�q�D�i@Ο��|���.o���x �'P
8l����@��,���,{�0�P���B��"ѡD1*3t��w
RQ7��=E���s����W�9���1f��E���G}�`���nً�dD�zdQ¡Gcr�kea���~��9b�8��4V�x8��IMƖ1PK�u@��	�j@:Hr6�)�)r�K	�qH�牪s�q����.Che� �ə\�.B�I	U��@sgπ`� ��F�/>��'� a�aA�Wl�k!j�X�S��mC�\s����ګZs"l�$�3�p?�aLK�	�b�X�R0i�:C�Մ-G��Zc���a8<%��0�)���ґL�>?S��:tj�,S��5!���ͳ�%�n��VV͑�I2'J�zA̀5K��'����əSN8�kF�Id}8D���I5X;�mbC�"�)ڧ~:�8�߷,n��˘%u̸Y�ȓ
�\zu�G��P�C�"W'�ႇ	@>���	�E�Z���G�hND�+a��
�'^�������"�R���+�,q�� ;�'fv�b�$]�h����e�y���dF"X) 
R���'�lQ!ІCZ,r�*�1!���}KS� � �4 (`Cb$9�'��%�0ɧ=ɧh�<��%�*����W�U�l��"OƩ�l3�И:���Vu��>q�]9 3���
�Ƕ)�G�Zj�F��0���y�@���2T�L<�&ܑ=b���L��^�Jĩ��L��=��)k0Hɵ�߈xЮ�	��L�M-�mG}2��X��ȇ�	T�Sឱ���ɫi,��mH5V�!�$��2��W�XF��cs	)Y�^���r�x�rrG���S�O���� P)p�z�C�k	K�f��'�&�@s�O;F�F)���.G����L<���r)),O��Sv��(*(��	 �$4���U"O@�ʃ��S2���(�ho�t�f"Oș���ۋ"dVPr��� ~�P�"O�Q)4�[�p�A���Z�$5�"O,0�)"<q|�*r�� 9�D"OV�� _��P��BEy"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��   �  C  �  �  �*  v6  (B  �M  mY  3e  q  T|  :�  �  �  �  L�  ��  ̳  G�  ��  ��  �  ��  +�  w�  ��  ��  ��  x�  �   [ � � ! V' q1 ?8 �> �F �L vS �Y �_ �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�'��7mL�2�p�)2N�&g]��*ϓ�Zφu����P�ݴ�����'�¯�'��SF�=�����df���'QVL{q�i��I�|�A�Ox�\L���5�C76���v�M�+���<	����7�'�l�� ԐOE�I�`AͶGn��aQ�i�0��y���ڦ�]!¶Ex�C,v�tX�کk��d�Iԟ@͓����ʏA��7�a��`��q�L�I�1�0��ǫy�͓o��z�����'Z>��$�R�1�&�8�o0Q'&���'��I��#�MӲ��Q�
wp�� �.2�l�3�\���ܫ��o�>���?��'��	 ���r!�G�{!��h�Č3���?i�ND�f0$�|j�n�O2$�,��H�
H�48c�+D�`�*O"˓�?E��'0��sΘq��a�L^�ke�Tk�'�7�M��	0�Mێ�O���$ƪa-čp��N�5,z���'���'��øST�F����'_%�T��VT��se��<3� ���K0��-%������'���'�2�'���s��y<�qw�C�]��M�!X��޴W� ����?�����'�?!��?)#�l�e��_�P8!�Z��	��M��i�O1���i!SiT%S�X�I��H�D錍n^ZDb�0O��д���V���@�d�%XM����W�0���/L���qk�6�.������	�� �����}yk�ޕke��O����ݪ1��S���s�B�qR�O,�n~�s��I��M��i�h7�Q��n1YP!-�"��ӇQHi��_�7�*?IT`A�J�X�) ���`�=�]#9ebԛ̊5��R��I]uT�	���	����	���D��q��`�#*�Fcj�9�
4��� ��?1��LśF�$��I�M�L>���<R��x�`[�aB����jY�'��6-N�� Uú�mZ{~�MK�y�8�CP(�n7�aq3�E����c����`�fS��+ߴ��4�����Ox���;D	��
�2�h$�����d�O:�l3��%Њ���'^>Y��M߹e��Ͱd,�;}=�@�??6Y�H�	�CN>�O�� hT�K�`���\7����rNϤF���*������޺k���O�k)O�չA�����!X��]ۥ� LFn�D�OD�d�O���)�<�4�i��y1�D�d�D]�3�_��~��r� ��'�7;�	���s�8��&��9o!�})2��"��|B�C���"ߴ_a����4��$�"!�q�'��S�z��`�U(�1>�j���� `��$�ߴ����O>�D�O���O���|2	ˏ��L���ًs݌�@��
?כv�CI�����,%?��	�M�;e�r��J��dtx����$4ȁP6�'��F@2����FS9�4O�uC&�ՀL�=��E�%�:u(�0O\	`���?	2��<Q5�i��i>��I�17$Y��据c�Ȋ욐6u��Iß��I�8�'1�6�K,ZT�$�O����T� !+�\�u�����ۭ@7�㟰��O�5o(�M#��x�M��\4��B�g��H��.N����'|�t��HM�H�S�O�譻KiT���2�?�Aǂ~�(�(��!p�����CR��?���?i��?y��)�Op�:��D9I����$�#0����o�O:�nZ5������ �ݴ���y*E'6 \��C���6,�Sa��y�eӈn���M�����Mc�OvT������7{R��0tj�Z!�m)R@ª]�˓w�F_������	��|�	��D�15�P�`uC�~JĤ@��iy}Ӧ��0F�OD���OH����^*"��I��
<�P R��S#y���'��7�]rL<�|c� .o��Y�!JT�}��҂Ȃ�WҎ���}~�%Q#K����7{?���M�-O��CE�?[b��6�,�,ȪAd�O���O����O�<QF�i�H(��';�P�dMU1:�Ra�N��J��'6^7�!��1��Ėަ!X�4K�V!�+zuDQa-��(Cդʉ�rAxW�iJ�d�`��TY��Ɖ^��t@�:��ba�� ,uJ�dT >���s�H����?OD���O����OT�D�O��?1�w�� `��ش���qI
0�m��?q�i�N�	��' ��'#�'б��%V7G%=j�EX=m��)��A}Ӿ�N���a��i�7l��6�=?��N��]N��87#Ƨb3�d�G,U�Q�
a����OP|".O\ynfy�O�2�'�� �<'{❑�n��&��uKaτBqB�'��2�M����?���?��'�� �Ƞ)�R�ؔfH�s��<�a��<�������O�7�K�A�´�%
x��ӏ��E�@��DB�N��TZP���*��'�T�]
+�\��;y���yW�� 7�\l����8:��@l=c�"�';��'�C�����aF�I��ugjêkZKT�WN^����ZQ�R���':��
~��_�擅�M3������V�F��em����W�<�6-]��B�˦m�'�B��EB�?����(���  0P��[����i2�/���'���'L��'���'���?k`���e�t��k�>���4&��(@���?A�����'�?9��?�;��5�5 d�[$�F���Yc��iq�7��Ȧ)���O��`�p�i��䙯`� (�P�ʿeF0�q��O�P�������k��k_�ʓʛVW���������p�R&��,yʔb�e[ןd�I�����oyR�h�R��C�<i�w�Z��o��F��W��?m2�3������O��'a�7���޴����.;���х�֗}�Q�mI���I�/��{5,��r&.�\^���b�>��%�?q�h��*=�h[C��R,h\���H �?A���?����0X%6��̴e������O���HR(3S��¾{亱��L�O^�o�5F�版)(f�S�X�'ݤ��O�;��� w�\+��|��1o�╸0�'w�7M�ߦ�Sڴ"��(�4��Ğ�h�����h="�1x0dB��� ��{ ��O���W�e�����'�"�'@��'V�	{D�Y�X^B���`܆!H,ը�V��)�4G���R�F��?����rƁ/�?y��y0��'Œ_A�i��f &H��QS�� ڴmj��	b�|�D����7����ώ!��q���(Mcw�����01t]���C��Ӓ޴���F<@�f����dRH�p��@��$�O����O��4��V�&&�)q4���:J�Ua&�M*�z��θ�y��~�X�h�/Op�dnӈ<mz�d��"�R��T"K8VV�ɠ0�3 ~�LoZr~r�B�ZԀ��u��Gź���*��5 ���#K�"T����1��ϓ�?i��?���?�����O~ ��� ܔ
ͱ%@5 *�\���'
R�'h�6��:�����֖|2cʌdp2p�Ҡ�-_X� ���PW1�O�m��M�'zh�	��4�yr��W5��@f����\�ヂ"[D�mk�-�N����Q�?>a�H���?1��?i��@�BƎŀu�&q�2Nн[7��a��?q.O�m7�B�	�l�Im����}>bԚ��,t�&��$�~y��'��V&�T>�b�Mh�xY;D�������+� .B�|Y��C����|��(�Ou�K>ɢaC~_|�ٲ-Ш �$���3�?���?���?�|�)O�xm�(���46
2 ���`t�PA�0?�3�i��O�'�V6��\"�L�7�+
m	(G@9n��M����M��O�HQ%"Q+�rK|J�&^k+2�Q@J�>[�L[�ay���'p�'^r�'2�'��S�c������Mp����*	9�^U�4�@=Γ�?i����<�v��y�h��mc����T�L@t��G��ϲ6m���0M<�|:�@K��M��'��P�U�)�b��f߲���'VZ�����q�|R[���Ο�CD��.brt�cdI6D���UNN�D�	ϟ���fy�
p������O>���O��##I��/�ΡT�%�lmQ2,����D�O���(��*`3�pQ� �����K�+��N����衒ԭ!q�r�&?ɢ��'�r��I�;�Rm� ��)7�ą�E��%�@I�I�0�������f�O�R/��lƼ��c��j�j�K֣�B�R�d� 5�G��Ox�� ɦA�?�;E��0��^@�ʄA����f��sț�OT7-CN[�6�*?q����J�)N���ǪT�F��Ņ65�>��M>�-Ol���O*�D�O����O��:�M�0I�M�C˅���h3è<�v�iZ�F�'E��'���y���Ra�Q�+JfT��Z�Z�
���f��O�O1���rU,ž5�$��G��1�h@jT)������H�<��O�Iu8�dͣ������7�<�0ag���Q1WG�=�\���O��D�Ov�4�n�c�v#�B�bE޻ N@)W@�9�y$lB58W�Md�⟬8)O����O�7��;L��h����60:�#)A�,��p��
aӺ�AR˖����:L~��d�E�v�K�K �<B�"�!j�ziϓ�?����?���?����OǢT�g�T���a�)�v��7�'{��')7�-��)�McI>�aN�7��k�?M���C!�'��6-RΟ�I�3¶6�9?�aN�7l
�U@��$*G�D�BԎrM��� �OhL�H>1.O8�D�O����O�!0'��~v����^+X@�Eg�O
�D�<�@�i���'���'/�������F�<���ě:g�R	���Mc��'U�����O��͚i�ZA��B��4	�2�kǋݐ9���A7b�.��?���'�Pp%���cHt���B�/'�������ʟ�����@��ڟb>U�'Zn6m8OS�xj�e�77C8�(!�5_�D�%e�<��i��O��'��6��x�2�KF��5|���JQ�&Ql�D�e�Mצ9��?���[�
�N���k~
� j<� #4��`BE&���;Oʓ�?	��?)��?1����iN�:������-�x�#�7kўTo�y�:u�'���)����݌� �
/H�JCk�f���4 ��6�'�)�"��m��<q��S#ED�hP��{`X��D�<yD����$������4�D��pĴ���G
�Y���-;~����O��$�O��	��f�ߌ	���'A�
+�Mq@�.qÀ$�cV�8��O���'�7��ͦ1�	ry"��Re�j�ŝ`v2H�iA����;��%"G��<n1��)��0nF��H����1�-!�ʭ�Γz��$�O��D�O��d/ڧ�?م��+f�D��P�I!}V֐���?��i���!�_�,��4���yW�ڃQJ4��e�=B��
�{v�<�5��Nc��dʗ"��7m8?�IH�ju����(7:1��
%;��=���)&&�axK>�.O�I�O����O����OR�钮�T+��(\�&����7��<�u�i������'R�'���y�ړ?Μsd�Fj�ZTId��9Q��c7��e����t�Ob̜����)#�:pYâ�`��-��$�6|8\�2�O<��`�4�?9e�3�D�<��kJ�&����Յm56�
�0�?A���?q���?�'��D^ܦ=��`x�\�Peĩ^�`�N�!������w�x�ݴ��'�z�U@�6MgӸHl���\4Lƌ]u� @�
��l2��*P����I�'����6���?1�}��;՘����޶Q'�� �U�#���?���?���?A����OQd1"��!Pk��b���bc,u�'�"�'v47m;h���&�M�K>�U��=Fc�Ỡ�[�!F���Ǐ.[ĉ'È6�Zަ�.	B�mZc~���{���b�N�"^�u�� �{zz�Y�Ȟ��)�|�X��Ɵ���矠`�:I�&u+�/L�g��y�$^˟��	fy"f�O��+�O�$�|�73: ]0�Δ�P�u3��@~bɽ>1��i��6��N�)P�F�\s�5��LA;j�d���O�9U������K�
4��ĥğ(hT�|2���4<��r`�7<ɴ%�q%l���'2��'���_���ߴ�(�����2��p���W�Q�؍�q�N������?��[��ߴ-���q0��U%���뛁�L؆�'Q��*L7ћf��(���, ��@Vy�f��\��cA��.4�ByYW"�,�y�Z����ğd���\����X�O�H���˛��I��u�	0�l��cSc�O`��O����d���]3����P1y�2��a��YR�شot�x���]�E��4O��1NR.p����������̎$-��R.4��Ɂ�y�\�O�˓�?i��e 4�X`Z:X.�zv�"�����?1��?�+Ol�?�N���ݟ��I�(�����L��"��Kڣ2r��?�V�(�۴+�x"�˚a��qȃQ�Fƺ�)V��2����,���EbT������e��$߈JE:�XӃ�tVddIBJU�E�����O��$�O<�D9�'�?a���U�LL�߈"�Y*�-^<?�rIxӄQ�A��O������Y�?�; �&���	�� �@l]�8�q�Qy���O�7m���\6�<?�`lL14�����'������sy� ���2�<�3H>(O�D�O��$�O����O����2,L�lp�`�"��0)f��<9�isX����'0b�'p�O2¤�60l��CI�!(�-nL��Q��[ڴb��x����P9/� 1L�bT�)g�ڲa4`���G�"k�kC����'��$���'����݅v�`��
өoj:�8g�'%��'����dV�����څŜ���ѵˊ bY�L˰&H<X�IC`gy��޴��'	��h�&O�Op7U�s�P�:�'؝Q�A��զb����k�:�U�����	���IL~Z��Z~��bԫN�i���bY=[�v͓�?��?1���?�����OSz��D��F�l F���j���b�'B��'��6하u-����MCL>�6@ô����_�܈��4�[	o�'g�7-_Ȧ�SQ�flZ~~2m@�i�`�����W�茠�Ð>Ѣl�0H�ן ze�|rX��SПp���ɴ�Ĉ(՚��a.])X�:�I�ß<�	Ky�kd��\�gb�O^���O�'z²�c6 �&\�ȑ+�cZt ��'Hf�$w�F+�O O�	���]{�'�Jd8MB�kݻ#�\��ݵzdy"@��$~�F��B�I�O�qSO>	3(Ŝh!��pQ��l��#��X&�?����?���?�|�)O�o�g �b'� �oh���A]�V�,�A0" �t��6�Mӊ�b�<iشs�%cg��4�"�"�K��{��&�i��6���1�n7�k�����:�0ݱu�O�|��'u(��G��	a_��� ��.5~U��'�I��d��Ο��Iğ���^��@C�<����	P��h��$x6�6�K�!�8��O&�!�I�O�mmzޱzR�Ý<�8:�g:,� ������M���'$�����O��ě�C�F9O̐K�΃��%�t�>������y�AN�BI�I�'
�	ğ4��_�U�Ae�4NʴQc����k�����ߟ������'B�6m�$G����Op�$��e�2�q'�*Jƴ�u�r\��౫O�lZ�?�I<q��>X�lZ@DK�jD(=��jU�<9��DT��bJ��T�~51.Oz�I(�?Y���ODu8�`�
(U�����Ⱦ�P��O��O|���O�}
��`T�B�]�ݲ�L�'��U��;i��g�#[���'�7�/�iލ� �_4m��t"�d�&>eD @,��xo�5�Ms��it)
S�i���O8������"�� �,A���[(M��G޵kzђ�!$�ľ<���?����?����?Q��L����Ѝ؝$���JF���E�%(`��䟀���|$?������y⭎�X��h�.Z }���O��n�&�?�O<ͧ���'Rಀ�qGƉJ��a	ܕl&�V�C>'wL�.O�W���?�q�2�d�<aqű(�B��.e�TڴO:�?Y���?����?�'���AȦm��'ʟ��󭞨]�B	���ΘI?5K��{�d��4��'�v�q���D�O�6B(�z�� �d�!c�����p�Ǫx���� ��/��S:�*xyb�O�h�Z���⠏�{'�hï
�y�'��'�b�'�R�ɘ/W�<�9�lQ�B9�%H'e�����O �Ć��5��t>}���M�I>i�E��s���i�L���P���'��7m�˦y�S�x�>�l��<�������'��G;x����X?&,[�E]�RwN�Ś����D�O��Oj�D��!�*���{0̜ёJL�p�"���Op�/���d�z���'mV>�*d*�m���R���+K�@��!*:?�P� �ٴ)��&;�?�	�/34�Fԑ��_w-` e"�`��$���|2���O\�+H>s��*"s���g��U� ��N���?���?���?�|")O�l
�����ΠD����̱oqj�pt��Yyr�xӚ���O�0nڹIu-#!犱7��QGb
��2��ܴa&�v7C�6��3���76��~�Ф)p֐��b5]� �7�T�<�(Ov�d�OJ�$�O���O��'.�ָ�0힎o�H��1(��(��S�i������';��'U�O9*`��n��e҈0�cH�(,��r�	̱q�&-n��M�x��T6G��<O��{��o%�1kB
]����<O��"Rb�3�?�Q�(��<ͧ�?��	�	�`:c�_�}_��g�+�?9��?q���dG��ix
Q{y�'��)�;Z2)�� �8��-�d�t}��~Ӵmn���@�I0���U<�[ծ�%#�u�'&�ha�17FL��� ؟d��'	m��J�j�nL�6Bɓ<�$]�c�'�b�'u"�'_�>1�I�^���J�O*wdA�D�']�(�I��M�Cb�,�?�������4�t�y���u�Td�%!F(��8O�l���?��4!!�"ڴ����YFb����Cu�	4|���T-�)82Hq�&7���<���?���?q���?�sV]`	��K��0��7O����ަe��-�����I�%?�1aN�R3-D��j=��ƌ0N'6�8�O�=lڻ�?�L<ͧ���'<n�e�#�]&F�3EM&#��m������#.O�dj�E�?a��1�Ľ<���̾a[����'Oq��Cc ��?����?����?ͧ��D\ͦ�[@/�ޟX[��4����-Q<A��.����ߴ��'��˓�?���M�4[z-H��4e����
�Y0ܴ�y��'������?qZZ�����ߥ���ɺG��Df����R��}��������	���	������JQh��H�7u��}��D߷�?���?�־i����O��LqӬ�O00)@F/;��[�k�� 5&��S�ɘ�M���i.���C� ƛ�=O����zd��rR$qa�hb�źa|̚g�X+�?�6�D�<����?A��?����j;|E�⯋�@�dP�ҰB�����4�'d�6]d]����O��|�`��. :�����/8���g��v~�J�>� �i�d �?E��!��>��x�*ހG2�+����jSO�"-����i�����$�|���;.�E�9G�R�'$VB�'���'e���Y�� ݴ ��#�@(NɎ1"���wG}��KĠ�?���O/�V��J}Riw��1�(X	C�e��h]	U�����Ɛ�%;�4?�$�B�4���ى�i��'��S�E��{�$��V� �����9Ќ��qy��'���'�r�'��\>��E΋W9JX��/�5Oٴ���ψ��M���	�?���?yI~��r������L�9ToN�Y.���eaC�B�i�"����jL�Q�g���	�'*)Ed͕���G�׊2�D��#PR����'-z�$�Е��4�'VfPr:z�<±	�T���`W�'��'��]�� ߴ/��̓�?��\�b�� `�0T�`Y�+݌{fZŋ�r`�>�&�ih�7�n�ɯ|����7h�m���q���⟄q�cڛ[B�'+7?1�� � ��W.�?����=� `�MX�r	�ț�G��?����?9���?��i�O��y����r��8�VB�G�"�~Ӽ�0"�ON�D�ڦ��?ͻzz`!�c�6mQ@Ff�4&�$8���?q�4`f��,՛gs����3lZ�t��Ɏ���:w�ʅr��x*�	#���$�t�����'4��'���'L���R��6+y���Kn�@�V�\h�4>�6\����?�����<��Z�1@ 웡pHP��a)U5/��|�'7�릅�N<�|Z�
��/��a҂ex2N��U��0�����~~��={
m��;|[�'x�ɜ(t��7�Dd�H�AMN(ޔP�	ܟ����i>U�'��6-N�AK��d�.Ep�Y��V���L�%[I��dXަ��?��W��;�4����iӨ]+-�=�\h۠�%���z�أ1��6-r���	�]t5�&�O2�����;[�8����k��A�B!0,�a̓�?����?Y���?����O:�YE鎷8�6�H�̩:*ʄ{�OP�$�ȟp`吟D�ش�����w����|c���Tw����x�Nc�P�mz>qIF����'@a�� ��&��5��ubem�+v.��4�K�?	`J9�d�<ͧ�?Y���?!D�Z0c"�9`eU�m~^�r��L.�?a����DҦq�	����	��$�O=���u�� �2L25EŚX��Op�'E�6��֟�&��'V`Шr� �(�DK5���t�R�*Q�eÅ�C���4�pQ����P�O�9���.t(d�	T�N��I���O���O*��O1��pJ�6�ɓ8�*��,X�p�az�I�$m[�,�3�'���q�4�8R�Ov m��dyd�yd��Q��<*�!A��	P��MC���	�MK�O�02R���z���<�1��43H]��FLj����U�<a+Or���OD���ON�d�Oʧ\5bzF#C������X�&�*�i�t4�!�'���'��O�r���X5�Ƹkrs�ոs�˳!��ilڐ�?AJ<�|�G!U(�M��'Z���7�����жO�$��'��PySJ�<�4�|Z�H��ΟT��G�iX��P�ظaKݩ�ӟd�	ȟ(��ZyR�r�`� D��O����O��z�L˕�$��ێ_L:D*>��=��D�Ԧ�
��ēV�����LN�:%j�b��=at �'sJYe!	1�¸ U�����ן� ��'�
lgd�.U����4oVU��a0�'[B�'��'��>��,Y�Q��ҹ,�h�c�
x���ɚ�M�AE�!�?	��!����4�ċ�+�8_ڂ<��T6�½!�6OҀoZ �?q۴���޴��D�N������"��}K�m���*���'�*��Q%3���<���?Q���?!���?��E$T�``�IgObtsd�'���9
R��by2�'��O��@�wIp�
�(� �Б#ݦR�N�l����O�O1���x�I����TA��a#��aL037�u����<1s,҆<���d:�䓾��F2W$f@�D��Z��
�k�]0����O�D�O�4����֯��2r���e�Ƃ$2��y��=��Aq��⟤{�OV�oڳ�?1޴��t�g,E�`X\�î� �� A�����M�OT$����,1�i���I�/}C<����>���O����O��$�O���5�N�Ta�/�R�rC��+�P���՟��	"�M%�R�|��&��|�`R���)s�X)Ju;��À �O@�d�O��$ų���$�ԉ���Ĺ��P'edr�����\@PQ�'Q'�P�'���'�"�'�!��h:���կ\�@�Vi�W�'V�P�(zߴ�����?�����I6B0�`#�W-
<u����:Q��������	�����S��kB
G�❹��  ��a�আ�5�&ds�g�ϐY �_�擘n" �m�I**DV�zA.m�w�	T�Z�Y%�����՟���՟b>]�'� 6�S2���Q��JK(�f)��_V��7C�<���i��O (�'��6�Y
~��!=9���X8ک�I�y��H��a�'9�1�pK�?���X��h�)�,��Y��U�2�8	�a�Ė'�R�'��'~��'f�&Z��r���Z�L��A
�q���4�ڱ	���?����䧷?!b��y�a�~X��@��_�RK��"U�I�6=�6�Ӧ�O<�|������Mk�'D���ݐNQN���J[/G@DQ�'
�a봄�ٟ�rđ|�T�����wmR�G!d�k N��Fr60�'H�˟������iy�ay��P��*�OH���O؅3b&	�C�^,��(M�`9�����<�����d�O6-�c≎L[�lx����f'����#�5D��A�xYf��"!�H�|�VB�O�H���B3��Y��7``� $!J�v'8�A���?���?���h���;3�"�"��ρ�
�"��7��d���]�$���������Mk��w��X@*�� ��)��7x�@!�'d�6m@ĦQ��4xʔ��ڴ��$Ҷ\o�\��'Nj z!نF�L	[� �`�s'�&�d�<�'�?	���?����?���� V�|�#�Zi�UqT-�4���	C��J�����%?�	���`d�!gK�T���	i�:� �O�0oZ=�Ms�x�O/���O|\�b��8��:Scf��1�H�8Ȁ�O�� �G��?��#�D�<i�ɇ�t��y8`�_�2z�M��I� �?1���?���?�'���Ϧ��oP�lZ�*X7^_:���*O+ ��I�'o�柘��4��'�x�vC�&-�O�6m��{؞y�SEB�"�"�Q�J�p�3�j�j�E�ʰ+�"���T�J~���0!T�+%�0e���h���2pҋu���	��`��������|�: ۴M��ds���G�,��cC��?����?���izf|�͟��m���'��	:�̓,��1/�8p�o��Ot`l��M���=�1yٴ�y�'���9!�ҭo�
�ÓuO"Y��h�78&��ɤ0��'<��T������	=I�$��_�VF�3�b�>���韴�'W 7�'Z�F��?+�����Ɏ������A��1Uċ6��$b}R�k���IE�i>�S/&������΂9 P����9b��O y�VD�CcGy��O���	�1U�':�]�6�R;<F�5��ò t�R4�'7��'B���OG剁�M����9�U�\�K��9�r�&#�-���?a�iQ�O8i�'D@6m��d��/7'��&!؉>�l!�MCM�M��'[BБ�p��S2	���5"L��Ѓ�
�1*@{�j�IRL�My�'B�'/��'�2U>Q�g�a)��ퟱ2 �%��Mcլ�?��?�J~Γ���wA�i���A+���$f�)Pch	��"��Iy�i>���?�y�o����S�? ���1�?7��JU�A�Dj�>O���wϭ�?�4i=�$�<Q��?��K��$�*�6�Y�������?���?������������ǟ��I��!ӬU�|۰lB�MEJ����o�$��ɔ�M���in�T������%���k��E4�еp�|�ɖ�d�p`(]2���j�;m�d8�?��OI���`?N&�#sJ�?���?Y���?Q��I�OHaG͢�ļ���X�9� �O�<o��
r��<�f�4�bpiÂA-7�,�10�Ԉ�2؃R1O��nڻ�M�$�i5,x�iL���OR�s��=�â�,/�Y���X��2P���v$��O���|*���?����?	�9=�0S"j�8��A"-F8�B+O��o�T,���ڟ�I\�s��R#�o���Z+Q,[�Ր���Oj7�o���)�� �j���0���:���|`�ه˘)��hr㘟��*W�S���zy��-�xZ�ɟH��4��I+V�r�'	B�'��O$�	��M���Y��?�F�F��E"�Iz�<D�+@&�?�3�i'�O��'��7M��XmZ����T6xB4�S�H+����צ��'�`��I��?i��w)t��V��+b�8���%���{�'�r�'��'��'񟰨ð�5VfDu�5`T.K'��O �$�O8�lr����H�޴��Nx���T��y�R��܇���गx2Hh��8��&m86gj�
�Lx��`�f���Tؒk�)ӛ�nZ0\�ն�M;RA"���<���?Q���?��l�M�ҵq�T?hv��{�k��?9���d���IZ��hy��'+��^E����n"k���'��tA�	��M���'u���	�e���	˖t�, S6��4����H��(9ͫ<�'t�h����w��آ.	4�4C/SCDD���?���?9�S�'��DZ馁�6G��eoJ=Ц*�5a<b�2@�
�$.6$�',�77�	7���Ҧ͢�aS�Z�Z<�F�G�k`����Δ�M�v�iD�\H`�i��	�[ZX�6�O�L}<y�U.A$�10���&;itd͓����O��$�Oz�D�Ov�Ī|2c-
��D���ӄ:&tH2l�-��6Ͽ2�'B���'��7=��H�ʈ��Ą0%�*�$sW��Ħ��45#���OD�%�¿i%�d\�}0^�HA,@X=sQiU�Z�D	Y$��:��T�O���|��)9�e��F�}�pyچ���h���?!��?�(O>qm��>��ğ�I0D��Y G��+fVmS�I6�
(�?��V��H�43U�69�D�  $I('��
g���R\�y:��O8��҉L�jЊT˧��d�m�2O����ZrH���~�J���6S:!�7�H�4�����ܟPF�D�'���j� ��#�&��Bρ1K�xA�'>�6M��n^��:B�6�4���h�� ,"B���%�<�8M�p4ON�nZ �Ms�_X�(�޴��d�7�|A��'z��C�ֻoE����$5E����#)���<�'�?!��?Q��?�s)�l�9��m�h�Zg�!��@���b����8�����$?=�	� ڈ�$m�/cn����[8!��OhlmZ:�?�M<�|ʓ��'0�,����l������O}0J#�:��/G���6뾓O ˓�X�B�,ݨo/�]�P��+� Z(O����OP�4�zʓ�F���@R�@�p�91���c��4�y��yӨ��C�O��o��?9�4=��`h�d�@ވIJ����a�sb����M��O�iS0l̰��t9�	���@�˜9)�!���ۂ<���&<O����O���O���<�|�!�maS�[ .�F�Q�/I"?<�����?���:��fdÁ_8�	+�M�K>�r+����u��̥�%)��'vJ7�����E=�6�&?�r+7'�tH���n�,�!.^>d�<p!�O&�L>	)O(�$�O��$�OX�F��g���IJ�� *�k�OX���<B�i����'���'}�7_�`��$d���@��c �8)�n����M���'������>�����d����U�D�`�@�<C8�t��Ny�O���	�s�'��Mq���p,�b�5� و��'���' ����O6�ɢ�M�cA��dVL1������b�#0P<j��?1Ǻi��O,��'�d6M�",�)�dA�7R�)��.�7 �	Ҧ��P��Ȧ9�'��@�0N��?�sU�h�B��|����@�.戤Z����'?��'�2�'"��'���,�f�*�LS ]A@9"��=8=��4q�$m���?�����?���y7 �	j�X̊F�LK,�;TMZ�1c�7m�˦�!K<�|���V��M�'ݴ9�!�^D�(�S�Y�<�Xhz�'��)B,A�ɳ�|2\��S���!�N�O�i����i��|�ՃL۟�����	ayb�l�~�"��O���O~UӤ^�N�fH1��v\ �f7�	�����ߦM��4Lt�'1�%����9����M	����O(�5m�#��g�)W��?�g�OL����AH� &�߮Dp�e��O$���O����Ov�}��&�0��5�^�(�pN״f���1��Bg�֪D2m�I/�M3��w��9�O��c� <p�f�Z�<�2�':7�@Ħ���42\��4��DL��(u`�'B��4��0��A�7q� ��JKDO���|���?���?��7���2�2\"���ʁ?�b��+O�m�:���ܟx�	o�s��)�	B�t��BJ�b��}�W�%��D�צ"޴K����O}v��� �y�k	�i7�7��
�t�
���|��ɘ����e�'�)%���'��wd�*�j����5�,�Ȅ�'{��'�����V��4D�`��qx��q�7�X,�C��<*@���e��V�D�i}ҭv��m��Mo�Ա�����F.;�}���vt�)ܴ���@�xN��ĺ3����w
��z�d��yHasd�˿v "�B�'M2�'���'b�'_���*\=��D=���QF�5V 2�'gbv��E��:�������9&��Ȱ� w�h�h��X7B��<x����ē>���j�O�	(=��v���Ȱ� �@�EZ#�E�H����$[�a<��:��'&X�&��'��'=b�'�������:l�-i���i&��j��'�RW�hXݴ{pN� ��?������٦~.Ri�S��1(�8��Ѧ��	����榹�����S�.��>�rQ���<��rgB�B����B�En ��pU��S�3"�G���y04���|���B��D��������I���)�by�Bh�$�:�A��Zt����ȸ�DP��ʓi����d�l}"&w���"�$O{
��6I�M��"����ܴ4��ߴ�yB�'�"�ٳ	F�?�h�R���J�e�޽��U��@�r�|�T�'���'���'wr�'��ӣ|r��6*�.LF�0�'����ݴF�΁���?!���䧂?����y'�K#<2*ţ�]�^4�@��7L��6MJ䟼'���?Y�s}\�P�i��$	��x�$F�W@��Z�D�%����IV����8ҒO^��?)�*]�`�vH�R�ur�G@	iK�j���?���?A.O�o�s�8��I���k�|����4�Ƞ��I�$� �?�T�P��4j�xRl^^�ʜi��&=�J��i���y��'_ �уe�*�X��X�d�ӑN���?�R�-���)a�<�pyJ!�ɘ!n2�'���'Z��'bT9�׷C�"�'PAͺҘݑ��R28�6�RP����qӶ��7OZ���O��D�<�&�	�8�(x#��&!wPd���,Rc�x����?a�i�x6m�O�pT#~���Wc�|�4
���lS��!����cA,Rؙ�Hˀ����4��d�O����OB��I.ddLe��@]+�ttC�bK�5/O��o��}*Z|��ޟ��Ix�ޟ4�2f��%�����[��O�0����?����S�ϪPhu�Au7�����>��܃҉ʨVh��'�`L�î�䟜iÐ|�^�D��dʧkp�bJA̴1`*�ğ��Iݟ���֟�Svy��n�� ��O�]A�D�I�֜0��P�di�B�O�!n�X����#�MӢ�'U���Q_�lT{���E$
Y$Н"����iO��1@���Cd�O�^�&?����Lo��$�\���GиE$F��۟��̟��IΟ��	]�'(�%��C�{�D�7�^{aPX����?��n��鈒��$�'X7�;��"ɂqBD&W�P`ï�/��)&� ;ش��'s�*q�ܴ��d"B�⌙�n�'K!�pb��Ѯt�J��H��?�'��<����?����?Q���P"i�7+�3lPh�9��9�?���d릹�g����(������O�|�&J9 L��,��)[�T��O���'��6G�� '��'�x��FeW�E�5��
�'/���Q�
a���T$[���4����k���O�L�u�Ŗ54�P9R��(d�@D��O4���O��O1�`˓9כG<V��0������֎A� �>L�qQ���4��'��
���b������4�X���G(�Dn�p�C�h���zrXhB�g���L8,OP�p��οM���ôE����K�;O�ʓ�?Y���?y���?i���	��z�M�b,�M�W�*N�R�"ֵicN]�'�R�'���yt��J%ee����kؤXO���ɓ��XnZ�MC&�x���@�@��?O�B�,]�3�N���A�|��b63O�U�1�	�?��8�D�<ͧ�?qBm�K��;􋟄�ށ!����?A��?	���զy2kb����ܟ�J�h^�$8��S�g�$<?�prC�h��yK�I<�M���i��O�us�!H�(�ry"�G�<�"�>O��đ�c \@�kD�E��I�?�� �'���	�#���n<	�Œ)����G��O~�$�O��D�O�}��?����v�O_���A�o�%z�`ݩ��qÛ�O��7�b�'�
7�<�i��b��)��}qP���w �B�(k�Rٴ�V�}ӆ=�`�
��ߟ�j��P���Ģ��_��(xWO1���`=*��%������'f2�'���'	I$&���x����|b#Q��Rڴ"�������?I���䧋?�G�>��5�ДLp�(a
]�	��M�B�'������O��O���1s֏M��1��"V�>�tX@6W��	�X��г�'�\�'���'��U��ƮEAb��_�wD�A�'���'����DZ���ݴ�$a��}Cj�iC���N�4q�g��R�����Kћ���u}Mr�
]�	Ц9Zf@�&%���(�@J3�F!h�h�5A�hmZd~⠕�y��A�ӫxq�O�������Q�aȊ��y�OV��y��':��'���'��)"[�8b`,�Y�BࣴlZ�Z�*���O������}>=�I��M�H>!��/k�/ѺL�h���@,2҉'Y�7-���)�	6��6m1?�*B�A!�\�N��SR�QxNHr���Oj �O>Q*O����O|���O�Y�íϒ>�8"�F�X��TZ���O���<1�i������'���'~�w�Xx@�e�0���L�`�g��	4�M���'̉��� B�y�"�h�N�ңNӳv�n鸓�ěO(���Q�(7����|JC��O�(�L>�����K"U(�=҃����?Y���?����?�|R,OTn�6}�20�Q�?N��Ď�Zmlɡ�����Mc�r�>� �i�8	xPm�ML�\Z�ʕ h�[�
�O�6�#Z6-$?���&)V�iH���9<8��S$�9�Ï��<Y���?	��?���?�)�"œ�S>SdI ���8=X�y�U��GJ쟀��ɟ@&?��	��M�;G xs��
?�,͛�H��{���r!�i�&6�Na�)�S)}���l��<����W'��hmp\P%�3�a����.�����b�Sy�O��(�� /��e�W YdJ�AK�����'n�'��	�Ms1�ج����O�с���t��0Pę?e )spB?�	�����ڦ�j����:������ԸM��d����6*ޡ�'�����|�T�C����Gڟ�CP�'D�hR�oG1ވ�
�j�s��3p�'���'���'W�>���P�3]	s8��B ʙ["}#C�'��7m+#T�j0�f�4��Ap�*`�(��c��u��:O��n���M��lì�Rڴ��Dh��y���'����ތA�`�f�Ƚ�6!V=��<�'�?����?y���?qQǔ3��(yH�}'80���T���d񦭰��������ȟ8&?�	=6��O����U�q������¦��4�?)��3�h*­�6�Pሄ���z��Y�F�"���!���A���O���M>I*O�D�M�^\
��@&q^�{k�O���OF���O�I�<�нi���U�'��p���@�4��k�4���'��6�"�	��D�O�.B(����t1d�&Ѕ:��X�$�T�8��iC�	�c+�����O�q��n͋�ȹDnVYI��"F�T*\��OX���Ov���O���>���(ᢱ�O5�dpQC�(b"x�����I�MS����ۦ�%����N�l�ꅛ�
V�Jm���ʟ�'�\7m��ӓ']|�lI~"b��:2��5+M $P����� C�b��`B2�|Q����I͟�B��	�W��	�V���U�c������`y�i�������O�D�O�˧"p���3��&vt:�q�m\ O�\�'��PM�VNn����C\�'BdS�D�$dx�P�~ؠ	D��#��D�TW~�O9@��	�.��'�ҥ!a�&b�p�R/_�t*⬙��Q���H�	۟b>Y�'�Z7MS�w��Q9���D<�t �U2M�DC�I�<Ʌ�i��O�t�'��7��>$fÌ�v@4S� 	���lğ�r�aI����'�T�A$��?M����7/6p^v�Z�-Lv�T$G6O ��?Y��?	��?	�����K*@��k��L�x!����%`�l�Ddt%�I��A�s�8����+ւ��;�u%m�5-��!�*L�2,�v~�^�d�<�|����M�'�R�R&P�B|���5��iƢب�'`�#���d�v�|�U�����DX��fp���!�5b��ş��	ҟ�Ivyb�k�@�Z���<1��c���6o]� �@�i��߶k��r��<����M���d |�� j�
+0=�@H�ñ*��IVvx`k����cLc>�s��'U���$B������1R�rDBփ�� �6��I����	����q�O��H�8U(��: �I�#��uzp����Ac����a$�<�s�i�O��ӻ5��0Y �\�n6�X�M�D���O�6�O��jA$j���"�(�Q"���`�WL_4�.\�V-�l����CÖ����4��b����O�d�O��b�A
$P<�0Q �5@�t�Ѡ$�<%�i1Μj�S�p�	e�'�`���"ݱ,r-H�- �zà@�[�\������Ip~J~�q�&8�$U��"�C�RMO
ϐ���iQM~� �9���u�'!�I�.�6�҄�:~j��.������I�\�I柘�i>a�'��7͎/VN���
�U���xA��MމU)V,2�D�ͦ��?Q'S�<ٴ(����'� u�g�P�X�[%�Rk��������Ju��A��t�9��q�� r����ڣW� � 7OJ�$�O�D�O���O��?�Ɂ�SHO�%��̟����hU�
ܟ|�I��)�4m��\y��w���OT!�wD�:D��Q��l�;!�a�Ф�O˓5웶Fs��I��6�5?y�䜑B�P�R桑�ut��CL$+�d�8e��O(�PO>1-O���O�$�O
Hx�AϑP0:���N-�v�p���O����<9Էi�D��p�'F��'��"ƞ\	��5p���b@]%�|�?�I�MS'�iXr�'�Zm\� �i.�i����(T�<���畗d�N�vc7?ͧ>�m��ʰ >Ɂ�M��!� Cg㙄@��hXV���o�0QgI9j
湨%���sy�[��8+$��Ŕs�8�Au��*��E�h�H#>��L���'-���F������죲I���#�J��SW��A�k+�&�[�
Z7C��)'j�N�C��s��%���S�le�vnɄ���tW-w��Uh� 
V���oA6e^2����ab���~��'��!o߲ѱ@(4θ�cJʠF��+���  xֈX�D(��}��Ӕt�T�!��#�\�񄑷N���Iy2�'��'F"�'T�$@@�Ιj���b�ޢZ&b��QN+>�'r�'K�Z�����F�����M{�� `�$o~�����M�+O"�3���O ��4p���8p�:ѣBf,I��-�#FQ�wP<��?���?�*O�PR7��u�T�'�:�Q��44ƴ 0��d(NT�V�|�t��<���Ov�d8�^�� � af�
�G���@,QW�%y��i�B�'�ɩ_3��(��0���O~����d�\�ڂK��V�K�;k���$� �I�C,J����4�� ���Y��� X�F�6/ڝ�M+,OVܺ$B���A�I������?��Ok̛ &Ũ,��-d
P�i�����'�Oа�O��>��D�ebH����M�I��c��4���̦�������	�?��Oʓ8��HH���
�Щ��K$@��i� ���'��R�O��?A�	���er#��,Ҽ,Q�'�/}�d�4�?���?9��� �Ifyb�'2�dH%X��TM��ׄ(ሊn��V�Ԭ���_�\��'>=�I�����,�lXKg��:m�ڣ\8���޴�?A ���	��	Jy��'0�Iʟ��
� ��e�U�r�-#��Bf��!�K>)��?A����%Lh�#��Ǡ{>t�P�eH����&Up}�[�,��b�П(���x��mj���>:�����JD�����g�	՟�����'|����o>��2cZ5���x5��%t"QeCj�l��?	H>Q���?释S+�~JGM=����U?>�����݃����O����OʓR󊹪�W?)�	Mh�`�������	���54r�iݴ�?�N>9��?yb�Ë�?y@i�Q}�A�$V�0�$��`	H��"J��M#���?I*OƬ��k�k�S�L�s�qb̀�[��uY��)��(�Ќ#�$�<�Ε��?�N~r�O�b�#ѥ�	`L�	�	�u`�l�ߴ��[�<I��o�����OZ�I�z~2�AN�RB E�y�.�Ɇ�6�M#(O2,z0��O�a'>��O��d�ZS����Ob��)j�W�5%�F`ݲ8��7��O��D�O��I��i>њ�c���@&N�s]�ɨ5F���M���?a����S��'��3��u.ݭ~Ų�$�ŤI1N7��O����O�U�%)i�i>���v?��k��HT.�1'l%����O\��+��|�'��sӰY	1ǜ�.����$� ;Eގ0'�i1Ҁ�s���>���)�	�9�Z�	�@�-�L
�@�s�Z�J<a��^g��?*O �$%+Zu��V�$|(���'	�2���<!��?q���'����;E�f���]*b*4I&,+v��V� 3�'�rT��I�E-Z��� Kb���ޅ�̜�2.��k�ʡn�����I���?1)O4\�E�iC2} ��H����fIռW��8L<A������O�ak��|���)�P��	�\�b�']t���qļiW�O�Ī<�%Ȃe�	�)�T�S����$Qʌ��%S��7��O���?������i�O��d��k�ӗJ�ҥ"����<W�}I g� |Љ'x�P��a�*�Ӻ{�ț2;�z���U�_�dk����}�'�erD�x�r`�O<��O���iz\<� o\�IД�@ͮ�h�n�Ky��'D�A7�i-��i0,��S-��@�e���)ݴ\��qB��i���'u��O`�O�)AZ���Ƭ�֔	��G��n�o��,����L$���<��c沜H��A�~H
lhe�Z'$����P�i���'��KGW�O�	�O��	9�^4��a$/��!�%MڞDײ6m�O2�O�e��y��'�r�'�^���'J�jR�\OpAH�)n�T�D<oLZ��'�������'�Zc��Yփ�)M� yv�_�G'� �O����;O��$�O����O��d�<�'N�j���"ŏ5��ͪ��+����P���'A_���	� �ɳ���4�ރ\���ï��tD^�C��w�$��џX�	��l�	By�XW���W6.��f�_�rl���Z&T�T7ͧ<i�����O����OZX@8Ox\���O��-���Y�!��RЦ������	��X�'RD9zt$�~������H
h���KD	��k. ���ئ��I^y�'�b�'���'�I6k*]i�M'\ ��b2��fm����NП��IjyRo�5��'�?q���:�H�\�4@��1(�0��4�S��I�D�I�(��*n�0��TyRڟNX�"��,U������)Z����i]�QI����4�?����?q�',Z�i�Av�sk���G�0u���#Wjl���D�O��?OF���y���9y�}b���(�P� ��۟cI���,O��7-�O����OT�	�s}BT�,�S�F���A23'�CJЩ!�(�Mk�ȋ�<�H>�����'�V$It)���6�˕�J�@lJ�A��~ӂ��OP���!B� ��'��I�L��c�`��윔c�I�2�_s�h�m��'��T������O��$�O`���8{�V���47]������M����Z�V��'Z�S� �i���F�_��.()tFA�����2¬>�ᮑ�<�.O���OR��<!B�D�9��hf�H�S��b��K280Ȧ���O��OZ���OR���^�"�$�C���8I:��g��2@�<����?�����۱b� ϧq6HP�Fΐ=1�b�)2��cc|�&�@�Ip���D���+@
���J�Q�2Z)f��#Ę5#�O@�D�O*��<)G�ˡ'�O��x�N�>�$!i6D�%lԀ��6 }Ӑ�?�D�O����)B���R�P��cA�;t̞TPv�o�f���O*�-8�����'"��C��6��udY�m	�bV��f�O���O�P52O��O8��C�$�P`l�/xt`��@!M`6m�<�"eDw��~��� ��`R#�?PG���`E�b
��b�h���O��@�=O^�O��>� �UqU��50[^�����l>��i뚝�vkӸ��O��d���l%�����R�8e �n�DQ���C�.~Ӥ���4&������O��ĸK/t8cPgޣ~~d�启_�7��O��D�O��+��Cv��ߟt��C?�E/]�*��;�Ɩ ^��F�HƦ�'��S�%n���?��?A�"Q"k��ِ��� aѢ�ʆ�Ƹ]��&�'jP�C:���O��d%��Ʈ��R�Ѫ´�a��S'$�h}�1[�|��Gh�(�'X��'�T�th�#��eʞ�(BD�J�F�c��Z�}��B�}��'��'���'L�h*4�Ŗ.u8�can�A�dh���y2W���	�X��\y��On��S��
�'��g �B	�0�^��?	���䓾?��b������\����E<%F�%J�K79�Q��Z�0���� ��vy����kL|�CC�)7��	ޤj���Â�}��&�'��'�2�'nD�Z�'�V�\y�HM�|�#3�XS��mZ̟��I~yb��8��������\B �0e:��S���^e���/[}��'���'}�50�'��'��I��L��>lIŭG�o���Q����D˘�M�X?����?m��O��*aI�.%2� �hƙu��LB��i$��'�f�y��'��'%q�b�`�mB�i��)��+#�T��ıi�&u�6�p�����O"�D��>Y��9b,�Q�H�jߠ�3s�	�'�&B�>�OB�?!�	�z�37*����5%k�]���4�?���?���W�E�Od�D��4�"�R�_(�1����#)�9�|ӂ�OR��5O�S� ��ԟ�ԋe� �uN�.!���P�W�M��j~��$�O��OkL�d��E
3��^�`�6�F-�I$K�ޤ�Iuy��'�"�'��I"#���V;1K�����7K� k�
Y���'�|��'��:C�$�[&��(J"�"�)��'a��ݟ��	̟��'z"�(҇q>��fǗ/#�(�3`.Ȳ}a� �w�>)���hOL���G����/u)�H��)�Q�#��>h��0m�ڟ���Ɵ���ZyD�B���He�P�i�Nܳ��GG<*�1��W�G{r�'�h|�!�'���O�M$h�kpxb�Xej�i4�i�"�'��	�{�$�	L|Z�����4X�f�E�K�����Zv��>��;�����S�t�?&X�\��G.ļI�* �M���?Aׂѷ�?9��?���:*Ok��13��L��Qp�}�r+݈A��v�'�b.��OB�>�X��U��[�Ϝ�+J�Y�d&��sr8M���)� �cԹs	���>��H񳄬�Q@,:2��"'I�ȓ]���Kc��m����'���f>X�BuOɸ>
�i9FJ�u��(	� C$N��|���y��!9����z4�M�2U�L��t���B��n	�w?*M2�J�Ck`�!��F�%�΀� �)y������2�;Cm�kz�rH�F��S�O�i82�9�Cȿx�Z!b��@2l�����?���?S�����Oh�Ӿ5��hC�R�	B��ࠉ�(;�,�B-s��-����;gF��)��O�%BWĚ��Z�kqeS����z7 S�=D��8�j��22� sIW�Mj���"������{aJ�s���-Q�qx���V�h���O��=1�r��n�\XB��4;�cA@I1�y���#�ܴ��@��D����Ҙ'���Ğ5dh2$�'hb�F�6��Q	pB�~�p��wF�F+��'�, �g�'w�4�P�c-��n��<�e��F%�6�8VND��G\~��P"��o�x"�ɃE:$KSD�/s}ʼ�B�iȼ8�b$��5�&���ꙹt��<S�;������ė'�xA�� d Y(&bY�|� �yB�'���!#ٍ�zT�E��w���9�'k�6��$1p�k�Ĺp�*�#�R��$�<�ѯȷ1��Iʟ��O�,Mqf�'�b<�W�xRT 5�"Q����D�'�"D�j�F�o�n������O��g����h<|�`���_�\}��KG��I�T��a�
�<�2�@^�O��Qѡ�SL�i`���@} L������Od��'ڧ�?�GG��5K t�!i[%��]��`�`�<х�@�6<x���҄r<��7�x�H��dM�<z�����^�Mr4�g,W"X��mן��Iߟb6��?��t����d���<�݋
Z(�#�L02�S�b�}��s̚��I�#�|����%�3���s$�W��Y�ȵ+��/]�bt�X�F0�s��y���?�3�/Lk�0�!V�nE ��4��L��b���<��t�g�ɿ���q��!>l8�Z�Ɣ m��B�	�n��\�M1'}���ӣV0��e���"|�0�ŕYRڀ��%+��Pq��T� �%���?!���?��'��n�O��$m>Œ�c�	j����o@�uQ���zR�,��ŁtŐ���Nx�`�Ƥ�P�Y2�	�)a�� &H׃;OD	��<#�jsU��Ux���À���͉J�:��^�K:�d�O���0�	_��~��d9��1�D��!�C� a���ʙ�� �gX��C$F	�N?��<��Y��'z����ab�'4��˦�eJCB:s�>UY�Mzr0O.y0�'��1��+ �'�ɧ� j��f@j>�Ń��͚4T��RC�'RvI��2cͮ�`���$J�]�jI��Q��p<��ӟ�'�,�d�	
,�� I�}-�9 �h:D��yVj�� s�G��ƙt+>�$��4ix@�U)$1x��dLA�!��)�<����"�V�'E?yࠌ�Ol�hэ�9Vs�(����}璘�Ջ�OX��N+���)�|�'�:��V�@53ʄ�5(^�`��M��pf�<�S�'슥�V���i6�!a�+�L�O |��'1O�LP�q�ʗ�.�P� �T��ɩ�"O*2c�=5B�UIǁ�I�����'8"=�`ĝ8֍��q���΋>M����'�b�':��ũ�;{b�'��2Og�ǵ(�J��ѥ�?{�Q��n��Q�1O�����'q2�(F���uT�@��(��]�{R(I���<�aAD�p�fT8��i�P��H�#��'�P��S�g��-|��@U����T��d��b�C��GalU�V�߷z9���0�{!��
��"|B�h�:�L�q��P�K�-�a����iߴ�?���?��'��O6�Da>�c������� _Fƨ�U�Fv\�B�	&&�u�5��D"�yc�O�<_ �s��=�h�5�H�P	[wMO�q�xu��DڜP1���6�Opm �W�7ji�6iǭx�FI��"OJ���"�=�P@q��%�$����D�`�{;>#'�iR�'�,�3�[D:S#Ąxl�pd�'s󤐙3>b�'���щmv�|�pz �H����h�����p<�֥Ts��M�.�ZEFI*��b�3n�����sx@��(��O�a�H�e(W�o�2Q��MӽUL!��T5Q[���r�I�hc�FӾ��sO��lZ$R:�QI!� TaN�SA�O�b� h�eT��M����?1ΟN�ڳ�'��Q�G�Γ���Z�řp�B4QR�'�鑱c���T>�q,x�;OCB1"g/	�P�N��O�8�)��.n4��	�E�?��%��UI��>���[П<�<�B�+�K� ��	Kr�T� g�\�<	d���Kj��4��R%<<"�@n�����$ab}��F�7�~`@6��El��L�	ޟ�)cF�����	�|���<���?��DC��R���֭M%ڍ�����{A�y��~�lƿe��`ʄCu�E0�{�牡��<�w�	�^��a�7d�![ 㔱�'c�!{�S�g�	�L~ɰ��
w,���m�B�Ɂ4p`��G�_��x�)�32\��JA��"|J@�=�Te�3��A��c�Α�N�ctLJ��?a���?)�D�n�OB�$y>!3�)�wJ)��m�#c&p=�7�]��C�	�  ��%����<R���q�����/����H&!� �&�B������'s��D�O"�O��$�O.⟼	TI�	�,����K�H�h+D�X�s�I��݊�O��J������'Mr���d9R���n����I(���` ��Q���D`;H��	�<!A������|Z�!<*���G��$/$���L��_�6dSaW���zc悧@���M*x\�z�-��(��xv��9=R��j%�&=7j�ȧ�ܵ�(������Io�ɽb$�AOX�Z� �#A&��;�C�ɧ_�m���3?�����jφC�	�M3��Mb4#���
)`ʈ1��VC̓gx�y ��i�R�'!��!����|2\0Cw�N�f��FEy�����O�8S��Ovc��g~ �V�S��� @b�K���	�;J�3o���!�*r?��QH��G�$\i�j@i3P<¦�"}��Հ�?��y���CΚp*����4{,`  �F���y�Â)g�VbၦpȲ�k� M�lў���HO��U��6Z�@�V,�X�A��(Z�����|�	���]��럨�I������a�RlN0:`�Q+���DU�\x�\f�g:p̅�ɶ#�L3��S8��!׍�A
�㞌��)<O2qP3�X�a�tq� ��p��R�7�ɻ
x���|�,��g���+!*�H��Q'��y��P&�Rpz��ܖX�4��o#?�)§�5YǨ� ¼H��jߡ"����כv�t	���?��yҰ�8���O�ӊk���j\*nH�6ОuՖ�: �'����� �@�s��q���1 "�J�$�\�s��9p�k�M²��	ec�%Ȕ�$"�O���h�e��A�R��� S"OLp�d�=��\���5�ԭ3��di�3��(U�i�"�'
�i8s�+=�f��aH،l�6����'��V!�2�'L�i�0�h��0��H��B&brӦ�7bګj��AŢA�����'��C�[�"�F�$��^��fb@/p��X�d߀=H�i�(O��p<Ib`�ҟ�%�{�	T�.8|h6Iύu�N���4D�`�'ڲ|����o�,�<��v�3��޴���$.	J����Ŧp�<yd	���f�'�2�?	����Ol����@*u!�h�h�����O�����U���/�|�'��hk0��ra{&�_?I�$M�N�0�5�0�S��IZ氳W�̆B��M�G���|��Oā�"�'%1O��	���U"�
�j޲���w"O �iTX�Pzv|ڦg�G�Pq��'?<"=y��G�	���"9ʦ��Bf��FG.$��4�?����?�a�T�{?�e����?���?�;0].@�FU�l��	� -ʖ\�21!H>���`�������$��9q�9`a
#�� ����RI��'�1��2dVU#b�I�٪���'�z` �%t*�H���]�s�N(��g���n�ʟXs��蟬�I~�'��i�'̀؋SMӡ���n®�B�'����J�7( ����煢R��9�O�o��M������?)�Z˧4c�-҃I�*#d��s�'J��-�v/5�������?���?ᑱ��D�O��S-c����I!$�	�BF�`��P�2$�+6�Dk!JdD��C�'%rd���Y.@~�	鴤]0�5�K��LXD}���| �(��_8�|	�͊��L����� *�(Pr��x� �D�%Rܴ��'�c?�8��7:-��V]X�,H�.=D��:�d�3!z�|�'�ӐP���Ǆ<�	���D9�W�ө{��=�g��,vYT�)�$��U��C�I+n�ȝ� G�u>}�� O \	�C䉿2�l���!�\���R�}��C����di�o��h��c���C�ɹjA�@we�*���5'�k��C�	0?����]Nf�hP�Ο�r-^C�I�8!hx;�oļ%{����'\XF�B�	�}�d�v��*����/�vB�I����#%/O��p	۸&�@���.,-R���H�`�h�ν^�°�ȓs>���Jf\��d�R.yʸ��:����Q�|�px ��TC�����^!X�J)"�|@�� :t(�x�ȓ�xIk��`129��+9x`f9�ȓ%��@%W6d�J Hg�R3!P=��.���(��H�X@G֚q�I��J $ 9l�9�*�Ö���S�Q�ȓHS�(� [T&tC��݊lKxL��QSZ �R��<
+&��Tl�n�⬅ȓ�T	S3�P2/(z$�uc�獡�KQ>��i�kžf8h�@_�c�!�䞷s̚�:���"x�:�5�Y�`�!�ĕ�<�^�BeqB��T�N�l!�$O�h�$���F`��Tp�ʑx�!򄀁���p�^�uب�q3�Y.Q|!�X�Y�$��o�0w�0B�]�[f!�$�.o*�s��J��<(a�޾H!�dH��� 3i�55��Q Ԃ��Q8!��Ȉ,
E����
���� A	+6K!�$�lπ����	�U,�t�M�u!�䍂F΅��D�:A�* ��n������=��z��~��Z$�J<�%�L�؁i�L��y��[,1�N� OO�@�j,����?Q�=����Dѣo^L�h�5Ad�E�`��N	�{_��'���D)y��4y5��-{�D�Q�'�D!�&d5Bђ;�K�6v�x �B�H��F�tC[���Y�f��ZX���
�y
� �A؂!�1bq��
ҧJ�C�҄��)<�=)���O2)+$�,Z���I�`)<dj�"O0}K��A�����ʓ��|@��'Q� @)�HX�|J�O�1@/p3Ǉ�!��a��>�Or�|������'t�yа(�,'X�d��d(�sӝ<��Be�C�9� �ȓ��\��L�f�*�B�P��D��3���;�C�2�xx�l�lJՄȓ=�p�BwN�#2����� ��9���dX SJϐ���_m�����91��)"��L���rK�����aQ��JJP���AM�k�`q�ȓZ��əA�Q�N.N��,Z'�t�ȓ!b��&Ng��p��ސ�ȓ0�,��O3 *Հn���!�,�S��4qwصi��[0u��$�г� ��h�:X�c&ʣd���e휅�J6 E�QD��1�6؇ȓF�Ԓ��?�.)R�N�;�>I��}�Pq+a&�TP҇A��"s2���� kl�
�dU��I��p1�ȓwCZ���!Ƅs��`S��D=1�T��:�dqqf��Z<;�9h���i�Z���NJ�cq�	# ϛ� ��ȓx��in�A��,{���&�~�ȓB�(��KJ���RDB>4h�ȓl�ٓ�N��^�:ĠD�jthԄȓ57�(pq�@�^�^	�Dl8ԡ�ȓ)C�����?D�0��]�D P�����!B��dA�軃���ꘇ�X�����p=��a�h`��7��"�ϖ�/�=���	���ȓ�"�А�K�n�� ���(=��a#)[�h��!��-��F�j݅ȓ
�%��А?C\`@�R�G%U��,(@�3Lģb>6�N'(|A��'C0(ʃ�A\�8�3H�jC��c�'Z���Q�������"�&$"��
�'��슐)Ӧ[����K,kz�{�'!���B���	 �}�bj�G2Je �'�p�'HB�p�����_�T�У�'�X�h&���c����Ɣ3�'�ni���6|)��0 j��!�;	�'6���爴O�q8�GS
	vH+	�']y���[G����E�lP�s�'���&N���Dٕ��e$ԁ�'��`��/@��ͣ�ğ!Yz����'t�C��	l`��O	=T (\�'d�X$)H2 �2�� �V��4��-2H�A�$ (KH��ě�]�~ݘ�	_G��a�I)E�axr��.H�"@x�m�
EZ�AN�Y���n�ER$�� gͲ����&�hg% ��d��O��|���'H���� w�8�{`�1�l6�
w��j%��8㣏.-����3��$�t�X H4>i�d㗭m�r,s�LH?��%�|M�c8�3�'0�}ڐBݱ[.X�P�g:\C�� #8�i�1bL[*
����.�ƨ#��$+�$�%����>�@n�ȼ�Eo&����g��b�Ȱ��,~��ITDG<���T�-���S%��gQT���ZF�!�DA�M�����P2wor��f��M��ɣ`��ĸ��W%��	H��i�Q�@���5uÀ����4[�!��>>U��nI�U��(� �D�/��@�a�Rg}�E�D/�]���y��T5N��E��:���0�F%�x"�PO���A��b�tD��*Nv�Pw�),j�h6�!�O0�kЂu4j���g�	ݜ�R�'� ���k��:�xl�f��>� �� *H.4TN@9v$�"x���G"O>�c�JX���B��2hȒ��$`!�U+>2D�%ą�ȟ ��Ċ*Ni��J)�1�j)CA"O`	�kW�\��@ǂ5��݀C��T�f��'0�Yd��Ϙ'^z8q���� ԈtB0L��h<�VX<�RÈ�&�¢W�:ux'�.
p^�*���%$�q15�'��zbTg�6%KS�I6X�j=k�_��c4)X�nE����[���Q懂[�Рf��ES<A�48D�p ���)B,��Wj��?_�i@��4D����P��j�kIi��d@v�7D�pr�26�x�"�A P	¤X� 2D������C����E�ߣG�Ҩ8g�=D��"W
K�d���1�b�S�n1p�.!D��x%��sКA�F*c�9��@)D�����	;V0�b%"\��d0�+D�p�畽Ms��ɵ��8i�� �PH'{qN���'�h�ӆ�'(vY+�aԏk���Cn��nd��H>�n��jl�(&����|R��o�b9�4��!IEl�QBMZ�!�p�"OH��F־?&��T�#ڬT������nϴX��+)9����ׄ3��rD��n>�3\Լ����FEj5����;612C㉕i5#7&��C�����6c����iA6뢹zbC�)��j�Θ�mc�&#�i��y��ƣ�|�{�,ݭQ"�IK��N���<9,ܯU*�i�O��ٷ �"���J�D��X�<q`���y�H"�D�`���#�7F����3�ɿ�؀s	Ѕ=��dyPcG:�O�D9�cO�'f�e{To,r���؇M�?Th���F 'k�\5��Ɯ2z�N��E�Ό���d���87m�-���[�c��Hưh�yk��}�V�+7��f�ї����F��4��y �m8���V��9uȎ�1�OT!$��bf�u�@Hɐo�rK�j�"&: �*`�C�oD��!O�$)�-a��[�g?a@� )*zr���^��X�
fN�Jx���7_���'Sl�	 ��+H��PtE8f��7Ɇ� �z��҅�9%�d�`�%�*����䞙$�j|�w��!EI����`��a�'A���'`�sܓ$���P6���h7L%��28E�h�'O��x�a�	\�x��!�_���DT�O�Ɛ���d�J�o�0T��=�7ʐ3|b�|�0��L���$k�O8��w��i�G4+����@.�xr�P�'��Y��Vk�h}�� _�����P�a�D�`��'az�2�O����sӴT���]�t�  �D�;M�Q�"O�M2Al˗
@ҕX�ֲp+&���R� KSj��B��T�k�0hAY�����V
K�8�Aw�2��"��,G�*A�ϓ������N�L���s���c�<rN��"��!L� |�㉵:p��8�ùy�h�x��!2�8[��"D�@]�y�ıe&W������"D�Xku#�)G��Z��U)Y&��>D�D�#���L8��g�5�`�=D��`� ���������8-�2�"=���:)���>=�@�Gu��ӧC���H�);D�pp,��PqJ�( �*Ls�<��:�I�#��}��ɭU�r��'�1Yʴp[C$�:�C�I�&�L���-M:')���c8��)�ȅ}<�Rl38F |@�dFU�Hŭ�Vx�\ 1dGF̓Ǣ�KEg0���� !�/�e��;���v�D����&by���$����b@�SܧY�\sfF�3U�� �ȩCX��&E��R@�r�h�`����~�\��?QSO�	�0<�����0A0���	&�z���!�Sh<��g�>��c���DRE�_�H��1�'^����F� �4|'l�����ϓ�$\R�yr��_-T���n�?d!��4����y��Y�L=�!�˯W ��ãE�0��S(������FKCh��S�*;}fI�7f���y"�E�g%�1�UjKr+��)��'�D`p��'����B��/(�P{OH2h�T�K�'�©V��9�BQ��3^RY"W/��x«I ������Ť|�4�Цן�y
� 0�*������"tnN	���:�"O�к��YD���FoL Q�08Qb"O>�S��ˬ]�W��%j�L��"O<��B��	WH�凅�H�!��"OP�W�Vfy��y��
&��d��"O$����Ŧ|^Dhf�֎H0Z�q�"OP�a�֤�|9;��Ѻ'PL��"O�����A�9�j=�"�Oʥ"Ola8�b 3":�]{U 2o�̛�"O �խ,��{cc5ٲ�93"O��4���O���M�7�Р�"O*Lز@�q�X�J��ƅY� 1�"O��a����ii�e�FO��}	�"O���
�
j����ٸ9�<��0D�1���j&��W��1;�)��B0D�� �m��4ے *���+��h��1D���X	�Mq�$S�H��Ӄ�:D� R�d�
{^ыѤQ8i$H�C*O�� ��'2��qK�G���Ku"ODAX�D�a�t�A�EP�M�ƕ�"O�tB�H�D��U%D(H���	D"O�yS""��a��«9�fT� "O6�;�S:9
�e
U��V�
�pa"O���@uhw(��N 4�R%��q�<у �^����s��j�gBd�<ѓaU��6�����zg��Y�<�t/�b�B}C�B?X���ID�Z�<�QnۓF���EߒZ�d�i%�l�<ّ�V�~�Bd�BE��=.*tA��~�<!��î%��p�ïP�����'~�<a(5r�	��A�?@�|��KQO�<��2���4�	5a����J�<�Âʷ�椐�O�.�W�x�$B�Ɇ [4lb�M�Jn��U�A4xM�C�I�I��@�O�+�45��C�H��C�I�e&0`�AIt"�*���g��C�ɇc�p{�^�%b���֪o C�I�x�w��n��`pw�	�?;4C�	NCʸ+��E3>�� ��nƎea�C�IxD0��k�1`e��$,��($`C�" �����9A�`�bb�.&^C�I�!�`BmC��n�ig%��nC�	�V{��UD�X�>@�U-%�bC�Zx��r��G-/Bh�4"��	�JC���N)!�:����]�8~؇ȓt�~�2�/Ѡa��*���w�: �ȓ0�zD��CI�N� x��Șn���vm�,��˝b�"��DkM�y��$��.�f�{��V5 ;���U��Յȓ{�șd	ȺR|\4 �gA�,�i�ȓa��(b�5[e�K�kC�Y�ȓ$�d�T�B�,>h����H�]����VEl� G�Iz-8P���H�r��/3}���|)��'ʊ�[�D�ȓ)i*�Sa��L_����IĞh8�ȓO�&Ay��{&�����7���'����D�� sv<ag�\�}�f4�ȓd�(�@rL����Iqg�$f�@�ȓ*�5��,*�ȳ*&��ȓM�B���A�9Wۊ��!�Ժ@�|]�ȓSpH�eBU�Z�x�PQ�؊X���|��ɦ�L*aU��Pf�}xŇ�(W��YoU�H��ѳ�U(CT,X�ȓKV��p� _���ۃn���:$��S�? *8*�'׉�
9AR"�1�"h��"OUyb�
���*�@�wy>Q�w"O�A���V�(l�P)��@��qA"Oܨ*uW.T��5Iv�ؚ'�>��"O*�R��pl`e�����ҴXe"OX����`�
\�t��?���r�"O	Z�ˮ�qD&X�8�8���y�U����D�؊�4��g��y�����ɉvT�w�\�he�v���`v�ـ�L2@u�P��˧M@L��YdP�8L��r}�H��˺u���D��橌�"��a���"0_�!��_��Lca� C��f�2���ȓd�D�C!� �,�.$���8/���ȓ9��$&£Ң���J�>�n���~H����^� ̱%ME�#����,����(�&�*��
\�bJf���[�r}��͔9R�-��C�J�Э�ȓ |�y�$@�-�.5��ɍ�m52ŅȓBPl;#)"�p�j@�e�L��ȓ@d��p��Qsp�+�ŀ!��E�ȓu�UZ��:"�,���'Vz8��'�V��ek�8���c�,��5p�̄�mU ��u@	]Z.� �bą~d�l����肣r}��fYHu�ȓ�x��cR83]�8(S���E5
8��x�Es�i��F7v|��Ȑ7��U��.jH�����1I�ĸ禎�+i��ȓkٔ��5Q)dj�5���y���ȓ=�ya�@�cmDѳE�BX���ȓ�����G�1cB�c��+1�C�	 �����̩tK��� �HB� yt���_,]���H-gTC�I�O�(�C�/w��IT*ڠ.�B�	�;!dD@��Y6�Ԁ�§9�C䉎ip2�a@W'Z8����e��sZ�C�#`�k���<M��Ţ�
ʏK�B�	>Y�l�af��-�`���ŝ�!�B䉸,Ʀ��E`%M���K��N0݂B��!���!��ݵoL�i��&�7_��C�	9I|l]3��]f��h��VfzC�=;St)��'>���b�Ԅz�VC�%6D60"�E%K���XVL�#< B��4}6�`F#�O\@��� 0;۾B�ɂ��(���B 	j��Nњr��B�ɿhS)���˾:�4I궫
6;u�B�	O�u��c�� P��fK�u�C�I 2l9��d�4,06K�7tk�C�I�}s�AV����K���t�C�ɮB��$�(ug2�PBG5u RB䉤V��a�k�8nL*P�UH�1�B�I'!֡��:�@[�/����B䉾_��s�f��3���hy�C�ɀ�`��G�)*d\񥋂�[�C�%�ܹx��J;4:p�C�[63�hC�0yjUP�+�
Z~c��3D�����T(�P�iR�]<h��h��*O��+@�g�����a�r�h�"O�S��Ut�B���S��C"O^8�tg�Vp ��`B��z7�4�6"Op��â�V��q��26�e"ON(��W;�N����F�H �01�"O�Xpv�	�V��$�e�a7>ݡ�"O0TZ4h�'0�pq2�v9P�"O� n����V e`r�cA@«1����u"Or�aP��Cj��ҠW^.2@��"Ol�p��>k��<�f��n�H��"O�Agm�)Luz���&�>r�
ЩA"O�5"5F�b�]�E���Z�"O�8## 0p��� $
�d��<�"Oؔ�K�\C�h��$@�X��Jg"O =Y�l�F��u�@��L��h��"O 5�f�MNH%K�T�y�5p�'��CC��0�F���zYK�'�1�� Y���uJaX�e�E�)��<٠�O0)NtT˅˜�($�C�@�<�d-�r���:��C�e!��ꡌv�<�Q��=4�m�3b�C�x�jҡ�W�<��Ґ.W�L��D?���,]U�<�7#X>*0�1�3-�<����K�N�<�$� Z��=���8���km�J�<��^
�R�����,!���-�k�<�Qϴ/�0�F�C4��i�3�h�<1C��- �%�WM�I����BA�`�<�$g�9nsF����j4,���N�Z�Ǧ�oZe�Sܧo����g��>jW,q�Κ#0�Ņȓ)fXa�'�0,�$�ހX��������?�'3�����qy5Y#��TB��'�`���Gr� ȗe"~�T@s���$ �O�i���#���:��Y��8ٱ�'6��&���	<N�y��h��\^��?D���2�ԛsj�H�j�v�N���)�I�{'�#<%?=xd�H1Y�
B��u��p`��<D��a�n]��4��q=5�咢*8D��9A�γ]Zb��'�N�Ȧe3D�`Хb�0F�r�����DM� K�l2D���3n�
%���h�\%#
��I��1D������"d�ZF��z��YK��3D���qK�?"��q0a������/�Ic���'@n�ЅK7O��
��IS>��ȓc��z&hH,�R�B�k�+Q�)�ȓj��y L R���a�M�]��,��U��Xq@��,bC�Tڄ�ۍKN���ȓF��<BQ'>u��]�
2��ȓL^���)���j����.58�ȓ- ���ÉP1��<��j[\T��?�b$��X� ���B@�po��ȓ=���R�g�6����,/�4��Ojx�3�K��I$�ǻL���ZP"O����ۇ8{(p�\ "Ohc!@�C�Z�	��:  �A��"O�J1�� R�Z�C 6g���"O�l�dT�*Ѥi��!���x�"OJ�8�"�%Tǰ��$B�9v�hd�!"O���`���g�ty)�!ʨ�]�g��nx�|���זijxI��B:���A�.D��c��6��L��NL�ݬQs��/D�<���6����/��}㊱H�	.D�����߂Q&>9�[���+D���7워vC��JgL_�2��bW�(D�8v�%|��`��?WC\A�Ѕ(D��(t��X(�0��GV}��:D�LA����.��j�g�8&M�� `�7D����%�I{J��D��5 ��
0�"D�����ξu��A%
H� �2D��q��N8+@a�1�\%=,��-6D� ��%:s��Y�Х1�EA��'D�H@�n;b��� g�/x-�Q"�#'D�� Zt��c�+Sw!��B��fR.�R1"O� �c��)���JA^�l� �)@"O@��v�=mz��` [������"O�M�T5HV
V��ō_n�<q���)@,8���aB�J��\E�<A�����*��IлꙠuWH�<9��@.�Ab�H0l�h��!N�X�<�2�Z��\��W̜�rG��"4kAI�<)Wl�v������l>^��'O�E�<�#��'����&�A�ySf�}�<i���!w�v�ӄ�
�H�j�q�En�<�`��Nv�EK$/4�@D��(k�<��i�L��k"�3�pu�_d�<Y��M7���Ā��Ĉ�\�<�#��Z���)^�Q�f�� U�<ѡ�$* tl���DrZ�J��S�<����TZҩ�v�1B��q:�]{�<qw'�:u�1�S�/K��;�.�w�<a�E��'O�A�@��}���J`Gv�<��N�!
�B�+�"�1X0`a�E�[�<i`͈��f�� J*y����b+�V�<�E J�)�d=yt��.�rPCf��T�<�F�@W��TAToaP�� 'T�ܢ@f��j,\��$�=��h�� D���aC�F�ʤ��ş�i�J�� D��SE�l���xFJ�� ��l���$D�HsBj9�v
f��^�65�E$D�|�	S
0<�\hBb���.D�Pɂ��%K�Q��JXz�
	��L-D���զU$'�Dp�O�{/Ԭۧ�5D��S�LJ^��s$�Q��T�SN5D����K��0,~ث�J�e�����2D������_���j�h��:��,D�,��D�V`4�J��]&JP�U�6!0D� �A�W�< �X8^c��h.D�0�� ���DB��D��)D�p��t�܄(�$���:-�'D��:��*H�j��~_Z  ��:D���ׁҜ~����ń�TX��m9D����Ę�{�l��ˁ����7�8D����EJ��0���e��X֞�915D�dz�O�%��ivY� {��2D��ঀ��I��Ր5�ݝ0Hl�8*%D��9����dh��p�`��J����%�&D�|K%�ɤV���J�j��FjE��	:D��s�f���z�&�[c/؂�jC䉳J�����XI5B�PG����*C�I�xJ���k���>��Q�$[�C�	4Zb�0�r�Ӛ,��|�U�� +��B��&>Ո}���#,3���R��eQ�B�	>m����G+m���kP�T=�C�I$c�^` �j��m5�ћs����C�	�g���q��&f�4�c��CU�C䉆@qdT�E,�k/\���ڳ)�C䉨"m%ZW)߃N�ճ�D�`�PC�I<Z��4i Bޔ\���q!��!B��%�9P�S�<���HSĻ��C�I?V'�0��
��S>�<:��N#�C�	�DFxMH��a��bv�N5�pB��Kf,��%W�ʀ�V�N�g'FB�I�Z�.2@ϛ=Z��B2 �6�B�)[i�P�,R.oԤ�+��·��B�	�OX���鈐rڽ�B���x��C�I�-8�w�
�N�l�!���C�)� ����7��ZD#Q�m�X8��"O�1е�
�`T����k�]"O�I��a��-�t�x0A�4���3"O\�S��J>
�X�G��u[R"O��7���m��;DO$v�"OХ�� �/)u�t��?����t"O\�.J�;i�A�m�(&��L�"O�0 ��h�X�K�j�)yd��"O����1q����6L�y\����"OZ@�pbgz�!cLV��҉!�"O HV%��K���� (r�(k"O�����ZQ]9Q��UO.e�b"O(��#Ű9]x��[�=�!P"O����E`�Tb�FN�f�"O@A2wg:&
��u��p�����"Oح���O�$lY���Y��8(�"ODlA���6t���?!��K�"OvT��]2!/x��TA�5o���f"Od��&ڗH�	uɁ$a��܋�"On)c�a\l�!���:1��s�"Ojm��f�jǊH���f���2"O\��c�L�j�p	�����;�"O��T��@��b�ژn,D��2r���(�$�#��H"�VA8B-D��Ũ�:��͓� ��o]��&�+D���UL��b����ܚf�k�)/D�4�R���w��S'f4SI��s"�,D�p�F�HCdÕX�Jr�y�`,D�� c�k[`�#�/^������4D�S�j(l��x 4���*�Jd�/D�@ɥ�B�ЮɒW�e�	�$N:D��S��Љ^�y���N����)9D�db�i
,C���g�V�>��e�$A"D��@��u�J��Ԁ
�+N|e�B� D�0�����^�B+J�yz ���I=D������a��Ȁ��˂"��dm(D���'�A/|��a�$J
�?��u�+D�P�0��D���nJ=4:��2��6D��2��5��pۅ��9E��� �4D�tȐ��0/X�UK]��ԠhCo5D����	X+b͚��X�lzs�'D�!�En�US��ͻK���k%)D��2FN=a$L��$�,W���R��'D�tQG��P�,l�� ͙jDPT�&D��X��أP��Qq��V�Y�z�9B6D��r�!��w�@aYiӧBD\���7D��`qJFu\epŎP�K�\)��6D��A���Rt, m~0��>3�!�_�<�|�`���!��D��LC!�D���t�5���j����P*!�d�,����C�&�AkT��#t!��M3+=�9;'-�;�I�f����G4bL�����f�IS�3�yR�+Up�pm�x�N|s��ݔ�y��Q)6$� �6IY��䥇��yB+��1Xh�,�.$b��H�h���ybo��#!�KG�"y�u�#!D��y2D���V���ֺN�^u�Ư��yR�@4(�y q�ʃ0[$�b ��y�"�x�nD�D�^�vd�9��C��yb�Z]�6�r��E��$��B���y2�^�A��e��_�t|aj��y�I
E� ��*<�UX�^(�y�I'۪�J�&�7�lp�[��y
� �X�n�7�䉄��č��"OX��%d9P�BU�g�U�ͱS"On���O�n�B����z�<"O�����T�����ƛ����"O��i@�G�WЌ`���l}�5"O��ru�߽9���C��! �� 1�"Oja��N�e0��aD)��{�E��"O�}���K>�ig(-h����"O�M9�a��l�܅��ɔ:�d�"O�TKթ��DհU0�XL�"O�-��$�����+�/
�(�*$"O�E�6��"t���U�����"Ox\��m>9"�x2����1�!"O&�qլ];=�\�ʳN�(b�L5�'"Ol��������ZvO�����4"O6�jA�_'l�����N<El�墀"O��a��6R;^ ��섨1/�P�2"O|�C#�O�QQM�6'Lу0"O�aS�N1,_xh�����:$""Oq30�^3>���Eќ+��5"O�q�`��u�j(�Qc�(%�lY�"O�\CBo�k�pɄ�Sl�\��"O̹ф��QQ4B�X1�hB�"O�����'"v|PK�GN8�䐴"O6!+׏�\���
7��X�90 "O���a�ǁC���%�G�85�X��"O"s��
<x���ȥ/�~$��kw"O��{F'���ib4��3]��q��"Of�6(�X���e�g�0�d"On����6��$	��=ID"O ���(-v� DC�0nb�!V"O ������4�2��Q�[�"O���I�2��l��W�&��r"O�1aǖ6(���Ѣ6Һ�q"OҤ�c�΀n����uj^R6��C"OB��������C���Sk4ݫ�"O�X�ʚi���`�0dlbS"O�QY�
'e*|9���4����"O��Iv�ׂ~� ��rP���b�<��]�c��t�Dn���UH�<����&(Q��<-��P�%�D�<���"ᾴ��T�J��@ R}�<��A_8#tVmK��Ê>a�A��%|h<)�c�(`��P�T�$�Rؑ�D���y��̊]�R�p�#ŧ5���ܐ�y�nJ�==6`�-���4�Q4�y�C,B�=.Y��P��IgZi��'�D���N$G����*M�IhX�
	�'�p��HV<��B,F�.��q��'2U� �ٯC3����E�|��b�'mȽ#L��X]0d�e��=bYRH>)�yC\ɰ$��,HA�&&ڝӎ%�ȓC!�Y�G��M��zE��tL���ȓW�`����=ɸ���@�,�nA��(\~�"�c�J��}�!
(���* ��I���,Nm�@�Q�q*`(�ȓi���
�,��J[�li�����ȓW���d�#I�o�Z�ȓ� 
1&T?Zf*QR0� n���[
]#�B#O�����جE�"%���
����1,4�9��`Zޙ��N���!S#&�H1��m_�y𲀆ȓ{D�$FˆYs�n9t�&����zW�=�2Mͪp�%i�=sE�B�)� ʍ �1{s��P��ƄP&�L;�"O��ʱ�ӛ,�x���jX�Hr�tH�"Oؼ[�G_�VG���ָ&�@�"O����僝�x������RT"OXx��)�0ZT|{�E�����"O��
�%L�D]3T�׀,��tX��'0�'�"��>��&PZlza�֎���傀�z�Ih���O+�@���1}ڕP�I=\d �	�'f����O�7k��yf��D5�A	�'Zid�F���Q��%B8��)	�'��KbC;tt�3�@���D���' ��C���#u �x)��
�'X I �DB`����W��xCb�
�'�@cF��9(��`��lܪ�B�xJ>	������O��10UE�"s6��+T"�|�8��'��x��5X5kb�ɠC�U �'�rL��m��8��ҍďB�RY�'��|C6�#K.�a�MT4(��J
�'��`�!c�$(�I�TEP$1�.U�	�'��k���.*�4\c7�Y�/S���ʓ*xAw"�]�H� �,L�a��Gy2�'9�Oq�����Q k���LA��5*�"O�@�#�"wm���t�\*�jh	"O�+�� D�	JS$W�z��`6"O�q��}?�9Hр�S�9"O��(�i�\X����ܮ`J����"O����L"Lh%�ѡ� ��њ�"OT�S��5S�X�2��:[����A"Oxh���Fd,0���Ά>ftU)d"O�D�$�
$k}Z����[�)�jԒ"O���fV����R���4�����"OnHa���f���*D�T�[�V= R"O����`���d���S�X΄D��"O~m�B�X�
�喡Y�t�{�"Op��BB�M��3�$5F�r�S��'�����y7�m )}����L�\����5"O|�js�ڷ^ܔM��6I�X	X`"O�Ѕ������љ!��͢4"O�AC��ap���f�9�"u@�"O�a�ը�/=v��"�o��)�"O0�{0��1�T� R8J��� �'�1O��6�X�M9B|�#)��ة���'
���O\"����(��QS�*Id����^=�H�7o /VV	Ѵ�8��Ćȓ_���%��<�̘��&��\.2L��~/� �:F-�!��P5�ȓ��X1�Y6~bN�p���G(�8���
i��$i�4��2�Ԅ�ٟ��'�,�˗*���0�@%�ve���?���?�*OD�Ә'r����ߴ@I؅ZU	������'9�ճpb�pӮ��
R�fa����'R(���N,3_p@SͼV#pJ�'�ȁ�U�
����2�Cy���@�'��AK���&����Ȗ5&H�'
R�RF��m8{���9:���ߓ��{���+÷.0x��ٷF��tz�0�d6�Sܧa�6x���DN $륇qKh��ȓn����]*Ed~��R��U�U�ȓgrй{1nd�����q���y�:��sBNSZ^��S��Y���7�i�g�ޒ��ؐ�P2)�����D�9�u��_��0��Φ~v�F{B�O���dN*|`���VOǇ�0�
�'/F�K&Ռ
�j�&�۽���p
��� Q�B�œ>\���#JЫb0�8Zs"O���! �|:��f�U�)2���"O��ӭMe{��Ӣ�63�l��"O4x �	=G3H��G9�x8"O�K��\Dl�*�!שn|L�D�d,�S�	/eb
p�+9N��&/!h!�]��dh��65�D=��D&6-!�˟4]�qh�/F?����+'!򄈖ʼ�R!F�R%0��e�; �!��A�TD�U�9%lUMG�+!���2�*�!"� 1&�6���!�D@ y�z��B�C�8��ű���<kў(��Ӯ{.Ԛ!mO�j���D�E�a�����O��OĢ}��OP�h�2�܉WtX�I��Qu0��ȓd�v1�0E��%#�U�ޙ�R�*D���Al�?�蚇`1v[�	kA�*D�@� �S�Nl�to�3�T��A;D��aD�ė<Z�`6+�+b!  ;D��ad(� �B��N����Q��F>D�t�6 @�������F�C[�qpV!�O8ʓ��S�4��3M���k`a�8;`�QP��Ԧ	�!��?hq����23Fr��!�P��!���O�8܉��I�'- ��)��,z!�ĉ]9�90% -,T�hĘ?<!�.	 }��iB
�|8P�F�3!�_�~�R����T��h�E��B0Ofq�u��P�8@��:P�\�u�|�'U"��̇2*gHq�V�C���*O`�=E��\�$�a��άX)0M C�����'#az���Ɗ� �b d�D�С����y�I�
'x���L�J\�i1�Y��y��E�|ؐYY ǽS�z)��8�y��\,ft�R�ů;����Y���xR홼$��F�F=`�(�^�O���$@֦ ��LXX�P�T�Ͷ2x!�d���l����`Pt`0I�r�!���:�
`y�g�X�b����.�!���)[n��0`)���a��*P61�!�$̻T΢�6H��F�����B��!�$_�4<��BFL?ti�����#K���Ą
^����%��jʾ�He��b�C�I�]ġAanB4]ŲX(�nߦ+;�B�I0@Ö=q䯙Y$T�`t_�vB䉋\��Px%�Nt�Jl�d��f�.B�Tg��
�3]�B��غ"��B�s�\����@<6��R�|T��"O��X�H�n�{��Ԥ+S�5�P�'�ў"~JԠ�3]r�2vΏ���! UEΚ�yB�E+*9��s�K�	̬�*fښ�yB�U?)=R ��g@'T�`C℗�yZe����C��p�6G��B�	��� ˳.�-&��JF%��~�B�%KCX]´o��H`p��7��C�	�i����e�A�b������̃C��=!�'A"P�0B��$p�H���%�TD�Ӷ8L��sgݼ��i��F#AhB�	#>�$�Z�,ĲQ|a��ņIWB�I�X0 �&]�L�6���%��W��C䉧��TQ Ա6Q��R�	��C�<0*��)��@�_NX�E�[)�C��Dd �T�xhr� �pG~C�	�#�"P����j�(�Á��@�O����O���)ʢ(����hف/�Pr��ה\�!�D�l���S�˞�.f�k�h:|!�� 0�*ҪE�S_�xO�2�Ƞ�A"Op��Q���Y؄hS-O�Z�L	"O������ A�t��+W�}�	 1"Ob�R�� �@Pj��Tk�.a�Ԛv"O\zg���o���˲i�F]�u�@"O4���C�+���"�և���a"O`�zS)�PV��W+H##���`"OH�+�I	y�����JܺT"O޽��c8o�d�2I9?<l9�"O��ʠ�L3����I �(�kw"O�i�%G&Q���id��*�J�y"O��Q�b J�&!ҫG#�j���"Oh�!�K�a����J�E��4S"O��P1�@>(u����a[)���"O΀ӆ/L�n����!N�}�4���"OT�rtK�̐y1u@
=J	>:�"O��H��]%��B�O,N�8�`"O��[1&���8e/ˎ9���T"O�`��BN��X��ƖJ�iV"O�PSFY-A� �A�0C�6�;T"O@M`$�,F�X0�.л^rbEb"O���BOR���jvm&9���Q0"O.���,�<:�.Qb��p�l���"O�@"pgW;#p��
��L�{W"O�٢��޸V��	�FXg���R"O���$j�
H�p1�kT4�r��"OJQQ���>L��L��D�0��"Oh0YS@�,\ڦ��֡D�;�p9Q"O����E�	V���J��QZG"O.�XWe�!l�,�̅�(۔t��"OX���R5'�BN��$l�"Oz�����?[���rb��;�}"O\�hwB�9BNѹ��81�$��f"O�JD�Z%:�t��gE1�P�"O���ț+P�v���DK�(Z)"O(�	���]�<pY0��[F�q"O���v��:
��c��G�L��"O��!rBցseZ�Z0��V���"O��2���f*>%�Bf�?>�t��"O���� �:j@na�ń.J�j��"O^B�� b6��͟�h�,��7"O���+
���P��iB��3"O�����m�����>>iHE"O2	K&҂y��XB��.��sS"O��2����*�����ڟy�h]�%"O�[�D������,b�Zq�B"O6�#��LW�С�
�-�1+s"OȼA����"�uag�(,M��c�"Op��W`U������bM1.1�)��"O��p�Z�X�<!cB��N�J!	&"O�!�gJM�A�FDy3��$�Ej�"O���L'(�4�a�(:0�`V"O¡�!A�0]x�	Âw/ �F"Of��.^/�f�b�*&&!�(`�"O
U�&䉇<y�ywi�i(x	�"OؙT��L�@`����f�6�Ps"O�͢&�1N1��@ ��1o�1h�"OI�gJ@�UX�@jg˂3m��$"O��C��Ln�V�8�Ѣ:@�hA7"O�A2��B�B1�&)C�^a�4��U�O�*|;�D�K9��s�F3��,	
��yҥ
jȡR��2O��J��y���]U6�:�V,�ޔ����D!�O�ԏ��a��p�G��}��Z�"O� D�[V�H�4|P83��@?�j���"O��:�kW*H��Œ�aĎ�~8�"O�����΅W�<�X��&*���+�"O��!�`�={j�S���)u�~my!"Ox�a�o�)d�t����?9z�wS����	�L�I�֦_8j�:��	���Z���Od˓�0=A���JW I[V���^$*8�7�A�<��f�-l�� ��c$
^¹��ď}�<Y1f Bv��� Ýd��;2Wd�<���L�@;�g�-f�򬳱�b�<��t�n�AL��dU�I�b�^]h<�@-��h����s�)z=VLZ�F���?�/O���ėCR�D�q̓�}�D	 gH�)Q�'�a|��Y��BTY1ˎ�u�uD�:!�D؞=�Xb�.Ͻ0��E�'-!�Pa�6�)3�Pn�"Q!�Y1h��bsLȞx�4�*��!No!�DJ� 0u�b�C�:�G�.�!�DI�W4Yeo�p������ lY��w��A5���b`�Ԫ�^�a���J!�5D�xc!�*|�jŭ�Q�2YC��2D�����=$��h��J\�+�$=�d�"D���r�X+$�IG�v) Q��#+D� ���Ҡ$�¬ۑM��\`��`�<D��S��Jc�l!ʗM���[��9D�2Í�Pi:����Q.���@�a8���䓘��@�y��<А�'�()� �	D�!�d�&eD40ڷN�Zh�|���ŋ~�!�D����n��mY����X1P�!�D]&6�D�l3sP�L��MR��B�ɓ>�����l�P���i��$�B�.G="�C�q��Ac�~�vB�	D�B\&N���$}�&��>8�
��D{�Os��B��e�G1,&�`�@�?�!�Ej�H�v(uʈ�W�
d�!�
5u�y҃v���/��w!�ܟ^����U�5H�L�6���!��U�y����¨V�hy`�.R$;B�'�ў�>����I�u[Px�q�T66�d���&D��h���%�\�S6҂$���U,#���O4��!�'�?�sB�<"�탵 Q;D+��a3鐴�yB*W�,��}�6F�,;�h�H�J�	�y�_0E�B��O�.z��v��
�y�ET9yY��Su/S;/�k&�P��yb�0��
T!Q�+K�|S�Ɛ�y�jښ �p7Iȕ&�D��y�!
�9��)x�F3>�5�A����O�=�|Z��T�=�B�~��HZD�y�C?}
�*@L�+^�!
r��yBdO�T� U�a���O,C��A��y�A�3�tI�k��P �a���y�N�8j��[4O���kΥ�y�D�C5��F�W?�@M��@�9�䓜?����^69� �%�Ƿovyk3j��xb!��ϻ&��`3�d�c;~A6n�>cj!��J�%6��KΘt/��H�+А+k!��J�:�q2���/V
Pb�钊t-!�D�18O���%�|�'Zb�!�dXc�pت�OҶr�j�t��7�2O����eԤN���B#
&r�򜫷"O=:��L%������K�@�r��t"O"��K*Z����3Ii�Z�
�"O lj�S�U���n]>� k�"OllIwP.Kt�i�D� =��(6"O� ��r� d��bBmմv@&���O>4#1�Q��}hdd�	i�z���(D�L�G�A�x�^�c7�:X�>@Q�!D�lzcb�)m+n�y�l�2U��P�N ��ƈ����AȊ)S�bX��N�,7XڱP"O$KE"ږf���g-ϓs:��p"Oލ2CU%���h���TZ�E
�"O�T�F��g4hN��[B��u"O腹P*������'D�p���'!��_�Y��X��͂���(��/sm!�D_�ʖ!&`̅;���QҊ��kaxB׎�?Y�y")ܙ�@��H-_~�a[6�n��'�� �0�ћ
Q0�Q�.1�{
�'��I�T�F�(Sw#�.��A�
�'��)��N,�T}�FkU*+=��
�'׀��Тn��`��I�	NfJ9�)O�����!I4K�,δ6c�Di�	҈K�}���q1�S_��X��w�Lz5"�$�<)�.�eW0(K���?��������yw�K$]�&U���ZUH�����y��A�@N���J�4�b��y≖j2����N3����:�y��D x��P�դ���f��Ү���y��P�e6N_�|���!3�Y��y��W�'�5�$Oۓo��#"�.�y2Jؘ	����Հțc J�S􏁫�yb*�l��͚����
��ၓ�C3���hOtb�İ�M�jr�����"����v�$D�|
��S�L�N�:A@K�Z� �%D��sf�ұI$�(�T
K�FQ)vC䉟]A�E�rK3_�N���#�+P4�C�6z��M����;Q�V�Z��C9`��C��6:f�	� �4\��q���Y=�B�	�Rt\��c)��G~��
��u�0E{J?��p�w�� �E�;$V���"D�TB�o� 4�ʵ�`�F�w<�R� D��*��؄68P}C'��%jA�(X!�$�B��@c��ԲrC$,��V!�[5M9$,X�j��tG49�4�$>rO���e	�]~RT��cC1�|�h"O�Ը���!��!�P�m!e�˥&�On�=��:p�O�C�(��I�#\Ty@�'=�PnZ'b�h�w�J�,gN<#�'ꄌr���&rA��I�M9����'E�:CB��Z\R����ơ(�'�:�p4�Q�Ӑ%��(����@3�'o@(���jop�i4HT_��'��=XL'm�m	�B2u:Hȍ��'�a��`�����E`�'~���*�%ۑ�yBEf�@���Q�xY^qQu&���y�� �\!bSJ�"ot@ ਞ�y2	��(����a�/Q�aiw�Ɗ�y�HR	T%�Y2e��HyTmBg�W��y���Ai╠���uV� �f���yr�Ӡ+�l}I�dZ�;� ��v�Л�y�� 8|����,8�]!�fU��y�B�	� L�e��p���UK���y���:!yf�#�aT7Y0��� V'�y"�p��[U�V/',�I#���yk�S���fB�&4"D�܎�?	�'�|�z�+�:S�r!!a�,?g�h8�'��GI^�d<ɲ#/�=?yF�B�'�\��#�&L����)3x�h��'$�#��1D��t#Q�^�+�����'Ҡ���b�)E�1A76~�Qc��� ����Ɖ(���h-X��p�FV�d��}��GSe������]J,0�C)D��&@�$F)`�ӔjW:6�t�S#�,D���S/��~W��2PI�=v�E�v=D�4��B���f����e~�`j9D�H��]L)p��C+F)T@6D����/�L\[u��'T�#P�3D��G�QA`����-�b� ̲<����38�
�,ٗ-G�����(����H<2i8bN����a%�h�/RW�<�U��QeL	�S՘0H��amR�<I���P��I�C\��,C%!�V�<�r%_ X}�
U�Y�|!!f�ɍ�y�F�1����6
:.��;�#���y�+?�FXч��/�N��̐���>��O�A�5GD5$+�:roZ6�M�"OzYhOA$L��Q�N�*k�0�"O��ٕB�Da(��snM�{�^X�2"O��Yw��a�Jy�Po%u��=�"O��땯V"cF� ����+����"O��K'�^�$Ҽ�����.��u"O�H;��È\�l���:PT��"Oؙ9���x��k�%x���a"O��s�۾ej��Ґ J7`�B��#"O�� 6�<9��H	OB�Xy��"O���W��*zt�Y3w+W�P��j"OvIW�D�+%>���A����c"O�U�#�6F���bBC�*z�!�"O�d[�j��8*��L�'x��A�"O�9�c�M:odNE+�i,d�T�&"O4ؓ��>$<R����ʏ!P�10�"O�� �jPc�FnT D�'s�����YA���ƌ9DI��/4D��#��O�B���� _wS5�ǆ6D��Zu�^'�� �L�uG6D�p����{�l�JTA��X6(TH3D��{�aVi\����_Z�(āW�+D���"	��
B��6��WLPРqM/D�h�!΄ 1<�1m�3k@E�,D��8`
ܥP��4�'B[�)� �Q,D�\�S�R�>��e#�F,��:�%D������P��`7��8q贡u�1D�t ��C��ܹFg�6xiv�I#D�,3��t�&a�A,.hNE`�;D��H �ŞZ���D!^n`�2�L8D�0�g��5�@5K�b�w�j�Qu� D�hcs��~�H���ڊe�-E�4D�8���ÂN�ة��!	:��fm3D��j�N�s���bbÐa(�;'N1D�Y�НzTB��P:L��F�O
��Or�$�<�O�2���b�(ӌY�0`Z!9FQ��.D�t!& f���%�V-��a��'9D��I�&�6 gl�V&������#<D��95-�)���Vg��sA<8��;D�pc!!�)x "4bN� I6�iW�,D��Xc� *JG<AȆ	����RB 'D�؈㡟9kf��u�ų\�ބ8�c�O����O2�O�3�	�$n��ΊG�R���2=tPB�ɫ��#0���F����>v�VC�I�xl�) ԩV�	0q�RFJ�Z�@C�I�Y��Q�F��>p"�#fe̥\��C�	-i.�Lj4 N4;���`N=
jC�I"gʒ��G�ƚ�̠��j���C�ɩL�X���U[3�X��$H�˓�?�����S�π N�j!��!,2���$�>ZEF����.�S��B&�p ���ԸkD�D�����!�D�}� ��D�B(�&� l�!��).4Q'Ϗ}����\�C�!�ĉ4f���;Op��;��s�!�$�q���ʥd�]���Ss'Qw!�W(:��L��o���f\� l!�$�i쩑��ӫk�2|���r-�'����i��I >�&\�Po�a��%>)4!���0�fȂCb
�$5�X���ݩv!�$�vX,Ax�B�$-B�gK'U�!��H�XԈ�eo��A+�Y���B!�ZJ��9V�w5DX���:)�!�P�e���$H$��$Q";�!�����Ij���	���e$�%�!��8]��Mʅ"0f	 �(����>�!�D�?)�xba�[>-:f
�
(p�'�ў�>�TH�(6J*=x2�?(W0K�.D�����P%zn�P��]*��8��,D�d��;���ř�8|k�O7D�Q!.	�飧�m��Q1�0D��%eڬb(���En�u["K.��-�S�'d������F l�x��E�J�00�ȓp�m��お�n�"��4)?X��-�Ԡ�!MW�P��!�)�(A1�y��ڙA�×UO����5���ȓY��ЈC��2W� )�E�x2J�ȓHY����9S���H_�P<���)D��!k��^v�:��x%��f�<y���ӂ���� ԫR�%'U�y�HB�Ƀ|����Qv�:�q%����B�	�"N<�ϋ�aZ����H�B�	�mq����#n P �Q���*>C��		�Uc�%�L?�S0���1�C�ɜe&P:�MR9N�����h��Hq:C��+��t`��\m�j���(�;k�C�]�dHC��ߢa`*�9�ퟚN��C�	?P��x�⢊%DC 	[�
\4#��C�ɣ�N5R���=f�ř��<Vl^B�I�� |X�I&Tr�2��'m�DB�I�Wipxzd�ǎpQJ	��
���C�	�h;d������w��� ��	*0���=�Ş�����|P�1d�/�Lb�	�3]�!�d���u��-5[�D��	\�r�!��+s��9�0�E��<1�ć�;-!��2�TR�p<X��T�g(!�Z�$�
�Cc� �%�Y�U���"
�'���R��dxv��ԗ}*E
�'\�Q����Gn:�P��q�,X ��?���O�лU�L��Lܓ���6(ກht�"D��e�qjR(#Q�W�FvT�Pe^l�<��*�%�����]!@�j���\f�<Y6@�PV ec�'��{ ���x�<��þi6�s���<g��=xVo�<5��Zx�b�G�JXJi�.�k�<���,G ̘EØ5-�� 9��OyB�)"�O����c��kQ����!�
`SB-A�"O��IF _|	�A�p:P�*�"O�!r��r������+RG��W"O������v�fQ�aNQ�4��-z�"Ob��$��^m<q�wMܗ� d��"O���Q�Y�Mx�D1�K[�m�-x�"O��w#-M�t �D��������'aў�ST�'����O�(#�.8�U抶Pd���� �L��D�%^�>�ITH@;X��z��	ßdF������
92)ݏ8n��I��yb��'�0�'���c� � �	���y�GV�R���[�hQ���ܺ�y­]����"�J6P�B��G�ŵ�y�U���dA��W�@zX�����y�����!���J������y� �;7&̀a
�4?7V�� l_��O����O�b>��Q�	�<u(6 ̢[�RU�	2D��:�퍚0Hx����x�8!�s*/D���ڦ�"��H�P�X1�sJ"D��c�ɊZ�x5S��+9�VM;�!?D�4� ���H���0�|�Äi)<O"<A�&��mʃ�\K�d��+^u�<�%�(��Eg_) �嬘|�<)7�L`�`�E�=y�<LCf�Uy�<AE�^\� [�nX�
�&�J��y�<)�M�>�P��3d�*iz���o�<MJ&2r��pv�j��z"Qj�<!�N�o��j���EFD��M�N��k�'71O��Qr��Wt0��2�=�|%�W"Oָ�����y;C�dv���"O��Z��
�JE12ĭ=�� �"ObH(�%�"yV�A�@ �0ء"OV�hϚ O�2T�vK���Y[T"Of���Ĵ\q��+��� y�"O|Q�V5�������d��`�4"O�B�`�8��b��+�ȵa�"O���dk#���ʄ�Բ䆥��"O>��D���0���ꑳq4hs"O�T�#(Ww��L�QmJxZ�"O� U��R�uc�kرCe���"O"����*�P��
�_r��4"ODZ�DE
C�H8QT�[�N�L	��'}��%b�ʎ,C0��, ��b��2D�����*Ϛ�@�&l�$��)0D��SQB_�{���Aw
R�B�T���+D����W10�m�%MS��,��+D�$�6��]� eK�(��N�$�a�6D���e��N (�D�ɑf� ���A*D��0�F7��qG���6I�a&D�Ȩ�b� �:4���ghE���#D��I$l[%�:���đx�Ez��"D��@�Ss$��V)��Ϟ1b��!D�lGIN�V� �+�hA.R���a,D���ІQŊd�fG�"S�� �5D�����^!�\�W� �^-�8h�n5D�`Ö.�,J�2�J���G�n���>D��e%W�6��e�2V�@Dy��9D�,�RG�*f�<`���;t���`*D�� #&\�vE����|�>-*��#D��i�&��}��b�B��%D�4��*��,�6��eI
'z����$D��Y����d�(�(0k�)%�ּ&&D�`����i*���GcA61z��1�a$D�X��k��tQ��j�%��V^��Qi"D�x���ŚlW�=2�e��=���!J?D��)���&y"�9��"��]Q1�0D���6�R
>{*�P��0� rG�0D��i���Eڈ�7��)���A��.D�ْ�Tr.�rdB���dz4N-D��( ��:o�`���*�~)����*D�\�R ,5���aq���6����&D�ēBCʤ�9X��\5R삩��b#D�� �����!t�	QG�P�V�L���"Of  %J�cuX]C#��:���R"O�0uC]�!�DAh��#�
)��"O��aS`�c�!��.M#x��
f"Oh!4���u��u�t��7f�""O����A
g� ءf�:lQ�
W"Ol��5��
A�*l�`,�0@G�<�A"O` S�-ܩm�8\��a�E�"O`S��D~���E���	B��"O�|Rd �&=F�0�	кMS��A"O�M�Ε�b4&m��F��[<DlA�"O��cR�	�?#Z�`�fՄg�G"Ox%����#5��}D� E�6X�"O,�9���:�N ���?�tB�"O����n��'�Щ�3�U4�ذ�"OtE�P��(��\���
?�Zu��"O<�LJ�Gwbi�[�,�`XZ$"O`���ZL�R��R
�	J��	q�"O���%��	[.H�j��/ Ơ@"O
أ�@"6l
�货\���\b�"O�za�V��yHWǟ��$�""OL��u

7��Y�%�X8YyݐB"Oda�ƛ�T�(s�Y�,xj���"O�!��䏫f��M ��@r���"OA�d��
;lh�)�� �?U��q"O�6���~�V�Z�	
HB(H�"O h�
r�b}J��*M]ȩ��"Ov=��"<��hT��,fa4ȋ�"O$����
�^M*3g�>Q���w"O,t�G^�DP7��h���"O����	ˡ��dč=L����""Ob|��2u�� �@�(t�"Oވ"Q�N�#�`���N!n�X��"O\�P`[�
�d-Qg�T�W��X�"O���		Jb�8��ڏJNP�"O05 �/Â{9�@R ��+��P�6"O� *B��6a���{�hL�p"O���3mDO����"E��D����w"O�t�UBK�v�Z"p��G[	A!��6I��`�A,M���
�u�!�U+W��g,�`��`�e�<X�!���KTl��C-W�H�õj�,�!��94r!ӵ(ʽ�Tz��w�!�$[ ?��ġqNӬp���x���o!�@$(k�tz��h�j��@D͂}�!�֯+�k���(fbd E�

!�D�y�[�FO�#X�M�4d�&�!�d�.��!�%E I����b�0�!��?��%5�V�gH�Y�F⇸*!�$�����xi�5,)�Lɢ�I�N!�[�1{���� mP�ڤ	��!��?d~\-
V�:e����gI�u!�:��U�D�D-7��� 5-W!�Db�&�J׋��FU�'�#QE!�D� �<��Q�6������O2H�!�A�A��!��O^�ˬ��7�G�C~!�DCH���B&$����ѵg�_z!�dR� ���٦[�}1e�!"!�dJ-%P0ї胻 %��Rpd�q�!� �Fx���*R
ޜ(�M�<R�!�M��U���X3�����<�z���θ4J�A��
NV�;`E�]�XՅȓz�D�q�/�W�"H3jKq$� ��0@�E�ߢ!x~%8��C�ȶ���S�? haP��9M�����ω)F`��I"OPE�P�������N�:["�a"O$��b,���SS�_8C]�"O���FY
l�P�{�[&=�ʽ�p"O(�@*ԏ����J��l�ђ"O4$�`��D�����(oM��"O��A�[�K��ħ9���"O�f#��rՈ�矼=%^<�E"O8j���n"
!�˜;)���)D"O���dbT���W�=�b�`7"O�� �"&���)ж)��&�y�K��W���)V�ORkEQ�ڷ�y�R�zW�9y� G�D��fm���yrͿo�č��+��6ھ �Eo��y"L�`�Px�4�VE\x��$��y2l��%׾��T5
@&�T"�:�y� c��uSį�-��!�L��y2g@l2���Ͼ&A:4�^� �'T���t抖[�z-a��G�i���a�'���r��.y(��x�.]�v$Ԛ
�'B�Re�iG(9���7��	�'G���
�;Yb�#ݿb�l2
�'�ա KL@�dA�*�3GH(��
�'B��r����qpW�JU�~xp�'���Ca*�;zI�g��bO��'�l�Ą'v@9qw�ɋp<�=��'�F-0 )�	���֢ÀW��q�'B0�����M�� ��MS�Z����8{�t,s���WҰ���W�<��ǒPqZ���	O�j��mv�<q�م9����ι{C4��HDj�<�Ǉ�+mIZI��әmIڂHe�<�@�ʯ$F����chB�����b�<���ߖ� dp�BBEVёC^F�<�PٱA��1�5N�#YQ� J@�<���ÿ0��`�	]�R���)�x�<A�oֺr�fi�p�J
�b����G]�<�vk_LP�����:���2NKU�<�Dnĭk��t���?Q�FL �A�O�<��"N���a�I�V;\qx��a�<A�A�y�0�Q ޲G�`���eT[�<Y@ޯ���ԏ�0�P��T�<�!�X�NQgi���5�S.y�<S�Yp�RD���M<j��Q�7�AI�<�Sj2���a�	6<5����dp�<)�܂o�@�(3.'{,re��h�<�Uܰc��h�ǉG }2)J��<	� I���z&͐�}��-9��Wz�<YRBŜ^e����mN���� �'�r�<�a�~rqsu/X�k1bшp�ID�<�fWKj�����$g���H@\�<���H�R� ��!Pi� R�<YUb��8,u�S�t�fX��d�<	�FD):�1S��� U����]�<� �"z9��)D�C��{aeTe�<9'��0��Dl�-T��x*6j���ybM��L��Xe8��DB�߂�y�/Յu���fB��Y	v%���_�ybL��=�d0�B]�|�����y���--]��HK@&����U)�y����C;L�y%F4�H�@"�4�y"ޕo0U�� ΟzU�����!�y�']�L�Ќ�tl0gAN!�y"�X�J�����
�����J��y
� |� �Ef�"�P�b� 3��* "O6���˒�)�f5c�����"O8���� %P�Qy���czn$�"O��P���I<4Ls��
|��(t"Ol����׆>�@vi�^z�UPc"O�IxQ��O<�;Fh�p��M�"O�C�i2z!	�]"c�:�7"O8���A�&^X+eœ�)}b�"O&�0��*�H�	�V�FW"O@�<��]1��w�T8A7"O����O�:�q����.C}R���"O���Vި�E�I߸I`r8ۀ"O�� !	��1�RU��MB�\e��P"O�ԫg�%3�]Ag핐1��
"OF��A��:8*	&&9(^�J�"O�;��@K�[i�NR"O����Ѫ65H����I�o�LlC&"OL��ꗍLZE�7c��;�`}QW"O.T;$��x���2��U4�zy)��'�Oڶ�/v�^�z������0f0O$!��ɾi���(ҲAF@��PCS�����ZV�	2]Fea�cL
��mr�%�zB�	�6����N�u�X�2ѫߨ2X�C�	�pҦ��ƠI�;�L��j Yz�B�	����%	�D�8�@�dN�B��}x�сn1`�Fl�sĄhxLB�	�_N�ВM�U�"<��� ߀˓�0?�3c�?N,��@�Q,: (���W�<q�* U�"1�H�	r�@�@FW�<����,]�6E[��=((�vM�T?a�����s6�4IO�; 4�0a��!�$�2u�rp��MZ#��A�+L�"=��9O��*%�`�螒p���AW"Oތ�6��<>5�D7q�"OT`�U��(9�J�f%6^��2��IB����^$WL�t�r"��P��ꃅ�!��ͯd5t��"�74g�����
o�!�dɆZ�U�VeM uYir���> !򄀵#i�!�5��.9t�@fm��!��(�d-
�kп)'���&m�!�dI�3��e[ԃ��)
��q�E^�y���Uf�����VM�i����1 �jpX�a���y����i$��!�H쀐P���'�OH-KhL���{�@�31��M�"O�(��8l��D�H������"O2e E�����86�_>L�nL	�2O��ԅ�I�Xt4�#!
	���N9pp�B�I;l�t-J�(�>�N	�Ŵ�XB�ɣ	�~T3"JxabT$2,V�1"�#D�Lk6K���5����8.�h�l D�x�7�ݕ16�kg�U!L�,r�,:�u؞h[��@�MrU�%�U$j��m��&,D���R�e_�-�#'���Y�0�<D�,3�Bŷ6��TIpn׼R���R��.D�,�� T�%_(u�c$��䊡17�-��`���<�Z�{�%ӄ� 4C�H�^��d�ȓ8n�q���BUJ �AD�h��]EyR�'qμ[7�V��0 �k��yPzڴ�hO�	,�Q�T��a�?l�De�
�[���/4f��LҎ?X4գ���m(FX�'���G���'>ơ�gm��m���ꝈG��F��S�W���t���ik'��5�V�hF{J?�k���	�,��iƝ|�`U�!��<Y���S���J�*[�6���PqE��;��B�)� V9�B��(. $I��V�@�
�"Ob����Ȝ{$T�)�
���"O����Ŭ`u���W$~�bSB"O�!���ɺfK4��C�K�n����'�qO,�e]�0&��#�	��&�&��s�؟�E�ī�'��iC���[Ѭ��t��*�y�.L��4�p�ץ$R��j4�O�y2���;����-�+�:#�hY'���ˮ̰>�"��b��ݑwB��Ju8<�r`jx���'h�{�Ӱb2��Kd�^�x��	�'�H�#���XD���%��p�9��'����M/%K:5�B��<c�~1��hO6-C�c�/|l�W�摩"O<�hOp�R5����J��[�"O. #�.H$���%$D	&"O.�i�*/�H�o
��"�IlX���O����W�0����"ٗt�#�O���T䖽!��Z�#R�0d���} �x��	�^��-"�Ԫ7��p#�[�>!����?�@R(�����Ĳ�C���06Z$�Oz�=�J��?-�
�Q���6nZN��n�F�<A�Ό�m�\1�Պ\5nf�Z�d�}�<�q����3����7��z�<�CZK�d�ңA��%+��EN�<9b!5n�"�
�CَV�mh$b�b�<�আ�X��!ԭ�]���a5�WG�<�@'L��rU���:��\��_�<qK�oY������i��mk ��}�<)��k���)�b܊Uj1� ��B�<�1M��BQ�B��	1č��FZ��p=qD�=׺D�3
Ős��ȢQ�0eV!�F7���mB�G�u:���
�!��1c� 5:5�S,!;�E�G/�,ax��	�h2��ץҵY��Z2���P�:b��F{J|�ν?�ܤSWnهl�Pa�E�F�<1cJ�-��s6�D�}�����~�<��(���JH�gz��Ô��Yc��K8�8�R@Y��(	z�ŏ?GԐ ʢ�9D�$����
�ȆD��G�x��BI6D�LBWJſY,�%��9+ )S��>D�8�<}��U��"�+D̀d�>D�@�1K�X���Aa����8D�Ȉ!���k��:�ȸ�7�5�$0�O�T�􎂉5����#�Q�5���� "O�E�e��7?p� 5e�5��"O1(w�H�U�\�J5,M7}�<9�"O ��)V�m[@,�^�r�ʒ"Oh(k�%�S/B�)�K4U���f��x1��)�'B$0t`��ע!��"-٨t���g<�/�6� ���'�bu�V"�V̓�y��$\��ēo1PyЕ��9alB0 Q�rj|i����?!�)��s0Ԉ0"�Y%6�P%��Q�'�ў�'t�����Qx�	zE��pS�a����t�&Ɖ+�n�Y��HB5���ȓ���D�ѣ_�⸃��Y�<��	|�#�Ű'��bR�ĈT��OET���OZ|8���/)�h�#�3��>q�����1Z��9:��M6^u��x�
"�y�F; ,�0 ��x3���y��P)w�Fom��x�`')Y!�yb�@�xp�dƂm�4}�V�C,���T���O��H#��%ոx�v��94�J��a,5�S��?a�$��%-n 	 ��O)�Z�,�S�<��iM�s��qY� �D�^���K�<� �x�G�M�.��sbJ�.��A�"O*� w �{YNu��I�&>`�q"O�\���ţhh.��EH��M"r�"OV$[J�<�^ q��c0<�YD"OPs���"��`X��5+��+b"O�P*�-T3'@��Y�C��h(�a�4"O��&I�B��ur��
�}�=��"O�hB��_�X�*�A@AX/Wq��i��'��ė�b�l�C��9�#� *���L}R��ӱ[5�R̚ '�V�
t�Ͷn_�"?!����u�����G^3h�,��A�>0!�º`\��1�R�½�rL�:8��A��(�ԁ��S�np�%+�H\�w�"1X�"O�Bv��P����D�+O��0ѱ�d"|O��j��x!���1'��JA��O�9c"�Ï]�����CC`�XW�F�<Y��O�Q5t}���0�<KTË~�<Q��#~�����	]�~5}�bT�<!g��##��1���G>5cXU����t�<Ya␺Ohr�V��[�&4�'��r�<��X�F&e�KB����Jp��p�<�BA	�V^��_2g�D�ŊZk�<�D�Z�o�n
����vo����Vd�<I�M��~��;��X	]֩ca�^k�<1FAFnƢ �`�Y�@�Ա�aHd�<��&E�Ĥa�I�`��؊ �`�<i<=&0�ʓ!Sc��Xq�MR�<q�8��	��_J��ɸ���D�<����K[��P$��� ��K@�<��͙�{D��eP�l�n��c�v�<�#��7h���1S��ZQ�8���t�<9хљ�@��Ь9A������(T�t��� 9&�8�	iW���v�8D���� �q.\�#��А[eBm{f�:D���p@�=t�A�pL:/�\e*E�4D��Kӭ��&|H�*���W�:y��$D�HP�ҧf=�	��c�y0"ё��?D���ɝ#�P["Y�]Y���J>D�sc�+H���Wf\)N�ؘ���;D��
7I��1�h�����C�4D�Xc3BÌ5�����J�aϬ���3D�̫��D2;�kU���\y�)0D�t���@;�tA�W�%A<7��V�<A�%�+�+��
����h��S�<�lF�4��E�d��#`7\l��Dz�<)��θV�\BVH9
�ԠPA�q�<�p��.E@=iD�51�Rб&�o�<!4섉� 婀"��R��ek�<�&�W.��=���� *(�&�RP�<Q��� H�D���H%H|�k���K�<����$Xv��:��>Dd��A	L�<�Q�!d�,��&->�̡��$�|�<�eˀ�RG`���ŕ�f�<Xr&�r�<Yժ^�e��l"���6\����j�<��A��F��ȣ���-!�4 �w��M���
�Wj�C'�$	�ո�I�#pmC2gԀ��8ǀ>D��AЉ�#�((WMS0��ҳ�=D���a�.��`,Q/_�ФP�9D��Q$�P#�X
S�B;~��(ӧ9D�|�צJ�	 Xp1��@�BЮ��Q))D�h���Ʊ`m2 �c#��y�nX8D��ufDyنp�J�b�R`)f�4D�� �(�4\���EDX�MFQ��!'D�P�����[l}���L�0m��d&D�� ^��LM$"�ƭS�EԦ���"Op%�w.U
@�H�X4Jj�$R"O|��ͺ"T`$���
�X�>���"O2�qu�Y�%P�8y3�/Q��l)5"O���I=�2����5w���b"O�)�cM�=^8D1���0s �ۤ"OnM� �ș.��鉡#S>z{�z�"O��`V؉ע�3�l��Q�L|�"O�5���>o��iY!�^��Ւ�"OДl_�jƊ�0郑��Ȑ"O�,§,�s���[��ܯ@��T�E"O��B�� ��ٸ���%RV^�W"O�4*0늎wa���+P~0]��"O  XR�	��:12kʃ6�8�"O<��an5�<�Ҵ�K�`L јt"O�����θV��hi���,2��=�s"Ot�i�N�Ze�C��/�
���"Ot�b�`�<|.�p��J���e+�"Oz�B�$ �naq7I�=/��t��"O�$j�!����g��Dn�Y�"OI�ӆ׵A��B� T
~N�]��"ON��HN=	�����X?�D��"O���qh�H�ܽig+K<`�P8� "O5!uX�Uw�RWcRi�,�c�"Oj���LJ4	I�%p7B�2sǶU`�"OZ��v֗gf��J@"֯+���f"O��«S�e>�{w��.�"<Yr"O�ĐS��~H��*�R�<��"OT�2��0o D�K:ln��7"O�X��"CڕIC�W$W<�T"O��y`��%:�p`PJ� �:�"O�ĺ .O�^Jt@S6dK���Q"O�T�ү^�Х��r�����
��yE1N,J�{�� wWt}��(�yr.��1���历>?�>�yЇ�	�ybb�w͂ec�AC%1���2�)��yR��1~�̜�ᓽB��s���y��H�$��g�<9��	�I�y2�I:0k�(ZJx���y����N���0!w���bFʳ�y���=JB����v����%�	�yҊH�}�K�:1�vms' Hv ن�}=\lx'В8��y��ɖV�"%�ȓ-x]s�BR�@�-o�g/�Ʉ�S?�=�eBւo�BPO�q,-�ȓ1�p+��V7Z4|�ڃ�� v�:����V�GQ�D�شj��9WΌ�ȓGKj�PGՐ,�$��AV�o�����O�̓WLY�i�2'���@X��ȓ%X���ԇX���a�ggA�k�`��ȓ@'t�Ȫd@"��%I)6u��/�A��)K6I���Ӊ�m��B/��kU�͠?��( �"L5���/�D��2Kc�'�K�:-Ɇ�<��58�ۀJ��� ��M~o͆ȓK���J�Y�}	&�x�L�����R��(���`��q��S `��M��@>8���ղ�X!��#O��܆ȓU����
F4d`:�U$�%�XA�ȓx��ʑ�ǣ�����据:����P�p��CY����� j��|��>��`j���;1��� ��Ʉ.��ȓ
aT����șh�={`S�C�8��mJ�=iC��p-��C�(%U����	=]In� 
�1��� t%���ĥ-�� aRz��!
7"O�!#�aK��8���P������б�����Y3p$�}��Ş�=�����ײa}�e�DI�q�<I�,�?+S��P�.��a,���K�2w̮��B�Kd��dO�]���?�'�8����ȜU�;D┾X=Ɛz�'��H���F�_ h�fR �(�I�J%�z\��A�(f.��Kʍ���UCd�lR�_*���@n�\2���Y  }���\�fy�� �R1�a��DΎB�B��xq��	Ҫ%ItH�F*�f�Op\����~!�G� y�$�����Ԣr���HV'T�6X4�чfu�<�C'�6����cG�h�y���=x&]S��I�8q� 0��u�����Ox5��BcOr��5���>]�EORl��؜rg��h���O�bTB4+ħ_���y���s���F$Ű<�� �9aP<�@�	���4JW�Kx�8�n���(r'�	�9�%yQ&X6]��*B�e^�5@��!��݊Z�OY�������
o|M�<�����jtY��b񀩒 �IU�M��5�LR���)C���^!!�I/uZD��@J�c�`G��`���r�5:�T�A��ƟT��<yҨ҇p�%Vm�m��n�}�<q���0T鲆$�g
�;���Gy�K��|=�ehPn�NX��1E#?�f�X��X&���`;�O��ǀ�eZ$*�fݫ,�����Y������e�"�Px�n �0a����`� �ES�H����I^u�` �_�'?����D�3> �z��Q�r5���	e+r\�՞|�o٦3�*axǁ�y�؀
�K���~BIC�9���=E�*�!mHZ�S�)~��3��C:�ēR�<��*�<Q����O� ��0�V݈�:d��KG(l�O��%hX)=�����*N4���"�
M��Y�����`(d�pjd*����O��"�E�W�b%~dVcGB��IQ�A �x2ş�V�F���$�����yp�1u��<q`o0_zX��P�(A��� ���?A��"I&&(���%A��d�!,OT�fo��M�P�&�X2��]��@��j�$���p���|�)����:��dZ��?}��i�NS���a�. |���ҡP�r���O�����P,r���t;2����:��+e��蠂KU�b�谨�m�:�]�z�2��F�@z�d��IzҚP C�ɪ�LTx�"����	�2���B!kDV)���)�S�^��#�->lJ��2��W+9�$�Ł{� ��A_hH<���+QML���¾X	�̒t+ ��?�DD<&�� O�K��d���TDT��PP��*�0�p�;�,#"^���˕��Ś�'�X��!���-`�{�A�"'�������RiB�rT�5T "tn�uK@j�iy����c����܌s,咕뜽N��+�)��'�p�%ʕ;�L���W�y�0$>�!�`�"�k�K�4=�����p0��Y�JD���)<O�}Ye��x�8�%ǁWU���0���V��Ep�6Ub H�O�qq�
��B甆>���"��K�7=ʹɲ+9N�Z��*-�y��S!����ɔIɐ�SBʒe U�ى�X��T�X< �8q��F@W-���I�x����rL��k����e
�q�r,�҅DJ؞H�s.��!Z�� !E����9��	�0ɖEؖd�ȔaXQO�"z┈3�����ɼD��5)����]��f�H�س=����'�~�pb�q4/�(j�
�C�"ΰwa��O?C�Q���jr틬wP���.�>���iZl��
�6@��J�(�HH;��ҽ_l��AS��D���E�q �����]�'{�ܜ��&h��`���� $�"�᲍�V�6��"OfP�ϟ)n�N��G	�<x�E)��E����̅�|�h��GY�A��n1������(΍9��#@"��~1��	"qB�W��+�=�'� ��	a��?h��P��Զrr�!0/�_��9!B�N�°aq�o�L�Q�'�<�1�?!�Ƒ�wA^��p�R�5h\s��;��E�rm,��v�֯C���ʅ��	�a}���7���Iw�帡H��-/e�ӣ#��ͩ1���t�r�ч?9lX9r*9�g?9RÃ�;p�0 �������m�'�`5�A�]�O�@�D�V�rlP�f���pB�'Ar0���(�mX��ώ&џ��g�<J~4�Ӆ�3 Nazc�p�$�۷�N����ħfB2��f�y�&�#G�d=�r��ECRQD��:q"d�	�h�Q"ц���d��#�61vh�'/<x��C�<��Ӵ� �H���FM>T'?I ��4O~N�z�2l�����=�On��g�:�?Q��3i$6L3a�9I�U��[ݟ8�f�%(�ご>E���²C.�dZq�Ig��`�0SўD���K�π i�!^�7� p�ҫK�z5t��>�V�h��$�~$��F/Đ5
*UQ5��'!���"a�� ���2��YUKϐ}!�$6O�r��&��"�@\{�AR&y!���Q�J}�e"��4�t�Ñ��8�!���IT��Cn ����D7h��'�������Λ/@�Iy�ǅeU�5P�E�i�!�d�(�R�8Y9Acj�,� �+2 ���L<��_�3 j��AnE�H*�$�4@RH<�g���w��c��V|��O�dR΄)W�1�OHd�����laT`���j�z��'�)�rH�s�I,G��\����a��X@�BB䉸(�j�R�lh.
�H�Y�N/4OZ�!n�2帧�OP�ESf�	|wjA�(��$�b�����3f"}2��^�%�v�RNG"U�@��X(¸'z��%�4�3��Õ<O��tψ�3H���B����]�B��+�{���I�3��L��e�(�LdRe/��(8�k+�����-$`Ê�x��� ?At�����P�{P^��W*�-9Ԅ�p�ÝL�a~��$u�,̃�蔚��@{�/�m�@r���yR'E?
��E�Țn�Bh!휣��O츸���8�(�n���J]�nQ��̂�$`��"O��E��9
�̬;5�9d@���v4O~��/��Ҹ����@�
\l6����S��=��"O��a6<����A^��	c��>$cC��=����6�0 ��J�A���ʸ�!���(zf�T#�f��d�R0K��!��@�&�~}i��rZV=9���z!�@!z��"��TM�����
m�!�d�$?t ����b7�3s�̆SV!�ę�L���H��0����Q�!�$̄8�|1�d�	h޴�a.xs!��D5���A"G�p��� ���}!��-�n�[VE
5	��$�v�!uj!�
�$?�T;�(�/���`�*>&!���[�:qX�DZ��2x"�o�>P�!򤐊pbx9aU.Z��h��I�C!�$���<h��H�2��=�ѤB	%�!�ă�k�ju�rS6&7T���cɋ �!�� ��'��O��"S��!�$��1z�+2%O6�"�bI�!򄁠NGzuq�g����$�á��x!��-Tz�blY�X��@��Ék�!�)�����4-ch����<�!��	ʕ��]*D�� ��.P�!�D�W�Q��$^�\Ԋ�r⯛&�!�$W�9�F5p��`,���/]8*�!�J	N���
̷�]��ɑ�I�!��J�c��`��`W+��D�j�����P�:��5 �+�@��������ȓf�f9�G��aZ�8�fl����a�ȓf���!�F���5�lj(�ȓb����Sc�4l��B�ό}%L��>�(2ϐ�m�����!����>\n�j���Ğ%�C�K��؆ȓaB���`^�Z���7��"q�4�ȓM�,�R�_�"�D���L2f���?:B�:��[�5DV���e�8KH��ȓ`Phe��"!(��]��'�A�~���TB�%��Ǜ� P�R2gM�����5K*��+�+S2�t�&��RP��ȓ^�9��AB�U�~��%��2�H��ȓy=ʴzEiM-/Y`�b��]�&D�ȓro���6��*��;A�D�k�J��S�? �Yp��`����7��,�����"On����
��Ĭ�����"O`ۃK�2E����$��H}x�p"OL�#��	*��I��-Z6d�[�"O�Q��N�j%䌜�r�P5"On�al���,k��`��D"O���A@�08,2�0�C<~vt*1"O^�ʆ���z,Y���!.�5�"OD��',�+sr�U�&d� φY�V"OL��5`�4l¸�ׁWWQ&U
�"O�l0���N*��)S
�)Q|v�
0"O�8!R��,F��q�S�"jh�{T"O	a��fƞ�1��4I䍠B"O���t�Ў}y��ٖ�2M�-�!"O�X��O~����a"�O+��V"O$���ѐn��d����i.�8:G"O�iPLR02pA#��� A. D�"OXݡ�j��3N��\r�(N״�y��˅l��X��`�6RFFU��k���ybI/$E�1��gݱZ����f�&�y.��}��c�%P"�j�$5�y"� �> �ePWfr �&m@��y���)�Fy��
�Vla����y���M��|`T,݉\7n���ˊ�y� ��6)~��5�Pi��y����yOJ�7C�H�gV�Q��Z��>�yrE�V��-"ՙ<+� ��yB&�=o CDnH�8��k�	[��y���v�jD�� �2�Z�aE��yBoN-��y�HZ˴�Y����y2��� ���j`��=Wa
�P��U9�y�C��-�H=���E���`R
���y�l�2:�9��+�j0Ȁ�m�/�y"A�<;�̀���u'�L�q��%�yr���B����ug��҅G1�y��{���Rj���:Ŭ��y�n�G�l�BFNƣo� h�u�O�y�
�d8���C��޽XrI���y"�%_*��fG��q�bM��yr!�7n��'��uȡ��H��y���tn{��ȜkdmHQo"�y�n�6=(`�S��ͣgiVٹ@"���y�(��I5�i�mܮkU��q� ��yR��m8T���ł4��2�(M �yr�w/�4�s��(�N��Ǥ��y�k� D�iv#�,uzV�3�Ǒ��y2�7/�B�8t�5H��Ձ�yR�;	�l%���X-=��q�q���y�lPF�1rT`_��,�+�M��y���1U.���ߕ���Ӵ�yRNO� ��d曋H<�H��c���y�-�=\��� Ix��q	�yMȥt̤��'��8W.���&�yB+�>O�l�d�4�<II"聁�y��Wg�\�*s+ϵ%�x��f�%�y�%V��]@���b|J�� �yBa��nOHL�1']�c������/�y�c�:`q
%O��!���Y�K �y��ý��bC`�Vu>$���ؘ�y��Dz9pC�Z��Ub ��!�y�DЖ���+��U���0�����y���88 A�ŬM����gU�y�I65-��,�����pw���y2 �Gx� �C�������L�y
� Z`���H��
������"O��G�4:�i��E�8y�Б��"O��Ð�VDp��KP�{7�i�C"O$e�e�ѣ~}&-��C�H�hД�'
`�@�@��#0!�J��񠂄��S��#�/��n�ډ��$0�IʐlZ�w����W�4&`�<��A>1.thR$�h��q�D͑ P[�ea�rҦH��"O�4⃇2M��(��NV*j5�V-��"9v��[N?Yq�7������b�&O�Te��[�ω|�B��4
���5��4_�����K�D��a�0�	_�*e�U�^�(�a{jB�h�R�I���f��5k��*��<Y���`���/�&�"<�v�>K����3�ϯc�̩a�O��y�i_?3F:�,	e�D��Ñ���d�l�CC����3DС"��V+C@ӾpN5;��/Dg�)�"OvD�рӎ"P�}cK�3Y���F� �xr�&2�@=��`ُ.���aO�� �ِ}!�$�v\&O��̅�{�2(p�O	���0���]�(`��� ��@*��]za�5�",OP�K�`�����䗼+�p����'���W�(�~��P��a�E:0��8���#	�iI�4FO�dH<IŃ�	a��3�F݈��M�3�Nɠ�EZV;���Ɗ�hⱟ0�@W'�	��)�Ul!V'u�"O�X�jĉfҨ4�TkU���]q�5@�L�8�K�M�\m��6Q>˓��� `�'UuT݂��N+��ȓQl⴫*Q3h�$$�a��$@,x�'ϨY�0,�Uh���ɦ�l�ã��9B]�W�׈6U~���W4Spq@j�%M���b�%2$���/I�HU��'l��Y�%�(�a���J%�������16��0 0�/��;k9 �P�F6q��!�G��:B�I9=jh9�`d�S��tQ�O|F6�I"a7��ӸF��� eʃH
M{�
�f�,B�	%H���1hD�*'�ƣG�c4؜�΂�0=A�,�$����uL �8DN>�O�08$���G���Wg�k��h��kҾD ��X���xb&4�I��]�C9t�*A	�hO���B�Hc^h`��4lF�B;Pa�R��U@@B��y¤�7+����̙1��݋#�?a�BX�Dش!�=}���+Y/�X���ō*�Τ�����BC�	�I�\�E���ʴ��CYD�r7z ��F������A�&PB"㎧p"Ҩ��,տ>����dW3V������ 
q^�+��P�d�H%�"�Q J��4�@�%$����Ȓ�/t|�ZA�F�M,��˃&5ʓ=l^��g��*|p�J��l���<2�%������J���y�"%X��xR��ѐi�+�	�%)�-fuy��N�i��)�� $��Z*\����=:"���+D�x�O��g���DQ�9�ڵ
��4#��D�!�����0<O��W)"h�`�F%5�b� ��'��<�A�ݙx��]����a\إׂ_А��\N�<�V�R�=<��ÈA�~�"�FK�'b����Ӽ94�F���>^��4�VP �x��&�yr.��q�x{�f��2�v`�(�S�@3�NJ6$h��!K�"~��
6P�|Z�C�����!D
�d9C�Ig���y�ڵS�D݃Wf,�P��{��;$���I�b�����L�V����&�����&����4B��l�3!ݮΦ	�D�[: P���ȓ�2{���!�%)�ąSqj�C�i���S:�E %��,9P��;$�:D��#�OX�#(U��,1��T�0�=D�h@J��G0�Y@�C�AqF��� ;D��*`��;Հh`��hY|]H�,;D�H�eV)e�\S�۔"Yp��,D�@�c��^�(1���s> P�E�'D��A`�G���o���M���&D� T�B>����8mb��ؤ�'D��J5�A7kT�CĸK�����o%D�� .@@Ku��% K'����"O60�̜�zȎ��B1d�����"O\ 0�C� 1��s�#�%Ir����"OX
E@I�e˘U"�ūk҈��"O�8A��R.h�����䁙nI�3a"ODL���L�~j�ղ��� ����"O��A뒭U�̘b��3����"O^��c�2q�B�+uA:h>䴒�"O���e��7���@�GG�m"��Y�"Oq��̾�Dp�&�Sh�ʰ"O*(� ��
R�L(�Cf܊.Ph�g"Ov��W��8��ĸd&J0!�<h��"O��
 �=�8Q�'�*�uS�"O���!��5O�����X@�"OF좒�F�e��z#MC�"�TX�1"O^%Bϓ1�4�k4��iI�=��"O!�C(�y��8�#'2U��"OP|�4L΂g�V !7*̵i.���W"O�ͣ���2�v�c�Iņ'�hk�"O��Y(Ԋ+�*M�����w��Ճ�"O���@ٷF����Ў£l���O�<��H;O&�JF�65�6����J�<�BڈZ��=)dO ���eB�<��m�0����������(�g�<a�i�,� A��6��� !
U�<�Q-�0�L���9Y�ՂAEi�<���H<^ $�dL�=�j��Veh�<	���;A�h��m�9A)�P���h�<�S�$8�@PQ��LC�r%�c�<��kH�T4��<"J`R��Wq�<i���=(�*�� �,���W[�<9��āS~�dsE�	�_X ��e�|�<�W�H���Aō	�bAJ���~�<��ꃓS�#Ɵ�݂i�qh�\�<ɔ�x����ŞN�F	�2�Y�<aţ��,���FeC"-�\͹IR�<��ct�h�p�� �n�!f��S�<1f��y�P��6W�5kaO�u�<���ȸl����LZ9����Zs�<Irψ*�4���8]2,;��K�<� �ۏ�F�b��A�����G]@�<y���XA $#'d�t���`�!ZH�<2'�Mfv3 �����b
G�<9���~&Ƭx�@ĚKe�Y!�O�|�<i׫R;{h��r��E$|E�el�r�<!6!�b�p�q�%J���8r	@j�<�4+�>B:���c/juX�kGb�<�W&6,$64�jR$��1����Z�<�aß�LtS2)P4�\����DC䉺S�Z�	�/��r�S, ~C�)v��t���H
u��p�g�Թ1�JC�Ɉ)+�!�+ݚ*z�C�k�+{t:C�	�lk� 3�6�Z0A��ØE�B��)^J ���u�Ɯ��@_;E�(B�I�oڜ��4�Q�kY�t8$� �+�C䉩?ؐ Q��?�I#*ҫ19�B�ɟoI\��g�3d��҆Aл!6pB�I�[�D�D @Z�&�{�&57�VB�	PL~���:n�Q�]�,B�	�u�Y��J�&�,LqB���C�	�>.�Q'U�Y"ɰu)¾J�C�Ƀ&蘴P��*������"T
�C�I��ek��A�S����tk
�k�����B```���6vӔLPe̌ZN�+�K҂= �[R�Ϲ!�!�� ��Q	ʝ��=i�̄5+�:Q""OX�Y���E�������g��Y��"O�Hq��Φ]L�H9��њ*���b�"O��(��ɜ@����͵(d�M 6"O2���+*��hH�ATvh�E"O���qZ('����fH2{7n%�"O�b��G1D��LhƌE/L���"O ��!�K�/�2iX�*�%x��iU"O�@E��iV�ǉT>[hU��"O6I��v�~�Е(��pO���"O(���NO��(�Th��D��"O�����K�xfSGG�q˞�!B"ODX�`��� &Y�v��q`5�'��0pn��eL�R�*E��,;���F� r�Ì�x��i�Ɩ�b�4��g�O z^w���
B�iΙ)�*}CB�L�vf9�ǉ�b�䘑2���$���d����5/�p��F85�tԠ��Q�W��]���>�QaU#d�P��I��f�x�b0u?�y�7*B�X��'�|��2O~�"�}��b�bLQ�CA�u��РCCP�'H8�)�b�N�S�O�`�X�nD1�h�{�����+�O������![�1��K v&�Zbɖ�ѲC䉃D�z�a'�#���B�.'��C�I�AX��A�˕)T��ys�IG�Y!TC�ɎY�$�Rb�_8�$Bse_8�"C䉬5�0���	�7E�L�u�҅|�B�	'%:Թ�7MF�!��H�є��B�24�:��2��A��x���,��B䉘�3��ÖTz���<YU^C䉡6��`�cM�*	������
�HC�	�y�`4JTȈ5ch�s�G}�C�	29��I�ǂT������fM
�C�I������ �:�\����*B^�C䉿GS|���L��ߊ�M(nC�8d� ���K�V�8!��ڞB�I�d����%�%t,�q�6;�C�l�D��"��U��a�䊙@y�C�ɩ~f�����7��Q�h�8\��C�I:S$|�e�s8tyz��ǘC�ɕY2�S��
�
�p����!�fC�	[�޸�,k�,��h i`4C�0m2���w�X�82�`?C�	�{�^X��낁	E�0-�7i�B�ɂP��Ŋn���I,"��B�&QP�i�O�#�T����
I'B�	�t�Xǆ��;�4lZ�oZ')C�ɤ:(���wA�Lf(�R��=@.�B�	� P���aD$,\2¦�50�B�I}���iBgҷ�!JfB�	�"���F�4m%��o@b�C�	%<|�1ua��P��гF��+�
C�Ʉ~f� ���[�d��Qa��\i�B�ə"���Qō�F��T�K�;@�B�<g<\bU���d=3�����B�I%bѤ����I�i�be���-4��B�	�z��t����b�:�I�I�i�^B�	*`t�P�S��&q�Q	C�Q,�C�ɜ	�~�xP��7i*J�A�^C䉏	"�� ���cT��U"C��"M��L����-����d��;;C�	;u{��фF0'b�����Z�C�I#�t��p�ۜ2X�X��N�5
�B��;q��u:U'�>^�NA@���:%�NB�!>�@�����@8���"nT��ZB�Ir��1�"׬_0�` �Jթya�C�)� ���PSJb�c�4��A"OT�i��l������L/ d��"O$Xc�[(2(H��K�u����"O���d .TǪճ�E!vH���"O�)[W��o���A��'
=:E�2"O|�j�&^.;��u30�e$�e�"O �NI!��r n�:E#�1{�"Oҍ�PÂ,'�B��}ȨaG"O4]9��$���#�L-���"O�\��[�D��,�/s��<��"Ol�a�K����(X�r������yBg�]D88�
J4���$-۠�yҡ͚"W��;�OB�7~�q�y�aGj��.��5���y2x�LA�H�X��T���yB&��� 4��A)��o!��	$@hЬ�Z'��;�� MV!�d�%-ΐ���X��Q��}�!� pGr� `��9n�
H1�DT�7!�S�S��Q�M�ʭJ�nF/QD!��΂Jq*�P�i�q{�!�.ZhU!�$<DBTT�pl�,J�n�bE�^.!��A5AҖ�k��N�X��-*�!��h!��K�P��q棎�V�"]: �/!���H��i�c�:h��RL�}�!�X	C �@�*^�px9�iݷ@[!�D�gcH4��FN,�%��)N!��
X��U�_*d_�h�ta�.�!�D�!�~����ͅi}�uI6� C1!��ǘ�
��f�P b}��X� ɗ/"!�2jShq�'ӓ	h��+��2I!��\'U��4�S�z��Q�τKf!��@�}C~���Ú��.�BC.��0A!�R��n�p !�?�D��f�-Q?!򄖟W��0��o'�*Pc�)��S�!򄁞?��p2�a�<�� �O�!�D�:����5E���"�S��Ww!�	%� ��H�Y�Fi�#�x�!�DیB�F�����W�X�7LCaS!�Jh���B�� Z��!���>8!�D��nŖ�3A�mb\!H�y$!�d
�7��5��#YcT~����@!�
�S� �Ж ��X�<���E�d!�4T��$3B��#��
E\/c�!��[ U����CN!L����Q6�!�dŖO� �S�ݲO⎤ �Ϋ�!�$�$l�P�����
pnh �̆�!��h�
E�����h���UIQ;t�!���{���1���g.ҙ��A�`!��̌3Z�|��B7�D���a�&G!�ȔM-�eGτRvh�<!��P�Zx� AABϮM7���P��.;!�$6_CF="�%b��P�4&!�M�Ԅ
�nJ$K���3�KV�vb!�ټbL%���[�|���*i !�Dk�V�<b��0 j���!�d�#C�T�%W	���si�$}!�׋v�h(�Q�ϼ}�����!��Z.�� ���_�᪔%��e�!�䇳0
��h�k�7y�S�bU�NS!򄞎l�y2gb
2Ba:�AQ� ���dQ1��c�lط09`��PBۻ�y�I
m�$�9�G�/����l\��yR˃6"���d�0�ցK&DK!�y
� �؃D`ٗo��� �ć�2�<XRv"O���$jIg��	��F>\��f"O�`�J�a"lx���9;ԅ4"OP��+*B�j��(��AT���"O$�f޻P64<;�G�jBXia�"O��!���8v�9���м%Anx��"O"�r/!@ X�-53F���"O�)R-�W���b޸X�bi4"O�y��9�(����^MR�A�"O:��g�y?� ���K�!J
���"O�) P,έR�D����8l�
�"O�s��ۼVR`���E/>D��"O�+����"�V���O-�nyi�"O2�D��65_�9��ӹb�Ą�U"O�X��Ė0|����A��q��"O�����(W�L�K��M6 ��Y�"O��r�勲";�q�\64�|k�"Oؙ@�hZ"W���cP�"h��E�"O����Ԃfs~e�$&\�{g~�a�"O^��b��?{�ziS兗:H��˗"O���g�^�e���p ��*��w"O.���!�<���#4,��m �ab"O�Aװ�ȑ�0ʫ[^�xe"Ob��ΐ `��Zg�B/+��p�"O��`��Fo���(�,)h�sU"OV��ŀ	R�$�c�3<XX��"O�q8G�F�7��1��G	H��"O��#r�E�1�N�A����]�d"O�0�l͎^Zh��!�ѤR۾|a�"O*!�!,�6O=������L۸m��"O<H�% � D�H��Γ�
ìhsC"Ofŉ5�M�I���m�2|�:��""Or��5�2&�m�@-B��-�"O|D*F�C9^&Q���Z�~��e"O�5Y��ɉ>�XPS�+ר@W���V"O�\����3�l��e
�$g@�i 2"O���V�®:�D�3�ȇ�i����"O�y�%G�#|ea&mN��� c"O�Yc)W�j)	E� %a�&�)�"O�(Y��?��9 u�����,��"OX!�U�2w��H��V
^fB!��1ik��̀�wJ6Mcߢ�!�D�%{�JQs�%��B�@�T"C�A�!�$U+�8��4n�q��D�O�L�!��0_CȄQ�ȘF�������%�!�D��|8 �*E��JEҒ̆��!�dM {=<Ó�>Tmn�3*��8�!򄍇,���ÂE��,��*3gUJ!��E�"`ak�h�30�x��@�0d�!���>}����دa�N���	�z!�dߴwĔ��S�w��0!B�ja!�*	~$M�#�ۡ��;�*W!�$�P(cE��eѬ5��I�6J!�$�;C�.U�5���d� !4bR�#�!����+��ř8�!؃�߃a�!�4��t�EN���|b��۬,�!��F���I���p��UqO� c�!�^w����t�\	2H��R�R t!��Z;\�� G' N^�`@�V�<;!��&nڐ��ڷy\:a�"��-!��=Ғd��G��M������?'!�$@�Su� K3�Q56hV��r�K5�!�ÏA1�ܺp��%G��u�+-7!�L�X���1!AP<R�r��G�Rg�!�� ��I@"ٜcLxA�D�?�պ�"O��3c��^4�ū"A>:�PȀ"Or�I#���T������^�)�p"O���B��9&"���ӎ:j%��"O�tVG�S,�9��/��H� "OH��f Y�j|"�Q�)I41��a"O �.�wƴzv��^���"O�p�3��7!STE��31d���"O�ͣe.&�zp�S� :�!"OF��7$��i�Ⱥ�M��B�8x�"O>��v�Bt��p��.�,�%"O��G��#/R&�S#�W�ƸX�"O8x:3#��8$�H���<a��,��"O��X�!˽#s|4��׿xR,��"O��ѡFJԑ�"C�1����G"Oz0�D�)r3�@3���X��|��"O�A��+�b���)�>5q��""O�[An߀�
��Ǜi�b�"O�}�G�[�G��|�. 9�r���"O�8Xwϑ�_<P�s�G�ʂ�
�"Op�"4iI �4u"U��v��c�"Ot�#��N�=QL�k�	��H%C&"Op�p� �,����gS�;J��#%"Ox��Tl�a��}�Q,-VӦ��"O�\���W�-B�k�>�6Ix "OH���B��R+���lP�\�2�Б"O� 3�֥^���vK� ���"OP݃ad�z�q���۫o�$��"O��a�   ��     G  �  �  �)  )5  t@  �K  �V  #b  Tm  �x  ��  p�  �  �  x�  �  ^�  �  )�  l�  ��  �  ��  ��  \�  ��  �  l�  ��  M � � p V �% z- �6 �= WD �M U �[ :b xh xj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>�z���瘝 C��rs��i�99�E��^� �O��oW��|��?�Q�952�b��d̔��&*�?1��MO��y�4��Dm>�������sXT�0�
L�VeF�˂�̕(�c����Uy��S�:��MB��v]G�\f�[ش0�M�<����Kw���?�m3Q�D��	��F!�X�$�Of�	`}��ʀ,r�F<O��(�_�S��kejC3&�	Ie5O��I:�?	a�;��|R�-�`�P��O�]F!: �y�,͓��� �$�զmp-1扉��Zj�{3. ��.H62uj��?aV��	�t�S�Fٴ(��A
���N4���������O\q���%9�1�\u���9����̨aSJy��[k��(ɵ��=v�ʓ���O?牟uhq�:)�J�ƥ�m8�扉�MC��i~R(d�N���,غ�$?Z~e��'ש/d>���H�	���QiT٦�'��K�?��@�V8]�|��F��mK^�SE·@%�'O�i>M��������$��7"�0������={4,�>Y�\�'r46�=G�����O\�D)���OP,s4�5ز�r���1���vdZr}��'B�|���� >-��N	(p����ÞE9���V�S0������^H���e�ړOZ�Z1�|�d�$����@�B|B�S��?���?y��|z,Of�oڑjv���I�.��6�$;ް�������x����M�J�>Y��?9�=?��+Ӭ ���p���Za�穈)�Mk�O˄����z����wYNcC꛳�p�ͥ6I de���I���I�0����
��7!%�0V�D�7	��?����?���i�H��ȟ��n�e�ɘUl���h���Z	���S�4�%����ß�(P`Ymn~"f�[���Ca�h���z�ֶ�N�ȐJI~?	N>A-O�I�O��D�O��ɖ�C"�,e3r���a��م��O���<a7�i4�aC�'���'��ӟY ��`��jx�q��߼^���z���̟��IN�)*f��_1��!�	/A��5x�[�3a�	�dd��:B��R.O��?q�j0�d͹Z�����Ǌ3�HLږ�ޅG*��$�O�$�O����<���i�+��|u��&�)��j�����������ڴ��'P���?ѢGG�e�v�����
!;�%E�?��m��5Pڴ��D��J$`�c��d�A�v8��;>I��4����y�Z� �	���I�����0�O2|�`���,��
G�)��	��d�LE����OV���Ot��T�$�����%n���: d~pٱ�T�,�*]�I���'�b>5qu�צ�MČ��L��tJf�8g�Ȼ[��͓
�d�۷��O���M>�/O���O���f�d�U$Y<�TQ�Y��<��ʟ���FyR|�t\��"�O<�D�O�Pz冁=i��M	f�1F
�h��J(�	&����Of�XBt�џ|yɵJE�dj���	6?�����.�T�#gS)��',���S��?a�/�;rڭ��#� =�@�vo'�?���?���?Q��	�O���1oni��(Ͷ`y4�{�A�O(�o�3Q�������4���y�g8wY���(G;���u�̗�y��'��'���ـ�i���"l�~�1�՟��w!�$T4,1�wU�+����!�d�<�'�?1��?����?��@�wJ��Ĉr2Y2�A�*���٦��$�����������gKCr�ZA����!ud�9"�&�����柨��Q�)�S�7H��f�Z#O3$@��BГg	2�ߦ	+.O�<Knֹ�~|R[��H$��	���X�`�<3@H�#��ş,�	؟X�����@y�NiӖAS��ODu��j̀)�h1�ţ	�Q}$qa�*�O6lZo�0�I�H�'�`ÈݾT<�pP�A�%iL�ժd!J)	ߛƛ�4�6�R e��/]�S��� �ez"fB�.���A]!;��+G9O$���O��D�O��d�O��?YȔkĘ�hǯS����R��ğ���ȟ���44^R%Χ�?���i��'�����J� $I�(t<���y"�'��I�F]0@mZd~�+�������H[,yb�O�`����ʟ�$�|R[�L�I���I�(Jde��2a�@�tÆ�;�ִ�ů[���	Qyrmr�j�� ��O��D�O�˧9�D����j�� �L~\���'.��?����S��DȜQ�,c3AͤK� ��EɁnK��Տ�5F�d�O�i]��?�$�0�Dψqԥ�+�����o�=gq��$�O:���O ���<�iz�JP!½!Fl)�w�;e��u�!��:r�' J6M;�ɶ��D�O�)0r����aQ�-l X9����O��DP��F6�&?��F�kGP�I:�dlL�|e�TK�v�bP�`,�yrV�`�I埘�	͟���⟘�O��$k��H]D��!c׳1��tk���ɫ<�����'�?	A��y�e\=2e�;�:����!�Џ9R�'�ɧ�O����R�if�� >��rEd��G�H��w ��]��DZ(MD��[�� �O���|��#���� �ʃLV��+�%N>��!A��?����?y(O��o�0w�1�	��ɨMY��(ٛyІ� �m^8cn��?�@\�X��˟�$�D(a���w5h�ħ��j��u'5?�gIJ�%���4ޘOHD��?��B���y"�&=w�萇�,�?I��?���?�����O|�SiE������/}U�e ��O0$mZ2���'��6-"�i�!��C�2!��m�ì*������f����~yB�Q������I�(��C�T%Fd�����]>�0�
E ��U'�4�'���'���'�'S������}$��.�R��T��ٴA�r�����?���'�?��j
24A������;o"�:�#����؟\�IY�)�Ӎu>�9��A$x�A(q�8xFE�2��3G4��'��E,ݟ4�@�|R\����F
	Ab�iTI�AF-X��]ݟ���ğ���֟�Lyr�u�vɨҮ�O���¦�P��L��&y�ҙ�S��OTdm\��h[�IΟ��	�����D�~�+2�M�%U�T	���.SR�\�+���RE���>��*ix����Ҝ]}�<S�%�.F�F��t���P�I��p��K�'s:h=�7�7y���.[-<����?��Hƛ� ɔC��I�M�L>)�BD�C�eK��U?h?�xRa�T��?Q)O6@s�r���+(��C�:]�����Vz6*XZU!��<F���@��䓾���O����O���"cfm �N\v'�𑑥Iw�b��O�˓;Y��!ޢ�R�'W�T>)�W�3e�Ĺ;��<; xH��� ?�PZ������ '��'Q���0��^���3HĿ9���eJ�;�f��˝j~�O(��	9Ua�'c��f�L(s�`���K>��V�'w�'���O��I��M;�o�`S6�a1��<k�.$�����[��u���?	��i�O���'�OP�^�>�����( Y�P(�!W^��'�LS`�i����~m�S�O\�:����E�E,� �f!=JCv	����O��$�O����O2��|R��_&&n���+�(oS��Sq�I
H���eC2w\��'!2���'�j7=�f��t"D!Ml�=c�����%s�a�O�b>�2���=�mDT�uM�w�ڑ���[�zA�1Ox]#@�\.�?�n:���<���?����%�=p�
A�K! )+Pf��?����?i����$A¦�Q2��@��ҟ����8�J�QQ�I�JD��(�"AK�g������h�eW���IŹ%�
��1IS��sK�$	��0�M�&��DKw?���:�I��#�;z���` * ��r��?y���?����h����7(�<`�2
�� (zѲ&�IJ�d�Q�$E�D�ɔ�M#��w'��C�*��]K7�̢u�X�+�'�B�'��)��]F�v���]�u�\��3)( 2�ƹd�%q&�[�5��Q���|rU�,��ϟ��	ğ$�	ßD@�Λ� Y�� E�3VDz����Qy"q�Q���O��$�O^����ɫ�����@�gO�ѡ4׽. f��'G��'�ɧ�OM:e8v�^ M��tX��0��pß�k%����X����q�D?��<q&J�u�N�+�K�"z��=��G��?���?���?�'��DQ�Y3�����q is"��E lA�!D�| 4������C}B�'YB�'��, A	M�@���"Ք���(����f���g��,%�4�	��R�e��,��%���Un��LI�6O,���Ot�D�Oz���O��?�Q�F�	�J����#�v�e@�ڟ�������4�&��'�?��i��'b��y���}����װ	����y��'�	�^�t�n�c~2���z]b�e�d3�U+_�)���Xh�~I�I�dz�'���ޟ���ȟ|��N:0{@BȌ-��� +�=7�M���x�'a�6m� �$�Ol���|"V&N�[�n��d*�4o��5KV~���>��?�M>�OxJ�(�*�����O/W�:B���!\��i����|�a`��l$��Aa��s���
,�ld�%%�͟��IП����b>��'M6��7S������Q�0EWS��\9uͽ<1`�i��O�Q�'�� �I���8�͔28f�Yg��G�b�'�҄��i��iݱ9��T�?�Y�W�� r�����=n2�q�E��rޞP(t7Ojʓ�?����?)��?Y����iC�^�����,�{FrEr�ߒuBtm��U�	����G���H����`&�=CDV(m��g��?����Ş��Y��4�yB�A�>#���Wd�)�j����T�yb��|U�a�	�xD�'Q�Iџl�IU���Z�$ɌD��/� S�,�	�����ǟ�'��7M�BG8��O�d�Wtڀ ��%<ޝ��lY�h( ���O�$�O֓O�Hsg�̡��E12	�S�,�瑟�ba:0��LXo!擿0��oAП|P�B�/�t "�iP>�l���ß������	PE���'����f'�#k� ���c�HȠ%�'M
7͚
1^~���O�oS�Ӽ3��$��h0�K[҉�����<I���?���J5�u{�4���Ӗn"�d���S��%�ִdI�8��,��o�`��,��<ͧ�?q��?	��?م��� Ƃ����g��5L@5��D���Ґ���	ӟ�����%�@����qc|�0N
6|��ǟ�	y�)�*�<  +�/�(Њe����Pyq�K����ٗ'dN�Cń���"��|�T�x�F�J�&��a�2,б���C �U䟔��ϟ �I���S@y"�b��)�J�O�d9$e^�z@�yzV^({[e��7O�o�w�|��	ğ��'sd�BC� �.�yF&,d����і8��v�����R��TH y����mۄn̻-l�;��_?8
���bp������Iğ0�������2K��ݢ0A���/q�KZ#�i�	˟�	5�Mk@��|j��9ț��|RG\�(	}i�< �����l�Vq�'L���4�����V����&J:mB���P��0�L�C�eԊa&(��v�'�
'������'v��'�R�ӣ�=��5��Q�q d�'��\��:�4I���I/O����|2ワ$.J0���T��j� ^~��>i������F��|���|�2�I��V�h��@uҦ���ƾ<�'���������zhP6o�=y�R��#'�2ߤX���?1���?��S�'����H$�O�2��]!�R��1p̕���D�	՟�s�4��'X��?��@�UV�����#V���Ղ�?I�e�R��4����T��K���/O�m)q�͏�hJw �k8�T�#9O�ʓ�?���?����?�����O>�\�8C�� CU$��C��m��\f
h�	ş��	]�Sşd0�����,V�̼��V)������Ζ��?�����Ş)�"�ڴ�y����Y�I�r�c�ݣ��]
�y �.�$U�I?��'���퟼�I�pDXxPFg�(Į��I_3�Q��֟��Iџ|�'a�7-�ր��O0��ŰX�� "&G��P�،W�-&�\�쨭O �D�OܒO=ke�0fpQ�Ѩ��e�ЪR���ԧQ4f�Vl,��'`�l���<����.bv��I��$:N&����R��<��۟���̟�G���'f���ҍW�:���E0���C��'�p7MW�|;���O:�oZm�Ӽs@�Y$I��;c#ڿ2XrxɇD�<����?i�����4����^�%��O���AVE,��*����![<(�ӛ|�P��ٟ���ϟ�I��+�'�L�L��%x�=��b�jy�f��$m�OZ�d�O���\��ތt�v��6`H�-��D�%�4cW��'���)�>�zDsW`�ek�|8#��p�l�i5�I�uV˓d^�����O�AO>�)Ox�xQ��)x�z)Kg@b8�}9GC�O����OZ�$�O�I�<��i�~q���'
d��O�_�d�8V#ʠq0���'�6�<��9����O"�$�Oά3�C �L$؃F����3��@q�6� ?qc��9�D��V��߭���&RZ�C�%ߟB�|��4�u�h�I��I����I����#BǎV����@�˽R��1$ߪ�?A��?���ikD	S�O�r�j�>�O��w&S�>W�aa�Ɔ(^�rD) ���O^�4��a��o���el���B]&/�T�H�/�8�:�0ӥ\"3/��	X�	Xy�'K��'Z�'K�q�Q!t+�8+PJt��Q :#b�'��ɪ�M�ׂ�8��d�O&�'���)U_���	��X@��'�2��?��ʟu����n4����	#X��(��Q�+{�}Hq��* ��|�ׁ�O`�HJ>�t�K�{��ːg������?a���?���?�|2+OR-mZ��`!8��#Dt�Ŧ5UhdQ2*�4��
�M��ͪ>��NR⊙�'�<��3Ӟ�P`����?I�b�=�Ms�O���nK���L?�HB"B�'�^�2�V=aȌ�"�l��'���'{�'&��'�哜3~�9��!�8��aB�I�D�� Y�4S�����?������<Q���yW�^�
3�%� �N�k@���w2��)A)��7M��ɥ���!	���-Y	/Ű���#{����3
�[_�	sy��'E�FO�,+��6�ψ]��Q6�N�8>"�'�R�'Q�	��M�W��.�?���?af�W'�֬�4& �A|�i����'#���?�����za6E��H@&ڊ	ѦD0x($�'+��Ԅ�;�x���D�џP�R�',5�TI��@��U��Ȯ0������'���'B�'�>��$XL�RoРʀY�F,]+]�@�	��M��K0�?q�x4���4�x�P��C�R��6���W���>O|�$�<Q"��Mc�O(����Й�z�� tqh�
� }��#b웋�l�9um>�$�<���?Y���?���?)2�	/͈	��Ƙ1O��7`���d���]�1��}yR�'b�OfR�ƎMAdTS�"֩:�Z�"��0H~j��?����DC�xY�%�%�C�8�6���;�(�94B�P:��$�@8���'	B�%�4�'-�
ƨ��jƁ!돴y�P��'���'�����T\���4u��LB��`=��`�#�h T)��)=��̓}<����O}��'22�'��yB�ה"E�Tї!͡�����������R2�¶w��!�I������@��b����+��<.n<�R3O����Ol�D�O~���ON�?3'��8�0���7.�f:�N��I����۴b?\m̧�?)0�i��'2Jt2A��id�̸ �Z7ze.a��|�'%�O�n�ʇ�i�Ɍ�L �dL�{>�b C�I��9�u��L��0��<�'�?	��?1 g6\&�Mq�mJN�����_��?I����DĦŠ�![cy��'W�*xr�A�Ⴡ.R��[`�%IPX� �	ş���d�)rE'���('	(�9c-VtFX�"��L�� +O�	8�?A#%������A��	�dL���4H�d�Od��O���)�<�d�ixV�f�"jA�%�K�F��-	Í�l"��'��6�:������O���KՎ
X�P!JU�rj��:��OP���<|��7�/?��'X�X)��wj*˓)%`SF�]�� po�	�M����O��d�OJ�D�O����|�W��o^����1�"�ض��b���lŞ|�b�'�b��t�' �6=��\���G�z���6 �h<�(���O|�b>%�DEئy�_���9`f�l(�#����0�f�0��&�O��J>�(O����O�@A/ j��,I��/*��д�Ot���OX���<��i���z��'���'��q�@F4��x*��� 
�,!��$�S}�'��|b��\�XT�g 
h��LJ�`ĉ���@.�b���oш\1�t����\����%l� ���Y�N�XDГ��70�����O���O��:���b��	V\Y�H��P�(����?)P�'�^����?1��i�O�.�6���&g��p�DJ9���Or�D�O�]�mӨ�4� 1Bn����l�v&Q��E�B�����%H�����4�����OH���O��D�c�6�yC&51��E[��]!P.˓	���g?�"�'����'+H�jү��t���5'رz� �ʹ>����?�K>�|�T)�
{�Z1��+Z53������n4p���Tf~���j��I�L�'�剆@�6)¥��;��iF���:pJ!���L�	̟��i>y�'
�7-��8�<������������"�/�`0�$�a�?QbX���I����I'`°!rCI�,�SU/ʍC�Px[@#�¦��'5�B�HX�?�E����w����gF��\���ȃ�(�H�`�'x��'���'���'��1�.\%���k�����&9�?���?���i&�Y+�O��Kw�$�OfP#ʘ+]�fHX�lĎk�Z�hcm7�d�O��ԟ�@"u�i���� ^D]kg�؀t�@�sRl��=Tl2$F7vR��~�	vy�Ox��'���Աٖ�jb*�F�ԑ��2�'���"�M�M��?���?�-���3�N)��y ���u iS矟x�O`���O�O�SKz"��Ҡ�5���ԁ�0T�M��"%�:��*?ͧJ����E�\��h�\餽�@X����s��?����?y�Ş��$��?�(boJ��Bԑ$�Ӭ���h��� }�F�d�_}�'�,�A���e�]� M�[�����T��r�mզ��'�TQ��?��^�XȤIK���H4ꂬQ!�h1�w���'��']r�'p2�'k�S0qh��\ vl����Ss_��޴"yV�+���?����O��7=�b�s����|Ԭ�[& W�h�J4Ѧ+�OX�b>%�g��覽�?��02#HI�
�K�$ޡ0�θΓ3�����@�O�BI>�)OR�$�O@��pF-]&9ۇOۭq�0s�/�OJ�D�O����<���i�v�ɗ�'Y��'����lϯ3r������1���"���HV}��'��O��	���G<��C6e�H6�h���@��oJ;d������k��8e������
�E
c�at��yW�La��U�h�	ӟp��ݟ�G�T�'���'��6EhaCu��:�D���'H7�O�J���D�Oؕm�P�Ӽ��Dޏ|�B�ʠ\'*Z��O�<����?���HΙ��4��DJ�~,T�{�'|?�A���04p����bTe9��<�'�?Y���?)���?���/'�����-UW����������,A`r�'B2�)6$��T��L�$O��r�.F�BA�h�'���'5ɧ�O8H�sՃ#�U25���(�v����(ؙ�O��V���?�3E �d�<9%с>�"�j�)8L!; kG�?���?���?�'��d̦)[f�C��h�aE��j9b4c�1u��E�o�Ɵ�ش��'�6��?����?Ƀ�[�>����YSM�ҊZ>�JA(�4���K+B�$�����O}��۸V�l�R
ռ5Xt�E&���y��'���'U��'�b���$L� q牕^ ���ҁ.�,�d�O@�ĕꦝ�a}>I���MSM>�PG�&o�����L��Ji-k삵�䓪?i��|ƥ�0�M[�O6ԑ�� �U�憎i �'���b�;`���?�6 "�D�<ͧ�?����?91(
?.qM�w��<?ऺAa�&�?�����Φ��ǡ�Ey"�'4� ��A��%�\Y�f�)��[I����8�	`�)r�"*J�~�HX�VeA�f+��ڰO9h�����@�џ��|�e�+A�H�vg� �a�H1NyR�'Tb�'��^����4z��\K�eR#He�<�4�3I����/���?���6������l}��'��-sq�Ƥ?[�h3fCR;VC�!fU�������'�h��e��?�c�P�ہk�5|��t;wA���M/t�P�'�"�'�R�'�b�'���w��|����	N��h��TX޴QJyj��?�����?	D��yGEK!;*r�h���&JZ�B#)ŀx���'ɧ�O;Hӱi��I,eABuh�%�"�Z�z��JL��T�&[|< �'�'=�	ǟ�	�ı��k�,:$X�P`
u��	ٟT��ß��'^,6��-ʓ�?a0"L S�<"&e�	-%���E�H���'@���?!���_c���'cת����j�
�@��Pi'b�5P�&Un��'`�F����b+S�6�"�oJ>��7��x�	矈�	�hG�t�'¤�	B��W� ����(h����'?�7�\�<���Or@o�O�Ӽ�e�L5^�0�Ǥ� &�� I�N��<���?q�HL�� �4���I>@z�3�Of�䒁�I�PJ��s�P+���Q��|"T�������	۟x�	��4�&Β.r	j����%_�:�Aw	�Py��j��Bǁ�O��$�O@�?1UF�*m�D��kJ�v7�:#g.��D�O�7���6��1���<DC%(���n�v�d��O��<'���'L��� &,��"^�~�8�3$�'j��'o�����W�T�޴x5Jz�� �0�Q·'a��駡M�10P���N⛦��x}��'���'+8#�ȅN0���BG!o��K���������Q�,�����	����:��e������g'��ȕ6O���O6���O��d�O��?�j@d�I�H�Z�v�� �l����IٴBz��'�?I�i�'8����B���x{wa����@ɢ�|r�'��O�:�葶i��I=hR��=��qs`�ޜ�L��ȥ���2���<���?1��?��&�O���y@*<A�l�'(P��?�������f`���������O��$��=*n<�e
wzD��O���'x��'cɧ�	���Ł��%3�F�U�L'(�2XA ���Xb#���S�(bF�H���
�����J�jx�bS���)�I��(�	П��)�Gy�aӼ�8�#�'v�n-a&!�A��9����#>���OlTm�t��fW����4k@CőXau���˲"�mh��M�<�I�r�.tm�t~�$VF��4�J�)�	b�0��C�Z|&���T5LR�d�<����?Y���?���?�-��y��KR�zq��y���;Z�hT�tm�ܦ��BNԟ@�IΟp'?M�ɳ�Mϻ`V̀p��P�O�!�"�Ҏcf�
��?�L>�|��F�M۝'�0U* G�CF|+'�^�'�A�'r�1%��{"�|rU�L�I�Q$fUh��Ŋt�W�'f��CGZٟ���$�	wy��V���k�<I�[0��F�@���*V���a ���>����?�J>i2��8[e>���;��q��~f�5w��aǓ��O���	uL�f�8Ĭy�
 	i)�Xyf�ܩr/�'���'A���۟�@���n�D���\5�=0���͟`�ߴ@�U���?	��i�O��(j��u�܏J��H�A w��O��$�O��)��s�0�4��t�ǥ?�Aq��-=�5�� u��N�Ay��'Zr�'+b�'RFʄ(���2��.��xP���@*�ɐ�M�u/�:�?q���?�K~z�2W���ԅ1x�l!�֜>�z�TU���	���%�b>=�`K���2,[�2���9��,7���Ka�)?�s�Z\oB��������D@&%�P�X��eDD 2r�٥ �<�$�O����O�4�l������f �I�����Bvʟ"\xF��H�B�x�J㟼:�O����O8�č-"h�����-�4��O$rr����u���=}0��s���4�>���~b$����n�:P�T�C0pOt�I�����˟��	؟8�	i��)\S勑�wP�F�-0��j��?!�vH�f�H����'6�<��'\ ��q� 0P$���1O��D�OX���}r�6����< N�2���&
��ݛF晫�,�!�G^/BN҉�o�Iny��'���'���T�;�T@փ�?7�6UIa�$:���'�	�M;⍄�?���?�+� ���+ۮ#�� i� s�hy����R�O���O��O���	ȚᚂN�1'� s��^�6 ����uS���b+?�'���Ė��`��� ��,G.pI��̺*�b!����?a��?a�S�'��d_�)rAmE�~�i�D.J�-�p\kC��T�Tt�'�6�;�	�����O�1@��F�\j]�`dƷ7&��QU.�On�d��
4Z7m&?��qBU���2&�L9dp�)�8��5���>��ϓ���O��D�O��D�O8��|�P 1m��E�.WB����N�9)�& �5m��'�R������;A�Tĩd>R٢��
E�9�I���&�b>e#1m
�u�S�? �iso�>*�l����>�Q��;O���G��?��<�$�<�O����CND|k#��n�����o����162�'��O�/�.�Ir�T�d�`S����s��O�|�'Cr�'f�'�p�1�6@RL`��� =|�5R�O����Z?Ŏ\;�C9�Iؿ�?i�c�O��˕
7�l;Tk�4�$�5"OH|��n:r7H��
²&`}	U	�O�o�s�VU���|�ڴ���y�j��o h�5N:���cf)I�y��'SB�'�F��i�I�5��	B�ԟLA'��gbP)��P�,��QJ��=��<q���>+>��Y�m�4y֌�KC�ɽ�M��O��?����?!���VU��D&V�q2�A�D��l��?�����ŞC��e�Qf�rY$K$�V0#����M��Z���,X$-��<��<�hC?� Tc�`��+�l�Fd�~��IٴW�$�3��7#�q2f�K�
!^T���
{~D�c�D���d�Q}R�'6��'�@�b�j�q�v��Ӊ�=�,��n,�v���� F�2��T@�j�S��M2�K��T��k��
�X;���Ro�|��I�?;���Ճ��O�xh0�	2,����ߟ��I��M��W\���s�@�Of�8s� �D�1w֕s����)&��O �4��kPCh�D�"Na�G�)ZD�kD��F�%2g�My��	q�	fyR�dl20���٩P�����͡C��XYݴi��q���?����򉎏!<|�[f�M�@��	�P�	����O(��7��?���/�3��+����]��L;h��y5BԦa (O�)Y��~Ҕ|��N�`i�m�t��1y���:��Np��'<��'���\����4	
X����X.���e�<��Ч�¼�?���{\�����W}��'{������'=���(�$8���ѷ�'���F''�V��4��M�6��)�<ya���\��dE��sw��g��<�-O��d�O���O
�D�O�˧(?t�:!�(} �S`M�G|[3�i�$t
��'d2�'T�O`B'`��.ͣ0:����\إ�S��2��$�OT�O1�f���ad�x�ɴMd����&yC�Q���X!��	*M/�|�w�O��O���?Y�6�څpLM�^0�IC�`ߴ$X�Y��?���?a+O�o�8hӦU��۟��*[L~�-�����aVcë	[�?�Q�$��ʟ�%�X���W�Qk��[4�W)L��P�P�/?�h�j��y�ݴ5�O�0-���?��o۬ 1 �k"��+O�@��1nW��?Y��?����?���i�O�a�%��״�xf)�>?3�(�$"�OP\m�2g�.���ܟx��4���yg
ٵ��9�#A�?T�K4mO)�y�'���'��ً�i0�	U��ڟ^�YeJ
�Rs�@Ȱ�9T�>����,�d�<9���?���?���?y4�֌A�E���P�~�@0sM�����٦u+���꟔����%?��ɹ"*];3 �^�|�J��آ2� p8�O��D�O�O1��ax����v�!��_Ҩ�ha��	f��7��\yR%D[�L ������8q�sV�śp�����ڊRɠ��O�D�O��4�8�4��o�'d���3�f�$��*�h|J����]�b$fӎ����O�$�O��d_�H����jM�'�ܑ��j�8.������j�x�y�8�z���?�$?��ݹZ����w$W4���'X d�蟈�	�8������	@���]Q� \jD`��1e�H���?������������'C 6-'� �Mk���j3Y��=0��R�A��O"���O��ܴ$��6�:?	@d�<B�IB�Y8L��ݨ� hѣ���$���'82�'��'0h)��گY9�a��/�D!(��'��P�lٴUb�����?�����$�fmQ!)YB�����f�4a@�����d�O��$6��?i:PI�8e����#�!�fH���Ŧ�d(�����1r.O��|~�&�4"��Y��1�O�+�2x�ѩ#��Bٴ7��ܺE��o2���`�
5���;#��-�?���f�6��C}r�'SLeK�A��|�-I��	���"2�'���{@�v��|�d�fO���<�G-� .p�`�M� ���0F�<	*O�����`�QH4�N�p� FE��S~�o�/I������|�	c��t$��w� %��E�O��L�6n� elݹ��'��|�����ʛ&2Or$q#�
W���I���(S`�[�2Oꨠ���?�2%?���<�/O�Tg@�� \l����x��B��'�7�Ğv���$�O���5:ة�p�O�p���r@���qY��<��OX���O��O�0*��H�,�d��Z�T�&u�s����/�,x�l���R��Iџh�3l�=*�H��^+�|A07$$D�Soԋd�jѓf	�vBE�E�p(�4~2�()��?��i�O�n�1�(p�A�Y�$���OOl^��O���O�(9Dw�J�H��s��?��d΀�.������t��m
BGn�y��'���'�"�'��9�xsF�òE�޸�� )w�3�MCcaԭ�?����?�O~���W�4zr-љy*~��V��y���\���	ğ$$�b>e#�L0� �!��B�l{����Js�����
2K8�I��>9�S�'�p�$�4�'��e)C�߼:}�����I�B��5�'jb�'i����TU�LQ�4!A"њ��f��r��'�ZHI$eL�6��b��L˛��DLr}��'��'+��ڱ�WQ�D13L�1���J��6�����JT�ޏ0��)#�	��T�fH�h�KF��e�E�4Ov���OT���O,���O��?�b�#��n��@�X
2��0)��� ���H@�4"%@�O8.6m"���"lnX�x���]����%��_o:�O��$�O�ɗ�	�7�5?���B�2�G)��C�ҵB�B��I �T���8'�D�'��'W��'�29�BEӿX��! k̶
֦����'�^���۴*yj]�(O|���|����7o�p�˷i�Żc@�p~RE�>���?aK>�O����&ݳ/B���c+w�0Ex�K�_�^i�úi����|"�ʻ��$�������5p�R#�Pw¡�Vݟ��	����Iڟb>ŕ'
06-��*����$Ȱ`�dr#K��F��r���O������?Y�Y���FiP=�#BZ-x:}(��T�$�r��Iß�bY���'���*�O
)O��2�	�a�6Ts��w��hv9O���?���?���?����	K�rm�����q��L�^��s$&k����O�O����O�����D����q8�e ��ԥ��e��n���IޟL&�b>��II¦�͓!�45���!%Fh��D�H`1ϓAX�r$�O�$XH>�*O�I�O�9갌�Jr��TI�+��+A��O�$�O�ı<��i(t��'���'�&{�EQ�n�6���fu8f�_l}��'oR�|")� zW�X҅ɍ=^ ��ߤ��D�zd�SU/U�L�1�@�{��I�&�d� �Ę�O��c�ö�}	��D�Ot���O�D'�'�?�4nW�j�L�5��� AX7�S��?)g�il��R��	ߴ���ygj�:�:�ze��,n��[� �y��'��ɯx�
|lX~�I
���S�:��-Q�*�Rb����A�������|�Q��������ϟ �	� ��fR1g$l���tjNd��Kuy.k�@t�g��O����O����D�3�xdi���Q*j�2H�'����s���p�
�Dn�D��?k� �!N�e�0ʓ*��!p#��O���J>A+O�E�� �(��|�ǛoJ��L�O����O���O�	�<9&�i(��PV�'J�,s��_=؞᳣
U0y��X��'��7M:����D�O��MTbY�畧t�M(W�R�J��@y'ʇ��M[�O(����R�)4������,[?�\����0���3O��d�O�d�O*�d�OZ�?U3�Ϛwm��Y�LK�M;(���D�����ݟ�ݴU����'�?9��i�'��������҂�!z/:���y��'��I�"_D�l�P~R �YM�\ �9�,QR��r����ğ���|rT�(�Iԟ ��؟���	S��e��L=�ي���� �	ay¨g�p�#P��O���O|�'oo�A��OBK�f�%N��:K��'m���?�ʟՁ&�ΓNS����B�� ��QsBܤ:�z;���|"S�O����H���x����V�`�3H�"�D��5�%��H���!�l�@C��Wwf�)��B*��z�M���К���?;�j�Jg�7ze�jF�q�d�ٓ'HM�l���*�HO���ιm5�ș�$�%B�8�2>�l(�!��ȷ(�*y�(��ɋ�B85��S5)H���P��!}����'�!�ƅ2�#�99����(�'BP(�r�H��r�(�bWΓ�C�
��ET#a�\)���)x��Tʋ�n
���u��B��}K4(�w��%;�n�	#3<$���#����3��4*���'�����&�d����x��� L��,P�kR9���bb�Μ]��&�h�	ן\��By�bh��	w>�P�ř�I �O	�K�^l�-uӾʓ�?M>��?����~�K��&�̳��ŀsJ2�����d�Oj���O2ʓ9y��XG^?u�ɝ&�P�����b5�zGD+/5T����$�P����\��LaܓtlpZ�ᇔi� �LF�2�lП��I@y�ꇞ6�>맂?)��b�	[=��� 'C���`dH9�'7B�'^Z�Z��$�?u��
��@g�H怟
jż�zU�`�X�_�rU�ѵit��'f��O������Q�a��s��� �c��9��������X����OW�Y��FN4��	�4_��} �i&��[��s�r�D�O�韄p�'���);��W��":2.ܐ��Y,�\���4^��y�����O�k��F64:��8��τ`0� X즵�I՟<͓� ��O�ʓ�?Y�'p���f�1]L��q�GYA�$�ܴ��u�`L>���?���f�P��}COX�gu���̦I���)ЯO���?II>�1 �`q��cW� aXcCO��bh�'<�����' �	���	����'0�y��cLT�Ȕq@`C�<���r� U���꓀�$�O��O���O��P����T�~9����~~�թ��WTᲒO��$�O��ķ<����*2�L!h���hC�R���:��R�\͛V]���	a�	۟���;~�v����K0R�@&ղB�����b �<��O���O��Ĺ<Y�#I�����*˯r$�5�#�QG�%2���M���䓆?��pD�>�U`b@�1e�&R��	������1�Iʟȗ'�@"0a'�i�O����lࣵ�ԑx���f��O(�@Pu�x�]������$?�i�� ֡��g�8Fg��aD.�
DHmCu�i��.�V\:�4Z����8����DF�i�xպCj^'��L(��ԑ%n�&]�4���qK|jJ~nځ/����OёZ��1�	�	6�GQ�$nΟt��Ɵ��S,���|z�O?2�n|��R�)0'M�jۛv�'�2�'�ɧ�9O���˭7�,�[�m@���T�l�g���m���	џl:������|����~2��:?�F0 gD�2~P|Q��V�M3������3?����~rm>,��e���=tG�`�tR��M���0mdx�/O�e�O �O�aa�mʹM�(��!,�n�HP��+�D≑m"�b����]y�'ӄlHƅ�gvh���Ԉ'�
���d]���	C���?i�'Q����#�=�����  �H�2u�ݴiʊ��<9������O@0���?�j��i|�mz�DH1 5/m����'y���Oʓ;m�HnZ�7�4��'�σ2�~��3�@h1H��?���?�)O�KA�O��5E+a�5\��p�EE�E���h��p�^�D1��<�'�?)L?��p��G���X��
�t�!&hm�`���O���&ex����'��\cβh���f�E
� (a(��M<�,O����O���������������X�Ļ� �>���4������?!��?��'���T%	���b̚8Rpx"eS��i R\�|8��$�S�S=^u
qY���+B~x�Q���NI7�X=*�lZҟ��	ҟ��s�O�N�C�ne�&�J�@x�a��Jw���m������\%���<��Ytq��Y�6��q
�����s�i��'!�.68��O��f�OT��T)L`�, �)?}Pտi)��|b��~��?���?��%���AC���Q0_/����'�7+�d�i>	��v�B#��Ӄ��<�R�ӂ�G� ��-�O<�����?q/O���G����!lS#|�B��c� ?-$�S��<���?����'��䖨S4�+DF	1cE85�Bɚ+����U��$�O���O�t,གG8�ڐA���d�2���C�8X�Υ��V�$�����&� ���4�'#^�9u�Ī>��#&G�c�u��j*�D�O^��?Ѣ�[����O����Q.2���u$@�xĤ�bA�Ϧ%�?����ğ3�'�A�r�X6U�dDP! �N�H�9�4�?�,O&�d��$ɢʧ�?������ph�lxvA��&����}�>�'�H�	wy��O��R]�t�� ub`��GI;\����H��&����������?��u���*6�<�� )W�K;������MS���dR;Y��Af�G�9�Pt{u	Y�i�*��'�iz|l�ky���D�O��D� '��2CD=:�l¬]M �
��Ik��K�4�?���?�I>��y�'���F�*�L ��)�-,>��
�d����O>���I@�$�����K��0q��Q@����%�4��ulZџ8&�먟��O����O�0)����Kp�)X.B&{9yǬB��9�	YM���L<�'�?�O>i�E�s"��	��ѫX����bs��'�BW����П�I]ybE��M�$H2֦Y��T�Pw(�<K�>1�� "���OT��!��<�;f�2%�C�/4�����M�P��8nZ�$�'W�'��\����/�����%P�1j\�QA�)?����؜�M�(O��$�<���?1�~�$��
c���c�-K�Hv�؂{IZ}��V���I����I]y���!ꧾ?��#%Yg"����b�����CK�]}�6�'m�Iޟ�����\�хg�ĕ'���1ƕ-Pu�A�T�Q�hR�Y7aӄ��O��m!��X�Z?1�Iڟ���Wy�)�L	:Ĕ��$��$z�O����O"��άw`�IYy�؟T�ӡDțm��q�j]�F|�Ʒi;�	��h���4�?���?��'	�i�]؇H�*������Q�8�5Lp����Ov��B8O�	��y"�i��|' �t�Ӧ^����E@f��Ac1�6��O����O@�)�]}�U�;Q�B	�� ��'�����G��Mc����<�H>1����'oL\#�Kюwq���Ƌ2!R���b�<�$�O��DT)=��\�'q����|��e(�kS=mLl�� ��sO,XlZ��d�'�$�����O��d�O�e���K�B����F ��f�`�æq�ɡP�
@�O���?(O���Ɗ
wjF�<\����X�<p{�Y���f�Ė'�b�'Y�O�f�;Ajԙo���.E�Tƨ�����*\@����O�ʓ�?9���?�FJ߄�bX� ℗�| ��f~�]��?���?!���?�(OT���D�|"t,�8"O�x�r�'�*H�F����	�'IbP��IП �I�Nƈ�	�qFE�!���'J4�b �-��1�O����O0���<�f��2R�S��@�1��
�yनܷ3/F��2ŉ�M�����D�OF���Ox��W:OB���Y`,,e$E�G��1�J2��h�:���O�ʓYmH(A�V?��	����5�����'˾iΈ�HQfF�Z�ڮO����Oh�X0)��D�|Z�����l�74��=C�V�caH�s��J��M�.Oȸ�QbB�������8�	�?�s�O��7���@D��A��L�ui���'RI
<�yҞ|��� ^� ���i�r��_�V����7-�O����O��i�}U����J���ӄ��:� ℎ��MSсD�<�I>q��4�'Nn� R��s N2n=��Y8i��i�iNB�'T"��1U����d�O��	&lz����ǵ"�E�t6�-��F�W&�?�����p��}���ᑫ�
	I2���ao�ҟ�j`�[��ē�?�������/�T�pc(OL�qrƊ�}}"o��yrX�(�	�%?��V*Ɣ|8���8&窰�W@όl�`�BH<I��?�M>A���?i���$����	ĳ.>Ȣ%ԫ)�V�H����$�O����O(�=޹�u=��$h FO�e�D� ��K���xb�'
�'r�'��`��'	���R�U?6�z��¨+T.QP�#�>���?�����Xȸ&>�r%/�?�PiCM���֢���M������?��'x�j�{RB�.:�P��q^�F"��VF���M��?.OviY3F�]��ٟ���*:�:�����c���@�L�c�̛I<���?Q���?	M>��OER�0(�s+V�!�%,Ġ��4��d��/Hh%mz�Os2�OL����2!�][�*Xۀ̎1�Fdo�����	4$��	I�	Eܧo�����/^�{K��Rԋ�?�o�n���pٴ�?)���?A��j-�O��J�%�	�8q�)WnX�3R ����"@��$� ����3'�ё��'@,,T�D�0F�L�3�i��'�B��\� O<���O>�	$� Ab6 �2M$��)֭��6M7��G6aF��%>!��ڟL�I.H�z��0-�����S�{���Rڴ�?��d� D[�O��$3���°*�Né4ʽ�]�m�:���R��s$��h�'���'��O`�'C�@�޴�O�G���p��|�rc����v�џ��ɸ4,R����oA��V��)�,��1�����'^"�'��V�������4���N�C��1��DX���d�OJ� �D�OH��9|���ʍcų�%��tmb����])N�LH�'?��'�rR�D��M��ħG�h��0e�1KS,]� f�i[W���	�h��TF
�o��X50Q��I�f߉0|��%��u|���'kV���"��'�?a�'8Q�\25)��@1��:�Ė�l��!&���	ʟ�ASg~�&����
�8Eے�>Qv� �̀�`0mZgyr�� 0� 6�S���'/�de ?���R `������"��,��IΦY�	�����"Z����OIX\h�OJy�����m{�`��4P�JM��i��'�O/�O2�$B�|c�-,L�H9�̲m��dlZ+���?���$�'�P3��01hr��Ɨ'uV�`� S�'i2�'�l%h`g �4�8�'��=8��:px�hA��<���ߴ��'���f��O.���oml�.�tdH��c]"yt\o���J`����|���A����`hY��\#6�X/b4�'rY� ��ȟ���ey2@S�H����b�ԗuX����X�lk:`��#-���O���Oʓ�?Y�U�%����8S�`��e�V��t3 �[d��?����?9-O�p��]�|:� ˟dp����ř<<l�M�U��A�'�b]�D�	����	.Uc�����b��8���g�63� ��'���'�Q��R%���)�O��Z���)>�6Tb�M�t�Q;1h�Ц��	Byr�'z��'H��'�哱SrR�	�˜9��	3r���c;�| �4�?9����5�:��O���'E�T&�/S����#C�	"ՅA
zwl��?��?Q ��<�+Oj���?q�p�C{ݬ	�N3<�
$+z��ʓ#;
�f�i���'�r�O:��Ӻ��� ux1����>2�{�ئ�I{tw������"��Gv�� �,m\��a��H��6�4�f�lڟ����Ӳ����<q�$����f��:I�t���ȡP�O��y�'�F���?y�	� ]�����Ɏ�5ڲ�3�'E�'ӛ��'?��'v���r�>�)O.�����H0#��{���6��$�8r��x�v�$�O���˴P�?���ҟ����d�B ��-��O��	�&&�Y�|�ߴ�?d�5=���Ny2�'i�Ο�����8׆Ӽ1��	1�$d���: �����Ot���OJ��t���o�S p��������af�U��	gyr�'��I矐��՟\�E��
?���٨_-|`���Q*)Γ��d�O����O����OdȪ7i�OV��@�˄��
W�Ўn�f�xR��Φa�	�����H�I����'����۴t�� �̱~Īer���UF��'[��';"R����X�ħl�����=xԥp3�Ť%,"-A�iR2�'o�OIy���
)FpI�.J h��tBX�z��6�'e�'�B(U+R��'"�'�����`).T�Ǣ Vp�X2�"D|$O��D�<��NA��u׺q����Ea��Z�$g�� L��v�'�Bl��"�'���'��D�'�Zc;R��ǲ�d0�4�B?p��Sܴ�?Q.O|��)�)�

�a{Ŭ��|���o�*-�6�Ȩl �7��O����O��	s�i>���A��z{�=��͝Bc䰫r؛�Mۧ�'��'���y��'����$�:L�F���̥UH���1�o����<��	���d�<����~�a�i��W�^ Zb�m�9B"#<ɰ��T�'�B�'}��ⷡ�46-������P���o�4�DQ خ��>Y�����sB5_q���c@�,�N�1��W}"���'"B�'mbZ�hr
� �u���?�� �[�iǼ d���O��D#�D�O��Y�31 EC��5�je����s|f�`���O���O*�@0����2���bg��7\R�A�ɨC�f%��x��'��'n��'ۘy��O�m;Ԣ+�<�r%�K3&��Q��Y�\���T�I�����|�H��Iӟ@�ɠ�͉5G�%K	6dc3�C�Q�q��4�?1L>�������$6�'u(�c���q��qy¯Ly�j-�ߴ�?y�����,��&>��	�?�c�mߤ�%b,�6/}�aW$%�M��2b�5��.��i)�ȸ�i�3Ċ����܏pI�1ٴ�?���j������?���?)�����;�l�!|H\mEa=7ڞ$��i��_�D*�&�S��J��\A��b�� ���*l7�<8��pm���Iʟ����ē�?!�ԩi��ƍ"���lɃ���"	�O>�I�4ϸQqs�E�%{�	c�k��A��8�ݴ�?����?�����O�������6��l�����\�dT xA�7�ɲ�b���I������>�Ą�v��g�Yx��̍�zL��4�?yD�"wl�O���?���&�(�A΋	�Ε�K�k��hvS����<�I�����X�']�ՍW4�F��t�����x��	]%~c���M���� ��0W\�pa*�zpd���k8ҩY��=�I�"�"�	r��i�����d�UP����A�.��0���Ӎ)�(�S%� Q�x,���ۖk�C�3fM�%Ǥ愉�B��#$��$(�	����ؐ˯68��-ƐX��x����rP(��L��,E�҈[�HHҮ�H��+pJQ�%� 1�V̍����i7�A�8���9Q�g���	Q��|�\8�'*H�?�Y%�8�dL��v��t��oE\Y-
����&`Jh�S���
hq���Za�-KQ
����R�[\��CR��'-�i[##�="�I��T�*B�vj*�̉��C�p�4lA��?K��[�>Yp�M�5��´��!&�`���4 k��m���<d�ҝb��J
%NL���Q8��#�$�OD�}���M���cb��xTK�,2Ĭp��g��S���a��B�@�0*K����I��HO���@;8A�x��j�;,�Sg.}��'f���@�d���'A��'��w,����*�%�g�� S� �+��&Htp�Cd�O�����ߥ21��'Z���#+ �!�,8k
ޱ�N�;SG��� Q�+�O@�j�	Y�����RD���
�a߀��CC�Uz������dF/��O�ўpp�"!�h1a..,ތ��%D�T���W.��L�	�}�m	0�!?a��)*Or�Q��ٖ	�:�p��1��x藯�9!!��Z��O0��Oz��������?��O�ZT������ �Ĉ�he�؉��~��B�ɜp"N���Hۦ0r�M�(`2$C��¹(�,�&��8�Xj4j؞����-ê�&��(r�X+��)�`���Op�=�"݁ ;�a`�,ٞ6�̚�Z=�yb�^���Ek�aKZ=���"J�*Θ'�j��������lZꟌ��t��p4�-D�<�2 j�2Q���<y������	�|J�e����&�|���U<,8���=9E^tC��#O�Mѣ��.1����2hT����k��xB@F��?�I>Ae���uc!��V^Ę �Ν4�!��d�������z	�h0�=\�!����m�CG�<9���hD�3����B.扟{�ع��4�?1���i�59Qr�5"#&DFIܯy���C��F8^�2�'�JA��'(1O�3?���	�{��L�⥉�/+D�s��Qg�$�;��?eó望Hz ���KpM1�	-}R5�?�y��$�-Z���з'�ft|��Dg���y2CÊL��k�\?a2IX�] �0<Q��	kw�Hæj��<��Q��YO��ڴ�?q���?��(B/"Q }���?��y�;E�&)�g�bE��C�/.B��l1�	�g���U�|e��ò�AzDs�cѨ�qO,���'M����2���3q�ž' (P�$ſ'��L>�7�B?�N���Q�`Q��@�)�~�<��f��^6�e8AȪ/(�A���x~��=�S�O(.Ѱg˃�^�ŁTi�FJ���l�=V�0���'���'���s���I����'B������ۇR�jy�u�;�h��na<�Rm�X$"X�q���F�����A�A����[ "ljkE�6?c"+�
�$9_.>��!�O�8f�\��ֱn�6 d�	s�)D�\��mߗb��I�v���f��('��9��'L���T�l��D�O�l�P쒊xR��4GڏAF` ��O�	�2s��$�O��S(��;��q�����G��ʕ���?��x2gr�d��Q#`)��l�U��UHvA��p<���B�`&�� xE�я�]E���oRZ(p�s�"Op��6��s�hP[���$E�4��O�nZ��q��S0�Urd�&%^^c��*2���Ms��?�˟��z��'ʬm���f���)&hO<J�	�'��kW�T���T>��H���#/l�P+�j>(�)�OV���)�ӈ�<�;��A�P�(���F�.��'��Q��ۘ��O>��2ˇ4K��e�t�E=�X��'r�eq`��6{���\75�u�Ó$葞�F�E/��X ��P&̙��C�)�M���?���o�D Ed���?y��?y�����a�@�����`���I��'V�9�ϓX-��!ܾІ�E��<5Z��=�PNYGx�Q�-��L�%��M*Ya�FHQR̓]q�)�3�d��T��h�T1Q�r]�4��;�!��U%_d4��r��X����&ɍi~�ɢ�HO>��4	�/g	��0��W$Ѣ���h�
�B�o�̟8�I� ̓�u��'��<�.�K�K"M��xs mUYR�X'fɯ[�!��9{&@9�M��b�ܳ�@s^%ON)�MOy�blTҎm�
f�п���'�xa�&J��V)���Yz!C	�''��R-�,@��cA�2%d��{�y�H9�	�~�~$Zڴ�?��v��b�&{�RLh�J�;�b8���y���?������=�?9O>�voǁI�����N?;�6���	F8��A�,�I������^�bz��zBB���d�2x���|H�Ġ�@H�r�`Q��Y��y%w�q�!�(}8�5AB!F4�x2bj�@���\$C+�<�$;r�`q�dŤev�n�����Y�Tj�%�?9P��( ��c&�9%l0 G���?�>&�)r������p	&e�	\.8�*&}�h2�7}�X+�O�L�����A1���=!T�l��>�"DSΟd�<�j7c�=G��#�ʓ�dnY��aW^�<�.�"����8 �qWDR�������iO��``�)L@�ʲ씂N���'���'��qѢ��'���'�r��y�G:cHH�WM]�nލ���6-޲$�c�o�}����qC����|���>i$�|��B�=7a�S�[%�rm���=b��p��-�d�P��L>��`D	�D�J�F�@X~����E��?!�O����|����@�N�||ʡ�Bi}���юd!��B0^	$)���=qplL9��ST����HO��sy�R�L|���㇌Aўa1"W�m�|q��GO�;��'mr>O��ݟ�I�|�7�#j�F���Y�e9��9  ńY������I��['/��q�*=p͎�}�"���Wf<ag/�)}zp�5�Fs��`
�A~�\�	t����qj�by�d��4*�0� D�`��2=,�AQ�R!ODX�sѪ(扞��'~�j�|�����OR)�0�D"o����t�=�]� ��Oj�I4�x���O瓳X�`��7�d�z�a��L<� ��啟��x�-����'Xfe����cHy6�F7{�4��Ǔ4��%�	J�I�}�� ��/�����i���62S�C䉽.���A���"Ĭ��#Z�DL�C�I�M{����@N~ seĨ>��3^m�%[�p#�iD�'K�ә�����}�,G��:^�� �d��.E����O���f��Ob��g~�Mʕ'~֐:���;9��K�����@J#<����UK&���E/1���[�CO�DÊ^f2���� |F��Y���)��/��KX!�� 4�򕆖�m�����-W9DaxR)�S����QC���Gв|�0!5�i�B�'��Ĺ���A�'���'���w�c0!/͠4�sOM����󤅊/z�y� �;ovR$2��͐:�� rG̴��'/N���3�l�I�W:
����
O���J�y�I
�?�}&�\�w��iq��z�j�tI�X��4D���$�q��@va�[��-�� ?y��)§*� �`���p����23�ak������?���y¾�6���O��SB,ȍ��ZZ[Ѝ��XYP�<020��a#�R?q
�:EL�z�l��F��6��C��> q���6 �F�Q&�@%�ū���O���� p�����z�xq�6�^��J��"O��bω�	>j����(w�p� ��UW�U�4�iŽi�R�'�)*K7}�������J�
���'��$�$���'=��,K�R�|���AK��тY#\����fZ��p<qt�IR����!��m��c�`	`�DY��\��	�g��d!���)�ب0j�?23��qpF�r�!��\��͚Bl�xzdk#ţW!�$��Q#��C2�SQ�G�B`g�%扴rQ�h
۴�?!�����L8���K7^�h��7vl�	]��b�'K�� �'�1O�3?!�ώ����'�A�YŘr��t��?Yc�ߥi�A��ߒX�(����3}�N׿�?!�y���g�$IV�"6�C2u�|��3g�4�y��ϼs�n\QQ$&p��Pe���0<�鉡`�>0��"1��2'Æ,G"�ڴ�?Y��?�-� CF|0��?����y�;2�����6E<��"E�H*LԘ�y2)E��<Q��8��afl	�HӸ���$O`�J�Ԅ��qD$`�ѫ�� �[bA�� �4�<a"A�џ�>�O6=��۬Y�qa�J]b=��"O���֎��c܌|H&@�5�Ը2�������5`/���7o[;zy����iT~h�9��ԉ|����۟����<�[w�R�'L�	�4e�ZIɰ�R�]z�#v)ךZ��J�O����ؑ]P`Q�NܴU 6�[�G�4!�Dؐ]>@����D<%�,y�.�*�L�à�'/��%U&BB!��n�'�<=ؠG���y"�2��p���!�F� d���'|�b��P*���M[���?!�`�)�+��D�6`��
h�9�?a�'ϢU2���?��OUX�
����3_Ҵ`�2&�V0Jt��g�>l��	�g�P� 	a��iִ��t �\��3�;O�I�2�'��'��	[ҧO58�NX���L�z܆|!�'����3JL'5�8��ڃ(p����'7-ȓ	�QcLB+~��X`	Mx1O����K�)������O���Y�k86��� A�e �0B�#)"���?�vĂ�?y�y*��ɵS&���@KE��jq	�|y�'�������S�b
0�G�TO�;H׷)��'�����o�S��ᰄ�F���
Y��AUq7���d�<l�ċ� �-i7��?l�%��'�HO�W�m����nL;	D�����Ц���ҟL�Iw��)R��ϟX���������B`���/�=
P�ن=�n��E�l�ݶ9�牀?b(�v�9��ݐ��!]�x�ԒAM<<O��{4B��crm���d1��.�I�����|R�� ��hx'CU{T,�$��?�y�a�M����	��P�F%k4�ݵ����}���Xa���_<�����b�4e�׊H3�ѐ���OF���O���캣���?��O7�}a��	�0�R�3'"��k����x�����b�@���Lit�7J��	x
�'���zgI�yl�h �ڏ[�r$�aݢ�?��3�LL[�`�]��H�g$M��m��P��a� ��ZHB���Ϝ�Ѥ��<q���I2n�ȟ����2yF=
�i@|�@���μGRY���<���������|2Q�M���'�S6E� I��9�mC�AH��$@-O����$^.g܀�#�
���I��e.�xr�̎�?�N>�үN_,�tSq��9.��)�A��l�<!%�@�c���6A�(�s��c<�ֺiJ��1n@B�r�o����юy���7-�O��$%��HП�ڂ]H������5ipxf%���	�}����IG�S��Oި1Q�U�1�~(�1��Fȋ��Q��ɔ'��?ŻDl��=��;�ET#��{��*}����?�y��d��6A��� �4>�����y�l]'eHN1q��[�;�L ʧI��0<���I �n�[d�X�Xް���ݭI�:�4�?I���?��ߓ@�,�:���?a���y��oa���u�	����̜�<�����y�(����<鳦��|������ϘO�TbծEFܓ,!�!��	�����T�3S� �S�	��<��	ǟ�>�OT��GoR:#SlRc�94�*�(e"O� rxSb0W�$�A]�s� L�ѓ�T����Ӥ)=�m��+��sW�J�4�Tz�^�����I��h�I�<]w�2�'��	ٛMFT��֤_�>aD��gϟ�p�8�H!O���fP�cN.��M�7u� a
P�!��P�c���CE�ѲzV�m(6�ІwK�H�7�'����H�:/X�'G<�R=�5\��yb$,�n�0�����,�1�K��'n`c��+�e��M����?�@D�.Z.��h�SQ�\iسa���?!��J��p��?əOh.t�������0�B}�♒wvD�#�����W&yXRH=�D�8����];g�xR�ÒOv�x��$�?Q���?���n��}x�`�.Fk@�G%�6L�.O��<�)�',=�,�Y��i�PgZ$���S�E��.�#q��z�H�	�y�Y�`TDA��M����?A-���Ygf�O�)!A'"�@�6�� |�����Or�/V�P��8�|�'	Ȅ�V��ň�L�ʞ��M�J�"5�S��=�c#E�f>"0�!N?y�P�OrT
 �'�1O񟰵�a�<.k�|� N�LM��R"O8��eƟ����9����?�����'�#=��Ԥ\�x�Pf#	E����p�e�<Q�
Ͽ&�j��hS��A�JH[�<IE�Y7]'�<�#ꕄ{���'��@�<1��vA��8�>e�D���DJy�<����� ,�����(F�4Ɣu�<� [�q쎝�0ǚ'��y�q�<)��عkp���hYi�N��v
�D�<Q�LY�< ,9#��#D�-<�TB�ɷL�^=��%�%)-��FIZ�Xz6B䉁~x�j7%?G�$ W�ԙ_�FB�Q�^�R#�w۴Y��a��Q�
B�'Qz� ��"p�ppɲfVOgB�	���ɱP�6�A��^"��C�	D6�[q��^�f�G$���C䉿�[��I�*��x2c�&m�C�Ɋ>r���0_��c�̜o��C�I�Y3h���n�,Z/�	*�I�H�C�ɝf����R)θ|VZti���p2dC�ɱ_hk%b��r(�2��{�8C�	,$�Έ�@�)r|\����1�jB䉵v��dѕDE	0u,9hua�y:B�M1d<i���9E�����Do@�B䉍7�Pi&�;B�ۤ��l!�B�I�TS VXMI�q.Hd�vB�	C88�@#��v�	�#��1t(8B�	�-�� �Ӧ��\��S1c�:"B䉽:pR���U]�(��A�1��B��4���'�]�~`�pBiϋ-^C�4�D���6!��$���7y!�ȳ'�a���}I:�`�@4i\��^��x�ؕ�ܗS�%�q�R0�y�\� �H8SiD����`!��yB�܇dq@��U̙��E��Ȁ�y�D?I0 1n�&H���Y����y�Ѥ ��5� 圳/�ډP�����ybcS�줬�ӫ�7TA�²K��y��i.�'�<)Fx�F��y�l��H~b�Q��|�Dl��@B��y�7D��	A�S5|\�qA��0�y�g�3=�4c�O#z���1�H˶�y�m.O �jamW�"�J|l�y�
M� �|��¯�'��l@�P;�y�kE&(R��V
jqzҡ��y�ʖ��e��A=[S4���L��y���/L�d8��3VD������y2��5s9�P�E(FTp���9�y
� �9�C�*��Zg�,w��y#�"Ox*��0`*��ꢀڧZ��( �"O�8�'L�Qp�0x �ʊ_�b�Y1"OvEa�n��i������N�9g��1R"O��q�ħc����o��za�%"O։��}
h4SnR=`gR�a"O��*��rK��� ��J�kK��"O��a*R���Ap� �L`�z�"O��(���]�t���O, O<)��"O5�S��)�P�2&IȞ��q�"Ol@kU��(Am�F�ʍcr	�%"O�x@g�� �A6�Wh�*� T"O �Y�
F2��4'˔@*y���'D�GIʭ_r�� �q~�qb�!3D��j�Ŏ�`�dX�+F
b&xI�1M%D�l9��1\���c����l8v9�-7D��`�mR�\?<�,��^��5�4D��)�� �<E�xᤌ���N�C&1D�\2ri�3?b���ηzb�d�e0D�L��C�:���u�J)Mr
m�r�:�OM����?5ԭ�c��O�� #�8Dw�@�D�hh<1%�C��,���*�2ՔA��Lm�'�\i���/<`��~�boU����#2ᕒ:��t��	�c�<��MW1Z���b�ؔV��j�J�۟4�EhQ�)��m��>E�TLM�c����qo�3H���J��O�!�&pU& ��B[��\�QI6���	ieJ,3�F&@ay"ɪo]9"+�crT{��tڀ��V�<§,l���$���'��4�iHB��ɺ=
�'���he�@��Lt��ўm�L̓RnHQ�%�1�u��O���&ΐ}�Y�U�'��Jߓ\ͮYb�L�>I�D��/g�a(���*f*eR$%�<��f�������8�7�۬����cdK:���!��dQ�<L�E��HϴBx�J��H�^(������$�Ǌd������k���T�'K�ɡ'-�H���Qj�	&P�50�~�1O�Z�OR��p�Y\%�b�IB�a�>Ȣq��2f��T���K,�졄�����u��KW�r��B�A4�(!�\Y��pMA
';*5@��2uJZ����9/���>�� a�3s�Yp1-QR`��K�!\OLl��<�剫U��pooK�,[��� 8o&�YCg171F��hѢu�n��n"�Ӓ/�4�&U�5CS$J���i!B�{�dL�=��!ԿA:6�E��N̈́JjFi�kN�U;,a[[a C��|�Fh�gV�5��`X%�6PD�Ї�	�>L�hH(� ~�<�s1�� g�q�[?1O��{�O�R �7� /7���!� �z1"��JRв��ƚz���e�m��i�U4Bt���Q8|�8Z��-AY[�#U�3���ɝ�U J�B���5��U�2�H
�\��RT�c�;/h�5��{ ��ʰ�Cr���������P��V����ְ;U���΢ʈt�g��?���U)t�^�[PH�?�����кCb/}B��4�z����t8y e��9��'��q�7�	O �3��;l�򴙇��z|�0��`@]�E��-_�9�j�����X����IAJ]ax"�#�T�5![�P z���N�qb�|��Xr^�3�BU ������' Α�'�+c��|��gl�4^��$ �ak�}��o��t��$1\OU1C��2"�P�Vnʇtp8�`�@@5s��a6�/e�}J�cQX$��)^��S���:u�=��T1JY(�#���2�Ґ�9p��IV��!w��c�P5Q&}e����>271O��� ��xr DQ�q�S����7-�!u�e�W鋰/	0Qa���J����56)��3%Ձ,*�awK�CG6���FV�d= ���;67��r�l��dTH����䖁c�hc�x�ׅ��f����)�h'�ɢ## ���9�̩�!�]��l�'dй�f��kZ��J�*�9m]���A�;P��I�Q��I��I�0$�2�d�obT59�h�:!+FDG
	SϦ��"NE�C���j4�|Z�%xmRpbgoG�C�,5� ߁T>�H�'�����9b$�3S�˙w�8|�c��01Y"N��?y��5|��(�	���T����q�?�*����]��@�� �yl9�O*��%k�."]�\8!��A���h���-`6� �MߧW��p�ϭvY���޴̪ɻtJ"�?����c�YDu*9��(ԕ[ن�	?{Nj����-!��pD��?Zz�B�)=:x���N�Vt�)���
�? �������UxH(0J��״
�̌����3<��ɏ)���[�E''�ʰh%�P�̧U�P0�}>� L�C�V�R��A�E�`���jP"O~���̎$�zRo��-pk�m���JǛ�guf�؆���n��b�?�	����0��+c�Λ�f���H2L�!��3p�l�k�G2Ҝ�ƯI�$�zU�.�]06!;�+ݙ*|��K6�O&��1	��Obd�'�?Ţai ��?��P��'��(*[#I\ �k�`��� ���WMb����e~ ���o�%�~2M�*�Ї�IѼ��$"z�(��\���'���U�F9Jd�&*����V8���*j>)2�o�z�G��)x�8g�ͻ�y�ř�6�ƀ�va�+%Z��Qj� Jڜ�h'b�,����p�b�VY����w�!�M��Nm����I�,e�
�:�'�=�"�D�]n����Y(�l���3h�N�Y��n��{򄂄7T��bg��TB�C�Ź�0=�7M�-j!�RTg���o�~A���$�:���R/k_�C�*?�X��#�8=�@�`�4\fb�@�h��f��G��>ki���m��r���2�$0�0B�Ɇ;�d�s)�2H�*}���)J:�l�'DV�ēt�G��O�Ђ��Y`HBv�I���4"OhШ�M�Q��a�$]�E��H���:��5��'/�M��Hڶ	�L��y���דC���pI<���Jج��f��o�%dH!��$oT� "�F���43ƀ==4!�]�V������ j��pO�f!��ՈUFR�Z�I#�̉b��Q&~�!�˰kV�ȡj'I�&�x�#س5�!򄋥R���pc��!� %z��Q�a�!�d��VdA�ƤD�[���c�A !�!�5V��4{�ՎF�
�P�S+&p!�$O���Ի$�;�������!�@$8pp�;pl�cb�џf�!�F���=��G�ye�9��QX�!�dţL2����>X�t��ֳv�!��4�t��B4`���צ�7q!�D�?Q��R�Ѐo�L@�FSw�!򄃓:�d1FE��������9|�!�X���0�G�+����ˀ�@�!����Xh�G�BȞ�2��O!�D�7L\�x��*_+���h�+Y?D!�d���0	���Q���x�+]�~�!��#"�*�ছw���ۂ�[��!�8�I��̺,Ąx��� �{2!�$�PR<��e�G�z$q0*+*!򄃔�������z�ڥHN8�!�d�0h_�,e��̨!gm�%Jm!�D�	$��y2a"t���͈�PQ��{�E����*�5��s�8�+"�T3F����e"O�)���%�
Aٓ���E�*���8}�W���O,A���B���ˮ%�fuH��ݮ
A
xz��ފ)H��}Bu���ظ�8�I8q�4�[��'@X<ibGװ/R�s�o��Z�dĊ��đ"~d-H>ɉ���S�H:r�̓!`TZ��X*>�@��=Yi���Dmt$�����'���g~��I /�0���.O}}rc�22b��'�8�&�Щ�.i����[y�L��4OsNa�g��<ɰV�u3ʝ�F�0r���B%c�<tI�|�`"��!{x�+�I�}mp�r������N�pe�[� �.IH�#�[���"O��RE����U����C΀����/aX����|r�����xn0��5b��4���03	"D�H)�m�;{q�!���d�J�3 ~���' $b��dģ`�8���bX�b�
@�a�!�䀣0�� ��S>S&� ��V=3�!�\0@$t�Cu��{q$���]-!�ވB��Q��ʴb^z)Vo·�!�]2[�QɡH���l쨃��,`�!�U�
ib�����@���R��"!�� b]8��ͦ>�0��ML�HŃr"O�QbtKԫC����nS�n�@kS"O��Zϋ`�I�U��
0}Ba�"O�8֦�)<�ȱթ�2��<��"O��jb�*p��``�i4rh�+ "O�EB�,3�(8�&�P0V]0�)R"O Q�aDC�,�#��;V�VY��"O�d�`O�^Eܜ�����p��r"O,�@e+N-t�:-��Q,S���f"OYH��7TM(���m��U����"O��j%"$+ɞ �w�I#8��U�C*O|!ʠe]�4d�Q.��>�|��
�'뼶NF3H��l�%F�aq��a
�'�f8he,��OdV�%���&�	�
�'?rL�r�4o�<H�)���8 C�'k�U�tAI�`�ʭ��#_���'�>4�rb��;��|�ר�0a�'4�	�cO�X2t��'E?�, (�'��pw��q�J���BH`�'Ov��(K/i�i:e䘿�<T��'�\�H�T`L	  �
#��@�'�R�Pd���hS��v��{{~���'�$3�ǂ1	H�0��m��Q�'R	�cϗ���S��a��H�
�'���!�E�H Q��KJ ��'p����Fb�9`B��x�D���'�N��n� /� t)`��#��Q�'�����'u�UyT��0@i
�' ��ufQ���Q0�b�6'���'E�e`��A�ud\�T+��T����'"��cRMS�8��_p�u���y҆R�[�^`s�.�r`�%JKL��y��+@�nU���i.nq��/@��y�$R&}�^���\�Z�ؔ�.�y׉Q�^�p��4R��D�y���H��H� 蓫g�Y����y2�W�\B���.�p���.Q&�y"��8׶l����s#ԥ�y�G,T����\�@�@R� 2�yÛ@^j�+�9���AA)�y�E
.����V �� y^=h�� �y���`�(�Yf���,�nT�ʃ%�yrk
r�
���[\��x�4��g�<��o���7�V'z�� ��r�<�@��=7�䔠�i&A��� ��\r�<Q�(N!o��"@��#Yxy���G�<PCO�O�\�9F$��paȀN�<YpK(��Xc�D34�S��	R�<A��V'.�2`��K�?`�N��flI�<)��-e��T���A�B�8��bF�<�@��S��	�G,q���a�F�<��)J��xBiے\*� �D�<9V$^�k$ҽ����M���v`ZD�<�@H�o���ʏM�F0y�o�}�<�0�зP����jÉ,
�	���^�<r�D�(}��F&{l�h�+^�<1w��L9>�Z�&O�R_�� �C_W�<�T	�|��I�P�������G�S�<alT�g����v��12���4��N�<��˄(Tz��zF��.�ݠ�a�c�<�BNI#a�V�q �� &v���X�<��/۲E��F�/#��3�d�}�<�D��z�@Y
�n�>����VF}�<�u㜱6��(��\�(](�� �A�<� ���!͈;ntK��]60.��07"O�Z�Ȗ�E�vyz�蟹s��q"O�1�v�&�$9���q,���"OJ�%@��.���`צ^�%����Q"O���Ε�9Q� 	v��r��;4�Ip����Mm�H5h
5kLЙ�*�!�Ĝ<?BV�"�O.p�Y���¢C	!�j��(��=Y�E{�鉹0�!�d�G�a����{nV$���˪vA!�D�~��J�㗯S^2h�(K�g,!�$Ϙ��5��S�&{�8�(�z !�܆X�Z�釂��7d0]��	�Q&!���-
�)9�	�*E��3&�%!�$�7Th6a@��$:�*feE24`!�F�)C yS'��l���C�->F!��RI.أs�ZRG�M�B�8T!��0r�r 9G�?b)&�IeO"�!�$_�-ްy�&ԒP��I)��ߣ �!�DVv��(u���Z`�R`��q�!�$�mkh��@�^2OxJ�z֌mq!���!Vv|-9 �A�%p��"!.$�!��J�� � ��I�@�tLh7�X<	�!�D�A8��X� N�s��	vh�?�!��߻W:,�Ճ�|`�@��
#j!�$̡E��u�!O>��d��8`!�$�p��1s� H�`㨎^_!�dʺ@��Չ�C֗I�h�p��JI!���7X:$����׌�T烄N%!�ʁ1$��ŕ2|�d�y�l�4&!�V0���H¬6�tqp��5w!��ϒ6ª���4C� y� �]�lm!�䏥iPR��k��ZD;��>e!��\�{���+��q�V0�dςgY�䓠>ma~r�qt���sM�.Nx��q�Y��0> �"}blD�9�F���X�B���:�N��y2%�p�X[�l!6C(�H�`:�O�C��O��볫�LOj���Ž>���'/��	>E;0�I(c�V=��%PT���>�b�|�mȢɦQ��*P�ȓ#����UeYva6����8�X��	$��?��"�#M𢽒�B��%�Q�ii��t�c E�N?���'Z���E��DD8�(�o�� >z���'�����SES��B�u�iÌ{�'��zc����X���G|�q{4a�b�i�"O�y�"ʋWd`� ��,Rڌ�C�n�'�"}�'ʰ�y��G/c���IWÇ��a	�'�6�с���K�d0��KЬq�
�'N:9�TE�9Ħպ!n��,��'IdѪ9�p<���+V�a�'�Hl���N�O���� U:A׸8��'�"�[v�S+M&M{2$B4?.� �'���X��Ѹ;Ni�QA�C��)��'@�᫑CE3�n���ڌ@���	�'>H�;��ɪu�\˃i=��h�	�'���b��.������/0h�1@	�'�p������^�
�5(ښY��'�Hy0�A�v�0Y�UA/z��ؙ
�'�A
�+̵�F�r%��!1X�k
�'��:��Xq�����)e3
�'�ڨ��LΒ+����X�Y1fP��'*���E�M�mt♂��#z�t��'�� ��%N.2>�����u?,�h�'<���7����rH%|2���'��	��L".Yf5��B�l��M���� F��5����V��O'� �"OV*E�;*�n���*g�����'#�$E�����Н[Ө�$��g!�D9|�e�Fm��+�d�hPMӨ1n!�M�mZ�*���;�B���Лe�!��y�h�եֻW�4��/�@!�䝧OGЁ 1��5e�@��@F�!��Eb<�l	�,,�0ϙ��!򤐳6��U@�5�"��=}�!�Ă7�FE�v ��?����k�:}!���hz�q���:}[�	��m!��,m�X��܊'e�iO�=e!��7��Z��n&p�+���5e!�F?;�dUX�� D'nE�-�!��D�F �Y1o�	D�(��*D��!�Cv̘�b��nd>��6
��!��~F]��I�`d*qr��1b!��*.����&[�uD��XE�ɗZ*!�d�9`ޤ�AO�;I?�0@F�1y!��ǈ4��XP@�>��Ԉ���=�!�D�O��Q��G�}��Q�!�V�qJ�����b*T!!Ȯ �!�D�.Y��e���[.��ұ�\�L�!�To�5;G$Q�H�0��*�{�!�Ǎ1g긁�[f����2$!�7dH �B��8.��֍�
�Py�B�p��@�m�t�P '�։�yr"K>� tRe
�)t �0�*��y��"Tք�2`�t�9�5���yҩ�#k��	��Ǳh����u�[��yb�V:���8%hB�5hH��샜�y",U�@d����u�Y+�L�y����H��G�~����yRЭil�@��	z{BU�`�ߧ�y�@ߢZ\��H���>2�py�����yr�S�&�l9w�7G�@S���yr�D�w�%	��=�VV�.1|���.�jĤ	�r=*�Q5�U2L��ȓJ�:��J�_|��sp��/H�&ՄȓL+��w���.�@���.e�,��T谨�,T�A�8B�h�3!���ȓ
��#�3<�l�br��:<�ȓ'��}2��݈zL&��O�in�D�ȓpi��kEP�x���&�Զ0�0\�ȓ!k���e"_�q�8Ë�0z�P��ȓV?�B�.J5_� �"t�4}C�U��Q �̩te��A��=b�a�
- H�ȓ|��aPK�Vg��	7�mת���;���� \�\U�I�΅�-[p��I<����h"�e����>�\�ȓ8~Q�ì0�����
�3=�2���9������68,a�,w0�����S ���9��I 7gӦNĄ��	a�'��E��C��&I�W��n�^���'����1@�����6(O�X�v�
�'9�t����&a�*Mt�H��BК����)S��u���ʝU}��ȓ+���萞M�|��%�Ix��P��Ѩl��ɛNy�`�C��T��]��F��{�bȪn�b���ϨyVń���-Y�)��iR.\�H�4�ȓD`-��].^���h4�5�☇�_���1��VU�F��?[�|��-�p�f^ e>�h�V,u�x��S�? ��B���?@m7���.OH�4"O���vHW�3�z�E/�046R��`"Ou2S� Z���Boөk,����"O�Q�F�'S��)Qm�m&Xq�"On�J �%W�1C��9Xt��"O����Ƙ�<��5z�a��N@���"O�x�(|�n�J�%HIM�"O� �a��8s�r #CCBE�'��lZB,V�!�Z@�#�Z� �zŃ�'l �� ���R!�E,^�J���
�'���	��ϒ0�&[�dǷ
'R)q
�'�fd�đ�UƼD�2�A� h�$�	�'���1`�2eٚ��V={K	�'ӎ4�E�@ȝ�@���v� �'٘���C��[�^�{@/%�r�[�'z���U`ڥ�
�'�Z�wp��'!�L�c@�.�p����j$�X
�'1���P.˓x���U��P���X	�'��k�F��c�V8��Em̤��'+\�а�M�7
h�:b���9Id,�
�'zh�R��4a��ĭ�2���
�'���Ye�Z(fnd=�D+��y����'@�˗d5o8�L��6�:�'��ir��/
ظ��L	e�B�"�'˰�"���R)�Hՠ*����'�
�<F 4�� cY�MJ:x	�'qt��g�Uq ���.|���	�'��AQ0���'��'�I�#�!�	�'�N��,G!�@��k,-o����'�D�0&^>f�Ա���Dl�A�'�*	�$ :LO
4S@�+�����'���a!��n�1���������'�ʰ��E��u�O�� �'�j����B� ٠�&-5
��D��'�����$�lq��":
!�'���ԏ��K9�����<-h�<P�'6l�R��>��6V17�\)a�'3����m�
w0Xi���/%�z���'i�͑t�
 �f4�C�#m���'2r�2�F�j�i���<n�Zi�'&�iX7H��T�#dE�<"�8�'΂��5I5nr�`c'�3:P���'zF)���޻{���S��4k���'R~�Vi��w�T$��`�:��J�'3<������;�`���B�d��'�,��@$J3ex���=B5�'����U/H9���B�a����'�l(��۔BoJ�x��#c���'vN���g_m0������.0=��3�'��<������P#�ַ!k�"�'��i��nO:`���`eN,�9�'J�)��ĺBE��ևծM݂�r�'v��"b�	>ML��u��L�f�p�'�v��&/O�&P���� PK2~��
�'�6�2�Ad �SCS<���'�r�腮�.8Z)��@��g�V�x�'�l���_�|f032��!dM��I�'qd�Y+[�S�l��B��
V�"��'jX=[�:w��|	��Y<UFV��	�'���v�A�N�3J�M�n3	�'���'Te
.` �o��{�nU�'ʲ5s���h1^�����\�3
�'�l�B#Ӵ<�<]X�kX�~#f��	�'�vLPSl�	Mު	�ʔ�qI�}���� ��ʢ ׂ�^a�7$ܶw�D���"O^ԁe`�*��,�1���w��P&"O�)aEĤ*�D9L\�`Ǣ�x�"O���$CP�gnbTy 놎g⚌�V"O~�AAa���Y*����sl`��"O�T0��2d�m�b(~d�$��"OHE�#�ޘj���S�o��IR�"O��v�ŌO�Z(�Mǭ?RL "OD嘦�H_.��b׫�82J2��s"O�ۣυ_JZ ��N���]�q"O
x0$	�)!ʮ�۔������q�"O��r�]��!���\�(�ִ�r"O�dQ��3b. �4%�z)�B"O|�ˤ&T�Ȩ�v�&�j!"O~���>kwB5��E�=%�ur�"O��C��*d6� �
(�m �"O��3���m���n6�#"O�Q�Ƞm���#�H7w����"O*�ҧGK�F�P�hF^�#H����"O:�S�,��? L��$ʉ4"FJ��t"OJU"LӼ�r����-k6�B2"O,�����T�^11��[4>!V�"Onh`Av]x<�AF͘c�� �"O���''��)J��$EǳlYD[ "O����+��w�($x���(�@<�u*O�5S�M"��!�ܝ5�,��'�2��v� �<g^��b�9k��Y�'`��y�S	����,�@(�'��`�W"�	4RH�1�+X�:��2�'t!����x�QV�Z�@a*�	�'��`�p���wB(�إ���@$��i�'^ӅBo�����Ƙ9��4��'��,Am�<�8�Q��[�@.�
�'�:�S�g�`�j�kq�� 2���'���b�I�/`�`���E�;dp�@�'Mxۢ�ım��Sa�G~�x�(	�'3dy���¬>���n��jvv���'�D��L�U���A'��d�tȳ	�'�1`�fW�N�Б�w-B�q����'�V�]�R����&H�A���@	�']�d��&]�Hx���׃
�GfdX�'�����d���(��GyVԘ�'d�\���/B�4Ӵ>�ji8�'��H��oT$�����?_��ч�\8�,
�c�;����5�����ȓ ��{Ԏ	�&�`����*��@�ȓ_l���gت3���� hަ(xD��h.M�A#'�X'�(v ������]�a#E
Ht�y3�&7h$��5�R1so�9�0�#$�_$I�	��0D�Ր�ѝ#c�Ļ�I�@` ��ȓ]~�I�ꛐ�L" Ћe8��s��CT��5u<��W뇄9G��ȓ�L�C�3b���*�a�>Z�4�ȓId���"˩gI�Z���:6�U�ȓ
	@}Q�%� ���r��:4T�l��<���g*D�ĥ)`���0fv�ȓ53�������d~�� ^[�<�AH����Y�hߩhQ�DӁ B�<	h�&\��U��]�s�����{�<1�Կ|
��"�*k�X�h��r�<$bW9cɜL �ѝEzL�C#Jo�<��MH5�4[��B0=4�В��j�<�$ŀ���$ �W#��x���h�<� ��0��ۑl1���i�up@�r"O��;w����}2�>�8��S"O�t��i���0�B� ܱ"OR�cw�JA�4���8�P�I�"O���aM�$�Q�aB�/����""O� @틦���#n-_�H黡"Od��(��P����-ɤ;I��$"OD����
`Ҿ��JD���|	�"O@� ��S�~4y��M���ɔ"Oڕ��/V���a%��"OP�AO�PPdY#��)g`�(�"O�yZ�I� ��`[��6hT��C"O<9�Q`�#�nu���='�i�"O���f��NЬ 3��Y�z�z�"@"OF�"���DśЉ�;��a�d"O`�X��]�$d:�I��#�d�x�"O"��Oؕ0T�10�͈�S��m��"O�|:r'��]� 1�'��~q���u"O�ݰ�� Z�6��6N	�`Y�Xr"OJPT	�6@���[�VK^s�"O��EBT��UZ#B�|&�$�"O�T��� 9�N���D�4)'"O�$�! �?8�\�y��@;Y'f!�C��F�O$|H)��>N��lx �����	�'���X7��A������Ǝ��	�'�"P� &W�8X�hI3 g�J	�'Z�ui��: �L���"~YD�ʓq�H��-S69�q!C�&}`ȼ��v�y� dW�Iњ@����(7\e�ȓz�hQ�g�`�J)�
0un�ȓc���A0���p�պEϮ=��͆�	2��wF��!��4��.>���ȓA�.��v�YT��A��z�ŌG�<�#�A&:�xIǞ�b��e�D�<�%��P�~�%���0�J��Ɵ��'aɧ��dJ��u
��@Ws����  �!�dȯi�x !-)`*E�c`D?V�!�d-������L�d�¬q6j��Q!�D�K/���,ͧD��`'�
l!!��*%BEY�C3Z�&m�� :!�G�.�&�w�э#&��:��Ͷ2!�d�E��%��P*M��b[�~ў�D�I��4��pr���<�#��k�'�a|B�ςs\dU��D�;w�h��(��y�ɟ?j�t 'f�k�t|rp�@�yB��|��|� �ʓRg�d0����y��R&�0@��Έ�?�1h�,�yD�G��<Z3@���:��ÄQ���=1�yR^]^ �
�nE�Z�`M ƦѼ��'�ў�Oi�ԑ�)�,�`qzE�[�T��a�r�)��È�[!ZM�s�Kd�,������0>)SÒ�^<1��D�vP�͌J�<�h�Ysj�z�5'<b��0*n�<��͋�����'|�����<���m��C�IT�)Np%8�ɋwh<Y�ڸ`���b4L@68)�F���y"�X�Pe�a�2��.3 ųꙄ�y*
	$�.�	!��Q֜A��Ƚ��'�az�JT={�
�ׇ�7���+�Δ�ybа�8����.��4x��˴�PyR���t��ĔJA"��%AR�<�ӊ\�>�(�G
�> =a��M�<�u�V��Px�p�I����`TGy�i>��<�掝�h�@���M5�LRp'�{�<� ^��r�Ap���R�7f�Q�]�8E{��)���}���Ϟa��L�c���!�# P�(�&�@�z����O!�ęw��;%d�5$k`�{��Ǻ?C!�d(��{A������N
H!��$ �x�sC�:�´�Vh�9!�UVo�����N����1�!�d�*J�:�c��זwu*L�c��2�!��N#� ��%��O����ue�N�!�DҐA��;%	��[R(3�Ꞿk�!�$�H�<�����;1�]`�&)�!��X�^Te��%�O<�M���ѕ!!��J�tt�Gτ~��|�qG	@!�$�g;�I[э�}P�}�U�1�!�8`蜥k�j̦]0(@!��f�!�D۠?3`�d��J,)�g��'Pt!�d�O�n��]��r�#�.�=`!��K�"��+ŬU�vCGd#T�
�';"�$�%�|�DYf�H�'���#%>�� �&M���x�'��걪������+ֿ9�����'
��!K>O�@��C�.#� ����xB��Qج�#Ѩ��Hql�0���y��
�ܼ(�N'QAV�Iu��yR�ߛKM���#���>���+�쇆�y2J�%~Un�@��A�^s�l�r�:��>��O(�s0�S6dD�a ��RE���""O$y��9;,qI��9=p��c�'�!��7lV�]zB����|��1��_u�Ii��(�0�c�))�`3u�M h�E��"O4��mA��lT��߯%:�a�"O�1���즙�en� c@���@"O�((��P9 ��@����q%"O|�Dɕ�F>�k���%{(�B7"O�%���-q�
���j�	h�}Q�"O��s�)^-cEv���α]�t��"Od ����(8t�Z�ϒA_R|�t"OP0#'-e%ZчLܢ[W��e"Oz��t��#3q��)S-E2�"OFa�7-�<U��4)��?8t,�V�	h>�1h��0;��1sD���� �d6�S�''��v�Iq�Ա��}�朇ȓw�X��R�ǐ5J<\���{��!��)@�)���oݰ򡅿A�.(�ȓp@@����T ���#e��A�ȓ}�2����h�*iK��Y�~_�ȇȓ1��d����7k�[�}�,X��7v$`u"��6W� ��'��_�<r�'���Á�T3�����Mp����'���0w�Hp��K��If���'�0��_�AH����ǗJm�܋�'�L���fA1��x��P� �Y��'��1s��;!��j��>���i�'H�-��ā<EP�X�Ïb�J�'�4���'�-jݸ�9� (x��4"�'ϪI"b�����4a���w��٫�'l�~�)�' 	:�%Ǩ�[tE5n� ԛ�'r��XeM�̸,�6������'EָP��R?N$���ku�l�Z�"O�]@�l��sͼU���
���rD"Oؼ����[~"�Q )L�g�Ne��"O�4��M��A��I��>5�!�"O^ �Q�]:5w�tqṽ�;�v8�S"O���&b]Q�V�j�A�M� sS�|��)�3� ��	C�C�L��%pF%��I���!"OF��ЧEI��1�~�>���"O�%�*����]ѵ�Р��D��"Om�ԏ�b�8�c�#� up\8�"Ofq2r䎌vN(<��`�<�"��B�'��:��uBD�#�L T;n��$�7�O��h�tC�f:Z�0b/Ɯņ�_V�U!$�Q������E�mL�d��w���h�B�������
�EbQ��C͜1�H��j�9g(��J�P"O��Y#
A:J̄��@�fi�W"O�y@D@�U�p�rA�&N�X�T�'B�'6+��S�v�X�ZW��3s�Nȱ��'$���tŁ��R',��e$�9z�!�DVO+pɋ�,�G؊�ycNY�F!�$/uD���G�"t���LIk�!�)V� ��&��!�z��jG�X�!�dĽ%�h��&��)S�vY�"H5,�!�O,D�u�`��2l��Ő� Q/:�џ4E�T�;j1�)�G��t�~�ʧe����?q�'	2e�"�A@�aK�gA�z��Y
�'=l(���`���Q����ֵ�	�'�@I5b�&JP&��d�q���Q�'�*��4�ݹ�~���f^�y���'�8\�1l�?W�4��I[
\!���'xz�Q�@_� �RC�� W�؉��'~Ř��^�ǳ�$kA/�^�<Q��V��H��G�	��jS��^�<a�gͨL��!����fT�02��W�<����!`:�%��M�61GRm�C�CW�<I'��|�8A�e'�5q3F��h�Q�<�U$@�L �ݩ�)ʳ/�	ۃNX�<�b �+N��ш�i��2�W�<��):N(��� B.t�܉�&��Ux��GxD'�P��Gɘ<P���*œ��yB�4h�%���D�K��|�S!5�y�b�Bg�PJc��C?�`aC�Z�y���#$��U�޹h�̡	��×�y��H�jF
�j�́�l��  d���y�i[��ꜱ��._�t�"J ��xB�9HP���z�||9��I{��t���ᧂ���r'p�йZc,D���GN�$:9%O�(V	�Ã�+D���p��:`6,�Q�T�� `g)D�Њ�g
a��������k<D�H:���=t�P���^1&��9D����L�u�:t`$�Ȳ\P�Q��K8|OLb���/��/�"�R)P=��H&K4|Ob�ф���G��$��ďoU���O2��k����եB�fwB�R�ˍ6X�
�JfH1D�𪶌^?5u���!k�
��c�/D���rC}��P�f/<����S�.D��а��o=�FjKh΢qKn-D�8�N1.�!���Y�l�(,D��
���Z�4���"x[Bz��)D��i���&�4,��M܏�� ��"D���C�$@�-�W!ږ?��� �,D�)`���Ɖf��po�!�=D���b�Y�F���R�&"Zd�1��(D��z0a��r�[��S�C.�sŦ&D��A1�{��5��E�&E�����"D�XOQ��tCf���H6�	�'�"D������Q��ͦe9Do�A���0=�t��1)>�i��Ԫ�]k�@�z�<� 6y�p�	).~U{�@-)��Y�"Ot}!e�Vj80��N��D�q�|��)[*X�`�dc�$I!FO�yL0B�	�4����V}�<�Վ�	�jC䉻5�	PRM�5V��������C�$9Č���s���T�53)dC�}-��d���`���6C�-�*��͉42�4�4CE�m�`C�	k�����ho�r�ñEH>��D&|��87��[5�5�T��8����ȓ>������r"�8+��GM��=��V]����3�t��pB�,'����&�>MsӬW.A���֥1�����r4��@��R��A�Hx���q��8��>�2��#��l��+6A��x�^�a5�γC3�`Gb�sbd�KE �}�P���*�DC�<1�PY�U�;|JH]�f.��7C�I#<�`�rȚ?�KA�F�*���"O"�ٲ�ײh��xCq��A[�!�"O*����*ɨh���\:Wl��"O�� ���mI�[5׀WF��x�"O�8���WL���K(=rDJ"O ]��˓�#�d����
�g1��J��'�ў"~�e�$2E^}�Ҁ�<�@�1A�P(�y"�O�K��PZwÓ9�����j\/�yB΀� $]��%�=^-Ԕ��)�y���wB&P�B��(�8Y�uƒ%�y�8h�h���P�W�QbE��y�W%QB	��(]I��!#��"�y�2���)�b7@�PX��L��yrL��L���ⱋ>iv��h�E�&�y�U$ܜ�yv�-��&�<��?ɘ'n�i��ዪc>�K7� Or,��'Z��x#l��B�>��n�~2}��'j2 B�d�-uh|*�a�!���'����D�F�m�hG����B�' ����OǪ�v#�<�"�B�'�T�g�Y�/����O� b]�'���(0n�x�Q"E��ma~�k���2�^$��h�#4�8�L�J�j��r"O�#����䩐j��y���S$"O�,C	�J�����E�����'"O��rv�V��p@'�s�l*4V��E{��T�U$+L��I�5h��,Ɛ E{�O���͙.
t;6��{�2��
�'��y-�$0��x`蘰}��	�'��!F�b�&��P��>nvRih�b�'���	�ƙ�X���WJJ���'!D���g�L�ZLa�%�J��I�'j��s��&%��es6�� >�|���hO?��D�:S �0��_�Bٞf��ȓ,p� CB�ɠ��,^.��ȓ@R̭X@DխG�`+�&�ktbmD{�Ot��)v.N&��V�W�u����'ء8��g�8�f�b�#cΐW�<QM��ai�,RW,L%���{�<��`L�i�R`;"gʎV���0t�<�S���B�c	1h�\9�#Fpx�4�'v �7I�0o�,�P�v,I!��k�<12���w�(�ӏU�F�D�
��o���ϓ�dH��~����Lզw�h��ȓCO����Ó:D=y�ʣ|'f,�ȓNr,�q��_��X ���
J�!��S�? �EVOX�0���b ��uv��R"O�X���0��D P��"]�5"O%��͛$#z}�S��9~��%"O�D�Ee�'`Pњ3(	�5u,<'"O��IGm��$�"�� �y	��2�"O��<mTY	1�x��
�"Ob9�D�*^^���c�0�eʂ"O�}���uu̐���C��S�"O�q���ۦF׸e�D��T6\�e�|��)�ME}� חd\��X@�I5�|C�ɔ$��)���:b�!+���p7�C䉟~T��W�.^����n2?��C�� dd��F�K.^d�P֮V��P��F�"�"W�
���(�s�ñs����	/��Y ,�n�x����T�ȓo�H�����N>�͙r�\�(L�i'�|����A�k@"ؚ�9��:��C�!E@|[c��b^h�{�ˋ�Q�x��d'�*�ԋ�*�X]g/�w����0�8H�sd�^�Pb� `�艆ȓ���sj��a����fOH!�ȓq��5���ƧyV�����2a�.���+f��h���R���/!��ȓg�2=�w \*����*8��t�ȓ#��H4 ؗ@֨qQcX�"��-�ȓ#�Ԑ�&iV�{�^�i�M�1q�؆����"JCv�Ε��c�V;^\�ȓ�	y�k��[ޤٹ���,�ȓl4R��GI��8{�E�-ED:��ȓ]m\�Y�J�B����F��ȓf���ԧ�H%�=)Q��M�2��ȓ=�40H�)�/�D!١挌Z�d1�ȓubX�-�!��Ȑ�TT�$م�#�mi�o.lhx�����m}�H�ȓM�^aG���3���xf`���&��ȓ\��bI9�t�b�č86䁇ȓkMܱ1bF٬.w� CJ:JM�e���v�yI�<Od��1�]�	�8��f�P�Hg%� 11��&˖�C�,��ȓR2j̑�l+b<đsHZ|�̆�<�z��#�()���`����1�ȓ<2�H��'�q��e��8p���!`"���(C ��� 8_H�r�)�$ã\ �LZ���L�ـk��yB�ޑm�� �cn��+��	�Њ ��yRfɣ:�*$��B�'V����-�y�C\?g(Pu2b��wȲ\��ϖ��?�'xJ�a��Ht`�!Kȍݴ�@�'����E�8P�E2��ˏ� Y��'}���A�E��`Q�(�:����'��M��I�2n?����[U^U�
�'i�:%��*�de�6(�3�E��'a��Ϗ�?t���vj� �2-��'��M���?^>\;Ueݵ��b�'M8�^!^�FU�'�z�f��'�|�`wEG-8�^�W��w02�B�'h�{��;	窭�d�l�ⴃ�'�.U��̌O�(��˘�4.�	
ϓ�O����N�bÔ��E%�>P����"O�H�5O�x��*4���VGHԃb�	R>yp���-0��f�1�<K��#D�Љ�c̚PM���c�@�p0|<��"D��Q���H�6��k�z6B���-D���D偡icb�� /)I�}���+��w���3� \��Sd�,�0��OW�|~"@��"O�����7��EH㨏�Pq�#�"O�	� J�����%�].Sa���'���C	(c��������B�;D��)��!*�d�q���t?��w*OX$���"Np�6�Y�\�q�`"O�0�� +���!�O�Ty��c�"O���V �o3u�7��Dy�Dr�*O(]A��9dj҂�	6���
�'��0"%�[=Νx�1;Y0�2�'���Y����k-8M��Mŷ<a���'�8�x�m�<��D�l�5�@\�ʓWT��@�x���Gƒ���]�ȓh�����&=�ru/�<t��ȓs���s��fh���>�i��QA�AY7.����E�â]�m=.Ԅ�/�kD(E�?��a��e�/��-��s�e`�ƞ��j���j�-i��ȓB��S"!	�,�����G�>?o~���09°�1t�6,���ضu�V��ȓ�v�*"�L�E�ZEɷ�]����ȓE��� �%��O&4��E$@0�����M�Ly�m	�	�
)�`��s̀��"4��2 [��t��1͍�b��ȓKĵb���qA��ѤkUF���W+��x�*
$ު��ݞVw�A��@�LQ�$�
8Cԍ�Y}���"O���J�V��	��
(2^�q@"O�󡭝+}>h�VN�>�H���"Op�!��N �@���,Y",��11�"O,e{�&�X#���JڵS�T�a1�'��Ih�r���#W�����8��C�	�"�����"tk>����K/��C�
7,�Y�R�-�
�Xf^�E�rC�I5l�(��J;�5��'^C�	5s���`�
[~eȂC˖PBC��.]��i���%}�H�	u�DMZ\B�8-*&�P�*�^�0��^^��=�'sZN�@
J9xeBL`��C6N����Qw(4���یGB���2NO��찆ȓs��0s-Y�8�� ��dG4N�ч�J�4��D\ ~8�g����-�ȓ$�밀�^p2��Ѓ���ȓNZڼ�@iܢ~�����]^�5��!뾍j']�-��{cS�*5��G�0�EB�(���ҶM�/7ՀT��Mk����/��;Kɹ$�� {��І�}=�����0Z�K�>����/C�$9s�^���Qᡄ�<UOf`��ph`�`�Ğa�yQ#�Y�� �'kB�X�d�$&���[�`H�j^���'�){�	�RBBa�nޅg���x�'+��B)ˤO�LТ���a+z	�'S:|  %á=�Z�A�W�V`�P�'�Fy�ӝ>��M� ���"O��B��b�:h"N�-�B�z "O`4q��q*�u  gƯ)�Y��"O�ca�L�g��0�֣J�.k�"O^���E8~��Cf �N�4�G"OR�ٱ/B�H<5zQg�8UJ�)�"Of�!�9<�|�:#�٘D�)؂"O��z����ٲ�A>�X��"O�mcl�{x�R��ع`�p*3"O�T�gղF�pm;�O�<�p��',!�� ���s�הq�Za)7�vT� C2"O �H�(/��%�F �|,3�"O��" 
d�K��O�b�����"O@`�q�%CsZ!6c��it�x!�"O
�����-<�QD�?XevtR�"O�M� c�!H6N��V
�7S:��T��D{��iý@���$$�0BH�ԃK�<W!���-���A�'6>?.����B�!�V4������$19L�|�!�D�	�8�v���+۲H ֪�+c�!��ܲ�jfF� s�@�����}!�΅* ��+Ti�â��@.x!��V�[��Q�pWk�%[!�Dׄ	�N}-���SN=&ۼa
�'�y��O�/
S�֬��	�'���G����@ҋ�Bl�
	�'O�\
4n�=0�iP�@�Uc�'���BÌ$�|T��(��0|`P��'ƺ8���;BP8�bT�#f:qP�'29�F�$[��:ٙf�B��
�'�ʤ�&#Շo@�� ZJ���
�'�L ���
��m��-NZ���9
�'����D.Ո(����� )��ib	�'na*4�3���s��kD��r�'Nذ�I�f�܁��KYOi��']\%2ҵj�*�{�)� �=��'5li��
�Z6����ޏA���q�'����Q$�,D2��'n�.��ݓ���/�z�!��@)P����1`�0�1�"O�A�%��<߼ ��@�W��$��"OX�9�݉Ϙ
я�7 �n��4"O��������z��`�"O8����6_<\�b�@پ���"O�,1`���*t�xt�C�`�!�"O0Y���=$��A�V#W�*��Ֆ|�P����K�
|2'MW�E�0sfJר84bʓ�0?) �5u��brj�3��8j�B	I�<�t���5��0�b�/9E䔰%�	L�<�*L�w�А��i��IX�V"\E�<�$N]�l��q��+O�
����^@�<���Q�d�:l˜}l숓&@�s��UyB�ONx`E؉W�Ȥ@��2hI�qsN>q
�'o(�0!�`*}��\�V/�I�'�a~bM�'�����A
-A楒En��hO"����\0���wo�� M�����$�!�䁔k��8[P��6)E(@���U6�!��0v�"���|>Z�� �{}Ȇ������/�fgإ�#�A+?
`I�ȓ<o@��b�u��@a��]#<:�t%���I�xV���iI�ZD� ��S>~B�ɯF�t0@D��7v�����N�g�>B䉼E�-A׍b�q���
��<B��e\`�s�˶a��Ҁb�7d�B�I�<7��Y�aX���Q�Z�C�	�X8��ӡC�\���6B��"��C�I_���%�B�de�[s�ԗZ�C�	OCL�B%W�(��R2M�,C��;@�X� ��i���[�-R�p��C�	�& `��指]Fe;Ŭ�[]hC�	W[�԰բ��+��k�B�)"�B䉀D�x`fϗ!�� ��=��C�q��I��Q-Pΰ����v\�B�	-[yx-�3��/>�e���ڤPoJB�	�a�,�M[♃U�Y�#$�Ox��� ��遊�
?���[�H"Τ�1��'�ў"~BC6,����O)��M���ͦ�y2-Q�b޸����M)X�@�Z�M��y���1qs`<��M��S@B�b!�\�y�%��lɀ �Ս�"I���ѧ�ݥ�y2Cw>X��썊Bڼ����
�yR�]�W�*���䎭?��Hg�=�?��R�ӫvhT��v̺@���y���3Y��i��	u�'r&0X@HJ�g�t8q���g�*5��'}*U���)S�%K�D߷^����
�'"�-�2�\O��p��N�O�=1
�'��Qm���	Q�B�K��8�*O:�=E�@ǫn�\�� Ƈ_���+����'�az"N@1�,�p3C���p����yR�D�M�:�I�3p�v@��y"D�;L��J��Q�}�h���ۙ�y򂌅nRą�t4	4m��y�E��5��y�+�:[*
��3����y���a� ���F�L���G�y�*�9\����!���ad���y��&�T@�(��/��ۢ-����?Q�'E�����^��!A��S6�����'���@�N�_7����a%� ���'�@�j�1U=�����>g��
�'�4A�Dg�G�1G�H�
d�b
�'P��SfI	!�&u�Q"��O_�T�	�'pe#1gV��)�G��Hr�9)	�'J����H�y���<����'	>B&(0 *�<�AC�)HFa�'ạ9�¤8v�|Ia�J3/�%S�'�-g �2���P�*��O���'2jl��W�$���g5���8�'
b��N6	���ǁ��*�z���'��9��H�-f8ef,X�8�lh�' b1��L.�����ҵ,%t��
�'���ӱ��,�r()R��+8<�J>���E�d#E�_�h�F��EG��'�T�d.�t�eE%c~�26��.��(D����霴x %A9���f$'D�����OK���G�
)�p	�c�#D���ӡ�J�Wb˂u,%��"D���3�#X�rɑ5)�LQ�p��4�O��!�bS�=� ��E"�/y�9��IX~"&�`�\@p.[&H&I	�y�hR)l����"�	-$+^�����$�y(ߙ��X[�*T#{� ��iB��y�b�>U\!�A�ɟ��4IDǆ��yBB8��m�u�@&uh�A
$���y�L�
� �y2�܉lք�bۭ��<A��$A�a��蓨�8��ke$J!>!��7IZD��%�)P��1tID!�D4u۾Q�mX)�,�Ѩ�;!�_!��[����UB�m?H�!�$ҥ@M���M�{��%/{�!�d�4Ra^@��m��(�ȡ�S���}!��L1g2�Qf��bN��3�+ܭ(�!��L(CG��#@�D�o�< &+W9�!���D�S�θ2��h�J�2;�!�
�Qf\!��^b���C#ǉ�!�DӘ-��%��*.] �{�oN�]!���B@���'�N$;�r���7*!�D��F�pb�	�g�*���B80�!�$*抉`�����|B�K,�{R�|B���qY�]"9�F��3��{+ўd��3� ��3�/X,Fuv���h�.�t��"O���q�
v^����cꎬ�C"O��J�� E��Y��Z� px�"O�Ik'ŏ�b�����1&�ҭ2"O�pg"�'a:8�b���1}�´��"O�9h�N�8g�^�i$�Һ��CB�'�ў"~Zw����љ@�	&7Yz�хi5�y��Oo��4c�:*h�m�&�7�y2%®��`J�<5Kޑsԭ���yBd�h��%t���x8�3/��y��v���P���V�H�B����y�8$����甪P0$�`�	 ��=��y�+�+?z:��+��BԾ91ѧ��y2�F'h�� ����<�[��(��>��Ob��H�oRrњ`"J�����g"O"e��c�x��c�5w��a"O޹��j��.<07�N�"��-x�"O"�%��h xb�0l�n�A�"O�L�3�0s��Q{V�l���i�`�'�a��D��)���%Úma���t"ʜ�yr�S:��Q�wo�k��"��I��yR�BM���f
�]�&�`'��y�� ��� �^�L���������y$�5GRD@��E�Da�UE��y2�P2~�d���Ӓ7�vY�E�Q��y��"��J����(,#��)�䓣hOq�%�����A�2Q`�1;�5��U����	1\N��p��M!5t�y٧ǐ'qQBB�	�[ZVq���иr�ʈ ֎NPJB�	Wޑ0DҬ6ޒD�G��[��B�	�e(ģ�N�������?<B�B�ɣQ$����b͟l��$Sw�I>VՊB䉸F_$��bY%Iu������u2tB�ɪ>}��eh�/;Uz���j��j�`�O��D?�6���k�L�e�c!��_+gT�� ���8?<���I�!��/�${ �K�_�Hp�q�!���)ٕ#r*(X�j�((v��t"O`p
!"�J&J ����&��+�"O�xp2��cF^�bOb���Y�\��՟h�?�}2e`��3ݰeK�M.�}Qa!�k�IZ�����y�[� X�70�S3E�4�y�H;i�H����.8*�}�@ �yR%�:6�r�[3ň(+�"r@���y�/� b*��̌�.l�����yҬ'`tV�L�-#�hGNL9�y"�!>����.E�2Dn`3G�1r!�$�c�	j�Y�6G�d��ΣB�!�P��wa�xQE�*"k}!�\4=�h�C�ܱv?ZXӂ�8l!�D�r,�"&�;n"��	_!�d�{H�$�R�>TxQ� 'oW!�dX������.1[~d��n7h!�$�*k�2<�7�U��x���ӭ%Q!�Q!6C�QD��M������}2!��:l�d�'��5r@��2�V!���)q0��4dǎpj�9r���-n!�$��O銙���|O����oR w�!�DF�d�N���ק2����j�!�d�+1\�Q�T��n�Q���.w]!�d�9HA0�(@e@�R����哪pX!���ò����H�MH:dϻ"�!�$ѭ*���a%����a����?�!��
�{^XiS�@
���r#7Xp!�� �=��N�^	���Tm�8�,��"OPmp�&Gxh��b%�Y���J�"O�mK�@܅w)f\ s�I�t�j��"O읠��71m&��G�88{\9hs"O��`m��f;؀k��( \l
"O(HA�-F�Y$\ᖪU1`AvBt"O�`q��#�`3ǈ^ x���jS"O>�KROРd��/�b}Z6G@�.!�:A�,�Ɉ81�O�f�!��:��0q�"�7d�	ǀC�	�*����M��05�-hC�I�^F���e�
f��ꔅٻSS�C�I�^������)�����G�f\lC�	�9Q����u�Y�� [�@C�ɰy�!�+-^���S4nR�e�C�	�ZՊ���#��戱��*eƴC��C�"�g_=T��zR�_��NB��n�PE!�G[�n�z����JB�ɠU:8)Ȁ"��Z����2,D.��B�ɐU��	H����s��d�4덐�C��a`����H.N���HBC��,K�2�F�U8`h���R�C�b#�(�̗�s�䁑�mѽw�0C䉛�� �7������� �z��B�v�1wB��6�X��� S5ŪB�	>M*���p��M� ���i�%j��B�:!?̂�ęA�,u��Ǌ�C�ɰy,�5*6hËB0m ���PI�B�I��!���U���%P�O�:��B�27�Da��#�[�d�h0mP�z}�B��+K�����[�R�rP���8 �B����4EFF��LYӇ
4%�B�ɿZ(���B*����ƥq�rB�	�s�~��& ܟ2AFu���^�M�fB�1"�d1z��ޓ0ze��.��B��/@������"x���W�f�B�q*��bլ�<|�9k%�2so�C�I�/��;�)U,v�Ѫ���_<�C�I�bd�r��*uS��B'_�NC�I=UD�c�)Z37���7�ޅ�ZB�I�#���jTI�=��T�e`[=،B䉧a�����E�detܲ�i�$�bB�I;�m�Peӌh�  ���E�6B�I6���A��1G���C�ʸJ�TC�I#a(h��u�R�}�>D��ǅ[�fC�ɨ)�H$�":�����!�C�	�"iԭ�&�7c�N'_���C��&x�^A4�͔y���@Ϣ~/zC䉖5��tK7��	��M"PB�B�,R���5 Gu �<�'��(V;0B䉀:��#�ZFy���Y�kg B��6 耀�CƇ.� �@�ڷe�B�I ^�D����)^#��hV�� {�B�	#�t �$̈�+j�HR$�6U3B�	�Cn�y�LO
GR���N�>=2FB�	�U�)`e ��\�a�P�^�u��B�I�u 2��^��x�Z�̝� ��B䉁fR�lq郴��YE��Q��B�Ɋ
1�̊�i�����Q�`[�C�	� �z��mG�Y����i%2��B�ɟ����A����,�$	5|�B�	�e�����FϤĹf(_�{g�B� N���Q@������ uEBB�I �.��&O�%����2�� 9�
B�)� ���ϭ�Pಯ[�B$�5"O�ɲP�+wp�<ږA����yK�"O4���E�2r�	I ���dC��'"O��9�'^'��ˀn�:{^�]re"O��	��M"Y�m�
�4\嶵k�"O�a'!R�l�0 B���mZ$"O4��)֊^��9�(Vl���"O��zS��u�X�ѣ�M�A�T�:�"O<�s�hR*)���Æ��!'D,`"O��0�O�*�uq����uf�� "O>�lZ/*<� V���"�"Ol���jM�T �P1�V�$"Oڭۢ˚�z�0�H�nI0�V�8�"O�$ r��sҒ�ِn�_r��3"O|X�A�(G�����^�����y�gCCr&U�ҥ̑o"`�����y"�L&(S^��R���fPJ�����0�y" Ġq����Ae�\3f�8q����y"fT7`�¤@�L[_��7�^��yh�
�`׍.�����N��y����(ÂH�fr���2|��mh�'Ƥ	P%L	<݌���]"r[����'a����f� Z&����dP�pdx��'�jA��A�錙��$uB����'M6���Ə�@0Q�� �#�t��'� @�.�5�}J�GɐN�ؽ�
�'L>A��U;BBtbp���v	49
�'��
!�ӧn ~Dl
�'�@�ڣ-��>�������z�= 	�'��a��
"y�蕊Я˥B�pdS�'��`���O�q���&���&F��'.$����M� � �G�$D"���'����	9�J�y�m�	��"�'TDy���O�!�OU����'����cĝ:C��LHG����	�'�0���ߍX�ɩ�k�r?jP��'N"�'U�.<�Ыk�	;�4���'��2���E��dbR,� .��1)�'Z�i�`�RF>��­ �'\bA*�'����f �d���q�\�����'�tB&ńwf�ʢ����2�'^VDX��݌Z�l����2�*�`	�'Dę��ᖎ��1!�Up�ݪ�'�L���C�X8�&l�Hi�	�',*%�g��1���sI?8�<1Q�'�6�*���%/�y��ʯ<��Q�
�'<t�$�� J���<�.P�
�'Z� B�63��*��vV�S�'�t@���H6aF�}ؑ��=�����'ΖhÖ�ڠu��-r���@)�'��(�@�Âp"�J���f���'���ʝ�'��{�:6�0M2�'S��*���`�"�blT?,����'Q��zU�U�7���8��0s�I;�'ޮ}�Ǆ�>l����ʯ'>a�
�'y� b���2A�Vp�v.L#Cf��'��)��@iI`�-���Q�'����D����"�B�X���`	�'�4�2�H^��;AeW�O)����'�N�#❦\��1���Z<$I#�'|NI�IX�]z��b�(Gt6�1�'c�t����By�LjA�M�=�|T�'��iڢN@� (���Ȓ3���Y�'��X1Ǩ����	�A���D��
��� ����aY05C�f���x4"O����w^B�+Pa�&  ��"Ob���
W�@��A�� }��)r�"O�`�%LUgE(��G�ӆ>��� "O��3��G��"\kE�&E��4��"O����Ȳw�P�����\�@(�%"O>�Yjނdg\@q���4}��!٦"OZ��/�9@��X����t"O��i]R������=���"E"O�H
��3*�̙p%�#U� Hx"OT|h�,�� �X	���Cɀ��\��F{���-ph��U&�!��T��2-�!�DV^u2�1#H�>�L0p�@@#�!���s�&�;f��f�L�%/�{�!���x� (��H�o�����Nĭ!���q�$9}J|�':@4�g@�������p�(��'�J ɒ�8O��t��G��c�6���4���A��@��!�?�xh3�LJ�",jL:D�,�A�Yʈ��an%d����c6D��C"��o:����Z,)�ps��>D�X1�؍cW(�"�Y;O ����0D�����][NT��m@hh�Ь�<�
��v�p��Z?�$�;��S>\qJ�G���h�6az���(C �[�H^5;�~C��4c,��%4��l��!�?5]R��ē���S�,fչ�#8 v@��`��m"C���q�CH�9a>*�s�b�@�DB�	?u` jE6_1
���C&�.B�'Z�D�T���m��щ��BdT0����h�t�>%?�"ǍA�>�ҽؐiZ�{+D�U�<�O��'v
�W�� <p����J6-�d���'�Pt��/`n�8���E5�L\���d8�'~����'�
G�	@Rc)�|��ȓ_�1��7n�4��IF�A��܆�,�©����~L�%z�`_G䍆ȓ��ȑ"��p
���c♄ȓb�e�p*�%&��f�Gd&0�ȓol�ͱ��J
t� j�KϹ���c��?,Oڬ���X�!8aU(A8vԴ�b�"O�,`"*�,�2�b! �1h�!�K�_�<�Q�Q�=OL|S�+]h�ў|��ӄ�zt��e�	fГ�DʀC䉱8'��+��F��*@BF�r�T��?�{R�	�'7�ppRN=�0<�0��%	BC� {Q�x8��g�܍�DZ�L���n�a}��G5{x*�B�#��X���<�K�ؖ'Z8�˶��(��TO����c�@��y2ʉ�������@�  ��(ިO0"�d@�0��0��"Kr��p���e�<�Q.ؐ\{��b�"Xs��h��W�<�bJ�()X0(q0,�4��X�SR�<y��	�V�f��J�T�Q�C�v�<i�ȗ5$��!�e�!�0%��aSo�<yt�ٮ�v���X�q�J�:b.�l�<��� � ��I�i�����h�N�<i���,2r]�tC߷5Ah�����t�<�����L�2���_ͼ�%fKX}"�)�'4Z����*���
�f�!,	����[t0�z�鉌0[de2�ě�r�u�=Yۓ{=\Z�j�"j@�3�ĕ�)���M���R:I�#�	ǧn�q"/�~�<�����B��N`H,��@�$0�Շ�K�`�Ѱ�)kp���m�.*3Ь��	\�'�8$���J�^(���
X�j%8�O�-�O� A@��!@�*P�RDȥO
�43O���J�S�Ov،�Q8��#5�6v%����'����B�7$�$����v=*�(OJ��$HQ�b>�@�ݣ!*���`�8ud��<�O�`�'W@����/YV	)%�	2���;��yy��'}x ��Z+.}9�`�x��Y�¼i[���O���H��)��u�׫�w@��z�'$�$����5$�1Ȧ"�@�"@�,�(O?�$�/�Ɂ
H�
{fY����?!���g0ڨ1�@<i8��Cʻ)���=O�i��&?�"ƣL��U"O~�@����EM�5)"�M��9�$�O���o�g?I�.ǲgB�������T��8���9�y���2Ҋ�`0(G�NZ �	7`#��$�<�H>���ɬl�d�y�G�KBPDsc�r�C�	r�e�EǗ�l� ����
ѧ�ē�p>�'�
SK�d�Q�P�C�ƞu8��$��'njI��d�%�f�I�^e{`�m�<yT'�(Qgx�"'+2Ƹ<����h�'� �F�4���3�h���`�N x�E(���yrÀ8�L�z���8S���m,�y��Va�T|�Ѡ'Q
���u����y�kX�/��i�̑#NA%��6��D.�OX�VZ<f�. ������P��'��	� ?>�B�+	d8��`�⎧�rC�	#Zb�ѳ�B�9(�����F�0"=���T?=s�B<Q����(}���P��"��F���'*JV]�U�#m�ƅx����( �H���F{r䐋`�Ё�'��=6+��ɥ
��HO��$�MSmX3E\�_�q�U �#,�!��hT+�H��{p�pwOX$��hD�ԩ+}!��zU�	 �b�ZG�S2�yr�B�PV6��c[(�Vl��A�y�l� %D��#ӌ8"X���O��ybJR�$
�9,�&���V����%�O� �\�O�h$3D�L�
i*�Hc"O���Ξ�G5 �����,t_x���"O�D��͝<]f�R�o�>1�R��"O�%���A�m12o��`08a�'Y��OLԨTM̕kJ��!N__��@�"O���'bD$s�tS��D�(f�s"O �r%�53��1ɖ�H)f$��"O�)b�	� |�`�P�u`��X�"O��{�$�
H�b��a�à2?v%Ӈ"O���	��gi�ۅő�mB�8���s����j�E�4�D�CR��sC�m!��M�oj�b�rY� pW⇤�!�Z$��Ձ߭@���p@ԡ~�a}ҕ>�E(�I�
�(�o^�h�s����?�/O����(l�x��/16�d�r��:]�!�DWPC.��#-h(��֪N�D&!�$�v���ۃ��\�"]�	��IhX��&
Y&�P<� ��j\���e+!D��Q�O@jA�pF#>-R�{�h)D�sugM8�lR�˄;&�h�H$4��C#�,U�����S�p�lC�h
E�<�¥�B n���$�>A�5#Cc�~x�TExB-\&U�͎�&*�,Z!����y�V�c�MX�Q5j��mS��y�� 8�9b�\�,? =�����xr�ii�i���߻>��mc��I1&X�6Y������'�v�>�w�ۉP�	�B�гP�@����'LO��#zyr��L�19�`*`@U�:!�'t����	�?��xJ�ܳ$��,S ���D{J~� �����{���W�ΌN��H��"O��p��� ��A�-�TyV�R��	}�'��ɳD��5@5H!Q�dis �N;�B�	�g�V	B������,�%h�B��rI�]#��N1)/X4�+�.d�B�w8�Y	�A�e�L,��F�X"C�ɉT/��Z�M�E,��j��"<q?�S���Y�IP���gR!P����T"���yR�F;/v|`�Z�_�*��7�=�y��)�	z�����X�Q�U[b[0��ȓK69!p�"��!�s��M��%��R����R��$�^�� �*a~�W�P���7
�xth�l+d`�c$D�L���:B��h�G��2��5S�$0��{���';wҥ:U
S	\zp0�"�:��ȓ6��4`�d֜\[��-��'����J������p}��;� O�"��w���1eU$f%4�Cר�J<���ȓ1p�D�5���+��%;:�B&"OI�e*
(7���$υW&��#�"O�8"S�&��р�0A����u�6D�X8��%U��PR7��I���S	5D�,r�J>"*  e���礜o3D��u�B�t]�,ID
<#*f cqa,D���WN6����U��/T@F$y�+,D�<d��)V���*uC��u��ɦe(D�`Z�I�
&@��5�m޵+�h'D��
T�R�_��)#C��3������$D����H�0uziƃ^_��Q�3�$D�Da�*I �H�2f�F�{�~m�B%"D��xE��C��qD�@C���Q�:D�����	B�|3v�
���Y��8D�c����%j��҄:h�A�$6D���� ��(QhU�w 5E�� �5D�����X��NF�`iz���'D�ԛ�&�6d���9���j+ qj J8D����F�agJ�ԫ�]���Ja)8D�����Wak���I��7D��sv�L�y�| �_#Dt�"�M6D�|�ԍ�0*�v��ě�Ql���63D���%̞ R���vE�9a�@���1D���w�� k�`��f@W*3��,�'1D�Ȫ1/J!�q�2�Ӡ}w����3D�PqQ��$S���x�+�-Zo�0c�,7D�����<V�Pi0��d<�dF #D��(��]�!��3��x:Jx !D���w��8�LR��9����<~�`�p
��]�#
 LOt��6MB/t2���I�� 	Z�BT"O��* ��2 �ɴo`x�"OEp-P�R��@�l{^���"Of�J�-ѽ�Z�CT[�[�i��"O��b("��Jc�_&P+qkP"O�Ջ��V3_�c���z3"O�`�n�o��U��d�7��8`"O�p{��@'H��́hy�؉"O����(>$���ϐ�F�$ڑ"O�i��W):�3�O\�1�6���"Ol�C��"K�q�7nJ�
���"O�ɐ��U�2QP���D�$��6"ObP�gL�u���3NBxvv0�a"O��c65"��Ȋ�PTy��"O�0V,$A���Q��=^^nĲC"O*M�匯Q��Y'�VATq��"O����X�b�jhQ@$�,X�l��"O� ~�ۥ`ƘF��a��	4$`��E"O�؃�?zt�t�6�D0@�"O�4��R�a�2!8�T�}�@�R"O�D��H� ����S�C��$q"O┐���i���K��Ǔ/ߠ��#"O�J3"�3Bhl��Rn��n�"p�"O��p�O�Y��ã �>&�Źp"O4�r��Xy-�I��6;�P�"On �e�N7k^e{`ΡO'xXK"O��DB��:�Pggø0K��S�"OB��r��H H;�L�+�J�"ON�� -"אm�b����*U��"O�@2W��gT)3PԳH_�}	�"Or��D��5�J`�5
�+f9"`�"O|��p�ɒA�<�P�V�W<lX�"O,�	]���l�1�s&��p"O$%�(S�k�ҹ�MZ�ic�0�"Opm��Y\�;��S7o�h(�"O����A����"G)�)~y���"O.Uڶ�m.�����g��E"O.����Z�k��X�2F�N�h��"O��`��3�d����Η9�b4c�"O�U�0*K��\8Q�dI�A�,���"O>��F�*kDڱ � �:YxhM�V"O��iạ̇̄
�"���ܴfh��a�"O^U���%4�ᆛ�[Z�Rt"O���&�g$� s���R�$�{"O>5�&&} hu��L,2�j�`'"O�����X��U���G����$"O\X�6�zW�-�R�P[�"%�b"O��C�M��1O,�
�I y���S�"O��EFN�$��&FPT�x��T"Of����M/��c��0�H�Q�"Ox�4nƧc�¸�C��8�l��@"O��� �U�"�@$����B�:1"O���n&F�h�h�>v�朲�"Oܙa��9z�0$�g�X*�	@"O4E	��L#�6aY��T:Eʶ"O���KȨ[Ѩ��3��m\��v"O�xh$�'K�(�+f�R���"O,��a��F����(9<��0"O�m�S�
-Me� #2#(��U"O��
�ER�x @�Ԗ�7퉠�@q���S��!D�](x*Z5���/+��B�	5md�%	bn;���i��P�f�!�`̡��0}���'�`X2,B�\-��J��[��U�'�
�+�n�<d�@\Y�f֛d�*�+�"�B�[��ĔWm`�YV�",O-���m��H[�.������'*m�ECW~� r�CĚh��x�ǐ�y���O��TԠ��
O�ة��˽E�qy���8����T�dD�)�2yGη,�8��-�S�sx�I��:A��[��6=HB�	��r�U��]j�SFH�,u{�q�G]��ðֹd��Z�'���v�M~n���&�ѿ]>1���^�,��UKw�Sz�<!�ތs�Z��4�)ADp`����:R���0w�J��Z��7Il�oڽ℩�)S]ܓ"�P�pT��%|�@:c!�,nz����I�c*��F��8��=YB�"��s�`P�h)� *|�5��a�WL88Eo#�����tJ��j��H8O8W�1OJ4:B��S�
 g� �Z�J�����#�D,�9`���	WqFLI#�@�XD�0��<�!�F=Z�&����Qe���a��{�n��u��+m��IՆOcf�JG>\�2��!�?��3�t���$Y�CC�PeeK�~P���-2D����(4~Æ)*���)\���a��(��t�g�##��I�t�ő�5zɐZ`b/�I�bPf�"3n�\�n�HE�����L�<t��!#�'d�+��]��8���N�3n
�y�"��*�b�����`C&љA#��	ӓP�X��&�	U7Vu���[
��'�j��DA��v�A�
v΀s�J�+O:�T�P� PH�u�	����reV�!s�4"O�D���K�o�$��sN�
az&1[��H'Z#�Ę	��=��8����g�X���n��d�b}(-k�1�l�́{�А�!�x R��'��t�Q�R��E�oάn�>��掟��]`E��+����6�n���ѡ�i�A� �^�_�qO�������u�!V8s���J��n�'��-��/��]�؉��j��<�����	̞�\�(�IBL��ٻ)�7&���i��'� �n=�p=11��0w�(M���C�b5�d"�BlyM�
є��ɪ�\䫕�\�H�vh��O����@kĽ^��j�v�N���L�$�IS"ON�s�;i:�V�Ѵ8����#T=3p�K�fӍb�Y�S�ً_>D�o"u�p��[�����/�yG,,���A1+��Hn�h�Ǣ���?� �	)cj!�N���@}���ӑ
%��(�旰��#q�7J):�@�j� �P��3�Ji���|��2��!9B�S+E�n9;'ϐ��O�ز�ȼL��Ŭ\�=@�u�P�̝u���{!)�-59q	f%�2;���H4b���ʲ(����Ĕp�Q��N��bc�`@eO��2��(Z�����Q85$\}��IL#��"I�*$�x�㑰J.�tfH�N�t���wh<���0df��x�.ǌO>��

F�'�Zu�& Ԝc��D{?�`�+)�	�sCv(����+q9@T�B(�.$!���}���R(R�O]H�'K'_L�7��(�:-Ä�d�p��<AǤ�n_H����j��]�M�d�<���]8.@���N{�0y��:@
���%���R��M���<c�� 5����4,�UZ�4����v���1)��-A<�!M�30�l�JQkB�g�N���b=�"��64�|�R.Hl���!���%�x%��,�I�x�ɩ��wF�xC�-��M��Ii萺G����@�8O��B�	�r|�5�˘t	�|Ȇ"M����J�A=]��G�B�$���(��I5 ���	�aO�IJv�Ih��C䉺o��6f´-ٖ�
C�
�$�����J��ji>|�2��1��z���)��)�E�Ȁf$DX�p�H��p=) ��\> SrLܢ�M;Wl�>��PFF)x;�	�V��v�<9![�ݨ!r�(Ӡ|�:�Ӷq�N�����l�i0|G����6~��ڂ%�8��[�ٶ�y2I����q�I�(n�^�iG���x9�!�]$���'�>�I,�����N�_�t�q��{�C�_�L�'���~YhP׬Y����D.y��|A�K��=�d�k����ɐ��do���0>� �^�^$��*dJ`�¾kM(�r�GZɖ%��Z���$!V4K � � ��N�QDy�	�[� �F�t��#`�L+S!^�FN���ȹ�y"O˿|@1��9H��xiq���y�E�E(n�j\��m���y�嘗bW��*㋃�Mf
�k�)��y������c�E�,�H���f֭�yBm��K��|�`('5V��h� �y��̀~2VD1��?#�@r�]����'C�r��K1B�4 ��m��L>�S,թN�$�IV|=)g!g<�s���;tP(�U�yB\�*�◂E�"p�C�G �R��D�.p-v!PϓEn衔�e��(��\�E��U��ԣv5�CƁ�j�!��U�^|ظЂC�
�]�w�^H<����?���(�OL�f�\��3l�Dy�#�>5�E2Q&O�a��A��5q=��~zDM�5 ]& cI'k��P���G�<��*���Lx&H�#e�2��C�����0nχa��-Rvi�
:h�h&?1zV�x�Ѫl�X�wfP�%��j ����?ك�Q���=�ɸ�NɩN��<A��$R�Zh�@l��螀���A��@���~e@9yD`-q�V*��U�^ >�?���W���;�(M<T�t��4 ޛS�M9�
�p6i��k�6{����&�1$�̋b���:�[��BqЉ��<��]&o���.�,_��x�G`½��c?�$�D�$����%CL޵��.4D��yw�S�+6$�	��W�Pc��$-�tA4]��Bs~t�+U&��CԌ��~�#M<Y%�L�X�� *1�SQ�б:Q+�m<QhB{.�J'�������9oC&�
�g(vw�p1JM�#L���m���
�EÒ����@���IIz4���_qD�
ۮ=�4��!R�A}��� ��U�ޑ10"Oȍ��B" /�L	�eQ3f.)�"O.@0�Ϙ��bd[U#I�li�@�E"O� f����׆1��+�W�U�c5"O�Q[6l�"#�a�n��C\t�rw�'Y��ˁ����ɵz�$����}˲��d�	�6C�ɴ3��r����S�*=@�)O$L`�b�8P���Ne�\+��S)p��a`P�_7�ҁB�&�BB��=�6����
t7���b*:d�K`�S=���e��!��L����������ا,�\@���/4���U�U�)�B�zo�uN�^L��1"�)�6a��D���f�$~dڠ��̓&_���M�}n�L�%Z��	�>��1/W�؂$�vO(h�B�Ie�*pZī��8p�O:J邏O�,HG!�9L༽i�"�f���Q��R< ��t!Z�+�Xm��g+R�jQ���B�|`Ȉ���v�T��B��'< D��>�gϟ+e�Q9B�N_��� �`h<a5$���<�+���,8���@�-TG^)�Ў���T��
�{4��s�ٯD��H�AɅ�z�牯E��T�w�	��~�ΓGk
�B3�0\��д���S�"Oȵ�#AY�t� �A*(�R�	���**�X�!� ����
ܩ��Bjx��ɀQc��
�'�Tx�fW?i��!�	X�fv.t��oDr�O,|��Y�4#7�Ͷeݾ4�5��&9:��!D�\�'�H|@��)��'8���C:D����|m�Z��ț �����9D��(�@/`�z%k��P�yP�0�E D��#f+O�?��ip�ѳ2 (D�V�!D��ÕJ�*�8����"�H��+?D���B*�1dn���C�ub�y�6�=D���`F4[d��Pc�
���p�<D�$�F�R!Z,ڥ�4�F=1,RPZ7,)D����-�N�� ��!T��3�	'D��bSK�n��  ��<K���$D�<���:A�J<(�ȑ)_`����m1T�P�t�"�d��F� Z���"OΩp$B�(g����x���"O�XqeN9]5�Eq C������"O@�8U�(q[xm�_9(�� #"O�$[�B�7?��01v$W@��Piv"O���f��	9kzy���O�x��"Od��#��a`Ri�b�;N��uqW"OH��#dJ$u̰S�R
�
9h�"O��!�R�q�,x���La�� �`"O����ę%Ot �d^�E��U�W"OV��$�4�r���Y�BK׌6�!��,�4*V*�*U�Z�Re�+�!�dk����D٩�6liG�A�h!�d��L����q���h�pp*�"λg�!�$ķLt�P����{��5 �=	�!�D\�tnB�A�:L3��ZN��!�D�5q�Z���ݯ 5���EN�R�!�䋺	̠XJU�J�d2�y����b�!򄍼G&yZEN֥B2D�o�e!�D�s�y�*�/w���YA���h)!��ΌX����ŏ�LA�]�U��!D���g�Ɩ7���^�t�2��U/z!�dߝCK��i�)�<�hm�č��!��v�1�$g/U�̐U%V�|�!�d�2dCD@���	,e\rhr�KA+�!�DC�J�J��ɪ[Db�2S
E	�!�d��9����V�JHr��c��]�!����Hf�$.I������+�!�V�b��R���\"Hx��iJ�k!�$��rY�QI0/���(C/H!�,sπ�)�@E(M������,n!�B]}�E���xZ�Y)���b�!�� &qS��̸��� $�<Ŏq�s"O=phρc}bU��A3m,m��"O �f�&*�}��)Bl�1�"O 1��LT`�t�5l�J4�%"O�x�*P�X��]"�b��I�Ř�"O0��b�X�eX�9c�Z
�lt��"O"���Ŭ&��B��T��9��"Ot��7.�p��X�I
~pp\Y"O"Y���ʒv�(��!� q��q"Or�J e�3z7��V��Ujx�j"O:��4.��a��<�b�ŭ0���"O���L�A�$S��CV�!a"O�AbZ-PX82W�S�J�ؼF"O�2p��n̻�
�1�| �"O\�9aꎩd�`����
��)"OX��ɏ�{M�ZA��;���P�"O�`�f�LC�1�Y�}�^%
1"O���lD�؄��!W2"���`"O$�'�P�q�$Q���R�ĩw"O0��fK�NՖ��f��@��JT"O��BA*O4��#l���d�;�"O�8"HQ(_�: B��P6r���E"O�)�h�)Z�@L���(+�Z�"OZ�����sp���T�����X�"O�I�'K�@�F�[rc\7[�Ԡ�"O���p�I2�@)$�.`���U"O��QD�I!T}��^�$�:鳣"O���qjS�:0��6�Z�\����"OL032-�!
DiA���6�\��#"O<�k�b��K���0� 'SO����"O��� 9�z!2a 
�67j@3P"O�1��o0~RS	�c�|��"O`-��锫4(.Ջ`g�*M�$�"O��91!�=~�������N�f��"O��@�׏	���*S�+���T"O�%�c��U��QP!AؠV��\@�"Or���*��w�	�$"4�"O���Y����RNE {��"O�{FK�i����®��:��#F"O��Ro�]���� �
3�H"O���L���P(���56�f	�"O"]Ck�%�L1y��)$�2�ل"O<�v ��\\���9��S"O����h;��9(�L2���[�"Ozy@�h��j�D�`���9g"O�@��*��$8�A(�.�m�H��#"O�B7斩Io8��-��s،b�"O��:v�_�T�ġ����+�n�sG"O����*���A2P�^-��"O��)���2<�hsD`Đ9�L�[T"O����=`wp����B$w��Y�d"OX-�CL�7#���A�X#.ǒm�"Ov��d�����2��/#��q"OLdJ꒳d϶d��F�5���6"O�к&+h��;��D0&�.p%"O���UΏ�j>��_�ɱ�ՔN�ў<���9>k�>���!Po������;����*1D��6�۴*�����C�6��ɸ�Jkӄy�eXz��O?7�����EK<!%��Y�{(!�,k�V�)�%�8
x��3$ӧD����).g�i�O�0=y��]-^w�Xq�Y>u�}k���G8��Q���6� [w+������V��9�fhS�K(q�!�D��BH�a�a.E"V��q�$�ΑR��a8����V �'E@��f!d`�'?��;q`����H�b="��]7G#�Մ�S�? ��ɠkSt���h"ǔ�k���ɳc��*ag
�&uD��O�`���B;Ubf ��y�m�qwQ#���40w������p<id��"����cקlGvh��L f[�)H�	C̾��ǨW<S�J��:rI4(6��D�azb.ű
�J\+&�*�E+����dP1Q�S��>�܍h��҈i��i�<y1��_)�(��P zЌtd �d��C�ɓd��H�����D�B8�b��i]d)��&`Baq�J#/��d��Fg��P����@�	�-5�21GV�@5���t��V��/��"�35M2�xgf'&��\"��V�
o�v�S��gi2)	�K����\�H��,k�i)�={�vm2����,��͑�Q�qp��?��)и$ڪ$���G�AO��I�/ީ\�V�H����o/@��^;���-O��h E��z��z��Gd�|y��V�Z�|���)��XvTqR�=E�<!�`�8[��'M���TH�G���[q�5 x:��Q�B6@)����'+bL*�I2'òA@�/�,.a܅J��%q�J=KR��������F�*.n6��fL�םJ}��e��c���\��p��o��:���˧�>�O��S4�7~z����cO8e�gɱ�X���0�a�� |�}ax��Sn���'���)�CH1�|��$��d�`p
���T�#�> �e��gH���id�^w����U��&�3tn294x��O2%�𯙢u��u�	�dm�:�`U l)dL��	��0�n��'�Vذp��L`ɧ� G� OfL��G�̣^*�0ZC��6tP�b�Y�Fw|��O��`��D��pA��h�8�@�d�4}y�HGl�8��O�1��hC�|JeȐ:�
HįI�O�:`C�r�<	�� �q�f\���U�ܰrMτS� l!���l;�A�'��XD�,O�( �Vm>���l_�-���5"O
}�rO���\�%�we���P�+�4����N')VZ�H�!<O\�	�f
�B�x��π'�P����'���c 	�.-�Y#��P�A�\���EF�:^�����w�:q�',�qS�jӞ Ȉ�UI�/&����{Fגz�u��Z�T��I���G�	%�p�'��_{�t!G[��y2��!������:%�=�7,+D�T�q�
X8[�¡[�'[R=F�,O��1�@,2��N]�yE:���"OhոF�
d�kt�+p>t��֍9gD�6gкC�ڱ
דS��(�T��w�t��S���&\O@�J1G^+��E�!
w��1��:0Fp {V���]~Dp�"O�D��@����Q�=��d�Bvu��	S�Ox�>e���]_�}2g���S���2D�6D�������TSA'� J�QRD��(w�1�J4��	o��~�éI�rY�%��0G01�g\��y2�T�r� i�I��c`r�@Ff�
�?qG�e�
�&'lO��9����B�:��w抱x���AD�'V���N#C�Bb�A����+�!d�������yR YjrJl!���$������(OȘqp`٘ꈟ��që8,�B��$遃�N���"O��bg_ċR������A`"O�E��̙��Uk����GLԩS�"O 	ʒ� ��������f�xR�"O��kN[� �F�[ōҟ;�}�`"O*A�wgQr3*�A���?t��m�"O�4P��  u�(u��'I�} 7o�to�pG
"Q�:|�
Qq�q��'W|P�G�&"&��2�N�4��'Vx@�$,�>F�Q�#�G�/�.x�$N��X���K� $=Sz$�H�&O��yB��c�(49q�K��2)2�k����O�e�� ,{l��hP/+|M�Qf�yP�L4O��xh�v��/02��'N����]C:4��Fа;k���.OT�P�D�����J��#��-+W�ő��O������!LB��F�ī3���;D��+����E�p�@�N[�<�y�hX�4�<b�2⾵����(�������K<A"͔7qS��)$��n��4��&�g��tjR��4\�!��@ʲR�45Z�Ě) �� ��X�0R rB��*��'�\1t�Еw�ҥ��(��U��J�����@]�*7jO�FXE
��H�7]����-}�z�����!h��pc�ɼ�xB�O��@#�-o���p큄��D�-�$��RC�����91������D-t0�գ�F+5_�0
2�y�(�0k����a�..��)����>G�<��m͝�b��"�x���KL~��<��,t>�;�郳`=&,�2.|5���[n��1�Jn͌X`��Q-\�$�A�Y�A��ȆL�6X�����<� r�!2��*sf��`���l1&�'9�ĉ��Jl�����]b�H���ޠ������ѢmT*,%%ZK�<Y�d`�]����	.Ļ�#�@�<!�2��a�iB���	`��W}�<e3ghB!Z�GK�]� Ly�<�o̍~����N/%0P�I�������	nD�'q�)Y�%=v������1pt	��'X�Ā�L�5	�(�V�J)t��`��yB�J�v��t�ƥL�O��y�/�f�Q3J�S����'�L��O�<��My� ��s�$��4�\��%�+O�ջ�2�3}�B�cd,Ōqr4�'�����x��vtP��ՎL.4w �sunV:Q\$!*�G��[���bS�'���q� �V�8�Q#��a`0\XϓS�𑣇�gj>HH�'�,�rf�]:&�*�;�mQ�^�a�'r>�!�)U>!�J�������zJ>��������ӈ��%��!'~��p��ڕu>*��F"Oؙ8��5|#~� O�� H�@���U4DA�R�(1TBD�g�d��|���C��XMf�R� �s%��D�!�蕁��H�uKd�ҰD*A<l�P��]���i�&�O���w�O�P2��B�?��@"��'Q6��c��<��T2�3O�Y�`�1Z$�a�D� s�+�"O�����\b�0��OǱ6f
���<��ݾY�HG����Pt���T�׾s7ƕ��]�y�D�Z�4"�@��^'\}B/[�$bN��e�!�ۭ�(��ɪN�㢋_(��Bq
�i#�C�	�T��a2�*΢F���BmS�[�TB�ɗo��QVb׺Bz�CҬR�'�8B䉒_{�]PT�L�!�ܴ��ǍG��C�|&��y��Y�vD� S���C� AA�T�� �= .�z�H�e*tC�I#%���k�1W�Ӌ�60NC��3�"��ř���!��2{C��%+�eʱ�C7X`&$�^Y�B�	����W�@�i� t����(C�B�	��	
�ǘ:m��������B�	�˾�90j�	i��i �"R;"�B��	&}X\��?<��@B����B�	N�t�n�/b�Q���i��ȓr�hl�e�B"G�R8��l���ɇȓ{N����*O�ab���Ԅ�ȓ3A`���:����L-����9B|9�&�D9���g�I;�*���Z�ĐסZt��O[���ª���%��oȀ���/��x��^ՠ���K��
Q�U	@]���ȓ��C$�_�!�L�A�#4�D��!��(wi	�Y�΀Y���xɸ(�ȓ-�
]�T �	���Vڹ|fZ��ȓ)*DB��G
.M�5�̶;�b��ȓh����O;4��D�$0z\��ޢ��`���c�Zq�a͙�GX���p��ud.�UE�99��XY��}�� ����c!$(��9Q���ȓhL��c�4�R}�!�_8�Ze�ȓ?)JE��θ:Um�:놀�cB�����S�M(Tڸ���Ɍ���K�E=[�O=o�C�6���h�Io�6���')+/�C�I�aVv̘0cǁ@~uZQ��0M7zC�+/
Hl�TN�����صJabC�	�.�����ͤW�R����{�B�	#r`��Kd�_�e��D�&I��:��C�U�%�[�.4Ա��L%xuC�]��7�
l�A�VY�t�Ny��'�L}y�����{�B[�'T� P��Q��0�v�OE���JE�H�%�>P�zb����� ��Y�F�Vst<�w����7��]?���>��4E�=�0|Z�E�XG������=-,��Ɯ�-�ˈ_�T����%2���)§��dŇ�Q��e�!�[�"(`���3RW~��6c��p0�b9���Yi>%���,F`Ԍ�$�;(���sF�M���jf��Y@�f'ő]}�,&>�}é�00�|��b�
�nh �8%�ڗ0���Y������,k^a�4��;DNXb,Ѣ�J̀��3w��	"E ����M�g��S�'��PQUh=)d&\�0��Y��m�Bz�M)#��)��O�3}�*P���q�[��f5#w�Z.�?	������"~e&٣#�܌�U��l���ɀPg�92
�'g
\��"�
���}j�*7H��y"�U��()0)��"�0�$E��y�ǈ�%���� �@�f� "B��y���t�hibB��:�n�b�l��y�o\�S�� �d`��Z�Ζ��y��I&O�QC�T�PD!�W$�yriP�Rkp�#PO�GoȤP�^��y�ŎW6�ÆE8c꩘s���y���|E"�'f�����yRȃ9(jf���K�ؕ����ybl�,����2I�-�jY��c�Py�'�-j�$=ۗMQ�o�$qz�@�<��ҸJ��]kfJ�>C��Љ�T�<���owv�X'f��#�pٖ�P�<AR�+/��v�[�'H��Z�Q�<)���0Lʹ%��eW�U�P*6D�N�<Qu�Cc%n�I7%��-=r9�nFa�<��X�2�-�S�%��)j��Q`�<�ы�R���(Q�CL�	ԃ�Y�<�2J��i��t$��
Oi�511��U�<�$ �%J�l�v�	���*�]�<�a@�@����+:�L�0'*�d�<Q���7F�P]৹B9�e�Ŋ1f�B�	�ag<}�%�]����#�D�I|�B�	/j��#c6Yu6� ��0�B�8�Lܛ�$G���������O̒B䉣;�b|�s�@�q�tt�E�A>h��B�I7D�\��#�J�^� ��C<.��B�I1d,��@�V�MvL8�uc��.{�B��.8$�� ���En(���$Ҁ��C�I*"Z��@i�}{"�X�AN#�C䉜JyȀ��h��RS8x����\�B�ɖ	����2p�e� 	3?�C�I Ӧm����iNܭk�%�	-��C䉓� �`�Iȹ��v �C��"T���`O�<�����[^M�C䉔D}�i��\<"�XH�vB[1��C�I9I`����J�g[�x�)!:�C��2��L#�`]�MB͡��
r��C�I�Y2+F��^�8SAF�)V:��'m�A�NE	�x��h�H��H��'f�����L�8�	cCP�E�.5C�'��q�����eF� 0R�:*_z���')�h�!�J
93����n� c���'���0m�m��y�@�V���y�'���KehO�3朹��F:; 9A�'���T�K8*FXD�҆,v���'���eW�H���bC邷T��3
�'+rx�"�)�����T ���r�'4�2���l�(I+6�ߍ_����'U��Y�a[:!@�+YT����'���3�@^��k����`A	�'�6�����O|�t��;�1��'-�ɠ/�%8�yP�nW�;�<���'�cSD�w��\%ޔ0e������ �͊A@�T�ƨ8CBT$67�`�"O�s���)R�j�� оa")
0"OL-��5 �J��N�
=��JC"O��b��%p�����"#�Qp"OA��GK�0�ݐ���zl�"O�hr$�<0i�U�H<["�X�"Oڌ��J1�0B��$ZP��"O<i�	@�>T�e�(at���y盇jLt���� ��h
0���y�N�d��pY� SG�v:gA )�y��q�J陲�
�2�^�����y"g��^���˘�W�)P���yb�¦���A���N]>��A�م�y�(B3��,*���>*��A��y"�_ a`��{�DI=V�����Q��y�J��3L�0�BY�`��a˜�y�ճ!\�(����2G��yB�Ϳ�y������,)dh�1֨�sRÝ�y��	 �%a�@H�, h\Af�0�y���M��P��	�8$�����y�aD�E�f�80BB�6j��K
�y�&�7hܤ ��e����pxW� 	�yR`�,��4���+
0��e�_��y2�ˊ~"V<����U���9E�(�y"/�$H��R�U� �����y�P�46�PAifI�L�0@E�ȓV����G��d�f��m��p\�!�Ũ�en�*b��?[E&9��uV���g�(@��rS��N�<�ȓ	P��"�]&F��-���֤z�D	�ȓDHp,	�  �s!�i��FHyz�8�ȓs)�t*�%��$K��Xc���G<��VkF�H"�`%����ȓl~,i��n�
�b�4�ˆ>;)�ȓ�&Yq�#�lA�@H+�$�&��ȓ	U\s1(�IQ �+�·{��}��goJ!��`@�F�I��Ǳ'"�B剐g�"i{dO�iִt1a�& æB�I\@H�4 ��,�XhrS.7�B�	�6#b��NA�f�P1萴.>�B��R���*��Ƞ$�7D�]f�B�	<���V�DY;���ӛw�xB�@�(�&ַkՂ��A P/Y�lB�əQX$K�cT?$���-��B�I�e�jl�W�W�#����V�T�t}�B�	�g���ꔧB;�Ї�*��B�I=etba{2c�Y�"�q hR���B�I.Z$��zv��$/��6�.<�C�ɯL�D�4�C�j�5*���DA`	�'�$l)�nȶK�E#�! tdY�	�'��\8��ɟG�f��Kt��	�'}�5z�'�*k N���N�2�
 �	�'�,=�OD�#��VP�SdP��	�'~����aI���f��R궜"
�'`ZEN[��^uL�2-��'�0��b[�n)L̐%���>�h�z�'+������8�H50��<XD��'����A��-u���/## *@Z�'����e��:ԭ�+��$�t�>D��{6�D-��|�cmũs���Bb:D��yP�Uv��@�"�ƎiP��+D���͇c�V]R�K�$VXF|�2�*D�T��A�gT!q��_�~�:�	s$D���	S86�f�afd�&pM�2c/D�� �|h��<8����KS�u�:�1 "OjMs���\cd,���!?��Q "O���Ѧ[�r���T)��|pg"O���BZ�(�PZ��84�@"Oܠʷ"$j��5ڒ��ܐ��"O�8q�Ɂ3d��x�����Iq"Ol�Æ�� @�$,A�w�$�"O\�I���9�p4��J( �6�;`"Or�y�Gˍ{�$x����H�N-9�"O���3A�,
��)A&:	��p5"OV�3JR�H`����G�Ľ,�y�JZ�6P���̵L�>��%��yB
]cqj�"s��Z���eH�B�<sZ$4�̍��ʝ�K���P"O��Q�_�Q�p�EW���� �"O֝����?C�j������@H�!"O:\�'��.�����->@k�"O���Y	]@�H0q�!z��8`�"Ol� D��!)hu l[f
@Q"ObIRp��f���hw	��Q����"O�E!&Y%��9R��>�d�@4"Oplsѧ	�. t���g��?Ƣ�ò"O��q��v�21��֊9MD���"O&)0�5 f!⤣�0L�Mj�"O���4�� ��0h���J6����"O4����ΦJa����[=)>��"O���A�ݜh��$�#�ۛ/	H-�S"O�yS�
Bn~<5����sd��d"Ox���
M����t�IM6���"O��Iec[��\���IK>����"O��`R�G�<��L�G��;���a"Of�×�P2-p]��H@{{�m�'"O��0�-ޝtЄ�ѡ��_hƐ
�"O���J�+�r�bN���)J�"O(�ÏS�^|���&�e���q"ONYЁ��h���֎��
J��"Op�K��F=cpL�Tl�h]R� �"OȘb��{5,1�M͍/3���'IN��s�N2lP����M�:��#	�'��h5��9H��y��<W�Pa�'_��9�/�0�t��<��
�'����"Ӗa�,hK��[�C>:�3
�'�(�#D+Y�]���0>� x!
�'��8�"�<i4&��I�i#�@	�']d�P@E�m(����R�L��'�j��QC��w����A�*M��S�'+"��p�-E%��+Q�U�5�:��'g��a7F��g8Erqك:T�%�'`��jw�
#P�&๠��.k�'�0�H��	�*�n��#�VeY�'�JYZ�F�tX�H
����t �'y~l{�'�39;�a��P�V\r��	�'�� ��*~���*THĄl^��'\n$r0kĩ\����X,"H`�'���3����N1M�*x��7D��;Ƌƙ�zIj��Ǩ#M�ݳ#�6D�\04(�8��-�A���<���t�9D�Сg�meX9�Jc��,�ӭ��y ��cb
�#K�<��� P$�y�K����"��EJԙ�r�Ҷ�y�b@�[�v� �I@�B8 �����y�GΫ\���"F�H Ȭs�I��y"iX�b��d�����>���.ʛ�yR"ԝe��	���E�����C��y
� ������d�p�'��1R��x�"Of���+�A3PY A퓭_��7"O,���	E�j�$H�E%�5/.5��"O��d��q���Pd��#E aP"Oj���Ӏ. �4�w�7'��a�"OJ}��BM��p����P�_�q��"O��T-�EY ��<z�<�U"O 3�c� ^|�Agk&KΪL�"O����@+2\IF�@�k��u:�"O�%�w'
:����2
v��l{�"O�-��Y0�S�Jh�`"O����GT"^�P�2Í�3A����b"O��{�g��:�&�y��ʦ����*O�y��JG���b/G'H�Q�'�ܠ6g�F�b��%X1Z���'g^�
K.'�*�`ܘ=���K�'�f�bI|�<���Թk� !�'������s��İ�E�^gB�*
�'����f�d�"0amY����	�'�bպ�KU��B�X2���V�Fl�
�'�jx�  ���   �  C  �  �  �*  w6  *B  �M  iY  e  q  K|  3�  �  �  �  �  ]�  ��  �  ]�  ��  ��  ��  �  O�  ��  V�  ��  J�  � � , � h �! '( ;2 	9 L? [G �M wT �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�'��7m�?3�p�)2N�&g]��*ϓ�Zφu����,�ݴ�����'�"nlr�q%�E)-`�����:�r�'hr��iw���|bA�O��)�t u=#�h���	W4+���<�����4ڧk���j���=3�6[��
b�,Z'�ie�,��yb�i�ڦ�ݛ,���d�!&�;$,A�;�R��	ΟDΓ���	�^46m`�t�E`�p��%]���2��t�P�p 2Mm�����'.�8bG�C�8 z��;1I�(R�'E�O�I�M;�˛C�Fmv��'֏el�C��:6\ui����>����?�'<�ɯF�*Iɇ��<Yެ��Zn��?���><�ޠ�|��+�Oܠ��l��|���B�`([ LK�2O�0�.O��?E��'Lt��ӯT�L����L�6LI��y,|��,𘟌�ݴ������V,ws��c!�ΗM�k��� �y2�'�r�'o��b�iD���|2'�O��!���N����!�6)����Gb��My�O��'.B�'���_�v� 1��k�/2��GM!n��I��M��aɐ�?���?�M~�<�t�*phR/�J���ӋU�>\�`_�x��4��6J9��	?K��S�%��"�L�;��C$$fx� ��= ��:'h0DrA"ŕ���<��*�I�rd�,�d�>F#�����fM�Iן��	����i>U�'�v6ّ��$��c�b����ѳp��h��Ъ%����Z̦)�?ѕS�T�޴c����n��b�bR?#�V@Zc��&r�^x�f(�6)h�7m+?Q�)��
���)���s�=�f"�|�Pn��hR�鷢�K��ן���ʟ��I����|����B】2`�M��O+ �&�3���?y�Z�F���~%���MsI>��_#L�x��Lՙn~=j6b6
��'K�6��ɦ�/a���mZs~�!P�FO����	$����A��TǄ�U%�ݟ�@Y��4��4� ���O��R�'X`��Y��X��C,�M>��$�O˓�����,*2�'��P>5�n�|Ot$�rd(y�8����9?1sU�`�I̦]�O>�O��ucr��X��3b��)G�D���&u�@(��P;�����{S��Oα�+O�T�4�Q� ������W�K�~���O>�D�O���	�<�T�i%��d�Q^S�D�"B�^H����M��'D26-+�Ɋ���g��,aG�֏%dݫ��ɮ|	�{�FҦ���4xɰh�ٴ��dhVѓ����S�?P���e
�g�Q;3��p����۴���O�D�O����O���|R�ݻsA�\S�@BE%�kB
�vK<k���ʟ $?��ɓ�MϻD��tH��(I'����S�f�I��'����$���tET?ԛ�=O*D`��͖7NF�k�>���S5O�h��$:�?1ᣩ<A��i��i>9��>G���JeF�}꘡R0�S������,����'��7�í3�`���Ot�DS�7���v�6 �Ed��?2~$����Ol�n��Ms$�x�/&|��Y�
�r��H�:���'{����FQZ
�O�T��#3��dQ0�?��G�	�dTc���*d����'�̫�?����?)��?Ɏ���O�mY�ڥ�p�z"����8��Ԍ�O�Mo�p�p��矠��4���y���c���׉wTP�[3���y�EoӘ�n��M��f ��Mk�O��³Fş�s��.�R���Z�y:�$�N�,˓O�f]��S͟�������|��#� ~l,���Բ#Z����Eyrco�N0�&$�O$��O���d�?!>��'G!�Uh$!J(��'� 7�Y릭�L<�|��F��'�2YC�%ۆ�"��͚���ȁh_~�׼5=��I&>I�I9�M�)O���,M00Ҝ3���#MdT	b�O��D�O��$�O�ɪ<���i�j	q�'wZŲ�$�W�n�jqh�,�rl�`�'7�6�3�	����D��͹ٴ<����7���8��G�Z�XT�"�z�. ��i��\�Xp`OD�n �iq�)�D�~�� ��c��PZ9V|��*A9bT�0�0?O
���Oh�d�O��D�O.���Y�� K`��b�X]� �C��Z�Vr��$�O����}	�ln>��������Wy¬L�zr��TOاW��Yd�\>��6m�<iC�i��7=���A�q�
�de��KG�P�A�p�R�ߌ/�h�1 gؑe� %
�+���?���s����uڟ>���O��8B��� ���3v�se�\(6v��d�O�˓&%Z����d�Oxm��?=i��Z��]Nm@�d�$	o���OH*�t�X����ūݴ��O�̄1��!G��BJ�_xP"�̝C}Du��A���D�ٺ/�6�T��?��Ӽ˕�S�\BI���e8X��Ȕ��?a��?I���?ͧ�?�����Pצc�j�����*�B2TV��d�6������ܟ<����]�<z�4%�@-�"�7B5z�C�L�7)��!R��i�P6MA�$7�.?Q���7S6v�i2���N>�HD���j�2�A��յl��6�<���?���?A��?!*��e�(/
����
~�4���[Ǧ��!��JL^Y�	Ɵ���/���i>i�i�%��([;ь����%"�Z��@U��MU�i�z7��<�|���1�M�'_"�"�oQ�k`x�IV��e���<��h�5!���_��������4�'�T��d��?�%��!#�D ���'�r�'rY�X�ش/��Q��?��N.\:�cڎx�a�%�,c��	�OL��?a.O��lZ�Mŵi��	�@��h�e�)5A�KuL��V�>?�抩�9���	W~�jmݕx��'U�4�I�x�P�`&S*�l�CQiշ#;�����P�	񟈗��)�O���O0TҴ�����c͌R��%AQ�O �l?Q8|��	����	ş�����w�~�Ɇ�oj6e� �ԒR�:���'�j6M��3ݴN�ߴ��D��.�@yJ��6x�d��e�V,��f� i4���E�O:�ĄҦ����t�'��'��'R ��*k{�U:��""�����V�Y�4!�(��(Ȼ�?Y����"��.��E?<^jla�*�J��<2ѩA�y}���'ɾ6M��	X�43��>Qr��P`�Ւ���fR~���,r�H�(?I2�K"Z��������'�8Ȋb��gh}Ү�5�*Hڥ�'���'������_���4|t��*�dZf�
1M��i�h-�v����x]H�/ۛ��$�ty"�'��fk�J!���	"��=S�#G�uw���K(m��7*?�"D\�C���+�$ehݙ��2ar�}pc��>%XȘw�Yj�D�ǟ���ڟ����Ii�'�\��(��|�T.@�7�҄p���?q��R����_��D�'JB7�5��ݽ\�����a��`����Qמ0��'�<��4h��O�.�
2�i�d�5��KeoǉBe�l�F�I�.�rŐ�I-N��TK�h�
�'�\��'��'c�'gd1R��6C���%��Iה��@�'��_��s�4.z-��?Y����)]9��	��+���"jIo�������O�7�Q_�|�Ƭ5Vh]q&:ȼ,���9n�U�ЀV�'r����d��`�U�|�
C� V����O��ج�vb�1�I͟��	៴�)�iy2�k�� ;���P, hq��ԦO����LK��I��M���j�>)ƷiR��1#��#"i*��U�L����!/|�R�mZ4-�n�L~��̶"D(<��n�)P6Z��Q��W�c�Dڴ%X�J*��<���?!���?����?!/����F�`��� A�Yl�.GB�7��x��D�O~��/�9O��nz���`S:L�3�!�#Po��P���MK±i�NO1�d9B��t���ɢ!,�z4(��ZJ*XӲ�����ɩG�@]�%�'�x%�L����'w�x�t��x?>��w��$h��!�f�'=��'�Y�X�4q�����?���Y��r��œ9XVM�RÌ�a�������<Q��?�I<q���)�2���E��ZuiANA~��J�咑��W��OP���	�W��L��x#�RQ�H5�.���#C�^��'���'����QEP�^���!ݥ;�b�! ܟ�ڴh�
��,O(oZL�Ӽ����_�H��ȌK:)�7��<�׾i����`���Ѧ@~� �H�(hWn�2��`DE��I�E(��i�x��d*������ON���O����O��D��/�� �Ac�$��I����wJ6ʓG�&N�"��ԟ�&?a�	�x�~��Q�O'�:��0c߻G���ʯO")m�*�?aL<�|j�l�6���� ��^�N���,<i SȈ����Z�� ���)�<�OʓV����9d����R�F�n���(��?I���?���|�+O�DovCF��	u�Q������$jɜp��	,�Mۉ��<����?��44� ���E[3v�X�;���&���M�M;�O�8"��?�r֌4���� �[���<!)����G]�p� ��s?OL���O��$�Ob���O��?{�HZ�Q,�C� H�H�&/�py�'��7M
�5���M�M>9⁓�
���C�y�RG�#�'g 6�Vܟ��S�H�R7M#?	⁍E�b��p�S�my>��
�`k�d����OՑL>�,O&�D�O����Op1�d�V�ߐ�S�!h��{w��O\�$�<1��ib� ���'o��'s�S�/7DX #��#����]�hF�$�I&�M���' �����O��``��<�F���ȓt��	e(	
���Sb��m��	�?�3�'��a&�pr§��u�x���D�\�|(#�#�����ğ4���b>!�'�6�Š����a��B�@��#��Ox��̦��?��S� �ٴv;���S��*,�C�ľcȬғ�iM2�E�(��5O���O�A}�t ����)� �p��ǳ?�����ϖE�79O|ʓ�?1���?����?����)G�|��S�XL"��R7v1
tl��?b�t�I˟��L�'|՛�we�P�� [l_v�I��B�0��RR�o�ioԟ<���OAli�p�i��D��f ���'����U��y��ě�z{�e���{�O���|���!�y�E(Ѻ^т�)�M�P$�İ��?����?1/O�oX"ެ�I����	��vT �F13k��*<p���?��^��	�4Rg���'��43�hLQ��//1�\H�E�!�\^N��M�Q2p��|����OB����+ E�C��w�֑�w�
P�����?��?���h����س7��8�.�G��H�2/�����¦Ey�Ĉ��d����M���w��9;��F�$ᢱ����,����'l6-��M�I+�t�mZK~b�H�,����ӵC���e!F7�ҹAĊ/4�'�|�Z��Sן ����D�	֟ �4��?@�ʅГ�N/}�l��[_y��g�Jmj� �O����O\����$ҋ�,٠�@�*o6�[U���s2���'�T7m�����ɿ�H��Mj�햣0 �C�O�TW�C�C�u+r8£��$+B��?�F�c�Oyb���v@�c ��,���AI�1	3r�'���'��Oe��MC����<�׾A�RUB���}�������y�,t�@㟀J�O�oڋ�M�Ǿi�d�'\�İzׇ����c�ƖZ��&���[ª�5Q������f�p�f�:��1�Um�#$�f?O����O���O����Oz�?�h�!V)=�P�g�B�(F�����$��6�MÕ�z~�feӸ�O:5S4��N|pU���ڒO�@qw�s≕�M����&��(�&��hj�MR">Z��s%�(�\�2p�_ 6���(b�'X�m$�Д��4�'��'���Gg��K��@�%`�mTh��v�'a_���۴S����'2U>�He݆	[@�)WU�P�H��!�8?	�^�4��4*��A"�?�s�A0|���QW�2{،ht��09�,8��>u���|"a��O�1JN>Q�	���	7�X�iv�B��ܼ�?Y��?���?�|/O�(n�0Y� ��R��V��(�I��	��y��-���<�I��M�����>��i[�E0��'_��9�h[�/�M`���O7���06-5?�rȂ�z��I݀��3@9>qRbH�,��H)���2n��<��?����?���?�*�"]��	~�!��_t���������� ��Ο0�Iԟ@&?=�I��M�;:� B��?g\1Be��W���MC0�'���O�И���i$�D�Vq��K���3R("�7�ǐ/o��0��([�v��O�ʓ�?���~�ViA�^Na�"���<E�Qy���?q���?I*O�qm�4�2��	ҟ�	y�.���G	,`;�H�+L�<�?	�S�(��4hR�x�Q
'J$�����҈�3e�<���JA�у��ؐ~8ғ�����y8@�$Ƙ`�ʍH���ud��E!8
���O��$�O��D �'�?���)��rgĔ y~��HF���?A�i�LX`_�|�޴���yW��0'VF����
�fV1=OR��; ����O�6��H��7�<?9�fG�1JL���uf`h叞�EO\���H+�,EM>�,OD���Op���O�$�OW�:К�b��Htl⨚ŤJ9������jd�����ߟ(&?���0rh�
��ݠ�&T �m�0C��b�O��lZ�?�H<�|z2��G��\�0��*8�����'w6U��H���$�3~��ȡ��'=<�O��x�D��� v��|�Ы?n��H����?a���?���|�(O�~(@��F�'$r��V���kfᐟx?�u�'�p7�7�� ���F�}���M�!B�sG�]���F���R ӭ �bŉ۴��J��H�h�'o�v��|��N�~x�h�FO47�6̻FFW/L�D�OD���O���OD��)�S,�I���#�l��TfL�����џ�����M�fS�D�i��O%1F�<A�\���"_�C� �R��/�M�����D���}ћV��0J҅�x��i#��ʠstQ10Έ�K�����'c�&�������'b�'a�8J���.���㐻kpsv,Tk�$�fT�\9�4��@1�OG�'c���wt=Ӧ��9$՚�{堚�v&���'krW�؀ܴ)��]�l�O$��˒�OH����.�)+��ذ��/�,��4�Z�iq���GZ���S�i�b�_{�ɂ0�By ɟ�|��I0$��.Y?���	ԟd��ݟ��)�Nyr�d�D���K�yD }�^-������bΰ�H��6��_my��i�n���啂#���'�ȂF�Ĺ�Hf�Ȱnڕ~Z��m��<��,��!����>4�-OpM{w՜A%�1`A�٠�e��>OX��?����?���?������Z�4�Ha!��);0�d@S���um� ]�-�	D���?9�O	���yW�74�bܓ|�f� �G�`��7�矀�'~�O,���OjPz��ik�dʢ��1�#�ܿK�� $Ɔi���Eb����Hr�O���?��^Ą��rf�Y���1�O�S�p�b��?��?�/O��lڊLGp0������I/��BU�SW���h��ًa?V�?�\�DaݴJ��x�hI)zB|ɲ$D>;o���č��yR�'r!�#..`@�\1\����S�2�T�l���]�r�������a�^�i%Tܟ��	�����՟(D���'��x�Ó 5# �A�8/JA���'�7��r�J�l�f�4��4a�BX=E`D���X�0����O*6MO����ش,Op�4�y�'�4D d�?�Q	� t5�A�9)bR�;p��`>���<����?9���?!���?�SɅ�Ls$4:ъˡCC
��G����dC�����ߟ���䟄$?�I$4hp	p⨗�e2�#�n�#w?���O�`lZ��?iO<�'���'N�Ct�S���!v-���[7禈r/O�dX��U>�?9"�4�D�<Y�Y�(�@i eꝔF��}�!߲�?Y��?����?�'���T���: F�㟼QP*��%��HA���Q�r�۟�ڴ��'���}�����O6M��w�X�(�,_<u>X�CM�R:Ќ��mv���	՟0CE,��Yly�Om��;)�D�	�9H�A���y��'9r�'���'>B��1]n�����0�R���jXd/p��?�Ķi�Dq�O�" i�*�O�����`ܴ�æ������!x�I��M˒�i��4��Rz�f<O$��ظS��)�DZ�5�uh&�X>$}�d2s��?��@4�d�<���?)��?�v� �X����U�ߦx� rH�?�������(T���ϟ�Oo�䣁Ş��V ��΃�P<��O��''T6�QߦA�O<�On�����0���1��w.n���(� x�&��4�` �?,|�O�ɗC\0+��왶�;�N�� e�O��d�O���O1�xʓ]?��Х����2�'W�^p�F�(ܜiP�X�P:ٴ��'�^�N̛��mZ`8� �@6ȝ�U�ףI��7��˦qz���}�'^:Ga��?����d�s�J3�:��׭��zR�8O���?I��?���?�������~�Z ��%q�iB �V�lںs��y���`�Ie�S��I���k5�h��P�7�1R澡Y����&R��s��%�b>���D¦��9+�+��I� �B7MwK�,�@�%�P��O��yO>�(O���O8}p�jD�_�z�`KȔR\���(�Ol��O��D�<QP�ih�`�EU����+�
u��_�_��Q ��I.`<��?��\�t�ڴ"����8��0�D�±ŏ�Z𶕨�FF'���'.���wl��,D�b>��'N���	�$)j��צt|�e�(ɲ&������������z�O�R!I�.&�xZ�(E�r�z���׶(�!f�>ĀD��O��DOЦi�?�;FBIb��6!�x;d�@�����Oj7m�)n�R6'?	T�^�	�����HVX���հb��ÔC0&���N>�,O����O$�d�O����Ot8�7*�x˒�	��|r�ϭ<y��i`�Ԃ�U�\��V�S۟Ƞ`ɐ82n�B�zn���IK��d Ӧي����|�����P	_�Y����2�"u
�d�7 ���N���Г}_�p�c<>�O��L����3��ʇa0�������?����?���|�.O
qm�)N�vp�ɝc�rQ:��܊F���DHDʨ��	��M���<����?!�4+�J�jA�����p��� V121cǫ�*�M˞'
�)FfH����9l��?I��W,\��iG)~���T�Q�>��şl�	��<��˟���|�'Q'��H�ܩN�.pУ�O�O��D3���?���">�6��:����'��7�(��[�"b��zc��28@�AvN1,��$���4zƛ��O��ca�i���O��%&
a�j�k�䙫x|�r�ǆ�C��H���N�O�ʓ�?��?��G�VM񑊘=�T�+���!�~����?q)O�oQ2���˟8��P�Da��K�h�GGP�r�P�X��F���d�b}�f�����Q�)���K�@쪙�������n/X��$>���+O�ɇ��?Ao&���T�X��'�3��$��&ԌFz�d�OX�$�O��<�$�i��!B��Z_<8�@�h�'gS�T�r�'%07m(����DB�Eې`�,]�IK��^�T8��\��Mۅ�iB� �v�i���/\��-S��O2�)�Δ��
L�7%�ش�΃}��mϓ��D�O����O��d�O\�ĸ|Z凁�Y��#qŅ�?��A:�d�K:���|&��'7��O��ޟ��i�qYCJN9:xx�Z�3YF��?�۴�?a�O�O�4����i~�J�U=���Fj�� ��l	����Ro�\����t�O���|���C������ :`n��,�r>�#��?���?9(O\�m�0j
�	����Ɍ\�7+�X�+����І�N��$
���M �iG0O&�����?>��tj%�;��xC7O���I�lP:���H�0����?�r��'o�I�I�cJ�EQ��(89�����*$�����ܟ�I�4��k�O��l��@�㎨{l����R7l��l��xA�O��D�ʦ��?�;��U0��_>a� ��� �:����?!ߴM	�v

������xJ������+v�٩�&R<$�Rɔ9D=<Y$�(����'���'��'���`
�k���Ń] L�|a�[�\1�4h��x��?Y�����<�(�>����N�/y$P�dI�V��	��M���i��O1�����AI���{F/��x!S@�4`BU����"� �/n")BP��|yҋΧ8����@��� � �D�
0�R�'�r�' �O��Ɏ�M��![�?��牦6"G��+=�:�l���?���i��O8�'�D7�P�U��4߬���_�&�`T��GW\��qZ��MK�'���J�?1�E�S���d��Z���4�``��C�<`&�4
$ӻ{�$�O����Of��V���'���\������@�p�Bod�I`�������M���A~� k�T�Ol)�Q
���(�H�EG�p0`��R�	0�M�ױ��tΉ~ɛv���R҆4� zXb� �zy��:����5�\@�d��%�?ٗ'9��<�'�?���?Qwj	��aPa��(p5X)`��%�?�������)�%��̟������OMJ��]��u�Q�j)�UJ�Odp�'��7����l&��'j��qA2��2y܈Y��	z|�ē�"[&��J���4��t)�"픓O��@��a�H������x�%����O����O ���O1�8ʓ|z�&-�-�, Jĝ�88F@�יyB<D���'A�ee�&���ODtl�%s���7�9�h`��*�{gh�+��M��Ύ�M��O���K���ɩ<)���-tN,��5��w�}ps	��<a/Of���O|���OJ�$�O��'#��iP���,Kv�p3oMI��ѓ�if�ђ%�'m��'D��yҏ|��Ζ� 2l+	^�iP����C�4,umZ�?�O<�|R�):�MK�'Z�m�¯��FF���G!��O `��'�
�k�%Y۟�K`�|�U���ܟ�D٪q��r�� ���*�g����쟤��hy��t��X���OH�d�O�)v��
-��=:�M�?�m��&;�����Ė˦�Y����O���ԅV["@�&��<Ge&H�'�D@&�B�m:��g���g�՟L���'��ӆ�W@ubus�׵h���Bg�'���'Mb�'��>��e��D��a�)�"�C:=�m�	��MSf�2������?ͻ�˥@�*�8u���)C�ځϓ|	�FA�O�7
K�\7M(?���)L���i:���@�h
�?W6�r6ǆ Kk��K>Q.O����O����ON���O�T�@<��,h��=|��q��f�<9�iDƅ�D�'@��'p�OAR̲Ek��԰1�Ĉ�'�'4z��?��6��O(O1��A�S" �VKf ��!�a��d�aH�,bn��n�<���!$���U8����DC%G�����K�8��#�P�)N����O��D�Ol�4������)��'�/�%&<i�쵢���T�	�0
����@}BgyӒ\����1�ZB
�h��<(�~p��JǄP��o~�E��`��+�O�W ��YX�#�/[P���R��ɿ�y��'���'�r�'���F7x=S���:�)���>T�˓�?��i!~���O���k�p�O�)�!B��>��I�ꂆ�H:`$\B��ǟ ��ffKo��s
�� ��A<Z�� 3Hy��ҥ��
M�6�$ל����D�O��$�O���H0Q  �2���OeTHB �L�T����O��,��V�ڎ R�Iȟ��O�|2�Fތ[Ќ�zB�^)Q���1�O~9�'ո7���'��'u�;Ƈ��c�r�@�УL��%c�0<V�|��#��4��@���\��O�8���I�8"I����q� ����O��d�O���O1�f�&
�V��&{���p��
�-$�����$	���'ODy��㟼�O�En��d�4�cC6j�n�jV��f�@Q���M{#G� �M��O1�Ș��
B�<Q��>d<B�;s�5����<Y.O
��OD��O����Oʧpf�q�d�ƷcՂ�[�D�/myN��&�i����F�'n�'��OlR+n��ΌG�"��SW
c�t�ԋF9�mZ��M���x��$B֬G���4Op��Kވ_�|	h6שy�Pa�d=O� ��T �?�w+5��<�'�?1�e��3O :���*~>��
�
=�?Y���?�������¦}�5E�����IџHj�'�#I�Ґ`uIՃ�.��d��e�
��I䟼nځ�� �~�d��6����K,p@��'i 8���]A\6����d��Ο���'bR&a�5�*-�w�N�>�P0a��':��'���'-�>��k5ʔ���YO���Ȕ� 4����$�M�Sm���?���ޛ��4���`-���Ց�,�:4���4Or�nZ�M˄�i�ؑ�!�i|�	't��-���O��y�/�s@$Y)	˼X�q�q�\�	|y�O�'���'_��)0�B�H0HB�њ�˔*5���/�MK�,���?I���?AL~��b�i��� !,�"���i�xy�[���428��� �4�|����\�f��?K^n��k�$�$�jiq6T��D��\�e��/�b��m�Zy2-S���IX0/F�3�d�	sj:���'���'��O��	<�MK@%Ή�?ae�4j#(�� [l}�vj�<���i��O���' �6�To��yXB,�k�1]���f		b����	����'"�i�F���?�Zf����w?�`�ή�R�S`M�$޵�'��'�r�'jR�'����*�G�A���;��Q�dV������O�d�Ov�n�6u�p�O���'��I�u�Zh	�|�����J��~�BO<!@�i,V6��^e0�y�R�I���Z��+~&��Q�*����F!H�YJ4�b��'�~�'�Ȗ'���'���'9����Ö8Xn&���4��:��''�S�̨ٴ~�D����?Y����3l�^��<2���X�JW�� �����Uj�����|���<�h\`T!�X22��>~�X��I�;q;������sy�O�ȵ�	���''�qs��F�PJ��4���p��'�2�'�b���O����M3�LM�0v�ms�A�*J`�)r�C:K��1++O`m�S��/J����M����j�A���/Z��TA�I�b��6.c�J����n���I��L���N���
pybg֥"L�k���^u���q��ybR����۟���ϟ��I۟��O�1����x(����H���4Ix���� �O<�d�OT��:������9Eq`��#DI�)��L�׉P�d�T�������|J�'��֬�+�M㘧� ��	t�E$��h���$*zHY�;OPDG��?��=�$�<a���?�ǔ�&��A�H�.����.O�?����?y���dH��%h��W۟���������P+U���k����� Ȗ�Z��7��I�Mk�iP�V�9�mľi@<�%���P�J���m����^D���A�� ����C�O�;�XF\̡��J1 1Ȩ�6�F`�[���?����?����h�n�DU�\D5s�d-@v@\+�F���䦑s�3?)ֶii�O�.<���3b�P:Kj���ЯJ�W��$B���Sߴu,��'_�gT�61O��$�!��`8���,�G�H2�u!QK4�~����2���<�'�?����?1��?��S�k+���r$�*��cw���D���[�}������|%?�+a�����d�78�ti���^�'S.O��v��($��i����I�A�6��fg���c��O��A�/� l��	?U��9��'��u$�0�'%�ૄ+ٴģ��e�����'���'B���X�� �46�Q���T����"�'T�b�Ұh�/`�TA�$��$K}�%q� }��Ħ�;�"�J��9BUQr�ɴ�S����n�^~&�N�D���.h1�G��.��E�Q�M=�|�h�A�yb�'�B�'&"�'�2�	@-Z����%Ѻ�K�o�?1n���O������$�m>��&�MK>����κ�Ҍ�
�{��O��xx%����4���m|��ڴ��:��`kө<���aa.�� �։���:�?�c2�D�<����?���?���I6r}J'�ԳL�8�H߁�?�����d�-�Ӈ՟x�	˟4�O?
���끰����`M��O��':7���4$��'l��M�g/X9���j��Sr�
i��I�*Jv`�կO���4��<��9X�Op�J��H8d!��rO��G��O���OL��O1� ���*H._B ���l�%�>��h��U���T�h��4��'�>��CX1�H�ڦ-���5�ԍ�6�i�L7M�p7M$?�g�2٨��#��D�=�p�8U���M�`$#��y�Z����˟���ퟔ���H�O�L��g*\�;�*�c㠍0����N|�<�eg�O���O����d�ݦ�]�f��q�ȇ:
J
5���\�@|�شJ�&�"���R��7�b��8��Br0�$��y"��Q(j�t(�C� I��`�Vy�O:� �"��q`ę�`��,�\1�'���'}�Z���ܴp�������?���N�Y�ꌻ;z�p���N�66&�q�"��>YӺi7�6-�j≹{�X��7�җS|���1�� $������9u.^�"~А
�B+?��$F������?����,�R�01��q��I<�?����?	��?Ɉ�)�O�u�b��	ʦp��>\�L:7`�O�mڒ~�x���ٟP��4���~�g��<�d��p4^��#���<Y�i��6��O�dKw-`Ӭ�u4r��i�����jʑI�P�
��g��TP��^9����4�h�D�O��d�O���=Ub\�"�d��R"�{W�8%'˓�����j��'%R���'��=�3
�.C^�B�Q	Z.h���O�>鲺iD��6��	ɡN�mr��ˊ*��СÚ�k�D��!�&M�,�h�N`�pA�O	�J>�(O�L��m�J�����	i@50�A�<���?���|j(O��m��6v6@���v��&���)�N�
@�)M��� �M���F�>�6�i"��e�ƀK���'�4�0��p\P���
�Ga�7�&?aE��=��)'�䧰����N�*i�s��:O��K�#��<����?)��?A���󉚢-��Q��"[�����Caڠ�D�O��YȦ5�!o{>��Ƀ�MN>�&N�:U
��s�B�h>�!��ڵlb�'�x6m��)�<eL7�!?�&_�U6����;󔴣Zat�0Ζ (���O�	@y��'LB�'�ꏶ
m��sG��l�.�{�M>�R�'b�	-�M��A����O˧#��%�5���7
�,AE��8�O%mڷ�?O<�OD�Qh�$G�.8|�D*~�1j��Fi�����i>��6�'_|%�L��O�xĞ����C�M���p��ҟL�	ȟ��I��b>��'o�6-V�6z���k��g6 �q�<C������O����̦��?Y�S��Xߴ�ؐeM(�.U2��S<=Ƭ���'S��J�{4�6��ؙ2.TG��$)Ly�B ?Q�0)%N>BަA�f��y"U�|�	ӟ���ܟ�����ȕO���!�M�(����x�D��w���˷��O���OT�����PԦ睊k�(�[��K�{�0Y2���GU�(��4K��֩>��i+3�27-�|�u�-r(�����U�%�P�K1ni��"7+�	KB�{�	Iy�O�"�;T�6�X��`f|e����/��'�b�'��ɹ�M��E��?���?�GJ^�q^ ��ԫ,�d��A����'W��a�fgjӢ&�C��Q�df�*�(*�e�A�6?9U
(n*dk���G�'c)j����?�r�T���!�l��h����3�Q;�?1���?a���?!����Onu�V��-I��R+ �vIΙI@��O��o��h	�'�*7;�iޡ���V$��Pp��?>��Cp� b�4}��o�Ȫ�g�Z�"}}h��柪RV��k��q�`��ш��`��h9��<ͧ�?!���?)��?i���5H�T[�.��f�4�������ha��ߟD�	؟�'?�� v�R���
,\bIM�5�ΰ!�O`�lڅ�M���x��T��� 
���R�vV�	��1�@�f��u!�I?�b��d�'�BP&���'���Fl��.]p��τ7� tQ�'�2�'�����4^��۴K�-��m�D	�OJ%�Ԣ���!k��̓����DJ|}Bs�Ʃmڴ�M3������j2Î4��¡e��J<�t�ߴ����x>������OB��]�2��JI�70Z ���$�y�'�r�'C��'+b����
�p��'K�'eF�"B n�@�d�O����ۦ�P�Iyb�p�>�O�Pc�Ɨ�D��Bd[9`,Y���u�ɞ�M����2�K�-�Ms�O�P㲦G1n�L`� 9#6�*�^"iNS��RQ��OF��?���?y��Z]$�4�P�"�l�Hg�S%0bh���?�*O`�mZ%�'��P>y�m�yb6�C&"xBx�3?�G\��c�4��xʟ�5�� O�֌��L/����� $�x�M֨b`P��|j�"�O��	K>)ԋ��H��D24���9��C7�?A���?���?�|:(Or�oy�y���8p'� �H�vK�QS'	�柀�	9�Mˍ���>��i��lWF�����@!�4Bv`lӠ�o��]��Lo��<��1����� �X*Oh�1�HX�gŒ����*��<O�˓�?9��?i���?�����1b�9�E��� �5�S/1�@n�=K'j��	⟨��g�s�8c�����$�?u���MB; �t��s��L��!�O�O�����A�>�P7Ma����g�$F���m���gp�8J2nD�Lf��r�ILy��'�"�Ε��5�e� �9�t9�߮I�r�'R�'U�ɾ�M�񡌜�?���?��_&���;f,��S���'E,�v��v��O"O~�(�V�x�D-�� ՈR̂ةE<O��$� dtx2���Pn�˓�j�!�Oj���fH��P�ݶ"�v�����T~Q���?����?����'�?����?�)�(�����b�8!��D�vmQ�?!��iږ��'���'l�]�l�i�咅�Y4z@T,�!�X�=��$���I��M[g�i򩎹d�F��؃��%���$z��#U�G�6�Zae��\�ZD&�h����'���'�Z֛&�D="I��q���+"%Ѣ}S���Mv��?���?	I~Γe���
А5�T� %A@t��#E^�L�Iğ�%���"�zR��z2�H
l��C��A5	S �;Ю> �ʓ�4Mِ�O�d+J>�(Ox�0��	+J�Y2�D�:?�<qr��Op���O ���O�I�<��i�^�1��'Z�$h�ib)c��Ǻ�#�
�=���Ʀ��?�4Q��i�4:�B�i�T�ʇ�@�8��8�l�-.z�i��6s�������������/g�S��Փdlׅ*G����$C�0���P�x�X������	ߟ�	՟��F��<D�X,��^�':-3éΑ�?Q���?�3�i��1r]�dKݴ��I�8�+H��4�[�(X�%)����x�"q�V���D��czӄ�K�(���,��9s��`��}������4�|�D
������Or�d�OR��	�\hP*�^�j`(8��ƭt����O����E�.s��';�S>uS����/:�j-"�Ȇ�:s�I%��������S��lA�z��a��?	��9D�A�0�V �
R?2����u^���J���k�	�,{&RD
R�pbe�t(�+)���I��I۟`�)��Wy¤c� �32	��bG���������$;�����O�!oZ]�W��	��M�K�q6!R�V�gϦ�ڶl��2�i��h`ֲi�I�9����O�xM�'Z���h� /ТeI�dZ���Z�'��	ӟ���ڟ\�I��H��s�����ݞ)�F�+���U�^�avNq�H�R"5O��$�O��������<�jI3�P*�� ����-|](A��4ye�&*&����<o��6�g�X2sg����bfhK�Q8�zF%q��� ��f�r��j�I`y�O���&(=b�/�ɚ!C0C*J�b�'�r�'w�
�M�W���<����?�K�<�Y�C��'��Kd�����'��L��dӊ�'�$��G�|�[u�B'\r��`${�H���U,ĲD�X�	I����t��O��A�s��E&4f���8���^<H���?���?���h����%wfha�j�+n�!!`B[������Ǧ#��`�ɯ�M{��w����U��
DZ싓*��P�Db�'5l7��˦Y�ڴ�:-�۴�yB�'���x���?��e��5�\H��Y�2W�`�w#�9r��'S�i>=��˟��Iʟ4�	;I��� ��|��/��!�ݗ'
�6�90�l�d�O���'�I�O�ܣw�(E�����ފO�4��vE�}2�m�j��Ik�i>��S�?Q# E��Aqa��^�tX�@W"m���h�iFy!J<]��}���Q�'��g���ihګ>�vU��ڀ0��	П��	ߟx�i>y�'@f7MF�?ST��]��\����M�e:i��LYD��Dʦ��?)R����4u�ijX��׃H�<6�2�nƔq�.(�"��8]ڛ6��8���
U��T&�_����SEM�
���k�f���W�c���I����I矘�	ß��r/��qs������L�P�Ӏ�V�?!��?��i� ���O���h�J�Ov���o��* ���n�q�e�X�ɋ�M�w��jVN���M��Oz�1���"v$��bF�5��D�,M�~�(���"f��O ��?Y��?��1g��)���R�H��55B(����?�-O�lڭ?a����@��X����k�2l;��M�\I�k��U���d�Y}�Ju�8���F�)� *�Ӆ��b����9j�H|;h=%h,ى6[�w�|��|b��O��O>���Nv��3c�ԣ-�%�'CP��?	��?��?�|�+O��m�(4��o̶|S@�I�(Z�r!I�h�џh�Ƀ�MC�&�>AѴi�0���üvŰU{��V�[=� �d��O86-	���6�#?9�a@�mކ�)׭��d��w�>�Ard
r���q�Q�J��<9���?����?a��?.�
�s��0J�:s��$��Zs(Gߦ�z�A�矰���� $?�����M�;iD
e��T�+d�P�7�H�n���c�i"�7�Y�)� "L��l�<�� ��p���f�g�����N�<A�iD�FkH�Dʫ����4�@����9�����_;���H���H���O����O�˓52��Cߠ���'/֋R�b!
�-�v���K㬊��OBu�'[d7��ڟ|%�pj�D�>��a䛌/�Q�1?���ַR\��a����']Z��$���?�QiH!+�)B���Ӟ�S����?i���?q���?��9���8#C$
�����\)_����M�O�Po�����I��Tr�4���yW/I%�G�#��a�P넩�y�&x�ȥm��Xʓ�Ʀ��'��9�p��?1Q�&�X+�H�7#@�x�)�
Q�Ii�'��i>u��ɟd�	�x��u`l�%"S'�zj� �C3�9�'Y6��6���D�O���.�i�ODk#�����T��on�aKvmLv}"*o�l�n��Ɏ���53+�!�D�b8@q��ayH� ��̡8�ɶ���a�'<p�$��'�^��!���Y�v�7R�"�'y2�'����S��Cٴ`)���sW�-��*
�o@X�yQL?�P�2�u��6���jyB�'˛��'b��ach�!aM´�T�?���:�"I 8i����l�� �h~���9�@\k�����T���9o���T2O���O��$�O����Ox�?�1�T>y��*�������� ޟ���ß��۴v̧�?���i��'����A��<#%$��Ѵ������'���+�Mc������՛ƙ�Lr�\{��Rg�!n��%���2c��y���'l&�|�����'���'^�!RuJ:Y�H tR1�䉺��'��^�@�ݴ=�֭
��?9���$5�Cp�tf��eٖv�ɣ��dM֦уܴ�?qt�铝7J�`��F�gy\�AP�E9n`4�ɳ1&!�!�6��擦cJ�l�k��(�e�0^��R��cY�H��ߟ�����)�cy��m��PK��D�^W�<��+�/	�2-�C�-e�L�D�O<�nd��8��I��M�t�ʟ5�̹`/Ч*��QAA�	:�F�'�Xɡt�i~�Ir�^8�w�O��,��s��]�R��`4i�B�!̓���Oz���O����OX��|�qMͅ>�:�7��jP�������V��x��'����'��6=�
���CӦ+�p���	k���g��ʦ��ܴ�?�)O1��a[��v���$g�����r� O�6B�?N�9���'�$l'�<�����',R	3�F�Fܫ2��@SS)ޟ���֟��	ay��m�6�D��O
��O�D2r�#G\�8�3�����ۗ�+�	����O7M�O:ʓs(���A,M36z󌐩t�
5�'�f4�OMjq:���-�̟:e�'���@��J?@���vN��:.>	��'K��'���'��>��	q�>D���,���Y�Ϙ_cq�	��MÑ#�1�?�����4��)�w*Z�V�>9zao~<[C�O���q�h�ҕg�86�!?������ܩ�p`�)]�9��}Cwj֜'�ҡ I>I/O�	�OJ���O2���O��sY�l���Cϼ%Zl��FA�<�պi:&��B�';��'�����	�,�`�# �UJ.� $�Aky�'ᛆ�'�)��_�t911f�OI�Z�����HVb\:>L�q�'$fQZ��D����|�^�T���M�x�$PY�.�+d�R�)ϛҟH�	ß��Iȟ��Syq�����O���HP�=��a��8R1˔,�O�unZ}�I��ɣ�MKҼi�b�ѦB��M��JoF&a���#bՆ���i��	d��Q`��O
q��N��@T��37���=t���b��e���OZ���O��d�O���*�ӤO�<!��8	�Բ�ᗼ$E���P�	 �M1��|R��x���|B�4@m��3%":�z�p��$�V���ٴ3f��O�d�i��I 3���c�D�2gF�s/9bd�R��?p�g�~�Iuy�O�"�'��P
o���6�^�)؀�������'��ɜ�M�ANɷ�?����?a*�X�i%N�u粸�aUq�HM ����0�O�El�M+��江(Hk�dP�p�n�f�� 3�&�6/��ML2�p�	�f��i>��Af[=��I�7!8A���.D�a1~�ؖ@֦^����E��d�5��`�w=݊�Z
ui���.��TX�-����o�8�%�R7B�G�� �E� �UBmБ��O�8`DHI!_��$rs�Z�FHVQ��E*e2e�nO�� S撶b �A��U;Ԯ��C]:q��R>M�2�kD4E,%A����&
���ڥX�< P�N�'�0���&��jdM?^�c��B	ܯL��D�Ђ��X��3&�?)�8	;W�E�-�&�#Ff��s�*,�d	�y���"�>�-O�$.���O�d�#M�8�"�۹{'Ĭc���k����#���O��d�O��+�b���7������̡V����6 G�7�<#��i��	֟�$���I֟ 2�q?-،Rh\*�� �a�O�>��'��'��Q�,F�����I�O�[Ս_e�Tj�Ǉ��D��EƌǦ��IX��ٟ��ɉ����=� $}�"�m�]���N<E���iN�'��I5<�
����d�O����(8@�U�E*�W�Z {��]�a(U%���	��@xЇ@v����$���Z+0,K2��(]A6}�fC��M{/O�Eۦ�D�)����(���?��Ok�/��	SJ�p��M�AG���'Q"�Ŵ�O.�>����Rt.��S�n� ʙ8Yh6m��A��m럘�	֟��Ӓ��d�<QU�.L�^���\�u]�3��3�&���L���d3��Οt{d
/G����6��q���M���?���Ie��9�_��'B�O0��iQ9��U�E�Y3�BE�i�����O�P�Q+}�П�������hT��X�r竇�h6�hb�直�M��(�H�"]�\�'�V�X�i���'��$S!����K�:�$��%�>�H�$���?)���?�/O�qʱ�� d�@�>_J�8��CP�Qz�|�'������%������dz�'ì?������u���c��'M��&�T�����oy��'vv&�Ӷ-��z�M
Di�'*Mഐ4�a��˓�?qK>���?�����~�ݵnAШ��jǖw�顳K.��D�O��d�Or�A�h蘥R?����n�Y�4��O?�	��A4�� ;ش�?IJ>I��?�6���?yQ��e}R��{&v�rP�ƱjW@1������M���?1.O``D}��<�s��8�`Č	Kc㗭q^�p��
9��<��A#�?IO~B�O�
����'g��x��
B�DQ�4����Q$n���s��Ia~�(�d��ae��N���C����M++O>�3���O��%>�Oc��Шs�Z,;r��,o���M�G��f*e��7��O���q����}�i>����3B~L��ɺ:���j��Mk���?���S��'R�ЍZR,��ѢӼgɞ�����)�x6�OX�dy� 
&��O�i>i��G?�&&�#rDH�f���h�y�̦���H�I�������Mۢ�Q�4�Ơ��F�o���㇞ɦ!�ɼe��Ŕ'�L�'��'�*x�@�-b)�xƧΖ"�;`�"�d�"R�1O����<9�n�45y���<���SR�E)̀���O��d(�	ԟ��Z3T�"R
���P�Rǔ�[�qlZ�%��b�`��Yy��'vR�KU؟�-s�L޽#n��	�ʊN�&k��iB�' �O��$�<� ͦ�[$閅l��;�c�L2�p2�2�d�O�ʓ�?q&��9��)�O�2�#X���=Z`H����{�k�ݦ�?�����w�'$����$�~t�&��3coI��4�?q(O��D<?
ʧ�?)����}E��)7�@�N��b%�/"���&���]y���O�L O�61�"��8M�L��J�/P���Y�� A �M;Y?Y��?�A�Ot�u�ՕM��ix�E
��``W�i��	�,�ɱ��'��禡���W�j{J�"��	�o¬�Q��oӚIaFM�ɦ������?i)I<ͧF��M���?�L�f�&`���i�i��'��|ʟ��O��Hƒ>#� :��1[��-�w��O����O"牉W���&����p�}�蠃��^�WO"$h�Ⴡ6� 9n�ן�'��r����O���O��q&B<`X��x��������A���T��"�>1.O��d�<9���'̙���\r톏9�4����Ht}ҡ�y��'Er�'r�'�剉9:B�#��!Vx5�1��y�f��������<������Oj�$�Of�Xcn��J�D�Y��6��t�I�W���O��D�O��d�OJ˓9T��)e8�깂COB%���b�T;D‌A�ix�Οl�'yR�';BHD�y��ޅZ64ʆ�nު���'��b�H7m�OB�$�O��d�<�cA7����֘;'C��@2�Z�Kf~�jݮ �d7M�O���?���?ib��<	-O�e�f����-��B&^��y��c�y����O"ʓ@���a�P?i����D�=f�TG:<Z,��"Z&����O��$�OЙr";O���<9�O[<5yP�%P�d��iتT�lZ�4��D�|°�n����I埨��������;gC�)}�r��V�D�i���''P$0�'�\��<i���bA�T��S�/܃]i���ȓ��M#'I��i�v�'�r�'l��O�>�/O����J/|T sf��1	t�#��֦��Ю`�T&�X���&��I���0?������T`8���i�R�'��˝GlR����O��	�	h�������Z�E�'�6m�O�ʓ5OZ��S���'p"�'hLrrN�d��4��,����AD~ӌ���eThh�'��	㟜�'�Zc����|�*Q�ä7%���+�O� (!?O�˓�?9��?�.O<U���Y��!��L��������>�����?���Ә��'&j��@#Zv*�A��<i*O��D�Oh���<��I�@2�ɑ<O�|L���/% `< ���]0�'+R�|��'*bN�/��ɗ'M�p����#C~ 0ke@�>���?�����$��q�$>1Q"��j����6f��$ѓ��Յ�M�����?���0�^h�{��I�f�3L����B#�M3��?q.O"0��D^B������4�"�j�$��W[L��sO<���?!�h��<�K>a�O��䋑�D�Tm}��F;G�)��4��DH764n�����Ot�i�c~I�0U�uX��Jw���S'�M��?1&���<�L>���  ��bc������q-�L����v�i� ݛf,r�.�$�O����|H&�t���������<N�(IvL�1���޴O6$�Γ����O�R��G��� P�[�u_��9 m]�7��6m�O��d�OTt���CX�ן,��C?�Ղ͞?;8�(�a^4L*Be�e+���%�Dۓcr��'�?!���?i��ZQ� �N2m�8��C��'��'|��J&8��O:�d&���ܴ� m �p�f��+��H ��BP�$�1aa�L�'��'""Y�02�cɉ�th:�,!N����Ou�|��}��'��'v��'=h������B�P��RŐ+ ��}��(��y"\����8��py�`
e4�S8=���'�^�8X
�j�f[�_�^듻?������?���N:���EP�,@3 ��I8���֥�7�( 7\�T�I����xy���$~7����F��5Y����ܖR����L�ᦹ�Iv��ꟼ��hˌ�	t���!"f��he�Xz��S+1g�V�'�rP��
�����'�?!�'*f��R��5O���w�ԆLI�L�T�|�I��`�I�g#���f�	GB�	�&�ře"���,�w&HΦ5�'oPY��y����O�r�Ou��2{�u��	�F�` 0G$����lZ��0�	�Z����~�ILܧ8$���c�ݏ)�0��'-Τg�Ԑoڑ[3�9��4�?����?y�'[?�O��0Wo��6�>�x��*��`��O��q5�YG���OzrA8�H�"s��:I���Z4�`7��O,��O�lq�"�l쓊?A�'(���H�{�-��X��쭪�4��t@��S���'���'��l�sIж<�yv$�����
��k�,��� �~��>������c�0I�< ����֜:'NR|}⮝'R��V�������[y҉IAd��H��W��stkT.)<�� �Iן�'���	ן�!��EL���RȊ�{d|��wE� �H�	my��'S2�'���;F|�O������~;}�pz�M�Oj��3ړ�?!�)T��?��aĬ yj��1
"^�� p,��GV��'
�'$�X��a&���'!y�M�rnY-AT�\�oH�I�Z1kӾiўp�ɐK����	韰�PW5�e�J�fջ�Ф^��4oZ� ��lyR��=+c����k�٣sR��@���ƅIc!Z�O��d	)�L��'�T?!����n�0A8�N�t����FhӐ���O�P����O��d�O��������Okl	+/^D�S�L	H��h�`	�(���'}Bm%�O&�>iH���:[0��d�-L7�KB̝"�K B�s��cG� �|N�i-�
��]qǀO�DP�qpKV(hF*i��*�Ua��
pI�I�T%Y� ��T;R�Z\��@�ץ��By��j��H�9I��!$�	dq�I�&^�<���{��_<�H`�%\�~�������X14�P�<@�����$#�@�T�3�� B'Y�j��!)s��DdA��	���e���A��hI�(C��\��A9Cж`����?���?����d�O�擓R���#���W�<2�D��o ��Y�B�5"ā��;U"؅�FG����O������H�@�"�$<ߠ�;�j�y�lKcL� L�����9�衱!����x�U����Գ��\�������y��d�OL�=)��DkB�Z4�S(r��qQ6n�(�yR!�;oܖ�Y�H\�R���q���'꓆�LJ��'!r─h��:��I� qC6b��'zB�'p����'3�1�����ڱY���+$�݄'t�7��3x��G��[t0�i
@�x�C�g$�Q��h@7qN� ��i����.��6�|y���3E��u��CnD�	��'D�{�P?z� p���ߦ?�z�y��'W.�3�:V���8Տ9��ě�'��7��^dJ�i7��f�����ޒ\e�<�B�y��	�0�OH
=)��'2x��AL�,�����;(�rЈ"�'}���$a���C��G�`J3��O��n����D������Qل���c���	�0�`�(�gJ�5 ��Q$Yq�O.f\G��7b�,�%�1!��́J�<A�K�Or��#ڧ�?�q���n*�ې��U��,��%�ȓ�{�ő-��Pr��11��	�HO�ștBʸD����1�ȭ6�,�Ĉ���e�I���	��Z��G�֟��Iɟ����}�a+х+,ze���Qul��W�(���ɑV��ӠM�+�<b>�OJ�RPLk���
qA���4�L�7�����O�HIC�3����N�8��6v��0$�O�QF��yR.O��?�}&������(�FuS&�ާa�8���9D��Cwo(s��d��!�)AX�:D�*?1��)§m�vdAP&\�=��ݣ���'a�V�H���2����?	���yB����d�O�"4�,�"���w�4FОx~���Bb�)"��z�͝�w
�q��	�-P���SHIu����W�s������B4	�J�P���-�i�牵�"Uh��
�cj��Ə���9� �O����O����b*��M���4��d#/T�iu�sФ��]� ��i �"+���D�<)���"?��'g���R=a�@{q��sFɄ�%�r<O����'�"?�܁s"�'{ɧ� �加��E���RE
V�����')�Q:�Bj�_��d��C���4����p<��Iݟt%���M�6@݄�ġ߹ U"�R�G!D����/�=7�DH�B��4^��Dy��#�@iش��-A@��8��MrvLӗR�$�<����QS�f�'-�?U���O� �CٚqY �aH��pV4�B���OT��.��d#�|�'�Ȥ"�T����)�#&)[�M�����+�S��t@�y�EV1X�Y���;�bħOl����'Q1O�\Њ3L�3[Z$3#&�.�13@"O@ӥDa��u��$�!5�$=���'�,#=���W(@�8�AD�(�
S��I\���'�'��RQI�.Z��'T�?O'n���x	P#��*\�i(�G�\�1OP�I��'�t���A�z>�$!R�Ɲ5��x�{���<�f�ųUb8�It�;�&��V͙$�'�.���S�g�u5����΅��J��QE��'V�B�	(�i#d(�4 �<HJs1�����"|jC��L� ��cs�A�� B�ci��;�?A���?��'6�.�O��$c>���˕8L�Lj�JZ���@ �
��pB�	 ~�k5�X�ɻ@O�$i�e;��K5&B\�<�g�6�*���$:*��#�O�H"A�V5�-�B8�}K"O��EK�9b�iS�P,?�$���$�S�S8���i��'�0ˢ�E3�D�V&^�i�氱��'���9lnB�'���TsW�|��Isw�ad��\@�Qf�W��p<�E �D�X%j9B6�P�Q"����G�#j���	�AaN�D(�d¡p����Y2e��Hó*E��!�Ĕ8P�le����F���r
R�:!�$KǦ�f���hM���퓚{12};�g1�əv{�e3۴�?y���	��E�B"V�	�p �L�Nip}���f.��'�@����'O1O�3?A��7�Б wk�$@����E��V�=���?iy�%HNc��S����Yc�b'}�'\#�?�y����	<d���Q傁kcx9Z���y"��,�P�Ν�n����[��0<�F�4N�rAXS��[��5
�� f��P�ش�?i��?�Ѫin����?i���y��7iL�)��9�PaHU�	o��dp�y"��<���gy�B
]7?�L�����<�`���5~I��O�a�@�$
���<� ���>�OR�a��!���'(�K�<�6"O�=h��/B9,�r`F>!�Z����i����*1�4ڣ�BjXK%C�o �Z#�͌<B*�I����	�,�_w
B�'^�)ǐWTE�W$�k���C�_�N��FO����_=yed(ҳA��]�\-2�*�a�!��=y;������z箙&��>G\x���'�"�|��'�B���-y�>4�6��F��AK��P�J!�P�66�]�c�Tb��݁�Ζz�1O4 �'���4,�RqHش�?1�\v�$��F@v ���w��5q��a����yrjA��?A����ԢMD����Z�N�<�uB¼I�/X����h�d��	.�}P��
�H��f�Ɉ���L<Q�J ��E�r�x`K��'�L������a�[]�n0[Ө�� N<(��_-�]�c%�.6��
d)ѩ9+���� қ�]�W��<��@�b�$�jD^���'A=�'.nӎ�D�O�;v�	�9��q@���v���FQ[_��I���џP�<����<i8l$���خ$����Ѭ 5�~&����E�;Pg�d�t�*�F�2iR��ΐb���R�k�+0��Oz٣��'1O��`�	 )R��M1����4���"O��x&�Y/WV$�KV��R��E�P�9��|�!�I�~�@�#u�'HС"V�S<<~L��4�?���?Pm��
zT�J��?A��y�;W��y���0��c�$��j�y�y�����<iG. 09�/@2hs-�/�U��N���	9QPxeS�������3*�!o���<�s*����>�O8,�HJ�c,ؘxRlͭV�hp02"O��e�ݒV"�P����xp�r������ᓘ����'=����ꞼOk TB4���}�	՟P�I�<\w���'���#\��S�J�P�j���H
�mGJh@�O&q� ԍr���C�a0C��-&ܨ��1��R��j����b��q��g����f��5�O$��ա�9Ybq�6 �m�vQ
 "O��7��n����AR�s�(�*�u�O��Xs�i��'�yȦ(� ��L�w 	B\����'��d	x��'���F��!�&��fg�i86|�`q1s:Z����O�a�jS��'��A 臶����"o3���N�Y��i�k�(m�u2f)�p<�c���$��WJ�Q���ѧ�Qa^��ǡ(D���(�!2�ޝ�È-N>����2�P޴)m0lH �r$��8�
��^��<��ţ.���'-2�?��V"�Od�Ӏ/�P�\da���k�H��� �O��ć�'j���4�|�'�~�b�&]r�-(�
W�8�~�K�D"�9�S��=.������?��㶅_]���O����'�1O�xC��$zB*q��n	29_��"O�8���E�1R~�Ň�
O�웶�'�"=1�Ê�0@IWD�Y��tQ)�'p��6�'���'P�a���+9?B�'���y�f��qΉy��L�7�"�s��?^	�'��\z!�$glџ(`Մ��"�)���TsDS�m"[r�^�(D�qAA�B��>1��AV���$�`֘qn!u��E��%�Lfum�
�M�g�8u��8T�������h�&E2,_0��%�N�BJ�{b��OT��ʜuqʍ�vh�1�4���فy��I��M�%�i��+n����|�-���
p�\�
4F1�m
�xs$\3��-Xp�jG��O����O��ۺ���?1�Oqjܠ��	��u2eh�b�J�`��ܿ�BKaEW�a�Ԥ	��IT8�hr��� tR���/	�
�qǭ�l��p#!���=9�̀C��x���
a�Bْ6�BXդs���	�?�5�i�Z7M0�I���OC@��&������� �bLK�'�X�i�.V�P��YpC�(%�B̒�y���>A�yҙ�Į��$���}����o���y��T�t[ȼ�� �4|
�<Q��N$�y����f�N��kZ@R����)�yr����++��?)�a�t)�.�yR̟"��m��Dؐ4n��4Mď�y���<ߢ5�FK74��-`�����y"�"w~f�{������C�O)�y"�,��I�S���^V)��_��yңܿ7>�%h�T5m����W�7�y"(UZ{tX@�ۖk������y�����u�\$d%�4j�)՝�yBNr���3�Y�s ��0����y҆ʹ0A�:eHȶpFf���y��tE��x�A��	�Q����y��+w�`�q��c����� �y��e�y����`�~����:�yr��)�DY3�I�VȔ�Ӡ͛:�y�c�w8��g�L$oͩ���yBo]	��2񨃻s�&�j���y-q���B !6��l�7�ԏ�yB�D�
���5��@�Q.�yb��;Dj$a�cK. �,�ъע�y�eT7LK@0�͘�u`�䀴����yrGτ1и@k�o�.u��������y�٠r���O��g�@�E�L��y�63X�x"0jk�NX�U*�y�A�_j���w��!��ʈ��yB㕋9�6 ��_#j<T��u���yB7l�.���n�>h	,����:�y�
͖}<vu��8����
I�y��� �VT3�]�6��z��ߏJR)R���3�g?��	ή0d��k��0~���# �H�<	��.ԱUaK w���Çϟ��a�@_a}�	������~g�٩�j���=��������_���l��-6Uذ� b�쐅ȓC�脲O�^�#"�D5s��0�?��N�"��#�a�1� �"��x�aّ�Y�<� >��ܪ_�DY���b��1��BXh؍�=����O�Y#�j�64��B�%>:��)�"O�a��/�8i�&'U-��&�'2N�Q��tX��j`�����sm��d��|�B>�O��T^d�Iюļ.M�Aᔊ��""O��ǋ�=S��PP%��K�l	R"O<y����
4%���D��U���J�"Oj��q�J���APE\�Z����A"ON�	�͂�a�<�B�
k�L9�"O���e�#՘��̅2�z��u"O�� �%D�uL�؁��#:�0�8�"O�Z�O<�D���)f�(�"O�4(� ۺ:�V]`�`֦}�y�5"OH|�bb@��h�B��\��)ð"O�5�ro��a8���O�GU|P��"O� �t��L�D��L�/Q�e�"O�x���P��Tk��]f��	i�'TƐ����<-n���[��`"
�'ւU�'fT�9 �����:
���
�'�*��O[����3���L	�'�&iY��������x���'\��JG�@���n�4l2���'>�ld��O8=J#N��c��	�'��7hǊZ�(�i2�;
��4 
�'0X�,\�^6$�s�hP
���k�'?�Ey�@W��ʘr�G��Z��X�
�'s���w�P��æ,�$�*42�'k`�
�4J����ԓ{=`�(�'j�1���-:4>�%�مj2�`�	�'OhXb0�I�pM�K�A��dP0	�'Ȅ4��"ހ�f@4��._����'���zp�;ET!U�C�V�b1�
�'gN�j$��$(��[Ĩ��N���S
�'����1S�<uDm`��HB���'ʺ���îs�t��w�M�58�Y��'[�\�
��V��
��^�v�K�'��Q�*Y�%�В��S8�����'�X�9 �I�K-�M�Q���	�@�X	�'&ܘ��ZO܀�XPb�|��qB�'z��fH�	޶����%w�Z��'c��9�k	>�<h�ፁ�"EDh��'	nx!5`��Z�PA��,�AxA�'� ���K�LY��J�t��'��}�4� ��h�Cw�+hn@��'V�c.�	��`�d&^��]��}�$��আ#���lA��nC�	�wx���2D�g��_�C�/̆؈���9��!�ujO> H�C��-Ė�1c��{�U��&ۢ01�$[��7�����_�ΰ>��ԎN'�u���טS���!��G�Tz�$A�ּ��	���L�C�l�"�e��KFvИ���uN��b���/�)�����I����'WF�) K�6��'�(�'mٮ�pU��>�&��Ȑ��ܩ��!�>a�L۴ݘ\��bQ�L�~�QR��Y��	��D
t#/�3�Ix����9��N4@��ɷDC��x�_1hFP� �;���ʲBJ#s�Xy�aX
�#*=�OL�&ēp�� H��T�I�\)p�')���DA� �JlfJ�>���G�<��ݠCfNj�j!-BA�<I�E�/)��
�g�*y�+D�F~���\�kֈ[1��"�&K-��ɑ+[#05j����E�<鴏�L�9چm͞W"!���J�H��P����	�| �c>c��qC�Zd�a�+R'5��4B�%<��1Åی@����`R�F��3�)~��HT^n0�)�tB*�UC��8�9Iҡ*r�H�ቪZ����H�
�@�#�O� ���Q�@�j�=��c̾�&0 �"O�����
(I��]�Kk`LRq��p�@Kй����$♲�ȟ�	�"G�
�VJZI�" � "O4��&lY��Ы���q����u@R�hʆ��'� �Õ/����Ϙ'O�u���Y� H-9j�KHf8��'G�U�q�ʩW��@"�!��M"��V$���:E���
,���$���eIGj��%G|�˄A�=B:ax�-J8V#�yb+_$R��4 LrU-^�r���G�	�j�ȓ:_*a���;���I���U���J�JΕ�Wp��ӭ:�*$�ȓ>��Eh'�&��`��HU�9�Z��ȓT��8 Q��#!����ũͦ$
�}�'����M�6$S��3�eq�(�5B��a��O�b����"O�0ۣ�
ڰ� �� 7p2i���}Z��	%h_���A���g�A�A�
�9�� �]���ɟ<�X�'��=MqFU[��A�n�0��@�fL����oE�E^��a���p=�֌��w�@l˂)�?���CL��	7�,�fbӚ����-� ��&�ֲA\�Aȑ� )I�I3n�3R�ؖ$� ��|
	�'؄tj��ůMG�I��CJ�z�B�MI妵���	S~iKPGJ�u*��PZ���DZ�~�R�Q�w���X��ɈQ�(��Aʩy�����'��A��$�V�t`ܞl���8�!:Prz`��a�mGF��	�w�!�&�u�g¡1��$8���<)�
(sW̩�G≃*�Y�To�`x����∁.��ɀ"���&�<�$T��F�NN���FZ�Oz�8��DR�
��[f�Ϳ{�$$���c�'���
"�۷HTxf=�\kH>9�À5�|�'_RQ"U�=H˞��t�YoU1�-ь	?e ւZ�Ae����_%�̛�+ �OTXS'�7U�jt`"�
�]×O�7��z�	:�FuT���AM�z�	�źi����w�(�����;ɂ�2�q� ]��'}��cC�FA��3��^���eT2�Āj�#�� ���O��#�C4�d�����ɍ3�L=�1퍃E>6����ݛ~���䌁A6&���O�x%*�7]���SCJ�S�P�xQo���?�։S�X�$�9#�w5�I{!"�W�';ณ' C�]��Yш��P8BN>IQ��{�@�&;r��?֠s�`,2�� �E1�nPK��\��|���JQ>�^���'�򨑕(�!~��q�e;LE�g..?��6xBf�Ȁ�E.Ur�d;�cX�y"l��l��Γ	4H#@l��;}� �p��!�*J��u �"�$���E�۹no����EG5R�Ia�e�>yG�l�*�1�D��r�����͙%hf�H3�ѧ*�Rg�;���]�H|��ص�ݍw�.y����}��6��3X;�����/��GǾx��T*�ͨo&�CM7n���Z�, O��
$d-\���'J{�*��b��XCR��l�R�2
��".�9*r�:�O&��A��ڐ�D�8L)r�	w�>!Q�^0R����ğ\z��L�<%?Y���v�	�e��B�>8�"n#D�����>=t�J�lޅ� lNh���ɳw�xݴp����~b���K���4�r �c�! �"�?$�x���Ŵ3��y��ì_� ��BE�^M9�����y���q�4��㉄<�R�pA��>.���D@(�O�����)�$)ߒT�����mQ�Q�n�����J��:$��ScRL��b��A�0����+�	p��X�N�Q����DS0]���{�۶>��ҥ�'4�H�Ѓ���V!Yw��3$���K2*�
5|���Zi�Pa�.�V"X�9!)T����{^2x�<�S�%��S�� X���\z�<����7�A���$km��;�Őu�&oe���?�}��Ԝ=�������Z�����x�<�̍�p� �SE�a�6IH�h�6�@	�{�^5�s�LX���I������Ɠ"�朙�I�]�=�A	�#MW`�H�oϛ�x�~���H�T�_��`w�'��<	��U�ۘ'q�yZ�(@t{X�2ue�_���#�'Ή�sd�3;��#P�V� M>��#Q�����O��2�Õ�hI���dQ�ɸ�'�HHBK���(O�=H|R�r��K�axr��0w"��)��_�Vg�41��Y��yF�,y~E�F`K�`�>�pVȂ5it���'�2��F�R��D�5LO!b���[��� ~i0�٬3�p1"��5#�\yA"O��R[�3�5���S��Hj"OȰʳ	�=s��sc��{�s�"O�<k�b�����$.$����"O2�0D��0V���%W1m�%B�"O~�2A":8Hђ 5NB�@"O�%+@� � �Hc�"�2���s�"O�)#R�ڇ��A(c��77ED1�"O�� ����&���Z���>5`H� "O��#g�گ4q���<o�h8"Oh�CR �uV�y�ڧ\���A"O��XI ���ՠ�7x�v] �"O� �"3f��8рދ_�؀��"O�}��h�xU�PpQ��%YÖQ�"O��(�D>[¤�a�4�(��#"O�=9���7�,كF�Y��P��"O�5;�g�:DH��en.L�:�"O�;g(ü{|0Y�U��,70�5"O"=���? ��c���_4�К�"Oހ!@L�x�:݃��kA���ȓ%�d��I>8���� >�|��ȓj���p� A�b�\��c�J2����*��"�Ӧtց�j�JkB��0��Pp�_�-���b򇙌h�ZL�ȓ?�Ƽ�F���(��ځ�4M ��ȓ}:�TDIܓYG6�W��c}�̅ȓH��HeM�M�l��ȓ2��ٚC��@�i�4옅+�d��7J�\j����򨪴擺m��C�	!y�bqP ��(I��xa3c�mhtC�'.NHP�E�Η2�V��ga�$�C�;Õu��:c�p�-�4�J���'�\�6f��Z-~�"�*���I�'�<9���"V�X\cGCD'��đ�'Z��`n�b����ʍ�lc��
�'y@Q��ٵ;��Z���i��Ur
�'xZ��6"�?�����%`�����'i$4{��;D�h0
�,K=��Z	�' �� �iI�Wj>lS+ʺH�`y2	�'�80q��L�4�(<	׮ծ���	�'��hsO�[�� �-F�Y�l��'��UUhQ1W1<q���4t��"�'�x����4q$��đ#tB���'��`��C��)�L�g�J�nVu�
�'�j�ғ"C�A�4��C�
b���9
�'��]*�D�(Cfl���F��YB	�'����5#\	�������=��'D�x��^�QD�U��<�
�'�9SV� ��3t.�<t����	�'���#eı>���F��gX&��	�'��p�0%GWCL�!�팉h�,���'�@ē�+:n��%� Ƹ�b�J�'���i�f��<'0,�D	����	�'��X�.�-Y"ܽ�3�!,Y�	�'RDP0%�X ;�6���%8%�6�	�'����P.؎oj�`R�bH�"`K�'�%�ф���\�� �F��t��'�=+P��h$��b�)|E�q�'d<ɥF�f:U�5�ʅ
��!�
�'<������5��6w�K
�'2t�%�5w�2�M�}��y	�'b��v�0I��!��|d�l�	�'6�}z��X1l�.5j �S�f�4��'�(��G?s�$���L8KP5���� ��H�%C0m��UI� U_����"OH�h��ۍ^a ���,�bh�"O��:�gS�{	Ĝ�a�_�+�1"OD)��A�=Mcr�c�i͉"ɴj�"Oj1��nɸ*ݘ ���YZ�8<&"O��=@D9��I�7�H]ٴ"O�a�e, �gv(!���#C��� 0"OF�{�/�>Ø5)�ɞ+����$"OČ�!J]�S���"ń���"O0��F�� �2���s�x�zr"O,đ��.��AAAW;1����7"O����^L�`L�s��(`�"Op�J�k�B	w�x]�a�Q�n'!򤕀<-��жm��5����r���5!��%
Y(y�� H�d�F��.��'w�KBV��p6nɂq⨠
�'2P��pq1S��l�C�'jzG/S�7���c�6g��t��'B������ X��Ǥa6m0�'�R���9d�3�� h�օ��'�^]CB+ٿ=~�s)�,� t��'�졺��?~� |:C'T xRt���'��p�0u�xI)sDƟ^����'��	I2�@e<�d�r��*[�4i��'����'�+*��̊Rf�� I�Z�'9h̡�셒Lg:EӴ��FMs�' cG!/	�H8���<#V����'7`��M�T)�8��O�6-�Q��'�ڼhT���0�P�DȞ;֍ӷ"O<�t��0#�&Ŋ��M;�4�p"O��֎�,]�uS�J�A��"O挹���l�΀��nVd@z��"Ol����y:�MB��FL�"O��`� ��~x�Yp*�^���"O"�;�ٴ*pڙ�w��{°!)�"O��2c'S4L�� rU�"`��ѧ"O�����<�� �޾\�61��"O�	���Q�������8>��9"O���j�VlH`V�O;*L@誇"O�`�!C)r�S�J�(��IT"O��!�_`� ɗ��J�Z�"O�$c M��l06k(��y��"O�)��%�<&����c-�:��5"O�C��
C��dL@Q�`��"O��&�X?��#ҥZ�v!(�"Ov�U-Ԅ,�x!J���>(j$|��"OzY�"BH�A����-aT �t"O8�&�P�8����ˏ:Q�=�"O�� "	Ӧ!���q��R=I��"O���qN�����L*=
��"OtH�'�,#��9�')p�8T"O�I�FL�L|�[wH	}�����"O&�:Cۥs�+���i��@��"OX��ՌJ�N�v����ё�2� v"O���$�=���{!�˪^�P��%"O�����N�/g��bTDڂl��m1`"Ovi��(�2f���[`Iʯ�ha��"O�P��L��N����ޕM>�P��"Of����tB6%�q�LT@� �"OQ���/ x�����:=����"O4�E
U%5V�e��`�;�$��"O�u�g��L9$��pnފ ��$��"O���6Mכ@��r2Hvs<UB�"On���§q�ĭxlד%X�ʢ"O� $�3�i�>7G���E_�\M�T;"O��0���"`1��d��2~�j�"O2����"`�t�h D�y(�La�"O�9�>g29P�a���A:Q"O(@�Q�X>s>������*6���	�"Op�����)�$��ە=�Ȁ�"O�26'] ]�zT�#\{J���"OB�H����a�#E(4Fѥ"Ov��c- 0l��1$�.��2�"O dh�o��?�聶��A�`�×"O*İ��"/*ё�Y�E��X��H-�S��y�O������W7f�d�'9�yjĈ'ټm�f^-4Z\l�4/�y�#NT��y8`�L+;�t:����yR��;|M��ӡ��Cg���\�y�]�I0%I�`b�X��J��y�`Hm��Y+U�
2���u�F�yb�>b.��p�@|r��`� ���y��N�g��x���v6���k��y�I�a����G�@�Ĥ�Uf���y"�)_@�-PË��m�f��V����M��4丧�Ol����O�q\��r�`?=�*���'��[�i�u�t�K��ݣ�
P���/qs(���O� YD�)N��i� U`|��K�"Od�SQ߭0P�� �.2q\��X</���X8�����)����W���.q���M)lO��JM>IӮ�u>���"@�a�v(9��M�<m���X�"I�*V�6!�f
@ܓ��FxJ~r�b�;z3�)��"�{��8{ͅz�<Iu"�++}е�צW8e���rǏv�<��KI�:�N�¡˃5�F��y�<��I�Kyty*Q�,eL���s�<Q��O�Fk�̣3��P�2͹2�T�<�f.ߔ{{�ݲ�2=���a*�S�<1��1�DC��
^}P���j��hO�O����dI.7�@���JŒ�t"
�'^��Qg 
��֜`�6wd�k�')��!

�~����"�ҟ[����'�z�#�R�R�n	XG�ܷr� ��'d���v�Žs�Y��B���9 �'�|�����f� Y�!��!��'���`c ^fk�h�X,��'��ܫ�E+M��QbL8jI��K�'�v$a��(�M��-��]�f�ѯ($��Se[4\�*�P<-���uc-D��0���C����t��\D1"��&D�L��h�$���6�]M�� 11�*D���b+C	
�,�Ӯ�Q��؀J.D���D�1�~�+1i J$1	@�/D�A�����P�cU *D��G�i�`�@�*�!�:�K��(��<�C͖;y�B���ǌ*���CagNF�<qE%
I"P$���	��[�DK|�<!!�
}0H��Cӂ(EP�{�MHt�<�B�
S�rr d�&N��!��j�<��� �6��rE�98n �
�c�<���8F:�0b�������h��@c�<qc�N�7)"�B#�F�}.�����`�<!�+ݳl`�*��՗|W��8u�P_�<�)�%/��8�k�8_���2�b�^�<�a�  \�"��H4`)��:%)I\�<�D�C�a���f�vB0:�!I`�<)�EP�o�h�
7o���j���u�<�7�\C�����Q�sb��n�<� &1xQH��_��ᗍʯ��Ļ�"O�iC�A4	�������m��@�"O�][Gaڤ((X�J:-�<�3"OL �Re�j1��B@�Q8^�̨
�"O�Q�����Py��
"�\�˦"O���$�-aP�S#L'�p�4"O�dR���Eb�$�ʏN�Lpp�"O��1ド���	��D6ZȁU"O(ura���hS�����n-T�y5"O<�5���4x�L�p���O)d��"Or����F�<F�+&�O���"O\�wI�&�(��Ѣӯ8�Hi""O�
�ܹVE���c����#"O��t`�@�$L�#�Er<���&"O2�(d�$c}�C�F'p,��c"O�1��'M)	{84c3k��l�@�"O�uH�o�,_*m�/�xvh��"OV����\~< p-L6rf�M(�"O���1�3�tA�ʍ��l[�"O 	�֍á޲	S ɛ�w��<�&"O�,RclP�M����N L����"O�����zG�5y��G����Q�"Ol�Y����|�&�zU�F7 �r"O��ٓ�:'�y@N�frY{�"O��I���r"��`����K	��k3"O�TS���G��)��Ú���""O(Tb��|���j
�x�`"O���\C���`��m��h�p"O)ǃ��F��1���m�"OP�z��ŕQ8 j��@�[ȥ�"O�Ȧ�������#ÌB�xɶ"O�0����=|ހ�r�`�z&�a�"O�-i�˛�Ľ�D��(��r�"O��؂�P���h�E��
��؂"O�᪥č�wS�=0���:)�
TXa"Oޡ�W�W�q
F�R$�)�(�h%"OA�3O��KN�����`C�xsG"O�e��/N�@��@���f.�;S"O�q���2j�t]j�	 �=�"OPM£�Q�\��3�&�<��d"OR	K��,��Xa��?(W$Ii!"O&u�!f�<Z���nI�l\B� �"O�$Ca%�u7� �G.��]�4��w"O���K	(t��ҍ�h�D&"O[���$����mB��ey�"Or�`���?8 �س-ǭR��X��"O��1�菮9���уm/U|��s�"Oސ	��[2��ό#Վ��U"Of4�T�3�U�̋8$�yC"O��b�)B�Q4�~�`"O
��0(+MBe�1O�'��x��"O,]{�cC�O�0�SD�"o��XW"O���!H�- C����̀�94"O���,���+�f��(Z�"OF�Q��Ȝw�(A��iZ;�Z�"O���&�<j�lbj�����"O�h����gq�Iu�	.i�	u*O��*���%�D��AΦAR��'�H`�GꚺM�@��nX�7u� h�'�"�PPFF!mH�t�3]�Y2�'�iPcQ$R�bM�
 T��i��'$�(�'��e�$q#�b4$�9�'�,-����<�$�3��N�L
4�b�'�FP�7�Ō'����ま<��ܚ��� ��ͯ~��(s��*n����"O��kFb- ��B BT�YR+�"O"���6�xq�`N	MR ��6"O$A	��2�"��2.��Oj0�Rp"O4��3J?7�2!�d�J�A\�$Rd"O"�Vg����|�`�$X�\�"O�4�6�̬&t��y���n೤"OjȠ�g��<&8�g�D�h�ठE"O�p� �݂I�Ƹ�FF�����"O4@ ,Ķ~N�P��"�+�^��G"O��@�kQ!Gf��a˜TZfq��"O�}��N< �X[4뛟I,R�"O6�yD.�=�}���I񀔩��9D��aGC�kxb�K�m�`L�v�4D� 藃Қ�А�f@�w$D1�g4D��"��|�Q%fI�򀝈�!���kG� �'��&�p񕠇��!򤁝%��m�s*��R��9A�n�!��_-Z8���� O�N�9v���.�!�DP�"mF �D���/��df�ٙ!��4V�#��ԠSE�t{7 C�T!�I���A�c��7)�A�'
�"O=!�D'GKz�J� ܉.Z�p&�2.]!�$W�O���Y��
D��W��<O!�D���)@�ƫ X�ȷj�"_!�d�:$kf�
'I�W�J�+��%\!��
9G��#�BM��rE1�h��Q!�8c)����n���U��"k!�F�v�L!���*$RȺ�&<f�!��,�*WM�#]	|�`d��']�!�$��Y,z���.ׂ !�]�%��!���?��0DA�f�ڵ�V�%z\!���3��Y�eo](�T��텥Q!�D��#���G(=�6h�dK ]!�ե��`#�/G�8�~HP���"&`!�$Ksj���#��@M��/��ea!�DY�$��+�A��N���B���d^!�D��[3N�*��5b��L�T-�2*�!�$.����%f�!�U0O�!����C��s��Q4OeܕP���Sj!��D9�4��S*P�xu������`O!���.oYP��B��q���sa�mD!�$\��BaD��	Vu^��w��/!�!���#��e��wfn��J��t"!�dڨ�h�s�^� ��8�A��4w!�DCs��F���S͂Tz�M'�!�d�'z/f����Q�
	;E�$Z�!�$P'I��ZU��LpG<G�!�dI$
i� H��
��$�A3@�>!���Ac���g�.��W�	c�!�Ke���BF�H9W��1z����Xl!��W���,��;!������v{!�䈪d3` ��m�jn|XdM"}A!�D�+^^$<3�@�"m]�Y��N�~�!��DG?Y���]�#$�m�FdY$k!��Ҋ��PB��_<7�8���'1�!�$�V�X�ҭ��u�y�@���Kv!�d����e��?" �0q���E!���e%�-1u�|�������%D�!�$IP�M0��(�n��#��wx!�D�'h�2�`���LѼ-R���nk!�d���űg��_�dm&fۀbP!��T�&a�vi�i��	���*o!���H�� �C����ud�*j!�� *����S vB�9K'�[�)�H�W"Oh��܆�섢�H�/#����C"O(�p�gҠ_;��G8���:E"O
%�ժ�1K�myae\0dàɉ�"O q2�\>�~T�A�И/�����"ON�pr��:x��p�_�^���"Oa�sNC�)�R�A�@�7+zT�Z�"O�L��I-�Ҝ��̋�;i8!��"Ol�����UQ�0+!�1d�~�r�"Om:B�R�]��{$D<M�Ƶ)�"O��2	�
<�X#'�W9q�U��"OH��j��bx���w)�@8"O��2�&żs�Y9sς&o>}Ha"O���o�v���ط�@5f��)w"O⤯���8M���ؒQc�`h�"O8EeC��e��a��[!YQ�)�"O��چ*%�B�@%�_�6촜'"O��5��$�BܱuJI9N�>ؘ�"O����&�8qj<�/�1 ƺ	0�"O�Hk�`�T����Ө5аh� "OP���oY�*=�$o�)]�u�"O�=���Y,����QF����"O��.�I�1fh���A^y�!�[��` yvhͦ9X$�3Q �@�!���B@�b��><ZL���3�!��
��Xq�6�TN����b/A�%�!��G_ (*� ��-�VIۆk߽Q�!��D}�ȱ���78wQ�Ф^8D�!�$Q�������6�`�b#�!�$� +����(��t ����!��[�iETz�BW�*��q �Z8RU!�$J2NA~�1%���߄�XĭW�ct!�D�)���P#,���0�Nټp!�d��8b�}I`��8��&LPv8!���/��������u&@T��4!��C�,Ѡɏ)�
���O�~!��
�,,������tB׉՛!�D�%�$ố������k�!�D��/�T� 4��s��C(�5D!��1d�8�R-ŭ1�bE�ʵD-!�J<>����$!q�j8C��z+!��BG���S �V0Q2��Ro!�䉝v�Z!{*�jdŪ�@�aV��䎃ft\T:�/�`"��3l՛6�0B�ɚ\�j�*b� >�4�1��X�+IB�	!o*8Q�a�A����`��8"�B�	'8�L�y2D�
{I��(F��N��C�	�	Lt�S-�@�q�LC+}�C�:P���
�M�xw��I��2_�C��0{��C�	�:]�L�񯔢WE�C�I�[��U�sf϶5�ڐ��&z56�O���� $F4=9��?<�B�fצ.�!��"@��L�L,(<"х^�g�!�Ĕ�W�Lq3��A	��
�'�!�䖉Ә��G�T`��d�Jf!�_k`pxS
����
��<M!�DU�^�28�.�!�4�J�I�=!�dE�f�N��s�+���z�"M={�!�՘O���� cOF�c��R��!�$���X�I� )�$�
��!�!�Dvwr,�jR'=��i��Oǀ9�!��V�H� �	M�dݺ!)A��/�!�$Ͷd��	B+�,(�t�[���F�'�a|!["� �9(8d����ą��y
� &Dԇ�&{69B�ZR38�E"OԄ�tN�������cY5K��a��"O��:�ə7_���%B� ��T��"OB�(��ׅB�X5�t�����*�"O�B��	����L���R�"O�C�I��|���ŕ+|��'��'"��>y�'AF��XJꔒ>�Ahg&�S�II���OiL�a(�)ry���q�̊q�<a
�'ɶ죓�J� ���RG	e�Z�C
�'�v�Bcʙ�g��q���.�:
�'�07 �r_�qCE�/O�Z���'�`�4�ϩk�nI��֑J�ʤJ�'�Z}��A�9~&N0��
�Y�6q��'�T�h���l��zsHՓdQ8�H>�������Oߨ�ە�ȀV�
�Ӈ�d��a��'/J��7�'D>^�[��R-]ђ�C�'
B�q�F`+I�f.)e�2!P�'k�����*|�8���g�^
���'�!yƩ���e�P��9�''�X��1(0��G�Y��t8�'>z�%)� 1�l�{�d=R�}�������O���>�IP�|��`���-0�hȱ�K7D�����3��`e͹����7�4D�pI��?7dZU�d#
c����M'D��'c��6�t�k����~�~�Df#D��:�%�~��01�7>�j'N"D�ؚ�R9,�¬����8�`Xs�2D�DB�׿�n�d`Q?.�tLs�1D�t8&�[J�xh�,:-P�ؚ/$D���0e�=Jit����7qW �8d-D����
!Kti/�!X�l��+D��cC���&I�ϊ	>���'+D��c�N�Nt�"��]�
���&D�<ЗU7+�j R�D�$�8��#D�8a��99ئ���]�s
넌�ON�$#�)�'62�����o�f`�wdȫ9�����'n���2�-�D��ǎ��~� ���'Vn� a-�;O���2D�
��#�'����y%R�r�����V�<�fb�G'�L�R�M�|N�P�F��G�<�AdJH�̙+D��VD�XJlI@��\�<I�iȵ�L]��kА+�t2t����x��W�S�O�bV��"A���
�i1 �����"O��	���0�d|�E� �j�Q�"O`���`�o���r��ݢ,H��8�"O�劰c�vP�i�Vn��S.P�u"O��S0M��Z����,*D�"O8}q��V$�4O��^	��'�"�����#\hJ��\)r��y�I�O<�D�OR�d�<+O�c��`Ԇǉn�h���_8@ �Y��#D�<�E*G�<�NLP�Q�
Rsc"D� ��L�,�9%h��ʼ��!"D� [�C��uQ~@	�
։.��l2�!D�xʄO�1Y�T��R^Nuz�M,D�|13�Z+u	���i��xDb��(|O���yrO
�YLν�A&i��H�C�W9���hOq����J^ �q����8>�|P"O�q0ƄԬ���d��ĩ�S"OY�&l$:����+����"O�xDD�v�6 ¤�P(��I��"O��)􄑶�����ډ|L�q��"O.IY���,E��6f�'�"0�"(��0|�Ao�8w;��bC㖁[�ɳ�*�q�<��O0&�04����'�o�<� �Q@�۠W�t��ӑ{��%@ "O�ĳ�$�`�|�w�5zj�id"O!ؑ���"�.hJH�v��tA�"O�h�gI��
V1�*�=і%�c"O$�Ʉʜ�u�\�*��m������/�S��_]sʨҠl���r-�B��%!�$�;H&���F!%�8�Q�
�u9!�D�u�R���E	z������L5d�!���! R�Qag��]�L�)]U�!���?,��J�N�-\����F�!�d¦g�T@1�"��:	�mE8$�!�C�.��ᣄ�=^5�6l҃�ў���y��Pyb�ښo�]� lS'�d�O��O8�}��+�J� 5/�)f�h�"g^&�昄�#�L-�d�Or���@�	ͼ�F���U�����ꕊ���/X�n���b�G�<!��P�O��fک	a����C�<�SA��4- �����p!��@E�E�<!��^�Q��SW��@Ul�A�<I��B<h���J���	ȁ�T����'gɧ�i/�	�O�N���)\�B��L+4G[WC�ɪi¨�Bj/t��J�MZ47��B�	?V��c,[����S5a�1KvB�I�;{=� �
S����A��:B�	qPN�G�hHl�e�[kPC�I�� �AG��Nbdz1a�Z6"��$q�$�q�	?j�D�V)(�j9�d�/��4�O���À�?���
��8�AV��G{��)��=֠�R(�?!:L @͞�}��O.��"r���:�`�:H��)a�!�d�M@|�N�+�8r�:R�!�D��H��M��@K�+n�ȊtÔ1�!򤑢D1�l��߂$Z���D�חơ��%���Ac��1~`��n�u�����*�H��%�ިi�x�Č�x�C䉱W�T��s��8~�jV�5y�C䉀;��� ��!Nf���Ob�*C䉡W��%���H�h7ܣ�Eݡ��B�	������_��L]�]�C��h�	�[(6�ty��V%m��C�I8S�ʉ�	G�5�����%^�qhJ��ȓ
K1��L&V�*�"��#\�h��X���xc˨Hd\��WQ��eRdp!L��	�wKHm�U��Z�j8a�PJ� ԡ���~L�-�ȓqj:���N�52�	��ۊ#ǘ��{�yb�� �xX�b� I��o����<�Fꇾm���% �.y���	Q"D�|���V�o��x���].���1b!D��I��JO���!N� �&�f>D��*��	�\���G�g�JQC#)D�P�b�ē�0Lq�"�!�Z|�eL&D��o^�n������� ���/�I�<��aϙj�nH��ƷP�ΤzԪ�D�'Ra��"�RF�$1tL^o�J[�����O�#~BC���@VlĻ炆�'�T����{�<��L�3ytr2VO@!��e�b�<qw��`pԈ���	�ø�Sp��g�<iVo�#\�&��v"L���a�<A%�=OL��@��ŗ2��0�t�^�<���7�&� `MDHY�e��Y�<р��  ܡ��K���V��V�	ٟ���C>A���)]�2b�W`�ajq�3D������0
�p�mI&g�j�Y�L'D�� ���#F� ���S��ؚ�B=R�"O�T��	֒@x9S�g9%�Ty��"Ov�*q�
22|�8�`L4nl�=�"O8�4 M9J䔥j�]�x�8%)"O�i@G]�{�:u�[�O����"Oƴ 䀏��D�H -0i30"OU^'Q
���ǧ�+�n���"OPt��	@49�:U�L� &����"OV�y�cQ>jl�hRR�@ ����"O�9I�E�#�8-����k� �+�"Ol�˙ f{�Q�gL�h���!"O�9����K�<� -A�����"O���ք�,_@08��B��<�1"O�p{��B�]�@���dJ��9G"O��q���#���E��^@ax$"O��Qp��� ��,�u�ɺO>{"O�����]�)���"Fܐy��
�"O2�A�D`�J���"G��X��"O�Ĳ��zĘ}��o��1U(y�"O�=�G�B;ZOR��p��6vG8�82"O�P+5�Q�!OHUJv씓{0 ts�"O�����n�y�R�ǜJ5�G"O�]�ԠM�u#�ċ >R���p"O�MKנ]�/ٚ�hq�@�s=��"O S�@���(	��ܷMʀ!��"O�Lz��&s$�DC1�\�w�&���"O2��P'X#�����<U�6��D"O��[Q��u�f����ͮ<�I��"OD��AO��X�.�1 4p�@à"O`2%�V���DY�9�����"O�{R$ %���C�*.�5C�"O�(Z�gC�Hu֍�ա�:X��`��"O8�Vd�/�����m\i�,�W"OVt1�[T�VQ�*@�k��
R"Oɐ��Tl��JV��`�@�ñ"OZ�b��ٳ�L�yCҷ>t�:�"O�z��̈́S�j@!�>54Q�"O�!H�]0��K��0n��њ5"OܐY�����B�OX�k�ry�"Ovͣ�@ ���œ����"m��a"O��
�����LH��ˣ*W&�(S"O�`��܃L��Ĺ`eǦTV����"O���k�.&����$0����"O���qE��w�x���`�U���;D"O���H��DҠ��ψ�c���a"O\H!�<<p���ytmQP"O~�(r!P��åM�E��u�"ODi�v!�y(r8�u.^��xr4"O~�!D�?|h�v��=0���"O�YÀ$�*p`r���b���:͢�"O A�
�
�f�C���" � �h"Otܺ6��:L�+d"�Q�,�"O�s�^�G��=�V��[��ͱS"Oh��䏁 U��1�`�3�D5r�"Of=ѠU:8,t ��/Z��6�a'"O��1�AQ rP� r%���g?�4�"O>8bql�(j��;��X�p��i��"O� Jd�̼S^�X���{�Ɣ�"OL$"�C)%)J�B�l�b����"O�U�V*	�*=R�ڴFS����w�OS| T�
87�P�C ? 6٣���y��.-��� �!lv�81HN�y���:�Z���P�I����)���)�OX!Ȇb��
�%[E患1]H`�"O� �`��$��eJ���GI���yv"O^�i֋	H�`�s�(�`a�"O�ufGUxl�tS;d)"�Qd"O�Dc�� �c�D����s�@��"O���� �?�b@@Gű�JdR�T�����l;�҃2�x�
�f��D�O�˓�0=Q�پ/ �L�΁$R������}�<�S�.}�<8ptΝk�Q!F�|�<��#�8A��a�� 6-���Aiz�<�`$ڎ)�P�p`�%����O�u�<�#���Y\�X��`Z$��aQ���wh<�UO�u(��@BޓQ��-Ё,��?9.O��d_�lì��u��%J ��'I�K��'a|B	�,�f���*���r�'�-�y$_�T�A��Ą ;����¡�yrP.1`��h�*ht8� ��yB�T�?x)x�P?�Da@��y"3sJ�@�ꘜ~`��X�$,�y���-�D�QiR9+	�$�U�� ��$"�Ox@�sb��
�b���5����U"Oȧa޴Y�h8$ �m�����"O�ͫ��� �p�+��ʂ�2 "�"O�\K��E.[� pV��/]���Y"O�*�1�| ����w�;Q"O��Zr�\58��D���["O�Tr k�0���d#�P*���D��r��W�D ��dY^Ȩ6lW�<@��	���y"�?/���G�5"�0�v��3�y�'�pN	鐌C�&i�ƌR��yr���h���}9�3��y��JpI��Bi������y��N�˂m�Cڀ��q�1�yr��W�L,s�F*!x��pjS���'@ў���<U-҆F�ЫVa΄���*ZI�<Qu�ہ��N%m�r�{�f�n�<q���i�f�ŖXJ�-��g�<��×�@N�ۢ���9����a�<�`g�Dv�}�ݐw�I�ƌr��G���O��:1)ǉGK��CѢ]O�(��'i�,
�[��	���0�DBJ>���?����O�+'Jl�*DM� �l	�y�,	��Ӑh�7{P�aW�D��y�ɜ��Ʃ��k5B��q��*�yB�i�bY�uk� q��Z%��y�� �P���ŏe���0
�y��H���	��Z �tH@���y��"'	(A�!ْT� X!�D���d�Ox�=�|��X�aA���
\�S/歙 ��y��[$���J�XO�B�7�6�y"���id���I\�5�G�ѽ�y¥Bd4��pK�E��Ɂǉ���y� �6+�f%�s`��<�*����y⤔�q�@�:7N�5D����]��䓖?���d/d���!'���P �&
��yBJH0�f��f��CWi��!�y�W*M9�a��dƼ9O�}��ȝ��y��[���#J�+�@�`�(�y���S!����R�/�>��n��yb�؎t2�q�M�.��Xib+���?��'j�x9c��n\<t�R�V�P��	�',ք��h��Hn�{"��T	t-�'$��+��O
q�NLQb��/L>J�k�'��t��cY7|���P2�H�R��I�'_t�������za�۶I`l�
��� |hpu�MQ���+
[�B���O��A��
�v���mu�J�)D�l������}xg�S����)*(D�h�����r�^`h�H�=�Sc2�����H�-J8���`��m� �D"OF4B"έiӨ�Jr �2V���"Odc�4
����c�ɑe;l��S"O�t���[�=
��x/�'$��ag"O��I���)������l��r�'�!�D�D����$˸j�(����l�!��8d<�  ��E	�-ۆ�Ώ+>�W�l�<A��@�O6e�UbSj � Z�aSo�z	�'���SQ 
�c�|�!�ށ;��Q;	�'cBEJ�	��|8q��£1#���'r6�1�]% ���	�Ro@� �'\�����yY�i�AĜ�^IT�.O���ě���U)��D.�9RU�J�7*!�d���0t�b��6U��� ���Q���|2�'���'����+ϾjO����I
gT�x��V�s�!�DY�-x\�h�{M�IiE�K?D�!�ă]L���G���fV��
+K�!�ňx�D��@�/DV��p�ʆ�!�N�
X���mF�O�4�x�4>p!�Y�?T6���iC'{Ji#tEF!;[!�$��O9�����7M�������!�dH�u��tphыn��ʵ[��'�ў��<Y�ęݚ\+PLːq8�HтD�R�<Ń�-:�!Kg'D#�i�!b�e�<)���ez���Ӭ��' b!��'�K�<���r�)5犊;�,��DB�F�<yr���U��4JE)�^��E	Wx�<i�=a�y��a��V��c��L�<�u 
V����7)�/� Ȑ�!d��hO�'Q�pB�PixR��jɅ�%��ܚ6�(�h�)��I�̇ȓZ-�ip�7p��E�>/C*(�ȓ���.L�o�����H�d��ȓeR�1�͉/N)IWf�7��9��h<w�Dl�FT�F���H�$��X�<��NĲ)���u��l�WeT��hO�}���i�Ò(7>
�����(�Մ����4K�*O�]:!E���Q��N��i!3�V��8�{fjͿz���bs��$ݚi�f�W���_��Ą�$l��cb��fՠ�HFMV�@0����M���١��&b���� �Z�-Ɩ �ȓ�)�H�-q<q���ɔ��?Y��0|Z⛫K�C�`@66Խ�hVJ�<��	AR�ƴb�L�)0�.�j\�H�ȓ�&maሓz���g��̇ȓ`�`�B��z����$^ �ć�D	:\ui�O�$��I" ֬��l�p��&H 7�"$��d]�z^��ȓ[�&���9mT�Q�j�0 *e���D�r�W�-�J];��24=�h���JH#���.XG:-+���Ht<�ȓg��ly�F7(���!�ARօ��=v��ב"P�$ �/Ԡ]�F̈́�RF��@������ �Y3NEv�d9��3�U)d�H�KԩJ')�����*+D� ��$����I��SԠ��0�'D�Pj0��_���k&oRz9�؈`	 D�ԃ� �j��ӵ��;��t�C�	 �����*ε��/$z��C�)� l��gՠN�fYH���R�UP^���	v��Vn_!{T��G�]�h�Z�$;D������)�B��`��Ӥf<D�(�`H�	$4�1d!� /��,�B�9D�@��MǲVb!�r�O�u�<ZP#$D���DÃ&o��,�6�?+��܃5h!D���q��,&���QTa�0/�,i�� D�lh��ˣX�!�ɟ�,����1k�<q��$-4I:��/�!�b��S�	>`�0`��B<�'�� ���	 �6(���{���F�<��̝g,�ъ���x�@�k�.\�<�L�3`�l4�p"�3[n`[�IZW�<�gδ1����B_LR���,H�<��F�k|J��f)L�p��EC�<��;�}�U��L���kv/[gx���'et%��f�$�L��"Fԋpb�)[�'r8`�(՗�x-�2�К��� �'X�)SD�2�Z�*� h,Y�'hD�ń�	p4�(�U���d�'nf�x��<���!w��~ٶ��'Z�p[�h�3N��uZ�͗*y��)�'2�8���0I"��
�/C�Z!�
�'�H����# ��IHj�	*�ܹ	�'s���pcY�gV�8b�It��I�
�'����nY1GT"3	�%�0̙�'<n��B܇ϸђeM?~�q�'��x��"'.�����ԃ;^���'����S��F�� Y� i���
�'�
̸$%�NB��C���d�,�
�'��VB�2x�[�h@�h����	�'�p�tąD_(�)C	�6wX0�'V�d��BN�rM�AbT�G6�;��O�x��&@22�dT�T�:It��"O�Y�Fو�~mK�B�LNP��"O��$Ȱd�V�S��N�8��"O��'ڥP|.�ZGI�|68@�"O<�˦`_8'�!3�'0l.�E��Op�XĝcC� �$/A�j�0�ˀ�<D�H�fn�:O,#1ɀ�c^:�z��<D��7�&�9C&b@�Q�$	�ǌ<D�ܣcˏ%{=<]�!K�%��Ѧ;D�0���2X� �b�<3�AE=D�3(I6^��	���(^��� =D���$!]�k��qC,��k�|L��9D���5�p|�s�öd1F�9�),D�h��͙)g/��Ȧ���Dr�@�58D�T���c9hI�K��1��i���8D�`�w��/Iz`*S�P�&�~��F:D�h;1�@���
v�M%CT��#�<D���c* q|�xRF�E��� F�O���O���<�O�"���Q慵z/���I�'x:��!D�А�	<<p$�O�4��p�!D��B�Hm��% t�#��#�B>D�dl	���q��-_!?Ej\ئ�:D��낭ޞQ�`��D[����B�=D��r.R�8
�xa��.n�H���/D�Xi%)N��!S�P>d_�y���O���O`�O�3�	$r$�sD��
xN9qr�� ��B�?u�f��G&��/�*a!i����B�ɄMے�b%$8��Y�1L�C�	;G���Թ2�|)Q�!ǖC�IJ��X��Ķb�Ј8&� "6�B�	�D�P�:Nf�ɦ��
�$B��8T'�(�ELw7x�: ��8!$ʓ�?�����S�π �2�NA$tP�h>}B�|�)�b�f����J��l)ˆ ��wy0C�.5�T˂�
/4L2Q�T&	"F"�B�	i|���֟j��p W"M�=C�ɰi���di2fH��3Eŏ/8K0C�I�uH��C�E�c��)E+ C�	%3V���k�]u\"�)�, C�I�
Vq{��O�`�B|0d�3���O �=�}�	Fk�e����R�{ch	N�<���ޟ=�@����Z�>��aj^�<��!��Hp W~�v=���X�<�IǠU���V�Բ3X�:���I�<��-f^���3��D������D�<���z���ѵc�O��Q���e�<!�B�{�tY`�@�cB��!6G�c�<��'E#K�z$�vdԭQɶ�*r�^T�<�r��j'`�v�S�@��bAƜX��n���OAd�� o�B��S�n��\b�
�'�����A�2%���P��4i�N�z	�'�Z�Ru�lf!���)A��Y
�'V�Q�&#á/�01@�@��8�Vq��',XL�C����	V�в7� M>����I0wL�� U�N�
�Ą�å]&+�!�Ӄ M�\@ �ʵ]�b���	X�	�!��A��$/) ���[�!�F�:_t1
$�KO�AzGV�!�D�h@�(a%ċF7b���eW|�!�Ɠr��P���܆u�4��ھX�!��x���D��N��D�h ���	P��(����3��%Pta)V���|Vy0B"OTd���p(��jӈÈq���{�"O E�_4.Y*}���S�S֛~�<ٓ�;n��1�Z�+�&�b�<Id�+m�Ti`�+%���%*�T�<q4�W�������5�2}���	V�<f'�Zqx@ PB�SD�d����N�<y�l�.a?h����$���J�<�q-ԣ�<�b�I�tH
my��J�<�ѫS Ijlq���\��pk�F�<a6f�?Kh:��r��>^0Xa ��l�<���_�
�t�P�W&$!!3��<��B Y��<���<5^�\"'@���lG{��ԑ�x��O�KlB�ku!ۿ|�LE�3�8D���Fc�V��`�K��O{&��sO:D�YF#7ypD��@��&h��+Շ$D�X���Q/FE��F�/1�$�v�#D�� ��^�ϐ����	k���ie	#D�(S���-A�=�j��fJ���B,D�(�kF�E�t�pf8M���0F�O��D<�i>�DxBe_�dޘxP���R%�(�AQ6�y���<�=J#n�P�|�R&�)�y"	L�()V�����Q�"�_��yR��>�l�f�A�w�8!ׁ.�y"G��x���h�-L�zO�[d,�y��\�)��(x'#pg�}��L��yrb��hq6P�c�g��͚�	��$9�S����lp��W� ��yCB�e@p�0��$D����b͋h˾�	����g2Ae�$D�`��H� @��h�I�T���hև$D�Q3�>I�$�R��<'>��'�#D��0dH��Cj�5�r������7B6D�HV.��hĴ�"%f�e�<���&D�h"�ԣ#�e��ҕR�Q+�-�O�=ͧ�O�m����H�r)[��H�6��1a"O� �R�%D�*�Dɱ�D0�>up���Ɵ�D�d)�*V,@9�R��D�� B�Ý�y�`\XK����5l����&V(�yB
�$�5id�������D��y�g�1����'`5�@�4	��y��"=��*"$��[�^5��ӆ�y�IN�V5���'`�(n���i���y��U]6�����"Vn(�镏��O
���O�b>�b�ψe��td�@:�Hi	O)D��P�ԵWp�e�J_�`�8�!��3D� �����.�2�Պ[�E���rm,D�P�r#�=>`��Q�m�Eܸ��J,D�b��YJF���ϗ X�r��&6<OZ#<y�Rf�H�⯒(l�p�F Dj�<�"�īWN�!"�H� TP��X��f�<�m�:zN$,�E�YO>\uKr��c�<	�È�=T8���ƗiZ:���a�<	�	��D���7�ߏG������G�<�-������v��a����F~�<i�Cߟ(���F�%w�!#�@�G�'�1OV����#�z܊�(�`	�pJ"O��%�=bl�� ��t!�̃�"O�)A�O�
k+P	y4/�".�,1�"O��: $���H,R�CD:�|���"O�9�Db��c匄9�(��'�DP�G"Ot)ffE>G� �ӤgN�0J a�"O&D��)bV࠘�Ɩ	6AS�"O�q� .�4�EB^�1�2"O@����0-���
0��K�<�"O���b4^J�<3uH\�+6�l2Q"O �АB��Od9+��4��"OV%x��Ҩ:�,�&g�
l� I�"O����kJ�8��f.T���P"O�,�7�B�#��a�!�� |BV$q �'*��R�nF�f���a@�:�d��&D��HbLM�A�\$)$��S͎ [vf/D���'��/(�p���Od����.D�@�q�ŬUA�i���L	�v� �.D�T��G�&��:�eJ�4��{�+*D�HCQĄm��Q茴:��ܒ�*O"H��,ąV�0H�Q�2�X"O�%� �����fI���"O ẗ�OײhC�e�l�DX�1"Od��A�L�X8��s�S���k "O�8s�G�SՄqa�cL�XE�"OhI�4� B�0��B$T�6�!�"O
	��NH�N�y{��C#:�<\+�"Od$���tEV��/"�R%p�"O B�_J�x!��I��:"O��
3	ډ7&@����-�ni2`"OT�GlV;\��)���@�:=�R"O�,�� �l�Q��p�Pc"OD����U�j.V���k�?r4��"O�4����  Ѱv��f�W"Oz�ό8�T\�D�+GL�z6"O:(�rثm� �x�&�r7vh
�"ON-�QAϖ*9�p��%��KQ
��"O$)2�Z�-W���*�<s18��"O��"P��'b��1�''�N!>���"Oz�b�½F'�Y�#G�;9���$"O�T�����?;,�Xg&�)_6��u"OvPx�&�,�6�A�� -,wB�"O�����ւ
�T eP:5WzQɣ"Ot媃I
V�x�	�*���"O� ���dm�x��@3cU�~zFm�"O�( ���?
����"a]�Kv�ç"O�m�L#
��` j=Ҍ��"O��8̊2��#�/0=��"OIpg��آX0T(_�S*p�+�"OP�{!���"z�E��>"��V"Ol�+��ɎWD8�.>k�E�B"OB9h#��	t�՛��LR5���"O����nɼ*�rp�"�AZ"O.ɰ��V�k�4R�*L\(�٨�"O2PY �U�C��D���&"x��"O�z����6�cB�L�!
�"O�9��d
�Ȁ5F� &���)�"O��"VɎ�K�.�Ӥ�$����2"O�P��&S��$Hj�V����D"O	 D��M�]�T��L�
y�r"O�Xc�K��c6<c�n	!*%�B�"O�@�C
�s����Q+g����7"O������x	�aY')I ��!�"O��+M;H�4��6n����"O"�IˀK��Ie��^,R�"ON�d�4D옽�"��q�P�jF"Or�-F۞�YŦ�� ��y�"O ��^/aa�5�gе��eQD"ON�2� ��C-�pЁvsZ�P"Oz{el\�Ai�����a��)p6"O����6̨\��Z�#�d�Jq"O�P��J�=r�d�`�ꀡSy�H�"O���S��63��P�J��Py�4��"O��X��ɰm�<���Y�$rri�"O��2�,4G?�t�4�L�_���$"O USv'�W�J0��Y"�Ȅ�G"O�S�	�	 \�h���_����"O�m&NF2⪐ѥ�ߟY��[�"O��r7�I�)�.M���/;����`"Ovr��&��l)4�Z����"O�!���Os`�
�$H�r� "O��1A���X}�f�S!mHĻ%"O��tLB�'�~�S3��=T��"OxԁM�Ơ����jɪF���y�E���(�A�	.�X��gO�y��H	w*� �ۡ�Rh�v�]��yb*YR��ш]��:� ���yr��=.��s��P!�L`2Fm��y"��'#� l 1��u!ȵ	V<�y���(|)�! ��n��2�G��y2[�(|�����T�~��4c��ە�y��ѝX����{�Ԡ��C#�y�ܧEF��C F� �6�j�k��y���tSҘ��KM�	1bi�,��y�$�Yh�|���Ơގ�BTD֍�y��Ȋ$p,��G�C���dA(�y���Z2z�@J�?����� �yB���
% ȱ9x���n�,�yB(�"3e*9`F�Ҳf*6r�$�
�'��j�f�g*�Z�G�N�d�;
�'4��P*ڊp�v�+��<J֑
�'9蘁fh�	V��	c���A��

�';�P��+g�*��=:�*�'�re��
��y�U�T��F�x�'��(P�ʁ)�v!�P%�o�����'$�)�#`� .����A��Vi�t�'����$�]GR�p��;�^1c�'2�S�c	�T9��@S�S�
L����� H�eP�$X��@�:��"O^�:���J$R�dZ�I�\��"O������~*�:���T�ѥ"O��#bp���ă:u⮨[�"O�e��������c� �x�"O����ʽpM`H������|t�U"O|}�oϿ*��T�AN��IR��7"O�4j:f�P��@7Ny�u"O�$��Ɔ(�HX+�$��v$°!�"O��(���+���&�G�v�Q��"O�-`u%F7;6�X�$�E19��"O��`�g[`������l��M�D"O��r��I3m���ӅC(cO��!D"O��2���+u �+��ֿ�2Ds�"O���-�&u/�p��ԏH�l
"O��A�*M�j��s��5D䠻�"Oʅ�g+'�J��)�a���v"O }�F\'B+�Ś���#$~ެ;""O6�[�)��59<lk�%.nl(J�"O�-��m%Y�2 ��zU�� R�<���c���*r�8evP�NU�<I�aȍ��B�rkb��@��,n!�Xi�����!l�hIDI�al!�$I�@���X�l�ee��y_!�d��N4:'Nt�d�ԙ U!򤚧/�-�d�F79**4�3���=!�ў!g����o����'x-!�$Nj��Dcf�:e���2bԲRp!��|S��
f#��y��1	��ш�!��?c,M�������Nҷ �!�dP� ᚄ�5�[�A�>{�K;D!�d���|����L��t�l�0!�d��tn����x(r�+wJ��u�!�ů\
�̀@�S�+���I���i�!�D��u^�	ʥ��+(��X�>�!��&12hy�8r�
������!�d�(Hv�C��9�FP���pw!�D iY.���KW4Y�d{E��hr!��J-��h�i�*u�+r�[�)�!��(^2E˥)]�	���8����!��(�$
��X#2��X�d�T�B�!�$��4���
^ $l0C�7|a!�d�����Qi�s|���"S�}C!�	@��ȳ!��F���u�ؗ�!�d�c�@�S�N�x�ZL)�h05�!�6&L8,kQ�ȝ|��U	w)��h�!�D޼l�6p:c�'t*MJ�jX�]�!��]""7�����<>b6ذ�҈d�!�$V��:��$���˕,]:H�!��˔y�mi���FYn8aUe�Qv!�$�3|�~����{W����d9@!�]�6=���כC@�H�d�2!���0��AL�m��Q��͞�!��[)+��0P�d�2�9�6O'�!�$\�r\�wc�)2u���`_,�!�D��eL�D�b�\�'q���ñ+�!�$ .6z�֨]�s�b�(R�3M�!��@��qǄ?-��F��7k!򤟚}�@tj!EOr�pe�	V!�d�l,��%쐁u(�K'W�N!�D�1i�^�'�9p��Yh�.d!���<�~%�� Z�F�I� Gɕ7Y!�ĕ�N�&����^�]���k=i�!�Ā+�p4y�b�;S����[,6!�� P�Y'mT�(i�A4�z�J�"O0�A���	N*��R��U��x�R"O~(M[*�<1���q�(-R�"On���t!���cf	`�4i��"O`$	'HT#����֡w���r"O
dzA�J�^�,x1��i��"O0ȓ完>"�JP�*��Es"OB���I#V^�(i��sG�� �"O��St$�P�F����2a,f+1"O���b�N�V��(xq�ϊf%~4�F"O�	��L"&NJ(�O4��{6"OX8��FK�6��9���+�P8�"O|i��ª.=`4�F�;�$��#"OLI{�H�����̕ �$��"O�|$�S"~5*=	�`:�Ġ��"O��Ӏ�
<�tM����(��"O���B>#.�=��#�1�:��"O�}h%�ȍ5L<"C��3
�>��"O@���N[�b�x��#B�rހ����'8�O�-h�-��iP�p�q�M�H��|:a?O����	 90f����0@+V�[�@n���Lb�	�`,��ʈ�aC���5.� .�FB�ɴ@}�,[�	^,sp
4�m� |��B�	�<�pX@����?��!k�oI�-��B�:+"�Ђ�F1&��A�afB�]w(C�ɏpV��[E�HA�0�����j*�B�	�k���A@˞�P#�۴_�0��ʓ�0?A���=��A�E_��S�b�n�<��T���r���7�H�@��f�<!�E4v�,����'��ᒄ��e?����$ɧB�h[�蓧(���� ֱB�!�D��00zehT)�!7�h��*��,��"=��9Oٚr(�l���#6h��*>	�"O��f �f@չC�ԃ�
<"O\qR�@��L�ڷ`�:q��Is���	:�~,z�Z�ؑ�k�<�!�$��L�`�e�	�1�ށ{�*��!�տR0SU��<f�F�P�K�!��Ŭt<��T"B� �Q�D�0�!���V�����k�3St�ur7J4z>!�$בO<-���2Y����Ѫ�2
,���Os������/ 14&�2��C�"�p��āʡ�yrlH�Z�0H�Q
�H����`���-�Oɒ�e�(<=�p���$
0�t"O�d'�v`�8�f��$��ʗ"O`,Q�M� ŀŢ�11� �5O@� ��Ʌhry+�N�xR�ݐ&(5D>LB�	�?(���c�~�9�([��C�ɐtlI�Q@�$4�������"EsB��.XT<U2�'��9�j�P���eb(B䉆#͠�ݜ��˅��}F�܇�I*!�h�S	�L�x�
����C��+ �$�@����>�1!�e�7հC䉔��	��
<iv�P:g	���2B�I�<.��d���z�+�]��➜F{J~*��S53N��3���HP��+NT�<��JШ\:�L� G��>�pI�1B�L�'_ay"O�$���P�U�P�N��M��ԟ0"<��fX�=px��䆥f�6��-�G�<fj�xjZ�csڜS�|����E}�]�4G{J|�r6��z��s=�h�r@Zz�'�?iW
	�hԔk1.M9cZ�	�:��W����.K�*y!�f@�S-87��<\��hOQ>]�F�ݹ ���*۝A��X��3D�� ���0�ӵ��h*��vc�]��"OA���\�.��� ��F���"O�@����5\?J,�2�]�&E �b"O���B㍏=N,y� �.Y�XXS�'kqO�0�˖�v
+7��Tb�	ޟ�E�ī�*���	paQ	��y �����y�u�䒐�ε8��Dk?�y2�{�-����o�%Y��M���$�)�>��M��[��̹f�L�U�6I�$oGUx���'
�%8��Z�"�|󗨃+Yy~Y��'D���d��, ��H��1W�@I�	�'��(�%�v#>�Sqf�<@�y���hO���U��bH4�cϏ0hV�{�"O�[�"|�rd�� TK�B�"O`��-N�~�E0�y1!w"O�(�Uh�;-i�D�aW�wwt��'��e��a��@�:�)12m�=������?�w&�)�N��T|0��YT��P8��Ez"��Xy�{ѯ�8*��c�!&�0<q���U�dG���fcH!u*�a ��E�>z��hO���f�6;��*���i`"O��+u�[�T̮��m�.M�� "O
d(�����Q�U�P42��S"O��J7$��J�$�9H�w~���"Or�S�aʌ
;��	F���7����"Oh\��Ç/5240��!�17��×"ODx��эM}J��AI�έ�"O~��uM�\����4��MXq"OP����8 �&�8��� '�8�"O��q2�Q� (���ֵX$\�A1�;\O$�(pa^�f&���G��*'������v�<	��������:�����v�<yt�	(bsL!p&�'{�V�[��o�dF{�N#	��Pգ�9B?�8���Y ��'Zў��<+h�^�����u&�	�5"O�M�QM]�n��)I�L7^#^@�v"O����'	�x�"6�ߥ;�d�K�y~��'R�ギۣ.��$�i�\հ�'��}p@��44ޅu�T%	m�<�'�^I���1�5�kW�S��y
�'��mc!�ˮ$JX�`k�
?y�{	�'��A�#�PdE�)�U������'�^qScB-$�.����ƴ:��H<����!���J�
j����fi��u��^O�H�� Y��H��D�nnB�ɉ6��iG'r�0A�f撕&��܄ȓG����M/��]���Զ~���ȓ6�,�pqE��0���6G����'��Ey��	Ρ!*���խM�L�2�k�<�O�%C/�s_��*�KKuBʝ��dk�0�=9�5�d�-p��Q�ŚnL���ÇH��d?�O �3 ��&���OB4kV�1��O�����7 �!��W��dE��C��O�!�$:M��-#���pӖ�a&�(�!��ߖA�B��w�ɢ<������f�a{����5V8Qx�F�f����Sx�!�d�Xk AX��� ��HK��I��O�=%>��4nǡoÜ�S g�9_���p��)D�<����Q��`�B��B��%D��3!,O�~�d�kM/b�-�gB$D��+�ѹCd4���P�a�t,��'}b�)��"u�|�[ �J�[��Ī�5}9)�����O�I��Z�����L=b��\��"O  ʷ m�$���`��E�>=j�"O� �Г�T�Y���[�J6z� �"O:$�u�/[Ƣ��+[�J�"O���`��.o�6���k�I��qR�"Ol�8��~��y�!��4���ʔ"O E�w��eL� �g�r2�"O�CbBN�M\R O�6if�=y�"O��&ÞH �@�2BrB� w"Oּ�SbԮK��P$%	�WZ���'��$��PAH�jԮ�i�d0�����	p}���S�JH~��G�\�p(j��P/G�n��"?Q��	�L��-�d�;k,2I�f�{X!�D)h=x!�.Z��|��]�!��q��(�4��g+�
K���R�3u>iD"O��@�K�=s�ۀ%�����d7�O03�K�)�����ΥxK6\��'�L�����`��`�BI� a��1�/1D�XA`(�06�4�agF8?�TI��3D�� b-�����3t'E.`��	P�&1D���hЪ�i �$|����$�,D���r��X�b�Ӄ��Y@� D��{elBTp���.u����3|O�c�d�A�H;�(Q��?b��*�l,D�x:r��s�:�Ɂꓝ\�t�#�=D���N�V������S�!�8��:D�|�s.C�	Ϧ���O����
%h$D�|�Uj����O��$�O#D���P�E��,bEm��X���(&�<D��93N�,]�g��d|b"�:D�<I&�J�WX4��%~D�s��8D�t����#�`"�O�n��Ak�,#D��C�K�c����bd߈\��%���4D�\0��%u��=b%�G,��c��2D�ċ"�ɻ\�X�uG�;,|�2f;D� 0Ag6��q�d焠(C$�"O:D��'��Z�e=V���Տ4D���4�K���)Sn�=��i�N1D�l�%O�?jV�O\���Q
f%1D��y�=�z����� ��g2D��#��LO��sw�W1	^(�a �0D�XIed��m:��R�{��Ab2D����'X�
���a�;v�d�(�.D��1�e�>l��2͵r�����,D�����li�����"2��,.tbC�	*�M��M��V:Bi � ��>C��c2ʵh�.�*LXޭ�tM�N�C�I�9�"����M���)�7�ܬ��B�I5J�K���6$��ڢN�u#�B�	n��}3&�P-Fe�PX`�؝��C�	1S�}u�_<q�}B$K.3��C䉃a�����g
)�e��ܜw{B�	c�Z�bTИ8�j0�#�)��C�	(hՊTA�&ۛ4��U7:��C�I�N�^%�2+�G��P+r/� hB�I5+��q�sMH,9�u�IӁI�BB�	�]�AK�*פ{R�CE�L����:&�Z�F
�nn�B��ƿq7�8���@5m2ȈrěJ�!�dԖh>,����,+/n�� iAc�!�bK6Mf�4]�A�P�!�$[&7���¤W9k��%�c�GQ|!�$W�+�X<�g�R�*g���W>Z�'����/9�i��䌆_�Fh+�'�NdP��҉q��-�a���U�z��	�'WT�Q�xlܠ�Т�}6�E��'��xfh�!��`�E�ԘC(u@��� ��
f9�
����͝Q�%Y�"OV�eoɯ
��u�Q��}Ӽ���"OV}A�B�I���K�oO����"O���A�]�|K
U��(U j��=�5"O�)@��v���G��x�"Oz��pbY���Tŀ$pi`"O� ��^,S� [ ��![st���"O�<���sy�X@p�
3p���W"OҼ3b�|����,L
�,��"O�]�^�0�h�C_�e#^��G� �y�H(���#��U$ĄK d���yR��<�� g�	7�j�d�ҩ�yR�AN�"X��L<y�|B�M���y�LC~	�m�V�I�"���`$���y�����	���58,X ����y��-��iج
�4��4hY7�yB*՗}Y��A�3R�𓭔�y��EP�P)i$�M�5�h)�b����y��V�4m��d��9z{����K$�y�I��
�(��-b���yc�5�y�&V�	�p��1j� Y�́�7�yr�ƤR֖!ۧ��?S]�xd"J�y��KF|(��G�_;E��OO�yR/�,��#��I�B���x��ˋ�y�gW+�h���YF���A�ʤ�y"��*m�V1ʧ�*�������yb)M�z��V
Kx�zw,	��y2$��e�d���`��E������9�y"b4j��4�蕶KR�TQꂢ�y�f�!U����ŧۡi*0x�hA�y!¿V� abY�{f�( $��y�C�:�� B ��{�t���	��y��X<�v�2+�%Z���Ar�-�yBG�6iX0ȶ���[e��&A��y" �*�����CRTjZfɇ��y�+w�$2�+�K�����y�		�x�Ȝ��CƚA� ]��^:�yRrW�0����=G�@���Z��y"�Wa��92��A�?Ǣ��R��y"
�2<�*T�2��5˲��y�
�6n��r�֯_�h�yr-�y��
^���/R��C��Q��y��Ԫv*�D '�E9v�����y2#�9Pv��dR�O�$���*��y�k�(�q�V w�MЁ ��y�V�aQv��a(�/=�`+mȢ�yҫn0��〆X>8�8�-
��y��G6HT�3��TIV�ҠBJ#�y��ȵ�q�e&ז+2p�V�y��Z�=F�����;�� � a��y��#>��PCAk�]q��z�GD��y�K^�vxbD��ń�#*���N,�ybď�a��)�e�9nP��2'��y�DF�~��r+��d��8�j@��yr�E�D
���ń�"���!I)�y2��*X�<��k�_w�@����y"�ն{tpB�P���Y�,Q��yFG��J\KC��!@[.���Kޢ�y�nW7v�0�+�N�!G����F���yb�����"���~��"���y�bC5ݞ�+2�^&N04��ڄ�y���!U����W$��N��̩!��)�y�D�22xp�5�Y6qk���n��yB���1��N�i��ޒ�p=����s�)��h�� ���%I"�Nz���<4�0�I"O���#L�؈�Q�+���
������*��c<��}���	����Ξ�yW�@a�F�<9�(�z)иKd+	��~ �
 �����ͺE��� =.^�?�'[����.o�ђ�e�Ƣe��'W�a�eΖH<؈1&�W�*�����bV�D�d�g�p݄�I�!�,�H��(��Bv��m��󄁩��"�m�k�aB蒠Ts�a�a
�4�JaQ��47��B�	%,���0`�k�~8��#%��Oz  pG� #�l��K�2e��uC�/c ^T8�C=ٰ��$�j�<Iwf���Hh�����5�*]�5��rk�(��E�j>�\HC�R5Z~���O�h�gFӓb�L��Z;n��O��HVgn� ���,e���E��9:������p��ܯ^�|��Č �عqt-�o4`(�����1�牵!�͸���'I��R��D.�έ�'[q[�0�)�	ɂyؗO0x���ݾ$��4��J�Ș%�$O�ܸu�C&���B+�C�X���d�T,��<�W˟U�44��1��q��YX�8P�g��E�h �H�U�!�EEM�7z2�F���7��4����<n���8����|m!�X�I�|7m��q�-p�\sU�I�?<�	r�P.rgay���,s�<�����X�HP9��>��и/���Ԛ-S-BP(�$ڦL��.��yLC�I|$<�����<��K���K�D���CZ�'�Dd`��	'Dx�Z(A��T"Hˤp���:�3��'��U٢��i��5oE�v�rsl(����]��	�z��s��p�h<���x���'LU�2�O��qY+����O�ƽS5�P+��Ȑ�"�9ˊI��O$ձqI�q ���D�8��$M��f��sR�;ʌ�(Ac܋��OJF�0���6ݑ5OH�7	T��"�(70@ߧ7�B��+4a���V[b�:�>p� j�&�*m���!���K��'o����KZa�<ҧ�T�>�f��qK�	��xh�N	���<�V�/�7�Q;$#L��t��6��$ X(#z)��� !r�He�K��C��RRG�#��)�'<�8ȳլ�U2��d%]�l$}�K>�T���m&y��=Y�RhHCL�˘O�"�j7�[��BD%��0��êO���G��-]���'�IzdE�j��1&��(@a��P$FRN|��۝Ae4����O�vXYpJy�0!����ʺ���$�?��"i#=n!�$I�����$�;x�y��V����9H����oQ6.�s5AȚ�����zy".UƼ۰�Ԩ-�j�S���K�(�ʤ�B��t�
R�Omp�0�)rvjV�5qĔ��+��G��d�0#`�``�(
��ɝ_��Q��I�**� �b۪fI��j�`P�K-B�25	�	y]F(�f�4V˘Ћ����̈�tIG ��p��4��J�'�~�ȸUʴ����<�E	ѝ;�`��B�q���߷]���!C_�3�<`�ߐ?�u�}��/��ɚԨN+X� %c-��V�����/`JpC䉂ztb0�͙�rat�P�t�J9�GGցA݌Ma@�F@�A'˔�p=(��8}���#�P�.�Z�*�[ :#
���GͶ%a{RD�tR���v��">Q!k�BM�����Z�����02,Ԍ�P�ڜb"�'e\�)�A6��Ol�2M^��49��⌅z�=����@gʼ�a�I�~'ZP�dB�1�O�r�""O��s�`	��f�B�
�[�OV��W�P�5yj��d�.`� ��E�����'ҔG�����&�9�F�8��|z*Ay��Ϥ(�DE�ݴ/�%��F�>(�Ha�@ jTDĆȓ?t°A`��+oi�P*��_3d�s'�cV��6��D�y�&к���(F��(�P>0w$�
5dʍ�a{�N�P��l�`ղT�p-�׊��6d��0I�p��V�� ������'U�D�e$�m�(uK�?	Ŧ��,O����O ���2|1�Z*BFтM|ʥ,Ρ
�~Q�mG�l`$��-fX�@�G���N���D�B+_2F�~�p���)r �@���D�>��#�떎t��:'B��h��d�9o �L�Sd!o�`�rW�ˀ(���Hɔ��E�>��f�ԁm<����G�x~�ӧ)̟�Ao�r�� �<���D�mX�D4�`T�[��"cי�M��I�"���M &��/1B��!!��=v���a��&d��3��:,/�Jt����
���4mD��L����[�A�8O��p��Y��![4!��O�nih3�K	w��|�!�/3tU��Zh��v��O�B�Dϑ]S68`V�[�aゔY�'L��C�g'��O?5�'&\l*��� �z�fl�G�'z�Ѣ�3� ��i��J>�(4�t�̹M���rq�>a6�s�b��d�- S�-`��� ,�*%�!�d�%=DZ��R�]�T�Ib�H�>�!�#LǼ�(ǆ��;�t�&H3i@!�$��}�8�b'K�P]���Gj!�$�80��(��ܙ]��%��c�*1T�'��5����i��@1��D�z�d��"�4I!��_�p<���Ֆk
M�'���U7���1�+����c��u��mL/&�\܋g�C	[���ēfڬ �6�C�}4�M�NG�/J��v�˲l�8��d� FEfᄢv�x]�#Cېayb,�B��&�,�2�`�n8�G�
&�!dI?D��鳠Ȫ_�1"&�W�4 ��k1�$��Q&|r�{��D��5q�dIvLX_ሑ��J]���O�Tc!g*�'#�r%Ò�8$̍�Lݰo�� �{��6G�zb?Oj�"e�>8z��2�@�M͚��7O$���G.���h�� �����U�P��U�E�&��D2�˲hLC�ɿd�0t9��ۈf�
���T�q�t�ʢ9�M$\OT��u� 3-,���NB
+y^`!�'+�<r��+"pl�Q���]�M��Ҷ,#^���'����-%�V���?-�4	�����0{߀Ġ��)�p���T �7}}�Y�Ú!D!�D�'�̽x��И.2v��eT�DI�
T� ���{���P"|���Ӈ ׁ�xB�C��@l!�䐳d�N�H�&.�|�P�1)P�M_.H�
�xd�ia"��J��ؕi�3��U��8���r��N�Y>����&��xɄȓSˀ����U�%V~8Z��Q����ȓb�A� ٱ�4�$oM�"F1�ȓ#�tʦ�U���z����yr��7L6J��1��M���	G���yB�Ü%����窞(Ct ᵢ��y�'�2�����I[�9�,�kE
כ�y�k3G�ܰ#��2�*�%���yb��h��Q)ɡH�eQ�4�y"�ئA:&�Z��� (��|���G��y�λ_GH�H�*ɖ&2��b�^��y���y�2�B&H�#fE4�eӱ�y�i֣D��� �b;������y2���х���7b��z����yj���ȓW������7Sl����H%�&M�ȓ%>��Ȱ�#H�\P3� 1�!�ȓX�V$�doɭ�8sWE��b$����(�Q�/��:��>~�H�ȓ_�*���c��]�L�bGU9Oj���7>��'���`h�lZ�LKz!,���/��4&Րj}�D���� �����x�A��.]@>�B��\�
�ȓ_;����x�E�a���6����/jB䐴MʂA)*1§hǤ_�Tt��K��أ�jP�V�"QX5��.xԨ��z0P2�ՓW��Ux��[�� ȅ�l�p\��JS�C&N �Q �܅ȓM�I����/��'��V�b��S�\� �(�
=A�xBR͚���x��h�x�A�dٙeX4��C1}���S]�f`���A#u&�(tֺ�ȓY�x��jU=*׺��Fb�(To�h�ȓ���1��Z�R�k#�M�`�,Ň��*�9��4`���"����P'����c44�P#�_��@z�*/}S�!�ȓ!�P4sd�Ȓ��%�É3AzU��E8�(��	!t�@T#d�z���ȓHEj��'J^�#�B��UE�?�ń�S�? vE@!n�^��-���+��lS�"O�P���C0P�)xeL�M���"O��ѧJ�#D����²+9�\#"O���v�"2t�P�b�2,>qh�"O��B�o�UX�Xg���WN��"O�k��M�`deXS��:��Е"O��,E/X�����gX���{�"O
���!{֩b3�"yƅ��"O���k�<;8j�0�c�I�ك�"OX��&)�:���q◆\�Ɂ"O84	��9��ܩ��\}�U�7"O&��cJE�W��)E�6IT�1Q'"O���Ơ��<<��J�4 O�"O�lA���~3l� �KV�1,�|�"O���z���!	C,#���
D"O���;0�X"����є"O8�0��8$�} ��^	'��	�b"O�PA�K--�4I9���/�84I"O&,Bwo�r	<@xb�/`�4*O\�C�ٷX�4�J��� {�ޕ��'z"! ��#����P�T`'ر��'��#�j�y=�ب4��0XF΀��'�bB��:����#�T+��]*�'V�L�5��!A���j�#n�9��'>Z���I1C�,�[!�j��<r�'�p����+|�*<���>P�|��'֌ ���)X���%D&D@T��'�9�V� 3��s 'V#'��
�']pq�@j�����2Z6-��'�:��v���b�@-�fk��)T��B�'�0��d�4��y��͍;Qƪ���'��m��)@w%x�`^'N�	�'�n बؾ?,q�����݀I	�'��방"�&ɲG����z	�'r�D�'A�;�L��@����	�'�=��c_"D>2,��/�\���'����,��u10�)􏃕_���'�n�
��W5MV�e�C�C�T��L(	�'� [WŞ�UMH@�S)\*v�S
�'Ln�v#. ���&�.r��z
�'슱[�MT�G�5��n���bi��'kB4b`�#$�\ �PJ�P�'4 ���VT��m1Vm ���'R��g*LZeTE�����A��'�",�Q"��X�[*K�V�D��'L�,h��ɮZX������
O�!�'�D!�l��� ?�A��'��a+�� IaL�ZM�6��' FlcD��!��1Q��D�9����'Xx�Qġ�*����@@��3Q
��'[2���ًRb�|؇�U�{1ZU��'����&�2S.
=�F�ο	����'Kx	�W�!W(���"C	���
�'游�u��-R[NP�U&�U�Z�	�'�)0ugY,�ܡ`�52FZY�	�'=�1PġD}�d�V#��.�E	�'倭1Q�1-��T[���Vx$��'_���S�$Ԇ���� xj�5:�'�sq��d`Ip�!��Ȫ�'��!��"R>Ei)0���.N����'��Hu.�"@�� '���@I�'8��`�����W�EM�C�'T�z�D�e�X�9L�&O�fm��'���+J	 ���hňMnA���� fC� M�RA� �tջ���"O*٠��{�8 Z��e� � �"O����;�����C�0}A"O*���D�#T��MQ��@��y@g�'RС00�<h�]Γ!��x�1� �f�\�@� H8NI��Ͷ���L� g�Fs�9g_v��<	S���eZ~�ـ�˸�h��H�rm"X�"C��L���"O�+�f��r`�D�t�ܰX�lep�Q�Ah�UWfd?�F�����	)FĹ��*���$����bC�	8`�ٚp&ߩ;��%P"!�3#� �"�m�m��J�'a{B(�80��q3��5�>h�u���<!�I�7�&@����1���C��
4�q�L�p�T �u���y�'^�-�����#����MH��"����'�i{t�����==񟪀@�OӌD�b!�B�4�Z���"O�����/̼@B��	8�.��A�>SR0��"
'!����O����&��ņTc0c�bT9|�tهƓ8j�8���R�(<
2o�'b#�k�ƈ�8��ayE�á%�2\vB1,O$��LD�&����h8�-f�/��<��eL
k?�5!-q�x)S&�YSI������*d;��3�i�d��C�ɛ)ϖ����W� (���	:�c�8�dS4>���R�X�-QrAQ���(G�j�X��+LRYH��D�yb"���U��;SL�S4&Z�P$�Q�a_�21�c��O����Y�|aӍ�*3lR}:�C,&M�L4K0D�(!dF��"���ju# LN�X,�<�&kՏbL	�"-,O�ؓ�K��K�Θ� �\���`%�'���PU�K<*�&%H��G�Y����_��R!BH<�2�d��5���6�6�x&�G�'�E0Ɯ-8���҇+8�d�h���|'�\@"Oʱ{a�K�vLA�غu�j��O�T:�#�����h���c0�eݘ���߁cc�؀"Oj\�i3[j�u��-O"[������R @���	������	�0z����̯�����L/��Ma�H��2�H
�#$=hU��
��ٳ	�'���0�I�;%�-���$�FIZ��$��&"�R)N��O�U�ː8G�c ��$�b�'C�J��YSP���P�ʩ9r͓eߒ=P�eʘ�ҧ���]$n8 ��Cq�A.xP���)<D���SB
�vM��n
����0�>a�-�4q_.�����EX����*#4e����ڶR�ȥI�B9�OH}��c~��2��-}��e�fg
�m5d�Ƌ�:h]C�	�޺�a���~��BD-��~~b�<����Ԯ�1G ���O{�؈���k�
�5�[,^�����'a��Q�!�_sT�T�<" �&��F:��g�R�B�S��?��
�kl��2eF'EP�lX���i�<�Q �tl�Q����A �40&�c?qso.
%:Q��qx�d�D6v�(	YP+��_��	9f'2�Ozaʇd��N�y1�Sd�5�w�]/5&� r���y��K�F�2��`�ӗw^���.ڼ�(O��+E�ʹC�>�È��R߰ՒD��8���,�C�!�$û��b׈ޫ-�aa�	�:2�+AiQ�u��ʒ�>E���8מ�B�T+T��D2��I/���ȓ$�0e�!n@G��0�P �8	�2��'&(�$����zr�F<��%���ϬC��-��M����>���
Un6M��A.��Sm�I�T)�*¶P�!��QKeĭ!�0��O�FL��'����M�o&��;���?�Y��'���� 97����0��
�'>�!4*�5F���biRd�����'x�qi6��`�$���O�Jm���'w|�[sӘJ/\�w��<��	�'�<�P�U�=�� i�36"�z	�'�ZpP$��1EP�@ՂW�~����'*<`��_
�0NC�m����'��t��`�- 2B�(1���oÐ!I��� D�31d�U�H�t�3�Zx�"O	��c
l��b�C�%��)R"OX����%��;�cPR�΄�"O�5q��L+~.`!pAEN��3W"O�dxDdأ ��h�A\�b�ĲT"O�d@�3L� xh���4����"O���F��B�ԂQM�+U9H���"OpI0ף��î`/A�P��-	�y"撟/��(f'Wbk������$�y��\.%]�%+T�]�I�Ej؃�y�],=נ���J��P
bYô!A0�y«��\,N}(S�D1B�bq�k#�y�oN�\@�f.�'NN������y�Lâ|^���f�3D��0���.�y򇝐?���(ҭ�?�t��ɂ�y�>')�4�F����K�ƙ��y"�ȒKI��xu&�I���l[��ybN��}jt��e ��B��8;wGD��y�Ӫyx��&T82`�l�y"�T qY� �)$-,��E%J�y��K�:���V�$Լ���!-�yr��?!��+�fD�
K�ؘe����y���n�݊��ăxق����3�yR#�	I9��)A��n��_/�y��<���.@�ʺ-!v���y��߄Q��� UZ���M��y���i�ȭ� ��G��5	E���y��h�|���g��8��෨��y2�V�p�ڑ�d˔� >D!����y�O�C��s�	�i`�ۖ���y����q_��R!I�!n%���h��yB�H�B�����"b��h�R��y2��3>�ȹ!�l�u锑k3�܇�y$��)z�q�"�O92"Ή�b��yB
BQ�=SE*ǔY�&hPRB ��y�F�}׊�pwf��V����&ㆴ�y��Q�4�� ���D���Z�o�3�yb�T4�y�DU�L䘀��'�	�y2,I�-�Pċ���?�lh� ��yҏ� g��P�$`������y���wT<�Ǩ[�}vɺ�eA��y� T�$[�	ԗ	7���Hߗ�y��T�Wl޴Zj@�YFZA�E�A��y� u�h ���Z�c�FD��3�y����������^��ˣ���y����Ȅ�,�� X�9C���yReE�JHb,�1��q�����K��yBJ�;N<`E�q�*zcEʓ㙶�y�Jק$Ǵ���ڂp�8 � �y�!��+_�P�hpY`F�y���R�3� ^�AI�x�7�.�yR`A,s?>@�0��6l�H�i�-��yR��F���,V�o�F蜆�y��Ɣ�i!C�(B�r��W��y�k� BRC�``���"+N��y"@�)8H�򲅘�nT�k��P*�y�cN3��=ʂ��q�D�%�T��y�$�\�����	�*>V�9%E<�yBb�v������bt�s%�C��yRGɁJ��`�߾d��(at$��y2%��D�t��A�_����8�y�1;8ԙ��oG�Vi��P.���y�EIP�.�P2l�8u�$b�\4�0=a�d�=Jp��[�(EܼjqnȒmkmjƮЀ����_�<� �,zƃ��!$�!A�Ƌu�Rܺ$"Obm!Ǌ-7�H$�ΗW�t2c"Oƙ���<�h�ul&~*�	R"Oj��a�v�t�_�:�	�S"O����Ct�$��J�!�2��#"O��0�!J�s���!�I��p"O��bg�T
܈�CU)���$�IV"O�Z��K�[��H�T(砱��"O
��[!(C���GK�W@lI��"O\P�VN� 1Fr!�)K)>,�5#2"O�@T�
�;_�Ƞ��,����"OS�U�]���W
�#�2W"O�@G���rP�Y���<�&�(��'y�ov��#�N[��|k�*�>bT@�v'Y�1�y��	 2gh>E3���2����[C�${�����	78���'>�ю��oO'fg2�� �ua ���g�|��pjfá�y&�-~|$������tM�oB�%�B �e7flZ�醓A�vM��O�,�!C��O6���S;'�a��E=l�6�J1��p[��,�e���
Q�
�ӂ�O~��H0/��ۖ�Ue8	�ڴQ�����r�Py+O�?M����`:�9��h�(N�HՉ�4z�=	��ڃ{��IO�3}�O ���m�?]�.�[V�%<�$ �ڴ��"~n����)V�Ixb�Y�bP�vtB䉤h�\���'b!h̹"FʲW�dB�I��� aˆ�m0��p	ǅ][LB䉸^g��8f �A�e��X�B�B�ɏA;��3�&�?hV��g�T��B䉸��q%�;o����7-�$u�C�ɰ
q\(Z�V1kq��B�N�K�C��R���g�NGJ@	%E��B��=s2�a��0
��"�9���d�0E\��J�uK���A�P/!�$]}Y��1щ{8�x@��֒r,!�DB�~�|���&E�,���nZ�e�!�$',��XyFȝ�1�CI�3U!��"g&�jA�֟@x�6��"�!���>x���[@�{Q�y�`C�W�!�4�"�UgE�[GV!QP�O�!�=K�����ӑ�
��p��~�!�d]=2@[�#� #��=k@�GB�!�$� |�>��/������&  s!��%
Ĺ��͂�p�z�J��C�!�C,dM���TKA23ؔ5�bCE�!�$+�����X��YDb��!�d�_�tc������%1!
e�!���~����ıB��壳���!�d�64z|jQA�bk$�YC�Ӌ9���B'Q�hP7O:2r*!r����y��܊1䶜��E[>zP�*�]�y2$�>@���wB�mO�ـ�$Ĭ�yrGX()\�Ճ��űX�D�³a��y��ӎF���yՀ*J��G�!�d��Xy��a[ ��[V�\	!�Ė�n�~!{B	�p�b�î$!�DE<L�P��ȝ!d�|D�1@.N�!�%k$�$Śx�t��;�!��W&k�^|;��P	R�ToV�g�!��˔] ��·K�X��Ō:�!��73��\����/�ީ��AU�`�!�$\)bd��0��T��#oYZK!�4 ��u*�&_�r��l�����U�!��B�7��2:� }@e��8vx!��C�ql�m*H�rc�Qc*C�w���߳Lx*=Ȑ��pF�C䉋w+6m8��D'vh̼jPd�5� C�)� �X��$�"n��4�b�1D����"OBy���N���z�aF0C32��"O4��&hҹ2�n8� ?w���5"OL�CW��n���k�H]�~e֍"O�I�&��� �v�ʜ>�\��"Ov��*��������`q S"Ox�0�7lA����1H��"O��Z��?jHa��nB�w20XK�"O20�c_�i��`Rl<>%ve�F"O@-PF�ԯ$�2�2�֤
#"�83"O8�� ��M�<�)D	M"-
�Ͳ"OR��u%A���80�G�-�ވ�"O��2eD�r�>T����-Aߌtx"OpU�n�4;E̬ڀ�X�!�܍��"O&� f1:�b�2%L	-�|�C�"Ol���,�2�*Q�����d��"O���������Re�ċq��M�s"O*�0�LY�X�(@e�`u�I�"O`�cׅ܍�}�s��q�=��"O�����V��>���B�l,D��"O��獊+{P�Ӧ�>i��*B"O(���4`�������n�Y�"OH�Sd�yL	����:���"OVb�H֪r��43���}߼x#"Oy�bM�@�p�"Z�X�v	�"O��Z� ��}J������.���2"O6T9a'��|.�jA/V'Eb�=�2"On����&sn�rX��&�*8!��i� I`6���0¦�B�%W!�$M%h1Jq�@>��`dU3Z7!�ā�d�{� '��5����P!�ҍ:�rPK#n�@"diAR�2�!��,�fQ`r��z�����ӏ]�!�$��i>0!3��������b�<]�!�d�>>�P�q�g	�a�P�YToc�!�lm@䀃 ��.W�Ԋ'A̚S�!�d]+"�H*X�:6R�JB�pd!�DXH�t0!�c#څˠ ��Rg!��p��f�v}0t�5�E�,\!����D����.\�N�{���B�!�@T(N����w�Xġ�-�<x!��_�h�X����P�3	.)M!��V��-�w�
0$=dXa���W"!��Ұ=c�� W�Ǻ%�J���",!��B&n�F]w��+�p!܃j!��ܢ:`Zq�C)�<P:�S��ԞY�!�0�nq	����HO���S R#�!�ē�R�4����Fi(�zV��2'�!�[�<e�h2�N�EOj3��!��<+ v�{8���
��Ql!�
a�ص�B"�T��5���ɞ&W!�2}:`�IqL�({���P�J�q7!�ޝ*#`L�whM,A�P��Ş}�!򤏒b����AS�d���r�!���&���R"��M)��X6B!�&+z�Z%$Cb������/!�$F/&|�}��yD�q�֥�j3!򤛞Bp��+E�z�]�^d)!�d�9ij�
Ad2l�
vI�X!�ě�TV�ݹQ��,�$\+�!�i!���I�64s��W�w�n�JC� )!�d��8E@0��~x�ٲ�+D�(�!��(-B|@�!��%��8s*V�A�!�߷[��@��p�8��L�!�� ĳ�EG� Z�����Pz��"OMr���0�,�r瀗EJ�<"Ob��RB��q�$�Y�/LP2DH"O����O��p #�oϏc��{ "O&0���ܟm]��ڶ��V�Xqʁ"O�Ӧ��~�F� �'^�v�G"O�Ԡ1-P�������q�>��"O��+e���maZ�Q呰J�Ti��"O-¡��i�}�vF��5�<��V"On�@aU�9���ӄY n��v"O�R�(�Sx� ��i�S�>Ԙ1"O��wOt���P�iqv(($"O2�j2)Y%H2q�);v� "	�'GT\�ԭ�&�Yt� /4��3�'����a'G<t�q�c���0&�Y�'��r���'��"	2Y�X��'��5��I�5�땟�(���'{r�jӆ�,b�j�) �N�|�F�
�'c2�;�/]��&ɀ�![��:��	�'��ZC	!K?�����61$U1	�'����C�7����N��~�\�	�'v�(���D8�kw	\o�H��'� H��g�^X��+ס�i�"Ȑ�'-B%	S�j62R�e̷w�~!r�'p&���M�?n��DY%%�~�
�'~|2��$E(�d���4��9�
�'����L�HV��C�D�'�����'�~���M�������('�Ɛ��'H�]�D�hrT��5*���'4�A��@rꀕ�Ԅ��>�Ԙ1
�'l6<Ұ�
v�Y{�;Z|��	�'�&;p�V��T*��.��s	�'
-���1=F�J�NG�~4MQ�'��L�#n�Y����k�^@(�'���"�C.J�Y���b����'�^T#ҩ�����놁�b�aq�'J�`�W��W9f����T5B�
�'rYE ^���G_�LE���'���C	K8_���)���Ah���'�������[�td��儙8��I�'$p��)�i�N�P!��Q`���'��3��T�V��mZeƝ0rx�h�'�*�i��̮""rŹ�ꙟ ���'�V<��W+�����b	r�'�̛b��]v>�(��S��PMh�'d, qnٺP*�'��&�6q��'8Ԉ����O
���v�X�d����'S��W�W*u�X�z����.u��'|��K���1k�H-z^nl��'{Q�ơ%!6�ȹ�쌮n��y��',J�1v����AQ�X�P�'Q����$5V��S��񈉹�'�hh�CLB1z}���S���+�'9f$b�4G$���Hx,s
�'Ø�[s��r`�����*��1��'�L��N�z^��A0,�Ԝ,��'�<z�.Q?ꉢw-M�!����'9�K�LW;c�%��A
���0�'�h)9�X/)�>	³Ëa"h��'�\�'�T"C;�D�2	�U	��	�'��H��[/ Ѱ񚵈�:R����'���2�̰:B����	¯A��y"����&�24F#���&�y2ǎ=;2Aq�6z|9���y
� �}�����Q���̵s�%a�"OV�k�F	�B�ZP!�Tx0"O���/���2	R�e4"3���"O�xy�Hޘ�d�F��`$�r&"O��
��a�W$
(�(` "OrY���Ln��)�@�[�:��m{�"Ot���J&���#���R����"O���w*�6��,����, 
��"OL��a��� ���[�
�-��"O�AaR�D@�ࠧI�[ҭZ�"O�A$%,z�՛�e��I�"O$]��o
v��3����6���T"O�(�PdՈ�4��e��o�8i�"O�k�S"	�
	5�H�"��Mx`"O�A��ɂ��e� \+][n��"O��N�0^�����nBVa��"Op��ᤏ�<T�F& �I/��2�"OPpQ櫃�O X�6�
/)b��"Ob�"� G�x�t��&��j��p�"OޔA����eV�򲥖�N(�"O,��v��;�P05� <�N��"Oh q�kO
L��T�W=o�T�"O�4q���9N�[���B"Of8��g�����âҨs��=B�"O�}PcMȾ2aP��٨Z
���"O`؂'"�5m9��� ��� ]X�"O^<���*��!��/R:<�ic"O��)D�1RT��ƠR�0r"OHD�   ��     G  �  �  �)  5  c@  �K  fV  b  ?m  zx  ��  M�  �  �  U�  �  N�  Ѹ  �  [�  ��  �  t�  ��  L�  ��  ��  b�  ��  C � � f N �% o- �6 �= RD �M U �[ :b ~h j  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>�z��&�A� C��rs��i�99�E��^� �O��oW��|��?9�h[%�`n��u&�3ȋ$G��'��񀕶i���|���O��'BU� )a��k6�JP%��0���<A���4�'uy��s�B�Z�6�w�#�`�V�i�h ��y��i����ݯVsr�s���x�PE�\�Q����I�(����	�f��7�b��a�J-��U�CԪBO�aj��i���a:�_f���$�'O6u�_/_��`˳ 5>;.��'\�B��M�"�^�JIB��%:O�A�H�V�|�����>��?�'��I�%�ܼB�a5������1"{d��?	 !@]D��|
0�O���W�B�����k,��􏊭x~p�p-O<��?E��'*l��,�[��� a��K|B��'�:7-Ai����M���Ow@!�C*��=��]c�E!?�|��'���'KR��N	�֐�ͧ���$O
*v^YH�? ����g�t�8�$�������'�2�'GB�'�0#�T�_���$x�@8�T��(�4X5�5���?9����<��I,*>p��B/[�����	%������	w�)�8� �+@�ЇB�tH""�Y;x��CC����w�<5&�OH��H>-O�p ׋�"ۚ�"F�(k�
�w��O����O����O�	�<q��i���1�'F��qC�1 uV�i�j�**�jU�@�'26�/�	����O^���OV��@�I4E�Xݙ%���  Nr�7-;?9��� 8�	0��߽����8�* .M�/W�����p���	������IƟ�����č�K�}s�$ �̌+3B�P��Ɵ|�	�M3bH�S����f�O�嘲��D�渋6FȚJ�����9�D�O$�4����rH~�.�c9�l���T����iƓ(Ȥ�I M̙X����@�	ly�O��'��Ё�2%ʶn�!x2�A����U���'�剅�M+A+_�?Y���?q)�J8�V�G>:`�2��Y.,$D撟Hi�O����Oz�O��f�|0�F'�.��<��hπA�"�aF�ǻS�2����ay�O�J�����'g,�[��)�ԍ2���b�T��'��'}2���O[�I�M[g�F�8��T��E!�p�a�λ������?���i9�O���'g�C_�e��j&���P��Xb ��6^��'���bF�ix�	*��u(��)^/wϘ���MA��A��S�;��<����?q���?����?	,���Ѧ�ğib����S�
~ x�A�]֦]i�k��p�	ßP'?�	��M�;:�91u�ZU�,B'��?�����?qM>�|�w+�,�M��'˂���.zu��l  A�.�'Ӫ�����D� �䓋�4���dͼ.�Hi*�l��i#ce�J�@�$�O����O(˓E��6G+]��'+�aTB��5I��:�$��BZM�O�\�'����\(j���I%B�c	U�0��ɓJ��i A�Q�~d�$?U�'a��I�Q����o��kҮer�7ܐL��ϟ ����P��a�O���R�g�0��.�N�����&�!�B�fӪ���I�O����䦽�?�;b���ʃBC2p��%�2ʮY��?!���?Y�N��M��Olqyqf�2��D� 3oNjH���ɶ@�xE(����'��i>E�	ϟ<�I��l���A?��S'��|_�2G�e� �'R�7�9��ʓ�?a���i��;%
]K�oרx����̏$}����?�����Ş9�P��VnѷFc���PdU�S��)�!շ�M[U\����ϕ���1�$�<��ƸP�j���e���π��?���?q��?ͧ���̦Q'�ݟ���I�)D���s�U�s.�8���h�p��4��'@�ꓐ?q(O^@�E&��BК�	��*њY�w@FB7�4?af�؁�|�	��䧔�� �5
2�V�N��R��{����?On���O����O����Ox�?!u۷_�Z��H���]��-ßx�Iȟ�ٴ!BZA�'�?���i��'��@�RbԯL��ԨO]6��y�'���+k��mZp~r���*�:d	��������E.!�Q�ן$Qџ|Y���	ݟH�I�lʕ��6!����U�G1M �{E㟌�IKy�lp�H� � �O\�$�O�˧{~\h,�6;�Xyg�9=s(��'*��?�����S��C��  0V�+Ȏ�k&��*;�(�#^Mژ�O��<�?a%&9�Z�1��T��m��}ˁ%�m����O����O���<Q��iu|T:��<�5�*����Ј�m��'�&71��+����O `����>La%��QBȱ� �O����]��7�&?a㱮 HA����ӷ6��pr!�8�NqQ��}���gy��'[��'�"�'�R>Y����L��E�Y���am�MrN�	���O>��t��Φ�c�ȱ����a��S�݂R�A�	˟\$�b>��f ���Γ2�2 ���K-����/�e�oh�Ԃ  �O��I>�(O���OJ��4���I&V0�BǃD�ʙ�%i�Ox���O��Ĺ<1��i�Z�s�'��'=:P!�Ȩ5����"�C�2����G}"�'C�|�Ǎ�m���@)��+�9��(�':8R��W�M����/�~��'À@��N:FZؑ"����=�~}
��'�B�'�r�'��>���I�(�QAσ3Pj,!��,�0����M3��?������4� (2!n٨We�4HG�K�`l��ZD8O���<�P�9n�e~�%�=6�d9��q!�I��[B��U!�'>�HY	��|R���	՟8�I����	ӟ��%��&t�.􋁅ڲ~�|1�"�Jyr�cӮ0���OZ���O^�dU'�v��e��f�r��1�3F���'���'�ɧ�O��y7@���2����	�i�D�׮�*�dJ�Z�г�^�3l�(�y�I~yR�4�f�B�H>Q��F��2�'$2�'0�O��I�M����?92����TE�k��;V�� ��<�S�iK�ON��'���'CR&Wg��a��˔^�ݪ�)V�X`��c�i$�ɧXub��E�ORq���n��>�F1�a�bZ��I�P��D�O����O���O�D3�S(�����f㌔�o�Pꢕ�	؟`�ɵ�M����S؟<H޴��*-���nA�w�.�����I"@�<������q?�6-*?��bY�E�R�hnQ m�@�J��C(���*���O�L>	,O$�D�OH�D�OBq9�c��5���zj�+�����O`��<���i���!�'���'�&.?�+�LE�a����͚e���4������{�)*RLʠ+X�HY�H��R��@u��#�"�+��<�`���D���E�|���U�}q� XX�嫑� ���'I��'���P�H�ݴY\�y�d �3�������)����L����A�I�?��[���?]
�±c]'D�f��3�x���t�F�����'�p�Y�(Q�?�@�q6�P�p�a��4���C�0O ��?���?I��?�����ɇ1=��0`��C�-�{������������ƟX��ן�$?]�I�M�;8{.pz ��:m��q���۶aT%�������O> �:v�i=�dL�m$!aƃF�|��ȢU*
�?�d}<z����X�0�O|ʓ�?���M�~4Xq��m��%�Rm(W�X R���?Q��?�/OV,n��_鐝�	���	�}fe���<o�&Yq��>�,t�?A�W�d���%��"�E�o�:h�� [o����1?��C�<��ߴ|O�O3Zi��?1%iJP?tӒ��$�d��机�?���?Q���?!��)�O�4�/֠(��
�DD�����O�n9E��8��џ�@ش���y��_�ְ"�D-vњK���yr�'K2�'I�|{s�i��i�mJD���?�����2:� `t���C �b$�� *#�'F�ȟ��	��I�����}��hۦJ�8C� l��T?��'�T7m&"���O��d<���O��)LD�t��]+���0&B��U]}��'���|��d��,G���WE�B0��'���T�qp�i���.A,�Z5�O��O\�FێQ1�J� 6��d�v���C���?���?���|:/Oȩo8��9��4��陷�͒t������/���
�M;�bg�>)��?q��,m��ؔF̷��iC�6rU����݉�M[�O�U�	��B����w���+�#�,PHfG�8�|q9�'<�'b2�'�r�'�ؽ���Ϣ-,�"1�D��.	���'�R�y��}����<Q��i��'��qJ�b�%b-����EΜu���I�y��'>�		4�n�@~�n��T&��$@�e{
�+��ʽ�6�i!���pX&�|2Q���	ݟX�	ן�+�kL:\l2=�c�ʎ4�TH��������xy��{����%f�O����O6�'h~�����S�@�2ȉ 	D� �:�'ݐ듀?����S�Te�?��HbV�Z�gU��bE 6HTF��3d�^��<�'+BT�	U�ɧ-D^U�M�"iXɉF�X�?�y��֟(�Iߟl�)�MyR�n�uj�� J�� E`�(Δ1��i:��$�O4�n�p�#��	��0��#2n�MٔnI58u�E�"K�8��*�8mZe~Zw4����O�e��� �qd&�cQ�af$�=�BH@>O��?����?���?����%:�ha��͛=f/HհWl�4X�,�n�4��i�����Ik�s��������V�%o� Paоo	&` vhJ �?Y���S��j�Sk���ɤ>�y��+JT�aKd��u���	9�ta0�'�(�&�d�'���'hMY}�l<�"́5R)(R�'���'oT��2�4Y��Aj��?���Ah2�=��5%��_^Z9�2n�>1��?9M>a��U�%R��H�l�Xj��yf��S~�,�$7`�\� �P���Ov�H�ɥm�٘]"����M&3���)0��b��'x"�' ��ݟ�Y��_�"5�$�-Z4 ��cB؟��޴
_����?��i#�O�.@�z�P��]P`lBD�K�rp��O���Od1y��s����xс*��.@�Ü�B�TF�7 Y�qaE`E�䓠�4����O��$�OR�d�~�p���ʤ:ͬ�j�$�8|�|�6���*Ѵ'���'���)�4/[�
� �٣k��)Q�X���u}�'�R�|��t��3�u��ȑ���e�POC$6R�cQcѥ���=�� Q0�'�4&��'�h�A�M�Z�E�Y0G|à�'s��'{���tU�	�4Ve���#p��Z4c^-X5Z�d���@0�n6����L}��'��I)n�9�֯��DL���� 7���I�˦��'�|�J��?�����wo�i�&��W�J��"�~Μ<��'`2�'�b�'8��'�� d�%Sp��h
�� ��%�2@�O>���O��l�--3@�'>7M/��G���yP�D7r�a��.U�B�t�OJ�$�O�Q�'_7�-?��!O�V�b�8A����ce��Z����Պ�O��O>�-O�i�O����O�Q@J�	�lU;%V� ����O��D�<��i���)6�'���'���p8�����6U ��F Wנ�C��	��P�?�O��y(�C�@�h(��B0d@��o�bՂ�p"�,��i>y&�'� &��� J�dp��`��	�}��<�	ߟ��	�$�)�Say�k��5�SkE3�Dd���*>�j}��%��G�^ʓg��v�d�j}�'��Y+hB�z&l����i��%���'���t��v���݃z"p���i��	(<�����bWH�%�t#Ţ|b�Hy��'�B�'��'v�Y>I��.L��Rਖ਼.�����:�M�F���?9���?�N~*�y�w(�=�T��l��Q���~-�Uڀ�'UB�|����F�o���6O(�K�
E!H��`���"O ��W2O`��bV)�?y�$9��<A���?	d	N�_�N�PcK��'�V<ᤍ��?����?Q������Mj��ß��	��'�&B�l��6��	ҌLaÊk��G'�������S��#����� :�(tYt� 5^�|�tzQ�ӎ�MSr���f?q�h���G�RH���g.رEt֝q���?q��?����h���E�~Z��+U-�6��u��{PF��˦A�`Ɵ�	�M���w$<ࢥ��*����زU���':b�'�2%
�"�����`3VnU*4�)�$�2��^�<1Ð+M�8g8u���|�[��Ꞔ�����	��`S���2�JLIP��?Ί��Э	ay��dӀ��E�O �d�O����_��MA�Kϣ~ l!��dC.BQ�'�b����GuP�(X8�c��	�F��t���˓'�1Bh�O|�N>)*O~�92�Z)=h����V�:���!�O����O ���O�)�<QE�iv�l��'iƥ�̇,<�B� e^��*�'�v6'�I3����O|�d�O|X�v��"9�� 8� �?�8�৥U8z�>62?�P����H�S�ߵ��Ƙj��'MA:�����k���I˟�������Iҟ`�
�M��yNA��/�	;ON�hW-�;�?���?92�i}�iq�O;��Ә�O�9����0k���Y)rN�bE#>���ON�4��4;rGmӴ�yΦ�+�	 x�퓧�K�/Ō�4��;���n�I\y��'eR�'KҍR,k�-�򅍝Ӯ�3��Z^�P�hB�4j������?�����I[#��m��) g"i��
��l�I����Ot��AFH�,��b#�� k�|� �� #~4�b]
6�R,���4̟˟K!�|�K�W����JV�dH�ly��J����'��'A���Q�l��45W�9����.bC(��)�b�},�\=�.O&`nZp��'���ʟ�*�;]�N1���O=���FG�ǟ����R?�xm�g~�N�S��|�}���t8`��3�)
Ȕ�It��3f��Ķ<Y���?Y���?��?�.�L1�!���`�h��[�}P*D�Ȧ�R�̟|��矄&?y�I2�M�;C�<��H.mJ>$���Ќe��X1������O:2�q�i"�F����'
�	48%�@g�D]�e���X��t��O�˓�?i���a����(8@�7mN`X��"��?���?�,Od�lZv�"%��埠�ɯ<6R�I40�ȅ@
������?q�R�4�	쟤$���J
z�0� �Y�=���")?i$�3���Cw�DO̧����E��?1�^	�%�v��7�������?����?����?ٌ�9�����\.~������B�̀���O�Unژ^��ѕ':7�;�i�)j��ޓ[��xp�hed�0�{���IayiĠe$�6��\�6E2���>� &���ڮ5"�T "�+~��B0B+�d�<���?����?����?i��;�Ҹ���^�ƍ!�f���$E�M�pIП0�	ߟH$?9�	�X�X��Dcۑr-45�D����O��1�)擮Lʌ]C僇9Y��x�d!6�P}i��T;���'��0Ce�Iߟ�@r�|RU�����\	�X��H'G��}R�%Nʟ��IߟD�	��[y�Nt�(E��O��F&(8@���Bq�.���O��n�j��B���ݟ��	ݟTxS�L�ANvp"�lZ��Fq��o�.�P�o�S~��ƮE�D�'��'��s$-8{0�5G/b����`�<���?Y��?	��?�����ɄT� T���H�]�Z(Q$+��kLR�'4�(`��a=���dЦ&�P�4�.�h�+��/P��ÍG��ݟ��i>�p��ӦQ�'"5A���8V�@�Fhƒ��	QCS�N��������4���D�O����=ot)RI�Q-6�لb�1R�d�Oz˓&���7���'P>��N�8�܁qIH�AAD���n7?YQS���I��$��'u���#���;^�P$�@�<-%ʅB��W�j��ts�OD��4����=2�O�Ⱥ��M�:���ǰO�p�e��O`�d�O����O1�&�(���Z\��ѫu"V8m�DSV�
��­��[�� ڴ��'`���?Q4`�:���J�&��g�살ƈ=�?���Ͷ��۴����~������.O�ST̉� Dc�'3���I0O���?���?9���?�����i@?, �t�	3	�(qc��ۄ�rDo"M� ���P�IA������T���4�!a���H����?����4(>=��:O�5�P	�72Zz�`O�'4�Q�3=O} �!�?QB�7��<���?ٱ0Y���;`���$o������?I��?����dV��A��_ܟ��	ʟ�����,5���T�R��.DH�l�����,�IL�	�w��فSZ�&���;��"�M:c�\�,2���|bs�O����uH��Ń"ήhʰ���.�&i ���?����?I��h��N���`G}{(� c�գ��[g�'0.�Ā�0�剑�M���w��52�� "ӮU(�	�3Qܢ�'X2�'���O�Wk�&��p��L���t�H4�b�s'�ʄ"EX<@$L�2#֤q%�4�����'Y��'���'�YK�M+לԒ��,BB��jfY���4+r
���?������?Q�HA�w�8��''��,'p�i�C,;���ޟd�Ii�)��\�\%�ˍ�<g�D��J�y��Kq��/}�4�?�]�b�O`i�H>�/O$�Q���	��		�~X��n'�?���?���?�'���A٦�V��ş<��铧q���.��*��h�ΐ�<3ߴ��'����?���?�2��Lꂔ�iV��:��[�
x�t	ٴ��dA	��R��%�v�����S���B@H�*hq����. �D�O
���O��$�O��!�S����p� O���攴A| H�	ϟ�����M��^�|��6��&�|�eR�W��A��% �m�̄(����T�'������A��M{�O�L��
[�#4���8�����7V����=�j�O���|����?���^I���S��D�d��Z�/k<x���?�-O�..ic��Ov�$�O��'3<T`�_�:�MBG��:��1�')���?1���S�D�G�Q���U.�z ����xH[�|_B9�O�I�6�?!( ���:̍;SJT>����QxD���O��D�O~��ɷ<�E�i�dXH2�˞<�<5�1��/>���'��$�B�'�7�&�	���Dx�h�'�C�{j�\bbX�>��ҷ�<�F���6;?�$��9���	+����2nj�!��<1��j�
����<��?���?���?Y)��9c�B;p:�YȷXh�J�	Em���)�Gi����럀�����y�&��Լn�? �:!�I��]�b��	�g�F6�y����ω{�윙��ǿ���1�Ew�����ΚX�"�O�I[y��'��Z����2noɳ�C�@O����?���?!-OP�m��2�0������n�p�n�F�qA�n�j$.9�?�]�(��i���n�$@�6/N�1���
��I�l��L�%j�%?u
��'j��I�z�8@�eË�:�u�ǌ<S�t�������\��T�O2k'/O,��d�'.�B|1����c�bGwӜ\�ץ�<yg�iu�O��^!j"C�VR�L�Wg�F����O��D�O�lpLb�8�0�\�y���q�u0&4�f*��>�!U��䓼�4�P���Ot���O���� <
$bC�x ��blS�{���Hh"Ʊ��$�OX�?�RխV-ʴ#M�R�n�P��������O���'��	T�=� �:��^2Aey�P�E��1�2�ըv/���:�Zk��'�^�'��'����
$��f���hH93�'���'�����DX�4��4>�~��g1���Fe� �̅���<�d�BQ���U}�'���'�%p�S�j�=�dE��qR�!�����tHa��D�t����L<�O�L�
1aT��-+*=Ce2Ov���O��d�Oj�D�O,�?i����L@9)��]�4��d�"��`��Пx)ڴT�u�,O$�n�U�I'2yd8A1mӅh�(В�� 8d&�(����擔ogNYoN~�L
�� �bG�ؚ�@��&֥'ʠ�"���?��,4�$�<�'�?���?iSQ't?�eá��)tXksP;�?	�������9R���d��ן��O�N)�@�8�� ��K�v��ѩ�O`��'���' ɧ�I�(oH鐤�5lFJ�p��ʡ#� a�f�7�HQ�&���S�j�Mi�	�T���G���u�"�?��Iџ��ҟ(�)�_y��p�ja��C��d�QJU�g�z�P&��!%�4ʓ~��v�$Tq}R�'p\R���>�nt��B8L�]� ��"@����'J�4����?%*�U�p�ͻ[�0��ފ(� ��g���'*2�'���'7��'�&e�x@��S� �d3���-.�2ߴ=�:y���?����'�?Q���y	�F4&�C&kM�+6l��?B�'�ɧ�Ozx�QS�i
�E�C��Y���D�8���%ՈNc�����[c?O>�*O����O8��%"zh6I;��يP�RQX�o�O����O
��<�B�iĐ��'�r�'�8cd�ԴB�&i�+�Z��\���d�P}b�'���|�ApQB ~�X����� "���ZV�x���'?����Ob�$�d�%J��H甁�'�B��$�O�$�Oh�D?ڧ�?Yt��!u�X��v��_���Ɇ-��?�F�iC��+��'�rMxӠ��]�<NP�?s�	"�þgl���1O���O<�dߩ`d�6�+?���+ ���&%���(`"�#��P���1W��M'�D�'��'��'���'l��	��F�p4�`XShS�$��x�%R�8�۴6{R ���?�����O��`C���5�a�@8i��h&��>Y��?!M>�|2�!N	r�}Yu�G32�Ȁ�蜥3�hٴ��$��d��H�'��'h�I) ��1���SĞ�h�'O-^�����ȟ8��ٟ��i>ݔ']B7���L�d�4�R|�b�þI�tp���e˂�$�Ʀa�?)�Q�h�Iݟ$��~$�#�!}�M"�+�Ҷ�s�ȦE�'���¡�?��}���#���5�Q^��a�$OD�F���̓�?q��?���?Y����O��0�De�2Z�����vK�iÑ�'Rb�'�@7m��l9�	�Ol�d��̘x��V�\��%!ס��(�%�$�	ٟ�=h�h�ld~r��+3"�����Q�Q�vͅ�LA<�;D�PN?AM>�)OR��O��$�O�ru-w�/E�	lB��A(�,2�z���O0ʓ��։O	k���'��P>��ҤF�(����ZA6�k/?�rS����֟l&��!
XYGj��mmL� %k�e�"��V������y~�O�	�	�s�'҄QA6��l΄�:sG�*0����'�2�'7����Oi�	:�M{$$K.�H��nH�T�
��'҆s��Q����?�w�i��OJ	�'�bB!>oȧK��k�D�a"N�V�r�'\L��iI���D7�����O��aL0���,Mr2��4����Γ��D�O��$�O���O����|�4S�7�p�WK�	-4N�V�X'V��@*.���'���'� 6=��m�@�Q�4 �V�N3 �d��(�O�� ��IF�MK"7M�;�ꌪM����qoϢu{҅3�'z��ڄk<�'j�	}y��'����*%������D"�V��s��_H�'[��'�*�MS�\��?)��?I�nB�z�C�]? �̡��*��'/�듿?������&`��R���Ԥ:��'(N�1G`�`�2\���4A�џt���';�5�
zx�
4����'V��'$��'�>��ɧv���k۷u��{�a�) �L����M������d��i�?�;=�s�ؗ>�\q; E.~�����|��������˦��'�H����x�T�_1R�qPç3���0�[��䓲�D�O��O����O�����ţ�kB�$x�%!�`J�n ˓͛�B�#PB�'����T�'�����Ɓ
U�hX��CR�q�A�3��>���?�K>�|�
X,JFR���4`~�d�2�8�f��bda~e2z���I
Bu�'~�	�RϜ�w
��H�u͉�Ӛ���矴��ß��i>e�'447mH+_L���тzj@(�/� E ��!dͱ��LŦ��?�Q����$���C6Dx�����2�"�΅.:�
�2�
�æ��'���+$���?�}����}���դ8b��AE�?_�L̓�?����?���?����OU,p
d���#lR��#�'��'�~7mH$J��i�O�m�~�ZL��� !�1�Z̒�'��8F�c����ݟ��ə*��]lZ�<���-��������h��b� 1���p-��X��$��䓏�D�ON���O���M���G$���ԙ�Eǋ+t�d�O�� ��ԽFI��'Z�S>-�hB/��yT$�P)���:�W��P�O��d�O��O��l���СE-"�LE@5'	$!�J ��M�(V��!2K:?�'[�F�$�4���(D�1�N&bn(�@�R�_�����?Q��?1�S�'���m����8����W�[>�:&(�$rN�����0�ݴ��'�n듏?�g��J
i���7AY�q�X��?��������4����i�g��
Y�+O ���ħ?�P�;��>� �y�4OD��?I��?Y��?i����5}������0��� �� <�oZ�:�������	h��0��w�:@*R�Yl2�2��J�+����'B�|����)���6O� �L�+�$$1���JBeJ;O"QÌ�?�4���<�Og�8�fT�U�pao��p�<Ó)��⒉p��ڟ�����rV�,iq��>(N�8��RN�i���,�I~�ɑ�q0�Z�1i��_y��/cf,�T�P1L8�zH~rtB�O�2��*ܐ�q� =ȥ�1ņ9���ȓe"��Q���#��-�N�	q78P��i�v@?Ex�'q�6� �i��!���9���3�$��r|�f�x�������I!Y���nW~Rk����I��,�=��@V�l����Y.z5�H>�)O"�?��R"C�t�E�ɝJ��0B��El~�cӪ�Ө�O��D�Ot�?!0�A+IrlSr�ߜ�$� 5
���d�O��d&��錞Ykr��qK$0^��pN�`n̵�5�}�A�';�r3�o?�J>�/O�h��բ,GZ�Y�+ɺ c�-���'s�7m�U(��$��ny�a��C�)c�*�
ro�5��T����?��]�T��؟���;I����G���[e�~�!6d�����'�%�奎�?������w�p=!v�ܹ��}Q�JGp
��'���B�#QlsGj��Vr(Q��ѕ|+B�'�2w�x\���?���4���PȺ҃�%ws�ٹR�֨z�H�sH>����?�'����4���04�N��E� 1� ��G�t�!�
�~b�|2S�\�?��U� F�ؐ)��$#ځ��co�'�$6MX�V���O����|2C�$Vi"�	�fi.�ɲ�Ji~�>���?QJ>�O:y���A8�j婦��17����7+
j�"�i�$��|�@���l'�t��F����2 �A(�}���|����I��b>��'�,6-V"�j$���W]����1�V35T"I*�Oz��ئ��?�rV���I�;��ͫ�!�>"��z##^����I����3٦��'�*e	�I�(O�L���7Pg���̌2z���2O˓�?���?���?�����BI�� Ť��j�{Ш�/�l\m����'I���d�'t7=���w��z��A�vkG��̽1���Oz�d?�󉜢I�t6�w�ВW��"k0^�kՊ e�\5� �w�,���<V���0��<)��?��'�>"pH3��Ϟ$�e�L��?)���?������æE�Gݟ��I�#��� �,�u��/�(�#��s��]��؟���n��a�~}h���CVR`��G!,��7�,�@'I\	�M�4���o�y?Q�cܪ��NM�e2d	s��)����?����?���h�����P;�P���'ޱz�g��:Z��Dަ�����d�	��M��w��S�
�9!��Q�×	gsiq�'E�'9"!E�<�f����e�ٙA^��" ��㓍�A�0����� >ޓO6��?����?a��?��i�H��+C��8��TCVA�/OF�oZ2'���I�����G�s�L�v�{���Ɓ ,pt�������O���#��iZ�)^]v�Y�K��pZt�+M��P�`k���'�X�i�M�{?yN>�.O���!��Y�F�`@O:��X���O����O����O�)�<�G�i&��p��'n�U��ؤ�lw�GEd���'�7�#�I/����O����O�tZ�fɾ4Xƙ�"�D8]<�F�-wV7�%?�P`�6���j��ߍ�c�I�/�޵I�,vż*��È�yB�'��'2�'v��I[�RQxl�q�Π��I!��·3����O��$�ߦ�)�Af>���
�M�O>���am� ˒', ll��Qoǉ���?���|���+�M#�O�yq��И�����VlB�$�t^5i�'��'��	���	�����	r<�0cB��y���� Em�m��ǟD�'9L7m�86���O���|��H\�kkn]�'aX�'~D���iGy~b�>����?�N>�O�z��f/��8sE���!R�ƅP��:l`���iL���|J#���$�Ĉ��Z>��hA
E�ma��/=�,�ڴ|��e�P-U�q���-��Sh��]r0U��ğ���4��'0���?����6ZnF cAF�[+��3��Ŵ�?��Ee�d�ڴ��䖛1�p�1�ON�%\p5{�A]1D� ��"�_Mn��	sy��'���r���:0��&ĳzqJ�s$Jl��@G��<����O-@6=���
�DC�&���	�٫َ��q��O4�;��� �F6m`��¤�3�����I�hpAHj�0�)ψ��S�	Hy�T��;U/��B���S+��T	�<OPl��\�:���՟��	;fNaS�%�v�"1#u�

z��?�Q�`�	��8'���'�>"ʘ�"�	�K��{�F*?�ED�$��%1�4��O^4���2ܴ(�:�`bRg�ܸ1�
�7��D�ȓns�d  �ٖ#�l	g&Y�(�e���L�v �-�2�'��6�'�i�9rE �o"���$O����"#f�(�	蟘�	�/}^�mZ]~r�ƭt����mB.YH�H�9�A�կ�j=�L>�-O&���O�D�O����O�����6"M�ȸ7
Ԣ=������<I�i2b��'����'Z�0�����#!�E��3��>���?IL>�|�&"C�? Z�jg��)n�(���ɚ{(���E��sR�	�5�P0��'�0&�<�'N�c��T8ty#����(e!��'2�'R���tR�� ܴJ���X��!�2��e�c�XD�s�[?^�h��@[����W}�'��'Y��k6����"D�#�[) j8���ҁM+�֔���B_�i���8�I�����s��fR`}	��H�9 P�t?O|���O����O��$�O�?���I�?0qJA��a�1w��k�E^����	ן��4Z����O�6�?����H>�����#,�N8x&5�|�ON�$�O�>B�7�9?�e%6��h�%ѱ<��9�&�����C�$���'1�'e�'b����S	FpCb�%Q���#%�'��T���4����?�����èU����)�h���hq�I�����O��.��?{VK5m��X"r��bU���CJL�g���ĭ	ߦ%`(O�)J'�~R�|��̕��4s��y����"�t(��'�B�'a��D\�\Q�4q9!c��J8$��Q��D��#�?���ge�f�dX}��'\�( eI�$vT4x�6+�O"��h��'�r��IX����T�"����I�<�VI��ղ�oX1�(�ψ�<�,OZ��O�D�O���O�˧ϒ1�hީYo�M�dA�x8j��0�i�>x2�'���'-��yªg����pn�5rr�����	L
7�0�D�OؓO1���ԍq���I:;!�k���j����dC�<j��I�v�Pɢ�'<4�'�ؖ���'u�V?w\���>�"����'<R�'��[� ݴ*6� ���?	��!Ϣ��7�G<��{!�C�1 "`{��>���?YI>�2bI
Z�v,�rn�	���Q��h~r����r��Om��	jP2DƤn�hPÉ�/��$bCʇ;gk��'��'���џ�㫞�����DM	$�b���ٟ ��4(�@-���?�a�iH�O���-KN"YP�g�*K�t��ᝉS��$�O�/����4���M�4ʑ��IN��gg 	dΨ�u�� j(8�I0�$�<��?q��?y��?!V��@\᥃����kg'�!��ĐŦu;��_��|��ʟ�&?y�ɚ	4���#�6,�ȉ��7��ܰ�Op�D2�)�$X��pE��!2�����U�tLn��T!:W1T<�'���ğ�Pa�|bR�H��Z�A�E�7�q	�&�ɟ����������S~yrL`�N�� *�O�xa��S�؉�R�]'~��[t8O�lZy��,�	ӟ��'�{�K&d����3MϏ<.\�3(ϓ#�ƛ��H��F���	q��ߑ����s)���#�H�x���w���	���Iϟ�������Z�˳P|Db�ƙ�C\mq%Iϖ�?����?I�i�9вV��y۴��M�Q)"	Nt�T,�ERD��<���[}	�6�&?ل��X�D	�%(�`XHd M=9�uJ���OJ]�H>y(O0���ON�d�O����	7$�� �{>�,���OH��<1s�i ��� Z�<��V�� V�w`�A#Hy6��O�����s}�'��O���mw�TzU�W�$�^��үC.zB����$OX�Hl[Jy�O�j܀�d�QX J���:�ji���I����a�K���Ğ^e�T�GQ6��E��$]x�	�L���dp&d�g�2���Ʉ�E��aPV�Ӊ@Z�z}C��ג;ͼ�H�G��HO��t�D,d��E눞a�N�Ci��X����*@�ڽ۳�� �`�)�Á�b�/߾7o@谌��<�92	�<l�
�0��4��x�7}���3��V���Y��
hxj�3Fh1y�05j I��w4��`F&=i�^���?�\��$DF[�%buIҔ/ � �E�"Q���%���� �����O��O����Odhc�H�L���4aL�y�%H�'De�~�O����O��d�<�D���df�iU$�ܠ�"#�:$��iN*]���T���IW�I֟���*D8 ��f���IdAB M��r�[�w����'"��'��V���a�X��	�O��Y�H$d�z�#��Y=����F֦���G�͟��	�����=y��N�x��)�R�̌<�lI�c��Ʀ��	򟘕'�LL��I�~���?��'*��6꘬l��i�p�ՙLX�D�x�'(�k�_��O"�S5,�1��&��E,���F�_!u�7��<!�΄7a����')��'����>�194XH�ǠK�\_�1�Ē�v�T	lZ˟p�I<H�D�?Q��H�����[Z�x��jݵ�M�@ʝS��'+b�'����>q)O�� G�#P�;5m�+(�p܊���!iDDv����O�"�Q&愺�E< X=�P�G>�7��O��$�O	���q}U�0�I{?�K�\�iKdM��w��I�C�覍&�̡,�Y�����Iҟ�'�M8�\%_�ʐ�c�Wzh�7-�OnuK�k�Y}�V���	F�i��#0��z�xz�(�9�fq ���>���9�?Q/O�D�O��d�<Y"�A�P��TP�+G���@[�I�*���K3X��'���|��'��nZ���Ո�e�)`,�#���������|�'�"�'_�I� �4x(�Olp��
L�g���T�@-
�P�#ߴ���O,�O����O�"�n�O���BL=�tͣ�f�^̴�C��t}��'���'��0g��,�����dL��P�02�ɴ=��%�1�պt�Z}nZꟴ%���	����6���^RD��QC8M��(�6#[!+��7��OZ���<�2� /]��O1R��56�	6O/n��P��(-�,a�ě�����O���:�9O�� �E��F8S9�%�@!20�D�i#剼Q�2�ٴE��韈���� �n�4B���VP�L��@߈ ���]�������xL|zM~nZ%+]���oBz��v� �,��6MW'в�l�؟�������S����|Rq��	_�NU f��eM����3i���'��'�ɧ�9O���Ц`;�غ��`�6��c͗�L�.qm�۟D�I柸ALԟ���|r��~� 	,!ʥe�;\��}��Dߋ�MK���� g�3?����~ǚ,h�5x'ͺ@P�"��M����X�Q/O���Ol�OfA+�LV�s�ѸF�C?=bu�qN�c�8��c����ty��'҆�Z��"<oV���h��r�:���5u������	j���?I�'�.��� 		s<|��NI�h�dm�ߴ-i���<	�����O�4K�?���i�2[>�dyU�XF��m	E�p���O(���IEy��5�M�#ɼ	B� ��+J�2
�@Ӳ��[}�'IB�'�	4yv�H|B2��lF�b�/�:>��tH�fS�����'��'�i>A��h�)�/~�$�F�� �Tّg]�2����'��Q���a���ħ�?9��s��ܲ.��p�$<�J���Ol�	fy��'�B����uGĐL��AѦa�GO��E����$�O|��AG�O����O���㟦�Ӻc򠕅RM�0S�#,,�PcbD@����IZyjŬ�O�OZ"0�v���)o�4�C�f��m3ٴ"\���iz�'���O�O����v&o9ƕ�G��s��IT�i�"�'ub�|ʟ��O>�ID�@��)��f�N���`*H�����6�i�*9��6�4���D���BTz�xp"��#.��P�a�
�6�$�C��'#��'c�BT�c�@�:@Y(kc˿R��L�ߴ�?!�M�}"���D�'��'�@�#��;7V\�SDF:A��!��I=�d�OT�O<���<���D��0�/�8]�RA�~Drpy'�C����O���5�������s ��9� X�~_�}���w}LoZ�G����?���?	.O 4���Y�|*�b��|c� �lBh��1jW�	q}R�'S�|BW��S؟ �p`S�j@$Mx��<���������?a/O0�dN_���'�?�P�gX u[MZ�[?h�:���nx�����O�$��<%���Ӯ#ߘ�6�4�'J�6��d�<���O�a/�r�$�O"���Nu�&{ҙ���,}|��c��x2�'���	g7�"<�;?��yH�n?:Aƙ�-7�Z0�'�2�@(hD�'�2�'��TT���<�y��K�$>b68���d��7��Ov�r�v�DxJ|r'���eԘ�J��0~��`4�զ�#f�̨�M#���?����Zb�x�Old�o�8B^�iTę_�" �h�����O���+��?������S�ۄ��i�ю��r9YD��:�M���?��Oy���x�O��Ol�X3��`�"����[����?N>�*���O��D�O�L����Q����O\���� Ǧ��	*��i�I<�'�?�J>i5#<J!@q���8TFhA� �t�'�RZ�T�	՟l�	iyB`~�X��NR<�C�.ݿZ�H%�a�+��OP��2���<��_�����L�1ne#Č^8���nZݟ<�'���'&�T�P bf������jʾ���'�3_&y'n޶�M�+O^���<����?q�$t�;�de�b$Ў{DT����;E#8�pAZ�H�	�x��Ky���8#|r맓?�b�F�Nt�`������&�� ��&�'����� ��П𰑥h�\�'0�at+W!!C PXF�H�+ނ�;6�n�,���O��5�~4��[?�������ө\<�09��Q))H�9����/_[��@�OH���O|��-UC��cy2ӟ�y3M�&<�l	�r'BB�Ѡq�in�B��49�4�?)���?Q��Z��i��4�
�1R����I)=��t@w���d�O����5O����y��I;��p�ۊ4����"`G�OS�p��6�O~�$�O����Y}rS�@����|�& �a<}�P�9����M�Vb��<�O>����'�U���Oh̡�2|;�2|��jl��$�Od��	�����'�	˟��z�4J7�� o�lk�ʫR�ftm�۟\�'_V����I�O.���O�4�#ž)�z�`����[h�6��Ҧ��I�bav5J�O
��?�,O����Y`�
=㡌��J ���^��#�}�P�'�"�'�O��Mj�)� ��=+�B=10�%�Ƥ�6eD����O���?���?	g"!4LY��N��X�����,A>Ɔ ��?���?!��?�*O�� ��X�|�C��=P�����uM@�괩��'�2[���I����	�^��牘7@�I�QL����)���WT!I�On�d�O��$�<q���4V�SПL���;���P�!���bE�D���Ms����O����O"pS�0O&��]� 8[�E8�HHM�V�rM`���d�O��>}�pP?�I�8��:�2���l�!�\i���<@��0�O�d�O���?\�ı|b�����Z�qS�Ƅ5�2�����M3(O.-#���ߦ���ßt���?��O�N�����H�F��� ̕�<����'wB�	�y�|��IT-5\�vd�.�<��4+�/x�6��9(�6��O.�$�O�	�Q}�Y���Ad�/� 6
i32��M�C��<)J>�����'�� $��嘃^H�C�t1�#��i�R�'i��cܴ����O���;^��}�E�4r��(�PE�L��7�2���"`��?=�����'C���k��[Ɉ!�h߶9�b}o���l�����?�������O�8D�%�R�.D>9�@�s}� �	�y�Y����ϟ0$?)9􍕗����)��L�P ���Z�RI<����?�M>���?�J��m���z�m�/
�n�Xq��<U$8Q�������O&���O�˓e�V�r2��U�� �=.M3U��	0���`�xr�'q�'*b�'vN�+��'yވ����o+"���+�:I2��.�>q���?����d����$>%0� Z�?�{�cđ�(e��A$�MC����?I��m�8x1�{��295N��e��S�
d�t�E��M���?�)O����JD\�Sן���69�=a�@ÚJ�pP�# ͅ�H� N<���?90�R �?qK>��Oбs�ٿn�%�0�VR�\Xڴ��͜B���l�����O��iM~2�K�r:��	֢,o��
P+��M����?���<�N>������2�D��%D�QX��vV�2p��V�~\l�����	៸��1��'�4$P���,Iu^�`3E�0]�x��y�\,8�9O��O��?y��;X�MX�do� �`cV?�BP��4�?	��?ɶAV��'���'��$��K�����X�2iJ����V�|R_
$�X�d�O��R�G���S��d����B�B:U�!n������R+��'�|ZcE�t� ���;��0��l��k�O|�@���O�˓�?a���n��4BD��������>.�p�.U�6 �O���/���O����g��4  ��.c�$8��7������O��?��?a(O ���oW�|���P�VQѰ���&a��R�f�L}��'��|��'��ߜ�oͱn�&lC��.tt>���@	�2�T��?����?!-O��
��G��	4h�ە��r|鹐fK%L��A#�4�?9+O(�$�O�$�E��$2}���*���÷M�R�|�ؠ�>�M���?Q(O��d�U��ʟx��*��xp'n_�p�|]"D��x�|TpO<����?��@��<qN>��O{�ٵ�� bz�<����2cc�m��4��$Q0�o�5��I�O����q~���nFإ+�����bu�+�M���?1-��'Mq�؉�t�H:^b�2��Y�1@����i�̰@'&l�����O���4�%�l�	�c�4U�J'��X�v��=��4q�" ��B���O~����ͷWKD��'Ӿ%����������l���`�8�M<ͧ��	�L�� �Q�P=������|7m1�	��'�?����?�tE�>Dr�tP�܌@���DD]���'r���<�4�f�<�W]E��Z� �U�荨%#KD�ܟ��'���'TbZ��C���;�|����$g?$03M�7�Nm�K<i���?Q�����O|�$U�^?`����O��T��R�e6 u��O�d�O��:����0�RԳG�ۊ*�d�;WaƱ�Z�@�i���0�'�B�'�"�I��T:G��@PEQ�t�3�^	%���ԟ��Iџ,�'��	�X��i�O�+�"0 ��怖��y��̦!��Dy��'���'�#�'��SwHD���[�c�Y2BK�4M8�q�4�?i����M7}%r@�O�b�'4�l��!���ψ1�\ aMQ*��?1���?I3��<�-O0��?1�ů�<K�b�A7 �-=��b�c���m����i
R�'���O���Ӻ�WFǴ$-BY2��͓�t��Z�l�Ο��	�l��I ��I�O��>c��׌H>����㒎>wq8s�rӊ}�)X�%��ߟX�I�?�p�O���"!ڠ�P##�0+5ȗ�f�L|1ָi�ԓ�'��\�`�����)�g�l�~p�w'W�X���(�i�"�'��nΒ]&����O��I1<JuB%����x���O�6��O��O�ȁ:O������I̟�(���>�l W &]�րS�N��M���MEz �[���'�2W���i���6`'g���/s�^t��I�>����<�,Ot�$�O���<'�w�Uq�n�X'�+椃5 G蔱�P��'!RP���	���
"�h53E�5o�y�Wm��1m��@t�H�'��'�2�'�"�ձF��閥Zb6Y������	���N�B.�[����Z�I����'z�!I�4M��8��a;K�V�@2
�2q4l,�'U�'�rS��ia,��ħ?��	��Y1���"l�n�LUmZԟ���U� �T�~:��Pi֔#���k�4p�L�ͦ9��ԟ���П��a���'F��O����2�]J�w�V�L��ѐ2�/���O�'�GxZw�x� �#�"���$��&�&�zڴ�?��]]���?���?Q������]`W끹e�6`���:�2�2F�i��\�,
`�+�S�S�$%45RqBN�(�P��,I� v$6M n+�mZΟ ��ܟ�����|ҠI� T;���� ~Ԅ��`?ӛV��>C�OV����O��8�G�I�~��DW@�k0�P����Ny��ʾa��'>��ן�V��l���B�.��d��m������i)$>]�I����I�-������D
k��[�Q�"A����4�?	G�2H�O ��#����)"k%1�|L�$�W96@� S�иá2�I�����ꟼ�'� � �a����`U2`�@��x��P��Of��"���Od���2!�L�Y�f�Q#�ېKB	;�6XI��D�O����O��]�.��W5�v�X�[��W ՌtSG�η�ē�?qN>��?	�+�R}R��eX���$�_��N�6������O"���O��$�O�) ��|��'\����N0Ktv�(�3Q[ļ��4�?�N>q����䘆 ��',�PZ@�W,k�"X1�eʙx5JA�ٴ�?A������>|� $>����?Z ��/��i�bK�(�Y��#�M{��c�����i_f�3�K�HU@ex��}�&��ݴ�?����а��?����?��'�?I����/�TA&U(�-��Fxs�B�����dy�-D�O�Oޡ��J��k�εqQ�F�aV
��4`M���G�i7�'3��O�Ob�$�?NLȢpF��e��٪n.<�n�I
"<E���'d�JǠX����#�|��cG�sӮ�$�Or�ĀD�}�>9���~�ϔ.*�����A�'Ȅ��p�����'�h̻�y��'�R�'���qb�͒]�&<��Ӻ�d�P����DH(w�l�>�����+B
I��i����.肁���`}��:��'��'�\��sT�ېC���39����a[�Od��"�}�'��'��'\*�āP/y%F�p���5oy���恐ܸ'���*���5����?*�vɒp	�<��p�cN�"-�DL{q�A�9ޔ-�����hr�+�'�Hk���[�����kn��H�{"�H�6�~���`�i�n��`I�1IH�˳l�C�M�+B��s
�'��#��>�pp�eٮ?�8a�
 *�@@�*~=[����Q�a��
��ЉQ`�4�� n�e�*X�4�I�^�Y��+��Q#��R�yczsSF��4P,Y�H�*P������1�?�s�"ZD�(��&E�:���ɑ�?!��zල�n�!;��(`�ώ� 4���M�?e�O
<��E'�X%��
+[
8�2K��3aE�a��苴b,�H�ٰ"�H�ͭ|JBiT�.��W���zgz����J�D�-���'{�>=�I�[sV��ģVWͰdB�ʀi�B䉫*K,A`e�B��xT�DkI�f����T�'��H2 �&!��1�̥ ���T(�>y��?1�*�?��%���?��?ͻ+7���2� p��Ua���]����:R�pD�'���������Imб��h���D�"P��Eo6�� 	]�>�:��'�da�^B�g�I�>�25@Я
�4]z�'��7�����O~��O��?�'�hOP���mi���W��b
R��y"���E�J�!�,N9xEpUŐ���c�����<��B�Q�F�J�"41���"�;׸LP��[��?i���?9�Qd��O���`>�qF� @�ZpJ�融CY���g��T���s�H���,a1ۓ^���(Vh��"��,qGW�D���fQU�vt!h�
@Ua{�
�rj����O�8�8,�!�њV8"}��?)��d(�ɀP|P$�d��S�����;L��B�I���l�3?���e�E��b�4�O�'B��z6�iB�'�4ث�
U�l���9�ON?$�"��r�'�������'��靻Z�2�|�����@�➫
al@`�d��p<����S���lTC J �w�;yeB���ɱSY��>���)=�4Q�PM�|�B�_�!�d).b-��. &2�<(D�!A�!���֦;��b��wX�`F��a�"�	(���4�?!�����T�2�$)dH!�,N�Syl\h�W!I��'�l8Z��'�1O�3?�aB�=`b�5�X�1���L[k��ƪf��?9�A�����BeN�x��h�i6}�J� �?i�y��t�C�C�˳��@����?�yr��bj1��i�4�4;�Ɛ��0<�鉋0P��bÉL.qdHtQ2��y"n� �4�?i��?�ӌ��Nə���?���y��J���Q���=[��-� ����y�B��<Q��RLe21R��7)�E�Sm}�7��u��I5L^Ds�m(eD�#�r��u�<�W#�ğ�>�O���U�X>k?6�(�.
o����"O��"q�B�� �Em�!Zϼ�ɑ������ᓗE��dRp	v�@J�	V{@t��������'r�'��dq���	��\�'L�L+��U�8A$my0E��L��0�b��m<gN�$\�!� Fuk4E1C��8<�N܇��_�a$ǖ		꜊�O�2�z��f�ןP��	�S���2DIg��5s��ժJ��C�	�O�����DmҴa��a\��c���}b�%t�7��O���R��L��kƸ��e�4�(�$g�cW��'��ɍ�Vfb�|"%R=l�{����0��T �$��p<a�jX[��`�}ʳh[3-&@�#��j|���	�oͼ�D(�� �0	U�Y���f�H�
 T�jp"O�h"�.��CC0�Q B�1 �)��O(��I2�ڍ�n�05��:үV�/�1O��&�Ӧ	������OJPa��F^��A� +��H��Ư1RI;��?1RK���?1�y*����r�#S����XZB��8xD|�'^<�����I�3}T
(�5CӶ-�N�:��ύT��n_����\�S�'+��ڡ�>q�ȠF�3�
M�ȓ6���93��>�jXЇƃu�,]��	&�HO�8� f�8M�6�r�ؾ1"
a�c�Ӧ��	㟨�	�dM�dI�NL�D�	蟰���k�Vu:�+�ՍI���aa��q�j�"��
N�|A�@�K1Kb@�c	H.�➔�Ǣ/<O�8�U��~M��giܴ}�j9�H+�	��b���|"�B?[�l �K��y\�l�J�*�y��E?aY#� D�  �����ęk���0ʲ�C�RĬ��#P'r�x���1 �<�B��O>�$�O@�	Ѻ����?I�O�^h{�iK���i#d�3kt%�gΣ�xbeD�;����&ت�"�x��:t��ؙ�'��p��h?2uJ��.�X�UC�$�?������D�K8��}���ׇ<*��(}f�S��I!0�vAh�K��R	�<�v���k��nϟ���A+V�jS^-U�М���� K�T���<i� ����I�|R��S���'�X!��?���l	('и�q�,Op\����*s�v�;Rb)��)��g��x�oH��?J>!�:���z����t� %�3b@�<��dJ�U��Sv�F/g u�5J�x<IA�i�d~JP�+�.a�
@9��ʲ�'�`H볊zӾ���O(�'i<�y�	�~~�Iр�ÁN^��H�%�9��̟\��M�0�<����T�|����%�3N"���H�&��E���Ex��dl[.Ҏ�觩�	:�Q��A���|�>�)��#���Ņ���8'k�.x�C�#c�iZ'@JD�"<��ѝY�t��E�'jn����L��D��,@�J)��Ʀ>i��?	��'E�
Tq���?����?�;@L<@�!��OЈ���d��N�kJ���ǅ�:�Yj�K�1��'�|@B�Ɗ{��}�#��-�FЂ�,+���W��={���v�g�-o\��Ckг ��Tp�|!�
�O����4�ܣ=���R��U0�D�d�a#pF�Q�<�$f�(U�b�i�/��*��A��O~"C �S��V�`84��1z ��U�D�Sr�3)X�T���P����I؟�Γ�u��'v0�܅�@#N�W��cP"O��!5k�6%P!�Ć�0�p�c��N�B��־D���bO`���l������U�g�������'Az���O�6��0(���86x�\��'��i�d�n��T{���<n
T��ybf7�	;c2,��ٴ�?���{C&Y�'�.vɒ�j�>$���y"	�?����T5�?�J>�����A�p㞲1�lk1�E8���ŧ.�I?Y�����E��@�ıU4`���>n��|�7ᶱa�?T�L���O��y2P&
t|�į�La��6K��x��o�4��N�{��x��� 8���f�F���oZğ���R�4��1�?�4���EY�tH�X�,����'HO��?Y��\~^E�������',ل}�My b;j&�b&�)}����O�v%�鈆y�"��v&�c(Z �>���Lß,�<���
�m�@�A!��- ���@�_�<!�JG�*\�0�Z!SP�I�  r�Ĺ���_*�)b/��5#�5o���n��L������j�?Y�2|��ҟ\�	�<�ݕ��\���C�=�t	W�I(t�jX�<1�ADqx�3�J�D�:x�5�ҍ"�`�u�$� Pd���0�6�y�gT�Sy��`@旟PG�c��@@f�Oq��'+���Q���5��"ҋ\|߶y��'Y�0j��Ci�,%ib�C�a��P�Oj�Ez���[
ZX@9�cR�}�Du�@�2G^���B�1$�d�O��w�<���?������
֑I��5x�!+>�"����?�hٸ�'�(�٠�\�zT.���~�&�ל���������@A�ak�M�T�;����KΟ ��)� �a����	F��RA����S"OԊ���l<0y`�#ܯC�H�����P������i���'K"��� Rk.e:�kZ
T�a��'������'{�)�;d2�|Bi��B�<b�"�<?5�S�$�p<q �R��1���qa�ҝ5��!�sH��kR���I�Iw���.�dT�r�����Q=�!�gʈC!�D��+<9�0�S)10x0��ɗ�+B!�R�Y�g�/3���r���(x� �bED(�I+Mw֩jٴ�?Q����i�,!\�&C�Y�'H[�}��P�c��'�:9�d�'1O�3?����1��LC�n]�Bu���,M�D�L���?��դC�n���e�W��-*e�#}b+�<�?�y���$�9�� ��pn6%{&-�e�<)�.�3[Ȓ�	�Ì�&��a��c�A�$�����+�$!h�g�[�A���0�d|lZ�0���� � (���a�I����	�<�ݤsk�X(V��5� +E$E	I��I�<��HPx��
N�:Id���4LҠN����8~6���W�PY��M�V�޸Ч���[�vc���!�Oq��'lI�χ*��0�B� >���'�%鐄�&'��
�;H�C�O��Dz���� Լ��7䙆v�a����$cc�l����C����O���i�����?�����ą1���@�Ǆ/k�Z|��H?+�$,��'�Ndi�]�B�N �d*ӓ���
���xrl]�R0��$#�yz�"��D_�E����?e���N�����"n��2s�Rr�<���2-Q��	�7�*�RvgG̓H �ON��sgR�����$�e�����5/7�t!�"@��(̓�m��ӟ�Χ?�\<��V�	7��eD^�wq�Q��� ���^
O��O���� S&�4�T	�l9���'�D�����5a��c�H֩ue���`�(@��ȓl	8I�"/۫l��Xe�9얝����V&Q'ߴ(��*�#�p��,���'� ��`�����O�'����I�m` ��f:X?F�҅��$'1���	�������H�<�����>ksH�3	f�uQd��_��!E8Fx��DN&����/�"���1��#��E��"�)�Ӎf$腪Eǘ�m�bl*�i��H��B䉅q߰\��dT�"�|݂r�
�v��Ui�'"��� /8"�!�cAu@b}��z���d�O�dR_�DD��A�O���O���کjB͞	Z<�\��P�F�>��7�=�q����$L/I^L��2Ԑ�ǭ́f�qO�M���'�����¨C��(���ҖK�v|��җK���L>):�Z����'GF�&��X�<y�'Ĉ�"��Ό%`Dbp��M~�+.�S�O��$��V��$�Q��?D�D�A��`9�q�'i�'���f�q��؟ϧwh�����K^�%K��ܟh��\�*�v<� jƀ|��� '�?T��u��S�$������R�낹.�칢�MՒ!�	cc/韸��I$#�R��V��<rF��7��ȓm�N!�pG�<U,�p��(�+����<QW�$u���oZ�� ���EӨ�@���v�B�B��`�`����<Q� �d���|zM矔&�����tւҧ��Q��6	:O^�jU����D��JRcT2N\<\�c�˵Ej�xR�I��?�H>12��g�l`dC�1xl���[U�<��	�l+��z�,�`��T�!��N<QC�i����GC��|"l���>c�����yҌ�v��6M�OB��%������KՅ�A?��gI��`�ÀH���0�I_�<���y�S��O�LC�GT�eLD1���%K�, {G�>���l���OPd��	�
� |pv�2B�u�L�\��l�O�c��?A�GiGL*��F��M����K0D�H��F�� �c�՚.d��{�!"O��GzrF�/��̀��(K�L!1BM?�b7�O��d�OZ�Q���-O_"�D�O���g��N�?tAHF�5�-Ҡ�[�Q׆b�0�c`7<O��R��%,D��J6.���!���ӌy��yr���|�������	Q���e�^�1O��%������ �_/��%�
�+z��t��S�? N��%dP	�y1�&\�q��Q"U���	���S� 	�,�$��A��l����9)I=�D#J2>�b�Iџ����<�_w���'��Iۖ�Ԥ�'�ҷ�l�L�U���OZ���x��9刎6]-l8���'P�!�$D���n@���K��8�����'��`��g�e;�OI��)��)�y�j@�&��N�����*p(�y�?��	H�L�۴�?��.Q���.I)R���A	7#$���?Q��>�?��������d�rQ�O>ᇇ�<xM:�#C
�`xЀ1`7,O�`Aˎ��'<FV�S�pPb�ɗ���D��NLTp�	ٟ|�	Ο��)J�f=�ݰcۺ:�@�j�aViy��'��O>�`��ܜ������?|48��>�$�۴"7�U�Ve^�]<vt�'�5S��͓��$�s�DHo�ӟ�	e���?ObȚ�m���ԢĤ9p�p�Kܒi���'=���@�'�1O�3?a��˟�R�꛱]�~8Ђ&n����"<�� �89��l�p��.5h��k� 0r����*>^,a�GǕE{(<�<�e"O�ųS�J#0�`)��i�*xj��'��"=i��X+j�ltc��J5j�`סFI�<��M�*+��SE�/w���	�n�F�<	e��E��ⷢ�Q��)%��C�<IRPP�12�B�X�b�R�� J�<�Di'eL�!k��a��\�z�<a�D~b�;��:7�(J�%�w�<i�F�'�:� �; ~L;"fHs�<)�ea>�Z�9J 8�k�m�<qd��	c�B���k�<t`��UO�<��#Өc!*�X�HU�j�tP���N�<�7Mͥp �Q�7-�*��aA�LI�<� dY^�Fu��H��"���0��^�<)e��fݰّ�$��V�T@���QO�<q�o-�PU"F��U�\-3�	YG�<��<z�r� @�Ѧ ��$[��AF�<Q�*F#qm�jU��/q��C��x�<�f#ޡ�l-�&��X��Bm�t�<��>[���
�aѝ;&�CNEp�<9СI���di�P|��"'�o�<9�����= gW�
Gx!UN�m�<)�I�k��QW+��.|�@���i�<��@ j��I����=�T����f�<�R� X������H�4*�A�mFb�<YAסFfd�y�h�5'&	�ǯ�w�<���n���D�Њ,�ǉ�|�<�Ec��O"�q�J̠O���8�_�<Yf��g,04ȕd���D
E]�<��MQ%o�vX�2cW�C�
��i�X�<�bo�$DE��l��i(��ԂTU�<�G܍o'l�Y�_0��4�A[P�<����H*ͨ�N��4TR��"��K�<�+�2-Zn!�2*��j<�Y��lBJ�<	�i֐�L�4��VQ�`��c�m�<��
�2U����GϫR� Gm�<�e$ �q~"�je��DN0@:Ӂn�<�hϼb��)��aکM�&�9ddOq�<� F���u[���%64JS���c�<�ĥǦh��	9��6KV�O�C�	&VdP��C��=���ˀ���x��B��gl�IKAMl��%s$zB�	�V��÷G.*��U��R 4C��'V�4�æ�%�NYB�,^&:lC�	�4�v�B&�%I�&ufa�Aa&B䉥v��yA�.hA�(YH��C��!|��eJ��P�C��1	Ui�C�I�|1
�I�72���&m�?n�jB�)� �d+ �H�Ep1@��
4W�^<s"O�h���]0*%�Fɓ;yrhc7"OP��b@=|:��EÀ9^^q�G"O�9�ӌP�NZ�Ч]�Fd4��"O^�9fk��Rg�	�O�BE.��"O���q�� �0FN�
`�
@"Of��$bA�:����ϲc$\��"O�IP��oKn�SpBƕNhFL �"OZ�2E���^B�HB�܀?f�9��"O�T�sdL�0[�M�� �7)~�rd"O>�"UCA)`�T����XYC�"O�i3�(�A�ƥ���.�i�"O.��hZ?����6K�di�"O&�+��#[z����4[��ܒ�'��i���L�@(D��cX*O�*��'��h��3ZQ�9z��
�EI
8:�'e��G��bH��ǗA��'A��(a�]�A?B	8�$�%��s�'�BȊ�+R�Y�Z	�WA�!���'r����h�5:0L9$���K����g��{�<�8��}z�9fBY5BL��	 O "T�	+;9��{��W^�p���	1�u:B�O�t���fб7��;)HzI�!A?�M��"O&�p��=nq� ��9ruQS�'�}�s�5z	�ɤO?ݙ� �<>xtMs6#�:��1!���J�<�d��>+��8�G�,D:�݈1��Cyb�%� ɸ�#�^X�����oJ;���>�d�C�;4�<��>�����4�@,Y�-���T�D=!Ɓ�u+B�	E�ؽr�{0>� !b ���)s9���O<� Ht���S�8K����$�n��q*��y�����G���YۯO2��L��ioP8���.���9�;O��r
$�)�'~�&�;�e�~q"���N�O�`��?�u�R�?A�`Ɠ�.�t`ZuL�������`ٝJ<��fD�G����J;��܇�Iue�P刣p��EI Q!���f�M�����/Ў9SBO�D�41GcE!���q'�f��%t�;>L���P!�;7��������y�|�6�����8@_�@�jI�g�Ч/��he`�A�d�HR���V�}�}�ش%���AU�.pݸm�Ǌ�N���&]5j��28�,X������c�+m�"��вU�<�3G�F |ƹ�r�I�'�F�'�̭��JɎ�r�S8�`\	�{r)�s8����)��5�|ڲF�a[|dr�N�C�dQO܇M�����_+t�2�B�p<S��#9���P�BB,�x8S(�,4=�!{�y�(��|:�k]�LE�E#�SMr�U��4F�#�fIu�j�cac_	f5xJe�0�����'ْujB�]��J����Q�Z�>P;-X�f��Hd�\�mܜ�����CTiD����ӎ.�F8�T@���!kKn���$�B�T��'@�qvJ���}f.?F:^�Bh/g��A�(Է���@�+h�I�,TI�֝�P|�)$N��`�:HK�
'�Q9fZ��?iG,B�p[1O$=(�$S�4�H���dȀ
�����~w����-Ά����O����q���~*`��Ó�\0�BM>yPӵ���@�1�A���O�!B$W��RW�_�CTt, �"��p���Ҏ�X�L�qo�$��n0k��XS%��m?9'�l��PJ���	)?bX+N�1w��r������v+��2`�q� �agPI���{�ԟq
%�J��=�f��
SC�У�j�����/R�t��'I3�NR2f�X
�D�Ah	��i�T̓D�h��'a4!�E�P~@��'yz�Q.n��M��)ː@�����'�P��Q9xxJG��2 �Tc��x�b��e-t��UɊ�j��l�N��W�6	Z�J�>�d��'�t�W	�bXy��锖SXB�j�r[�6�낧$kD4��&e�	��/p0����([
L캅AR�F*4��
c}�b�/�azb�Մp#
����\�Ɇ<c��o�ZL
3�@�ʔj�d�= �y*���)�!�[���od� �bd��[�B䉁F���`�b��1��cv`��JR�j�����'�O���휃B��� $jr>�ar�i���;n�N1S�m�%^��hc��������.N�0DT��\��t�=#�922kI�K�D�%�W��1��c3�7m��V��"��D"mQ�A8T��#?��
�J &�axҁ>����D8B 0s" ��h����Q*�~��=BVI�F�JF��O�w��!�0>y�%�&C�*��ǝ�&}B�y�/�k~RG�����HO$����`�D�M�S�Tz��`:�� n��Bn j�ԉ�`ɐ�-q���"O�Ȓ%�BHӥ�E��>}s��I�2�(pI��^�J���g���Ґ�?�Γ+�(�]5����v�W1�4ta�F�C�IE3�	8t��4 �!Q�o�^�{�����Q	�hψQ������<y���t��"<���Κ.A&=��!�z�h�2�SU�t6��NY$ёB����Q�goݠ\��R!���l��E��4a���T�EK��'��q�쇫q>�e�q"�3S��kJ��Ɇ�T'&=9��@w���r���s��ػ���F�*R""׿��^��y2Iڤf�E��Ƙ }�����K�O�LXd�J��?�\ؤm�@����w5���bj��55� ���O3[l�I	�'`�@���z ����v��QB.O D_.����Lx�{��̌������Gol�07F��0=a�囃w6T�'�Q�<��Őm�`�c�c ��A5)�d�<q�#Bq�Q;�D��7� )D�z̓[��+@�'�"�~��S�S�Xi�"�@R�PO�<���Y<2J��cg����2J=�D�'�x L����	�_�F��c$�$l_�#r��W@B�ɚq�΄Q";5\���m�!NP��\8e�అ�I?rA��;��#y�Č�% ����䁜�ƍ�N���A�TE������5�j!�`�)D���ĨqDM�@�Q�L$Y!Gd=�I�N�$"<�|�G�љti�u���K�Hd �N�q�<�t��͘EK��U7�1 �q�<٤mO	$HfE����+l�H��Hk�<Q&iV������u7�XG`�j�<aӤ�'��z�E��M9☘V#�d�<���� �*���mI�]fL��m�z�<	)��f�ƵTLߞL��h2�l�<��A��$���NB�p�\,��/Di�<�6d
V<���R"@�z~�m�j�}�<Yw�Z�)�t���w�6�S{�<I���9_B�q�Y�V@Ru�w�<�!�Ԏ7e�Ī�$���1�t�<�R˖+}L-Q�e�8c:5���q�<�k��{Ȥ�4$؋w�0�k`�C�<yф��T,��Đ�K��KRD�<	�C�;�ڕ� �H9I6����kZQ�<�%ҞQ1�dⒶW�m�x�<AW�њM>��@��m���x�u�<iWDD�B\r����`���q�Bo�<��bK��!hGB�q���@�<ѣ-�N>�Q��Z���i�bT�<���N��T[��TiY�iGZ�<q0�D�J4��g�H�p�\���
W�'�P1��%�R�x��v�#e�u�RK�@S�Ԅȓ0�Z��Se��0HLqЄ�u��
ӭĮ9]��=E���PoH� �=̐������-�?1��U���D�d
�8������'=^������~�&�$,Ʌ�qc�yc�΁� 2�B̾w^��P��5��O��>9�f�9+��$�zh(�+���^jl�S� "�!���1%!C 2Xl�6�F;o����T"$bU�Xk�H��ا��غ(�|a)��O�N:�Y��n`��{"��,� A�<OЀ	�� N�H�(�G? �`,��"O����K��!Z�F�I?2u�q��F�j2~��So0�'!��Hy���D�yfߣFVJ���ݔ��%��>/���/��i�p݂PMH�]ZJ�'��F��'~�e�[�jl2!3W��.=Hb��'�����(�����_�"=r���'�9��)@��0>�LF&8R���R?�bu��� p�<y冫8V6mYt�܁d}SRf�h�<��kù)�"�����e��M���[�<!d Ui\�!���G۪t%��l�<i�K	�+	l��T��OT��"i�<a�M�H�-(0���--&x�p�Xe�<� ��f�߫}�8��V)��"Ot�
�dC�e�a��6fGȕ9�"O�9��Ț �A�'ǜ�@�P�V"O�ZG�O�>�Ȭ;6��)�pa��"O ��V�i���a�
�Vu�(@"O��b��=7���)P�s8��"O�t[����T�Z�Yt�N4%�s�"O<]Q-O�5<�H��ǹJm@}[ "O����8'=�K��o��#�"O�3�K��� #�
�(��d��"O��eIG�Kf�apd)�4f.]i�"O����j�eV��ȓ8nKZe �"O�$p�h��hiBƃ�P.z�H�"O�Y9&��Bp|a+'"�A�"On\�d�ȦE���He�[�Cz��"O.i��Oi0N��I�5aP��0"O��P��jw���dB�k�q�"O�Ӏo�$$ ��1��i��"O6���E+��/Q��ܳ�"O܁��O�p?L����6u�(���"O�mBSE�[t����%-A����Q"O�l�PHͼ9���4n]�a��U�"O
A��3a0�E �l��x�"O<�+��ѡ- �ؚ�霒 &��:G"O2A�B@�|~M�
eA����"OL�K�d�.� ���@�*����"Op�b��X�-8�\��Ǉ�h�z "O��I�Y�"��gΓ%�h��"O��E��|�@Ӕ�o4r��0"O*�B]�	)�q�+�}H|sU"O�U����#ZJ<(�
��~����"Oi� �L�Y��
S�T�c�Fk�"O��$]�i����PG�KȤ��"OD�����4h�RdĿ{��"�"O4��C{��hGd�++G*����>D��S YC�}{g�@�nAL�ybm?D���&��;|N͋!e=6�d���8D�pkv"@X��@�<s�{f�1D��i�A�"p���q(�) �b-D��s�(?yp]ɣcK2]�Y:q�,D�d��'�{��(�\�
�`�D,D�<�=\�l�B�ژq��Ƌ?D�trN��<EY����l �T�=D�tPA��Q���jw�^+{�@Y��:D��Pd3���X\�"7F8D� ���!�*��o�"Φ�SrJ:D�|�pݳw��@Q�K��|&D�0�-D�<���.�$=@c�U�[$RERk D�x�CC:(PQ��.�yRp*$D���e�K�k��Ӏ�]{V�`r�%D�l�2�	'CBh�Z��ƖbD@�p�7D���AaEt^�(��ȝ"��P�:D��9�k�e���*f��* �����8D�d�d�@;qO:���c�c�􍱐.5D��!��35�F��$��v��n&D������v
�	�F�<%x�i��"D�(�?[���{��Yg�X@�$D���N]1v�X��+}��L�AL!D�4@�!N�%Kӌ�3��xz�>D�КC�<VĴ�ЗE 3T�����:D�8�%��TؠX��$ɨ5�J	#D�����ǃC���刮z�|��3D��a�KP�r���1�=J���6D�XȦ@�-]��	�ǖ�A��9�m4D�� ��0��+y�z�SNo�jM��"O��� e�W��a�D�M�l�T�Iw"O6HZsm�\hL�-�Cm�D"OP	Rv�X"���Q��@���"OT=�k�=�h�cRd>�A�I���鑪6z"hH�D�j���bK�+i!�$�m6�q���@���#3e!�D��B̤��^�i��H��	��xV!�D�
3�Y���-� 5Q��N9Z!�䑢B��{U���uƈ�1aN�'U�!�ć!L@���eBD�*��hQ��>5!�έ~6��Yp��9Y�6�&b�p�!�$R�q�I����^�jH�����!���-;���!��`d�b�6P�!�DL�^���C��j�H0 תI�!�$�n��]��g�2a.1D�K�!�d�._��Z��K8Z0QK�$_'L!�D�&x 2E�1�Th�3a��r�!��w4͉���5vZ�,Xw��.\�!�Dߍ!�h��b�ޔ�kw��!�D�&u-<���b;i6�H��&!���W%�1�@Gۢ���Z�/�:v�!�$�#ߚ��$ ��٨�.G��!���:�B��`N�e���e��DL!�d�wf���◡d��as�B�g�!��Ɣj����@�B��4� ���!�d�*Z&dXƎ�y�U�f��u!򄖾w���j�bwh���Ҧ^V!�X�j���3		%ut�Ɔп\�!�O !��|�I:{�l�t'ΐZ�!�D|P�q� �^#,P��C�
7>�!�dB�EΥˀj)�a&�Oz!�d )���XDC	^!ր#�$L�#a��yCa~����c��ź��"w�	ʱ�͎�0>a@�>}RF��ZH`-8VD�2� �A�B���y2M�0��!a�Z�X�����c���O��93�O��� �rقi8�J�I���'�b�+R$�&+��`%��7�*��g�u%�>�kF~�q玠MO�1���ξK�9��V
�My���<w% QX�#M�WI�I��?aw��~�N��`��$e�\C���V��X1�e�����'7j��S�^!�����P���xq
�'Ը<@�� l!�5DJ�^���{���*�c���b������*��гj\� r�G"O�����M�/�,kp��35a�w�'�&"}�'�Ĥ���Z;�t�4�Ѹ*.>�{�'������Q�6��5�����(ڐ��'
ʈXB��^�8	��;&0�L�'12 G�u�~���$f���'"Q0��U(s4Rx�A-�?#ࠑ
�'�d� D\
)¦y��eЃ���!�'����3�
ch|	�%`_:g����'�����Fߥhh�tZr&�� `�
�'��@儍TڀQ�a�+T��S
�'!��C%��5#�tH���J"��	�'&,zš��6^9h �0Z�1��'�*��FO$�����&
�P��Y�'�@�����I��5���?F��@�'� ؁�'�+ϺY��ĹC�.$�	�'��P$���,](=~�Z����yB�E�,ʜ;�E�-Fe���	�y���������J�	�z�Ysڞ�yrc?��0r4�|*d�y�&���y���y%"xX'/�?]�(�����y
� �Yx��uپ�ڄ�Ok��(kb"O��17fB�~��tȐ�ً4��M�s�'X���s_�Qr�ɑ=7~x�lցk,!�$%.���B�΀mu��`�X�B!!�T)H��r�L-I\�|:�<>!�D�3!Œ��Tխ[����sk�o�!�$�g�:q)Q%Z=;���	�-|�!���.,E8%g��������m !�8(�l�h�Hr�r�)D(U!�Đ<�p�Y �P8b���bJČ'C!�[�5K%kR`��9S�����&&A!��O8t���.�X��i�/H�!򄗉O5(e�$ �,WҔ9���Ft!�Dԯ5]�
�	?t:��1�啈po!�́(c0�(@�A3;�n���唁4�!�D�c�,}�d잸=�f��g��/�!�$�X�� H�"�O�T)�di�4�!�D!::4�Q�F 2�0�B�]%�!�DR�/�a�10+��}�N�!��v�t���X�V�%��� h!�D(E���ҵN�RxJ0¤�)W!�P�D�LI3Ĥ��M�9!�d�G�8��0��%IS����Ô&!�DX�ȼ��ǯaO���U�U�6	!�dGA+`��y��-c�m���!���%�v)��Һ\�~ Dm�3y�!�df�Х�8eҜh�,ޘ7t!򤍿P$bq���";3v��-+�!�:%e��e�߲W�l0BA�A�!��t���B�Q���pOݺw*y�'�p� ̑/m?`�Ѱ`�!X>a{
�'	9���Y?���<���I
�'^�l���Ͻ	��AqO�]��%B�'��H	G)��X��}x��D-Ӫ���'��"��R�i|��Q���p��Q1�'�J���K�7r���"�[�<���	�';���b��U�0 �wh�0�$c
�'UI:��@<� ����$R� �	�'{,!�����@���x7�ܠ#���J	�'��0A��1�6�����0����'e�A����-�0a�@�U��P��'�E�T
�	��,#�(�O�h�8�'n���$3�\U3W�<C|\!�'�P����Z���{G�:+����'�������;�x�{$h=8Z�pS�'����ǘ�^�����L'+^��'4�e��7ԾMH�O��%����'��|YΙ^L���O�
�4 �'�4RmD�)d�����j$P�'5�Xǜg?���g��V�p��'�X�r�J��<d�t�V�Q�f;�'�P�����.2<�!�#d�	D>,%{�'~$}B`�I�ؘ�ìF�'KPܠ��OzU�w	ıCV�!�eDM�I:�P�"O"�!S�*�*�Z�g�)�r"O*@�̈́5x������
%���"Oz��F=*������>����"O�1�C���Q;�<SU��i�H�"O�,�K��Q$>����#@�� �"O<�x�ŜZZH��wܭg�Ld�!"O1A�&iW������2I���"O��z�끅q����rMH�8��X��"Ol�R���.�Ruသ=�>0��"OzH��g!;Ѣف�!�8�T�Z"O�  "�'� s|}(S!E�DΘ�3"O6����-GJ�x ���H^�졂"O����4�� ��1����"O�e�Wn �_��թ�OeT��"O�xZ(�.;�Y���I [ҹ�D"OF1R%D�su��A�lK�#��2R"O)./t,� ���"T�@"O���,$)i<���$Y�k|��"Ou�P�f2>�S�fS:,r���"O�AP���P��P:�V�5���"Op�;B���N�����M�&J���9�"O�A��&9ʌh��N��6L�q�"Ox�@�c(^R�D�.�� Npb"O�0*�b�0��y���H"O�u�4CH�iS5�ީl���A�j�<	�"܆k��PBAC�4��@|�<�G
-"{R9;�ɛ�+�tC�c�n�<9T�֙�
	��%�Vc�
B�<Q \e�:	�@H!<�F��@+�|�<�BBS�|R����.۵mpȩ�2!�t�<q��\PB�)�лXX�i�O�p�<q�g��!H�!�S n~����o�<��n�2LA$xZ�d��=[P���j�<�j��A�AҊ;@伊�ĉj�<�@�E#?����C�hB�:A�OM�<	K^�uy��;�ܵba*�O�<���j�B)���Ǌg���]>FB�I�lx����Q�c�L<Xq(̨i�C�I�`�
�C
x�rE��K�W�C䉤a]t؉��Q�l�ni�0�NNa�B�I&
�B�E-[�<)�pj��#a�B�Ip� �R��#N6��t�J�[�jC�I�dEF��hA\���#�Ǡ=3rC䉟Xݮq0s�ԏb}�dp��C�ɋ&�l(8��1x���!5�ĉ��B�I�`XP�DOɫI���a�2%�B�#4�`|r�,�:I�=�bKqn!���OU�([���8D4�QA	)[P!��Ձ�Ri����v�ᢂ�'%�!��˵-��)H�*��2�X�0��"�!��--��ĨC� ��1k�ʔ{!�$V8^^ҽ���6O����2�)pu!�q����LG���P�Ɔfq!�$�<���b�N>k�~!��a�qQ!�$��q�����T���J��;%!�dϳ,��xT��=P�IQ�8!�!���,�ᇍB�dtD�"&N?�!�D�]�e#�b _(l�p$?v;!��[L|ٚs��`fVL�r��:!��]���l�
+wp�[ï���!��nl&�P6�hN^,x`�N!�Y#s$h��7�4nB������
-M!�=a"�R�V$���v�u���'L^$cb�8K&�,A��@�{` �i	�'BΔ�U�r��5�7�P�e:!�	�'��ȓ�
0j$��
�	��X���J	�'�Px��=E���[�LF�P�~���'�:E�V��v�^���nQ�EwFH�'_�t���R">��xz��D?��-[�'�X�U[.c��A�T͟�>b��Y�'$�`�Bd����i��ɗ0�<�K�'E��)���B�69Oy&I��'�}�`��S��:C�s����'�i�+l����eƞ_`���	��� �(����w���B��:����"Oơ�ʾhHx�'J�FF<(`"ORLB(�0�*%�!��0	,�@�"O̝!"�*s�`p�&(I���`�"O��2*�J$�*fPE w"O6� ��GQ�4�(�G~�PW"Oh�0a��!�^���/H7���"O�u��B��O���8<*y�"OBP2�=`Z�Aj&M>DڥH�"OhD!��H�Cc�`׬^�[=>x��"O֤��M{��P�K�8!7��k�"O2X*���D\i�1I��H%�E�2"O ܂g�;��P@��W9��F"O�Tjg.^�|I蕈W�1(�D`�"O��NLKچA��}"h�c�"Oҥ(��4�D���]�WyL�R�<��#�$N�.Ek�,� ��-y��XK�<���:x�TiԈü_��iq�[\�<�Rh��HS�f;IO�Ċ�B�^�<9'$Օ>�,��p�I�05��X�<y H�!�4(��C�}S���`��h�<�㗼\"��� !օH2����{�<q@o˪n�R9�B)�y���O�v�<ل�ٻA�<F���]Z3�t�<��E��j��p�7Fӭ, ,�񆢂f�<�.�!`=�-	cN�)I�!��(Mf�<��׊&�:!S�/�(H"�L[G��W�<9�Z�2&5Z��B# ��e�t�k�<��ǟ;�\�'��5q�$ WF\n�<�B��/=
]p��ګi�f	` �c�<���h�E� *;���4KS\�<�cȒPi��G��0~��q�%I�T�<��ϝI��[ Ö_s�#�N�<�➱<����%��V9۷H�K�<��DV�;�X����0&dP�l]�<q��.}I�T	6�H~� `G�NX�<G��.ݼ� `i��D^�e��hBP�<9�ՐiSnI
��gl�3pELa�<�Vn�!r�� �K�R�d�5�`�<�v��b�L�憕X�*��SR�<90�K\��"SgW#��0A#�y�<Ѣd O�pkpX�(�(�'T�l��b��Y�f��7�}���$D�@S�T�܄)�V�v�(��%#D���F̬,d{"�(?�`��m!D���	(��A��#�'�\ՙQb2D�X�����M��4q$E�M<D�8�RhǍD�	�N�J�"q�;D��s��ۊ6�@�@"O�#7)��	.D�L�dD�La��bk?b��iQ� D�h��&ٯ�H�Pm/ �;�/=D�q���-�@�Jj�h��u�.D��Ц_�+�ͩA�I�d`�ZP�'D�X�2�Ӿ0^,���'��u�*}²�9D�8:wE�_����F�Ř:<�|�TJ3D� �V�Е/>��*�D5(����A6D�@s2.�(>���5(6n?��k4D�d@��1\�ru������,(D�HI�JC b����w	�-rrm�'l(D���ǣٟ2�؝*B���L��\�5�)D�̩�
��qrvD"��:�<D�xE��+r@(��*�:}���o9D��q�Z(Uۦ��X���+�6D�ԡ��6X-8�jN��pDe�/D�� J����'BHi�D�" '"D�"OP%� ζ� �m!N�n����"O��`��K�;lAhb�
 B0�2"Ozyj��m�&���i�/�	��"ǑJ�1{� �JŇ	=S2n�Y"O���� �s"a����M�xX�5"OVH�aaS�M�ڰ��E���H��"O��!aA�"��SeM7aN@�E"O�\� ߩs���xg�ُDB6�C%"O�@�4fL�-���E��@(���g"O���S`;����F`�&��"Ot����E2�·*e ��"O:i���/⸐@V���w �}�f"Oz%)���]� A��f��I�7"O�[r�ރ}¦�`t+��c�&1�R"O�q%��%"V��*�,
*8Q�"O��j�G
 ��T	�3F� (`"Op4�Ǎ���&N3��=�"O0�2���M�u�V�V��<<�R"O 6��r>��e�.�6E2"O$2$�	/	��p��?�FEBg"O4���ʆ-�X���˼���*R"O�}'�9.�$tA��.)�2�����R�Or�X�#��H*Z<�Ul�dR���'�z�p���(3
���O\0e_�=��'���郯� t�Zi�D��uU���
�'��<�h�=6��4c��X�b)�-h
�'����U��;]~�P�+Υ*��a	�'ɒ�0î�Y�؁Q�>v��4��'�L(Q�R+g3>4�p韘n����'��e)R�9 c�=��T�ت�"�'xܤ�S�
�v�ce@���$��I��B �p��iB�I�a+>���|`�4`�J�?s �H�j�NU�ȓb�<�3��T#tA��J� �jh��oy�|ʟqO�M� (�,���#Tm�a "O`�A���Z�1!�E�ba*H(�"O�\���T�� ��1o��e����"O��s��)gk����ޤ\W><J�"O���f��\Ȓ5�L�W;�yj�"O�k�����i$�H8c@�A�"O�@�ЪHE:LB4斕*3�@��^�'��[�$��v���s  ��)&�|��'<UrTAߨ�H�!S. ����'�L
r�M�)����AAO��t��'��Qj!�W�n)���p�<-I�'!����N� ��t���jG�:	�'���6G�� ѢG��q	ߓ��'Q�, P�C�2�R�R5��s��!i���)�t��*�� ��K@"R�%XfJ��'�ў�O�%���'S�]z�䑻}¤�I>	�H0����N� �R}�DN�s���ȓZ�@���bJ�0>İ�&g�,�ȓ;��c�	��&��!k֡7WJ��ȓ4��pC�֨t;�rS�S\�RH��b���³���4Wv����LR���'�
����W g�����K	J�����'3Jx���*\��/%6l�b���c���0=�Ū_#�
��@�Z$�p7KFJ�<���������(=�|��bO�P�<�S钔R�A*� �:]����U�<QD,����@LG-oC��7�|�<�$	^�J4��c�(�Q���ӱ
uy"�i>�<	2��v>�1�"%�T"�[ {�<� �a;�H�����UhE�o٬�8�S�$F{���Ł��8:��_�T#\��m7V6!�{%xr���GX)���-�������:�Å�IyX��A��h�1��K�8|��c�D)裈�E� ȓ,^���%��7j�lA"�Čr����|pis�	ϓ;�j��S�Q�3�n5�ȓ`��U�AC�Q>��;�O��x�D��ȓ8��a�$�Z#^�p�`�E�I?x���A��z7k�=�8��<C�.h�ȓ��_0Q�%�0I�Ĥ��iZ�<ѧ�|��<cB��84��$�a�<1%�B�.y�8����24A��Dh�<Y���6t�>D����K�D��rC�`�<��Gܸ[\Aza�� O􈝪��	g�<�5���:���p���R�Ce�<9a�8\��B�kc�Mb`�_�<a5��@�vHӅI�zU�8���[�<�"����+������Ë�T�<�T`���4�6�\!.K�0�Ug�<i��7�h$��9i="��I`�<P�-J^����2��w�ǟ���@��(A�(�(%���V��kH:t�ȓx.�}��ʂl�v�h�&��yf؇ȓ��t�0�*�P� r��*���ȓa���FػGp���٣6�����	`~"���z�X�{0Eǡ�.��ӊJ
�y2����wN
�������Z��?y	�'F(��`�h$��@b�|��L�-O(�=E��Ł�C�\2�5r��Pp���y�X�M�r���+s�e�f�J(�ye
�|n���Xg�4	�̬�y�Szց�W��K	T!�����yBH^;>�G*�����R`Q�y?$sLH�'��
a�&�!J[ �y�C!e�<x(H�	/v\����yb�7U�.�`�ӧ�*(������yb߄$9�uʷǃ�`�5��yBC�L�F`���xn�����&�y¢�M�f�Ċ�z�:9����hO���i�.r�ڥy�J�9�i��có:��'3ў�>�	�I�=#8\cţ�jjr$�!+?D���P)P�%	���֮�+�n\(e"D��g��6=�;7n��-���k�$D��3�␨O��c���-r'*uK$.D�4�A)��9�r�xU�ׅ	�!�V:D�T@��K*?P��S	�D�
�kR�64����	vnͻOYeNx���HD�<)&.�쮡�&싚v`�X�C�<�&)V�~�: P�@�Tt5��@�@�<Q�ɼr��-��m�p�h�'�[c�<�u�p��Y{@։<I���u�`�<Y�GT�uSֹ��V��	���p�<	��Էz��}3�l _�ΈfCMo�<�4䄸hNz����&��v����x�m	�w�z��"�F!_>,�(�*L�r_��$�"~�5��'���%��#dN��g����y��> Y�}�ª?פE�gI
.�yrhV�F9���Ȋ4��|7E;�y���t���1v��+�
��F"��y�k_.c��HBܵz��I��H1�y⡍8'jz!�3�Ot��p�Ղ��y2FR"dҹq@��n��P払�y��?3�8�*ՠ�<{���0�����hOq�� �Q���ߛ	@,�c�;?+r���"O��:�*���`Ŭ"n  ʶ"O�a����:} N�0�W�Ph�"O�\q���#9���aj�G�:�"O�6 ��wܸD�Q�Y�.�Z)�6�'��X��΁ �`ʁ@��ؕ3S	0�OH�y�I� (3DNm�g#<=h4܅ȓ'kX��d B.�>dde��7����ȓ$2Yi"��b�B�҇�N6P�����F�lH��C���b�BKKfP�ȓbs@tё�	3o��U�Ǧȝ9BՄȓy�ɫb��1R��)�O�N���	J�'���a6��)l�� �ȿ+�`��	�<��D������b���@�S�!DF�<�$����@�� ӭRy6��PH�<��A�XE:y�a�-R��� G�<�&L�'h_d��碝1 Ǌ�1v#�F�<ɤh_4e��!�����I�Z~�<)P�Z�s�0�s��"~���-I��?���I*u�$�&N�_d�
��յS�b6O�\���JM��-�+G<#q"O�@*��=��%|P<�#�"O���K�nh6��怄1�x ��"Ov�*VMT�`�>\��e��7�̡Z�"O;V䋆f�J�0G%��њ�"O����7��d�E03�n��"Or�A�5��rB��K��:�"OҀBOT�5� L%	��`w"O<e���*(|� �F����f"O�XD��']�a���Y�|�~q2�"O��RŴJLX�'c �7�T3��o�<y��9 ��	Wd�v`�d��F�v�<Y�������P	�Vm����I�K�<��Dݗ�8i O�'��mF�^qx�hDx�� ���eh
� ����m�y�@�*[��ѕ�§B�X��-��yB匙`Li�	��:�8��p�ն�y�
�C���
�@N�=0ry�,I��yL� !!�bb ��,�<е��4�y2��z���#e�_�Y�&Jɒ��xBiC�O��,��F�(z@Q�h�%+�B��$Q���3�n�l�Y��;%h�}�<9�nא8Q��k�d۬pG�}�DE�b�<A5Nّ@�<�*0���a�fH���t�<Au�Y*YR�]���п'�}`Q�Z�<�hJY܊�a�8옽y��Z�<q� 64\���2"J���'��S����<���׬D:��@,�.2\XRQ��N����<�[�D�`�k"�P�C]�����E��0=�`�ژG�Dh��^�o�f��"A�<�����a� J�q]�{��C~�<y�=St�\�L�V�F����r�<Y�Iĥ%��Q�#־U��ѻf��S�<�U�C�J�
�z$�A7*x��C�B�M�<)�J�H�(%�aH�����F�<Y�>y���R4�K�o���W�[W�<a� E�a��0�D��?��u"��H^�<)g\�Y����刣�|��֥�u�<QDa�p7�Ḃ�� ��#�Z�<	t�J�F�^���#+��ԣQ �R�<9`aQ?$rԕ��"�!Y��#��O�<��.�0|1�2�$gMR�(ЀT�<q�W�_*�AC:py �0by���0=�!H�W}f\�ë��_�L��h�q�<� Li�cF&[j$y ��B�(q�"O��T)t�%���  �,y�w�|��)�� AW�1 +�Q���Ce[b��C�	:G��P"���m��U#�a_]��C�	�#�2�k��ѭ1��u�3�� ѲB�	;x�4A�bc�	��q'�]<C�Mj�Q(7cp�ZD�\�M;��D�,E$��h!��B�x���϶'�!��2'��$���&0�x �BOX�r��y��#6��tHm��*��c��ܖ%$�B�ɴ1��(37�>TR���ٓ�^B�	�K�9�C�íL�y�A$U�bB�ɯ"zЃ�l�m��9{�F����B�I�k����߷G�#R�]�h�B�	54����.'�~y��	��B�ID����Dj��ikN�뵯L k�d�?ш�	�^v�x���g� ){б<!�B?3V<��*Q�@��E�k!��Ȝ �.A�E��O-��84��=`!���;v�z�Ύ/�M�7dC?C^!��D�w���+P�`&4丵ҼI!� s����7HB�q& �D Ϩ9f!�R�c��qB�^��`�%.�
�!�$��w���#�ݨ]�
5�m�s�2�)�R�t��!�M��K� �X^q��'�\��@$�����`�>%m:���'�&���C�<��Ǚ�M�ؐ��'QA#�	?'�fTjP��BJ���'t���錳K��1'�ۓ�h��'��)B%�܊!�fL�!x�b�
�'��ѣY�	�M�d	@e��}*	�'�H z�I\%k'���.Z�V9�EH�'<�H�!R'XM��q@.�!C�|3���y��S�sK�ĨPBH�(Eޱ��� �yjJ<.���Z���('G��(�'ÿ�y��d�Z< 0�
i��8x�G���y�B	�o\$M"�e���f���y�	�+���aq�.!�"�S��y�(;:!�Q�0j&j��ia���y����Tq�+�*2r>U�Q��hO8��	�EY~|�� �;7aP�R'@Ɠ"�!���@5¡�3ǔ�bU���V�I�W�!��ٯ[�,PF��g�@����99�!�D��rE`�(�&�*%�4��� o���C��(�� #%�2v]^,��
���2�p>�ɵ�ٗj0ę���*!�B�10e-D��؁&�y�<0c��j&4m���*D����� ?�<��"�ea��[�a*�	[����`ԡx0��6
�"]>�؈f(D�� ���?BT�d�I2�B%C�)D�|��`%
����F�=���D�OV�=E�4DǛ4��E\*#�H��� `E!�d������1u��I���<!�$�b�h��e=��i��Фo&ў4��S`U� �$&�<[�j �C�2q�:B�I�b[�$���Blp0q��Z��C�I	4I�L���^2-�D�M�&]�C����)��ŗ����)E��XC䉲(n1��&P``��oͰ7�V��$&?E�Ϟ3^"MP��.-5jt!�U}�<)5HN�V��i�.C�?}H�8S�v��`Γ5�����@���k4�\����� Bakp
�"Ϊ�{ B��(.*h�ȓT��QW�@�~�|�W�V�3h8���S�? �k����<���rbAH+�#"O&Xp'L�Uh��b� b�j	�"O"딠S 1���g��@\B�"O&��Q��pFn��c@SDA@t"O�<�6EC�c�ε+AAŲk@��7"O���ϗ"T\h�SI�^,ء�"O��jq*7Eܜzu�<Y&�� 0"Ol��ڲ8��Ѣ� |:�k1"O�U���@#v�q2��#[�a��|��)��q�:�JV6 2������x,B��(�x 
񏍍*��s A�w�XB�	x�1t'Y�u"��ӫ�6f^C�I�DN�ٲF" x�QU��IJZC�I���������Q��%H�zB�	3_�l$ȱ�[��0�Ɓ��B�������� ܤu:T�A�m���O���D�7���+�k���R���-��(�!��%V����W�'枵�-�-e��yRቸA�n���ō�v�P�E[/&�rB�"z��PTN�|�����mӚV(lB�ml��H���1a�l����).�dB�	�J(���G�0�JHB�&�,\�B䉍Ggf���CJ.@4L�"q�~�^B�	,��Y`�gT�'�"L�Rf^�A�,B�	�R[�qQ���#�4�GH��C�	�r�r=��	JU��R��{C��]2�I
�@�yg>EyW���O'�B䉖R��铁Ƒ8(��.ɶb�C�I�Jא���䜭`��7�K���C䉀g�6��3�%V!�j4��r��C�	7W��(��*SL��8��G�*i�C�	�C�td�3 ZQFM�u�F��jC�	�i��HP��ø�2	����<�B��"f �*�bՌ0�@dR�d!4�C�I�+��U�w����!��2l�C�I�d�𩛕D
2��i7!A�G�pC�	3&`a9�فQj$��ɂ.|PC�Ɇr/���Nܛ/t��H�MկtC�	+dWj���v��b�jҲs�B��n��3f��_d`}�EcR�b|C��;J:yY D4B:��e��-&B��56������,�Y�&J�hPB䉕 �`Q�q)B(��ѡMȫ`(�lD{J?���퇜"�(T�U���Uh|X��-D������M����*�U ��c�(D�H� ��Y�fq�PƘ�1p��yI,D���
zҼ�3���6��}�we�O
B���2���0�1K�&�Sd��IE B�I" |����3Y.\�En� �$C�	�_R��J�#]���"�@��`dC�I�n�.}���1�x�B ��K��B�	I�$ʳ��7B(y;P���*m"C�ɔufj�0�f5D�ؘ�&�̐.*�B�	�[�H�܈1�s割ۅ>D��;�-���j�����N]@�/D��"$^�+|�[ѫ��X�(�:.D��Y��G�VL�E�*F �0�h9D���s�Ϊm<��#�cDM�����)<Ob"<���S�lQ9�H-�b��	D�<	��;U<��Q)�xY
��5��A�'ia��
�-#���dܥ~#*9
uj��ybI٣G�����Q�oP>i2C�] �y�@C�R���}�~����4�y�c=p@��ꊧo(V(wN����'�ў�π �HY3;!���O�'(���E"O:d9!
�?��t��oŐ��6"OF`�0+�g|
IȲOݳj��1��'�xR2�7,v��y�+\�b�&i�cn+D��9�*Z�Z�<�k�iO(�Dq(�`>D����&�M�t<���?Ujbx��1D��+���;��qÒ%Ձ(����+1D��#�D�l�he����?q��P2D�Dp@I�Zs���"�iPļ#�@/D�,���]$G9>���ގ���*�O2D����%p��D�E��4��1�ҁ*D�0!��hOn5�#�S<��P(D����T�g�f�A��]-<��!3D�h�e'I�2���j���*�B�;"a>D�����L���H��	1�4��b�=D������$u��Iqˋ"1.%�3b D�8@­�f�P�`.K/%���?D���jƈGr�\�+Ɨ2
�LJ��<D���a �	�9��*_w`���5H<D��Z��ZPH�'�j@:�6D���P��
K���õh� (B4z�h4D��cQ�^�<R���8`j �"2D�� �ȗ8#���B�o�f� &O5D���@[:�D����3:D�9�4D����-��,��ˋ]�p�A� ?D���R�vNEs&�>	�`��p�;D�T)5 �4j]���Չ �y���9D�d���I��:A�+kr����=D��Q �l�Р��vIμ�Q�]�<�4�Nbf��8���\�`,dUo�<iS��R�>�W�X8#�ڜ�&�ZQx�\�'0`KPރ���wl��v��
�'{r(�3l��;�Ĩ7�gg�y��'F�e�"�_/ƌX0)I.o]�:�'M�����=�B()(5iO����'�r�[�@��{���:7Y}��h�'vⳠӦ9���GV�}@�8�'�����D��$�UHڒr@ƀC��$+��4�0��fqr-`rʀ'KҾ\�c"O��K����K���(P���0"O4�j"�ˉK�����f��^����@"O�R7�,�,�PC[�<�~� 3"O2�(�)ǒ�� ���3~D��"O��Ǌ���l !�	glmA�"O�U���4��(q�  ;5=z�� "O	��8 R�ȰwBR+22i��"O��8��Νߢ�ص��0�h��"OJ	`�6U���FM�l���3�"OV��fM �~,��hY�J;ޜ��"O  #�jA�Nh��kbm�����"O:��wH{�v8H���5�B�"O-�UlQ�@�Dȫ�.�G�按�"O�	��Q��T�V�j�R9�"O*1=��h�W.�c���"O���^Yb�P9s��0'n=�u�@R�<�Q� $��蠁N"J����V�<1�(E�U�
�"���8f˴-�q
MO�<��j��eg�]cӬ����L� �G�<�i�u���C'� &�H�����F�<y�T�`4h)3M��h�B�
��Pm�<��@�<L�`��i
H8l9��iP�<)�'�,z�^��AÇ _�\Tp�WK�<�G�L �q�.��4R ���bG�<qT�5^���@�n	�~(X�a������S�? p��0gU"f2�y{��^�%X�'"O���#4	�ȋ�Ϝ]��]�c"Ox��ݍe�R̡t���0�W"OJ`����7S�$Ȩ!oɝX��)"O���O�)r�N���m�y޴���ybf����ѶBLnٜ�81�P;���:�S�O���8b�	*TF�re����4q��'�Ҽ�Ae�0^ࠓ�@p��#�'���s�ȎG�H�s�+a��'�Nta��%��m r���z�'�\����]��(�� P�Y�.y3�'�aiV��7�̹!�G^"Q^���'������-Z��б�Ð?P�Z03�'�1S��Z�3�t+7��JW\Q��'�lx����D�!���V�*�֡��'�r,9��� �E��ꚹ*Nx0��'� 0�g���Z��!���L�V|��	�',D"���]^z��g�B�Qn�P��'��49�f�"H �')��DXFx{�'e�p�W���4���/�-\*J�'$�1V���԰\P�(��ɛ�'/V����,�@���
��n=	�'���{ �܆�R �MG�e��'w�E�\B4 }�0₞8��A��'�8��l�`��!iPjO@E�@(�'2��5�.*)f}�t��<a*6�R�'.ΠbS�n��Фm�]�|���'��"�,��r�x���������2�⤀1�E�UKJ�ȵ瑖Z �S�"O��!�bS���tjQ�\-�x�
S"O�А�M��b�2q�v���h(��9�"Od\�7�QH<x\k��Y	D�b(�F"O~�[��B���)��	�"O��Zf ���T���%L���"O8LcFD�; ���tm��#dC��|�^�x��S��0�R�I�(�|����>����0?��MQ�O��Dp��˕="$1��'x�<�CE�@h�h����s�[�<Y$G^�[�i�լ��U\B��D��W�<���7C�� ��,~�������R�<iE癌Fߠ�H#��d�-�f�R�	[y�O��� c�i�� HԨ{��	I>y�d�2�!��Q���Yp%��'>8�'�a~�FޖN�&l)G![�1lJ��U��hO����#@�9�	L�qL~	���p!�䚛?��j$A,� ���!�D��OA�� ɦ}�s�JK�!��=.��,�"9 6�3F�ىZ�!�L����ҳK�Ѵm��]��'�a|���M�T��a��!\q�kB��y�&O�@$���\���AS�ɠ�y�GԤ
Q���jعQ�:e���C��y�S! wT$������҂�%�y�h� Y�ō[d��ъBhъ�y�EC-�R�0�ǈ�Z�~R���y�(�6�z<k�N��<�$ړ�y��T���3JL����5%�;�yr H��j�@��P�
��ˤ/��y�O��*4�r��t�"���-�yB��u��i��޵s��K�Iɐ�y��͠���J�c��^��<��͑��y�M��y;��HP*�(";v؀��� �y��*5|�)(�
Lw
�R��T�y�c�:B���j�(>b�eӤEJ��䓘0>� �TJvh�&l���	m������'�ў"~:��J�PЦD�5F7	\V�`�Ҹ�y��7`&�M�f�5�`*�aW�y�'�&L��F�+~���!����y"���B�|y�ЄL�(�R��	��yb� �.pR���l;Vd�ӂ���y₅� (���dK!T�
`�"F���?ɉB�S Gw\�Ё��k)T�2�fRL[� ��I\�'	9R�IɌt��*e�'!����'#Bm�4+�<��/�r.�Q��<D�h��@�&+��x��ծk�ؽۑ�8D�tk�*A��26⒠n,��JՃ�<����&s&np���ȳU>"uIs�
/Z��`���(J�ʃjR�p��0!�-�v��C�	�B�.�ӱ'�4��Xq%l�nC�Ɋ$�؉p���6o�@�E�A��<C�	?���x�h�%�^��VDA�y�C�	a���h��c�B�ZT��uBC�ɺK�(��bA�#u�,�zRm�!�HB� Qh��N@!E^�,K��1�B䉥e�~���‖qKM
g
�"8*���c���c��d��8I2C�G�8	�!�+D���V+��)D]� `�[_
�Zb�7D��rr��G9:J�
:zДI�(D�d��k�?&i���ɧv��HK��0D��I���D/ڕ�)�Nu��Ȁ�:D�@�V1)đrE�.��%)�7D�(B$Z5����F�M�#X�Y9�h D�Ti�]�<t��㏂u$�Ur#'+D����ė�m���
wJ��d�X�SW�*D�<����2L$� ��*�4Dy&��eG3D�h�ANE�ب�%o��U0,�O/D�LIT`�A����̣j"̙p�:D��a�eV;�v�����ʁ��5D�����К޵��O�.HP�xa�4D�lZ�bU���HQFg�%8N�s��2��,��_�O�N���K�� r,��$�!F�Q���xB��4��
�B�(XԊ8�y����qʀ���l�2M/p�C3���y⁏�y"�9��,Xy��gU��y�*��)w$��7A�5S1nY#T�Ǎ�y�ϼn���b�En`��O���>9�O��
�l�A�\�8�i�S�9��'I�	7'wb�s�ȗe�΀�&�T�.�BB�	֠Y{�J	w�~ ���Ra�C�)xz�]b�%[�d��5T��C�I�7H��LÄg����.ѱ#�B�Ɏ!;b�j�B	Q�����@?@��C�I�g�aJv�?��$�UN><OP"<YF�X�fM�$(Y0G����Mv�<)b@���9�,�!<R��S��q�<��#$��3�����`�HKR�<�-�r�B4��J=�[E�R�<��ǐh�I�`�0M�R4
qAZX�<!T���1����M���E1��U�<	C�I�ZL&q���+p��Q��om�<�� �}o��f�1m^��k��g�<9�"�.D�� KƬ
!C��cGK�`�<���Ɛ@J� u� !c���G�Z�<1�3^\pa���&2���m�V�<s���^��A�ºxB4S�NS�<�� �?mzM�"n�j7�끃WY�<ygϊ�����ȥ}�k�S���&�d�Ca4r���K�
7t4c��Q�'6a�� .U�BK�>�+�Pb��`"O��E�6�r!�!�V�2�(7"O^��R$F�eӤ9j�ы[�Ԅs"O��� �"F1�`��:u���"OP�J�ŉ9$��1ؓ�ӱWqNP�C"O���e��<7�S-K%O2p���'wў"~�B�G 2�|I���R�L�Ӓ��%�y�F�%>�l��#ν~	�h]�yRb�*!��	�D��i��Ѡ�����y�'R�z�⤈�J��0�0�Cj���y��8;4��"��N-*�.��L�y���@�nC�5�%aAi���=��y�t.Zpp�D� Wl����J��yB�æMCaY|ƶ�9��>��>��Oĕ"3�
�g&<�en�[�i��"Op$0����l�r@�`(��|��`"O�	�0�� _J��7Ȁ�p E��"O0�!@͟���J �E?_����0"O�d"�A�-l"Y�Q�;���G>m�c�)[�JX{ā!{V�A�.D���C�3Z��˳m�$�~�W�(D�P)��\)���6�T�|UQ	)D�,kq���܉˕aY�pb�b+D��
2E�K��3��K�l��B�4D�T��-�0�1�J�:izf�Ԁ4D��Z#ɟ%C��3��$��pWO1�$ �Sܧ	�:�J!IX�ൡ��0r�`�'9a~�N h+� KvnՏ��as����y�!�'5Ը�0��~9if��y���8>dd�M��i�0�e$���y�+F�X>5"�CH�:�J�����y�,�w��$a�ċ-�`8��ɣ�yR���i�v����R��'��y2 ';h6(�F�S�(�=Ca�� ���0>łި;"0]�PhE��dY���
|�<0�	x�0��fnW&oS�g* P�<�$e�2�� �5�._��UW�@W�<0j�U��J���J�������x�<���A�l��� <TOp�b.^v�<�t�L�y����<�~�y�k�Fyb�'���	üX/r�A M�4t�I	�& $
�'�O��Ot�	�lu˃#��V=晊�)���C�I�-9�Ӳ�ئ.r���,ði�C�	����Pe#Rh�t�L�aK|C�l�!�=t0�0�ܹmcpC�I�OK���E��J��ڃYB�ɀ{u��� �^?)Υ��b}B䉄t ��wi�i�Ҩ�Jݫ^[B�	5av�@�o��12�(C�6�C��FA�҄���p2,��Z�DB�I3YMvhR�)]������(m3B�	Cy�c1.@!D�y�`�F9b��B��W�rL
B��io~�r'e2�B䉷Xn�H#k��y�"�� (QtB�
�T�v�( ȍR���\B䉈S.��l�#	�^)��DԲɖB�ɷx�`G(�/,�D��S� 67pB��V�P���b}&�� �Η=fB�+$$��c�ߊVބ�d��2=�C�	)�ʽ�Pb͔Jly�C��\UbC�I(i0�CT��"/�4��[z�4C䉽$�xmbK�`�,!�.�1;<�B䉂w�1j�lI&�d�EGVq�B�	�E6����w��#q�ҿ��C�)� fq*c�)��CB�Vmx�0Q�"O�S���I��(��G-p�Q�"O�����,�X���;��Q��"O����M�/16��E�fi�F"O�P9�J�/쐔!�$K$dӒ)�%"OHi�f�
*ܲ�
QI��W��r�"O���F�� H}Z���8a�@}��"OnmP���g}�p� ;k��`�"O4����^����I�)wȄF"O���ġ��S��M�2��jcNyBd"O�%(�<b�0̛���9T[��W"O����
X�Š9
[�i�r"Op��CJ��bݬ *��Ft�x�@6"Ot�1k�n��!��f��j��̐�*O��hr�W��Di@̓���Z�'m2�Q�lP(&���'�,@��'sb�:K�42,I醊S�Gh�Z
�'a���GH-���I@��PR�<Y�+�}�V(�'� (hs
hK�<�($cX��nֈV(aG��\�<i�D�/4�I&*�6[��`sa�U�<Q  �|��E[1��T�dDZ2�YJ�<��T��&����ؽ^�t�!���l�<1��L	YUE{�朿6�� �6�^j�<�hH������< �v��+�b�<��/�"#�M̡f7�%���H�<	U�9%�28�FA��64�uc�F�<��aZO���3��[':Z���@�<!G͓F��d����3O���b�<�S�޶�&h�3bΆzG��Q��]�<a�H;`�r!���MuFI��X�<�4��W�r�z�D��a����Z�<�.ݫK; ��6�_H���LU�<����2&)�"��W�4`�x�p��Y�<�4o�
���e� �D��z%EWX�<1 �-�)����U���j���Q�<�b�M�"�q��ǎ)��U����P�<Y�J�B�,_0�4١�,YO�<�U��7e�F� FZ+SWX����a�<i�J���Zx&a+/tL�3(�\�<I`C�=
� �Q%?r��X��CD�<� ?z��@�{N&a �%j�<Q�6�J�٧!W1�̭���CA�<���p��(H���aKXW�<ir�V�*��M�D��sǞm�R��g�<13O�$h0 i)� ~�h����~�<)��M�v�+�o]*K*�bˑu�<��N�3zgL��w�]x�"�M�<�ĂؔtT���	�8[�i����<9pk�z��]��*��q_�)#O�d�<�W	�#x�TCc�Ѥ6:�Óe�<���� s���S�Ɲy�,A��j�<���� ]��A�" ��%a奅B�<���ղu��q(� ��4�ʶ/�R�<y�/žH{��bc��"+�%j��N�<Y���S�Xmi�A�o+���MTI�<�4�B>DF�r��p�H���Ϛn�<�c�FS���"�I6���d�Nn�<��aسL�-kc%`h����[@�<a��Zވ<����~����V�<��oЦ0�,�(��c2�	���Q�<i�� (6,P����m��y�#Q�<`�خ=`X �"A7��1���N�<Q����g���ʎ�-�p��#�q�<� �]�e���\�R��D��A�"O���f��}`0eÀ,@9�8C�"O������1���a��+eJv�R�"O<�83�:5���b�f<dt��"O��%��1� ���ʃ�`2����"Oba�aک\M��8p��5Qk�"O��h���1G"l�"b�ٶ,,�	�"O����\P�Q�q���H�z��p"OX�`b옌& ݃�o��"�:i	w"O"(U�l�t�DΓ����"O�}��J��,�*.�����"O�4��Iܡf̾H"ƛ�r�(y�"O�P�p�aH>@��4Y��B"Oj��&�9U�l��tÉ|TD���"O>����DL�ᨠ�ͼ>���"b"O�$��qY:ke���9B:mr�$D���/P�W����ŘsJzf� D�<��a���L�0o�=�ʙJ�*=D����J���8����6!���fJ<D�pBcA���I�#�z�biJ0�:D���'�!*�4�ps�ߊ_��Xר>D����H�)8k6�0h �ݘ��DF D� ��
�*����$+ -d�n���(D����ʛN�b�!PE��#�D9@�#1D��G��>����0O��gP!�Ѯ9D�����VO.Ȉ��B�u4Q[E�9D����?t���f)Ń�&�� &5D����J�8�u�Ae�*U�ӥ/D����`�OI�]�T�0Ѭլ y!���@� 5���$�r 0L�%u!�%!]0P�1k��� a�	�x�!���;[��`҇��t��@`&F�+�!�$˹)�h�Ib��3��y���r!��vXJ���0{h����%RL!���|�j4K���UG0�0cMҞlM!���50D�H��-T(N\A�.Fh!�$J�a��0�b�f����7L]!��-M
�E�� j�jK�GX!�Z4{4���$�� ��mb�ʌ>:B!��5 � 	��T/�DX`�ʉ''!�$B;( A�w�G�T1�ATf<!���%Y<�d;�R�U�\�!B�"!���5OyB�CW��.l��χe!�ƭr?v��F�\1ބ�	Џ��`z!��W�t-�AE�Ϝd9��]�8g!��j� ���ױ�esE���I�!���]d� �E>i�����	�h!��%\� �
(�$����Z:!�]�d�q��]�@�T,�!���'�xE���=j�RY��摬_t!�D,C������z�P(B$�0�!�� �f�Ӑ3�(iz�c��!�D�a��}�d�
(��,�@��)�!�$X'a��)x��
����~�!��8Ke.��Aٜ:��#0/`Q!�䃐w��ze�Ä�2}���J*D�!���,�(�󀩛�@��b
A "�!�M0H��B�,<�6��t٠)Y!��QЬ�{�&ƥ�̱�U��0!�-8���a�!�.d�����@5A�!�$N�#/�`!� �8Y.yk��/h�!�"w=���@Q'	Y�(c/#:�!��ލ{uR9�\1T<�` �́9qw!���E�85!"/�HӐ���Py
� $��5��"�p�Ć��aCR"OzX��ǉh����U�S�Ő�"OH���k���ܣ���+,��aS"O�틑�m��	��-@#n
Q��"O����K3�4yT�%'~ޕ�"O�@�҂�~�r�)�K�.x��3r"O|My�EN6*x�7d�c�����(D�x�T�AD(Ek3N�@7ԍ���%D�<�cF<V*]��a��!>��;�!D���P;NJ�9��d���3D����N6P�
�0���wID��<9����+i�9p�P�?E���G�"B�I���Q�F�A~v�cSO��2C�	�Z+ ��Qy�@	R�D &)^B�I V�HZ# Y��H\�C�\=����U����O�����82�<)G���Vپ�	�"O\�#�e��0�M!���i���=��A�{�}`�F*pHvnJ�<����;Ȉ�4��Q�9����Z�<Q�#E)_K2H�h�B��;q�X�<��ES��Ur�����rv�EW�<F�V�?8Bdّ�CG�P��"S|y��'��u�6D�>�8��N�E� mڋ��+��U3�j��T��1�t� K"�ȓ:�
�+֌;�z��G@�;���'I�'�)�'-�APUo�<'��\"�-<����B�\l�w����f�q�m~��ȓZ�<ѕ��?I�䕱7`�j��\��DA���$̗���e�lN��'<�I�<�}J~raj�'�,�F�R�mҔM�lX�̧O��bLJl<勦cS�.�ͳ"O����l �J�N��VB
2~��5�W�	y�O~�9�FK��
�dQ a�Ή[@R���'�t�����s6���W���"����'�����ς<;6 �Îʕ�9�'ƴ!��շ׼܉�.Y*���'Ԑrr,�Q#�}Zv���~��m`�':b�g ��\bf��rGu]��P���dX��j6��
<�L8���sp!�r�;D� +�I<9�胡�+Up�ؑJ9D�(�m��Y�F�S�̟%i]����6��0|Zů�?t��XS���	Q��)e�X�<�� �`���X�$�Zy�	S?�'qO�#=��7L���B���<e	8��Q��V�<)�c�6M���ȴC;Tw��f�j~l,�O4�� �\�F�&�b2����'�铇�$[�ax��T��p1I�}g!�����jcOP<�v��a�$xKQ��F�4�@������O&K�L�yN��ybo@��
��6f���퉼�y��w����r�PoEL�����$:"!�$�J�8)p���x�c(Dl!�$�f��aC@܉1��sj!�b��X���e0iJb��7Z!�I~5(XתZ3
�"�C���'�!���Qb.Q���X�
���+1�!򄎗<�p1Ɓ�@���(��Ԋ*���m��H��ԑ��<<.��U녣}��۴"OfmH��^�Dh�Ǉ[*q�������%lO���e�9�/G6J���b��Px��itAc3����`�'�:GN �q
�'�(�Y��Kav�P�n�:��A��'h��ّ�ݏoX 5��ۏ�Y�˓�(O>�I��̀cFfٸ�`L.-��S���	N8�� ���p���,J�ݣ����:�0��2OV�	J�S�O&ƹz��ʰT��i9�J�lK�|�	�'�D�ƢS�,������,v80�)Oh�	�Q�b>ɚdDڧ~^
8��t��E;Eg#�O�U��'�$b��^R��<�sDƶL�F=��AyR�'� d9"χ� ����J����i�����O��PŇ]H=���R�H���'���bWa��L�ze`�D���A)�%�(O?�D�5i��e �d�u5H�DC��!�ā�TK\k��4~�X���[���":O�� #�S�(ڭ����2i��9�"O���AL<m�nI�'�O�8܈,)�D�OR�|�g?!Vm�y�½�D+�`ɖ���̈?�y���% !K��6#uصeO���<�J>�����UC)"Sl��p$^M�^B��$x�ƙ�e[<^���SR��)Z�.6�x�'��1�D��*Pl�m#��ř&T0�!	Ǔ�䓸��&?"L��'U'0�Dy4Þ�r!�䉦c��5�$ʕ":$��aA��; ������(���e�2o0:��� A-�C�I5h<U�ͦa���PujJ
wvB��%I�a��`�._�8�Ư�$`.B�ɻRV�L�)$D�����ʉj&��p?q���,:�`��E�B�x� �b�C��0�'ۜ��bk�@���2�U�8�Q	�'G��ҳF��Os|J��R bN0i��/�S���܈b��2AνI0�ŀ@���'�ў��)�D"T&~��<#f�2Xp��;O!Gz퉉k�pKщ>�u81�ߐa��#=��l�p�e�ۙI�����]�l`��������r�O�H��!dDA�Zjn}E|���
@�.5ɆmS 5H*5���&3��B��!]���-O<D
��#��DʂB��7S�5��g����jS.z�,C䉪�聀wH�J�V�e�8%���p?�T��(��iJ`�,9B�9%GWX�<D�M�|�ӄl�њ��.�\�<�'�۲-�6a����`�
my0c�<��t׶�BJ?F�P!��SaX����t?���M�#s��H�F�J����V�<�T�A�u���Ĩ�/vZ��F�Ii�<Qf�0�&�y�g^� jF�� 	d�<�⟫kQ|I����_�2x���k�<�$��#>���V���"l��U$�f�<�v�QIt ɱ� �$]�r�Dd�'ў�'b,\�r�A��R�� [%�����#�V,����J�b�;�M9^�8���ܭ�&�W,q�j��� &5"$��I_�V�on��I��Ѕt-����s`���<A�i�!3��0;ۮX��1r�ȓe�P���m3R�#C��kJ�=�����# �&&3�|4$ׇi �Ey2�'Բ0��l�,�rXa�W�}K	�'ANAɔǅ�|�jLIVo��N�q�'�ZQ�w�J14E�`;G���5[�'yb)��F�#�$��CG��xc"O���DL��B�����X�.��Z �'=�����S�:S/F�R� ]���&D��X2���&~8)��Q�M��%D��ѵ�YCհ���N'0��!Ն#4�H�E�
3.gj��D�10�s5�˦U�'���D/�����O�8Q��eC�V.�����v�^Ј���'dq�"� �F��T@�:j�D@�J>�V@.lO�8S�	�!�`( ��|���0e�$ �S�3� ��Qgj��/��<B%�ڹy��+"Ol�䡈�U	6��f��|�p���	p�'��I]��9	��\�L�:�ʏC�FB�I�0�(�2n��s��y� L�@knB��p�(8�q&�|������˅S�>B�	}x�����E"�FK�2.E8B䉴)�@IP��]��
���'"��"<���5�S��N7��l��C�7ھBa"և�y�
�-+ܽ��G�!'M2`���y�)�'�&@U��2͌��HҨ݄���`�aƩ{����T�L�S��y�c4����?���Q�GQA�,����9@ a~�^�YBCWc����V�KrF���:D���˂�Y\�8�-	9 :��S 9��V���'Z�ٳ��>h����	@���.lp�����4l�N�8 %	�Z��ȓ0��Aq2���N
vL���C�����{�谅�8촘��
n}�E��Z�r���THF̺l�
S��m��}���dJ�7I$v�*�h�S��܆�T���Qf&��*|��as&QO8�ȓ?� 0j6���W��i����.�f��>��	jr"_a��� �9�Rņ�nQ@��#�E���T�f�	Ȇ0�ȓ?{|yqe��5��D�#�g��	��VE~�!C(�\Fqr��U�]�����z���� ��zz@1�e �#@��ȓk�u#7��_AB��@�����(.y`'5{���� � GL��N3�A�p��' /u� ��RP��CBD��Sឌ] (�ȰCF6x�>e�ȓ^*(a�/�	T����,y�H�ȓ_����τFblM"�H�����ȓJ�0��w�ܚd]l��7�\)_ȁ����:q�
�8H�홧���[��ع�'���@�q���扆(Ԙ-Q
�'��ȩЇ�>`<��n�49��'d��J��lA�`N�\\@�'�0�B�CC�bZ��b��!]��'�� �^W�4��Gω%]H�Q�'�����ڥ�8�,Z�ߺ��
�'�p�)��\e� H�\�1���	�'N:9�@��-!H��{7�ĬЊ1�	�'�$�[�N*�~�2�(�{z��"	�'̀ɨ���=H��ݢ$N�!�|�'s�X��M�	*���r�%�8����'�:!g�8����3"ݩg� 0(�M�1wɒ��	�)9,̡ӓk`ѣԪ�_$��)c�F1O�`��ȓG��y@ɞ37l`���D/mhb���bL��R�<�H؛䄓)c�Є�ȓ\���""�N�WAށw�,��$�Y�B� ]Z���%A�|��م�F�T���S7+�A0�\+.�����pJܜ�F�8&	@�䟧Og�]�ȓ��F�ϯ(ʴ�s�)N�^��K�����C+0� Y!�D��Q�ȓ}���b�oG�E�I#�[�5��n���``k%kP,�� �Q���8��O�n�ʳ�ղ)�ܵ��
9�b��ȓI�<iaЯ�B,��SgO6r�����8^R�����8� T�FZR@�� ���
�� 4���U	��I�l��g�츋G�Y.B1���f����Y�ȓ{��h��9?U@0j��;��<��S�? *y[��ę]���B�V�v���k�"O��C�_;bh�Y�s��m�(و�"O��u�W>[����Ўܵ�b�("O>�"�!Z�{n<9����\x��"O򀋱��7L��%D�:����!"O�Y�t����x��9p�H�"O�dk��R>y��\!�`��"O�M+�)����(�d�^� ���b"O�<�5�S��4��#�
N�:�"OB$Y#I��o���2^��f��U"O)��hӺE������HB�vؐ�"OV�cD�vo^���D�Z��͉T"O�|A�V&CM���f⃜[�Z�A"O�i`�I��v.h@���m�Ѕ��"Oޕ�4L55��0i�`[�Q��"OJk�"��dT���@��\����"O~��g�	#M�"��D��1�P"Oȳ���9|<qw��9(8lbQ"O�y�H$��Y���{�"O8���@�8hvz�y�/�VWh��"Oµ�B
�$H^�1�F

(�Yj'"Ox�4dD�Ҽ"�늖p�.7D���u��5dj��eϒ
enƸk�'��� ���#j��ݘ�*�\~����'-��c�W�!�`jdC�|!r�i�'��t��'�"}���q��u��'�~h��
�-"쨈¥�V�[J+�'������P�L[�4bE��@eX�'a�eۆ�?�z�#��y�ʘ�
�'Դ)�!`� Y�|q��3B=L�(
�'` �Z��ď,����:�(�
�'��9y&Ù&K��m,a�x�"O�1 �'��A:`��go�=wTpu3�"OƘ�!�1s�xhkΠGZ���"O������M���1�*��ji��!0"O��:�ۣU���S���P�$�"O����MА9 � VÖ�^�0mB�"O��$�I�R�R��V�~(��"O:l+�T�����G�W���qn<D����$Q�n�<��*.lUN��@6D��0AP0�d�W$T�	�@�5D��`1'�Αj�NX�U���a�g2D�t��	T��g�� �$3�LFY��H"�'GG���@��'�q�7�ٖPȓ\<v�We��~f����5	����#ǉpVP���!Vi���O��Y�O� h�VQ��Sú��v"Of���^xFTSs@,�X� "�'��͘W�U17cȪ���HX��a�)P�u3*�2��&{���b�6lOT��T���U[&��(��e@*�/I�v���{�f�#|5C� ���mN%if�R��2r3�1��5���c�Z5(�6:�0��1�}�'qu \���[1@-k��'%���K����ӿ>;�)2�b� Uvő	� 	U ݫ���#Q.�h @%�J�������4�y�/�#g �P�kQD񈇊���y�iݷ{��-H���[� ����/��u�7�^r�.��<r�����4n�N�cP%��'Z��&J[9 +�L8�+�o#d{
�I ��� ����R��bk��S,�$�ڍ�bE�i�m�f�=ĆexbM9-S��鉗 Y�E������q��^`hb���1+��Zi|TiRe��zX��hQ����0��Ƈ�#]�u��B�s��ң��S?����E#D�4ZD�J�<Tz �T'�?CB������A��t���M��d�IMa,:�i�6?Q~�'��Dλ
y�Q�p�՜UU���EnP$݄�R	����� �&�
-1�o� n� a ��I�o| �Z2��u��,؆�҆R
������ ��<1�n*�X4�G��f=ZKA�Z8��s��މ%��8լX>g���*ÕNx �㭄�)�� � s}<H9Ѥ� 8�^����=az틽�NPQ� �B,H��������#;�x����:u�M�7aV�.B�;�c�H}�-���� �!K6N�?-��mX�g�A���b"O�����1&b�M $ �uJQ�aB	*&�!�f�fF
�� g�$����"_0'c�d@�rDM�2�,bQ�X)/�DTB7�ذm�,�%�'�4"�O�/'xz�+���*��p3k�C
��:�g��!����@H�4��m)��iF�ܚ��DTZqO�%�IĞ)$ �vO�=��H�%���|*���<<v�p��͗�m�hT*GNM:5}&J`�
�%ndB�FI�p�Р����8K��&\O�d�5�J�,\�"�큈 ��q�gZ� XE�I5 .�Tcgi+!�l%��U����4s���z�ɗ F���@�)��V˛3+��X�ȓO��2Ch�=/�v)�搳ds�����[/0�8�Â�ע<d	+�KM�F�z_��3��en�Y0dL�BlvU�ˑ)n>-A�.�O�H �G3h��}�!Ϝ���%�U�� �:�&,]'���B��؃]&�i	�'��m�qo�- ��5$��r�2Rp!8� ��Ĉ� �7�;�Bu�� 6$*3V.@^�������I:��\�%��y�!ɡ���8-�*)t�����<�J9��k�$���r`�\q~�M0-��i�B�B.Fd��S�S	��S�"�p��pdӹ�Z]*kʱ!�je�O�hrE�LM�U��!�?R1�|qa��ߩp�����E�E$.xB"�OL͠Ӆ��|�0!��'�x]�手C�, b�Hi�<1��Y����F�`i��1�'�# 떉�pl@9Okz	�'|6-F�,O� w�E�^+tU��T	^Q����"O�Ѱ�Ō�A2�IS�P��Y�r��4���A�c�$=e�!���
ux�d!GbU-&�RmÇϒ���\���.\O���kC&;[b��3���W�0`� (K�V�j�%�{b�$�cO��Xuʐ�1���YF�{�*x����<~��*CF(P���9�铦fuj�PȖ�"I��6��YA!�D��1F�eID2\��hx��}= h{c�U�N4�U�O��Ӊ�Y�����0]��ܻ�ɓ6$����"D���V ]�UGhE�� Zw��1k��pׇX�N���IBa��P
 o�x��A#���!QR��4\O
-�@�Ȗ6��]i`����K�D,J���b�ya�A�"O��6��L��̀�M�Y �Ȇ��ǖB$�8$O�xV�>	р'C�woDu���+��0Hi>D�L$�˚Cbu�5!��n��+2&�%B���Y��V����D��~�D�/pF�w�4y���qv ���yB�I��yh��J�D�^h��GG�?�d�%~��b��%lO���	3���cd�c��E�2�'�d+���`�B�"d�Q�� t�5Y�o�&�yb�Ĺ{�E�V ���d�X��(O�=�E�D9����0:5H��r�*!��ɮT5�E��"O�=�C얮Z���B�ϙ&�L�"O���o���u��x��Q"O�LB�Q6�l�GL֫4br�	u"Ox\H�]�@Z���+	�'3�a�*O\=�ĨN���MIEf��u��#�';�D�F�7"���Ι�n	��3�[�Oh�j�ۺA����?����R���b�XD�"���>��P�������2I6t�P
��9��A��l	����A��X�
��<9�܀,�8@��3���#!@�e�'����ٱ@t´�'�����
g@5@�m��#q�(�nõL�T�ēqF�๲͕�"�ܔ�@"P�Xz��'D��2���D�v�9"��#r�D3$k�'S������p�jU16�(c�A�ȓ(/��b��^G��`i�,A)q x��2bܯ$*�$LM�6��r���J�4̉'sБ���Ц�Ql�H�t���qv޹�%1K,�q���s,�#OOC�!zCD�$M���@ 8�����JG�\�� }ѲlCsG;V�џ�	�l��u�rM��L� ��H��T�Ń��S+%�(�l���O0�PI��s!�S��1|u+�W����N����,�u��N�|��݉>걟H�aW��?jJ�ԢB	$(�\�"OZ�F&�!p�xB��̙	g��CK�>baf	�qgL&G�ʌ� �Ϟ8��O�Έ%�H�c�׉�L���1�ʌ�b �L�#W�M0��_��K���g����DA�?t��Y��:f���1q� �ɥ	�$D��l�VA>x����&���	ۅ��JG��@��p+�&^�+J�|ѓ�w1.h��'��"�Հj�\T�P�w��S�'�`�*�
Q)m�<P8sE��8�X#��� � ���`�ܬ��%�;{��3'"O61�� Y]�a�ƢC�Q~���'�����Ŕ!���o��(` ��m����c�LZ2B�ɀ�։A��,����+;B,>b��鴋E�@)48!���CO>}yu5�L��2σ�>UB�	�KƘ]YdoW������n�8o�R܂lYG�t���r��L���ӄ�Z�vD`A@t����14��8!D�.7[��C�o�,*:�q���D$�"��;`��Y��	946��Kf��9)�b�R�f�{��󤙸*�z�2 �'x���Q� I˒<�i�
|��B�ɂ��"!�Z4ל��2�p�O��㒁v

� )�'7���3&>J����'<p$Ʌ�[��|�ŏ$5dx]x���r���˔X��I�'Z��%��>� �#CwĨt$�%$ٸ5aZyh<iTE�(=d( ��Z5�0�x���&kQx�q '�E��i-��g�4��yPf�Z�C&�M��5��eha��@#�I�w��P�&H4���QnE�V��ņȓ0M��X��*`�Zm�Î�\eB�<�C�<^`H*�D>�'840Dɵ�ʷ�%y�mIr1D�D: �VTǀ�*!��i�č!s�Ф�jIM>)S�0�gyR�Օ
�v�x2�P�C��@�AB$�ymU�}��x���*UN
�b���y����,#�Ђ�� }�&��2e9�y�+ɻlS�a�0�O�hɸ�1ㄮ�yb�ϼi�f�k4�	S4   !Cȑ�y"��ph욱���T0��C����yR���5��ኣ$ٽ~����c�C!�y����l�<(H�(ã[)��H��y�Z�2��L�S�Y��/��y�a������!ذI��4�eC1�ybnN/���Ұ�Y)}4� ��& �yb�ُ~���0R#�0e�Z��7,Y�y,��Xe�-���Qf	�k��y���+B`��-,�&���y��	'��s�Nͩ
l*����y���0Yfm[FnO�%�u���y�f�4e9p�'��v�1���:�y2���T�t���ڑ�����C���y��ڻFW�\{�B
�wp��� ݀�y��5:���f`z*m�K��yFk5���d{���;�R3�ybO�>_hث�$X�i�P̳�����y"m�>]��C�U6ve���t���yBᅸ43�u��H=[��0����yr�R	%u��[b �ONL�Xv�Y�y���V���K#�Z/�<��4Ó+�y�mګ��a$D
���Xc�J��y��ۡf����`�
�|�HI�g���yBL�a��'�#�|�[�Ͽ�y��5��)g�%�pk�'��y�C[�/���e��#'����V$�y2�Ĭ0�l9��N�wpM��j�*�y�
�Fk&Lrԧ<Y`�3�!�y�X�R)�#�&M��R0G��y��#[L�C�¶�v�^=�y�˕�_Qn�`�P��*�'f��y2#Y�4��5�����,�� ���y�·7�Ptkta�R����� �yBNA=0젅.��O�P+F&��y��UQ1�������B�D�[����y��
��@mആ"D��x&cI.�yr!�h�hD�$�A�27l�@u�I��y���z���@oG�e���M��yb��~���K��Q�+]|�cc���y
� P�Ru��5?��A`��%_�1�"O��xa�� W��rAJ�;k�E�"O0 "��n�!��oˌD��mS�"O�P�˛iU���G�D�����"O�����c��	�����+#\XS�"O�=Z�l��TU�0d�)U�=2�"O�X�s�ؚ�|�SP��bx�S�"O�Y�����CUś�$�"i(�"O���tC�I2��9}�`��"O��kS�	�A�`���Je�7"OBq:�ɯ@-*ᛑ'ε0�2yZ�"O�	��k�gI:L�(�I��آ"O60&�Z&t�Db&�4
���x�"Oִ��KΖ79���Cھ!�$�G"O��(�4#���$�̩@l��"O�"1��m�L���J�A"O�Uh�$oJRʄ����q6"O��+P���*���+r�8D�S"O0i���L!a�D�$i�$���s"O�(q"A�Tɐ��.Y|PP"O�� �.U�mLI�Z�=�x�	�"Om�!
S b�,�3΋:'j(S�"O�k�"Ϊ_n�08�L�Jz8�"O�aچk�^���k3f@���"O���L�.�B% /+Pwn�cV"O�f��Y��l0R߰P0�(�"O���'@�.]ǊQ���``٠"O�@8��T?���3�U("�K�"O�p�|B��dś���:4"O��F��*ׄ-c')�1_B8q"O\�x0��^ 
Щ��c8P��b"O���V
F�6�P�@��]#(�L�"O.�*�I�� t�� q�91�d�"O�qK��t�iQD/��E,�� "O�iz���:xJѓ�9. ��Q"O�|Hp(�34r���R0m�"O�[�°���@n�m�E�v"Oh��(V6$���N/�H*�"ONh�`CBF��$ҰX�P�z�"O�%I�C\VH|��IǶo�&0�"O��3eMK����tM�)sȊ�)"O �k%��a_RP�� 10��b�"O��j�aЯd	���B=u��q�7"O.����ߏG�ɰGB}��
�"O�jwMݤpI��0eL?lr��"O�@�Wn̰]���Qe�: �ܰ��"O�=2��f�ua$��'�F$r�"O�ܲ�GȪ5SΔ��c��+""O6A����E\^@RE��/���#"OF	ۦbP�k[�X0N]����q"O0\��.
�HC�tIQn�7(��q��"OZ9
�$]��.�,ى$�i��"O��#AĆ8�̱�)�IW�$� "O&�	�nG<Gq��S�h�#cFH�@#"O�A{�WW��PY��M!
B j�"OXP�H��Vgv]�"�e�4��.Bt�S�g���U��:� Yq�T��B�	(%���:�bD�X܂���$ ��6��P\X��(=��s�.��.�� N$+`j_�x`��)T"O�YB&��p��p:釠c��+��O܈{ue�K9�ӓV��
���7�>x�#��<#�Fe��	�t���K5a�a���Vi?7�๧苳�T�`�"O�ؓ�U�l?JAz�ƎL��x���=x~T����Tdy�a��+����[O�Sü�pj �� ��!�ǖ_� #e-Br�<� Hi'l5$.)��n�r�����t��ur�X�$��O���.Z����"�yr�\&^,�QuiЮA,`0����p<QsU�@�����W�#p����W�y��d:6��P�Bf�5�~�I1k3̵��'ĕ0AazB�$ �\��p͇��j����Ĉ�4L9
R$T&6I�ʤd
z�)�<qtIȧN�Ԉb�.��{����+O�bB䉭`Dy9�Ɛ7	)@�aFě�f����5gQ��b�dRN�)P(,gJa���B�	�C4��
*@�lu(�`�?*�)�g�H��D�+D���sR��D<RJ�aUh��5 �#0��T�ģCBi��Q����!#�=��(�=[��W�ћ3��W�'.��J4�@A Hq؆/�;PR�8����z
�!P�ԏ"X�Q�/ΧM��	S=�hQCd!\O���dY�%�2�3QQ"�R��\�T��E�Cy�,
�N��>5�v�Ie��hŸb����$LҒ��%�h��=K�i6l�!�aMB�m��s����Ii�F}	`�G�*�(g阻Tq���&	�צ%�Ըź��O�A�;L�-�Em����R%��ZĎԄ��N�8W�). ���$F�f:j��'�N�vi�2�Q�Gd Z���<y��ʊBg"<��(9�D��r����tr$(:r�9џ��q���݁��H�~0\� պ��8�8KR�Y�O?`�4���P�P��ϙ6q�$��y�C_�S��O��$���#wJ׎��$/L�mig�4��OH�qY��h�s#jS9"����4!�q��M(�2C�	+����7�q���ʽ>^���f%���p��o���7*�Z�p�OY�t��%[7>���� ہP����'����:
0�}h3�I���U��*_ |����4q��5�(��iI�W#�pԥ�6'�ܴ
�"O�qa��a����71	�t�%����	K��(?�9�`7<OX��d���	xr��4b�hr�p@�'�0��Ũ�A%�3���i6�Ranدa������R��qW-:4��J�
�j��I��sR�A�48�I�+´EbǌW�eP�M��.�S� �Si��| +�"�� �3"O�`1��|QZ�9���D���r.��p�gE�����(���_� *P�C�
�$S�� q�bB�;:�V\��8-�8�Sl��^�(��#��iR �s�͢<��z�?y0�Ca�$� z%�;�p=9"�ɀ4�F5�Tn��MSO�{�]BV�	��ʙ���}�<d;!�IH3ό;Tdx�@�U��9 ���5�Z�D��G2�ހ�Daŧ>�!bP��yR��,ҨIR&R���-C���'wAL���a��'a&�'��>�ɉh%�A��@�"ʲ)@� ��)utC�	�7)����8
���J'�.�4��_-,r���o,��=��۲8~�Zw�.mA�r�I_�l2H�	H���I�0H�x�%�P� m�wh�G8jC䉎D����)Ҫ?��eoL*���T�e
�	#�?m��M	�I��������>D�T{ �F�h�%��KJ�0a*���:D���c$̺dO�i���%J��dI%D��iU�� `=�����Z6jY�X3�j D��A�ꐴ1tz-��Ι��\臫+D�0P���;�pA����s�p���I+D����U�9�}r�%�i���A��++�Z�P�#]'_P!��*YE��>�O��a�� m���gH����43�O��1���z�Z26�<��J	�+�,��a]�C�-CSm�-����O/ph�!(�9ؐ�x0f��*9џ���iG!u�|{�"�� ���X������RG,��q)�-���?��x�1O��x�n4b�X��G��>���0�Z��B����?q� ���A*|!��ˠ�+T<��D��U%��4Gy2BK�
ն�["O�|��@Ùx�;&��2�ҤIi�4=	>�ه�y�Nx�Z�2:��@hN<��'ߜ[��!��$����e�W��xɶgޟ^��ze�õW9�!
&�����o�,P�(@S�C�"v�|J��'�>�Y�FW8��Sl�T����$I�7D��"O�C�\#4�ŢIp�����7m>�Dʨ'���1���ِx�#�*X������7�Lys�,=��޳}.�0be�L�)�\�x�㋔"I�=���t!�<||�p�E�{A��@#E��y�Ł;8I�l���f͎�I�FDX���DH�_t�I�lx�Ҕ8�����p�	�D�*��7�If���z>�9���"6Z���O:F�.�)䭝+k��d�k�K�iBB�ҭ��(͆��<� ~�� �� ~�]��JX�0���'��iW��+`�`H�n��^|���F2�a��H�`W���*�Y�<��*tt��&(�!���@@%y�<��0eLm�ua˪t�n�t�C�<)W,�u,�!��R+=#��q�z�<9�F�I�
	±���P !�q��(�a+0DL�'��R����I�e
�������'H��!�.�#��� {�2Y�y�Κ�y�8q��]�O��cV�u�9�@�ܭF	� �'K<=8�%��m\���A��u��$P\���.Oҷi.�3}��?�Եbv!Z���˶$���x���4La��V�|�������^� �� x=��'F�ҁK�8@��ܩ�E2[��3�A����!�1]��#�'{��+���#"|�]Bq��.�5��' ��a�NH`�#E
?.�Z��N>1@��=(�B���@����.���K�f�!��S17g2a@e"O���XK�1	�n�I4����ΣW����T�ؘ�B�t�g�dƙ��E��DJ$��tW�&#g��dT�:�Ա��Y/�f���K�P���
�9=���+&�O�����eA5�O�s$0�"�'��qqEH�p#$�2=O� �B�R<,���(���7|@p��"Oޤ*B恴Pm��8@D�*k��0�d��(n� �`k�*���8��!ƃ�KX��Y`�w�%b�"O@�jv�*N���9�@�-@�4FĮg%��&� ��<!!��U�1����Z��1飮�T�<I�� e��RM{}\` D�N�<��Ev9Ҭ����P�Q�m�\�<Q���f�`{CAA�Q�� r�<�!�Ň������c*�s�Gm�<I@�1M����;â	1'"�v�<�'IeK�`���������@_�<Q� 558�1���-<�썈F��P�<�D�S�r�61"F�5���_M�<ySą'6�p,�Ï Ϝx�u�A�<I$/��HB�:l���	���B�<�G�H�ҕ�� �l3�9�r�KP�<�0� E:q�(�{m�NHW�<!����SH�eIvcE'y�D�#�$SF�<sB�|��5���	�[��_�<q�A��]B5a�U���H���W�<��$�{���C � ����a)JM�<�q���ugR��DK/�lh�!�R�<�U��	J�V|�@��:>�Z�H�n�P�<�7�Ć_�j�90`�����N�<��C;J6�*��gV�����J�<��K����~|�D�e��jE��_����jѥi��i���r
 ��ȓZ��0!T�˔"t��h���?� ��!cvD��K:��ݠ�A�)B�ȓ
.l!7j�(a:��Tc��<�J��Z̰q�d�F�\���߀_�0��F��� �G�^d󤍘��y��^Vp��ē?[�e3���?4�r�ȓqiD(��1>�h��4 D4eXXɄ�+I<��!��/�:%ئQ`*L�b$Rmd���J�jɄ�	-0���W�g� �[e�	�{_lB�	r�@�j��ԕ+}�i�Ǝ�n>�C�	�/3.ب���?
Sz�1vFz��C��*N%��0a�"P�}PD�>f��C�ɬ@:X���+f�P���/x�C�	����z�ɛ�<�+d)�5w�`C�2� �7&�i�����5!tB�	� rc�N/0����ǘV�>�I���V�<d��aݝ��+,�
.� H"A�' f���� W%X�H�BI ��҃\Z�hI~��� ��hA�J<�(b���(�J�2e�YI?	G)P�u��AiE�֩�0|:�!�0 9I���I\"�:��ܦa�F@�'�R��#�Z6�)�'������k����F��<b���勄)���� �:l֝�3�����0�Ov:e��I޽"��0Z3��$I��q��n���#b�N�ѓɗ<�O�q�FD���ۿ`lDL؆��T���sB?���'cRmxf��I>�	ӋF��lR.����N_~���q7�[\>���&=�-�alƜ:�d��b��4��N�c2��y6�|ʟ�=�Н����>�(�+�%�����x :l���өnQ<Q E�K(g	CK��<>d���S����u��4�d�S/��U[*�A@(A�TͰ�h�"O��҂��]U��(a���]!���"O$�K4��W=n�n��(M��"O2�Jbn�!~bMn�T�5	�#D� C���5���\�-�x�rO!D�$Îͭo���� �Ja$u�>D��Ap�×t��c�ժb�VU0#'D��0�˟��b]���T�9�KU�9D���ӈ��:�|�"-��py�Q3��6D��;qG�2	�&�{1�OzY�1��?D�h鷀�&lɊ%��hٲ��i��B>D�(�vg��s��Y���Y�={�%Q6�<D����KߞCv8�Tʘ9PҌi2��&D�<����"h�A�ŬE�(I;t�/D�P���
	nrm�qG��aJ���"1D��C�
�*K*50��O_H�	fn-D� qV�̙F�4IS��zW�$��c8D�$K�g�y�<tC��?�U`S 5D�Xb��U/=�2<�k-l�@v�1D���B"�^�*MK�-�p��M1D��3���J߆�:�Ĉ %����J;D��;��#G�(�8�C,39�
��7D� ���޲ys<�"�莔 t4D��8#�ߠU��9����f^f[�=D�<(���a��!�!��P�V���7D����>(Қ|�Ԥ[$luT�Ť2D����!W�B���A�W>{$�#�+D� 4DĉG}ޕkǎ�,L���AG"/D��K ��4{�(P��E�ot 08gE,D�̣��m5�v�B�k���xg�(D�d�d�@*/M�<q���$FB�+b�&D��h��	]"5����0LS�!��($D��i��M2L�>}a���|���t�!D��+�J�n]K�M�bM�VE-D�(+��	[��k�ǝTD�5�tN-D�L��E9�;`�*K�)х D�H"��U�$����#��A�yI?D����@�OK�ЙgEٛ8���`WH<D�\:��:LDK����R�����@?D����$B�Y�jK� �Az��RD<D�t�EW��8pd��ހ�ra@:D��*���sX���ЂP~��	e7D�h#oS�V�D�f�	�S�dC䉴"��1Y�R$	`M@�A�x)�C�!/�@xy!gDtX*��Q�yR�C�I��@h��#<n,�۵�C�30�C�^U��x�ʏ�(��ӧ�?f�~C�I��^�3�\�#���h^F�|C�	v�j(P7�� X.ڬ�A�o>C�I�Bf"�q�I a�L
f��"� C�ɂ6����F#2�����T��C��2c#����jU&��WB԰|��B�?s��)�ˉ����ʀC�I)
�H1��=+� �%΄[�@B�ɝPl��:���.P�zt����z�8B�)� ��s�d�?h�LH���/CZ���`"O��[&]mʠX6́=3R�4��"OB��+ �y��q�P%WM^81q"O4�J�JR�s����1+�$yG,��"O`���ҷt�0����4���@"O|�$M3�T1�*N H��`+�"O�)à�	:E������ɫ[���b#"ONA�"˘n8�uZA�T��EP1"O\a�
N��Y��LZ V�޸�k�<�ĕ��P	��Z�b�I�OQ�<ihR4b��8t�0_q0P1s �E�<��#�u�"<#C�σ�L�A�B�<q��
[�V�j�V�W縰I�G�<q�h O�}�'e��f�f2%��l�<�$����1n��W�I3d�^�<����Qo^����8�%k�B�<i��ܩih����ĒurQ!�&H�<9f�G*-�Z�5�Z2�DAw@i�<) ��-��8��n�&�H�-@y�<��D�[(�!�χ^`֨h�/^r�<��G�
��5*�6l@���g�<�R+d�0�"Z�P�pᥣLK�<�MG&����Q�Ll�<	��	��	�W,I�W�>uʠ�B�<A�z�6��СP�@�N��łt�<��֦E�n���lH2Jvd��L�o�<��+�?v������E�Z�1��g�j�<	�F��Bm�])rͮrht��#�d�<Y'�9R�l}!���~�TM��_�<� z��`kQ$8��Y�]	!�].uw0��'���T��)'��g7!�Z�e�����+:����\3#�!�$^'f$X	�GE%P�ǎ��!���E�ҙ����G4౧�R&t!���w8
�'��Nd�H�W��hK!�gĴ���3AcRY�fFN@!�D�<X�`����a�naad��Z!�d��,k�|KV,(5��
P���9A!�DX�!y�m�D��*�!�b�*!� <|�J��>�Љ�+ۖF�!����tmc�c]<O��4YPK� 	�!��i��	�KB?�j�Q�	��#"!�DA�.��`��~�R��5�Mr!�Q)O���A�E�/��U����A�!�d4cMp�!o�3���-�<�!��C܀hK���<�|��"�\!�T�7/��7!	�v��1d�J� \!����8�JՒc�4U)�$}7!��Ɓc����°-d����*I�F3!�$�=7i����f�;[���	���*'!����~��3CE�u�hء&	��j�!�d�� O�ڶ��g���ѨN �!�D�B���t�_��|��]�!��:z�TA@6%.I5v@p��"#�!�$�)4�c���}v,=��F�^�!���8K�쫲խwuԽ"���&	�!��	���+ 	�gk�tR4!A�]�!�H�^)��ÒA�4?L����Ə�!�� P�Q�Ԡ�($>���`��Et!�$W)q� �����|tO@�SR!��RBX�q"��>rh�y ��N�k!��u��Q�'!B�?��	�B�ԧ1!��>:�"18B��P�JA���_�7f!�$W���)灇�J�9YQ��;!k!�� �4��'V Ēl�E�I�Ҏ�s�"O ��g�E���p(@]>1�hL#�"OT���k�5=���e�M/4<��5"O�*�6�z!��N�K(�XP"O�e[�ǂ�X�lɲ@$+vQ��"O�ȩ7�%�ҍ��E*>���"ON��_?�<���.��U�"O����B:l� 9��`S�n�zD�@"OFA��H�*���3��_�>��6"O����g�X��'�7q�8�@"OJ�� ^�I�$���_2P�����"O~�#	��^�P�F�r���C�"O,|G�ǂ{LYh���8b$H�"O��j��%�txq�տ%���"O��3�B�2f��(cD�[!&��v"O�K��h|
y DSy�-�"O������2j߸�����&n� 0��"Of �g�͙;�c���.Pz�鑇"O�I�%�3� ����`ي�3�"OtQC���	�|I�������ؑ�"O�E���
 }�`y����z�¨�W"OVpbqo�2\ʨYg� n���s"O6y!�!�.#A��c�#](8�����"O�}O<��h���C�kuZ��"O|bq�U?��}�����\N4�F"O�}�Ң�\�l)D�
����"O0�+҄V�QJ1�2d�(VQ`��"On՛�"aڲd�����(��"O�!�tl��]'qk��C�=�> ��"O09e@��k���{�B��\�h���"O8$ʐC�V��他��48�>5��"O�=P��o�.Q���5+��+A"O��w&�%͒ {��K�'4��"OV[�[�0Sd�pV�l̉�"O,���!TN����V4��r"O��ч'��[������R�ij��C"OjAi�*Gs���'Hï^�4�S�"O>a�� ��!a�W�3��4CE�T��y�HX'2�DY�Bђ)��u�s�'�y�,�b��}PV#K^
�Hd��y��܏l�1�P�L�>==��$X6�y�h��J��u��E]d�Ձ��y�	��Ai�u���>>7�i�����y�Īe�DR���/?e�qQ�bK5�yB��TG�� R
O;z��2dJ��yrF�5�M�ɑ�U6��c�y�΃�-$�xc�KB�x�h}��)��yBd F���w�G1#��j�JW��yb慖J׸��v@"#��}�ń�y"��_�<h�$�ϨC<p�˄�ǖ�y�9k�0��i�V�Ʉ�]�y��,��]	�
�Z� A����yrfԐw�܍@�C�VKHU��':�yb�g�6��0�șK�KB���y�
�O(a�!-٤���M��yr@�_4��s���t�)�r��y�\��,��rd�1jG���솨�yN�9wh�ʅ	�f/nh[����y�� �-xc���6�fL�a��y"g@�x~��@�@��| v�"�F�yb�̉�x����h�"��3퍻�yR����>`ˤ���Iط�y���(b��]�#�V<G^ISA���y�"!��,I��I�t�2��C\��y
� �:`,W=:�rHC�,A+*�ȍb"Oح�q)٬yU2��pMV�����"O ]�G�ŤkΒQʗ�'�q��"On���à_W0\����k��8he"O� r�@36��7����D���"OJ�SE�O.����A�W"Z�f�"O��EPQ��-!!!ގ,͎���"O>��"Ǚ�q(Xp��@' ����"OJd��e�<(���O
1A�c�"O��s/�7b���3�`P�U3��#�"Oֈ��R#T��P`�7L̰��"O��@"#��x�@$�&6�@��"O�e��M{<�Ҕ�-x�4"Op�J�
��팑 �A�=Sb�aYr"O�L��B�K�R�I7A��a�(Yc"O��d#ݍv�@��`
A@^6���"O��JL	xix��0^���"O@d�˞�-F((���UZ°�5"O�<��c�H�xEH���0D�pK�"O�Y��D�H&L� (ǰu@>h��"O�\��   �<� E5_�xH3�ǀ>�yB/B='�BtŇ�I�8���+�����ʎd�fA�a'��O �c���4:x���@) �F� S"{��E���Ț�~"⇙��GxR�\�~��u�mL+ R�i��R�	NVi�W�w�̼F}2��ti&��ĕ'{4ҍ̪�x�!��F�'�V�0Ê�z��a�-c[�O��:�슎2E�����D�'h�d�(�2w�N����90��+�8;vY���B��"E��c@��ħx@)�V@,@'�Q�_�ES���l��RԂNv��ӧ����`���2r��K$�����F(^
"�$#�Mѻ I�	;�k�j��OC�!{��LR}r`H�Z�Z�i1��\�E*�+���DƱ4/���4�װ��O� 2)�u�Y�k�H�L ���>9 G!�#���4�DS�"��� ���'pr0.B94�\�ȁ��y�gn�%@��)R��o|���!�v��A*�M�7�H�q`�jxf�zƄ �G�r��E�T������	�7���8���C�JJT��i	"2�<����T�LY��''�ܴ�`��Ua&y�p��(D:Bȍ�(�OJ�*�/̓S�LTjB 1�4=�	�'p��p�D؛z*g��$7	.q����4I����gR"t�Ls����'q�l"3��>	A*GѼL����^�:�x��R��$�O��
�L��׈�|�ܱ�u�X&��� Dy�<�G�]Z�yjA, 	������R�{ �d�Q	�m��ɚ�H#O8�#����HU�|���%E���1iD�l�>I���G${0(L���ԼtLP�f�3�O�PF��7qW�,;��� �␘r�>QV"ӕ@>��	Q��)��|��J�d%4c>�W#˓b�pmX��3G�l���9D� ���\�-8F%0N�,R~�b4J�h��=��T��	h��~2$V�nø	�̡f����Ɉ��y��O,[:��LI_:��uـ�?��#ќ(ǌ���c,lO2����Q�y�\h����W��@�%�'Є(U�
�\�8�n�<��I�ƙr.�W�P�{�TB�ɤo���h(0��@g���0⟘�CBǀO��-���ӾCr*)�w�[1+���p1�"O��Bc���9��qC�1I�*L�F-0\����]��"�g?���".2P3�c�/*s��r�Vo�<�Q�K�\�M;P��%^*r�F�`�	�Y�Q B�$_+a{�?w�j�
"d�z �0P���0>	��r8n  ��\��YA��8d��3͝-rc(��ȓI��u*��ީ_����J�}�B�Ey"iԟH��qF��GQJ�@)G������!��y��5
q�4�e��H�ƛ��yb+ߣs���:$�PX�r�a��y2��R�r��GC���¢���'AZlq�N}����+�f��<B�K��B��Ih6�9�����.*#*R�)�	2żI���[7�h��r�`��� ��T��H�*a�LM�I�6���	1S�.ђ�-V14��O): �F+�*R�J]8�E �W 9��')�઀�8/���5i��K ~�/O��ҶbU�d�"��M��|�A%8AnTt�	٩��`��u��\�ae�8H�"�����%0��35���&���>�7��7ET !�1�\Lx�JΎ���+��b��F~�_�Rw|T�土��Ė=E�ތ: ��YR-Y��Idid*�)Qa"���Qs�(z�.�V�I�X�j���5���� f�:ʓPv� ��1 S���pYC�4ttf\zOU�$Z(��"O�(�-?h��ٗ	7D���0�Q�`�V�^=%���GC�F�iȿ@�	"�Ϧ>1��έ3��<xv�5,�@ +GM~��i㏉�=��4��iJ�+0���Ԯ�s�����Ȓ*����v�����_uF�"?q���%-UH�B0d�p@H��g��X�'�"D��eU)Dܕ)'���<Ha�Z�H����_g��CS�S�*�����@���C�
P\B�[c66�*)�.���:����9��ן�p%�K/"±1p�i�5��ĳ�g?l^jH�E���:�.,;�O�̓��ԃ�_ {�h  cZ�'��Qh�"�O����0��bO��"�t�<�l;�#ۊ"��`���IZ!wL�YH��b)��D�g	k��-�6a�ڟ6���S^�,��坾{d᱃��*� ���xQ��S���9�����C�fQ6���d��nH�`r�ǃr���pu ��	D�����T�^�)�����d��n#V�%E�t����#@~��;C��Jm�X�t�&�~%*��'}�h)�I�88��f
�E������QDP62X�E���!<Y�$�d�rNe[c�^�$ϔ�;&��0rV�Z~����ՆH�0؅�	�$�� �wKp\��2�τ;d/�"�B�y�H��刯D�R�;��d �IٷԚr^�SF����'u,�aS*}���F�$:D��J�'n@92#/ν����'�ޤ��"�/�j-Z@��'����G�*��bP�V"����ѻiq������{��(��ŊH�z�Ӈ�L�w���/.1��(0����M��9|���JW�]~�9cc� #)Y�}8���;��t��K13~ �
� ��M4M��x�0�!x�i�f����"|�Y�枀q�(�֪��s��9�G
i��%S���*!e���^��pL�S�B�I%R��\@�¤i�~���KT�'nX��I��6�(L��O�}�NR��ey"��fd��su/��X�����\���U�PbP�y���1q}�x
�͓:8-rał���'(pxJĂ
*�ax��5f��8�ӁN�ﲵ����>�y�!��[����@{��Ԋ��yr��X�|��w�.MgN9`�O��y��8 �Tʔ�E� ]($��y"l�=]U0����9=�bipW���y�F-0��|1�h��7�R5��P��yRi�M�����"�����Ί�?y�dЌl����|;��7�ϸfnޑ2�C�%�a{ͺpF�h���O��e
8%90���N6p[���p"O�\��_871��!PNІ@�1���DÌ"�]��E����jM�)B�K� ɐB�J5)���"O8�j'b�6X���yV @���cсҭs(p��>q�b#�gy��ް4@�� �G�dkr�Iqꝣ�y2�D�Mzt5B�@�%�� ��kK�{J0��V r�hA
�iktȪ�x/��P�#Ϲx����Io4�а�n߼t��$�(�>��U�_�"!^�Q�K_1�!򄓲=$ұ�2�\�o�Rm�����qO��x�LT�r���1��i�"(����5tPYw��'s�!�dX�%!ԩ��k�$h�`�DL׭[��-
�B�(��Z�D�|�'Y$A���ҏ޾p����#f��m)�'�ʤA��'Z��0+$'�SL�|1ň�
�a��i�3�0>y��܀�PKV�s)nx���A؞�z3���Mpx�tG|�ѥX�/�h���!7mr��ȓqP�]���b�1 Da�,M�?��âh�"B6��	N4p!�@�LOD]0%�Fz�<q�&�LV�ԑ�P�1G�\���u�<a2�D;^k���)ݺ>l�)�g�Wv�<�U���B����DZ�l���(�s�<�ǩkIz �q�Z!�ӕ�Na�<!�Ő�~�hb3d��"���2@	j�<QP!��`�49j���9B�lDZ���L�<� h �"@�!�����٫Z�hʅ"O4i �I@�]���8����"O:���	 ?~1���2D��w?ʉ`W"O$� W�7�<���7^�Je�u"O4���jЀ[Jlp�sɳ+b #�"Ob�r��	�=���K�/����t"O�%��RHu0�@�%%Ȁ�J"O���($'�1Y����^���"O��(x�p����E;!h�\��OSb�<�F�
�7�@�1n����G�<ٖ�$
���ퟙl׆(6��f�<q��T=/�bL�b�	�F�ܻ�CS^�<)G�R2�!D�)
%£a�`�<��R<#C���Ac^�v��1j�X�<�PO�!e�*S���d���b�R�<�4��-��UPtd�R`�i���N�<��kL/:L\�`�?�0��RXF�<��ǋ�{�"��%K�!w�T�1��v�<����"�^����B"�m�u�ȓ��:�� ��i��"�$ǖ��E�dt��E1�n��S+P>f%��R��-��Ȍ)A��hjP%�sFf`��$��@�đ�\��	r"�ڦFa�0��t�ܼ�S%�8�c�!���ȓ�v|B�. <�r��23�z�E|��5����Z���Xd2���H��M���>D����.�9T�B��.3��!��Njϸ��CĔ{-�B�?ئU��ӷZ��u1�m�#�DC�3kT���I�PL�qC����b%(C�	3T$�%���)���N���B�	�W>�<!Hm;�%ʝA��B��^�h� E�R�J���F�_�B�	��Jx�B���PH�N�B�əx���sM]������,+�R˓m1B�<E��-��(1̕��\�"�"Y�ڱ�?��<�S�OQ���m\�z H���M.�bܨ`��O����8,�B"|�A����s�NTNU�|�qe���%�x�aE_s>��0`ݑ��y�'��><BS�2����<8JC�2��La��?�) �øo�$ ""O8�æ;�Q7��L�:�:�"O8v�׏xꄋG��rN� A"O"��l\�zu �H׀�1�fB�IP8�L���<�Rn� x��)��#D�TGQ�X��)��+ܳ	�����N=D���-�[��@cj�3i�J����/D��KdD�0o�1�W����(�҄�.D��Hhҁ^�8�G��6<s�Ɔ9D�̙���ɪD���5It.LBBi7D�l��-] 5`to�(*�A��0D�<떫�7������}��Iza.D��SC�:�ԥ�0@F�Z+�)���(D�,��"�S~�]���+n0X�%D���wm�'`kp%8�KC��4���!D����.��b�����B�	�����*D�@:E��^캀�u%�=iL���E'D��́k�4y�\���+d�#D��;�C"H��	1�� ��q�M=D����k�Z�~Ţ"c�3D��	I��>D��A��C �U��#�7{��
@7D����mʕ)�N�b�MC8��I#�`:D��0aG� {I��+q�_1E�E�6D�������g�"I"�J�+:e3�o3D���D�Q4� ���ئ�*A�`2D��U�^�"�\���<h�)('c*D�� �H8Ə��Ib���Wg0`��%�"O�\9D�9B��8�f̅U��T*"O��c�ė�>��6�w���Ҳ"O�����7��9K�㏇c�H�S"O"ux Ă!o|h`��"ĵ$��1#"O�E�r�� g
$#T�%�DI!�"O,���0�@�
 ��M;�"O��X'ʈ)VѦ�yb�Bى�"O����KN�fj,\�qd	��:�Z"O�1��@�=+j��@d]�8k2"O�DÁn� g<��9�CU0MB
!Iw"O���b\�*l> x��L+g9rᰰ"O@�;�-��/`6,�QkC�9�@��"O�m��kZ
G�00�0��-J00�"O��Zv�͉1������]f"O"A`���4Ǹ�Ү�9�l��u"Oԇ1</��O.X��"O��2ȕh�`K��X�ڰ��"O~ �@I�Y�4	RQǹ*0FthQ"O<�������Q� 1����"O�u�We��*���H�G�5^����"O>-Z�k�<�� ��W�R�4�w"O���5��P�Hj0��'x�`�f"OLh��T Ev0�#G:1W��y�"ODћ®�C�xMx�r̹�"O�}�,�,����\X�Q1"O�-��̭i5�-*[e�B��%�P_�<���$2jb�W	
��āR�.D�8C6���Q�4�A1��1XE�(ȃ�9D�8��M[�T�$�VC�Z[��p�b8D��w(�`8�e�S�8>�AH��4D��R��Ș�ȁ�`*"
�U��G-D����nB�S|<�0�
U�3��r +*D�pP1�	`��5)6����m)P�-D���⋗G0ĺ��`�F!D����"�� �2Q!�M�|�l�C�#D�{�5�H��&��QZ&K/D�t���׍_�2�Ac���V|���+D�p�VMֹ:y�A��	PC�%q5'6D�,K �T�Z�Tq����0	�f�5D��+#G�'��)SJ�.&���4D�D(��D�>��|arI 9I1�H.D���֩w��+V�ܰ�$d`�'2D�4Y��G�[�ڼ�P��c��
&#0D�����7�&%! �m��iۖb,D�D+ ��b���@*րBB�;�i,D�!� �=~�������g�(D��P �� $�A�K��,־��B�;D�Гd䙦St�(��&L��&D� "�ʓ�!@�����%o�"�B�"D�H��� M��q��^/TG�S��?D�t�ǭ�@Ȳ����+:��}%>D��s0!�I->d�ق)���I��&D��y׍����S�� =*�� w�$D�� G�#��1�ф���K>D���u!�B���iROLp%��M<D�x�!�ϩR�橒�)�dx|��n>D��.��yRZ�@��$K� Y�f'D���T̛�Ū����>�:�0D����A���l# I��T�C�� D�
��־,K�T�	�91QB�<D�,��B��I�g�.!?��!"i8D��悀]c�ݫ��?��lI��7D�\xU(ĭO�D�+��<��w�7D�� z�ďx�!9�ǂ�x�PdA"O�P���6�R Jcg��0��a�"O�U1��ٓ��X��fY��"O^��� wN��,� @m��#t"Op�e ��5l
��+�^���"Or���H0Z[��R��Z2(��3t"O�Ms���0�jݹe� �n؜�#�"O.�����9<ExvF؎o��TH�"O�8ĩ�u��[�DM�i��� #"O�ɛ�-ˊ!�r�۪)��`1"O�bt�A�1Kڹ���ʓ%�����"O]҂�+U`�l����)��3%"Oȡ@��7b�$`s"�P[D��i6"OTI1R���T��B�|���"O���c��>��9���5�`��"On�f�[����I�
�hX@��"O�� H�-� ��6)��dB:��6"OF��`��2Hv�a#��=B��iZ"O�`#6�ߚQ�����oº:����"O�er���05��x��+9�ޝYA"OhW.�IF���-�4v%���e"O��+VJ]�_/"M���$Q�"O�XHQi��*KXQ��H
R���t"O����w��E��[)��=�"O6a�F���ZU��'C1� ���"Ov"�"�!}�e�  �$�tl�"O�x,�t+��ǂZIfT[8�!�ҏ7��#Ԭ�>A�!��ͯ<�!�܇p����iS".� ��ׅ�!�:5!b ���]�4��c�%��'$Բ��ʲX����I	�Xvl��
�'��9�+P����:M����'ҕ��C2���K"2�T���'����A�936�	���*�6,��'�|ʃ)N2��J�ɖ"rfy�'堘Y���G���g������'c��ǭŀd8aq抉��
�Z�'���;2a�a
y�5/��T�.9�
�'
p�a�L!6��{��F#��
�'�h�s�ыc1x��� ,�B��	�'(rdRE���������S�I
�'|�}8҈�-+�ڤ�'S�!��@�	�'`�
#���a��<��Dq,Q�	�'�bm����Pm���p��'),J���'P�q�fhI=�� � ]�|��'�]�'�	�V���١d���i*�'��H����)'@�i�.m��I�'%¨cP#�(6�>[(��w����'k���M6+,����ѷh�uB�'�12��ϛ2������ڤ�	�'V�q�.�af-�D����~���'-��4LZ�s-:� ǌ)�0���'{6�rqF� 0�!�D��9)� �@
�'M��R��,V��m��a�<�t�C	�'\���-O Zۄ�H4LG#
��@��'�4ʰ��^�i�3.�}H���'04X�5.�	R�nx�g�V)*׎	��'ʀ�J$
D�
n��(�`M�%�-�	�'�PR'�â[L�����ž!~�s�'�%��!�+">euMA�&"}h�'�H�ʵ�/)vؙCSw~pz�'�F4��݄,{���e�DL��'�ViqT5�6H���U�6����'�dB�-���5
!'섥���� p����+U���D^k����F"O�0G�`+dU��DZ;Z�D�b�"O<�Xd�8Mf�,�֣�v��p��"O���kL`J�|9��Qu��B"O��QЄơu���Y��`� ���"ON�����N���b&�X�~<X�"OT���I��
�����j��!!�"OE����\X�$YT��;c�6R�"O�]"��C�<uk�3:�d���"Op(;�����"1 �*F_��U��"OL���C�?#>F��bÝ�0ĭJe"O���O�(q��1��"%����"O�GN��ˬ��� 0n�v�0�"O8�*
ɍ>$���pB�^����"OJ��bA�*Ǌ�Y�.�!gѦ�8�"OL��3���D��	�Ѭ��z����"O~0G-�
Z_z�k7�'c��L��"O½p�f
�|n�&Ǌ(6����"O���� ,~�1B�%�%Kl~�"ONISc�ǌ'�\I2�T�,el�Q3"O�d���I���q�6Ώ�e����q"O�(;&�+F�L��+�r���c"O�����B%_��(�Ӓ9Z�ȣ"OTLK姕�X@l<1p�]�$Q��hB"O=ZR)�H-љ& 6ך0�B"O�E{��B<�y�% ��q9�"O��+�̗�T���oP�a1�"O��"�/#�2$�#j�<,cH�j0"O��Y�Ē�s���e	S�6���CD"O:,��-�f;8����=:*	�"OԴh�L(aӲ���fK+Y�p "O��Ҕ�7\Ř!SP�ұA:4�zu"Of�qTeY3\ވȀ5��0yΰ@+�"O��c�)WC��iJ�$Ū[����"OԄ��*�"�����#џ'�"X*�"Of��fe� �=Ec��#��p`�"O$Q@C��)=���\�)�V��t"O^��� L}�6��T�O�?���
�"O���M� Cl�c�"߭�<5�4"O��j ҫA��,���سkX�Xن"O�|yq(��"��}ȵ��?c��}��"OZT��ʘ{F�$��^��`�"O�̣э(��m�t�D�T�j\��"O�,�F�$��h2E�!V���"O�����?�P����']�`�ʗ"O�����F�a���B��@b�i
�"O }���?�Q)�I�C��!�"Of�@�"��~�6���I�F���0�"O�p�S/)8�6)9ba_�hNyJT"O�p;5j�+[� !)S`H���"Of��6&��D�qi<bE^� �"O�T�F�� +����H��Lx�"O�sB1S���0&V�%�B=I�"OF�2r	�2�V@a��Ϲ{��ದ"OB��A 
  ��   �  C  �  �  �*  _6  %B  �M  iY  'e  �p  @|  %�   �  ؗ  ۞  �  _�  ��  �  _�  ��  ��  ��  �  K�  ��  R�  ��  D�  � �  � Y �! ( 2 �8 +? <G �M \T �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�iӸT���_�6HF�Z��
/��A( �C-)l�	9�M����y��'�����"қy����g2-m��Z��'9�훑u*�f���̧ca���~�6DI�o�P�YfJ�z�����ND��?�*O��}2'�X.xȝ�����\����X�jƛ��!��'���nz�]8�"D�O���3CmX1'�̻%��՟����<a�O1�i��u����9o���3B��\;�슰�"����<���':$F{�O����>��&_*�xk��Y��y�S�t$�0�4�4T�<��f�5KQ.z��N����	��A���'8��?y��y�Y�ЫIX�cHp�s`䆵]�>L�p�6?1�T�q0�j�'T�����?�ѐpI�Q�Z�$s.qR�����D�<y�S��yB@�#�B�a4�Iy�Ą �y��l�ƽP3���b�4����T!�#^��rd���k�f!z�$�yB�'�2�'߸r��i����|��O�x!*�m�E]Z����gA�4HTb�IBy�O1��'��'��ݥk�, D���-��H�銙r�ɽ�M��"�?����?N~��JGX��7h�|l��q�V!{CҠ T��2ش?1��(��i� ��B��;.��q��ѭng^��$,��[>�w���~����:3��ɓl���S$��	-Ix��P)L�9=(T�I韬�IܟD�i>��'B�6-�<>���F�H���#��,ƚ@(V"�%����ɦm�?y!R�4�ش�&�}� � J"l2`sg 3ܼ;�n8f��6.?Y󎟺�*��#���}��]	%�� ����6�� 	0F��I�������h�	ڟl�IH��eq�i�@ۺ,o�	��*B�S�A��?���q�6-1��I��MCO>�T�������4�)�x(I��-N��'L�7-�Ӧ��b�x�on~��I�@;נ�'m*:�B�MO؜�� ���P�VQ�,i۴��4�`���O$��>N���fo	4˖LQ���h�����O �����V�'�r�'@RS>���D��1���]O��q�1?�7S�(�IƦ�RL>�O`C⇒TjZ�iQCǩ}��@���-6�<	ꇠU���d��֩�O�Ġ)O�ѐ�y����e�dDIW��W�,���O��d�O��)�<�u�i��	cŇ�F�RI�%�>����	�����?Yw�i��O�D�'K����DMfu���J.�}Q1E�W`\6�즭r6�\Ӧ��'@`�o^�?U������K�)��$�sH��%��	Ϧ��'2�'3��'��'���?.�ҘieȎ���s��G�1��4,��)/O��?���O�!nz�m�珄2j2����/\�`�Hq��?۴4ɧ�'�(�4�y2�9!�1��,��V|�5���y!�9�4U�I�\��	�M�.O�	�OBaj��V�=@����́�CF�ya5F�O^�d�O*���<��i����f�'��'���:g+ƣX!H"F��G{����dU}b�f��l��ē1���Y�ala�&V�@�������Q~�o��p�`�@�-��D�ںc6��Oxi�@[����㗬�D�l[U�py����?����?����h��^����1�x�ؐD��t������M�G��ϟ��	��M��w�n���;#�]�����DQ�'�6m���Q`ݴm�(�ݴ��$�zJ��'V�x5�F�%_�pW�K�a���1S��<�ҹi^�i>���Ɵ�I䟀�I�j���C���i���"�Ȗ�rTT�'�.7�M�e�r��O���1�9OT�a�.v��($DA�[������D}r�q��l�=��S�'m��|ad�Y5͠�!�ɒ�ZH�"�冤u��%�'�$�*�I̟4K�Q���ش��DD�E������@��l���N�8�8�$�O��d�O��4���<_����	w b�?�^�p�Q�������8�y$u���{�O��o��MKղi��}B�*�'�^P�`��cҬQ��ƛ1O�����L�#(�k�ղCN�OcP�=� d!�%Ȋ��2�� ��N�l@��?O��$�O`���O���OH����Ӊh�Xh@֊�i�QȐ��~���D�O���Ԧ�#�*�ݟ���ܟ�'���"*P1H%����(_0,p5H��K��M#.Oj�mZ3�M�'�@�ܴ����Z�`ٳ�ϙ3Z��G��y�j��qER=�?i���O���M�����'"�'��I�wa!C�f|��X+W�^����'vRX��Z�42Q�����?�������\e� �LM�I�Ҡ1��������?A�O��$l�Z8oZB�'Bq����H�lRs�� ؘa���v�8�W��a~��a�=���'o��Iğ杘}8� ���A�>�@�bЯ^�+��q�	���$�i>IQ-^A	�4�'Q~7͖;h6�q�ƨE�c�phUF�41tc�<�����?�(O�9mZ|�jT[��88r��4�Xyp8���4mɛ(ġzě���|K�-U�9>���~�qi�7H�%�A�ީr4*P(��K"��Y�����4���,����d�O`X�X%�,Yz�vO�,`�ĩ6m�����>_(���O��i��'M4˓�?ͻ:��dcF� �PX���x�+��iAj6��Ȧ)���O�x#��i���k���vm�4���	4��O��č0b�q�LSJʓ1Û�P���ޟj��O/R�L�C'�*`r6�xT	���Iϟ��	AyR|�L�o�O�d�O:��"
�0��5�ti�40T.�O�ʓ�?	�P�D��4Tϛf�rӀ�z0���paA;Br�\
 .	8@R��'���Ta[,
����Oͭ��n�$���?�0%Qg	x4�Sj�^y~Рw�N��?���?����?��	��\�ɹ�ztIc,�/X�0 �aE�b��ɘ�M3Ca_�?����?q����4��/U�`@փ�	~�i ��\���Ʀ1*ٴC؛�
մM������v!�<��t���Y�B(��wa6K�BR:�0�A��� �	��M++O�I�OP���O���O��)\���@I���TdC��<q��iA2���B�b�'����p;��'��M�%^�
�S���	=.9�g�RH�U��vHr�Rhm��H�B��l^O�Lhx��ͽUl.�&,�+ ^8u8���|PSmؼV�)�Iy"am��� kj@2�B�;f �\���ƨJ�d����?���?��|�/O>t�I2p���=^̱���H�U��rB�}�Ĉ�!�?��Z���I����4Q��BD Iz<��TiUjF���l�?�MK�O�m��P���J?e�Xw�IGp�x�FI�&*nxӢ�C��yr�'�2�'���'���Ӆ6Wؑѧ���MF��;�O�cP��d�O��릙��)�qyB�o��O���R���Vƪ���"�~�p�X�i�I�MÕ����眒N��&3OF� ��H)'Ģ(Q����Zl~�)���S�,���IZ��P���.}��Ryr�'R�'jb@Q�w�
�;��^�z'z�`���i%2�'[���M�6 ��<���?)(� ��vF6���G�0}iVH�7����+O ��e�v`'��'Kly�G�B�"��C����,�ʰD�k�(L�"��~�O��q��<~�'a�-³"�l	��C�ҹ\���$�'��'�R���O���Ms�āY ����9Q�*�:�L%�ƌ�'7M0��*���S�Ar ��"2�å���`�!
5b��M��i芁�Q�i���v0u�%�O��'#� AQ .e�\(P�mYmB�͓��d�O��d�O���O���|2��Ʒu\�$�5h�?0G�Ź񧜜j�����y"�'>"���'��6=�"Xq�W�$'�!S�]�_�U�D&J���͒O1����!q���I�s0���ą�Π�2+�:1N��ɿ�H���'�¬'�蔧���'�2������r�\0��4���'�R�'�"]�d�޴X+Y����?����5h�a˭b|`9��ƻ�C��<���?�M<)ck�?<x,�'�^ 8��:���k~RN�p���&c[0Y-�Oj���I5Yd"	2m 4��Bk@��d�#�i�K�"�'�r�'���(
7�M;z���s�[�6U��JQ��\�ݴL�$����?�q�i��O�N��3%Ba�Ei${�E�Ȉ^~�$������M��m�M��O�I����S���QŐ���ԕOp�ac���C�z�O���?	���?����?��Rqa��P�*�1���H2�),O&�o����T�����j�s�Q�	�=}�p�R��pk�����N=����Ԧ�*���ŞK�\+BMïzm�Xfo��U�������-O�u�P��?�0�>���<AF�Ϩu��7�<q�|9��j��?!���?Q��?�'��$���	ccm��dƇՐu80���;UlX��럐�4��'Jʓ�?1���M���W?N82.R��2�(p�	�#ڀհ�4��d�!_,������������� c���%Ɂh��,	�Ɓ�'��'��''��'h�P���Qd�(8�!t�a�R��O���O� o�u���|.�� ��4��$��hN�u°�й+��O\o�
�?�(��lZs~b.�� 7^8XsIA"�Ju�e�՘~��"Ɵ�!b�|�R�\���T�	̟p�`��^ٞq2��W4_���x��ޟ��Ioy�`y�\`�B��Op�D�Oz�'`�z����)+����ذ\���'�Z�l�*�O$O����`<I��ц{�$x���h��8G��<)���G
�7z�z������O�U�K>�c2#�JG`�7Rp� .���?!���?���?�|:)O�Hn�?af�	1���_خ$��C�!H���vCV[y�F~�
�d��Oao�m�h�
�D�x�n�1�
�J�.$�޴�?q!�_��Mc�'�"*D�}��y�-��� �I�ƿE4�ݪ��*cB�!0Obʓ�?a��?����?Q�����-��\�sH�'���7%����oڢz*��'a��)�¦睙V�$릆_V3"����F����{�4"ߛf�'��)�әY�Dm��<)@ON~�N�%A�D�{���<ɧ(֭@X�dW?����4����җH��M�#�I(t�VE0o�%;���D�O���O�˓\����/f�"�'��@g%��"�؆W�:��fO�V�?	�S��ڴ=����' ��*_Jt������"SBߴy���-(N��@o�#W����|�q��O��S��?�J�C���qH ��%��¶T����?q���?9��h���dZ��~�������� vI.���@�qړ%VSy2�m���]�YO�y�7��~z
q�'O�	����M�ǿiJ�OG��v��<q����de�\�FI��g�����ae��]F�T&�������'���'Z��'L�0jpjўVf�-�Y�Ԛ���ݦ�S�J؟����%?�ɬV'.ْ�Ә���4�[vd�X�O�l��Ms���>���,�N�Z(8�C��P�T,�¡\.MZ��d/&?q�E�O�*��]������F�
|Ke�#n#�l��L�v� ���O���O��4�,ʓ!��)��y2�E#��uhZ� �5
��y�i~�㟨��O��m��M�Ӳi>ΐ�����"_d �'T$m����	xț���h�� �3,���i��^�����t��K�톰^�Z���>O����O��d�O��d�Oj�?9)"lY�N4�M],&H,�W}��	�BشJj���'}�6M0�ā<\��D8`@��w�4��59�
�'�h�4՛�OX����i��Iy���'���v��䇙�f�-b�Qq���{�	Ey�O'��'�Nޑc���</94��ҡ9���'9���M;�G�q~�')�S�>s��9��N�Cpj�+E�U�c���t��I��M��iqLO��#O��I��
�P��SF�ԋ];�p0��(;����#?ͧGwV��ԇ��>��ñ���)G�yЂ�҉O�"�H��?1���?Y�S�'����?Miڈu����F��8��r��
�˓d����$�l}�Ns�j@z+�r�9r�L�dߞ�֥�䟸lZ8eܘ�l�p~R�E&9��ӱo��	n�#BJ@�|} `�[ -���py��'�R�'���'("[>A#g�S�L+���|ɤ�'!��M��&K��?���?YJ~�'盞w������:d*�jV;^�� �{�����e�)擉G��m�<����h���!*�Z�&��ˇ�<���̀�L���+�䓔�d�O��d1(�b��1B"���I�?�2���O��D�Oʓ["��C�V��'�bF_9 ���K��L��X��Сx`�O~�'-�7͍� %�pz��Ead��Bϫ$)*���8?2F�\�� �	�6��Q���䏶�?)��2U�� ⭝�|Ip���Ջ�?���?Q���?�����O�4�&��+[�%S4�Պ2r$ԃ�!�O��oچ҄���ğh[�4���y�Β�:�Nh� ҆ڤ|c�Ō+�y��dӄL�	Ԧٸca�ڦ��'ޠ\aSdL�?u��*���и���	���aD#i��'��I����	ޟt��ܟH�ii���?�v9�נ�6]~����<A��ie����')r�'��O+b�'q�,q!1��}�Z�0)��-6b�	�v��O�O1����m!a��*��<&>p�2�	~@j6Ϲ<����+m��Dؼ�����٣s~���C��W�|؉�n¾(���$�O��D�O��4��ʓ2��*Fd�2�i�p��L�#uRl)�#��y"�wӐ��­O��n��?��4w<@��:��XS ��B���P"�M�Mc�O��⅜�:�'����T��6F��������d��0O��D�O`���Ox���O��?�@�G�#F� J�{QыS؟L�Iϟp�ݴN��u�O�7m#�D�PDn�#@�;{( ��G�`6t%���4T��O��0���ig��-!;��؆h��O;T��A����D(`�@l�CK�IIy�O���'	d�xov,��f����k��K2�'"剣�MK���?	���?�-�z�s�C�+\�!�,�~خ�U���q�O.nZ��?�L<ͧ�J�2=��3%*���BT&��\� "��06Q�Ѳ-Of�i��?�F�?��U�+V	 !@�c��+@��]S
���OT��OH���<��irjB�$�h4h���B"���A!I ���'��7�$�	���i�.D�3��'l��"&'̬lv�z�aŦ�ܴl�Q�4�yr�'�81c#���?5��[�S%�V#T��%�
�DM�P�Ghc�d�'q��'�B�'���'Y�,�@q�� LLq ���X��c�,ţaD�O����O��ɶ|Γ�?�;.gH�	������6�K�p�z��0�i��$�>	��|�����S럹�M��'q� ��˷�P�Y�ł�j���'M��(�͕ڟx�v�|�]�X��֟�� &�I��t�ȼK�j!n�����Iß`��tyb�z�ZP��O����Od���hͼ��IR���"t����&��2��d���e�����-�Z���K�~}<� � �w����?i��͌�\C���d��n�C��>��Dmc�4ڣO�!t���E���@�$�O����O��d+ڧ�?��JU$OT��X1�ȘY&,a���?y�i�,	s�'mB�u�Z����d<��*ñ(`��0.�!UVf�Iަ5�ڴ�6�Mʛ�2O��$��	�0���L2�  ���Q)C��P"�����J)�D�<Y���?Q���?���?��DÙzАPcR:F 楫�+���$Wݦq+f]ܟ�����8&?���.rkd���Bр3�l�B4-��sb�(�O��m���?!O<ͧ�b�'4!
-	Pf�scr��6I^>^D��㨏Ge~�q-Ot����?Y��<���<�R���sބ;gJ��_1�	�pi���?����?I��?�'��DSݦ!�be��<q&m��S�)%%J�k�~�kW�z�4�ٴ��'�j�rԛ���O�7ԗ�x�€ͣ-?H��b� a��g�eӨ������"C��,;��YIyr�O�G ܶ@��������Y8�fO��yR�'�2�'{��'�R�)-0zx)��ʬW! 噃iQ-)�Z���O���VϦ]�sas>��ɹ�M�M>��ǓK����2O\�A�bߩ|��'�6mX˦)��i�.o�<A����=��
�}ڨ:AhϺ>(��Q���+@���H!������O��$�O �DЩ�"t(��{mtزF��E�r�D�O��n��̄@��'1B^>� �R�P]^QL'i�XԐ'�$?!�]�T�ߴcf��l4�?m0�
�I�Zh�v�	6X�xa��s2 ,� E
l}���|�T��O�HIH>�,њ`��k �^�7$�Ay�'Ɂ�?Y���?	���?�|�+O�,n��C���#D/۫v���`A�/M��1�Ϟy��c�n㟬ɨOlZUl$���G�
2-Z|�Rh��uΕ@ݴכ�k<$̛v����N��3*���~z��S�Z��]����2�v	���<�-O����Of�D�O��$�O�ʧ��ko�t!��<K�%3��i�~����'��'2�Obb|��n 9���7��<K�9�)��J�ƕo��Mkx��T�SAU�8O*1�S�[@i"w!Nx�*7O��ؐf���?��g*��<�'�?���ɣA�Va�5�F@�� �?���?������Ҧ����_yr�'W��$��A�~���`+=�89�����f}"�aӲ�l��ē����"�A�]� �,��T9J��'&��r��_<r�`����џ�`��'���Y��,0�&t�V�VPƤ��7�'��'���'��>����gl�$X1�H�g��1���cƥ�	��M+���:�?	�)ɛ��4�F�R�H�A�@�<_��s�3O��lZ>�?9�4Lf��ٴ����D_����'?�<���Ʊk`�rgG�N��ru�*�ĩ<����?!���?����?Q����C��!&y�O
��d�Ʀ�"g���t��ß<'?�I�p��i�[L�$�!��rK�u�O��nZ��?1O<ͧ����I���ւLZ���#� >m� +b�$�@]�.O��Q�엉�?�u3�d�<9r�Kh���'#��g���JgCK��?9��?y��?�'���Y����П�D���zD�a�¤�7��V#����ߴ��'����?���M���u�XKgKB�P�t���`F�,�۴�yR�'/,�b��?�
Z������E�F�еPZ���R�Z��Q�ѭ~�X�	ğ(����	����J��'K����0m�<&�h��
��?���?�ôi�I��O��z���O&��U���$�H�*��E[.���n�k��;�M�g�i%�+�^��f<O~��B+#Eƕ1��]0TBmP]ufy�b.��?qE!*���<����?)���?`jO�#b|�J��9��y�3�?�����S���Wߟ|�Iޟ��ON��Wj�
�@����������O��'o�7�U���$��'g��qd��/w���G��%K�@ց�U v�N���4�b@���0��O�$��L��" :�*A(��\$��O����Of���O1�.�9M�)]�%�Ri�u损|�R|�#胺z���R��'e��e�㟨J�O
�m�$3��A�NǖB�=�2�`��YPڴ0���LУu�Ɩ��Q4G�C ���~B�AֆQ��xS��k�˒��<���?����?���?����?1�⚐3��N#�,� �@B+ir\���-՚t�y�����?���?��i��'�2^��N�K?�K�CM�Z3<\1��H�?��426�U"��Y��y*���d�-S��7mk� ��k�q#ݨԩD�J{�a|��W�PK�"��@�	Ey�OG�dܯ)�:ap�$9 ��ji��'k��'*�I��M;����<I��?��lť"�HK�ܞO��bT	���'<��BǛ�Hh�x8%�����,��x��@�02�H�?<�'m�B�5�JT��,�7��埲���h�
��Φ@��8
�zP.lA��Y-Ӣ��O����O���*ڧ�?Y�ẺeJ���͝�(r�Ip�,�?��iw���&�'��k����]
^q�I��@�0�d�2/�J"��ğ�m��M�d��MK�O�A� �%��SMU%\	��+�7�:��*^UWV�O<��|B���?���?a�I�*Պ ̅�3�b��Ǭޥ{=|=�-O��n�&�,��I�h�	X�s���yp�(Ku��d��P������D��aY�4np���O�Ji�'�L�`Q�5�*>΄� �#+ ��*�O�	CE����?AU(;��<�SF�5�0�!)�'�j(Au�;�?I��?A��?�'��d��ө�ޟp�ZV�lk��lұ�cC6�<��^����?9�]��pٴmۛfAj�pɡ�ÖC�^|��&2�M!��
Y�~7|�X�	�	�d��3�O������;:N&h����*��� ��C=9�DUΓ�?����?����?�����O�
812�N�G��y!��H��O����I`d,?	�i!�'�̭�d挺DdH{X{3dPK������,��Fm��)X�k�7m"?�d�g�? �������<� � �@��v��;��?��- �$�<�'�?����?�%�+#Z���򂀾E��0��͜ �?a�����!���ڟ�	��t�OT�����Z�d�p��ϟ1W�T@�O���'��6�Z�%��R�����d\�9�b,;F������.W����ĵ��4��D����̓O�d�'D؉��!sN���U&�O��d�O����O1��ʓÛ�Ǆ�-ޔ ��B�]�fRbG#���Ң�'(2�v���L��O�o�:|x����i�3)��t1*C�En(���M����M+�OpX@������<!��׎mEl��!6g������<�.O��D�O~���O����O��')�H!�.�
�y)`	
�xn&s�i�R�QA�'��'Y�Om��'-V%2���aO�帠ϟ�N���o�"�?9H<�|:�!?�MS�'H���F'׺@Ä�W�v@ !��'m����l��k��|�\� �	˟ ��ፊ}".�9S!�n\�(H�F�֟�	؟���Ey�wӀ���G�O&��OR���ND�F�.5��� "x�#�%�I(��DP��H��ē�&i��h�TȊ�JS�e����'��� 5M��oȹѳ��������#�'���1O	h�T��牌�S;�j��'���'��'��>��r\��Qb�5�ι@B�Қ7yB����M����9�?Q�&㛆�4�vU��E�b�dę׃:,�r:O4=m��?Y�4Ns�4�ش��D�:,����w]p��a��WD�|�"�-���S/.���<���?A��?����?ys��>:!�[G�8)vb���O�6��_ͦ	�E�My��'��O^2B�)Oxpn�bd�� "b�h�h�#��F�O`O1�t���k���uz�/�>R^2�ܮ`!�����<I�J~����:����d2h�t�P���#m�b��������O����O��4���#w��А'��^�^:����!8{������ry�jcӰ�p�Ovho���?��44���"c[�[��	�����$;&@��M+�OX�˗��$�z��?����
*�e�B��.�5av��V;O����O����On���O&�?��b��z��h���sG��ٟ@��ɟd�۴l+"��'�?ᴶi[�'H|{p!��1�pj�H�$�9+��!���O���O��Ԋ�i���/���͘==�X<���Q�hTr(�߼�����䓙���O>�$�O���r�+.�e�1���e��ǟ��I~yr#i��
E��O���Oʧi��8@��'��i1.��T�d�'��d�6k�OO�S"e�މR1m�4t9���r���m�n<R�] ���AׂX}y�O��Ib��'�B@����"�٢��~���v�'R�'�����O��ɼ�M@FXOA���$�R=$�nU���Y<u���,O�oZD��!�����MKe��5��P��\5C�JM��o�Rb�i�2d ײiO�IK���%�O��|�'�ީaOS�X�|����U�&��K�'���8�I�`�����Ic����rX$9DI�B $���T#�6��+�.���O�d"���Or�mzޅ�B��/@�|Q��Қ^n� �N �M�յiW�O1��,K�Cp���IZ2����K��48tL�<Z��.>D���p�'ʹ�'�������'�2	�3n��M���LR�if�'\"�'lbV��!�4qL��z��?i��r�}�rhU�r�����oڃ	��`�2
�<!��M˱�x�%H\�b!O��w� c�ֽ��䞤2-�p;deK�~#1��|��{#��$ǸP�v��ƕ4^�4��A�žN�(�d�O�D�O �$"ڧ�?)4�>j3@Qb7%\\(ma��?w�i������'#R�l����'X<x� ����w�h�0*�H4Z�I��M��i� 6�W�`6$?�G�h�f��	�ѩ�B�
�+��٩%���I>1)O�i�Od��O���O�P����;OO�r�ܪ
��A�	�<ҾiHĸ���O���.�9OZ����Խ>I�5���Ӱk*�Б���X}R�y��o���|"����Ƥ� Lv����2Ԓ���T�n���a!V[~�]��y�ɮ6"�'���R�nlI���f�:ADGB�_��H�	ş$�I��i>�':�7�hf����%y��g�N��a󪚀h�������i�?9�_�h2ڴJB�i*�`�j˖ Wb�1(մM3�	tK��b�֑��`�(��	5��$�G��߁�c�'%��0��u4aC�ko�|����������I�T�����+�,,�����:bHQ�`g��?����?qb�i�dY�˟�8l�џ��'��I� ϕ�b$���B�A��ъ �8�dĦ9ߴ�����MK�'#Bʘ?��h������
�8� 8�P�Jϟ8z�|R�|����Ο���GN= m`G�[d�C��<��Syb�dӴ��1g�<����i��S����eP�5���8.@�Ɍ�������������|���?��(�4�$�a�ʷx��qa�-P	4ƶ�Ѧ�����D�� k�	?D�O�)�0�U�?������Y5Uh�H!q�O��$�O���O1���a�V��>W����e�\�9C���Fm��z%�'YR'pӚ�;�OZohن�YuI�]��@M�n�1��4%��6�'n��f?O�D�3J�����b��w����� �:0O6�1V�ٴ�r�ϓ����O|���O��d�O����|��2DJ⬒��ښ7�dJ��6A���U��'bR���'�r7=�8	�bO�9r�$LD�w\�<�p�[�	*����|��'�JQ���M۞�� �Y[tfT�CɈh5인Y����;OJ��l7�?9�*2�D�<���?�D�^4%�Q�e+K2t:��H(�?���?!����d���I�f���X��� � ��D%:'��H�)���`�2�	+�MKS�i�S���B��99=��0(�G;�Yi��p�x���𨳐Cи%2�bV��Oxdj�L���BWƎ&�t\㥍C�=������?����?���h�>�$U7{��80 �ZbĜȠ�K44�@�ČҦ%���8?ɰ�in�O�.
�4I8�AvA�.����*^�?�ܦ�!�4;e��-J-%�V5O���I+�����'3I�h�C޶sp��)A W�u���ʷ*���<�'�?����?����?	P/IY�!���@$���[4C����$Dߦ���c|�`���X$?�	���J�ٸ|V�au''1�3��D�O^7��X�韼�	���-S��)p(���Ɯ6���͜oؾ��P��d��&�9��FN�IQyre��G9
̃4��halLq7�WlR�'T��'��O�I�M#F�ƫ�?7%�g��`3��]�wʂ�@��?��i�O���'��7m���Dm�^V���Q�D@s��őp����	
9t�7�%?��%���I��ҘϿ��-�i�m����Us�BV
��<����?���?Y��?)�����[1vAٲ�@y�fԈƥ��$HB�'��n� R�4�l�dM���&�t�T�����"G����u���A'��!��O�O��k�0^�f��d���֘5#�$9PNL0�zEp��� G���q��'�� &��'���'4b�'�(\�A∂8���,g����'�P�Tbܴ2ޞ��(O�ĵ|��$�E��}z�
A��N�8i�~�!�>90�iښ�3�?�"`N�y�TlP�9����(n�tx���H�>喧�t@I����|bn�{`dS�NL�7�rh)!�W�c���'�R�'c��4]�T�ߴl�$�����>DTh(@7e�:�|��taʪ��dJզ��?7U����4)d���+��0ًCJʳ*ઉ�U�i�x7�_�U7m:?��K���>�	+�Ԡ����Q��t��udX��y�]����֟������I����O�P8���U�Z[ވi��[��C�mӬ��G�O��$�O�����DH���݃@N6p�pE@�W����e���$���4>���5��	ɓ}��7�s� �S$n�XmHB.�7�6I�p�P�ƁU %��i�D�@y�O/X�)����O ?F>�x4o�1<�R�'���'�剩�Mk2���?a���?���� ��Y��\o>�Ec��H���'��� ���gӬ�$�؁�/��Y��H[q�<E0@It� ���l(hK+�|������O(���D��3w,V?6����/[�BՒ���?����?a���h��ė&%w�M��<t_�RV�[�C�\�d���=���KUy�sӌ��]�ecέXcK��W~p11�@�a�b���M��iS2Q8~�����X1Q��0`���眠a�J]�ri�2�>@����5WuF&�P����'52�'�R�'�Q�4��t쀰u���q[؉X]���ٴ�f�����?�����'�?�D��
|��+Rk��Y���C��"�I��M���'����O�� �e*�l@�e�i࢜HfKZ6��B�_���r-�*j�
l�	jyb*CV{��kU�×[���T�X�y�����\��̟�[yBxӞ9� O�OjP6L܏���8 ��er��>O��l�S��t?�	�M���'�L�=_p�;F�Ĺr"A�1G�	l��0!�i�����e{U�O�&?	���K85�F�L	[ڎ��@�=��	ß�������Iʟl���Oc�\;�mI�$f�I��J%W�0��s�'���'� 6�xp��kț��|�b��۪lb�O�!vP����*2+O,�l�*�?��7���n�W~�b��a�R	�CKZ�!ĩ��PRTq�G�ӟt0$�|�W��	��	؟�3��՜`=`����0qS�I����Ify�Ge��0����O4�$�O��'J(�X
�V:�L�!�3k�u�'��Si�FE�O�O�S�C��T�탚wq�yQ�ǂ�rw"�8����z�ǘEy�Ok>��Ic_�'�|(V`�q�V�%��0
!n��'��',b�O:�0�M�瀋�Tb��U*"�(9�p��7��P��?���i�O�p�'��7m���Qk״o�B��f�<���O�7���6M#?�2/U-Q֠�隁���x�ɻ% �@�N��`�<f8�D�<1��?��?���?A/����I��bܩ)d(طG���!]��D�C���	՟l'?�ɻ�MϻV�x�Ԃ�'��H�!oT�R�d�h��i�^6��|�)�l��m��<I�h�
\C@�^��&)��<Iq��5	��$��䓈�4�����L8Lx8E Y1,�Ęh�T�/K����O��D�Ov˓Z�F�H�zA��'Cǂ�i��p6��,s�h��$b��s�O$U�'��6m�ۦ1�M<��̥k�܄p`��Dd�DOZA~� .zE�}�t����O_�a���1�Nų\�]���i�x��[����'��'�2����J�n��L�p	9���43�`�Q�^��4ufr�.O<nZK�Ӽ��T���*���+c� ���<A6�i��6͙����&�DĦu�'ˤAB�A�?�
b�K#��y[����R� P� $� 1�'��i>�����T�	ן���;�vQ��$E	jpH���� >��ȗ' 7�G�V]�d�O>��$�9O���⥖�aD0p�B��it��`��[}"�aӴlm����S�'O�L�� <i�5H����|+%@Y�<�ZH
�)�Y��ɳ ��݈d�'�>�%�Д'p*@;��({>j�H�՚8BE$�'A�'�b���U�|K�4}  ��8,��@g��a��I�!��:~��͓)0���d�M}�ijӪ�m�M�%���+�(�0��ݸSJ1���k޴��DN�P\P���øO�wNqe�X+F)�Ir� ��a��yB�'�R�'0�'O2�IͬW��$�6e��:h�NZ!Y`���O����Yr/l>e��6�MsI>��DY� �!��G��ZE�\�{H�'�r7m��I�	;Z7-3?��DʄLR��w���I��'��� ���O0�J>(O����O����O�}�V�X7d��l�r�Z .Ŭ�2s��O���<)��i۴D"��'D��'���U/ݜu���хL�M�a��I=�M��'�������0Q�a�cA�O�B������D	�E��(%�5[d)�<�'x����%��Kt�����=NZ�l�H�r������?���?��Ş���֦�pDС&iQ6Ĝ�tTb���훲b�'�7�=�I���DE�EA2쏕�`y�3&��\�6�Se�=�M��ir刖�i��$�O�h����ڴI�<�Vl��]�B��&��3E�iZ����<�-O���O����O����Of�'&W��X%� ������X�h��3�i/.dKB�'���'M�O�@u��΋�'|��t.U�n��a#����,�|�l��?�H<�'���'H��H��4�y"f��Hs��@H�w����f��yRG������k%�'��	ɟ8���/xv ��J�=L��@�Y*]���	ٟ`��ş̖'Wv6����&�D�OP���1t!x��������P$`�>����O4,l��?�O<q�FK)[���h0J�2v?t���D��<���4)� Z�9NL�3/Op�)��?�q��O���s� �Q*Ď3e��;�Oz���O8��Oꓟ�ä	U���ښg��Pb�]�k&�R�o�)^ˈ���uDMğ����	gy��y��Z�q��K���4Z�
�
�*��y���^�n���)�ܦ��'�
��H��?�"ލ"�t(�7+Z��Ha����.a!�'��i>��័�������"'�ܱz@NM*LaN(ТJ+^�@�'��7���:TR���ON��5���O,\��\4z�D�3�^�&S��T�Tty"�'|J~�`�A�M���%�;\@1������ݣB+����d�3;����O�˓d ����:g��TI����d�VLY��?����?���|�,O0�o�32s����6|؀��g\�C�5�ca �Xǆl��6�M��F�>i��i�d�D�v�s�g�e���P+�+ڐ��ь�ze�7�2?a�BW3Q������ܿ���WD��Ř���.p�ȓ`�N�<I���?���?1���?!���@��p����0�K	[Q2ؓ"�,R�'�B�k���@�5�H�d֦�%����d�8P��ӿHy�q�5��ē���k�O��d"E����w(h�̌`6�(hEN��sg��f쪶�'� �'��'���'K��'�H��f��x�T��3�W�
}q�'�B]��
�46�nm���?A����Q�D��pb�� ��i�#��I�����������S�dj�)7�p̉��Ƿ3װa�R�A�`���pc�R0N|@��Y��S#H>�m�u�	���F4]v�(���]K~��I՟L������)�sy2-m���)��ÿD�Ix�� 8�uW��>�2�^���x}B�u�����:��E����F-`�S���ܟPm5K��oZL~2�
�KĨA�Ӡx�ɟ����S&X��Z1BŘ[X��	`y2�'}��'���'�"U> 2
ڴN���k̆692��E��M;F![�<����?)H~�9t��w�0�+��`�M�b,��<��mc�2�n���S�'D�ta(�4�y�_3�T`��KT܅Cp#��yb�K�&ZQ��;6�'�i>��	`�`�x�d��6�X#
޴+٨�����Iß��'9�7-�-]����O��䑗Q���A�ml�ja�ԍo'�P��O�m���M��xb��M0N�"eѡ/��1i�Չ�y"�'eM��8kZ���O���?�?9���O(����
�o|�Q��R�e�l32h�O<�$�O���O��}���+t�}�@�2s8th�d]�� ��#�> r�'��6$�iލ�$� D�Ȁ[���L�P
e�r��P�4@ɛ�os���P0�vӺ�	�$�$�&Q��$�Pv��A�?46����R'��%� �����'���'�R�'� �+f�m���h���BX`�!]���ݴ(z����?i����'�?i4[=T���:��%7����-����ɹ�Ms%�'߉����O���X��pi1*ȣ5�ɹ���8:$���B�	��剳"��0V�'\b�&��'�"�pR����7�.����'qR�'������V���޴%O�;�bך��VJ�&�҅�`�Y$��3��7��v��[i}bCh�&��	��MS�F}���{!m��0�lEb��ɢ1l|�n�x~r�Y&�X��ӻ��O�+�d"��ցBa՛#�^�fL��Ot��O����O�� ���d<�7̒M"nY0�f�P�� ��	�M�`���|J��}��V�|���@��a:W�ǗK�����M��O�l��?�SO�v1l�b~ҋ�=@@0�"�ͽ~i�T�����'>d���蟌��|�U����ʟ���ޟHx��_�j�2,,��2��ɣ���ß`�	dyr�^��Џ�O,�$�O��'i۾�B�C�2��$�@ܯ#���'Ք�l'�&��OzO�3� 2��!Ĵn����\;5����㓊W��A�C/;�P��|�s$�O� O>��j��%�r��.۱S���R'g���?���?����?�|:,OԤoZ�$��*�Z|>�i�nݱn�D���HßD�I�&�#�R��>�u�ih�p�3ǜ"�ly��m��$m��O�7��>g�6'#?�SN�k���C������D�k~�b�[�m��$�<q��?���?I���?�,���*<+pb]�@f�_,�<P�Gɦ�s!�쟼�Iџ$?�����M�;4��8ɇ�̫\x�h	�lށ�N�Av�iYT7-�^�)��\���oZ�<qρ����҄�:5s^�l��<Q��X�/Nf��T��䓭�4�6���.B�li�#ض<��+1��8�~���O��D�O,�?����q��	�Z/�E:6�
�i"�Є��`��[��	
�M� �'G�' ��h�L�:F�*D�&#�$7:j���O�U���8M�ո-�I�?$�On�
[v��F�D
h��I��S>B���'���'�B�s�a�qB�y��8�h��D@ -<�ݴi�)s,OP�lZB�Ӽ�g֊*��TY��۱@L�庇�<�f�i��7��O��	�o�n�EL�᪶��T���/߼�i2N�� �bЁֆ����4��$�O$��O��$��fyi�����6?6%At^�vp�N�6��7;���'����'�R���U*B�
-�Ә9���>�v�i�<7M�O��F�t T�=w��X�K�{��E��9Q$�Ä*؉��$
&fr�D��w>�O����$R�S�9X��V(C=o�����?����?���|b)O�o�f����	1`J
�tŔ����0�R�a.批�M��b��<���M[�Tc�<af�]�X@ʭ�gJ�"�l�/��M�O��@�����w�X��eHBl`иJ�E�,�2�'���'��'���'%����n�����f�=.��x���O�D�OBplڌC���':V7$�$V�\�ED
� ��բ��k�|��<��i��7=�ȹy�`h�*�Zi\8��L�0�0�Ҫ� �JIh�!��(ɸ�$�1����4�0��O��
5*
}ɕB�("u���ǏÐ@�j�$�O�ʓǊ�?9��?�(�H|s���[7��R"r�ȤJb�����O��n��M��4����0S$�*zO�2t�Dh����e:D��z ��O[�i>)���'���$���Sl�}`��r�iʲ'TXP����㟰�	埰��ğb>��'�~6�_	o��q��۠n%���`��>(R�Ʃ<�ǳi��O���'o7�V"#��,q�)�;	���-�,�Gq������B~6-#?��ۦ1��	%���)`�t�3�K���r�*�y�\���џ����� ��ȟДO�� ���=H��Ē�o�7�
) �gӀ�)�O��$�O���$��睥=�h�̀<�Xa��m��� ���4?���'�)擰d��m�<��H�:����mA,'��s�kY�<��Cۯ��������4����_��ʇ,�X� � v��S6D�$�O����O��=��VIƹK��@I@$��@��3a͂�8E&�h��VU��C�����lZǟ�'�P��йv��5j�h޹�LS�O e�����+��Qf�G��?�f��O(�1�a�0,�t|��̢a`�B���O,�d�Oj�$�O��}���L!hA� U"iWܵ��AI=q:��I�^I2���$�ɦ��?�;4H��0�F�k�Vѩ���ʰ��O���pӴ��KY�7M&?�i�;y� �)�^ ���d�؄R��aw"�!K�p�M>i/O�I�O��D�O��d�O\A��a�9���V�U0_z�}�W�<�ҿiOƠ�3_�,��X��
�h�pl��4̸M���`�T���P�4��ߦ=��m~J~*A�;�^�9��\����07K�(�t]��ˆ_~2n�0s<���?��'r剅��R�!Y l�^�J!;��%����d�	���i>��'��6���{�(�D��){���	�{��Y��D]7!���ۦ%�?�V�\��4ܛV�'�\�jT�2
��薭 ]���RG�{�����`��#�V���9�p��lI�R��E#P�2D����3O��$�O����O��D�OP�?��'�Y!^�r4x`��hq����Iǟ� �4�x@-Oz%l�I�R?�1�F
 -�nmBG+��Icy�G}Ә(lz>1��LA����'OH� ��th3���:e^��KՎ�	��x��0s��'��i>��ퟔ�	�8�YOK�=*R䀠�U
���IڟЕ'�6�!7����OR���|���7I`,v�*����C�w~'�>���iV�7��O��~���!34P�����ą��N���l����;��������';��2�gۥ
"XH�T��M�'�Y�w��ZQLӋy
�}"'.�g���ئثш�ye�1^�>��TL�E��[��|Rn��|
���̅धB���O�J��HQLhpc�ҝ�J�KǄĸXBޤ)@ə/�A06!\��}k�gK��ĉ��ci�H`"��߲Ljn���̒Hn�q�

;h�&��g`D ?�:�����6}T�q(���1�^��,�E�ݳ���(� �#nW*+���)�I�!RC�9�GA���QCA��5l�� 4�O�@Y��:D�7Z$��ZC��>�*OJ��0���OH����^�>-��Z� ;d��W#8XÀ�3���O\��O�ʓg֬��W=��tKw�{ �S�@O�Zഅ�D�i����X&�\�����TCQg?�!M4vhT	��F�$sQB@n}��'�b�'剶3ذ�y���M�O<8�:R�S3�*��+��j�nZǟ�&��	ǟ�#l�d�S�? l	�m:�J��K��I��R�iF��'�剥SO��Ү�����O���O�y^�\�G
�9�Lm��٢G*Z\&���I�j�OCS����)�	!��[D��:�M��e�3�M3)OV��H�ܦ���ȟ����?���Ok��p�1�BL�^�pQ(������'��h�4�O|�>�ǉ	�(;���#H#i2r|ЍqӸ���������͟p�	�?y!�OfʓVLK�-yޤy!F�4\I�e�MS��Y�?&mYT~2�	�O�l��)JLv�E�F��lňQ����ϟ����	  ��Otʓ�?�'@�P`�蕍	^r��[�pm"'��̦��f*?	�/��w2�O���'�R�Ō�z�{ū:(��$Z�ꚯ/7V6M�O�}� ��^}"S�4��Iy�Լ�Ī�,�R$b���h*�Q���G}���,n�'���'wBY�4q�G���<4�J�"�$�s�.5�$X��O�ʓ�?�I>I��?	Fb�7S��a���>4�Q��e O��
M>q��?������ ���'+�0����w�*0H-�S�ao�@yB�'��'�R�'N���O$]�R�ǭ�l����߃ 98e��U�$��ԟ���Oy���3X�>�'�?�R)J�Nɚ�x���&,�"�+�`�	M:���'l�'���'�h���'��1®O�ˀn_�/n��!�9j���i.��'��	6f��[O|B�����@H7'
�L�LA��ӛ<�N8$���'��M���'|�O$���1%��BA����[�D�-Y$�6V���g]�M�DR?����?eK�O&!1d��	k`)�bN�ըE�տiG�ɩ(��5�����'�򩶟T�̍c�`q�gC�`�N��s�l,
g�̦Y�I����?!�I<�'gnRy�@&U�Xi����J�B �J��i��'1B�|ʟ�d�O��Y�I'��1B�]�ū���ܦ���\��

��K<�'�?a�'�Ƞ!!���z��2q�V8��P#۴�?�N>�GV?���iZ8�����VH�QC@(a �O�zc��<�*O����ȍ_����cF�.�Hd���3 ��<�����O�����$FF�	�aӀ;Ǆ|k��NBظ˓�?����'Ur�OJ��)�B�4��p�ƚ&�`��i��+�y��'��	ǟtBv�_h�UA�(Y8M�QG�5"��wn�Φ���⟌�?Y���P1$�&�A1�,�2���k������	���?�*O���B�N�'�?Q���Tc�`*F�Aq�1"6J�)s�����O��>��%��b-7LQ��W��fu��j����<���`XJE�.���d�O�����U�3G� �������-�h}@�x��'[�	!F5�#<��!q���d���!�h�j��Û'JH�l�]y�,��7��6m�O�T�'u�4�-?�/��b��X���S���d)�ɦ��'�B�':L�������=���򋛕k�IC���M�	^�ZR���'�B�'9��%*�4���a�$�/0ǀ82p��6)z�HEA���۟`�	o�)Γ�?��+
r������6P�����bś��'x�'襃��8�4���ĥ�,��OF���$��悰v@�ԛ�yӦ��4��s��'W2�'a�OƟ{q%C�'W  ,�a�@���7�O�iۖ �D}�[����|y���5f�і~��A���Ɠ�yؤ����DA�r�$�O��D�O&���O0ʓE�"5P�ă��H+�`O
5��p��d)I�Icyb�'A�	㟬��ݟ���*�5-<M���(�
��f��k �I����	����	ßP�'�x��@�e>���d��O�j��E��8s�51)bӌʓ�?!(O��$�O��d�^�ȼrd �p�ՒKc����1.B�}m�̟P����|�Iry�E31���?�1Ul&e列(
0���b��-pb�l�����'�'�"���yrP�00G���1�~d梇�US���O&�	��'[�����~B��?Y�'#cj�����U�� ���N�`0R����П����0"���'���S�6�4���*�!$2�1�nM%\��V���r���M{��?�����^��ݖJ�.�9�f�<R�Nh��J[9+�@7�O������:OP���yb��U	��T���>iN�8v��0����
OX6��O����O����K}r\���J��1۶�2L��*(!�d��;�M�b��<yK>)��T�'���ru�M�]��e;�Ȗ:�-��zӢ�D�O<�D�]�2P�'���ڟ(��z��p���>��N)^do����'t�j�����O��D�O�`�KS"&��DG�<Mpp!eF����ɈP���K�O���?I/O������e�����ȿv�L��d]��Rh���'5��'��^�@�Y?��p{���q"�M��d]_�,�*�.�I%� �	�8"�,V�l�ѢₜO�����%׭
���myR�'���'��	 )p}��O�,�ZPhX��y�e)K�`�ؑ�N<�����?�����(*��Z���勤K��k�]�i�^��[���	Οp�	oy��E'{�$�.xIU�QPg��AT!ġ`�9�weW榹�IQ���)D~��=! �
+`R��c%�f�΀0�)��)��ş �'�:I���#�i�O8��ExXA�Ċh�4��ϯ
k�D'�p�Iޟ �%fm��$� ��!|�H�ʈ5�����Л������'m�,�dv�@��OT��O�`�Z�H��Z�7%�$�oռp���lZԟP�ɳ*���s�IU�g�? �Ų��2�0�yF$N2W�r��5�i�xJV�s�����Ob�d�t&�����,�L����S� B��f���ݴ @���䓘�O@R  �?4���%�A0�6HYU�T%#�r6��O��D�O�vĎN����P��Y?� C��~���2�J'~�)$��ʦ]&�<��t���?����?����"?����1*�M�T�@τP&���'��]�4�0���O��D.��Ƭa�jL$p0�����q6Rt��Q� ˅�h���'^��'^��*6�  ��p�E��f'��q���%���}�'��'v�'a�� wX)�V-ٙTha���yW�\��韸�	\y�B��=Y����}�E%ЇZ���:DV�l6t듨?A�����?I��ZSZh���K�{3�N�zj<h8�Ǌt�$�A�[���Iџ�IZyҌ�������#�)o��𑳰
%o�$A�n�ןX$���ןP�D&l��O*P�ǁ1~��8WDۖOth�K�i�r�'���@O�]�H|����z�AB���u)r�X�\[5�w�R8/��	џ��I��h3��x� %�|�� հI+ ̀�G�~��ƒ,��nZvy�ǩ0\Z6-Z`�t�'��D�%?�5	��c8E�Q.�}���VE٦�I�4�6�]���'�@�}D,{0
݀c@[�*"4��Ԧ�0�*F	�M#��?�����v��8�HY��*ƞ�^u��j�>q��=m�)x:��?)����'𬉀eC�&]선�o��{�����i�����O��d��Y;�5�>���~�,�X��=Z��g��BL��M;N>�qE��<�Ok2�'�R,V�y��X�U*n�R�	�Z<7��O����Am��?N>��Lv��aC�
�-N�bP�S8:�i�'���c�'��ܟ�Iϟ`�'MVe;"��l�p�B�S�_�N�@��O%#:�b����J����	�=���3��H9IĂtc�	ӋO�9q�������'��'�r^�*������*Ԝ!�8Ɉ�H��Rs�/�5��d�Oأ=i��?�z�"�)C S�N�aH(@�a�\�c��p�P�iaR�''2�'��	� H+H|SH�#
� ����z���4B�f����`��H�ş��	Z?��e˛caj�3�E�/i|m9���ɦ��	����'����2�-���O0���$�%�D�Qr�hQ�g�<+.̒��$�O��sM�O�O��
z.����o<X��!���@d7��O����C�<���OH���OZ���<��O���D�T�_��0�T��-Kn�nZ�������""<����J�<���Re���$��<`2C |4xHj,7h�t�ѬB$������Od�+�Ɔ+�A)�U�i8�-W"O`X��"�GvN��ү�>,� �c�:w:��5;xI�zSt����5i��1���6Ś	p��&3&a߃�*��wD�2(3��ґ�\�#!.m!/Нp[�|#r��"����Sa�	�z��F�<4�}�[�7	~�H��Տw �8�p�hF.y�%�٢si^Z��uG@���O����O�8���?�����X�
(���f�1L��ѻ"��/\��s�G48�=��R�u����8�QJQk��^�+Q�dZ�I
F�4�R�u�t)��?E�*	���Z�M*�̚K�'��Y�lY�e��ɡ�ǃ���Lۻ�?����hOL���4
�xp�ph	�tK��Q7$ D�����2xe,t$5E��a3W�<�Ɋ���<Q3E�����p���TH��a���ڴ�_��ɀU���쟄�'0{��!V�T�*� M���߳�M���Bk�j��q��R��D��d�6"\Э��Ϋ~k�-�a�<�б'H-^����Ϟ�5�����'�bxa��?�+O�4�ІE�	�!���0��h2��$#|O��� �R�2t�Y3$�*
sDi��ORPn��Z��;�m�=H�Nh���J3<ư�I~yr'.5����?9-��؂���O���ɛ>H��+2�`��mKT��O^��(ǲ�q��S�T��i�C(�'�򩁹���`�E4������@OX1��+9�9����H�0��V�Ǯc�l���	\�0��}�>qG����j�O��"�tN���ED��Jz���(O��y"��]�$((�ݯA&6(�C$���0<)�鉥/:��I7�����6�س��A�޴�?���?����5Kؚ���?����y�;$-��q&n�bQ�u8�˅q���3�D��W�d�|AD*�aZR�g�;����(��lC�%��FT�R�T7[���	i�0���|r�� g��+V@-�#0<\d����"08��L>B�^@��"�A8$��	i�<	���P�@���ޭh�� ��e~n4�S�ORbY0���:�ֱi��Z�g��p���|o��c�'�2�'��xݩ�	�ϧY	ucC��/Z͆�K`�G���9� �, ��A��n�#4�^XHϓ)�x�He��*`�H�JΎ�\��T&��b�.3���2d�> R�a�.UR� %�US�b������������?9��tc� ��m U�1P��h'���y��Ř"�TT���t�@�S����'�x����F)l�l��4�ɾ&�u3�e�R����f�0eS�a�I�<�����$�	�|
$�ʟ�'�� 0A�"HS�}8��[([0(��';��،JO�~�l��ʃ45�E��e��p<�.��<$�t���4���C#���<ލ�6�8D���"��1���Q��"MU|�X��6�dcݴf�1��$�2&�d�C\�z��1�<1Ƥ��y�f�'�?U����O^tQ�$�5�8u�Fo���� ��O����&Y����.�|�',���3a�1>'|9wj��V�>�
J�$��h8�S�'l?T�8�([Bp+f)�{�ŤO���'�1O�>l���]�BD�2u`3(���"OJ0����N<�����`���A�'��"=�fD�g�D�z��23��T��� nǛF�',"�'��x8�-XR�R�'�>O��	�_�X�c��2A,<C�L�-
81O��"��'t)r��]Vl{��N4P�0YX�{����<!�-M5@La�a�21*�%S��;��'-�%s�S�g��?q�lbfl�	n��C7e�$��C�I ��S�(4Y��*�@:�#<?y��)§?�����W*]��mA�ō�x���,�-&������?����y��`���Od��!�5b��B.��/��'�� ԭ0�(W�\�-1R]�%��`�,�ƇN,e*C���/1�1d#S�.y�q�,��J�NI���O��$̮mj�C#�7�F-�R�5g�!� -1_ƈA��J�V� a�e�Zc�1O���>A�۸<���' ��O�2�5��׫M�^Ar�؃l�b?O~`�$�'��:�0�Ұ�'��'F��1 CH�jp�� P��Z*Ǔ*�H�?Q�����e�So��1��}X
�i8�����O��O*ESsL��dfl]¶Kں-()�g"O�u�`�kLι#�+I|(�OJ�nZ7KB�D"�`�
L��Q��Xc��b+�3�M���?y˟8�cu�'N�� ��Ҳ6�zKDᇴjQ�SD�'2I_�rp�T>��tH�V��͑�$�-�re�OH9�`�)�S�l0��2��.J���x��V�8�d�'�(�������O+dm��������RN�f�	�'n�H��I�9��@��IЬQ�ÓG���|�7��b�ܣq�ԅ�͒@eZ&�MK��?���sl��� �?����?阧�#G��8Lxd� ���Lv8�k`ژ�'1�Jϓ+nX�{����o��@��#�Cr8Y�=���xx�(3gG�#d*%B ?��H�#�z̓<���)�3�$J�ue �`�@�0d�����
�*9!�$'=xT��Jp� �3G�͔R��I��HO>�D�H�`��0�c���8`�.V��,VOΟ��ȟ����uG�'L"4��YSa����ޑjC�x�F�D l%!����4P�!w�K�ah�P�u.�	h�ܫ3O�!W���`d1��I
%Ȉ�7���'��'���'��O���W,ʥ��Tn�s�2�H�"OliJsHC?lX��l w�j�4��_}X�����M���?��c�iG�Mc��U+PDA��j���?�'���
��?��O t�BŊF�'6Y
1�|X�e"!#
6���![f�*Ԛ7�Ky8��K�K�[iF��1�Ї��L��d
�tJ��`E�tj���
��x��H(�?�J>�ň�Tm�A8ֈ��~K���LX�<��=ge4G�ń8�`�B�LOQ<qw�i�� a��7�Jqn��JwT�y�gގtqV6m�Ob�D.j��ğ��������!zU��&X��Y��ٟX�	&t�R\��X�S��O
l(PE�-(�f����ݎ=q���!�>3�������V>`r"~���
UBY�P�����/�o�D\4:r��ɑ+@L�kA��nw�}�= �!��kz��t��\ъQ��k�� ��=ͧM���tA	���	��.;*�>�ZwHؖ�M;��?Q�&�����?A��?ᚧ��pdA�)�ř��"7�$���#��'�֔��HW�#Ƥ�mc�e3@#_�L�=��&�vx�� ��,�F��g*X&.�x�å��I̓-�x��)�3�?�$`��9B���
�*E�%�!���_#�����PXf��v�-C�����HO>I��U�a0����+#�����PA��+v�ʟ�������u7�'��>��5�dI�
�>�q`���H�B��1�Ĉc.!������ �@���
<�@���E$[=.)+'�\��*ߊF�T���b�$bȉ�6��A���d0�O�U{��S9Kf���@��̬Q5"OH)(�gG5T��b�����C��d^z�2�x����i��'��dPäј�d�X!aU?�F���'\�ֱr�'��I�-�j�Zp�Y�Ɋ9bw�fӜ�P�#��s�8���VD��q�'�-�q`���~|`f(J%D�cؕp;l ��!���үZ��p<�A�ǟ�$�PZF8l�5YQn�?z�*D���G��������9J}C�)�l9�4'||���L�x�΁��Ń��U�<A�k�D�V�'b�?	�P��OD�ZУ$Dah�@��:ֶ�Z��O��D�Qa\�D+�|�'�"�;W��,�p@�1yX&�;M����:�S��`L��6@>N�T0��P9�2��O�	� �'
1O��r��u��-*�"��I��X��"O��#�*P�		����#>��(��'~"=aL��r�Yq��Y�v� ��)W0@�&�',b�'��aYD%�(Y.2�'����yg(
${���(�5{�������z��'�vP�EM׻C�џ�_(��']�+�qӣ8:C����"���3�#9�Ջ`�!�	.�E8�7O&��4뀇I�l�s0�X}Z ZG%�ش�?Y�C�?���,O��U�r�(��&ɯ&��4x�[=��!�O��%��0}�����Z(����t��Pkܴ|��v�'��6��O�˧��i���d����Y� y��WK���?�؄K�C�O����O��NȺs���?��O"К񊓟t��`m�U��x�cY>,��aH�	�:z�y�.Ek8�4�t�:3�@��5@��oP\�bC�B�!K�8lo�U��c�2B�x�LA�3��� �I<V:Ua���21�����b�F�k���p���$-	�9��<K�#ѱw��L����y���	;�n��(O j� �e���'N��Ә'�O^NH��L��Z�pB�W_����'��U��ʖk����ĕ�'dfL��'ȽJ�HKl���b�$!���'P�;�M�� ڜIUKNN��b�'����D�xς��T�MA�x��'��"&��S�ȝ��e��D�j���'̖�#�JZ����kvkR�5�@�'.v��sI��d�m�Ba�:@��8C�'��uj�b;��S��D����'\e�����
��iѨ�;��S�'�)q@/Z�K�6!�׈R4� 9�']l]��������f� %��<��'d�����üG�� 	E������3�';b���� 
)�)��^	����'��1:!)Z�x4�d�d�i�`�
�'� ����G��!�f�V���'�"��v��N���[��X�'�.�WLD��Q	
ARd����'#��eL�9����V�	9D��}�'�|M��NZ�\�Va ��܍>b	�'��`��F���$S�M'����'v��0�F�t�V�9n"j�t��'�P�Z!A@��=�W�Q:��Y��'�Ș��Ôn�h��M�5�"Y1�'�-Kc��(R�.X(�,�=&p�`
�'����{�p�'�J���	�'c082ՋԦk�J���cQ?�Q	�'�BD��Eʀ���
.b(��'vra8��A�$��ri�'���'������-C��a$�p�h98
�'L�;#����Ypf��vla��ռ7z�Oj�}�'ui�u��H��9�qL]54^zM�ȓd|p}�fE[�d��S��2E���ɵo^�E
�'<� ��S �����\;�	X	�_�l�5#�>	��I�8;��ED�1s��(2��Rn�<i�	��nE�����c��!oh��?(�mBU�2�'Gq��0# Ag?8
''ܚ�]��S�? �:�
cUN�	&F�P��$C��ͣW����=���O6��EΏ0$� �`o�wn���"Oƈ�d�Y�Z�	`�ǨA<�����O\�1w����>1ufUiJ���tbWHņ��7m@l��l�'�8u�s���o��!��lJD��'�X�t�4b
FX�t$�7jEnt�	�'���5�� #��JQ�@i��e@�'��ᇄO	 t�H`�dU<D��'w���A� �D�ˋ��2���'�6b��E >d�H*���.�v��'F8M��A׏(��d\��ht�	�'" 0�Ǚy��q�bo��[�rġ	�'�Hz���+O��8��@��X�<Y	�'���	�K'h��P�*��Z�ޅ(�'�v��4
M3)�V8�pė�N \��'�t�"���u��#�,9�y�'A�V�O�W
@Dk���)6>����'���x�J
!)��1�EH6i c�'i M���$_��H���^��\��'Di�U��b������1!j�m��'L�(adAHE�a)Tn��*|���'2� $F?Jׄ���B�f���'�� �e�&E�Q�E#�nX��'Fɢ��SU��H��I%��=�
�'d����%v�@`ÑD:s
�'�V �G&��GR܈z���(z���(
�'�20a���(PP�0ɳ��i{���	�'�b���H% 4�k�O�h�ʁ	�'1� �O� �����D�\����'�l4AkV
D�r%���X�Y$�A�
�'�� fh��t�~e�7.�$CX6AP
�'V���'m@�b���b��18G`ܠ	�'��Ij3@�����3�A�1�ĭ		�'@ě��Q��1�ƅȼ*�����''��PW/�3D2�MI�E��Ęi�'<�a����@��y���xmr=��'�  *Q)L9���u%��Gj� S�'�H1�p��p�$$�p�Y@���*�'ݺ9Jㆄ�r���
aDU	a�][�'�� �E�M�VZT��U�2�2	�'X��Qj�D�l��
A�IH&)�	�'ޤ<@����k�`H0��"@D�a�	�'���[i�8���W��9Z|��'�.X�q�H�zF,L��`�7DU�	�'9��A�ƍ!6ʥ��4[ �0��'Jb�r2�A�W���`ǃ[�R���'%R�9�nĩg4�a�IوB���'i���Pj�.p����Ǐ��}"�C�I�&�(�`���r�)��Ɣ�;	�8
`�br���矰۰>!��O"�a�ΉP��oQq�XR1�	9{x^d��$*��DV���`n� ����.�'"�!�$3m���vНP�ZTM��]�	�?�5���_�D#���ەo�"Ё���6?RFd"B'9\!�d^�z�0t,�;N�[��X�5��u ��B}���̺�����yb��J�$��7�OtҨh����x��N��m�AfԙS5H0�ag7r�c�,�lV�yՃ%�O��&�L?{�`���p���+��'n��k0B� ����>��+�;����3�E?�v�	�$_x�<	Q�� 	:UP3�S��P@1��t~"f�|?����bm)�#bs��T���S�!s
�q�'�Bp�<���}��`�Mߊ^z �����.Z����Q�Ԓ�H�
/fc>c�X�0kr�F0�qg��x���E9�x��kB�w����#bƍA�@��c��z)f�:g�(=*v�X�o�9�KQ4�H,���ּC�9���Z�z�I�b6��X�O� �̲wN�)�x5����+��EK0"O�q;Rd�#}�����$���`*@t~�ލ"� ���U�lԨ#��J�K%�xKŤM4pl��G�e�<y'2�2% ‗�#�@Z O�y 3 \�<a��� |Ҹc>c���Q �Y5�X�j�j����;����%@���B�Q�����A�^��` �>�:[�`���bc8 0�y�s���-��H��	���!�Q̚�?�dM��O�0����+zU��P
L�D��h"O\|Ӳ���X�lI�%I�E(>�s�"O�����9N��
�d�Ȁ"OyʴI�)Yp^��n�)R�9
3"O2T
�E�5��1�L��Y3�i�P��j�L��r\̙�B�8�0|�gF�#sR@����J~���,Eh�<IVhD�Dq0�`G��>t2Ĳ	]�E�K�']v��-��((:��O&M*A�3hP����Bɠbm.Y�u�'V�2��&��	۰���N��Ur ��c�>X0x�a�M�����(��y2r)�,�8��қ��'$�x@�ә�Mc)H/�������u�x]y���!bY��2�͆Qb��:@�D8f����rN$D��`�����횤�?2i�,������f�K�=ST��*�%�����H��(t�1AI%>��QD��߼ G��<\���.Ɂ
�BP��`h<1�k�������؞h�`����.6@�WハY��͈DޮA~���pk���ٯ;�"P��c��/d*�I42��FHJ�=��-����v"��DK�9���'<O�D#E�I=R�ѹE�ݒ�VT@���\\�"���?�^,jwa\7 ��]���Pr�.">a3$�a��d��g��^�\ ��aO`�Z�L �'a�<єR�=��p���]AX�D��/(*�[��
ZcT��d��;j��򆪂��a~"�]a
*�u��.2:0颇Y"��E�' :��ƨ�,�	p�M��JpB\����N̪�!V�i�`0TiC"F0h����C�̤ԡ��=� �{����	�Uφ(��̓5�7����Upl����9�0������	��<	�nE-O�^�JG7 ј���QPx��X�JF5$��ɺ:p"�:�I�!tL��@��:Kw�C#J�X�G˜�m�J��pO�d���9��dV�+< �K��,̴�X�a�$��'Ĥ�a�f~�)�(Y�h�� �)����s�-EW��cD@L'���C�f�$��Pp������dX��Ԕ����7Mn�s�k.k����'��)���8�)��q>���ٍ2�n-��wޱ�dƅ�p�up�ST���%9D�L[��G���f��m�$�#�k��Q���4h�?,�m��^D��6�����-Rz��'ɠ%3$	��H��@���x��'I�$1p�/`
� ��ګ>�����e�%]����*Bl���� �Y�q�?����LF�{�l�C%O�B|�u��	Y�����,
��O�C�"�A5�
/~�����x��!B9è��ɑH=��Bq�Ɇ3��(3��Lp4�OְSbK�B`h�9���N9�t����fi���ؽ�-��A0T��'y>����Oy����I�7Cb��p��S��?�c@�;
�y3 �^n�'�����T
�Ж	�XG��N2�!�Yo|
����M?5V��D��v��$�¯��.��dհ)�$(h�z����e�L9�p�c�ͯ2��h&��#,�S����|����!&Fe~d�`b.�K��ТF�{H<H�\?�5 �'�1o���@�ĞV�� ����'���<a�j�MK�Jg��*��x��hh<�eK��}��}[�#	/�! ��V�E��h��'@�C�D��Iז��U�	�&�jϓM߆���y���&�~�O3P:5���"�y"(*�X�� �_K�1��씩��[C�����doW�m��\:��$	��}Yu�	�y�ѓd�YC�#=V�-�lU�Z����'*�*dZDL���/ޠL��E�	�'�Fe`7.,{v$��Ȃ�,���$bUr�!���?&�d����*���hN��y���"1O"-� OK�)B�� !H�t(���"O�r�)�-���j��^�`��0�|2�_�h�Oq�,�&�0��]��L�
q�B�"O>���9�BbTkœtfF����͊U_0��DA'�h���)>\���!��Z&#��BF�
�,��eH�üEr�O�����3ye�����ɛ0�*I��"O� �2�$��E��4�w�+)���1"O�ɲ�g�>o�$3g�
��2�"OL]� e�bO�#��-h��L
�"OBI5ĽAZ�3!�Шa�&t�"O8�X� +&��t�0d�6w̜�I�"O���gYl�����ϜN����""O�ԡ��Τ!n�!�)O�!�"�6"O�i1+�	cp��E�K�kI�T)�"OlD+M�ll��gG6,r���"O����f�gR��^�8$B��V"O(��읮u+8�2BbX�r�"O�d[B(�-~�F�˶ �U�"!��"O���&�'k��y�a���:���w"OP���\�sen�����r�ʥhV"O�	��΄�"{��S�<:rF�c"OhURnx&P�*��xx��u"OL�de"&��6�W�/�����"O\���?�zL�#���kЀ�U"Or�����	r����+h�=`q"O�H��m��	&ݠ��J�$�� "O<(�Cţ\큡�ǸB9v�U"O6�A
��7�*m�Tj��Q)4�y�"Otha�}T꤀#(L�Pɀ"O$��P�^�+K�2�ȡ�FKZp�<�a��"6�����B)i^K7@�P�<Ydf Ti�D�!Q�	����J�<�t.�\<���(�\g���5OF~�<�"��S9��*����9fT��v�<��揟V�D!D�D�:���2#B�p�<���@<1��2E_8
�d��.j�<q���25�4�w�µO�vㆨ`�<y��1��	�2(�/9
����F�<����ic4�3�ǧV,Ա�Y�<����N�R�Q@Aj �z��p�<A��?h��"#!N�<���BB�o�<9b������sf�5u�J%��o�<A�d�-�T��"&.|�m�@#�i�<i�)��+	VM˰��9�ё�	�q�<���T�x���jN���`�l�<��
�-=�tur!��=(��A��<q��D\�0-���]�`I�s�<��Ɗ�.Gf���G�6+D��*
v�<�1��� �h�p�A�:ƾ!�"HMr�<���	(�u�rYl��(���X�<YG��-#�x���#�z���"�p�<�4�U�_,��8 ���8��Ee�<�s⇫c%ju!��@�ƸM���c�<aa��N�I��lX�W:>�`�Kb�<1�k�8ՐH��݆+��8yr�O_�<!b�3O��\�gNV��<���aC�<	rJ��	��i�g�
�xqJ�����f�<ɕ�_�H��R��T �i�<�%l��b��L2��D�&� pG-�i�<��Δ=M�@��K NbNa��"�h�<Y�Er��Do���1)c��e�<��6D�d�kE{o��U,h�<�2�Ҋ[?8p%��E� ����j�<i'���m}l��cOɊ%��5
n�<i�˝�7��\���TY��d�g�<Ym�$]P�d�7��2zD�#U���<���ʚi ���%��jK��B�hC�<����^��(@#kY�;Ĝ�ʢ��z�<����p{B�j6�����TM�|�<��`����S� �R�A�*B`�<�  �b�Mм?�>=q��;[C���b"O�Y�N��N���!�+<b� �"OP�Ч�Oz���C˃H}6A��"O�y�Jܖa���A��_��d"O��z�Ȗy�)��ڲ(�����"ON��#XwA��⑦��U��-�yR�ɖE�����`Dք��F���yR�
"jd呇.T�g��Lه�)�y�;��IÍ��b�3'��2�y%��1j�Y��Х]&��Q`��y����_���4��s#�=�����y���"1�a��ǔj{�Y��f�y�D�s���R@=cφ�jG���y�GP�-��5劈[6N\4���y�`�rOm3F�Wdl=�V���y2HF�-|-�׊��^��D�f�B�y�S6�����ݟC���a��y�� vۼ�P7n��9����e�̱�y��Q�z�K�E�(c}�d僗3�yrA����/D��ڬ)���yr(��^<� �Ѝ^�*�v�3�y�=hڐ=��˂��TP�l���yK�7�c������$j	,�y�@��^�^�7���`����e��y�*�S���S�F�i�b��㥑��y���7>�S�kקh�lL�-� �y��"�.�Igj��UF�}!g@��y���X���!3�ոD?d\r����y��a��`J��׏8K���R��y��61 rPk��@/�thZU
^�yB���F-2)����U�Y+"�I>�y�@V�yK��Zc�����yr�ߌZ0		S��;Tp��C^��y��� ��`z�Z�b�]�ф��ybc��&ݸ��D-#���Ѷ��y"I�>	:�P��L�� $����I��y��#
	�A���tf[Gf��y2�B>�D	6��HfԪ�'Ο�yr,.\H��"���("b��b�	���yҫA�F�d�W' �d0�(1��'�y"��v�Cg�WC��`�
��yb$: ���1��Lh��i��Ê�y��I�B��(ִ0~�#�I��yR,�;FX��e�Z�� �ũ"�y"GL�'�,h�!-�) ��"uK��yb��$8g�
hJ��#�'�y�c�Hf�����)1��c�?�y���8v
 ̉�.W''�6#҈[��yB��- ��bF_5vǼFq��j	�'J�r��I�L��
J7�|]��'|duK�+a*2�#�|�:tb�'~JySfEbˢ�8���p�=r�'m�h+qBΖU|�(80'ͱQkL%0�')�p�WFR�hyq�*J'J�u"�'B��pjׂp2�@
W 4\IA�'��)�2D�Iy��C�*���	�'��|r�H�#���`-��)^��	�'��͹t�0H Dk'/�+�$(�'9<���i���蘘�0��"O>q�q��#p���dg��y�͹5"O*h�F�?r<b1  <5��"O��፱]Hp�#e��0T2�"O��tjޗF��aqSD�i�|�`s"OP�FG�5hr�5�ѥ!Z���"O� ��j!'�`
"u���I��5"OָsƊ��_��L����5!X]kw"Oz�0t��\��<�'��W��a�"O�1)&�D\�����&l���"O��3SdȰ4�Z������"O��bfQ\2p�_��hME"O�M�)2����(�l Z�"OhnFOI��v������&�(D���7	Z�h���3�	F��yBd�'D�SW�@//��Q�ӡ�*1��T%'D�P�f COn1A�/���M�q��z�����d^
N.�q����D��8c�J�H�!�-���e��@z�8賩M�#!���'
�#��Fw�	�VZ�!�d�<29ny�Td��0��ZQGT�N�!�d�4yT�`1����ش���4/�!�ªt:��*�K��&����d�9$�!�I�*j��r�bC<%&�!ƈ��p�!�$L�m�苗&ߝx�P�gۛM!�d�E��)��� ���+L(!���wy$����ƚ�:(����6�'��F�iDqOq�RH���7d�y�.U6l`1b"Op��H�Ep|x��,�w��%����IܓQ��I���L��2����[u,�xSG�<?�����-D� ӷ�F���a����΀@��/}����p>�o�:l0\tsp�M:m�,�%�^U؞x�T�|r�_�OA�6m���A�*	��y��f� b0��e&	�ò��'fb�q���� PL�48`!S�Hr�P�3)�y��2�9	$GD�8�2����yL���@;� ތzK�i�R���y�ԃ���"N�	<Pa���yrɏ�j�\��G��$�p�劷�y���|�]P�W�(�8)J���y�D��s��[欖�n�8������'ў�Ԉ��W�kEB	sF߁f��!�F"O�#��]q�ԥA�DH�B�1�"Ox�A�fȨ#�p��7����5	��>D�DC B�Fd�A��-*rD� >D��4&�� �У�lp�C�;D�����ƓZ���R!�4jz&��B�'D�tѓ�K#k�=�%���2����!�$D��)`E�J��`;�FP�:b�!D�@p��O�`�n��$E*`5(	y�� ��xR�ҭk��A��J��Ïם�yҏ͛%FsQ�ߕ���%Y��y"�ցpQd��U{1l��B˴�y��J�1��'��6z��0�K� �y⦁)C�����,m�\�ڠ�ܟ�y�Q�n���h����ś�CB��y��
�lbt*r��<�|�x',F�O\���ߺ��t�0zph�'��!�$�9&�1�$�*�42�/Dy�!�$�'S:�D�qď0��Iv��G�!�HuW�}(����Y�P�C��V�!�ć\�`���a)� ��0R�!�ErR��b�̚0y�� $��(�!�Qi�0�M�C�2��W�O�i}!��7���1�摀+�T� A�G'L}!��b� H�AqUVŢ&��Q!�_��H`@g�z�n�6��
�!��p�jD[�( �T�Hq`v�^�G0!�^�m�0pӀ̀�wqLA�Ц�t!�$0\�H�$oP4'^�S��4 R!�� N� ��"��	�&֘<��!"OP�!@��$c`0�#f�a�tȢp"Oԅp��$9�$"�k�Z��`"O������x�n�Rg�-]�V���"O<�*W�_=j��xGNs+�[�"O\�0�E�7� g䏿Y�� �"O���H�'� u���7 e.-�%"O���3��O��yУ�&a��i�"Oz"�C�.zf���%�"O�5�S��K�Z�&A�t4�I4"OL�3�#��h�����cU;%����"O<H1-��@ԞC
���a	�"O��g ��q����n�����"O��[@郐7x°�@���~q(�"O&P+��F��(�J�G	fy�T"Ot�� -S����ޜ9���K�"O@�0�"-�<�rWL�	y�a�"O�ĳ�L<�*3k�E��Ԫ�"O�:���;���S�i�>�@�J�"Op�R�k��"D��"��#�ȼit"O�ܚWL��8�D��5@��U��}q�"OP@��`'2wv$�`�T/�Ta�"O�i��˘k>V�r���f*v(@ "O�\��"�!r�T��m̸M"�y�"O��@���7nk�5�6-�LB�S"Oz5`E]Z�{5�D�D����"O�j��O�8����,/j�Xp��"OZ����������<s�"OF�(ga]t�.��>*fʐd"O<|Z'm��e_.��&,�?c�K$"O4�ڡl�#_�e�W�TxJa3g"O�
f�Z+h��x8%���fq."�"O�Š�&9M���I3`�t�"OT\�O���������!"O�|��!��+2���"�zѪE"O�4�&R�z8�P�p���h�~���"O��A��%hvk'���f�8�
�"O:��D��9��<Aa"%Y+��Qa"O\�)�����Q��V΄��"O�Pe�4�|���l��yQ^݃@"Oj-[���9���i�[?Z�k�"O�!��H�VдG���v@��C"Ob���Er���)�^�-��ٙ�"O$M��R���Lڗ(�ҭA4"OP���HG�Q���P�Fo���"Oة�kĈj��=�4�˃��	�"O@�C`Η� �|�Ѫ����E"O���N)h�>]QFl�B"m�W"O.`� ��#c<�P´ ֙{	&�A�"O$���S%�����_/#�Ruy�"Oƨ!�Ȕ 7S(-ѓ]Ty��"O�9�ϗ�V�X� �m���P��%"Odp*�@I�p���Э�+}*YP�"OH��a�:?-\1Q��HQ���f"O��x��FGz����e���R"O0���ׯj6$�	����>!�L�"OJe�k:��(#��A��# "Oμ���JI���BL��Z��ԃ&"Oj4��۸Bt�3�	!C���"OZy!����~5�3�ٌm�r"O8�0�Y�-l(e�b�G3\r���"Oni� �?@*,��B��6g@r�"O@02���iup#�ѢWK0MS�"O�횔#��sr����I�5>4�"O� ڰ�@XT�0�aJ�i��87"O0�A���A��*D�-=���"O�-��mY�dU�8´/Փy�(�+�"O���%Ė]�X����,a�* 9S"OZ�@Bn�1��l@���UBX�S0"O�Y�  Q�fw��p��U4��"O0�
�Ð�uT�P0�,ƍN#|5p"OvUk���
	_�t�aˉ:g\H*�"OLX�p�����q��1j��1"On���@�|%r�it\ ZP��e"O⤙�MK��A���Z�0C��"OB���H#S��Q�c�}%=�q"O�T[��>�
d
�M���X�"O�ГQ�
iox	�� a��5�s"O����'.���z�j�7�pL�g"O�0�$�C�KFZ �� ��b"O�%᫔�7�.\z0K�r�x�Z�"O�Y��D�*�����o,����"O@Q�5�B7�T�O m��@v"O�q1��	x���Z@hďg ��"O�%u�2Dᩤ�����܁�"OPHQ'��	?`�t�wFJ�2h�lBr"O���$�ȭ<��r�R�F�DӶ"O��(D�X&U,�Q񆝌)6R}��"O0ma��D���ah��}.���"O�鹁��K��ӡ�5d��P"O�l9p���IA4�34���u��K�"On�SƋ�k����T$6�$Q��"O��p-��/�l����# ��<:�"O4�8���,XZn�(�\�Y3"OZ):�H,�ƭ�-�[��aAd"O� ����H�i��i�8��"O�� BF4?$�����l<� "O*���F���A3'��=i��ӳ"Or�iWdE�S\���TeE*J��+�"O0�1�㛋���X����b�L|3 "O�蚱���su����߲R�z��@"O�PVM�;2�l5!F�C,_��A�"ON Q��.}��2 ��R�� �"O��Q	�n������w�0`"O��&��:&�ӷBS)N�l �"O� cE���Dl�!��N�%��"O��7G �r)�e����ne"�	"OЌa�����r�
7`�:@"O�{�̃g����L�$2AC"O��ᡔ�6��A���lH��"OdT2�b�
##�A����$7�%Q�"O�8P�E7 �@�D!��,�ؘ��"O&�q� ПOư2�I��3�"O6D&�t����'H�=����"O��Yvۂ`��D3����~�V��#"Oؠ U&_�Y9�颰*�
�~���"O��0��*�P9�c�цz��rG"OH$�S�1?�ڔ�'B.N�T"O��8�ܘe�n9�Da�P���8�"O���Qb<yH�9��"ў����"O�Ɂ�I,9�UA ��3!5 ���"O �J'���e'�|zU��;l��˂"O�wn@>QL�q�pA��g����"O~H�%��!(���u`���T35"OޜkB�̀���:��P���ա!��Y2Vd
Pe-y�T�Y�"�c�!���D�J�c�A�J�6��S��+?�!�d�i�2���h�W���w G�"u!�� n|c�)Ä,K��гgL��"Oޱb6��	Z�x̹7'@.@��{`"Op�
��ͦ}-FI��ߊ�#"OL���{J�H��4h��0ڥ"O ���!=�:� �����2d"ON�!E�� ����4��&0��<��"O�!R�C�>٪l��H�l��  %"OV1C�ꅯT��� h8kB��A"O�@���RJMJWFA!(N(�+�"O,q"6	Ҍ<�	uE^�m?�d��"O��zB���*)v9��s�`�"O(�sK�p�"�Gi�/��,u"O��ض&΁J��Q3�-£\�$"OV�:�)t
p`׋� �@8E"O�ps�f�9
fHx�)��{O��"O8!q���88��p�Ё�.)�"O�!BԪ�*A�E�T�b�b�hf"O��5F�)vER#3	�,O�d�"OL@&�4gX܂�MЧQ�zL`�"O<� �枇0F�"�nO�C��۷"O<�:��C�[۞P0-ʼ$+�ŀ�"O<�؃&�)(�baa�,�$	��d�t"O�u@���j�8,U-��v��u[ "O�9�bBA�v�#���@�����"O�0kD�5?W.�d$˨9���"O�Ś�+V(\yP�H��*���yr &%2ܭ����:9�f=j�lL0�yr&ފV&��!m�,2zP,��+^�y�F��%�����#<,	K2n��yO�.\gRP#�V?;����6��5�y���.�2@���1. �X��y2H�`��ң"4*Q�Ř ͪ�y"i�nq����^�K4@Y��ڴ�y�g��u���Pc+[1I ����d�=�y"	=f��I�⣄2F���(N��y��@��ruS��W� F��"ħ��y�`Oɨ�Sw�~I�xp Y��y��#�
ĨTŀ1x�ؑ"���y��W'�}r�΁k�:K1����yB� �`��1��\�f/��W�ħ�y"ˆk�<�j7��d�p	٧o�*�y���0=b@
ŎZ0Z�X��A��y"�#p�1QRhQ�d��2W�T���xB&�29DՈT��\`j$�W�+kr!�aGh�+����s�j$�Zu!�Ě6�J���"�7<D��K��F�!�$� q����k�	 ThZ�`X�!�ɤ}Jٴ	G0)� ڧM�<�!�dL�x�Q��$�10 rx�DbX�-�!�N(~P����10:�IP ^�Bu!����
�Aveޒ^������v�'a|�ˌKu,�ӡg�:.��Ff�.�y�+�"F��lxd��52�,��j�yb��Z���6��2�
#���y�2t1�B�"l���ɢHЅ�y�C��AZ�a�W���Z���\��y�k�9A	�]�e��P0�*���yB%	z�9S _�
5��!V��y����yhZ!�A�����ȍ�y"�]"D���i�7rY�� ��y�)�����)ED3z�H!c	ط�y�
����/�� b���IP��y���$:�t��X�"��<A�F��䓑0>C��F�jy�ԡ�a� �Ȱ�=T�� ��B@5��xK����^#����"O���dj��Eh�=�e�# �91�"O&庀�C�f�xA�QJ��%��T"O����O��F�iY1JG1�L�V"O\Ո����̱A�h	+$��ӓ"O� vd��8\�hH�/�����'.�'����>��"�?�|=�ݚ�rQ*�#y�	A���OP����ИP:`���	5u�T,��'P�+u'�e@�� ��gh�'d�y;0E �?��y/�����'c���A�=>���Ūjyr�'�$$���\9i�$�*:v���' zM��e�Q;�E`$i	�b�'�L��T�ȗ#�҉�S�µ��M>9������O
�L�E�=zB�<@R��}!�8�	�'�j����::p�1���sʐ	�'E���CE�iv���.��d��d��'R*(�1�9��e�'@V11Мx2�'P��[�NΒ2A�4�	@�*��]��'�ZM���X/�$x�H%���	�'ܽ�ao�$[���M���08����O���>�B�Bũ\�`�� �&p�2����3D� ����	�~�P��1lQ���b&D�8���4i���F�p���A$D�ȩ��Տ�0t���N]��G� D��[$�&%�r��6�M���4D����I��.A��V<N<�P�1D���b'
+�~�:a#ׯVt���2D���3`��f* ��t�Ҫ"��3�+;D���A�S	U��IF��6J��@��5D���+�<����a�ݜH���H`H D��s���Y%���B`�y�$,ِ�>D�DSfA�N/�y3E� V<���%0D�@+f�@J��k"DèQ)9*C@:D��㡭��!32�0ӫ�%Cep�O�O|�d:�)�:�|l葤���"���D�>�"���'�u�A �Y��8��Y72�9R�'����#H�+@��Q �w���'!��á��<����'B�g|r���'�8���
켄���o�H��'�|���6���/��j���xߓʘ'(�P3�`�6�)��Kƴa�(I����?q�����"�����PSii�/�? �C�o�BE���^�� �)�!�D@�v���C� Ҹ������]�!�� v��d��'GcɌ�{�ʃ6�!�$�N�.��!f�*TW`�Isk�7D�!�DL����z�GG�j8�)Kªܔy�{2�'��	������	��NnT�i�L�\����O`���O�˓��D%�I:A&�e�t��5,u���!3-�B�	;U�`)��D�W�.11���l�B�I�f��'�>b~��:d�L	C��C�I�������:u�j�QŜ�b4bB�IP°tEV;D�0�`ږ��B�IDnLQl�� �&��_�
��D�<Y�'�|��#�s�[e�ZF�KK>����)X�^��u�`#��k��p���I�!�D���Ԝ9�&�&��ҷ�ʘ�!��<Y�Y�%�R�:Z$g*[�!�d	l疱�	���Y��ɝ.+7!�D��度H�"��`����R:!�Z&-h��1�X%m� �	�G�>d�ў���S�)6$s�g=�F�37��S��B�	'j����*C1C&A[�⊊y.�B�)� z�b劘4�h�h� �NRr,*B"O�����$�2ag��@;f	�'"O�k��%Co�q5f�_.�Is�"O��˧ޒ&l���Z)Lp�6"OaY���,2ҵr`��d��jB�.�S���xH�P@��?ڔB�Zf�!�DW�8U7ώ�p�� �!�[-3u5ɐ
�8
A�Ġ�9-!�wӬ�e���:�A��g�!��q�}�W���.��0$N�E�!�D��I��!�IȨ4���#�+�!�� ,�ej���:M������
Zўȅ�ӛTb �f�Ŭqz���V���Oj�O �}��@2l�rؙbU�b�*P!xɇȓA��!��%^_|�y1_�j�쭇� ,^�sGAϑ@i���$�ڕD�<�ȓzI���"o�>X�"mH�<D�ȓF-}����)J��UKr�QpNq�ȓ1�p-��ʭT�޵�� iB�ȓ����A+��B(.p��W�^����	hyB�|ʟ0b�0��bݹ@�&�)%1K��e���7D��@EŧU��h��hA�u=��e�+D�<G 
���HBO�*� ��2%*D�d@bY�5"��+W��8��E5D�D�����5��G�+I�6T8��4D��Z�BA��T	�A�P/ZL00A'�OD�	W�.����4nY`��74|r�O�����.�-�V �8������'9*�IX��(�0��v� ��6��3���X�|i#���2LOB�[��'ra��x��{�˘�y�!��<N3�d�a(�p�	H�!�$׼X�xؓ3�^�P�*�h�"s�!�d��YΒLI�,I�s�:���E ġ��%SH�O�7�(5BcҚw��T��	��2��O��X�<0TH��C�I�s�xXa�"��J��B磒z��C�	�m��$xnԻ`�n���� \LC�	���!J�DǙ-jV�����C䉪t���	��]^|  ��6�$B�I�?�E+jN�M]F�@D����C�ɥq�Vm��Ė�q��%���Y�t���7^D��U΀3 ��ÒA]�'�BB�I�f�l���H���	�"ɩ9��C�	1c���)t�:Y�p� L��C�ɓsKD�� �nt^!��3ϚC�ɳD9~ �'ȗ�Q�p*D�;w�rC�;�P��P�*�.�P-޲�l�1�S�O�F�S�R�X��a����f�¥!2"OZ��2)�,T����B�jX:�"O:����$;!�L2�'
�l�� ��"Ov��6�	�G��(�$�crh�3F"O飦��2,���%^5�Iq"O�<�v���>�8�Sbԙ �@u��"O�B���r�ś���te�Q�	Q>!
M4e�]� �N�h����q�<�����4]��KY!y0ei��@�=2��"OLp�a.=6P�����&� �&"Ole�]�4G�R���R!D,ч"O�lp%�H-(�t�H4e

J��"O�ܑg��-.�D�B:i�(��"OP����x��A$�>�J 2�"O�h���3v���V�4,�}J��|r�'�
�'J`��vb�0h�����ˮ""�����xL���^���`�a��+W����S�? ���Ǎ:���#@A�l}^I�"OjH�g��#a�xP�%(Q�-�XT�4"O(��w�8��1[��	nU�i�"O����D�!Ih�HH֠O��т"O���C��&~#�4ɡ/�nE����"O�bi�1Mq�ђeD�n�D "O D�T��>���D��0*a"O��{���^2,8q,O.~��I�"O���'�B�o�.4�"��4*�|QB"OHX	�k�8W �X�!�ޒ��ٻ�"O���4ˊ�sw����W�h�2p"O�Y�ao�w��VI(��.I�
B�=M����g���F1����(d4&C�	�_�F���"
8�8}��M�6f{C䉱��|�D�N(�L��1g�1��B�I,��ꉢJ&�B�e[�J�B�8��+�O��l�6���N�5�"C�0�����V�tS�G��l�C�Ʉ�d��0�K�R��W��]�B�I
`Ä@1gł�c�ҥ��hM�B��3U\:A�"�R� ��͇r�B�	23_z5aК�!���ƩM�B�	�>7��t �u2�-Q���F�$C�I�N���P!IҾK^����c$j�C䉮\H~,K�-T�_��A�)o�B�	�F�f��dE�j��h�rG]�w��C�	�R
�E�0��6�@Z�j�#��C��oMМ�@�S^�8�J�U��C�ɓm7��b�۴[ .1��	����C�		{]F��A�(�&�:���"qЀB�ɒ$ē��@ ܰ��G�F]�\B�I4?CFl�&E� �v��DkF'(�B��}hx�3�ڋ<'j����ś3��C�	�I6|h��8x6T8e�'b�BB�	�ELj�;��׊w�\��
�DW0B�	�}<�0t,��1K�i��`A9Hy�C�Ir"f%�`�Y�j����@x��C�,N�L�!��.Wӎ��e��B�Ɏ�����F���%kW�83C�	�k ����e���;�хn��B䉙,|l-�1G�?��ś�ЮIm.C䉲DU,��g�ۙ}��,�*��B��B�	av@��Έ��J��F�q�|B䉆q���*ƬÀz�.�����Q�C�:P����A��
���
'��^�C�	�Q�������
�eF��'HC�)$��	�W$�6?��樀�<C�I�t5�"w����"��D�!9�>C���|�GE]�+�Y#ĥ�2!VC�I0�\H��G�r��Dr�^#S��B�� [k6�AIY��H��ۗGݸB�$Z�^p!D��2@���3��]5��	�'��"���>�H�!��A�W3�D	�'4��b҈��:H���դ�� ��p�'Z�US���&0��R�*S�Kn���'d(%H�-K�bwR4�+C�Ɣ�Y�')�@r�[ =$B���*� �H��'� a)�R?��i�G@�,1���'y���鞽;U8E1���S����'ײyX����h4ps͎�Y&�c��$2�	or�7C%XL�9qS�ƫRt&�����<AD�)r�8R�ތt+�)��"M|�<a�/�<(��pC M�z���l
yy��'0Y�ы[4F
؍i���[�-���� P���M�>�e��2(�`%�#"O�aI�#S�-=��$��!T��P�U"O0�j�kJ[(4���gy�8�"Ob��,��\ٔJ�1l~��p@"O<)�צ
�N9�)��C�xq��_�H����4 ��������i�e�����O���0=�Ǭ=� 1cZ�X܈�b�M�<A�'�b4u�6���P1A"�E�<��%�8v�� G��d�L��jx�<)�%�f%����(w\��E�Kv�<1�&Z�p�����a't���@�Pzh<�v��}(Q��@[�X+��Xv�=�?�)O6����4ʘ� �F�wcp\V���'3a|rR�[n��������/��y�#��B��]9�OA� �1p#�y2%�� /��2�	�nx�y��d�7�y�k�+c��ҦǼc"���Ō��y�	GI��a�W�N�\P֣4�yJk���@Ϧ5�뢇_,���2�Oft� �H5�I��ENt9�!�!"O�R�f�yA� �dc�$b,;T"OdI�B��_��l bT�(Ʃ�&"O��@܊[ɸ���@�3U�b�3�"O�RB��:E�q�#��X�6q�"O`,3&�,8_J$�Ə�AЬ@q�"O*(P���.-> Tk�ώ,q�\TR���|�Im�ďI9~[<]�B��G�����+W�y�'�3��\����DiȀ�+�yY�THtA�"Kb�Ũd���y�o�W��ɚ4�Y/S�޸y��Z�y���
gH��e���L�0 Q�U0�yr�^/:;�)�Al0V�H��̶�y�K��`�P�x=$�|��ФI���'Fў���<ɠO�;*H�@ɝ�%���wJ�D�<9�%T�P�����5u����UA�<�F�˕x���ŨԆE+��c��|�<!��59��T���?��A�b&�r�<y7 ����C��}��PZq�	d���OO*�0T�O�M$�	��Ϳ\/B5S
�'V@8kU�^�L����R]�a�I>A���?a����O��P�Y0x��������*!D���"�<{[�ઁ#����:D��QU��-%��|:c$��F"�B�,D��3oDI���C�	j��њ�)D�TI4$ҹ0������̱1\Խ���%D�DĂ˳@�[��+�X�˧!#D�軀@�-%L���%�	>|�L��<9��hO1���Z��ªRɨ�c<��e<D�p��I]��0���˰= 	��;D�{ ��;�$�e�J'L��AP�'6D�|�"b�Ls� b�H
7gܢ]b��0D��CM݁V��h�d�/j~y�v�/D�$
� 2Ei1"D�r��5iԌ.���O>㟄�<�w�\5>����JŇ$�RQZ!��D�<A���D�QņT�MÒ�і�~�<��#�����mS5G��a	a�^x�<e��/iҥ���JN"݊c$w�<iQ�Cp���'x�>��r �<Iã�=oi�0������hk�П<���n���Q@�E�r�y�D�z�̄ȓ4�=*�A�,k��!%@.xX�ȓ�(���0]5rgE�%K\����x�1��Gܗ���⦐�Q��ȓ�]!�F]������̦|_ą�S�? (h�%�N�B'Bu�q�ՊZ��("�O�������`���y�1yw+D�X��ي2'��0E䋨~��`�I'D�xq�F^<GT� R�l�S���I%�&����T�AT��0s�0(2Wm�6if�2"O�`����kDD�d�8)���*�"Or�{ӄّD����V�J���R"O�\��nº<��y�ARCP�D"O���a��CB�( %d���'�!��	_���AI8,��Lȴ
�/\!�S:�	��ǌ�c`(ʥPџ�$�$�O�p�тG�|^����K�K3��	�'v�I�,\ 8��4+W�+z�	�'��-��Ί�4(���F��'`��'q��z���_-D��W"�(�'��x�D%��D�b�+t��,O����4� ��0�P�N����@0��<�	�<���ÉdbL�`&i�7���%�H{��^y��'5�O:�9��1�gKZ+L "��K#"J0�"O�x��)� i��	r�p:@"OJ|Rh8��Z ,��\�Vų�"O�񥞵I˦�10ꆗe��5P�"Or
b��V��(2ъ�ͪ!D���3��`����M7:�e�f�=D���&�]�I���D+�'&��3��<D�� "K�|4�`��9�Z8�)'�D*���'�[ÅY�@�X�	��6�c	�'RPD����c�f���Oɫ2[bXk�'H�p�T��	�c���+�Q��'_I D��"#���B���v���'�����AN ۬���㑬Q�	��'%�C�� F��C�-ޤ�
��'��i�҂�<=�����]4�[���)�4aI����|͂p��M����ȓ6��9B0�L=K������;����4�P�%�;��DҲ�Q�|ڂ���:tb,q�+WB z��ΘJ1������0�p�آ7�*,zA�U�<���H<�Ac�9�.��pɀ��x�[�l�i�<�W��%^r:��3�d��`C��hO�'�R%��:a��BpmQ4l���ȓj�ryӊP ^��J!�N�Oޤ�ȓcd�*���n��8���Uv(��#���(��Ԍ5���RU+��ȓCT�� BW�V=|�(� _Z.�H�ȓUʰ� d-
�8����M L!���F�8�@�]�MY�Oͳ2��0�?a��0|�򨗑|.ƀA�I0 ��Fx�<iqՆqRUȷ�M�t0�EZ�<Y�ۤ}J�s��{bB� 5�]�<��N=/-r0B��΄\s&Xc��\�<їHF)2�6db�&قJ?�4`l�m�<y0bD8ZD��'琪9/.�8V�A�<�U�H�0r�*� �T3�0��<��BC6��0*F�]�;`(�ð��P�<�J�5+��Sb�'��l��V�<!2`�:V��Y�hU	M����JS�<�D��0x�@������T���1��c�<�p� W�D%z��6 4}�$����T=�=+m�*p�|�@�&����7[ʭ�7��>&t�C
�rnŇ�%E\hC@/v���d}䔇�Q\d%P�����};���i��,�ȓ`�L�f�!R��I�byvm��S�? �=R����S�X<�^0��P����h��k�#$��
o�;@8��g�;D����P�c׬]K�a��T҆\(�,'D�<�.�*;}�E3G*�@���"#D���G�^.C j-���V����"D��*��K`��q��B@*���.D��h�� ��5��Ĝa�H C�+D�db�b�;[B8õ��DVe���<I���1A��ܨwI�ж\�_�&�Ԑ��o<���[�#jtX�e&+�,t	֥�o�<�F�E>ex��I��:���(5�Dm�<�ሿڈ8�FF�ul��D�JM�<16�@,�(Ыǉ�ܡXT�V_�<yg۵$4���F!�x�dm��C	A�<���ɸu:>\���QI��E�{x�(�'6Z�rb��h�2�;�aW� �J���'� Ph'��
4,�؃��t1�U��'Qh��Q[	-�
\����t����'���p``��jTC�(�f��'.(�rG�H��8�a�����:�'���Y�OǊT�D��(<5�3�'�v,#DMG{!)��vF�c�'V	�� �$	NE��oP�{{����'�0 F���*H����	ok��I�'�X�` T��vH(�'�`L�k�'Z6e��,{��L�M� Q�(p��'d�ibE)ׂK��6
�-N��@�'!��1"�h��MeI�E+��	�'Ì�7��
 �B�)�(�=�� �'*}z�n��}��ف�쌇 ���
�'�p�����5��/�#B����'VH�9P�ۓTs|��H����5Qϓ�O�����ŤuL���b�G�@YZ�P�"Ov�c&��]B�i�P�E�(T�"Oh)��3-���ZP��PH��+�"OiphB�m*i��\44��S"O��z�[�I@e�g�9Q�>0�A"O޴3v*��US���D^� ��\�"O�,�ш,X���%2���"O�d��[$$!����+ڀKij�"Op���*��),�",�F��!��e�
����]�<��bL�~!�ęf�F���
K�����Cq!�׋E�B�P���5 i�(���k7!���4[Ek�F	:Ă�1n��h/!��1A¨1&�PP�X��+�)4$!�DAS� �kek��`L��s��U�@!�$Vˤ�� �7��A"��B4!�Ę f�,ZՀU)K��d:�Eݕj%!��&� P9'ٮ[�����I��R�'���'@�)����O�n�����m_�1����5N̜{!��?"X�KR.��p0I-bq!�D	�;9L�Q�m�	t��e�ӻ|g!�$�$���-�*	R�Ұ�N�i�!�D��6�<��W!�43��y�F��b�!�$�5P��m���)��U�!�d&H�8b�N��U��ֺ�B�'v�|ʟqO�c��&�4��
�66��"O�r�ڛK��)���A3f%X�"O6i�ƈQ�kٚ�@�jA�u����D"O�-#2B��s�zE��j�P����0"O����M%E6L�p4cڱU���cT"O�a{2�%+��ܳC�:8���;R"OX�$M��Z�@��&���kи����O\��;��3� Px��jċN�	�ƭ5���j��d�O����P-���RQf[�##����  !���'&Gt� ��N�g�N�I࡙91Q!���n��k�UQҀ�!F�.=!򄔖_��� &΀�4x�)B Ɓp%!�D#y���J�c��g"�5;R�@xw!�dK#��ܹ���1���F��-�!�$�1�r��� :��4i���}��'�ў�>���j��O�fa�A�D�ze�v�7D��A�`nHD�g,I<xRI�2J)D�$`�F�(N]�"�̉Q����9D�衴mZ�f�KB$�m?��۴�6D����V�en�b�)4�b��v,4D�`Zrm�@&\!A�F���Rf2D�h�Q�t���Q�6o<���(.D�P+Wi�%T��*���|�Y&�.D����$*N\�b��=P��c /��9�S�'����L�B���d�BJ�-�ȓzeBEɊ�-A��M��L���c�*P �e��[��C�<��y�ȓz��u�����4~�GF!Rq����3fI���(�*�z"!+3�'� F{��d		����M\�W�L�p�a��y�@ȗk�y���:�z|�6�V��yB�4�
���1>��i�&n�-�y�h���߶4�v�c�'
�yR,ݸf��;��+B\�LBl� �yB�I@����,m��٣��yC�'�zY�v�}U>��d�۷��d<�S�O<6x��!3�����W=5t��
�'+�%YU�W��I�Nҕ%����'@D��1'�1�X��KȚNz,1�'4\��a�ШW�IS�UNd�E��'��x���	4�<Sr/�	u2��'�\�BG�1"��!n�YW���
��-���L
���B��ZQ�(#
�'f���K�/u�m�>h��q��'�(-cA��P���`ӀL&3+"��'�PM�Vg�.v��Z��L�;-��
�'��E+�'�0XBڔ[%*81���	�'T)r�K���'�/e��|�	�'�1u��-y��\hb�W��}Y��hO1�J�O�JY���y��(���&J�P��'�&@��"�O#u �,P+�<��ȓP�@U��G�1s��P��)^�����Ųs�ܿ,���0�>
��ȓu�))�$�<�h`��%1��ȓ|��B�
O�Mw(������>��ȓ?�hsj�����Q�-�2c���ן��?ͧ�O����΄�5�2��&I�����"O"@:C�5]��� k�.�'"OL���n�j5�L="� �2"Ob�8�
�2B�
3鄲Au����"O�PցT�c�L)sp'^�v��"O�	���M N����&F[H�t"OH��_�H��x�R���*U��Q�PF{ʟ��'^2%�ujF�[�F�NF.cj�$��.H: @�_~T���$5����#�I���b��u�&n�
3h؇ȓ!�l1s�[��)�@M�5Kj9�ȓ>���A��/r�(�%
2HGP|��1�q+W�3ͮ��o�YQ�}�ȓs3���F#J<O@U��*Ѵff��	k�����	6;\���+M^��a`��]|��B�)� �4�uH��%����`�u�b�����\F��ŧP��a�#�ư%���у�y�f%x6�i�Pjшڌ���`���y2��+a�\+R��e��;aJ���y哻<o��H���[��qkw���yBGB*g�TDr@�ø N��/Ǌ�y����/��P�AC�lBl"���y�,�1#�H�y棖"��`wF7��O��D�O`b>�ദ͔C)��+��+����"c:D��ce��%%�
��A\�!�~-1Ɓ"D�t���awh���]�:۾���3D�H�G㞝=5�� a$Q�<jƁ� &D��X���ӥ��';xZ}c��jXRx� Fx�k��I.������/=��R����y"�D)
t`�C �/�x��S��y�d״?p���,<�k�)���yr$�O;	�g� �fQ�N��y�ǺV��ɻ�0c_��f�@!�yҏ������(�A8DA��yr�_�w�ZԳEN=����D���䓗hOnc���T�Â� X��D8v>N����&D���3��Ti��8��	&��sc0D�ĘT'�o���u���P���2D� B!��.je��Bu��2����L-D� J�\�^�Αpa)W�I �R*,D�D#�س5�\l�Ħӌ�� Tg)D�p��c�1�l��CD��O��  ��2D�Р��_3M@p��Hb�P�k�g1D� p�j��!����҂�!E�<	�q�0D��H�f�
D�Y����ʲ�/D��xk_�XQb�3�y���.D��{AbƂD&��0�%����L-D�����Lh��D�0 ��&"��yD� D�p�BON�=���D��<:?T�`�o><O�#<)��6 �s���&H`|#�GPr�<�a��Z��	6�Ј�d�"��i�<A!ں7��mi�hW�Fm��GO^�<� �ܡG�h���f��qA$F~�<����p�e�X�H"�Ls�<!G�L
[=<l1u�R�H�ʼQ���c�<���M�8�ш�B��q���_�<���׍H�1&'H�[�Q�^p�<I�hK<&NP
rY�#��@A�h�<�㌖D&�P�󥁐c�`=ɴ.e�<���&����d��,�� �g�<� ۵"[���P�?(��R��[g�<A(y��:��I�@��*
�_�<�2Bb�bPۓLܑ/�L�Z!��]�<1b/�4�A�(��h�y���U�<7*�%���:F�_'o^�uKh�<��!������`�<� �D�c�<1t��X�^@ےdO�N�Aʄ��`�<�&��9nb��ee�(
u�@���Qx�<���Q�JS� ��!8�Z�ˉs�<�hD�2��G��(V�1���k�<�𬑰d���@b�((�g�i�<�; NI5���7b��T�i�<�ƨ_�����N�.�\�@sIEb�<����cNt�BC(-4��9�(Dx�<q1�. g�$2K�p�9a��i�<���
{�QGŗ��%i���c�<)� �;ˀ���\�A��x�A��D�<aw�ôx
��ȿ:"tI���j�<��C��D��C�/�2+���I���i�<� �A�T�����y��A �ih,��"O���eF��D��A���҂M|	��"O����o��EJ� ���ݺ1IV1pc"O��3��\4f*��1�ޢ^9,�P"O�	8�,�W$���4�@1��2�"O�ب��YЄqF�6*�k"OС)E M��x(�҅R<=%��	�"OB�h�O��F���bЄ7
����"O��P��3�:8ڇa�;um�%"O��B�ӌ)���JژS�Ȭ�C"Oz<�`S?�v��$�:g����"O�3�uZ��Ԉ� |�ܜJ�"O>�+�mU?B~1�!�
;S�� `"Oz��"9�੢�Y9"�.aQ"O�	CW4;z$+E<�2�$"O�K`i�PVP��i ����"OT�-T,Πhp���ck��"O�ę'�ة}�`��'֪&BR�"�"O�MH�%�#0`N��'��U4��"�"O�=��e�0b6��s0��Pn|k�"O\�3�H�,p��1���|���b"O� 	p�9!�U�A��n�1�#"O��q��:�`}�BH
G�Hm[�"O���r퐠|���%�C��r�T"O"�u+�.�J�����p(i"O�0"�h�@*e 7_��T�6"O��
P�}V�,Ke/L�9.�Р"O4$�eŧ0�CrMR*���"OF��1E�'Jv��Elڒ+�ځ��"O�q� ��� ��B�Ѣ"O:�&��3l����-�D�t��"OjIۗ�F2�ZYy��
r����"Ob@r-\���ѻ&C�3\o�`�"O�h7�Z�]�J�-��rr �"O�f�Y.2�,���z^� `!"O֬(�>n1�a����^:�X�#"O�ݘ!Q+�tx"�̠SV�:U"O��C@
��=����ba[3'��mZ�"O�A+fm�U���H5�	�-j6A��"Op�&aɝ0d4���4.�U�r"O�Ű�%غ>�".O�I��u(�"O���w��/�6 �Q�9w�
 ��*O`��3�W)@�0S��X�PZ:��
�'Tb)a� N�Fd0Y�HX)���
�'UJQз�ц�~�i�D�T�z��
�'�Y�0H1=S�i��+�K��L�
�'攴*#��r���('�N���
�'�9 �\.���W�Mn\XT�
�'�&�5�M� 8�) E�a�D�
�')^����\�I�@%Q$dL6R*~1�	�'P�ͲwU�����#.�;	�'#2��e�9.x�(�9���	�'�F�0�`K�M;F�ѱ!�n߮�X�'����B�5GuTb��O$gт�Z�' IcZ�#���dc�-9�'�"����T�D�6��(��c�i�'Y��z3 [�b��ŉt(E&��9	�'�hK48��AX�b ,(�ʨ��'���r����X�Ė&GZ���'+85HqdK�/�lJ��|4, �'��aQ"F�AshO�Y�T ��'i�5(�T(M5&�����h��	�'} H�#k��6cdXt�H�^
�q�'e� ��N(�F�ۃ$V
�!���� >i�`�\�l����#t�D"O�,R�N�Y�*%AEߺ""�HE"O�|Q� 5L"Ա0d��;Ȁ��"O윛1�/K$h��O]d����"Oz �tE����Pt΂-M��c�"Oq� ��W��A�t�Xw��aC"O�]9��u��B��3b"Hi�"O63 ]�2�Y�Q��<�~�
'"O6"��%gƼUp�C��je|0�E"O�Iۃ`�6��1�#>\y�� �"O��!p'S<
�����D��T)`"O�Y�Ch��~A["aҹ$���P3"O���Z>^r��!�4�|p�"Od�h��U�w5��r��}�+ع�y��\)]q��b�fԉ.:�A��U��ybL�73��,��Q��E�c�U#�y2�X�%�<��s蕂N�B�	�O0�yR�Ʃ9�I����Kx�q�+��yr���>M�du�A�@����`�A�y����E�5p�B_��d	ޢ�y��S�<�<�:���'1�И�ϙ�y��+P�.��$n��{,���Ğ�y�I"z�	���F����ND,�y�$Dv�Zg[F��i�tK̪�y��-�j1��W8>L��{As�<�G�l20��qi��3�D��k�<�5dL"� �RAڞ:��� �a�<�ć۝k���fi�����_�<�`눦6��r��_�~N�H#D��Y��71�lZf(Ӌ$�����4D����Q�s�d��?C9B���*O�QJwc �!�c� G;(�D� �"O���d�@��I3�̾{p1K�"O�I�a�0
>��sfG�(n:�"O&�� 晈;6��I�KL� n��C"OPѳ���<iiFYe�ϮvX�"O���C
�B\��)�i�~KR���"O��V.�4�&�[3�L+A�T*c"O`Up6��A!�\2��.F5�Zt"O2%`�cP)[d�4�G���C��t��"O��2�fڃh�r�2���"O�QKr�  \$tI�Yvp��"O��k�K�?�m���ށN��G"OFa��j�����K\	 b� �"O����n�;4�<q�D�[��Y�"O����,%F���h("���"O��mK�y��;�H�mP� �"O:�)u��A��]h��KY>��#"OLQpV�zF b�c�Y'����"O��ZĆN9g<ti�)�>���"O�!%@�d|��tǗ%p�F�jp"O��ӓ
S>�Ĩ{���OI0� �"OH	@2דW�(X�����$�D�"O�*���qf�����;$�JT"O��C͆4�z����B(
�P�v"O� ���F�jR�''޿5����"O|ȋ�i׹<��&,E.3���9�*O B7D��%x ��v>>l��'�,+��
�\�,1q�m��={�B�	�"έXU��7DP���FaİY�B�	-S�4���|al� ��5��B�Id2V�ӡ�"�D�jvME�)�B�I#8>^d��_3g����#N�ND�C�ɢ*�|�Xu����L���!�lB�)� ���Ў\��FT1�J�Kv���u"Ol5z�G�]8 �Ӣ�	z|�!P"O��J]#!��:��4d�`ˠ"O�]h�ȡw\, �C
�(XBd%�"O\���CK�o�Ƶ��#X�� I�3"Ox�s �ĒR��(ҁ�7�2��e"O�����<���Y'_�Ntl��""O�P�C/	�<��H�Q:jD��3A"O�) �hCP���)pU�4�f"OP��1e�F:��C�<B��K�"Oݠ1�Ȓy�^�J�h�� ��b"O���g� ,�\��նSB���"O��҅�͗(�"�I�&�a�b�c"O�@�c)����A��)$�uP"O*��!ω��Б�`�t8,q+D"O�HrB���4�*pz�U�M�)�"Op\q��(������%7@la�"OTu�#��<WH��A�&�C�"O�H�P��,"I(=�&�Gnm` �5\O<c��� F\ΔDH��)ls#t�����-M�Y8�h�'<E�=a�" �n ��	��ē)�tT�X7�L����22��+�"Oz����Xj��ʂ���D%*1�%"O�k©w���3$�����i�"O���Ř�(�s@_�n�PH�"O&a�Ƣʄ(��� R"�>I$)w"O��I�$[?&2�����.=J`�!]�L���{�dIy�,�;+$���$?@�B�IxI�D�$ܳ�B1r�n2��B��0�`Yz�K�P
ŚW΄;'���e����'p���>(��Y
�h�����'� a����-�,�sx�xCA�	T��y����"7'�2Y����I
�yb���\l5-�1�<�R�M�y���4^��``UVL�@��D�O��=�Omh1��ށ	�B��┑t�՘	�'(�0�OE6J�|!3��o���'�8j�J�Z��`�ҋ/m��	�'	�ݳn���r�g\.g�H��'��<bF��;;�yB,�����
�'�~hz��M9)����tL�<k���4�6�<E��4��X�q���ap��w�^6�b���V��Ṳ��tw�ɩ� 	�,�� �'w�~����'�ġP�D�*�� �ti1�yd��LlT�W��%3��S#m��yrf�%�P��O�
���ɓ�y��d'O2И�Ӣ5 ��c(�YHhY�U"O�삄J =\��jw��8��"O4!��폝'�t���?q)U"O��:�	� %�$MX�E��7"�p��"O�bq��Jh�-��O"b�1��8lOvIf$�1ی��R��0_�>�:�"Oq�7l]�r����(ԓ�l��"O�+ql�8b5��\�	k�lST"O�0X���� �ah�@�&n�Pg�$)�S�S�H��$�'�Y�u�L���d��-w�B��%7=D�ic$��|`VѩǢ̤V�$�<�˓;���aI�!k�����O�X~��mZr�����ɾJe�̻׉��L_t�M�*T!�B�I�i��'��:o�N9Q��'R������&�S�/&7��Y��M�t� &��c�^�?����đS��%.�0U��HdAS=U�OȢ=���+��F�F���9�,��;��:�P�@G{��Ʉ�n�}���\���੗)W�!!�� *�is�C 2v�a�C����H��"O&ݡ��1j��u����Q,����"O���'ݘ!㢝!��ĳ&~�0�"O��ą��&19��P�ep�ِ�'QqO��b7�#*{�I5�����I�� F��-~�<쓶�?2�̴Q`+Ă�y�˄�}Bh�; ��U�E(nN0�y�DM���}*��TS�B��m�:��d/�>ɕ(ȉ#PdH v�w�t��!Rmx���'6�Q#$m�5'x���ȗ|��
�'�n�9�̏���g�S<�-`�'���bN0N��V$���
AÓ�hO�Y��I?ߔ����L�N��P��"O�8%��	f!j�x�)Zm�J�t"OHI��� bJ��b.�,�x=�w�<)��3^z�<�jI�>�h�d�@X���O���6���*�O���0"�O���V0^�. �&���RDKe����x��I+G�R$�ǃ��rf��Pօ�
f�����?ړ3�"| d��X�*\��O�W�D8�O��=��Q�Y��Se]�wL���im�<@ѕ<�&��/2za��)XQ�<4i[���Ț����X�J֢�P�<�ǆ0&�<X6��9��%όF�<�4%֫_�
�Xm��\5�YK�Ɨf�<��Áx�:�$�خk�d�@�DDg�<	G��r��غ�o�d���h$C�d�<��MP�u�r	�e�"0��KS�Md�<E������9i[�|@�U!H�i�<�e$3d�pu���Y?܌�l�_��p=��l�"P,RW-��@�����P"m|!��-2ަ��@M�\f*M�7*ڿf>!�$�4��!!d�YO
��'G�u�ax��ɩRW$tIv�)/\�P�0Vc��E{J|Z�N]7
U�Q��Lt����g�<ɥ��q�!�����l�z�&a�<�g傆(�ĘB�Ol�p�S~��a8�X�0�����1��_F9xfl5D�)���J����!)�L�]�&D��C2*,F4��f�� �,"�M%D��s@�?��ئ��\���)��!D���B�Ȅ`�>���<����� ?D���A&��F��`3a[�L�D�(7-1�$=�O8e)v
�Y�T��I�A��@�b"OL(⧏D�t���i!Ņ�oG�rE"OͨG M�T�uX�L5���"O��Iӳ$f�Re��aD��"O���$��5�]���SF�ⓞ�����)�'P@|+��[,Xz��"�H�n�$`�IQ<��Z�J�{�v�Oq̓�yR��˽�����N���qP�ոj5����߰?QK�o������B�jQ����'�ў�'g,8lZSC��h���EA	Â	��z�r1�f(_ɀ��0�C� �]��aB2�b�_?t-Ճ^� (����Nܓ�2�s�	 <4�"�R�H54��ȓ,C�8�C]2p��!� M�wh� �>������Ĺ%���%���v1�e�T4�y2, �u0Z��e��2pt��'�Z��y"NM�b�)��n�c[�RP���yRo�!πAC�BQ�\2�=���۬��z���O�X�;�a\90צH1��?v�PA wI.�S��y��OR�(��o��o࠱� Pp�<��	]�^�̐;�Ȑ��oZ2�y
� @��Я�`7d��2�E�]��`�"Of
�
�v]��i��?�"���"O�t$��?�D��"�]�2p�t"O���EJT���e�B�<���"O�� �h��N�����/_2-�"O�i���,�N�@K�8�X3�"OJ�(�(��Ea�t�G͇8��B�"OV�P��E�a�H�`D�R��D@4�'B�$MYM��
���P
T=��GQ��	C}��� ܮ8�*	(k܅)d�
�"��#?����9�bq9Bh��z�n�JP矋D�!�DW�a�j���B|m��X���Ik��(��᳴�}�`i�7a�N�T<ɴ"O٫���$5`�̢7K�e&q�V�$4|O���qIS�z8�$M��1J�ٻ�O�\jf�֥����Ι+�\y�V+�q�<���	W��]�0��?I���@CBw�<1�HĘ=�µCY;4��d����q�<郩�2nO�q�G�m�:�C7̖Q�<�snHb!�G�F�I�f�L�<Q% 4<����%�\8e�^�p�f�]�� �<��B�#�l����� aωZ�<�
*q��5��D):}&��S�<�c �.O�B��i��;�Az���S�<)&���v���c&C�Y�V��M�<��d l��C��W�_k��j`q�<)d�FA��ɰ`�:,�"B �j�<�`iR�Y#b�[���q\z���Bg�<Qd�N�t��U�l��B���|�<��E�843vE8&HS�dx,(�@�|�<�#,\m��M�
=k�
Sb�<��͊6��Lx7�L���z���s�<���ܓ����h�6k�P�eK�e�<�W.V�0" /]�ءRTa�<�Ũ�:@$���,�$py��F_�<�,�%-�@�c�%ӥgth���_�<)"N����X�~�]�%�@c�<ɱ	�^ �h:G��,�������a�<�`o�{֤x4��e�a��_�<�&'�t~�u@`�sJ|�� ]�<i�ٕrv(���0O������V�<	q�J�4�����FF|�����[�<Qɯf�ze���Ϣ}��!OO^�<Q&�ӎ"�٨�Ϟ� 6�y��[�<qc5x���E w��E&WV�<���4&�AAԧ�Rf��$.�I�<���G�.fV���'�sB��Y� JC�<�B���J��	�F?\�03���@�<�V�Y*w-�q0�f�^)z]��IF�<��@*n# <q�%I9c�.����@�<!a�V7Bbl�t��7\{r��PGD~�<�����ؔD^�c�Ґ��"�r�<���.Y�Z@�$�A��h��Y�<�'A��v��t�R�������E~�<���Y#)���'��[�6d�ՀB`���� C.s������A�A��$U�/y�tEo�vD|,�%c0D��pTm
�%�!O 	�U�L;D�`!q��L��=��n�l���Շ4D���7M@�!㢼qc�7d��H�p�5D�h 3F�+\�%�Pʗ&@��t��a1D�(Y�nK�@�\���KI��m�6�,D��Y�A0F�B�G*`��m�b�!D��� .�]_�x�GG:R�����!D�����j�Z��@�ŦMg�M���"D�� <�%Ă&9��@S��PR�,T"Ol�'�ɂK_�p���f�X��"O@��f�.i�-u���t�[�"Ou�'��1zB7��>7-5ch<D�p�d�Z���P��F)x���4� D�X�w`ZJ�6�{��P�eh!���?D���I]�2Gb����<P�"g�?D��h�ň�G*��k��H�<)���=D�LrV
�;�j��3J�-~�8Y� �,D�h�6��G��x��ɉ
�5�tC+D��J�;�D i��ҿ7��H���,D������ �l��A�ʔ�DN-D�����E�@!�{���`9D�`�!��f���K(1KxT��4D� �7A>z�dx��:`:���*0D���ׁ���qr��@�PP�E��1D�`�L�
��d�/R�C�`�@#D�|aE�T6[U��y�cѨR�FoH_�<!�N�-�R�8�K��6�ȉ��_�<�p���	U�t�TMԩkI�qh�b�<�c��2lݾ-�E̓�os.i�b!FX�<AEڸC(b<R�٪]��ђ��O�<I�
@�b��\�%ګ%E$��E�<�%�ٯ����WbZ�r���KR`�h�<�	[n�<x�e��lT�i�0� k�<����I�fA�5��G�p��b�<Y'�J
Y|���RA���A�\�<!E쟒K���7R9�N�j��C[�<y�n�%Hm0@�Ζh�T��g�Q�<����SJ��p �N�n���*L�<aŇ;M���Vf��L~�u!�L�e�<����t���U�J�DMPSa�]�<�u�����'�J��z1��[|�<����I�De��0x���Bn�P�<���[�	�f�t�W�5b��S�<Q���7QVh3���$.�H,2ap�<��ƪ
K`�r�N'4�F�$�l�<�q�\>O7����TV�Ԭa6�Ak�<�ЅՎ
f ��̢lv΄�QO�f�<a� +>�P��L�X��H2�T�<y&�=8��rO/tA@�W�<�r�#Z[\ոf����-�UI[L�<���=t������;Р��L�q�<�v.C���Bd+Ĕo����g�F�<����1O���)J�Q2�A��F�<1�^��miA�R�r��q�`h�t�<��ˎ�F(��.��A@�����~�<)GBZp����=�^=���u�<c�
_E�ń�tХ;�%D�<�φ8wV������  �>����F�<�Ŭ˨J}��R����"i�ت }�<���&M����gE����b%�z�<𯈆D��rl��Z��*礝r�<�׎^#1cFT��K:;a��za+�i�<�CN���Bd�� Wm5��f�<��H�V��cA
ʊ{6�4l��<���U#	φ�@�(��i-d",z�<��H�:I�=��	4�pxA0!J}�<��k��CZ1#ӏ�dp^�#�$Xx�<���$wɰ���I�1e~�\�b��s�<ِ%ҁ$�R�b�造h�l�$-�@�<��I^�2U�܃�a��K�6ɂ��B�<��ˑ(�Jrf��lS�0��Ww�<Q���L��i!(H.F+8�3!�y����Q
O�H �T>O� ,		�/�|�����D<4[���"O��x����Z0�%�a�ϑV3J�2#�O�T6@�s���E��}z�E3�I(�%�;#ԡ�#�Q�<�2�ξt.��{૜�Jh ) ec�5-���s�b[���d����?�'R�1jdM�6j]Ju07�\�y�p9�'�"���ȕG)�y���MC���F�B�JĔt94%�2D��	(S�Q �>d���bZ�;d���Dſu|��q�[�=n�$�eO�WtI e���n=�ĨţgC:C�	�k�`�uÆ�z�f����
��Ob���L ������A7[3h|�偠.��3���'f4�Lpg�Y�<��錸zZ0�W+۴'��ƍ�?�ڸ{a��2{��Y�`"Q+h����O��A�O��9U��=Kk��1BOLT��L,x��q$��8a�� ��*S�ƠY���B�*�CV��ٰ<�#)�{�����:WK��U(ax��A Y�TL��%h":�F\	C��?3�b��T��eC����1�':T;�㊗[�*�s�Ȋ\z�њ�y��^���@÷U0�P���"��~ b��ܫq�~���C޺;0B�W�V�����,EA.%�rCګH�P`�*��f��2�#�?��!�gy"�U:���qw�L>E��aY3%�)�y�� z(��iB�a����"/�4��V�
}��"
��ٰ<1e�D�#J 0s��H�;��"��Cx��r/�P@�Au$I�6촥���K-���"��V?UF����B��D�E��w��̣���),�}�(��J�p����O��x�2@P�m���J�)J$Q�(%�˓[�>%)��3�dת��r⩃25pj�c�H�I���N����{��	E G��q̓�6a"��6���dw�'n�lHэ�C�S�R6��5M��:�1h�HI�}�t��'ptK�L��i��y"�!��X`�]�{�ҤF�O�rFqO��G�x�6�K
�rEn�9���9�h���A i�VI�f�Zh�B�	�:i�]��ʊ�L��h�b^��5^���<�u�^��<� �$�S�zǰ���"E!7�|��֬��R*z��Ai����ٻ���Ho�}�iB�}��	�u+��m�Z `���C�x���O?�Y��^0F�q�g��0`���gb�Y~�X!`ò5j�O�2I��G����9�����ǕdZ�@jV���D��?�p��G�2 Gay�/�$褐#f�h��QC-��2���Aq�Ί�?���N7�ȼK~n4i��)ǆ^30+�E8�Iٙo�Y(��hE�vL��c�~��؅a��(2��ܔ������ǣI0��4� ��U���)��O�S-���ˌ}T��S��-��"ж��)G IU@ �&����O����ƁM1i�☙4b�����q �o�����h� hl��ȱхW�.Hjp�� ��)�����eB�-�t]A���r⬐����>y�kJ�%޴C�������=ڧ34��r����`��Ƞ�C^o:%���h)C%ć���|���j�0�q��,'<{��D�Kޡ��t�H��P�ñk\��<���'+ܤp�	�4�li���լ^dar�G��9eC�v�����Z:S��<�����������a����L^�@�!�j\�<u�	N��8��	� ��S��Q-�΄Ӥ'̺)���K�,(ҨO���	L:Hqژ�h۾a����+qݑ:���	K)�J�(ɘ|z����)�r����-&��ҧ���a�D�GiպO���g�:�~2���Ť� )s�!0�Pa2|��IV�-���DK�@u�=�r��([�I$[�z�㬙U��8�CA��#e"��Z`��B��y1 `(�N�1R%
͓��N*�T�O����+�P1��4c�lk1�2V�\=��B�#?��܄�ɫ'3�e�#��/T�3Rl
�X�%�t�*{ر�0�D9&̶8�% R؞|��϶9��D��Ń�U��C@�%��x�#6S*�)���<qXt�Xwh��r��&�*@+��5c�h��'��"���"x�&I� aHf|�ҫO�s'�J�Kp�V�U� �[w��]�p�	ٮ5�\����k
�l����	�a}2�ö$)��o�=���)n���zSn�O� ����"�ژ�vH��5�Ju�t1��$��äi!�&sL"��P*V7x������Ybѱ�����u�h�j0)^	�f���^�)��Eak���``L&�O����f͏Ln���a�+��пi�Ԁ�!)qܓ|l��Ф��;[|��������7�MA+���k!��8	�!�D�%d�����
v紁�1�)Y�	�]t@���܌k�@���Rr?�����[���{�H6'�U3F�25������fm,8�U�'�����S�dW�S˃Yg�Y�\Np�J��Uf^5����ݪ9��`M���懬�, F{"(A6k?�  ��5dW�?�Ą��@�	@\�q(�_Bt1���m(�E;� c�d�@#�@�9mʥ�ȓ;���n�=�H �b���͇ȓ}�i�2`_"lP%Sǋ�"��a�ȓC��h ��IWR�qm����E�aR�ܢ/rm+$e��ni�c�d3d
r�S�'O�dx�2
�9'刵��'3b����J�J���[$4��fb�2'tԄ��{�Y�9mHc?O�KcZԩ��9�T1�DO��Bb%̡e����H��Wy.�3g�!]� �	�����E�D\� ���2P�^��	0��T9��|�Tz��	i�(�<q����/۱�yB+֑at:���۾Y�:�f����|��YhW�"�)�Ӥ)��48���x�,�ԯ�=M�L�>�b����H�Z9P6IvC�2�\v��;��5�	�9��A��L<)j�%K��Z�,��>��=;���<�4AZ-Fʖ㞢}���ìb�.L��؏a��x�r)J
?y6�:�'����F�.R��t�`�/�����O(q������=1A*L"lD@Ae+&��X
6 <�O$C�.LPa,�z���t]�a�� =��`S"Oȁ�"��$=;���
��A�T�Q�ɹ3[2����S�8���㖫D0Q�&�S4 $��B�	&>��I�:8}� ^`p��&D�k���Ӫu�tDb��wo�0���VB䉂H�ԔyDM@p!�T��)�%e�'�D����'>��A�΁�V��]�/��9�'U�LK�ح�P �!ȣF ��'W"��"*�<���Z)DR�'$|��F-Y4|���J� ,B��
�'M���iE 8UL��)�-����
�']�n�|@�pF���.���A
�'�@Uĕ��0\8E�@�	�'���f�
 Yֵ�'j��`̈́	�	�'�(���HѢ8��E��ɘ6gˊ��	�'�V��A��/m��}`@��+X���'�~aV(O�#���T�"&tL{
�'�R	�a��&x6��P�T�Od,�@	�'c�azcW�$ڌc$?g���'�%�bnZ2Q���!��УF%���'pl���&KDi����Z�M��-��'\��% �F�j����,1`j���'���h�ꅀM6���@�A21
�'�*���I\�zP��x`����'hh�	Ѷ&q��fO5m$��'Z��L���T7��~p���'g8���Z�k��H�N�I=|PK�'���q�VNi�� �\�K/���'!Y�˲XFI�u�+���0�'���2�g4<�����7R�����'���K���X�9��Vx��	�';�S�O��!��$��E��D�p��'\����%�HQAD�:iĽ��'4^�*�f�%��`�d@=��c�'�h�2fʓ<s@8ԃ&`B�*zb�0�'|�xx�m[�`�Fe&$@�}�
�'�J,"4	��T������zH�	�'�L�"�,&A�M��>��`	�'� y���S9,x�J �S*|�n�#	�'�4Y�.ۂ/[CG
� �jݸ�'��=�_�@��ܓՌ[)�T���'#b �1�L�����(}�X�+�'U���"��b�AH!H%p�ɻ	�'�J��C.��	�ZB̕7���'�u�d�(qR����
�?�jL���� P4Y���z� ��*�4�c"OX���Q|�@�q�gOF\�"O����'(4�P��
Dn���"O��Q��k' <蝥x(˖"O���0h�;A�rQcPjS�f"�q"Oh�M 0��4;qIü�f��"O�U!�FA�����x�(���"O�;�E������p�P<Ye"O�i.E1��"`��i��(�W)��yb(V�"�Q�p%��eG�P��*�y�#F>]O|�X$��k��daY�y"��o*�q�����q�	$�y�G�:����H\8�jЁF)���y���9S���@ @D��yˉ9=��Hj�A�u���h�� 
�yb,G}m�|����m�y+�j���y�DQ 	�:�+� ���@�2+�?�yR���+��9)e�Ɋ*�Ѳ��8�y���L@��$��_�������y"�� N>x,&�81�� �y� �R����&h*��r%�6�ybM��a�z�	�,���
�M�0�y���001��j �ɩ�Ht��^!�y�)�.L��7n���qvY�z!��� ��&hI�Dr1@���ڵ"OD �uDJ��n�rF��D9TX�"OfIA��G�n����@�9]B�5h�"Odi �%�_f�5���6I 9ht"O���S�	V�`���[9���"O�`�����l�z=���;4jjM��"O�D�q�� ����'�Q:���"O4���FصM{��V��Z
<�"O,�abHKs���`#fA3^D�9"O4����|
§�?}T�|:!"OX5붍��*� S��φ1��	�"O��a'L�V�8��wb�
#
��T"O��0�ٲj�����U�_ê�y""O��y����/����"��g���"O��.�in� ����2CNԣb"O��Ґ��c�H�Je(G� ��"O.�8���! ���*�g߀2�"лa"O���1��9{��i�R��jsL�x"O0�)Ba�w�l�X�+;hL��"O�В'��=w
A���!N�q"O|�yB U�Q�µ���ОJ�=�0"O(�{�ѓ�乢� K�0:�� �"O8Ȫ�.�01��ba@]�u=� R"O�4�۪,K�l ��Q�8<)�"O@���=xTD�R��W:,�h�"On�z��<h\^�iꁧ_�`�"O�� ��)2�@��>	�$kD"O�q����?_�����G�BZ!	"O��rU	,��@y6ӳw���Q�"O�}��b�+o<��oè>���	�"O4�z�BO�-L��ò��1(U*m��"O`%���%k&�fI	2�l���"O�HJ���l4�2aȃ��bIzR"O�TC��0yQ�z�
��-�t#�"Od��r�ћ~xd�G��*d� Y�$"Oָ*`'��vY@�E�m�
��"O�x d�\)��$�"����2"O��Y��AE���n�B��5h�"On���a�Q~z��5f�Z��<�q"OX�
 |*B�B��[�(�nq"O� 
�����a_Z�I'
I:O����"O�I'��Q�D(�tlF�{����"O�D8�j�*��
_ �qR�"OJ0�R*ܶr��H9���&	�J= v�'S
<��	��S��Γo� L 5�ز ��U���O����ȓ;�
���_�4/�ݢG����<�gٕ􆕒)@.�h��U�P	S�=G�aaI�,���"OTp
B�I�y� ��&�2��¨Ŧ#c�(��Ar?q��ė����	�(�"� � �?��s�)�5Y��B�ɄR�Z����w���k�n�T$q	���/e�h�)w�Y�4�a{�d�$g"p���`���B�ʋ��<a�c��f��<ʂK	 N2@ )ԪB�L��,2��Yq됷�yb"�A�~e��� y���S����!|�̻�#��)� )DIW� ]��ș��+��\���(`V�mӣ"O
ذuFG�48�@YV�D�(�6.�^kld�Cϕv4d1I�+��j��� *�xEI��84�U����S���Ɠ���4o>1�D�rD��:kʽ�u\E���C�
�(B~^���<,Oғo�VfU�3�;^v��A0�'WbA�C�U:]q���"8��x�oū?�<��Ff
!Ap@���	gH<�%(X�s2��V�HI'D�9'	R_̓I%L�w�\��U��g�o������!;H��d�Ň�m`7"O������N���D<��l����N���i!Ď�HCz����8�Q>˓?��$0v���� C�7R�R؆ȓL�.��u���v� �Ȏ,#9�	�'VR����	 ?����I�6�2}bT�4�
�{�O������d	*��hS��=�%s5B�AP�w�D�M�а��'"��Oǝ}Qf�7�T�YK`���������*�S?Ct4�0���d���1�̕�X(�B�IA��Z`cP)2��a¦a�95�����N�����ӵw���@�@D�I&
Bz�C��.70��ʴ8d5��P5��ix�BV�!��<�Ԥr��q��'X��a*U�HFx�d:-��KJ&(��ؒ?\0��	7]��-���)�!�@/hjX�Ɂ!"Vq9���x�ў0"�ۅFpR@�iD;$��
R+�v�-�P��Py-ߔS,{���u{�����?Ya%³q�pa�g.}��)�-�D��4fѪ}�	X�a��NB�	K¾hj��ˎ0ӄ�1q.�Q4*�7]|��欏�v����I&0�q���[�dy�c��Kr���)mL�Q�� p�T�
��?@|nA�%!ԸI��5$��Y%kJ�z�����X���,%ʓM�^�	�+�O�v� ��cCk�65���ϥA�Ʃ`��A�yb��j
e��J��-�&��w!]�a ǢV,�P�Tk�<E��{��2@�O>i�~:cV�#�:E�ȓ��)�d�
V�;��P�`b��%�0x��];�� ��	4S��|I6Ū�z�s'냝'8����-|��h�->-�C5e9z��4���V#����'`�q��H
`�ҹk�7J��d��gh�Y�F�H��ЁȖ�R3�:���aÕ�
�bU"On��bEX����F ��P���,S�<���_h�S��?�d�
��d��n�q� ��$�EE�<���D"02�[zZ���/L�2�f���+P��p=��N;��h4H�!8���I4�^}x��Y��=+ ��I��3���sPk�-m�DۇFC��yҍ�My2�x�M�-y���#ϔ��y��,�e�w@
��HSJ �y��N1\�RѲ�+�� rU;���y2o��{%IQ��ĉ#Y(�
���y2���m���Ƒ'��r6�A(�yb�ͪ��Ii�CN�*hF��y���!26����:�^���_��yҏ�7V�0���"<>�����yNA
E�p9[GE���X��Ѭ�y��fyj������������y
� x�:��UEBXS(��%f�A[C"O�i���0t����
7�9��"O,�9w��a~��1���7.��S"O����E�kA��02���hj���"OF�yC�O��@����i2 �b"O��)�$ӿ8�Lh��)Τ�v8)'"O�pQ��>P��-P���v� ]r�"O���5��{R���(�*�Г"O
iE��1��L=(n� ��"O��'c	"����E�(S�`"OZ� �ɥa�금�Z'8��aH�"O�!����8�p
׃R�G�B(��"O������<#צQA���x�|e! "O�ux�oߍ�.=�t
@�҅1�"O���ѦC>b2���I� ���+0"Od9��M�faSëQ3AvP�U"O�Y�7��M�P��ɗ!cHFفG"O�mz�IZ�hab��'H,���"O������?xP�;�$�~0X�V"Oh�+5��& ��=iƪ�;��!�"O�Q�L�&S�H ��pC�-"OP���1 8a�TM�DVqa'"O~����Œ�@!��˺2;^���"O*\!���(l�h��6D�]F~
r"Ox�'�3�ƌ�a�϶?$zDi�"OХ�!B��@$#���ΩH�"O�ЂvC���#f��2R��Ա�"O�z��K�g Ir���0���"OH�c� �$F�FE+�\<`�Px��"O ��&��'��dT T���ӣ"O"�K�#������C
�0x��)�"O����ō?!��z�L�v��iʰ"O� �)w��p2s�F���,��"O`,AtJ�s�fX�e�؎D���"O�Q��'���R�J`�q�"O����Ĕu�B����' ��xQ"O���eD�M��|r�$_W�S�"Oj|e�CT��L�0ZQ�83"OF!�R��ba�=���Ӛ=율�w"O01�a�Ϟ�Q���X�-�2�k�"O�-jpف/�����L��&AD 0!"O^�PE�(,j��Eʑ�qZ�cS"O�	���m ;���gJ�p"O�l�j��76�#�ǌ�^����"OƈQ�KG�8�Rw� z����D"O���͌=���)�Rh��"OjtY`푠Fb�i��<Mn�!�"O6�B���Ij�	C:R_��3u"O b���-���a�BXP�"O�h(����'` ���W3�x��"O�a8�D�N4�<����5N.��"O��0��
�/�0��-M�7
Rl;�"O��;����]�H�갫ʿI�ԌA�"OHH��D��=@y�ə�`��9q�"O��#2�$H^i���#ZZ����"O�l7K̝L�3�DTF���A"O��3&a�4�&I��$��9����5"O%ۖ(��kF:�7�Y՘��"OPU�t���d!�,ϔC����"OV�G¨x&�z뎶k�`PH�"OxTr�<x���z��Q<A~r��G"O:�e� �jlj�Ɗ�S�b$	G"OD����r�R(��dҎG��A�'&�y0�X�r��y�����o�~�E���)T��5 ��� j�P0�Q/*�t��E����k�"OPm�^�F�����ʰ�Qˑ"O*�ki�Eپ�ա�4ug"O�ze��0B:� �t�g0��"O�k'hU,�*H�e��O*�1 "OX�5̃�+bl�aB�A�p%�He"OH,���Wa۳O�4*vX��"O*;��D<_ |`֭Y/��E�"O�ضd�+\��c��Z���9��"O֭���ƈm*,�d��7�nt��"O�I�r�Y�-��H�#,�Ӫ,	1"OP����S^H�)C*C�G̲ ��"O@�D Aff�Z�������S�'5�Q-�2��ԃN�Ʊ���O>�����3]N9��y����c�=�Į�а)c���%(|%1� ����I�KQʧv������t.B�%�7N9\fX��hW!� 0Xa��y�@ƥ<�t!������ �EŊ�pP!D�|���S�D�$�dS�O��\+k�̫��Oy�3�"���= p�T1w|��˩O�� 5�A+����s�N>ݢ�.O,c�<�(!���6����c�e���u�ا$��[�ƴ<E��?i�B���L�aN��H$!�1j;P��FĈX�Fy��>%>O�ΞuC��г���6Ԍtb���1
��N(�S��Ms��ߤUO�m�����wG��s��S�<�AG�"���Pa]�jl5�D�<��� %3�hda�6hn(4����|�<a�� N�m:�K�6�D\�$JQv�<���%<8;��4�ș$er�<P��	^�r� C�UB�B�z��j�<�#�7Gu
�\�OB��r�L�g�<y KO�b��U1�K� X��Ȃ�d�<	G�~�ܸ@,_�} ���GCb�<�a/�z0R�6
��h"� �V�i�<i��i�tA;d��Rt�B�g�<�p �?:�J��%u��"�·I�<�����$R���<�� pS'C�<d�WlQ�q�%��&�т�F�<���2w��$+ch�	H��0U�n�<�&�"�,���I�0D���-�m�<�v �%7�e�DX�<�(�M�<y�36>�`��*��4��$��gT�<1/@�q��p�L
>��Z�
R�<��l"��P��
��0���O�<f�65r���3��X�d�<�`4m�D�iZ�7�nl�V`�Y�<Y��_;X�r�b�_�M����!z�<	FQ������C11&�3��t�<Q�H�Ft�,ц�� \���c��W�<�ĵxq(�k5�N#v��[r��T�<��� ��D	C�8v�����PM�<�蔋@ Bi�v��2��0��`�F�<�p��,�����eN�z�
�]�<�DnTO- <�Tg����%�n�<�1�%@T��u@ϟX�B�4D�t�<��dƥ(����jݗk6Iba�YG�<�/_5�LtٔFUV�Vh�u/�h�<q�JL�[�4��bgNw9*H�r�f�<��"�pPx�#��6|Z��f�<y�$`ɧG�	TdX#Fm��&GC�	�H���a��"|,��u�V�!h�B�N��i����7�H-X�BT`��B�	�Jڙ��)�>{z<*��\�b�B�	���y;��ώ���p�؆h2B�r�ȔC @�G������V�8C�I����5�@B��X`#/�C�&��Yy�ќ!���j�nZ�6B�)� ��A�+� ,�tz���*��e�2"O�= �j�*y/^1zSB��,�Iu"O$���$T��yGǪ7��iR1"O�lJE�8fY��E�A��x�"O*�S�h�0r���#�-ն\���2�"O�eYW����[�@�谹�"O���p҅j%�Ask��r"~=�"Op�4D�-Z�ri)#��)=��(q"O�e�b�6�4H�P��JW"O~t�p�J�`:�G[?)���7"O���%�[l�3 HT��n\#�"O�[օ<$0�p�#)�(w���F"O�{bNݤX�*] T�V"v�5a�"Oƭ���ˎ~h�Q!!��Ш�s�"O�у�'�@O��� ƌ�Q�p¡"O$�@ ��4�p�i�d�C'P���"O��䛥!�,�!D�f�,݁�"O.���A�C1VB�)6%��"O��҂C�37h���߬R5F4�6�4D�8��
W�=#Dmk�A=pr���4�4D�\��b�?lv�g��A��R�=D��8���)Y� ��- YVe�O;D�d�w�Y�ІP2��*`��Jg�%D�h!�(I�4d�C��J5j�sB9D��;�J��N!`�*0*�F�!�4D�$��-�0 q���"͆2U�X<2��2D��A�Ǌ�P�Ӧ�Ĝ9�U�2D�t
���I� ��;jZ©2D���ਆ�U�cW'_K��px�H1D�xK��1t�a���Z�g��d�U�-D���VG�#/+Y��(�f�t���',D�`��!"�X�o�o��3s�(D��!�Ԏg�	�i߆\��H��#D�*�j�:56x�9#��/G��!2� D����鈂S���:�J��>TP?D��0u�@�s���h�@�8J�4��n'D���P�2p�,�$�ɍ(�ihw	&D�\R"-^�9����,�/w��y��0D�<��BH68��5E��+l�6�,D��(��D8�����
[A�A`�$)D�|J�m�$TZԃ0�M`�h���*D�@!2H� tT��ҁo�3-
P�p��<D��C�ȅR�D��@�$�^��=D��Cf��>0`���oVI�,��ă9D���R�zH�ݘ�bV:,Z
H�$#D���#�P�5���I�f�yC"� D�� ��-�xYÒ�)V+����?D� ��.D2L>~0�	�t��lI��=D��$����)Ӕ%A��!��.D��@	a쐍�щ̙Ld��Ʌ/+D����bW�76���I^E~�9��)D�L��i�v�4j�3�B�3sl<D���pKI�[ $ݱ�(Zi� 0�Q�-D�L�bܳ�Px�B�`B�6�,D�[#��?\F��Y��ܣ@��i��/D���mӖH��I����qW���q";D�P��.AU�L���Q�g:r�ҳ#7D��@v#�z�f�"���!�@@�'4D��Pb��� 닚Ah�8�d=D�Pi1���1�j΀L~��@�5D�4bd�|��b'�f��V�(D�|�v��p(�K��@�~��x���$D�� U �h�0x��k������>D�,�œ�>�X��T�]�Z�:�k'D�� �4�FfW�Gb�q�P�6�~�"O���A%r" �Io�ȭ��"O@�@����Y����`IݷL�Fl��"O�x:���5V��xi�!�FP��0c"O��tB��{VcG�
?Q:��B�"O� U�X�I^Aڑ/���}[�"O��S�M�WR����m��
�If"O����b��R$��7�TG"OJ-r ��X���㨛�>I�C"O������'g�$H`j�:]�P ��"O�9�`��0��d� *��\"�"OF}{�`D�KF��B(ˊb��`9#"O�����V, �����l���ea�"Ot��taXiN���D�|��"O^��Q��6�:1�m��P��`�c"O��BvF007�$д��S���a*O�̰D��_(��A�ř��� �'�t�x�Fʛ��4#.E�NH!�
�'1�Q�%I�b3�/L*2�vT�	�';����3:�q#EL�5��!��'[���԰\�<�+�C�1�����'됴c�䛖?v��5D1q�hk
�'E�@'�CK�8��^2%>�{	�'����,
�REQ�,ϣ�LX+	�'%ҬSA���!�R�Bf����H�	�'�R����:CFe#V��LE��'�z5�u��3\*����I5���x�'\���M��)4�����4` ��'N<��K��K�Y E/�+_�͒�'	���WZ�H�d�^%Ge�@�']�6$/Z4�KWc׿�((��' ��H�J.!H���FH��>h��'4��m� ���~"�9�'��t�DC�{�&�p��D��j	�'ǀ5#�/��hph(��L-*���'`p���j�>����ޠ�0�*	�'����"Y %z3�ㆁ����'Sp����"E�8��0F\�x?*lK�']�m!���RT��w��#B��'5n|�d�2N� ��1�H��p�'��ũ�C�lX��Q
�k�'�Q�#� u,`A���(p Z5��'	
�!��G�$#��)�'��j���
�'Kr*��N�̘0�p>��y	�'��D`Ӏ�l0\���m�����'Ry
Ug�F�؛F���j��49
�'�B��%*��M�8��fZ�2� �	�'H����V�r��ȣ��^!+�.�8	�'W2В"Ǔ�X��@��(&xpɫ�'���8p�׀W�b; ω�����'����q�P����Ȓ�S<�		�' �U��A\+�1�7".Z!�5��'��a$̒I�b�����GQDu8�'8I�G�k�Je�d*[�T �Q"�'���0�ꋘ\E�l�S&�G;��!�'���S�	�/�1Y�
ӥD|xd��'.d���,ڮ/�I��g9Rܲ	�'�R���>L�� 3+Z7*)i	�'r�B�hUJЙb�ʏUz�Pp�'3l�`��	ht|���N�G��	�'��p1��D�!(�QJكE9�e��'
4�©�9"��,X�'��]��'�6P�H��
"��@��%����'�hp�ŲP��� ,�
������ P �b�A8�=���� O���@"O����W&�x���~B(H�"Of� f��hz@���凈9�ݛe"O�q!����`R�IQ�5'�I�4"OHـ�/@�vIͻ��L!)��)A"O�Eh0��=����%g��a��]�a"O���Z�F����%FT;�j�K�"O	��(0�ڴ�_���"O��j��mir�c�C͗����"O�xB�`""���50��A"O�M�Řb{�y�é#m�T�"O>�� Y,l�VA�6�[�s�$�"O.-�� �p="�"Ҩ߶[�^	�r"OJ`S��% ue\Ӧ}��"Ovi�	�a� qYE�Fˈ0�""O
E�P��ti{u��.s���d"O�)�"�G
LҌ<��$ٲd�z|��"O���u� ����s$[�3�mf"Ohi��.�54�j��B�.0��؃"O��V/U�i�Btb�K�B(0Xy"O�PE'�;E��`���85#rp(D"Ob4{QJ	9||�E�΀���p"O�1 ����؄L��B3v��`�"O(��F��H�J����$\���""OZ ����,�,<s�ш�2�Q�"O���"�=V��I6���f9"��"O�)��n�fv�R榘�.Y3"Or�b��@l&e����2��K!"O@�ҕ   ��     Z  �  �  A*  �5  �A  RM  �X  �d  p  s{  �  �  �  ��  *�  ��  ��  �  Q�  ��  ��  !�  e�  ��  d�  ��  m � > � n  �& - f3 9: �@ JG �Q L[ �a �j �s �z -� m� m�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��'��:�aɤ,��`vcء|�~Id�=D��Q��ˌE��z%O/Fs�mQ�7��)�S�'XM0�UhR: t�3��UU\`1�ȓ���q���*T <Ia�?c�ؠ��3�� �W���TCԺ����d7�-{G�0R�
Ը��̳c����N
��
����J��8�2qz�=��wYu���'R��r����e�4݅�u?��+Qœ�M@\
1�W�1�؅�h�eI�*�~UZD�����ą�T���Q�dD������(m��ȓ	��Rr+���<�Aj3\�Q��I�}Ru��4y�v��`E��2�b��ȓ2�,a양^�d� �N>Bņ�Q����$�Go 4� ��@>j�ȓZ�X��%G�,�Xd��غ"t�5��W# Ct`�A���X#��rg�-�ȓnV�yC�U���x6k�[K*��ȓQ^@d�p����sVl݁oVr���b2X�3SMD�=f8a!���t�ȓ0����I�<�XXC�
�Q;���ȓ�"��w��7+�dȘu�ȷ���ȓ;Ҧ ��B��IT��(��D�꽅ȓ9قu1�f�y_t ���7v��P�~- Q&�Y�F4���-wq�(��@֚,@�ϔ.���V�`'p܇�l;��GD8!�,�w-J*�هȓ5��S5!O�tk���f�<z6�ȓ~t�i1C�M)><)��EJM��{�R} �L�j
�*3ѢM%r�ȓ"��\��o_�4�WbD(l��@����<��;-o��P��&>�����C �3�^�A� ۤO��X���ts�*R)G 0�pHb:�H��?y
ӓA��Pq�*K<T��@e.�'�r5�ƓydI��C� uj���� �A���'7�	P!H�a�������far���'?(��]0:|��F��6��
�'"2���a܋,��aCN��
lL�	�'�҆�;V1�@&� |��TP�'0���"#�"�d��e���'xv%;	�'��$�߸s-V�!K�I�����'i�}�# )�j̓��_�@2< ��'��p`��
(两j��0=l��'Z��)�� �K��{S�L�@�u��'�J�#��D3.��i���ՋlG�
�'�x��&d�0:Ȗq�f&I�a�fԳ�'�\1Z�M���h #L�	a�9a
�'����'�<�,��#��I�*(h	�'�X��7gNa]r(Kr��F^���'-����;�t��*ԑ6Y0���'���t䖓e����FD�y��X�'È�r��4f�� Yu�
~�Hq��'�$3`�W��б�1b����C�<�AW�Zo�h�5˞1M�xS��z�<����6 x�y�� <�|���d~�<��"J w��@Z?&�HP뇦^z�<�0!%B/���� ��X�'��n�<�DD��c����-�{���1�E�<����;-i���g��n&�pT��H�<)f�<ؠ�h�s���sb\F�<!ң)]ݬ1A�m�$gn��P ��f�<� L0�i�3:���b1o��O��郢"O�A��M��]��8�-k�l�v"Ort��
D8g�\T��̜�f?���"O|��V$�9m���a��%
6�ɱ"O�Ī��$$���2���D�l��"O��)�ce<H=b$ٲ+�� �"O����Ο�t+���%�5}ò�ڗ"O��4��M��A�#J��t���(0"O����*ٗcJ��p��d���s"O
�5����6�h8Wo���"O��A�&Jt�H*�%�"j8	��"Of�->5���Th�hC""O��w/�p L��g�
M�$� "O>�`U��c����g̈7�v|x"OƜ�� :�)�k��E���"O$��0��<,��H=�� R""OX ���9^�H\h`Ȝ4��xIP"O���!�Y5�`��D	�6��V"Oй���X"	"m��AI���"OV��Z�SA�!�Bs��"OМ(�F�����*<���x�"OΩ�X�ޙ�4gW*���Id$PU�<�V�O�~�	�d(	�3Ѱ�Ɂ k�<vCʚQ��ݛyu�#Ak�i�<���<&�8a���yf!0���@�<yG�t���b
�S��U�<V�['g�Ȝ
 ��Z̐��FT�<�Rɝ<Gt$�#͈[Wꭢw�v�<��G%)�޽�5�ϊj��ⱍ	v�<y��0E����i�{��pZ��s�<Q�W {�j��B��y�>(aFU�<��Ɩ�5�"D!������ÊW�<YGF�y{��0���8�ɡ�i�<YU��%"
Й B<!db�hD�e�<���;1A��ӑ�ɸ�@ݓ�JI�<!��Z2q�@�D�$I���p�<���
�T'�ٓ�Î,B똙��N�i�<�	A�sP��Sũd4����y�<! �v����L'��5���O�<q����BB���j�v�"a�K�<��#À:�Z`��dݙR
RIȕH�<�e���#��8� ,��`q6��A�<Y"ݧS�i{v
�D.t�B�NA�<!2��>$R8�'Qx���
��W�<IB�֏}�j9�X?f���JB�Q�<��ȏ%ҭ���O�d,�Xc�r�<�e˔.ta�'��!HvZ	��S�<QP�_�K�B-�W!ٝcD�y��GL�<�7���v'ĝ�%�ΩGwRB�	Pd"Lq�J�H���k"�� :��D�[Ԝ�yP�8v�T��:x�!�$�'9]�a qHС84]㷯G�	�!��[��� �fK�56Ͳ���H�!�$�����P������p��܇r}!��50cX ��!�=;	��ZUM�g!�D�%!Z�u�����)ԭ��>�!�D� w#&4��ȯ�t��D��!�$��]���ȵF�? ��ٺE@S<!�d��Qj�%�E��(f� اF��X!��	O��C�A�]i��q�H�<�Wg"��u�ͅg:�T��g�o�<qGO�1�؃D
߷2�=���j�<�b�l�N�L4`B�Uç(�f�<��Ά�!�������8XN� mH�<� �s���Z|Ä�R?T���"Od�ڳhL�,n��֮	&V�&<pW"OX��@�3�����n�,T�Bw"O���w,K�]�P@Q�,жx�2�PG"O^�B��D�L}�,>����s�'���'��'�R�'���'���'��Y�̊b��D"a��?�@a#�'���'��'��'��'���'�F����)�� 	�!�3r,|��2�'�b�'"��'Dr�'���'&��'� x*4m�<$��B�i3�'���'4B�'t��'2��'���'=��I���B��q	�-����M)1�'1��'���'tB�'���'���'?r�
c�KX�<��k��:��M�'�'���'��'E��'���'���'����g�6m��@��եO�A[E�'��'`��'�"�'[��'��'I�0�� �w;T�S�+��I)���'b�'���'�B�'-��'#b�'�m� \<~=3�
;��c�'/�'U��'W��'���'���'!f��HU�1��}��c_:�~���'���'!B�'W��'���'���'�ˆFQ��Y��L@�8�n!�e�'W�'���'�"�'���'���'Y6���NL-+�V�z�ɑ���#��'���'���'+�'�"�'�b�'�\sD�&d�c�\�e�l��'+2�'���'7�'���|Ӕ���Oҹ��ܽ�6	iT�S]!b< ��Ky2�'h�)�3?Q�iTе���z��,�d,����,�C����d����?��<���}��i�
�b��\���یJ�4�����?9��Ѫ�M��O6�.��N?����\ ��Ȩ��͞3�p�+Ql<�ޟ��'4�>�-F0�l홗M�rXP٘��Z��M�&�m���Oc�7=�\�{��͝Z���O��8�2&��OX�d~��ԧ�O��D�T�i�󤙑D�D�y�,W��y����v���e��z�g)�=�'�?�A,îu@�,k�^%l�p�`����<Q/O��O\�mZ#7�(c�����	��[���z��h�n�����ݟ���<y�O��`0��$�Ȕ;��Mol�}Z�����	�J�z$���(�J����ߟ|9�
 OD��4@��Z�&�Wy_���)��<	d��Y�0|+F��=$��xpr��<��i��X��O�-m�}��|��kĿ�ޘ��-p� I��+��<����?���A2f���4��$>���'�hacG
�u# ���۠"�]�D�6��|�*O���H�.��Eu��YR+BT]*Mᄞ�48ڴ(u�q�<A��d��s�]�D��:L��(�K%A����?���yr�&zs�T
� �y� x ��R��$Z�BQ�������U&���?i�o*}�gy�� �&�Ƞb�1V��/�1+"\�\�'*�'S|6-V6c�Z�:���#�ڇg�D����6s^���U�?��<��?)��L;�b��Jr�=�Ƅ�)��y��_��M[�O��$�����)g�����h)<a�6��7�TP��i�D�IFyRQ�"~��n�?b�� w��" ,�	�S"f̓�ƣ����$�¦$������q����2�)�@��0�O�<�O��D�O��ΓL�66�9?a�� �G��~�P!�VǞ#R�訉@�Ox��4����?qTa��:��Ab�/�h<n|�WA��<�K>�u�i�ꀺ�y2_>ia���b�"MbC��\F~�D�"?1V�����|ϓ��O�� 	B	L,C�T,�f`E8I2�1��'@LPJ�M����4��������O����I!H$�q��;"�R\�5l�O��Of���O1������H�+�N���6�LT9դ�
i�`���'��keӜ⟠3�O�0mڣ!tz�x�N��Br �i5���,Z�Rڴ�?�iS�M��O^<��� ��H?)8&!_� U���q��2���bs�Ȗ'zb�'G��'/"�'��Ӏt�>$��ň&h8x֙��fґ�Md��?A��?YH~Z��Y���w[���gg�*N����2J��tM� ��|�,�l�w�)��]e��l��<yW�^�J۔$���ƇU�u����<��-�"mv��W7�䓂�4����
2�\a��d
�d�d�i'j�e�6���O:�$�O0˓l*��
���'���kx�i!�$K]QST@LS��O���'2h7F��q%��J��]�u�``QkP�L���1�h'?��DY |��*`��]�'d���D���?�!�&E*8"���$��9r���?���?Y��?�����O��RT�=Ft>��d-[�Abfh���OoځT�u��̟`�4���y�OFW�"�S������92EƠ�yB�b�V�n���y��㦍�'��(B���?q��ڿ`	h��f�*	[3х��e*�'\�i>���ϟ��IßH���}�$�r��u�$�j�N�j����'�7�
:n��O`�d+�I�O(�`�ǹ}�L!�@+�R��J�Q}b�i��mJ�)�&��Q�P?������K�H�%��`A'!9?�ta4;����D2����dX�dx��>6��\�4jZ�f��$�O���O �4��ʓ��F�
�� �p� t�E��z�̘ �I��yb�aӲ��O��m���M�d�i/��jfnș;�Z�A�8���vMWL����O���#�H?o1�����{�v�N�� ���AL�Fy`ek��תRdnH2O���O����O0�d�O��?icFkK�M�ѡe�,���{�\����	ޟ�P�4'V��'�?	��i(�'�0\c��>Zv$jU���x� Ȓfn#����	��|:���M�O�ax��Cb�\]�`*غd�֭��ǔzRt@�� �O ʓ�?����?���./�e��\��	2�G�6{�H�p��?i/Od�o��3Y������(���?=��5��T���@"Y6�T�bT�0|P�n��I�M�ӱi�lO�Ӊ.��E���n��x��'g�6��B�ؒ5p���&M�Gy�O]����2_�'10r'��;84`�̆.cՌTy��'aB�'�b���O��I��M��T�)*�]��ӗC1�8�R�RLPxP���?�ƳiW�O��'ئ6��;�t@{�� N_X5r��E�Q:ʱo���M[���M;�OjL��d�����<��e����LϺ}�|5�r���yBZ�\�	ߟ���L�	��P�Oז@�F��$|
h)2k��N���07)o�6Ԩ���O`���O��I�|��^w��wG�h��֙	D��@�9H�P�sd�Oh7��q�)�	��4�07mg��XW�[�rh�Ss@J�i�^t�v!q��*w�<7��G�	~y��'��
dڹ�p�*����p O.Aj��'���'T�ɚ�MctF��?���?I�B�TZ4 ���	�i� ��s���?AM>I�]����4
���3�$O�T���d�����X8V{�	w��cb��p�l�$?�C��'�l��I,,Q$Hi )H��3���RMX0�I��0�	�d��x�O�"�*e1��q�ǚ�-�
 #o��n"�y�Tx*���O��������J�i���4��+y�5j�f�\F�<`����L�I���ݴi��uڴ����./Z"���'��X�/>2,�wC�{���.9�D�<A��?���?����?a�.($R iB��xT�������Iڦ��/��h�	џ($?a�	�J6���� ��L��Pb��)�Pd��OH�l��Ms�x���h��gPAcdC�$���#q-(��<)1U� �	�H��J3�'Ђ %���'��L��l��F�\���iə��\��'�B�'�����t_����4d/���,.��z4��{Dy����w�V��k����d�h}RE|�^qo��M3��;[ϊ�e�ڿ�Q�X��9QR���-�'�bͲ�O�?q1r����wk*�1�)=C����gD����'�r�'/��'?�'Z��T!���7B5�Ű�*�f1ۖ��<i��͠�a��d�'� 6M#���s��p���r����.��M�=$���ݴ@���Ok���b�i��$@��)6\���h�fU�q���#�l�:Q�I�f/����?q��?���d�H#͒��2�S5W�1 Ql�O��$�<��iKFD:�'*"�'�哣>[�I��ªTQn�ze���	L����ş�m���S��)#F�F���	��w�bbƇ��x��Qj���7� ��_��:>�"O�o�I�B�|��򁀓B'�0����:H ��I����؟��)�My��v�l	�U���|, w�U�5=�a��J�N˓z����Tm}b�h���jM���,Ð��8N�1���ix�4g5��4���Ó��<��'4�˓Y��{0K�;I����@́\m 8ϓ���O
���Ov�d�OP���|��;6N<�R�F<�����-+��-/gC��'�����'��7=ﰤ1���4�����Tް}Ғ
�ڦ���4;f���O�~0���i�����F�z �ƸO&��rT��<��ĩq@����K�2�OP��?Y��V>xx��ѫ
2�x��'%������?	��?�(O�nZ=dD��ǟ��	�'�D%����bZ�yǊ��x�̸�?��_�$��4����=�$�2��0IQ �J�L�#A�m���9��zF
(�~�&?]Z��'�~���y�b� �g�����N�6R�la��؟<��런��^�O.Ҁ`2:�ڒ�M:�u�0�ιO��e��s��O"�KҦ��?ͻ5_�,a�GZS~�+%A��.��A�F��F�j�ZElZ�ƴ�o�A~�*��C"-��%*	Ô�\,n	�7Aí[
��AS�|�Q�P�I�L��ȟ|�	۟8X��'K����Y�^���H�VyR�iӠ����O��D�O�����C�p��MȲC�?�fy����=*��'�ұi�O�O��WC�!e`t)tJ�;^:�Q��Ί��|�RR��(�eI9'b�
Y�IUyr�[Ol�ԣ���8��a��+��'�R�'��OW�I4�M[2i��?��l	&y���ǋ�9?fq�R���<Y�i��O�M�'3v6mB�uQ�4h,u
��8u���a�A�:�(��re2�Ms�O�<bD
�
1N5�������c�ɀ19��#�EJ��E0�2O����O���Oj���O2�?�a�m��}6���Я�:X��az�kZy2�'�7*����M{M>�������J4i�y�*���J��>����M�Ӻ����T�P�����oԓ�`1���ͦ8���d�?�d�a�'5�h'�D�'�"�'M��'D	!���b��F�i��'�2^�4�ݴ��I-Oh���|�S��1��� Wi��~
����SM~�>���i0�6mh�i>�ӗ=O6�Kt�Z�麼qPI�$�8��sEC=/�d	X �Ky��O�<�I:n�'���1d�c�(��{b�q��'B�'xB���O)�	�M��fW�+��d:B>1Ș0�5,$$@�����?�Q�i��O� �'�N6͛�+`�A��]�FȒ���ҤnZ��MS"�@��M��'^`C�j�(���|��)� Rh``�2m��hs�+?:ī�7O�˓�?��?���?a����3X��� ���Yc��SaC�d�o�8{<t�Iޟ��I]��ޟ�j���˄��2z(N%x�`ݫ]l�T�L�F�eӎ9$�b>-�p�¦�͓�Q�G�Y�:w�͢R♱{����zԪS3'�O��M>Y+On���O$ z�d�8'/�5��
M�ZTr���O��D�O��$�<��iB�{��'3ﬀ��&׾/�j ����v^B�za�dkyb�':�6��O^� 蜁#��]�C�T��H�ol�H͓i��xTL�mTI��·�?���T=+�KZպ�p�'&��p��Z�x0ZQ2�ז?`<���'���'�r�'~�>��I2L@ʉ#7�,:VŹ�bV���	�	)�M�M�*�?9�N��f�4�m;�mP,S��c�_/�$�Z>O�n�MK'�i�p�Ȧ�i��˼ ���\�%C�m�w�RTc�L����{D���y�����>�]�<�	ß@����������Ic�c��Da���H{H����TyR�ӔBW:O��d�O����d�{ؙ0
@�+Y��r3��CŌ��'�J6M��$�b>�� �K�a��IJ�k�^8�cI;+v���6+����`녱*����&[κK4�>ɔ�<�'��Xx�51���r6.�^���'���'��O��I�M��`�<Ʌ�-$���tO�5hv�D����<���i��O�ė'sR�i��-ϙ,f2�2aհV�D48am��(��Y;��i�I�Z�����Og�'y"���8 㝱np�dd�9�ԡ>O����O��d�OJ���O6�?�G�T:zNR`9��0jt��)�-7?���F�a����¦&���@,�?JHL�cI�m��I�v	�j��M�Ľ���'V�v�v���� 	ߣ3�t��$N���|�*��W�>4J�2�'�T��'��6M�<ͧ�?���?��&�1@��)(���
s�x�D���?�������m�#�x� �����O�%�w�@|�J�f�/c4>�h�O�̖'�i�1O�S�g5�x��k�N6 �d�V	4���xf��@���*?	����@�'V�Ӽ+���()#El�@�F��V�W��?1��?���?�|�-O��n��j`�[B��qo@�;
_�U�n��(&?٥�i��O��'Ǜ�D�0U�m�%�Wt�q��;PI�6��O�d`4�xӆ�,��z����OXѪu�U�+���S����	Ν ��u�"��?���?��?I���)�Pܨ�qD\�Z�r�B��%t��m�"~���ΟX�Ij�s�(�������[�U5ڥ���эmb��C�B "J�i]1O�O�D���i��$�e�(X�pa
(0^�R��ܗ4���ƕ ����y�˓	V��W�����r�ԣ{�H��G�\iĈ$�՟��	���	ry��xӰ�`���|�I)P}t1�Mǭb�d�i��
1A�4��?��X�����%�8@��۸,Gd�7c���L�d=?�!j���i~�a~��ۆ�'HL=�ɨu98�+5�q��W2]>�hR$�O����O.�D�O�}�)��H*N�l�)�q`�?Q'2��@қFe܆��� ��?�;Wy��G�ъ{S��9��(3,-�`�v�j�X�D��U�z6�=?YK1>2<�iY(~!�0�&fS�����!P��/O�ImZ^y�O#�'H��'�R-�=��}�0��%�챐�OԚ+���5�M���<����oZe�s�D�§_�B~T'��D�.���������j�4��Ş&
V���ĕ;AqP�K��8(q��:k�Ph�'���x��D����`W�@B�4��U?q9� ���;'� 2F/ޛ*���d�O0�d�O��4�`ʓ'���(��l�R�ُ��%�"������Ѝ�+D����⟬��O�mZ�M¼i8:]a񆐐TJ�H:0��X�hEٿ>��F��pѳ��	N_�d���1��׾8��	�P�N�N���8Oz���O����O����O��?]��>� �ಯ��?� ͒EnNş��Iȟ4hڴMl^�ͧ�?��i�'{U� ��04j�	S��1EN�q(�1�Ǧ����|�5�Fβ"�%?��(�Zd�@�JXa��I�&�x�A�O,Q(H>Q-O��O�d�Oځ�Ĩ^$:2xT�CE��O>B�i�A�OX��<)��iJ�tk��'"b�''�2h4��uM�`����"'��3��|��i56M����M<�'�z�㝪@w�TP���jT���@�8?���t�ߔ^6��'u�����<2Q�|��P� �@��6Z�`�ゥG�"�'r�'x��T^�x��4z���sa�z�M��Ԙ>�q�u�S�?��-����G}�t�$|��Z��c�Z�k �p���J,'��.f�A��i�"�ܟP��&��h����+?Y3��:Rr����HY]Ŵ-)&�A�<	-Ov��O����O����O��' xl���D�r��A����X!��iG$�hp�'���'񟮸nz�킒�]:A��c�߄D����6�MK�i��O�I����逼+��6l�X
�f��,���!"� GX&��U%o���K�"j�dB�	\y�O�R�ڜl8��K��92�h��h��f52�'���'����M�'�U��?I���?iEi��9�ݑr�\�R!^���'0�o��6�m��U'�lq��5_�� B MƑ	��g�o����.ldP��]z�d��zB��O,���Ae���AJM�&��P��ղv�8�����?����?����h�����P)vT���*? NH�*4���d����S#Dɟ �I��M���w����-�'�^	 N�3E�h�@�'z���eӤ�l�pA��mZ�<�q3�(:W��X�� ��1�)��sA�EZp%�/���<�'�?���?!���?!e� ��0Zf@�n�vA���H����ͦ�K/��d��ϟ4'?a�ɱ��@R��ۺ7ۈ4CgO�(JIҨOV�mZ�M��x�O��T�O"�Bʇ1ʐ�2� β`y� =a8|8x�O�e!��D�?��b9�$�<y��$G�
���_�E�:\P$ ��?9��?����?�'����e�&�V˟!㮐S.L��)VY����џ�Y�4��'>L�L��Jgӆ�mZ��B�$jߜ!(&����E�m�f�faK٦�Γ�?��mΌ*����~~"�O�) c��d�5��mRx9�.�y��'9b�'���'�r�	�52�F0Xč�ZBgbߨ+q����OX��m��n>��I�MKK>QQK(T�$���W�����H2$�'�D7M¦e�-9��l��<��%��9�a�f�8�H%M�jE\	#�%����䓌�4���$�OD��P��T��Lε1U���$��Yw"�$�O�ʓ0�����Vb�'��R>A"�*9�x"b�H"�FI�ѩ(?Y�T�H�ٴaI��j.�?ŉ�"�Ձ�ֿ;y�dIԢ�ubU�g�o�l���O��?��/�d�#��S
Z�D+�%���-9.��O��d�O`��<y'�im6��LF	bFH���@�4l��j���>�r�'R�6�>����x�����S9�&�;���Z�,�H���eٴ=�����4���g��{������_̜ ��
4(�xdH�ʖ�bb"�Iay��'���'�b�'%BZ>���ȗ�Gr�+d�
������Q��MS	��?a���?9I~j�9���w��Pf�E��P���5e��i���a���nZ>��Ş&�plZش�yR��|sR9�T+P����yr'��J���OybQ�������'�FtY�M }�) �S����r�'���'�"]����4g�4Xx-O��DO!V�n	�b$[�6.�A3k�WA��X��On mZ��M��x���U۔,�~����(����Y�������E0
/1�����/�ʢw��,�`B£(�ĝ��)@�L%4���O��D�O��,�)�Sf�9�*��2b-	�}K�M��ly���U��OFn,O���՟T��I��֟�<s=&M��Ń<����Ǯ+�l���Mw�iO�7���F��6�{���ɟ`Dx���O7&���
_�P�Daz���?�,���z�Ay�Ogb�'b�'��A4b_�m�G�E5*�����e�.��	��M�$k���d�O���d�Ҡ�k��� 6 ��ч��;+�9�'d6�˦	ϓ�H�~�(�K"�:9�B��(�y��C�~(��`㝟��t��v�B�g�JylY>u�L8�cH��=iw�1��'�B�'��O��	$�M�`���<aS��k����5�W`�����A��<QĹi��O�E�'�±igH7͕�
�P���;��@���#��퉳t�F�	̟�p�ݠ8�T�=?���տCЏ;n����B�/���1C�<����?����?���?Y��4��� �	���E0d�%�C	A��'u2p�t s3����E���%�8���2\��!�"$x��	��'�����f�j�p�	%"p�7�s���"_�Y�j��>�j���l�:��i0�M�`����M�	By�O�2�'b$vD�8��(��j�a	��'`"U�(�޴_8�+OL���|2���N!fX��
�'���:7�[~�F�>9�i��6��H�)r �=IAF,�0���G���^�R�B�!��1?�'/���$����rj��'�n�,��Ռ�-y����?!��?��Ş���Φx���y�'�Īb�F�"'�lJ�{ț��DTq}BO{�h��(ݝ >�F@։0�&9 cJ榉�۴R7����4�����
?R�H�'����Gb��,�:=�|rA�?f0��Xy��'���'&��'��^>�:�.A�p#dܸ$%ʟ��a$fź�M+d���?����?I�'��9Olnz���H�8�����+��ł3��!�?q�4YZɧ�R���ش�y�#��.��zP ��X����u�P�y���#%�	�_�'&��Ɵ��I�)sDh����+T����w�Y��՟x�r�̟��'�6D�Y�Nʓ�?��I�:��Z��ל+P�*� Ķ�?�+O���By��'��� %��%����U�)1>�8�	̜h����OJ���#ʵ����f����j4����g�0�9�QaƦ���H�����������	̟�G�t�'�`���gX�G@IC��Iq2���%�'>�7��5.)���O��lO�Ӽ�R	Q3T��)�E��o7�Ik2���<A��ie�6�ͦ�������'�ht����?j�h�Dg`�k��5�҈`��'���h�Iꟼ��՟��I�OZ�OW�|��p
�b�p�')�7܈9*�D�O��$-�9Ox\����:X�d&	"i�/�F}��b�Rl���S�'0�����*K8t"��O�Z�ph��I����'��e�M�ޟda��|B]��b2��=ir�P��?QI�i��F�����Iߟ�����Shy�r�.81��O>I���·o!����[9�|�����OXHl�r��<�I��M�C�i�&7��:"�`�hfd�;�Z�q��?�@٥�c����� Z 쁬uL���(?a�'Կ�Q��[q��a��[$)�pz�*�<���?����?���?q��mJ-q��� m)>�jp�E/)���'�R�`�U�15�X��ۦ�&���`k��N$�3̚�+��E�����%V�^<��O��	"s�i���)�� Ԅy�YO|�����3:p"��I�?��d>�$�<����?����?���mKp��fI$�pl��?����J��%b���|y"�'��	d����ߝ6�N�rgJԮ4<��`���M�'�i}�O�ӹ5˨�bEN�P@��+�ݑI���[3�k��x���ny�OC��	��'�t,�@��*h���9�LN�|$l���'��'�R�O���4�MK���:[��P�@�]��ǌD�(�T|�+O�@m���]�I��MK���+��K �R?�b�W���t[�F�cӶ�i��yӖ�)��Sa��|�-O�m�ʺ`h�)Rb�fr�Yp�1O���?���?����?	�����gG���1�!(�zSe�I搨lZ$ �d-��ğ��	@�s������k�E���J�g>���KF�V�vjѵi�
6��D�)�Ӳk�XqlZ�<YqR�e��Q@���y�h|c�N��<i����dǷ�䓔��O ��ѽ%މ�`�k�X�k��M�`V&���OH���O��@��F�Y��'�rm)G *�s�VW�����_'-��O��'�(7FئU9N<فHP8*.�(��Wd���CJ~2��8w��@,2w�OR����2:ES�r�8L���.�����(~�'n��'nR�՟ 
��
�&h���S��@�P}�ST�P��4Ul�y�'�X6�;�i�q(�A&6��xU�ہO�>M�$s��z�4_����s�:pQv�uӀ���y��K��4�N
�%V� U`�+=D(L�Tg�#����4���$�O����O���֣E���
 b��/��:AE��8��˓C���%��yr�'�R���'&�q8p�I�Qz�\s�خ!*D02G�>�շiq�7E�)擘`ZB )A�^�ZX�a�BR����H�a��v�!�Q��O���M>a(O�U6L'0AT"� �D��!�O����O����O�<��i��5��'�4 "g/U5@�,�#��Hr�B�'�H7m2�ɿ��P˦�c�4{���R�$&��BV��(��#M���3�i���B�6���OJq���NL�j��a�)�
ˤJ Nݵ ���O����O����O���'��_"��+��"����H��I���Ɍ�M�2c]~�"d�t�O�9
%����!p1��|~I����c�	��M����D��Is�撟�sT/��l&�@biZ8m���Jw�_�9���^�M�4<�d�<ͧ�?i��?��^"�j`��Дh(E�T�P�?I��������:Dl�(��ǟ\�OFLŰ���6 c�B;V0�!��O�X�'��7��A(H<�O�J�kt�P��ÕI��a%m/S�J�b���	>`��O�	5�?��3�d](^��8�j\Ėc��Q  ����O��$�OH��<y5�i� ���\u��b�gRVʠ �G�y��'"<7� �ɝ�����}�G�Ǜ]�Dd84��kOjM8��'�M[��inR���i���]YD0��O[�\����.Ց[V�p򁠗�2_"H͓����O���Ot���O<���|򖠏7o��d#KT!bNz�"�i�)M;��E lFr�'(���d�'q*7=�<e��dd=\т�)C3��l+�������4U����O( B��i �;j=��42k�XQ���5���1�$��/�^�O���|j�HM�T�t��4LA8�a�
 3��i���?����?A*O��n�NW�<�Iӟ���w���F��U3�	�E��4�}�?Y�Q���޴��v8�C�D$�@�-�`�`9��N��I36}`%�A��*�b>E���'�t��'>%�<��8�N�fCJ$��(�	㟸�I���	w�O�Bg�1{S&�q�Y]�����1}!d�dm������ߴ���yG�˦8��$�ӇD�S��U�F�Q�~"�''�FN|�����{�x�q�PK�(�(���]�Yq�9�D�^�GSv�r'����4�����O��$�O��dO�18��c���8G�y�&ʙ�u7~ʓ=ћ�+	��y��'�����F�$�;#j�&B���tm��
z�ɩ�M#�i��O����Z�Ӆax�b掍����gc�6l4����.+�	�m�j���'RV�%�ԕ'�����:���e�7l84���'�2�'����^�<��4'
�T���Y`=��4hS�"{S|d̓+{���D�]}��n�,AmZ�M���^@�c�A?5}�`r�J�Z��X ش��$�� �������O�G�Y�Q�f0�0��� K%`����y�'U��':R�'�"�IKD
x�LL�<Υ��� |��$�O��D���YX�f5?��i�rQ�D
t �ZZ�!:�C��Y��Y��D�&��M����o�H��Hl�l6�e�����@S�lk!�.HrR�QU��?}�M0�<��'UZ�}y�O,�'���A��6��%��hO��(��'�RX�D��4B8�Γ�?)�����Kn JN�/Q�Ԅ� ��I	������4�����O�����C�+%8�s"b������A�K�v�Q��������H�8��pF�Ox�3���Nr��A!�7J)F�E�O���O��$�O1�l�|r�&��O�>��FC�~B�p$MC1��E��O<�mZt��%q���Mc�e�3V���c��*/��i��N:Y���j�
��d�r�|�	۟��B`�C�dd.?���ʧPl��'�ě.lHi��<9-O���O��D�O��$�O�ʧOV8p&'J�Uܢ����ݎ�Nڦ�i��C�'b�'���y�Ev���dopy�	�HS��qU�(#JX��I����I>���?}���N��n��<� �<����N�ܨh��q�!rp2O�H��Ȋ�?awa?�d�<�'�?	�?2j*Lh@�N!t�x�c!c��?���?�����֦ys�0?�������F'S<�,i��ݿ2����C�>�e�i^7��n�I"Z�����s1�!kEÌ�I�v�I� 1W&�4 ���>?9��1��Ĝ=�?9���%�� z!A��ް�4�V�?���?	��?���i�O�1Ov,���ƌ��Y��`xr��O��mZF��A��f�4�0��ě4O�,�����B���s�8O�Loګ�MCd�iG���i���Od���<��D�1%��qB��.�l�"u�^֖�O`��|
��?a���?��aܔ@�f�x<}�4�9�X�/O�(mZ�S�������D�s�DR��ťP�ó���U�ָj�����@ަIPݴRL�����O���aڍ<�.� '��#�*���Ξ(4c�!�����$�={i������O��{"H����Q�i{*-�m[(�DmY��?9��?!��|Z.OԌo�Y1��	3!$R����*4�B&H9D*~�ɮ�MS�⎷>��ie7��Цq˥�32fV"��-L���;��
$�$l�Y~��\�*�p��SZ�'��Ѿb���G�N�Y��u���<!���?9��?y���?���d�/IR���p�JQ���'�?�yR�'��g���iӑ���ڴ��1���
��.b�
�N^!�"�@�xl}�`eoz>��� ��!�'d⍊���1t�;�P 8b��ïJŎ����3m�'��i>�����\��Y2|:��VNu�DC��r4`���T�'�7�����O��d�|brG�Ԉ��
Nyxq��LD~Bʶ>q��i��6M�F�)rc�/�p��%DՂE���)2
Ϳ56l��P8B@��4B�៨2��| j�C�F5�VLC4/��#��',B�'���4Z� �ٴ݂]�墕�.8*��Å�iO2��L�U~�fӬ�PکO�%oj����i��d����i��'2�P�޴9=���vl�f����L�2d��$�~BB��!�Ľ���T�6�~,��Ǝ�<(O����O����O��$�O˧7l��Ȓ$I�4���9�h	�'+,mX�i�~��V��	Z�'&��w��Y��CR�,)�=b��R�>�Ν� H|�4@n�
��S��".AӦq�B(0���!��!�(aj���Po�R@��O�yL>Y(O���OB`��`�v�xC�Ŏ
D�4��O����Op�D�<�Ĳi��I��S����c�(�:�iY�r�l�h�hG:^�I�?�R��ڴ"���3OT�0�ldqn�;y��|zww�L�'������#�����ԁ\؟P��'W�A����2�@c�N����r��'r�'�2�'�>A��+3�T�Ц�Y�T�̌3%��`(����M+�n���d�ڦ��?ͻ���� C��]mXZ��@�0"]ϓl1���m�0n��R�vs��F�b�a�O�|���)B)�h� ��/O�0 �!�Q�ny�O���'���'i:㢒:'�\ <��ŀ��<1B�i���ؤ]�d��C�SƟ(g×�\�.��w	L���P"E�P���������4H����O��X�$���7$Rh�UH+5���굪�L��y�O�MC���?Q �$���<���_
q����;PgF�Z$�'�B�'Z"����Y�x��4wb�)��:���a�/��@I咥c��0������~}Fj�Έn��M3#���]��A���G6%'(�	�G�;���۴���Ԟ$Z����'��Oe�@�{	��ud�Z�8W��j"��	��������П��IB�'�X!�gA���mzF�Ö}�r ���?9�FV��a��$ �I�M[L>Q C�u�jd�3#S L�2� &-32�'x�7����
Ux�ns~� FN��̑�,))W��Is/��O@����ݟ��b�|�_���� �I��x:�莰��(C��X�.�Ґ�G�����ay�eӊ��f�O�D�O~�'n�8�P��K�D5����%�=i}V��'�p�|�ƣqӄx&��'!'����h��b.��%5�`8r��0@����Wk~�O*�(�	�VU�'︈����2�y�
S�&� 8���'�"�'�b���O���*�M2튚M�x���!#z�����w�����?�p�i��O��'���D0{� �X�N�L:��m#`H�7M����A�ɚ����'��Z����?����-�3 ,L�X@ɀ*5��h�<O�˓�?����?���?�����)ߩ��U���^0�s���xhzUn��K�,��ǟ�	|�SǟdZ�����΃�x;�L�� Q��c5���(�)g��9$�b>���^ߦ�̓�h僧	1~�(@�!m��9͓z����ӧ�O��N>�+O�	�OrUy�D�=$�.��u	�+t���O��d�O��Ġ<�T�i�P����'��'��\���Ң�2���퟊A�Dh���k}��r��`n���ēF����7%�92:�1��jm5�'vdjca����� ��$��'�8hASȝ�WB����@���̓�'�b�']��'��>��	���
Km�N��gC���=�ɳ�M���)�?m~�"�o�q�Ӽ�A,�1��	���,@!��#���<A��ia�7�Ȧq�����-�'�FP��&��?2��������ڊW�����m�=h��'��i>�����d������3B����V8W�nux��ۋ/]�ɔ'�87�U�!�X���O��D<���O>��� �&Mf4�����Hђ�M�y}��x�^�m+��S�'
�<8� �!OK�.��!/ɱ
�<�+W�T���	�c��P'�'#~m%��'*��27%w���&��e~�dy��'+��'�R��dW���ܴJ 8J�����@ΑmL�|`C$�N��&�$KB}�f��o�M3e�
�P���^�<�Xz�J6��iߴ��DI�Qp~UI�'��O�_�DH��Ķ8��ݸFJ�wl���?����?a��?Y����O�Fu�q�Ы�p/�
߲� Y������M�����|���6�|���xc�%�"�S8ym!�NADJ�O�$a��i.t�6�(?Ap�W�6-zl��FM�s"�8��G���B�O�1O>�+O�i�O���O�����Lh:-���HB�����O&���<9b�i��s�'���' 哉v|&��̈́�a�c���[)��O�����M3��i��O�S��.Ls��A%-�D��
Ԓ:p炜(���p'?�'7R ����jn�B���^���(��"y�@����?����?)�S�'��D
֦���A�
)��1����GW�xa G-vTf���ݟ�ܴ��'.�J�V�C20��r�(0N���iȧh�86-�զaj&J��m̓�?�a��J�8�ɖU~"G�QwHK�F�{��,ñ
���y2W�����`��ԟ�I���Oo:��FI�J�"�b�Љ2p���e�QE��O����OȒ����L��睾xIDiw˚�2*�[�,U�4P�����M#B�|�����'@�#�4�y��cn��qI?��˃Nۖ�yR�����	�<��'��	韴�	*?�l��f,:v6�rP��	>cn���ş��I���'S 7�����D�O����
%�lM��1b���邞,�����OlHn��M�x���`7:P���\0�#)���y"��5�J�	�� 	�I2?!�'��D���?�ֈS��:M�v)�fm���FG�?���?9��?�����O��Ia�9�fY�C-��xY��ҷ��O6yl�`��Ea�6�'ɧy�LX�U^�,��:s뀗"�|)�'5Z6m^ۦ�2�4A�v݊�4��d�D���'%	����w�U	ReO5K=`yB��0���<ͧ�?���?����?�6!�6&�.q �%Jp�$�%c���\ۦH@x�H�Iџ�&?�ɊP2F���c�a�hQC!�q���a�Oto���M[%�x��T+�}�*8�dV!d�|�� N:V�إ�B�����^�t��g͚�Ox˓X��Lqq��/�H}���I$�Ό����?����?!��|:(O&5oP�D�	^s�A�A�Zܹ`G�]?扽�Mc�2J�>�P�iqr7mH���B��$��Yyf�ƹvX �#/��3`&�m�i~R�)|����p�'��6�K8,+�!�G
�XH�a�C��<���?����?y���?A����F�\b��*�̢@�"N����O�oڒ3(�zd���|��M�Q<(z���7�����	�>H��O��oڿ�M�' ��#ڴ��d��v*
���Я�X(���_lD�ȕ��?ё�%��<ͧ�?)���?��hѮ�. !�
����p�ئ�?�����H馥ʄAw�\��͟�Ou����"�M��t�����,0��O
��'��i% �O�S�K�Ĵb�hTҞ�P�d06���m%i�X\C�M0?ͧ_Ӱ�D� ��+,�y@�η�-yԉh��+��?����?��S�'��d�ǦI{�A�8y�� � �H(�88J��<���~����A}�Mo�@Tx�6k0h�#�E�1�<��"�Ŧ�ش+<R	q�4��dXjjl��'��S�s`�l��Ê�S��->Lɜ'��	ş �	̟8�I˟��N�4̓�K��퉑1*�Ȉ�Q�X6mi]��O��:�9O�-mz��+GC9r�
��	&���Ѷ����M+b�i� O1��sr�s���	��N�8��_�F4I��]�[�z�I�-�)���'�!'�0���t�'���� ��LѤ��d��<2��'r��'	R]���ڴa�m��?��f]����]�&�����ͫ%�%*�"�>���i�B7-�F�I1+Ŏ�x	� ��� C���2������"�_�z!*��$?��'7���	�?	$C�y�I��bφT�V䚐`͎�?���?Y���?����O��!2gFDU*��HE����S��Ov�o�2A�6�M����4�.���޵#d�C�鏭}�&<O,Uo���Mr�i�ܐE�i��D�O��ze��Ҥ-,:v��!��Ztɠq&Bt�P�D�<�-O�	�O����OL�D�O�t(�/� ;Q��@b�p3��<Q@�i&���'X�'L��a5�y��'D�A�G)Ȇnl���2y��V��/Pt�jٴ	���Z���O*�t�ҶtY�`��*���89��Ɣ�r����Ӌ�%���)w�j���L�Z�$�<�-On��@��^@��!��,��X����O�$�O��U�"�H��<9ƾi ��w�vt�'�G�,���hʞY�a�'*6��O���|�GQ�4��4Ư�Ig�Ez�"��eQ<0�H�UQ�|�rh�
WX6�c�4�	�O��t�OĢ�b��l�v��! B<#�]u�܇y4xU��?i���?����?�����?�F矪#��5;%�@<(F`@�%^K~��'�6M1,��O|oE��[W�M.|�����!܈�aI>	�4d/�v�O~���q�i����Oʴ`.ԫt%��K��%��C��K+sS�
�3!R�O��|z���?1�O�а@w�|�L��3BT(��@���?I.O��oڳv�Z��'y��O���K��]�|��c�6h�m���R�yb�'Qz����n�z�$��S�?� t�2,Ә��X ���3�Ը AeG�ªLp���'��	�?��`�'@�E%��[�H��2Ң`X�����	������	ȟ`��֟b>ŕ'�26�ϼ"���
@	�E�d��C��!w݄��������4��'�z�Q���T���o/c\|��0��,>6-Pզ�#�f�u�'��@��M�?���\$����$P�T`�����<��0O$˓�?���?���?i����I�p���K�
��.-&��m�<hmMg^��ş��	T�ş�K����pn$-szp(�Kӄ7.�dΙ=��i�~�O�O�`�
��i���Z>tY@A)a���.���+����W�I��
!��O���?!�Hi})]�f	���M;��,���X�	��x��]y"Mt� ��6O��d�O�0���>E��%� p�(�`,�	����ڦ}��4{�'���G�_جq١H�<<�t}9�O�YC�C�8:it肢�iߟ|Q��'���y(�8#~!�1	@zV��86�'���'�2�'��>��I�ch�1
rN�S�>����ܕZ��e�ɲ�M����?�� ʛ��4�l���_X̚� ?F14��23O��l3�M�ҿi��ɪӽiq�I�~0b���OJxX�w]>"xĀkC
��$��2��E��Uy�O�b�'C��'�	D� z(�
�E1j���]�w��	1�MK��>�?I��?1L~B��t.��&I*wD��r�	9�JU��W���4[���`4���N�@[���U�mª�A���9=6@����V�	$8�z 2 �'�0�&��'��-��MH�l��+
��5^�t�I���i>m�'�6�S�V���d~���j@�l>ru�B̘=�����M�?�W[�d��4ab��b�R)D��5�L%
bI�"��Z)P3��6m4?���V�[K��/��߁��nǟ0lp%I�mB^F��r����֟��ԟ��I۟x��概�}@�L�A۶"��8DЦ�?���?i��i�:%�̟plZ@�	�7�5��G}���KtĊ�GU2��H<	��i7=�n9�%gv�(�T鋀��=2�<�1�*L��g �>���#�䓇�4����O6�ē�u�^c��Y�9p��"
��t��d�O��
䛖g(L���'mrU>�R��,n�L�s�!R�:}�g&?1"W���ߴcțF�;�?�"��/&:I���p{�Yp�FW�!����e�S�N����|�c��O�՛H>��9v�8 �A7���2�[��?����?���?�|R(O$�m��_c 18sgL�TW��J@%T��|��#�CyR�`Ӯ��J(O��$�1h�%S��B��d�'���f6 ��]k�`Pܦ��'�IQeg��?M����0`�7�1kPEڲI�\��3O*˓�?����?!���?����	�U�-�ըŮK|��`S��XHn�n!�	ßH��Z�s�8������k��tNR�fm�k9�I҃���Ҵiɮ�O�O���i��Ę)y>x� t��*��4 C�Մ%�d�h������5�\�O���|���a�vXq�� 3����CdX�)� ���?	���?�(O6(lZY���	ş4�Ɍ�,@�E�?���s�HO�|H���?�F_��K۴j~���1�M� ?���$v��!�R�F���9Hz��ڱ����c>}�1�'����ɫ6I��آ 
<D���Q@��`����	ߟ���؟��Iz�O��M]�#fnH�DOA=2jY(�bCx���`Әp0S��$:�4���y�jl�|�Gw}�X
Ã�y҄gӂ�l���M�Ä��M��O�L���Q����-�.~���E��p��J� �O���|���?!��?��ux��`1��'BM��k҆P-}B�J-O��mZ�Y�h��I럀��c��̚���2�Z}Y��K"���3�K�9���O�1�4���OOl!bv��!X3hT�2�߳ Rm)"�X.
3:I��O�:W$ձ�?1�O&���<A��ǧT�qP��ӣLD����W5�?����?9���?ͧ��d�ߦ��V������$yK��@�ᑆ�O"t�����Mۉ�I�>�Ǻii6mX���٥�\�[�rh9��ςF�	�H�����n]~b�SYktI�|�'��;��by&x
VbJ�J5H #Q�<)��?���?��?!���kQ�cZe���
���J �
)k���'F2/i��,zw=�>����'�C����mtB]H��Z(��������t���w��)�3j��7*?���"�,Kbk�^0R���h�i�2
�O>��O>�*O�	�O(���O��7�ʓ,�|�Hv�ιg"�� �c�O4��<�U�i+H���'���'��j_z%i0G�:*U!"a@�e�P�x�I��M�f�iMO�0TަL�3�M+�l�i1�
�*C%f�DT�h1qj/?ͧ>���d֞��"����C�E� -�%�2E�? �<7�'?�'Mr���O�I �M#U(S+/+���N�	�-#�!\b[�����?	b�i-�O(l�'�6�����i����n=�M���%.w�	oZ�M�'��M��O����@ޕ�"H?	�gMMɒr�W�-��O?u���<A��?��?���?�*��Q�g.p&u�6�%5]2`��զM)��A� �Iş &?%�	��Mϻ	�*��Ӄ��R�1�A��>n4�&�i�~6-g�)���eo�<Qs�� ^ �0c�
��M*h̔�<��3z���$������4���$S�'�$�X�'	x����ݕH�r�d�O����O�˓{��H7�y��'�"j����(�>~�Bezc#H&H��O�0�'?�6���1M<� @��^�ty*�OB�-j��@�����X��<y1!1�ӏX��!��B�D�d~���^_An-�W%N��x��Ɵ������F���'�� Bs��8yt��ᦝ�[x�8���'{l6�Z:�I$�M���w�̭���H�h�ԫ]L*fc�'�7�Cͦ�b�4wp�ڴ��$���J�'�$!{���3�2y�&Eѥ6|	rn2���<�'�?1��?���?�c�'*��q*�o
�P�����(�9��$�ubWmm���Iן�$?牟z*�8rNJ����sȗ�S8ڬ��OZ�lZ<�M�f�x�����@��N8�1��1^HV��P����JI�¨z��r�O��Y,F���`Z?F�r�8���z�,1��?����?���|*O�}o�"���I�7��z̱7`$@CSF�H�I;�M[���>I�i7m�ʦ����3O���+ާ� U!W�1?d��l�R~2�\[�t�����O��ʀ40���V*b���(��Γ�?����?)��?����O�䠈&R�;.LS�KI�Om�	��'e"�'��6�H����O�l�~�I�M�� ɓ/��+�i��\@*u�L<��i<t7=�J4ʤo��.���IS�ǱK+*�����+��eh�P69�l�$���䓻�4�f���O����t�f�A-Z9n��q��O�)�j�D�O6��V"�(E���'��W>��Q. @�����8T��Yp2f)?y�S��z�4*?�F 0�?�I$�
 (f`	�.�C��A����D.�}��©0����|: �O��H>��(�@%S�h��v�޼���S
�?q��?����?�|Z.O�m�*^����UǁWS���'�B(f�LP��>?��i��OZ��'�V7�
K |ܓbm��)Ӗ�1vɥ�>�lZ�MS&��e}���'2���m��?%���� ��L�v ���ؿC
`���4OV��?���?A���?9����d��UFT��!!T/Y;um��7*����� ��p�s�p�������}ˎ�)��4T�~*�-���i>�O�O2��F([��y��DK��٥LW5�t��Ë��y�aL
]�vu�	8?9�'��i>%�I*�����i�z"��t�7T�D��I�x����'�L7�θO���O���99��5�w&[�R���Y<�����$�V}�i�r0m��ēzt��Ќ55\��i�)�/{(�<�'m�,ړ�P,[�R@��$�P�|��'��2F(FND�]�.�`_R����'�b�'��W�"|r�\R��&��>4JhJ/�9��N �/@����IԦe�?ͻw ��0w)�5��)�(�&�X��?y�4w�����"=�h+�O�5��º���"ȫx�"��u�[=
gN���.�OB��|���?���?��*a���ۥZ���)�� 8���+O�}o#CJ��ݟ���m�s�@�r����,��^Z�e�@�L���O|7M�D�)�	��i��P��2֐�ЅkK`<zЙ�f���	�,�zT���'0'�@�'�<U�1d�>����˗��Z��'�'F��'�����TW� cܴ,�������aj�؜"̱���{m��K�zݛ��$t}b'g�n�mZ��MS��A#dB�b�	WkZHU�D�`k&!�~Ҫ��R�Smܧ׿c7�Dh@��ʴNث&RjT*1���<���?���?���?	��4k�0h#N�OґPs��1ck�b�"�'�|�L�R�?��ܴ��K8X�ru!^0���C��>�$���x�fs�\Dnz>!ÖI��crh�I8 ���B�:N��d��N�/�0��W�A3D*$�dL�����4�����Ox�DL�[d`q�ɍ?E�D�#�)���d�O��u��Ɓ�����O{�̺���96*�����>>Q8��O�`�'�:6m[Ѧ�HI<�O������K���V#6��(H&�O�(2K��P���4�d`B��^�h�O�t�Íe���wŃ=@L�kRO�o�7����������d	�
-
Mð@˟h����MS�2F�>���i�p���hCV�R�B\�/�Vx��dj��l�$`Ĵ�J"?Y7`K40�f������R�(�㉃�#h���S$R�$h��<	ߓ�p�Ip-�&z|*����@	��i�B�t�'���'/�@lz�����5|�Ѹ5n�8Q��ɻ�����M���i6hO1��P{si�-\���^ي &c�o����R�D_4�d0e3Ѱ�+�֒O ���K	01��q�� jx�y�P��;�ax�i���ђ'�O|��Oh5�a�O�D��Q�q�L�cMt����7�ɻ�����ݲ޴2��'�i�s��g¢9��_��e`�O�E3R��0��1�?�iʱ�?���Ofy9�/J�\o>��Ӧ	(��C$"O��CL��4���>#��LzR��O8�l��f�^1�	ԟ���4���y�
T���Xz��߫G4LzG���yr�n�R�o���M��OT�R�)�'0J<rwFZ�?	:���d�:����?$D�bgl��5�'"�	͟@�����	����ɨ(����)�+Tڈ�:��7w��'�47�6���Ol�D5�9O�`��ޜNēkR�p�8`�3�Au}"h~�&�lڅ��S�'hH@I�ل�D��d])m#�����_�y�'�F$�%�ߟ4�|BW�0r�i�w���g+Q(S�zu�0.埈��ğ��	ݟ�Ryҏr� ��3O��@qc�U�Dݓ�� �g�4��8O%nZh�m��ɡ�M�i�T6� ���`)֊r3|lcUD@�h��J�g��:�x�(痟*Ջ���i����Bd���_kt��(U��H56O��$�O����O����OF�?�s�H]�p��2���-R�b��3�k������4Il�q�'�7m>�$Z�~�X�CTC$=���@a�<3��%��	����7LhEң��X���� M�x�D�q�V���9m�6,P�'��4$�4���4�'���'��R��=�	�ֽz4� S�'�R�Aݴbb|�ϓ�?�����)��C`��d`�t؄𣜰F������T𦥫޴]㉧��Ws<t��lڗB���GB �p����U�f�y���!����y�-\��b�T�Q����"Dur8����`�	���)�Siy�nc��#!޶-���v�@28���ܺ+�	�Mˈ� �>!��i\dQC�k�5?t�(��������M���i~��٣�����D��AF�(�����"!� "ԠW8B���C�Ҥ~�0�cyB�'���'���'��[>-�À1rb�憎d�5�Q�ӓ�MsE'��<���?yH~�:��w���dGر W)+�O��$�@!��p�lo���S�'nV��
��<YQ���lz�a2H�^��I�b�<�W�V���������4�f��ٔpD���Xw����o%?�����O����OJ�@�6fE��yB�'��,�vk`]��o��o|���a� �[��O�)�'�d7�OȦݩJ<i��I���n�0�bhs��x~�Oݵa�Ua�%�טO*�u�ɵW�B�?;�L�N�?]^�� �]�X22�'��'v��Sٟ$I�H��BL�D� �J�3.�;�Sџ��ݴx�Ty���?�@�i��O�.R	�rY	�+Ĩ+B1�"�5�$�Ԧ;�4�?asAA$d�'��(P��W�?iPT�ȼR/᩵Lژ-P�9eK$��'�i>������	ޟ��I�#���C@Cy�4�&B-6��'-h7��)�ʓ�?	K~���[6��R$�^n�Ph�v�l�`��S��ߴ:C��=Op"}2%�¼D�:T2q�-u˴�@�B>j@p��t�v~���6|���Il'�'�剂A.U�ȚO�b�("%�[��I�I韈�	۟��i>1�'(�6m�A���֍&�Yؔ,�#J..xY��_	d8n�d�Ʀ��?qdQ���ڴ&��'X��P�� ������NC�0��yʕɗ�/.���O\œ�K͖����k��ǏN�k~����-�MX�p��du�P�Iߟl�����П���(]�iq�9tO�.X�1��!�%����O�l�u,���X��4��$�T����8�uJ��G�r�':�I��M�����N0>r0��O�H2���%q�J�J����LU&߿R��(�� ��O���|���?Q�wN(�6�-^b��%��J�%9��?�,O��m�)^�0�'n�R>�x�HF&P�L��KV�(�r��)?1`W�tX�4Lj��9O�b?�i�@��FذI^'$�h2Aɚf�6j�/��~��|����O6��L>Q�\G�؋)N���T��DP:�?!���?����?�|�+O�m6M�.%��J�'$p�$�p�<v��Bs���x�	��MӏR��>�жi)��wo�#yK
e �X��l���j���dϻ9^��@���[!d^A��ԓ~*��N�15fᲷ��2=� ��uf��<+O��D�O^���O����O>�'P;�M���&��'Ů	�����M��hI&��D�OF��t�d
���5Z�� f�=A|�KB���ѸݴgÛ�7O��S�'߸%*���<�@�Y2�bb��U4ҵ����<a`��?*�$X�����4�����3J���C`�� b�c��P(_�����OR�$�O^�p^���� k�	��H1�Fњ_q	p�B��$��Y�T��T��!���*�Mְi��$�>���R�x��L�2��0/T�2!�Jp~�e�aN���cXƘOz��IF�/��e)�1��n�_.x;3d��?���'���'��S����j=�D��EJ�3+bBUNݟ�@ڴb�n,�')*6$�i�)�c��<>����b�C�8E��,n����4���p�8�e&�K����C�:��C�O��UzU.�1����J�f���e�	]y�O-"�'(�'�Dˁm��+��/zl��X���1u�:�M#p%��<���?yM~Γn�4�j�)<}�")1C�D��At[�h8ܴb2�&�;���9��0��n�2R5�-�`L�o�<_$�4�e��ܘ�y��˔V�Wy���@th�G�I ������ѹ?���'A��'��O/�	&�M˗���<A��5N^���C��Q��0����<6�ix�O*y�'�X7-����ٴA����J�f���(T�L��p�0!PM�'�h��' H�?��}J��}��i���+���Ъ˝`̎͓�?����?����?q����O�B�uGH��a䀍2
� �O����צ����(?qd�iJ�'T(���B�Y�8 C��'@vp4`%�$J֦����|:�m�#C$�'Tx����sk���M՚W!�H��ȏ7u�Y�	2z��'t�i>��	��I�<�$��� ݩ@�&��pHI\3��������'7m�"e��˓�?*�DY�3 '+�d�R'ׅraP��4���ٯO�m���M3�'�����ƈP$��Qb��(^�0�H@��\)�!l�i>ur��'
�H&�4X7�ӵ&�ƨHS�	�O��Zc��Ɵ�Iϟ��	��b>ɗ'I�7�&9¶T�s�Y+�l��#Ϭr���y2,�O������?��Z��i�t�? ��6)��@%R��E10'�S�JΦ��ɲ?��(F-?y��	�M�n�	)�d@��!�И����"��
�y_�0�	��H����|����x�O�������?k�@��5X̤�U��M{T$�����O�������̦�]�Y���Ig��AeBEb$�;z|���4r�F3O�S�'?@FPV���<Q'f��\=�2��M�$}�o��<��O�5��D׷����4�z����LP��;��4��a�1��\����OP���Oh�pɛ��ڹs�R�'G"��2W��i��:�����"'�>�G�is�7�Lr�	"!�>8��IV�H�1s͂5	���c�T%�F�
zj� N~���Ot�H�H�e;��	�LZ*Q��Mp9�����?Q��?���h�&���*���@ş6r��I��G��$�D�yj������ɒ�Ms��w��Y�7 �'�����;�^:�'��6���u��4
t��Ϛl~��;�V �S�X��h�X�x|�3CO�5�h,�&�|rS�������	ٟ�	ğzd��

��9�p,� !Ӥ@9�Lry��d�4��2e�O����O����$�9U|�Hd���i\ؙ���UJh��'�@7�ɦ�J<�|"զ�%�, [�H���Ъ�oU!%�ȑs�.C���d�Q���k����O��-$h��Hֻ7���tE&�<���?!���?���|"/O�mZT�e�	.?ft���-D8�!ËR0#/��	��M���<1��Mӕ�i��Hy�)��&gx�te�@�����嗺O� I �O�]g)����d%�i���!R�Ȥ�А����k�f���7O����O����OB�d�OH�?ii���<��HI�vi�p!��Vy2�'��7��%3l��O��lZg�5� �R��5&a΀BjD"Z���͓�� Ѧ����|B�M�xM¨�'rր�oD9s�M���Z(���K�$�N��ɞ��'��i>A�I��T��,;�I�N�9�:l� ����I�l�'<6M�*�˓�?q*������^6�:�AA\�������8�O��l��M�'���
���#�2k�		s樻B�A	w����ˇ�%��i>U��'c�)'��M_�fy����gٴH���$�I�����ҟb>Ֆ'��6�K�]�pPK�̝#���Y���.l!x\ޱ�$�OF�m�N�{n��r����Ɔ��w�`4)����M���Vy:e�A_~��a��u�H�)���(r�D�%���Ҡ�ݾ���<����?a��?I���?-��aJ
;>����jG���ȕʦɐ�DAGy��'��O�Ra����R���R�`ͩ�6Y��C!5x@dnڋ�Mk�'�)�Ӎ{��*��f��u֣T�-����pl��m�JE�>+���V�I~y�O�l�]�HU�E�G0��рO�>���'��'��	.�M�!�#���O�@CR�*U~�{G���̀�K.�	���J��p�4�y�S�\�p,դ(X�ݫ�%��0%|hb��=?�WA��y�� ^ḩw|�Yv'T6pfdu3&"Q�;��q`P��N� ��>uJU��
�&�ࠇ�6mV\�!V�/ք� ���8 |����(Af���� T�q������O����e��&>"�b��ܲ,q�Q��(UԺq�|�W#UU��)�M�v�IQ!b�eK- +$������xł+V�Ou��s���?xQ��
T+v�J�[�@;s��Y@��6��@�L �vi�Ðké?^�}�eR�l��V%>�^LZ"��&J�a�eN�bA���NH�	 �C�c�d��EԠ{�B]kD
L�i�HE�i��L;kuNO����O̒Ok��m�*(�'	O�K�����׷���'t˞'Y�	㟀���`��ʟlA��hPYZ�ǜ�F�x��+�9l��'���'mҖ|��'lb��?���ٍ6T� $hȮOK�Ja�(!2n��?A���?����?�QÀ��?%d�*8,�s�a�;,o Mӂ	ϭsћ�'K��'J�'J��'D8�����M��d��s3LP�4V�3`ȸi'Gt}�'���'8"�'�|U"[>���5E���h�M�pt�Ү��yߴ�?�L>q��?���$�%���f�M_H\��ǎ��Q')x��D�O����O��م��O��$�O.����L��u$�!�&Tp���v>�+��i�I��$�ɘ֢��!�~JDf�.VƘ@#�߾N�*��t�E�	��؟��m�����qy��O��i�q�B�[ ��hh��6��qӊ�D�ON��V�|�1O���L���'��$a�]o���ij�l���'���'@��O-2�'��Ӻl~f�[��
 ���=B#���ܴ�:%ȴ.�{�S�OCBmU00f�`�RO*�iO\%e�"7��O@�d�Or�P�l�d��?Q�'����ƃ�!5P���B@�%ڔ̀�}�ǁ�Ԙ'F��'"�"c&8(�Ɣ8Ga�H�U	X7M�OZݹ�(X}RQ����b�i�Q!�GƲػ���/�
|��>�%��/���?���?�,Ox,굊�4?JV S��ݿ~p�c��(t��D�'��˟�%����˟@����^{@I{��X$Ew�a��� Fh��%���	џT��ty��A��)��B\�	0�]�O8k���}n��'��'M�'��'���[��Oj�2��N�&�ꗮ��7!��z�V���	�����Sy�̀1P��'�?	2N��H�7��.��E	�J�9`N���'��'���'��ycF�'!�Bp���X	Ir )f�x��@�Ц)�	���'�$A���~*���?��'h��R���p�J5Y��$;��i���x��'w�d�KU�O��������d��n�#�kU�
�|6�<� �W97����'���'��dj�>�q�? \I�h�$H��	��L�W����$�i��'��Л���7����hց�%[l��4@�no�7m[�G��}lZݟ��۟l����D�<ф�F�lbY��7��i�����RÛƯ��s��O��?U���?"L\����"Lh�A�ִ��4�?y��?ivm��R���Ry��'����j�`)�fbK14�Nus��^�#��O4$K$)(��O|���O����Ɵ5������a̺�*�A�ߦ��Ʉ:%B�J�O���?�L>�1O̘�!<ܬp)s��*U���'U�Az�yB�'gR�'-�	qBBԛu���ZE��/�|:�KvD����<���䓟?���Z���R���o(�}���&�ڜзK�4���?��?�.O���aB�|���^��x�_�k��8r��͗'B�|b�'~r쒘��	Jm�TAR���F�� j4�US��	ޟD������'(!�S��~��Jm���$҂}ڜ=! �ߡ'�xqe�i:��|��';�؇'�>F�Y�u�©X���������צ�I����'U�*aB>��O����F<��B�8��Y�[ N��̙��x�]���I�p%?�i���M��}0t	K����i!����EӲ˓hPHㄼiC��'�?I�':��I�?BUj7cұ�`šԭZ���7ͧ<����?�����ܴ;ܨ��4(S*En�Ԁ:Nn�o���Pݴ�?���?��'n����dM�;�Rh���u�h�q �"_��7-�O���O�O�s�L���� !��� 5ڴ�Y�e�=���"�4�?����?qC�޷)牧���'P����H@��
Tpr����(���'I�I#@�<�(���I�p��c�~��sl�U�HA�n��9��ao�꟬���
Ty2�~R��K��2���c��L��!;��O͜�9s� ���v��?�)O�����D��щ�:f=z�0ŀש?�N̂ao�<9��?1�R�'g�cԤB��܃�D8eJ�B�&�?"0n�b�����'hBR�h�	/'؊���x�`0�*�Iʲ�Q`��[�<Un�ʟ$�	f��?����8)�����! 1��H}vAZ�eK7 d�H���>����?	����{Jna%>�q�Lѩo�����N�)�hU1!�1�M;������$Q�{C
��/��f��@���)D�{��h��Mc��?A(O0IR�`YN�ɟ �s�as��Z�~���3!�"*p��k{Ӻ��?Y�"������'��1��ys��]��5���ׂ{W��d�<���Z�&U>����?�[�O�L3С�&	���N�5�n4���i剁&aT��&�ħ���ݺ���n�H��K�)x֍x�!c�~�I���O�D�O����S����m��\3E��?Q�@���͸M�,6-Y2��l������"SC܂x���J�2=>\�Ƌ]��M����?Q�����b�x�OO"�O�Ղ5bO�<6�93��> yq�i��W���w%����9O��D�O��$��XA�fn 
��S�%"�oZ�l�'����|�����Ӻ[q圼	 �*��
�m���sr��n}��J(s{�U���	��IWy�ÄB�tM�B��^�@�a�7c
�(�"7�$�OD��O*��?�М!��Ν�d�����-=�v���/�+�?�)O���O˓�?A��C���d�(j���H�f�1`Z\]	�lԻ�M����?9���'���D0�@ܴrjn ����$�0�r#�4b��i'�x�Iryb�'��y�Y>���$�,��ci�H"X,N�.�>�a޴��'fb�'*�aA�����[~�`�eF�/~�P5��@[p�Xo�ݟt�Ijy�K �?�����$�kl��s��z7@�R
��ucT��'���!R�n-�	q�SGj`d,n�X@�@8ѣ�ZR}��'4��x��'��'PB�Oj�i�=�!�/~b��㯊7�Y��@fӆ���O��i هT�1O���A#j�}	j^�9�R�pָi�j�aTBu���D�O���⟚�&���00�S�L�!>����P��гܴZ��|K��?�*O����I?U^~� 5�� `��pqm�Q!l��4�?���?y������?9�O< @���0.p�C�D
���(�#\~̓0�����O��	:_:<��n	�\�.H�Wm�h7m�O�9���<YE[?��?����1O`q�E��^�! �/X�L��	�lr���>?��?I����dצ0i�ŒBF��T��l	�O\?K�9���l���� ��C�xy�n
�/*֌�Ɓ��M]j�Xen�aL� �b�'7�	����ҟؔ'>�DF�k>�H�X�B0��2��+yY@��>����?�H>�)O4� 0E�O�S���&*Yh�Y���=T�e�@[M}R�'B�'��	;Q-���O|r�	ڪv:5�.�%�~��Q��*11���'��'c�I�2�4���D�I	�5��A!A��@|kq&>oЛ��'~�Q� ���=�ħ�?���a��!X�@Q�o�a]&DtDp�hyB�?�Ҙ��ٟ��y%e�+/�2䙵K�T����i�剚7��l�ܴ0���ן��Ӭ��䀚~)��ׯΌ1�H��jW���Ɵ��QfO�Ot|&>�%?7�$i1"y2��7�����	�	���CʲO�7M�O��D�O�i�b}bU����o�\���+���;�����_��M�$J�<�+O.��"����e���R��m�Oǵ6�|�#F�0�M����?���wp��R�l�'���O� ���B��B)H��@G�~��S�iXBX��K��}���?����?�BA�>@����^'|�T�B�
F9��'M6����>�)OX�d�<���kR��)��Z2oڷO�
�!%UO}R�����OJ�d�O0���<9�%D�{�|᥌]z���'-ɰ5x�]�Ԕ'i�Q������8k^����j\bQ�"�	�AC�|��e���I՟(������Ly�L�.)wn�S2��8e�O�X�1c'�)��7�<1����$�O���O��72O�)�B,���Bc��
!j��4!����ПP������'��ɸD�~B��`(٘v��(:��+B�D��9`Ӻi�2T�$�I۟��I�u\�c���*W4�@v��f��{�I�����'��\�FD������O���|!����;Y�\��e���L��I�@}��'�r�'�Ұ��'��'��^�>�^�`r��L��2c��h�i|�I�a�2��4�?����?	��!c�i�1��\�v<EPl�LyƕP�~Ӕ���Oޝr�?OZ���y"�	�g	�R 
3$�J�:�/ˤ]�vBM+Q�6��O��D�O.��G@}rT��K�c�7z���wH�#nP9����M��Z�<�K>����'���x!.�RPv����Hc�@2'd�N�d�O:�dW�4���'P���h�2Y�$�k�1�YY§�5E�H}l�ݟ�'1Ș˜��	�O�D�?�h����z�<�1b�3CN�4	Fe����6���'j�	ß �'kZc���O˻%����T�'��,b�O���$=O��$�O&�D�O��$�<��l�m �u���.��tSp)ˤn�$�1R�X�'�S�\������=��Qp�F<|,�̑G��+@��P!��q���IܟP�	ڟL��yb!�
2���{���1>Ȱ%0碔5�t�ٴ���Ob��?����?I���<�w@?
zZ��(8ထ���׬w!���'��'<�^��Kq,&����O�(�Ө	7ZJBT�V �5)жj[<�6��Od��?Q���?q�.Z�<�J�Dʃ��[�T)�,ؖQ���s�~�"��O�˓b���Q]?)�	�t�6k0��k�j�91������*B�zD�O���OT���/f�D�OD������kCt�8AFè'��cjQ��M�+O�<���m̟���ϟ��ӣ����4M�.��80��͓1�j��q�iT"�'T��'<���<���$���v@p���a�x�9-O��M�HC.%���'kB�'3�$��>+O��k�&A�:��hʅ�N��A-oܛvn� �yR�|����O�DRdNW����c)zK��-��޴�?����?ѥ��&��Idy��'^�ğb�����/��k��Ŏ#ǱO����$�O���O�i�ׯ�w���w�8C�l��%�զ��I3H�� �O���?)O���Ƥ���8 >� #�MA�P��Z����>?���?i��?-O�����ū�B�ãǖ�W��B҆,EY���'��Iן�'���'\2�ϊY�Ń��5��T3%�#�4��'4�	֟d����Ԕ'��Y8� s>�' SD%� ��/'� ����p�ʓ�?�-O���O`���s��A&1���s�ӓ<�)���P�R�m�㟘�Iߟ(�	Jy�ňz���'�?y4"��8E�7h]]�E
�bL����'��	��d��۟���f���f?�҆2Ml$ b�t�:�Ĩ��M��Ɵȕ'��5`C`�~���?��'~�t��7�L�G�t|�r�D�z0kQ\�8��֟ ���|3,��ĥ?��a�b*�8AT�����p��mxӎ�FV�hX��i���'+��OӶ�Ӻc�dF*P��E�!���`�������Hp*d�D'���}�w×5�H�����)��7����c� �M����?I����7W�L�' ��i��)%��%o����7�p�t��>O�O��?)��*2(�R��Ũ3�K6%��M2���4�?Y��?х��Gz��hy��'��I�(�Z�S���&��Q*� ��IQ��'���*u]�)����?��OK����ń�|����h��p��ڴ�?1��J(���syr�'C��֘���� U�U�O�.�E��Γ�?���?����?.O~����?5�44�C�]*5���i��W@���'��ڟ��'���'kҠ��07VUcb��+�P�Ӓ��
T'#�	ǟD�Iɟ��O)���0����2�q(�*�Xi�q�xB�'�'7R�'ih���'#t������3� n��ّ��>q��?i����dAt6$>u���3O�1�����l��D��M����䓾?���C*D+���I,[ԕsO�Ie0�
aI.M&�7-�O����<AhA�Y�Og2�OK�E9���{||8��J�
0~�@m%�D�Ob�D�',Mr��/���?ͣRO�9_����썁hKP���mb��˓f @[��i�&��?i��9(�Ɇ;:���H�*$@���Or�6m�O��	�6��5��$�	;���1gR�MCP�KA�U6��1�xAnZ��	՟�����'������@��<Ǩ[�ʐ�r������O�O<�?�	  �ʕ!��:򎝂�	��8p�4�?i��?�ӥQ{��O*�伟(�%ˉN�P��W��4Ug�@�6�c�`�O�ݚM�G��ğ��Iʟ�rBC������ɞTn`p�����M���3���s��x��'�|Zc�2E���8��u�B�>	h��O�8���ORʓ�?���?A)Obd��$4C�k���{;�p� �D�IbL�>9��䓮?1��b�� ��C�Ɋ&4�¸+#�Y	T��4k�<q+O(���O���<�c��:��i�m�މX��)_�pz�h����|��O���x�I(i�@�	�e�8{A$Z�Xh��7�Щ����O��D�O��<�w�I�#��O�^ ��!oM�LU-.,�rb,f����+���O����-$����#}�@�PȌ�C@M<f,�T�0g���M;���?�/O�t�2�h�埔��P�NL�RL"`�&�"'�X?�8H<���?A���<iL>	�O�mPu���j��0�%B�L2���4�?Y�������?�(O��)�<���.�Jw��_ш[��R:8�o�ş4�	=r���h��8�)�CДs�T��hE� �T	"�72J�z�n���(��ȟ��S��$�|��89�n��T�#���d���sԛ��43U�O��i*���O�Ȃť:��m��`��
�hqC��������I9N`l@�'��� �v�d�#�JÜP�8�����c�2)����K����&>M�I<�ɬ|�0E��ɒe��{�� 7�P�4�?�����?�o�����'�@����j��t��N�J�P�EJֳ��DԊ61O@���OJ���<YCD)�������N�q�Jр6ײ���x��'�'��	�4�I�G�br�	:������"#H�I��b<�I��(�Iry��'z��Q��d@��	��NB���m٬FY��B�i��ş�&�p�'���+u�I��Ms��
4]u4q:3�Z8+�A�l�~}�'�BY�X��Id�~�MY=y�:�	�	#B�1��ǃ�M������׻o���5�x�jE�$c�,O�$&X����į�M�������O(��R�?������j���2%���HF1[�G̥�I<i.O�sӇK�K1O�STݪj��#x�V��cɴ6��O��D	�<;J���O������?��:�n%�P�Y����QAW�f��Um��4�ɾ4,�"<!��/�'�mb��?]���P���	�M�An7�?Y��?y����,OP�'Q����.m�ժ�8q��ictl���?�Sݟ؂Ǎ)
F<T�õ#�j�gù�M����?��h�h�.O�ܟ�3z�8�u�^���I�&g̙`~dm�T�$\To��%?�9�@SnpH��i[.��w�
���<Q�l�#Rpe:
�'�Zx�ա�$+ �}@c�[����:דU�T��n (m��1ɗ��TXni���TXf�!ѩMO(0 �c��p<$������Q�  tV�h��Č�`0�`R���t8Db�P�:��d�V�]'C-����`F)�re�iJx��d�
�f^�"a�U�[` �I�0sLD˕�J8(,��l�q������&n��Y�	����c����,���|z��U�h����l�:Y��a�a@Ly��=����ㄈH��?������	�Y�i$���>I!�͉>����@F��<B��)��i�&#�>dԉ�N �9Rޕ���D�'���؅���!J�ѩ=����yr�'� ��b	��O��XK�52�z���'�6Mȥ����tEQ-a3j���$�0��D�<)�I��"���֟�O�Y�&�'�q�n/2c�|��x�Z�'�2g<%�d�FK�A������O�@��d&1J0�!�(Є[�8�ر��I4>kd� 柨s�X�����_�O׈aP$��;W� "g�����T�J��YD��Oz��<�'�?��`H�+� �-�cwɂ�}���ȓh��R�.�%4B�( �ױ%w ���I��HO��H'$�<i,���+*J��	{dDIk}�'>�B_�`Q��'��'9�w�"ȣdL��0�4�a�B�m0�1�莴l�x�C��O�hx�e���1��'�Bm"���0��H�)vΊH6�خd(}��E�O��tJE�����LR�!�&�E0Y �'��|g�S�����-��O�ў�R�/YD9����-L����8D��L��?�\��)��{P��g�;?y��)�-O� ��.е��(Jq*3L9�P�JQe��(����O��O4���պc���?A�O%Jik����Db�"z�L���Dې�x2'ʜ�]i���g���*�f�!A9�]Ru"�3j:����15��#�!�=bFa{���;���M�m�:�c��U^2�����?y��$=��%NNz=*@+�	L���X(_��@B�I�a�JMK�lM0���Ѧ�]$0�c�h*�O@�	>z�TZ��	6xݢqZF� LY�E���a��M�	㟠)@�������|ڴaT 5�ܹ��G^V��u��4r������u��c�&�)�H���0l�#Un���+#M�)�� ��#��=�4��4\�DQ��+O��
��'�bR����I<H�@�23��M�+,��b�4�Z@��n�.b����)�_xB�I�M�`�W(+6�$C&G��)L$)����<y����_�*�y3#�7Gg���*�I�&B��8���A��-�rHS��f�C�I-��x
C��%K�f:��L���C�
`7~�;��GL:��A�)�!�� *�CQ��?_�H��c��l�$"O�(iVi\hX��K�$�2��"O&�)vk�"��l���&"���(s"O�����[��a��d�Ҥ�ʕ"O>tKFh_X�𴣵�J&4-ۃ"O\]�P#Y�4�N�H@�� �rh�"O� i�dϭ.�,�(�X0��(��"O�pX�N�(��Ȳ�Ş�P� A�"O�`���Lޘ`��]'e�4�H"O�@�Bb�j��XtI��8�|5Y�"O:]C��m�����e�(|R"O�P��50�s^�� $@1"O���f�R�5�>��C悲X	r�j"OF�c�k�Z��P���+h�i2"O"�ⵆ1h�
r3��L��KE"O`t�ԌJ93�ԓ�팚#LE�"OT�!�i�-0��)�W
�+_��"O8�0�l �J1����S�"O0[#�X%4�^�!����1E�hs"Ot-�K�:Y�4�kc�U�fX�"O��w��14���ztF+_(��G"OT�`���U������U�9@�%��"O.e�0�2Ρ��C��\��Ĉ�"O��p�#F1��Al�I�HX�e"O�0�ۈ�Z\9R���*B��ʄ"O�`P4#S�hV­��OC�M��].�y�
�8x`��/Mv˶jքX7�yr�J�a~B���Xm5�<��l�-�y҆\�(�B8%HY��Xǁ\�yrH\�E`|y��2�����J�y"��Y=X�g+���Q!f����yb�Jj:t���U���]��y�	�lm�-c&�ڧI��T �-��y�˓2Yf���E���q��y�)Y�td�@�Q��=-��{��V<�y���9D��Q�%���\���	Q��y��ޤz�u` 䊀r�DKp���y2���~��T�%j˞��T#��y��I�l��Պ�Z��1o=�yB(^v�z<�sG
�t.}�U`9�y"�۸F��IE���(�r�el��y��A�~��s�J�/(��tB5���y戅�<�sB�,�<�T���y"���>����f�r�����p<����&�qO���t���"���+�%}g4H�B"O�-)$˝;�&ip2kW+~ZP ��^����ٌ-�b��|�䫝vgF�j����t��<�@�Ju�<1�kY�-ತ�l F$E�q�dY/FY@�J"� N8��#fȿR�����ń�HR�7�O���q��`�9�LbH�3PH�KT�є��'(ڄ�0?A$�¢? ����nOX޹	���x�'cȠ�� ;�:����7����O�Q[��1q3rڦ�L�
�f�'n-4���d�.Z؁�0J�	y��h@W
�O9⦍8O#t���&�&4%���g}����o}5C�i��o�*���I4� ���@��X Q�+>?�y
Sʛ�SZ1 �%Reʰ�'JN8j�P?7��/%�J��
t��F��r㯁�(�b4���=�O2�j-͛nX��oъs�fx�Ul�]�>��Jڼj{�:�g��?ّ�C{.�����R^���ME�HMiԮ��OQ�L[��	��^���E6XHLkЦ��S"ku!��%�f)�Ӎ#)50$�
�'B��ЗM;d�� �\0e��X !��)=Y��A��Q�Nr�Q�e�%P����#&́�&3��Dg���
'ʓk�`4c��S ź�;2�Z�J��D��
'l���V��Y�	X"@��c�����&^$
*�%b�(�V"'*�m+�&���|�Z�� o-�c�b>�K!�T_;��ç@K���3S���77�����CŴ�85FPs�zw+�H��:P��� @��7��p��h�J�v1��p��O֠+w%Fq}��	P��̱�M�k�����M,���#��yHV�V�M��y %�>��8��捅`�x嚌��*E5���}�0���O�H,�Fj�1?��m�0f�r 0�a �\H�2��זw���OX�p&�ƴ�ywɕ��.i2���d��fR�b�b�<i�/�'S2Q?a� �=jLl���n7��&Y�@ܡJ>���	P�3[��kC�˭F�r��w����艀G�m�V$ X��N��(�>�~r�I�%����C�Dԫ�J�2W�b%t�U'�N�{�@U�~-�-q� F �Z�s�╾Dթ��D�7=��HA��:z�du�#�";��DNV���'�]s�+	�p\,��SDF�{bz ��'�����X 75��Z�i��?�X��#`/М%0�C��O�Ⱥӎ�}?a�MO�Tu$�z���0�Q���Z?�'�g�j�	ρ:i��c�E_��?y���P8����|�M��m��V�BL�3�MP�'��$ATM+���)��ؐ<��8��܆r�����!�;�����Nm)U�	��	�'^^F�݉m%�@C�w�*�K��O%un���I��4������@&�t�>E�T�F�))�d�T� ���s�j� 'Q��Pd�X$
T*�p�� �I�e�D`�'
L��&嗧 �>��uH��z�����'�,%�t�7���dT���q@��:��ӣȄ�)~ ّq�\!T\ա��y�*�+��=YإQ�e�'ԨOX�G�?��R(����Y+z���!ky�ɓ4b0�K�<28�@��VW�6�^>f>`��>��`�ת)�2�1��	-n�<���	�aiV#*��a�)��I�1|8��4@��0�I��}T�ÏÚ
��X�C�g~B��k����(UX]i�"ٿ[D��H�~K���7�BV��]�E!
O�"e�[�n�Xs)�l�頔��p<�DXm�,�0v�vl���Y���Pa	)�q A✈eBB�#E��v���煐�J�$�X�	��	#C����$��C��=���A8#��5 v�ɖ�1Od4C��Фp ��8G��H��1Ο�X�(�.���D	�]L�Z� "@�`C�ɸN�| ��
�	F-�`�d�\�7���r�"m �c�J�FΕz�!��l �W
)�'>���gHK�X>���Ta 	̄��"Od��ň۰q�}Aq�\�90M��E�:L8M�%pN�+��$����O�.b�(qe���[�$�s��BZ�h�{��5LOR��c-�tx�x�F�;Vܐ��D�<aj�v��DΈ��h�-���]������T� i�����V�(��)�8~�qO���m�ezJUH�U���O�Z�K�=;��rޠ�Dt�U�*�!�1x��a/ܚ�Ĩ�v�]�V��I�q�r�1�>���O[�h�¢��$�L�k̘֭G�P�0�'��j\!B��aQsN��*�MH�yrF��n��l

�ؾ ��-�6Eg8]a2˞�z����RP�EQ�v|�Y�&�x刀Sv[�����O��cf�T���s"�h�V��㉻i�B$
��ĉ�r�����E��|t��bFO8�!��5����U�՘K�=@ '�\��'�,d; @/�)�ӠF� �n�>$~8h�5+έu�fC�C2�` @Q�M������Lj^C�I/C2�5J5��|�ـ��;�FC��%
�����CH�C��Ⱥ7�	�h3(C��4K����CE���թB6k�B�	2O������Z�<�h��3u��B�	$;�����8��1
���&i��C�	<n�.�YRlܳ-����u�ڳ^��C�ɬI/�Q�	7���{2`*+APB�Il���D���(�,�x��
G B�	0c�%ʲػ>�h�0��-:C�IzpM�%*k]T���GP3>� C�ɛX�t��s�Ѻb�.�ハ�VC�	4`���L r�ԙ������<C�	�z�T�]�i)�E��c��B�	?|�F�:b��+�Ϟ�c�C䉝nCr�㬐�xx�t�W�6͚B�I�c5"X��B�v%
��ՂR�|�$�F8tz��' ��	j�����#v<	�hIh�q�aƁ�y�O�
0�ꔡd,�#i�R�١�ԓ�y��|�L��둈.D���虨��'9S���?-�?)Sbэ[;t3"�3���P�4D�L`Ȓ����Iv���K�'ǟ�y2rbx��]��~Ҡ�)c��&LI�:��`�����~��5eB���� �HC�	�LbT��DhG�2u���'�����F�)L�Q��k��_�~�ĮH���e(�*  Lߪ=�Hi��DꁯZ��	2y�撟����'D 48q���	�t�$��r6�ʊ�dB�(L0D�OQ�2+�R��:�6ͰC	�'Y��j3��)!&8��k�?�0YҝϘ��i����)"s��>|����ځk��H�� �ا�:t��7�ۃo��� �?W��N+%w\��f��=!�Q��t�1g;qa���'Ϣ���B�=�ȩ�$�;q�8��xX����O����U������J�9����9[��B��O��+D�f��$�r�S s9ᚰm^�fHD@(�M0)?���>�(�Tr�I
�T����D�f�δEy�M,�D�~
SN�^��0#�l�R`Zaht��4�Dm��I1&�vM`��D����F�R�bXh1I��
��P���	l�8���T>y(�I����p����?UR&��;P���ar����0z�C䉆s\�����ݒ6%��C��L���	.熔i���Hl��6N�;*�D�9O1�j@w�تf��i �P,G"<���'�T<�p[�<��-YB>9�0��;5@�%��kΜ?т���8��h���E��O*0�O%u�Xpc����5�yI�剕Pa:Cs�S�g������ɂ��L��U:v��T�)��A��(�����ئ*Ɏ|���t����M����ا�	��d0�`@@A����e���
7��y��
<�\�ȕ"Of��D�S����[Ѧ�@�� p��'L(�Ȁ+ɾm:9Ad�
 3�v����yJ?��Վg���P��?3��)ά>%N�8ӓx�|ÔgW]?���,�^�(��<~�*�΍�2P<��6U��ϓV�̨�g�'�D�wi-f@�*gA�?�4@Ӎr�l�(�����ޙZ����S�<Ҡ%BV$�u����(]�:Mp#>٧B�@��� K��ȅj@��&�*��8S�L�J0�ˉX�b���O�m�Ն&u�����
D8`��aH1����4> �=�l���$� h0ܹY�f˜ �]Kf�ߔ!��Ü�g��IR߷`n�mY�*�"�����禥"��!QO�� W�ʊ/�NUA��S�%jL���ˈ+�^u$�OҼ�&#Q�3�X����+�(l��"O�T�� ܗ(�ĕ���Fz�!��	;l�x�a ���0g�-a`���@����ȓCHh���J�pLБE�	�����9
�閯�:jL 	 ��:�4��z�6��� ��{Ծ�x����E`��Ql�Tp��ǫ�(�x��C�1��|�ȓ��I�� �FS�8�<!����"E�	+��O��B�ܝ�yr�T59}n@��쌥z�D4crAB��y�	��0�`c��fD��*���y���1���l��cS�Q���	�y�痤2S��q6i~8����I��y"K86�)��J܅�d���@�y�DIS^������q�@�K�#��y���!��(��C[/oՒšAf ��y�� *wx9�t�H1d�*�q��6�y��_�n��&E�D=�����,�y"D �*0��P���<Ř=� �Ī�yB�K�~D
uL�41N�P��y"�Xy���� T8_�r��)�y��Δf�L0�k�8Vb4p*w,��y�.�(>^ֹ��Ԉ�5"aU��y�ϱ=���-�0E�rͱ0c���y���np���O���mI��&�y�BA!~�|��#��u��Y�yBm=WJ�U'�(���a=�yRcH�b��Q���N�6%$��y� N�I��ٰS,A�^�v�H���y"ϙ��ޅѲfW�V�RA�7ؖ�y��Bs���	[�B���l?�y�,�0�
$Ђʄ�ZT�����y��1?Vl��އ��кCX�yR��a��Y+��	�v���ԇ�yb$� pޚ�J�	��n�S�L���y
� И��(� -�=Kw��:\�X�"O��Ó��7���Rb��O�>hs2"O>-�"ͿM�D��� �`�;�"O�ɠOѻ3~9!c��-L��m�0"O�LKA�� x�x�!o��agd�H"O29�ׅ^�0R�"A�՚d`|��"O�E�'eܢY�:�Ag-��qs򤰤"O.�1nZ�9Ij�:���H�"O4@u��$Ed�	*�e�x�v,�d"Op�a��qB�2�ᑹ��5�a"O4�L�?��a� �9T��B"O�UX�F��v�V��Woۃ{V ���"O����W�N�{3�]
E#F9��"O:�zTK�B1Z�c�ylr�"O\� #ɋ�'pm�DE��1���S�"O�xX�ˌ�}0�]C��Նv�(�u"O�����?��H@�B[��-�f"O�T1ԏ�	uM������4�a�"Of�S�]�-���*%�0*��Q�"O�uy�l��E��E/^�4u"��"O�}3u�_"Vd��#$\C]���"O�M8b�Zo�q)ǎ�62=T��"OܙB�+8����ц{"�\*�"O\��)�&.�]�1hڏe"U�v"O�Iv-O�U��=��D��s��2�"O�Iz���
�H<pt�̓\ Љr�"O��p�G���A�鐴�"OP�A�A��m_
�y&�V��X!Q"O�4��F&�щ���>p���@4"OFи���rĒ%o�#b�>�B"OL�7�g����W��� [3"Ox��T��h�Cv�ϝX����"O�\���!�e�GD`�)�"O�P�̇,B�ʳǓ�v��Y��"O�4!%��e��6'ާ%�����"OX�34EWT�A�HȚ+�؁�G"O��QW�C:Vp��F���"�!6"O��0Ѫ_�H��w�9k��2w"OrL�P�	�бs'���\0^ثU"OJ��Q�\�{�<�҂Kߡ)�8��e"O48��V�7X )��i�@Sf�A��|�)�ӎBL�s�3@�@"G�Vb���ȓ�z��a��yĮ�>$�ȓ]�03a��U��ᓧi�d���ab>�R�e�V�a`�JЁ���� R�y�ǚrxXY��G�~�q��w|��7X:�*@&�D���]��
!|�`lA=%Cf5@Fmɍ���-fH}`g��" 8�C���w>N��b6�1�����-�5@�&N)���ȓp��]�a�Ɋ/j"	0��КE�ԆȓKn�����Ϧ͓�/�=�ȓsG|��Q
5o���YV�Je�t ��X�x�0vƋR��S7�8&�\���@)<���$�� ��5�J��.܅ȓG�PȚx6�S��v9*E��6�&��Ř�#�$A�Q�.$�d`��&�<!�V�̨��x(��=�)��;������#ai��hQ
�R�섇ȓY "H�'抓�&�v釾Y�r�ȓx��;�/���]��ʓ.n�1��-���@篖�s~J�)OӧQ�ɇȓjE5�3n�p�!��M�����(YM�D&�г��Qn���S�? ���KJ�@�r��g͒O8\KF"Ob����D%: �Q��,��t�8�S�"O ���U��6�q�,Rp���1"O�Xˆ���`�q�+?RZXX��"O"�i�GH�HHS2�5(A�!"O�� 4"�;(n2��_
4�j=pr"O��鱄E��3G�_�X�,�zA"O~�+��^�O�n:�G˛W�4�`�"O�y��Gϱ6\<�5LGH����"OJ�C���
�41�H�6<��Q�"O��yC��zO�x��
9T��"Ox��M��I7�}ˑ'����r��'K�<[��T����O�� �b�(*D��ke��+�m�̉J��jD*D���&��"���(?K��!S��)D��2T�\�=Z`�c^Q���4D�h*E�1<I��E��S��k�N5�$7�S����څ�	OEz4���ݿ�N��ȓ;�6�R�X�驁6)� U�ȓADN1h���;,���A#$�/vq��ȓV��u��(ֈ{�H}���P��!�� 6\�s�A�b򔵰��rC�ɠ+���V�MGl���ї`��C�I�6�}��%��Ik��N� ��C�IBdZ8�ë�%t� ���E��C䉔+B�#�\9!D�*Ʀ�\>�B�I�VXT(����\{lHg�C�_g�B�	6�J<#Q�W�y�J	2@����B�I�Bu��8tF�[\<����&8ŘB�I�f���b@�"9���
ςw�lB�I�z+ؤ��/�!���uN�qb�B��4Z-P<+�Aˊ	��/Me�B�	$�4YI�1 
��G��X<�C�"g����ʋ�w��������;ͲC��g�lH�S�s��\�&��l��C�I�X]�x�Ek��"��HL%6^tB�I�'	2q�c�w��D B@�\�jB��$����&ś'4��F�8�FB�'_"Z1����0-9*k�L[�<\�B�	o��p%&�\�x����<�pB䉫&�򈚦��-}p��7�� ZU:B�I�K�j�U�H$=v�	G��P�fB�	<��!�	B��.��f֥\��C�	�;�BTs�&���j4!bHڇi��C��2\�PD�dB2���چ�W~�4B�I?^�,�P�ޅSG�H3�٫WMTC�#^
I�C&�'st��4
��S80C�� v� PY@�ݠK(���C��,WP=���N�_�eS4��U��B�Ɏ⬉7���zC2���Y�",�B�	�3	�p+f+�(j��(#�[�|�B�	OTp
@Z�ax���j�AF!�dB=~0P��.G:&g��J	_�n6!�D�Y���Β򍒶JR��b�'��$��D!B� ��2���A4�'a�M�d�ߍ1c �Y�G��9!�T��'k��1`L=e>:����՞���P�
���h^8q�:X�ը�`���(,�\��	�
v��u,�>��ȓ6�b�Ӏ�\�z_0 w,H&�LD�ȓ$	��w%I-1�ɳ
�s2l��p�E��l�6��I��iY�6��<�ȓ���z���5n�Y���P�[�"�ȓ040��G�?Įi ! �&8 씇�S�? �cp�Թ{\t�8#B�C�H���"O��K�A
=)�ԐK�I�e�M�0"Of	FO1�4P��FL=c~�h�"O��(S`��,���S� �Q"OTqJF(�&`LR,���ʻ@;�x�"Oh�� �C�<��eMK�?􉐦"O����`�}4���N��a�����'ޱO�xRE�@a�92'�
��]�"O��ZRDY��*�3�4L��"O�a�R��5`�(��P� ��Ad"O"�!�$�(����p��[�"Oj�!&���r�xع�]*@�
lA"O^@��ˈh(���\����"OZy��h�b���3�M�Ht�"O`Z�̈)FKr���ިJ�Z�"O�Đ` �	?���ʕ�_�ZB���V"O�@0�M��LI�p,�W!�%��"O8��&���0�Y�f��~�Q�"O������W����$˃�+ȉ�"O�U����>��)�	ӈq�H��"O��IfNG)��1����|�N�*�"OJ-�a�J�uax��a��Xˊ���"O�9	�*�z�t�M���"Or��s�M��D7�����!"Oܭ��A
j\�m'�ϽAϾ!��"O24�F��*M���85��h��"Ob=!ī�6�	�	��N��[�"O<t��kZ:����D���1d"O��k���)���SǕ>�d�ȓgǒ�@�Ϗ"i�@a%g(^~���%(1�����l
��I�>��I��LZl�CsO�.7n���
4�"e��}ה�Y�-�l�b�A��Z�R����ȓ3��tYKؖ4�9@�C�����=�$���F�64�Ā�<�8��ȓr�22��Q�u�(ib&�-Bq
%��?��ȓ��[jh�b��wY�ȓ�d�!	6��k�͊(C\���VU`%�bA�S�����&
�Nq��y��)hG�ՑC m��]!c�",��w�z�֏K?SY��J5"�^�V��ȓ?}�E(3F�*��������B�]��b(& r��<Q�S�ث,:�����ׂ;�j�PA��8N|��iǍ�F�<�%f�9���w�ϝf���@'c�y�<	�9Z:��6��O
�5� �x�<�"��d��P�a�7T��@A��K]�<i�IT#İ�2�L�8]p���W�<iuf���<�ңjW�Z��� ��~�<a!����ѥ�#P8D�"2�S@�<Q��=l �e��/�(=���z�<�CB&1{Q�#%�5ߞ��`��_�<�V�A0�D�(c��c����1 FX�<�6�Y2-�{�d�7d�	Vʏ~�<1>��K�	�1eA*�q �y�<���O(��@�a�(W��|a�$u�<ч��+LQv$����xyyU�m�<�4'��0Ip,��x7q J�g�<94dĚD4���Q��>L)
0�V%�h�<�bN��W_��h6�O?6�PX�jIN�<�2���Q�v�c���#w֐���FH�<)��#�6p����+�\����Y�<���1. `y�C�RNh�o�A*!��ҬLVhy��c+d`�-*���G!�� ��@�$�8��1��)Ԥ�8�"O|�i�k̆J���C#V�'�bH��"OB����4���`� 	�S��!"O.l
�G�o���("J]!%� �"O��KD�q�!2��[�]ĐHw"O�L�U �2�=��a�I��Ԙv"O^c`l�$t'Z{��H��X�S"OF�b�h߶B$`���΍4Q���A"O�����I�5z0��RN�1oO���"O��r��O8w��ȃ��/G�tj�"Or|��C� D���2L�pԜ�b�"O���s�ԲS��|BQA��yK�"Oژ�f��n���@�?U;z��"O��@�E��Wb2��v%ÂA*�X��"O�#�iT�Sn��#E�\=�p��"O�UX��/0�0��QDTa\Z�ؕ"O0�y4���,�h�mMt�b�W"Oȼ�"K�2��Th�6A6T��"OP����/G3����,��H��"O|����r�赪�(c��	�"O� `� B5|�L�Y�&Έb��K�"O���DǨ����^���)w"OH,���74FJ�vj��X5PP�U"O8����a�z�c��-)�k�"ORĳv��
o��Ѡ!��wF��"OJ9����
��3
��o����3"ODd���):�pD�6I��`�t��"OrA��T0	*�����2$�H9e"O0�!#C�eDx9�aKƟ]�e�e"O�Aࣄ q�|�&j�	>Ve��"O� �l�|���8���{���c"O����#)��C�S��m"P"OJ���4�0kp���tE"O¹Ir�<l8$�	�̈�k�I�g"O88�V����i��E2D<��"O���w��K>%�7�i�UJ�"OMPԆ*�t����2zzLa�"O�zGr�^)�GA�c� "O�qj'��`�&i[R�[ib|e{S"O��򕦟Q��Ѣ�_$k�j��"ON�*S��|5l��RÚ#(��r"OF]�̍�ƢuS�T�c����"OJ���"+p�2'HU�{�0"O�!�̞�0	"T٠��j �!9�"O�eA���.�����'
�u�. �'"O6�hf�)t�
�u�F"{)ND��'���#a��C7���$��	��|�'��\�D��n���
I��|{���'��(��&Bur ȵ)ʇ~M搀�'Rĉ����?h4���v��3�'Q���s����E�0Aq�f1�
�'b8!Pb� �M;�X�`+�7}G��'7긒�GF���UiM#-ehq	�'k�����62M���Ef�+G*�0
�'���u熺T�2��`�K�(�@A��'=�!��Iˋs��e�2�'j	�'�m�U�e� �9%����'.(`�4�Ɔ ���I����,v)��';�!��פ;��X����6,|��'� �����,g`85#M�����'��򫘅+��i�c�:�dj�'�� Bfa܋L�z8�v��,�u"�'�D8HuK�VPZ�rV�δwݨh0�'��y��7BFDP���<vޮ,
��� >� $�"���'HB#�V�2�"OKg�$V=�� �-C�1�2��4"O�0AC�[<�)�%b_�a�����"ON��U���5�P��qQ*�""O���AJN*,�@a�r���e����"Od)b��uN�� �PZ��"Obm��.��vD|��.E�	@6IPP"O���#�H�^-�<r��_$*=h"O�(�F��_E�a�"�6I���"O�5��J֬(S-{Q�:* ��"O��0��]5:[(��M$G=�1�1"OĤ2��:Z���@|���e"O4X�Câ6���K��ȳ7~��Ӑ"O��XCݺ��0���N�Vc�q�b"O܁ �`�{�e���[�2b�1��"O���Cƽ	�f�"��2t^̻r"O�X��[$��a�F����6"O�iKń��Q���s�$��]��I�s"O"��+ >��3�$V�$�w"OVyم�I�M���
� ]����� "O\��F�: ^H�1Q�Z�fh �"O"��#q���t�[����×"Ofx���H�j�y0 %7Re����"O�i�nަ0o�p�i��4Q�C"O����E�&�u�G�C9Da��"O04�PL�I�Y�0��1A؁c`"O�)P�&��A	�e.F��P"O.�H� S760��ǲ\'�
"O��(U.S'��� P�<!�"O�84 �N��9��h^�9�"O@x� ��2%>-�����&��"O�0�C��60�$9S��~��г"O
P�h��0� H�!��$"""O�1��¯]��'�.��y�"O`�� e�-$�2�)WdL��4Ia�"OZ���GUC��puB����A"O����W(\ΌA�
�S��da"O� �O�Eď�l70� ���"O�h�dMS.�b�z���zy�5�"O8�mš-�ȩB@K����mʳ"O&�۷"�5'h,��
�1�f�p"O���'�o�&JDǒ�8̰�q�"O PJf� 8�:EO5OrA#@"O�5"��q1�x�ţ��Teڄ��"O�HB�Ǆ1)-���1-[�-L8Ԙq"O6s�O�=S�	�7��-8|l�"O�zGi�j�D���*7�y��"O8�Ѵ��J�6�vǘ��Ի�"O�
3/�8s��J���p�V�a�"O�1Q�k.6k�LJ�Ƽ+�6t�b"O0���+'!bej��޼3�dT*�"Ol�1W�ɨ~R�<�GT$Z� ��D"O^��Ǝ]�)��i��������W"Ov��ue/^xb֦\!����"O.I$�����J�ʹPq� k�"O���CɃ4��q���o�ޤ�f"O~	��\	i?<���p���B"O�e�?�4��͖ �<���"Ol�C�����8RbG�_%�!��"O��Z�:=�L�9���7���"O(	�5>�j�A3͙#<T�ԩ&"O���D[6a�*%�"X�SbX��"O��t��2D�l��`B�[0����"Onl�e�I0.A����II6#�\C�"O� \Hz�`U�k�`���2���"O^�h�P���4��M�d�Dp�"O��, �i��T9�Z�<D����"Ov��wIF:�L
��S	2B�F"Ojt����	Wc��P4�0��:�"O���"C�w��#�Öw�N�%"O4�[��۬��=P@#�0F9җ"OX����=�D��#��f X)�"O~�q��Af4
	�s��?Pd��#"Ox��C�_l��c�.�''
�����c>e�d���x�d`�.�\ytЁM:D���&iԒ`σ
Ǿ�� S�y�!�d�2!x�r��/ �d`Ѯ��0��'�a|�d3Lcҡ���7��-��BU�y�ImD�II�Ϝ>y��p�c�.�y��ӈ/�<`q�C��T0c1.��yr��2W6l�[���)�l������y�WR^Q���2?2�B˔��yr�M2S:��"��	�
� 3aN(�y�A�l�*�S�,��eO(҆� ���0>9`P %;@m���6��̨u��d�<) �
�N�JUDH�7���v�_�<�� {ʦ\r!��4;�\��d�<����~4x �Y�Fo�3�Jx��'5��H��ғ/-� Y0Yȥ�	�'z��T����^2z�ɋ���$3�O���M�;&�H#��c���5�����2BtXz�a˭;d���#�O!�$_�d����$
?'Pʑ�5gɼ�!�D�Du��٥�U�~�N06�ΰ$�!�dZ�:e&����2L_�� '��x�{��'��I�m�j�j��ȧ�b${e$I�3iPB�I�~�v1Hb�0"Z�9s��6�0B�IO`	Bqn!/<"0�C�G�d\�D1��]�O��2H���ږ�];�i�g⍭o!�D54�f��w�þF�R0H�6�!���#��x@���r$�Z�/�!�d�8���z�k�&a�xݙYaصϓ�?����d�#p�:�/�SN��EQ2 ~!�J�T�Jͨ��W�\�t��f�`	!��]�E��!SmA�v0dQ�-�!�dt�N	��3s�@�k�A�!�Σ~R�rvi�&D���8g��*�!�A�\���(��W�pؓю_Z�!�Ęqk
�p�f�v��Y�e��<�!�*_���"k��U��]`��܄?�!�$PS����6A�����	�M�!��ͳ"�E˃� �+V�5"@�!��$w�~����VVP�a��&}!���5�ȴcE��:r.V,q� �%k!���[���J#�Z1'-�5�ǜ53p!��Ćc�=�D�?�<A�"�	6d�{�Q���L�HP�c.o��ܑ���
=_�8�ȓ�
�6$+t�h�ӧ�օd�nh�ȓ��u1����k) d�S�Ţѩ2D���r�� �4�BQe�l ��l$D� �4�5$1L{�7-ʀL 5�<D����E*wd�4�p��I:D�t��-K T3 �R� E�af�
��$D� �T(�D�6M���B�d�^�pp#D� ���׈a�=��K6�]�(3D�tH��"$
r�� \����>D� j�`^-&)��́y̤��b�<D��
iٿ:�F��4&^@�>Y���;D�� h��34*����l�?4�^I8�"O�5����%Ǡ�pq%H#_Z!�"O~P�RB�Cq���qĄ�pL$A�C"Odz�c��p)q�Ӛ-$� �"O�1c�B��w~��uaFPp"O����&��x&x#F� �,��S"O`y�!m�
W��C�g"E�I�"O���U'WqN1� Y>GW�ű�"O��qCɄy��(ha���y��ڵ"O@5�G�1�MH�	�f�򈢲"O�ͱ҆ɭTa�X��gŊ`UL���"OJ������څF�)X*�Qg"O|��t-IW؎�b�D\ L���j"O�`� A������"�u�:i��"O���eA?��6e�/F�v`q�"O�(w��X>@b��D�d{ � �"Ou�4�)G�5�,�$
���"O��)�� ?<Ĥ�	�#c����"O����$ɇDf ���hڍ 0��{ "O�	3k�k��q�h��g @��"Ol���!
|
���d�R�̭qQ�����!V�v@{U���6�����a�4C�	<<��� A͟d���%�V�C�	�7/A�F��B`�)H�
VӲB�	�}sԁj��\	�Qʑ�� ���`�@�xdʊ$��C��F�-���D�:���h\�A{e�W"�P�ȓYuƩ+A[D�^i��)�I��4%�ԇ��%;��0a�N�V��}�5���Q�bB�I$i�P��W Z�p{Ul\�J�b�?����ӫ��yg'������-�'��{b�$dd|P�F�(-��9�!G�_���IN��8��eT&sgbd-40�`��ѭcUB�	.1W(�!'t�e�VI�"S����<?	s��v���0�e�6XR�W^y��'{f�KV�t�\}[��ѱF��UK�'P���C��!ub��JA+ �+G�hA�'�����6����%_(�,��
��O�d��G�1�b��5�ށvk�U��S����	�6�R�A�-�W���ɤ�ť8[,B䉡n�b���1�l<���&cf��$$?Y�n�Rnj}��/ņK�DpQ���t�<��W&H��u�d�(��uSFk�<ѡ���SԌ�T醋z��5QFg�hx�dExO�5�C��D���sD��hOjʓ�O´2�˃Q{6`q��T�5=h�_�Ȕ'waz"& �O-Z��U��B����[��y"�U�7u t��nC|���C3�Ԗ��?	�'
�$#������})��D38���'�.y(cʁ�X�����8'��p�'c��ٓֳL��d��fD�1���3��?a�y�(��*���+B/ۂx�ިsCɀ��O�#~��gL�>̌Q�;t���s�z��M�̺�Z�28Z�l�M!b�q��/D�8P��]	��L�ǫE����#D������~�0���	�-E�i0��"D�4Yъ�]&�1Wfć`AXDF!D�TAu�Ѝd��	��h��^N6e�č4D� �@��6}?*��H�/�K$ �O��0D{�O"���'���Y�s+�5 HA3L>�	�A�X�Z�F8x�b��d�ȅȓ*��i�,5���hw����\����bXA�o[�JD tP��Ғf ��t�$D��X&E[�2?x�C$�ó�*\�d7D�� .Ys"��>!��abbŝK�p���"O�,�Q��_�z�s@j��Q$"O��+ �:@h�J�,[:z�,��d�Ir�O��A� �A��D��"L� �'w*e	���%�ջ�� �\Æ��'(T��q�?��� �S��Y�'��]���T��แbN��a��'),�c�DATG�D1�	Ħ7�`%��')���-].+f�@��.j(���d>�"���j���E�&�\!p2�X� "O�f.À[㐄ɰ�� t�n=y�"O<���<�� ����]; ɓ"O����!�B�(�����	7��zc"O.P���a��)1gP�g|�(6"O�Us��L#_:�Y2 ��f����"O��qH�x���B/C�K��'"!�D�t
#��2{���LZ!�R�|���AZ���A,�5!�^�V4҈Ȕ�B)�du��+*(!�� 2������u�Fi����.w!��z�N���'ߗo�~�3P��?�!��+m��}��E�g�Vz��Y�S�!���\��(3(:��%XԈR�zl!��$L$		�!���9��B�Q8!��
@B��E�Α	f�h��Ļ+W!��Q�F��ƊL9fW=9p�H�	!��El^\���W?bTr���`ǀ^[!��,�L�s�]=0���#;�!�D��J�tp�Q�ď�a����A�!��N�����J�^v�U#�L�n�џlF�$E �b����V�B3Pzx��cҪ�hO���i�!E��c�C*XF�����!��>8�P�ф,�0.���N�h'���'�����Ą
�F�h�ů5W�e�e�'�!�d��=����4K� .T"��L�q6!�$U'Xꚜ3`��;="���u���x�!�@/Z�쀆����8"ś�z�@��?��|���4'�J�sT��P�
_�����D<�'Z�8#��N� ��-	�b<ܘ�ȓ}�]䂅!�d��U�����	�<	���#o�Eɦ#����Sp�� ���j	fL��ؾ�2`�p-]�DjBP��Rw0%�1�A)(�L�I3*�2xb$���;J�ɡ2�������GV�
�Iu��˟D�?������R4�P�gC�aYU�`��ԟ(F�tIG�--���̊�4jx���E���?����%*���%F8���Sh�3M�����r��B,KN�Y�,�b�> +��؇���VY�2�F
$�U�����?B���9�L��%�]�{L���aZ�b�M����<����32;�E����l�vI���ny��'j��b�	^���f�\x{��$�O�"~���#�~��򪁌_{�$��
�i�<qvė�A4��ab�Dq�c!��c�<���'`��/q�~��2��t�<Ag�W�)�H����'\VQ�S�g�<Y2�1C$"'N&�����c�<1FA|fh$:p���",<��'�]y2�'�B�K��q|��X���*A�Q	���5����re�:Pc��L���{<a`A��I�H�YV+[���9g�N�<�P�]Bn!�p  ;c_�@1jQH�<�FZ%*��݀���9mМ�V�F~�<)1ȝ��x����5hǤ��V�Yv�<� D�԰Z���@ �0"J!��"O��q� ��vt�z�F��Z��=�F��ȟpE��	�.g����5�Q3���҃�]��y+'t��X�!�J�e#�E���y�����k�醦H�����Hٱ�y��^-Q0`M#��J$BFI[����y�ϖK000Abȥ3s�8s	��y��Ǻ��!5�T#$*�aз���yҌ�$`l�BP��!���J6�)�%��g���Lȕ<!���]x��P��V_���U+��0	!��\�nqf鲒�^7RE���J�$y�!��:����g�a3]!�)pq8�'��l�+\�P@j����>��z�'ޞ�k�8`ٺĢ``-] e����'�ў ϓg�v<����w��mۣd>TK�=��e��˓'\/w8���۶7��ԇ�T��)S��5I|��P�.,(���iXN�(�A�v�:q��l�Z��ȓ������(�i��\({P@4��>=��+7K���C#
JZ=�ȓ<���;���a��tufB����ȓ �M�6H�9�h �d�۝9�.؄ȓ��E6Z�J!R��G��4ȄȓYv.�3Fŉ@�:�����	r�q$��	V���(C]�k�L����!"�L�&�"D��eʆ;Re�,P`�
��x*UL"D���*�������@ e�'B$D�l�d�atR1��ìd"��C"D� �*�:��c��*r�@��ì D������im��+�BC�_\(�7�$D�#$�'o�l��C%U�d9��$�$�O�����hb���!�#O�dY�� a�!�@��Bp)�"$WP����_�M!�d�t�2�鷢]�y��B����r�!�dȡ3��a3H���d�ɦC�!�E�gh��]�Nm0��@�:�!���YNq(t,ۗ����*?;5!��uG�bW>_��p��^5/!�ď�vM���a/ T�8 �7=_!��	�b_��1��A��dd� \l�!�ߺ_v�����C�X���=q!��]�[��z1/֧'���h�/�R^!򄒝l0�ĉ��ؒ$�NP�p$Yq+�}��q���p�f�SG��#!N�B4��OZ�D��'􌘛wTFɄ��퐜"�n���'�Z�(�A��,�����I�z���r�'�ax�
C�z7 P$k�>y���PH���y��.���-_�o0�#��%�y�k�1����I:�@�@7�ʋ�y�6��<��ڌ68�5h�K�7�y��ɚ8ؖ�s7���/0�b�G�#�?yI>�������IG��\��	32�x0P'j�-cfC䉟jev����Y.&F��0�\6��C�ɍI�F��&aX�wx�) ��]� B䉉\��i��f@�HB-+�B�	B�.|�I!r(<�:�&�F�xB�	 e��x���/+����,ݤm�NB�	�B��lQ���="��������B�ɋ1Z����?r�D;����B�	�.'�,{�L�5U����ϙZ�2�$��I6>���R3/�!��s��
/<U.B�I�X:*�xSEӎs@��`jԯ2�B�ɖr����aE�;�X��$��B�)� �� ���&  ������Z�T��4��p>�9�k�1�PC�%R�N%���5D��Em?&|	`D\ryء+4D����IN�Bt��3[zi�u�O�=E��$���xI�Q�¹q2��#s�ЛS�!�dԅk(,"�A��$+~�S� A'w�!�Кg^��D�:��I{���
�'���Rj�q���[���YvZP���D8�K� ��g��=U$��FiJ�~r%�I|�����	P(�|�v��.e�#ס��^��B�	:R��t�XQ(E�R�6TLC�I�5i<¥mW��<�[R�ћ6݂C䉀g7�1i����	I6� ���}xTC�	�p��3�G�Y9�abc Դ>�nC�	�r���j��x�ވ9�͵)�T���7b^ze�Ch>	Ñ���ee�L�����*4L��T�Zf��2z[�5�ȓ\*4�j�-��:���f�(P�J�ȓo�*H�C�܂ ����Æ�PAL���x�$ۆ���]r����Jb�,�ȓT�!Iœ�a3|<��IEML�ȓz�T|*Q��� �r4�A�݋a��5�ȓ,n(�v�4D��`��ET �dI�ȓr.0�'�Ή'�������{b���ȓ9r�� В<\�l�POg[T�ȓ�RɈE�^~��[�-�=�n��ȓq	�z�A^���k�)]F�(]�ȓ_?��$d܆S� IG^Id�ȓ�: Xw(�fu�Y*A�6yڽ��Ie�'"�]�`�_fn9�t�G5h��E��'�N8����4�D9�LD#*�V���'�X��W P�Ҹ��V�4HJ
�'�Y#̨~�Pw�G���y���g����E
0� J��y��M�2L��㥡�?��p%���y��6*t���珖n*���߰�y2�^�!<Ȍ�K��e<8Q8����y)MEl����)\��]�դ�y`�U�U�1J0R
Ta_?�yB��CLf�B!�ĆX�\s�H���yb�_�x�4� ��:s�������y«�;�l�x�C!2_���允�yr铭=8�e锨ִ<�����&��y�&(��\��I�;pA؁��8��'az�CT�}�@�8�(��]@�1�-O#�ynHA�a��/D4����6�A2�y��ρy���%)�ҵ�����yr,�nl&���gp�XFh���yR�&h���[g�N�an��ӫ�y
х]���H�χ�f.�i��ʖ�y2(ýu��*��i��i#sdձ��'Paz	)p�P�Ɲe�hL��n
��y"F���Lr `�3a��
QD�y�0�����욵p���8`��:�yr+�2�4��j=d��P��ڣ�y2�!	T����"ѰaO�u�&(B��yroSz�x��!�/"`b�a�mG+�y2GC,N�di��˕�����$H"�y�@&�HAa��HPfh��P#J��y�� 5,/~<q1��PR�Щ�)�(�y��I �<I�P��K]��r��Q��y"�Y��R�׫6L��p���X(�y�Gԫm�rcHҲq��{%F!�y���(}���R�\�J H@-�y
� �-��`��ijz)�eQ�w.��"Op-{����+�P ��)m�H S""O��y�ݫhX�04�����"OZ�20�ےWBj]㖪����'"O�+1,ƞmũYh8 \��"OpYkP�9W����� ��ۅ"OB�K�� �C�9!���)�B�(v"Ol:E�<7�X [&�"����D>LO��P��ރm^�Y���  ��M��"O��q�]��θS+�&Φ��'"O��"�
L��2��5G��4rf"OV� ��i������
)u�� �"O�5ImC<��R�f(8	e"OU���(i�B����9�DQ�U"O�I��l��/a�t�EK��E�Ґ��"O�Q#�LQS�Z`�j����A��'�r>O~�1C�ھ`��9�	޷/�<@H#"O����1o��A�t��m�����"O ��F�R5-��=� � e��#�"O�/Y�(s��9�-��qQ��"O
5Q⧄�$ߠ�� O�<�yQ"OT��RDҦ#��EH��������"O$j�i_�3,�a���6!��щ��'�85���[�"��,�/=49�'r�a�lG�rf2�h�=w:��	�'��t�4M��V���ZSCO**&�PC�'�h㶁��W.Tq�&�r	�8��'uP�	�@�#24�� ǽn(�L��'�rMѥ�*�I�W���T+�'6H4�R�R�y:Z�;)�� ��#� �^�e2��_{�a����+��B�I2!�h#�Ə4P�޸`��k�FB�Ɇ ���fe��j|�sө�?�DB�I�U���R�ڒA.�q�&'֌)q>B�	�-�`$�!C&4�����!
��B䉦B�>�C�!]�>0�H�E�*xI�B�	:��8�ǔ-X.j�ǪF5�C�/ �KE�͆s�D8�!�)[�B�	�����$��"��VB�=z:�B�ɐ_�Zը�� ,F�$ �럂<=�C��>\��]�"��4�#TE�7:#�C䉨#���yc!Z;�`p��ƁY�tC�I�z�2���j@�c}��rG�P3
�
B䉵�����ŘGM\���&�f|���?	���?��'6�~�Y�F  0� �ЙB��4��u�j�QgG~�!���e�4��*��HZvd̸<��W��� ~L�ȓ[����"H���Qyɛ2T�n���C����֐��Ip���K��7rĈ�U�8D�,��ȭ[����fZ M{�(���#D�t�H)1ժBfY�H�n�#�&#���Ov��>�+C�+	y��E��<X�{�� D�\x7"�>`Y |(�$ �G�&h��	*D���DoS6b���;&ȈR� �D(D�4���~��8c���@�r&�%D��[V���Ki�Q��Ņ����D�8D� ��֘L~^!a	�c2����,D��t͖�-p�P�C�jhd�0h.����G����		�䘑��"D�<��1"όUl!�$Ru����$�-s������
b!�ʵm���K5B�Q�Z��w�+Q!�$�mi,$)!��nQ� ��:<!��0I0�@&��08 Ud�<V�!�=�<�L��I�P���P�!�� &J��J�)Bth�(Q�9X�3��'��T6eX�H4\��"�N+
��-���;D��)!����I����5Q/�X�c�8D���A
4`�-X�O��JКq�8D�p�B?]v�ZF2j�P��ѧ"��O���J㮀$R�]�q�Q��H$�+D�Xr!�3�&�c�õ/��p�F�)D���MW�lB�4x��Dh^"Ppv "D�����
#xyF��D;V,Ru�u&>D��0�ֱe�fIXsf��	�Xĸ+)D��g$���,iQ�0u\�I��(D�XPWM�j�FM�a�v_(�ҁ�$D��a�jJ�L�e`� J�H����<��	vBH�#\8��fdӄԤ���I�<Qb�ҵ�7-�h��! %�hO����Xn�0 5��%���C"��]K!�ā'����o͈@�l��F˙�-�!�$��.v��JC�S0�
e�'�]�5!��˹t�m�р#:uhwH�j!�D\�%j(���h̦"@$h�jQ"z8�O���)���Q@nd�2�˰�� h�j�`a"O�Dx ��JP���Õ7�Qi��'��0��IT�|-�R�'`Y��r��<�M�B�Õ��I@T�`����d��b�h��Ť�
Y^�� ��WфĆ��ß��bk֌9;tir��9��IA���ȗ'Tў�>�a��H�s7��Qo�_��<s"�<������(��IX��2oT����O: 0y�"O��Ŭ�!O0x�����1v���"O�y�$'�
�ƥ�DF �t2���F"OᘱD^A�N�Y���9�ȼz"O�D��lY�	�FD��7g�8d�c�'��$�IOH+ѡ�0X�����/ln�X��D{��4CF> 9��*'��p�e�J��hOp��	@�i0��!�f�)4*A�� _�:2�O`��<ђ����}����"OR0�	,QR���D��ȥ	3"O&1AB@Y�^@�A�F
+���@"O­z��խb��x1�ehM���'[�,Si��\�.I�b��x@VB@Ht"�|��'�O�v馭h��P�+~��¢o�x"ą�g�'  U[��Hb����}����r�'KP=3�� ;:���ʶ]'����D ��M�%끕Bj��c�*8�|t:U"O���:*��+�eH�G��%�2"Oܬ��̙�=�Ptb7�� �:hI�"O��j�/6�
�B!
H�dU�ɳ���q>Y"�U��0��1dP&Wǐd ��3D��RQ�R'}�F�!��M���c�`2D����X�eJ��Wɇ�7�~�@P�,D� 0Fm�s�X�u�
;P�p�6D�`K�iL�,�>QkI��)�@�B"�4D� �G��H��[0� K*��3D���BB���0 �0lƻD��q!>D�Ԉ5n�)I4&��!�0�����!D���'�k����5M�! V��<Y�~�&\���ǈg��I��q��y҈�z�\�����9*�X��ҋ�y2B@"��]jN*~�6m�:�yR�8r�j���G�f���h���y������ ����cb)�y���c-���DQ(tV�ac�hH(�hO.�𤒘>���4�,>+*d�ux!�$(�*����ܷD :����)8�!�� 3�i �0CeQTֽ�$"O�}i@�_w�<�Ӆ�w :M�"O.�S'�����Ƅ5��E��"O�Qf��F��MS�����8p"O:D#UN�#;�����D�4b4���@"O6��N7t�����ӡ]��6"OR�I&�-V����/�&dA�"O�S@��O�����8�>-�q"O6=jDG���B�]04pYj"O���BG�	�x�qpb"B�p�"O�c��ۙrch�@p�J@j���"O��x1�s�"h�r��,�ʓ[�LF{��Y$J�𸗃 ����9C	ȴU��D�O(���O����O">Y���hS��(&� �����e�<i!�C
�֖��R�Q��[�C䉛[O�|Kr��m�
�rS�:�C�	<o���-���xIì��<~���Ofp��醤HYҭ�r)&]�`�HӦ7D��bX��ue�/k6\X$n�O���OB�O?9se闕h�Ro�S�tБ��l�	����	��x�	P�'�Ѱ �W�V��&n����'v�R�
�1V��2��'q�v���'��)��#��إI�h�q�l��'"D�F
�c�%��+)R�`�p�'�6���Q�?64(X��E�X��
�'VL���E�=�ba"D�o�l��)Oh�=E�T���S)ĉ+q�;l0���VdW!&fb�'��'er�'4��sW A2g�h]R�lQ���1G�:��0|2r��.=Y�97H�a��9�c�q�<	�_Y�=���G#E��l�FEJm�<)r`��5CBHRa��!-8y��N�<�O�7{��Չ2�U�F�P���R�<�wX�猉\ĺ 2*�w�<A�E�Jc�9���	3����%B�W�<�KN�[��U��1U�<��*�[�<�bhZc��J.	�1[�:娇Y�<�SfX�Oe^! ��XN�܀J�Q�<��ʟ��l���ݽCMzp��_�<��%�p �r�'�<�>�7�t�'�a����=,�&	jd.#t�F�a��O2�=�}�3�H2�A�o�l�l#l�d�<�fO�)[Q)3(u�S�#]f�<!��H+v�T���Me$��3�j�<1�KG�����K7�<�Pb�f�<QR+�� �4���G�;�����e�<!��&]\��B��9Zx�3P�X�<����GV���$&��8��+�^P�<�$m jb�+B4P�-���ҟ����S�Ft�R�b!"�;�A�Cyp8�ȓ2��w�8;V��Qʂ�s
���itfq�E�?7t�$M��X��E�ȓDD�!�͆`���� B:4> m�ȓRSЍ��X1Sq~ #`D �pلȓ1�����䈧vB��j6 W�F����ȓu�.�R�H͍����#�V!x�
̇�b��L���W^U���O�m��L�ȓ$8�Qqn +5uX@�fe�_��A�ȓȪe+��MH�psc�Ԭv�ц�Rh
��e%��	Jn��@�{����ȓjIn`�	P6 �� ��\,Z9��xl���Mݛ|� ؚ^礥�ȓa��H��νfYh����m� ����R�L^��<uq���/F]�-Ro5D���D#��u;���*S���!ڐ/5D�� �D���H�,=�����d��Ä"O�0'L�? 咬�ק��x�� &"Oh����ɳg��'g��N �� �ICyr�'1�������2��`d%��_�R�2�"Or�
c$6GY���CϾ-~pyJ�"O��@'Xኔj�$Y�:� "Of5��ȔP���㊞.���[�"O����.Y(P^p����I�T�p�"OD�A��Ú�p�P%e�����"O���k��Su���`�Ȝ	<�9��'�X1HU�H2N���dDR�O&D�(�P��li0 �@2w!JP��A#D�9�J�]�(1��*OP�c�+ D���fLG�s��R���(�j%�C�<D�h�A��Je�Kd�:_��"�:D�0�G& ـ�3�n�),Qz����9D�p��!@&�j��&v���d�8D���&�!6,y�����o���8��6D�|z�eܽf:�M�b��f����=��0<�!Oy�9P���b��-��!�b�<1�_�^A�8��6�zd*@�9T����i׀2���/MFt\Ly2�?D�T��+v��˰���Drq0D�h!V�J����1G�|����.D���D"|~�-S�gݚ%�l��5h7D�8����hۖ-��d� [`EА�9D�dx橘�H˾𠔥��M�� �u 8D���V���0 ��%f[�<��5D�Dx�L�/N8�k��ڦ5c|�"� D�����ƹf��U�Ø�1t�*ӄ9D���H�Ǝ��i�� l����$D��K�c"Oj���$��h��=D���c'Z�"�⦭ΌeJ0�B�.D���0�z)6�`�͎' ܋3�-D� �U���V�����(7������0D���ڇ1���%�&G
��:0�-D� V�m��F��-y�|S��,D�4��F�'I2f\�p��.㘼�3M-D��0k��H%zH�4��N^`�i"g7D��9SfU⢵���J�s�R��5D������C�0��S!H�K�b�i#�7D��)�%�#/:~P��M[�r� @�w�5D�;��ҋI���J?Z����5D��3.^�gE�8��g$f�42D�\��D��TX1dZ::�H�h�,D�tQuh�3,����Q���I\28�UL5D�$s�䞙I&�A�g%ĨX�l�@s3D���WɎ7{P��sK��l�P�*0D�$`%i�����S��� X90�m-D� ��J7|�f0��
]�TY0Մ0D��(5KH+p�0e�@�Y#Z�"틗c/D�ث4��]_����K�e_�P��!D�T�J�-�N���ʥvT�Q�`2D��Ţe��C�%�@*���b 0D�`�5�R?@$��Fk�:� 苵D+D���7$^�9Ũ�"�'	&>�^]���>D� ʀ��Z!�a
jF�`�@-xO>D�p�L�;X���=lZ½2C:D���U%ˠ7I����MS��jw�7D��2"�*���3#�3�jA�Ê7D���0A��`� G�M���6D�4s���6)��I�Z�؊s!D����JΚlؒD6�t�Q��2D���ؓo��)�RA���j���1D�� D��sE�#p�0p7���Q��y�U"O�p	���9�qaօ9s,Aq'"O�93��-����q�07� �"c"Oآ���hD)�,�5`�.�c�"Od�jTIg�'�Z
px;�Ñ#�y�@Ȫ.Yܵ!��2��5�SD&�ybB" ��G'6.z6])#�2�y�"�H��.�6��3f��yB�J�oS@|��g�J@���y��B{�&��_��tx����y��Mm\�r�J;lm�)Q�y�D��d�5K��e)T��_~j�ȓ?h�H�A� Բ���E�ڨI�ȓ+��<�3'ڴ�(�qe-̫Hr���ZK��@�-G�z��3g
$)Id���_C�H��X1�P� t���[:.m�ȓ1̌17)��4�E��ǋ2`�bX��4�<h�@�L�y���"���؇ȓk|1�cj�Ĭ!�,��	掅�ȓD�t�c��4hX&,i��v��ȓX�$ô�O�'�"� �쀲Dך��ȓ��0�É��J�%)U�;aP��ȓE\�m[�k"�MP���MZ�E�ȓ+F��)�#�"�k���f�:|��V7l�u�خOg�-�0�-�t��5��4	R$8RY�G�Υ;�����Y���ǋ]3� ��NN�@9衆ȓ�Бv� p��5��a��V�%�ȓd��)�Q��&��h-�}ԅ�:5h���K�Yܐ����N��ͅ�6�h��]4�=x_c~Esw"Oᱡ̅�B��iqV`�iOH)s#"O����L�b9����8B\�"O�T��l�T���&/]�g'���q"O\(����V��d�V�W�Ƶy�"O�`��BO���1wo^=z�����"O,-��&�+6�*�@\�3֖�CA"O܌�#�ތER��1O�I�bL�F"O8!c�	�!���s� � ��%y�"O�M��)�o�|���\����#"O��Q�4hx��	�$�A�"Oz4J#kj��͠#�B�%�q��"O�y�_5vbX�SIN,(�@���"O,��b���Dn (�P�ۤ�~hBp"O���v�4�R�Ӆ�z��pr�"Or�0
X��'� �Μ�"O�yS��7 ��@���3F�\!`f"Oh���9�$q�[�l!�C"O���%�C���;A��'݄���"OT���f7Aw�M��B�g��b�"Oތ���^ .��|��	�w�P��$"O��{7c�x&B�c
�	>�P"O.p�t@�M�Řņ��4�<��"Ol0�S!�����r��
T�4"O@S�qO�����[��E��"OL��w,_�#�F���	x��B"OZ��!�S+&e	lˎE��`��"O�I+�B��y�EY�j�,!L�`"Or�ر�ΰ<z^Iŧˠ8{
�B"O(�ɦ��-:D�:���(H�t!�"O��iF-ŉp�da��g_����"O�l�e�]�Sq��+cG8%T�d"O������/!0$�G�^9���C"Or���'D�3��r%��=�D@b"O� ��22e�!V��Q�R5}J��"O��r�n̽A]�M�&�}X���g"O�xC*.�$�x��&[Tz9#�"OXp� K��+E �Jç� �"O,Bw���{^|`�רQ�6d�!�""Oʕ2T(W63�q��$��3/X�0"Od��!V�Z�Z�Edr��"ORq(@��w��m��DQ�5���9C"OT�Y�5���8�� ��a�"O�D��q&��Պ�GkJ]*"O�A�a �B�>�TC8�i��"O<��� P!T�\H�EB��NӴ��"O�A�C�Z�N���Z�ȵb"�A3"O�T�5�S�H4���C*	@��G"Oi
�j[���9CQ���s�j]��"O���qh�����(6�I�"O.�;d��!~n��
`.	�o��<G"O�Ƀ�E�o� �9��G=!��$��"OT�Rk��P.�У{�RVp�<9P�ӷ1%�;��޵}�Mi�%p�<��l�:8�x�;+�}��Q��T�<q2/��]Tj5 �"ϯ%X�)�N�<�3�ǚ*�=P�(m�>�A�kFH�<��e�9���`�K�f�2�o�M�<���.R�uJ𬟝!hl�j�~�<��?��T0�͘i�|����e�<A��7vg���r�W�yV9CEn	]�<ɥ��Tf�A��^�=���"A
�M�<�����@ƃӘ/,ѱ��G�<)BEMQ\�y2�-"j��!!IG�<�g���C��K�HM7q(�(���E�<Q�*-	)�D)3 �>m:2ؐ��El�<ya�**"ʙ	C��X���<ɗȼl :���g$����hc�<��J%|W\9��Y�:�㔃_[�<y�BR�S�9���B�:hKQ��[�<q�gT4~4 P
�ˇ�}��ف��M�<��D�5D� d"�F�X��SA�<!���5\��"A	�Qv��g�|�<Y�/ʆT�p�K���,��u#1D@�<	G.Ŧ
ά(
���H�.ia�<Y#� 3���r�V� �[+g��[�<y�c9,��ͨ�LG4�R�����[�<i�i̩5R So��&��Tx!B��<I��� ���	�U�rtDig�<�go8y^lIɷ��,w ����H�<A5`�C6~h��#�$+WJ�#K�I�<��.�qP�iw!�	#����%�Zl�<Y%+U�@3*x�`ɱ'�@�<����� �PJ�	��p��q��Mu�<�7HF�R-R�p������V�<1/��*�Ұs�C�n�<=�eZmy���v��J>��	=q����G/�<e����<�S�G���$�j�cۜ�S�(f�����H�8�I�bC x3���t�G���	��p>�Co��A7�� ���2T� �Ơ�R�d.�S��	�>ᷩ!/���񌅓ښ܈�-N�<i5G�, �"E��zed�qV�#Ⓚ�\��%�.��x3� 
��`W"O��bEe[.�Qj�+��L�P"O�E2`�,U��%���Q:H"D[`"O�Dӊ��9�� )wF� "O|�g��K��D�Pb+�u�'�	_8�(ӱ�͸ �l�:T�K�`��;�7D�� �q��k�U;w��(��u��iQў�E���A�a���Ĺ"=��AD�����>���<I���Dz[t���nJlB#c�F�<�rG��9q8!�CC
�#&h�� ����P�=a�Û����'S��	��:@�'*
MBلȓN�l��/֧

v���]AJu�d�'��O��|?L<i��yi<���D6�v�#3K_�<e'�h&�1�&���u˂��~�<��!���zg �,%����#φ}�<�%ɜP�F��C`']!�x����t?���'$��t ����K$�X#V`<	��(`��� ��de��#��"\}��8�>��G�Q�� �to�:zP)Fz�'(����[�g<:��ա24�	8�'gdq���Z ev�W��7�%��4��$1�Op�p��0t��h۱(?Pz5�|�|��'�.���fS��&lC$��Ĉ���1<Or�bpG ��>9
1���cE��y�On4׭�	��3�¬Bv��H$ˏ��>��'�	J1K8d��b+��SLD9�S��Py�F�o��U�P��*YxZeX`��\�<�N\�~�JC�޺Q���{5�X�<!��/��e��
N�Nj�X1�i["fў"~�I�j����k�A��f^�a8J���>��@���.����f	rf���0=	N����<^����T�r�
R�7�O�O�Đ%�C3�l���	�={N�;d�I|���i�*!.��`Β#$��Y�&$Ä1�!�d٪>I���Ćl��cG�ў<��ӭa�̫���L�@�õX }�,C䉖!�05�b��2"��(�Ⴠ�UIC�	%J�����hN�\�".˱3��b�L��	��![Q	rn��:�Ȭz��B�ɹ|��+��� ��{������O���?�L~�+�^@���^�fyp�qt ��]�(m���t�O���F�ΏHQ"�#��ۯD�p|��{"����<іƑ��:	>R%P)h�&t����?��A�j��\�AH9	:n��q��x�&R�{6�g�Pe��1h'O���yB-��l�F"§Hk��v�Y��y���
����CE^�U�����T"�(O"�'���d'P|�9QD Y�BdR53} !�d\ql�+�*
6�zQ�7���!�D�?pj���D�%!ފ�#�,I�n�!��?dQɃ���!H�Ȳ
<$/!�D����ꧨ�c(�!�^2OA!�DS�K�$d-�M�y @W/q9��x��8�PJ,+>��6mB�~�(MC";LO��O���Ϭ4��	�Ko���U�2�!���:�L+��D�Mm©U�L�9���3���(%��B��^Eʀ%WoB�8e"ON���O�mNq$��4��+�U�D��'��}h��h���	b�@#�4����N�J��\P���m8",#g��`�V
O����X�J�pT#�*|c�����'�������(P�@c�ġU��@�/1D���*��Q�b'B�My��i�L1D��P4	�wD�݊�C�,/ܼ�C�/D����'Vg (]Y��E2e&���V�,D�x�V!E�H ��A�4���&D� �B�ƨ4�D��K�9H��Ѫ%D���Kр/iv	#ݶj4QY8D���SjG8'H����/ip.=��N4D��	�ǝ(������A�X��(p�L2D�� ����^�`]�v`�<EZ�@��"O��c��I�G��0ȳ��pH�� "O�<�4Ξ�K'4Q�#��]H�)W"Or�i���v��Yu Ǜ	�cg"OFcE!Z=D��ѪQ��=@����'��	V��R�^N�<p�ʚ/��">����,@�ΩÓ�F�6*���� 1%!򤖶y����j�� �З��I�5�S�OJ�U�!+Y	t8\X�' WX��'���4�۳(4bIx6�
x&����'��d�,/KP �5`C0t
�(�'f��k��^E��#�I�4�]���D9�S��I?S�53a"�;\�&]@�㉤�ynI+S� ڳ���jq�a(c!�9���p>!��� /��ZQ�(gT,hǇ1�D5�S�D��O����<�-�fN�I ��8b"OT�2���(Ue�/z8 ��x��$IJ�'�0y3��	��q��߄5u(�')��`�&���P�I+l~��ˌ�;�	V�4MQ�g-,��愙��T�v���yb�6_(�)�����А�H�?�y򋈝f��h �K���ݨe��1�~r�|r[���ʧ#�t!�枹v�0[�͆�npB�ÌK��������#7ޅS&EY�_�`��FLE�p��L��?�"5��"�L��&S�[�� 5Fw��B�	6w�JL
7N��J�����l�=���q\L�q%˞Vg��'ʛ0�ў,G�T�i%��s���a0b�:�뇯I��c�'�4݁cm^��m]`�%C#>]<���2�S��"�# GTQ{E�" ���؃J��y��Y�R��v��%a���� +�5I�v�=qF�i�����C*Q��@��XӬ�V�<I�L�dS@ SUgR*�2]Pր�m�<�ざ)M�<,vL�����a�<����9�4���$8��3.QX�<Y�^7f�였"���	�2�i�<�!C/]�*R�J���H�`}�<)S��>Q� �B�����u@2Hֻ�hO?�I?	>��g*r/�|r1�C�	35�� P�Ž.g�@��^+Pp��P����d�����eN�3}�ak�(��0|��E8I�c�FH�p�F�H�'=�xr�4>�$�JF��5gjmYN��yr)żo� �V�ʥ����A��(O���$�M
,h!�,L2=�7�ޙ3�!�D�>a��hh���9����C-P�!�}���h�Έ-Ҟ��˳z�ay��	,k�A�HZ�PeK���9��"?�q�?�'�X,1&�@�9o�����ڞg�l��3�t%�W��M8��R�;���'��'U�?��WN	L�8����ǻ<�|{&�"D���-X�I�.�� F�[`h�
�%D��� �"���N� Vu[5k%D���t!<;�0g�׺r.�IG�6D��Zud�,gd��k�?n��$�*D�(�ʟ�����)�4d�v�z�C)D�@xOT�\���GK�c�R`j�m%D��4ł�R��`Cg��CNPz�-)D������S�|��ՃS$��ׄ,D�H�bA�f�T@`өT�<(��+D��gO�	�a1�㍣��q�6-D����!~��3��Ԯp�a5D��P��ŉR;�b�C@���%�5D�����gX���6"č'��QCH?D�� .�A�狒d�| �D!ɌP]\�"O��j��%

�u�� �@?rq�f"ODp�M�/"��w�H(78�@�"O�x���58�n�IE�ۄ(0� d"Oޘ C��P��Qǁ5;�U��"O:M�u��\�Psd�E�jH
E�f"O�D*��J5AT�]�׮�f@�q�"O��r�)Ƕe�y@Ӯ�,c6���7"O�\"Trf塡���1!J(J�"O�`�2��0�Y�P,�+T����"O�M�c���*
�u�$�ƈ��"Ofp�fj��D�fa�IH����[!"OF�ҷ�ē�pxPM��Iz���a"O���_9�"��#H8+�.r�BC�<!T�W��|�;`�8_��Щ���t�<)gE]�p��QׁU�t�h�7��l�<i���#Fʨ���'d����o�<�t���f��q��%I:\��)�k�<���34=�� �^�Z���i�<��\ ?�j�8W��:
��Б(�e�<���D%9�|��0E+�� �$[b�<�ԀB7Ɛ3C��&gJ��#a�Ra�<i��޲~T����ޥ0�\�3GOw�<���Q�j���d�D�L����F	p�C�ԋ��3O" ��F X�KyP��<��%�on��r���Ҩ3r�RG�<�"ڮT�Dd�O�B�
���g�H�<���ԫ���c�R�D�Qe�Nm�<��/(<買�*vf��7�j�<�qW=�NpR�h�!u� dV�e�<y���+
�l��-��=o��І�Ay�<Y��٭JA�Xx��4H `2'�^�<�W��mZfL�`ԬH���#�MM�<�A��h�������{��-�AK|�<I�F��&�t�%#�5'T�4k�JQ�<��G\%2[J��S$�6��!�$h�z�<�pSr����R��4��A�l�<	�+ѶtU^12��ߋV�(����Ov�<Aԩ�pv��R��A��b�����q�<���J���\R�M'<:`y�@,�h�<1���G�2X�6���9�D�sq/�i�<)q��d>�M���4X��K��M�<!U�'>Ѩ����ȖAEhȥh�I�<9t�Y]vԑ��_	V �+�H�<A�m��
E��&I�:i�1�eB@�<9ń_4v`�U-��;��[��@�<� R5B6=���1,�j	p�A�<q���U9��u��h^�0� {�<	4��# NPQr�,d�� �l�<1��&<""�E{!ŏ
3��-�ȓ!m,+U��yW$����Y-8�؆ȓ[��iI�/X�O�M�Ŋ��!z ��ȓZ�&���b�v�Jy��ʚ�U����ȓ17B����ȟ��Ia�F�!���ȓ,Φhx2A�'�%JBOQu^؅ȓ88<K���<�)a����ȓ?�Z(�G�����!���]TX9�ȓ?WXa�)T�#���&�LN@|P�ȓ B�L@#gͣ5�=[$��I�6�ȓMc�K�&(1�j@�#���P���u��+��H��ԑ{������6e8�9/l�9!���3.�(ąȓDo�� o�'�i�C�I���ȓa�ڙ��A�w,hDP� �#�܉�ȓ5�5+�M�5`ʈӱ 1bhh��S�? ���iE�;g@�a�m�,= L� �H�p+1��� !���1%�*o��H��G�[��B䉏��U3���"ؠk'ł�,�찠���P^,�O��}��a����*N)S������	[��Ą�3T�A+;�JAz�$�`���l�q$|�1���J��{��I%od&x�!o��D�"�;�%U��=)��tl��:�!�O\��ri�
|
)��|b��U"O 0J��φ����Fŏed�92��٘8M�dX0H�/�h��A�gj�
�)��
ϔz�\$�1"Ojћ����[�b  �ި$� �����>\^�e�U�&}��?�g}B�:,fb4��.��=�p����(�y�FH^������.����Q����M��+0&@�e2|O�|�3��'��X�D_�!$|qF�'����E$D� �b����Љ�KD�X�dq5C@b_�C�ɠa��£m�|�@҅�@�++���7�0@�.�G�D�J�V�.��k2��'H��y�!V� "�pq��e��x�0�Y�y�m�5�* �K�B�>���ߛ��'>�$��&Qv�O�ވ��͕W�n��HN�.h���
�'C����HʾzgP
se���b�J���O��:��Y�|q�K�l���a�mN�(�lp!"#D��;ׅU�8w�<�e*9�2�I�&�rXT�G��Z��|�%ˡ-�FE�T+L�-K�b�ć��0=�Uf zj������,�8_�����˅��c�<D�ԫ��l�4�4ˉ<:�E�S�=�	�8�uɓ�<8+Q?ycC�ނT�(U�%L�`�J��=D�ۅ��9��hhpgF
8P�(f�T3ZD|��a�>�,k�����/dFD3�j:WK
�JE�S�%�!���z�zTc�G�1N!��.�8E��-F6p�~��1�3!��O�.�y>p��i<l��<���8Z�޴x�GI���r�'�ٺ��K�'�Р Q�ÏL����J�.��@��:j]� "ػdH��=!l݌0'�D�5I&>(��I���0s�L�?�0��������G'��,F~���`6�	
.Aj�� W�aK�>)A�@T�H@���艒6���
�A�\XU�td����0As��Oj��Ǫ0IHS�	�'t	H5�҆;��5�R���;�X�g*�cZE��ڢ(G��<��OA���Co%}b��7hBd`Ã�7	���$��,�vć5;4HA��K�uC��Aq�A�iAlp�フ5��O�8`��fC� a�K^�pW*��$F�$RVd�g��IY��xY��ș'�v��nK�z��0$���-pQ���"&*���NƋE�8�iN���`HJ�BR���'H\X��K�����5���a%G.�Z5�ЬB�iMT]z��h����,��.6�(Lc&-Al�<^��B��6؀��Զ�upb	�83D$�j�h��8�K��ğ/O��pR�'d�Tҥ�QF�% 4�����]�T��Y��n�'}���Y��J�X��u+Ŏ\��`�J�'<����ڟ.�B�F?[Z����$�0�@�G�z1�í-M��O�2ǚ�۸��S($2P��>^�n�
@A��J���Gݒ[��Ė�����_r�%��!
<[�|�Z���\��`�!L��u�W�R%8���II�u���`B�q$��?K��]j2�ć�0�� l<�Ð@�CW�ejrї.�� j2������0=Q�bǶ[�T��"�,{�#1+I�b@�@�>,J��2G����D��
�]�
@ã��.y�Ak��-�)���6eX����j���*�U�ay��ˀr:��&��)v�ߢhک�喾Y"5�`�� [s/Ё7�\�2+_
,�����26��SZ�\x�t$��y�`��y�nQ�,p��0F���i^���H,�)����"
��!�>5���E])%ђ��hAK��ӑ�ߝB[܍�mȨ:���d�=>���@�)+�=��n�ֵ��C�~�N�T`�q���M�s�E�"vnu�R9P��w:�"�ժlba�ܹk����&�#)eR���F�5������Y[�uH3/��p@}(��_�,��y��1��*ψp�"��A��4��&_����p�(��Iͧ
@m�t���1g���PH)ι�ȓn�j�R�bR5����$ߍs��<����,Q)JE	%�M�F��P��a�S�Z����.�>y%	_�g@\��sG�"K�6L���[���ae�߹&T���g�=^_�A���$-fxqraT8w��ەE�yl�h�%��4x�i�Oh��+s�ޤz��觋&�i8�aBO���1ZT��u����i�uӱ'�~��*�*"�T��fj1�O����O3K,��� �Q�P����\:� #�ЙR���A�t�y&	ä@��$?%*��T�m�I�٨R�L!F�#D���d�2]� H9��	J���� �^�Os1˵N�#[J���-��	��c>���.?�d#*\u�a�Q�('�b��U��P(<�D��vht��ԈV9b�^���)N�nZuq��G�I�n�3��5�O�ez��#Xh��&��1h,���'Yl�,��&�r}
� a�ӳ&�d�	��6V���B�O�=+��0>Y��6��A6�٤oY��v�,I�C;扷-i�#���w���2H���r�Ai���5D�p
pb¯&��"�G_<D��i*3�3�I:L`
`�d ��^�>�" DJ��P���+�h���#D��X�J�w�)-��P�6��]�z4	,9Ҝh�O��}�M|��:4+:�����ț�<켼��	�"������C���h�H'_��xS�"-��O�@�e
w؞8SA��;!ℨ�p�+-�4d�� �I4]
�
�E]~R/Um�0
5`ʺ��D�(�F�B2OӾ "ɫ�@��<�sLX�Y��)F��?�@�Z4=��{�N]y"��l��,Cf��V�i��@3U���կ�f(h�L�8�!�d,hD��"T
H���P�>1��F���bU��ڤ��̃�Ę�-��$i�ᚌN�ȹv�FN��z��~����'S'b��I߫|�|Ԛb�K�&�jh��P��?�Wo�,*���C�&lO4�PG	!а�@d(��cu�pR���09�@I!ĻX�L�l���1�Bɱ��b�x�(P���G��%���"1�B�I%��H�	/#v�;B��r��}2)�r���
�C#p�g	����@�I�/"t���9H��!VYZ$s#לOH�:@��&ta|R�Հ� ���'f$݉v"�:W
ݛ2�� �3�Ҟn%b�ɳ�Q�,�A!pK�.3f ͹�b��?_c���!�(y�֘�g�͸
*����/�	�V���ɡ�P���ԚrZ((�-��>�i���(~�A�e�L0����L�W�d��BR2`�$�'��ы�O�_q`��!)_i99��j��@�UGf���cђ<����1�U�^ul�ȁi�o6���|��YW� '� ����C2l?�����*D����N+�\mcm��A��I�"��L�n��B�U�5��0t���B%��T��)�D]bÍ������w0��c��L�@$Թr�M"��'FH�{��''Z�l�Hcb$I��N�D�j�c��?� ��Ħ��C�� 4��28�ȣ��?-���`���͉�	AY"@����#7����?i���:#�C��<��M�V���,N�P�h�`�U+$t�0Fl4U�q2G	@'H�"b���=q���	+p�(�J��a8�� z\��V� ��	���!B
�\)���,����GG���2�<��6��-T�&|�f�E�<Y��Ю+�l�I�.MA(�1�BG?i&#U)K�|i*")O��60k��g0V��D�&����V��qa��&|���"r���s:Ĭ��I�bh��a&�3֦� pG�s� .
<�{ulu��ҁrC��'�Zs��P��G�(:�:@�7X�X�s�l0ʓ�@��'�Q��!)E&�Z��4b�"'�u��Sf&x�e�q�<%%��H���0�)P�e\R�(2�6D���7� i#�Ч�řZ�XPie�5D�L��i�*Ұ����S���5g3D���'.��Ua:	RIè�@���2D�(
Ң@�8�P@��)5NdٗI*D��$��7$8<�s�]�4����%�O\��(�H��l�^�aؒ�u��
�'�ڵ�BB�:mٰ�ςB������/b<��I+S���A,�.�>�醤ڔr�C�I<+�py���:*X���Y�RZ����<�A�򍍍y��{>��������4Y��(��D��Ҍ~�[�cZ��S�&a� 
 �˙
�hx�O�&5x	�Am?}��3I`4�R"Z~��1�J�6�$��#��Z�=3׌=ʓr��!�A�*�	9d��x��ST����F#^��0�;�P2V�(�h�OأeA�[5D-��"�[D�G�A >Q���䀟.B�ʁ��������ee�9I}^��&�ǻ@EF|��"OvBB!�T��y����7G>Ax��Oڭ�	�ک)J��s�aZ$1��`�S-,,� ��o�z�L����'M�q�o��<)p�#-(%+4c͹�D�����C�$ƛp1Z�8�)���0<��'����"#�=R��)�#K�Q�'8�[��d�!�^ �D
�s����D�-�n��e��.���3�'�XQP3���ݣ�[<�dx����C�"����>�Ӛ
��z�jM%p�^�Aw!�87D:B��!'��b-ܷr$:���A�@��p�Ι���?�)ʧ9��A�Ғ"*E���*��9D�c��>6 ̓ �`gN4���7D��rTǘ4vE�P��/_;�6`y�I3D����HO���-#+ݢ\e�T�q;D�� 
S)��
�B�L�2)z ��"O�A��F�q�� ���3)"(�"O̠1c I�DO:l�� -x�v�Y�"O��  ��:u�񯃂i��=�"O
�6NF)y:Ĩ{�#I?5b�h3"O�@��D��v�E g �z i"O�}���?.�V��!+���"O$5K�e�[Jt0���o�9�3"O�0[�IDD�h��#.&����"O�\���WX��i�F�H1���{�"OҜyv �5R�RYu.�{�ZQ��"O i�C�n~0,�n�)b��͸�"O�dB�Ɋ"�lݡ��8%U@�"O���$'A��/aCf���"O"�q�NUH�x��c�۲h�F`8�"O��$"�R��m��m׫=��I�"O��qB�#<�LdK�f�>v���"O �A�"�~�c]����"O�� oO+J��ґ�D&QӘ5�C"O��Yw�5O�X����;n�$ha�"O0�qdԺo]�u�0�v��"O�Yʴ�N�m��i!g�;�X�A@"O�` S��I��8���N�%��ź�"O0�+�����;�!@P� IE"O��sG&=��[�S�V�@|)�"O \Y�#�=OX�Iģ�cߢ��"O�9#���y���Q�a����"O�� u�/���vb��v���q�"OZ��ƛ�LVFQ��H)�*�B"O\�����8:�B���� O`>��3"O�u��B�~�td+@-PW��I�"O�5�B�Ç3�>�� lH�(]p�Q"O(� �+R%heB�%��9c����"On�aF�K�Pj@x�TJ�3�lͣ�"O���l�=>�у�����"OX�ۣ��"��Ā��B�z�%"O0��*b�`��<�C"O�Qr�e?F�Ddq�"�����j�"O��ǣV�/��G��f�4@��"O ,Ȁ�C?{���S�\.o�"�"O�16#dY��E��;��qB�"O�t!T@Z�m�8!{�g�kQf��"O�z��!IzZp ���_���u"O(]���ޣT��B��_5mE@@#�"O. y��Q���5��cU"OnX$D�~��XB���]g2�ڰ"O�mDC#%�H�hGLȗE����"O�ē@-�0X���& �<:ѐhЦ"O�`��#Gk�y"u&͖Rd��p"O��0D�\��pQq�K�!J�p�'�,]y�M��g��AB��(0�v�j	�'d2՘�H��ؒҳ:Q���'��=i�n�)Z�°�Ր6f��'�V�c��2MƖ�i@K1]���{�'f�����`�d��d��gͲ�
�'����%��>��ᛓ�\�H�\	�''r��50C<iz�
��FV��;�'BV�Ӈ� 3���b���h���
�'��y�G�T�*��!�P�Ģe��9`�'� ��A�8K��؀G��P�:�'j�Չ�A�I�l��Gh���`��'��X�r�Q4>�ы�f��A3��)�''8hqA%ßj�D�1��˙���)�'p������h$k'�������
��� J����_K���QM�m��(+�"O������%5И�1K�%'��X�"O*Y;�CÐh?����������"O��U�&)L
0��p���"OA�nцv��\�bZ�(���d���>����!P�%M$(�6�ވb�B�	�?��������R�ޭ]Z�����H,r)4�O��}�WF̓���>�Vx�6��m2|p��/}�Y(�BŔ~��*�K@����m�	@��b��"XG�{<	0�b6b�Ry��ZG�����=� j�1]�v�����O��Q�(-�VQ�BH�|k�5�W"Ohr#�#�T]�EGH�f��{��$�,=����L5�h�X���iN2m�TX0 �N��kU"ON��a�1� { iE����d�ş1��I3�(}b)$�g}�̆/kި�vh�!�����F԰�yb�!.tJ�Ќ̚y���M;��AD�J=�a�9|O�ܛ�HVP�4� SH��v���g�'f U��N�"R��(�ɮ	� 9��!V��a@�Y>��B�I�o��Ā���+Mʨ��w�⟐�.B۴�E��c;"���8p)S� \N��DHT#�yb���C���P�1Q<�D3�B��y�H�%p��tDo؃z�AT����'zݰD�Hb�Of@��ޢ������PѠ
�'�.��T�P$~�W�ʅg�x�5NH�ȒOpٍ�Y�(��.�!����A�����23B D��чI�B�,�T��5~j�!��^x��
:@�|r��=O*~M���t�͙5��0=�DW8d���*2��t���4IΎ]��+]�Y;6�:D�`�b��-et����"fUyJ6手%re�
ׇ.�Q?]"s(@�*� P�v
	)Gp�uY`k4D��eO�1v�����JzX,K��ճX��08C�>I�]i�����Zm��	�-�dMZ)I�n[&8�!���f��YJ�	ʙ;P�c�M:,��P�I��b���i���#l�i�fh2Om~�SG��?/�x������?�����'�qY�c�O�'�vТAM��:�����.9�qxG��'>(X6)C:Z�AExR�*Xx`ˠ.5N�,R>q�����O�\궈e����6cקb�~���y��g�f���I@e�O�U��*ɃM�n�ơQ��h1#oЄn��$�dmX���0�M��
)��ټ�q��>�ċA#�/M"�����,͌ȳA-}���6���I%d(�	����Z"m�P��6\� U`S�v��5`S�	pyӅJ�,�9'�A���' y�KSwL����ǶWq���A�]�:�A��o�'>R�6�Ͻ'�$x����)��*G���
��ѵ&�<�V��bO��w����@ �X�� 03��Ͷ��dK�k˼!��?��L0wD�-gU�O���E,�ݎEC��1~�}��nI�]Ĥx9Xw^�4Zq���D���A�$�X�H�}"Ɇ;W&�|E�4FH��p��0N�'30��2A�.$f��zю<�Q
S��-!~�2���-�t�>)�;B�%)uO��yQ�4E`�,c�BB�	�+x���ˑ���k�&ޱw�&��Ҁ���$)P�Cc�k�-�|��`�J���'�R�wgM���UCGg�|2�l�ߓtv��W�H7�\�+�K<da4.�*�DU!�I�}�P�+��"g���a{B F�BN�z�f
�i�xx���O�4P�- �H�2�Z��`�@Ѡ��
�I����xqхԟ�rH����4+!��� {lV��P�-�����Ǣ\s���&E�
W*t�"(Q�9�~(��M zmQ>���R���Bc��:Pw�y���6y!�dX�0��A���2Z�H):�.X	U
�m�O��b�@ܲ���qO�:�:DǄ�
�O�:^6�q���'��jǮ�;zB�O1u�@���'_�R9�ӇDo؟#��U�!��9s��&g�:��4�W���gM����­�g��!2�z#A��'�)�g"O]���F�,�|����C�2'��q%Y���k�	iހ>E��m�VO���Ee��}��]����y"�+ڸ��J��l���+�d�'34���@�S �ϸ'>*�IG��	8 Qp�$�0(?�%"��< �qs^*,O�-�ǁ� x�rd�ۊ���K��?���d�Xa�%�+yH���'� �BH-�X�'��R�f^�/B`(�k� iQ�9D�� ��*�E��^���3��B	-��	��>�G��X��?q��e�h�d��T��/ ��  $%D��!��JN��@J�7���B��$D��x3��nT�P"�m� /��zs�&D�Q��l�q�v�?;0��&,��dSG̓��a|��ؠ�A&���,��.ר�0>�FIL.r�N��8��� �L
_��Ȱ�%/�J���{>d�0�C�G���'�"�e�?Y��#�rИA'ҧ{N�Mr���j�r�ZW��X��ȓ�f��U�0|��0bݞ�nIJ�kG�ZO��g�>����O ���ߤQ(x�JR�!y\Hq�'$4$���t}�i\�,��d���R�[ �a�B���?ٲ�(4̓U�:lO�a@V�A%*���
խAK
y���DP�@��<�g $?a�
V�#�$ui��`ݹH��A�mM����F'Y>� �/#D���%I��	s�ĐX��A�^�I�$��<q!�'��;	2�針�yW��d<̲ KI?Rq���R�y�x�\Eh��)'����`J%h����Մ@Rƈb*O,����)RY	�}B�����O�(��ċ0�p=AVA�L�j,�r��-�Mk�IpZYb�@ʟ]��H�m�����PgU�e
���u�'Ab���]�y����ڝȍ{�JH>z�P�ZbK\�zG�	.UC��C7b�?��� ��`�Bݑr���ವ�j7D���#k��~�P�%m%p��D�;����͐��?�vB�L���C��~�@%ȹ?q�?�h��ï��N�lL��莌l�>9#�'v`t��i�	�r�̖
w���c����0�s�Qq��\�Pg[>;�ly
��
�=FU8w�̗	�Ń[��O�����D
FL���Phh�� �k�q�'�S	�?�Ņ��&�0�&\4}q4�����N4�<чK�.T4D@`θ�b}��c�{���RۓA��-����H�vL�1?�m:$�] Tq�@a00O��3a��D��B�
�`��ʲ8�y2d��b�e�]�b��ӓ�N�^�~�[g"O걸hJ�~�mk� gc]��*�=�q���<h��TC�&���э�n#��v�A���w�F��2�2yG��x6��j��H��'�м��ȉ:\L�o�� ��D`4�ˉa��%i%�Q"3:R�k@J�A-��X��X�U61
��?9:��Er�G5(%�@�Y�f=
�����#MQz �?i����rxrB��<�@G'+: �ai�<�Ly�sFů/���ba�`��+�O��>kL̚2�Q?��=ѷ-��y��Y��m���yZ���>�� �	�k����y�s��d�iۀ�D v��s��_�c��^���'%ѝr4�x���F�<a�ED�D���(��;`)bV��B?ᶇ�k���a��2B,�B�U�oy\��&h���*l#t7m�� ��r ɇW��I�L4��¨@��D��\�>9�ݰ6�(c:(x���Z�¡��#�My�������ɜO��;�	�%�����!܀H�H�<���D�N�"~J�� �c>����/<iT����\�d

8+�#I��	�"m|�q�+U���5�ʎf?^B䉰-��=���MK�@���3�*B�Iu�<�QwƠ����2Ʌie:B�ɇI\~�*��D MUV��䃝V�C�	�	h���/@a����8dP�C�	�~{��:�Љ>>ѹ��^�4�p��$��y��!2H�7V,�A�#E-f��z�fI���xb �� 8� K�"��p
���O&�XW���[8�>ݸ��V�72�{#;2xl�P�%D���Go^��;U�T�ND�������׬(yg��f�>E�4�@/U-�Z7fR4L��F �y��U*
.�*�۟QZ���2"���=��CUe�)F�axl"!��	���_�N�Ā�h��p?	 �ײ����2�ݡ��HŊU#u.rPQA��/�C�	.g���2CA��r4p����Z혢>aVLʼ/<,bpj'擢:UR���(�KdYՆ�W$�C�I*s
�r5�2V�c�e�b]��	+C����h޲/��S�O%��;��ܹI�P5��@�	�:̈́�Hq4�"FNW� ��yǈ�;��x�O&�sΐ	r�q�
�HV�����2X�&)�Q���$H�4��I�ƈx�JO�6/�����&=�	�C&�C��)�@��E�+��A�Ęx� ����O��Y� ��0��>1���#+�8�kج8�My�l"D��P�ܙ;�h�V�D���DK3o�<9���4➢|� `�@�EI�M
���2��joL�B�"On���&0zT�8�)*+�q�"O~�j�ރ.�8 �0��O���Y�"O���a@ݬpz�y"��Y�%p!"O�-���1_ʕȲi�HI�` "O�1@��]�T��iD=un؀�"O��知&�B�+2���LG�((�"O���w%R�r]0���ۄS醰�"O�ѣ(��3e�y6�����"Ona�`��f�\9ԧ��h�As"O�	��
[P��7��(�r�6"Ox��
3�(��d_"�2���"OR�+2�в."�X1G"�L8f��w"O�I#�]�=�8c5KB3A.X��"O�Pg����Ѡ�+݄(�d��"O��$�X�~0��ϓ�9�t9�"Op@���+��"R��#�T;"O	�� rA��+�O�ru4,[�"O� #C�K�M����1+U$`o���'�y����l�h�����**ze��'������>Z�A�L�2 ���'edlp#'Ѩ" �X��b�$����'�|�ؗHǺ�r�������'�<h��ߕg@"4jr�B�ﴼ �''y+c۽Qa���|[z,R
�'{,1' F�}����o6c��x	�'pU���*�����C�P����	�'�b�� �>�����,G�J����	�'�d�rU�I�G��xH�a��T�X�:	�'p�]�j��j��T�qE�{*���'`*����	T��A�W(֨p�����'|�r'�#� ��fZ�>vh���yR��9yv���!F�'x|�Ir�Ë��'�|]����!d�X!Эܟ��B�'6�@���
�L1W�OO2xy�'�:M�ՅT%��t��G�{|�
�'�r�p��]q�(V%\�!(  �L���'B�*ç��q��-N@�����s<���qm����DV�z[e����0|JGA�>z]���OԐ7x�U��E2t�$��o�F	q��%{�X ��ӷi��i��I�`�$�P�T��74 L�5a��`���
w>y㇩Gl���BBN�8���jϧ0|�r�f�(&p�?O��𩉑R�J0卍�pF��U	�|�!����S����'at@��'K�B�kU#Źq>�1JB��,⾈�T�=V4P�Y�y�'M1�,�r�I�$$Lp�kB~���>��L��&���ç1�Zi�c�-�e:E�S�s��'�N C��T�OH�A�OQ>A9 E7��I"lQm�DHT��Ovt�L�$���N�"~ґ� Hl�bt�Ӫ:�n4��� �~�@V#{��O�>)p��͞	N �̏�SŜ���"0D��U
��W��DJdk&o|Z�0�),D���a��s88��,� 2�T���,��9�O΍Jt#�uX48#�Or�(Y"Oh1� ǒ�c����P��`<�\C�"O��!ѧ8�r� [$)��"O�,Y��#��0x�.��)�c"O�yؖ�V����I6/͙X�P4;c"O�qy���$	��1z�oU�$}�9p�"OD���(4�QA� s�慲%"OI"I�b�6գ�FA�2Y$T�""O���R� ?�i9��UL0@�"O��9j��(@�\3�钾�Vh"�"O���J�=@�@�*��H��!;�"O"���,:�H#�ְ~:��"O��كa�/]���k\�T�I�c"O@��#Ƨe��+$G�l)7"O�dÖ2R���
�K;*�\4�0"O� ��h�f�	w��5*,���SQ"O��ТmV���� �4+N���'��`�U˘!�HEK�*��V�0��'b*�QC�ؓI��J �]99���+	�'f�qI1/Ūo�^d��'��*��H�'dr���˃2�v�QG��� p���	�'�,�{���~M�V ͉�hH	�'�Ԡ"��_�6=����^�p��'����.�2��qa�R���b�'r�-Õ떖���a�gT�{�x
�'����a(:�ШA)�!E5�h�'����AJ�%\����B�x��'�2�qB�D81���W� .��i�
�'�8R7`��|:ta���B'6��
�'�.�KNw�Υ��R����	�'_�MeO^��
��4�Љl͈	�'=8��'�s�,,��jû	1��	�'S��1��S4P r�h4�H���E�<ya+ʯF�xؑ �Y�	 ��A�<�!�̋|h�"	K�vl9֌�a�<A�cѪD B��t�<X#�	S�<���
^2$e!f��SA��)$i�R�<A$b�1}�p�Y$��=k��	ɐ�
K�<�7���R��$��=B<���jn�<q�틧W��+��F�����֣�j�<ys�z�(���4�]�Cg�<���U�uHb��F@��T �)�Yz�<a S��j=�T`E&jBz��&)Zy�<Ia��LU�U�A	r2yy�B@~�<����,�t,Y1倠Ip4ab��`�<�#K�r<9�4#�����x��B�<��m�!d��%�����-�<�@���A�<�d2&���Rd֋P��Ի`�KB�<A��T 0�L��'� ��$�E&�A�<!E� �C$,JJ�Z�XԈ.s�<�D�$��<cS��(G���!O�k�<�s�;�R,���X��P;'Jq�<yaEЧ!'� Q�៮#4F�q݌�y�f��dln��ۡU�>%�5G��y��8(��"�(H��@�� ��y��IԔH���/���4��.�y��O3{���b��V����œ��yB(�4M��T�-�Q�$&��y���y� X�4�	
Of���I�1�yB' $p�qqv� �FĐ��$����y�BK�u��!���&D�r��4�G��yrL	�%A	��Ά��<ei#d��y�-�Ȕ�A^)1g�c�@T:�y2oIB�e�E��&��(�;�yr��??�:�`�G��ʝ�t�6�y��A<,��(w�ψaݸ	r�Ǘ��y�+F���u�^RൃƬ�y�Í2�H�!�ō�X��e��U��y�Ƈ��t���M�N��i���;�yҥ^(>���6�ƩE���2��ʙ�y�ˋ�.mx�a@�=� �`�M�y�HN/Q�܍򔫛5��!���y��Ȃ ���R��۪.Vr�J!H>�y��ެ_Gt��`�'tܹY�X#�y2A_�g����-W��P���_��y�Cϭw�DӞO�x��$.�y�/�4�P�1�/M�6�уSJ��y�%�f���S@�5�~�p㮁
�y��+lk�}�@�1x���G%�y
� lԣ�f�(I�AӥDG	=I��y�"O<�*у�I�RՀ"Wg�B<�"OmѤ%�c���� �$�,�q"O��dd�!u]T��� S�" �sE"O��؆�j<P:��CF�:�R2"Oqg��-����S;)5�1
�"Ox�B���A()���>C�lj"O}	0dHi/vY�m�73X���"O�)b7㊄��y�D��i"O2L#2B��`j�KWP��e:'*Or�7T	A��)r���B��\��'g�������d�$9d&���'�.i��B�2�H��[�5%�8��'�p$ٖ��Sw��k�名.�*�Z�'dH �I�-J��ٴ�hh��'��xX�,�6x{U&�r�d �'�����Fڷ"ۮ���d�'xj$��'�j�0!�Y�`����	K"oݲ|��'�hpQ4g��x��9z�g�b�H���'��(e'��5�N�P�T�٫�'-�!���< �z�����)N�j�0�'��a�I��_�n��G�څ�حr�'v��Ko_*'��h��(� cz��[
�'�ެ[��؛b�J�	@�l�:��
�'��3��J�H!�D��f�p9��--��e�I�b���y�M��k��Y�ȓ/���(Y3V�҉�@ �1l��Ʉȓj��7�]�L^FX��*-l�<���	�zse�sO�m��F��@H\��*�#0N���@� �) 2L��ȓ=H��)�㚏i
�1�k+��X�ȓI@��b�X�m2�J�A$f��ȓ(V��j��BO7�a�i��;G���W�>4zՏ�yt����B ]��	�ȓ|�Ja�4�R�a����U*�L��{U�9�B�S�EH
,�ք�"|��Q��\�n�a%���G3Ry��g�(��ȓi��D:`+�{�t�!@+���B����ii�N>�x谤�>h]�B�>� �!�,�0~w��9t���?z.B�Ƀe"ةQ!cG+\�h�g�&d�2B�	!Fn�2����ZI����^�"B�I� ��S�o�'q{�=sqnԧ6ưC�I)O���2�F�(d�����P�S�xC�	��k��[8��dZ֥�$0vC�
"٠Ĺ!�9���Kf�ק-:C�ɍ
C(�xbh��{^T�3�c�RsC�<!��8���9o�D��U�Q @�C�I�Hb�@���)d���j�	>��B�2^T�}�o�	�ƫD��zB�I�9���+�+��7�ޘQ�� -{n�C�I�#nĔaT�޲���2Ѝ��F��C䉢&�ta�D�\���]--JB�4��	3F�=J��$)��M�C��%P!�\���}$��H�$��(��C�I�}Ռћ,��!Q|�C�?msJB�ɑ6����29�PX��	KR*B䉑<UT�ի��9�(S��L�0<�C�	f���3��<Ϛ1�.�C�I�-�x��qbߖM����Dd�lIa"ODcg��%z�(�����AO��y�#�5f�u�� Z +�U�2
��yfӪ�����FK�x�x�81���y�#�9<fT�H�G.wZ=kʖ2�y
� 㕥̯[�D�ьPb�I"O�� ��^�_1�[�( 6��:1"OҜ27B
u̓���=)�@��"OhT4o��>\l%i���o�
��T"O"�&�\�<�DHA��4���q�"O����c���p���%=�ֈ��"O��'�m��tǅ�4XH�"O�pѪ�>0�5�QF̝Vx.P�3"O�x;vC�<��D�0w@��f"Oȸ(Mɤ!Rb�Q�FŉE<	�"O�u@����dAhkP��x�"Oh�{�b���X ��BI����"O����Cp��X����'H8V)	"O�)���!� ����l1��SU"O %)C�-n��PE> &�y�"O8l���^ l��� �h�*��Ђ�"O�i3t�>I���1��*,�J	�'�+1iZ/A
� �æp���`�'��@��dӧ>=`�ʧ+X�~ɣ�'ن5����;�)T#�Y��'� ���U��=�@!���� �'}��k�G�20�BS�Ł^�*�'��� �ei���3���	z�s�'�E���<n.�҅��6{:=��#܂D���.i�@��
�)&@@��ȓ^��q�e��f�4���@st��ȓB9���S#��`�:��J�KJh-��Az�����0���d� �ȓ=��@����<H�獁�P� T������������V!WN;f݄ȓ\T�2� v�x :$D��1��,��,�*���t���Uͭ}-���vx��U�M�5����	U�g����ȓ,3��.�99G���$�x�� ş@�<9EA���pXV�*Q2XW`~�<9 j�;�b�3Θ��x�[�c�t�<�'��:=f�*�%F0uY.�C��F�<�*�)<��Q��-
4�8xD�B�<I�hU
[�\@�AY�f2hPi�dK@�<��~� ����W�
��rϋ@�<aR�ԿjT��Cև}ºm)A�He�<�c�¦*Y�����i��)��,j�<�0�
pHr� �/@��4+^�<�+Q'|�\ 0�I�D:z�+��V�<�q�X�]�d$�J��HP�#Ff
V�<�6�jo����M��k��Z�<ᶋޫ��)�N�'q��D{�j�z�<Ƅ�F�@A)%_%4[�#���x�<�b�Ό	�T׏��Z8�t-Xw�<9�M��1Y,jᔄ�Rp�<!f�8^���J��	 �����Vl�<Y��AS���Ǧck��M�d�<y�#�N:���-´e��y[���U�<�P��Jv0@C"��	E�%3w˒O�<���C#�T9�6S�h��)�ĥMH�<�V��p�lxW�5�t$��F�<Iu�6�(��"B�'���c�[�<�e��o�&\)v�� ��}I��	Z�<!�_�Nj��V�
�"�e��&V�<1���H�Z@A�Z�.�B�O�<���ս8]��ȕ@S�Kᄄ{��M�<i�    �