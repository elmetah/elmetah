MPQ    �g    h�  h                                                                                 ��N=;K����+�0�D�E���u}q��䌯�u�ۥ����sM�=�rk�F�?FU*�$���u3�2Čk���7]˺塚NрQ�d��������.�-��h���G� |�uN��u�UD�Ѷ�#��!G�wL[bJ�i��I���ƍ��/�@̂zg)��yMm���`�óI���ߨo+�=9
�i�ȶH�4�����U��񥿅 +�"~$qO?�!w?��H�w���.�>ɥ�5�&U��:�ܟ�~�\C�+��&am3ul�P��]����'�5��7��kO�CX��5�sN捶%��!�����nE2Q�Xb�DTʯ��۱&�혆�F���ď�2h]J��y��ZL��A1��5 DӴ��Xr��7���89�M��'��iz��v�PJe.+r��<A��(���0��,�!���8y"~�q�Ǔ��4fX'�"�5�Q�����k���?:������L�{�ׇ�ٰ���U]��G����RN��5��=�Kq[m$��h��K(��:-��s�>'Q_ŘI���kq��>�k��j�R)����OS �eaW���*��p�\�_;�Ƚ@�q5����]z�* ϥf"�V63��ck}=���e���>�LK�~�)�A!�4�CLz��� �[��{'�֚�WOO�9��1�b�CH�;�7ɿ��d�aOA�<����V>�(��=,�=Cc?,���-�!ѽ�uo#�/7�٦��q�/T����#�Te�ٰiwe�/���C����r ��_��mڹ���NU�#�x�{ah�k�]?���8Q�}.|Ȑ�
����E����E��ѥx����?Fi�U1���d�O���+C:�ET�|��[�V������E3��@�u_ٟ�Ep��g���B�J�#�F*�U��h��d��*�.Ec���U���B�����Z^�Ӊ��('���ߤ.@����T:��С�Կ��M�^����97	��XK�%~�u�KB��k�DC�-�W@�S�<J���X�����
أ
Sv�S�2o�aj��AYE�&�*����,�kҨ� �P(�����m@���b���:�MU��k��k�J�%Y�\a����>8at��Y��;{
�%NA.�
��9PS���h���Oq|����N�O|%o��m��E�bs�hY:�r[vW��%�CK1�{X���!��DX�����[�I9�P�1�ǸSjK&���⨍;�K���hegB�LIIka�Y�cX���G�*���.@`e����i�N|���\��*Sn<���uZ�0=~�f=3��f�	�n�+(������������g�f��?�V!�k�ɪ�0'I�S}g0?���_�4"��q%&���Ք(	���+����K�$ٟ�� �PD���y����C��֊+#����\_-�~�����ŌA�L����Wa9U�7�͟�oS/�¨"��ݚҭd�
˓�����e�xx �MtLk��ݏ�w=�F��e�Y�Jej;��o~�7��9�'Q���!�d�fP�
bT�-��-���K��Gz|������o�<yN�fL���2�=�:�P$��L�}ѻ�?��7�D�o��ކ�uvB|J<qˢ�ӧ����ש�"Q<I�J��Q�����|}�5N���r��7�_�*].o{A�޳���-�(0�$R�]�q��i|ɳ�ä�^FP�,PI/�:�?��� ��-�������>ݺb�U�B��6�J������5�PS$"�S�O�~v� DO���ZfkǿINdxA�G�c��!6�S4��!��X��W�wU��Y�ڨ�p;�h�̷W�j��cr�-���"�`B^����+s}c�.f����_f0�wU4C9�!�_���;A�P6��n#*��S���POқ1����]@F��/ՙj��GK�q�e'�G�6^J���L(j;�靈j����լx��������S���S������g�ъj�o~g�'�A	�z���鷨ӽ�e�#��������+fc�Nǽ�/�����=R�u�E���}��Z�4���lͥɫԙ��N����z8R����G}������䝦thcO��2��nv=��͵� �W� �]V�/E������g�7�M�֥`�5\l��˾K;�1o.��6�9<��Y�"R�zs������L׬����L ,��F�9��DYW��ޑ�/jy#���g���Tm�ҋ
��� �x%ӵ8yW4#�=�P�ځ�"�ysܼ���n��*"yY.�����co�&��$��Z�𢡊���'�se�A�&`Z�	:�!hrEu�cļ�n����z�c��r�{��HYӀ�Q���s=PF��,���1ʢ�ϩ������iSsh���Kx�޿g��� oB=����?l�2#��n��;bP;8U�s�U��,��讌��E%S��1� �)[�{KzGg�?%�+X�	nf4���J_�2�A�.��w|P�:�?@�`�����^Է���
u!�F3sF�b��[ڿKb��e�׼wЯ+6�	����F�#������T��h�����W+7����K`�O�>(b�n��uʈo����5t����f͒���'#�_��И^���N����၆g�b���whb�^���U��͢fW�����	c��/�/ =� �fM�����g���0]/�d&���;ø E�u�#]�kp���l-nۡ<ڹv|���dU��{�D��b�Ð��K�/Uh���H�V�\�2��}��%����JE?KRh���G�	[3}
Ń������5@�QH.�YD���cܜ�s��>��9�~2ut:�>�iM'�0����T���a4�r�
�ş'c��<Nu�,P�w�j}���A�UR�'s6W�����8S �T�q�-�wix��a*��0��V(�/P�A���ژ7��eyu��d��!�wuj�սd?MVf�ŪB�~�~kr�-�ȲK����O������
��`c��GA���9�4=[�z].&����폒�)9no�oQmd�����`�}�O�E�Ϊ%I^O�'ӴA$V(���2�#�=�[�Q�b=�С���i!;ٱ3��3��3~a{,����G��d���"G73�)�Er�
�8�m�')6{��k�|���8��\�.�O�YX�.k3�N���j�-�������E��:�9�1��9{9��`ɬ�Eg߁�q�O�n���M����]��ոk w����#in��2���mӑ��q�mL:h���D|H��R[��RO��t��n�OrcfT��;�?FZ���<��>Vl.!��jN��� 51!�����OLlm����ގ��14���e��6BE�X]TcT%�ÖpJ�/"��i���Mi�mhJ<�`y�m]�ʔ��zh�P��DNY��3�ٯru�b��H�'jz_�~�k�Le�o���V��0��,Df���7�y=իq��`�yT�f��t"�	Q��"�+k
�N*���Qv$J�Vօ��%嚓d]�`1���R	%��P�=)�[�L;��C���jA��Ck	�s�?;Qz�,Ii�kL_�>�Q���)�VvǪ����_ar����Wp��1_v�H���5�+׸%*���f=��в3m��k�9����`��ܙ�jK� �)��-!I1$C'$��y��u��=��1�pW
|�9�����H�r7�V�$��\�L��bu�y>2���@�����C�\
� �ϸ)���o�#�rt�0O�
�+�4}��٫;�w�\�/tN����� �j���muT9��<��~���6��/$3�ز|㊹��Dn}Ɂ���Õ�cE�����`2:� غ���z�U������OW�>�N�`��|e�F�1��7�E�`(�;�n_mò ���3��x�%˜�pUze�h�=dV����ɻ�����d���5����Z�4S��ܞ'�%�_>����T���|���S�/{���:V7d=����S�@p�u �ܓ�P����-3��@��=<������"�������Lvߴ2
�Ga�)��^��O�ҳ�,7��;������;�m;4c�.b�0۞Ui8MМ*ks����>�\n��\t�E�a�YY �4{�4KN|چ
#MY9K�g�K���k2Iq�+�m��*�OoA�+�:.E��/�i�:�O�vrd}%��C&x{�v�ݼ���?�q�Z`�[t�9�10
�S���&���CL�S��peg��MId����jlX���G���[8��x�Yx�lN�� �G5�5S�!�����+�k��c�3���(	H�+�A�OpG�l�,��S���x�?��B!9��D,0�d��X}Q���ʇ�����i�*&��s�����v+���f�h��M�0�����[�g�n���:1���O��+_��'9,V�_���Jk����{�U���͚$�o�cy�c�z��Qέߙ}�n���EeG�_x$/t��
�\(I������+.�@Im�Cz�j��Q�j�s7W�r��&����d<�f��0�h�)-��F�:G�1�eu��5EQ���^�A7��y�=0HqPWoL&^Q��+b�'N1��l��k�����'B�q�.�.�$ǔr���p<Ė��h���F�����}����Aro�Q�z2�]��{���PW!|�(+	�$�Qn��q�>Yi�p���;�^W��`��I*�o���N�D��<STᏐ�.�,��U�U�˥�:��J��ˆǱ:5�uS����H��} ?���;=Dk��IiIXA7Лcق�6��T���!����d�w]8Y٪���Hh�AW	H����-z1h�y�"���^[�oǺ+�`�c�׃�~x�ZJ]�Ҹ�C�ۙ!_"z;8���	_%�	I���	O�+f1�R�ċ�$@!̲/Y�&�FV�������+�6y���f�R�0;"Lm�#|��~	u�q\n��������g���0[�j�хzio�v"'���	�̚�3s������eh���� ���ދ½f���Ȥx=xu4�������-����ч���& �빰 ����z�]�	�G����t.���vt��!�n9T�p�=)X��<�Wf�ת}��JCD�n����r��C�MMj0`޼\�{a�y�u�LX�����������RDy9���Mߨ��g\��YL��a�!��!g���G��.�/ŵ �Rw����m~%ȋ�V�;�`%n��8��4~'� =��jy����w�QnR+]*���Y)���Z�QA�A�$[��6|�7���-ue�?U,�vZ�r(�<�-E���c��X������a^�h=[u{��Y��HQ^às��2F@c>f�1�6����Cu�in��" �x�'dgU$�śZ=��ߚ��2�n���Ƥ;I�s�����詶4���SG��1�L:)�?�KU������ 	i[�#t}_=RfA�E����Pj��?{��|��?���
0�FNu���'j6�8K��� �������Һ�+��	��gVג#�mg��0*�Wkg��9Jm�7?p'�#��ʨH(=�T���ue�2�̏�_��Z�������`�##gB�A��Y���������4A��!��R	`Ι<6������YxWy>Ig��$�U���� �2��-tMV���ę0g~���IB����E�Ó���c]��
p�?0l�Z/�\������m����P(�ub�H푄c{/�q�Z���qf�\�=�����{�%O���-\?��[�U2��$� }�����	��F�5��!H)65Doӳ���D$�0�p�F~ms�::�iH�b��>�t@R���4�\h��k�b��Om~u�p�=;�jǫj��G�U�J�sP����4� �c[^����N�i��va�#��D�VcΧ뽘A���5�ϗ�R y#Q�z~��pJw��}�XֹM�.��	�BAN^~�9-s�K\�ナ'�����`:�T�}c�YA�<9M*J[�	.a�=��÷���o���Q���y;�`��|O���i]�%Ddǂ�Cñ�VC�u��#�8�[8���Z�Мñ�SZ�;�������3Y"g�7�d�.�� ���G�!)��Ҽ�+�8־x'd�u�����wDa�1�LnH.[M�����	 3��[�n/N�(&�Zv���ܑ���{�t�-�ɧ�8g:�,?Xj�ٔ��������`}]�%�ճ3Rw�U��2պl�<��l����m����P|i:K�_����G�t����Z���dr�p󡓙F?�w��m�L��_l����7d�5̖��ɏO���xR.ީ�bͫ�c�q8�Eh�jXXH�T�v^�QO�#��<�ܻ����&J��y�,�i-Ϸ��k'+D�e�����D�����C�'n3�z�j���e$*~�Jͻ?���|0�7�,�Z1�K�AyXLq1��T��f��Z"�.�Q���	5���N���1+d�+���5�+]�K��<j:Rĺ\�k6�=�7[�L��?&���g��6�~�sM`�Q��I�!k'
D>�W���z�)��P�t�cN�a��!� �/p\�_��\�v>�5�f���*v�fX��,�{3H�yk�U���*�[�W��zHKW�<)��b!�M�C�{2��ґ���3��� W��r9*�E�X;�H��J7?���73W�ԯ�_�0g�>Mp��Ӆ�Cٙ����	���+��#i��'. ��L@���oS
���K٦~�w��//<�m���0� �fb�H�m���JÇ�N���2EJ���SF�e�pǢ�}d���ۜz�j[����U�{��ћ�	��5�Ƶ�Ղ�2���O��r�@�{ i|�^�X�rbEi\��6C�_�U���F�N2 ��� ����U̔h�Wd�oeӤn����#���AF���Z�K���'Q�6�nJ�0�T0�"�W5k��ʷ��
7�j�����[��u��"��U˺c,-Ά2@{iX< �\��Dى=����+7��I�vY�42���aA����\ؙ�],�"横����t��2�qm69���bg��p<cMKӯkN�3��K��o�WjqWؕ� �5a�}Y�fZ{�� N��
��^9F�צ���&�q��T�sĀJo|�qͣ�.E�fH����:IL�v���%�C{�X��W�:��\C[:��9/�1�l}S˭�&p�ޖ��{l�]��g��rIH�O!XhE;G:���2V+���A�3�jN�N���-����S�"ݵ(+��&�5���3|��hl	��3+�9(��~�s����އ!D?R�!Tд���0� &�}�����̗���$��&��DՊ���~��+Bۍ.���7���-Ʒ�� \���9Y�!�� j�8�w�}V_�ʯ���0K͌7�KF$��͵�U&�͕١o	�V���)R�ZT|�I��(N�e��x��tJ8��&�����
1����~ʥjq=V�e�7�,����\hd��H��]ϣB�-�B��A�vG0Ϛ ���P��2�[�BW�U�y=�u/P8�L�^Q�q7b�B�2�:SǳFf+�8mB�[q��[��`�O	���<?�"�C�r��d�P�}��_.�r*0���']�{��H�������(&K�$���<sq߂dir8/�y�^�Jc���I%� �gxß	�l��k���ΐ:g�q���1U�������J<�!���H5�PGS�����X�� :u���?bk=;�I�N A�xDc�:M6(���K�!�TY�N�w�5�Y����f�har:WU�m��]�-uj���d="V�^76��c+�nMc�5ŵnc�UN��-<gC��3!1�6��J;��ƾ)ʤ�X�U�=āO���1���8@�/A/K8L�J�\A�4��L�w0�6�bs����%�;]6坾��yn���`�)�&�哀�Ij�B_��kPU���р��o4��'g�9	?윮(I�aeI��eT��j�ҡ���腽�(۲س�Hiu�
��mb�sE���tѢ=�ɡK��k#��ezn���<G3�Z�@0���Nt^p �I��N��=�f���W�b.�����ea��閐��-�pM��`��+\"���4�t�ga������5���RߗW���/:ڬ�"{��7�KL�����ȷ\���������/ �_���cXm��I����vD]%	8iD4ٮȣƒÁ4��yi��Rpn��*X�Y$,��H\�?��\�J$�`y�����r~�]�Ne�]h���ZO�z�W��E��c��d��]8�1ƽY�K�c�{`�FY	w�Qٱus���FS�-��1��A�_���ai�?���9zxz��g����6f.=��5��`2�06n�f�1KE;�\xsZT��b�� )�^8@SM,1�?)QmK0��!Tr�a��	dp�~(�_���A�|[�m�PE�?��ݝb��E�l�
�DFi���X����KؿX��f���B�-ŋ+�s�	˔�ч#�-Y���S����U���37�P����E�>(P
�[9u ���]��뿞�D�K���͈��;�#^8����Y�T�l��^�;�C�X���-������V��0�W����?�e�%f� �M��M�c�ſ;�gr_X��V9��N[��*��n.y��U�]%�}p��
l�fW�L)��zܱ�)�Ӹ妺r\b,���/�!��Ɍ�j\�����W�G%����0/?����B�?�} �;��!<Ӂ��5vl�H$�Dʫ���-����n���{�K�e~���:��iC-�J�i�/ԡ�5�4��i��}���>����u����mj����m�UH4s�h��Ϗ� ��c�͋�(Si��Aa X���^V����lA~�ߐ�G�Q�y>M���Έ�ߥw��F��g�M�s�6neB�=�~� �-�=�K7�A��|��/������cu�A��9�?[���.�~V�>u�%��ߍ_o{��Q��y����`�=QOA�]�0�%?����}2~BWV^�6�i�#�S�[s.���kЗ��̮j!;O�3О6x�D34�X�|G��3.�ُ6 �G�`5)"[��l�8�/'�.$��3�r�㟌�����.#ē�OQ���&�3)]��	���#x����1�S��0Q�/���Y`ޯ�@�ȸKɢڧg��,��͔	D�M��+]>zծ wC=�ʙ���N����G����[m��O���|�L	���]���X��"��r��j���?����(���Pl$)��/A�r2L5g,\��O�3���į �'��������E��XS\�T�	��N~�>�љ�|C�d�,�㴙Jrt�y��k'��rn����DD��m���3��\Y�>I�'�"zվ:����e�Y��%9��z���R�0��,,�n��W�ys��q��7�/Ȧf	�T"S��Q~N������_���l�I��r�f���Т�]�V9����Rpm���=L[�lY�PZ��Pf�\!�s��Q�mI_}�k�>7~��;h�)�x'�`4��a�	~��Gp7^�_�-��45���nܵ*1sFfs���p3#�k.��͵�	�V�O��Kĝ)���!?�C�}�mB��,���!ß���W�59E�����2Hj@�7zV��Z�#RVدM�\�^�>h_.�6U���SC��V�۸9!��~?#$XB)�&j��Z�˪%T:١�iwv�//�Ib�2%��� �ު��m����xć4<�ڬ�Iedz�����@ߴ!�}��h�֕[��s��=�XٖH��d�u����&�1��PSOG\�c閆[|[b�������CExL�1�_#�I�vQW�i�8�n2�������U�R�h��%d	��_3��Jɩ-˝G�>-�Z/�����'��i�ս��K$T����2�οS��eG���c7�\�H���v��uL�~zH��#�-iNP@v$/<[�
���J�X�)�옣�0v�U2@+
a�4�R�Q�WMř��,.Ҩ��K���V)m1��|�b"ޞ�/�M�)Ak)��,,*x+R�o�sW���*a��Y�{���N�R
Y�9A��\��5�q͝c`���o����>ׇE�����:i�v��.%~J�C�E�{	[_��g��5o&�y�[��?9:ν1&�S�i&X}n�yK5}�ï���gs�I������XCµGuS��-?Q>_�.���B�N��+�=F���;SF�õ�!w��w~A37VV�Ȫ	>9>+��Ŭ5��h�����w�.?rF!o_��:V/0�@;_}8�s��,�E�8��-!&�>����Y+=�ߍ��I�6^������;}��]~,��5�;�ɒ�����_>��T�KWm��I�!���'U���͐�$od,4�����. ^��.�$�vc��e}��xD�t]���(�ȃ���V����$��:�j��`_N7���X2]�0)}d2X������޽�-R%P�<)�G���ۖ��k�̅�KD��lWېe=f��P9sL�~ѻ,c�]t<��Y�!<*�?�FBMq����)=�
��m.<�Ѹt맼 ?�è}�����r�DҮ�]��7{�����4�Wy((!�$ct���	�q���i��T�l^�����1I �M��D���6���9J&F���p)݋0�U��A���J�c����5u��S�H��+�O� 58���a�k���I�spA-A�c�[6cm���<�!�⣿�ߩw�. Y����jh<��W���4�-pÀ�/�"�C^R1�ed+���cJ�{�Pf�PrԈ�pCj�q!L�6uUG;ү����?6���0����OP?G1ըā��@׳�/�7{���k<� �v���2Ux6�z�\���T�;�@Q�Y��t�'�'��2�� ;����D9]�e٢�=��{��o��R'"�	!��)�tz���me�:����ŕg�\W/f�\1#ۍ�s�uj����S�����eM�ѽ�v����oF��TTz	�Ω�T�G��E��4�57/t�&��$%G߉�=_ϴ���W^%��*�怟b�d����P��K��M���`�*�\}�����7�����|4%��oE�
r�Rz�́��m�+������R��L��.������(*)��Ȉ/{���fb��b�mt�W����ñ�m%���8%44V���%n�O��y���-M�n���*��Y����.��\��w��$Qٺ��&������ e��W��Z
�1�rH]E�_�c�����:��T�*�u{Y$"QT�Vs�v�F�R�t�1���ϺA���ҏi����SxU�g�LE�ёx=�%��P��2Tz)n��O��1;ɐ�s�f��!��jy��S�!?1�)���K�\����	_�ħ���_��|A�Ӕ��WP x�?�:��������
���F�َ��O��K�X�6>���A���Y+g�|	���LXV#���1�Ѳ���
�  ��7�Q4���� (��/Bu�1��"�F@���QQ�r�a��-#�)ąwØO ��_M����l��dE��k���&�o��'PW/������Z����bD ����T�M�R5ź�g�`Ӻa�����;r�Ie��&h�]�ip�9al>���W��)��c� ӓ������bǱn�z�)/f���4nɧz�\��Rذ�ǒ�+%��*��S�?\y�˭&�Z��}{�I��YӼ�45KH�D%Y����F��������&��~��Y:p�i>���Y���١���4x�w��f�؇��.'u�XG�!�j=i���U�=�sǡ��Z4jk% ��7��^"�i�Ua��2���V�l!+�A
����D��<�yYi�p�&��n�w&IՎM�4��BB�Mv~�'7-(K֯� ��������m�
�c0oA� n9Cuh[d��.�������ޠZ�:h8o6�Q����o`��uO|���"/%:�M�8��9�Vy}\k5�#e��[���3�Вű�	��;
��Q���3����E�ꏑ[�Gh'�)+��w�X8��i'�چ�����mr���kj���.>M"���P��b�3d���L�ꛤQ�{���x骟��@5��a��c��ɝ�g����nH��K+�ߋ�?��]��թ#�w�DH�T�%/ٵ2��"��"�Hmy׀���|��k��,���j1��|
 � c�r4湡���?W��㶘�?)l�+&���׭  5⭭�{�O]����Y7�ߺ��6������
6E�qXN�hT6�q��l��Y��26ֻ?����J �y}
����-����vD�%����#CB3S�9�'$&uz����e�:� x��т'�V0�A,U�A��[y��GqFu�
��fD�b"Qy���<)ӧ�r�.�A�tK��4���ڼ�k��]��W��^�R:F�0=�M-[{�`�������<�R�|ɱs��Q��YI���kݿi>r�v��uF)}9�ǻ��ha�l��p��_'A���5�^�����*��nf�JC"��3��Oki��Pg �QZܪ�DK���)+�!��C�i��������C��B`!W;9`���NjHEש7��ɕ���MCX��X��v�>�n@�G3��%COt��E��ϴ�5�#��P]����t�G���C�����ٜd�wѣ�/�wp��!H �vCKO�mF�
�ơ��IT�g���4��I�%�"i=��}�R9�Ѯ8� �E��8�ٱqё�����++����ﱸ4�Ohw��d�,v|����i!��3E��2�,��_~R��1�,�4����Ļ�6��2g)UK��h�+�dg� ���j����x�7�y�Z�	���K�'s�ߐ-e�f��T&��IB��sp ���
U7up��FƑu�᳓Y���0,-6&@q��<���D0 �s䏁��ƣs	v�@02�}/aB��.�^�#�[,~Y��`��<Ag�h�m,�5tobݣ%��B�MA��kT<�6.Š�M/��v�a���Y��){v��N-�F
��9<�+�\B+����q��lj��+�o�y���8E���z��:��7vÀ#%��xC��{D}"ݍ���0;�k��[�k�9U�f1��rS�q>&���� x+��F&g.b)I�S��EӎX_`G�KQ�RmLq̿�F�� 2N�Xm��~�r7SZ�Q�^`��u]��;3�O�H�	��4+��E� �ں=~1�NF��љ?�e!��T��$�0��v��}�r`��&����Gꚬ&c_Հ�0�4J�+xꗍ7�����AZ�<���V�����K��A�v(T�nZ����_�}`j���f�u�-���AQ�C�^U\~�͋�#o����I7�P)���l�8Ge��x|t�����M�ㅐ� �����Ȯ�ʶj�L��[�U7h��hs�KZd��q�v!��YO-�'ĥ7�G�m��W�ֆmf�('�ҷ����=1�PZ�L7�ѻ��x7N�0�O��1��zz�B��:q��}?���Ŗ&�8s<5�������{�}}�QX;�r��8�˝D]`�{�����'�(/�$�5��I��qk�ih'[�/�9^�F1�IB��1i��Ɂ-*y�xs�����M��&�(U��y�K�)J�f9�`]5�k�S��E�?�2��t  0��L�^k�6I���A�)�cj
�6�`�򁗒!��ʿM�wAG�Y*�l�\I�h�}Wˣ���S-k<ϊuh"�/L^mL����+{�]c��U�믁�K����C%T!g�^�p;���<�w���g��G��O�]1/Ɩ���D@�W�/�V~����7�h�Ѷ���6�����\�n�";�j���pX�o�;��ɥ�D�N�?�H�2���q�;��vjo�d'�[�	<�����LU����e9���
#M 0k�=�/e��q��hX�)�GuP���Y��)��� ����-7ɗBW�JA���s�z�|��%�G鐰����P�tT�������3=�W��氬Wwy��I� ��-�߹ҳk���(bM� `ϑ\��[˪Ҿ���"����åk%�E�R5�����ט�{�m�gLJ7Ȳ��ҍ���͍���/�*�����|m���v���>�%?�S8١4�ԣ<�<�j�ay_R͛J�n��*�7�Y2��� ���󑒖�$�qȠm�͏�l��e��"=��Z�lL��(�EC�c�O͛Z���g�^O�NԵ{�fUY?�Q��Csst;F��W1��1���t�bi��2��Yx0�qg��l��=��߫%'2��n��'�j;��Js���՘ؕ��%���Sx61��)GK�j��ڗ�	Z��4�_nqA�JV�c��P�!�?,j��M[��(�"��
a�.F�;��N���m�KN����5����1��9h+"T	n�Hj#a-�l£�(3��^[m�7pr�1l��;��(΅�ZH[u6�M�?H�������4�1�~�Q��#�:c�AD�Jl�����8n�����N6���y�J1���}��>W��gzL��u�]�� ��J�C�M'aŵߘg(�.������D�����$�m�a�_][��p��3l�ߧۍۈ���-��n'�n���0�Bbb���uk�/���狗m��4�\ֵ؋�g���C% L�ɖ	?�����N�u/}�&$�_�2��6�5���H �D�&�O��ߔ��v�h���~.9:Vi9�� R?���c�[4󗑰v����� ��u���NE�j��Ȧ"�U>g�s�����g� �P(o�)�<?i�j�a!����uV���AҴ�F�ؗ��*yt� �\�i-waӵ�)��M	�q�� Br}~�N-�2�K�/.�;�.�ey�	pq�e��c�)NA��9��y[?�,.���t��;���bQo��Q٘3��{`d}�O�2�:5�%56�Ǔ�0��V�ej� �#@�[�j!��s�Ѝ���d�!;�`D%Zn�3�v�"�5�u���֓G#I)F~��OI8gqj'���S5��h9��B��}cU.Y���E�����3��Q�?	�|��k"��x��"9�%�I�G��%D���ɘt�gK��]vc��K���r�k�z��]t��դK�w�k��U&����c��Gf]�im�x����|z�E�	��G���)G�W��;f=r�Pᡄs�?��������7�lo�u���.h5�����)O�Mâ����:��|�h��"$ZE9TXI��T���Â�B�t�!�������YݛJ��yx)�!x��Ჱ�ʈD:+w���S�^r��i'�4�N'O�zKH���tge�;���'��]�5x0��S,��ɛ|��y�q6q} ?�廘fA�"��$Qt.���:[�Ih7bz������*�2�]��1�M	�R�;[��ݹ=��[V������R���h7מs~�tQ�}�IU��k��$>�*��q��)x��v�sa��N���p�7_b��G��5�
I�$�*��;f������3�UCk�j���jo�L�1�cK��)+��!5c=C�uc�0��bp�������qW�n�9{�o��1DH ��7�Zؕ�dmHPT�Xa�->����,ZdKC�L���G���<k#���xs�vT�� ��[�?ٗw,��/`�� ��	ʻ [.,��m�� �4[��v;�"]�$b��������x}x}5�����{F���������?�`���f�ς\�ű�8_O���Ҭ	���|QU���".�#�E:Q�'P�_� Ѳ�$��偝d�������mFU�qh��~dN���)ct�";�S���Ze;�װO'bw��K�����T�k���ƿ�hk�-b��:�7�:�����Ƭx�u���4$[�k�-�=�@l�<k'������A�����NTv
L�2v�,a���:�͎˙>�,��n�;g:�wWl��m'��ϼ�b�_��uM�6�k߹�qOj`�-H�h
��1`a��Y��{Q��Nh��
�[�97֏׷H�W��q�HY�/���o-�;�t�AE�ܺ���:ziv�t�%ttC��{���([��+����<[kS�9pl�1T�S\�#&��h�s�F�nͦg�ԺI�����GX�;G룃��́G�����'d�Nw�3�=Mi�S��	��*�����-%3�G����	4`+o}�;i��سx�7t�-ڄ?�yZ!�U#�0c0d���15}ne���A�����UK�&0٨�����S+�n����_���8��4�qY�Sg���ֱ���	� ���_��%?����匨�t� �~$�U�_X͆��ou��O!��dn��C���hs��e�D�x��t���H������{�۬ܜ�/{jB��V�7����ν��f#�d(���Q���T-�J�2�SGAGL�Q8�֡e腣"ڣ�"����=��:P�gL�R��{��h��ƥ��G؆�K�B��vq��8� �ǀ�ԩS��<������2�l!k�}�(�p�r[(c��V�]�<�{�x �<�I���(��$E��q0�i�N�
��^C���vI��x=<�:F��H�@@�,�_v�K���YU��M���Jm���3�c5k)�SkӋz�m텄� +��=kn��I��A#2cE"g6�s �&!�^Ϳ_�w��YE+"�ל<h�Z�W�j�-fՉ��->"���^���[��+VX�c���ņ ��F*�>�dC�V�!�ޮk�;���w���u�C��D��N�lO��81J���w�<@��/��U��2~�,�����6����RܣI�;���6�j]ˬ�-.Z���6��i��L_������q�oE�'�ּ	WUќ	�0P��^�e���~�{���BaJ���R�}�C��d*5u�"T������T��N��������%\,���z?F!��/GD���q#J�k=t����ڐz����=� r��l�WҴ�X?�{!�Z�5�F����M���`��\3U��e
��<ԡr-�À�Ֆ��[R���2�K.N�SQN��'�L�!�ȍu'�0�^����/1��>�Ⱦ+��mj��Q���'��%��8��4�
���/����yڿ���f1n>L3*)��Y���Y3~�=�~����$G*��H�ޏ#h��.�e�w���Z�U˖�(-E�F�cd�)��h��'�J��<v{��"YZ�QJ==sN�^F����1����pHև/��i�a����x��gA���I�=�Ø��*2�m\n-J����;Xls�1�3��蕞.�o��S3+17=�)�=K������2`�	Uo���I_)�A���,qP��?go0����^�}��
��F����}����K����lM ��߼>��+�4p	| BYJ#<-���ɲõ�� wx�7+�kL�[��V�(�P��nu�����i����u��O��������#l����ݘE�e�����-9��'����7΅m�\A˹�uW�װ5.�E���� �Q��ʊ,MGŰ�sg��i��<w���U�1a���2����]�+�p���l�K��HӾ���"�YA��I|�k*�b��P�pI/��F���.\~���f�Z�\�%��%���?ީ�A��ΐ�}q�ʛ:)��2��5G��H.=D�ڳ
���D���=��ܧb~Y��:�Zi4�)[j�`r�2�-4n���Q���Nz���o0u��x��
j��0�=�<U���s}s���<��� �����w��u[i��Sa��	�w�VO��W�A ,"ߡW񗂥Vy��f<�D�Xw�}[���TM�*�G[�B-͞~�o-	]GKȩ��v<�� w��`���4c��AEt99@7[�.M_��l����|�o�t4Q��<�e}�`?M�O��}��g�%0�����?��V�m`a,S#dB[$AɽikЈG�̿[�;��!��u53��]S������`�Gr G�I)a\�m�e8BB'P�h���c ԟ����8��.t������u:3������L�.����b��=����7xn��`Fr��5�ɓ��g��%֌ה}0�Mc[��լ]8�՟�2wT����&�A#�(��������mS�����|�C��K�1�b\��`B��2:|�v��rj��Q�?-��Y(u�Rߓl����_Hv�#]$58�9�㭩OY�d�P�1d��\ϫC�D�]]EԴ�XDX�T��=
������(	�������!+JCw�ysh:|"ϣ�o����D�o�z������i���/!'ژ�z���re����U&�+f+]�0��!,lR�7��y�h�q�ڔ���f���"$�'Qo� ��G����g�dJ�ݟS������{塩x]�7����HR�Q8�ת9=�T[1�_�l���r���2��s9#}Q6�I�OLk��O>�#��)s��q5�O=a�����
p�a_��v��`�5���^k*b7�f�F*(X3���k��͆���Gh��`�AKC)Y)F�!��ACn���D����盟���W�;-9�]N�D�H�d�7+ە+^�C}̯^��e>����?��C�Ύ�'S����1#U�6�V����YQ��[�H��bVْ�w�Ȋ/3;B^���� 6e���m|9�����EĂ��U��4��?����"�[�}�}�@��|��n {���hчp��;-ơݠ������\O����R���#|��s�x���^s/EՊ��"?�_4ϴ���#��ߖλl+�E�U��kh��d�\ӐAԱD�a��.=���Z �ۉ�52'���m����T�����Y�~z6�S���7+���y؜��
/u�l���,˦$�-:e�@g<l啫��7�����톣)I�vEw|2�a��7�cY�����Y|�,t�B�������� m"=y*�bS;A���_M7�=k�?����g�Q�C��]����aP�Y���{,�XN�K
*/�920�o����q����@�q�Toh:��3�E��C�0p;:5~v��E%��Cmz�{�!�����&���!��[&[[9�kP1�6�S7�&	e�J)�n[r��tGg�gpI���;�X��EG&ꥈL�B7ۿ?˻<
N�H��OJ(�S�o��^���Ĉ�3h�n��	�#�+JE$�v���s	��@����?>�*!� ���!0?z���}	ԁ�ݮ��V6F�
�&Ko�vaM��;�+�%�mA��9��6g�3錠 ��oe1���f咤g���d�_O�����;��#�Z�ߨ��ީU�aó�ouI��
�K�Ų�F~�˵��eN��x�tn�/�~��>���Vۇ��jK�j�ۘ�Q`�7O�3lсPld�i��,�/Ϗ�-#�4�-� G����9�ּ}R�>������A�H=7l�P��L�R�]������&-��}���<LB��q���˒�;�&�n�t<+�丯�u�m����}����r�Q�0�]�8�{c޳w��(�o(�A$tk��/�qKӢi^�7���^~��gfLI<���i���6�ch��}r�:X�Sh��\�U�C��c J(��Nt5�FSF������� �� &A���[k)��I�qA�Z�c Ze6��򷬑!}L�����w���Y`���R�h�=�WA ����-a��@�"B��^���?}+1�c���!q �A��ԙ�NC��!�$'�F;c���O��iW��)����O���1eK���@h��/7� ��G�-���I�c�6 ���{�$�;IN�*���eB׬8��r�Q�;�5T�����Weޢq3��l��o��'Sq�	rGÜ�>5 5�eoq� �y��2ҍh`e�d��R��X��vu;ǈ��~�ߚN����pɍ��� ����zڣ���'xG���,_�� tJ
��vl�:V�=0�t��HHW-˪���=��\ų!����`�MT,/`ſ�\��� V���͡����[�U��7�RKRA�|�P����.���$L��h\'�H�������/����=��F �m�1ʋ,��b�%u��8�o4E`���F����yUM^����ny$�*��Y����e'��uN����$�H�#~?�^K��b'e�N�v�Z;^���HqE�ic?U���V�����Ey�Ŷ{LntYu�QūBs)�F?� E�31������Z����i�W��_�x�s�g|�>Ţԧ=����a��2��nH+��;Z�]sF�U�Υ��h��ʝ�S�_�1R	f)=�aK���}���4	P���9|_��=A*�q�Y�yP�թ?��ɝ�ԅ��z��=L
��F�_��Dc�}wgK�����"��.H��.E+�
�	7	[���#mA��D�^X���ln��7��g<�1�O(�;AдMul��ퟡ��W���0�zj~��tT�많�#J�]�H��@dF�p
J1�#{��D9�������<��$͹��VW@��/6��u� _=���M]��ū�g�$������ϥ�����"��^�]���p��MlO����������3��$Zy���yb����k�B/w�#�����j\�0��As}�C�%V���|�?m�ݒ��jΫټ}�=��i�m=�5��H|eD6!��Pu���l���A~�JT:A��i/�Q���S�Mb4��,u��#��V@�uۤ;�)jnu<�XF�U4�sX}��X;�� ���%�����;im?ajg�RW�V�Jn�.A������=�fy�}��;���tw�G��_�'M�`�?�B�<9~�W-��<K�C[�����9��oM���ca�)A'��9�ՠ[�75.�?��S��ѿ�K�Cog��Q���]�`=�O-�0�p��%+b	�IS�j�nVʕ>�W�#��J[_7��Ѓ����";;xe<+�d�3�$���N�k��ŏ�-G�;�)|Z�貮83|'��煉<e�^'G������2.��~�;�8�P��3�o�u�� ۤ!%2�[�X�_�F�S�Tޛh��4��Ɏ�=gy����K���)(U[���]��՚�pw�
ʅy"\�h���gӳa���Gm�׿��ޏ|0ւ����}���z��������r���zO�?h���y�m_%lV��:;h�^�T5��s��v&On�n��#�0���+.�9}㘶^Eo5�X?�jTG��������S��"���"��υnJ�b6yn���`j�^���,�D0���U}��0�U�*1O'5�z�Qd���e�W�����f����#0��k,f ۛ� y��qs�v��/�f�+"���Qj��M���J��LX�Y�x���R+)�<A�]~����Rk�Y��=��[,W�<w���������s���Q�IK+�kn@�>#W(��^*)n<[��uL
�aV@�! p�u_�2o�}9�5�� ��ɒ*�f������3�w:k���!ҵ�BEܻ*�K���)a��!+��CI�cY��Ҙ��zi��SD�Wl(V9��̿ H�[�7f�ѕ�w�>�����S�}�>�[��"�wo�C ������؄��#����]� N,΋ڪ�R%ٍ��w�
�/���V���z ���Ȓm�u�pb��1*ژnE�d�ź㬪&�Y6}kC{�¹��1��)Ď�����I�{�����幱���Oya�H�?�߶|G�g�S�W癇;Ep&6�N5_��X�bxE�է�Z�E�G��dWU��h�YHdx�J�K���_�������	���*�Z��+��ڐ'�5��<,���-T���О���?����ݕ���7��i�43~��;ub���M.��d2-լ�@bP�<�D�u����[s��-���v� 2�5�a������CPb�t&,��<&�����9�m�}0b7��;�M���k�偣����ڐ>6�!���Mha1��YΫ{:�Nރ[
�"�9-��m�&�ͼ7q9�OR��L�_o��<ͪ�\E� )���:�xv�r%jh�CH!&{��$�^�2�!�a�|*�[�9���19�S&D���])i#:�$<g_JIܶ[�X���Ga���#�=�|�����y\N9���)�"�	Sw�/ ��/��3�3#��#��	*�+%�;�������ić�J�?� !��ش&P�0x�'��}����آǗ��5���&f%�������b+)���h��rP�R�Um���A0�I�r@�F�'6�?j���_�yz�������Ǭ��<����U-���|B	o�=��� ���<߭�ثː��O��e�=Ix�Ftɦ�㾈��4L�q,��bfծ�;Wjx�5�LK�7y`�D�Nќ��dZ�������i-��0�(A�G�+��Yb�׵���y �cX��|�=�9pP}LLH@ӻR ��@����v���Ɔ+NvB�67q�P��������1<��C�������jW�J}�6�&�7rы�)�]yU{>����<��7(u$�9q�z|}qf��i��ǋ�dA^�C��I���.�⟰�s�~7h60D�Z�������U����\ڛJ�.�i.i5atS!<~����� !�r�]+�k��IHA��c���6O���Rg�!xZg�U�wrQ�Y{+E�ͣ�h�@�W|^���ٍ-\g�ϛ�i"��~^�]QQb+�/c6o\żd�<B�����CVT�!���a;�;>S���3ʫd�����O<�:1�Y�m�@C;/rt��Q�(�h�����(j6O��H;U�O�;����ŅY�`G_��V?�1�l�^�������p	�gzo�r5',	�Y]����9�pSe
M���*1���H�����H�����`u�'��+,�:���QХ�)����T���b�@6�zu!T��X�G�!���p��t�@�|��u�=˱���D�W��B�zi��׀�Pހ��S&�7-+M�
`��/\������n�h�7�6���?R��w6��o��*���/L}0��Cc��������|i/����?�a�/m`��̤Ý�x%&8���4�3֣m����iAy����� Bn�W*_�1Y�Q����b��5$=��������N��d�9e�ӭN��Z����ވ�Ex�3c3�e��8�@�_mw{"JY�Q@:Ts.UFz���	�1�Nl�&����in��9rx�|�g���=��=��\߼�r2@�nc,����;5�s� N�i���RT�%��S��s1m�s)��,Kw?FH7��hCA	K�N�E��_���AEp��ԁP���?��v����>��3��
�l�F�!!��h*X,K�a������ym���+S t	R�}8�n#����t��X���@l��7��f�Բ��m�(_F'�u("횂����K��������:��D�#�.���X�;C��:���>�ٿj��tn���E'��(��C�W�d��Q*��2�� :I��@yM�L�ŦE>g9���Mvj�!c��'Сõ�e��O],��p���l��!۾"7�3&��OF�������D3b3��f��/ҫt�D�#N\t������~��%�� ��T?��Q��$_���:}g�{��x}Ө�f5}��H�iD�N���)M�0|��7��M�~��:�E�i*
v���ֶ�h=�4d�'�������0�u֨_o�j)d�spU��Vs3Ŵ�FŇ�� ]�0U�JI�i5sa�>�-��V�)����A�?�W���Zy�&\[����w2���sM�x��C�B���~(��-��K~�	����6�~���%�v��c�AB	9/��[М.�?
�E[I��Y��o"��Q*P��[^f`�L)Oh�7�-�%&( Ǥ�~%�.V��W��#ѹ�[�Mu�����~I��u��;�3<W^L߂3{����B�_��HG���GT�5)�x_�c�#8�C�'���$���YN��S�9�xG.��-ݶ���+�p3P1��ݨ
�R�|V��.��s�'閽X.��֪��(OɉKg\h��͓+��s�Agk�+P�]E�Օ�Kw
�5�@�w�����ӎ�Jm�7(��1|�������ɘ��V������/r�Ph�umW?������و��l��S�N�י�5n����_�O����z�K'ύ�����E��/?E
֞X:�NT��ó'8���ƙ\ڻ����

fJynyiF�2����5��oD�X6�0������mq�%{�'���z|��(��e'Ńl��z��z�0��1,��c��U�y��3q���v��f0�d"Z�Qen�����k퉚n	�J�SȌ���
����]ym)�^��R&ݾ���=�O�[�랓w¶�#��j��ޙs�ĺQ7�I�&xkI��>^��B�)i}�'�w���a/9��hAp~�e_��25���5UZ*�zf�±+�3j8>kU�?ͼ5��=�(��>K� )|O�!��/C$Y�����3|�u���%�W'5c9̅C�:H�H�r�7�Ѽ�a��971�����>����Q��0C;�P�]|߸���MS#�Ŭ�*�����;D�Ѥ��,b�و�w=m]/�nEq�l�z�� ��7܎m���>����1�S�>�
�5[F�m�)xC}),��R����G��&�0��}��������-6ر��O�D�9��r|±��.u�Ի�E���}�_�˼�R+�𸌝���"�����U��gh�S7d�����z��u@{���\�e`�Z6��ȟk'sDi�|,���g�Tk�y�z�l�����27���ףּ����u}w��`�Ŝ-p�@]�f<":3�0�����u�w���v�-2G6a������C���9,jGD��Wė(Z4��JIm�����b�Rm��M-��kp��"s1�f9�y\��b��aL,ZY}�{⪕N 
`69(%��P���qTk���G�'�:o�H{�EnE�rj��r2:��Uv/%�?�C#�`{0F����:��f���5[���9��Z1�[�S�x3&�w′bd��#�g�GI!<��1�{X��G�lS���J8}ڿ�ϣ���NT�D�����`ESF�+��J ����>q�3ޡ>�|	�
H+ ���s���駲�>�F?�tW!�������0���b]�}?��Ӷ��=���A&��u�lt��+d�����S��P����(|����Ĵ����b%ǒ������_cCV���s���jh���/��U���w��o+R�����ӓ�<S��kf���e��Yx�Clt$���y�M�O΍����=�9��KJj늙GV�7����~uѷ
�d�jU�����-Yr�#�GR�*���T��߅ե�>#�۷�h=m'�P��L� Ի�9���Z�hI��f4BT��q�����Ǳ1���<!�θeؗ���w�U�}�m$��+r�m{�7B�]���{|	��Xs^"X(w1$*{W�5�+q��2iT�ċ���^�W�yaI�u�"��kʹ��&�����{���ݒ8U�Ss��qWJ����h5�!NS���+�W�Vs� �����Xk��[I&[A��c�)R6�ml��A�!s���pBYw-�Y�۲�HW�h�cEW��ֵ;<-W`����"���^����S+�a@cq���W���7��O�CF!��܄�;��(X��F�'����_zO�b1����&�@'�/�ԍ�4�#,!�=\����66����P��;�S��`w��[lc��������^J�+��dZ[�ͯ�����bjoVb~'��	�����	f�^�?�e��@��N�����+����ó ��נ,�uqZ5������c����D�JɃ���l&�{�z����GU�]��6Jἶ
t@�6�k� ߰��=f�µ�`TW�&Z�5t����h��$�r�M��`�m�\DH�˖Y��	8������Ɩ1oR��F�r�	\��ׄG���L�g��������/Z����/B��om�|>&m�Ӌ❿�س�%��8�8�4�zl�(�����yKȟ�t}n�47*��Y���j*:�nѹ���m$���٭��q��W$e������Z�Ϡ���E��c��ߛF��ӧA;�K�5�{���Y�Y�Q��qs߫(F�0{jp1��bρ�D�`li+�~�2(x��%g�a���K5=� �߶2��gn~MXG;t�s�O����\q��Sd)�1��)3�dKR�o��<���	F�g���_Z�}A`g��O\/Pg	??8������=��\s
M��F*�:�O3�K:�e�=T����N�O�"+\	m�h�J�#�L��X�4�������ǂO7\5z��:�')a(:q}F�u�u�핃���!��*���jAY�]#����~c:�6�[�&���S��Yw��:���O��6�Ŋ-Ly��ڇW��f���᫮�1Y uv�{ *M���š�-g�G\�C��<�����ÐW��M��]Ǹp��WlQJ�yzy�Nu2��x���=��b�h�a�
/-���wb��.]�\�����SǹT�%�����?#��r�����}∆��P����E5�wHxJD원�;"��K7�bT�m�P~
�?:w�3i%c�ls쿑:���8�4�Qr�ⰳ�����Asu���Ij�r@���EU*M�s�����jq�; zL�����HiP��a3�?gV )$(l�A���߲�{���2y��ך2��}wM<Օq6M��>�Xh�B^|z~C+�-z��KY�ȃ'��L[������c�T�A]��9�`x[�!�.�_����z�篷�6o�eBQE���~�`�|�O������%!���}��FSV F��#���[Ճy�:�#�y�m��l$;��r�Z9�3Vt$�¡�&���XG�!)��ؼޕ�8�tN'�����T�៮��ij .��$�1<��n�3��ޕ�E)�'�ק������W�U�	�o�9�j�QɄ(qg��I�V'*���w�ޘ��f��]��Ր+�weI���~��f����i�I��m$�H���4|�Z��|��ɳ{R��K���q߶'��r;;�p��?����®٣� l�������ԧ5	NЭ�hO$/��V�f��	(��Ԟ�ɳE���X5tNT��n�|��_����I����E�J�>yd���=]��H?�(�D&����ϯJo�:� �'�46z7�ѶCee�v�G�»�4O.|�0�
t,��h�byCqi*ߓQ#>fk��"���Q`n���N�& f����N�j�.���ȫ �rп]t8�����R�Rh�(�i= �[��6���J���� �C4�sj��QRrIAB�k$6r>���ݙE)d��ǂV#���aJ<R�}�npY�?_N���JE5��(א �*��f�����3E�k��o�W���8�H�q�]Kt��)�(�!!�C��ύ��j�pͱ�	'uW�aT9�IZ̵�xH���7�㛕�
�4��o�OM�#>
�����3Cv�ϥ�@B��h_���C#�������;��,�͚�Ǒ�ك�Bw��&/L<?�q����� �M�r�mM�J�,ڇVl�� �%Ű�\�bP�d��}�.Ր�P��H��kB�8���K���v��RY��Ȧ����O/Hc���8KU|=���	FB�pE����̭_E���K���u�P4��i��Y�URjh�m�d.A���o�������h˿����ʤZ�A5�Ä�'�Ȝ�7<p��n�T�U��T*v��} ๕�:07<8���H���Mu��ⓠ���WE;-�@X&�<}b�묉���H������]v���2���a�_��t	�������t5,�����җc�	�o��mA;��b��I�-�rM�ЧkK�+�]��KT4βԷ��_ag��Y�p4{�;<NT��
�i�9#�y�#�9�C@�qo�)E�=��o ����E���A$~:f�vJ�%`7�C�΋{k@ݔ������2��[W2�9�(�1�kS�
Y&�lO�'4_���*�g��iI<�ܬV�XeO�G�DV�Y��3P��P�PU�No"o�y8�H�S��4�e�E�K�ę�m3��Y�+	 .�+۝��'b�D�F���;2?o�!®�\0����VT}��h��꽗g���Ah&��_��-C�{�2+����>_1��O2�rs�����'�?�^���֝4v�u�3��b�_`l�R���?���F�C<5�j��Uc&��rLdo��g�;`-�ЊЭ����FP.Ų2e�x�.tE��4�'�jp��g��pή|qj�"��B��7/U;�T��җdd��� W�@A -���/G�\��=������P����*'=5�P��!L��T��	֙�� �� x�C����ІB�Xq�>���l����a$<����@1�J9�9�}�ĭ�
�rGo��R{{]o��{�gW�(�~�p�(��$����u�q��i�,-�vrL^/ʯ83�I���䮉�&����5�,���˽��-,xU���)3JYTm��5W_�S���f
c��> j���7kZ�IA�{A�4c��@6� .�<�!n�q��O6w�:Y����*�h^�OW�z)�ք�-Rym�QO�"sB5^���G;P+�O�c��E��s�2�ԪS�C��\!W��;�d�c������@@���O�yM1�[v�c�@�j�/��������5��d��ѻ6Q'-�>��$;�����]�V��I�PF�U��ŝ�Ӑ?�$����BI��]z�o�q�'�	�݉�������e@����)��?Ҿ������>��ۯ��P4u�0��W��j}����_�����D�Z��pz�|g��<G�"I�]ҧ���t�j�F�����=��͜W>���2#�"���FA|����%�M%�i`�to\�.U�Q�$!k�^�	��6��lsR�́m�p���?�����LLs�����Ƿ��������B/��*5Ǿ���mV�)������v%F��8�74V�"��5d��tyƵB�On*mK*�5�Y��ż��)�U�@�$3L���B�����e��O�Zl8��i�En�`c��������n�f6ty{}�Y��HQ6��s�I�F����21�Vu��թ��iF�u��K
xw�Jg-ƍ�s7�=��r�2���n��e�j�;�gs���՟I�聆���y2S�f1�-�)�;K-]���ڞ��	A�����_�#A{~��V�PBS^?S��T�O�����7
��F&���� ��Ku�������o켪�q+�K�	�p.��#�������/ ��y"�$7���d����(�C�G�u=�2퐤ɏh�w�a8I�gg��g9�8�#�p,�<4�1Ȑ���{*��t%�ٵ-R�*��q��ȏ#���zWQqV!�^��D����t ��	��&M.��Ŝ)yg���/��WK�����kN���u_]b��p�'�l`=s�4�i�G�E�~ӵ�ѦW��bi�5�\��/��v�2e��I�\j�������<�%'����Ň?~'��- ��H�}]q]��H���x5�F	H&DG	��:)�fEډ�K]�Hs�~E�c:��i ܲ���L�ӡ�S�4Z�Ȱ��ٟ:���'rdu�-�Hj��8���CU��s�4���1� u[06�2���uik�a}GI����V;H=�r�A��p���n��y��GR���giw�f{�0�qM��ﳬvBL!~^�A-�FeK4ї�bQ��l)���_��,��c���AxMb9%V�[��*.9�X�{�c�"·\&�o�K�Q`j2�Q�T`���O�jB�Ar%��ZC>���V�IM�h#��[���Ǧ�t�T�+]�;lv�$�� 31��?���<P��`����G�o�)�z�Y��8�ſ'<���Z���O��	2��$|�.�#dݬ����i3��ӕF�ͨ 6W�25NH�����*�I��L�c����%Eg�s�BIW�iz����J]{JqՋ��w��ʶ1d���
��D���Zm�V!��7!|AM?�7���pW�L����bV�r�EP�k	>?y��E��پ�Jl��s�����V�5���ϑ�Ow��Pp�ށ�Z��V���҇�I��E@w�X0hjTX���)�e����/�a���rqJ��y_�X���Ϗ��C�D�����w��>?պ��o'F��z��޶^�e�%��"����ɝ)0�_2,w}u�#5
y0��q�e�,͏f�{^"�%Q[���^ȧ�
����uu�	R��j��G]o#{�=YR��U�C
=|3[����2�Yb�������s%�QmV/I�}Tk��]>�	��xg�)__����N;,hae_���T�p4�_�ҽN��5�Fg����*NR�f0����3 Vk˷S��\D�3��̭<K/p�)�!/!��MCڐ}
��iy�k�ƟdH&W��)9.��0��Hg J7o����/q���B��k>%i�퓖��fC�c��%=��ප"�#Ak��~����4�tE�Gɪb���~$w�0/*}���p�� ��i�b�m�cy�:���9a��x]"��+b_�=S���}<Tv����B���Zo��S��s*5�$Tƍ­�c7]��,�O�k�y6��S�`|��K�䞿�J��EA�2�;�_�HŲ�eC�&;��˨s��mr��U��h�)d��U�|�O��k��˚8���TlZl��')m���k���T`g�/�J������
�7���e��3�Rus��{�S˒�-�CD@S��<�ѫ��׉�_�k����H(v1d2}�a�����.��tb3��\,`����P���S�
&RmA��sb?꩞HU�M#�k&�أ��%g4Z/�u/3&�ء�a���Ys�{��N���
��m9y
�~H����q����W��raoT�t�{m�E�v���:!��vek%�N�C�զ{���/��Z�썿�[�d9���1� uS���&�Y;ⶻ�Z;:�5Rg��IW�'�'�X@�RG=���.Cʿ�T���N�wa��qu�P�S����  C��x��Kp3T�^t��	�qZ+�P"�bpA�ߟf靤���?*��!,���80�1C�o�}u���>������D2&�r�b��V�"+�㰍�
G��n��cp���������F�@���c����L�_��u̦b�,1��+�����U��|�mLo��E��?���a��2�&�!Z� �je��Cx�#�t��(��h&��2}���]��$��V��jIz]�=��7����uJ���D�d������{�y-��6�#LG2J��{e�(�
�t����-�Y=�bP�LY�U�I��jc�����AmB��q���a���'?ة��Y<�h�zz�YƮ(=}�;s7aTr���m�^]�j{�su�cG^�ߠ(�ڑ$�]ē�"5q�#ciJ��Q)�^j\��WI���?[]��C��d ���:?c��pPU���m /J䆺^5ҼS�h����팲r ��n�Vk)I\�dA�<>c�y6 �C�#W�!iD��&}sw�{Y̛F�>�h9	�W-9�q
�-M��Ϭ��".�V^�"�yY+�]c�j�ōs�-����7C��!	}��w;����D�|������KOm��1��ޯ�@���/#���"�w@������Oֺ6l��9��[;5������Qତ�����Ly�!>����Cz������X��o�p'?�	�O��T{w�! ce��P��$�Bn��y?�QŽ��Tۊ�p30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮs�
օ8�9�/���q�!:`r����"j�z�W�V>�n�/�M6�
6;�?��%<�0M��HPn{���wLD�����,6����8H�g�,����I1����#������8���'p]�DK��1����m��""E0+�O�zݾ˺�]-�+"���/�|<.��A7�#U����b3mO�����Q��DI�e��f7�uk<��҉�E���٨g:����5�ou��,f�J�e��B_2W� Iޥ;��j��'w|�vq�=��� .�h23����D_5㭵R����9#z�ꄛ�"�g�:ȪY*��Ǿ�1�1�!����N�J��G��Y�^b�z��+*�?�ը�3���4o��n��Nϔ����i�@�W�ᑭ�3�֥��Y�CQADN��7�NB�@�MePY�Ҹ�w19�⚚�{�2�:��r�3
��%���h��2�����P^K %��D�8ư^�@`��`9{=xHxU���ڂ��7��Gb�x�����e>�NF¯���a����b��*�2R⛯����bNR��3� x`�ZBs�� KIր���� ��-�Ǭ�R}�u�M�4g3�����|�<:r���gN! ��,u&�:��G[$sF*�MO�/��Z�b�D�g�;��L��+]\T��}�q�O+!tT����<��8��)����w-=\�S]"��X����󣶱��˨)G9�n/�3�x�qz�!	D����_�'Ȯ����Y潎���n�?u�=�UJJ��g�ݘ�������j5��� vjq=�K�H���Ϛ�B%���W��F̷�B+8���j�aF�	�
|�a0�i������.��$Cļ�E	�«H�����ήR������i��V:-�5먔���������1�{c�q��:�kҌ l�:i{��E~0�Oد&x���Q5k��
�1c��z�|��E��`�i�{x�� �%/
5��i<)��wx����Eѻ�
�������A�ʠG,�T�7���䔘���,ØfMB�F�$Uu�qUFe�i��ڸֺ1�,�˧�u������i݌�ذ���(��a��>�B]ˇ��J�B��Ʒ�h丆�� k0Y�����2-���-�C������Xj%)%����S	���B��" r>���r�:n�íN�`r'iq3P~v̇2]1f`e:@�<�J��L���j�"ȁ�W)Çg�S�[���(g>� �a(\{">�x9��I&M�JX1�O�1Ta����7�3�N��g;�`=<?���?�W�@�J ��c�qRH��v�G0Z;^���(:��dCL��%Y��V^�nHB�km��ڷ��9y��{�[��n�<����$F�X����"c�p��Z�����ς�S,���������q����Al�=�ZGl��Xˊ��>�˙D�N0Ў~`�m�D�V�=�����<���#8�V��Dѣ��Ϥ���VS�;��5hD!��7*�cDQ��ͣ_�(W�(��]���}Ϊ���a������{gB��/�6
_��"�4}� B̈�O��2N �We=��F�
g��oK�v���d1��@5Wj�\�cw�*�z��1O��[�gd�Є	cL���Մ��ZΉ���1R@vv��6f�т��X:N<��֠����AU���ћ[4칠{�'
��~G]����#�u&� ��a=�����ҷ	�(r��S����f*�F�˷w�������A@a�r����A�ʒ=#��e������/{����R�C��P�6����Z��̊��q���^1o�=�)m&f����תk��b�k������sQ�Vtb@6&��)�Z8�tW�,j���!��Ls��1���w��H�M	rَ���=��"�ħ�q�t<�u0����M���1��������'X㶨?���M�<?1���xR�Sk4 ��U��B'-m�,�o�y֐��������`�4����NRƲPb�q;"���?��(B;�Fp����'R�ؖۺH���S�-��s�Ɖ��Ɉ�����特��e�`�b -*�����õ�S��*������z�=I���B�:�#�솵Q��z����V�A�����y0���:Bi������T�Ȃ�Q���]�e��6��],��$~ |��i;J�*��Ҝ	7\A@u�.�C�����D6WN;i2���U;4ܺ!��C��@D��h� ���"?Z�Ih'�Y�Pᯨ���Cŝ��p�?��G�T��_4^j��PϠu���5=A�Y�L�g��hho���Uc��m��V_�
O xL�2�����ɝ��![H'7�6�%ReA��������IM��\�X�(fE�%���w��O��u��^(�2�ɋ�c0!5�h�"�<����u7(^D�ZCӢ�p�#A��j۸��Y���g�0��Y�dX���څ�3Ƽ�n4#�H�J�.��/ۇ`gY�D����/�J���W�D&V�d_���z�Cw��$ $0�jx�l��ύ���_��d�%�0P��9��l�/ilHAY,Z���e�m���6['Or�9M3D~���C_�
j�Ã\���u«�	����ţ� �Ba�����c���3�e��m$�W��q.� ~M�EEZ�I���#z��r[5c���@��:���j��1�}�?H�7z[a��Oz��o�+�@N�݆��z����%i�NA���Xm��S��b�1?��Py�df��E�<�./�����}�-d�Y*�s����{���|�~0.�k���@bcY_���WLF)+4{�0J ܢ�ͷ$c��=UD�Ŗ�>����X��hbC�uy"��։zÕ!�Ug˃U��'Tfn&?�/_ӧ�'���6�)G�T�:���� �<-g�]���/�W�4E�X�G[4���5	�Ҿʔ��<G+��1���=��i���^��� 	(�^N,R5���Z�T��Y�x����?�{��=�o	�����^�d�t�*o|h��53	��v�9��SN�����	��bᢌ/J:G�+f��Do%�ߴˏ+w�1���w	��@J������0\ d�q�q���~�c�d��J-����zv(>&�q>2����\Iƨ�6����4���_�R�q�önC�e��/�)Kc�=L����p]����F/�z�X����W{K�Ш�A�H\XS�%���ff�XL�}��ꅡ�I��Ĳ�/��@,%����ٻ��r]��7�0�q#����=�[�F��5L�cT����-�����/��Q'`�N���[���7��E����|c}v��f���ǐ����R�!«�2�*[e����U��f%�rK�@�xځ��������gaX~m�}�H87-Yz�D� Z�tt��s��h��ȼR��Q:*�V�y�O��RDJ
_*�^ܲ�g�4s��%�i[R�%�,�� ˦��t�h^��3g���l�	2�1i9��c�A�?��'t�O?�)~P,�4,�|�/�;�A82C� ��x;���mlF0��d�%I��7�}���(	:ɜ��O �5�mEG<,Y;���q6�ɰ([|�M�d���#i����cwl�|3� 8�Q*���H9�D�8P��R�b���Ԕ�;3i�ʞk����A��~��!�h`�S�����j��R܄vρ#��n�NQMC�6�O�ѩ٩[:��~{��D/u�>��^!6\�x朇H`Ag5���1Q(��WV��Հ���]o�ɞ=w�
֝�_�P"��5�\Q`�'�@�e]]}5"i}�/�PS.uB37V�q�����V�Ou�u=4���1DJ�?eu�G7;&g<�JD��œ�O�TY�Ҹ��D�n��w�������Q���}����sm�V�x��>��b�֞���O���Q����q�B�s��Z�hp�uǅ�A-jp�2�=,�t��Ŕ,J��)�l��K+��"i�R��)3�h�' ��#b=��̯�i?��R� �
�R�׼��%Pdk>M�9�Q�]��@E�;��� b0��y1�p:C}��ÜOQ<�;>" t��i{gҗ�y8	�J�~K�\�-�WS"(TO4S_�붦G�7Y��`��A
<�Sc4���٥G��d���-*6�nRX�`��'��m�TQOQYP����o�xh-�\��MNZ�g>j���'�����UB�v��Q����"�kPQ����5�1�~��BɚY���0�r�~��=q���p�H���.��#�n�����W~�m�t&-��-E�2J�����ؼ%�n� �Sǜc�\��#����ki׻��@��@&̚/d�/I����ȸ�6�ԗZθ����M"2��Y����2�Z���gOE�f��7o*^�Z��"�V��4�#���l�|h-J�Z7�oǙ�t�/�"M� ��aI<�p
��|�{!��wn�.����7�s�I]T�\�����@b#偀$l��	 �G^��M�^�q0Z��т��#�V	���,u��4����>'|0(s*U15q·^!����k��n��!y��Ϧ������XY*+����Q�1��3;�?�^����׀�ܞ��)�_�h/��i5�r�?��馡�)��v�,qU�>��u���5�(U�AWU��e����n���"�>��#8��P�po �Q'�9gn̋g��\\4�9��۩�e�I���r������"*�E��"u�h���i��e�ʇ*my7n�o6���?=����������W����ac�'jELW��m#��?���D�j����Б�1\@��9TL�����ǳ5�)b��Lx=��V�^t���[�wj?~��gl��HV妀�����&�]��"�� �<���0��H��xj�Eُ$� ������ W�Z%:J��ڷV񒇣Z,��;�G���R�Wɤ����C����{(�| Z��;���l��	����v1�/�q�C�Ԭ�h���>8�#���bB��´��AY�QjFI�z%�	Fk�o�*���$���SK��z[����K�<P�:(0,*qDQ�a�O��UM�=@�L@�e��'D�2��&��9s�?x7���L����4�z UU58'Wj,A��y¥&�w2q��m���*4~���GWcƞf������O�a�9��FܞK����RA��ۦ[w�d-k�Q�sN�~�x!��$y��s�%w����S`��-r^�A��������+�!���z�׶�~�B���# O;�=��z�NއBTn�����e�Z��BU�1� �\Tq�����{�����"�t�w���A� �N�i'R<*��Μ���A���.�a��g����jW���iP���; ����mwC�E;DkR���bێQ�Ʃ'�8Pͺ%�Yq�C����晕��Tjׯ��^֥�P�צu(,z�ׅAU���8�`�0�z[� ���YW���9��2x�~��l����v�[���{�%��Z�������I9;͈�v��v���ݾ�������u���^ػ��7?��Qq�}��N�"J_��P����^0�C?�gp��%�W�L���Y��e���B0;����^�������(��Zskݴ;�J��ߩ��PL<?�"/���>J�IWᯄVr��_��v��U�D7wa=$�����l�B����_�d4e��2:�J�9r����~Tl4��L���݈X��ߏi'��99wL~c��/N�v����*0���`�_�xذfU�1x �]P�pd���	w�e�~$&��).�S j��E�~-�5{�R��zϦu[��2���������)�V���i^�H���zG8�9v2��cG+i����%���;���/̺��p�+X�h�?�=bO�����yy%�f�(E�/�.UZ�cU���x�����sޒ��w{�KF|.YG��*@N�K_|=�Co�)���{��N H�ͣ��f�U0]��`��ڂ���/_oyx���n��� US�`�bl'@�&��/K���?b�"��G�*��&���k��<�]#.,/�i�4����3���	s1	}�5� ��<3���!�ε{ ��ƥ���4�{�	D�N�#f����Z1~�E{��@r����{�Ę�[�w�6���Jօ���H��h�5�s�k�b�%V�"�x���ڞDa�J�y��	��F�p�)<������%��Eh�6�>���%	��N��m"4Z�D.����T�t�
r>{`��BmǦp��ϑ�����hf$�5�׊�۝[����/�]�H,Cj�����~0J��	+BAH���{��Q�������tL�7��u�Jޜ���f\\q��Mqc�H���?G��Q�ܜ��i�֤i(q��l2���J��I�$
6G���&�QU�_t\�qbz�J�C�qe���K�m�L����K���	�Ij+/чX2���_sKx��Є��z�\4��%�a�fB��X�=�}�O���l`I���i�5����%��� )��=��l��t܀pks��P���đ-c0Cx4z-\ ����^_%Qzq��*u�ٷ@@���Pb�������}R2<fݢ��l[��@������f*����8 ô1�/f��KK��x6��kF��:2a4ځ�ٗ�8���8�����-���D��wT��r@�R+u[���?���2皍�D#R 7�_�A�^�Fog�C.�� �űkG�,7[L˂�Mt�֕茰g��l� ���[�����AE�/�8t��c��ڗr�g;��}~/ՕVA��T��l!o�T#�"��H�B�d�������ō�uL�(q�x����a�E�m��,5�����6�BT(�M����>�ﶂ`kcS���؜�����ǭZ�̄>ϠD�P�5��``��sɌ�L�3E���&ks��,�ϝ@:�Z�z!�`�9�B�jjzX���ޛ��nK>�M�v6D�(���A�y����{K�t� ���{ɰ��U�6��HºQHa9Og�9��8�	1-�E��~)��Q��O��ߦ]�Y����f�;��"j��8�{ꃭ����]v�""E�l/E)�.Q&�7� ��I�k��O�����Z�w.D�n�eQ��7�!�<��9�6���l���ҔU�DHQ�S�y�,�x�-0�\���<��RV�	��f.b]q�D i��e��{�����o�ڮ��o�Q�Q����p^�=��:�����I�������(H�@�����?�Rf^3�3Ń�ϊ�F��LMn�E˭�3Z= ���R�%<��?�d�`�N	��7	�-�8� �t��	�g
0�+y��::���U[QV�>~?O��k�#g��y��Ⱦ&��KZ��	��S~��T+e���j��L��75K�`�
�7nS��`ج�n���d~%-��,n.��`f��ą��dUQ5�w��G�T�K-���)۾��f`���%�����|-tk�, �k,��e/5z�$�'���Y;�S��>�ڭ�ƫg P�LjH�?����n&����Q����&	ڶ��AX2&Gֻ'Ru��'nR�QS����i-D���?�.�i귊�P,@k�/���va����`�������W�Z*tP����"��D5���;nZ�.g��f~�o����6�".�\��#�4��Ӯ��|ę�6/o#��t��g�~� �K�I��%
�y�|!�!�Bq]���s�Q�7o�Io:s�[��)����p"#A�F$H�$�er�#����:ze0����^;P#R���E�u*�4���� �>��0�O�U���eg!��Ɋq��k��S�K���Ι���H����WvX5@��2n�-�,�G��;�8&�s�c0:�ܳ��z�)2B2h�\���r^T�EW���vdQUǺ�>�9A�w�p��ڶ����8����M�ʩ݌�?�>�.#��P�9�o�L?���9Cb��!A8�]ݕ�ڜ�+�e�Ȥ��BF�c:���s*m׸�x�I���R�E$�e$	*I&7ʳ�6w�?�V������4�W�u��V�'L���m�$�?<	D�)�Uz�m��c�ڨ��L�B�����#����_��r/�.&
�^Pb ���j�������$=���X�t��a&u��Ə �^���@�օxF9Eq7  ���;`��f ��j%��6k#�n�Z���;vH��V���3���8��˧J1(���Z���W�l"|���g�ҕ8��S������օ���8n�V�p� Bc (��SY~]�F�3%�|Jt9po����֣��S������,[-�\�I�@���D]L ?,�?���h��	\[��O���C���l��5�0v
�Hhr6���a�o�EYբs»#����5r����'0��l=���G#����'w5�Է
Ts6Kb�n2iɸ��o^>^Y�Q AM���6N∗������{\�{UX�j1Ѓ�����E6�L!BCH�qg���BY�1w�݃v$�Jb��?j�'(]U\ ��C�p7ȵ���"��}���G��-�] Ә"��/O��.���7<�������u �O6lV�[�A�D�g�e��q7!��<K�]�v��E�:���^�DR�+靉�ֶ�w��.�)4�?�YU�V~]�3�b�|��7z쎎ɞ��&�<%��(�Ϥ,�y���3��',p(@�=�kv�?���z ��������I��1�*�ȼ�R!|b3.]��z1��Y�VXB��7��O@ T�RR�ҷ�dQ��I�����w�2��ñ����q��0W�y`�:鿤�)4hQbg>	v��u�<g���y���bKd�j�S@S�T��W�?t�ܓ��5M7��i`!�x0L�SII�v�襭��d�N[-N�n�l`��D��:�]Q�G��$n�����-��������V��{�� Јr�ܺ�x�w��̶F�k��$�V�5ē�d���L�YE�V���d�����q[���&ۦ��d�?n0�� #��S�C&�%���2p�]�����"n\%�S�-������$��8�i4���EU@5^�9K�������֪�������.Z�w���B�"��9�y�x��Z��g�8f��o��� b�"8\�?��4�k��x�4|����=�o�d=t^W���i� o�I"vz
N��|(�/!;Z'����g�[:17��`I����%-�3�b���7#�X$��o(��m���'w��0���ѨG�#ܳԨc�cu4?�4)�x��en>�sC0�d�UWS��!�Le�{
�k϶����_��y��o���v�X��|�'>�wd���.;k(g�\"�:v�fi�DQ�)<��h'|\�O'�r(n�O�(�OQ6v���U��>��������C��˵�Bo5�+Y�T�T��X�>��#^d�P~�o��.��6�9�jk�M3��ݟ`��I*ep�I�_ڃ�m�*�#�v*���B�����ӏ��e��(*�;7Ԯz6�]F?#<��m��>B'W ���ʣ���L��SmI+�?�lD���_Tgз���q��r+L���ӫ�ޭLν϶���:����c^�����jeX�M�m��Q'��=��@ָ�~d��0j p����\�.d"xGgE{OJV�Ţ�bX� ��a%`������8�Z�;�����Ԓ��l�Zɞ�oj�Ԓ�(LJiZ�
��8�wl��6��~��v,�U�ç)e�a����%�8��2���_B-g���tY�	F/i�%~c�~��o"�{���ƼOS�m��A�[[�&�\�Z�J"���q � q?S�h�޺	�[��-���ƫl��5�?�vԍ<h|���*���1Y����!u�`�!5���W����zE�������!i'����A��s�il|b=�f�3�2��a����((x�wSS�W�f���,^� �卜Ovii��z����-.�t�5�:��ÐC>ċv�[ϛ��<��M�G�=#q���AZ�H}���o�*�ǝ��޶�Ы�(�([>b����u�B*i�jq�ǝ���b"�woʐ2n~~�w�t �Xb7*�$O��,<G�t۔���k�l���	w��s|>��i��	�2Qe*]��
�Mɐ)P��v��*w�Ħ0?C�MQ��4�Q��#���J�+ځ�,l�`��Zm������.8����~؀+s_ǰ۪�}�,�<ÖBf�kF	��8K��]�=�ʼ)�F�|DCs�0�9�e�\��Q\���{߈?�`������V�!�%��n�C���ڗ��ߕj��TL1M��pYɼ��,z�Ϸ�FݑEx~~S�])f�F�Q��{�ӹ	g{�C���t�
w̟���o��hF��+��BX_]w���7A��5����]�H�ڤˎ�m{�ʮ˺$�Z��űS�2F���r�u�����>�m6�526�?I�>ך�G�p�%�{��s&_�O��u]�I��T��u��G﵉L�и����;1!��.�v�Tl�1��#]���ŗ�6��	�$��!�f����+Prz�����>�5�7��0�������.��0�����%�ŀ�qMT�oD"�� �����D�-=%�?����ib�\xCBX�գ�B�!)���s!�+�ů۩S04B�b��$�BW�t�e.L�p�	If�#�7��"\����d׹@J�j��ǓJa��a�a�hNF}M-v�rwo�w<������x3�[��Y��cVE�dM��d��0[a(��RG��%p�
���c���iz��t,�=�<~�8 p��R�������a/���V"�m=�6<�c������#-�r�����x/�y�ܼ�e{���$�IcE����P�8�i�y����z�I����$K?ɲ���gb�ă�~�"L�����y�6���}�B�/��_I��;��~ΐ�c���)"g��;��2ھyp}�˘�P�R����܄���[2���b�(���F
j�y��5~2*kIS-��N�j���w�`�v$OK�Y� ���2���#X!D�㠵،��ŭ���਄Q��:�-��VY�Z��
�b�1�{r�������G��Yru�m+}3f��w�3َ�4����A&ˁ�����\mP@?4�D�3���Ct���DM��1�N5��@��e.
��1��N�m��{)���m�/߆7����f��h�����{���꬗�K������y��q��T�9N�Mx{t~�%*#��ː��ՙ+u���@�e�4�N�%q;����o��@�2T�µ�����N%��3�"�`t�kf�U�q��I�d��l� BcJ���\��quvyg�'_�7!k�/��:�q���vF!o��#�au�+�:�� G�#F�maO�Oe�ͤ��7g��&��ų�O�\�lT}u^�O>�aT�����%�k�U)#���j�f\�d��kz��O�=��L��9�)��n"i��˳�z��^�~�xŧ��ј�A*y��F9Is�=��쩈���UG�.���+�����5�Z��/b��jD]�K�b'�V0?�5��EŖ�aB�Ҵc8��j��c�<��|2���T�&C����7��1|�	�(|H�w���/R�7�HCid�VMe5^�`u�F~͑/�� b�pa�h�\�k.,dL����a_���C���/�Xe���IYKk����If�-��\G� %n�f��X��}IqI���=Iدk�ѷ��Q�%a�/��'�|����+��|����Lp��֓���c����y-����| �F��2����`��'�}�u<�����|�r�B���i�:`�7JR9���r�i�zh~_�퇊�x���:�Y��gtLR����-�z緵�3��� ����kـr���a���"o�͔lo�9�t&� ��	���e�OL�Xa� ���{3b�[�;fh<��}YӘ�� ��U�nH4���;������<����L����N;V���H�/�m����]9qه��-Y�*E��a�����:��3e���1�pL�R����k�ɴ'��S�U^�I,�l��׺�)A��������=�؊�N��#�롦"X�֝"m-�V�G���NɔY1xr������&
�ݳTV��;��h�"%��J?����Qwߣ���(�D,�� {�T�P}&�E��e��	���B��B��ơ�X
���z�t}��<B$e�O0aNx�W��s�J��
��o�D�m�ٻv��d�^��D)W�N}\��w,��ҏ1k��XdK�	�N\�wL��ܯ������d�1�yrv�������m�_����.|��	_5Йf��9
��!���i)%ϐM'�][7�-�S��&k���e5=�ڪR��	�{r
��S;���᪞����ն,)��tF@�qr���K|ӄ",	#ل��8F�4j|��'5�f�����Pc}}�PZ��u���Vq?�+^��m=2�&���epU�/�.�%�k=��P��s���t� �&"��j�8$7WTy��ʖ!Mjxs
+��[���6;r�uv/Mak�m4��89��K�{��qa���W�k�YM�f����;yQp'�����ڥ�$?d��G"%��??4X[�UA#�'�,-�y.��c6G)¸��4�6��3q1�
�%��SS�9��M�%�F�y8�,�R-�>�_��P�㎅߂s:-נ�����+X���3���[��`�*g-���-޵&]v��^J�����M�zU3��jr<B�#Ƶ�۱z�凮�a��z	�����B�(�읢T݁�����꽽R��~��c���1�c �ZIi��J*㪮�a~�A���.��R� �$xW���i���:m�8az����#��\�b3i�Ը2y�:kf��E�&.XI��@я�kp����[s�]��o�{��q|�K�.D:���@��G_�ͽ� �M)��
{�ْ �h���y�`�$U����:����@�z�H,')y����)����U��ް�'��&'4/H.��0T}�_QSG_ڵ��L7����<֌C]���/���4N]Áp-���	������<�����RβJi�ru�J��X�	�I�N�؈ۺjZ|�"�B�L�<���C�{���ػQ�S������y��.h�M�5\&��HƵ���D������W�������!Jc}n+��F���B�h���ԙ�̨�����XJJ������\i![��"5�����,��ޔ{�����j~(���q�*�2x����>I��6�
L�9C���_���q&�F��mCJS�����KL�LL�����
�=�tVQ�/~P�X���L�lK�.бq��G��\�k%�f�#�X�:}��u�nO�I�.�6nƓ%�FZ�b����� ���Z����|��f��@�uĞ�c��/�	-I�l���+�M�QG%���������B�������Y�e�?}��f�Ӟ�٥��+���:�I��*�SO����^,fN/(Kv&xC`��=��fa!0��f�58@u��C�i����?>�q����_3�R�ŕ�(Q�z�$�������R��_�[^��1g��B��_���|�,D���/�)tdP4�չ�g�k�l�<�Z���}�ARF�}m�t6�Bx�g��`�Υ�./B�
A�͇���y��{�A�m���uk��1QU�n��ࠈ��"q?(���e��8!�>�;mn&�,���"k6d��(�wM�%i�q�S�I�-�Oc�
M�����sM���ƹ�y�-@�Pʢ��-s���5ߔY�3����s���F�*y2ԇ�y!ޒ`��OJ�j'��-�����nسML 6�֗R����^��{�l���	�|��Yr6��/~Hnj9g��ܐ�FD1tՃyn����թ�J�g]��5��G������(�"����e>��P1��P��]�9_"��>/���.>7?����=�8�%OY���Rd�$�dD��e>)57$�<�)��хb�h)��!�AcD���@�-ֹy��Z�V��V��b���4�Va-����bJѮ�� _��K�H�_$���lχ/w��F3�>{��*Z_p��B=U�h�b����m��*�Ҍ�5�x�41O�+,�R���3Q1�Ő�;�������D�2eV��1� ��'R�L�A�d�6n�媬�����������Dg��4v�09�y�^�:̎��l��Q*/>��ن�8��g�y�拾�K�8���!�S�aTXŚ|���3�Y�@7���`d\��E�SLwo�ٽV�p��d�a�-�Šn���`b�'��0�=m�Qb�,��;����-E���C���M��[���a��稺�Y����9dxkٿ�B�(5gfMg�%KT�Y�yY�������x�9�I�̙M�ǧvn��!�Cc����&�Y��ֶp2f���N��.��n?S�΀v�d���o�{'7i�s$��e�@�~��w���K~���֍��ag�흰�Z��Թ�"[�����05Zq��g��fk�uoi��c��"�k|�bH4{�[��|c�#��o�}ot��W�K� *�I�XG
1�:|k��!�Ѩ�3��%�%���7�sKI|f���v���=|#��$un%�2��������F焒0H��K��#��j��޻u���4Lq/���>�?t0Ѭ'U�� I�!R�>��k���X6��{^��OT`ί����.�Xbh{�������T�;NZ�P�Pqd�iܧ��)�w�hJL����:rӢ䒫(��z6v���U���>��П�����t���cŃ�8�H��W�M�+*>���#��P�o��=��]�90zX�P7�e~��bq�$r�e���B���W۽ƪ>*�)ډ�=��Ӳ�~e&�z*���7��6dS,?&���2�y�WC�e
�꣰Z�L �>m�"?��D�w��"�~��6�p8��U�TL*��v��ް��2���]�_��^�k���j'��P.y�QU���v���d�n�׫-3 b	o���X�1Z�xs�YE>�_m���H�E�(  e%e���+��x,ZU��;�Y��c���Nʞ����.�(�fJZ��¿[�l/x�R�����Iϧ, ��b\���8�� �}��Bے�1�Yk�HF2�!%���A�?oE-A�M�ƟK�S��#��x[���\�;���� L_�?6�h9�	I��[��r���ĭ��*l%��5q[v���h�];��r����SY�G)���_5��:^��KP�������$���;�'����tos����@&=u��6���a��M�K����W�:`�؎��Jb�#�q��!v,�םL�qW�.��-�S�:1�!Ó�3��y�v�.�[�g����!�0��Ѐ��q}z�D4�H��E|O�Mٴ�C)&ޙ��������s,b����\*,�@��.ʚbm�o4@n!��w��#���*T�2��8�<�zn�w�������a��w�sl|�F��,A",;�Q�ƽ� ����)�A���C��-އY�?f�QGK�4##^����+���,e���#��â��Vv�R�88�N�!�0+v+r�>��}pu<懋��F�d08�yh]Xpʿ97)F��?0�s�a����?�הq0֕x�ߋ�`�?X�O���D���?*C�F�@����ߘ/��\1��p||�E��z�.r����L~V��]�~�FSv	���@����&7q�bB^
c������K��F�ܫ+��X���wu�h�_ZA6��TR4�����1�m��ﮮ�ꠝl�T��2IU���j�����U�m�l2�`?��w>z
�G��Ȉ�1���_٭%#/�,\�T��u�d�G�l�L>h2�c�E�<7n!E�YD|T�F0��y1��&��w���0GM!Bof��`�l=r��`��?O���?���]�S�	�!�߿%{�����~�(N��KpHM�gw&Ճ���7E�-�k�B
y��&b�,�Ce Y�&�������l,���/���0�XJb����e��tzN/���L�����n���u�4�''��@mF��P:�JD៼��a���NIyu-�v�:x�w_ܶ�g߽�ڄ���G�l}�L�`������n�h[�R5$�m����j���Ĳ�]�69	�]���s�<J+X�+w��u�!�0�I���M���v�a�wB�Jsp��si\1^�°��]�B��7������|�i�k�g(OW�qog�2@��_q�IW��6�k������Jl_��q�궿�$C*|��@wK5L���������/F��XG�9��vK̈́w�y{`�6\in%�f�ѰX��}kԾ�6�_IzcƲ��h��u�%ã��*y������5��"�e#�.Z����f�:c�%	� -o��O�ES/�Q@��_�ٌz�
w�w�]�[�-��}G'�fr6 ǡa��'r�=�*��e��O�&�Df�K�ywx�,��R>�.��a����.L(8/*k66�1�r����9�,��4��'#�R��`��R�B�L�g��� R���_�f3^mgT��évZYw��Z,<}����t,��9*gi�l��1�"�1�ߠ�A��E�/t��O�?8/`�u:H�m�%/
��Ai����\]�ϒ	�'w�=����v�6�D�h����6�(�:e�-� eݠb�m6ɔ,jģ��w�6,�I(̎�MTř�9���1!���c�N�����oɸ���Ɓ��� P��ɂ��(��5�!�3����;s6��7����O=�!�`Жѩ��j��5��+���n�$�M�;6�U���m��N���&(�{`S'�Փ���4P��+_6Mp��kH6G�ge�Muc1�{ڃAoUu���qi8�l�]�����{.V��Z"c�e�-����a���]K�D"���/Z��.�x7d�Ў�� ��O!=`��.���dD��e	�7젬<v9���"�0���ė�	��D]j�� ց��"�q����*]��y�V)�㯖�bA뙉��Ȟ���''Ȱs2��OUo��%0�3=��
pS��=���*o4��z�a0���������)���=BR�"`3�l�X�2�t7��aLv������rA  xR|���	��d����㢬�{���M��U�b�	���P�0E�yb�:��ڬ4�`Q�u>�a��p� �Ag�gyiۗ����Ko�ʾASӟjT ��DR�����!97���`,����'S�Hء7\�8R�d�mI-[JMn���`*��y���Q*�Ӻ�6��i-�������^S�z�3���g�b�N�y�k�m

H.5/��/��YЎo�A=������>|'F�t��8��A�n����.��f<&~������2�5��|#��c�n�Y�S��I�>�N�t��CfOi��D��v@`�(��̫��`#l�U���)�A�exZC@�Ї�"#�ej	#�í�Z9Ýg�Pf3=o�	z�+��"�^c�*��4�?��#�|����aoxf�t��(�
 � �Imer
�o�|3��!�	��d}��џ��5p7�OID���Ѐ$>�z�g�H#��6$= ��~\�X����LB��0�6�m�#�������u��4���ե>x��0���U³8�hR!�s5��k�T� c��C$@��
�w
�׬X*�j�����b����;h������1���onY)�bMh�o���7r�(7�Z�G��b7vg��U���>�꟬l6�Yy/���MZ�dxދ����k>~aZ#I�P��BoYk���w9�����-��*4~�썺e�q�
9�x>���j%*�☉m+�Y#c�z��e���*�l7�*?6,[�?����!A��ːW���	��x�L�M-m�c�?[Q�D��ّ�8�Т*�8����L�CQ�>r�x-|���w���C%%��@[^Ź����j�����GҦq�F��,�6�>�sÑ *X��L����zVx;7EE�5���'�f� Ȟ<%��Ȓ����c�QZmg;�m]�+�6��<���Pτ����(w0�Zu��#�9l�L<K�;�����IЧ����t��},�8����E��Bؐ���"�Y3�F���%�?�	[do��Ա&�gI�S��dҬn[�D\�1��ާ�y� �?�b�h�^	fD[K���刭Q�kl�Z5�epv}�h��`�w�m���Y���P���K{H5�[��4��ړ���	��Ş��d'��Ԍ�$s��9wP==c[�A���Sa�ݕ�b���ʉ���q�f��B>��̍��v����e�7�9l`.zPf���:�=�[�Ķ˟v���[�KT�a飧���HOJqE����ZH���O����|�a�ж�'��Cbnܬ��>�*�8\\�����b��<o�r�n�EwR����*&����<����?v�vd��)P�ww�`|i�r����>Q�CA�r�Xa�)l��M=H�U���OLS?.3�Q���nq#�te���+��,-�A��ѣ�jl� �c�c8 +�����+>\�A�}8�<�c����F�R�8V �] ��ʇ�)��(��sܸa�K��F�\`��]@1�Sr/`�&�����-Cb�D��v���*�`8���+1��epDǚ���z��� ב�s�~d]T�[F��f���T=��D9�*	(
���^�U��F��+�}XLP�w=.&�'�A����4��-��䤶��mƚ)�vPe�e�:� �2*��@��z���(�m��U2�F?TCt>B�rG���Pf�����_����)���T��}uR$DG�%�L:q�+�^���!�!��!��Twu��d��_����4/�V���r!
��fQr����tr~����?�i�8��:������߇+`��;��w����v�KM߂t/�z�K?����屳-�K"�
�1���b~W=C-����0��=��������� K0_��b^U��-^xtBJJ�f	�lݎK���4��!�@5Z���J꼮_Va��N*7-�@�{�w'8ȉ/���#�I[��Bڊ�c!�yd0��V�P��b(�{GB�Tpƾ�w�\cr�&�����Z��t�?=A�~K�lp�R*�e
mt}�aZ ���1����=̡W8p�i=[p`��D��=�ʩp4/���f�{i��$Ԏ�E;Ə��c�,i"L��դQ��e\�f{�$V_L��ж2���𧻓~Pc߯����=�6fS�È�GB���*3��f�0~Y{c��֐t�p�l��=��y��c'�P�p�F���o𥥦$:�]��3Y����8jM��`��2��,>=ʥ\=jQ<�w���v�\"�D ��2e�ۗ#GD=���K県��W4f6)�9`H�ō��Y��1�w�m�1"���	;���+G�ĕY��y�G�+�P���5�3�4�#�����l���aO�7@%7��x�3�ٸn򅡯�D8x�|��N�I@e�enbҖ��1�}���^�{�-�oһǒߑ��3ld���h*�Ӛ�oq������UK�ʂ��D��5�i���:9��_xf\��p�kZ���֙�Z���ӣe� �N�b���?Q;k���PSy���y�#��N�m�3���`��\kj�|�I��T��5 mE�lƬp�u�����רB�͚;>:P�˙�S������u}_:�zGG���FH?O�N��|,�\g�U��1��`E\�s}�j�O	>�T6\��\	i�V	 )nZ���\�W{Y3�6�d�zjp��S�>�)%�n�Tv��z�_�-&�G�����}��Ȍ�o狭�D������V�ێ�U��?z��v�l5��s57͢y54�0j�K���ݡ#���P����uӷ�U87f+j7���'�0|}���s�1��Ls�T��\10	P��H����1R0W]�S�3iϛ�V<�5����*�1��z8�Ϯ0c&��Xhk���l�,w�7����0�i?Ovw�x{���x�k�	𹗕�S�|14[E����Q�x�Q�Ch�
�:i�M�b/C��x�E�
�քX����Ρ����ҲB�7�-�r޲�5��,!��M)�LlK$��q�����%6���к���,+Bѓ���i��<B�6�_��d�?�$>B�����J����Ƙ�����%kNјw幷�hl�"�ρa*�Ӫ�X T%o'���T�1G��I���J6���r�����:f����,�rſR��p~%��X*�}:�`�h?ZL�Rh�G�蔀�εu~��EĐ����ن��Դa�%"�q��r9�jV&+������O$�au�$)�3th�!��;�U\<�d��w�^�� ����!�H:{��e?�;<����g����L�:�7�LV���H�іm�biڕ�[9��M��bԃ�i��_P�綂>�����q��p�^����1𴭰�Sʚ�O,2���^��o�?A�a��xoY�Ä]�z�)5�l70�\K�mT�V�����	;w��������ݣ��d�#�	V�st;�F�h"I*��A����Q�W�=ʚ(�n���s@���}��3�C����=�Bt��hj
����@K}w<�Bj(O\%N>�FWC �ؐ�_
Ů{oi���컼j�d��x�^W�WH��\V`$�}�v蘕�1�ng���]dQ`>	�����!�"rӾ����10^�v9����[��{K6��Z��4-s��0��q��i���乾��S����]a���.p�3L&����f=�*9�ث$	T�/r�Sk��DBت��ط�
���9�����@��r �������#���>�����s�qwĬ�>�P)�>����ZD�8��@xq�x^BV=aX�&Ċ��+@������k�kC�.�A�s/�t -y&(D�0&8�6W�8n� r!�s��������<vg�;�M�$��ټ�>������tLqJ�P�ӬB�1��M����.�/Y��'6�g���eګ�K?*w��͂	��4^�{U�'6�,sTMy4	��)���k����4�vU����ƐY���?�����MF���2��R�y�ۘގܖs��X s ��j�B�$O��Y2������'p` �m-�����ӵ�U�%h~���v��Kz���ٰ�?B�#�h��/��z)���h��S��W�,7}BǓO��i:Tc�M�3g|��s߽�N֏�˔��6�7�� ���iF*)ft�g�,A^L�.���.�>�*/����
ĥdfe�wj�[�3�>�!d��?Ei�Xd��uLb!�r`v(�}�j	��ۢw�Z[dn�M:b�6��뗈$n��,^�L {FPf�{-��6B��Ɗ63���H��g���3��1�[3��C���W�3���']�󞴉q�a7ε���"ɹ�S������˾4�]�Cu"�/@�.��7m�и�{���qO�Y��@���D�)e���7R��<��W���֬��m2�/��DC��
^���H8��gi�з�
)�VO��㕷Yb�~��{���XD�������P���/�u���j�ϙ����X4pyˬ=a��U�+6��X������M)�b(�	�R�R3�~ž�i��%��G�b���8��v&ԯ�K���5�9�!��Of�	!�Uvh@�#�U���;��"�u�8y~ ��V�Ç�oU����|�'<k&1�H/��0���T���G1��lxA�qZ�<�·]��/�s�4�N���K-���L	÷���<�$��#!���k��ۿm�����p�	Z�N�/���I�Z�Vz�Q�����`T�{v=���f�<;���;�H��\��h�I�5����}�k���τ�?J�����Ƣ�wqJ�v+X�N�v�U�Q��ݸ��������7J4aC���\2�j���4�����U1��'Ә����,_�(0�qpe2apt���-I���6�C*�)��3_��q�J��ڒCS]��!ܵK��GL!�@�c���z���/g�$X����uGKN}U�����-t\J�o%�k=f�B�X��}�b�qjI}.��Fԓ�{e%�e@�K{E�$��)D���ﰀAײ����S>�g��cƸ#��p-rN��Г��jxQ��K�@�?ٍ��+���wj��˱��i�}�sTf3�ǂZ���!�����R��*5޳�z����f��mK��#xcb��$�oߍaJ*R����8��,y��s����{�Z�����F�R>n��ҫK��H����zR���_��^��gՂ��d:����,=��Utmݕ���g�U�l:p�㝪��.tA-�f-�t?Q�1ֱ�²���.�t/��Ajm���w Ւj��T��P'κ�<����i���� (�jɎ ���ؠ�6�m�1s,KEO��6M�(p&M��캺�Lx\��,�ci c���򺐗?����℄�vG�P3�\��p��`�"�C3��,�|�������s�(��D8!g	`�
^���jǮ�6 ���n!-�M��6����2��Ow�G�O{��
�6�߃Q.��dU 6y6���H7�g�\��˴1C�V��YU���2�ܔ���]�W���U��56�QJ�"�d���q�ً���c?]LZW"� ;/�Ba.gj�7��¸q�&���/OF"��,1���D�}5eg��7m^�<�P�Z�'���Zl�* D��,�iu��I*��=�u�����_VJ�G��abst�)��Z� ��Ka�#��t���p���šșg7��s��p�f�=�k�����c'�9����^Y��}�����Rm�3�r=�YI������*ٖ[St�	��  �yR=����d�f���
��CŸ������ܑ񽘓0�|ycG�:��T�uQ.JN>T��BU
�#+g���yj�¾��K�pP�[�ST�5T��������"5=7˭Y`m�e��S�>�B>���,�d��-\�n�a�`k��ڛ��={Q��X�pBG�j�7-�a�{���������>��(��C[���k���K�d5�������Y����"c&��Ȣ� �����b�D���0��n|8��줮៹�&�J~���2<5<�������n�)%S��?Y���UaȄ.bi \��&S�@����̌ ��aX��v���jg5�Ʊ�Z ��qO"��Ksɕ�S#ZZ)�g{f���o\�b��0�"��u�O&4�V��D�|���L�to�?t*2�ԝ& �,pIn�K
��|tr<!�G�펂֧�I7���IE���A�:�Ȣ#"�$��gֻt��9i��̶�d20%U�t##(	r�/��u��4�ۻ�ր>���0ڂ�U#;���Ŧ!�W���nvk��L�!��d��X#���b�-�X�Ơ�O��C^��MR;7��Y� y:;ײ ��t�)�h�����Zr���l�]�v�&U]�@>C
2���{�Z���������C܋��:����>?}�#*�eP���oz{Ϙ�9Y�?���\�@��뀝��r�e���+�������*C���Y>����[!�e�Ë*ߞ�7 �V6���?o��9|��zW�(s�l�����L	u�msj?�L�DgEf���Ѓ9y��>�;L3������齛-��N�Ng��|^���j1��������ۦ2か����7�Qה9� k�8��<S�zI�x�էEǷh���N|.m 	�%,(�T����Z�H;��R�,2ϒ�ԭ�W�.���v� �+(�Z6���Oyl�Uil�	�(=�!?ͧu���-F��>2�8�NׁFE�B�J��:!�Y��YF{~T%J"Zʑto�'�՜ƈ�S�KD��C[ȍ\Q%O�F_�Zv@ h??8hBIrn��M�S���Ia�V�8̢&��"�BA����p�Y��IFÿK%��9EAo6Dr�B����SEcI�U��[K�5\�W���.�Z� ]հ?gUAh�(B	���[���b�Z��l_�5hqv�Ȧh]�� \���Y��W�Yi#�t�5"���k�-G��i�����O��_'լO��ms��� ¤=�^Eǲ�h�a��ޠ<
)�x �k�7�^�@������p�v��q׎���R�.��һ�"�:�K��$��ğ8v�rd[�%눪�a�L��d�q�[���P�H�ȏO�>���T&��Mg�?~|�<�b71_��,�*�����۝?Hb6�`o^z<n��AwK�lӵ*%����<�y4ۨ�9���@���ew@�M|RX�����}pQ�FV�'��ZC)��O�>4��X�9?W�~QXL{�e4�#t�I�^��+nh,t��` Ó�$�g����8��ْD�+N'��k	}A�<�����Fʦ8߄�]�}�P]j)��+�|}s[5�2�p���=������;`���� A��5��P/�C��c�nͷ/ع�)U �hW#1�jTpm�W�V/!zwO�8�i�Y4�~���]=w{F$�����ٹ��5�W 苳Q�
�\r�'����F�,)+�GX��w�b���ݬA��P��|��n���l����9m�K���Ǡ���ŋ�2�*���Z\��ѽ��`�m���2-�?��Z>�/G����9YX����_Ff6.��]�TN u��G���L��4���-�!$���R�T h��c�( �ūٺ�_5�8>{!S|f�c��bir'��Pm��Rtk��u�D���2;��uHZ�+ ���|E��p�M�aXhՔ��)�n½-2mn��9��H�b��~CVrW�74q�5��DEY�?���o0�0H��bg{S�VE�t��`����n��7��L������$@^Z/�a��Ju��7۔a2�(Nګ-����cwPQމx��Ό�J[��d�3;mc���d"L_���D�o(@�.G��vpO,+ �c;�����c�%t@/M=�=�~�K�p]9N��=*�aCF���4F�&/=���J��������\Fʲl=/`��P�{�f<$]g�E䯔�#VL�i+A7��:�����?s$߰��)ն��@��|�~&>���_=��6�p���[B��G����O�s~b c�ik��ƞ��r����qy�ɸ�,q�P��O��ܘ�p��*a���ؼ��Z*rj�}�I�2��[g7ԥb��j�dRwc"ev8C��= �= 2nk3�76�D�#��h������ � /�b�"n���X�G�Y,O�����;�1��7]���y�֏G�	�Y���z+�Ī���3m�4��T�Ձ˕:��rCp�'@�P��X�#3��ǸW����eDa��NI�@��NeF&�_/�1��К�{+o ��$y��_�����*'h������gW�+�
Kb��+���KU�H4*�hi9�Rx���4��J��}ԙ?	P��We�xN��Q�9���M�[e������+�V u��!N� ~3�t6`8�z���I����_+D V���u�Ƭ�(u
b�; ���~��C�t:�љ��w�vI�7��uMh�:���GBՆF�Q�OU����ݖ5�gؔXAV1����\;r�}��O�^�T��e���a.)����~�\u�$�������c}�Pz��)n)�n6�K�_a�z�a
��,�3Ͷ���{�ն���e��J��QF��1��S^U���BCݿ�|��"{K�5�h�B:1�V�j�\oK�Tc��d��I_��n��u4�f�8 �Xj@���P]�|�-I���ĺ@R�������$�E��	Y�LH�\�$��R�s���]�ixv)V�k5r�a�poZ�e���N�8$%c�я���ky��l�.
�v{׭�0��O�EFx(�v��kR��rܽ\�0|Zm�E�>(�px8x��r���
���i���k`}���1E���
Wb�]sj�T��Ƞ�{�һl�79a�仮`��Z�,��MM��5U$�{�q�ư����˺##4,����<2\�2����z2�?�W�D`��=�>�K�n�cJ��VӲ��K���kw���`Ƿ9M)�)�
�T�s�X��N%x5���ϭz����D�)5	i7(r�J���{:o!z9�ƭu��r.V�XB&~�ad�����Y�:����@xL!yF�q��	�ϵ�ч�:��%�ُ[��1aO�E"���t�9qq�&��J�X���O;Wva��l����3�B;��j;\�<ƒ��b@ӇE �˭�H��V�x7;�Q��n��k\L۟_��)VeNjH)��mU4��^��9�e)��?,���c3{�����?���M�:S�p{��~�Z�ϴ�,�S3�$��̎��p�W״�XHA�0����:h���w��`���b�%}�m=�hV&�]���"�c���@~�=�W��u�@�<cV�4�;)�hkp �>R��J�Q�&��nu(ދ��-S�C�.}�0ݾ������,ձ��BHa���^8
�[�i1n}��_B��RO�kvN粹W6��yT�
�Zko��<jw�%��dq��7W�a\?���6����n1:z �b8d�ag	*�K��e���3��z��/�1y��v�N�MI��SG��WLô߾=����2�h�M�菁B���gx�x��|�Z]j~�����&�Kx<�=~(Ǫ�^r	=4r�S*��1�M�b�^������M
�@�.r	E0�:C1���#�Ï��Z^�2�:��ĕ�����PR�n��SZ�+��qq��^�s=J�L&����T5��V;�ԓ�k�47꿢�s� �t霪&1�)Y4X8��$Wu7��;�!��sY<9��$Y�E�C�d95M0���o���ť�_wk})q3������Z�.M��68��U��'�o���̷ڴ��?S�p�Q�Z��4�)�U��)'԰�,\(<y=Z��Rv��f��g��4y$٢?�YK���F�H��<v����Fw�Aӻ�=R�qp�a�T�������s)k����S���H��2����۪�`	��-���Ρ���������>g�z�]�ٙ�{B��#�>��x�Fz���=��T� �HCB��ק�X�T�����B�v~q�,����f
���O�@�	 Ô�ibS_*�R��%�AA�.K�lfs�3O�W���iY\Ʈ�D�;����S.C;��D�;��g#��i���I'���PȌ��^ClPZ�����L@�TE�+�^q�P�t�u�h��M��Ap]m��1�������\���T�y�X~'��o�x�£�[�G�|2��=H[O��v�T%d��V^��8�8I�s���s�O���,@ؼT�۴䖬vAu� �^�[��]*��.�D�ڣ��"��W��D+��1�^��MC[p��4��PG��YY���d�0VU��w&x�����+"��p�Uқ�zJg⣩��Ǡ,�Ʌ#_J���W��5V��f_�I��kW�w<�i$'�k�q�Rl�7}�u�,_@7�dO|)��,��z9�8��6�l/�� ��}�dݣZq�Z�r'���9t�~�RV*����7>S��^���:T������ ���m�q?�͘$O{eZ�$�p����.�� e�,E������my�zJ͍[|�O� �u�A[%��閾����$5�H�6�z��� �+�������A�Ǚ����!�X���zqrb�����*y��f��E��.�\t�>L�)K=�`�s�߆�m��{g��|9�e.��B�x�@��e_���>��)��U{P�: cH��{��^�UkEL��O݈佲�x���#y�^�=W��ܛU���\�5';��&K�/�ڰ�o=��G]���a�
�`�<�6]~�/c44����7����	�^ʛ�&<.B-�����p�P���ۖA�+�V�	OX�N3�����Zz� 5��1n��_{�hU�����яS�E������I�h�5�)��F1��`�C�Z��ӋdUc�S��)SJ�ޕ+�Z�k|ǂ�f��jb�ʀ%�W��-(,J�ܯ�i\'�c�x�N�����*���JŜ2�f��*
b,��p��Qs�׶#L(C����$�lK��L�����p�i�}�/��,X+��x8aK������#��Sh\ͦ�%���f�PX���}υ��f�I��;��ߑ�9�%���ꎥ���}�,\������.��4l���J��c	v�q]Z-uh��3��}Q�n��!	�p��n�{[�$��8��wd}�-ifV	e����(֠����*�u�q�
���jf�P�KJ��x�їD{��aM=�^28l}vOQĕO��hlΝ��p!h勬dRdd��T�B&�q�˷��d(oR��L_��^ѻ�g8\��'@�>�N�,���[�Kt,���gM��l��H���C��A�2V��$t�[�45�����QZ�/nbAM�͆��ze���m�b[G�����������u�LM��N˱(j[�ɑ%��NŠj�gm�,�l�γ�6��c(�S M�&�$.;|h��)Nc����v��ӥ�Ǧ�A��/���R�P�
W���c�Yؔ��3�S������4��w�Գσ!���`4R����wjS�w��ܢ���n���MxC6����FM�2m��p�{D�2�9����R��'61B#[�H��g�n�1nW1F�M�%1+ٲ��U4��v��]�(��X�_˖�T�h"GEA������:��|�}]/^h"�l/>��.j�7���4�����O�����c�P�D���ej�B7�N�<څ��}g�Ȕ+i�V�m�7DA�X�l�o�e�,��M@��$ ��-��V�+W��bv
��}�������%��װWz}ϳ���h�˙j S�֤�p��/=Z���n�ũf�Ř��~("a�_��g�W8�R�i�3}���<؊����Ee��^�!�lT4 �>�R`�ڷm;%d�ϒ�b��8��F���9{�pK����#0e�yF�:���?�Q1�>��}פ��gG��yMWD����KS���"�'S�m�T��P()��+�	77�!`�5�r�S�I*��k�ͮdE�-?�n3G`Y���r��+�Q�}M��Uӛ�dF-�y>������`�^��耺K_�ƥ���hk���ܣ5��'ANw�Y�������ᓻǢ��``�e�h�xH���n����o��Ⴚ�&�gҳ���2?��`�x�ZƘn��S<v�"����'�ji)л�� @�.�-����D�ֹ�������Zc1M�42i"�e��!���Z���g�Ef�"^o�����p"��͇���4�#�Ӈo|��۝O�To\�t���H: V<�IQ��
]��|��!
7~�>�Q�����7�gI(焎4)"v%��J#zb$�:���_��8���0���w�\#��$���u��4xd����>ܭ�0}�cU&M��L�!K� ���k ��{f§8.��s���ǟא�nX�xT�r�ƌ� L�;z����ը|����u��8%)�y�hv�W�~P   7
  Z  �  r   �(  �1  58  v>  �D  K  �R  ,Y  m_  �e  �k  <r  x  �~  ^�   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl�&X��;O�{�'�jn�!3� ���ٻ�
��3Y�"`�j:.5Z͐�%F!5�̢�(w��p0��?U`���?MR�*\�!��y��F�]O�y��Z�LA6�ݻX��$����*�@� ,��냊�(���*��ea��)CN�!2EcR�b�L�ps��,���A�'���Ё#[�H�2��n�V����O��d�O���O�"��G��"H�J��UP���b��O�����%`D��By"�'�Hp
��O2�'~<��%kJ^�#�A[�>�q�P�'�2�'��'8�;b�'����O��I�{�
U(#�S /� Ҧ�� f`C�I�|��TO��}�N���(�F��O�I<Utȡ��?Ū��"�|�+�C��NȐ2	�O*�d�O���O���O8�D�|�w4cpd�5�Da[�͔�Z���;�v\��h|�V	oZ��dզ���4˛F+eӮ�ğ�����{E�%
�����UEz�ʅN�>Q�ӂ堰�7�J.�N�
�/�3�*�s@\�}r�<�	D�B�oZ7�Mñ�iA���O9�U�N r�
���,��"7D!���X#&d�3�`ӴA�"%���k[iv6���E��E�,@B��ߦ��ٴ-���.K�p��@i��T�n����p��4@���@��v�l�o�M��ׅ9VR���Ɵ%?0�X d�ե!�)���|V,�a`ɟ�<���9q��"k������2��.s��n��>O�$��$;�6�@!Dͨ
��T��&#V�010��$uǂ1[p�	��M�S�HRĸ:��0J_L=a7�N��?�2f��qt��C�I8$�<8 �*��.�B��O(�D[7*"ilk��<ႃ	D�:��!��d��?)O��$�O���z�8� -C�~���x+�ҟ�J��ޗ��)���P�g�t	[��.O�)�Ȕd��=[�m�	8�7��5R����m��j]T�1��@������M�2���O|�6�r�g,ͦ::=J1�9���	П<��f�S�Oޞ��vM
 a6B����U4}-�p���!�,
x��-�We vxxؖ�Ϛ�?	�����\�ݳ"!l0j�E�>��Pq�
AtTB�	;LNtL���ܹl:L�`F�1B<B�8Ic8�ɕH�F
,[ 6�B�ɮT@�x�ݝSN,��-xR
B�2+񐡀"ݾd�M��B��$)�&�J�A�j��<�R�&{����{��"~� Ò�j��p�3H�;K=���&�yƈ)�a3���@��`Spc��y�� =��k&��C��A)a�P>�y�il���ڨ6��<�U�@�yB��S���ӎ�4��|�T�ŧ�y'd9tL�e,"�8�R׎�2��d�+bO�|��٫|��[fiV��Y:m���`�'ަ�#�d�1L�5�	+Zi��'�$9�����_����D�=B1��'r�ɲ���}�h�S�ٮl	j��'	�hBF�|۞�qTkƚlCX�ϓzXu@�i���'���K7!�+c�PXň��R��]:�'�$޸U���'��)�62(Eb$�e���s��O�����?�p�`PF�<��<s��'�E�ׅ�
J�Y�d�X<�&l_�
�29�4� U>H� �ߧZ���a��dӓM���c��o���s�c�j�^͓!8O���s��ty��'��OQ>ŉ	K'��h��g�Q��f9�IB���㟔XKK>es�d��aV&�\ ���O��O�\�g�6JO1��v�IGa[�f�����Ѭ(Į��2D��c$�ۙ� �)%Hѿ~�^��*D��K�� �B�@��ٷT�E��+=D�ӓ�I��r}����."VI �:D� P�쇰;0��qQ*\T0Q3�:D�xzbb�	�>��֋"\�#T����$�r�f��?����@��ey��C�ve�G#Y���	�g�X�6��Y�*Y�J[\7�ު3������|����$���0CN
;�XR!�%@,��]���$!���&�T"1�zVг�'���y����+�����v
4��i<�>����IC�矬��˟�� ��.袸��*Dt���}x��Ɋ��W?DOb�&8jq9s"�(��dBܦy��4���|��'����B 2���9P\rԳq�F=K������xxn���O2���OJ�;�?!����4�݀ ���R5�ȗqZ��+���8-�ba
�'�(s�DU�.Ȱ-�w�V������x��U0,< ���~o1��]�2�������2?n)m�X,Ew&�{�ŉ��yb��O�����
?IlabB!���@��֔|��\��n7�(?��$�2T0$q��lw��5�Č��l�'y��'��l�y:��#���_���;O� d=r���s��yK8߼4���'}����SxRT�%�ĄU��q���=(%. ��&ŏTӆd`q���)�*T�ŎN�'R�����қ��'Q2�FJ]RRd���p`�Ca��'B��'$2��4��=y�8M+G*AqLhT5�_'TV��
�O5�wm�W���T$��I����'E剈\�j��޴�?����)Cg���Dۺ��0#�������6+���d�O��GE�nV�a�h #<Ɇ�I�(����d�?M:����m�V��S,A�x%�R-?QA�
��qRt��z�ܐ!AK�4����`�Mѕ��b�+@�jf�� H'*�Oȍn�/�H���)��N�.�P���& &�9U�6GfC䉃wQ��:T�ƛ�\�bu�A�D�"�?��S�����e8O��(:�Ȋ���4lZ����'�%Q��a�����OB��<��=2c��c� ��茁��+�?���O`�*���B����$�-@ODx!��þn�H���
�?#�\z�B��/�HJE�Ã`�
̀�����	;:�.���"�8�.\�aCR4H�8���O����6���*�<���E,8��l��i�Ǳ\�k+OD���	k̓Hގ�#�M&"\�� ��@��'���C�~I���?qDd��8�O|�a+��ÞGJ����ʜ:��ݺ0�4oZ�G@��'�"T�4%?I!˕�\��MJ �B�PC����J� ��8�,Vx��L,��.J2���#ХB���F|�^4SQb��zV�ݢG.�+@`��I2%`x��\:�8�+w��0��H5��O��d"���O��?�	:uONy����P�0���I�Q�e��;'`DI1	R�-O�c�B���zX%����O�ʓS�i�!���_"w���Ɗ�� m� �*�?�*Ov���O���	W�fC��J7P�p�1�-�)�M����6C�$�X�XK� �q7�A�T��ȁ���{�m��n��H)U`�'^Pm��O��M)B�8EL9ǔ}�r�	':�V���O�X.��L�/Vs0�0��G�JNU'���	X���; �ǲ?%���c�a^J��8�Or@�I�m.�@	g�.4�L�;�e�&:�&��<��N����):-�<�0h��C"�U�.�D��B%N.����O|	�Q�Y�t<��qf@)_�
`��t�O��z�� z{�×"h��m{�O�x�̊4U�BM�����i&x%B߸O:FP�Α5��tP!_*I�L�Od��4�'�b����<�URwH�j�.��De���ce�w�<� ��XQ*X�E��%�r�'�~�}⒨��iش�31J�q'zɳ�ă���<�&�������?����ّ	^�1��oC�IS%͚/M҄�aA%%����b�~E��� �3�	""� 0���
���4�[<;3*�#�Me��4mZ��|��a�~̧���'���F��a�fm KѮ1���x����V�]C��'�ў���H�I���R��59!�K�<AE�M� � � ��B4}A�,Py"�+�S��U�����5TzR�+P�G:M�CA:��U�I��,��쟤���O9Hxs��I.OD�)Ũ.T<���Z7.@\��Mt��eC%�4<O��R&�I� ���h'	A�j �as��Қw�F�	�N�P��0���r�DU�`�		4!��H��E�Z�v���&L&0U`Isfe�O<��!ړ�O�i�A��m�����|�TMpf"On,r5e�nwBU1*\�0�
��P�|�ţ>a�2F��� �-:d�b��:Y:x59��M�y¬̍�-*d�]�HE�B3�_��y���Nr	�"OE�ĳ [)�yb�_����"� ,	ݓ��T'�y�*��:����o�z="}�e����y�&��Q?���4� G���R0�hO�A��S�?<�GcUW긜��.�)
��C�I�*�� ���J&[��x `�zh�C�	�r���X�X������
��C�Ɏu�DY�#������+�"&�C�%�
EG��_���d��*�hC�I'TE�[���r
X-?Q.����"~R%ߥl��l��&<:,Xō���y��+`�P�z��W�l��ĀF��yr� �6>6܂`(����	��yBⁱx�x��(G'����〴�yR�͇G��	9t�>{�� ���'�y�hE�F�fL[ ���n�FaVD%���'}-�|���%�
����h�0�YF)��y
� "���^$/�(�1V�2��P"O�T�UB�F��p@��A	��P"O�(0�`�9 f�)�� ��!{�"O<� �%[�g�-��n�1c����'i	s�'��Y"&�.P�Yr&`Ӡ>�H�#�',Z
	>��b�v�b���MJ,�yB��<a�('W���hB"���y��U~=�d�2��X*���y���|h��ېe�9�$Q����y����r��Ŋ��{�"(�@dC�hO�P���&y�NX�,E?7~,��m+[�|C� N��Y�a-J 	��#�:=z
B�/[� ف1^�7��}���K�N��B�Ibw�%w��2Yݔ5c�f��[R�B�?_9���T"Q>�T�BtI
�}{PC��8l#V�k�m	-<���3UE�<=�>��
)'�"~Z��Ŗ'��$�� <X�Vha��6�yb��%t�p	�3g�FTaD��yB�X�����K `�����y�m+&���W���ܴ�0�S#�y���5rt�ɢ�ᇱ7���Y�yr��SV�݊i}��Eҵ�L�����:��|��k�~����n���L3�y�%��8�TI!m�6c}p����ɔ�y ��>4\�k��52K���)��y��)w��H�`��%�Z����y"#ۗIl������&��,�1n�,��>AƁBS?��L��v���r��{���a� b�<q�O�7!��� g�-vu��	c�ZF�<���Y�g�� ����`��I��A�<)di�<$H��q"L0̴����B�<����&FV��0��d��WlI�<�"�L'�6䅕F���҈�A�'��]3������В��]s$\c�
�#2�!�d�r�FBeH�8�z�R���7P�!򄎓I4Tp#h�3~&���ņ�nj!�d����H�h�%e�()=E!�d��[�^��%$[�:e�9`�-C�<6!���9
���jJ\a\��l*��N��O?AH�g��c�f����Lh�G��m�<a�9|n8�|'��"oAi�<A��K�4tx͙�9w�D�f��M�<� e�{�j��'K7k��PC�G�<��j߅W#b���o���$&HA�<��困S��" B�-)^9��gyB�W?�p>IdV�U�r8�B�C4��Zr��f�<Y�G�3���lI�VxI����Y�<)Ŀ_�cF�ՃK�ͺ��L�<9�JF�I����l?�i��
D�<��&Ƥ��@j  &ڶ�c�&[x�h�Eɹ��R�#�i��yUe�eW���d�,D� ȑi�1&�#�i��~��{U%D�<�C �*	���#��.T ���ċ/D�@;�p> -���Z @���&�-D���W�ժ&*1E��W (8�%*D��H�m��DU�AA��l�.9Zan"�vЬ�D�T�1<H���.�$i�
�,L��yb#fQx����r������yo���D�C6j�X��zCc���y2C:i�.4�5�JMzr��SY��y
�+� ܪ��1���c�@��'�`���۞\��b fY4-��@+�C�NFx��)O�,���B�*b�
�-�7^w2C�Ƀ$eV�aš� /�
�p��M+Eh,C�)� �����j�C��P�@c&IP�"O�A�`H#���v�pX.�s"O���O]:8�.�%��v�0"O�tIVEĺ	��D�T*T��l)£W�$9�,�O�<b �Ο�]��/X�ʼ�S"Op��O�g0$���+{�P���"O����I�LY��H�N^4=�B�
�"O^�����@&1h��P�C��mBw"O��g��[��K��pt�!�1�'���'���0\e}����V�~6�d#'�4D������	M�%���Ԉ)��1�(D�t�r���@��kT�/�8b�'D���tL��"0#&��5d߮�S��&D� :�朩 �����ԣ&Ԏ��0�0D�h�$;;k��!�R�\�l���!-�K%��E�tiۃtE�$�D0E��u�!/��y��ߏf(�E���p�.M��X�y2-J�<�&�B��J�j�(�q�O��y�愰aל��Ei�%fQ�Yk�I��y¢�x�l��Q�5��L�4���y�n@-]yzq����4�^93h
(�?)bH�X����t]��`^�B�2d��	��D�8���<D����(S��c"=d���:Ac?D��Q�G"3�,L���	� �;�h!D�h���6���Cb��4oi�];b�+D��[w��-#���)G�{t��@�(D�k��z
<���C�2�|�1�g�<��d8���6�R>
�x�����_�nijci?D���bN�a�Ҥ����#4�:RM0D�Lr�%żxH��K�.�JD F�.D�H�E�I�fi�`�ը�0�i��+D���):sizhJ�=\j��*5�+�Oj4���O�m��bXvS>���:B_@H"""O���F�D�g�d����>omĵU"O�4[SB	P�I�Ըk�4�t"O&���oӴ�48��
���i��"O��C&z�|���D����׋�y��Q, \�9j�8ِ5*����hO�U����	T`A�B�>>R�`���i� B�ɑh��qHb�"��ɪg��0<�B�	2��T������x�� I3ZB䉥S�x����<�~��!���C�+!u#�I� �l�8p�[+j^�C�I�E{�Ź�B �ZEs1&��veX���#t��"~&�G�A��(�&ϨT��dQ�ψ%�y�֒!��a �'H��`������y��̆!�کz$I�0DV��B� �y��ֺo��|P�C�r��bJ�yB�
5]	`��Dk?�t)GOY�y�+�Y� �Y��ZY��� �F������|bE��9<
0��������I���yE&.�
-r�ڈi�)�"���y"�K�i�ǣS�^|�4a�̃/�y�Q�RSLPa7�� [8=���A2�y"!Mw�|mӆĽO�ƴj0K����>�ǤOp?y�@��(x �G�ON@%�!)�g�<15��6Vr�:�햂X}8���IPx�<���@!(f��Ek8>����1�Z�<9�`Н^���3aJA�$�`��AMT�<��J��-rB鞴[l0��ff�P�<���H5|�Nɀ U�:@Ш��v�''�ۍ�I:X�v�
É�;�� �0ꑧ�!�$����I�z���j��B7w��1�'�q��92��X�A��n(E���� 
	kC�\.*\^}�����o���br"O�Z�����\!��i���"O| �c��/���I�<XpZ}�B�'Ũ� ���/�5q!�1+x��)�->��L�ȓ=�`�%g2	Rp� �c�e�$�ȓ W.���6_E��#g+�*F�؆ȓH/.�' �T�X�R"�
U����~U=b���\b��J=z�d��ȓ$T�I��$�������7]�F1�'m�I!�V,2mX�K����`w�Դ]��ȓ��ĀV��(���[c��5砐��^�i��.m."|K�fC�>��d��D��u�T(���A��V`%�ȓ4*�@SB��2�����gT��	���I)n��q@�U�&Y�TV��l��C䉹 h��q��M�4�H�*�[��B�	�D��`rW�,�X��!�$ UB�ɲA����fA�1����Ro͆Y��C�ɤGX����|t�h��&JQ�C�	��f�3�A��u�����Ԣ=�t�U�O�d�@@��
�:@��(ɮ"��j
�'ȼJ�K�3q�^i���{>Ա�	�'Ҩm���;R��[��#;����'�BY��"--H�Y�ڳM��	
�'yJ�����9�ޅ1׆�8B` %r�'�����d���g�̬Y��~@mGx��I �V�jm*WiZ�c��p�Μ(*�B��5V;���B���*EcP�-�C��9A��#�J�HI0Pq�LT�|B�� QgPD�0��
��Ha���5r2C�ɐ�P��یy��i�a�P�C��"(!�h�P�ǥy�t����
	����Y��yy���:1(c�,)c��#&��ј���!e�N��%���d�O����Oj����^q+��U�%�d��i>i�2OߨX0=�&OW�?�~���$2�e?Mb��4�t}C2�^��MC���"}��t"I	�xYdEs� �W��������Nc2�'�1�H���F�3:�&��S@� ~�@`W������DQ[�/��B�"��qL��A����NRyBgץxP-Q�ꈓQ�m��cS��D܋_|D�o��ؖ'�����I�W� ���Y�\!�r��U<g���	�' pѳ�2D��Qz%o�;�?E�D*G�X�����'5O��`�Iޮ�y��W�
2R�*�B��D�<I�0�i�����鏴5?A
&��}mdP"����@�$Ф`���'��)��9?yD�aM���`�(PU���j��-C!�޺5�ZX���Ӵ2❋����ў�y�����#����P�B�y���t�����<1 ����?!��?!����ԟx��n�L.D�zF�P=��%�򮋛}�x�Dβ]��m��R���3���}�o�;f
�@��(�2����S,�M��)|w��+�$� ���S��'g��"�]1AU�xKV�
W
���O�D��'���	�<1���qx��Z�Γ6c�Y5��g�<�qEʉpLB1+��D3C�
�P��O�`��4�����<�bɄ���9y�FNi��*�`I���2���?����?�)O1�@(*$��9Qn@���.A��UH�&W,g��A� ͸ ds���\x� �C& �8 ��q
�>*�V��U�qst���@�g��i��¦�"`I!�P�ɳf�� c�R:cJA��ƐC4`���E�'��J�h�0*B��$j|F�ۦI?D�{Yyl�ѡă�'I*����^���d��M�	Ky�k�5j�7�M�P�S�~�����XN���pL�,P\��'M"�'�"�\Ix�1'B�N�����O�)\'}��+�愳g�(MS��\8����J�qwHZ�_#��mZ�p%n��ƃrb��	��8f:�B��RF�'�~p`���?q��Aʖ$x�Ó)�4$�Nt���d/�O�C �`�R���� Ӷ�`#�',H˓%�T�2K�ko�$g�D�D[��'�����,|ӆ�!�a�<�)�X�I�O��h<萍qC��vK�E�O����) �Fij6��g����)��|`��B.i�`�R`[/������@�U	�16� a�T(S2�M3�$�[�O��t���-Lw`�T#���П'�v����?��O�OD�)� ����I�&Av ����D�@T��"O���A�!m
��ŀOuD����ȟ�P����/�(�*�/�5����Ǻawd˓Q�zQX��i��4�'t"[����H0���,A.+�( �fT�/�6|�C"��?)0�̹'	��o�n���	cȐ�	&M�i�
0W��'�X�ye�e�2����UP��-�E:ҡ"4�)r�^��
"p*PҊ��i�N�G�P���� �Ik����T	�)>�������*.fH����yB�8D�xtq��W�JD��g r����HO���O�c�`��_�	\�`Ib��vvԥyk�O�a7�' ����$F������a�����'���	4�ť�h99u�I5i��d��'�t1�BK� P
q4e�a����'�l<��茈1�thk�bD�faFI	�'�HR��4�"���i�\���)����#P��n�����	�|*1ƒ?	{�)W�L?a���G�L�<Y�Șҟ��I�ic�"w���(vE�!a�"����|2�:u�J���N5�J�y�cEs�'�h��� g��iEC��F�X-[�栋�JG,>�:�BG/�8g� #1�I�t���d�O����O��22��X��]�`Y�eA�ĉ�dj���O��"~�/�,ʢI؇KKp���7ƀ��$7�S�ԁ�<�� �-8���A�y�XkЅ�oyR�'��5s��'5�O�r����g:��,:�,�H�`�f&O��=��Zy�p)Pbfە��h��Op��O�U&�T�f�'��Ӡ<��� �, �9�8�c����AZE��4�?�3�'�y�H+�?Y�������y�	��C঩�f���v��� 7i�f�a���i�"�^^��<O$ASҟ�^wИ��s(�����5�� ��.q!�T�'��w���o���Iן ��⟀̓��m�	�fQ����O�b�@ٟ��ɖ^�<��	�<	�%�pnz�r����sc���tu����4/u�B��'3�9���?�R�k?�ޟ(���?��ɘ�.��FZR��e@aj,ƄЩ��Mi����ҟ����ݟ�̓P������]��u�φr{:`�"��	��HW*
�M[�'�T�0���?Q��[���'�R�Oh�q�'���r�q:G�A `E��ߵ	��D�%s���'���]��͓1�<�禍:� �?�1Ԥ\:(�T��de�> �� �4�y"E�ϛ�Cf�| ���?����?�!0�чF�� PV�������Ǖ�M��Ц�y����?!��Z���y��Z��ԨC V:���h�8���򵨖�Iy�6N�\�W� �	�b>�I�Y�Ŧ	'Da9�oָ����ȓ:��0�� [��h*D*#$�l�'q��IyB�'�U�P��&�\�`�nU�-�j�p,�I.%!�4�?Q����D	Q����i�ΐ(!>�>aCj�Lf�i����3�S��&�P֌���@�|st�+�/��y��
2R�Е�ټw �ջ�MǱ�y���7���{��V~�af�;�yr퀿X���J-|�h8��Љ�y��ˈ0ٱF�Ǥv�����H�)�y"��+ �̵ѩ�^���fؘ�y2A��4U��gM���xFL��y��"�yr�_ 
�PxN��y�Вs�jA�f��G�(���j��y2�V(t�A��햀S�z������'=�"=���d"wb��"���w.�A@X�"O@���ӭR�%�Ń�71�Q��D i4!p��J�R-�fLT[����GBKR ��i��8ǆ�BuO�9S���p��@^��+3�[/Z�,ȓ��A��@l���V%�I�'o�&��Mj��H�&�f-�f!��r�x�8����e��y��b
*܋�Րԕ�e�Q�+�v��5��F���OԬ��Կ��)A�S�(k�!�G"O.ab�>=�� h��w�H·"On�($�X�p����fIY\�c�"O��0�hYj�&���ŭ_(�S�"O�,�EBƓ�6�H$��-`�xx�"O�pk�FO�9��1�"�V7+�N,u"O�˄�]~�ؠ�6ff~��E"O����1k��yC�	�%|&��3"O̐R���)w1DM�%�==��R"O�1�NQ�Zp��RFC@���"O�P�C�"��i�4�N/뀍3"O,�K���([��t;T$�V��1
�"OFT�i��]r!FT�z���"O� ΁�� �/Z,���� Jd��"O�Ir�-]1&�����B"O�e��*�a#�K�D�:��8x@"OXt�nX(H.,c3�Њ<����"O��q%h�d5��ygJ�BSFt#q"O��#���aж Q�N�_ti
�"O=�����k�-2MPe "O�� �C�I(��Cg�Jj	J`"OԌ����%>:=�e��&3�A�"O
��U�{���R��нl9`�҆"O4��0ؕge����; .��y3"O<�GM�37�L���,X��;�"O8�Ȕ�����r#�5H���"O" �-N9|���)�a�K�Ndʀ"O^� �i@<�q���@
{� ���"O�̡���+8踴����QЦ��u"O���S"M�q��IS�S�Ga����"O�z�l��bZŐ�c��XO|̙�"O��c2Fjr(E*3	D>'&0��"OЁ�S�9z6�(A��N
 c�"OĤ�uc�7���*Tƙ�^"���v"OL� �`�8��#����Bp�"O2�C�ԕh�	�D	�5.��]�T"O*}�@�*oF�����^޴e��"Od	�W�B_8:uqe�\ G"�0{S"O��֢��n�H1!�"=Q�"O������^��d�ՠNB��Rw"O�ب��65i�Y��M-c�|
4"O<��%L-�l傳�v�h�r%"O�	Pĩ]�?v��R��1(���"O��ӣ 7&y,4�&��?����"O^��"C�&���pc�<h�AP"O��s��7sM.`ׯ߄6/Dy+w"O" ��f߻�8�0Ձ�=t�`X�"O��BE�pP�������o���8V"O(�`��Vg����Ɔ�s��Y�U"O��2}�	r���3��!85"O�P�jHh�hB�6~:��"O:(���(za��H�ɇ	rkdY��"Oƨ3�LO�9�4�`UhG�qp���"O����e��|y;"�^Tuc�"O� [d�+S�V!��H�r�2=�a"O�@�&��&oFa�qg8o��1��"O�Yd��!��4s`��3\d�|�"O�������z��A��I'~|ha"OT��U�/Yqr�Yg�˶_(�3"O�|��ēvN&=*d�[**r�"O]�%G��_Vmj։�" �T��"O�����>t�4$	G�h�r�"O����ijdp��jƒW٠=�D"O�P�>�X��I��i�w"O@��J!rO��nw2�"O|p����`��њ��WaJ]�"OL��dךa&�ȢgK�<F�x)"O.����Ǉ=J4��e׽Qb(�'"O��!U�������$�t)��"OZ�!�J�PD�*e���v�"O���P
� ��p� ��|"s"O�� �cڵ5��T�v٧Y� ��"O6��V�A������-[��X"O������_� `����=�l9�"O�e�F'Ӎ�>%�A��*\�dő�"O4(��\�=X�P�$�B�8�"O>�q3�P
���jV��P���8�"O� ������MS(԰3��0�&�
�"O�,a��8 ���Ł<<��C�"O�e��e�F%0��Kl�|qje.�k�<y�G��P�h��)� ��!��c�<��G:���c�?2��g��_�<Yө�n ��&C�t}��QW�<����{�H2��Z��e��#	W�<���D|.-��Iː�V��)O�<&%��[tBhsDM��"c>��.M�<���y}�E��'������J�<��C	���9�Q�9��H�A�E�<���އa��f�:/D� ��\@�<Y�H�tgX\�Բqa��a�Xv�<��h�"&U�ӷ�4p'�T�J�r�<Q�Gx�1�Ԭǅ.m�tˆr�<��e��/v���l��z��7a^�y" ֞6�z��W�8CZ��bTͫ�yr��$t�9Z���@�SW$��y�J�Q��=�' ��ly�e	7ǖ�y҈�=6y�T�4��j �KL��y")�O�e��Ț�v
L���ϴ�y�'	�TK#�Àr:�U���*�y���4=��9qbk�)�n�i4c^��ybɘ*-k(4˰�׻z��Z���4�y2�ֳmQ&�7>+~�q�R��y�*˿Y���p�Ո0�=���]$�yMe1���5�ۻ,��Ca�ʼ�yR\�xb%.K�VcF���ޝ�y��_(����!($��B�䘳�y���N;��Ȋ"�6y^>���ȓ� �c�%��ҢЫ142�|��D�܀0��ƛ1��;�%B�*��e�ȓo|��T�pe�ȱC/�"#�����|�F�pp�Z,c�)t�R�1��Ѕȓ��۰�W6(,q�ܶ:���ȓz���d�{�rE���ޚ]0ꍅȓ>�L��w�K7>[|h����~2��ȓX�����9>��Q�VF�h���#-na��"'w���#B�[j*Յ�C۪ �G㢉{B'�#�@��"���;�8�9��r��@��Ic,��2̛�N����+�G���ȓ9�`Ö�5z�0�E�-.��ȓ5����C-YJ|��6&�y�`؅ȓea�t�4�`����f�z�\@�ȓC�\�C�!�,���թ�? b�(��~V
��(.���T�ۄ_b�i�� 3:�@��J�k��Q��'�>=lFM��)�遠H�?<��(  ��4;����\{�m���%��!(i.,��x����u+O�9�8	*��&6�\�ȓm*�h�+�h�%'�C�`�ȓF�B�S �>m �S�E�%��d�Tչ���>��@j5NSV�a�ȓ	��@2G#֯A0Zp3E�ȲT񺠅�4j�Л����<HjX;�n�-%$��q�pX�)�r���"łħUY ��ȓ+���$��7KbphKaK%g�襆ʓ&O�ca�\)$�f}1��ޚp8C��"D�i�P�YE���`��C�I�Rpx���G�[:HC�	���d�=r\5�c+�+l�NC��:E!�l���D�0�*�$�X�1�2C��-r>ށ���9��Z!Ζ6"�B�)� �u07dLV��\)qgX�c�����"O4%y� �,f7���5�AC�挙�"O���U�Mbi���ˏ��e��"Oh-�q�]�s�؁!�(`��
�"OX��Q��&k��x���>K�"Q"O�l�6��:n#�E����/)��"O���Ӥ�咀̖7�d�25"O�X36�����	�1iZ���"O*�{��
�F���R<.Pę��"O:��p�.��X��9IDh	�W"O�@�ݱT�D�#"τ0B=ڸ��"O�A8�� Py ���#�=��p"O>��EK�r���dd�:dݣ�"O�
V��#}�&A�A��$"O���p##��X#CO y��02�"OF ���/lɹG"���8��"OV��SǘU�@UÔ�M
!���"Oʴ"����>�ZEnQ��!��"Om���y�� �AS)m�*��"O�@�d� a}����F�}qP�{ "O��z�`��:Z1�1�4jq��R�"O�9��^� ���)�,�z^`S�"O���@o��)��8&�,"t1k"O\	jQb4v���t��)Z����"OtQ��F�Oz`���
/(��XD"O ̠U�ך(� 3���1����"O TaQ)<��@$ͨ��0�"O�|�S��3rL���	��a2@"O�m�'���h8�5p�˞<Urp1�#"O�ei��\?5Lf|�e�/6f�1�"OH�6����|C��dY�M��'�vU)"�1Ҷ� ���{�� ;�'��Ms�#��0����&As�� ��'DL0!��8AF���+�B� ���'�6!��Oƻ�:��f49�b�'��I�蕏!jLcG�S^�):�'����9?8������!g�4�P�'��0�g����A���U�+�''&��n@�_IV�"R��#V-��(�'<*��w�� {3:Y��풛U���C�']@�s�C��(�6�6EU6Na��'(����FFC7���f]!t�hr�'ӌ�8a��J��h��e�@�~=�
�'�$�r��"���SQ�/$��	�'ǜ�� �r�0<q��:l�L��	�'{H6��F^�I����Y0
(��'
B<J ��J�:%n�%O);�'���D�t)��J�p:4c�'�t�HGON���;Q&�2V�\I�'3�jJh$�@��(~Bt��'���P�n[8efPiVn��#ߺ�'\.�hd�"�
3 G��t{	�'D��B� E�r�x�%d���!{	�'8lE0�h��Ś��ɨh�U+	�'Q
D���M�@L��	�d�s�'�����6p�b�8i�C�'���0g� ���HI�w���"�{� �+f�����)k�� �4jO����6E��{�>�q nƦMX>E��\�$��#5D��<�2M�+w�`��X�80B1᜘J~�"�� +)�B���y|.L��D!f����R��C�`�� � L�Si�8/�T�p��QU�؄ȓp���	2Q/:�����BZJ�	�ȓ"
�#6ϊ(����N�t��S�? 4�(��M�{����A��U~���"O�x�BCXt@ x4JLZdH[a"O*�PkV�1鵧�Z娄�"O�{�K�N�r S���<�jU�"O��"pcԪL�`-�E��F��12�"O=(�#��r���%�\�'��!k�"O�ZB���6��< ���4)��<@`"OdHJ�%�!z���Q8;*u�s"O����ʦ;t���/8&�)��"O��9���rjVe��4��p��"O��Ig+�Z�48�րj��ٳ"O�л1�S�v^SGB�'�8�%"O�X"EI
[L�P����|���"O8�ru"A'�4���ړeX�"O�Q9 ɕ6Auz��4	F7�ԃ"O>T��<�<x���Ҵ>0܁+�"O��@�������+�� ��:p"On ���»	�V��D�V�<ة�"O��Afޣ:�B�`�B�"����"O@}�Rƌ�,�l�xD�˰HƩ�"O¥��ȳ0A���E��f�p�"Oj�3����^2���t�J��!�"OF<�B�ۡL:��1A�2��D��"Oz��w��L��\��6�B�Ip"O��,8$T�0�J�8X�����"O��ba�6���ȓ�=Ϯ���"O�HvɆ�*��I���Z-�*���"O�d8��ѯ~��
⁚������"O<�eJ
���)��,����"OMq���A:B�i�+�D4u@�"OX��$4K Y%��8�HA��"O�(���.�4c_�mS\��A"O�Л&LBx����G$]�6�@�Z�"O~� BH�
�tʵ���F
$)�"O�8��$ӯ~ۄ@��0y�5�"O<��c��<w�| �C�� �i��"O�1�.��OA4L�RA�5�*U�"OF��s��)Kv��@^�h���"�"O�հ���"ك�mg^y� "O�<����jn�y7��3I�QR�"O�<ZфA�C�> ��!Ɠ�F�P�"O�u"r�U4��< ��
=�4$�"O�	��G�;���g%����e"Or$�s�%�d�j���!n���Z "O�( $�3Y@�K�b��oĚ)۰"O|A����[��	k��F }&~�HC"O�ن��#"Phy�Go@�BkP"O�� �lY�B	�
"O��2{� �"O���@.J���.�����"O�x�S��� ��y⁤?1!jay�"O4�p@�P�D*,���G�bcq"Ob@ABb�G6Z�rhف<���4"Oޑcw�Jr ���W<�P[�"O��҄�F��Z%�
D!�l1"OX��E��}
��',��S�"OP��+
�b�[ �R���"O(�x6HM�>-��ȥ��~�.��w"O`5���ۘ~x�P��� ���$"O���5f��0��5�p�Њ�*��"O�qCo�1@O��^���6"O4���T�[����� e�HY�"O2Ũ�L��pvl��	�1�(�!� �jx�!�I���!��.S�~�!��6�T	ӣ�K>to���t.A�~!�� Lqv��n���c�k
�5� q#�"O��9Q)�s���X=(� �!�"O�)��oZ�=tzl��$��bY9�"O���͛0(G� �aM
�`���"O:|�6lS$w*���G���{�(y��"O�ܛV���[�ͪ�H����"O ���a\�R�x����5,�H��"OZi���^�t�V������s�\)�""O����&R=QqW�G��Y�"Ox����c480!��U#�8�f"Ot]�gU���{���.�(!�5"O������,=�r���R	^圅Q�"O��Yp,��f8F�#a��Q<��0F"OR��Sb�El ��!Һ_#��b"O�t���̔2k��Ӈ��S����"O"��ꑢZ��EI1AЬm��Y(�"O\��R��ed�$@<Q��xAp"O:�U�;=���uL_���`�"O�h�F/�6*�r���ٸ)�z���"O��Z!�BX�����3<�X5�b"O�ə��G�]@ťO�=��H�E"O������ў1��E�&7lƔs "Oj��Dʏ,^���#E�tFR��"O���Ki��.F��U۲"O��30L<�A9�׬�܅ �"OnA3��ň36���Gc�!�
��`"Od1�)��WݤԂ"���b����"Ol�3�N�4��1;@�K=���j#"O8���>h0�yPQ`@<�$P�"OT��- <]���V��@"O=��.W4�\"6f̖yd�"O��D�Kb���N�28�q��"O� K�`��P�( �s����DA�؟H��I��.#���i^D�:�%ԁ��5��'%��0����{�Z)j%a���(����Y���p�&�26��;e(��Y,�!`A��j�<B�Ɋy+�#�JG�A��� #BN.TR`7m7!$^�
3��?V�D�S��M�w�C�F�|DR��W!0.z,��J\k�<��
N��p]k��H��0Q�	^}��J+�򁒀&��:��x��Q�&��Li���w&]�w��0>�7ႜoI��G�q�RlzA��#�Buۂ&��]]�X�&Ն��?�F�C L�x��!��|[6���I�'���3��� ����KTWx�O����ڴ#g�ԛ��[d��@��'��M�B-uʼh6��O�qђ�Ȥh4��P�ě� �h�p��h��$^�v�}��0M;~=�� 
?!���1P��@�G�)����T??�`��,4�pE�6H��>�L����ϨOv}:$#Շf��Yx6f�6$l�� ��'O�Mӂ��T���p@2!W�{ 5ӄ8����Ln� vA�G��~"˅�iv�C G�W����X���'��x��WΦH�AU \^�p�~���K4�.�*����e�a���w�<�eI
�Jq�B�˟iLܡ���і�r���l������:;�J G�T�O��Z���+LO����3[R�9�1"O|:- �-X7@��_Ũ�j���3Qr!F���5�Y�Q��&��<�`D�#���=~a��K�!	�<���,ut�2 ���@A��)��Y1l�����x�Qb&MY�<��q���h��XXԆ����#���Q��1sq�'��&�������O��<��OX}#�O/��$ѷj��e�'�&^���'�D���W�B��ັ�� �l!�O:��ǭe���hi��~r�LM�AQN�؄XE���y�MO:0��͇�%��mh�	��MY��Xl��.C���'�X=:��VZ�xXF�W6\s��#��=b�`���99S i��)V�'xP��
Ԍba���7�f���"��W�4��V*Ž+#$��'�7�"�~DK�@_()%q��-���5�*QW�B]*z��g"O� �-����yYh ��8P&�OT���R;@h��&��}�ԣ�X��1���($�5Q#�	f�<� �ߒIIDH�l���MA�eC���$��jra؀
;<OX�ha+P"Q���Z��h����'������V�M	f����!�� �Vg6J��B�		H�����"VF��pl�8w��B�	�b�h� ;?�ȥy�eՉv�B�ɴ?h����$*G������9bg�C䉓#�b��c�� @��9��N�x��C�	*S*��3J�,2^�����Up�C䉈x��)�qk�"l��逫�m�C�Ɇ�B;s���OH�Q�E�;"�C��G]�qg��v}��0+�5/�\C�	���d��+ �x �!�͋?�B�	EO|���*.��I�X�C�ɤl��	�����T�X����W%BLnB�I�z}�%sC������g��+�B�ɺ$�hq�W+Fy�L�� R�[tC��6n�&仧E���JՉT���~*�C�I&!�4a"�ǆ4�4Yh�j�8M �C�	�Kk�E�ś6��D+q��l��C��3#����r���|�͍${|B�ɵ^'z�1T��*#?*Q*���HB�	d����'Udiq&cɒ��C��/
l�%���M��*�����9I]�C�	�BK�!SO]�/\29z�A�pG�C�I�U	��c`n��]'i���s[C�	�r@h�F�8!�u�S��^��B�(:"��%`��IR�h�%@��C�ɝA���s�+�kJ@,Aw)�6Hk�C䉡p5̑����R�F�\>�C�I�!���pϑ'\x�-*��	-��B�	:)U�   ��@;���ƈ�q�B�?=����A�R{if�CW�F<rC�	�*�xܢ�D�'N�T��Y0�2C�I�U`8���/M�c����;6"C�I�hZV�q��]�E�bYY��EJ
C�	�+Ը�TjJ�x�p�+C�[�K��B�*l�P����U��XE�
hlB�� \�,��%m��=
���FV`B�	;#�^��4�W�Qy��҈{�&B��3I����Ԕ#W�IP��  �B�	�`n&�㵌J; ��@Bf��B�	Dt��# FӔ�^�Hā(K>xC�	1+�h6�R�5����f�"�B�{DR\����дp"�F�lC��8I`	���J���h #�̩za C�I�W
��XD0�ȰKr@J�lZ�C�	�f���H�cD�L�f̓!�(ZݼC�	�Y��D���3'��j���\B�	�̫B��)`���BB vB�30�#���J�-���h�C��#�`� ��(�|�dʇ4��C�9����V���"�VE�5�jB�	�@):h��ĈA�r���@A2Il�B䉈aB�蠅�s��I�2K�oZ�B�Ir�����gN=}`1�����
�hC�I�h�����
�
@�+J�2C�	pO\���
����T�H�U�B�I*��h!$$�Iqԍ��1D��B�IU$Q��a��!�DB��O��d#��ͷ/�J�� �0-~
U
9�DXyѢ��6�֔7��� kƷ �!�d�&d)��@RI�XZ������!��K�m�|��'%E	M9�SSh �T!�� ��%�$��ղg%� :mpI�"O5��ǼJZ,�֭,]bR�"OX�'�	?��L@0_H��V"O�9Ʀ�7�N��
��%.�ə�"O��X�l�1y�Bx�ŊŁ0���{"O20apM1H�بke�7<����"O�  �"T�Zj� O�!s"O���tO�X�r���� -��E"OMkv���6�15N
�l�0=��"O>�H2�E.?ɦ��1H�>{x���']ޱ��% �p9��V�2C���	�' By�rO����(sɟ�}Ī�R�'�4
���R?�����֒`b���'��������2���Pr&P1M�n���'���{'�\Hڝ� �JJnI��'�H0'�M�%֦���Ɣd�c�'�V5
��8P�c2�H��Ͳ
�'~���G�+?���K�d���Z���'�ȴꅄ���ݡ�h�� ��':��q�X�1;�}� m-_t;�'(`�V�)z⑌U)���'���L�PF�X T�U�Gj���'��R�+]4Yy|��scvf�[�'��:CC��#^`�R�ƍ[��8��'gn�q�(ٿr��K�F҂W��
�'S�(����6d��1[�H"d`�'���j�Z�����v��0(��'�*4��o
ryЇKO�K��a�'k$t0�'�>Ph$�LXv���'�X0��ti�� �˗e޽��'Jl���`��f
�}f���'�l�f�D�P �a���W<r/�5c�'J�}�A���b�T����(p_��c	�'�.Hk�
[�_h,�+��&c�L�'~��ӭ�4Pt麤�^^b���'W�zW�<`mR$z$%.S�Z�'��P��¾jX�	t)O?f��#�'��;�G$ p����X��'�vh*�$ƀ6�����ފ@� C�ɴ�v1:�#�Y�lA�k���
B�ɟ8��������=0��Կ%T�C�	7,xYB�%ڋ'�,p�o!GC��&~Ej��e#S�4u�4*L<W�BC��/�nYj��|��9K�"��
�C������&KȞg۰�1�%�7]|�B䉀Ю<0$��#�x�q�S�B�	�,H�J3e�3�J�i���H��C�ɩU�R��pmC,/l���רB��C��f���)� 3���+��U�w�C�I�+���F�(Δ����G�@B�	8c����������PG	�� �ZC�	e�0Ya��#@ƒA"Q��u�C�
e��%i"�ԃ'F\�Pb� S�DB��3m;��Bd|$QQ�c��G0B�,mENݩ��Q�R�=."�z1"OZG�ѐD�䔳
�1<�yp&"O"���ÕM�-���в`u�tz�"O,���đ	q@��	���1~���"Oz�B!�> W�!je`4����S"O�x�Ѯ��= �4�o�6X�Z1�2"O��ѱfF�R��h�7L��0�"O�ب"�X9�.-��Y�:����B"OZM�cB��&�ȇ��Z���f"O��p�Ӌ���3Ai�)V0t�1"O� �<�h�?c�dٺ��Ƀ	(.��"O�UH��W �Ƅ(e���m&�QCW"O4uQ�H�Gˆ܁���=�Z�"OAB�k*9�2H��Sꔱ#"OXTZ�E�&c���H蒷.�j`�"OH`1��z��L�'�G�%nܕ��"OfĹV�ú5���å�Z&�2�� "O�L���mW��6�� �h���"O��@� }9���!�.+��b"O�,�eoJ3u+�-A�AB�Y�a�"OxԨ���9T¸����l��"O��k�mѡi�0��ŏ!f�%��"ON�[v��\~mU�І�!�"O�I�B�4<dh���k(��)�"O�����N�=�^�+�LN���I�R"O���$+Pr�|�Q�GP���5"O�l8`��ƊBt�����"O�*��B�Zz0�	'HĢ"���"On�B��
�`���iS��.�,-�0"O�I�͎!@j�)��EƸ	TPá"OP�b�Ķoj�xR�\>&��Zf"O\�0A��e��]�F��#��t��"O&�@c�N%l��`p�-�7z8��V"O����zJ<���{~]��"O\  1��% ���3���q� x5"O|���EP:"���RĆ�*x�f��"O��P��B�M�D+�+	�yz�<��"OV���홨e��M���+�x���"O�� /e�^�*Á�vvR��"O q)'��6s4py��ߘDt�J�"O����Ɉ�8�ԘY��?v}����"O�ȴ��UP�K��ǺGrLH�"O�RN�.#�F��ƌξg�8�"Ohd��c��[0�k4�^9J� ��"O�4ȕG0m,]���&j�$�"O
Pg���� 7�>M��"O��pH�ivi���ф_I(X�"OlTs�+ɪ��)Jd�M��(�"O�	 0���}��c��-a*l!�"O��Y��#DtͩDDO�DVm��"O���A"
��Ѣ��8E��"O�c��`���+A%I�P�4"Ol|8��L�£��u�8��a"O��J�":`s��5�>�C5"O�E��%�-fF��pCAY{<q� "O��%���=YG��,��4��"Ob�s�F�b��4�N�Bt%�T"O:i×��"�,)Qubߺh�h�1"Ox�+W��50��\Q��5H�S�"OTݘ�Ǐ�	Z �Z�H��s� U"OXȠ�ƷF�$�J��"�<��"O�U�r��W�ځ�#,�#�<�z3"On#1��IBf]#���!1���Y6"Ol8��)��6*|9��\�T�&|��"O�ij7�G	�-�lJ6���XS"O�=�'��?�ȀJ��kr�l��"O�E����$iМkD� ([������ |O�`g̀�PEl�Z��V ���"Olp�CMG�c���*7���0����f"O���r�Ղlx�5	!��l!03"O�A9%�_�3��U���γ�ͫa"OL�ч$��>�z�S�'̓P��4*$"Or]x$�|vPd:F��3/8Y�"OB�`! �%e�UXӄ�+X�X�3"O� ����_O�1A�O�3�6	c"O�ѡ� ����C���:�"O���jS�*��!+�oD�y�n��"O��0ƅ��n�@��q�P/c��|�@"O�!c��o�F����ʡ`f�y��"O�%b��?| �iw��;���C"O�!p�ň&�8T(Cּl޲5�&"O�I�P[�f�~Ax�%�v�Fi"OVi߽sG2��5�Єi����v"O.�f	(n�]ѷ�%*�଩�"O�9��h�E��.Yj���R$*�y���*Ȃ9@�L� ���ɂ���yS�e���
7.�7D�H���y��5k�pv-Y�X�ܼY���,�y2	P�B�	V�Wu�|6AU�y��Z�dZ$�3���I��ϊ�y�'D�3�&�Z�CM�Ph��
2�y�*ǠL���3T�=4�LI�B_�y�T�1쒌)E �.9rΙ(و�y�
\**zH�i4N�/qh�p�f���y�΂GK�т��Ʉ�Y��y�c���\��_�zGй@���y� �^N0H#�(g�,�4m�"�yRjC�b�����2�:m9�@E��y�� �~�����~�0\�����y2�+ ����&I	�h���D�R:�yb���@� |9 �Ӭ^�����yhH` �ɺ[�&9B欋��yRЪ\C�КL"��5�W<�y�È�8ā�F虽I`�R�U�yR��@�,�¥�D�<8����y��1*��y�`eP�A`�@�5�y�L/YZ��b�@B�=�fH�Gh^��y�g�7BtB�
ؼ�"&�ܫ�y�+@"~���B�[~��8��ٗ�y�`@���`3��q`F����y�fI'{BR屗n��(���y�C�K���7e��� H2����y�B�S���2�#� wl՛A�ɹ�y�) �?5Ҥa�Mޘ<C�9�@@ �y2��(�^�ȑC��.��Xea��y�nB�G��#���t[t���y�Iťg���`�#	UV$`c��yb�K�oE���G��v�1�y�f��Z2���-�)��,i֦�(�y�+"h���ԝ-Z�S����y�"P��8h��,О�
Ub��9�y�R4K����,,(��/�y��#7"b8X*1��jT�ʋ�yRL����a��'їv-J���y�����P�GU�FXR�o֩�yR�� Cx �%�U��Q�����y�헐%�dlq@�P(��g�C3�y�'�
$L�� ��F���F$�y�Ď����S���o_T�RB���yb-��4Θ��`�&d߰�iP�@�y�[$"�Lu��OB\�\��M�y��u���!c��-C���M��y"�%0�������0��i�M�3�y���P\��0�%7�a�&��y���l\��f׊(��� ��ʝ�y�)�6�*dI@�L:%�M��T��yB�g�~p;%,M�"���h����y"H��h�-�mS� q��	qnְ�y
� ������~��Q#@��`z "O F�1L�����ϖP�
��1"O�Q`��ڬe�����X#��E��"O���p�DVS42d��h�l��B"O�ly�C�
x�0��e� �"O,�c�ETa�Tj����OaC2"O�DH1��1�Q�X�S��+�"O���KB�`İapMD;@K��""Ox�â�X�ޙ;r�U�>�P0t"O�}�0�n'\9� בj#�Y�"O��U�ELߐ�J��ɓ;���f"O6(�.]��9b��%P�4�"O<,�M�FX�Js(@/x8n��r"O�PV���Dc�d���87$0" "O"���E/] P���tq;�"O��y��<����ƅ�<#�%cb"O&87�Q4�X��e�@��2!"O�!�e�D���'E���j��"O6��e�Z� �2��F)P��9	�"O��ɣ� `�:���ݠ���P"OD��r�ձ�N�9��W*�(�9�"Oҕ���2��qH���%)���:�"O�Uad���"��$=v�R"O&�;�,Ʃy��̀�"o���q"Od�`2,EN�f��ϐ&pZ�Y��"O	f��˒��Mʕ<��d" "Oj��O�K󦁡um���t�*�"O�UQ4B� E~̌��Z�L�Pm��"OjY8e%��+��T2���V)*%"O���&���rVJa`��Ř8$��S�"O��C�R�aU	�h�
i8p�u"O�؃@���y�:C$CJ-�Q�c"O����r9.�$�-*�4�c"O�-��e�0�`�$�ˮ����"OL������c��9G$\'Y�p�A�"O�R�(O�-{h�0QHI#��0�a"O`��Dؓ1F��W�@u���U"O�}���R�~��M�(��p"O2E�[-vI<I���p,��"O�؁�g�"J�4(wlM7c< ��"Or$�W-W\&4X��
7Qb�8�"O¨��3��]��T�?D�+�"O�r��
x���]��\���"O��`���P�m��lY$|q2�"O��:�GY5��[ье ����"O\����|�z���T�h�\r�"O2��we�>G"���R��AI6P�w"O4,��
U�f��Z�Ș^<X�a"O*@J����,�� �ڸcB��I�"O(գ��6x�� ��|7TiRv"O���4���:��gT=O42-��"O���/^F�2��q��Q=0�Q"O��AʤlE<�I�E��3t �"O�䈥hR�X�J�(sfޒG��i�"O�h�Տ�<`��ۇ-(�d��"OtqXSL����ዑ�ֿ|%��`U"O��3�Q�6E���!H�,2,���"O�`���3  ��J�.p�Xb�"OM�`��pk���H�.T���a�"O�03��"[	�	qg�#r�Lr�"O�x��i۽Kz$I�,2ѺUC"O�8������m�#($�*�"O�D�p
��`^j� o� "m@a"O0���!D�Y���e�H��"O� T��6/�n�*{e���S���"O���@BW�d�.0Xd)�1Pf0��"Oj���`�;.d�S�燲p.�c�"O6e*B�6ea� �%f�0#ZD�"O"e�W����Yҡ�tJ���"O�����/1�X�E���
4Y��"O�LH��(s������?X���r"O��I�e�5���
D�H�=�"O(1��� /�n��F2JK����"O�Yӄg�-�B- �0?�T5"O~�;dd	j�b<���ڃ���J"O걪���<-"=�ց���9d"Ob�ؗ@�k�В B,+a�Њe"O�=	e�ս��btN�,�\���"Oֵ�Ł�*�TH��������"O��ɋ9�謰3��(?~|���"O8���e�%J��=�Į;8��`"O�U�B�	9�x�(�N�z���"O����원Q8=h� Q(��jP"O�=��$B�.��}(�9r���U"O~�Y�ޜ(7�[�M�8ek�APG"O�bW�I(�S�A�~W82C"O��"�5��8��<O!��ٴ"Oȥh���6l�T(k��фb`�"O��(�"��?�����q��IY"O>,�G,�)}��D�띄c��3�"O����H�?M[* "��+� �"O�{���u��噠	ݑڤA)e"O,����
N/���7. 7�$�k�"O셋b�Y�nH�����x�"O�0�B�3�auǄ�x��a�"O�Q(�S�hs��"?�Ja�"O��Fc��72���S����"6"O�4��²&5�u�P�=�p��"O������F�Z��׺
�<P0r"Oʀ9�FCw���X��B>a�(ɑV"O�,��+�C��G;%�2 `�"O�t� (ٌ�����Q�:<z�"O.|h���1F̠XAˑ����"O<|��e)'��$s�H٪�޽��"O�D3�B:����6!��� "O�!���˶G�4�3��)>�XKQ"O�q#rW�=�d�J�i�f/y� "Oh%Q#]�-� ��!.�[�"O�����/#��(��(�PX]P�"OۨCO��]�ӂ7Id����"Or�7nO�B��H �k^�f�!��ɮ*�Vx��mZl�{��Y�!�Zd�
�1Ǟerh���f}!��M�.n����&P�N�"��ޝ<�!��P�h4Q�*ԋ	�T`�C� ��!�bX� {a�r]>d��Ğ�!�D�|�cf� HV�C�-#d�!�Q�!v��"��-\���)�!�Sy_�:�'�BU�mjg�ǺL�!�ͩ,t�<�d�X-,õd�-�!�Dʿ���y��$��0­�s�!�V"�������(dw���V��.!�D�^�ب�`o
 \�5�ŊL�?�!�/O4hm�1��[���ELT�!�dC�����D
�`�x`B�*�!��7p�4J"@.I~< � iV�!�ĝ:n���OT( ��зH��!�D��I���r�)|aB���şW�!��  5��ӹDp�mB�&���lإ"O��	pH�-g���r��O��0"�"O�l+�׸���.���=�!�T,="qG��c:�ܲР�9'_!�$��Zۀ���!�,:~4���#\;!򤚶Y#�h*���0br���B(!��/ �h�k���7p` ��!D�W$!�D^;JX-��] 4����!�L�H�!�Խ3z%� bK"��c���!�T%MTV�Q��c��ԑ��h!�ƣt4�׎�l�b���a��!�dŏQ�b8#�
�8	�L��g���X�!�-7r�U�$Í2�PP4��,�!򤘁T@�5�t��B|���9�!���>
�ӱʓ��J ��F�2F�!�����peį���Q �U J!�F15�P���䙍D?05�BQ�~3!�X�Khl��I�+Dժ�G�'!�DΜZ�h1P'E��n �4KE�C�2�!�DR�a:x�SE9���R��=n�!�D�4MV�����^��3Q
��7�!�D�Fp���s�I�b���P2�!��ӿ�n����ԦI�RP�q&�DZ!���-�Qp�O�&����6���/C!�䟊K�V}�F�ٞU����v�ǴL)!�DB�b�c�eA�����F9!��Nޠ$�D�Q�B׬~[�9��"O�����S��17!Jz)�x��"O$�Ac/�0ZKF�0���^mZE�f"O�͉�јBDr����U����"O���B�?$���R8A��i�"O��Xs�[��-I��Y<�P�s"O�E�C�=HR`+b�9I�.�"�"O$���)O�+ǀ8�E^P��,`�"O�q!FI��S |���H"����"O�qe�<3bM�\�*�����"OFHS-�-7E8;㡘�θA��"O�p�`�l~�=�b���2�X�`�"O�(�q�n��1�.��g�l�"O�C���� :28혶j��R�"OT� �'�72�Q�@�o�rdv"O�	��ʞ��^%��#%�*qs�"O­ ��+ui杺�%@�JA)�"OD�Pc�/H�T�R'�&}*MѴ"O^ar��ُv��TbG�3Sf���"O�8����&K7<u+4%��DO2�c"Oz���Ƌ�Ā�.�JD�!�"On�9V�ڂm:b��C,P�"O<=J���9�6�'Z�%Zv"O����oP.Cy$li��S���Up@"Ox�i�	��  +�=b�"O�p�C�(T< �®� Hnb(��"O�q"���,Pޠ@C��&���"O~K�mU#/
��@��:SG�Lq�"O��ӑ/_�maz��eΥ :���"OvL�g�� ��݀L���C"O��H�Q��Y�"��X�ܒR"O�Zp�[�,A�)�g˼s�(!�s"O�0ⴅS!mW�PP���W�f�)%"O�1Ğ�k�"��'�<e���"O`���	��D�T � �Q7"O��"0�L�s[6L��ʛK�ޙ�e"Oȭ+@E�� ��so�p�f���"O�j� I�4F���H�
�:�ʗ"O� �g��.e��R�nM�B�<hʀ"O<T�%ERT��D�Æ�3 =��g"O Q���Ӓ#mҲc�/&�	�2"O��sNFRfN��@�_�)���"O�L��B�w�|z�B��'�壓�	����Q	*>���I\�#�����ń�^9�t'�4_�qO��DZ�y������	�>tN�ٔm<�tE��O��\#B�nD� E�{ A��dʻ;�8�9b��zRb���%)����'OS�0�S��Ok����͝�vҖ�Ez�L�'�?��gg�OU�vȍ�e&�%��m��_ ��Ӫ���$9�)������ª2"�5��K�\��p��$}r'7�#՛gg�v7�\~�F�a�c�4OPI�P�K����0<僧l�՟d���i*��W"E���ұ!�2R=jt��"@~!�&oG�/ B��J�}�aQY_�ʱ�}����M�&@� d@љ�'�9�pl���s�"��1��3	�Ċ2%T��P��k���(�k̗-;ɠ�7�É9��4��a��t��v��?1�/�V�'�?7�,:2��V�ȱ'K`1En���O��=��}�(�.������^'�@�@&Ό�(O2�lZ6�M�K>��'�u��!�L�FlE7^g�1Q&�!w�����YF�i�ay"O�=d�������3zI �� H$8�� aT�ol�);¤� ���)'%����7��h`l��i&
����۵s ��Q�&��9����:*��2�V?1��D۫K���p��lܖ�{c�W Oe����
6�.��I��M{��~�'q�tY��S��@��5�vg�hy��BF%D�Ъ�T�K��C�*L>G��T��-5v���~�V�O���˓2Kd�딄�57�T����I*N��t0���&�vY����?	��?)5È��?i��?9�eI�dGF�B2[�K��R�A�p�p���e��Т�#��شC��*��,Lqfb���r�S$I��YnB����2��0 ˠq�(�/1�:���@�'�%
���Ms6.��� ��0r�И@@��2g��O��D�O��ʧ$t�3l�.�>MpGB:,�eFy��|����"W����"D{��W�����	�M���i��I�fOU�4�?�O|²l
7�j���п38l�{!e}ܓ�?���Q�e<�8!4�*�E�eіd4�=����ᒅ+�Ѝ V�YT(�#=كjɇf�!�sI�F����,L�#��	S�4	A�A�+�9�B�bɑ�C�O %l�/�MS���	p�X��񈘿Y�8��8���Iry�T�"~�	<E�y�ć��Y��u��]�J2���Ӳ!l��] &D"#،[�n�e���Ѫ����S�۵�Mc��?�/�j�q�E�O���t����� �h(���d�a�b�^�x�ʔ�a�V�^l�LA�*9Q05cFٟ�ʧ�"]c�~UZ�MY��~Hӈq$L�2ߴcD~��Ї8�����ȰP�Y�W�s��ht_�p�m��k�,Ȑٲ4/h���k��']Bι<��y��M#��2'<@*��ީ)��W�I?����>a�EҀF}j��Z+���+QC?H>9�i�.7 ��ֺ�uB֜{!�x���d��b5KցZ�'Va{rήY   �]��"O���ǉ�r��	 ��wq�%�"O�eK"��,-�jgK��3�8�"O�d R�=`�<��U�^ . �4�',~UXVbB1{+��t�O�n>)��'��bfFH
M���C3v¦Y��'�"I)�0�ȼ9c�H)[�z���'^�p!��)z�P�3h��RQB�'��4s�*��kk&y�bң}q:��'�d��U��"~�i���@9u� ��'4�p)�䉣	*�	p���qu�YR�'!�0J�雵Y����d��d��x�'����oBR�0�A7gZ7J����'��1
EN��n�����>�<ĳ�'�� a�ƒ>q~*=h�%#RZ���'�D��U�Vj&�@� �J�K�'�p}ɰ G�(∑� �M7����
�'�b�`�^�q�^u�U��WP�)�'���%�e���"��S�����'�阒.*Yc�����w�����'-P}��ǙD&l(�B*�6FRRT��'�=8���&�#A)F�/�`@�'��A;��͗'1�T��]6-��,��'vB�z���UNPA�G�-H�ժ�'��5Ə
ls�(JpG�5I HS�'T0HW#ڼ�����Y>�Ę8�'��h��M�hpL� �n�"�'.n�q��gtA���4	dd���'�(� �l�.%yl˕�כ����'I pS0�]�>k��
�^�Pܺ�K�'/�BC��1}t�Cc�]�6�xk�'ì���,��w��Q҂�1lj3�'@)��1r�|���˄4]�F���'� �A�nF�V��;R慺[�zI@�'C��kQ�ϳ���I��#�'��BP��8kT)Bt-̻p����'
��9W��/
XM���n�̴��'����2lR3^B�`ƃԟ9�ɱ�',����eP�8�pucN�1��
�'b (A֮!m����əR��{
�'DNI����ڠ;�gO�����'J�02�BlJ�QAI��v��'�\�
fKL�3ŒDq�N4af4��'�ԉZ�-��(�`ѡ�P��&ѐ�'n�!�f�gO^d�A
Q �,E�	�'@){e)Ow�"������(t��'^�P��ϨY2��L�vzp���� �Q#&��bS0�R��[�Ԕ٥"O`��͔>�� �#L�����"O�M[Ď0N�n����@��qh�"O.����B�_j�#NK5_���u"OLjD��8G�:=a�MԈtN��t"O����s,��e�ÔnV�I��"O�qKR�	8Wu<*#�Z~����5"Ovx)
�y�@��4i�+]��<�"Oĕ��!h%���[W� `�"O���V�4�ԇp��"S"OR%#N�1i�	zjrA[�"Ob �u��#k����H�>f.\�E"O�e�#�f�R�!fǝ�	G���c"Oh1���hy>���y����"O�AS2���rG4��dL�y,Q��"O��;7H�m�^���@.g��`�"O���B���Y��5i#1�fMSD"O^�(3�W�&,��+��̫?�|hcC"O\ءU�4^�\ HRI�D]3"O��J�*}Hd]��G�8XD"O�M�F�H<*������1���`�"Ox��NՈB�����8Ү1r"OA���
�,C�ɱkZx`�S"O����g��S#�#�ڌ�"O�����+W¦Б�ݸ'�<�h�"O�y�D�1�$QrAd���e"Ol�bV(�Q�\��!��U(�"O@�I'�6PBa��ŲQ�i�f"O��kU�Q�C(4,�#@�?Q
�"O�d�5�[�:
4�FŢ!7ȝ��"OtC�o_u���х�W)^#ĕ�"O� ��#L'.���Y��p�
��"Ov��' �;���iw��<�,�r�"O�ЂdN��Cغ ��m���	�"O0�Ҫ��vHa��Gֈ=}�ّ�"Ofdȥ�P�dV����g�1:Sz4�"O|��`�\l���G.Oh%Ѧ"OrL�w ܳqL̍�3��.j�,��"O�t��)\��0�I�Zڨ��%"O����8�P���źS���"B"OD8�B�	]���d�O�H���"OL�{�Nk��)��IJ�|hBQ[7"O��vc����%'�(Y��"O~1���*OC��Vd�}r��)q"OVq�5�΁l�P�a⡄�S&dK�"O�b$��x3	�����#URh�e"O�R��9l6���+W�2F4]Zd"Oj�p�mɛC���BEZ��%����y�$p5 [�JR�ċզ�$�yrC�v�l��0��@�`m�W���y2L]��mPD畋6�H!�6�y�nG�N�����Ð1�0H��,��yR�N�9%X���"y�a���\5�yr�T,�>}��/$�R�%'�yB�ú���A��	f�:թʛ�y�eճT�Ay�B���b�D��y��Q�[E�D1��
y���d����yR^�҅��5���*�εy��M���]X��h�@�9>��Ú�m�(C�I Y���&��"C]8h�gg")xC�	/}"�N\:R@��W�RպB��;���q��b��"���e��B�IƦY�d�� 	�4����C-.�ݡ�)%D�xP�+z �8�@�l.�PWE D�� �d�ѠA3yG��qǮ�3\��Y�"O�܉�'Lݜ@��Q�>=<��t"O�j��(N<��Q`��=#�mA�"Od�)��@0�>Đf��v�c"O*�!6�]�Z��[ŭ�<t2�Sc"OX4��/hrv�"猟> ~��#"OZ�A�fO]!$���-C���p"Op�a�bOv1"��X���X��J��ym�1&M��Z���<]=@�o��y��8v;� [u�PY��iԭY9�y��1�8U���ڝC���3J��y��%$x� ���_n�0��KK�y"��~X\U��AUx�t�����y  k�j��P��wy�����	#�y�
��4�@A�߯9[�0` ��y2L�_ѐ��"$��b#\��$&Ԩ�y
�F�.���eA#���e��y�n2zX)��)^*�����y��\�XϮ	pU�ӄ�ih��S#�yb@�.G<)�`I)!�$�4���y�G��a1�aP�@�F�����h��y�e�/ADoʄ>� �C`�Č�yB�R�1W��R)�3�8�Ѥb��yR�-c�d�2�(�����.�y��Q�L��Q1�@�0L^�S����yr"X/x�L��IJT�I�#d/�yB�T��$(�oܾEK:�S⎒�y����n/;�X��&���y� Շ0:4	M�h^�Z��� �y�l��)�$��TB�ZK.L�@�:�y2B��z��$�	;T.�`{wKȱ�ykG�Bϲ)c�MЈ�&c	�y�b��d��I��3m�X�Z�"V�y��&���3�5j$�93�̈��y���[�J�c��]� C:}4����'H����D�0�%;�Q�pk�$��'�j��$AΔ )��@,[cQ���'�|��`�v�M����׬q�	�'�HD:��	4D�V:�D��%
�'?���PΛB�ᚖ��8i�<�	�'�*���@&?���a�FI�Br��'ɢi#���:T�%ٲ�D�Bv8�x�'���⣩��F����`�51l�ʓR�PѺQiK&Ld� 1���?���ȓU��2t	�EB �li(�����܀3撁3.���H	}~U��/��ؔ�O���`�˗H����ȓYbJD�1%>q=����K�=���)d2$�#`�*fd`q��G�
��P�ȓp޹�t�ײ>��LHAiJ&�I�ȓDMbpX�gV*i�� b��Ʌ�R�Z���6;�N���.�kX
X�ȓGR,���)��D��I��9��I��f�E�gcֈL�Z���`^�|�N�ȓ{��В���W���W�͆v�H���~�|yI�.V,�Z8`�LLj)4X��'����3�K<�s����-�@�ȓT5��s�![0��܋����(���ȓ0���s���)2`*��v��܆�H���C53�:�v&Џ\��4�ȓ9v��{��H'q��sJϷ]Y���ȓn���Q%�
�v6, ����ո��ȓR/��B��X����(������5Z85�V���z��������4Qx-��S�? �D��F\�a��Q(r��t.n��"O �'Z2���(��P ]=����"O�3�DW�j���kɞ�*OB#�"OdH��tEzI2	ʖ_0$9P"O���,W��e3�M�uMx$��FN�<�7h�W��h7�� 
7�J�<�	��~�$Q����&J�ð��G�<�v�Y�O�<���i�O����P.Iy�<���]+L@�EA6�L"�v\{S&�o�<�aNQ>+�h����e�b$��Yg�<�� �B]��ZQ)�,�^�*���f�<���G�%�q�O��īFk�K�<�J3M�����*Q�p�� �F�<��O�{::!��FR%#5�0W��g�<��Jٸf���d�[$h{hxU��e�<1�o��Q��{�g��i�䁋�@�F�<A���deȅ!fZGp�CÅ
�<��E��@���j� ��u��|:��{�<!B�վJS��Zr��1;�\�`�f_�<���D	;F���*<<�<`P��r�<A��WcX��:Ӎ�#!3� H�n�<��M+FV���o�!?w���ᅝt�<��K�,;&m1�K��	ː� �(�G�<)'D��R��	$�A
`����Gm�<Ѡ�[� �{��ʍ4�^�:q���<�тʡ^D�UCA���5=&�Ҕj��<���X,�8�R=1���x��Vt�<A�G�o��(���K��<����T�<R�T1}�Lu��;Y�(�+GEQ�<���J%6k:��EG8&02��P�<�&��8�^�����.0|2<���L�<�fi'J�%(4�--u�4�S	�K�<�ҧMb�l�cCl|���	%��q�<Q$'�������o0
���d^k�<�UbڜI�F�Њ��	��ȃ��1D�����"8��Q��F�1���.D�,����*qh$����>V4��6�+D�@ a��~��IQej��.����s�)D�P+0B�Út!4�)���uE)D��9@d��kW��j5ˤ����%D�dr4GF�0�b���E��a�b#D�lSucZ�/x����k�A\����%D��B���B��$��f��Uf��+%D�*c%�.o�NpP���V�fa�C�$D���FmSn~}P���6{�h����"D�ܫS��:%�X���R�9Q�q�%-D�L5��
����
j��e��f+D��yGܴ4v'�*pC�ѲaE)D�,U��
s6F��j�=Oa�y�g9D�L�&e�+8Da ����JI� `�8D�H:�JF��C`��fD&�y��:D�������<�U) f�:DYB�(8D����� V��K��ТX �8;�7D��G��	u�ʹ#��L��`�c�8D���b�S?v���AJ�hа�1I7D�\ZA��%�f����p���+�?D�l��'�Y�8����& ��h�w#D��r��}��0zwG�:�x�n#D��8JW��q���3�R��"D���+�o��P��.}b���,D�� �
&(gXt��/
(��%�ve(D��2��re�x�Ώ5bK���>�yB��1?��y�7.V/BE��B���!�y��1Y������D?eRtyओ��y
� ����E$+����4D���"O��b�G:�|y�	W'G@�D:P"O
a�t�XXDB��ŽVxl��"O���+�? ��#ꊡgM����"OB�����_�����ȈL/��H"Of���
k�:phǇ6-����"Of�i�Ȋ�R�������O�D*�"O�\I���1!0��B�)����$"O���n^�#��I2i۬�{"O*݃WFO9>�����k�6i_�l��"OPdP���FY0lT�X�v�.ّ7"OB%�b��cT�(�d�Ƹ��"O2�@�EP��7�}��`�E"O�4ITo�q�^�j�Y�a�����"OFAn��}����@_=zX�x�"O��r��)KiD��$o\���\�"O�B�/_=2D�JB�_, A!A"OhUQ�*P�$apY����u- �"O^MB�&D�c+�)��)h��0"ONU�pfަT8~��f����Lj�"O�5Jl�
B�H*��N@N�QW"O�l��ח�Μk�Hў���"O*i� �85g��g�ڳ>%�"O�I3�
]
���2k�p|,�"O8��E�[4K�D0��L�{����"O��X�g��Ptsfi�$k�<m��"Ob8�@kP���Je�]"X��i�"OVĻ�T�B�����:!��"OPA�zz�p��1.d-�"O��p�KI�=$�Ƌ���K�"O>m�%ΐ�S^��aɮ
(Ļ�"O6|�7O�g�&u1�S"�i(�"O1ۆĄ,l�����++���"O��b/� c�5����+2�N�Q2"OL]���>���x�J��?x���"Oh�q �=8�+�'��,q�ٱ1"O��
S(�)�L��F�����[E"ONM��l�(�^Y��&�vZ�#e"OV��NP=�*hXa� \�"O���smV��v��fț�1�"Ol�+<��y{�J]j�D��"OU(7�f�)��ѹ�DpV"O�Ma�-˄N\��fB;0�� �d"O�x�&��,��9�g
�����"O>@Y���N��Aֆ�2�≛d"O���A��0�y��G��>a�"O �R��[�/�h<�M��m	P�{4"O�9��_�9�L�A�	�q|i�"Ol	�Ql���<H���U`�Y�"OD��Յ�.�n�Sbf��e�ذ�"Ov�k b���l�c�ܓu�le��"O�)�P�� ����c�A��my�"O:܉0�� ��HC�J�#bʬ�2"O��Y�C3"�dP������i�"OP\s�P�&���(1!ݞK�P��"O�C4C�V��(�r��+�bls�*Od9!U+M�+o�i�E�:?�S�'�d�yD�X'Omz���j�5ŸP� "O� �C����&�!@
���Ջ�"O4}�uA�P;BD8㨍""�h��`"O  C�_�x;(�c���y,�)3B"Ob�RsE��Jl]KI]�j"v�"O�AJg��=O���p	Y��5"O �l�C�b�D�@"Re<1p"O� ���H
3p�a���D�-al}�"O�m��	�JX|IU,Z�M/�$�1"O�L�k��Lq2=+��Ww+�i�"O�m����>}Z��W���>�xy�"O����\-d+d�A��$�p#�"OZ���
ۇ�8�#�Y/��z�"O�H7I��q��E�^�x��"Od�j`��7������.|%��"O�T �N�B���"�I�=����"O~�q���߲E���nF�[�"ON(��*@�&��]�F,Ƃo\,a�"Oح��� W�İR�E�BU8�C�"O�0s���SnJ|�I�M��})D"O4�G&��o�I9�H�'L���b"O�<I�]�P�@�ف���pY*@"O\<�b�06�
�
��A�r�Q�"Op$j ��5s�u���m�1��"Ov���#�(>1�islY%!����2"O* ��V�/��)�Tj�'j���)�"O(UQ����l��@�G�C�(�b]!�"O>�#R�ޘ5�u��E�V{�k�"O�ժ��w�l��B�5g^us"O��@w�ċ4¢��@��'yq`i:�"O����Y-f��R�˜�WW�5
�"O����囓0�z幱��c��)c"O�5�B�p)�d&`�~�jE��k!�d�!��-��k7ܐ�"�I�!��ȁ}��cv"-�����'3�!�D�-�!"Ǐ[##�ޠr�GV�'Y!��ąx���$�ʼ&��\�r&�#2!��z�\U:��"^ވ�)�"
u!�$˞b5E��+>*b�he�8>!�_*j*��Z�l�(��Qt!��u�R�J�L�5&���+�;D+!��Y� a�e����<&0�kӈ2�!���Ak��":�V%��!��?t<�4�	.�.Ȩp	�-!���WWzA�"�ې:U�d	$��i1!��_�Ku�i��(D�8�n��O!�$B�i�I:�,o;��Wo�G!�Kh�j���p3b�I��+!򤛩|0��$,�-j�tt9�P�
!��[<	���b�%��|b��E�۬	�!�Y�0��:s��g`�yۇ�g6!��Z�>��M�#�J6M����T�)+H!�D�2<�	+J�&��Z���&?!�> �n�����*��14�Q�!L!��4���!A#�ZHy2҅u!�D��qOH41fU��8��%��|!�D���v���n͐$��`ǉ�Y%!�D�� �6Q ���>�W�"8!�
�%�f(�H�m� �(dh�)(�!�C�A�L�H��ᖩ��N�!�D�?g��� P8z��1�7n��^�!�ę�Y$�����&��ܓ�џz!�$�? 5jX9�������Ӕ�>5�!�d^5U(>T	��I4��d��<!�$WA-�p����Z���8C!��ƑlP�R��J$n���p�S-!�!��6��0�� �iW�����#G!�d�(a��="�j!L1��{"�O�!�^�eb|�� �ְ'l��!��To!��4F�> c�푃"�����V��!�d7;��x[3烿$�>����\��!�� ���ZJ�\��RNX�HG !��"O�hKbN�w�LD���AGB�)`"O�t�`薡c&�����D�)H�"Ot)1��L�.�d���h�;�����*O�� GE�;n�xz�[�P��!	�'��|xW�Y8o� ��ڥMM���'�Q�c˜��F�C�<EX@��'����v)�:r�9�+�@eP	�'d�my�o~�ĉ��;��IY�'UV��T��9h����3��5@	X�'/R���Ǜ�5C0lЂ	w��D���'{<T:Ձ���5է���E�is�1Ira
h`�`���h�X��!
�l�U��JI�a��
;^q����w�!�!��OO0$�!mT������4eZF )���UvK҆����k7%`�F�a�E7�\c�P� �ޮN�����)j��ڴ��!�I��M3 �i��s��(�A���a#T��W/�;���4�O���%�O�eɴ����f/�bGTt�P�O"�O��lڭ��O�2�̧a�֜:��{n����7DpY�(��E�M��9F�m2���d4J�Jg
�lڱ! >It6�xu��dUxd+��P9G�ԁ�U�';|������"�K�m&����C�2;K�@	�������"�����I��e�&Iį���V0Dt� D�
f
�d��j�-~��!�\���OړOP�D�O��A�"i��&W1s,����G�d��I�4F�Obf��<x�*Q��ʶF�����CP�M�����|�����$�-�3�g��`y�'�պ_RUE�%~�����OrVB>-L�0"�J(��je���:xK����5�fd(!.V:f�KCU�'��a�7.
BN�&�fU�éU�a�8ⅭG7%I<�i���ZZuA��l����=��F�@l�����A��o�R�!�Вs�K��xr�')�T>-�R,�95�! C�ŹK�QХ�ޢ��xbiG$)^.A����F��������~�pӜ�lKyr��	m7m�O��į~j�`	'k�6y��ĝ}8��@�&0��v�'q��' �p�^ R����D��I6�kR���|�BC��?���T�g?D m�v�'�f�b�ʗ>�B�w���@�E�v������d=�8z�+Ɂ� 5ZAe�r:��QU�Ā91b�'c��6��+qfꔐg��f֊�z� ����IM���h��׮#�ْ�L��h�b�v���p>qB�i��6�w��x�'M�5�n�9P�G�_˚��~bA��e6��O��S��x�ϝV�\ݹ���3�4�q��=Sk� L؆{�����G"1`d:�!��OU���1pأa�IN:���JqH!n�Af� "�C�&ڌ���E+~O�`���σ�F�Q��~�1 /��jA�4�Y�1���E*�QoZ�U-����O~ԕ����i�*��d`�����Ò��4��J�O��8���<y�}�
ǣrִ���M�u�~��	��(O��lПd�I�M������P�k�NE�t �Sx��@�n�
��'֤s"n�<-8�'1r�'��J��
Ta�|�u�E�Ro(���"@��]���K�d_���c�*���4���$X�l<�T�1��=Yb��+.SUP�����U��d�8B�2u;�S?��ٴk&�
�-�<у����3wJŅ�g2X)�'l��S��?���x��'�X�L��AF���<-��4
+�	R���'-�̰�!�Y -���0J�+5�����/s�l$oZB�i>���L�I�ɺ�j   �   ]   Ĵ���	��Z�t�ʔ*ʜ�cd�<��k٥���qe�H�4͔6Z <���i4�6�<�TԇK��,���I�q,�m"�M��i�F��D�J���PEK�=������0��1Ï���M�A�d�2�O̨ٴ4e`U�5��nzneP'�R(f9�'���1�.���q-O��qo��k�<(Oh�:���*soұ �dV�O�r�2)��P��-O��I�b�[%�?�ɤ3eR`�W�MW�|t(fNM/��`��e��'��u)����4~ �KW?2A�1P�@8RJ/u�u;k�E?�eeD�P�?}"J��l�~	�M~��
S�qĢ�x�-[��n1����<�@�5�sv"<9c�Xb\uA��B%N־t��J�~�T�%ቕ*C�I�lS��Hi~�Cd�!K���'-: Gxr��xܓ~��IՄ�4�!����FG�\o8V�h��� �Q"q�Z�	H���$�,\�28ya$7�	����a���1���;P�:0���H�Œt�<�H5�����zqO�l!�,�v��)���[�"Ԑ�x�	4/�����y5	+�PB�K�Ϙ'hP�Ex�
�u��%}y�9����	�pH  �?�*�I�5��hE�xb`��l[7(2[��Q󴅈�^p@�(�OP4�-O|�雡4�1��q� m��~�MK�j�*���wv*8 %g�@y�2\>�� 4}�i��|��J<�
/�����Դ4�2���"�0TH@"��s�	 7T�"-�^���/y��DM�]_�����b��B��1kp��  �OV��?1��?���ܠ�JaJ_�*����u�P{� (����?�(O��np��IƟ������a t[�HS���X�����$�g}��'0R�|ʟ��2d+[�p���)>ԑ�U-({A��3$� 
I�i>��7�'"�D$��X�#ف:E�T	T#�^�9���Wşt��؟t�	��b>�'7-�4�($� !��"�p���V?��E�!��O&�������?��^���I�O*��K��LD ��*E'���	��@����e�'�R�q�#�Qܧ
NDR7�Z�D� �s�g����$�O�$�O����O��D�|
!$Q�!p�)���U#2L��hS�n��������'������'7=歷��F��k5�墎�\��͉�e�O��1��ɏ \մ7�}�@)C���X�s���    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   

  �  t      ](  �0  7  _=  �C  �I  <P  �V  �\  #c  ei  �o  �u  -|  �   `� u�	����Zv)C�'ll\�0"Ez+⟈m�R~��8˔�DBA��a��/60yfN�%w��U��&��*ADu�mJ�+Vi6�;n�$QA��<�Dћ��n�r�rgȓ��V�J�����l t�T�-�O
+~u�7�S=3�̬�#��L�s����<�D�{G�4ӧ�4��r�BL5i*��DÚT�z �	��:�dIM�0�R�Kݴ�|L����?��?���T��?�~!��ˑG�Z���?�ȭE<��\�X�I�+F� �O��D��$��A{��
2�� *!��ln��d�h�����Oh��B/[' �	׾MD���?zhȞ|lE�Ƶ��5�QjP+�!�7ns�JvB̔T���C�x��I�<H>��'YREq��Q�d䏰�Tu8R��w���qAP6�?9���?���?���?�����v�KhR�kC$��m֯.�^%2�� ��v�h��!oZ��MK���&NnӮo��M��W�����Q��`)#�1�L��#�	^>u����\Oh݉Ƅ_�j)�a��>~M ��(LV�����m@ܴ{��O���������X��\M����5,���� ��n�1�90L�!?�S��LYr�̛)%���۴o�$f��t�_�e�t�#d&F9h���r��R�<(�7�¶Zg��o!�M�Աif���E�3.P���Δ$Ё��oȿj� i`�%�@��
Q��3��٫FM�� ��k��,n���Mc�E�����F반Q�+S5*��q�ë�EM������(�ؔ0P�i� �%�!GL4����P���';�O޹�`�Q Rn���tŃ�x�N���-�O���	۟����M͟Dѫ�
D0.����̰v}rQ�6�'��������������R�@20�Tl�p�*��������|9Hd��蒥)�����5W�hX�B�N�W���)BAXܟ|CS
�)Y>�A6�øt��l��2O�@�B�'2���#�h~d8���9#�1�?����?����)��.���'$�*g� �s �<Z�R��O����gט(����'@1]|��'�'N�OX͸f��Լ��LW� �yQkě$n\ɓ(�V�<��FQ�f��\��(�o���e�[x�<iA.�5?5@��Q�s����a��O�<�&�(��B�@�'؈`�KPS�<�� �$4�R���7�>��'*�X�<��e�TԈR�J��`�F�Vҟ���b7�S�O�R(X�&�[����GJ)T���"O�4��I�>
���f� p��x"e"OR�����Q��@3���	R&"OD �gď)`��у%��P����u"O��S��&6B�CTTM�P`"OL���-�=l�t�r�̸1=�(T��(��4�O��zqj�$A�q�����e"�"O����j�$= L�9n2Ջ�"OZ��P�Z�h*�1���7?V\�(�"OĸjP��7����� e+Nh�<y6����,C�o�r1�T)�"�Jx�[2����M��O��D� �^��� %NJ�u�f�2S�'%���|�Iɟ�x�nZ�N�[s�ft{���O�a�`��Z�Jt;7G8�cA�''�m+�0 ��\y�hR5�BH��08` !  ^�j��w�ӿ�0<��؟H	�4Q���'d�̱Q�A>lZ����DN23.�P����Y�S�Op�\s�`4i�
U�Փ�YC���2���Q��Z��X��:���6�?AI>����6�T��|Γ�yfN�Fh����(I����4T��y�H\�}�*5���߹=z5jǊN��yB�6P�,�*���4�p�9vɄ��y��B��x�@�ԅ8��hUҕ�yb�.	��G�Uy"dhJsn��y��xc�HS�pbd0��I^5.ٛ�|2%��m[���'��'B�	
�P����M��)&g���)��͎ xX��44,��cg�����f����XR�	d"С���
G7J���O��5OZ��5��� �HdWŖ
���wA����Pk�6)��ٓ���|��6nM�!S.O>�hV�'G1���'d�	@2{�,�x��o�ذ�А<��	�ly�O*�k6{�@��E�߁/p@
�Q��ٴ}��ƒ|�O�DQ��P@���W.�x��@?2m�1
�e�;j�0�IU�L�F�
[C�Ҥ����k�,� �C�ɟl/e�T���$
�.��`��8�s(8�x�TAQ�vT-�E�%^b�q�0L�}��$�r����`�:k�t��b��O�� @�&D�d ��"T �h�3ǆ:w@�!A�#�$YŦ�'�����2��h��s�H�
�� �S��Q�H(�I}y��'���'�z��a"45� �r��?(Cn�n:� �E��j��T��4��EM) ź�D�'`�l;"��
%�����P7-���4\��j��H��0� �]axҁ�?�?������Z���9�ɛ!�`$��FϚK�'���'hR� ��%*�ʹ�FA�5CA���
��V�b�촣��h+��� �ͼ�?�+O$L
"e��$?E�O)���=��,��#ԥU��4�G!�=6�2�')��˶JA(i{�\+&4��n:§'��Y(�$˘��"������'P��K��փ!Cf�:��\�?l"}�0i�.X#�5*t
į9B�x�s.K}~"��?����h���䗽a�=�F��8$!0��]�C�	�v�]�3j�;C�n1�g%^)A�V�?Q���.i:0p�6��x�JY�&��lǟ��'	
q�6�O��'��Q�p �OI�@ڌ�cCD�Jaj�F3��y���&=���O�xb@p���y��i]U�M�`Xą��;��|acm�A��ߴ(�P�ATH�g�n&l��6��%r�l�bb��`>h��D~�����?A���hOBL�$�S2F�+���cF���)D�@���]�����Ӝ�`]�Pͦ<���i>y��y�a�+
Ӗ����ƦB�`Œ$���u��=h My�^�D�O���<�|BL�]q����^���T�KRҹ��!M�y>t�2��9D/���ĉ�z�Ɒ��G���D�	u_|���ϓ;����c���N�T���I� vh�᧤ϔ]ƌ��$K<J���g��O���*ړ�O(7��1��P#���,E�L� D"O&��F������L�|�VX�I����u�6�'��I�B��K~Js��2M&����L�2ND���R�h�'r�'��LYJ���wf��7��d�������7
Y
?�ŻuB��W5�T�=O�Y��S���=�bnļj�$n�Z�rͱ������	T4���N%Z��'N�	�t�^���ƛ"D�]��3��O��эs���q� &�X��t�� t}�"��O�܉�C�'k�P�2Eg�;SH ����' 剟Y�%�	C�S]���'8 q
�ۇP3z�� gP��A �'A2��5���O�'�����٦#|��(4��Cޛq���Y��n~��!�����Ϣl^�`�)ҧ��p"�ȗ- $,L�P�ѣ}
B��'GNX����?)��)v��㡌�O�R�(@��l&��È8D��r֩� ��W�ٺ@��%�gh7�%W�>��G�ޭ,�f�� %FQ�g��ۦ��������)h(��1������Iߟ��I�c'�ϜU�Nhz��*,��M3a��9E�lXP��	=�?AP���$�
$�|�<�F<r �@����a��#��9]pT*Ć���?���ϫ	L\!�|�<q�._�����J�h��:�h�ڟ8�'�!����?����ǘP~��CN�V����	P�1�B�'%��p@�oL�����3��A�'�T#=ͧ�?�)O���ъ��!�`sv��
(sL�iR�ݶ+���cP��OJ��O�������O���"�D#��!d��w�daT#�>J���R�i�1)�A��w�	�%K�;tӌ���@L��p�aA�n�r4o�) a{�훠S,=���ȸgإ�E�͆ �q���?ُ��?v/r��cK٥|JR�Ir�Ė:��͆�p�i%R�+葒�!E�&�li�4�?����^���4a΍4���VO3��H����yB��]��ъ�F��2�N��مȓn�d��V���hh�h6�*K��х�3}�̣$/1R�(d  "��Fa�ȓL�J���@ug.m�� n�Ʌ�PC�u#�ƞ)cQN`{�E��[�9D{�����r���)�ĴC�\�g.�u1�"O���h� �RIc��Q�B����d"O�����ſw3ޱY�B������'�Vmے�կ~~B����s���1�'�B���&YXR��!ޗ��
�'���
�%��ah�.C;}��9��_��Ex������LS&�ֹE��dc���.�RC�m�I�� �Z��HЁ[�0C�ɛa&v�Pw�ćC,Ҭ��k��k��B��[�0�)#���j5�Ј=n�B�I�m29��AAb���C�uI�B�I���d.ŋ&�*��n_�C���k�d���	�$j~�^b;�����C�bB�)� FlZ���):�Qjg��2�2�"O> A�V�8��6fC��h���"O��$��:z �%B�$��q;w"O��C ��5
�x�E�$`������'b;�'?�)�Q�5v^�q���GOnͫ�'�@9�S���X �ݹ�e����-��'a�2R-"!m}� !^8t����
�'�\�[ā_-?�P냷�VAC�'5�\��
۳1�Z����&Pr�'㰐����qK�0���d�SQ?��qT�/�v}b�A�J�JԢ��&D�̉ѣ�Y�����k36U*��+0D���E�?.����.G�����-D�����%[d4��닆o����-D��@S��TFh	� ��6����'a0D���b,A	N�>��֪�i�Mp%l�O�i3�)�;�Qd"ќW� +�L�#�����'0z	��T-p��=µk�:!�n](�'��R�ډrl��8� W �	�'V4E:ȋV�D��Ч-�Z���'A�\�2ß͜�ae�W�x�65��'<����JI?N0��qb��w�р.O� :��'E�Hڃ��4A�j�����in L��'Q(t{��1bz��#�ΣX���'�1f���)I�vV'R���	�'��a� �$�9�Ḿ6^L��'{�HA�n��Bi�W��6j|9��I�����\(⁼{PuC��ڔ"�vԆȓ&��0K⨀�^ٜ�	f�C�o��T��jbN�Bc�(D.8�  ڊ`��مȓ8�Tq��.-Y>�
v���	t ��ȓ>�*����Rj��:�I�)bH�ȓ�QXe%�S��8j�DNv%&�G{2 _����@(H�AϯR��kS�@,nM���@"O��"֠ފv���aU��rCr���"O�x;AL>lD�h۲�X+�
�"O ��HR)YSh�DFS�,��qB"O�`c6�؅D�p���+[Jƍz"O��(�
P+K��("� 	d,p��'S�HI����;|��J�e��S�%�(2�ȓ-���q(�<Qe��[i�1@8t�ȓF/�` O��R���ǍX�7�Q�ȓ8�~080lڿİu:RfG�f����u�[0l�2^��ae.�G3D��:k���T�	<�  �#Ʉ^o|��'٢�5G���0�F+i�$�4��)8�N�ȓT����bA�;ak�-�$�=����3J��m���������11`��ȓ/���0%�$L�x* �H5`p��ȓjȘ����Z9~ $�a�X<?�΄����@0��Fw��Ǿu�~𚳡��|B��h�TT�``�'C{!.�z�� D�PY�
��D���[[�(U�#D�HkC��.W������6O�:�w�4D�s��S5���5�K9	cd��0D�\�!��1Ͱtcvʎ@�i��� �|蚵F�Dm�~fX�dǗW�@pȓN[/�y�B- f<���gV�@涀Ȓ@���y�BY!G�>A�%Q)M���3Q���y�'��;s41c��.��\B`��y�Ȉ�|���o]�s����T�yb�G�0w�9�-��]hU�G�P#�?�hEL����¸9�E�#d��LK�AV�{����6D��2��6���j4m��$4D�� ���� %�����+6j40	�"O��J��X+��,�0��gh�IS�"O�I��F�Y�F����Mt�-�D"Ov	f���вG'�Qn�Ш�[�(q�$!�O�����0� ���B�wz��P"O�!���ґo���'P7
~J�0"O�!#�,��`6D%*l�"Ď��u"OT���o��AԱ@SD�w����"OZi���?�*8Z�a�t,��v�'��<Z�'؞t"�v�Аe@�5q����'3p��T�Y������.�LM��'fJ5k�m�V*�]�s�p��EK�'�*��Fe�F��l8F���r��$ �' ��z�Q�X�ce�ޫAkĈ(�'S���M׬lR�-�8w,����d+JzQ?�X�
�>)�ݡ�F�>�U0�� D�@s7@��l��ʇ�(}o���* D�l)��=q�`#ՎU� AxAE�+D�Hb6'NH[�m1��؍j�����*D��k��G)v�@i�#�(��P�t�(D��zw� ET��!��VZX�tQҬ�O���)�'
�@���|X8%�!.�8���''`lA��"1��w"��6|�x��'���!	�՚,��+���p�'9�pbbj.�®1(�h��'� )�Q���R���J�Q�'�������<P �a���W��0!*O��Cp�'n\%̆='��h�@�8�p���'��!�
A6y��� �Ց.�l ��'1(:Ŀ��S,@�p�Y"H��y�㏓���M�&4as6&­�yRǆ�}�� �� Δ`@wg�%��>���Z?q3 �����H7V|�iæ�c�<A�N&!J���^�*��T��Ny�<��H ��83����g�a�U�x�<��`���\��"P;a{d��u�<��g�4���ݴC�J��f�r�<ٳW�f�Aӡ��Zy����kC�'��:����
=2V�2���V`�e)݋\!�D�k�N4`
]쥹pn�4[�!�䕤d&(���-(_p���G���!�$��1C����/��T^<1�A�K!��[d�� e��!s�58Ո]�-�!�,�EP��JlH�Q �0vk���O?Y�f%���CAHXom+M�`�<"V��B��M ���`�<�u��Tw����^q��u��N�V�<�dȃ�y�l���,T��X,�u��H�<AP��,�t�����=�H�b�F�<���;��FC�hu4�ACCy��ǲ�p>���Zd��!���4�s'�e�<cQvo��q!c��f[��@�,_�<��Ԉj~��P�b�="l�����AE�<ai��@�T�hR�ĶT���2�HW�<��')P<Q .�6-�F���o�kx�x0�����5Ő�*�5�OW��}b D�L�b	���
!�S7W�vi�`?D��*f��_:nt(r�V;d9�G�>D����@�w�ų��40�~e�C�7D��A4�J�?O؁���U�=�8 ��5D�����($��eSV��!g�l:!
4ړ/�^�G�4ƀ�,OA�N�D(yH�8�yb
[�	0G-yR��8'���yb�I�[�`��I�5xl��6��y
� ¨��*%���®�X|~�{"O�HU�YB�<l"Í�lx�j#"Omy�D4:F<F�T�f��J��'�������SY#���]%6v�X��1k��%��o�$a�q�;�f`Q��Z/G*I��_5t��H�<.�<��*�*=�� ���A���"/�B����(zm��ȓv|�5ѧ�68�qeF 4^�-��sD���5FF��(�6@���0�'K�Ly
ap�ӎ{�}�L����.X8�3���b\4�b�Ύ�|���N�p%R��ʃE�R@�螬7<�܆ȓ]�sg$W
/��m(�l�%Rd2���
<x���1M*� ��cZ$0�!����O�b���8`��H*x'����JR6�
C�ɔB���#+�=S�)P�E�"B䉧V\�xaP&�f���B�n	�<�B�I,w�©I� ��@��;�a��rF�B䉴m*��s@ţgz���F�.C䉆'Ex��dD�Iv)�s>\��=�S�n�O=��Ȳ
L?��V�
�3���c�'��{C�Ǌ>�Νk�W�/ںܓ�'n^��A�	&�q���K!)а�	�'�� Ц�^�m�r��hESp����'Q��*�=������M���'��Py���<#���p�ŕYd6l��h�5Dx���	_t\Ȃ�G@��<)բԟ^Y\B��[Gr�C��R?s�,-�/ߵw!�B�I�D�(�%צU%ș0�)
�;o�B䉴E�P��� .,��9%L�\BC�	�giN�!g��%�YX�l��^�C㉋i�B�ʁ��Ir�q��oL� �ĝ�I+����#	���&K��I�B��4�@P80Ț�B-�c�ɟ����O���O��!�"'4�g&�O����i>q�2,Y����Q�Nz�8af�)�&>���ƍ���H���Z���)�?Xn�bcbXB:��yd@�%�����O(�!���bx�glC1�43�	�$b��0?��BD�&u&l�u�j�0��FNEx�`0)O��� 91��T[�n�א%��Q�`+�l���X��Ay�Z>���� IS`��,�ĭ��*-kT)A��0�n��y��U�2��+v��,r�S�O�2"Ìҳ&�0�8�AD�WQ�x�'���"��tP㗛 ��?�p�K�'3 Լ���g~:xQ%k�`*B�O:��5?%?y�'�r�b&9�(��@�S|8�a�'2FDЀ�6u(.�a� �R�b���dXs�O�q�5Ma���+J*Wjʈ
��'���4N�)ڴ�?Q��?(O�IS�p�l�!�Ҕ]r�t�r`�L�U���O��H��G�>h�ax��Oq��=1�G�x�����LD���A�O�Vɱ��0^<��b�.�j���O�Y�P�˭:{X�{���Z̨�@ᔟ����O��$�On���'!����'H\�0�F��T��y��Q���ʷj��]�e�"!P�X����	�HO�i�O�
6(��UΛ�[�BA�(�1"-���
ɠ䛦�'B�'�)擇+��A$K�\8DigH1hh	�A��E���
Fꦉ(�.�8��u�Ζm�����ټZ�P�r
�>H�@�8�d��9�Hu�ϓK�@��	�=ƀP�`M	TJ��b� �;O��������?���I\� ��s�=|����2_�C�I�:���BV@��aXY���o���'��I?Mb%p��D%R�C㒌�����t���o��!�I���I�\fd�"��.�m�tܣ��|��'Q�G���7(�[� mp�h�J�'!*���ܖk�Fźq�^�:��?Pi"ڑ�F���%NV�%#�">�7*M�h�IW�'u@|ꡩ��L✽�&GϨtY��'�a~��4C�Ȍ2`���0# 9j�� ��>�Q��0��?,� 1S�Gެ\�ި�&��<!�̌�y����'P�I`���'Q����c�����8���15�[�A��B�(�"+Bw6�8�'�O?�i �M&)�b]����x�n�3
a�$�q��T���H
���4D�4同>,���b�Ri��
�Ʉ�y�B)�?�������$��� �{���I��KňZDb�iP"O������,�rQj�g��g,hy[�퉸�ȟp݊��ΡD����hK���� �Ov�C��X����?���?�,O���8S`p:�B��C4�3"�H�wA����O��'�N$3=B$x#�?#<� O��/�h���䙌)k��aq`ؘ>� ���7 vm�Q��%'��O�u��\�g���h|0�V��,����OJ��:ړ�y�D2G�Z���+B�q'v�"���yb̟�S��Eˑ��lm�=
O��?���i>��	pyFO�"��mC�O�" �j�kӷ>^���'�2�'�bQ�b>�CM��]��EB N��%�pP��%p��Ag�7´R�炜��<��OF� ���ñ��=��hE�!A�\d�G/��H�����<)T�G͟��pJ H��j��n� �'&ZßE{b��7:��d�¨�8>1<���I�
B�	�Y��!i+<�����`���"S��'x�>[x���f�$c>�+�śj;�%8uJ�'&�:��OPФ��Ot�d�O��R�/�z@�9�nK���4�,8"%@B�#�-BE)�#K�F�q��p���t�	�U���qO|�S&�4?v^� ��,�
Ѓ�h�'t�D���?ъ�T[�JIzI�5�ʙ�7�µ��$9�O�u`r)�!�t����O}R�a �'���`G���
7Wa��A�K�",$0�'�R�'�R��8?	ǌŖ\D��ۥhN�Ux�r�C�~��F{�*��!�T�Q� NYE˓�6��'|�v�x��ģs�T%'"@k�z#=T� �'פ�I�T�lӧ�9O��W%�(���d�6a��6;3��lR�{Q
�O��'>U�r�_-\�ƨ!Q�\�,q�%\�*��:G��=��<�w�A<�t� V��8fײ h4�P�b8�O��O�ۥ�>��[?5�F�5Qz$qA��H��C�O|�Y�>��
J�O:��RF��=8"@(�@�ղB��%���'c��{L��#M��H�=}��h�4����	M�~\)��P�V�v��t]��aE#})%�'��*2HL3B!Z�<�H"��Q�S��[�
.�S��'��,P�Otq��m�,�t9� ܾ)�!���${�2�q�X��'�|�D����:����tE�$oY�a�K��?�C���`�L3?��y2�נ�~��]2vR�`���_�/G\ԋ�����?I�.�O��`�K�\Y��gG8=UjE�"O�]3��Z(8�0��� ��6iXL�v�i*��|r�~�'~�s�"��A�&@��"o��
d����V��$�,F{���QR"j+w�4��R�S�aOly��"O��1A @�A-2�#v��;�ܠ�"O>�zC�����B79g!�"O����>0ߊ���d��iG��"O�Q���}`�=:��	+:�Q�"O8i�!"ζv�U��
�i	��Q�"O �a�䵩w��)�P5�"B���yB$G�`򕇘5W~���1�D%�yb@�P�� ��
�QGҀؒj�y2g	,Ӿ��g=_�VHJ�!��y"�����S�I�(KF��6G]��yr�Uh��4DD�+�&�f��y�fS�|�ڱK�"��#0��i�����'L�]s���Z��G��+WVD�;���0I�� 
E.Ⱥl丩���3@��Q�A[-$��k�%B�M��N�O}le�A,ìX�h	�a��)|�l�Z�FT3�
�*�)�_���2ƍ��ܐ��؆H�Q������bF�
\�HE'\�4�9��MT.5W� [K>amU-,`���C+9(��KB�<Q�\�/�(<��H�2.��1OI|�<ɵ23D<�"��R/6}Bt	�E�^�<����$�r�@1��6+��b��\�<1���1iHmX��[�D��T�YR�<i����.�2w�+V�h����s�<����8'�>̂.�#y����ao�<���޵c�Qe��M�l*� VS�<A���.�ƬI��0X=��qE�X�<�t��Z�X	e�N�?�`���XU�<��LIq� �JÄ��mq�/�T��L��8�Eʋ�SNzQ��a�9/Z8a�ȓ0�6Q�Mܤ6�D��+2Q�=��S�? ��	� �񉄧�-[�ya�"O|�2���"��]S�6/[��q"O ��Vg]+<y�tRq
:���"O�����;	�r!�R).�6	�"O֌���W�Od��)�3ژ4�T"OZ������@C�%
�'�@X�v"O"��r	�$;�nX�N�%�����"OXԥhD�&��$�H(��"O�5 ���T�rC�+��d1�"O��
���("�a���b�P�0"O� �5Ƌ>m{>麂���,�"O��	s�\~Z���Ň�+; F��"OB!Ja��
up� 2�J�Xm4H��"O�`�dN�,P�En%XkZ�"OB�;G��e6��9.[%qw�iX�"O���t�6X�����-ݸX���@"O�<x�Q-���0J��W�r�Q"O���#I��S�� ��Ì��\+Q"O�)�m�/h����({ߨ���"OLh���|7JP�`� ��"O�賔m��GQ�� �K.�,�6"O���ѠM&pa\���*Q��:�P�"O��E���E��D�7�[��T��"O؉H )�+��Z��[�4�
yy�"O��� KG�48�����c�>���"Ozt/ץ �P ���;4����"O�P2�G�W�&��/WX��-�"O \cEHJ����6��x���aW"O�D��*�	3.ā/��"O<rtl��\��!g��Tˮ\�"OT����|2�%؃���ZA*""O�!B�������B���� H�"O"���J�rf8� da��M�\U��"O����$��
FG'~�Y�g"O(IբO���R�_C���"O���cLB`El��T䇀	Uj�`3"O�5c�5����֘h���s"O~A�� �#���.ʛ]O�tS"Ozl����sҠ��f�(FN8T"O�ܨ�# �+�*��KF�45<�g"O����c��bdt�ȧO-�%�"O����R5���+%�A���My�"O&$��/��XQ������&"OA���ړ@���� g��!�q"O�ԛ���9��#hֿz�����"OJ`�D1VB��BgΌYЪ��"Oh\�6&�:�$SV�@7n�D{w"O|�I�'lU~���.`�4#"O\LRaEX�["9��Ć&U_��b"O�HW�s2�;t#%r*`��"O����֞;�6�@4�P�0e��!�"O�CP�ɀDK�(xd�ӉB���K#"O0����>3,l<��IĥJf���"OF0�&�ʝS�2uP�)T<�`�7"O��z6#�=��a��f <��UR�"Oؘ
���?rФ pgF��d��"O�}낉EU1��1UH'��H¥"Oڑb��B�d���-I�nqɵ"Oh-ё�Y��9��J2� �"O�,X�k�A��x ���t��Y�"O��7(��W��-Q!�J�9�:A�"O�aߧGK:���u�b�p�"Ot=`�Ǒ'Q�P<�!hM*�Թ�"O�@0WbLN|�R�銺DzVh1"O� �+��*+HT�s(O�o�D|"On|@�ņ	�Vh�&

�F9"O�4�3Ɵ�v��D��.��3��[$"O`�rAd�*�z��I�	o�x{�"O,�Yf.-�f�2��-g:�Xf"O�����ҡ|`�Rc'���p0"O
d��C6(��G �B�q"O�`I�(�3^+ā`��X5u�ꘓ�"O��Q�)��=
�n�H��C"O>d�C$Qٚ  R��+B`]�r"O����9~���]#J:��`�"O������43Z���"\3hh�"O�y���M=i%�	:d�ө:V��r"ON�8�DM2T���U���,�"O��0@J��b9ubdQ��#6"OP�y2b�bZ���A!�*Jjј�"Ov��T�h��t�M�U)$���jĖ�yB�� f����(9c!��H�h ��y�-�?����hV2Z��3��:�yb.��IaQ0/��"&t�qꅘ�yb�R;���I�L�/쵐��Ӷ�yr'�>\)D��5mI�f�hA��3�yҠ��`!�
�яul DT��y��S�a�~� W�6X:�TnC�y��L�E��90�L�s
��s�6�yb�@3h���!�&���ȕk�5�yR�#b��	��~�X�um�*�yD]���22��A�䜩D�P��yR�-O�v%Z���	*l�j�o��y�I �+�q�M� Xݜ�1�d��y��<Cx�\ؔˍ)8�N���C�y��<in��Ú2#����+�yb���vB���'*Q&3F@�5	��y��
	hy��/Z�:B��%��6�y�	�2��RC�=*��3���y��O��eH�)g	��.I926x����|c���	�Bϛ�ɇ�pH8�gi��RO����]�b'�`��\}���]$e8��&�5M����ȓ,�z!�Fa�4'�@T�J�XEz0�ȓL�r�ۖ�W��`,c"�^���ȓ]I�2��
&qG�Ia�R ԅ�'90m�"�L�t���N"���ȓe��X��͖4^Ǿ�U��*C�t��6!N$Y�NG�=q05�`��H��܇���q{�Ƙ:;�$�å�4�^���.~�x���RL�(�.���9D�0Xa	IIw�y��L�`1C�$D�,5 ��ED��!�S,h�4���"D�be)nd�|X�R&<\��?D�X #o��;��X�`ݖ	����o"D���"�R�e�X4�'#�aǸ��ӆ!D� �eþT�b�%����#�3D�HA)?mQV ��E7���B�2D��zƥ1��Hk*C30��l�P�+D�����
'P�������(N?�P!�*D��"Ԃ�H^:�#!���֨���:D��Ð$<�r8т"�"�X���D=D�H��
���pr`�P�5�|� �l<D�lȒ��%o �}�E�Z����:�7D�p��L�>9������}t�Q �'4D�ȻP�G^ak`?���ӥ-D���v-C�\ɖ��Q�#lp�SV�8D��j��7�x�kL�G�$D�� �z��O�"TQ1ۇK̄Y+�"O�1� �tG���1��*��1ر"O�]3S �y�`���x���"Oa��$�:9�T�,Y�X@"O�U*����J����唉]��"O�y�����i�D]�B���ʂ"Op�:���:W\3�Dֶ�bhq"O�l.`.\�)O�!��p�D"ODE� I
�+-l� HʐfH+5"O�AasGA.e��z���4�x�"O����iֻn\$���Č�=�c"O�|��P�����.ʊ1���"O�a�&j��8Y|� 5V�~��@"O(���VT\� ��)Rm8@"OB��R�Y�w>آ��K<r"�0q"OLQ�����
�[DF�s|��sb"O<q
�k��H�� �ΚSi�4a�"O��цhӵg��=z�+σ)i��j"OF�X0��8��@l� AQ�؉g"O.MᷥU4���!e�FF��	�"O��YT��_�vH��
@cx��"O\�w��	f��5"D�)��"OHк��p�F���ȏcM�!��"OJ�1$`=LefKS����9�r"O���oK�z8��	^; ��"O�p��h�5rN����H�R"O�����	����C��T�~\��"O^�3�I0K�̥#���u��$C�"O��č_ɔ�B��ٰ/��1��"O�H��#�L�X�ɾ@�0��"O����G�%���C�uʠ�9$"O���TSZ�	
�832"ORT���'IV~��c�)N��D"O��x��P���̀�d�����"O:ݫǎ�'9S:�'J�.7�NA�"O���� ���
Y-M�X�+W"O4�7��s�R�Y�(c�)c"O$����+yE�;W��	�Li�"O�	�0�)`��#'��9�tի"O�E�� ͯD�Ys`�������&"OJh`@�"'��訧���6���"OvPP$d���`���`?+���"O �a�+{&TȒ������"OT���Ɩ"q}3���Y	�(��"OXź%� ���s�N;Vd� "O��� �<GP)kE�PPըiy"OB��⛜tcxm���0g��JR"O��`r鉗/��ՋZ�J`�� "O���c�?n9�zp\l����"O�hB7g�6&��{'�ճ �
�W"O����舃`(��@H� $�NՃ�"O���6�X:�,d�$��'��I�C"O���2�H���)��+2ݔ)�"O0p����`���b�Hu�B"O���%C�p�������n�4i	�"O���Zk����`(>?J`z�"O���Ӊ��u���U��%.�H�h����@d�4�B��nԔd�q��"��'�v�jŁ�>RT�����@X*�H�'�b�I�/RJ�r�ʄ�ހ
t��'�"�����/��
d�Q,z:^	8�'�pB�O�$[�ŀWBT�q���'�"P�!�����[�?��	h�'�Z�QD��6A��!�Qbذ<0�'q��ࢫX�#T�b!��K&�	��� �5I���.i�l�%���"��V"O���2�ɋ4qZp	d�χ|dj���"OV�����8;�2&�5~>����"OM��J�H��
/..^�a"O�A��F�Ik���@ߺU(x3"OQh"'Q
*����G��	�朊�"O$Y�LS$*G�4�G�G�\�,��"O\1���$4��ڲ	�G)F9h"O�T�%��6?RJŪ��>ZT�U"O�|ӑ��387�C���B���$"On@V�P�1�,��MQ��(�FJ�<��X����f�M<�2K�)I�<9b�&~ǔTk�C@0`�>�ȅ��}�<��]�v~�9I���1D���D�<I���<��u��O�i6�����_J�<ѵ�N1����L�J�ș��Hr�<��E�c=�����v��hЧ��O�<YS뎘oAZm
��ECfA�d�@I�<!tg^;m��m��Z$db�FO�<M�;���IH�Xp��FJ�<Q3+�7F.��C�U�������@�<���ވ:`����W��F�<CL�\n�0��q�
P��\�<	�b�'|h�H����>͒1!f]O�<A����x�d�o"P|��
I�<��_�9;�D���zL2�� ��G�<a��еBe�������)#R�@�<!�FώB�@D"R��4/�Z��U�<�7B#b�=IRϔ.u/D�&#^T�<��%F�D*��E����	��H�<�'�@�|0ITf7Ji�U�;T�T;�GA]�
��e�No�����5D��be�D5�N`����"n#�x�3D�����'�x4�P�t�B�A�2D�(�����8���U�����c�<\j!�d� �\�EŎ΁�d��D[!�d
𲁋���/�L�T�dV!�D�&|i�f�Ox�H�Ԉ�!�d�d�r2@#w�LHB�#!��<&��a�*�9H���
�B$�!�$��7(�H%Ƅ� ��}�'d���!��%gJ���G����d�$x5!�d� ���G�
�lz�P�a�"O��@ߘx᠐%
W�Z���q"OF�1R�
	(d���IA[��-#�"O.���F��ACǯ�S\<-"O:1�-	
!'*DQE�S��)2�"Of0�2�S�}�h�*q�D"&�$��"O\ K�f�z��q�!e�nA��"O$�  �B
���X�LΤ�+�"O�uYv�� T.�`�.�&WP��"O���B()D�]�3ۈ)�䊲�!��,����2�L���1�V�w3!�Ğ�A"L�yb�Z:}��z
�/!�dZ-9������c�z=��c�"OZ)�7-No�XE9�o��+����"O��)��Y����`'I>�����"Ob����>e�h��U(x6�
�"Oh��BR�eӎ�0��W�x��.�!��� �2����f]�l� ��P�!�Q�|�Hբ�jíY*Ua Sw�!��`ĸ��u��@k��#�C6�!��]�L�:T*AU�Kg�&�L��!�D=� Ȳf(P2[�d���%N!�� ,���-H�����ZcW<Ͳ�"O
<#p��&y�:1 �+:�a�"O,����4?�x���ڥ9DĈ0�"O$"2P�4�40�UG3r�X�cG"O\��t̉�k�ʜr��ѴN���k�"O�tQ$�O���y��ѣR^���"O�A�7%�!�I��L�1x��V"Ob�b�n�t0�%�޾g�r��"OR�{҅���S��C>蠁�"O�V�d�"y�	ʺi	�(;�J�<���Y������7(t� u�HP�<�$Ɂ�G�^�aO1o$��0ABo�<)$G�*TJ��ߊi �0��Vd�<�#��@`�=��Ц�(�MMZ�<�4(ׯF�J�S�ˉ$���r�g��<i5�[�_�����ʤ���<��ٜ����<x��cQ�~�<Y�ڢvt��S��[��ċ��C�<ٶ$�?-� x��K �>4НS��GC�<��ޅ���a��:��aK���u�<)ѪE�(E����6&1����^s�<9�M�{D�ш��~T8�E�U�<rÈ:x`�9�ǞWu��c�%]X�<�o�8�<�Y��-6�0��m�<��C�$
��ivK����� (T���2恧~MbAFM��bu���*D�����(aT�Y���J�\����,D����O�-4����e�+���y�f�r�E��ʣ;�L�CA#�yb 2/����Sd6��R- ��yRą*�$q�ƯZ/9:u��@��yrCE�&��x0�kY�4,X��p���y��*V�TCJ�`���@FZ��y���aG
��1'�.6`������y��b4iW-C�8?���UF�y��8RJ�a"�fz�@�mR��yB�V�,G�xW�#lu��$���y�K�$@�i�P)I	ke0;į_��y.΁ �0L�&!Sn3�`I7��y�кD�^�����=.�ǬS(�y� �:�|�$��#쉡F*�y"ǁ7X)l�3��	�!C|�"FON��yRWI��\bQ�/]h�3,N��y��H�s���@��M�b� ����yB���nm20���R��|�q�m��y��Ύ(0�E/E
wZ��J��<�y�E��Iؐm)����p���x���	�y�C�
+�bmC� �pt�ȣB��y� Μ.X"�۴��g~�8B�ʒ�y"K��\I�2�A�4�>M�%���y�.�%6�pT3F��'�V%P�C�y���v�"�ҰK���5yA���y"��7~��H�$��	���F��yR�[�6b86��t��0YP��.�y"�;B�L<ӄ���䦉��J��y�c���Ba3��S��@x�3���y�ǁ�U �ؚ@���@iyb� #�y"� U$���!�.Ҵ���_��yB$F+
�q �"9ԅYBJ���y2�
4]^R�  #�l��cBeN��y�&W��� I�v� ���M�y����bԘ�ʚi��,h��Ϡ�y��.,PM1SW��b2�S��y����!H�t����+�֝�����y
� ��ñ�S03M�5c��Ʈ�@T9�"O�0@#�+A*]A�M�#�t��"OH�/ .P�Ѓ�@���ڢ"O���E�M�c��q�4���#�"O0DbWj� /�Ra�"�����W"ODX�ֆU�A� ѩ��+5�8Q"O�-�o�5.�S�*�?�L�s�"O�bg��^��B�(B�xT�v"OP#lȁ-�Vm���Ʊp;��S"O>���;h�����%1۲�z�"O�ܳt�\�'Z��3���(�r�%"O��I�BW�v��� �՚V�\D�"O��0ӈO��r�r�DA'�C"O�ih��ݨ#l���f�#&�q"O���F�F2�rZ�D�x>���"Ot��s�ǣI���FD߽ Lҥ"Obt�䢗�?Ҏ��ej�z|d�A"OR2Oړ k�["	�xJ�8"O8� S�Ɓ<�:�n�#��)D"OF��c��JL�'� �!b�w"O&az���z&m[���*R��С"Ot�Q-��m������e&&8�V"O�y*Abǂr�xH� F�u%�8�"O8�d㝧���(�S�\�"�c�"O`v��d�D�U��t�|��"Oi��	�~0D�R`	��p��"O����a���U�Ո���H!�D/o�2��AIZ�!	��+��p1!�D@"_H��d���<�e�+� g!�D����%�"���lġ#l!�D%R_����A��g#��*���m5!�D��$�X�*g��Y-"8R%��.'�!��8`Nx�!�� x��2L4K�!�䉺c��h3Q�6+��Y�rmK�&�!��ن&!Z����U	A�L�����'=!�L&hP|[��àQ�ఁ`��z0!�d�G���Q�NC�nU�pb׫k!�$�<�x��蛃�@}(fh��.!�$��C�*��MH(4��3���	|!�[�T������D�a�����M�??_!�4ܴ](�K�4]���[�#��;[!�$�>
z	{�X2.�dY��on!�dPo�ʃ*�̾Y��-�jk!��Nwb�i��L	 5�`S/�f!�^�2��pR�L�_/�<9 	;O�!�ā6 Wؕ[�kZF|�O��!��ە�.��V�/9�\�(b�@�!�A#!�>�:`G�A�"�8��Ō3�!��
}����n΂O&���Bǟn!��D�G4l-���C e�iѳK�@}!�d�kT]�]
A�Z��0`��w�!�$����k���i�dqł(D�!��Px̱r����9��	�!��-7�`��e�2�J�3����!�X6ɨ�?m�i� B-2�!��φ%H�����5����� Q�!��Qn��-JԢ�S���g'P1p�!�$�qJ͠p��]���	�e
!�!���(���b#L :�*4���%}!�S��ճCl�V�C���G�!�V@��a!F !����dW#�qOH�p����q�� �
!20�`b�|2c�v��P,�8FIPC؉�y�n�'![�$�DC
"��8�-��y�-@+aV�3elI/"���0�y
� n��*�/H��mc�%P6Q�� �b"O~�iF�׻`'����T�>|L첶"O�`I���.>| ��!���\�Nq�"O��h1��D���A�JO�h���"O,$Ȳ����W�)8X��D"O^5Q���J�AMܫg�)
�"O4���'H�4 "�Ī3�z<I�"O�A���C� 50�hp�6X��"O�D�w���V�T`�
�l#�Ѓ�"OPػVJ�?b��c����R�"O49�#a͝>y*�z�	��3�ܙHG"OP|"4씦~a�ֈ� @"O20d�րl���(�a��A����"O�M�'�	=ͤ��e̝Yy��b"O���Df�[�,YQuN���Dq�"O^,Q��E��Z���&Z���"O@����y
��`�"OTP�ƣ�#���$�B�r�����"O�%c���rT^�*"�H�0R��t"O�D�7*���لCCI-t�"O�����(Jb��@$|�4��"O��ӡ^���#կ	\w�e[�"O��7Х/m�9�w�ӊ1���8�"O!��@Yv�^XjG�A�D�bH�"O��k��.qe�Q���:ua���`"O��1�R�ap�Ñ!B�.J63�"O�lj�H:N��x�FF7��@P�"O�:���U��	�A�O�(�>T��"O�'�Bf�5)�oܧ2w�IA"O~y#1%��r���� O�(@]��W"O��J���)�����NI(I�S"O�XS��=��p��7F��"OjY0�
���� Kwkb�д+7"O��	C��@����dL�5_<�9Q"O�8cB C�x�6U�J�q:�G"O�´EH*����i�	�^��"O$u(��=�x ��= _:u��"O����B�;���j> 8�"O 9j Gч{��<$h$FMa�e"O���C�a�N� ��L*se����"ON�����;ah�!��H�^be��"O�����bC��ʀ�-���7"O���ʱ_�䁛�B����4"O����%1�����A$c%�g"O��AgB_W�fQ�V�z���a�"O�i��
T��b�eݍ.8�9"O����	��R�CW	m,�"OD9k#��+�BIS2b@�x�
�"O��8��"-�9B3 G�3�ƹ*�"O<Z��S�>,��O��<�tx�"O�tS����`J���&o�`�"O0��e+=�t �m��!�x���"OI��*���q�F�%����"O°)W��A{|���D��\�7"OUS@��9Xw���ΑV�~�Y�"O�=�P�����MJ��Z�xQ""O�HʅC�8�jR쓼t��p""O�k�Av��XANNEȮ��"O",�'*N5ev<��,���\�G"O:y����:��U�G��i���1�"O,�P��Z�p��ݫ�#��2��Q"O�1!�f��_	��EI�:a�<(�"O�q�D^�C�����Е"O����Ɵ6}1H�#%�ܯsA���"O� 2�3��	�V���M."xq�"OB8f*OX�����>��A"OZ]S&&� wb]0gς6:�e�"O�hs��@�h}Zd/ǌ$����"Ohi;G*H!k�>�'�8R"��3�"O��)RH�1��Ȅ �9�0��"OT\��-)I:��ӧh�;��Q�%"O8�v�	pe�Cr�R�S�j�B"OΤ�P�کg@�cԥϥI����"OҠQoQ���h��6��̚�"O.]Aqf	I*���QAȐN�:d+�"OH��J8w�b��Ə]�L)�"O
������x�'nQ��X�%"O�4Rt��J�� �@F[��#�"O�� c��HC����ٰ��"O��b ƵX^\�Ja�<)���"O�)�b��2�m1B����G"O���B�L=^�R�Q��S���m�"O�u;���~�8lÃ��8��yBd"O�4I���1�n8����kNve��"O����%مa!܄�K�
6L̛�"OƤ��HŎG�B �R7�Q[s*O�jS��5�2s�@����A�'�cc�߭>pF��A�[�z����'��{1�ūrb���5��oA�x�'&�*5#��$����d����'��I	U�	�$`b5�O#I��) �'�.mk�"l�fQ����:B��3
�'���K��E b#���s,Y�4p�XK	�''�Zt(h�@y�+�!u�[�'��=��(�SJ�S�S�g�4h��'e|�Ct�/n��)�� \�Q��'��$�w$  >t����n�Ѹ�'!� 
_�G�B��2V6}�'g =QEdY	6
x8�e\�.4H
�'.�	{���=�@-x�H�%v,�K	�'6�L���7:��Paf杖u��'�������l�j��a�xͪ�'���$&����\�AF�-bqb�'�.8q@��.Lg���M�7&�F4��'��J5 ���{!�"�$�A�'�8Y#ǝu��$kR�8�,Z
�'h�Eٷ`�}s�M
e�0Ӷ��	�'�\Y��/T�B ʡ��vF(���'�Z��%��֭ ���n�� �'RX�22�ԉTh}	1k�`j��'����Z�>�4K��	^5z�b�'Vz����!Ax���ǯ\�^�z*�'5<����J�c���a	Mdwzȓ�'O�5ۅ��/g���"��\3�'��x�ӭ��Dx"E�1n���'�$8�1�	?�F�1��5��'�T������3�)1!�<��'^��;E�P4Q�=c��0x�X��'kظ(�ZW`ʜքE�+�tp�O¢=E�T+$b�L�rD�ӐdM�H�g�T��yR[��� ��Rk���u�ȓpڙ����t{���-�9MxA�ȓw�fPi���7>�j����ӵX"z���+S<0��U�Y�*xҲf��,��5`V�I�A��yF8����ܭOwpȅȓ.~�C��/%�Ԙֆ1z�����wb}�hڨw����+Z��ȓ*����`��@�i`�Q�$SL��S�? X�B%�(-��4A2#��P�"O6�٦.�+�d����Q��Q"O�	�dlZ����Oz*���"O��x4�P'A�2������P@"O^(��FSM�t��2��h��lS�"O뇃 .V����͉E��t�"O�P��j"6�>]qEL��}�"��V"O\ixc���^���
H�2D"O�X03B��بƮrjJ���"O�5Z���� �.�sEh0+�p
�"O^Db#�EM�.��"�гi&H@3�"O�EuB�=b���r&�K"X|��"O�R�^�I�}qQ�	V�l��"O�e8W��'!��U8����""Oz��U���:f$9i"��V���
"OJ�i���,�č��͖)��i��"Oh�`��' �@	av�Y�*l��A�"O.QY@��L��s�+A:���"OdP`�X��l�1�c±#(���"O�90��.gP����7O��0"O�1�H�0�Q�t��>�" �"O
��q��)T8�����+3��'"O>�%[�&���V�H��E8�"O���cș5�R�H4g�r�dx��"O�l���h��u3�FRzp�"O�� �B�M+�A�ReߏHY:X�"O�%:��͕f\b���dx� ��"O�52�J;x9�3!��-jX$"O>�KH_�`:�ա2�D�b< d5"O�}h�+�yd��*���,YȰq�"O� �ٕY[,���֔aM�\��"Otp��l�j�����G(����'D�TH��ؙw��9
��]�p��9��)D��H�υl�����o� �I�'D��{E��::��D�n��9����� D�����u���!g�V|���rd?D��)wmG!�tC%��n��pH�c?D��`f ��s{�؉�D9A�g�;D���WJ�H�<�uE�.m�(xPF/D�<�TC�gB�0�#�"W��R7� D��7�B�(����kI�%^�C�
2D�0��Ϛ�r
P��ň� �S�1D�j��՟ul�U��-΢<� ��G�#D���UG�>��z���}���q�f D� ��-I��%"P�5C9��Z�=D����E% hc�)��S�Z���&D�T �D�i�ZՀ��W[��IKA'%D�����Ua08���R�*��<�Qn.D��xË�;o���C@x��j+D��"�*�u�J<�1o�s C+D� 1�m�T��It��$��l9��6D��j%��8�@�؈E�lip"3D���" �@=�"��@���2D�[�J�-̮)�qh�!j)��*2�/D�T��ܲ���߁e%2��&�-D��;�ø* r��qk^|��*D���fc��B~N��&O޽ ��H7#&D�4�ԂA��f^�I��$�r D���udP(�'	��X��t���<D�8�dՔ4��1(���4C��C J9D��1��9@�P�ӰaX�Z�:76D�𓰈��#�b�*h�"MхN4D� ��,?<��� u�aR1>D�ԁp/Q��
��a�>$q�C�)� �*5��i<����Y#2Y*=J�"Oz�1���6�|y����3QVZic�"O�}�O�+Q��p4�RHs��"O�$	T�Y�阄��'�,Th4�"OxQ'��/tNt�򧖐S�nTɁ"O8��F$"qo���fF<L{��D"O�)uN�a*�;C��<wpv�0�"O��ҧ�={o�e+d�>R�^];�"O�G�SW~t�RF��Kрɡq"O8 �$�N3�)����F�)3"O~��Z�O���11d��Q�F���"O�`�@Dʙ�
��#N�v� "O���,�^iQ�lվif&�"O*ݛu�J46���r��-M��)�"OJ)p�t�MY�S��x�����y�E̎d��+ .όB�d�*נ�yoB�,a�q�$O+�(�ZW&�y�̊DG�	G��~�*ٓ�e�>�y��O :X�@��@�|�H���yr��&��z�'\�&7��S��F:�yr`�x�h5� ̐O�@�3�_2�ybO�F��M�c�	���F��y"��I+�USa� tL8a�lJ �yҎ��EL����Ѫf�@�tMC �yR���>p1p�ބ\���g�5�yR��U��H��%��^D���1�Z�y"�D�=�=��"�&+� <c�N�0�y��}�F)�(ΓX.b����yRo�1��82d-X$���q/��y��[�!��8���$�W��~�C��8Y��, �]*�3��v�C�I�cw���VgD="��'����C�I�T �5��@�&vu�7
��!�dB�	~ٞ@;�a�.�JI8���5	`B�I8�z���ђ1�F9°��(B�I2Zw 0Y���-L�1��*7B�	$tAk�6������j��C䉜���paL�'h�q�-E� ��C�	�#.����j� 6ŝ�f�nB䉭8lp���]�t!V)�'�i`FB䉔�`�"�±h@>	���;R��C�	]~��JDώ�/�6��`��S~�C䉾�tU3��mx"%�N�F��C䉧c	�� �H-b���#�Cͫ(I�C�	>U����F�����lʻ~��C�I�s�HJqA�w�ܼ!r�\-�8B�I�dO�)Pfӎ39�C�l�5#�B��0=%�Щ2ᔲ�D����	�"O ��8B���*��[�R����"O���f�t�ʽ�$΀;>�(�u"ORYhq�����2�
��"��X��"O��h%n_�V�,�◯�0u�^�h�"O*	[���	����&O�	Z\)�"O��ےkI4l��x3�Mʄ&ٲ��2"O�}#r��W�𘁡
��E�8耳"O���V�H�K�<�X�3�Rp"O���B�#"����F-�t�iE"O�0S��*5�
H� �Ӷ	oh@ѡ"O&]�mC�I���k��߰tO؜��"O��9�L�I��m`Q��&?���"O���f! 4+�f�H��ڸ���ó"O.�A"�T.�m�Ffr�l�+Q"Ov���.+08��D�#I��С"O�92nH��I 6���M���1"O� lD9�n-Rc*�3z|�D"O��9��>&~��)I�[Nt�B"ODd�e�W�f]D�����3OX�I�"O�@T� {�Y��k2_*J��'"O��au��b��� ��l�r�"O�]����'����K�6��x��"OJuP��1r�b��Cb!g>���"OzP�Ư� }3(:6k�u6Qh`"O����Ke����Ծ6l��"O�Xc1�ɟv��h�G�7���'"O8p�A*�`�x�'K�7�6y(R"O�U���$R�~���ɑpt�#�"O	�GE�~nPp�Ҩ]e����"O}���[��6�(wh�8cxdk�"OhA�գ9NUf!�#�V���|��"O<��C7l%3�'�|�0)�G"Ox���Dޥ5/�s�)��X��"Ot`SE+�Eg���i,?��zP"O��3��/f
|R�AE�|�t5Sg"O�| a�ΑJ�p`���"�(�14"OB�K�Oݳ7.ؓC��Z�B�)�"O4�C0(h�N(���#f�D��`"O�l(�"��6pi���oʈ���"O2���K	\��4�A�F)@�^ ��"O&�Q�C�8c0�T�0���jt"O���6$(�|���2fIv\+7"O|���ѹ+jԔYp���$~�p�"O�]i�"��g�m�f�&*l��"O`��SE@D�{V&��o&iX&"Ol�G�P��8\��&�0��K�b$D��K��Y%��ӳ�WJ/JJe D����GM�q��0⥄��GQx��K?D��ڕEE�'�8ҕ�(�t�)6A=D�`y�GQ \�Hʀi���X�Q�g8D��8�Ȳ�|�홌~�&����5D��I���&>a�e!6��h$�?D���aI'.hx�s��$�*���!D�D���ސGG�Up���2���A��3D� ��L��[�6iWG�:^�r��?D��1�GF�O��i�g$�oĪT��#D���M��tf�m,�8�D�>D�4a��K�3��`;�ٶ�J����;D�����4<���r-��@�"K��9D�P`�/S:Pu�uC�AōP�
F�$D�paH�&�ft9a問D��Ѫ��#D���c�&P�Xڒ�ԜI�6�@/D����/+fM�58�%S�MJ��cO(D�4�A��b��Ѐ���S&)D�� ��1QyHhda�1Q�����&D�T����W��ǯŧ+���W$D��p��P�u~H�z�!����(APj<D�t1��^Y|h\iץPQ ����o8D��`�_�yĉ�aiۍP���%�1D�� -�~C��;�'�7� ��*D�(�g+�*���A����J�*D��e��.< �$��q/� ��&D�"�NF�/�LXc�j�=+�f0B��(D�l����\�8���� (�YO'D����y�5K��>%��(
�j7D�P3���ZF��hB�
J�(P�	6D�PA�*]3q��dH�^L�ೳ�4D��;���"�P)0�?H�D��8D�lpT��/!ī�ׅJ����6D�4	T��
��U@�&�:=�n`��l5D�� �` b�KF�=�f���x�U��"O��3�	���4�C��	b�BU
t"O�x�"7e�tN�o�B0"O��#���d".j�����f"OJ�3���7<Wf��oR��t"OV�j��)x@`X��A���L@�"O���OɌERF����D6Hْ1�4"O�|��Bٴvl�����/�pq�W"O��h�&�5g�zx�n�;*��M�Q"O�A�̑�|ZBip�l�>���V"O* �b̯3�vq�T��,Q��S"O6�����6+<�� R��l=pDۂ"O�e
��<�~����O�H.4��"O�42(H<,.�k��#Ct��#"Odr��[U��	U��N^��B�"O�ɣ���K��\B-�&�b���"O�)�&$��}��i �&Z%p����A"Op`S�!^�Q���Eh��� D8�"O��K��G�$LC�&ה}����w"O�QCɟ)�$�[eZ�~��P�"O\1xI�<� �j��B�vp"$"O��a�-���L��%M;|�C@"Ol���#�?�`R%N�E��Թ�"OH�їoQ�k_�)P�%�a���{B"ODY�u�E�
�&�*�΂:,ई��*OH�r0����|)�&ٹx��K.D� X3 ؐF�iK j�7Wۮ��a�'D��P5)ש
��Y���Y�q4$8�'D��tꛋt�̉��؝340���/D�h�aF�3D��00���N�<��D,D��0�F�Q������`�*e8��>D�̹�{�T�i3�۽>��(�Wk8D�`�`É�W�KV_�v����)D�T��iZ�L��Ȱ���� #G%D��� �	E��r�WS��'@#D��93`?r8*�;��T')Q�0�?D�(Y�O�4|'v,��됴-j����)8D���cچ&�ؑi$�Й@�~���i9D�xbJP� 8CV��	J��$	7D�ȃ�E�<��0K�
) a5D�j�a�N�x"0�̠B��(D�r�
�#�~�h�+�-cc��K� D�p�ٸe
B�[%`.|�`���+ D���@�P�
2RQ��j�i�(t"qJ(D�\:PjT.=�֡��eH����#D�(�Dą���!�t��):`/D�d�1ƒ=��T2�����(�ק,D�Tj��O�& �*C����X�(D��3j�&�Ɯa7h99�f%D� 0�e� s�&�Q+R�?~�AB1�#D�����U�2��QF�,I�tXɀ�6D�xr�I/ �rd��!¿"���E?D���	\�k����3N��R#��t�;D�����:V�6��g��	~�c6D������{��AҢ�
;%�����'D��9�B�63[h���N�@���5K#D���V�ȃ �>L�GDM?��YY¢?D�l!wjʮ"��l�n
�f0��b=D�X�%nO.�@� ��{C&\��!&D�����]�*d.�Se��4%+@��1D�,!QA�V�����3��)D�@{����
z!���N"	86<D���P�=Q8I(����6�°��h8D�\Q1�����2"LΝ	2�9D�� �,�$�2%� Z�ԒS��h�q"O��a+!2�fDI����'"O>�92��9n[>u Pa�0��|e"O�E�"ŗw�E��S�B��P�"O��B(��`��܈�#}�"�ʗ���p��sɛ�'J�_?���e�"CŚ��@���`��7�+[Tv)R���?�w�<$+F��*r�ڹ��
bo*@3\���l\$%�N59aΥ\&D���Q��HOֵ�e(q�|�S�V4:r������|� N��QBB(��at��ǗN�'�pT ���?9@��D�i� �
���!��}��.*Cm[���O��"~j�4c��p��a���t[A�����ˉ�d.��O��6m���oZ0j���3Ѡ��\f@����A�H֞���S��X��iQ��']B�O��`y��'�·i�H9$�̢U!� �5! ���x+ѫ�u��[G�XA�h��,"ɺ�H�O@�S�?Ѯ17�
��$˵����td^�ﶈl1p�؈�@'+�f�k"�+nr�s����ޙ���Q dTFr�D�4�1��iy�8����?I�i��s�$e��I�/5����Ũ��pȻd�ON��,�Of��rY�.H(Px�I�)Hҍ���O6�O��lZ��H���]���x�0�Vp�$8�'
@#L5���?A$,^�_��p@���?���?������hӄ�I��S�6�n�E�/D����F�3_��r̚�nԜP'��_���4��@�)�/y�q cAU����`�ĝ`�8yD�:x��C_-��'"�����ޅs�2h��ސQi��9��C�\��II�\��Of�&���	Ο��'�<�R*Y==���'\�uے�؍�$=�'&�.��A�{�Ɉ��8<�
�b�qӠXo�r�	g�X��+���O�0��5jH�$����3nb�H&$	ß��	���	`�� �I��$����Q���E�#�ݺ�e�iF��K�ˠu��U
�rX:�uB�&#���	�k4a�2]�A�\������Av�U����-f�d̹�o=��yPg]�(˰#�}�oʲ�?��4J�(P�@�V{�\c��ȪI�$���O���*�d7��R8N��]zcaIf�~�aǙ*�qO�tK�)�IYŪ �6I��,� ���y�]����M����?���M0D��i���'��;�4��� (O�̥:a�2A�X�n[�'p%@(�fD�v' f�q�B��8D�̧%ޠ��4O/��(�4É���Dz�K
?���4H�	H��S��֎5���Ӹ&Y��ھ_�8�3,V?J�#=Abl\ܟl�I��M�����T~1��@��a��ǟ9#�6�)Vj�O�"~�	��̢CnQ�>�(W�W2$8`�'�7�\���lڊDt�(��L�[Qn�rdE�*B�����jZ�ʒjW���	r��K�]�R�'�Fń5�U�ө�I D`��Tn�X@�iz�R5Kʑ4y�)Cė���|��'�5֧�J��5a"FS�G�n���h-�M�Co9*����א)��u8�B5��>�X�cm@)Ë�k��i��-�&uF�7-�� >��'����"|n0��%`Pl�Yl�	[�Iق��P��jX�D��*�>8o���*R/��Ps�:ʓNT�V�'r�x7��[;�$���C�D[�D���љ>�J=$���퉟t�jp   �   \   Ĵ���	��Z[vI
)ʜ�cd�<��i*<ac�ʄ��i�)m�@x�a�P�mڙX"��xP�MPy�p$eb����4\ ���b��p��IhPY㒩D[���1�N��z\���SV��+<�ɋS���{��i��,1Q�\�n���۰�Թ�0��O���A����M�]��P�#6B��A\�0q���%y1��̅g̐��]Jʰ�P�T��;��|9�B"ΓN:I�A��؉ɀ�Y`����nM"v���O�@��f"z��'j�Ea�DN��~BF�:��\S$�5���#�΄ �~�"ș�y����Q�<�Bf�,|F��P!$�<�L�BPD��<9`6�&r#<���N8b!Yf��oP�AbJP=5 ���W቗>
�	.� �1!	�6�x٢�� �'�nEx2GR�=� :���Z�prHͬMj�oڿA������I�5 ��P��`�x9��KrCr��0K:�	�\D�l�e���Kצ�>jslY� 	�?(��bl�<Ib)<�FI��) HΟzEV�y��*;��L@6*Ԯ�x٥�	/Db�d eh6��#TJ�A�	�Ř'�Fxr�V�ɲ~6M)L�r��r3勺o�
��`m����x�M��\y��R�=�-� N�y%�����O*Q�ṟ��pN�$}�b>JTe�'e�0�`]��*|h\��@�P8g�4`{��Iq		��wEp�S8�:m
�зϑ�4�n�������s5#ݏq��'�04%�݉��'�H9�6�����'ڼ)���S?�!�dދ	 �  ���"O���t)!I<(	�@P�N�N�Xa"OH1B�ks�r���-$THpH��"O�X("͇�%��$�Ɓ]tބ� "O���$B�D��O#�>���"O�B�O�;���9ǌ�<]�Lk�"O�<(Ѩ��\Sl��6�L�7y���`"ONH!E�]����Y�끹���!"O���M�
-��
Y�md����"Ocf	%X$�ʦJ�6l<P��"Or�;%�ݔR�y��n�	�`"O�GEC�.��V(H4SV$<I�"Oԍ��(��ialT
QS�q�t"O�5`C��0�< k̙P���C"O|QX����z|����O��9w"O�Ԣp�L�G���KƤ!K�4�"OZM �'�{1`��6#�l�j"O�m)DO�к ɍ�dc�Q:c"O�YҒ�E    1  u  �    Y!  �'  -+   Ĵ���	����Zv�Ll\�0R�PΓ����I5&�H����O�����a�B䉢]dx�󠩑9b��)ؠO7)�>��F8�:ݳ�i����sboѥR{84�+�0q�N��!M==�N�Jtg���X	B<�,�(ƧNR�jАeL�O��t"#O��hh�d��)S�l���I*(�|IhG�KF�0P�O�A�l���H�)�0�q�[:e�gʉ5,,rP����%U8����'�2�'lR�b��I#'�0�P��$!����@�S2�x��7�B9;��[ lu��2�)R=#��3�&#δ@ �~F&e��`��<q����M[�������E`���(Oj)��L>�N��BQ�*�X:bU�8#e*�Ob���O�㟌�'9S�P�ȅ���	�jJ4�ȓBK�hʣ���rx�`�)�%P�mZ��HO���O�ʓ~a�� ���m�0A�Q:��iZu�k�`���?A���?�"���d�OP��b6b8@��ֳ����ʣ6x�;%���j5)���)v�|��
˓>T^i��`�@�S��	r���`V�
�0�Rr,]8{d94�'�a"��B5�����,���r��:�ժ��i!���&�禙 ��5�1�����Z��/D�thug��2t�#S�EK��0�>�a�i<"Q�|�v�G���	�O��S�.���͊*a�օ�e�<��6����O���Yν�CE��%n��ԟ��8Q ��#��y��c̜ct�LH��	�^P��ye
E `ִmy�!�D���̵"9�D�R�G$��Ѣ�*�hO:e1s�'cB��ҊU��<��CF�7�����<R���|��� wщk5h��`�S�P��Y4I3�O�l�'���r`̶n<ցyAV�k ��O��a;O����O&�' ��r���?�$M�L��Z3bӿ;�2�8p��!"��h]�db�T>c���p�**�yj��\��T�SJ�O�ñ�)�J����}ܼ�f�HD���je��	��S�O��y�s�H'�L#lF쎉��"O��jS�4Ӹ��Us�*��b�	��ȟ�* Ǟx����&��6�p ��"`��h�Ó
:*a}�o�o�jH�F�2ւ�y�D���yW]@t��&Q[�":�yr�̽N.���L�,ov�j�L���yRô!�����0xdе3�!S�<i�'$R�$x�5��l�( �N�n�<����!��%9S���c�*�/i	JC�ɵ2�Y�o�0��%q�	^7+��B�ɗx�8制�/Vu��F���#uvB�*��j��Ł~�ʕ�h�'q.B�Ɋ�^� l�*¢iYWɇ�DB�	eI �
"��T��I����@¦B�I���U�)	+^m��pT��#a>�C�*L��͢�H�>Kn�ٱA�D6��C�ɹ>��T(EJl�3}/�C��1\�FM�@/C�g8�)V�V�j$@C�I�!o�\�`S:^�X虃/5k�bB�I�EM��q�߅z@X���G�?'�C�ɽu,�)[3חnU$t�"�/M	fB��AP4��+��9�ܫ&.�)�,B�m6�]��H�\.N�+$�l� B�	uT`��Z�2�uS3��ZS�B�<�����`�Rb���Gb��
�'�6�8$/U�$���s��:>2u��'�NL
u��fS���Ҩ\1HӲ��	�'���@7o�9�\�8"i�3���1�' \$Q��<;�1��K�&�^��	�'
������(3��D��ǟ[sE��'w���H�N�0�1�̃R�"=1�'�<�#+5kv�۠oݺI�9��'�*I�t+/H��x �M6��H2�'nz1E�Θ�L��c �W8�c	�'ɮ��MW�l1T.ߐY*����'�P�����d,�͂g��.Wf4��	�'ά��Sǚ=C9X	��J]>W=6�r	�'㈘���P�x���	W�,� 
�'�t�cLM�p`Y��մS�tĲ��� b�J��ƾ-��k'���v�BH��"O���i��4�2dաQ�@�
a"O~��pD��%��tӡI�%
$!��"Oby�sς?���9F��#҈�"O�iҁ��0z5� �O�`:�i�"Op���Z��)����+*"�P9�"O�us�[F����p\��IJ�"OJdq���*/i&}SBL/���W"OnD*��	9<�5�v#E�C""��0"O*��pK\��䰳�
T$h�0"O���j��r"��CWc�� PF"O��ca�[�YK6ҥH�}�x��"O2]�S���M�nU0O�~}$ `"Ou;G�L"w���{���VN���"Oj���Ԣb����q�V��"Oh@�5d�m������B�6�8�A"O��i�/�HR�4�� �&�݈�"OZ0P��K���qyv�R�@���+V"O<��`E$Y�u��Jxi�"O�t�s��X[��Y�&��� ��"O�P����'(��U��K���8�"OBQj��/\��pԄ193YH�"O�Q������W�6�te۵"O��G�5��`*g��3�ؕC�"O"�R`��">R�٧��_���"O�|1fƥxƲh���K�.��܉$"O�CRN���L�D`�3L��aW"Oj����L�d�����]8;���a"O�pP�\�a�r���O��!���&"OT�6��$v�0�(!mѬBb("O����*�:����[�����"Od��#��4Q���7b�} ��"O�M���s�����g��e+"O�A7�C�@�%�qI��z�%�"O��p�e��2��JC�R����"O
�Ta M��٥�ٽC��4b�"O���t��z������_�Be���"OPx���^ 5���%@ւ-]���"O�ɢA������H��=A48i�"O����M(0��$CP��Yr`�w"OZ��g���V��H8Liڵ�"O� ��	,p5X���E�t �9 �"O�0�c���ܘv��'9a���"O�` 	�� w���5J�:q
�"O�8��#�5�T��C�u�bH�"O���agɈa����.
I�f�;R"Ot)����^t�<�lބaL)��"O�M�b��[�bUꡪ	f4h�"Oh�)�7!�6�*�L. A1�"O���@KΞ�Pm�f!P�z�DX�"O�D�M��C7,��p�Nꄘ�b"Oh�K�@V 9���;3*��~(`�"Ox��7�B�K��@�/�dcn�$"Oδ!R�PP<AB��v:�1"O(��M�H�:��c�]-^>��u"O�1S�I#t���u�τ	K���`"O�̹�ڀ쐝���1 ��x+"O������{��}��n�_�<�rE"O�����"O?���eM���0Z�"Oh����A�҈e a��K�|H"O�â.ȁY�,`�P�&MZ�j6"O
�BiƮ\d�!��I�W�\���"O@��� ǰ(F-��Ҹ�j<3�"OzB/C�d�dZ�6J�"O� q����}���Ud�=n�P"Of@��Å�U`"i.gdb�C�"OҘҁ�K9&@��soD�dZ�z"O
 �UNW(a�B���YT&��"O���v�P�,P��1"��� ���&"Oj!a4"v���$�ڒ�0aa�"O^x�J������a�B5X��A�"OD�3���{���c��[�8� ��"O��BE�Ԍg&H	�V��g��Y q"O��(�%�:Me�C4oU]�^�w"OX15������-�k�蘳"O*�SDd�ZH�����Є��g"O
i�CN�R�ؐ�bB�l�~a��"O�ؚP+U�m��A��h���s"O��`mU�4��9@6�* 10� �"O�a@w"SP}�u��k��#L۲"O��q ��4mQP���Q �m"O���c�ϬLoΥ� [�sj��"O�E���֫>���h��Ø�B�Ҧ"O�	zs��!6�PS&ٟD1t��v"O�i�����%U�z)`t��"O��y�g�}�:�u%��y .��c"O�}k�IU�H8�x�≽�"�"O�af��!Zȁ�O��{�(A�"Ot@�E�ҿ9�B- Q�.��z�"O8�BЌ	B0:H�"�=(�l��"OB5�����H#�(q�"O��pJ���`�l\a�d��yBD��>�R'�׮)H�����y��U+1lr�3c��Y4}*�K��y*��a� � ��nI�%��y��^%X�aC�ń&�NT������yb��=O�]T&Q�%�|��@i���y"�Hf��s�]�,�l:3@�5�y2��	2r��I�,/!5�Y��J�(�yB�_�P��R�l�&V��+�E�y�n��L�*}ZV↸`�H�z�k[�y�@�-N

���!3h	�#H�y�
�p�V�C 	<0��Ń��yB��&wy�<�e�q��yDm�&�yҋ�9+3|�����7K�y���&�yV�/" 2u��n��r�Ȩ�y�c0D��!��)R���p�� �y�A�a�`u��OX�0(.�(�@L��y�+��Z;��qB����B+��yB��d�nܓ�鏢oҼ �I�.�yb	Y*�C� �bH�M�r����yr'Z&jK�#T��ض*BH ��ȓ9�8pq� �7��)����\����3��X�HT�q��y��&֥�ȓrц�+�k�6!�&�Q2(5M�E�ʓsl��Ks[0��J���hV<C�Ia�8HK��ȯ�	��k�j�C��fZ��Ћ��P��1A0.�< �C�I�]�`ȵBɨ-I,l2���00�C�	� �RlE!^x��"��&��C�I"] �R!�I<S���ɀF�X�bB�7J� �D�����	4�>X�B�> q���"�Ӏ]�� ���:DB�ɗ&B~ykf�'}���@/^�O�C�ɘU�j��wL�.?�,@��zXć�dҲl��C8ˮ]��R;U����9\��4Ô�k�9:��6>�=�ȓ�h�J�)ҞG�!R�a,Y�8��S�? �I[aI | �  �
�����"Oҵ2�1�0x3�^/.��z@"O&����I�3P�y��H �q�P"O4�j�m�+DI~,+PL�*4?^-zD"O�a1���c�y��, ���c�"Ol���P�X���s`,�1X�P��"O*	w+A��j�Ag!�FOV�;�"OZ)�E�{����bၰN� ��q"Oⴢ��Gfz���JFiP���"O�X�v`�+$x^�����4)WN�U"Ojy���sG�i��جtL�m�"O��B�ʫ3�1Jp�z���U"O�L�p�#���bD,�:��X#"O��R@B�q�<Q��� ��T@"O�ar0�N�*�y���u�ؐ�S"O`Ļa��>t�,��/ )F*f%	""O�@�`��Y��{�nC�](x�X'"OP����'SVX#���\F�$�"Od!(�c068��׈�B��Z�"O"5���W"!����Ө	rB�\�"O�� &��Cr*T���̂ܬ]�V"O<���K�<�~�;� 1#�� �"Oz�+T�s�<��U9��|�"O��`�c�/]��ʑN�3�`��"O���mP�K��ͺu�O!��,0�"OryT�\�4`2Ӡ��,��y�"OP���-
��<�"�"m"B�J!"O4x�C&�Z�d�k" �	�e�"O:�Y��-2l`�u�W�E�*�"O����n� �И��F��"�.4��"O����#ԙW�Dx)УT�~��$@�"OP� ���o��VFy��A���%/:h�$|X� �SŇ���I��
/�:}���%D�L�	G�>�Ф��gѷT�!"�)D���1�!�����ΒVz��)��1D�,�� W�B�+�ט� ��.D�3c���ga�iy!�ũ/����H2D��u�;x��c��;N�6�[I"D�{���vԀ�4˄��P$ 7�>D�����H��� *F�zD< E=D�a3l(Y�����Ŗ H�q��&D����猅+Т�!0'�0#8� D�DQ��ZSFJ�1��0KP(0!֧<D���/@(ȵd�����Ԡ.D��� hM�L%�)����	^���@�m9D�Dh�M:0��Ӏ&ɵa����r�7D�0&)�X�$3e�=U~*��!D��(p��yMٸ�T  �6<��2D����	�G�P���)!�,TC�//D���
ʸ1���I���.6��u�'.D�舠bT#'����qV+.ܕ3f$.D���@�0p��J0NS�i߲�1q�,D��؁�]�Z[���� &*�YI7m)D��k��'A�^�z�*a��)7�&D��,N|�>E�t��brEK�7D��3�F��c�>)���²B`�PJ6D��{�ďdP���B�2�m�" D��eX,2�"��1cUz���=D��4'I):,�p#�Ҫ-���m<D���cD�*r*Б��쎞p����b5D����Ό^���4��^)��$�4D� K�FRx��Tn��mg����1D��E�)Ǯ��W��|��R�0D��2W*�V��@Ă�;VyBć;D�� �@ӕ/�i�XY@��D���Ż""OЅP�.Y5I�4�S�ٖu}��1v"O:5�� B�)�x�ycO4"q�Y��"OJ�g�=i+��"w��8~����"O�$��ƕ,Ag��&�<QBT�C"O�� sj^A9A�Q)J �� "Ot�r��OrB�#u��8C6n�7"ON� �L̫]�2\��
�;.e��"O2U��Uy�	KD��C�=�"O �zp�Q`0.ECr�G�A��Y!"O`�u�5�F91�� b���"O���+X�P����Ǐ|�>c�"O2Q��^��fH�vn�>Xi�p"O��ٗ����|�L�]#R��$"O��W@?&(�=x�阄!����"O�šA��E֬z��]W�=�C"Oذ�_Y��*S��2��Y3"O�Ńd@
 �|��B��� "O~ɲ�m�r�� ����tS�B"O�yy�+�����u:d� "O� j���}i{4�L�Q"x:�"O0���'Cԁ䣎= ��� $"O�L1�Ƙ/�pAH-ܒj��Pڄ"O�s g d��؂���Ip"O��аƕ:t� ��Y)I���[@"OB�Z�$Y&C�(ᒀ��	�d���"O�SA�}�H�S6�	Y�*���"O�� �0eZ�K�(��~�)�P"OV�ziT�c��P�����\�B"O�e)�e�\4���R"9R��"OJp��Ƙ''�D��CD�:U%�B3"Op�4)I޴!�1.^�8��#�"OF!�4����좦�����
"O��� ��`"$���A֏ꈑ�"O�x����<P��Ԙ���L�����"O��{7΍"D�Y4��e��u�"O����#��p��y�S$WP*�"O�E)oնI��x�P��/Jڑ�S"OZ��dV�4\*�3'¡P/��Ɇ"O�%�֢O(Ap�PU� K��P�"O�+0AW�yL��B$�by`Q"O܅J�i��U�-S6�I�\�4��"O�UQ"(�
-cAݑA�L�"OP蔁]rJ�	3��U)*�r$!w"OLIR���8DX��
JƌP"O
�qP�V���P�q��>��"Ox)	C��2��y'd˾} �bS��O��(O�'<��1)�kq(9d'Ze��ȓ|a���ՊQ�o��ER� 	F,��)���T.Z�e;��S�&JR���;D�H��C���$Kѯ�.t�TF�������gTuiЁ��fn�@`3`�2!��C�I�eX���������	βB�5�jEJ��G�<��B6�A�7��B�	�jT�`1P�*C�@�3�ɀZibB�I9b����P �:S�*�R�.	�~VFB�IFR`嚆e��1����!�T*B�Ipybp�W�ͥ8�����GE��0C���>hK�*��]�BT�����>�^C�	��x�!D�f�xD闆�e�@C�	(#��rc�ݮ6�f��
�brC�I�D�����8!L8P� �!�C�IB�^M���_8oN�#�"[�2�C��# V8x���<3�O���B�)� ��as%B�[�0�Qƈ
F���D"O���&B�$�8����F�Y`��"O�H�c4 h�`�� �[Hh��"OBP��H�*���Z��E:=�v���"O��GE���<,8���,K�֍G"O,0��M7�6yP��*+f� T"O�!��*�HxH�s�, _��ʤ"Od$��,�v��H�cC+t&���"O�}�cÎ�Azd��� 	�"$ �"O^u�4?V�t	!ɟv�K��yR���n�0"�Mu��ۼ�y�/�}�d:ˁKp#�lƉ�y��6^��(��F.��8�֣�#�y" ɁY��dw Z�)9ix�IŔ�y��	��L�c2�H%�b̹��y�+�6��i2C��8�|a���yBkS����ƙi]��xb#޲�yҠ�%k�T��)� b�F��Ĩ@��y"�C�.�E��R Y����s���y�)M�V�~�ʗH��=4��A��yB�DUH$M�	�>ߖ���+�#�y2��%K��D	�\�.aa�B�W �y���8c��ɩq�0}yR(���:�yb�Â5��dC��X!J�&�x�����y�ͧ$�rA�"�K0C|zԓAh��y2�X�6����G�N����ዦ�y�IڲR�P��]s.��P�ʗ�yr��r��Uy$�� 4�Y�T�S �y"gؗЈ�1,Ǖ�4��#��0�yD	��f�qw��$z	��C�?�yR��kcf�a���a�`xæ�-�yB�[�^��P�
\���3S�J�y�aس�����+6�8�f[��y�I��N���CU��|���3����yZ���@� ���$�1ٲy��u@Ò���7C�2R|�� ��RJJX�6�%hh�(�gN�"XvI�ȓ4�j1� �eU�"סЈ� =�ȓV\�5�±?GnM�'�N��̽�ȓ	��m�q�!O�x���g��E��h��_��{d�0"��0F`�:p�ȓ^%y�\�.(���5N>>q�ȓ�2�I7k3]?���/ֈ�e�ȓW����a��1֖� ���l �Q��x �}C`��V���� |g���ȓ{��d��0��B�K6| ��j��#�:Gi�{���fnP�ȓ2�u���آ����"��N$ḃȓ`�r!!��:=�� ��0wŇ�-6��Ig��)��%"�׊bޔd��-p09q,ΞL_�9�q��;D�D�ȓZ����v�X1=����磓� �ņ�^���Ѫ#a�4�#��)����=Լ����,a[v`�S��cb@x�ȓI�H�[3k��e_����#�T���ȓE l$x�$s� *p�١j&l��C>��� ƞ$������8gp 1�ȓ`�*9F�4�����A5Z��t�ȓ���)��*=�@�6����܇ȓ&���`lY([M���� '�����@j�1P	ܶ5*��E���#,���jِ�D��H���� v�xi�ȓl?��	���K���4�C<e���������I.3n�) �@<1�v ��S�? ��S�kF� ����#e�"���9�"O* ���@�E�\8wB��A�T�a"O�H#ч�Cn���̒t�2)
�"O���%(�J�9R�͎)_��h�"O|M"�oT2� �Z��ܙ$O�)�"O�q3�)�97�^uI�Oȍi9B�""O�|I��!��$ ��%9�t�q"ON�����8XN2����!o���yb"O��xqL1d��+���\�l��"ON��0�ڇ!$Z�:b+�;&��#!"Ob�S�ާp/���TsE���"O�<a�%ޝoZ���.� 8n�h�"O.d�t�To�8�Q3Q:h��"O�E�gJ�� �Z�GB)P8��"Or�9"���ZK�%�C&Ug,���"O�J��"#�.U��%�+���"O�!{��ւ"<^ܫ�*98|��ʇ"Or���
��Q8��	��Xt!W"Oĭ�vl�}�qXe�:��t"Ore#�I�9Cڼjp�J�P�.��c"O8��ώCq�ԣ�E����@"O^5�BÚ�_/����X%���a�"O�qNݦv6�@a4��v���"OࠈW J�T � �1S"��"O�[̊1\(���4`$p���"Oru�v�]5MEP�MN6()�"O��q��(;L�Ƀ�ٜ#�0�A4"O�<��n��JB��"��U�a:�mb "O�B�)��C�돪-�)�"O"���N�!�^���l��sN �"O�Y���R<Z����"�_4&p�ha"O�1P䙲6g4u*jm��Y�"O�I9��U=���i����)�f"O��P�W�x��+�Z@��"O��x�n�+<f�@�c@�Ch$��"O�s1+ՏhL8H5BD9M��@v"O�%���  �P   T
  9  �  S   �(  �1  �7  +>  �D  �J  Q  HW  �]  �c  'j  jp  �v  �|  Z�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl� Kp8O9���'�t��oŶL��5��m�-qbK�qU��� ��)U��ԑ�C�4Q�H ��Fa�U�@	�?!�I�?]���ʙN>~x�*�32���D�(����j� �5�@L��@u)�F6�]� �������Lre��r����%��Jް�
�"Z;X�P%%Ɉ�?Q┕d�\Hh�n
�*S�f�ɐ'!��'�"�'M��S*�4�t�7~�Òǎ&L���'0V6�J��v��?�U�ڿ�����?���L/O����t��&Y���QU�?��F��Iϟ��������,?�'ǚl�t�ؙ]qx,��#�dz�z�'��l�5"	�f��$�¡�2��ҭO`�U�Il?ѓ� ?r��'rJ�ZՋ�/�"%!3��8|)�	矐�	֟��	럄��矠�O����7=z�T���H����D	I�M2��h�R�m���M�w�i)��i��|l�M�q�iyr�O�}^���b@?<�v�I�K�;md�"=)�I�O��qӅF�QdYHcn�:���cs�\7Q�9�SB��6����i�(7M�Ԧ����|�p�/�i�fB����}��X�ݟP��@�P� �3��˷(ұK&m�zıQ*¼�M��i�7�B��1�m�,0X����a,zo8i�t�%ژ8��Ř��m��4��vi�m6���G�����{ÇY�/�1�v��7iؾ9�瞁Lb����L�n��X��#ʑQ��7M�Ҧ۴\�M�Fg�(	�4`ҤE�TӬt���U�AE�u
�Ũ};�8��0L���C�6N����o�G��`F��(?�d�	a2�@%��#�:|�� S�=���$#�	����Ʉ#"m��4�?���� �	:V#����  |(������?����?A�����kD'h���x��@M(V���fe��1�R�Իr�j �g(��0�'�Aj��H��05�� ]�j6��/#{"uxk�&J����1��jUaxR��;�?�����W	e>4�V"̓0뾴б��GKb�'1���#R�P\�wi)?<eX���E,���Vܟ�KM��D�P�B�yv�4��OV� s`�%§�y�ĉsK���NnDl�9E�-�y%L
i� �
�jj����u	Ā�y�g�v�ҭ�U嘰PI��{UK���yr`B)$����1�f�;Vk�y2�!����J�K��J�cԔ�yg
.*�H�7 M��R�(�ü�?U�T{�������tK?�8!���T��&�s�)D�@J7�Y�K	X� A�P*H�
�0�'D�����ۍL����@�M$)���bp	;D�@� `�Et��ّ�Mu%�����.D��H�ն�٩��-Y&f�k�o+D�l�S�]3)8X(x&�>K�*C䇳<�VF{8���Ü1i�%SV��..���E%D�\������J@j���b��#D�HӐ�3Ӥ R���)��] p�"D��q��C�?�@�v�&;�Ɣ �?D�[fcƚ_:ll���M�-�XiQ -:<Ov`�uEMצ��'� �F�ǕqK�,�cޡO@�e����d�O<��O�1H��	l X��.�S�|��I�u��$	�NC�d�RX�#W�;����$ �@n(�"��0)�Bm����O%CpB�1�}	s�#���"�'04����L��Flk� �D���h���iX	�(��%���?!���iU(�v��rE�~@����F�����O���#�&K���c�B0t���Iz�I0W�Q�!�1�s���;M�`��K�&:IƬ ��9D�JŇ�l(<	�����╘�A�7lZNȅȓk��u���N�C�|� >n��\��7=N`��S=i'p��1b��q��ȓ]Bp|�%�Nx0Q�.ڶso䤄�>
��k�m�4K����G��o��Ţ۴��k������?����?9.O�9�T��3EG`��U�'�Y�"fԣvh�R��惡ʠb�(1 �O��\�G�[>l�6P��F�\��U0iݽG,re�e�O(Xl �j��!�c>�[���)����pN@;1'٫<�����e� �9Z�d��E�	a��t���L���ߢ�&�0�+G/d�@-;�c�Yx����O^�xX��Њ�%V�x��`����Ĝ�Yߴ���|j����d�by ����:~Yj�`�K�xB�A�w'�E<����O����O����?Y����4���3�p4c�;]:�J7�ߤy������(%�T���3�0=y�f�$�����ɕ� 	@x��b8&ixq�{֖�k�I^���0ua͏av�L��n��	��D9���64���Ԧ��'���'�2�'w�?����]���Ì��\m�GH D��z��V���@�+V
y��JR%4������Ly�#ܾyO�7��O��$ ��=���Ø5Մ�QD��X0����Ox��T-�O��$r>!�W�O�b�� ��qbm�
Wa�,¥#�&rp�����'��+���Ղ�T�#�JP�k�<��&F�ax���?���|�oʍl��A+�i��^N�剳'��y�ǋ<_>Jy�`� Z��9��
����?�'{Vq��瀆SR(P���7���I>A4��4����'O�Y>���˟�	�
ׇ�>D×מJ�0��QiZʟ��I�U��]�'l� %�dm	���,�.���'x�)�2��q��A�ejU�'�~������f�P;��15T"}�ϕ/Og:P*P���T@� 2�X~�7�?y������O���c�H�I󈞆UF��J>����0=�4�O+8H�QB�4��d�ŠMZ�'R�}eHNd5Xr��\=r�'������O��$[���E5$�Ob���O���i޹�C�%j!���G;,j U"�<��*�����0<��m�<�x���Z���SEED�M��P��� �� 7̏�|#�|�|w� }R��k*��"�_* �l�Pd���?����?9���?���,O��Dٸ4��!ף߫6
�W�Է��˓P$�G|��d�)T��IIA��2v�-�Fj��X��I-��$�Nf�d�OF��Q��O��'0o�Y2��ԹH����W/h�Ա7Z#.	������?���?!���.���O8��X��Ã��=�4�5�C�$(.�(BL0��ʀ�C��b�&)5)�)��O��B�I	
�k��T#~��a��265\H���OP�6�d�O^�?�	*85h�T!��|���M &a�ȓ.7h��T&�d��afЊ Zze'�hh�4�?I/O8��s�$�'�|��a�%a��x�!Oާb��Kc�'2�9���'��	V=X�&(� ��/F:x��*����s#`ٰiҪ<�7%
N@@s�*O ��cܥ9>�8@�'9>]lZ* n�D�㬞���QbA�6Mt���g�"�'N�I2R�&|H��0򔙳3H�iO���!LO�=���=,�e2dfׂ?/^ [��'���9[&xp#d,��I�=�u�O�Y��W�p�&�X��M����?A/����0�OVL�����i�2-�^�B�J���O��$_��|щ�쉷t�v��$@?�M�O �S3uX@5K�-F,V�xP�/{�P�;��2�Bm��1CE�E�UP�>]�e�&j�(��E�u}R���O��zP�'�����T)�*�h�q@�&d�^TK�ǄW�<q��Y�z1CV�V$;Ɲ���O�'���}�Ef�� �X!�d��	0I9���M����͠lB�i�O����O�ʓ!a㐥Y�w���І��N0��bt�T�<8B���'=������Ϙ'�2�b�B��4x�1�0��	�Z9,��TH��:��'���#m���Ϙ'.� kf�E=�48k�/P�#����ğ�g�'�ў4���!��݀%K��U���V��l�<a�.�-�P�÷��.O��A���hy�� ��|����DKeh��B�F<x2�t�3|o�� e��O����OH�d�<�|gf��#/K�F��3)��D6H��*\��b�IW���y��Q�2K�����Ԡs��F��T��G"�
�J?~���'#�|���"Ġ|��螩p,"b!EN�?���hO�"<y���
|������X`<`��Ey�<��Z/|`�y �+;@�K�Er�ɪ�MK���',x��OU�C ����+Djݷ;�����'�l����G�#Gϝ�2y2dk�'y Գ�ᝨ4 �q;�i�#։x�'J�Аd��6m$��e(�*�� �'�x� h~tzeC,
�E��'ނ�	�� �R����8b�t���C_�Q?=z[)C*��M=ê�����y�[�w���C#��>�tQ�"���y��ˈOr�A��'ր1�� 3ß��y���
�p��ଁ,-:���Pǿ�y"+N�6��(�	O�7���!Eԩ�y"��c^l�1��\��� m���?�*Ya�����u�&ݚL�jp!ӧ����+,D�Р�`D0�|@�5G8(� �2�5D��qM-�9[ �B#W��a��4D���$ �"f�0��5:��v#3D�8 `�ޜ%�
��2O�	�*�*�0D�D[w
�:z�d Y���/���r��<i��B]8��j�H1`�$93�ގ8CXT�h*D�� =�qF�$��I#�Ck��it"Ov�pҨX<S���y�-��U�� "Ol��*�pN��{`.��d����C"O:(��G�T��=@'���^��b�'�xI�'f6�q���.���z��l��L	�'�|�2��܀o���,×]͒��'ʶx�W�@�|�[�LQ(PI��'*td���qAlyh�iQ�t�f�Q�'��ႃ�l,���@�km��
�'D��Qˮ&n(�E�ŒY��M����.�Q?�������!ӌ�^�!�H#D���1o�,�9ڤ/ R/8�Q�b?D��
ï6ڤ�'Ϛ�X�h�Ce >D�8��)?;׎tٓjW���� 1D��KG�8��M#�  2D����O.D��C�M�@�l�b[/j��l�O&9�#�)�'6�,`	@a�;r:(1����iR��'J�C���3���?^��	�
�'������f��-Z�$c0�
�'8v q�Եx��@ƃXF
�0 �'}S�,X%A�,i��m�E�$9�'���S���5�Ш��B@�8Wr�;,O*U�T�' ��j����1߀x����0�¸C�'C�I!� 3z�`��t�	3 R �
�'�Θ�W�M%"XHx�Q�q\D 
�'�h��*�;.�	qd�Y�j32M�	�'x!2%)o������|ݲ	�m4� ��6ή�����83O��لH�h�ȭ�ȓaݴ�G�_�3�X���ʂ`����ȓ�J��AӬFw�u�©�4^�ȓ.��RO��~�bmi`H��a��d�ȓLyF`@F+���t�b��T�����~P݋�FY���E2�8_r��F{d�����(���!T7b���Ř{�j��b"O��0��PhJD,0�%��	͛t"O|�q�jڏ"RZ�P�� AR1�"O��s��ۄqW^�rw釫a�y"s"ODh�&�b�t�L�(N���"O$��b���(�4fCy'��c��'�x�
���F?d0u�Q7[b�`f��	,�<��7ֺ��(�0kvnڠ͏%m� ��|0ݨƅ�s�vh�ըߙ"�f��ȓEܔ�#͘It��th�$*T��ȓK�&8��ʖypls�$�z��ȓ
�����l�j]�`c�,��\p�ݗ'7T�r�Y��=��,�d����v����l�\����f��1p�ښj����vQ���'�:d����oR�g��I�ȓIZ��S%GLPP�F�W��\��cX�: P�1�QA�̛:�����	$Ecx�	�;�! %K�CX�T3�J�mB�	�Dxh��%�DP!"+�*chC�ɄA\�@��͒�u���Z�(D^؜C�ɞ_��Z���!P:�+ ;_�nC䉓����ț����vIR�B�I#4�DlCT�U� Q�L�چ��=�'��E�O�x�"�M�9�f��q��*�c
�'uP���aS1;�Z���=2�JT�	�'�X$��oAXl8�$D~��	�'�pt���мƭ��(ҽ���J�'���)�Fن��q��L�;m��m �'�@�IW�,`)�M�F�H���Fx��)3�n$�3!Ȁzʠ�A��.YC��1:��0cR��X8*�OD�w��C�)� �1��Ȕ�f��%V�$UX�@�"O������gl�X�������;"O�(��/\Oьز�n���h� "O�)���2`�4%�����Ȁ�S�)c�(�O�x9�� ���O�aJ@m"OxQ��C�Cq�Œ��G47��ZG"O>y(A	 �&�|� t��!��i�"O�4sS�W8Ħ00����W��P"O`�G�ܪZY��`��Qv|-���'���8�' �܁��]*{�I�U��8.����'�R���nލd;rx���P�9K�e
�'�8���Ǎ�r�.UJ
�1͒�9�'�HQ�
B�
|0x��  a
�!�'\�	�ՠ}E����Pl�u 	�'��4ϐ�w�����ۤ8�05[���>]Q?=@w,ҵ<c�i�CdͲE���1�!D��B�H��ay,�)l�e�j���	*D���㭜*gyr����_�)�h�3�J;D���
� C�bp�f�+	d����<D����FY�Y��d� �[�L�(R/&D�0SI�Ƭ�'�S	�!�Cg�O�}�G�)�'Wt����?7Z��;3-]8r��Aa�'���jьP�H�K�O�H���
�'x�5[�h�%Ym�"�J���,Xk	�'��� �PVT��i_1�A)
�'> ��e\��⍙v��?Ѹ$J	�'��X��O��s�\M����;�Dm�+O0؉��'�∫V�e��)[�N�9�9�'; %I�ǌ�*�d�)ǨQ�;%Hԑ�'�xi3��&8�1@��75v���'�LXxW��"2�ٕI�:8 ��'�	"4��-+�h��J<N�|�	�e�<��{3ᐮ��t�[��B�Ԅ����P�ǌ�=j\�(��L�6I`b�Æv�n�F��vӢ���q�V�!	ϏO�P���	�A����ȓe�dD
�I�Zp��g_�x�ȓԞ�
U���>#8��Ć=s1G{�C�
ب��I@0	Ȕ&`�峁-D�XQ\�%"O��x�(6on�d��%I�s+恈"Oj��""��(�2��C��#\��q"O�YraZ�g�2��V��%XF���"O�I�d��_���+㟘hc|i�!"O����b9�Mz�"ٮT+
��"�'@.�ۉ���/:�u �i2GT��`��	f�@�ȓ���qNǝB��l����B���ȓ  9��K�8����+&�n-�ȓ?w�=h�wNm#¤��_?���ȓ`�6���Ń�!{�Bf��%. ̈́�A�����g\Ȟ�Bw���&��'��܀	�d>\�A*��r�$�Z�,�[���}
����:�|E� �y��<��0iv-�o#� ��QD�
\>��ȓ*�ʼht�^�1�"ȳ��G� F����K%�|Hb*޼-�"٪�A�)/�؄��8V�F��>U��t�U�¶	d�bb���#YLB�	&k�X��mB��tEK#O�&��C�	�{�h��F�4�ifb
2Y��C�4	��l�W%Vh��*9Z�C�ɏ8Ar�6�LaNy��O�B�I8J��
QD�8'���83��81�N�=�f�Qm�O����A�^7�v�����"Oҕ0g�G�EY��9�"w��@�"O���s�\�>m��{ ▢q�BP��"O� �%��"��iQ�DR�㙪Θ��"Oڼ�b�k�z!����7TO�q#�"O��)H@����1k�1��P�F�'n|�����S�(��9K1���v���"	�ȓZ��$�g���A��8��ʃ@H�T��������V]Z� �En�*)���ȓF3��K぀�4O��SUb�NZ���l��Mkr.ьP&h��$\Z�4�ȓjc�ӄc�:��V��q�x�'��k��%�Pd]�iaH���%��lp�8��;�����6��I�����g2D�ȁv�Y�>4�y���D��]j��3D��Z��ҷPZ~��щw��UÕ�>D�8"��E:A*,,�s'�30��p�g�<�O^�R��O���w,BJ�\!r�LC(X�\ �D"Ov�4�
m!`��G<H�l��"O����	Q�ڕ�"����{�"O�՘0�ͻ5��H��@��Wn�[A"O��AC܈h�0��B9VG��IW"O�p۶�]�oZ��jal��Y����_#H�~��S�r����� N�;�|��%�c�<��c�H���	�(6E�X#��_�<��	":��L�Ү�`�RE��h@Y�<�a͵R��� eBǽh��哗��y�<�G�gf���EZ��Q�U�t�<�sE_|D�ݻ��ل%.`uRv�Q��;��'�S�O	�@ `���'<�(I#���t:s"O|5�'�Vh$�(R ��(�<pC�"O(�C0��dBq�@��n0r`"O��*qL_g!.0�J�,d�m[�"O�99��
�U8*(�B��C���0O��[�NO� ��a��#{���m�O�'�����'�y��П�ρ!�VL���"sv��2������gb��l����/+z�YB��Չ%���#͟���i��ک.�"YQ �%��#>���W�Z���
��G��/�6|RvCU�\6�� �I
S�lI��	N�.���OXc>eBƭ85$b�P(͢�F�<����@�ɰP)�EرJ����	��$���4�B��ɒ m�P@��P#��I�e�氩�4�?�����;q�$�O�Is��H���ΐh�,���O h�ǉ4<���j^�IV$��|���� V&�A��
V7uZ1��B��yb��{üe	0�x�� :s�+T�-	&cЬgA���  Q�>�H�	a2F���Ov�S�b~҉��/�Yr�$���uc3�y"��P�b��@랲�xY�����hO`tG��_
FK�4^V��A��Ys5Oɟ�'P�9u�'4B�'��P��� �v]۔G_4<����7�@	��#��� ��H��`�4Fx#V�R@l9��>����d�FwP�1Zv�'A�0��� |p(�Y̟����gC��N�)?ve���/?%���$�	S�'O�D��n{�|��@%.�d؃�)B�x5!�d���~��G���DT��eA*'��8��|������ʌ=[���(�����c�'#H�t�Pa�OR���O��d�<�|�e���<k&��⮉5%��H�CΔQ"�8��*3��xz����y��ַ���d�� `�#��_���o��s*�h1�['5�y����?�CL��VDUa�D/wѸ�@ա�?���$&�	�6I�&#�&.`sBU.CTp��=g0Tp'��OAb1#�c�A߮��'��6��O�ʓ^��C���Km���45�B���� KZ��?���?��_
��fK	�b�XKG�����H�(�"�ȇG�B�t�)��^��O~���ݿ�<h���
�\�'�ɑr� ^�t�B%͛t�,DD|R@2�?�����O1H��lOW�@���L�b�d��/O:��c� G�Tx�d0��V&^?�}2�<���A%{�ޭ�d��8
���Sy�F�hUf6��O�����O��^"+�4���S�s�jHS2.�@�D�D�,O�9KtN-5�(h׎���"~R �mYʁx�l҇_\�Dub��<Qd#R`�f�����aK��i��)���`�d�v"�(�g�ʨp&���/K�'��)��8?� (�	@�6��\�5C�p�F= �"O,˙
n4�w�F7H�Z|���ɼ�ȟb5҇F�
�v�CS%�3��%�3G�O�ʓ|����i���'[�R��WU�x���'}-� "'�%s�N�ƣٟ0��E9D2��3�H8Fx��.`0^ԻÓ&J���3���Z�fDsu�'c���'NF�T�\a�Ο�|;w�ʨ%2�F�!{�� r�%?���ϟ��IT�?�O*D0��YY��5�<Ӛ���'4j� �ۈDz0�Bp��<�����O����|�'ى@[�=h� �f���(��ё&�J�r�-g��'x����'4ᖄ�Vk�|>�= �)E�1.�Y �'(�ČZ�ޑ ��`k��'�\v����ԢÜX�y��N	��`a��|L�h���'��`a��e��2!`������1RΔ�0���hO(">!���	���p'�]5o��s�j�<)w�����r_
(��Y��IEdy2�w�P�Ĺ<Y��@9i����a�� O.[4,��$E�o,b�j���<���?��>�.�PMz'�h�mV�_��O|1���\�z�D� �+U��l�h��dK7p�-J����9A�C��|�`蚳+9�ĺW_-[�p`��n�'
]{���?9��4ȀH������=&�l1�6K����O���d�3%�Ҋ�P\��q��}Bd�<�� ��qY����*h����d_Yy��'��'2�^�&��*���!�����B_^"���	A�'GH�@%N:�v��,lQ��cí����O ����>DU
����ٸ@��O���غ��O�s�\a�Z7m�P̋�j��l��xC�M
����'��'���N��PJ|�S`����`�!��Ra ��nD!9X�'�`��b��yR@ީ1�UR ]-i�`�Xb�0Zd��N���I���V�>}�|��/؞	��0�cY5g`�h���O����>���IQ�O�F �4��// �� l׬RnjyZ�'���
M���K��p�#<}��u���r��]0p	q�C5�t`��R��5$.}��3�rP�	*��G4q�Ph���N���ep��O��#w�>��y��_�;�"�'�f���ߌb����S@�(x.{���^���Q����x�>e�%�4��T��N�~����P�OZy��'��{�O�s���ׁ���Q�O�y�nY�FZ: 帜��+�O^]!�j����n�3���qď�݅ȓÒ�z&M��d躣���"��'��՟$�'�b�'B��O��a�&
�bF�Q�![� ��̋T�i)�|�'&�����Y�0 �>w�HmK3 ޸ ��2A��(�S�3'p��C
��ܵpp�\pCfB�ɢuCV0��[7`yR�H�/�BB�ɺ%�l��$e�E*<�cT'C nlB�	0JCV�r�F�v��ġ��<)�C�	���)ƀ��(�6%�B��	��C�	�Qc��Z��N�`�s���S�~C�I-���Ԩ�,E��dK�[�ZC�	�'�z@�%�T�HQa�?ZW`C�ɧX%�"�f�̌��"Њv	"C�3P��M"���.P�t��H.:"�lZZ���S�b�D�:07-����߁�B䉒>e��@K�K$Ta�r�ވF��c�h���mL��1� C�+�0�إ�p54�:�Ly��骆��+6��#�B�'s38��'��`�0ɂ�
8(?\�S��$B�HI���1j@0�1E�9OK�=¤��T�d4�5�T���x`�G�T�`�u�C&SWde��24�$E�.<b�Դ�B_(!���BïJ5b���Ql����X��ɠօ�$C`���Ѩ�ڟ����K<�IJ� �!-�z=��-K��?�O����r��K&O�f�hEy��ͰΨO�U�$ �q`P�s�ӁW�*�|z�"\���r��.)�mT$Js��\R|�D�OJ����d�D��;7��q��ʒ��N����d�OH��ďe�<B#�)V0 ��C�Q�~=�x�2ʓXC�F�J���h`�J�.�X����?��cZTx1��O(`h���&y�ȓbS���d�A��$�u@����ȓz���ɑ�/_"��@_*�E�ȓ�f`�$�ރK���j��?
�@�ȓ����r\�OG�!�Q+¸!=����b��CC� 7"����� ,5�����+�&�+E-�#V�e��N�3�r��S�? Ȩp�Qm�RlHd�K�\��"W"O��8F�ω'�I��A�}Z-3!"O��J��t���Î\�fT�D "O�p����7m��kG��vFj,�"O� ����
����9XE��$"O,����Q�h����,L�Δ�"Of�۔l�������<oyȄK�"O�8����@�FE��ˁ\�� C"O��%M��ʥБ�':��q�"Oh �嬖�W���bgc��%�����"Oz\�� Ŕ�<��a	AF��1#"O$�J�$,/�� �	�
JZ��5"O�U�U`��b�d��♽*�,�yV"O���v�W�fXX���J�gF�|��"OB�V�ϲI)�Lcb�yCvaY�"O�����Z�<8��"L�x�l) �"O�����Cx԰Q֤� J� �Q"Of��RKǛ�L��F��y�B��s"O����]�()4 a+]W���(�"O>E���w�Pz��T0\|�K�"O�-��\��ұ��2gfމK�"O2��w�K�1��*i<\X��"O��X$��b�
A�A6��"O�1Tl&��!mӋ&t*�"O6	�¨)D��a�lݵ0�t�R"O2��˜/Tsz̒kX�2�b �w"OD��5F�z�yQ`ܻ�nՋ!"O� �Ǟ�I�iq b����93"O�|�1�T�y���R�1�"O���uh�������.��ι��"O�-��L��t��".)/حS#"O�R�ɢ4bU𰋁�|y�y��"O�T,t�z�D�\4f�a�"Or��p@P�wu���WF��4,:�c"O�=�@�S�}P����H�Z����E"O�D�P��((�^�۴ǌ�	�İ	�"O4X��Q��x���η	�n�X�"O�Dy����,Od�9��k6��r"O>5�'ʇ b���T�0\�;*O�m��' <FFK�mC�����'��T�v�̨V�xP�-��D�'�4)d�L&�V�Z���%2��+�'��\cd��q�E�U$Ap��}�'Pn%8 � �T<���BϚS�&9i�'�H���BT�YC�9����J�d���'��a�'�\X�F#T��,��'�`���o�=> es��Z�R��	�'Zy�,]  ��$�����$�tl��'�j�(��&'�V )�������'����A��4*
�(�hK���5k�'���S!�0Sԙ���'"��
�'`1[�G��l��cDΖ ��d�'�8ya��S��8:t&�}�:)��'K��sE��o!�l��ƲGCp���'�n��b�q��!s
�B�¹C�'��P�Ŭt��Ӆ�*e+f�2�'��xK�B���~�S�"nn����'͞�6 T�D�:���]v�V�K�'\֭9�)���̄�$�K�tZ<|��'⚜	b�K$�B]��K[g�DI�'#��e�J�=�-�sڒ^���'#6p �i��U�V�r�*��=ΜXb	�'�n!���S�\�RP�RM�8;+&6D�X�c�� }�0!I1@2�H� ,6D�� ����Dͺ,)D�M���bp"O�Yb���8d����Rd}�6di"O�0�C�D</$ k��� /ZH�'"O�t0��ڸ\�v��[�r����Q"OJբ�Cә~Rf���
�K'"O��
��5B��l�Q�^&��
"OX홲K[9~^����k���"O�d�ċ/�k񥉜F���Q"O^�d��
ζu	/��	&"O�u�C�ùcZA��KH�"OT�QubBh���,� �&�T"OP(�S��v��h�a+C:�6���"Op 3�O�3�b���6�)��"O�܊a㒁L�N�+��ʌў���"O,��Q>=݁Fj?]ֆt��"O� P�J�k�f��CJ�(Ʋ�	"O�9x,ˉR<<�Mk����"Ov����B"-��ݱ��U1W>���S"O"��'�8t󾨻����*!t0{b"O$x`��I�I`�����G��)T"O�ч��<�R�������E"O�iC%i7�����@��@@9f"O�&��jzX䩏W��(�'"O��p�ԣ((!��N���C"O̽12�v��#b���R��w"O���${�8�U��UyXh��"O^��S/h4��2�Ӌ#h"y�"OD=
��ڼ����`<]��XT"OFXQ��:'�I�d���dj��U"O4�١�#)�p$�U��Zxp"O��1�K[�D�����.K��rD"O��eaX����T��$K��<�7"OF�CU��G��q�eHX!�H �"O�5ɑ�	0Ts@ۆ���[��@��"Ox=��)A�m�4�V�ՋH�hP�B"O���'
_��%"��1�U{�"OD(�D掝O��ݻ��Od���"O6e�cH �N���sm�}��8��"O�`��J�9�2�
�9]D4��"O�L	�$��KI��K�4�q�5"OL)��.V�gj�$+T-V{�(��"O^M�C�O��t#��������"Oz���.@�A�N�r"��
�*�9r"O�{��O�
vd���׫)��%ȃ"O�@��:��QP??�l�!"O�� �>'�)�fP;8�ܨ��"OqcBi�$F
���B�e�����"OB(����X9:3�ӣB���"O<9dF�,^��Vl@� �(|I�"O Ћa�P�p��֤�$�R��%"O���U_@�qaDБE�vɊ�"OP����
��i��N�-) bI�F"O��[4��*���� G_��h!�"O�0��M����SF&S�0I�"O�Ա��X%\�! �ȮT���c"ODA�AY�2��B#��~�օk�"Ot���ms���R-їk�Ę�B"OhaBf+�$��m�b
��MD�r"O�u��I}a6BU�<�����
>e%!򤕥Gh5z�H��1�h	x�/B�Z%!��0!����ކ}r �t.V9:!�߰$��8�K �?<�K�cF��PyB�ٿhȢ���OY�~��`{q ��yB���2�P`�_b����D���y
� J�`�jG��%�f�@m��"O��K�v�̡	�Op�}Y�"O%��4hD� ��!+�0�"O�K�*F5Ʋ���U�#)h��"O�i��I2]�e��័^�؉�"O�qx��ǳ63 ,"��f�Ƽ�0"O��p�c�9�AOŋ[�Jh	Q"O���BE
rXT�.	>^���Pr"O��qW,C'�.���,� �ꘘ"OH�#��ٻIJPйK��}�N�80"OR�#G�9bT\�J�3��(��"O�J��jZ��r�/�=0���4"O̔�熎�S���[��/OČe�"O����	�\�9X ��.H���g"O$i�υ-�m��o�!�(�CA"OƼyM����	�#� &�>`"O�\�k[�T�`��d+� �A"O�t�`�5���"Ad��+�4C%"O��!��:c����:+��A��"O����^�0���ԕs�x(0"O
 B�KZ1����Kߐp�1Ar"O$ B�K�>lq�1�댐)�@4S"O���5" *`7�R��4s���)�"O�aZp��mQ!�2�����"O�%+#
O,>]h���Ք&RQ4"OR�jv#��o1����Y�MY�"O>0"��3UE$$���6���"O����'&~x1��k�g�1qE"Ohc�b��/Y��"˅;6���7"O(%i%�Lyb�=I���?�8p"O���$G�_�l�p�D=�l$�Q"O<��É==:�R%敁gs0�Xr"O ]�	���pq��D�%q\Z��"O�4c5 Թ �"�E ���"O4�*� a�V�`�a_74^���"OnQ�A �#Z5�I`�`G')B*|��"O�\�a���[�2���h��h3�%�'"O.Yj�n���>��AOB�*�Z�"O�@B�D95 ��Ar/�u��P�7"O�鴋�Y	�y���,[Biyu"Op����K��, �H�h4�e;�"O���B$��`���V/֝#"O�a��D�������
	*���"O�1���i��e���C<@V�hV"O�T�fT-Ct8k�@
�l2���"O�����D'*�-����4�j8�1"O,�Xdk�Cc�\b�e	���%��"O!��ݪJ�Y�u�Y����1"O�����4#��#�B�7�-�3"O���B�U���s�A�'2� ��"O�Q��C�^���B��S��	J1"OPepČ2y�5{�������"O���MY8-z�j��Պ�s"O&������h�%	$uy!b�"O�`�S/҈$�h�`�'�	@u~I�"O���M¨1F��c�戣F`��p2"O����"Y�(�&ջ3��@"O��ۇ�ݧrQ<�j�CжP��psT"O�*bHFe��s�Q�_c�=�1"O<t���'�Ν�@�)��$��"Oف5�2 �1)���8W`��d"Oh͓vkۄT�<رW�	+F�Z�"OZe��cP<S��T;��a�	t�]�|��2��F��h�T�&<O���0���3��ܱ��,�(](�"O� �!&���}
��q���"OĘz,3�
�S�	�q���""O2}��Ŗ�ޱ{9B�Z��C"O����喋:�������|%"O�e��ʟ|k���DFO#�ɚt"Oj-��A;+cL`q&��>�ʴq"O��2'��!��-cE�_'\yF"OZ�#�10�E���Y,>�#"O(�,46}(�hc�A�pzI)"O�k��0�M����h}
U�"Oּ0�B,-&��sg	,OW�ZV"O��Ā�%r8Cs�[2%���'"O��A7�[2i����?F��2"Oh���˧#g,]:�cM��E��"O.y���״^j��p#A�{
JU�B"ODa���G}���En����3D�h��(�	G(vs���v{��.Y/!��_�{�L�Nߠ��R���]!��>b�i�W-1> )3�\�8!��'BJq��������6!��s��@J�;<��K�NB�!���&@P|!s��;y9� -�{�!�$S�{��myC�U4o{&�{��1e=!��U:+�$�u���F��8����.!����\\c�fӯd<���Cَ#.!�U�E`$�E1"����L?IL!�N8[3.�p�+��s#� @�k@!��үk�L}��Tx�a�s'G�o�!�DY)Y{�9�7���x���$���!��
5.�h��B�-7��lKQ9�!��C}�X��e�2hhM ׁ֜I�!��"
����%j��CLR}�Ӏ�+�!�� ��	áH���Ub��� #�!򤓺%�
`���1�6]��^4)!��X&2$�圹V�;�c��	�'���f�м.�}�@׶IR
�
�'���A�R�2��@�g�(�f]�
�'���i���c��`��_C�q�'jN�zEn\X�9#� �wN��h�'���ȦM2!�1�KEB��(�'��	�׬�t�Mp���i5�!�'�0Y"���1x�C����VJ�
�'���d�*rdQyW��>%{����'�(�3�@]01v��lٕmyz���'Й�#.\ $N�L��)c�a��%D���H�;f���GLC�v�����"D�J�k�j��=-�0"w�.Z9jB�I=U�y���_	(��,����/+�<B�*�P�aۡ"�܁C�ߎ�B��D_aP��� \�1��3NB�ɦs�x�aq�����	R�\C�I�<'��@u�ĵa%���*`>C�ɒNH`�bA�i��2��^Z%>C䉦
6 �a��1^F�E���8?��B䉐Y�-s֬E]شգ�"�>LH�B�	`cڤ3��ΰ��	+a��3B\B䉝Ġ	���u�-ZST��VB�q���س/���h��%��B��$����T'�C�rpY�A�g'�C�Ɋ#�D��h�>;�-35Ā3vgjB�	�=�HtR����:�*͑�O&��B�I`X�����_��*W(L!)��B�I�9(�sDEu��0{���@zC�I�$ t�[櫐�y�� ����NazC�)� f��I�&`��ޟ|���"Os�éH���b'L� ����"O����4���Z�Dc����"O�a!W'�N>�����8\����"Oh8�G"E�B����WL���G"Od�t�� +��t���CZ4�r"O�I���'�"� A�3	Z�$"OpU"��%+�t�W��4L1Q"O�(���|]�I��E�h���f"O��r3��c����� �{Ő��'�H9��
ٽh�Д�F���)��'K.�)�@�*k�8@�6��/Ϫ� �'Y�EJ� i���S�P�����'Ό�Y�莚%�=6M[	�A�'����Pf ,.��0H�-6�@��'/F0i�R�|K�E¬&��b�'�*=j�ѵ��;E�ٟU�4r�'GM�b���7[PŒ�!��RH���'ښ� !KT	N��-ش-�Sd0���'(�æ���M�Բ���"��$�'��%J���2P±�^6�:�'�N��ǻPc�c 4o ����Ѻ�y�g�!?L��3#I=-�HP���ƞ�y�(\� �*���D�,(����7��.�y�k�$��a�(��m��� g$2�yGP5 D��5��"�810&*ɔ�y�AӷP84��WI�0C*tA*f��
�yb��:��FJ�:sr@|�A�
�y"���
�4��f��kU(X��!�y�P�D%R�JJ�y;�*��K��y��4&@� ��I�E�y�u���yRKF�q��P�×#p:�ur���8�y�Ţs��4�Y�q�A�vR�Y	�'�`�ф4m��8��	80.5)	�'�DD�6�I|�F�IF��7��k	�'��]�!	��+,����LW0%'��*	�'���do�i���[A��^��TH�'54)rU˃�'���g�T9Z
@��
�']�}��*,�Us�ƻX8v��'sFܑ���0<�~h� W�f�z8��'���֩ME*T)Ѕ�H5K���
�'Q���3�J"1u�u��,�wFJ���'?�8��ꟓs�~�
4g�?p���b
�'>�HT���%�$!����jJ���
�'/r�5e��U��LB�`	����'�iR�E���V
�Cf ��'i�(� �{xR�x���3H�aZ�'LJ@���n� �[F�^�&V��	�'�|8��,K���9�d�R24��'�=3�[�V`�]WoCӜ�#�'�)�tj=-�E��T�z� H�'��}�u��z���NL:�xT9�'����H�5W�ZD��cI��'�
-"�hQP�X���(�tN�[	�'��m�W�U�+@�t�O�$(,�	�'����1Ƙ;J(H<)獜+U�©�	�'���*�)���^$��!�'�
F�M#���v�X\8�1�'!j5Xt�Ɍ Y�1�3�H�f����'@,)�񯂟Y����[:�V���'i���	�2aż,
��߄;�}��'R��eE�b�p*�eG�d��'��%��X%F<+0N͹��@�'D@Q"RB�v�܌s��5�N؀��� f�S�غw�^)���!p��!p"O��fAS���w�Ӭ;V�Q��"O�|�6��"8@��E�̀?KT�p�"O�4��l�9q����ĹD"O��Kv#� lL��QkN%�|E2�"O\Qs���	yD��%��e3�ъ�"Oʘ#0Ĳ>�^�����b���"O��xq��[�5k�� y��z4"O<������wĮ��S��bibX{5"Oz�c���~?6Ղ�B�)��$� "O� �B��x�F�����I��{7"O�*U��E�6Pf�CO��"�"O�$;GG׍x,\2��[�p�1�"OR	أ'��$�r��$
���"OڨY�G]I��x�0ϩ�|��"O�D:g+
�:H0r#�+^ ��7"OL!ICH�(*��`t+]�� ��"O��B���7R޽�dH�W�\1h`"O�j�H_�)5J����ݶ(���'"O|,�E�
9n�ܨ�aoՄ^���W"OD-����.��@��"v]c!"O�gA�4)�P��n�;䲤�@"Ohq´g��-�q�fS�Hْ$"O\$�D,ۄ? ��f%͇1 �"O��
W!Q�5jE�S䗊&���q"OT�8�*MXA
Tj�$t̴(P"OLq���5_r�y�*��cWLl��'l҄�tJ�*L��S�S�;�*��'d�tb� �\*����;�ޔ��'�(�ˡ�Y�U+"���)��x�	�'��tG�ޮnw:�z�C�\Θ���'��y�Wl����Z#�1Y���'��ȳ��F��A��>��1#�'4м8�X/_�rm` G�'����'S�����Pi'������Y6`�A�'3�803 �99�($���O�P���',�eR�H1~�( DݧB�=��'�`%[��D{��y��Ld����'�$\P�#� N��<���I�rR�Ԓ�'���B�+��{��$QRN�i�*�'v� Z�"/#	�l3c@W��H�'d� �Q�ZD:S�ҹ
��͚�'�4Mrq��)x�cM�0
r�d�
�'��+RƖ�-��]���ʧj쐙�'�`i�%O��+t�l�b�.A�0�'�X��U�f�r�eК+���'����խ[
4I%�Ÿ(#��I�'����U��|B:�SU *Is��'j��!���;+���r%�9�.	�
�'y�|J&N#T�̅�L��.��Y�
�'�`@�qM9p��P�˄(ސh��'h8�S�jǠ^6d�H�BR�7��L��'.�$r��+�~�2��Wd�ui	�''�캥f�A��	AC��M#J���'DZ�+̂�ZE�"^�A�.�:�'6:8�`�,5�6�(���H歫	�'4����#@�$w�ȩ6�d�	�'ĸ�b����`�|Х�:28��'�PYu�PW�(�A�Ȏ�`��"�'�8�2q�!�y�#�#:`Mz�'.��Õ!�|D�bN
��X�'�^�K��[���Pk��3>���R
�'��@	d��Tz��`��P�
�'<����	
3R� g��������� ^M������k�e�$�"OP ��� R��4�"
˄}
�ۤ"Ot8i�$[ ��x9W�7=L�`P0G��2cc��SŰ}���$<O�|��V0�Z4��KRs��cU"O���b���dԸ�)Aş�n0PE��"O��t�UW8��S&'�8(��[�"OnmSÃY�u�D+�.s1h#"O�#��S:V1��N$�:]��"O(=�EBC"c��ԑ�L�D�Kc"O�<K� �+Hx.e��fG�*�=�C"O�#iɱq̝�S��?ʔ3B"O��2J
���Ĕz%�9�D"O>My'C�B��)�cV�/�]B"O�a�H�!h���� c�� ~����"O���e.�*.�맡�<'�����"Ov�)��	�Uk�ݹaA��:O��b�"O`0�A�	���#'(M�L $"O���+E0����AG�9�"��7"O������z�5D�&a̸�rF"O$e�c�Ъ��
t�*Y��г�"O
}�	O&C�� �� 5�f�H`"O"�`#'ްJ�<qeBV�e�����"O��ء�˦|[�h ��ą?���1�"O���o�)����B��1"O��/��R	����#P�7v��"O@����[�&����\V{�58g"OX��Ǐ(t(��WbZv9��"Oډ*�l
"�R�ꤧ�bI����"O|���$<DDZ�(94"��e"OT��ed��0˰izs�RK,���"O���!��3<�^�;ń�j9��9�"ObT��z�� 0a�Z�Ϻ���"O*-��J�� "��#^$���"O`����T�:=��q�֕v�h���"OX89#ə�x���Pa�)H����"O���b��U�h%�T�V�(:^���"Oа$�cT�����q���"O�0�m�m�vY���^�ޤl�2"O�\���\��x�j��ăTivyʓ"O𼚥��`���G��#S~u�"O^ ��)Ż:�4nP�8ZuB�"O&Yh��
�!J�=r&푊����"O
��&^�9J����.ȋ�"Ol�����9�����M�>��tٗ"O\\"�"-C!!T��:-**��"O���D�[6Rt�"G%�t�YS#"O`r�͂�UsW!9EF���"O�����=O$���o��q5x< �"O���P)�r.�·�-�h�"O��b1�RO���!�����6"O.� �߰	�����V>+�4Y��"O4��´`���FI��r�0(�"O��HFn�/TN�󈎷E{��q "O��R�ڣp��L*G˳`��#"On����@�N�{ D�>'O��A"OL�ː�41�� Jr�Y�F���1"O����N��OT�H '[.8q�Y	�"O`8�VoZXfҁ�p��"
t�L۷"OZ=�˅�(��i��f[*�(�"O�q�p��V�b��F���n*2��"O����#߽6٘�hH��$P�q "OZ9;g�G�,#�u*惽Jq<��"O��B�y�&����5Wtő�"O��s�2^5�$L�\ߜ��5"O� d0Y�HЅ"�6�s� X��+�"O���A@A���S2���N��<sC"OlTCuMԶ0�Ed�)�P��e"O����fY�B����ᢑ�d�� ��"O>P��*�#� �woVf��H�"O D#\%��Yb��͸y�xQ�t�<�Ĉ�?6��������p�<!r��fJ6BC#�?�L����PG�<	e.��Y���shW�o��=�@y�<���>�zdAAL���δp��x�<�F*	&&�Lĳ�#��Uֈ�a��O�<��E�Ma��� �%����'LA�<���]����뗱4p`�1P|�<ٖ ��![��P��8�lQ*�w�<�'�L/L��u��k�>�t�!�Po�<�cV�zq��Ө�4i��Zcg�u�<9�N�hjY3��� Z> �a@��X�<�`"��P�pe�F�#����"AX�<)b��Q�9C�����6��m�<B%��8���Q����M����c b�<q��=x�t�h�T̤QbgLy�<iDh'��ɲ�TX��YPp�Ru�<I^���2��N��5k� &vo�C�	�A����a�(|
+�Rf�C�I�3-h���I�NL�9�jK��C�I�*�~��fcC*i�N��@	2w��B�uKԁuǉ�+�9ZU��@[fB��>(�f�36".�|�C ,V�0B��&|p�Y�L�#h�˳���Z�C��>Q��� ��	�Z�
DiK,C��C�Zv�	�AeX.]nK�g�"��B��?@�����(?*�v������?W&C�I�ΰ�Kb�٦B�r�#�+>BHC�I.�l�X_�`8��B�8iC�I;+���'�1\� �Pe�B\�B䉉��pf��/]VH;��O�lu�B�	�{�j��d �q�B�1`%�	@��C�[��y10)�MH�I�[2�C�I�T��Q�A"T98���'�S)ƔC䉦���z%�T�y�zx��n���"O��R�۞D�
4:W�\�	甘*G"O�s"�����)6���pu"OE������̌�"�<
���"O�=p�%O�h�����
�n�:��D"Oȹ@3��(VvНJ� <� �ɰ"Oµ�W-��XH��h��3l�8�"O�e��V�>^��Vb]�sO�q"O���קY?g�d|�9f+��D"O��ODG� �ccֹ|�4�G"O�<�L��*&���`f�>b�`ś�"OH!�'T�1����dƧt@�%"O�b%w��ٛq�N4oe�@3�"O�qcn��T1+�	�.I�M�"O`l�T$]�\�
aȄ��E68���"OӀd� � I�JS�BB�� �"Op@P����"��T�BA��"O ��
8k���E��!��P"O:���)ȩ|��l�A�_}R%��"O��L�$I�
�GlZ�H5"O P:�e7P�� -��,� ��"O*�
�)�z�F�+v���"O(�Aw�]��DI�%��x����f"OR��AE�kU-�	_�r0��"O��A�% tԝ�@@�Bp��S��'[ў� 
��QV!�,�`�3gv\�"O�D�"�����-�!3N.��"O�B���{iL�����3�q�#"O|����(M����O�F�"O����`Y:U��J�ע���"OZ��JF��]�p�ߔ+Y���t"Oj1X��H	B7�JՋ]�z9�	��"O~PPAL��ӺÃaމ:j��B"O�	�焎O�ʘ���< d^�;�"O��!q&�eT��B����as�"OȘ�Em�*x�vm���&C���ZC"O����e`z����
����k�"O��x�hZ
��l{ӫW�F��I��"OH�3�!8�P�7"٠L0"O��%)�>P��e"Wʟ�(�tH
�"O���e�Dt��"��J�ޠ�4"O�H�To��V����E�.4�!`"OΙ*@Ǘl��bREg*�8�"Ol����w� ��O[�"��"OfJ�e��8���ĪOh�"Oh�B˝��4����%x L=�"O�9�4��*P������ �;�"O~��Ā�2�Pv�5���c#"O��
� @fߦ��U�Ĥ+|�=�%"O`u�4�B�� @��G�Pj�3Q"Or��j^F��l���+`��"V"O�,�w��;!�i!�^1x9~��"O�5�>DCGe��xʂ��T"OZh1�'�'w��� 0�xE"O����,Αdi&��A�f�*��"Oa� B�'�^�2u S5pd8��"O�a�ĩ�^t�-	�I�	e�#�"O���ʼ"H@h��P�WF8�Bw"O&��-�03����GE�@=,А"O�jUŝ0cBj�맣=��+6"O�}���M�KN���b��b�T##"O������,>���`37}���"Op�kQ-�DU Ya$OW�|N�()A"Oy�%�	2���s�͟�IBK�"O�s��gZH %M�4c0�"OJ0Vb��2j�kP�c(�K"OxźV��16�V��C�Ι�rl��"O0q���	y� -Sd#��H�#'"O�8��^�QȾLYbE(y#��җ"O�0Ƞꏀt��`��:2�&eJ�"Od0�B��s �Dڵg�|<e2�"OмH�E��)�xeZi�4J��$"O���b�:�|�0ը��G]�Ԁ�"OƩS��+��8X��ZVl:�"O�a����m.^�[@�:p1����"O<�``\$z�0u$){�͛A"O�]�,�1V�T]�c6�i±"O|�H��0S�p�R�B�p���r"O��뵊F�vD@Q�G�(sdT� c"O\��� I��`(S�)yx5��"Op�𤧔0}�x���ti��"O�#2C�.,�9�懚�
� 5"O��rc,��k�x��UB^��|�f"O>T�f+�.n|�#A,���hp"O`U���J���J��/q�V�H�"O @�:3'f!���يi݌��"O ����d(���5���T"O��9�B�$��-�d�̐0`����"O����kY�E�)dW�4K�,�b"O� 3�D]9g�@���+X[�2�"O(�"���W�HU �a��Wl��s"O �ѷ�Z?,�q�FD�6X����"O�X�%KO eefL�WEF�EX8M��"O�Hk�͝�"|��fL^9D<�"OB��gP�s��L�ш00+!"O�̓ ��_��x��J:���$"O6�B1�́,��P���"Cbxb"Oa���C4̰�ņ�w%D���"Oh���=؈�� ��bִHc"O���dT1Wp��bա��Z�"O���I�n��%�eeڕ[R�p��"O����oȚ1�p� n��J��"O�!�՚?�V���Ԫӊ�a�"O(�
��)0��#儓C��	"O�)cc@[�k*��壒�%��I[v"O�LSG6r�dYQ�m��n���`"O���c��0i�Z��M
|�Tc�"Of#��%9�1 ��S),��B"O�\B���y80���I,. ����"O�A���T�/N N:J��"O�P���¢h���09b���"O��w���P�|�㐕	dU3"ON5�Sg�\>�p��b�*IV9`"O���KˬWK@�G'ܫ7G��"O�qK�dM��JA�%]�@�)�"O������1�H� ��Q_�1��"O�{u%X2 -����4CO���"Oz�����oA��Q���'u&d�p"O4�Y�h�A�n��th�� u���s"O,����;����ħ_�79���"OrTj�M:+{�8��ƒf(�yb�5[������Kw椩U���y���+��E��p�"TZtj	�y�G�ar$0�ϗ*k���{ҩY3�yb"�z�Lmt��K<P9b���yr	q�"q0"/@=Zm��yk�;vLV�!�Cр5�xj��1�y� Y`f���.�8S��-ipϒ1�y"�q����,�L�H�QQ����y�Þ�q��Ĉu�Ju�@��A	)�y�\+>T�)V��`��� t"Y��yB��`��BE)�fQL���(��yb!U��Y*�Ϭc����gd��y⨓	c>H�����4E��(�<�y"O5ay�8���M�,z#����yᛱ�,�e�N�FyHj��y��]�d����	L�%�u�I��y���`Ր�vÛ�?5�u���yZbX���ԈF3�!8��c�`��Rg�B��Ef�8��@�6��чȓK��y�3�
�48Y��ĿtW�M�ȓ �	#��Y?JF�B�h�vH�ȓ;T���B)��v\R�Ї��J��=�ȓ.]�x��OF$`�Ԃ���ȓ�T�:�$W/5v���S��8�ȓ[1P4�r�]�Ľ�f"+3D��/�� a�]�ԅ&g����<D�h��C�gVt��#�n~(���!%D�T����0Q���#��ٴ<��#D���'Լ �d�E�^�[�����=D��$(��{���b蝵C�z<��N>D�TpC��w��@�����."�r�")D���aa�*L�xâ���f��*T�2D�� v�	/Q�~����h��l����"O��9%#®S���������
�"O����B�.5�؁i�(��|��Y��"O�a��\�>����)�.0T"O�� �	چΜwhÏ�r�rs"Oh��s�[�]
�:�L����Be"O6�y@�ʲR��<8���e�t�"OܙK6� �����e�	]�Dx�"OL�1V�8u�QjD
�=��h"O|\J�F�U��!��$#�f|�#"Oȥ����N��8� W�^�6H�W"O���Mݔ	A\0�%@#��@x2"O<�Q޶��f�������"O�x��E�'��`��Z�!*�"O�\Z$&�n�x��r�P2�
�#g"O�Q��_�+z�%��n 2��xf"O��4�Ӝ2�I�`�:��P�"O��C�O؃`�8x��C�U��]�2"OL�� �� �x@stED��|Z"O�г$��7^��� �'Ŗ�R"O��˙$,&�A��ݓ]���
6"O�zƊ	�P.�u��!] 4��ɨ�"On�*�$��� � [�D�4��"Oj�_,Q>��ǮB�R{��AW"O`B�҄a���$�!OPt�$"O��t+W�,�N��eg��'�6@�"O�i;�B��z�a�����Is�"O4���oD?'��ċ?C�N��C"O�%��f@�/��$hb#�>}��A�T"Of��ٜ%�py �6Nf�!
�"O�"��e������5�7"O>d���%i��cSkT�z�C�"O�Q�U��#Ja���Ӈ������"Or�iA�� q��x��ԂY�2�pG"O�]Z��!Z���f�Z��,i�"OU{�]��Rȩv��-@��xI�"O���#�^n�!Z�\��i#T"O�$���J�9*D��D�M�"3u"OJ�q"nB5g>P�b�l�-`����W"O��I(��Q�����j�"\s��Bb"O����+9{�I�wDA .MfH�"O�)�`$H�nd���+7�8��"O쬡�L�>����6�F! r���"O�8�K'n��	Ra[�y]T9pT"O�!9�� (m��d�R�m>�`3d"O5sqKT�,R�d��޶m��Q1�"O�|Z5#�3%5�q��B�X��q�%"OP̀ao�U���*Ҫ+��!!%"O�I���+3��)H�	3dM2�"O���գY0!XU %��V�����"O�@�j̮@��%�ĐX�� zg"O\IȵK�5�҈���A1yQ�|�p"Ot��ՋġrN�ѻ%�-�����"O�����;���C�I4��A`7"O�9�b_L���B���w��	Z"O����l�$EPH���q�4X��	]x���i��
�h�1�d=�6�  �.D�T�`/��lb�
R�i�@�k!D��xe@/Dr�Qb�d��NF����:D�Zp��P[h�;u�L�c�^����8D��a��&$�F�p �L�$V�!eo+D��j��/iP�IF̞Vzry���(D�lgś�5T�k�	�S�`I�g+%D�K@c�8|p��G�~b]��!D�� ��ĩԒ_��	BW[0��q��"O����Ի-�t9��ž1k�t9�"O����lޮ5�t� !=^v�)d"O(I2Ɯ L�f5
��U�ixP�9�"O��'��/X�\�T�4u8�G"O�e��̆N;�T�@Hkn)a"O��T/&EP�'lޢB_Pt{�"Of�b�g^�s'���kH5\(ҙR�"O����'9;L��q���B�X�"O�����Y�a�f	A2JD�୻�"Op��bÕ?&���1,B>!kJ��Q"O^8g�هd�~�:��AS��v"O����'[�	�$��r�H�,M佐r"Or%���?K�T�� W84L�8�"O��:�4	��!r�UyDx$�w"O�����t����@n�<@/�yI"Ox	'I�R'����- z�""O����a�f`����k�����"O���
+e��4�deâC>��"Od����O1	���j�� �MN�ȑ"OH�+B-�8-x5*U�и+̀r"O���CǶW�Q�U&��/4H�"O�-��̏�W�DI����6ܸI��"Ot��M�/���Q"}�ޕs7"OxH{$(J�'W u���t�څ�w"OMz���2wz5��L2��2�"O�]q�ӒO,�-���7b|Z��C"O��+%-T�lN�BE�yd1q"O^��G�9[������4Fl�چ"OJ����c7��A�n��(��D"Od�W�D��1�G�ޠ��j�"O�u;�m^4(��AT���\k�"O��ؓ�I)_k����M�a ��f"Oܠc�@U�?��cr,Mi����"O�h���Q3H3uk�9��K�"O��1�$�~�@�sf�K lN\��"OVaq5��R��0��|,��t"O�����A��q� ��<fX�h�"O�!0��cJ�8��;7HX@��"Orx�!	�,^�x�ѰN  �j"O@QkgM��c���D�6i,Y�"O���Ɵ�	�椸cW;N�D	 "Ot����M�`}ˣ���W���{�"ON�	�.P�2!2��J�����"O��%�ۼ8�t���J�&�@e"Oċ&�u��p	/�>%� "O��`��^.��
W.\�-5� [r"OtY�-ҏM5{�MG2J��9�"OvhR�Űy��0�w|-��"O�E{Q&q�T��w��59��"O��b�l�Pb@�q(�.%�uXq"O��ꠀX�1�2	�Dg�u�$}I�"OT�
���4d�"�A&4�xDQb"ObM�fJ��0�PČ(j��Dٷ"O$bG	I�S~���`ƻ:���"Op��XI� x2�J�s�� !"O�Y(�F�&+�,r6/ �\���z�"O6��h���@�qNB�P "O���R+�!�ƅ��c�8TD��0�"O~�fn��a0p�a�Í|3��`�"O����۹ r���nҔ~#ZxS5"O���B�<vKP�R��"2V�b�"O�pq��M(t��+\n�L: "O�9{cC�1���$
b_�@qB"O� ��� �8�6���!�T7��v"O��4 ߚG+.�2Aߖ[F��"O�=�S��U����v@@4���"O(��"H�y.r<���"]c
9c�"OD��B.��Q�n�h��!]Im��"O�#v���v�ؐa��F1�L�$"O*0�ש��U6<y�CҫE%�0�"Ov`QD�݈@�C$�����"O���W"��X��e�ƉE���pe"O�E��' G�ʤ��aK�� �e"O8@{�eʥ�����4N\�ZL�O��y�
��M��O?�	}�>�RE#ݲ�B���KJ+;b��7��g4�a22h�;�Nl�p�I���>���� @f�d�@�ٰ.
�d5�k$�i���"���8	kE�`jJM��!�j�*� ��gP+����� &J/�(ً�GD7f�ڗŁϦI��e�O����_y�'�����y�0 ��_N�P�d1�x�D�O��O.#?� ęS_��J�B-u>�dTL�k�'�Z7��O��?�oڽ#[Vl����.���ό�B�[��?DяB4 �H���?����?�t��p�$n�h�;��1()PP���SDp�� `�༒�B��,���f�G�h����F�X�p��v� ��f��/Py"���.8�9 -�lH��J�f%M��P��2�) ��	�R��|@����&�9Ї�s_� �A�b�a��|�f��c�,O���>�bhɛ#!r�ԗ\�^H!"��\�<�lP*�dD����@�x�RoC`3@7-�O8�O��	�O4˓J�Z�(�+��!PK3Q`�+aKN� 3ϓ�?�k& �B�"ф"�Fy�M�o���%`�����)��:3��@�e�"��"r���Vd�e� sD�5�Q(Pq�˓�h �� �j��!��������F�ē*��I�=�4d�J�@*6���7)8	���3D���'��Işp�?�Om�� o�p�2�)+}����']aR���Zep1� �*�\�������I��M�i�剄$�x ��4�?����ID8Cbr��a�UX�,�V΍	?Dī�)������ʟ�H�dI���<�C.�lXn�UN×+Q�M�]���A�=�WƼ	7�ɨ����q)ލcj������#^��X��,���[�)P/�����EW��+�
$L��c��)�O���PA�S�"P��[��hW嘦f7x,17�G �?I���T�xbC���`l���%s��h�����p>�ӳi��7-k�ޘ��ij��̳"�L�8�Ḱ�O�فPb�צ%�'�ӸB�p��ğm�2��` 	{�B�.�!(#$,{�ć�6� L�#A�:f�ڽ�AD¯#uz��D��O.k�q�����N����'<Gp��$�3Zp�C��R(�8(��s0$ cC�,���kl�PF�B�DT'F�����G	�����?9�����N맭�s������(W��:Sa��6�m{��Ot�D4�O���/(x.���	hH@#�ɋ�M�i��'�����0��N� sȥȵ![=_����ƍϟ��	l�СuJY̟P���� �	�u�'���Hg�H�p	/W \,���GJ�R�p�f��8d� H*s������L���d��x�d����(��� 2O�v���GP��C�Z��G_?�I�J��hx�p;�OL�(�B�>H��d�P��C��7_�X:U��O�nڜ�HO��	�m����2V<T2C�(-HQGy� 0�S�$�/�zؓA �?������'c�mZ��M�J>�'�N>iڴt1� @�?   d   Ĵ���	��Z��wI�+ʜ�cd�<��k٥���qe�H�4��6X8$<)�ih�6���#�t�`�ÞP�nѱ�%��>iD�oZ=�M�!�i����B5����OG�wo�[)Ն �eaB
��M���߆�O��#ߴ7��z�fU�_��d�!�^>*b�]�'���2#O�)q/O��2�����h�+O�=�v�.)��(u�u��n;YzRp�/	�){�f�M���M�j1A�4-��7����T*��[Z,��/s@�I��hΏD2���E���F�;\ �u�i��˓��I�1)�~?!p	U43���a��;?�̘��NL?�$Q����<yP�ܑ]Xb���W*B�4�>9:0 �T+:���`b��HS�;��hq��� v��	7y��aX �O����[���$X$�d5���W	�R�"jE�Ml"<��=�	:^a 1sAہ�d<�b�S��6���O�x����0��񥁂5`b��WB�cn2�Pw���O���O �Ym1�B@���VK���	�T�h��I'��O��]����@8x����+E2\}ExRGFT�'P�4�	4e�b)�P���q�&lk�$K�<�c��ht�	;r�'��|��g �4X�Ǫ^ ��(�'t��Fx��h�	��~� ��\��JX�t�z��@.��?!b���⃋=�,6�(}B��9k�$�����t�v��<�R�:�*V��0t�'@��Q�����R��xY�lk�IRp0D�ǰ3��ȵl��K=�ɠ�o\CB�b�D PG<�Q�\	�L���4�r�AU�f�TZ5�:D����)   �v��요�C) (jC�I-5�:��$͐%.~�Q�k �w>C�I[�|���u�\���;Z��B�	�aRDl�QF](C�*5�PJ�K�B�	*!wN �6�R[X�0թظ+�B�I�F��i�EQ
~$R�0�ɷ�lB�I�d��H���'H@(G�GJʖC��qt5ض��w�`H6 �7`�dC�	3��b�Ď%��Q�q`I�4(pb��QrJ�r��R�茰5�xCgL�/���ᦏ*z
<�����b��V�J�Y��t�`%�a�0hȖ�Rg�D�/A
0"���5���V�����E�e�:���#�U����S�V�r�Tl@W�|x�):3�ޯ7BE���#K���4'�>� -�p&]�v�[�&Z4J
!poq�ZLխn��P�J"h�����Uҟ\��/)dd���h�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  3  v  _  �)  �4  �?  K  ^V  �a  �j  q  �x  !  d�  ��  ��  =�  ��  �  A�  ��  �  h�  ��  A�  ��  ��  8�  ��  0�  ��  �  �  � � � - �% , M2 [6  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6#\���<4�d5h��'�B�'���'	�'/�'�B�'���$��^] ��/U�Z�3��'m�'�r�'���'K��'r�'cظYA��4Z8�xg&�=�nܳ1�'�r�']�'���'l�'���'��41Cl֝wMƩ���0���4�'��'[��'D��'[b�'���'զ@�R��}�[�&���Ģ��'Z2�'�'���'x��'��'T��s�D
����c̚�	P�'V��'��'2�'��'���'X���EAO91�(��@�{�x=���'+R�'6"�'���'���'�R�'%l$�H^�C

��\�o��ص�'���'@��'���'��'��'��12����4��x�Rk��'n��'�2�'>��'r�'�2�'`P��6�.&M��;�	�:�d2R�'��'���'���'[��'���'��u��Ǎ
���z_��BT垲�?���?Q���?q��?����?���?��O�1^�����*J+Q4	zT#�?���?���?y��?a��?)��?i%��=�61Tg�y����ڟ�?)���?!��?Q��?��Px�V�',rl��~
I�"�m���rR"�U����?a/O1��	-�M#�  �Ќ�EKB�[�L� Ӊ^���'�R��<��k����@9;LU���x� P���?�p$#�Ms�O��Ӂ�zO?y�K�(Pd́�蘽,���;��<������'o�>�RR.�w���Sɕ���5=�MQ��Z���O�wL]�"G��9&F�b�Ya.��*��'223O��ŞXZ:ٴ�yڬu͎P)TcR?�eI�j��U�di�P��T���=�'�?)j�5c�r���&��nM�U��+U�<9.O��O�o�+E@�b���o���mɺz��(�0.^������O����p�'���B�]l�l,����9AXѪ�O����/ m���5�گ�?�5��Ot\S�j2f�ZŊJѯ|2�"c�<a-O���s���� �?��Mb�
I�J<
Y�y�%h�ָ������W��|��L$�	kgF�	cr��r0�S�<����?��.b<h�ܴ���{>���2�ZIs@׏��E"�� %��hԁ5�Ĩ<�'�?!��?����?q�f�8��J����g4��bS!�����P��}�.�۟���ş�*'g��0�	1�\# ��+0,���$�O@��!��)���Z�BE�>i=T�[#iI$ھ���#D*QB���>|�U9Q�'��x$�@�'��`(�O�J�!E�F�<����'���'�B���_�@B�4�>q���` ���Ѣ�D��rSL�+�� ���?a�BS����ş�	#_)����P%<�$��4oE��:h��/����'�J���WK�N~B��O�����F-^_�r7�ۂX�6���?Y���?1��?9����O� !�@�1g�P��4|�3��'��'8�6-[U'���O��&�$ȫVd�|As�D16`�c��:4���O����O�L1c��i �ɐW�Ȩ�afW�lrN�RSKE�2K�T{0c��i�_y�O�b�'i�c�.�p�`��06�lXR���Mo��'��&�M�q�H���O�˧&�\�8@�Q�ev�	:���6gm~�'��۟��?�O)�k�dߧS�^�K�,�*�����Q�f�z5�E���i>�i��'�>,'��tX�Ϭ|eF��������ڟx��ٟb>1�'��6mSv��A� Y/3u�tµ *���ՠ�O���O6��'#2HE�*9@��Э��-)���4K���'�,D[��i��	PM0Hc �I �.�,�w�ޭb��r�1-�Ġ<����?i���?����?�.�
��D`����8l��J�f�M�Qo�6{g�U������c�S��`�i�*!F^l��T��<0��d����d��U�)�7�� o�<��HAD��Sk^�$S��0p���<I$ς�M����S�gy��'�"�G�V6����o��I׌����� l��'���'�	��MKs����?Y��?q5��#[�6��0��+��8�g���'��͟d�IU�`���3��7 V�IsJf5��o ���ç�"�M�����OZ?��ӂl�6""0J@�T�Y����3)ب�?���?1���?���i�O�y�r�T���0���OnN\
���O�-mZ�����	ɟ$�	z�Ӽs�E�
1�9G��*E&��<!���?a��T�J���4����D��e�� 9(FP�L,�%���J1�D����:�����O����OH���Or�dςm��������u��,	��}�dʓ,��Vͣp�'Y���
9�~����_0s��U@���/n��?�����S�'`��E��)4�Ӱ��`^������M�d[� �� |�"���Iqy��T2j�&�kO:C}��A'0�	ß �Iɟ�yy� wӪ�)��O��%	Ōr���q$j��)�f����O���>�	Iy��'S�'a�P{eĨ� J��f��2 mH�iɊ7m*?�cʊ�:����?���� x�D+*��]�)��7x��>O����OL��O�D�O��?��B�țs'��0�+�t���!ڟ��Iʟh�޴M��[+O��$"���C�x���꓏#YfT�3��O����O�)�p�7�-?90��,tЙ���ъ@3��'@�L!8�IJ��~��|bU���̟���ڟ̀m��)�hʴ�G W�t��-ޟh�IuyBn�O�!��'���'�哅/�P�s�߷E�v�xV�	=j�����O��*��?#C�8�����Õv'X�؄��0`t��Pm�$FP��|z��O���J>qr`A�uJ^ѲF�U���Ru0�?���?����?�|"(O�l��\�N9"٧9˘��GJ���ΔПl��֟<�?I(Ol���Y �0ᤔ�d�U&� �D�Ol��SJeӦ�A#�8�u@�?E�'1���#���[�4y	F�H�(��q�'��I��	؟P����D��h����#PA*4��Fԯ��i�фM 7��� �����O��$-���Oz�4��y��ζ]ot}B�.�-RH�����O��7��aNz6�{�z���3$Z�5`�@�V����{�0C`^7�� �[�IFy��'��eD��AP�.����b�P���O����O�˓#^�v#�G�b�'M2d6��#��4����V�jG�O�˓�?����;R��0�E3L��p���6S\\�'���ql��v����TM�矸q�'h���K�ꁳ�A(�H��'j"�'~b�'/�>=�ɝ! ̹9T��=QR��懏1~������MS�*
�?9��?	��wp�u��+*%i\��ЌT03��$b�'{�Z�D�uE�ڦ��'�H�33J�?a��QCT�Ͱs��M�zE�צ��&f�'���ٟ���۟��I͟\��M�������[
jE���Κ(ޒL�'�7-Wvw����OR�d2�9O̍�*O AU �j��Fk�&��U��<���?�L>�|rR�J����Y�	;,�T9²��+
��pR~�e�$]"��8$*�'X�$C��)R̎�_Z��
G~�h���ڟ���П��i>��'X6�·l5.�$�?d�&�H"��_;<L��,=��O�|�'���'[����6f"�����L�&��5-ο$�@���i����8��a1�ݟ蓟���ȶ,Dhe�������t�򠕰L[��O^�d�O,�$�O�$(��-aK�)h��9%� �
�)A�M����������MˣET�|J���?�O>yË�;Nb
p0�AR�:y�2nǋ���?���|*���M[�O��厖?,*�*��&¬��V>.��?�
)�d�<�'�?y���?�2k��I`
�pJR,(S��##�/�?9����æA�6ETay��'x��^�^����B���L �,�P�h����O(��.��?qY�τ�Q�6);�$C���` ��5�L���hP�E��|bg-�O��J>	�@�f���b@!&,�\�`����)�I؟��	ҟb>ݕ'.h6�'�$�0T��;yN�+��C
��M����O����O:⟰�'(҅,@5�hk��� }�{eL��n��8FVtmZf~B�����W���y�n� -C�LY�%*��aaZ�pyr�'��'���'�B\>��u�pj��g�i�2�P��#p�xAA�O����O�����$�O��L�K�f�Z�'�i߰�'oK͌�d�O��O1�x���No���>�J,��[)8��A�� '�t�I�Y>�Ɋ��'�	&�Ė���'-�eY`�	Y����
16o���'Q2�'U�xڴ)��u����?��5ĐPc�-M+ Q)1�8�*�x�"R�(��Ο�$������<����U6$�H�C� ?���(wT�p���L�'.v\��͌�?i��
?t݊��)A��P�'��?Q��?���?���i�O�� �hM�`ւ���(0�p0�#��OL�mZ�6��IΟ��	I�Ӽ��*S6BR�I����E. �*���<!���?I��X�>h�޴����Պ2k�&e�EZ;� z���oU�1�wσ������O��d�O���O�����]�V�{���P���P�Φg$�˓XB��
u��'�����'.u�%�	��D��]�p��U�p�	՟T%�b>!���B\�$Q��A�2�&}i�a�5P9� de)?��b� m�z��������4F:,L�F��NH�p��*P����O>�D�O��4��ʓ���(7ҩI��ش��"BE�x2e���2�'��O�˓�?1���?Q�YKL0���g��ot\��d

U���ݴ��D�):(�AK�'��O��+��\��T�)w|��4&�6�y��'���'Er�'����I�sZY`sK�
%M>= ��)0�����O��D[̦:F�Sy�'��'�����\�ؤ(�"�'N&v�Z�|��'F�O�hy!5�is�	�30 2d#U�2>�Pf�Zg,���IˣC2��a�Iby�O5R�'��`@�� �2�WG��RĠ�B��'��ɐ�M�(��?����?I(�`U�i��݈�86̢ ��(���\�'���?i�����L�7)L.���c�&zoL�@��}��������C�L�B�dB�*�J�
+{��"s��q&��'��'1��tU�iٴd�
��ł�1��Ă!�-x���@�����O���'!b�Ҷ%y�P�U�˘?�d�,
�;v�'�4�	��it�	�4`n)�r�OM�g�? �գC	֔B���Ч%W7���HU1Od��?����?���?A���	Ť)��<��ҤE&��̀�pδn�+�P���,��H���?�;`��d�d,?,r<�	�C�C�¸���?�J>�|@.�9�MÜ'�ap�� �&�2��P.ZTp� �'�~a�!(B�̢Ց|X�p�	̟$��f��w�����b��P+6���������ٟ|�IMy�$z�5�n�Od�d�O6�1E�#ɸ��C+�J���h�B"��ay"�'\��|��-Xk���c�;Q_(�Ң�����Z�tɩ��|����^����y�"�d3.k�1�B���3�fIH!J�^��Of���O���$ڧ�?	@E���Ha��4���1(�?��i�vm���'>"�'��O�A'pd���H�������\���O
��O����e�"�l�&p�qM�?�Q���P�8M�!8^�%�&�]��xy�O��'��'B��	��t���6[2�����9!��?�M[��/�?���?���I���d�Z��0����+b�	���	P�)�S����f��p���F�U�=8dI�vkJ�h���,{��m�O{I>�.O58�/1?�>!���>P��h��#�O��$�O��d�O�)�<�T�iö�۱�'����q�ˊ$�6ubէ r�:��0�'���d�<����?Y�*���#�q�tɓ�g2A���A�\m]~�"H�{[��S�'���2L�%�D�1��޴_�b-�Ä�<Y���?!���?!��?���b��K��р7","�|z�ki/��'(��m�Zx 3=�P��OڒO&b(���֍�%ؔ	�BDh'�$�O��F�
�+�4��D�!-�,X���9��E!��x2mqb"��?��9���<a��?a���?Y`�kE���`��@j�SL�=�?�������*�+�0�	㟀�O��%����.�Q����$d�d��O�ʓ�?a���S���	=@%�I�m��,�*�1�k�����)��ƾ<ͧ)h��o�)ȴ�)Ϝ5`��P�n�/L`���4�	ş��)�By�e�v�QR�O�OZ�9�����jc6�E==d��d�O���6��Cy��'�"�� �v_��0'�/����R� �n�ЦY�'�uaW���?�Q\���#���g��D����3���qu���'�r�'�"�'p�'��2J C�K�q��� НK���4\�TyQ���?����O$�w� �T�I�B��(�,_����'%��|��T�?n�<O�����9������)oC� ��$��.����'��'��i>�I0��q�F��"vF*QpPJ*&��1��ٟ��˟��')�7�	24�V�$�O ��?9�ġ𭔠A,i��L�"Sn�ؔ'R�'��'cء�L�&� ��m�D�I�O�M��?�&7��J�S�~,�D�O�i��ߏ*��A����^� � B��O���O����Oģ}��%:�q��N�u8j�铥�/U�Pl8��F'�vDU�7y��'�4�^x��V'[����p&R6#�����0O����O&�d�!3}86�#?�;��ɋ��(���Ò� �`D���9{L��7�'��<����?����?Y��?��N��2���~�𢔭Q���A�����w9o��@�IQ�':_����%P��i�	Y��;)O����OX�O1�xt�Vo�v�+D��oJL�;�9=�>6��qyr�߁��������$��9-��;���Y��ؓda	��d�O��D�O�4��ʓț���rb��Z!|��7C6�q��@�8t��'��OZ��?���?�DC��C�9K挛�l�Mr��L71n̒�4����"(M2�p�'�O��S�v�v-����2�z��gK��yR�'c��'@��'���ɓ?C]tJ�ņCk��S�l�<�:�$�OH�$��-锧q>��ޟh$�x	��|�b�3����@i�t�U��h�i>�2�����'_����n4q@�`�g��mΚ 
�B5e�DQ�	6~�'��i>-�Iݟ������DЧm�Q�8��eK���	՟ܔ'c�7폷pO����O��Ĥ|z��S�Jt�M+��^�G�myR~bQ�����t&��+��ز`���2���+ȑOD�t�2��| �Pjb~�Ol��ID��'3.
&EV&h�BE����� <�4�'q��'nb���OO�	��M���ĸ�"���ρvB��  P�tԈS���?1���'���Dp��ߡr��BW�ۋR�$ z��D�<�I�z��]lI~��9�ҙ�}�c��"=C�`��l8T���<�+O��d�O����O��$�OX˧Xz�i:C*W;%���Ť����G�i���c��'^��'��O_��y�-P�0�E#�#�>B"�Qs��0���'=ɧ�O���a�i2�dٗR�D�4l�5Co�Z3��[��Mf�D\��0c��ON��|*�|3&��H���@���Q�vm(EB���?���?�-O��nڲAk�`�	�ɀϺ� ����P�<
B��=u<,<�?!-Op���O�OZ����Q;KάA��@#d޽+Ĝ��Y�
C<!vTo����' yJ�	˟0�4,�L&H������B��J�����I��l���tF���'B�xC���{N~E_�4s� �\I!t�\�*�O�$�O*��]�.�bɺ4K )��z'k'_N������� ���ݦ�'��q4)W� �M���,U�l�0U�A���8���<�'�?����?Q���?y$��}���@�Xr�!�JC���$�ߦE��.̟������%?�	�*�c�d\z~��k �W�E�
��'��'�ɧ�O�|�����I6Js(��)Z]���;&�VJ�<���J/D���D��by�G�2g�� Cf�++��!���Y8a���'X�'�OQ�ɣ�Mc� �0�?I �i&��qiL�pU
�@&	��?i���'��I�P�����ؒ�:'�a3�h�7J������R]E0UoZp~k
�K0�t��@ܧ���Al�=PHU˒D�=*�`��<	��?����?)��?9���C�֘,T��=\�jE�ԐDR�'i�oӸ ۀ8�����O&�O�X���ܑ1�Jd 	W?^�p�w�+��O��4�hFoc�L�-Ψ�s�4_���v
���q�B��7���D��䓶�4�\�d�O��$W�TA�!	ԄT9K�x�sF�� Y����O�˓nț�
* �b�'0�Y>�y�#E�=ڄG�)@��M	�#?�)O��D�O�O�ө<y�		��ڳIL|T(��0`̘�ӄX�.�"��d!?�'\��	��tRڴ�àV�%䨡���ZH�����?����?��S�'���ۦ�A�d��#2Zr�h\*D�]�B�i�	���Ig�����O�{���,9^�iI�
�8/z�:�M�O��I�B� 6-#?&K��n[��i/����$nYȷ�>D�R����C(�y"R� ��� ��Ɵ0�I���O��mJ3)J�R���4-�x��R�y�vu+Gj�O��D�OB�?I�iމ�3��q>��P�8��Qc ˇ؟ �?�|�%�J��MC�'{�YP�=�zU�3�S�e5����'�<��3��� ZƗ|r]���	ҟl
1��)6`i�5��d�beX��B�T�	͟��My�Mj��t[�e�<�����Y$���C�&J�l7 �"c��+��'7�矠�Iw�_��\�W@�H��q�lV`�#�����Τ4���|զ�O���Y/�Z��%z2\	�OZ*f�>�y���?����?���h�`�d�, Rv�cCM�P��I�aI�ls�����	��n����	���?�;ˈe⣈�="+��1jԵ��?����?I�����M{�O��;h���Y�8k�yڔf�\o���#~W�t�I>�*Or�$�O����Ol�d�O��Z�cA�}���C���*�k��<9�i���s�'�r�'��O�E�u
�� !E�&oR�*�������Ii�)���6ŋ�	T�8W��GP/,��Q�h�,�!^�,�+�O2Y�J>�*O��s ��0�Z�Aӧ\�a��H�O����O@���O�	�<yS�iŴ�R��'��`�I�04aSɑ%g2�� �'���d�<����?��6�J�S�D֎/Xa)%�Кvδ�A����Mk�O�9s�f̵����wTa����)zܴ�S��=\Ϭʟ'���'S��'@��'��Hx�
C�Q�j�fBߺ0����Ϥ<���^՛F#�(����'�R�|B+Y;T��' ���mY��z� �|2�'��O���D�i/���d�챣&�!
�$r#�A�nE�|2�GU�;o�b��[y�O�2�'s�i��b?ع"W���,"8����{�2�'��I�Ms"���?����?�*�њ`h� Z�\��C�]
Xp8�cѝ���'<r�'�ɧ�)"E��a���x���Φ!�޴hѺl�uA]y�OݦY�I=�'-B��應�z4���b��}Bd�#�')��'5R�Oe剘�M��nߪij&��u-S�N�=#C���sK��������?�,O��d@=J:M���=R�.��*R�}2F���OuQS�{�2�Ӻ{ō[����*�<i3��))@���*��$��A�F��<�*O����Ol���OZ���Ofʧ��2�?n9��A��'t8��R�i�����'%B�'�O'���y�f��9�ĝ�e��t�:�s���l��'ɧ�O�$cR�i��D��!���x&��:1&K��B���d��B���?Y�䓬�4�F�$�5��9:�΋�0�l�@�"��"����O ���O$˓g����Dh}b�'�B��N�N��R���4t���L��R��O<˓�?)����Aڬ�`� U�<���P��Q@�'{6]��8O������������5�'b6�z�hL��-�NT=Ae*0(��'���'���']�>���<F豩ħ��6�0y�b����t����M�U����OF���&��1�b�W��%A��>���	ß��I��<bEg���'�Dh�Eo�~R��ȱ/<�TY6��sQ(��1B�����4�����O����O:��Y-7h��т�ivT@�U�r��˓sl�vʐ�:�"�'�����'	v�K��/#�,��3�lۡU���˟�&�b>�RmP�K,�s�[.C�`y���<��t�d"�my�啐�`�	���'��		&4}zUK�)\eĄ��_�9�(`�����Iן��i>��'�7-�?e@��B�t����у9i���ٕx���O�,�'H�P�LA����,���0�I�B�*x�sV�Ϧ��'a�8��E��?Ţ���$�w�8����g�<�F���H�'�b�'��'�"�'��JĦD�8��tq�d� b� �J�l�OF���O�n�'��Sȟ��	c��\V��P�bdCDP��-%���Iԟ���m�A~"���� �� ��)u��A!�fz����_ �~��|�_��蟼����P�f��v���ڳ�^$!� T�g��ȟ$�Ijy��x�d%��o�OT���O>�'U��ყ��v:����.W�,E�%�'��I��(�	}�)��-i�TY�7C
4WhH�@�.Pz��B�º^3�����+IşH1��|�+�$Q[D��t�Кl�\�����+�2�'\�'����Z��{ߴB� �BE+�!!�h��T�-����E(�?���?��"]�t��mq�\CRn��0��,��K�r������ؖE���=�'ѐ��c&��?���1 �O����'E$M`� ��9O&��?���?Q���?����IL0H��H�"k�F- C���Z�o�`�"����$��Y��X�i�e��"A	2��d(Ι�>8ydJ���Id�)��.H)n|l��<��IY�m��0a���J��J��<�fN
�r���U����4��D-�½rŌ�SC����O�?����O����OXʓH����%!���'v��t�$��O-h�(�ē#5E�O8��?وB��*�i�c.�q��(C%(ش���\$#�Ay�
Z0k+����IQ��i+*�䃯����K^!Rfr��j� X���O��$�O���*�'�?���ՔZ��L2�"Ъ[�ND
k��?���i�dSU�'@��'��O�.�y�q����l�Q�s��D�Oz�d�O�P6GoӞ�D�Tra��\�yӀN�% �=9���7���q&!�䓶�4���D�O��d�O������ԥH�L׀1�d�ٹN�\�/���ӵC���'
�����'�����F��rL،�&K�H���c ^���	�'�b>E�I��Y��T�u�_�i=F��V�-8�5�Kwy���X�
��I�.��'��	�nR��x��8�>�fX�0�0	�	ɟ���埸�i>��'�86M]7T����Z���*��GM���-�S�����Ox�<�'M��'��IJ;J5�A��)ޮ�׎� 1�.ȃ´i�	;R,�L�����i��N�bbI�vF@U��N�eV��O~�d�O�$�OZ�$"��>��Y�Muv^���O��J��	ܟ���?�M+�I�4�'��'���+@ς4j�
YX���:���r�y��'4�I8E�6qoZG~��M����(c�Ɔ,^����$��i�7ɋȟx�r�|bY�X����T�I러8��Cy�ٕ�
_9������IUy� s���w��O����O�ʧ1�nA+��('��u��j=�'�I���q�)ZC&.�
/���p-:�j�(E1Ta��4�M�WT��;xd��!���Z���@���HrȈ�@���d�O����O��i�<�i�E��ʣN;�X�vJ\�q p�c@T��'�B���<���'
���cΊ f�ph$%P	n �ly.Ory�s�z�&�9��2F ���,Oĕ�Eoڻ3��� P�R1=����4O�˓�?I��?��?1���i$A���a�����H�&�H�n��uN�I��|��Z�s��i�!��lS#���B��	>b�@��ʟ���`�)�S�G�$�m�<�@
N�`�+�
A#V���+��<)F�9I��d�=�����OV��ɾ9��}a-�f��l���U�'g��D�O���O˓F!���Z3@k��'d�+�)6��Ń�4qNIj�Y��O��?�����@6T��.Î�9��y����'��#�	��/�re���t)��L��'����gڝ}جE�!��-?k��$�'�R�'�b�'��>���(`�tlbP��C��h�ፆY���5�M[�#ӟ��$�O���ݹ56�d.�!g>9R��Λ��I۟������例�'��ԫ��BjY��a*N��4C,���D�b���$�����t�'x�'�"�'�&��U�3I�������3z(�	"Y���4jg4��+O��d(�i�O��	f#�|���QoY�}aP)�<Q��?�O>�|��U	��q�6��f�as2��@@��CI�j~�d:%����	>U��'���4�"�C@��"?H�{�GD�1������(�I����i>�'�"7�gm�č�.��A3�T/�
�H%K�w��d�ON㟠�'���'mª��q�<Dh�CT/r��) ��I�
Ξ�cT�i[�	*&y*���П쒟\�nT�"��yѢㅕ {T��$��~V��O���OZ���O��D#�S08�&Tڕ�C�A~����;@d�	�P��=�M[ֆ����D�O��O�����:�()
G�1�T�rT�+�D�O��4�����Oyӌ�ӺK ·';�M�cÄS���7n�{�Pp���
1��OTʓ��'|z͋a�%������ϟf�e��D��b��̟���ПT�O�<e���Dg��3a�VT�x�;�Ohʓ�?���S��+��><����-�؂��H�\�rz�n�9x�<�b�T���$�r��A��H�4eh��
�h1�Y����n�$C�	�M�B!�A۵IH2VM�I)�-\�@1��?�����'���Ο��P�Ϛs5��"V�C2j�Tj�DMş���3��l�[~Zwo��2&�O`�t�'@�
4�!Ѡ��6��2�'+��~��[�cR�m-u��˺Cw�Л�Hɢ�M+�$L��?A���?a��t��y� U�dW����Et�(��X�r�'�ɧ�O����i�� ����f���}�g�ۉ!�y2O2pZ�(Z��?b#���<�(Or5 I�Iw`s@^&;���$�'��6��	!����Oj������HR�L�[PP�G��b]
��'�R�'*�'t��i�\zC�b�b���O: ���Q�&ڶ7mS�'.I���Ox���D92!��%N�77x@#�"O�9x���]��M�k5cmJ!����O��nZ8xv���`��v�ӼC��D�m�$-3�O��6�! ���<����?��^(�Xٴ����-k D��O���� ��i�5@FB+���RB�|bV��F��Ɉ1r�(�P&P1qp�BQ
��D�說K��Cɟp��ߟ���"D�0�&�Ö��6&_ڡ�D#�	���O��3��	_���W@�?([EMW�:�8�(CaM�3d�\Q^TK�C�O���K>A(O��!+��W�"�Z��e�J���OL���O&�$�O�<�ƶim
=�W�'���9A��"�� �5Ή�U����v�'l���<���?���+H��7�4`ڵr�c���F�;��1�M+�OT�j�K��(���.�W����:]}���A�$��$�Op���OB���O��$4��.��IIsm4�8�ad��b����՟l�	�M�g����d�OL�OTp�3���Z"�����շY��,��E$���O��4�z���tӜ�\�L���3p�<1R푮�4��Lm���Q��vy�Ob�'�B`X�Rd zSo�4bt�� Q1��'��	��M��g)�?���?a(����G:f Oӓ48"񕜟��'QR�'�ɧ����u0D K/a�̨�D�1O�\�`oA 0w|6�;?ͧ ���Y�Emj�t��!fƮ�Ѫ»i�\��ӟ���ٟd�)�UyR�v�Xm+��d���* /ޠ/�8i7��%p�˓�?)��_�@�I������
"8
u1AG c&^m���?I�eM��M��Ob43�bIøO�
H�D��J��1 Ւ%�$ٝ'A�����I럸������IJ��/]0"�ڨ�H�@8B)!]��7m42���$�O>��?�i�O��4�pá��6+v�����*f1��	�Oz�d6����s.7�u�Xj�єf�Q�B�)ac(4���p�H9�$�+7��)�d�<ͧ�?����c���:�ڇ;�>� w�4�I��@�	֟��'�~7��M��D�O����6��@8�`
|$Z���4+
��'6��'6�'	p8*��	c9	st���M����Op$b�N���7�>����O�d(�
]�#�zU���Q��5+R��OX���O����OF�}2�:@X��Ǆ�	\3zT���%J
z���Zr����j�b�''b�4���� �,7dd����U�Ht2�=O��D�O�����86�&?�����
�e,���Q�[�2=Z�  9��$������'�r�'E��'ǰ� 穔�]p�U�Hẘ�1X�H0ܴh��D��?�����<1dnL�'���
��ԿI�mSP�ɱ��$�O&�D ��	�<H"�]���]{�ѳ�� $����kpӘ�B ̘K��1|�2Ѹ��كW�NhZ�f�"��A#�
Z2<�Ag/��\4��S�g�=��AF~�h�a��N5 ���ㄉۧkP�d�����Y�،*���	8�	��MUJ��O$�zqiV.I���I�H��A�"�ٯ�^�r��Y�V������>��4��L�c!R
�+�At��
I6d��[դ[�z�J������
�H�"UK�_Y��K-V8z{j�;RG�8�LP�D,�?��5�v%Ľ)a,��M�B��Ii/Uv�*q��!-����wE��,H07�De�(��c�t��v ��p���mZdy��'C�'���'���U�Oe�u�՛G��k"7}�<�:#Y���������Yyr���s%D�'�?�u��%v��p������'�&-���'s�'M��'	2`���Dؙ�P�
��S<V�@�Pf�
B�&�'��Z�0	'�L8��)�O0���R<���}آ����:w���T(VC�IğH�Ib|n�?��O�B�q��1�x�4�WU`Pܣߴ����i� �n��������������J�Y�
-r4���B Ѡ�i�2�'�XC��'M�'�q����`��-"������=E���s�i��ͺ%(dӤ���O�������'��I�p�y��E����:�HEO&JБ۴y� \X����O�<j &�0S|]�@�Ų2l1�N�Φ����IVFԉȩO~��?	�'���GpT6��FK��=k� [�}r
"��'QR�'�2�����ӌ$^��1�!��X0X7�Oj-��ks}RS���	x�i�]q%	B*5bq%�����:Ѥ�>aco׋���?����?�-OԜ����%�FAb��6R� ���֤[*T�'��I͟�$�\�	͟��Dᕅ6������0Xx�Q�c�B1�A$�T�����qyҩ�1d�=�&�R�9M��h"�ވ��6ͻ<a�����?i��U �'��x��֭\���s��߈m��钫O�d�O��d�<y���M��x�g�
g.� b[�o���	��M����䓀?���jW��{r��Lz� E��' +<uk��W�M����?�,O�=;�c�f���'��O0���,�' 9s�/H�c�$���O8��?k���T�'a�$��,��7�����I�(bt(�n�dy�IB�O@7��O.��O����h}Zc��Jta�>{FȨ��&��zNY��4�?��/�$aɊ��� �={���7Qm ��5�?�@i8%�i���m�N�D�OL���f��'剿?4�ar�C7���25��7XO���4(��a������O���I�J~XH�WIq�T�Sa��rP6m�O��d�O<�PPC�J}B]�|�If?aU��"B�T9uEOZ&�r�FH���&�8A�lÒ��'�?����?a���'BJE
W$���� �'�)0�&�'�|�2� �4�"�>�$�y2��� GM ��%��@	7Fu�'n|��'X�I��
�
�4_�썁�A7��\Xaʆ>{�H�'.��'��O4�D�����@�=�0�H���[ 
����{����W�����̟ �	wy��&o�瓛r���K�yOj�;��Rg9���?y�����4�*�$�?p><�S'V�E�pm�ׯǞ3/<�&���I@y��'94�[>��z���j`�X�#�6�#�C.gdp	�4��']�_�(�C�4�dͅRl�	z��Cz&����I~���'��	�l�q�i���'�2��5�H�$�  �Vb_1K|��!.����?�)O�����i�Q"t,�:L���%��}}n�˺>!�EP�C���?���?�����n��d��u�D`�F��i�|�U�i��^����(�S�Ө{@���S m�x��WK��a�7MƫQt&|n����	Ɵ��>���|B����hǨ\,y�N ��I�A����'���'�ɧ���X�F�K4Q��Иg	��i���.��M���?1���Xa�+O�\�$�&LR��g� b���TD�̼�Ex�o&���O���O2I���M>-�XX��N'�J �B�̦��	�6��p�L<�'�?�L>a�RTv�k�$��Gc��� A$�'���|��'���ȟ����ތk~B�S�˃r�1
�eX�6F�ɔ'��'��O�$��0���<7Xݸ&!26�٧bm�h�{�D�O�˓�?хm����d@~/��Y'��I3�Ic�G��M���?Q�r�'+�I�N��6Mܩ44�٩�aT�>���#��_-N�'C�T���I-�`�O6B��:��=�硖5|��@���)�uӖ㟼��ry�@���,�B�5�U�Y��K0�vd��n������Uy2�؟XIj�b�d�k�F�n��u@��	�ҥ	�D[?��';�Iߟ���H�s���{��`ǋ�}�H,x�Oә_4��?�r戋�?I��?����-O��]�\3���E�	 ��
*���''剿g;�#<%>QB��-(����z�D&�aӠ!���%�	�L�	�?ah�O�˓|�t��D�-h��ؖN�9S�:����i�:�3�'�B�'����O`"qM�B�x��#ʵd�0c
զ���ן@�I�n<N���O���?��'�F���ƙr9`G��,��Hy۴�?1���?	��N�<�O7�'e�п;B&�\Q�fͣ���+@�6M�O�M�0*l}�T����Ny���5vJT9j��TaΟ8&��=���/��ą-3����O|���O�D�|Γ&!���%���H�t�SuoF��c��%a��fy��'X��柬�	���Q�����mcC�;���Z�f��,�r������I���Iٟx�'<�P�Dk>�i4��,d�J���c��$k�ؓ&ejӖʓ�?�+O����O���Y�C��$I=On>`!u$Y��`��h@>}Ohm�ǟ������IMy�ʒ`X�맞?�1�v�P �To[� P�M�3c֬]o�֟ؖ'�r�'[2�ʼ�y�^>7�D�J�p�k�;�uض+Z�3��'�bW�؛��L����O����
�ʦ��������P&x����2�s}b�'���'m��i�'��s����� ��Bȴ+�ru9�&^m�.�nZDy��7<6M�O4�d�O���XC}Zw�X��1�˩:n��B��~X!�۴�?1�tbt������O��衄!�X���vDO'x>,eA޴ua�  '�i�R�'X2�Ob���D%�JX4�Q�@.@cA/<F�� oZ�T
��ǟL��Ο����@\9B'��fAha���3A�X!�i�B�'U�V�+�������O��	/|��1婝o�z2��Z?A�6�<�$�(~�?]�	ן�')�����H�q֪��W�Z-f�`oZ�<���Z��Ĩ<q�����Ok�='d���c��X}�Ԫ���$����`m��ܟ4��ݟ����̕'�"0�P?@h��gK��0�ji�bX�������O�˓�?���?f�=�I�פE���U҂� 6M���͓�?����?���?�/O��M��|R6�ŵ"tdi�Gͮ<6h�biC����'rR������(��
o��vZ�	b��m�:S'��@d��'��'�2S��"%(�(�ħTh�1��&�Й0���q�"�)��i?ҕ|B�'>��Pk"�>y[7x�(�J]�4�H��6�_�Q��Ο��'��ف�;��O2�	Y�z��Q1EX�6��� ��ǵi�P�&�(�	ϟ�F�u������->�r��c	��Дz��0�M�-O�B���Y�X�d���'X�8��#>���GL��I'��۴�?y���Xx͓����OYt,Y�D�.hv1¶�V�D戴��4?�0� �i���'���O��OD���*#�
��b͔+\5��Fu�xQo�&w4��	j�	a���?�B#z�$��� %�؀�Ck��-��6�'b��' ��;4J7�d�O��D���[�U�zi�I��h�2d6��#DyӢ�Oꀋg�r��l��W� 25i5MS"+�,3BJ�����i�b  �@OX���O�Okǟlԅjri�!��J�O���	�|&�jy��'�r�'��I�`�$�\V�����V�����&���ē�?������?�� =��v�M�̴��| ��r�#�?�)O��D�O0�$�<AV�Y��i�o���S"H̛w ���/Œ����O�4���O��C6��d�$A�*5�����D���k�CX�1 ���'��'�]����X��ħHM����)8��X(�-��,���հi��|��'����y�>9tJV	3�"�3 ���T���Ѣ������8�'rZM3��$�	�O4�IT	4��-�c�d,}B���>j:
%�\���T�g���&���i	F�9�H׹i��5�V��=@X�l�Hy���!j��7��O���'��d�>?���5z��L!:<�{��ɦ����P��Jǟ'��}�3�:��Y!�Յ�68�!�Ʀ��c�ןd�	ğ ���?1�'��"u�%��. .;�T�+�(W�P�s�4u���Dx���:��&�N^"�1��?e�6TCdl���y⬘ �x���Į^x[f�1�p?�tN�`G�#�@��Vyh��I�u��0���;H<��萌|�4�&��Y��l�eC��&�(�L�a�DL�v��-dB�	�&@����婆3h�q�#�'a|�O��	R@;��(13G�;�XdP�Ο'[��m�&7n�yXN�,w���8���@0N�z�@�1d���O����O\��c�O��r>�D�رN�Qs�p��;@��:"4�1ƃ8*�4�"3 ��ۈ����w�ѡ�I(_$hZ�敭^]i(�"��@��t���Ͼe��JF�]�'�����?A�GD21�jl��a�;^x�K&�hO��?I6c�.�f�C�̃?���e�L�<i��/N�	�R.X�@����1	�<	[�`�'D� *�>�����i�l�`@���+V�.�0�g|f�sA(�O���O���@[& ����BI�3`�2��|�#�<1�Ͳ�h�0S僒]�'n�	��僴�N훓�@� y�O��ځ���(F�W�J=Xe�'�V%~$�����*ԎW�D�-���ɥC�,M�wj�<Q��*�8��E-���YG�VT���	����ԪU�	#T���5�W��dϓuE�$JW���M�� �?1��?��a���1��K�z���֨�5WOH�"i�xܴ��d�5X�*�<c>��@:a����T�eR�0�lU�A��jU�C66\���Ђ�e����)���bg&M?� ���I�Y��"֬ue�D��ޟ���'��?BZ�¡�bH��e��4���ȓz�<��#гq��y��1!�|Fx��?�S��a
�|�ۄ�̓3�$Q�E�$r�'�b�k
Z"��'�b�'q�ם˟����~��7D4����悌m��{��ǚT7����+B{fx�a>#>9s ЖlG���1N�%[~���'�Ea@M��n�*�#F���0YП(�t�*ؘ'[z�@`mV�?���jPN�0f�a��'�bQ���'e�6�������X�	ڟ��i�ey�U�0�
H�cBR�J�v)��0�E����'l�a�F��Ei�aR�H��1����6�ii�6-1��^����w��QAf�� �����X��u�
�'�
Q#��Vx���S�^��:
�'���u�/{��h�F�I*hOR�h�'��m��M�1`ĝkg�V�6Z&}��'d�\)�H(F j�`CB;~�(B	�'�|�R�اԴ��|����G�<!�FZ�F,����[�Uiq�KXF�<i�LU&Ap�$r `��H�������g�<A�� pZ��Y�E�!D�@l��l�<Q��֔5����@aل{����k�i�<a�ښ��s��OAX�`r��L�<��.�� ��dE�9q��Q�<QAL�)�X�aa˞}�����Q�<�"��y��X<e�J�<a�F̎&��0�0cF�,p92�KI�<Aw/C ����m�[Ă)��L��<1�C�k/x�6�͔*�b�0�Vv�<�1��84v&�X Y&.�u)��Iv�<!DG([�&����
�h=�e�o�<�ǦO�O���6���h���hdr�<�OK2^܄�SB���D�$���D�k�<�X4JK�	�b�4N��4�@ϟM�<��%�{�T,b�M-�Z� ��IJ�<���H�d�*�I���+T*��p2IJ�<� vd�H�0p�ڐȉ�Y�i�6"O´����71�C&�>���p�"ON��V�Dwg8p��+7S��[7"On�1�bS!y.L�W���n(���"O�����	s��Y���@� 
 <��"O1b��C�0�tq'��
�hPQC"O�%��gB>��L���I��"O��z���gp�aK�"�bIR3"O��0 l[~���	.͘͡�"O�����Z�3z��k���L�2�;�"O�1�0��9���iK�M�����"Od$"�d�3@�b��7e�@� a"OZ��W�J�iXt�4nA���
 "O� &�V(j�,X�ïnU pJt"O���S� 7���v�'0���a!"O�5(��և)w�!hE�Q*x&j��W"O�(�Ȝgf�5yc�Ώo��p�!"O�܋����(��6 ���:5"O,:���F ~�Z7�[�(\�T�`"O��P��I�4��A��g�5Z�����"Or����ҷn�@pRB#I|r5��"O6��Ԫȃ,�n�㠩9iPA1"OR)��Y�4�$��a�"O���b�PA.��ro�=�l�3"Op��$�"]M����Ɣ���"Oą��C�6F|�r�	�9��1d"O�-Z����=�񠕗2�:���"On	��·n'����&��)�R;v"O$�@"EȞ2J���Bmn=��"O5��Y>��=�uh�0N��Z�"O�:��S#q%�QFI
�%(.p�U"O�D��'	�T2v��V��"O���C"B�tD�IE@�D` �.�!�ĉ�n � :2jˎW#�-�U�C�Q%!��r[��rB-^	��f��s!��ZXD ȣ��O�}�&�A&(J Fo!�� >��kE�A� u�4��!bt!�(��Y:D����T�?0�!����D�$�h����a+J�N�!�D��Ȋ�k��{|�DRT�T6T�!�ި��|E!QMI����[�!򤅿��-b!��6UGT��@�!���e�d�*O:03$*�J�5"!�$R�0�6
����J%r�X�
�7�!��08TZe�� M��P�js�!�D�pʘ���6Cg�Q!�n� :9!�$w��q�FB�aIE�u͒�$!�d�&3��֬�
1ND�+ׂY!���wcTXU�)O14D��ޘ!�d�*#*���B��&m{.��5�!�*o~��j4�P� p��3LP)}!��
�8yb��PO�%9o�$�e��%P!�$OP�d�g�R�x��p�Sc^M!�B�R֜��t��0$����"��d;!�䐾�:��㊀��|�
v�W��!�I�m(���ŅK�x��:ԌXJ�!���+��e���=�^�&kV&r!�Щ.�!�ҍl�1XL��!��i�p�[ra@g|�	�uKY-2�!򤅻Q���E)F�>�9��J��_�!����v|�B�ųN7���!j͹,�!�Ȟ�V�AQ�^�S�\��W��5r!�d��af��Ib���]o��Zu'��l;!�dN��~L
�`��cp�(���V�!�� m�P��=�fY��O�C����"O��Q1R28av �F�0���Ҷ�'@��'�%��DV"f�Ԩ
%�CY�`�(ǥ{Q!��Fwj��T�ȥWI�dH5	O,?qO"��'�?�?B�!^�SB�$����	$��P�Š'D�$['F�!	Gvi��N͟!?�8�[�qj49�<Y��:�gyR/S�Fd	�b~���@W/�yReU/.�Nt[!D��-4�$2`c�BUFբB�E�J�}�Yb:.�w �,g�1!�`���p=��ʛsD�'��P�	��I����v*԰)��h�'<����N*�HaB��W���{�Oũ]r�r���=#� �_BfČ2!���wh� ���<5ƜD؞�ە"�z"��!%I�n}��jŽY!�b���O*���U�#3�Ǟta��!�뒞�(�gc�_��M��"OP���O��r(xm�� ?��Pz��>ٲ�%d����� 5t��U�*a��6lwA(L�dj�RH�C�	�v;���uB�6%>1���N+���i��;��h`V�3l ze�$�5�3��7uP������Qx�B�A�&AFC���*���HQ�U��9k�M�Y�J�HG�xD�c���"�j��'�@XiqO\,<��H���r0.%8	Ó;"���d_�`����%�92�,��!��d���i�#��b��US��Z�<��W"�B��Gh@.{9��!+�R~"�Ȱ<6�NOAj��)DhOh�O6�����@[�y����z��u2�'qf@ˁ�ۦJj$�!�F�ƤX�0ăaaK�g��۔W�ec*�3�	#d.arH0;����6��/|B�	î�;�'Z
a- ؉D�>8,�����C�"�SP��,d����'��pJ�gɎW���@�N�-�nh��|����&	F�ґb��{��Ȁ�%YK����Q� �\�ye�ȊiLC�	��"�Ic-��6#H}I�
y܂�S�Ƒ�� u28 w�H�P�,�|Jwbɀ!B��H<��09�	�E�'/�,X�d)ʧb֠mS��Ȭy���"� ,q��+`�5͙�9n�^	��DL�g�:hx�a�C�p5� � _$�����q9�)�'t<nU+�-�.c�E��I�ZR$Q�`g@�"��4
H==���S�,�z�E/M^�H��h��#N��O�x�d�� �0=�2�ګU&�����aP�àe�v��H�7�.n�R�h��N�qCh�8��+��eò"O������/�YCUb�+ۆ����	��\���	K�C����g��8 H32L��6�!��R$䠲��9fA�ɃM�y�!�����
��˛C3xXul��]�!�TY�a�%cZG�X��$^�<3!��[�����W*,[:�H�JH�k�!��Тh���`L*;&��)��i�!�䄜'p�e0���pM��A5Q�!�dJ�W=Ɓ�v���h厴���W:D�!�$��>�����8���(Ce��\�!򄘬 �hYZ#��E�N���-Ρy�!�ē(D�(����4>�2�9,�
m�!�d�h>���G��fJ�qe+x�!�dõ"�R�p!g54[F)�T�&�!�ǔgAQ����!?H��i�:x�!�d��kżIi�c?6Q(��l�!�d��ܸid'ա\Xu�昉!|!���;����w�]�-R��БŖ�Kw!�ǁ3��`����q+x��D�f�!�ď%B�6��0��iuRʒ��B�!�Ą??FpZv&�=^�pK� �
�!���0�z萄`�2MuT�J� Ρ�!��̥w�b�b��E+fY\ܚ�&Ä?�!�$�_���(Ԫϝo\�9��JN�h!�;t��¼nwB�C�)
!�䋚R��B�FO��-�'gֻz_!�$�6()q�A��@�Q.~n!�}Ʉ��?B��yke%ۓXm!�� ��.�cJ(0���:+D��"O�x�cf��!g<P�(�H�
a"O6�h�� ]n��V�F�6"OL���� ����%�d�dĘa"OT|#����|��FGNv.ݐ2"O���9�@��/f�d�0�"OJ���g�+�.�)fFD�Ry��K"O������7������J.`*�"O�Z��X�!s)V�6,6�x�"ON�3�	U�^���%�ߵ7#j�b�"O�1"�e����Ψ
@�p�"O�	S���;V�攠��l`@"O�9��K�|�F���GL3 B�*�"O*��g�L7	;R`�0�����Q@"O���ag�1M��U��Hˡg���%"O�-� �[�}8����E<|�<|��"Oj�Atׂ�b��Q�^0��)�"O��`��/ HB�D`��-q!"O2��a�͸HL^������1�2yK0"O`=�+�$!qL�3׆�+]��U"O����D1^��E�@�Cm5=��"O��޾V_��0 �9G/���5"O"����r�ֆ/&���w"ObQ�$�As.ٰ�C=*�#�"O�a���8c, x��,z�p�"OH�Z�k�f��d;E�+_����"OZِ� ����Q��=����"O����[�P����_� ��"O��IL7)7԰��ad�ȑ�"Ob�;��4�`A <����"O�p3��A}��E�##��� "O�xx �%����c�ch��S"O���A�>I�psC�
��+�"Ov�qELIV����jؐa�B"OޜA�坣}J� CG 5�vճ�"OԤIAn��L�U �.L�a�]ZP"O����ְ
�T���� $|����$"O~ �2 ��+��@<�
�C�"O�ӓᗕ]]��S��S�V���"Ol4��H�"K��t��K��@��"O�X+��G)��a֏����u"O(i�g��s�-�6/Q#yBPѳ"O=���űO]���e��Pt(��"O��C����8d��v<���"Oܱ��MN�w��0��D��r3fa t"Ol�I�!ԥ;��$���-,#���"O��K0M �q:<%H��H��Xi��"O� �Q"��I����C���d�F"O�+�G�V�m�q��4�p�PT"O�̢�/Pb,uq��/&/�p��"O��z�l̉��t��2�d1�"ORY�*ɑ�= g^�	 ����"O:| ��UA��L�D�R���p"Oh�#�L��A������8x���"Oj%��
ѿO~@�Ƨ�  �V��"Ob�k���2V43�ό`"]-x!��y��f�B�IAnΕ!���j����楁 -��|�"���7q!�$߷(��)�gB�?j�*�b �ѡT!�d ]�>�c��i����a�Jq!� ]��M0�D�.�~�	�a�NY!��d� 3TO0�v�X�!Q6t:!�׏P&p����a��HC A��!�d�j���G�ōVw��r O���!�� D�Bl�q�z5ಥ ��s�"O����\?"�p�󔄌v8��"O`�j�$�����t����p�"O�b'�'��kT��?	Ǧ��6"OƜ[p������1ʈbfM��"O�qyB(�c�H�1Rp"O����#N(C*ȁs�ƽ'��8G"O6�;�U	#5xt�g�Z���"O���$�"I��d�4i��R+�d�"O~�H��֑_���`�nd�6"O�e��͜&SF���ҘO�P=Q�"O��`RB��on��x����l� "O\a!��1s���i��<y|\�5*O^�(@�ר���bqC��9؜�z�'��8J���xP�u͞?=��c�'�Ҡ��B�X��T/��/pl�
�'��dZ ��>��u�&�&*���''6P� H(|氝
��/�*� �'�������R`L�j�&$v���
�'����F�ڃ'��C��ֱ �9�'�е�wjʤy��2SaQ����#�'�ƭRB\ ����� �,�A	�'TQC҈F�	Ś�%1o����'��m	 �ON�����Ƌ�~2�\�'%����T@Eb|�2�+mJ i��'���Y �v�4Y�E�:y`����'���*��	�e�R�Ȗ`̧j��9��'����eI�r��0i�U�h+8c�'�D���j��i����/�5V���'<�$s���[(ݨd�]�5�t\��'A�! ���9���p �v�u��'� 9� 
Թ=(��� �x�hX;�''�!ag�*b�R�1���? ^1
	�'~nT�j��Bg>|�L�.�E
�'k���e2(e����H6-R|C�'7��)�Z6v�&�⌇<K*�S�'ŞY�G�n��!�G���7��ٳ�'���,�^(
�])�i�'�rm�l_5xm~�����
 �����']*s��ZZ������`�'(��0�
v���`h�7[���',|$�S��.ub��A�|t �'̢X���;Lu� �1��i.�-��'�hm �f��qi-�C(�	a�$Hj�'�0X�7 �`�b`����@��'F �����9U8�ppg�^��xd��'��ۂ�;�xiw�z.���'0\y*�+W�!� +�K��>%,�K�'v�Yy���pKRQ�3���"�>��'���ʣNַ*xU[�Ӝ" J���'>��SR�^_�؉�┧E� �a�'K6�����e�d�3$��$lbjق�'I��{�l��-��cd]�_l�	�'8��ʑ6zW,:"Jn�q�R^�<a�
={=pd��%&����m�p�<c�W�Ud�����D����w�i�<)���-#���iݛT�*��U��P�<���H�@�	��S�>|X��a�<y��Kj��x�g�653�x�A�U�<Q1��%�~��� 6*����"�RJ�<	�l�"b����`��.!����O@�<�����BǪ����'a��7�Mx�<�7�ϑq�x��}gT�����w�<����)l*�$fB�K��eӖ��J�<� �I��H�#c�XX���2��"O
=Xǃ�d��P���!n=�Ñ"O��kゝ;a�ڔ�K�4R@iF"O�-c"��-|R�����Tu��[�"O��!��?k���@1U*�0'�D-LO$�Ʃ�bH^�s�`�BN�h2w"Oh�K&�=J��ip��IJl�!"O����G27��h`엽G�ѱ�"Op12@��0U�����J�-i0j���"O�1E`I'����gJ�2{ !�"O^���M�+w;4��c`��}�0� "O�����5:ڬ�[w/A�w��q��"O�p[���C4ʑ0�G �v�>tBA"Op���/��
5D�����>za!�D i �uQ��ܓw@@��V�W/!�D:8ˢ�[�[	�n8�Cf��!�$�?Z4�x���R,M������-m!�$� LNn �f��8O�Ҵǋa!�D�(#�)�Vaõ0_�0 �g^!�dM5���Y��8U�q0P╯@!�$��a�>xq5��JS8�뇆˼N>!�G�}�cC� $9�¥��Ғ�'�v��YMg��!$�T�s���@D�HC�ʹ*�q+�OA~���>Y������:E��T�����fKl%�2�Q�yR&P*q���ڳ 4�ZA����2�y��H"�fĀW�By�����/�yr풊=j\!��@X�s��)�@1�y�O�!b5�u:�.¦n�T� �6�y��pk�	�f��W=��J�区�y����lN}򶭒�;����� H�y�kQ!�zJ�$�� i���uʃ��y"܀m]\�eGI�u"�����y�Y�r|*�Jͯ|IH�bK��yb��w!p�k �g��r�+��y��I(v��M�1m[]Ԝ`pmT���i���O��	�`��nҥ�%aȜb�jx �'���j�΅�����a���WֱZ�'�]�wf�,u&rTJ��ʄ{�b)�'d���b��zT!�0�	�]�X��'+$�SL��V���z��לJZ���'h~5 &W�g/N�Q1��.x�\LJ�'�Q0�X�SX�8�c��j|�-��'���1G�C0!nxtJT� `֨��'�,�j�� m'Ԅ���!Rh���'cb��
�m�����T���'CH��PE��G�� IѩN�H%��'�$�pFS�\��"` �>8$6���'en� !���y�"�9Ghߒf����
�'��8�gn����D[�ǈ�Z����
�'kjC�LA�f��݋��& � �	�'�H��1�=��d����x<81��'K|E*S�ؚo�\ѐ�Q�u�V=��'�N5u�A�Bi�t�6drl�D�'�Ұ�BeS�� ��a�p��p	�'�>�铪X+���hĤĮj�.P��'p�|{��P�V��]�D*dM����'N��"ˁ�>1r���Q��I�y��'��q�Ј�Q�������JR~)Q�'I���v�DW�H��	�xH����'�"�Y��=��!A�������'v$��a� �,���\ tYq�'V�}AM7~y~�i�Eʈ(��'$�pʖ*,6]�%Ȕ:���
��� | {��
Y5�<pGL�1[�b1�"O\���-EP5��ߥ:�L��%"On���+A�3�qC�+�O�0ёR"O�a�F5����g���X�|I��"O���&D(z��Yx�^�|� �"Op!p#�Ϡ��#�/kb�3"O��!q Ɔ�����b�>o��K�"O��[5�H��A8���H���s"O��06�H=z�9��A�*�t��"O�h��Ô�>��R�I2q�d`�c"OZ�ے��<��$�M�J��4
�"Oi�q�:C���̄)��%�u"OLl�w�);�0xa5�ǿ���;�"O�HE�֎E�q*wH�1(~���r"O,����]TP�#�ܠq��\ir"Oܴ���@�:`�P��u��|`"O�����K1�iCa��>�r<#V"O^�������\bU#ג\�H�"Ot�ss��%?9�i:!C�.��9�"OBuZ6�B�M;��'AǄQ6��"O����#�=M�Ν�)l��p�7"O`�[�hʊJ�(���>M両!G"O^@��Ʒ(�4\S���-}юT��"OF4�u�+}P������*6ն�y�"OR� �%��'�(_>D�f���"OҰ[���	� `�4MR-]��H� "O���Hܣh"��2�K�g�H��"O��o�z�����e�%�"ON��d�L+��HB�թ�*LK'"O�p�Јĩh_ژ"bH��q�Vd�"Otx�f�����fU�}:�a�"O<(x3NH�^�� se�GP)s"OiI�+��х��:J
j��F"O���'-Ipp�,9�c^�"R�帣"O� �1K u{���C�ȄaZ��"O�a��#�?��𑲡�&Q�
�"O�a�ǵI�j�K�!ճ@�����"OdYӶ��u�f�I� ���@Y�"O�qB��>u��Ԑc �!��3�"Oz%
F�	�T󺨑�.��o��Lcr"O�KgM]@��	2���bh� �D"O��pA"�����8��ej���"O
���Ap:�IS��Ý#�~X�#"O�8R��<qR4�w,�#�x�'"Ota�G�X���f��|� Ux�"ObaB�D�!".�CG"͟p�颂"O�(a�aصR��4��~�X��"O ��	�F���1�/�	Up4��"Ox�h�ár�d��5� y�p�@�"O���ЅLE" "�j�RN��A�"O< �&�+\S[0���:�"�"Oq{��#nJa�V��'&���"Oz2�X4+�AJ�ʌb9�"O�� �2И��1�ݰ}�1�U"O����Ť`I�1dq��9�a"O�,IUd"$�cf��L��e"OȬ[c�8X�DPbÊJ#�EI�"O�U��e��U:��Em�ڼ��"O�}*���]���PH�#F�Pdb�"O�l�W���:x�p�R�U��+C%8D�Xh��
�mk�T�D�+b\B��S&5D�D��W9a�Vu��N�v�XP��5D��d�.&$� �Q8�k0�2D�\��)*���cS�d��k6�0D�� (9"e	�3�l@X��#閉�b"O���r�äSO����D6 �	�"O�%`�ק7��{@�vvASC"O��˔ثUJ��9��J�g� xc�"O��bE�/ ���%k�"8��"OX]��"�9"�$(Є�Q�m�S"O��̂`p6��&#�-��QJa"O���S�#uw ��4���O��l0�"ODi�I����������"O<�J��٣+=p�˵�@�w�^�@�"Oh�H�޺}x.x���.y~X���"O*�P$!��E,$�C�ƴ²)�D"ObMKNłn�������;y��0�"O�uQ#$G�u?le��B�	==BEk"Ob�"���
ܐ��da��%3�P1�"O�h3�oW'HvA(҉H3j��]�v"O���2��7)�c胖n��Z�"OB<�� �--���!��+6xr"O\���!O�lP�d��~ �8�0"O�Q����S2u Y���)u��X�<�'ȝ�U�^4+�`�Yy( Y�<�ԣO-trP	b-��Y�V�XRkS�<��A�'�1ԇ]:%��h���O�<�6�Ab�B-*��6F<��f�G�<�B�*0�|[��Fmy�EE�BD�<i!a��}b^�2� H�����@�<�ac�Zm�����>)��33Ç�<�IW.S

����C����D�e�<�Ɣ�\H5�r�Q�~��p�H	k�<�a*/�8�R��D�t��a`0��g�<���Y�tN4
D�Ȩc�5��O�<��ҡU����D�
�78 �3[t�<q0�� I��x 4�ğJ�����
s�<QE�Z?j��o� Ud,t��G�c�<y�ЗBO��ڔƎ�f���(_�<	�ǂ+]u͊��F�+�,(�d�\�<��B�6�a!�P\r̄y�l�~�<)0�^�V	�oW�O_p9&O e�<a5iA7p���5���YK�ՋRP]�<AT/�-Z��z��Wd���s�<)J�F(Y[��P���p�<�FN�=ZH�(6̆�,K�T+1(^t�<Q&�]�E� Y�Ѩ�ucd(� p�<y�܋ࢭ�%D�#Q�lc���m�<)�J�&t�������"/PX�d�h�<�Eꈖ�p�P'˫u��E��Hg�<ٲ�D�,�Ie��&n��9Ab�IJ�<)����nX�恜�x����,[�<����Q9&a�䏑��*A�	W�<a@G�l�2}��`C�H\���*C^�<�B�U4�89g�;���KE�<i`,P?莁�W�N�pX*0����C�<ɒ&Ǹ]�sM�L���%�g�<A�ſ�R���Ή�H�:	@De�n�<Q�J^�v`p-�a+�;5+3Pk�<)H�=��9 ��T����JPi�g�<�w����]�U�	32,!ՆDx�<qWGѯ)I���V4�l<0f�Ny�<�)�(��R�$�@H�#/[�<�e��0�t��B�81)��X�LD�<Q�Q���UJ�O[�7@��(kE@�<�e��#�Hdi
�9^Q5�FhQQ�<�Si�����(?)�2�Ӑ�I�<qᦌ�N޶�"Rn4ܒ�SG
C�<� ���g�.i�@�Ġ�9|6���"O&<u.� R`����#�2�23"O�m�Ώh�m2�o�8�l�+�"O�	Z���$�`�ƌ,�����"O� �Ą��/��(�nИe��	j�"O�����!�d(A�*	��c"O���aS8���4,�0���B`"O����2k�*L�c�8Nʸy"O�lAe���cV4��%����G"O�	��88X:���J�����"O�������(Q)q#�_��"�"O�U��M�'i�"`�6��� ���{�"O���F���@�@�	)����"O>#3ퟩ�2!psH�>���S�"O����00XR��6h�Q�&"Op`��芊���W@�ut䥡E"O��qO��2x2{(]kC�h�"O�!I��ժ � ��腶9	t�V"O�[$�M(5/�p���X4
z��"O�Ѱ�K�y|��a#�Z�P�"O�-	�lf��nNuz¨R��J�3!��ϩy�*̩���4o� ����Ӄ2�!����P�CK@7|y��0$�!X#!�DݺJ�B	���V,	��yDC�S!���ؙ�(�0: ~ū���J�!�d�kMZ����T	�b����!�$�=��HZ�A���!&
�Py'�T���Ђ��75x�����y����5xD�H/x 8���ǣ�y�L� ���@LR$�pt��*�y��R�Y5~E�栒k�x��0��y"$ڷfM����(��yEF��7d��yb�[�no�Q�*Y�͂���D1�yN]�Q��L�Ei*�Y#7���y�
;U2D�<x�� ��:�yr��%|2�����)j�l�����y���=[X�0S�K,Zpl�`\��y�� �yAr�P},�P�'ش�y�搢S���Gp�ș�`�F�y��������i�`��b��H)�y(K�1�
B�k$aȶ(��yɕ�e:��Ă��-� ���?�y"�F#3ȺA1�� /D������hO*��I<p� �cq퓓i�$�Ì˳'}!�$P06=���'�|e�����!�$�!u��B/>(�8��c�-�!�$$�tuy��UK���`w"J�{!��")�x�pE�0:N�Z��3!���*֏��~ X��V��e_!���#gŶP�[�g��[pLڰ.wў���������ʆ;�����X"'��B䉓HU-���K�!���#C��M��B�I2I�);ע]�z0�����П]a�B䉜i"����?p~V!��I0�dB��2�n| �!ϬTn}�#�Ղr�2B�	~a�1e�ҟ���a��,/DLC䉊|M�9[7ď�5w���A����B�	/w�0�U�&2p�����6w�C�	�b|�@)!a]�0���Ȇ��B�ɂy�4]��
Ȭ{vHa��<*��B�`�`���� c� u���@�`V�C䉘*�\��ŏ�G��,A�K�5)��C��0=DQi$���#`�LS� ��C�I�ZL�`f`^�:`�QX׫�	d��C�)� <a�"�T�:����T�D�2lV��7"O�0 � Ed�����T�'"O�|�e��_.pX����/ǰ"Ox,�����x�x�p�gW z�� ӳ"O�	ٰJ\3FT6T������T ��yR��7ۼ09���*,�0��s��>�y�eӬX��H�F��%��9��'�b�O�P������c��G��	��'5TIb&��{�v�Z*ܸA��89	�'���R�+�1�%��'���B�<qT��:_!P@��e��*�����y�<��͍(úi�ȓ^'8��v��\�<C���F���q�!�v�Es�tx��'0 ���Ʈ:hD�׌��壚qx���'+�9k��5wD�r�c�>��!�
�'���O��5�|qƯ�AbD�	�'������k�ꉻ�Η$���)	�'�Py��d�Oj���kG�E��E��'��ekA�A�h候BsΘ�;-.e��'~ K&��"��z�4\Bt��'��}"��طpᶼ S��2�Z8Ј��!� -��9E���`"�ΟM�Ѩ�"O`��	��+�̓<B:D��"O�q�tN<	须� M�A�$"O��y�$�a�.��� ���P�"Of���� ;x�� ^#%ژk�"O"��h
�cYJ�ko����u`"O���䍆FpvARp�L.,޼ѲW�'cў"~z��E���K@�Ìo�	���G��y�, �p��|�����Ę�D���y2&ʗq��iP
A4� �׳�y��@�Lθ��O�s�vE;G
�;�y2�K�~����qM�?e��q����.�yRn��W(4h� �ӄb�4A��ǿ�yr����U�3I�P���a�( ��y�	x���Ez �zD� �yR���w>P7Õ�:�R���S��y�l·SI��K��T/Ԉ�ѓ���y2�A�_�N������7^�IP��E
�y��4��d�s�T� }���P��y�K\8�!fî/�J�hƇU4�y���_X}���0\xBu�%����y�o�j-6�8� �����
�yGC�4
5#3!B�B�ܝS�.���y����$�I�,�9��}��BQ��yǊ+����$�ȴb�dӔ��y",� |.V`B��]�ezԅС��<��Č�>��PJ�l�,:�4�#s�%.!�d�G���:�&*���@�b	��O����IP~2��6T =4��rGn?6X��Q�u�q�Y�u,�Y�._��q��W�xtmG"�Z�j�K	��m��B7&	[ I�I�D�J��΃�x��"�|���K/��)�!�v����!��w�ĦSb��S(5�J���g����w���*d�T5)˰lO�y�ȓ4��%�����Q�9�r&ѐz�����1o,�6
��K�$ez�؏<��	�ȓv�|��B�L�~n�uh7"֔jP5�ȓs�֭"լ�n��Ӈe\�@�ȓ��iїiF&v�ܩSЯ�j� �Ɠ.	`�\<>����֏��#��P�'0$��o� �t0�A�n���'+�Z��O���x80��q������ 
��`N?92Q��$j�p"O��d�2o߬8r��	gF@�!"OR�|�>L�g̀Sf �"O��0&�R*M�Xp���OW&婡"Op�s2�N�Z�Ε����
i�! %"O(�K�m �aΚ%"&j� l͌���]���	lR\��*�-�`d0� כvU�C�I)/��D2�d��0��"!q$C�	� ��`�d��R�$q��/XC�	˖�㗩�'}E�P�B	�7FC䉖aP0�V�����:�Jڗj�B�I!�ހ�s��/OI�h+CM��\���'�j���r��^����J	�����X<��j��w
Py�W*�=�|@�U��<�c��6�:pɔH�
+)`��|�<�F�AA򩢕e�>�(u���u�<ѓD�W���$L��N�c��[�<��N��Q�\��iN��(ɋeH�|�<�	���2U�(o���M\C�<Y��n�d�����z�CԭMw�'���ӢW�(�S�O�)jZ�� I;rH�C��8+��	��F)+9J��Y:V�C�I5���t�`������\mH�C�	C����&�(q<���Q��,]�C�I*b�|@�-snSW4PZ�C�0q�u3�I�I�S#
V���C䉢�a:�C�(u�a2��%�h���<��-(<��o������KmbC�;&��wD�#-��=�5�X�R�B�I6�n�Y�DTz� �	��C䉝i������2�y�fӚ6/�C�I�lhå�'TA�)R�I��_��B��ML��2�=i��ykr��=�`B䉪b=�)j��:Z$�È��C��'p��$���r�.����kNC�I�5>pH%W%7|z��Z�w�B䉛q�i��A�y�����"�bC�ɡ$e�4iƃ��\pkG!�$Q\C� ]T0#0��+)3p!b ��FC�I>:� H�e
#P�h`a���hQfC�	�w���{�B�t��g�Y�V�b��p���!�݃fi���ÀO7�rѰe�8D���ҩ�i	�}�cM�
�2!�Ո$D�p !�47@��9��	4`q�}�A�#D��`�%��!����ӭ���0��!D��s���o�x�C��/|��� D��I"�G�,���D߳o��XX0d,�O��	�_�j�2uDE���8�S&V�xB�'s�y���%"����v�Í�C�	[~V��I�K�9a��Ǵd��B�ɹ|Rp����-n��c.-�C䉺�P�I�i_8�Z���X�C�I�#��1cu�èD�dQ��&,B䉰7@<���0s�6EJ�,Ջ�C�	9���8L	>�1�e�W�4C�	/lTf�8�V�(�hCT�Rg
C��'n.��J/n��dږ(�p��C�	�>�T `�J�I��@� Ɔ7��C� Y�l�����/34��jđ}�C�	Y�T��ƽOE\(Ir.A��C��>x��1'���$ԫ$��*@HC�	�N"���3��CLp���3�"C��?
H�⧆�*b���#M�.5rTB�	�+e@q� �.�p�
��Z<Z�XC�)� F�9A��@���uP�Ȱ�`7"O��9�I������KR�I�����"O^(��)T�X����g
�%��"O���Є��V?P}��w�x�Q"O0�BC���h3`T�`#J�3xZ��1�|��,�'6I�8����!��tx��N�>����%S�,�Ђ(�hI+\4h��ȓf������K�TzA�)$�|p�ȓL�:��"LC�,\4͌�7Ĵ�ȓ5�>�tM�iVHZ��ݢYxYF{��O�D#ƀ^�#<j�4�S�B��`��'(9BDM�H�aeG%Ag$���'�Н�$W��ic�g>;)(Dp�'����0@ܲS��Ź�C �3�V �
�'`����P�h�\qA5�_7*ɶY�'ι�p���6f��TY��y��'�6�
��P�Q�$ wa�!gy�M�J>q����_�*�x5թʺ_��I�yM!�ğ�&n1ˀ/f����M�+1�'��IX�������R�(�5(�7]fl�c��2�y�d�9:�T�A����Eh֙2!��#p�68��A�h�`S�\'!�dB��.�J�	!M�ΥHAj9(!�DM�l	S`왆0�^h��;,�!�13A���-BE�8B��!�$
/>�ҬZ��R�&C�M�#&�C�!�X�֤(so��Ǩ�� �]�!�Ĝf�Xc�� �d���ˤ�F	!�!�$�X�z��$��d��e��GC��!��:H����č��[RA�Ռ� �!�d2A�ECB��:s��H�i�}�!�d��@7L!��L3kf���e�v!�$@�%���8`�A�/�|���\>_�'�a|2g>v�Q�nڨ>7r��ϗ�y2o�	p�t��%9~�ɚ����yB�F�!<&�DÙ�,��t�eb���yr�_�.��pp����*��Z%a���yrǁ|�����s�4��)���Op#~�7Ú w%���ǟ_J�J3��x�<qAmC~e�Ci�<h"f�u�<ё�S�G�Vis��"�HM�UF�<�"�2>3*M� `�Gt��Ņ\~�<qU��,%FN�ᵏB)oW�����\D�<ɶOQ�I.�X�'#y���ACw�<�4� 2V�%���� �0-Hv�<� ��tq�	th�\�	� Fu�<���ȓ5F��������q����(D{���ɺj��H���E�8pI�<^�C�I�=��;���}mj�P����D$�B�Ɏ-:��?Zp$�q�ܑ9�ZC�	'5)�uQEcA�?PP��]�2C�I�;cF9���9��e�1P9ғO��=�}�W�Q<zFJ�U��z����a@M�<1(�d<��ħ�%:�li�NNGy��'��i��c[6��p��eԥ����'|
a�_oJ��ă�:�F���*fųc#�t<"qH#,۟H?�,�ȓg���Q�BH�"+���L�Ҙ�ȓ܂-�a�-y
�@�@��@�`���tM�¡�?Q�d����8Ś(��@��E@�䖶sI�	��B ,{�|�ȓx�J���D ej6I�e Q�D�,���h&dh�q�c�� ��E�u��_���Z�l��QfF����=�8��S�? b�cT�K�p�*M��!�p��"O�ѩ@n�~��љ!��8Ed��"O�-i�� i�e��[�5x�"O����I�-#�A����$�U2a"OFdb�-=:�q-��`����"O�	sE�F6Bвu Ӣ�[t2$�"O�!�C �̈́��dV�(r�{&"O��J�8l������(ydb�"O�i`C���\9zxyF�C0eA ( �"ON$aQrAL�{��62���"O؉H�!�^~@�aM�75��Z�"O@%��
3�D�S�J#
2�Y37"O�ٙ1��00�0hg��2a��&"Oz� �I��8�9jp)Ţw��:"O\"�mU�]	�����);���#"O�\�4"͛�:�)���5^�p9�"O��y �ΦF��s��#�ޱ�@"O����C16��4�3��#r}І"O�`��8J8���ɽ"�е�"O�u�^3P40���?a����"Oro�2!�rL��$D�_� 9�"O:�9  �"K��[1c�"ʜ��c"O��a���!U�	�BՐ}����"O�l�k
�6��Q���Lr�tKb"Ol�k�A_�u��@���&P-�"O��kS� 	'P�`M�N� �C"OaEP�o�\ ��lE)r�j"O�Mz��ڱ��T��_�_֜�	6"O�"V-��m�1C�3X�j�z�"O�aU�>F�B�y���M	 ��"O�Hjw��:]�L-�w�M�}�|!���Sy�ӕU(�50�OF*L��1���9'��?����;k��D�B�
�v�J��%k��i!!�䐉!�<�a'�S���jq	K�!�d��2���GF�l��0��ږc0!��t�����ʌ��$���(Y!�D�j*2��AU-��ҥ�{B!��-��h��Z#Ђ�k��|V�'�ў�<IN��I�F�St,�	R�m�� S|�<���-[�`��j�9�A�DA�x�<q�#P�P�y�/�,1��#���Z�<� �VҼ���@�_�T�R� ~�<9��S�f]� a�X�\z�Bv�{�<�!�8Y����fL�(��yh<!� Uo �b�H�t�I��K���hO<���O�
�A�߸6p�s�-\�z�'�(�@;~�%�sh#$$8K�'�b�*�����dPӃ�St��'(H�b"��e����oŹ:*У	�'j�"LTI�p��%k�d��'dڵ
7��.�0@��Ŀ��C��)�DNƱ.�FX���ħ�n=1�,���>)�O�ٗ#ãZa(��U���;�x��"OΌPR��Hrh��Z�I���D"Oz`�aK͏dڶ:DB�?\T�j"O|92��V:z�}kT���i@F�A"O���&C���|�s���s/��a�"O���Ӯ�&ذ�a�#T!Z��F"O~�ck		m'鋷DE�8\d	"OhH"T/w�f��#�a���B�'eў"~"�9m�F�C�P_��+g�ׄ�y�B�:w�zxK���&��HK�&B��ybᔄT!�Ȫu&&���r܂�yߒ��I�h��3�݋�y
� � ��	A�t�PQ%�˓W1>\�u"O��CV��9$�I�ӧިn�H1@"O��H�l_>u*شxV�ʹ�p}�""O�y�B/�3bTf�0�ݎ�t�9�"OLЁ���E���2���g� �/�y2☀.#�+A���5��hr�@��yR���BѾ���䚩bE:���`۳�yrGP�3�,�KVI� �pRe���y�L'�d8�El�
>�ZIȄK���5�O8TЇ��hG�08C!<V����'D�Tc�f�ul�"�A��u�����("D�T��DԇC�Qj��_�BxP�	%D��� AD�"=@����f�Z�0�$D�$R��Ɗ�F�N�1U"�IeJ%D�@�n]f�qFǅ�-����"D�l����L[�a�T�Ĩ�0Ta�/"D�`RC��:M�MXbD�!�I�b,"D��avl�J�|$���'q�}hE� D�@b�Iˡ=ٴ(ZE�?DӺ��e!D��;�-8u�FhR�e��q���=D��@p& �1c��KR�Qg�Y#0=D���rL\�e�r��h_�UR��/�O�=E�$�K$N�8���չm�p�RČQ�!�dז&�#����I��L�c��G��O���d]V�������R�{u�p!�>=��m§aH�I`$�[�iN)�!��/v�͑�МlZ�Ah��)�!���!�f�����`y��N�*e�!��G�"��rdK�)^hd�'DX�!���:r^��qb��*Jn�B��e�!�$���6RG/f��&n��c�xC�	9#D��
�%*?*�a'4vC�	O��|��@P�+�����P�`C�	�2v6h*�"ѳ�px�Q���6�2C�02M�Q�d"�g� _�B�	�t^�e�A�|^Z��s�"55�B�I
A��!W�]f<��2M��B䉗U������P���4JA�=+J�B�*[g^�b�U!���qD�[�B�Ig�i:&���P٥o|�.C�I��0е��v�,dY��5�(C�IH��	ۈ?Q�eZ5$ݴC䉶H�Xr�������;z˓�hOQ>���Mq��7Y��S7�Wq�<q��7E�
�#d�Ѷ:� �7*Fk�<�t��T9�u����z���� �g�<ybX 3����}�-����b�<I��@^2<*�-H7	� �YZ�<����Jnx�*����s)�@���T�<Q@�ɥ}B���E�.d{PTkpT�E{��	�>B�s�	�Y��ӄ��W!�$;��`3��y#Tȁ#? �џ�F���`����+ ��8"bV��y�JF�n@4�)�/G�����c���y2 �X���[�C%AD�0����y��W� ���i�0��O��y�M�=�,dS�EB7�����ʰ�y��̏EH@	�hN'u2�b�)ħ�yRm�<X���`����V-V��U�B��y��þh	�J�7�PM�A&��yb�\�:�p)��='�>Uj!�¼�yR�b� ��s"�8�P9�� ذ�y"���x���'
� 8�Tg�V��ybe�^w���2��@EG=�y
� ���DN�<�B�)0�X���J"OHa���C�&C� y�˖�9u��Y�"O*�8@!�!o���0���E����"O�E��AޙiRHAcG��g����"O �k��F�?.P����1��D"OV]����BVd5I��_�V�.�`"OH��mOJ���m�*I�����"O����ME��˕Q&!r@9�p"O<��#�"e���u��:mt\�q�d*LO�����0=���7�Z�EBT5"G"O�P�B�!G����� E�e��"O䁲���#,������˥V\FX�"Op��ՏK�K�j�	˫^`��Q"O~%D�ѝC�
�aa�%WF,5K�O ��)�%�ƅ▂�|TTX��f'D��22��Q�0�@�/L�"�k''D�p�S$C5%�V`�e�%P��@��%D� ;@�I,�԰���O�mx�GH$D���6M�A����$�u/�Y�"!D�x ��"��҅H�P�ƑʖN>D��C����1�еiS2Þe�P�)D�)!,�.C�X��b�{$�A((��Y���XS�Q%}�`a0��°��DK!D��ƌ&u(�p���S�p䛳�>D���c[�ff4�� @�V�.u�Ď �Ib���)�g�6/��	��@�#o�:7c"D�0��XV�4a�)ެ# ր��2D�ԩq/�;�ѓt��F���/3D���gG�#l��-`��8.4����$$D�T����hŐ� U?,�d�"D��`#[;(1��vkT�V�<��"D�x�ҀS�h�|�Xe�;e]��9�c�<!	�L�m���/T��F&g��ԅȓTK�P�G`�
W���"�*
v~��ȓp@�8��Սm�@���ё0+��ȓ�%�YYl|���C�n�*��ȓV�x)D�9~����@�<%6 �ȓ�P%y�� t����� ���?����~r&�E�2E+����2`
���q�<I�&�0�i�È�!D{R��F��C�<q�m��*�v�r�E�F���JRx�<!�ۯkgb�sRl�3M"`��a_M�<1�%Yv�艈& B�o�d� #u�<����j�`0, n:�pB!Qsy��'�~�a�b��(���G�J�h4Ƭ��'�$�j7��bd&��O��"�	�'X��2�"MH�d3��H�7�����'x0�bw䅐w��yI�ځ0�*�j�'���V�S�$ͨ� �I߲ �؊�'mV$�1뉳�L�ȁ��
c���	�'�N�Ps$V�5��8�3���U��2L>��J��'f20�^(J#�'E����<9
!S�g\)��i4��#O[h���,U>�"l͹0�9d"Ş�:U��E&�����$rf��wb�?�R��ȓ:�L�@�Ѽ+S�AY�'�3���?����~Z�J̉�,�Xq5@h�"F'-�!��2ɎY�b�2>1F���&�D�!��e�
�Kת�7��%�u�/'!�K7����*De����O�B(��m��r����N�n�7嘦H�Vy��zҼ :�ΝC��]@#�� <DԆȓB)��;g�&Xx���]*q~�]�ȓ&Z�q���R��.�cé!�D&�T��)� �4��hڇ9�BKL�Vu��HF��g�OCHe1EDJ�"P��s�4J�6�q
�'��a�U⋼|����&S�H��
��xBO
/1�048�aB�m��0����y�C�|�֨ɴܡ^{� r�iժ�y���&�԰�q�C�+����R�4�y�/�n�Vq�a,�0*�ZA�A(K��hO���$�<���B�.QčI�!ڣ<"r�)�'.q�� l�T�Z�	��F��!�'(@��T�>u<�á�X���HB�"O\�s���/��Y�6'kn��""O�E��/�:�[��0V���"O��r�HX �&h�d�@��V����'��hr�e@j�`90� X��M0��,D�8G��;}���a�������6�Ix���O?�H���O�F�I���8c�0�j
ϓ�O�9¤��2v�=˴IЀG����"Ob�цG^	Tڜ�1�G�?
����"OXx��"�|E�)���i`��w"O�=��	� LI�F�$R$ ��"O�P�`^�9�����5?Kj���"O:�ا��/�%�T�*|���a "O��Q�E�>2Vh��AƬU�2���|��)F& ]�"M�8L�
��Zo&�B�(9�04��Ŗ�0	�͢�Ew�.Y��Z>���iwhdv	I�R|T���'~������F\@apEi�M��d�'\�b���rWBMq�KP�>�q�'��a�,��6`��R5 L���'!6�#3 J�dQ�����,�0���'���P�ͥ~�u)bN6SVH}x/O��Dφ����CE>,I �B�hW�u�!�ā���kn��FE!iN!���~�<��ҹ2�h���#��oA!��n��RP�<z�N���ʱa��{��$}*,�ժ��<��(�R��{|�yB��&ib�]�b'�g�P�ã�����B䉏}����  �&$�hH˰a9/U�B䉅�
I�u璯0�i['OP;}^C�	�7��)f@���
�#*�B�I�i�ݫ��H�xTH'��q"�C�ɖB��O�G��T����(�jC�I�� �����=�D�K=���O0���8F�@�*��0/��0L<)!�DӄgK��XԮ&o����T�"�!򄁯|�Ne
1h�`h��LA�8�!򄙸B3p�X��@>�6��"+&!�D��g�ɇ��
G$��QR�e+!�d�nVvɣ$��r`,p����P�!�$�0F%D�q��=+���i� f��yR�Nc،��!��U�2�!�
хP&�B�ɀ�x���&X���ґD��*y�B�I�>4>��7 �IP�)!w�z��C�I�Px���Və'D��1 #߅e��C��4xق���*F0Be3#P�FGZ�$)��hO��2�-��NA1V�A���+W�'D�`�5+ �tXE抛Բ�ѓH$D��C�P!(ͤ�dΉ�1X\d�1*=D�p�Z�A����V�E5"fx#�9D�,��^�9AB��X*4�c�F6D���x�@�j��֊f���XF�2D�8ZFGU	ofh���A�M��I;dN1D�|r3#��$�5)͟�Q֕�g"D�xᢡO�k>~DC���z~йS�5D�� ~�Ȑ��iEx�2�e��"�"O��(��=_�T�FHJ�o����"O�Pô��d]��֦Q�n:JG"O��� �BW�԰ԆX�W�⌓"O>�9u�[8A|>�c��S�q�εӑ"ORK�f�Mn�Y��B�1�b��W"O��y�(�� ��I�FY�z�Y����G>�q�L��c�B�E*j�)2$=�I��G{�Oa�	K�$ƛN�<�a��E�z(��'��ٴ��"h=Ҙ�S�L4<� ��'�.<yU÷�diҡ�C8��
�'϶���+��&�h!�mA4&Hh�X
�'���&b.�X��#
8]�4��&<O�"<�.Z 4h�0��+n�<�իAL��S���O3t�W��x~XC"��,$@P	�'V�h�n	p6z��b\(3~P��'�V�0�j�!Gȩ �l�$W��'@������bT�� ���VEyP
�'���г!kLz$���Z�JL���'�̄rAl+qf:���G�<�8�j�'����F�.|?��e�1*�``C��hO1�>�"d\�؀	����x���މF{R^�,F��A�� �&p!��҄G��Y�bU/�y�.��D��Y!M�="^,
1��yB��n�t�Zre��4�`�����y2Nř��u���uZJ�dOG��y�W���P���@�"y��?��?Y�'4 q���E�����ԃ�,9EV�@�'�UҳIM�~YxT!!�l��'�=jT���5|L�V-�SNz}�	�'}�����>n��9�hI�8*	�'�NDE�ڒ!�x���ɖ4<� �	�'Hl)���$������:ؔ�s�'p1�h�<I�>@F)Ө$��8�'����i�	!�ލ���Dut.���'q�É�*,��f�gW�|��'L@�c�k�`�<��dK4h��ٚ�'�t4ݢR�ȻcH�^�HX*
�'O\(���
Aؤ��h���d	j�'y�m�Q��+L]��H�2�@��N>)�i���ءa68��aAbM�^��ɇȓL��Lb(ômo�T�&�I&g�0���o 艹�&�����H2�ޢ3��L��n�����4kȶ�KQ��9K�هȓeX�����V���u3h$���B�LU�%g+����N�9�Y��o�@�T.ՖWbt��� 8B�܆�C���i��NT@� đ�H�XQ�ȓl����!�&�Ȩ"rA��R�X��|����`1I�J˪x�#��F����M D��QB3T4��߄W�����<D��H`�L�F���sf(	�|��u�9D�P ���>II�ͳwǅ�%��ZcN6D�ț%,ۋ_�F����9B��&�(D��A�����D�@.$	p㳊'D�<��='��Do��@� 8�$0�S�'W� 8;c(��-$��3��	2ip��ȓ@
*	x���k�N1(s��h���ȓv�t���ްn0�( ���v���ȓkf��E�4(���ҩ7P��ąȓM1��8�ƣC�zQ��I�B>8��w�u�"/I* ���\�8ąȓy#=��NX�BƸH��\l�y�<�Ì[)Pz��&M�^���B�B�<� �9��b��+%�\"B�]�~xP"Oʍ(���"�A�ذ)���"OD$)��� K�$	m�A�Mf��"O
��a�ҳg J�"����1"O��C\������Ä�#q�Qb"Ob����f��vL�8B��	C�"Ozh�fʜ)/>Y�6?TT�X�"O*��eW*`	�&@�->Ե@�"O���ȋs�Uz7�Ӧd��4"O�h�GfM�v�N����c*�i�$"O�A{��W�R���bB���|l�t"O��(��T�+�Buk"�²u�zTb@"On�hŃsxU�Eͅ�H�"��"OdYg���L�6yȃ	�_y��"O.�&(#\B��Vi�'"s�	c�"OZ��f H\u�-{���E��9�"O ��BM�5g���۵#-�
\��"O�T��� Q��I��'	���"O�D�1�_�n����#�s��D9C"O���e�.yR4ᑆ��#i�l�s�"O���w�-�6���]Mq�q"OV] �-�2d]P���G�Wi��Q�"O��3&N��Z�@���.��aV�)*"O�yE��^������ջ�(Ұ"O~Mq���	?�}�d�C+l�� ��"O2�R��Wv�`��d� �"O�rv�Js|�s7�B�p��d�E"O$�3 ����z����Y v�� p"O�E�a=}ptJ�<kv
Hق"O҅�qN\�c8L!���)e>�""O0Pڔ8��9��j!�`6(D�`*�[�%���x�O#��{��0D��0��4�`����>(pG�1D�|KF�F}�٠������E1D��q �V�8��ъ!`ԑ�"�"D�@C6	} �Apf�,�~�!��?D��k��A����bg��PQAv�0D�gD�&o�U�!H�fX�}���.D�x�� X8 ��6c�7�pa�'�*D���Ђ�]U��pdg�7�X1h@�*D�x�
��-	"8�a�.
�L�P&
*D��:�^�5:Tt��	�@cőS�<D�����<Q�PH��sM���p�:D��R��>{�P9�U�� MJX���f#D�S��9G�����K�&��Q�"D�(�ʂ����s ޵R>�.2D��Aq�ܶ2����%��/@L �c>D�p���^�!V �#��C X�(�o6D�Țш˦`w�CmT)!̠�!�?D����aҦg�^]x�"�;2x9��8D�Dk��P����+�l%Z�م�4D�ta�Y�f�	�S���|�A&�$D��b�4�h�Q����P_n�#`#D�,�!l�J+ڤAw��a�>�ۅ"D�`@�A��F���z��L�,���u�?D���@3No�� ��i�ҨKE�;D�<�b�N�j<�E��=P�TTՋ/D��X��J��(����GL/D���3gD&i/@��$M��6�̹�0!-D�ШŉP<u�t:�c�ew�hBC+D����KQ� ��$�R�2~f�e�T�<D���w�ݙ\�hA�X�`aG9D�$���>J������ �J!�!7D���ҧY�b�R�@�J!,�,Iy7�5D�� "y�j�-U�D��FK���h��"O���rf�� 4���3|���r"O�1E��*�]��94�*9Z�"O.D�#F�L�գP�1����"O���9#��	X�F�"r���x�"O�i&"L�O�4e�EǼu�̼3�"O2|R`�rD�k�	nΜ=��"O}X�j5QZ.,� �S�#�,D�S"O�\KWFB�isrѐ��Q����@"OV١F��m�*y�Cޅ���q@"O$X�eϏ7�01��mĻ��e�1"O�=#�f]1]�T���0>��H�"O���5�0q�p�Bcʆ�R���@"OL�P�,Ć]l��q�O�jF"OZ�"��O1W��t��#V���q�"O�B`O��OTn�ݑqO�-C&"O��rd��)���&ɧXVb�j&"Or<��ǆ5o��³��ؐz6"O=�W��1-�^@S�/�4s����"Of�p$�N0J8�ͨ6ɕ�)���)�"O2ݳ� �
aT�#��_W�|h�f"O����$ʧRi)��э^��9y "O̼ #f�F����->v��ai�"O��"�D�Yh8��N�D��"O\���Ֆ�6�#�-�
V;�"O�����T-	Y�<��,�c����D"O$D����?r��EĹV�ڭ��"OzTb 烢=D���b�͉�\Xe"OJ|��Mc-�=�v����ě�"O*����ՠr��0ɓ��Q���X�"OX��vP��-���#M�ĩ
1"O�DFO��.�p�v�?9�+`"OP�;��3d�ޠ �*�3m�v�� "O�����T�v����XP��e�"O⩋���r�u#���yX�LO!�y��Ҋ
�\���n�0�N���H��yBc!n�U���F
-�\���'�y�,��WG♃WEݨu玼h+�-�y�G�|�0����
}���׮�y�M1��	3)�sz����B��yb�L��
��¾o�Vz�K�#�yi�C�bE�S��JN��dP
�yb,���X [H�����#���yIޖ*�mF��	
���`��'=�p˰ ؓ9�fa☹�L8c�'ZL� �[���A��u�~�A�'>й���T��hBpdq��;�'f,��J,����m<��'�D@ӑ��cZ��qEۧkm.�0
�'�V�v��#68�X�/ץ,v����'8N����C�<5�!�N�,��S�'��%�SD�;J��L�C��*k���'< �  �UT�A@��0!�Hɲ�'[VBk�Uq��q��_7+9�p��'"��"��N���D���ެv�d��	�'~�c���2�Fm��ٕk[����'mp���=,�t�!����z^���'|($I6�L�Hda�a	�7|����'Ʊ���ÍP;�Y��'x���*�'Ur��w��(wn!���x�|��'��r���k��L1���t%�( 
�'�������<Nvmpd� =<����'�&ȲWEO2ӆbC	�2n0�)�'(��r��XF��x�7��).!5p��� X�H#̛=0�&%�NCvV
�;$"O@�W*�8H�8$adF�X�5!S"O���d�V HF�@'%j�UPL"D�8�HAb��S�G!}����>D����GϓN������A�om�}���;D�$;q��{'�ǥ�]�Dd�Ԃ;D�d��'4�ȩb� Z�G�&`��.D�Hrd)!@��=�S��$8�2pY�!D��A3G�WK����K�>j�FA�$D���e�ZNƖ�ZeHT�I��)
�A"D�\�U�	�ikP�ȷ��!ʝx�� D�D�tiŁE�����[0#�x� d&)D�|R�����	x�o�9X�vey�+2D��"��R�_�4QW�;NoFb�,D�p�!�B�p�����o1ʨJ!�)D��sO�� Z�(��8T,4D��:rKB��H���?I��e3c&5D�8K�/�-0��lC2yvzU��2D�0U$ ��J4�A�x�H-٧)+D�\	�oʥ\��*�-d#&)��
*D��hpÓ&.h(����� %ˡ�%D��;#J�ki�H���.���b>D�� c�9#ю|j��]
%g����8D��+E1�
h�ģܘ$a��I�6D��ɷ	�L�йqGN>F`��/3D��B2낹*�HS�Y*.���{�B1D�(��
��b���ꘒt	�� �/D�lq"��P�x@��T��9"4�.D���f�+q��xS���$����),D�t��"�0a�K�OF�a &�%D�d��	e�)J
�0!Ήj�+#D�xK݉ s$(�&	),��is� D�8;CM�bt��+)��P,ҥ)D��*SM��c8� �Fڞ%�j����'D��*5��:|�B��b���4e�b;D���f�-cH~"u��\0"��� ;D�<8��݆5�7�S2vH ��&D�(���þ4������N8�1�"D�̛���{�͛E-��7�0q��-D����N�j���z1��{$��a7���<�q��*�¬0a��P����D	B�<�0/8*���%�u��9�k�}�<���H���I�������$��|�'�?�����=����eG��pA=D����Lۼd_�]�p��W҅�,���F{���k?�$�fķ)XPJ�JW?u2�z��ĕ96JY����/+eA�
L,!�Ĕ*K/ �u�Lg������u�qO���TX���Ȗ9���X4�%�ܬ��"O�H�d�D]֖,Y��D�c'�&ЈO���F�L�Nݨ����$a�MI`d�b�<D��-[2&�ƌ��S�V���&�O��*���sӐd0�)�7bf!�&�Y�?�41�"Oʀ��d���FY&���U"O^�y��Rv��� ���0K1"O���0�N�s%���v0m�"OX��/��_s�h	��V�d��X+��~����bYS���r��qE���� >D�4�d�sZ�k7#ɢf���!=D��Y�c����-��;ܼ1�#�'D�p�U��:1��a[���q�ݹP�0D� �S�}���Wm�#�(`А,.D�����T39�̭b3P���b�j�O�C�I!U��B�A��9E:e�n[l܀B�)� �`3 F�R�0��g�ԸB�^���"O���PM\"UN�����r�iB"O�҄JJ"y�J`��UW ��b"O\CtFT6@�m��】bLPm��"O����(��jݸ��Βih2��1"O�Pv#�)��]9uM�`h��ۦ"O���1f�:U� �
zP�B"OU`BaP�<Ƙ֫��6�,�ӱ"O �c��C`��D�J�\����t"OVqa�eG~u
��#i�k�I+#"OT����28�лƨ��f�("O�mI� _'�
|cƄ$W��E"�O�%ȣA��e�8�2T,^��@C0J�<��e"Xjn�W�ڨl����)NG�<�n�>�ش
��#N��tDh�<���)B�f����8=�1��i�<�c!
$�k Ϗ	h������d�<I�e�!� t�����	�*���c�<�G%�R���A�
�_������TJ�<AiI�wH�s��_Y>�xjXC�<Y�ؠs�����h�6H�p�!�H}�<�Q΂!�l��Ag�XY�B��|�<�`&`a�e�����{vƃM�<y��֞om� ����K�$���S�<��[�w�|8ѳ��eHL!��O�<ق�ĵ
�AI'@�9js��5�p�<y�d�#VLV�1"m��2�@U����E�<ɷLX��I�����CW6A�gL|�<�� آK�n1C!#
6D��Xw��w�<�W�484�9u�ܱ-���։�n}b��>�g?)�jʕU�%aU��)@Ԏ�R7�s��8�'K���4�Ʉ^��1[M�9h_ ՠ�O���6�Of�2@�M�j�q.AR�Ÿ��	��M�����O>��ň6;$}㇪@6r�=�'8�}� ��,�$
��R�7\�'!ў"~2��,��p�-J&�H�Șg�<1��dy�fg��DF6�*��Gy2�'�V�	�������քN�D�K�')�X��N�
p�N "�m�.G0�\��'��1%��
�!h���=@D���'Kp���h�$+�֩9�@M(.��[
�'J�6�D>_ς���$!�&�p(O�MFz��iX�`ܰ5����&�LE`�ۙX1O���d��'�鱦e���.��D,(m�ĥ>I��'x�U�� o˄ᴇ�3_
U�
�'�
�V
M4�b�i�:%���	�'�؀��ߗ~���CH�ڄt�
Ó�hOxZ�Ô�'kn���EZ(�i��"O�Y�2N5��X��%,��x��)�'Vr�i�s퐿\(�t2S��$�4m�a�d!|O�Y��d�{;<��4�Z�_(YR�"O4��3��a���V�5}���+�
O�7����ı�	��m���-o1ON��-�)�S(fA�Q�B)X�.,$��FH/vf�B��at({��0x������ǟZ+bB��Y�h����F�@�Ҫ gB�++va�S:4Y���É5&���܆��E�4$;F�-C��*��	^�pC�ɩ7W �*Wm�$rjڙ$��.B�	cMҠJ ���9�+׹;�B�	,[��+�ᅢ)X�	q�-��X��C�	!@q$����q �-ř&3�C�	=W�N�SSj>l�ذK�ˀ.�tC�IA1|�A�߀ �u�Ukߝh�4c�Є�)� ��i�Ԁ,��`C!�� �f�#u�'gqO�1ZdT%!������
�ku"O�Б�㋥(:$3dC(y� q#��	~x�(��N�	�(�"e��:,��E�D�-�O$�, ����մ>ʶQ10LDx��	�ȓ{�1CĆ�(Z�P�A3�' �8E}B�SϚ����1`�ë�I��B䉍]p�E#r�]����`�*\g����d$��O�1����-�)T7�̠1��~�8xQS"O޼���Bx&u��+q���Aë��	���S�'��9O0D3#O"I��胎:��"O&�;#I�*��0��Dà"O���1��Y:0���؇Q�N`"Oƨ��.H4-�B�K��F;53P�J�'b!��*djJY�U�3K\��!B�	�
1O
"=Q���D�<Zl���V�'r�0�F���Py�BJ�X��'�;GC��r��W�'��yrgK���	�a׵o�&��uɒ��ybcH�j�J�X�D�-�J������p>��@� %���D�B�:�,�YRE�'E�O.�ODr0���I�k}1���M�|��[�'���q�A�[���SGG��n�20 ��d.�S��˙s֐U����Y(؃�Q-�y"�ʑX/�����Y�Z�������~B�)�����r1��fG�I����|؟��7k~�ȕ�4����q0:֠���4��DL �T��|�7��<t*��ȓc��|3Q�J�b5��j��/,{nՇ�Z��|����J3��8C�-4����Op�=�
�H�5��1�m�h�
��^u�<y�ե$f��Q4f�!�=�򅌹�VOj���ٮ+~<B.�z<�������i}a{���#4s���4�]���A��!򄅑4�xi��#� /܀�1�\ Yl!�d[�tR!9Ve�� "�����$1!�D_e�� �*�!*���j�!�dH �B�s7��Yp���CO!�dK1n<��*S��>@wVA�S�N"!���0	o�He��v�h㱣 �!���	3�٫�d�4u� 3�b��h�!�A:�y��C��N��L�@�Ӏ):!��$�Uc')�2dľ�	&�^�=�!�(y�!;�N̾	����U���%!���G#6��d .t�슧(H�Z!�J�1N�U��-Me�IB�G?M!�� 8�@b�X8�`�qC��!��'P��	�&G0���l̩�!��'��*TĞ��R\��/O|!�M%]µ�+�, S�ؙsʘO{!��f1�x�0�[M��xА�م`!��\�~�B��� a.�8q�Go�!��W'Xʲ�x�g��.����Ɩ C�!�E�9�0����9P��u`��5NK!�DL�7�}�lW��,t0BFT`�!�_�n�R@�Zh���֫Rj!��Z�B����+Y�&����=T�!�1y�U(��Sb�|�#��2D!�S>9�����ȓ9��ôIL��!�d~h8��-� ��9���H,8�!�E;GΩ�bC�к͋�e�"�!�D��v�� ŗ��$�²�nP!�D�uBPh%��;���h����Py�k����*p��>�Ba�A��4�y��ƽ@S☩�iT=|H"&�=�y
� �i-� D&�YH��5� `BD"O\q�Ֆ��B�C�7N��"OZ����y[*��לA��s7"O�����!yl|�.Z0�^����'��@5��'x�� ��1*���{ �G�q�z�'�:���������͊q�ج�
�'_Z��@�ǧ's����`h1A	�';�iQЪT2�02���aۺy�ʓ5��a�k3^T���F�m��aT4aR�9*�p��AkK�-����i��($ѿ1���C�K���%��q��Pah8x9l�e�R��ȓe�A�i��[�\A���0Xꬄȓ2����P*W3[�.	�$�ı�ȓ0�x|�5E�#c@�H�M���$yn�!R�C8e��1�eT�Zn]�ȓ'��8i��.�`]G/�/ ��E��w�̘��8?�֕x N�g��\��R�8a��I4t�&�rŉ��$��),��  ��NA����Ƃlf�ͅ�mݔt)��Y��%�t�Z=���ȓm\����=q�n%[rj@?^4@}�ȓ/�N��^6Y.�aF���Bi����D�$��Ĉk$�0��Ɉ�|�>���0�@+� ��`��\�d�ׯ]�-��S�5j� ��Y�=��$'+�f	�ȓr�7eMdr�x��$CdDDp�'�����Ax����t�1M
�'��RV
,p��)dL�$!q��`�'A��;!�8��	6�ԛ�\��	�'�v��D\v�f0 ��+
>-A	�'�\�yAdBSx�6�K�)���9�'Y�|�+ݿ`n ���Ұ'�6�R�'!|L��HTt��� m�d�1
�'���2|]�.��YWx%�	�'_��B`/c��q
-��R&��	�'�,�%jS�0ܔ����!B$��	�'o���FiVŲ�$ۿ.V�*
�'n������@j�$I���2���I
�'��4;(�,>�#��_�Ak�A	�'�d��K��x ��-`&0H��'F���7�I�i�VM��.j�\��
�'��))I]�T��y��Қ3r��'������a� �#E��/e8n���'�©92�--��c� �h8݊�'�����L�>V��x���
dՒ���'���{s�R",� �D�8,�f,�'k�T铤�r��*uI��
�'���R�������H7\K<ň	�'sv�1���
6� ���.JBF�@�'94�9�MҫE��jD�ݬU�|�
�'� �J�#΄GU���D#Ve�us	�'�N�;ׅ
��� 0��]��y�'��s�>K��9�g�+W:"*�'o,m���*"x5bp	��T�
%��'���q��ã��:���=K&&��	�'��`�&G�L�1�� ^�F��	�'i��k �w����%b��2 �5�	�'�|����F>n~����䘦D,���'.�T��*=���EÌ�=&�٣�'�@T9�h�s��U�R0��S�'��0`�ʻ )`9��e�5$��'�nT��n�o4��f)܍w�]��'�hu�7� ��hx[F+�5Wz84a
��� �����α�v�˯^����"O��) ��u� �I�M��F�� "OVô�ѽ},��K�Z�x�"O<� 񂔪i����"A�\�H�k�"O*ᲀA��R�>�Y��õ����"O�)8��ƥZ�"TPO%{�nqq5"Oxy�G��8E�p:�o3�����"OȬ����,�~�ӫ�:�Q�Q"O�-�ୌ� �q2�P�O�(X:�"O����H]�p'�YͮD�C"O�����y�|�K�a�����"O9k���ZS�)��@�[��t�F"O��1S��-�|L!ƀ�v�88��"OL-��J$ߜ=�N��/{����"O�0jt*Xz�Hmw,��5
r1�"Ox%:V^Y����5�j)��"O.`�6�Fqp0��"�T���@"O0��ץ��6��RBaC%#}dH��"O��;��̵hZm�f��-ZT"O��鲌̝TfQk���0�8C"O���EM4�`q���ht�w"O����#M�A�� ^&>�0��"OX-��+.6ql���%�5��H[�"O���ƪW�Ҥ�w���p�F�Bd"OB�9V�ݷu=�"0�Ogp��ɠ"O}ӐO��^�dIЀ�>Ki"�04"ObP����"G4�����WH�*�h��*,�=y���OPx��o�@;��]�3^� [w"O� �/X�
�E���:>��Q��i��c���)�|B L�`������#})�p�$�p=q���7tXk$�l��j'�	g�0��G�, �͒;=!�].�����]�-₨R��O- �qOP9�r痂��`1���D�p�b�(��.����
i��qj4�	�A2vx X�9ɦ�� &I2XA�J�ㆴ�}�O�8�M|��%�faDK�O�P�gԁi�P�"�BO�|��"O�Q���O�%M�Ӳn��R����&o��[<�"���/���:5o�l��I�����~���$]�g�D�p��2a�1WC�?�p=!�XG|�����a��9���8=h2�p���
K"��I�.�!.`��ӦS�&�N��X���?�'Clhi��� ' ���'H�uX�e��{2$A;(�&|[��[�Ol�%�r�]h������R;�3"j_#(�F)8�e�����C0<O�84��qJ@ps� .�tx��I�B��\
��>���~�d�ev�-�aB��$ d�֖ũЪD�;���9�[(`�T$��y����%��$v�9�k3\%po�w�PY�$ �;�~�Z��f���ѧ
��u��)�H���A��c�bmxG@�Q�{"lV�v ��'�<�@'P�'9(��d�9x9�C����RӞNs���ǃ0��OD�'9�s )��m~��c�ªrM�h��'�)��ʵz��x��o�1\�k�5r�x�_'�����V�E�4��I�/Iސ*dE�W�qZ��t����gP�Bt�P%m�=��k�4I��b�m�si\�.�$vm����D9$�8����'��#�a��1�U1G�5?9g�C_i�5�N�( �Nh�QD7q&���,��&݊3"ZĨ��ɟ&�\C%"OVt�	��J�ڼ:�ML�=��d�SD�I��9�d)̨f�ʨ�JL%=y�O���$����%Ƅ{#��f���RPB�e��G�);0��ɊD�Ҹ2�f�q�L#	���P�2%�|���I�ayr+]�v<1� �k����VD���On�yPD� Nض2�F�T��*�E�3x��Q��5,��a��9�,��'c�H��d�c�N��i�;��.O���N�'�<4�Z�.Z0��X���O���	Ն��ب40�Z��ܽ��'a���d�@<"���d۫h�p\�d��>H�X�S���H��ꆉF��'	J�ODQ�$֚
$�!ĬS!��T�'�Ld ^"��x���P��ؗG��/�B)�EB�D9�)9u�X�{���DV�%"�1�p��	1.� Ŏ�h��`>T
!�<�/�0�@�� �؅*s�\sWKM���49��G�V�"�+S�4)���n,$���#*#�����_L��y̂oy���:|i>b�0��h!�	�x�:�M��QE�b�� ��A�G�!+&��'��P�)[B�'��q�燿,*�����	'$�q�ǽ t���B�(O��@r!�VLt�  G�//���OD�'�6x��H�<k
��]��0���#f�`�y�5��'	���pn��%r�1���3k}T���1q�a�tVZ!���'��A����P��.�К�0(OZ���θz9T{f� ���O�)����$�D
�a�"=a��ԦT�D
(�Q���dH<�"
z���3�K>�ٻ�+��(��D��h���#L�>�v}�B
���#�>�w�����Ȉ �J�[Q� u�B�y��f���ɦp>����
e�^�{�)�1;ǡ�?YI�@pf�5}b��|��D����d�V�Ƭ���R�U�pq�#c�	�џ�:�N��O_F9�eM�q�.�Χ*?�H��JH�`|l��+�,lڄ�'6���"�W1X��yÙz�4���+�3��0��;��/1¬*P,C2t�t�� �>�S9v4�h(CO�,n�S�`N�|=�q���=!��2:�%2��.=>й�Ċǳ$<ۓᛳ"��$O�r(�0��͑"����Ο�h+���'@6()����kf��a)G�Ch$��Ü�2'hQA�M��j�X$�B/�0>Y�k��DZ�yz#�@5.�*�h�fBF��@0���5ʸ��1O����N������E�A"Ob��`�,�~Mz�&�<p_bأ��D�8-7���q���~"�A�I��y�O��d;AN@�1�LBR��$5�}��'�*<�#�PD�Ī1�O�(��<o��v����ӆ
'$�mG�A~�y ����j��`^�~�4hTj>D���᨝>\�.��BA�&��P
Q�H.�����Қ�~R��qC���n�'xh�r��主lH�X1��',֡�ch�!q�@hhD#=|q��睻?��1R��FX�L��%Ķ]�4�#�F#)A*���-<O� ��iG /K$��O.�*�1z�Bed]�ʰB!"O�1�"W�"T.�#ǡ��r�t���|�K�w�j�Q���c�O���I`f܀p5:	9��e9��	�'�>MQe�P��� 8 ��&\O� �hR�V�
�'��PQ���>qCR�0�`s�p֤�Nh<�#(�"�*9�R��#*���O����p�등-a����֠78�	��ID^>A�U.�&2�y�	|Y0]�nZ[}��I�)�F��D&��~���B��y2���[\DB@$[5P�d�"V*�'Q�t�r�V+f�?���.Y8g�-����6.��)V�8D�,+���.R���*Wm�;IF���X�yJ�xpP�<1G-��!2$�L-uLJ�藨Xn�<�A��F�1	�U�p{�ΐk�<�A�̂#_�r����
��5�g�<)�)�"6�^)�E��*E� +���d�<9�߫@�p�*R� �n'�	{�`e�<�4��_�j4�H"ya�Hj�Yb�<�Q���)ؒ�1 �
V��� l�Y�<�'���qP�D�T���=@�P|�<Y��W0�Ћg,��2�8E�ǈ�q�<��ƈ4R{��I��пRߎ�3a�`�<�`M��=�hP���7G>��(u�Xa�<I�+M�WZ�"痱yS*2R�_�<	�#�9e3�`/d|B!z6AQ�<����)�n����
�:)M�čCT�<��蛧N���{���l
]1�f]�<1�I"o��k"%�:\~�QHL@�<��2nv�q��lU�M�z�P@�f�<!f���+>�8c$�t*����d�<��Ç�/*��#s�Zj��Dc�<�7GB ?��03^�R/tM�f�Q_�<�ISy�ј�eƱv�E�"IAA�<�"]�,%(ոE�ȬdO.�@��Hk�<q���~��m{5k�6�d�HA�	`�<Aϔ�UVh��@�=H���D&�a�<�U�_3T���Ap�,�����aMb�<y6��::�=S`$ۨL�L��4Ze�<���#�갺��O�\Ԫ�᥍y�<� �������=
>��pH<zmx�"3"O>�x�"��VJ���ND�Z5����"O~�eۂl�I��� 2t�r"O�i�bf��{kL��풥l�В�"OT`#���X5�`����<�"ON�	�^k� ���=V����U"O(�	�%"y�Xm�_�p�A"O4�ɱN@��L0��͛[�<IB�"OL�a���0� �wƌ>ab9�"O��1�^�8�r4b�L��W�e�"Oh�2�/Hg��ɝ�^��P�P"O2���ӧ�8=s�Ͱ8.lT�"O4�����0�̊�b�Q�d�d"O��ˁ���(��Tz@M���3�"OV ��� �" �)��� ��P"O<術/�=g7^IR�K�Dװ��p"Ot��]�:�8��-9<�*�"O��m>6b�yR���9����e"O~x��#��"�8�B��r�z�Q'"O���E�7�x�fM8g��)U"O�X҆��'؁�D����.XZB"OF)H�=Z���U��~Cj���"OFPk���n���u��pD�Ug;D�꧃ʯvj��I5c,N_b� @4D�t���)6�X�b�,�,��0D��󵤛�1��ӵĈ#R�&��a/1D��h�dC�8����8Iol@�02D�P4�(M�a�Udƣo�R��0�0D�`�V-��N�}�K�$x��=D�0s��!t)���ȵ�(��K:D��zak��>O��@a��= ���E*D����se�qB�F�>g�-�@+D��c����).�dX�$Ům
c(D��#J�	6pɷN��jXd�c�%D�@S�׭]�,�+	�>`W@q#�>D���W/( a �?�N	�&D�l���ѷd�TX�aW��� �A*'D�lA�DʷQNh��U�m���"%D���`�Yr��s�P�}�|�(5D��p��Re�јªU�]�l��3D��0͚�y=�ČR��\dp(<D�Ps@o�99��d��K�TK>T���6D����
�&Δ;���Y���ȱb4D��1�:nv��p�A�;><�H9D�*�K��d�@�:���Y�^�A0D�0:� $:P|�D�\.��a�#D�<j�x3��HC״����Ư>D�4a��*C�Ұ�0W�	�ҹq�K?D����g$�(�cb�=j�5(�?D���E��e{������:���rT@1D��c���z���@��qA�	,D���Vd@�Zŉ׌fJ��379D��P��;���"�eJ��v�8�/7D�Т5�*iй���y\�53D�\�πg����c���>3�3D��{Gi�z��K��<}Fɋ�:D�\� d���GC�P49�Ǝ8D�P�@�X�qIZ	kJ��A�7D��Q�%������R`�JD>1%�5D�@�bjߩzv�p�dC�i9
����/D�@���۴fW`=��"
�Z���&D�,��,Z,6�h��@ަ72�$�8D�l�A胴eP�㱋�z( e@��;D�C���
J�,HBÅ�+e�X�A�O#D�� F��듽v�0��Ȕ&`d"OnMaԨ�0Z@j�PA��0�x�e"OHaP��13w|�
�J�&�p4��"O�bQ��V�c���8h��`"O��0e��0��m]&vl�"OX,�A/��)�y �jC.Yg�8��"O�)�/��Ң�Ӈ!Lt`z�"O\}:«̪"��)�$Ö��>�Ї"O�`��A�?�M��eL�h3��3"O����YmL�01G�-�cv"O�H�M'�f���w���җ"O$d���P8#�t�Ă
�Q8 "O&��.�
=ߨ%S�N=�p0A�"O�q�Ƭ9�*DC#l�p�&���"O�M�� �R���eғ4�t[�"O��J�G��t#�	ஓ< ��(E"OԐ�s��{��YómĈ1�N���"O��K��s�����@�O�&�Q�"OR�Sse�R}|]�P��N�"���"O@��G��>.�>�h�̆�� Tz�"O���o�e�pջ��(>댬Q "O����B�'� +S�+Ɉ�J�"O�����p��3���f�d%�'"O(m`�����*�&թM}���"OR����rP�!�H�
y�ݒ�"O�]rd(D�%�� @�\��X�"O>��ol���qò�pqB$"O�@!���"�2GH9��,y@"O� k�@�&��uMR%0��e�"O���"ט��8s��miʴB�"O(�A�IL�7FXI �F,�p����e��`�=ي��O*E	���/_�@x��8Z�HX��"O�`�`T*v��4͕!����i��b�NA���|���+X���a`m�k���㵋�p=&@Z;u�v�
��s���s/S��n`��G%lӺ�ӢI/D���䟜- 8`S�B]1F�*��

��0���L�"�?=�A�9B���U���4�1�(D���aᖐ:�t)A̓a"E�H*v!��7}��Q����		G�LRF�;Y2=b�ǘmJ!��9�ܲ��?D��aT��$R#��{�����k�'�,�C曩y�dwa�:Z�Z	�1��uxt��R�ɿ(�D����{�U(�R6\>�I�����S���_���9�T�pډ�$��05�\��h�P��%�"t�:`X�����ط�N���.Թ������<��6��t ��[�8�v	��:NTP�mG�$���OBFʒ.���W�;��R��b@�v��mH<QB��&J���rd
�_a�u$Ŧ1�� Z�H�'�!"I�#.F�>�';�J��5�˸>�R@�'��8�X��I%|p��_�$��K�]r�� R���q�x��ò�����$?�
׫�o�4�?�'�d�{�B��|�!@ɆL��+�'�����>*����@�*�i�ߙ"։���B�#�,`$I��<yF��U:T�`�A�(M(�1SEx8��@�BI�Rp� ��g���)5c�7h8�١�N�-i:���&ԭ8��q�ēh7��PtfW�j� �Y�A�:5�'	d�8�ʌ�!��ezR-�������@6�-\M
��4jK�$6Tp7��;V�C䉄��(�
��
|�q��m��`��i�	Q��`��c�Dɸ)*�I��ēe��XE��G)��%� AS45��ɓg��p�����`�*U�DoG�@?��)g��$_6h[�ҕO�bDs4cp�ayR-�?lb�5 �o��HMzM��ԓ��O���v ���:�e%�PEjd+U"��:�	�,fx�D���-9
�'��U�ȉ4@*���#I�^`8�B-O���(��"n��tK�x�"�͐���O�����$ڻ!�J|��$\�F���'Y��я
�Q�Ӳ�[�\�����Y8��� aN�.���`���',��O}�� J,!���1�^���i���'>e�� 0���#¨v�a�fbS)D�]�%C�,<*�B`�&n#<�aD><O�u&ͮA�9@#�PH����>y�T#/���3k|��(��S���JbG\.�R�C�ַ ~�!hF�UR
m����q�lC��;r��QR0�Ny P���ǘi߄��'4��hՂ@g�m�N�(a� ��~ݡ�G�٦���4*�;�N�P���
#��b�ҁA�R�$�j�и*x��3'ֶR�t@ӵ�R���" �:tha;�	�4\j�G�x���x�?MI�m9�jЕ(T�4���	���O05�7���D_�@K|�P��4fs���ui�^�<=b�@y��l�dţ�(�`X�\B6b�S~�r�(�V��P��<��*١jdB�RC��O���>�!T�_�M�R��%b�K�\�ViQgti����] !�B����82G�.{��9�gC���  ����yB�]�}:��	`.°���xR�Kn��|�1�ލVc ���P�Cs$�&�'�O~$:�)�=GҰ����A�
�9�_:gf��s���.���,@��U2P��aHA�t��E7F�/9ᠨa䇝CDХE2�\}����f�|	a�6��(�Z-6$�����f4�p��L�E�2�l���!5��@�J����1�M�=q�˓Up@0�/G-5����ר���Oz��+�f��f���µ
�]6uA����<�ȓd�S��Q�}5�	�gO�*i6���&L3p���􌸺6�J@�g̓��`��
C����գ���!�Rv�@8�n	�gJ�XsO�<'�bQ�'˃�R�(� E	6����$,pڍ��H30���DE��z�$q�y�!��<!ucLV�6U�rj��@`�M���G�<�ǅN�	�.݃�A!��!��Aܓ`B��#��,v��8R�r�?u�b"�g��x�N�_��	�$%%D�tAB�U)����3`�ܱ���B�&�V�r�O�	��.�<��|BQ1���+�*�~�4���BV�� mH�"O��)
�mM22S��&y���/>m����d�`?� d����4�(�D�0P!n�ky耂��4��+��ܚ2'O%E�%�B�шu0��k��ȯ,y�tbT <�O�y��`׆t~���q�ї^fL����'|�퉱DД[aF��'SP}�d�/�TI�(~mK�'B֙�A�L�B͊�oV����3J>���ֳ���r$=�����eN��ۈ�b0�(%<C䉳g"x��!�u��m	TO<�	�b����	�z9��OI��\�"̸-��L�E��9�OK����<�r%�t��yӄR�G�0�b�3ɜ��� �sԁ	�"ɟ��ą�I�r؝1�≞��	��$�fL�!	�E�&��#��C�"6�@Q!q��<'N���GKI��Fb����	�B,F���ɍr��97j��5������5�y"��5L	�6�Y�'V
y!��3[��Uˌ{�m���ګ�E{r ݣ7)�9@$)ʫ�!��V_��'D�%X��+@�!�D��0�	X�-]"&f&�;ЀW�6�!�D ?o�A	p"���ʠc�K&_�!�P�(�81��ؿdM�ӱ�T���ȓRƄH�	�x��(8�eN�;T,ԅ�a=���C�a��#r�]
�Jy�ȓr��V��L��k�S��� �ȓVRΨ��Κ�`
�8�	��G��U�ȓn���e��8r��@��3����H0�X�r�+F>��i	0O����1��+�n-L���df��j�b,��hp��6�xx�Y	ԟn�� ��Ak �a�,S?�< '&J�c^���%�~u�"N�()&��J �D�&�ȓ,�h�Y=e:���m�0b+.a�ȓ�&�cϓ�3PI�],g��l��l��uK!�
l�^��i�+�b��m��
��Q�3%zM@#�Q8A^لȓd� y�e$/f�d���`N�H�$��ȓH>ʼ��ˬ.@B��եLHDF���!�|���G�6U�lO�8M��8�D|��#�V�x��>3"|ه�S�? ���2��LA!7A�6f��"O��S�
�5����p��	�����"O�-�g�:z���6�$a�d[q"OK��.eT�#G��=}��3EC"�y�+��j�P@M^9Z�9�bƐ�y�ע�y���Y�_���PbNR.�yr�V&���a�C�T��0��(���y(�
�&�����V�8m��GP��yR+[<�L�E�I2xtB" T��yr�Ȯn-�����S�MO�8P�#'�y�+O�s�xA��%�T#���!��yR%E&�x]�rcA�@�Xt;�D��0?1�!�!-&,�P�L�3�<1��+(�d��Ù^�<���^V�����ѱ~�����Z�<�b��G/]�cJ�(X3�I]X�<��Y�6�J"@O#o�-�f���<�Q�]�Y�$�ul��3���<��ȮO��D��ǻ#W0S���~�<yF��=�8���-��4{��o�<)���(�N���e�Y�<5���@�<�c�ІGL��4/�/.DMP5��f�<)g��=Y�@���P�V<s�Ag�<�#.�97�+��ǳ>ː�$y�<aUM&n��)BE��x0�M�7�|�<���!ef��Z���_v~�%`��%�M#V+
���	��uw�7����-0�CҨ��8c2e��B��~��^F�~��	Kw�퓓<�� ��F�~A")|38�c�H2.N8i��7}���_*2��7gR����Tm�?%������
zr���0|2T$܊XB굱&�K�c��h`�J��CD���O(���Պ�&����iS�@�ZE�҂�94DZ��'�\�O�%���qfLM����&H���*OF|�B�F���a' � V8X�X�'b�}*�K4u\�����F��� 	�'�jm !��,��@�Ԉ?�R��'��P��	j���8�� &t� �'&�8+�Xl�԰��5i��(�'�:��wc�<GB�����.��Q�'w�!iQ�˂*�D�B� �~Ġ
�'��pBǙ\,(z�������N��{����%������.3��ȓ�f}��ӳ!w��õ�"ݺ܄ȓB����^&L�<!U�ު��1��_vl����=A�Fl�*_�� ��x�F�2���%j���u <Y�h�ȓ �4�n�6+�`h�S��/ͅ�"z��$@Yd�Bt ��3:����9�2XʂʭP���j��D�x�����~X%'E!A�Vb!���:�q�ȓPCH���X�2d t#ė,"���ȓb>���NԪ_{�0p`��r7�4�ȓ]���r��B&r��}J�/¸;='\��D�/����ȌZ�f	8�	PQ!򄗄3jd��֪H~�Iȇ���!�÷d��e𦭞#wx���AZ�!�D4����&XU�ĊQ�Қ7Y!�d�X�ۥ�B�W��pq�ƘCO!��X�"�H�z� +�͚p�!��*Z���a���,�9�r#�15�!�$�1jQ���I� G@��`	��y�!�$�����'d�c�H��	=�!��'@��Y���ɯl�x�Wg8`�!�$dJ34K��}�^�'�bi!��`-��M�7Akؙq�ȍ�_T!�d=��ъ7���9�r�^�]8!�� ȐY��6IJ�(G�ÿ*�����"O�����$w�qA���2�D�"Od<B���}�Za��ƥ1r|$��"OL((J4������Uʰڰ"O���Ke40�٠d��Z���j�"O��$D�4>���dD`Ty�"O�h�U��)P��4{с?���3�"O�tUfJ�kM��Y���23."O�|9D�;8Q�b߆e#��"O"ٴ�3�4j`L�"�$"OR�V�Cұ�*���pKd"O}{ (ZV-��c7iE�)�D��"OP�K�EUPt\Ec��[��q"OxŃ�M=gV�,{�eM�5�L�[�"O��I��)6Nm��eЁ>�)(0"O�a�X& E\�`�ق0xk�"O<&��_m:|���ԋJ���"O@�v��.`"��TM���
��b"O�i��c9�6 Y�Р�!��(_�l�3��1Ҩ�cΚ��!�:*l����M�N��r,��YO!��I��~,���LD���H��͝HL!�dCq2`z��#v0�j��!�$S�~*�5j���jZ��t��\�!�Ĉ8ܐ4��G�&cE�i6)Q!��Q�~8T	�e��k^�Z���9I!���p� dq#�D� �E�Bq�'�8��ف�d2�lǄ7h�x�'��y�eC9#�d#��@�,�+�'p���ÿg��1�G�ƾ8 ��'���6C�v!�`�N�\*X8r�'�r�3�'��h٫��ٳO|�l�'��P���hm�\(�$^�NG�}c�',���3OA��{q@MR*�b�'e,�U��@�	�
B�.�{	�'J~Ha�a�c��Ɋ�
>$��B�'B�;��*	�E�R��%D�Lk�'� �[�$^.qD}�¬��B����'tV��+E&;��1ڡ�WLH�0x�'�f)r6�^��`kV6���
�'xB���B�d�xu�2'ߌ�����'���:��Y���%$�p�S�'�ʵ����^)���v�V/)�9�'�`�b�O��4�u�Ɯ���H�'3*��[�<��t����A��'�V�a�`�)T�K1"
<�'�`�BA�5{�~��B��t�q�'	�m;��A>@y�у��m$�b�'��(%��9���&�/lg0�
�'F@�U��l%섢7���v�p)�'����u,*��A?��p �'��b�PJ:0�YQ�S�<+��
�'l�p�x{��S���7�B���''d�
�C�Z��K�`|��''��8p)A�Nv�+`㞣+��|P
�'�.y��.("n�I�g5(��H�	�'��]��ț-�\��S�#���K	�'V2�0�%��	��Z�F=!�8�#�'I�,ر烣}ښ��с����\��'p*RlY2F�������L�2`��'vj�r�V	!Ϭ�yUA�*=Ƭ��
�'ZݱR闑*B�h����<e�`�'{6�R�r�X����!H�|�	�''Jly���hzT�4 M�BY�	��� LMc(Z�X���s Ịk�� "O�-��4;���S꘳j��P��"OĜ�ƃ������:���i�"O�h��)�IrHM��Ň<�$�"O�`����0� Qz&D�-�n�F"Ot���n�4U�w�$(n����"O��;gɤj�x#geA=YE&��"O<��b��6x�L2�C��Ө���"OR�i�H��(LXc�(/l�`$��"O*��b��k.�Ag��J3:|S�"O^�` J?�	��+��%�$"Oh���Dr5����V�x�#B"O"E��	v�j$��c�h$��"O���
#�XC���O��d�"O\x���,m˲ ��y��"O0䂂�T�Т��/
HH�0"O$,R�h��8~<�*fk��<Q�hW"O�!!`MR0~rF��%���"@(�"O ���bئjwv�������b"O.IѷoZ���3��,7�ft�7"O$�Y�d�/$9։:���f��1U"O��`�Z��������(�"O
,x�y�x�j��23�"OY[���=<S>��Bq��}�"OtL���^�r�H���/uZ��'"O�$���KJl9P�_b��`"O��a�C8ː�3��S8#PN}C"OZ$ �I3@�ڕq�N��cW���"O$9����1�`�@$	7F԰�"O6Q�rfs�ְj�S#Id%�"O5�.('��a0���Bp9�"ONU2⡍�V
t+'!;��9�"OA@F�ψ:��ҕ�ӘTtI�"O|+���$T���1�#w���T"O�)��Y�P>x#Ў]�I �P"O"����R��Y(BR"�m!�"OX	�1N�:N��($[Ppw"O��yd�@��t�"C�i��ЁQ"OP���;|�>i���0y�ШT"OB����!Wj��Q�܀L�ꜙ�*O��ď9~�T�{'V�fI@T��'#�e	B��$X�� !/� EK�'\�����#������)�Ȝ��'�
�[�i?I'HUz��N�|����'�&���K
7l��@�ǇM{�� h�'h^��Ӣ0�^S�GǶy�@��'/R=�%+
_<��sF���b�p�'���#@�s<��Y����E��	�'G�\{vdI 180�բ�@�H1C�'Q����X�YyF �4�� �'b���-�5m�6c�eܩ	r�i�'u�I�ص	+^�Q7�^�g����'\�x��g� J��X���]��,S�'Y�@CfѶMK&�	|�92�'����\�|�t�4lU���'0\�Ǧ����14���,���'r����D@�u:Cɛ�?!�h�'tlɒhU[�z\�R�̜O\F���'��R����Tg'{�&���"D�$ia��P�rA���I��ܑ��2D�����T����9Wn,�f	�Y�C�In.�=�磑��h L��C�	.G�:�u�e�F0˗I�3�JB��#��B��A5`I2�#sC�+L�C�)� Z�hTbO�vY�)��ˉ=��r"O´�G�R�6|С��_X���"O�\�"�	NP���N�C縕)E"O�T�S��;L5�Z�-9(/���"O8�� �W�rMSS��1yZh�"O�\ف�$B���􄐠w��b"O$�ᇆ�s��� ��x-�A�"O:��w�v��ЄB��P�"O�����|9(���G�0�	�"O�*2���������5.�y"�"O �a��G2И�M
�,lh�"O�P+�!�Cɀ5�M5|��D"O���Qi�����rz��"Oz�9�EÂU�V�K�!̐d��"O����
��hK4!H���2"O���f���q���+��)J��h"�"O(�ɔg��/��Xw�ҡm%h5��"O&)����%k�J��!BԺ!�!0"O�|S��I�u�T���7�z%��"O�+!\�M�iPLҦ:��i�"OR"Ƌ�;.N�P�J5GRXH�"O\UǏT!�	��� I����"O~|�G͍Aƒ0	�'�2C��"O@��^�y/��peW�h;���"O	*tÒ
�$=�p�Hz0z�"O�p��ؠDx�"C"/*�H�"O�\�!��;A��A�K�2L"OD1d�P);�tiP��T�%��IA`"OJl��&�	R�*	*�]+�V< �"OD�p4n�'R�Jq�P�r�ЙJ�"O�������܊ mR%I}��9�"O�<���<H�����ܸfy\$( "O&�S&V%e@��9���!` U��"O�I�����V�B�@CF���"O�0y�&Ogj��#�\$���e"O����-L#`=�{�A&\��"ObHH�� n�i����;�L,��"O���$��sk|ᩖ�ƫ?^�9JD"O`PtO��|'4;�� =cAiu"O��qT'/no��:��(@B� �"O�{#��:��-@��tXf�r'"OA(�   ��   �  >  �  �  8*  �5  $A  �L  X  �c  
o  z  s�  �  8�  #�  l�  ĥ  
�  J�  ��  �  ��  ��  F�  ��  J�  ��  ��  �  `�  ��  � - � � �# q* C3 �: �A �G N R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr�'��'���'�*��@
X�a}�(��MJ��j�Y��'��'�"�')��'k��'�B�'�@i��
�-���Kd�@~�@l�6�'���'���'�2�'��'���'�\��Ǟ3tK��ШV��i��'!��'�"�'k��']��'�b�'a��K2G�3e$���+�d� �c�';��'���'��'R��'��':�x�l`�.=��W�L�p���'�R�';b�'mb�'�b�'��'�R��tOF
z	��
���i��'�B�'U��'���'?��'�B�'�H����ܠ4V�}���
t�>�RW�'���'���'M��'b�'���'��Z��Q bVb���Ȍ�qn�[��'h�'uB�'y��'���'{B�'f��ZE�[�m��12Uf�g`A���'+��'~R�'o��'�2�'j"�'%S��?c�\RtIץp��q
2�'��'�R�'t�'��'���'
��:c�Rє��ɖ1F8aY��'.��'C2�'���'���'L2�' $X����7M�8�cûΜ�0�' �'K"�'�R�'��HcӮ�D�O���!j��EGV$�b�*T!���,F~y��'��)�3?��i��$
�.66�ҍJ��/w#8M��e:����䦉�?��<��:��Q�G 5/����9#�^�����?����M��O�����K?Aj�N"a�PYp����P3��K��1��埬�'��>IS5�>/� ���<3�<)�'%�M�`̓��O!�6=�tip��.�1����t��装M�Oh��~��֧�O�q�d�i��Q�?���z����H:�D�{��Dk��3��J�=ͧ�?�v�Z�8����k�4��q��)U�<�+Oz�Ol�oZ	,�c��r�eW�4�r0�3��[,6��q�Pm�:�I֟0���<��O�p�T/�0Wa�l�%�*|��t����x�I�D�4�`�.�S���'7��	��4(�udV�y2_WZ(�@_�4�'[��9O��õ�N�b��9��4;H8��c0O`�nZv��0���4��բD��!s�	��ъ	^J�%0O��d�O0��OG�73?��O�@��9E�n=BG	����@i(i.�hYL>����?ͧ�?)���?����?�2)
�S7�+�`R��"�Z�i�%���.6BP��k�h���O��oz>��>6��p���_�M`D��3xTx�	�����I4�Mk��i7m� y 4�'�B��yϺ|P�SWp�5k��I�L���,J�K�T%A��S;�p�to_ 9ʺ�\wI^O ��'�:�3D�.	�:��o �����'g2�'�����U�@��4]�D��V��9����V����� �;�0h�@��dE~y��'��j�LL�"n@�v�e��N=%��]��Q�;�>6M!?�w:P�������'��{�F��Vqɤ�ϸ��YQ5��<���?����?����?��T&��=���0⮟�]��L0�f�7Yg��'��eӄ��4;������%'�PB4o����c��U�j
!�n�%�ēԛ��g��IA�3�7:?��(͖R����"��Y���K�i�`��|ɕ��O��O>�-O����O����O��q�摿����7�Hz� E#{"�'��ɒ�M5O��D�O�'B3SB��LI94C6X��'�b�R7�&�o�Ȝ$��
���9T�/FS 13��_�P��`ɚ2i:$�4E ��4�����4ΒO)Ū�6]�`2�#ίd���sB��OP�D�O���O1��ʓe����8�=��e�b;X� �(�&?��ɀ��']��t���`-O�7��$$���8t�>͂Ԫ���l��M�e�^*�M��O(�C��Ը����<y�=4����bJ�)
�����S�<Q+O*��O"�d�O����O�ʧ(/�,A�n
�a�T�.G�o�Pt��i`�|��'�2�'R�O�Bgu��ȉ|��a�̇]}���
�lڨ�M��x����^.%u�v?O�p�Uf�>	�4� 昘5��$=O>�C�ΐ��?q�O"���<���?���1�hzR(ϊ2xZ�kݲ�?����?�������ߦ5�PCELy��'����hReSn�CC�;O��`Rv�|��'��v��6�f�p`$��{a�۝x<��wk��"�0��+?酯�o=������'a>��d��?Q�A��+W����p6���Ȃ��?���?	��?Q����Od)��ۭ^��ȃ�M<1֌B��O8�oZ�P5���џd�4���yG���B���m�*{;ZA����yb�x��inZ��M[��M��Oz�R&����_w���{�R:�M�6O���y��=�Ļ<a��?!���?����?Yf@ႁ�T���R����U� <Y/O�Qo�hk>��'����'.P�¤�.�
Dp0�N,Lg�����>9���?)K>�|j���ki6#�Z�
4�Ӧ!G�ZN��&����1�F1���M|ƒOB˓|h��b%�Y8���E��
趥����?i��?Q��|�+O��n�$>�P��I�k=�"��ҡLY0qb8��ǀ�O<9nZR�����*�M��iV�7M��:�S�
�g��`Z�c����E�k�x�s�
�K��� �H~
�{�? �=`sl�z�v��  �n<�dЃ4Ot���Or���O����O�?�҄��3���C�ޘ%N�)���0�����(�4�O\�7�$��ԡ2��)	�����˧~J�Ot���O�I�U��6-2?��ĩ��BΙtM�h���3��1f�:�?��!�ľ<q��Ϡv��L�kςAW�@�4�O��l/(��	�	�h��A�$Hϯ �2̠�E�26F��fBL1����I}b�'��|ʟ�i1t͉9_w4=ZF N���!�m�n��e�F�ã`xr��|Z���O��K>Yt�U&3N�� �/A%� ��n<i��i�.p�r�D���cq�X=XR��ǲ/S�'��7m'������O�� `G 6�V�i`-Ʉx+��Or���Ԋ�ش����l��F�|$S(O���$�C�)��'-ڋmݺ)09O<���=ie��h���� �WA,x��ԝuț��q��'Q����Φ�9C�xD�4)�.;��5'�L��:ܴX��F�+��)t!�6mb�H�P��Gt�A3!I+њKE�l�@y䎝��B��b�sy��'ar��g��h��O�9 eJ}���̂B���'�b�'k�	��M��lY�?y��?q��*T���ُmހ"�L��'o��j�&K�O�O� QaR	���siU<O� \
s��(�s�%'����fE�ӣ%�fAן�r��ǐ#7,�Krd�l�I������	��IɟPF�D�'�L���[�0ؑU�X	{��
��'6|6�#���$�Opl�O�Ӽ#�DY�n��	Jv+�d(^�/x}ϓ~����vӖ�lZj�oZk~�LEw!D��ӳh9�b��K�V�2S@ҼmT��7�|P��Iޟ��ǟ\�Iן|lD�u�UZ�� )���wy2�d�d�.�O����O �?���_��]�!ږX��yr�����O6��JP�)�Ӽ,&Y�KG)}w<0فc/�HAj��K���?^ԑ
�
�Ot!M>!,Op鹦J��7X!��
#�����O��O��D�O�<�!�'������8B>�R��C��0էܹF9�Q̓VE���ĀS}�'-�ghӀ�X�VA�.,��σ�D���@.PN87m=?G`	9*!���1�S��)��Í2
��PRjX"/��R��w�,��⟬��柠�	����j���|S�U��)n�XmC�	4�?���?�t�'��Dk/O��o�f�y���23.��bd��A�[��y�O<��i�6=��	�rcaӜ�
�}qq��#!]�����R��<����eb��ѥ����4���D�O��d�.V�p�ڗ@�~ĺ-�!��������O��mě6cҾnh�	��|�O���!֢���$L�|�0�@�'&"��>����?!I>�O�ְ�o̚n�!u Kr��*�j�-^���9ׄPlO�i>����'G�$��A�/(>��7�X�)�cER�����ş�����b>��'��6M>�<,��7�.l���Ԫ��i���<��i��O6l�'��6!�
J7�r�I�W��Ӧ��t�6�Gæ�]̦��'<�s��?����I A�%G�1P���,��P4O���?A���?)��?�����I�,X[,���-�$Nz)䋓�/.X���2T�����O ��=�9On�lz�=��M�H䅀m��z\Xu�����@�I���Ş�8�k�4�y��	Gs\3sL�A�N�S�f��y�U'3�0��	>Uj�'��i>�IEJ��R
�<���!N��6P�	ܟ�����'6:�d��<�"�'X��˃v0�����U74�X�Bj�$.�O`�'���'�O��Y�
 A?$٠7����)V��D��j�I�i�,+�S	NR,�ݟxrq떥A5����KYz����I�p��� ����PG��w�İ	s�A�Nq�2��'l�̝c�'��6-�)HQ��i��4���)��>�v��`]�X9�;O����O��d C��7M,?��M]�P��gP��rG$m;���P�3W���*<��<���?���?����?9��hz����@.�4�#�D��Ă��9 ���ޟ��IΟl%?牺w���{��;(�,�W�Gr�!�O�d�OޒO1�f �@�����cSA�q�d�[��)8>�'̣<�q.�~���䟰����d�g=zYbC��#�,��d#�"˸�d�O2�$�O��4��˓(�e�-ەOg�2V'�x�$�zqj�2�y��⟬�O�Ml�!�M���i��\��R�8"���W-<�<Y@�k�*��֐���	",��$�)��֕󆊨v*��رN�:Oy��r3O��$�O��$�OV���Or�?%R��\� �J5LޡbթE�����I� �۴&־�'�?1��i��'�v,F�Ю;l��);*D���M'�$�OF7=�f�tDg�X�i;��2n�;F�ඁ�Kh���F�"�h�Ā�����4���D�O �D�?h�le�!J��3�ư_����O��8��V�Ӣ{��'�2S>�3�b[X�R���#�)h{$9�bC??	�Y���	ӟ�M<�O��Ā0��h�bAX�k�?��Z����l�/և��4������z�ON0�����p˂�+�ʈk|!�ƃ�O��D�O����O1��ʓ0��蛯D@L��ʂ�7HD8��֦�x�C�Q��Kٴ��'DDꓔ?�4c��":1��Y3x����E��?i��ix� +�i=���ǘ%J��O��g�? �a!O�A�����{�@�&>O�ʓ�?a��?���?����:�P0eC�0�B�YS[��T�n!R��|�	ȟT��Y�s�������BO�FtF'�9�d�15�޲�?i����S�';�.=�ܴ�y2�з�<A���m�X�C �yR�M��d��
1M�'�	ӟ`���`����Ƅ8��J8/NB���ʟ���'l���(1R�'k"�^/�xTZV�$�TW�	�:��?�Q���Iş�&����Q���ȓx����1?�IH�53���i<��'>1��$��?�m�0�Z��҃�^
�� c;�?)���?���?)��9煮� * ���,ۧ�ݕx"V[��O�hmZ�q����'�X7�(�i�I�S�T,#����b��#Ev<�3n����џ ��)!`�l�v~Zwvl�C�O�N�ᄥG<�Zl��A�P��n�L�Ry2�'���'s�'
�FҴ;>���V3P$ ����!eH�"�M#E���?i���?qN~b�]�B��f��\T2 ��p���X���4C ��A3���rުH8��K�"��q�c�.�a����*�	l�Y�Fd�ON �J>�.O��b���P�@��X�N��.�O�$�O���O�<!��i�*Q
G�'s�)�7Ƀ4^2�j6õYr��&�'4*6�*��'��$�O�7�������l��x��X�(��ʲ�Z�	��1m�K~+K�k�z��%)�O��F�(!����`G�e��$A3 T	�y��'-2�'%B�'����jب<�/�5ky���%n�n��O��$�� �r>E����MsN>13ER0?�v�!���%j�c�F 2Q�'$r���t��&����� X�d�x���JC�+��`6F-9e��J�h��my2�'w��'�	�`]�Q�DfV3ۮ���)K���'_�ɷ�M;��$�'�RY>�6���I��g5k>(��/1?��Q����ԟH$��&��A��:D�����9�IyB�l@�UPB��'��4��	��.�:�Od��ψ�o	z}s`��  �q�C�O����O ���O1�`�zO����eR��x3Q�F��`�g��J�(-Q�'�B�h�4�<j�O��~�X�ń�)Aڨ bt�^�i@��ͦ�YA��ڦm�'�h�c�T�?���q5�ח/.)i��CSɒغ"5Ox˓�?Y���?����?�������5{J`��D/�,S*�r �£�dnA�����d�	F��_���w:�<#7�)e�=����&HP`���'�r�|��jfD��6OL]S��N(d@ L��`NM�|գ�0O섒�@�?��>���<���?��%��qT!�4�\�4r�����$�?���?�����Ʀ�:��]ܟ\��Οt� �!���%�<O#�-�Og�P���П�n�<��Tڽ���_.ͬ��$$�3%`��'X�1�!³o8�z"��@��z��'�,x0lκ.��}� �b�X{�'���'*��'��>!�	�t6�U�ٳ;T%�5��r�б�I��M�@�ʪ�?���E6�V�4�6����R�r�j�Ҳ��.J�E�E=O�oZ��M����E'��M��O��R�Ę�����M&$5��M�gh�تa�ɷ."h�O�ʓ�?A��?���?y�!Ƣ`霓><�e�qMӏvGX�:+Ov�mڣ!�|���؟���^�؟̛���r`������*�6�z�����Ʀ�ڴW-���O��)�c�"v� ��%��2\*�w)�O��5.���C%\����D�X�O˓s�ℙ�돸��1k�N����L���?��?!��|�+O�n�H$����]����2�@?xϠ\wbʔ,�����M��ϫ>����?���a�0�BU(�4^*r(�Alڍ^����P��?�Ms�O~m���ګ�!�>�	��~$j_
t�
�ٰB�r@�0�;O����O��O�$�Or�?Up�i1�^���Ĵ
���5Zğ�Iߟ`��4�H�s�l�ߴ�������V4�8��sdP�q\ڠ*H>����?�'j60i�4����t���<wW>8�b@�Y3 M�a�ٟ)-$���������OD���O��$
�ϊQV��5�����7V����O,˓$����gWB�'q�P>�S�g�?w�J�M�X�����@.?� ^���4a��f/#�?�Bw��FzM��
ʳ8���D�/t��X��Rm�X��|����OX�pN>�Gn͇�ȱt�T�'"�=�F���?���?����?�|2+Ov�nڀk�ɱB>rO���Q�֯Ae|��%Kџ����M�R�>Y2�i���N�5Bl��`N(a�T���`�z�mZ�L�R(m�o~��ί5Dp�)a��	�Zd�$k&m�u��A�G`�z�	syb�'G"�'���'m"T>�Ed[5F��X�C�T��������M+��Ȝ�?����?q��D�v���tL�eyWBͬЈ��ҿ5k��$�O��&�b>�r�e���]��H�@ȃ
{����	bb`�;0<�G�OƐ(N>	(O�	�O�%c�/��qo�1� ٬<>���m�O��O��<i��i8>Q��'�r�'R|#�+�6+�d�����������zy�'��ƃ>��V E����/ɍ<�P @� ��#��I��(�h���B��'?�p��'G���I�]���d�M.����܌a��Ο�����It��y�Lx6`�a�-c�PɈ��ȻO����b!�w��O���L���?ͻ�$���]�b�D�C�
�ވ�~��VJc�$Yo���L�nZ]~b��t������� ~��s�?tFV!��2U�� �>���<����?q��?����?��H	�u`����?[/`2��P��d�����5$qyr�'R�O��S2��wЀA�6]:�M�yj��3��vLsӾ%�b>Z�k����+A	W!"�0�C	L�H�e��lyrg�0�$u�I�[��'��IJ3~�b�����T����$3$x������ß��i>A�'Ib6�Q�?�$��2p�6� L-ņ
����SҦ1�?�!T�(��ʦ)��4|�Ԑ�åͨ`u]!�����Z #H����;?)!�-v���I,�S��E ���15�$dyC.�< &��-i���ܟD�	ڟ��I�������J2z�t�j�!b^ĚQ`Ƨ�?	��?I�i�Π�dQ�dR�4������S���Aק,}hTi�x��oӴ�mz>Ya����=�'+>�(�}�2WY�t�Pa���)��<�7�'g<�&�(�����'�2�'�`�7���ڶ���ІvdxT0s�'*�_�����iZ��������Y�D-�N��uc�L�x�V�C�nȔ��LX}��'tB�8�?!x���F>��u�$n6��j�	˂*�����_���|�A��O.	�L>��% ��1�Q��D�������?����?i���?�|�-O4�mڐz`ȩ���&aE����sAn�!"Fܟd����M�ҍ�>��7���u5vf��EHX�;Fs�X6��+����̲���:��Ԝ~J&�=P�<���/Hv0���<)-O���O���O���Oʧ)&�<�)��d��@�GZK�����i��I���'���'T��y�`��nֶuy&�ذ�	�hLhb4���9�&io�,�M+��x���c�T���>O`� Ǥբt�ziiS�(��8O\-�ŏ�?���.�$�<�'�?�a�$4�â��S������?����?�����֦%�U �柌�	��am��[�n�ʂ�<��lr���o���˟t�������XB��8����n��%\H`�'sE�͇n�� ���EƟ� ��'�.��1�F��@S��T��M��'��'�b�'��>睷+Jp��sj�܄�$+vi�Omm�
g=�|�	��ڴ���y�K��RI
<FH_�Ș#�@��y��'��'Uv�Ѿi��i��"T��?*�e�e����G���8Zy
4L�0=�':��ğL���(�I����Ii�29��̕&u�HE�&j�޼�'�H7͑dl4���O��3���Q���(d+ݞA�v�N$xǰTC�O�n��M�$�x��Dl��@v�L��#F,��x)��^�� �4Z�t�C�L4zB�z��ty��M�q�E; %�{�����@��R�'n��'u�O/�	�M�7���?��j�0}V��: �K�]�s�&��?�ҵi�O�Y�'�x7��ۦecݴ7��`iB�� `ջ�O0)Ȫ)2�큐�M��O� {�(*����*�����9���/��, A[*`�|�JG=O����O���O��$�O��?i(G��t_TS��<cjSkƟ �I�����4{��iͧ�?��i��'�ޤ�KD)T�41�F��;gy<9B�-�\ݦe���|r���M�O�9;��!P"Pn�(�̈�w�́�B�
�?)�&�D�<����?���?�@��z��ܐ��1i��ʷ-ε�?������W�Dė���������O��`c6&�D>DȦ��R_`�S�O�Q�'�b�ia&�O��U�����^'7DF�u�R�?��X�݋/n-s�[by�O3X��	�o��'XJ�ʗjGl����&�ďRj͠b�'�b�'���O�則�M�`-�
wp�v��t�~�����vBz�`��?q�i�Oʕ�'��6��#�|��D"��1��Vz�lZ��MS�b��M;�O�tՄ͢����<��I�( ��*Y��,Ԉ�K �<1)O�D�O����O���O�˧F>$8���ڍL�L(��݇` Y�i���'�b�'��O�km��nD�:=~*�N�B�c��ÁSd����O�O1�
9��h�0�I�%��+�n�04�J@:b�X��扸r��US3�'���$�X�'<r�'_���`��$Q�0�i� N*5z��'\�'�R�hhڴ Y�`.O�����)���g���{��� ��W���O���p}B�'�ҕ|Ҭ�1P�4Y�ЍB�o�&�B�ρ����9ߘ�;r���?
������?���Ȓ1�R;ab�}���#FJ�!�$���f9KpG�9{��� �ڜ3�Z�d�	�����P����M���w-aL����" J=u8`���'c�i�@6m�7�+?!:3x�ɑ2ˆd��ָ%}�e��;h| zI>�*O\�?��l�G�D�5&T\8h�q��G~��e�0��WN�Of�d�Op�?�d��&V?�uY�$]�zz����#�6��D�O�7MD|�)�)��D�[��\�z�����T²a�a��07M|�|�f�	�O�4�O>9.O0K�b�e�8թc��0N���Q��Od�d�Oz�D�O�<��ih�u�'� �3��
inN`$�%F�P���'X�6�-�ɼ��DH����M�C��DԌ`a"�R���]�5���4���_�2e����$�ғ���ným���5�D4ݨ�Ss�-N�$�O4�D�O����O��d"�S4|��$Ѵ���!���;�U��ӟL��=�M����|r��Y#��|([L��U��f�Nb�y؀/M�-��O��o6�?���F(X�lx~B([4̀ � B�H�w�JP�	�3rJ�TgJ��?��-��<i���?��?�H�&�b���_i�p�(���?�����U���ߟ��I����OI"и��<�fy0d�� s�$+�O���'C"�'"ɧ�i�1!U�Փ�T���5�����SV��X��H���<�'/
�� ��\���{��L�x�28��S�F)hx#���?i��?Y�S�'�������l�>	l2p3��Hq��Il�+Z���'�67m,������O L��� G��c��,�h�Cd�O�$�l�7�=?�;G��[�')��˓
r��`�l:iV�3)�yx̓����O����O����O&�$�|R��dy6) @$��AQʝsr��*F��+
� ��П$'?!��4�M�;���t�rL�!�oP< |����?�I>�|��"�+�Mk�'�^��caW�b�
T83.�?�:xȝ'v�*��ğ@�|�\���I����i" ���C�M�Q��
B�ӟt�	ß��	gy��a�X�C�F�<�?�rtb�&�D����ҧ�#>�p�K>��p��	��MC0�iP�O:쩖�ҤV1�Y!�D1(N y��ZK��tW�|�6e�U��4uPbeǟ,���	�6|z����'j��X�g����d��ϟ������F��w���U�ڸ~Y6�Bq��!E�q8��'�27-Ŭv)f���O��m�d�i>睔�@b��ߟy�H\� �[q<�	ԟ��I՟T2�����A�u��Zv��͇Z�����j�6Ǆ /oFX%��'W��'R�'�2�'��;���V^�Cu������F]�`�ٴ3�di����?1���'�?���n.��p#Z�0Z��F-�t�	�MQ�iЬO1�-��ǛLA��XWJƅ�xE��� _2����â<��Vr�$S�������j�p]��j	�/�p��IH&B{��d�O����O��4� ˓ *�&C*=rb�?!�d3s���V�|���#�y�#g���L��ONem��?1ܴ^��})���y�<� ��B|Ш����M3�O �����:��/���﨡S�'L���	�(��� �c�=O2�$�O���O:���O^�?��qE�uXE���;FYR�s�����T�I矸�4"=���O:67M5��P'V՜`@�a�O�h�@b�}&�T�޴C��O����i3�I�N6�=�thS2]�����T��̐��^�M�b��O�Idy��'#��'����"";��)��Q
SB"����ܫo���'�I��M��T��?1���?A*��Ha@	�;*bpi��95�[��h��O~	o�?�K<�O>��#U�/������F�%��Xʥ��R��H��K�&��i>%K��'"��&��*��
i���³'��//��z�dV��L�����I�b>��'�6M86�P}pG\u,JI��iʼ7PT �!��O��d@��I�?A%]�(��(�0T�C�S)/8�i�f�%1~��ş�BҦ¦��u�S,~(�f�wyB
�z���υs����(�0�y�P���	�8�	ğ�	ٟЖO�vm�A­,�{1dD<@x�P)c�~Ӹ�a���O����OD���dZߦ�]���Ap`��V�s��N!!�`������H<�|b����Mc�'~�@r��R,�VM��`_�}[�xZ�'�.���(��hۧ�|�X���ٟt0�/�!g]�hTh�)��	�E ɟ|�Iϟ�	~y�p�ʼ�& �O���O(�:U��hJm�'��*C���" 2�	�����O���v�	Ez��4+�� ��5� e�����v�["�]%<e�|�.�O"e���.�Ee^�d��˗f�s��)@��?���?����h�`��Cs��(����+�Pi����
$�D�� ���jyR�f�H���?>Gz��v�E�Q�T��阜m��	#�M� �iݨ6]�*7-(?�F�13��	I�I0��kFi�#7v��ǅW�]����L>)/O���O����O6��ON������P����6"� ;�
!�b�<�iri��'���'��O����1 �5�@�8s&q0�7U˓�?�����S�S�]l���3/ͺ��i�� ?�9Q�L�?�*��'|�z7��̫��|rU����#��9���Śt � ��S��I���ǟ�Oyr�t�|:���O�',=���iv>cn.P����O��lZ]�u ����M�q�'F�挞�k�(Ak���6T~Ei��ڍf�(�'�iQ���k��]���O�Z�$?1���v��|ڗ)�7��#��Ү;H�����I��t������C�'AꚈib&��+̘�Ia��"B�P��?���2�F`����'��7�-�dȧ"6,�!��-RI�aS%A�{��t&�d�I���S '��lZM~r��7��联C�$B*^Ay��74M��kJߟX"�|�[����ퟀ�I�d ���,�E�$�(8<�w&�ßX�	Qy� w�\��e��O����O��'oJ����9_ڌ��n��;c���'����?���zA����I�h,�E�v�[<CX��(/��tYĂE�
fչ��S�e���B�#�t�A�
��W|fT�B�7��Q�	۟��	�4�)�cy�i��PpW"H^�0r!�.0澕r��ۖ(�v�;������n}��'2���V#ǻM�����4�$�'�'=p6-̄$�6�"?�֦����*���F:LB���PɁ�Ts1���5�yT���I۟��I؟��ԟ|�OcD(z�'�H�c(�>^�VjW�m�F�
��O ���Oޒ��D��݌NwMq�5�I�&N�<v�������x%�b>ᣀ.��u�S�? n��p�Ⱦ��i�#�A$�d��<O��+e(6�?�g$�d�<��?)��p�~��6��|R�y���?���?A�����^𦑹B`��8�I��p��O��li1AܝO�"�Ұ
�L��	��M���iu:Oʕ�fD�ژ-:��ѽ, <Ԋ��� [�-�40��E��k��57����ɜ,8��5`�� 7���4jRҟ0�	Ο����E���'���HE!1S,���F97?��j��'��6mXh�����Ov�m�s�Ӽ�T)�Y�u����4$�H�JuG�<���?r�iW��i\���2��W����&7>	��.�70�	O� (T1O>�,O��O���O����O���� ӊ`����a;D�"EZ$G�<��iS�}�T�'aB�'��O`�	-�i�t�
h�e*�T' 4V듣?A����S�'m��\W/�,\���`��T��`RWꍾH�v9�/O
HRh�)�?��,7�Ŀ<qF�)Ox�[��9h� ��&O�?9���?q��?�'�����a�3�A�`؇F1Mr�����D��0IvD�Ɵ��ٴ��'�p��?a�	����= p��D��i�DK&�X"��C�i��I�vT8zw�O q�<��B���%��8�B:ъ�$�OJ���O����O���#�ӹc� K��֌+�c��PP&��Iޟ��ɠ�M����D�Te��O�p�ï�-0ڄ]��(�:{�ؠtb�W�I��M[D��i��M��O�p��/ڈu?L��씜CVX�U�
i�� ���ܓO�˓�?9���?a��X#�iWIO8&�$ԋ�	��-W�a���?�*O:dl�t�4��ԟ��	T�����	zv��lѾ���"�����c}�fq�84�	x�)B��\pXI�d�Y�"t��gAR&	�$U�H�vf�%k(O�)��?q��(�$
0����$�Xf�<"�ϛ(0*�d�O��$�O���ɦ<�`�iR��z�ʎ$fd�)z2&�� �V���Y9�R�'��63�ɛ��D��(d�9{i���n�9<��P��M3G�iU�}��i���8z��r�O��-�'i��`�]"\'�չUʠmߒ���'��	şL��ҟ�	��`�	�����P��g�RyrX�5"ՙg�6��:{����O^�d(���O�nz�Y�֖^�*�ЌQ3m�$i�����M�ûi�O1�v���Jl�@牭{x���A�$EU@ KԈQb^�I��=J��'�D�%�4�'ir�'�Lx9B��q�L	ӓB��xaJD��'%�'"U����4 2�����?���	��V(��d�Q�b�1�d����>�B�i�7]K�I�t�(�آn$���P�g��'C�
H�����I�%O���K~"�m�O�����s��Al�#�P�&��NX,����?���?q���h�����7o��<�aE��/tt���%S�@�G�)���Οx�Ɂ�M���wsXZ@ν���A�%ֹf��'��6��զq�ݴ6��Jش��ˬ>��!��I��r$�C!f<�rD�<����"$��<��?Q���?����?y% V�VLؘ5h'rXS�\��^�93G�؟\�Iǟ�&?Y�Id)�U2����œ�A]��˩OҕmZ��M�x����½;�Ѡ��0�*h("�X�J^���Zd�剥c�*	�s�'4�m&� �'G
� ���?\�x����$@SyRR�'|��'�"����T���4m�-)��#�r ��#n�6����w�h!1��#{����\}��kӞAn�M+S�
�z�B��'��
GS���A�PR"�Iܴ��� `����'9d������v4�i��K�^���F�8���O:���O�D�O���3�S8n�E��I]t��	�c�$#Ѝ�'!�i�hh{�>�����˦�$����C/(@`��&[|���\.�䓈?���|z�M���MS�O~���!I1j�b��O�^u� c(؝"֪���)��O���?���?!�k��jvaЫp�Ȩ�F*�?D,a;��?�.Op(l�F�b��I��\�	_��(�#�z C�DP.*��뒍ΰ��$\b}��n���lZ���S���V.��У��p�����\�ڹc�O�� �-@RT��ӹ e� �C�	#F���%$�7K���1�\�Mh�D�I��I� �)�~y�Lx�f��	��R�"�nɂu�|;�fH�j�H���O�lV�#����(g�+
�ȐѰ��W���A"��쟸�I�>��mZg~Zw������O���'�B�2S'��UZ(��&�'m$�B�'v�Iڟ��	�����ğ���X���ĞhC�0�`�Hf>[fG�D��6mD�m��D�O���7�9O��lz�q�C��uڞ�2($ S���uo�ɟ(��n�)��-S��n��<�c�<�:��V�J~hBQ�]�<!��Hd'��d5����$�On�$@���E�/� h�-�M�����O����OʓTn� ��?	���?a��ʕf�������:��܈����'t듖?���>��'�!�1�=j-p��IE�#����O\��%��)SPK��i��?1�,�O�XD+�6*,��ʾ[윍!"O��ū��U�C}��2�b��'��i�"l�r��OP�D���?�;��9@��y���@#I91L�$0��o�.�lZ�
�Pn�\~2�ƴr|�<�4�Z�K���22,n��#)�jl�m���|Y�(G���1�0�#��4�q�f% �����黎Ra՟<�	ğ���b�A�%�^�b�oQ�سԨټ~��	��M'�i�O1�ء	'� b�Ҡ��;Z80�5��9��Mƨv�˓5���L�O4�!L>/Oxu1 ��ӄ٘C�ؑ��HD�'�6��o�p�$�.]����ũ��:�Ҩx��,¤�$��-�?�Z���	ҟ@�	�`�i8�$ՏQ`��Y�_�Sf�p�c��U�'�>$��f��?	Iu����W�U���sad��uM��c6�֌5�`�ȷ	:Rn�&3p������b��p3�g��iu�`���ӆ!�0�6,5�@��ƪ�&��X��b'��!"$Jӥt�V���ʉ# �E3�9�V�0Qj�C47|@��fl��D J"a؎?34Ӄ��{�����:.�Xr F>+D0 �o��5�
�c݄k�T1�؎S2��� �!'|0�n5o���e��ج�#C��N�c��݄O
�x��@0����f�c#Гw�܅�LM{�7��'#�|�۴�?����?��#ܯ$~�On�$�����7m���������b��/�I�M��c�4�	���&�E��@�4ɘ&��^d��A�-��Y���$�f 	N<���?AK>�1')��X�nH�\� }��ђ�:��':��=����?�����ۓX��CՎ�`wl�!O83�]��M��Iڟ��x�	Zy��ƞe�Т��
uT���v~�p��y�'I��'��ɗ%Y:X��O�h ѦI��&5 D�@D�2+�(�O&�$�O֓O$�Eb�'(F�t.��U��,; �]�v���s�O���O2�D??�����ħ��!�bH����Y��.Q؜iKB�i�R�|�T��$�=�I�(zڐ��H�+5��!bU�YI57��O����<��bIn�O���OZ� µ�[� �ґU�7�T}���*��<)���f���)_�R��sV�C$�� �����P��iUGP��M[UZ?1���?��OHMu��"ň!J�W�Ƽ� �i��I	����?�g�%im���O-"���0V6MȒ�Ddo�ן���ş���:�ē�?�CN�A�(2t�ʶ	{�(qc1�v���O>	�	� �K�i�I�`�	㊏�@�$��ߴ�?)���?Q���{��'v��'�����	�v��!�(�&LJ%��ʱO���C�$�O����O$�à��k("��!;���ɦ��	�&��\+�}��'�ɧ5�#S	�����*f܎�h3jE�����(z
1O���O����<���\�ml�nM�g�Bu���� b��񘰐xb�'D2�|r[�ȊF�O\����-B�ĭI�f��&�c� �I��	]y2F�a�����BǗc����eT=G=ɗ#�>���?9K>�(O���\���"���a��"N,̤���>����?��?���t4p���?���@�V�ڤ�	�~�Ƥ�pƙ�Yt:!8`�i�Ҟ|b�'�b��7^�0�N<	�a�,����j='Ęp�զ�	̟�Iӟ��$C����џ<���?BSNG������Xpb�L��h�����?���01�L�I�S�T͞�M��؆�E�>�����ז�M[���?q mڑ�?Y��?	���)Ok�Z +eL����_�u�P�Z;f3�v�'��	8u)$"<%>��p$�:ྡ�'�	b<�0Յe��Q�P��O��$�O���J˓��)B�{�P��\�+6��:����Q�|��*9�S�'�?�0DJ�cTdR��F-}�M!��# ���'��'��I��h�>Y/OZ�������Ă �RU*��A��X��+b�ΓO����VD���<�	�4:a�
�|)FJ�	I�ZE�U�MS��;���qY�Д'�Ҝ|Zc�~@Rvb�0+b�b�V���H�O�msQ�6��O���O������AS*L�R46ϴnh������H��qy��'��'��'D�C��ƺK��A�5	NGw�\a�jv3�^���ៈ��{y��L�FEP擾!�� V�76��%����6M�<9�����?1�y�(�'�Ȉ[��$�����@����O`���O���<A�C͑j���[��6��A4��&`�h9f���M����䓴?��b��쀋{�)Z�t�ܸ���$�˵�
	�M����?Y)Ox���z���'�B�Omҥѳbޙ"�J��p���.����&n�>q��?���90��q)��Ix:�-�#'�0����5U�"���ߦa�'}��ӧ�x�����O����$ק5���8XE�$:�`S�[ބQ��͂�M��?��I���'�q�Ɣ���5Ng�i��) �m�D�R�ig4D���l�@���O����F��'�剳V�@�	(�:�����L��P �4��X�"���OnAx�!E(|~ �e�V�$뮴a��Ʀy�	����3���ڨO"��?��'T$ e)�*r! x�cMUs�a�}J��'�2�'�" �S5X����[obY�	NV�6��O�P[�͛l}2U���I�i�Y�ց��mZH��W�2�`�3�>!F
��䓖?A���?�/Oj����xB�)`b��3ކ��Y�����'��IҟX'��	ҟ���� �u�XQh��2���"ƚi?>@��Ny��'\r�':剤Ob`��O��qBeMG�4 ��K8C^\޴����O��O����O�7F��� �(�_�<Z�#U/�2�>���?Q����PTJ��&>!���{̻���>�6�&K.�M������$��L���D=�Ĩˇ��xk�U�D���
�^�Mk���?!(O@�[����@�s���D!�t�0A"��<d�)(e3�d�<���5�?I~��π <�Sr.�3we) � �4���ٶ�iK�ɝm �޴{��ٟ����d�Z`�`�LA+X�0}��Y9�V[� 3�aPğ|�K|�M~n�t)n=s2��l�h�i�A£1��6-�AO��$�O
�d�O��i�<�O(n���Ә]�v��&�P� 
���0�b���p���.1O?��Ԃ��,o:�Q&�/1�K��ݾ�MS��?9�ꬹ�/O�S^�D��2���ЭII]�A9�k�(4����<�@S�K����䵟0���X�q���-��5(@�\_�&�'�vѸ�U��Z��N�ૣ�Q��k�$��3~F�"�������_1A`
��D�Ob��?�5 vb�Dp���ft��Ic�B�lB��i/O��D�O0㟬�I�أlҾ:b����7cx��JC"z�P�I"?���?����䘄1����'m�]0��ڒ<�����Ε1�~L�'���'u�'��I�0�M�ɸ0@䡝�~�
 �D
[�(?�Eq�O ���O���<c�p��O� ���3dX�G�π!0�z��s� �$#�d�<)� ,�?�H?	IA��X�����o>x���u���$�<��q���.�n���OT��Ɗ)fLO
T+RɈ�V43�6��s�x�'g�K��:r��y���	�$��Y�$�C�j�*���#��i剆j�Bp��4S��S쟨����䕵h�<�kC�~�`���B- ��]�L17�����L|�O~nZJҾ`��!6�25'�]R7�ŗ�]��ԟ@�	�?YIN<�'h_��q2�n�+�N
�7#���i�j h��'h�V�4%?�9Ӹ��L�CA:�H���;*K��Y�i ��'��	&4*�)�N��Ҡ�U<�p-�'��-5D�i�n���':�}�3�.�I�O ��O��JԮ�3d�.*����x��G#�y��)"�U�H<�'�?�����3��YK� �,���(��97�o����IR��p$���	ןt�'�Z�⠥�y��Q	7 ��Y��B���\O.���O`��<����?�f�A�wN�y���$�𑁵�U6�����ON�D�O�˓0�䑁�П�h!@H�,�6�`��ȕl�����4���O�ʓ�?)��?q��<�B�߼}����Ή�1Y���ˀ⛖�'92�'��S�@;��"��)�O�r�ᇦ&2hHd���9���Ȧy��Iy��'���'$��y�}��OJ*�YYP���텂$ZՒ��4�?����D�~"]�O^2�'�����=F�f�����-h�}��Ƒ�skN��?I���?1��h~�V����G"� ���[��ق ���R�lZXyb���P-�7M�O����O,��v}Zw"h@"G�/]��1���j���ش�?���~�t�Fx��)޾-ڸ�'!��$�x�mT�, �f���"6-�O���O���D}"V�h�H�V|��Z6��ծ1��@߬�M����<Q�����*���DhƊ�x�VL�7C�"pyЃ�M;���?��v$�4"4_�L�'�r�OX�C�R/zutA�B+� )ZF�jýig�'�"@����I�OB���O��C�
.J�%�JT,S pJGO�-��Q�@i��O4˓�?I*O6����(���(m0u1s���* ę�X���'l����̟��������IyR!B�[H��4/� MĈ�g�]�V����>)*O�d�<!���?I��T�è�x��|�炏�v��XH�EX�<�/O����OF�D�<��"ǅ`\��8L4��u�4n��9��O�@C�6Y���	uy"�'���'AĐ��'�h��X�<
��ҡ#T�H�m�p.f�<�d�O����O��mm��&Z?��i��˖�P�T�*=��Q
�y��aӐ���<9��?I�u�ϓ�?�����q�(��tѓF670i9��i���'{剃 ��q������O|��W�~tp|�Շ`��Y�M=.���'���'�B*���y�'��TҦ,F�f�̩B�A�h��@��d�ۦ��'��<�obӠ��O����@ԧuw�
�x� �� %�:I�V�ђf��OP��
U���Yy��Ɇ�[.<J������l���7�ˎ$��o�ߟ|�	��������<y��B��L8�lL4I�Ʃk3�W!ϛ���y�Y���a���?	&�V�>:��E���7u��9R�HcR���'���'��a��#�>�-O,����L��_n:L�*�J�� �<���d����<�#L��<�O�B�'	��_�-w��ڇa��v���ä�3.�6��OPA Ů	p}bR�$��Wyr�5F�LL!��ſUn�$qEɇ��$W�4��O<�$�O��d�|�N��vKp�����Cj~D�#����Ny"�'6��Ο�������H;YhS��ү0�&�S�mǢ������������8�'B��1Ff>�S��r��i��"�6KF��'!�]����ퟀ��e}0�I�R�P�aP1��;a��9҂��4�?���?����8bl\��O�Zc����K�%��,�1�ŷ@��]�ٴ�?1-O����O���W&ft�;}�A� Nu�<ɖ��VXc�#G�Mc��?Y)O��(2k�g�4�'�B�O�8�1�M�[��}CW�R������>Q���?���.�j̓�?�)O��?V��CƊѽlV`]�AB��6�<��)A8_!���'��'�dD�>��i���P�˗.hfH���	n�ҟx��0?Z�I��$��˟��}��M6��h���":ܸ�d��;B�>�M��?�����R���'�\@�D���Lk��O�p�)��{�^da�3OڒO��?a�I�� �E��K@��v&�Oʴ1yU�i��'��"�&W������O��ɜR�%
��A?���"�!}K�7��O����OJQk@=O�s9oZ��h�I�dq��d��r7:Л'�]<b&|��4�?�%'��'=��'ɧ5�7
v�
7�G�i}H��������!:�<����?������ΠG��a�"��q[���'�,R8~Xa�W^��?iM>	���?I��I�u���?��tc��n�T����$�O0�d ����9jXΧV�)`��l�(*�
�sC>&�8�It�	�<��c��	#ѐ��giK32�̀d�ܽP����O���OJ�d�<)3U�m��O��)	vf��
�Z��`��� �����Oj��3�$�O��}_�0}�	>V�č ���QVt��.�M���?�(O*�9��k��۟t�:V!(�Ҕ�*Oy��)�P)�U�M<����?�B����?qM>��O�"|1a@�x%����@��YH�m��4��D�#۔�nZ���)�O�I�l~bGL�:�V�j�쇩z�;��6�Mc��?a��N��?�N>9��$�Ȏ"0R��ǜ x�P-��M�$�*w���'�b�'^���.�d�O~q���2 J�<T	�����`7-O'l3�D!��'���|Z��!4��AǄD�f�4�C"��M���?i��x=C��x��'S��O&�9t��Dr�:u*K�s� с�� 5;c1OD���O����h+��!cɷf�(a�\�'��Yn��B2n���'�җ|Zc8	C�K�#�ؘ��Ь/���O8�f��O`��?���?�-Od��2�!�J�0�/ǲM��	頹2�\�H<1��?1H>9���?)�d�-x��Be�5�t���\,y�v-Γ����Ol���O�ʓpi��p<��u��gf���E���D� 8c�Z�,����`&�(����<i�q��:�
�Vh�ы�¼
J����	���D�O��d�OZ�b��E�`��T�1Y4��f!�])�(X�ȋ%:�7�O�O�$�O���!%�I3,�����gX�3��p�3�K�b��6�O��$�<�4�Tu�OgR�O�����%G�6ͻE���p��s�)��O���F'2�$1�Ķ?URj�*CDV�SB� *�p89�f�H˓	_�T���ihj�'�?��E8�I)R~��阂U�4=�ѧ�?jV6m�O>��-T���-��|Z�'KrB�-�(�������;��y�4�AJS�i
��'c"�O�lb�BW�%���1�)��cB���5����M�N�<�N>a��D�'Ӗ�ї.Y�? �9�X��p��}�B���O$��0U�r�'��q�d�|Q�1Rdk��=�@�"�N)ZЛ��dt�Sӟl������0�Q��Cz*��$GL��M���޸�T�x�OuQ��0�m�$Y�\����M�4��i?���O�ʓ�?a���d�OP	A��Z'Jo���#	��9y��P��¼$���D�O&���O���:���O����.�T�趫�3��r��6MDj"��ҟ�����'gz���o>�B�h�:"�4����&�@����.��O��Or�$5�	�V����)�W��C���F����?���?)-O�����p�)vj����'c4�I�i��}lz�4�?aL>����?Y�%�k��@E��CJH�"x�C�E�"1oZ����	DyB/�cH�������`Ey�� 7�����
�,9c�l�	՟\��#:w4#<��Opj�cCHթ�N ���D�ag0��V (}�o�<��Қ��{�\��� �{L�\b��y��>- ř!!�?F}F���CQ$����!�f�Ô旎5!<�1�X6HQ�P�5RU9�RAV*��5@lӘ,_n�k�KЖ�P�b�+��]h�bˣp�,=ٱ!25��j؎ ��6N՜'��`�7���� aH���媃#��$�dJŢn7ء����a����D���{^Tl�Iݟ<��ɟ,�Xw�R�'�IR�"	�@�0�91-��4���ȆG�<C�D���΄�n�!������7ʓPTD�c�M�8�z���-��RT���RCE	��T�Po��_�"| �c�x�7�I��Y#��j��Ɇ�L8D��	�0<����O��=*OJ���� �~ဗ�e[�
C"OR�8�(w86�����/�X����v���I�<	�H\������kKV,+��.O�L�V��n��'r��'��J��'"1�r�2E-���ԍ�	q�v0˶�/u�8�Ӑ��+H���+<O�|rM0X�؜y�bL�6�[�ʕlG��G�nI���?<O̘���'{"��E�n���h��i�JU��JLm&ў�D�C W'�ɛ���gN�] ΂&�yR
�5R��%�^n��l�/�y�j�>i(O���T��B}��'���Z Z��F�B9a�d�
�%Fc��Jb��۟�����DE;��E��Q���2�S�tC[�7vI����)k1蝄�(O~���ֻ'm�ɱ��.���@���Ǘ 4h,9���/ ��2剚 � ���O�?��&�}|�9ʣ �b@��ne����I�1@�Iw@����ūn�*����R�.Y�D�8'i��&�
t�RL��7����*�h�O��d=��@ӟ�����pH��߾Q�����8V,���|�IbVO�1Bk�jd��?�O�1�
� �y�*��G�8�Q�H��8記�� � d7l^u�^=�HG  �&���hE�q�q����4�bH��
�
O����6!��K��'Cҗ�����O�Q��	�"+{�,��f�w���a"OHy��d�� ��S!���n�<���I8�HO�S*@��YbG��hx|�)D�R>P����Iן`3�1v�.��I�4�	�)Xw��'"�է;WܦL2Ԭ�<�8� �'}i�ţ�)Qۤ��$G+O�qۖ�ѻ�LI�&ɞb-�;��O~	����,Y�(�c
�A8��3.ގcO�쫢�N�L�#�ĵ� c���O&�$>ړ��d�*ȶ����\��e�Ƥ֮>�!�݈aD��Q�'�b� ��*.pGzʟ*˓)à�`%�i�^�Uh�PM�	͍���s��'�"�'�"��w���'r��+B�'��H��hA;1n@��T�<��uI�w�<dj�#٭��d��˖�Yz,�r�	/���0�O�D���'��J9�X5��Ȍ.i��z���:m�6��O˓�?i���S�t�jӶ}"�d��,Y�	!W��'�yҥ�mx"	�v�	�R*��A��:�y��mӦ5may䉍~>�7M�O���|:��^�=����#��>`�j|xJU�?*T����?�/����iv�'_哖-6����IX�i��)ha,�:D�<�"e�A��4§)b�k�����C�(�df@Dyr&ā�?���iT�7m�O�˧"$epd�|���ED�-Tn=h�������Ğ�_�@Q�/UJ�.��d�������A{ش�?�a��-O��ed��:�JL�����<����\G
���?+�t}�c�OZ���OdL	�ސ
�i8�k�=��H�H�t�ݨ�Q[�|����Cz.A3A��H�i�!�A!uL�9���/*�|���|���'?�Kq��OH���i��6��l#���r�'���';?�$�4��e�CKP6�ڼ@VD_����O8���s@���x6 	�M��c��J���?�bA�F64Z2����|d|I�S�ݟ4��r���J7������I�h�I�u��'3"��I��X�@L*{F�j�.\�G\t��G.:���F�H&P��y��hO+B�X?,"2d������2����O\�.�� K��p���xh��%�ZID��#|����n�"��c؞d��	E�W�L��::��xs�a$D�,��P>R~��� ��2Q���� �HO�	?���Hh��m�>WjI  cN�c��x`b�H�[`���Iɟ��ß�0u�
������|Z�Eן���2rCx�
��,}��b�aS�[����dQ�{U�I�MB�M�f�[$T������`�������'��t�Ϗ)�$��f���X��'�� �(_֔ �qmǋ�J�I�'r6)rR��7G��pr�Y$�rHk�'�v6�(�S�O}Z$��O�1�T4@��2 
� ��'|<	��`XV��V�H'MF����'%4�)���X�M��ǝ.<ET�i�'gr�AlD&02(K�#�D+P��'J]��
F�&-�T�ٓe� A��'RyY`D4�rs40^ɼl�ʓQ�1���,yT�l� �[0xJ�y��]��@��
���P@�*(|l�ȓtzF�DD��PA�&1��ȓ�  "L�*i��d�4)Pqq�(��;�����0p�n� �	��4o��`r.�KX(����İEN>������@� �	0ѡ��)ȁ��X�t��ch�*�G��}Ot��ȓL��\I� Es�*�á�4d�`U�ȓ"�}�	$��̲B!�<�|��ȓ3��ŌF�\ z����ԅQ�8�ȓ�
H9Pe��)A��� N�>�r1�ȓ&���i�I5d@��.H:l=�p�ȓWb�yӥ#,a�R�Y ���A�e�<a�95��lp
_E���:��N�<�I�:F� Eŉ6��8�Aďn�<)�m��x�dȃCΞ�2ҁ�F�<���H>2����眡� �ab�Y�<a�O�l��N�?�(��oFT�<� �`��X��.���,+lD���"O2���H�7*P)�� xX��"O�d��!֏N�ȁ�Ԋ�| �i*2"Oj�9'"ϣ7�n}rah�$;H*dʁ"O���I�p -��� ,�%��y��)rv�KR	B$5ֲy���	�y��='�V�:�eP.;��7����y���sX�AC�� �腒�M
�y2K�5h�v(�� �E+�B^3�y�䏰r��T�g� +_>�J�և�yҪ�,#�0��@�
6A2�Z����y2ԇ(u�Ū�`b(9��# ;�y��Bk�@�HP	$:��X�M���y�g%��ˠ��|@e����yR�N�B��e�v�,R��\��yD�#��(pdF��PtrW ��y�N� gdQ��`����	��y򧔫v������/K�x�XqN�F�<�NC�DJ� ".�bX`, �Aj�<�'��f�$!�3�ْt���
�Q�<��&-���A��
g��DHp��P�<A��6f\���#b%\{��kgRq�<���F�?�6h���}�ze�j�<񂩀{4T�!i�~%��a��X�<�b�K?�� ␁=f���`D�y�<1 �Z���ʃ� ���qS�_n�<�&
�jf�]vKD�
����D�b�<	��Z�DZ uYi՛Z�V�XQG_`�<�L�,Ω��I�%d�<Y�j�F�<a2�ϾD�)8jM Lj��E�<96H�/_`���GM�6�����l�I�2����9Oba)  �1K_�zT�ͣ4�"��' rAi�`T:S��mc�)O#%:&��X�V�s�O^i��c��v��E����D�	�5�n`��
V̧]�IzqC_�	H\����=(�8�ȓ;L���O�ќYڃ#�4�*4�'�F������|������tw��/ ^,��A	�Y�!��03YD�{�#�'<�@E�7'J-Q��'�Pe�'K/U�ax���N��P�� c����?����l�H�!�z��j��a#p4S�nɄ�x2l�T�3�Ҵ'4,��Ti<�0<��F�e���<y��G�AK����C�h�A�ZU�<Ѫx��}i������UWfS�<�b�#o�R}�� ��t��iC�L�<��@;^�-��n�E��p1�	E�<YG�f�X�Z�� �L`��C\�<񵮞�)�.�Z&;�d�B�P�<ٰ�F�t�	�ufѧ��0`VFPJ�<����$!p��2��!ظ"OI[�<��o�s�`Ճ��[$�BP�Kn�<q�d��]�̈��PI
 BA�<i4		���|�����,�V��x�!�
�d�����+O�'�u��-M!��?!�rt��F�0殽��*-@!�d�Z�D�s�I��9s�IEC4!���|<u٥DF��Z�;��U�2!�d��s�����O�r�8� �ND�!�A ���T���x���*� ~H!���<���f���ju,��D���7!򄊯HZA��(�gfz�y�H�$�!�D�%,� ʅ�ӖlaxTE�5�!��@DV�e`v,Hq1�k�DҧC�!�_�~�D������Q��>p�!�d�#@����!��=:(9�ւ��Qm!�� �}����~�dUD�m0Z4Y�"Od	��8Gv`�͉� �~�`t"O�Y�e^�@E9��M�=�n���"Ox�������$eY�+��*y �K7"OTy�g�10�R��f�B-i9���"O
�pIݴ(�(c'�ʎOD@�ñ"O$���MR.r���0Θ'
���"O�Ic��ՑPZ�P[����!�� Q�b	��Dλ/|I����!�D�eq�PkQ�#j2���DӒ'B!�D�:{Wr��hF�*���-ւn>!�9o7�8�6����y��m��9!���^�~,���	AM�� 3����!�d�?��x��P�F���#�!��G?G�*<�Q�Z>���BG'�!��ȩ
6�T�>�H�1щM�q�!�d��(�0�c��X�x��?�!�d�V_����ϕq�q��F�k�!�D�ѫ3P�l�DQ! �Va!�U1 �1�`E�O�9R�F�+�!��72<x=0�nG��53J�d�!�ŧj"���"�6>�p-�N��P�ĥn2�g"0�9�g?�d ߯K���a�ѹk_�)��p�<�QML�'�rI��!�<�rdZg�ğ�;�)�6hB�p�'o���4��T����m^/L>Y��x��Ղ����yg�6J/68tÐ<�q��M�%�!�Z�'�����}�c�(c��O�Z�W�HG��{��	��P�"�# D�*5���"���	�!�$*���e�dU\l���7��:�HO>�h��Y��b�Ffʼ7�t�ID�rG�5�a�'�=ːN����"��g�1�}���'��Bk�(y6�8*��  ư	�FIS~�$k5I��<�a�G�i���0u팣��`P�]#^&�'��@��LA�O
��i�'�-�e�=0��4N�80��I�'���g.�_�TD����N�1dfA	��DU���Q[�Gn��c&�M����FUt�1�K
Dj� A�`9"ayb��T�EC��>�%`�4SMR	+fJD�BM��)F����f�Y
!EL�jR@Ёi12Ć�Ih��$)���8V�d���� v��1,��
�Al"����L<�N̦Q�\���̎F�ts1m��|��m	�'����b�M:�ܠ0�V)�����}�֌��q6BI'�h�Eﶟz4�~�)�1L��#�L�f�K�zQL �O)�5DQ;_}�2!��;Zt�$y!mֈ �(�O�%{%�O����π)��РO?版"�J5���X誠"�=N�?��"żn�0�a���� V���T"L ���F�g'L>���L����'�� ��'焱��ߨO�>�ya�Q�5��,��'�ꭺ��B�S���C�*g������� �:����5 �(A5OA�R7��{�9%�S
Op�;G�%��
D!T���@��S��R��0�@4����\p�]��S6��4XP����N��Ι&+`xY+�!��鶸�@�фF�a~RhC�h�$yA��=H&�Ȓ��06��!&�%s<���O0L�%O]�����ɐ��p�&դO4ݠcE�z���P�.�e�
�A��������䚦�K�"�(H����-���c��K\���)N�W�P`���Y?�za��mڝ�%{��'Ѣ��o.E�.\�Q��iW�5�'�����Ӈ�<�rMM#Q��c!8�]�W��#����+a*�x��XZ�Vm���	37o�!��2��yC�_ �����G0�p�@�l^�w�������@a9 �v�PG�]T+:�H +�7�DD��O�kz<����}r��Y��'��9�*�? YAS�E����yA!�?f�2�x�&��$�*|1���܃h���&B�&7����'}�+H�]9��;s�Єo�ɻW���Oh%�3#�1=�0ؔ�ڒU �q|�ړm�'s�^��#J�A��Dj3N$f|1��M+}"�1`�\�vc�@��	2�*�I.�)+tn�&H��牪ā����o�l�0`�)BƲ�)�E*Nr�((rb�>1��ӜO����t��&|��Z/D�8���'a:q��OF�<�Ĺe��]������hxd��%MQ�N
��g���$\>I���pTĐ^C`�λ]��%㕧S�a��Ҕ�'�DI�5#S�x��!��H����Q,D�g
H]�2��#��N�0E(#sAӈ�E� *
j��W�>��$X��d��ҒH��b�'W�$K��g5$AdJJ2A��[��Q��� ����� r��\Sbj�>b�h{�f���"�c�e&�|�'.���p<Y7�| jx��
�{K��;�`�͟�������Csg�0g-��fu8�����%�I�W.VݸS	�1u�%��Λ�k�^�z	�'�
��熔��t��� ��(Q�����(9�H��!LF��M3-� �3�6 �Z�Z�p�*�fE(�����I*���o�a� �̾|#����xu$)�N�! ��@����W8�0���(Jgd���P�~���W�'��,���Yn�3��+��T�'%�*<��	M�h��� L@�2@��V�B��&��x�N@A0��!H����ɘn� �	4D��0�VB"~Z���>Ә)������Vc��y���@��!��2,�)[����Hhq	c
r�DQK�>���Q��Wvp���I�G;v��ȓS�I��Ƅ"� �z���%s�D�n�i5ܙrE$�O��xce�<#]�q� C���8Z"O���@�4:,BCG�
I4x��"Oҩ���Z!H���A�l2��
�"O�h*$J�$�ء(�.əC�F�g"OX�b��/9zP;���;z�2���"OJa�'��Rv2�S��V�|�)V"O�-9 ��2��8E+�A�܀�5"O��&��;�8�P`�o���2V"O.(�q�C< �H`a�#H������"O���jM�G�ݐ �ЋT!�ӗ"ON�!@��rT����(; ��б"O������DCBd��΀8W���"O(��)L��� KA]Ӫ	�4"O u�Ƅ�sz^�0@jN#5kz��$"O����-Nf�ɩW�@�!�|�C�"O�����6n�~5#�f��Hp�c�"O>U�`o��p�VEЫd��1"O� �ă�,�#㮒�U�u�s"O�t���E�N�[��4!�@��"O������V4<ȅN38��0qa"Op�k6M�-J� ��B��s�X��7"O��u�@'Gh��r���C�ZMx�"Ory�e��1��5r`]�b�ԡ�"O��b���M�00��$f��p�"O>dK�dNt8���oU.H�<-��"OJ�b)��[�$8� )�PW8�bA"O`ă����
Z�eYg'@�^%�q"O�e����^�������;:
(*�"O��yD��|j���MZ�tZ8��"O�7�٦'2˒,Y�0:�"O�pI�NB,
v �`"��a~rA�"O*VH��������)S!Yk�<q�g�%��%�'X&��{��M�<iD��8I�H�#��D��!�&�M�<��F#(4�ӓ�[vh�K�<I�g�x��t�B �Y<�D��
I�<��T�Ew>\Q'�gDLU�Rl|�<!򧍴A� ��AH�%�&KJ�<��O�T��T�q/�؅���}�<�gN�j�h0���ϸ}��Ia�y�<yu��0(>@Q��>Iծ�aciFu�<�FEQ�Z`�T��g�%I���J�m�<�r,š:��h��CL-j"k�<�F�ܮC�@�����`��{�a�<a��S3�����i5p9[q��_�<��KI�nݦM0e��-6Ūdg�`�<�:p�0uwT� %��Z�<����|�)A���E�`t
��5D����Wh����}��=1�7D���̍;q�����_)���c8D�L:��I��(��#�3�V���*D�� ���L�9\*d��'��(�� ��"O |��Yk�a�`�:^2`�u"O~p���cI,{�oQ=Zt��"O����+G$�P��Ζ�<�,s�"O~$Pd��?���q%MZ�u�� �"O�"gg]b��Qc�MZ��!"Ox5Y��0���Yf�7Qj5{�"O`���=0G0RUi�#U�I��"O��P�H-U�����ǭHA���2"O@��d����H9�nˆd=L�)3"O �y#J��
��ૣ�.k3�(�"O���Dɛ�~�h�GB"w#�]�"O(;c7?��e�w�= �"O,@�B�Qc�H�F���@ɓ�"Op�2lˣU^�� �K�d�2�:S"O�Ȓ֠ۍ{���Be����p��"O@]P劍*p��)ꡪ
�?ڙˠ"Oޱ ��T��Q@Pd�$�"�"O��Ӧ��6s�(ѡ��H���ȅ"O�����N��*����Cy�!�V"O��2̏z�T���Aöwup}�G"OT����:\�%���>id�<��"Of�bA.I��m���H�Mm�\�"O4 ��!��MΨ�U�:iX��у�Op��D G^f\��'�,�c�:z�!�DX(7ᾬKa$�i޼�I��*>!�$�����ϐb�"�G�4!�$�L0�
 ۔4n���P��!�*;'�y�f���0���S��֌%�!�I#9<*�Ҵ�уN�����.�1�!���9�x@��ƻm����tc!�D�� D��Ib鞒���ۑ��(~�!���:>��$�;��ȓ��..�!�D�6��PA	�b�zTi�(jp!�^�\y�Ybs)���>�G_&nY!�$O?�AqRS7f��q�&@�.Y!�AQ"`��`dӳz��9Hp:!��Z��1H��<X�F�A�:!�ˬBx2DX���-`�E���")�!�D��f%���Q
46����]#�!��n���S$w)���S�Ip�!�$Z�:�P%bJM���5à�C�<�!��I(:F�p��P'*�]b��T�
�!�$�)��Q�6f�D9$Cٷ�!��?I�B�qB�|ڲu�)I!�D�;$j(m����<�(i�$"�bN!�D+e%:�#��	�h���bg/!�D�]��\�E�E�q,���&	L!��]=����Q��S&b<Ð���*!�w?��[ ��?h��������G !�Dd)�Uq�c�4� �)�kG�U!�d=��eȨ8�$Z3j�:V!�"�*� ыߩE>EQU(�6_!�Z�_�0�1Nkz�y����r�!���><�ASd�CD6���Ɖ+F!����5�pa��J�<UH$��	@!�dg;����I� �P��QdR/L�!��[��� ��y��h���-.���mݱ��R�OCő!)�9�y��
� z4ږ���TJ-Ʌ��1�yb-��cg���D��*$h��ir���yb���|K����j�$+���K�����y�oؕ`����
,-1F0#�3�y�m��	�\ xâ�2�ݘRb��p=ɏ}
� |�'�ؐ��l#�ٱ
G�!�"O�A8�n��o~$�9&�ɪg��4x�"O�Գ���s�\X��Lt�ł�"Ob�Jd��.2�<9���}g��A�"OZ�u�-�6T��ՀxVyA"O���ǋ
%a�mA���?-�Q��"O�IhY�����L�K��`x"O���e ��K_��R��*P�x9�"O��Q�ԧ�T$�aE9P~6<2F"O�qS4lZ$�~-� fz8\��"O@�I�1�9�v���m>���"O�U(C	)Gńqb����QU�!`S"O���a����A#����ճ�"O��R�hs*8�!i��*���u"O���@��Q���r�ū*bQ��"OFԛ���\�i�dLN�PASE"O.�gNƀfX��F�ϬM���"O$��DbF�=����'ϳ+  ��"O��bG\O�q�D�J�ze��"O@�a-�rvIYb�)����"O��	b�~k X#G��
'ѲY��"O�`�/��T.��8chU�%ꀔ��"O$
թS��>)h�!�,ָi�7���OIJ�*1e�/M�p��;^�Z z�'U���C������P�ң_���:�'N괸D,��q��%˗i�_�~(R��!�S��?�U�I�S�:}j��Y�=1#�	n?��]t��m�$dN�5�ʎ�za��	,�t:r��=�f\�vݳ�^H��CI�E�V�E4�#c����	�'�Ѕ3���MCj8"�X���k	�'�"�`�O},�+�)Z�OU���'��2&LA][L��Ƌ:Ju��:�'�l�p�	�^��;0�̖?�Ý'��R��lR���0��}(�b�1�y� A �t8��AIq���c"��,�y�$��ms�`�㋂o��HQ�`�3�y� �l>�jw Fj�vQ�&]��y��\�][�j¢�a(Ґ�m[�y"թ(p�ģT��-��DY��yb��f�p� ���*���ұ�y��ǇCH$0Q�ϊ3��H�E���y�#�?&k� е�3u�z��菀�y�Q�i�#r�'l �F��y"ԻK���p�b�4t�4QF Η�y��S0?攈ǎ�< ��1cdnF��y2Bc��UK��Y2#�ق��yb N*��y�3.a��#��S�P,�C�ɭ'B��S��C\@<<��oP�i�ZC�I�#h����ȝ����A�6�tC�	"xΥ�G�Jh8y��,�J.B�+]4ReP�b�9�ʀf�Q;"B�	1WvM�5�4��L�Td#J>���r؟�k6j�	C�̠���X�{Hl�$!,D�(H���#�8Q˕�>p�3`�)D��T��e���79��)�1�'D�<�0�����B�"E}��l
0� D�x�q,V�(pI�JĊ+u��95�>��MdJ����R�T�~�y`Gߑΰ��MpЌ���\�����0(ߎ����r�|���C�G+�	*�C_�v�1��dR�r��;%'�e1�X:\}�ȓv ��.�:1�$qQ�
L�\��K�'��I �c^��l���b2S��� (a��f�*k���&$ڱ%�(A"O�s��.$��#�=
:���"O�tX����(���ߗ9���<Oj�=E�dB�g��`	�AD��ٲ�͔�y2φ/]<�0��-1�\e˕����y"`�+B8pH#�0{�$h�@��y�./v%��k���36��#!@��yr�!6ߔ����Y#>���ה�y�o�e�>�z�b�� ��0���y2B]�4{�!��k	�:��a�Z��y��T�L�&<�������fė��y҉�4d����ª�lڤ��@6�y�b3OABd�RB�1j/f5A5���y��Q,ah$�bpa3,Ř		U��y�C�s� 1Y�./f*5�t�H�y¤ƊgGCBg�<+I���JM%�y�lR�S��B����8�!�X��y"N���z8��(L�,��I��y�.O��� �ޚ	Y�������yR`U f&�����*.bi j��y���r
<*TF�Ud����y2��y�L�W�Z�HV �L[�y�-�I�|�
��qDX� b
Ɂ�y�E۬7ꖑ� G��y���ש�y���3(��Y[�BR�4)�J�"�yblw3v�:􉒇>�0��$@��y�A�8s��DTNQ�2���� �>�y��W%=r ��ߛ+68�ŉ��yB���C���(����)�9�y��Cy ��� ��$
�@�T@�&�y��-Wn��C��VlF�� ^!�y�,�1X�@Hc�K
2=�P� ��y҅����u�	�"���*$�� �ybϞ�x�6}��l�>���f[��yRH�%��P���onu9aJ���yR�V~`�&�� /��}X�O]2�y�o��Q^��R�Eֲ:K�\�G��-�y�)	/�����*+�Td��T	�y��A���MSD��)���˰��y��T@��8�'#s�4�:E�]��y⢌�,��.�z��0I�E!�D�����b#�5�$�(��H�!��G#Ĉ��_!�*,��ҩ#�!���t�8]B���j��4+��]|�!���,!u�\r	̍P��b�b��!�Ė�I��i!h:z-N�����!�DW�iO� x��;"?��Y�Y�4!�d�WI6�S�d��J6�(
2���;'!�$�nB�y�1㔼`-D��sb�/!�D�_��)y��v����&˛�?@!��[%�r`��`�8}���	��Ղ9-!���1Z.�5a�!9��i5�ϵW!�Ij�E���3�Rx��CT�!��J$�0y&�G�`}�`���F2�!򤈝"����,L���u$
�d !��Gp#���u��:� �ţ�?�!��i!�Hif�{� �k�]�!��H5���'+��S�0�C��K�!��.�Pk1��.u%8y�_��!�$�?Ä����?����uωT�!�$^�3�V�qI*ц���Qq��,TA� �ʵCx8)PB�zJ���ȓ]r�L��˛A6�!��\ B*.���c�F�`�)�yR؆�ے4Hh��S�? .�5
�t�v���;� ���"On����Ն�ӱ��,��"OTh3c�Q���sV�(s��88a"OnD3����>���U��:D�YJ"O$la!cE�X����Bl�X�b"O�-���6!�d��.�m���"O:�DƗ`x��lJ,h�yq�"OB����[�p����E��=���"O҈��e^ޘ��Þ3���"O�s�KK�{����chP.m�J�`�"Oд��@Vh���sP�;&~��۳"O���g�8����&xc�H��"O^ʧ
�*WJa�Tb�#w-��څ"O�3C�ކu9P""�&exfh�`"On��A�G�q4T�x5a^���"O�<�q�î!�D�B� �Z�(�H�"OM���<�U��Ҁj��)�"O���W�7�E�"�i&����"O��j� �s�H��a�$20�W"Oj�@P
@�)��@W /hi"OX馤G$|D�����V��� "Ol���ò]׈�����
�@4"O{v�_�ML�1�'V�b<�"O�=� �%��P�C����"O>821(U01$��X�����ͺ�"Oh���G��:ULܯ]�>�y "OzɃe�F�?z��P��@/#\>���"O6���NA
;��Eqd�5ϖ�y���s�e�j��B�>��w�V�y��� �"�Ư�:#X8�+�yx~���^ܤ���H��yB�ݍ���Y0��Xd�ћ�N��y"��42z	yVFQ���1f�I��y�lX�&PD����,A��JҀ��y"e�8R�`qf]!K1��H�����y2(;r�ЁH&���I����l�.�y����J�~1��	=�~�����y")���@���H8 _�R���y"�V$s*��df^�r���[��A�y(�P2D�#� T"|@j��P�yfE=_�@���o�+8�B3L�y�A��D�,���ͼ��c���yBk[*t��u ����h21���yr��R����^�t���;�y��X��3�	����h�T0�yRɉ=���7M�t�$�{G���y��'��5��L�m���Hף	��y�����
ͤ\��qh�D;�y�l�;���!�_�<<Փum�y�
��.Q�҂~����3��:�y� �$*~e3�]5j����M��yr΅�,�����;h>�A[����Py�,N4h�:�P� �d,I(&�o�<YW&�v$4	��!YvP��&΍i�<1a憺N��) �N�E�$��Fd�m�<i�'��a� �1��*��N�<YA��F��	q��%��Q%"O���7�Z�hp���Ø0�@ya�"O�M2�a��k�2 z��@$,�@�"O�m+��AmAI�c��q術`"OtY��_��<q"��&u���W"OhQ	�K�XBt�6� p��1"O6X�$�}��5�f�ީ;XD��"O���6@J��HM���$>�ܠ"O� �D��f �-����Ũ\0V P|(2"O8Qs,���&�W�	�� "OB����ݾN(��Ɵ 5S�i��"O"���ŋ�Bv���C�͒4i�h��"O�4�'D�v���`��(0J|�"O,�X��F�,��yh��Zg5�"O�I:��J.�d):6l+o�i�"OvIY:a���
�@�Q��@1�"O���vA�	�4��
*M'�ݲv"O�4�����k8�,�@	T	D�u�V"OB0�kݞZ���:��]S�"�V"O�L�dB�,s�x"��`��Ѥ"O��A�̞�A6���R�ʵGʬ�ӡ"O(��deN�;B	�Q��1Z"�t1�"Or�8���|������P5i�� �"O�`q3�
��`��+d8u"O�|C1ǉ1FC�r��ՉU+�Th�"Ob�"�K� ���Q�,`�����"O�b��]�WĄ�@�R L���{�"O(��+ם[�X)X�Y��)�*O�m� ��|���2ю�,z b�'�H��½1NLȧ���F��'�,��.�!�r��v�)1�X�!�'���%��I0�Ц�ֶZT80
�'��6b�8�Z1v��a>�8	�'� W�0�
��5AF�Qn��'d��	 b#4҆ a��ǘGS����'��xcr�H<.w�L�L�(=� ��'�Lm*���[�BA�bd�$�(щ�'o\uY1i�mmRB'n!s	���y�IL��d@l��j`�2᫝��y�U��am���9�� 0�y2��!|lH���P%Cx!�1!���yb����P����4R��!�1Aϙ�y���rj�c��7��hj�!C��y���������*r�,S�l^��y���.���x��s�F��tbˉ�yRBY�AɃ�Kh�FM0�
���y�b�#���w)%vQ�	5#D/�yBfկ}��,�v��� ����y�h�L�R(a��X��Z��yB�DjT�"�*EF:0�+I��yRg7y���kQ�I4;���p��ybcȓ,d���,/g�3 �_��y��0�&��`7,:���%V
�y�J�C%TQ�3i�/(�(0��mÖ�y"H�<�Q	dˊ6'����9��O�"~
eOǸ�L���CM�8���]q�<y���^��y�ċ�	(��(y�^o�<ɣG�-N���[E	ˊaH��#�t�<aC䒡x^�M��CNRL`ԋ�H�<��?f�"�2�k�sr��%i�<1p�֨S�Dxۘ�(��EE	�y���!�"	idBhI	����y�
Ì)SP5��z�ʬ�d�ژ�y��[4�T��,�jx���)��yB��@�2��S-rs�i��M��y�,PW���4�X'YV`�{�։�y"A�#D���3cڗSO�]�g�G;�ya�e�,�"�i�>A��l&Ģ�yB#޵g������P�7�D #�!0�yn/(Ҩ��D70z�������?�
�',f�!T�Fhޥ%�E<okX�	�'��*��݆%��-JdO�k>��"��� .��Ő4Tr �����16Xc�"Ol�A$a)$�WF!ޥ��"O��R�E�RH�-"� -i��L"O�����B+/}\MÕ�$u�"O�al>gn8�1,��V�h�Ks"O�Py�&	0)�� 0��45j�q"O�ف+І6����Y��4"O���C��'?B00�jE&�8���"O�%�v���qi�g.n�h#"O�*��r�� k�^'�U�"O��!��́L�z���.4G��k�"OP}�smL4qɂp#���28��Z�"O��ӏ�7]� �]�8&��!"O4�p�A���)S�晭Y�����"Ob��N���Ɓ�!,�/9t�"O���rC�w��e��n_L�bB"O��j���V�v=c��Kf)�3"O�y�q�P%V��b��~��Dj�A ��ϟl��	2Fe0����ґE�tyԢQ�hJnB�	�Id�a8"�C�,�3bMZ/A�BB�	�'� &K%e��苲���@�6B�I2���!��=��x���<B@2B䉮0�"���b �=�T�!ˀ�"0B�I�%`�:cA�w� sf �Rb�C�	�O�A�HӞ=�D���h�*��C�	7?ި���ސe(s4㙚NRC�ɼK�����5��ɳ��@2:C�I�)p$3'�ÜX*�9���DQ�rB�	)����'��$�h��V�dB�I;*��r���`�"\*D�;{��B�ɝ0i�Dh�(C��SQ��"(�^B䉘h���PrƐ�����r�+rG`C䉵f��Bf�ͮ[.��d�J��XC�	�;dr033#_�~�d	�%�
~��C�ɦ<@z�R�S*�tiVjJ3��C�I� �@�B$�w�Y�S�M/v[�B������dL�g����熥��B�ɷ	~���Jǩov��Uh�(\AnB�	�K��������V�� ֲ;��C�I%V	h]ؐ�0#���q.�9�\C�+(e2�Jŋa�q��&��e C�2Dl�uE�
��E�"��:(�DB�! ��]�6A�<@�48��b-vB�I<2sBi���x�nh9��Y��B�	�^1�}��o^>&��3��+��B��7p�,�f�H2,��! Q��B�ɂL����2+Ƒ'{�=HW΍oi�B�ɒ<#�E��ļ-��8�.�;]��C�I�y�x�����3���b��)��B��	=���H�ɛ4Z�1�숟.�ZB�	%>K>��f��68ĥ�dAE;C\B�ɨC�XP��H�blv��@��C䉘B����C۲�T$"U[���� �d�]��YBʗS�N ��Ƹ-+bC�ɡ{�����ZH���6�Y-RC!��;����a���?��k%D!�$�n
�X%��&u��pe���!��8s�dL���N�C�U"�_�r!�$�$b[�Hc,c�	���y5!��L�P�f�acÉ<M��@�V� ��:OΥ�@�I� />����Mu�H8R'��F���(@�3�0�sAEn��A��"D��ʤ�ϲ�l�� ߟC�x�V�#D��:qh�<��أ!k]�E�)��3D�� &��C��_܂x�!n�,kS��Xd"O���$EU�F��U�@ tJi�"Ora�Q Y,��Z,ƂuG����'�ў"~��O<ZHDZu$�+Q� ��6����'�az2�H��Fl��G�JT�]s5���y����Ek��%�O�w殜�4hJ��y2��)^����c�{Q�I�åS��y����b9�#��,B\|Ȫ�"͸�y©ZD"�Е��1g�����y�Z�x�v�H*j6�P�F��y�JC�J��Q�Z5��Į�hOB����5�*y�m���A���#a!�{���2��6K��������!�d�>lR�*�h�0X��ƤC�!�$әo��A6[��ڰ�!�dF8#~���DR^���sh�0z�!�DJ2g��⁉V�d��psHFx�ў̆�	-������q���õ'�m�D�d;�S�O�����
�a���(�S�xj�m�"O���Z�r����ˁwX�t���Y�'y�$O�Bo:��DE�����ƣ��-��O셙A��`����+9�d"O2��H��	�
����?40b3"O�	[Mq)���)�� n����D�OJ���Q=A��`�7��E�T٩�۩�!�X�iu�0�!�a �C]�!�@�/g�p`��x\"��wC�,t��7O��@C�:~��8� �I'k3�MS�"O�8�2��r<����,S��۰"Ob-�h�4�i�CKL�"�8���"O���`d����
"�Yc��IJ>#q�)^g$���+��A`��`f	$D�0 ���+�|�T,\�" !F D����G�DJ���r��(\�T���=�O,�d	%,�����֔@��r%X����$#�����[GnUIB�	��p=;w$=D��z�3,�L90 ǻ_j|](w�9D��I�H[�-��!�ɝ�j��t�#D�<14��3w�6}�ר,	�ӂ0ړ�0<��噀V��E�r	�+C^� ��KQ�<A�O�ư���5�TPs(Jy��)�'/Vq� �$�Ḇ�E-��ɇ���ط�~�����i�Lm��&A��j� �,Uw�%@p�H��z�ȓp� 4)�B�#��#�F�_�4Ԇ��^,����Ȣ���Q+ Q(�	ڟ��'���>Q�+:<0�TϘ� J�_�<D���t/\ɩ��2A��w(^y2�)�'7� �q��:�@]Y4�=�Դ��o��I�4&T�p|�\�1I
:���ȓ*�|d��Ձf�>���)�h_Dԅ���q�2��6fV��P���/R@�ȓQ�$;G�_4�:PC%b�:p��'ў�|��
�<m� �!W�u2t1��,�n���0=�D���<n�h�V�ޔ~�:E�1@�l�<�ga�@C,�(s�F�Tٞ���Ng�<�a+ϱ?k"��(݄N�ʅ�c��c�<�7�/K���%oԿ]�ĐS&,H_�<�0���8%�B�&�(�a�FYyr�)ʧ>h�آ-�WҼ����!���$���I�Sܧzk�I�T�-~bLQ�G������4�5a��+.K@i��]�5p�T��^7�1�`j�.u<%� � .��$�ȓs\���.n��ӇU�V��!��S�? �����z�H����7/�xK"O�]q�M�x���5�h��g"O`���6#v%Ӄ���:�0�["Op]BԨҎYk�б6�FB&69�3"O$��bfT�t�x���<�D�IZ�87�&F�oX�vZ���#�R�<��� ==ڸ���`�<t�j�i�<1� \�R�`q���2r����F�^�<��Ƙ�1�z���M�g�ti���YD�<1�lާ5S*�"��#tIҵ;�P~�<Y��7HP䨥��enb�S�B�<��	@E X�q`�M�a���q��d�<A-�
�nEQ�(�V�<����Yl�<i�����0�����w�Q�<�$��,��Bڹc7�	`��N�<���_%B��c֦��	HAb��H�<a�$α8��V
�| \)I�aV�]�ID��t�����Œ���$(;�A��?D��Ղƛ.�l��ʖ/��E��<D�X�V�g�AX��z��A�Q�-D����66-X�K�Bӯf��e��6D� C����y��"5.�!/�!򤉚b�f�J��0m�&Zo0n_�O\�=��:)p�,�/*t���ΒiO��+��'�!�Dh� �d��&u�<�Q�CR�Q!򤂄 �Y�u%�2�r�U�zU!�$��L����)ިXkT���l�7!�$�2(�H(��M!]d���ю�Y2!�˨Qz���Z)K��1�-B��Py"��5[��m!�.�	M ��X��©�y�O9-V� �!M=l��Bϔ �y��Κ\�R1��iK��f\H,�;��'Uaz��	�Z�تtJQ�^-����y�f�F��@�y�pḱ	C��y"K�]�рMѱx�`��e-���y�BM�e��(=T�I6퀗�yb Q��:�a���V��a)v!��y�c�(a�@!�eN;B���O���y��Kg�h��Q�+�zEå�E�y�K�jxE:v�&#� ��3�ԍ�y�C�*O�����֋F����y���H�#��ΏU��qoQ��y�b_D�T����8..$�w�K��y�W�'�vYp���}�(�Rwh���y�b��S�d�u�&t��@��	Z��y��:jؖ��$�Ѻ	xݺ�)���y"�^(a~}�#Ě7a^P�JFC��yB��j�9��C�RInM�RE��yR�Wd�p��k�B��Ep��Ϙ�y�Ѵf�.����A!|1f�\��yrU4�}R���"N��L�@��y� �s�R�ˍ�fY���yb'J9���k� �4XE�[��y"��j�2- �)�>~قс7. ��y��B�t�ԃ@���w�>��՚�y���J�z�����h�F]c����y�$D!��=�#�1HZr�y��b?D��b��ŤX7Rىqi�1/�`�*6 #D�\KI^�,�8]E(0N�BV!>D�D��N���b�Q��LC��dB(D���@�<d
:����3b���j�c�<a���Qh��U�P;^Ul8�Tl�
B�	�U�A����$y>��ȩ)(�C��(�"4�d,]�y����T�4H�C�)� 6媣�ȅ��]�2oZx"�7"O��H�i��Z���M�\���"O�� A�$���J��ؔN�<љQ"O�D(1L�$R4�Ҁ]�"���"O�S��ƕ[&M�L�/�@��"O����ʲH��4K��/�D��"O���A+�?@`�c��A�S��r"Oh���Jʪ)��Ι:+9t$�v"O�Pp��5(q!�MޯyE�$�u�'�Ғ�����2U�����mNqc|$h��-D�$�k���q"���h�P�c-D�`�@�L*Y/& Iec�=8\����+D���a@
�g,�[�Ox���)D�p� $��Z|�[�C��]�Y�L2D�81�]�*�����iq4�.D����b�1+Hl�Ɗ�E༥�j+�Or�q����fj� @�BԢ��7>��%��R,H$P���8zb�J"*��g괄�:̬�5�ч�I:��Y�}�ȓa)@�{d�V)Y���*�{}����Tq���>)���g�!w��l��Qj�Թ7���-��I��*�
!Bh�ȓB�Mp��6N���N]�f���#�>|Rc�	W�Τ:e,�{o¥�ȓ]/Dy$aݩG(Fˤ�R�R�JćȓK��Q0D6g������|����+q<��"�̡v�&|��JQy�d��1�B�c����$UV/��`�2���Z�X�a�ϓwjHb�#ӊy9(M��D��Pp�/~���1y�&��'-D����H�rb��E�'7� ��b)ړ�0|
E�̋M��� ��΀+�2��`bGo�'�axR��@?�0j��7w֜� G�Ö�y"���+Ң`�A��)u|�������y҇�/��AO��y�D�)�y��1/��g�NG�,�u&K��y�ʊ�vQ�NÙ9�U��$��yҬ�!���"�I>@��X��@��yҊ<2�^QsMO�6��������0>a$/D�7䕢����N��$l�T�<�F�	Hd!`#ʜ�Y�|E2��Q�<i�Ȏ�$ $e�u�@�kA�=��C�N�<Y�(^�y@��i��r<��y���Py��' �1qwO3l�a�('8� � �'�8���#H�ŚH�Bh�Uk��D%�N��R/Cn��]�#�/J��L��"O�r�/�3L��aT��z�T�3�"Orػ5H�!0��x0B�U�x �5"O\ի���f�@����E��)q�"O Q�Aa����q"_��c"O�I
�I˄5,��uK�I�K��'O��!3��#Q�f�OV��@Y�+;��Y���� �!j��F�5�3 �v}�C�	�(���C�*B9E�e���=X��C�	<@j!�mWN]N��_>A �C�	�=<� ���2���^�L�rC�ɜF?:ȹ��U�P>q��.�0w�B�I����aVGu��m�4��7a����$0�ɏo�����W0D��Ё�g�
J��B�ɓA�9���RP��#M�
�pB�	|�`YK!D�_�N|�>7pB�I�>C���W6C_:L�e�ШH#�B��-	�tC ,��V�5��/TPC�I4��@���=RS+FM~˓�?q��?YO>I�y
� <�Ia�V�2i��x��E�'��(3-�b*�!��$��1�5�d�Oz��>Q �'�&��d�7�?U{"���OrB�ɢ=�5j���F���4�M<C��69���S�LQp���AaK�?8C�I'�(�P��BK����N	�36��d-?3%�|�ѡ������oJt���?���On������ �I�6���q��3�S�i�	oPl��!皢y����eo�m�O��=��P�!��2��	�Ճ��p�z*r��F�Or�`yv��>�8��!c�7Q��dx	�'�
=���s��)a,X�Yv�1X�'N�dI@ 'U:��� #B:Z`�9��OH�:�
����cfR�k�
!�t�'��[�)�'U~�u�C�=`^Ժ�>�V̑�' )qdN���VȠym����'8 Dyw�zd>�9���p���'�.(����!u���	b�I�'H��x���$pTܐ���2f����'��"�#�5;dx ��	�W ��n���$J����e
 &l����!�5�_�R{as��ܾ'�v��ȓ(�p��߀n38�
�X?�l���/�J���`��	*�;I���$����ɐ|��p��ˇ=��'���H��C�	+�xih����G�U�C�ɀ6�����q�T��JB 5�dC�I�h����c�%ZնxJ2�@���hOQ>�8 �\�[��x�d�J�wI�5�,�OP�	(�<��C(,e�7�Q*��B�p�lm	�'Sɶ`)��B�/p���0?i�N�<$p@����U����?-M.-��4���Ŋ�NR9B�4b�xń�	��m��-�/4~���Aq�.��F|
A����$?�t\)���U��m���+!I<�r�RįW%#�(G{B�'��>��#�W 0��@���V�b��k�<Q���N�𑹳a�㐸���i�<�2䊸N~�bU��TxV�13�\�<�v�U��Lx(�h��^h�p��V�<���Eô ��#[T� 7�V�<��(N=| `\��*qQLu�ALR����<IW\"���B�_\�@f��'Nў�OrDl��
P���G`�5sMs	�'N��M	�s0�xF&:�$ta��D,�'rPșv�	1 �.x�c�t���:�d�!A�&$q��ҴDS�p[f���^���8�kȤZ�|`؃�S�
@�E��A�d��T�����+Q	m�zԄ�	F�'��,Ti˛xf�(y��� ��'��B6�M�{�4�A����~�f X	�'���*̌�բ��d�|Z||��D�O�"|т�rCJi Pg� @
h��Ӭ�B�<�
�=�p���/ʮ�5�_c�<P*�5���Qg�����i*���Y�<���� yL}� � d����/�l�<aV��� ����W%�zn|x@F]h�<��!�"q�B�Z���Q*t�a�<��Q3%I�=���1��1"��D�'a���ܭq^���Hˡ��P��A��yfR�HQlD�M6d�!�D��y�����n�Y���.54D��L��y���9��l�v��5.�2��e���y�_$+���rc��[쐰C�Ȕ��y
� r!� dKm���Іi� ��ٰ�"O�����4"��E;�ιOR4 I`"OPu�� y	�I���)g�D�"O�H8S ۇ%� �C�%Ҙ<W`��"O4ij!��kJ���K�!i���T"OTe�!��:+$�Mz���n��r��k>1�2�F�{'܈��nW�/(v��7D��CG.�}�Li��O�PJ�Y��(D�$�+�+�@�r��L: �j�+ړ�0<q��Wowd[�
��<�y��L�O�<1,߿�P��@��.bN h�m�e�<����	e�U���A�f����Y^�<�K\�fð�% ���&��G_T�''?}�%�xw4y��P+8�� Z�	*D���� A*N�������nu��'D�)2g�-#����$n��tJ�J2�7�SܧM�����2a����2��a�\}��_t����ӛ(tސJ�cXQ̰���ޤru��<LQ�	��[u��Co�����X�<��Rl��s32�&�$G{�����M��aV(E��i��1��x2�3S�KØz�
K4HP�2�J��'�>�!���u9A1A�T�%+�1�)O(�=E�t�	?(�Jq��N�j��`�ݖ�y��j��s�Ƒ��ڳ���y�`�:Jk�tt������y�ȏDJ������?�^��cÕ���'ў�O��T� 
�R��GY�0/D8�����M:�����B�mM�4��\yG!��6��1�)���6DZ� &'5!��/bq��bȃ0w��ը$n�0_D!�d��@�j�����x�Q���y/!��Z?J��KC�h�:p�6E�$!��Ok��eʖj�$QJ�a��af!�D
qjJ(р��LS@0��Һc��'Ja|��O�U�9�'�F��n�n
+�!�D�O�X�pT	�%��ǭY�!򄝖���2Dk�\$(Cc\&}�!��	'���RC)Ս⹨�Gʴ�Py��ۅ~h�A���9RĀ�4/���yB`H:~8,��#=����d�Ȗ�yr�����C×aͺTa��_*�y�C�-$ܠ��o��%�&`��ybj��&�[FȔ;d.�X�H�+�y�$���T�?]xL��UmG��yRğ0Rf�%��E�br ��.@-�y�/��D���(b��*�����y'�;i�N%�C�@7��-d���hO����F7SBdt��gI�z�e�a Ց,!�:|�xcF�^�0Az��J�;m!�ƽ>�����#[REB�O�Df!�Y�'U|������AI���)A�$+!�A�s��@#�BO"|V� ]I!�䇔	H�Ӄ�\MbYk�f�$!�
 D* R��G">$��p���S�2�)�`~�17-*�UHa��"�����'!��j7��42����^F6�
�'mȥZ��
a��:�l�	����'�`�W��n�����*��~�C�'5�г�Eֻv�!zS��r����'c
0�$C�'���'��>�0|�
�'���`�7D����v"��5�d�	�'8�L�梟� ��"��'��e��',�0��"��~���0��#i%�y���� �ѱ�o�)aZ���G%q�v��q"O>3�"œb��-�΀��B��"O�� �Ƚv�$�r�]9L�v�Z "O�y�f�B�4��6�ֻl�>��"O���ƅ�u4�D�ƋwI80����?����CO�9�C�5�b�B5*ȿX�|��ȓ}��ԫ�� �4�x��AO�Z���ȓ3p~Lz�j�->�4�+W�S5J����8��]��c1N���!#�٭!nV)�ȓa�a��%8���2���fp�d��'� ��3b�t��q�U #jh��.�n�S�cH�m���KQ� $��&2�}��ՃDN� ���@ ����|"�1�%{ܽ�'텔h�2,�ȓY'���U�4���Al�R�\)�ȓ �lX�th�)i�È.�­��n��4RK�5�FH3t>�:�ȓ>� �d�
�����QF�lh�ȓa�Α��+B���FC�����'��=+��Z�s�l�H�	Z�}dŢ
�'݂MH6��3-���G�%r�,�h	�'��|����Nnx�r0����	�'�L�wnW3r6�B���T��'A�LCv�;�.݃�c�	O,��'�qp�l �~�ā�& �Q��5�
�'�4�s��N/)L��D�#A��a)
�'p ��*3j͸�%"3t�p	�'�Z�9���4rA�H��mG92)��'Y8 6�I#/_j��s�)��Hcj��x��i�����g*q`\h�˟�yR+%�h�'!�U��ia�M���yBI�T� m*�B����;S�ۡ�y���Tb0)�qOז�¹벌L��y2�W'$�l�j�Oؑ�PU��b��y����OM���G�=	(Z�ࣀ��y"O�S���i�!��^����U���!�O�x@S��I�p��3@�x�0e�"O���p���U�	9�-]�8�Je"Ofx	Pl�rZ��a, ����"O�|Ѣ��'��驅@�̊��"Od��e�J�T����Qo�>q����"O��x@�U�*�����.�&b���"O9���Шc^P�9D8����"O&m0D�G�"��
 ���IQp"Oܰ83nVNЅ�Y.[�n��2"O"삠l����L� Jг�"Orda�+[�'�{���"�x�"O)Q����'���#7��""O�����9R%�0R�~|��"O�(�9{<z��&C"�$�"OԘ{WF_�gy(�P���i��!R"O��R�@�#�Ҁ��d=�d�x4"O�ݑ�l+-����P�m=�ʠ"O:a`  D�0|r� ӏh*@�Г"Or4
�BI� O��['��=wdi�"O�9�����U,�y* �Y�Vt��k#"O����N�� B���sJ��"O�1A��J�o~�ƄR
6�̌��"O��{1+� lQj��s�D�\��ܻ�"O��0 �!B�x�XE�  ���°"O��0�lK�z6��8�G�<xR�: "O���-H�|k��dg�n��i�"Ox	0���?M� �����m��13%"O�9r�G�X�B-z匂�'���"O� !�C�3t��1�O�H�]:�"O0ɛb�U2�j��W�,I<8��"O���ލe�~�:ulv%�d�"OFݘd+�4(i��$�	�Z ��C�"O��p H��n�+��v�	�ǋ9�y���<�<���nޜtW�9�/;�y"FWtYn(�A�:6ذ�Q%Y7�y��T�H����n��4ȮA�э��yçL[r����
y�nU	Do�<�y�iI�aD�i��
�o�49� �J��y�E(kPy�!�7�2%s�c�3�y���6@DuU��j��c���y��L9}�}�ԆG�W<ܫ����yBg��H\���9JF�����yb�Sw�h�Fb�<��`�g��y� G�?9�֎H�5sh���P�y�[?" ��XY�zT���<�y"�
�9Ă����U?O�M��!��y�c)�U�] ��� ���C{^d��+P�bB���u��	�6)��g}��ȓ���"�/a��adm�V30%��3�>�����>1�<���1�q�ȓVd�����[=�,��wo�0�ȓ��]��0J^diks�u����ȓb��4�����%�D�I��ߢɮl�ȓgH����J ��#�j�a� ���3t2�,D!"V$8k ��}t"���<��,SD����0� D4�ȓ=�l�O��2�&��ƒ7i���ȓ8:���q�F @y!�w-�+d���	4��pA���p��H	&B&|���ȓBry�k�y\��(E��
p���u��ٙwg��'"d0���+��h�ȓC#VYj��
�~Q��rCM��K� @�ȓ!=��˴��G��Ы��?1�ņ�ʆ���J���.�%��4��4�ȓ����,�c���!������ ���fJ��4�U(.��\��M}b���+Kp����$%d1���iqe�ǆrT�Y��[�ӆ���*>��޴]�q�	�e�( ��z�B<���	sv�	�0a�g=!��j�>��C�(7rą#ю�:3Q�ȓY�Ȅɰ���uh��Cu�*TSz���M����&�3��#!))����r3��v��u�` �BU&/D�y��A��y:�GH82~,�
�) �e��44��ѧg"Q��իK�!�ȓ\c�A��MZ�>��1ra��Q��l�ȓB���ac$]�	���IFN��=V$�ȓ+Z����H��t���\����8�d�2��Y��ma�Br�0s"O�T�3*S�5�ã^QLĤH"O�9w̕�\ȅSB	� m( *O(ݢ�d�(A����Մ17�,+�'c���$�E7�R`[�!�'�&A��'�8q�oɆh���ТZ%U����'H��Q��"Ӳ�#H�($ �9 �'�آ�аN��x"O^��n��
�'P��)Z�BiI��C����b	�'BTT҃��<`&!B�EC`$p�'K�1��Y��b�P�-w��|��'B�}(�,	�9�Yh!��?���'h����T�N�vPrņ�5y
��� �u�0D� M�� BQ�[�8[l��""Oh���ȓ�,( ���3|Hb�"O���3� �	�3�' "pek�"O����Oէ/ x�G'A2&�("O�m�E�X���D&H����T"O!�E��Q�xu[��)�I�5"O�p� A�8B��`&ܜC�){�"O�`" ��
堡e��S��"�"O�3�ڎb'�i�$�[���(@"O�U97oĜ,�U��˓&B5c"Ob�05�;�ΰ�񃓽d�&]�5"O
�9�E�Ma�%#!$U��p�d"O�4+!(��f�{�#K��2V"O�=R�oD���飔I�P�d=�!"O�%@��'4RɊ2"��	���s"O]ҡf��~���$D���T�!c"O�����E���7M
?�}�"Ovu�T���s3L0~���x�"OP��VRv� �jA�k��Qy0"Ol�D�K1WJ*�H��+4�6-��"O��Kת"S�"FJ��v�ΠA�"O^)��B���~mp�� ɘm�a"O�l����s�m�V��,-Y"O��{�O�/H�s�P�~ق`�"O�3CJ�Yx��5 [:7�Ω��"Ob��0�
�}�vx��(ѕ��ݢ�"O�ղ�e� &�h��!���?�8��q"O���t,�6VKV�S�왊��}Q%"O���D �h{�j���j��P8�"Otty��BE�Dk�J&��b�"O�����b@�����?�H0�"OX�vO�.2*u���״pIz��"O�d C�_ bpV��L&eQ� ��"OD�k��5����.R*�"O��+��T�s�f���)êDG���"OXȳCᒤ#��Ӷ������*�"O0-����0pp��*W��"b⸁�"O4xI�ǘB�U�,F��zs"Oހx�ܪ�(�'�C�o.���"O�H�2�#1�$1���*iR�G�<	'
N-i��@��	'
 �q�n�<� O��#��@�*VrgD`ic��g�<I# X�d��@����K3@����Y�<pCL$:�M���N0�9+��W�<Q@�Ƙ>Y*@�+Ȃd,d C�DQ�<a�W�<�0���$��C��zDA�I�<�t��2=���녷wR���lOD�<���'�2�b@�F-p5��bsf�}�<��N�|�2񋲋�?���"��Fv�<I�+��@5`�:u W	}B���J�<��A�"UИ�0�8pVM
��D�<9�ѫB0��b,�28j �+��~�<��
��h���.hL�SQ�`�<���
�/C���sJԨ(�j��B�<)0kN�HO (A��%����AS�<��ٺc��ᢑ+�#S���(��HO�<�B��]�E��$&c��a�hf�<q#��}�,f�7�~M@f��W�<�LQ�D6=*�m
�@\X�vny�<�:h2�T������9��<i�!��I�i�8����ߐt�p�3ԣ�x�!��L9h��3\�\�r�Y��n�!�S�d��u/۝j�r���Q�i�!�$a�a��,tX0`�~�!�� ��Q J<��2��	�l�B"O��v���mG~m���0M��!Ya"O҄���	�,�)�F�=�~���"O���*�"b��<8�۝h8��"OEAͲ���+Q��4Y�Ey""O�@�Q�GXh��c�.1x�1�"OԠӤk�x�-ђo�	@b 9"Ox�B�^�L�:D#��T�/ű"O.�����(Ya��M��q��"O�yJ�+Θ~ >�rӎR�{�hg"O�ࣷ��+0����˓�s�a�'{��C$�ǺP����M8zߐ��'��TX��ًDQ֔�s
��&V����'a�ebѦ]�d�ִys��"��i�'\�iy�O3�B�	ѓj�H��'���hE��*E���3Č�a�"��
�'����S�ɣ1%2�:'�Wzΐ�
�'�(�fi 3h$C��I����'�Bu�Эژ� ��d�LSBn%��',h���O+
�$�z��,u�q�	�'���Qg �'%����F+m��L��'�J��)��F��a���s�`A�'�p<p��H̒��#Z$��]��'���SQ�Y�DV��r�m5��'�  )��եC�.y`����&�ݺ�'80�# �@��dG���=��'��YPb  ��|у��	�yC�'~������(F*�'��-�X�r�'�L�ӔɄ���1#�Ś(�X-k
�'z� �dŹ}|���1��4��'�zmA��3[���(��$��I�
�'��]��ŝ*]b��d-���I�	�'Pi�+�w5��pdc
5�t��'�L�����j��qz�69��!��'b�!�Qȟ�1u�C�+×)L�� �'φ,���"��y�(y!(h��'�D��fdj��U�s4�̣�'��x�MM$���pUȔ�:��!
�'��䂢iN�q�hq�Sl��㮤��'��c�i�7���#A����'!�[�U�8p����(�:dh��
�'��8��H6}n���� B�0/$�(
�'��=�f��L@@���=-�V�q
�'Xb�p`AG0r�(j��U/"�z�B�'a@�B��P�$�����/*�b
�'g�,�*Z�g����LH�#�j1��' �0��^>y7N��	����@�'`���/���9CW�Fq*	A�'if ҠO�=e��9��g�=<�&�;�'ޔl�@��?�pH�5��
9C��`�'a IA��L��@D+u�<���
�'�0���Q&u:w倲9��s
�'~f1"�Tk�ea�gȲAݬ�0�'��@�1�S(^�A!R&�3��Y3
�'� -B��!vQ&̐B�%"�X
�'�x�'�7<୻����Ot��
�'7`��$ ͗R�.����ŽF����	�'c��aM�66@����G�/8�!:	�'���H�&6=��:�Jȅ7���H�'�9�Q��4aN&�Q��_8*�����'�ĕ���#g>��$h["`�4�'�V���X�L�5���&ȥ8�'�p�B�DJ�ȹ�\<�݃`��{�<�F�W�w�A"�o�*� h���n�<� ��A�\�/#����ƀ#t�V(x6"O������-P�-Y0U�gT긠�"O�i�&�ϕ]�Dm"��M1^?Pٰ"OR�y�	�@f�� S+g*���"O �1ʊ,~ƾ�Xtأ3��!�"Oji҃�+2j���qbϐ1�H��"O��BbZ�����߮���"Of�2��E	�F@dǂa%"O��2eK�}ޱ���Q��V��"O6�:"l�&0���qG��n�dAB"ON�#�Ⱥl�~}s��#Ti|бr"O츑�@_�F IX�K=d�����"O�)c�!h<|]�w)\�L��a�f"O�}��L�<�<��GۍQ�
0a�"OhɲC��}h��H�ѯ%��S "O@r6靻zZ�I���I�x��"O����a�&��Z�)�����"O���BY�{
�4��.D#j��A��"OtA1��9:����G��Ez���7"Od�ir��"@Ȃ��Xit%d"O�1��ڿ.��<i��	%]@��"OT���Hm�2�RQ��
yR	J�"OtԻ�$���hq��.�6ɴ�6"O��q�fL�H�8Ej�o_�Ld!R%"OB��ѰR���Bn�T�At"O��D�(O+4b�MD^��	�"O���A�lW~y�3�
D��9��"O LC�`Ҡkt}kpl��\�z���"O�q0��ßH���*F̏��<c�"O
uk#�p�΍ZAl��o�DX3�"O����l��X2-BCk�o|p"O�"��H�3�xؖ�ߣOr�('"O:��a�] f���*�N���	�"O �#�0u���N�#�`��"O<��Š�
*r0R��M>L�\2"OVt��씅A�l=ZS`ʦ�޽Sw"O��ä�NNq�TQ��I�����"O`HO��U�S�6� ��"OD P��2��풤M�"��=X4��\��I9:�X}ƮۀnmD<�@�P�{�nC�!< �X�4K^�����Ȑ�1�6C�R�� ��$bk�E��2P���D7�0�&�$V���N�(tΨ��2D���Xa����ѮG�CnD���H-D�ds�J�A2X�K0e����/.D��c Ǆpgxu���d�
ٚGH�O�B�I�{��(!a[q頩2B	'i��C�1:1��&K�)Ȧ���m�/J6tC�6J�I�kA7>@|�Bu��(K 0���>�-[&N��р�,�F��CvfDF�<qVł6���*��L	Z�xg(�f�<I�o��m�A�3*�l��Rl�d��hO1���x��@ B܃��=� 8�i+#=E��4I����5t��ز! 	f��'����)�|BD��d?Ry�6)F���d*�<Q�)�O�����
JP�x"c�=�:a�N�M�ax��I4)�T��BN*G\�n�$5�NB�	��m���{ax8S�U�[p>"?�4L�Q>��jЋ:��A�ą�:M��Qg� T�`s ����@�qCa˦37��""Od˄#�%�� B*�@D�Q��"O$aM��eԚ�q4*O�=6t�s��D&lOJ�35,�*�.�Bj�G�|i���������S�
�;!FP�/�X��2-Y&oL���D~�� v��e��'��\)Kݴq&60He"O���c��0PJ���w���-��5���	g�OY�ܠreL�6Y�:�տo�24��'��|І��"g>ZL�#i�!l�T�	�'-<h$N¸��U
��\�Mo`�	�'A؜3��L�4U#!��OF� �Ǔ�HOvQ�kb���2�`[,��DR��'��	�2��|Ze��UfD�j!��6��C�	�Wr�y��h51ҸQ�.�B��#>A���$d����Ƃ2.~�$��.�I��C�I �h��#eQb��$���k_��IJ��h�9�.�?�ɓw�F@DƁ�""Otp��c�CِE�d�;4;��1#�>�	�0�h����aKD,LSm��ȓu,0����K�qy�D˔*��q΄��ȓ.�� {&Eϸ��e�DF]{k� �ȓi��Dۂ银Ft�[�lυ-�v���'3���"+S3��� ����+��<X�' ��r���;fKXU�&'H&&�Vai�'9&A�vL�:Z�.x6�S4 H!��'�ў"~��2�2]����?�$Hٗ`�j�<�1`ϋziD�0#蛰j��!a�+�]�<y�f�(����/��A��	V�'�Q?	�t�K�58���Q!6��#Wn&D��Ҡ�C�E���;��>�H���i�O7�<�S�O��U��Ty�Ić��*�R#c"O������N ����	�]6��7\�����8t�}�sd�
�	��'Ľ: ��$d�d�3Y@�*���䎊^��d�>D��H�kڽ{�`Ԁ�],��qa.<�D��d/>�N3"˼V�� E�A8�!�<OM����D׺d�jq����9��xR�K�'�"d9���9��Ic&㇫y����'	Z�a7�֝2%���Es��z�'L�'��)�!�-ؠ���1����<�����W�DS�dq��� �L�x���?���CA����K-	��\�BD��a��KF�7����$Uv�ڡ*�7�K�.M�>ݺǪ>�S��y⮝�4�����.cY�tB$�
��y“.���H֢]{�8 T���x��'/�S��)5�{��A���*�'�(@���^lDb�d��~of�a�'��qz����K��i�T ͖E��e!��)��<9��H��H�OW�3���١�	a�'�ўʧP̱sS���&�ؙ ����4͓��'�ay�Ē�^e� (���61��U!ӎ��yR��-fi~�Z� O%ㄘ��K�y�F:;��l(�KT�8�Hr��F����hO���d�E�Po��P" h�m��r"O,����N��e*", ϞI"O~�c���6U�&��ɅR���[��Io�OH@�{�ėEW��p�ɑ�D�<�Q��d:Or9Bo��rT��A-�^��`k�"O�Hr �2��8cpΘz��8 �"O��H�.�A�������y2`�UP�p�vOǋF7�`�����y�`F;�v�`��"�RH��yR��24��9DM��Bw�$c��T��yrg�#BZ�(��ӭ�@�@A�8�yBd�<G�p$&��
�J�;Ӯ���y'Z%V��2���|���,¡�yB�	����VM4&�����^��hO����W��P9�c@�2rES!DG�	�!�āi�h���	�*jZ���N�{�!�� >� c!Z-A[,��#f�8۔ȺR"O� P2f�&��A�E�"����q"O��K����3C��PZ7%�\5SОx��)�Qj��S �F�*ĺ��%RN�C�	�|�c�IH�a�$@�����x�B�I
N���i����'��%	�`�.lY�B�	\��m�7e�p��J�k_�l1`B�++�+��B{���� +_6B�I�w
�2�G ά�"��8.���s"O��m�t�@����R�O��Ec�'	���k����7X(]��FQ8�H�C	5}24O���D˝�Z���Q		�d�ZrK��N��	"FS�I1�H��7�`��)peC7�P�b�O^�\S"On���B�}�%�1�G�5��m���'D�ꓑM� ����'�t4�gI:|pN�)�!]�>}��T��f�6�FԣcH�0v�Dp�@G��'!��Iz�`C�Nӝw�:��"hj��rq�6O0�Iu?��'&Lu#��ݠ-��@�U��iM2�Xw�P*r�!�L3x��S��e-J�9�BƸ6��|���?�J��S/U�c>�$Y�3�����:+��A�c�Om!�D���N��n�,3Jy�@�ء	X���,E{��D���
��Α����{ŧ���y�:$�x`�r���4�D�	�򄬟����-G:��#Q�]�,czy�Ơ͸w�>��d�����q��i�mȶ#b����1D�䲤"ԅ&_A��i\�
��%`��/D� h�O��3)�0id@���U�V%-D�A%��/	j� ��	�7�E��.D�XN�.��Y��H*lٺ�A D�@cӣ"CQJ�{�`\<#����Q�<��s� fBR���9�s(��?OR���Ig~b �%FM�)p��٢_�.�!i�4�y�HS�u��P�%)�>Q����fn�1�yBJ��D)2@��I�f50Ƭ�y��B=z)["LӲCr@�B�T��y��
�j��@#3U�p�@� ��y���)�qul�;{��3��X�y�㖢��-`RbɌ�H[6�K��y�,و Z�y�U�ժ.N�Ҵd��yR��?QnxI$D�)�p(�M�=�yb�R����#�hO���ge�,�y�-�?���brEˋ0,�G�Y�ȓn��h�
5	��qPgߍ[J���ȓd�X�[ Q1]~�PCB�<y���
b��T �'X)s�
�!e��e�<YT� �VL��Ȩ,I�E��v�<�bM�%w� ��!��.��YF@�p�<��(>,x ��Ҝ1k�k�<YѰԑa�At�B[$VX�LC�I#e��Qk���8f�*��3@�/�B�Iu�!0�
�s�l�Ā
=�B�ɤ	��xsSdM7C����7K�B�	8hľY�U�ߨ������΁W�B�	��d���{J�`X�lX;��C�	"AF�����$⨤��M̹<�B��TYd	�)ޮ<��L�F�I���C�!C�8���h �)\���� B�IcԽI�ă��N�S����k2
B�	(:�)1UeأZ�jM��=2��C�	�~8q�E�"@	0��eB�L̶C䉗t���J@�F0 �����b�C䉐M�,��E�d'��I��͔v�C�ɏ�J�����8��,��lׯ��C�I�K
f��7M~�f�0�I6W]PC�)� �� �V�,���JS-A_�M� "O<����l�0A!����(�H���"Or\`�E�.��j��	�"�*F�#�Ԣ�␛T�^�	�A��Q�6�ɑ;���'$_	b��`���+2YC�Iq&��$1z1�% QK2�B�ɦ6F��@v��q��\��K/�dB��%�h|��̛{��!��]��C�I�4��M���ȣi8�),Цs �C��BbL�@�M"Ǯ�p���<l�C䉢%���q,HG��9�bT%K�PC�I/0��Pz��Z��N�i�N'8�C�	�}�$Q&�t��f�ѕv��B�>Uq��i��i�^���j�;.~�C�	�l�t�gk]2l�\D S�]�4a�B�ɴn�L�HgA��<`��D =:rB�IR'�m�lB�	�(�.Ao�|B��+*ɨ]�� Z��������5�C�	.)�у�.%��y�gi� Iq�B�	�j�R4��f��t�d!7��i)�B�Oe"�i��	?b���Q�צ,��C�	>�Z� ��B?#����3s��C��C�A�Ƒ��̂#MFj�@C��;z��	����OK�ݡ��ĸ��C�.c�y�HU�Ybb�[�kC�Z�C�()XX(@B�%�z�s��́l��C��5��a��}�"]c��ͻX��B����9`#H|�y�J�;FB��0g�z���#J-B�lk�cȵ8B�ɏ/�p�&k:̠�IՈF�#(B�ɐn���k�M�x��'9�B�	!^�c�/_�a2������ �B�g��11�KJ8|��L۱�ܧd^�B�ɛP"����I6=g���E(�x��B�	�Y�x���F��h�Q��k�C�	�f]���%!�� SbG7B�9Nx�i1E�B�s	΄�	Q(2�C��6: 4e0΄�S �$�!�N���C��F���J /Y�^=r��+B�" �洲���p�(�+���O( B�I�8(��f��12�H�dϑc��B�I'`�*4+uj�|��H�7L؟H�B� 	�FeH���AR�8ХH!@~B�ɋZ).��ō31Y�}�B��`�>B䉪cBQ&��!�`I[!n�u�C䉩r�����%A#Fy�7G�m0B�	8y�v,��L�8����;
�C��.	<(��@b�	�R����L9��C�I�̡B�F� qV�Q *�3Jc�B�I2LOZ<(D+]�Y�A�4n��L>�B�ɘ	�\՛7⁶p�M��ʺZ��C�	&~O��"#�-g)�	����IR�C��W.�*�ʰ*،�SFMD^4�C�	�8��!��f���~�P�D�?����D�;sɓ�%;��4�F$�zT-������x�F��7~=����n��8�����OV�J!C��
�b?5C�n\.-`�����	����&/D�T�d��! wx9�"�zW��� �n� �@ *���g�>E� JcB0X�pD4�d�����(�yB�܇1Jh"N�&�8����/��DD�YE�Y����p<a�G,�Z�x�䙓�.%y�AW��4�P��M1v��K]��6E��DJ45���H��D[�QL��ui�X���Ss'J�Z>�`�F���:Q� �IK$3�B,�R`�?;־0D�1%!�d^�^J�}I�D�>��S����0)�D�@h�c��9��)�g�? ��C�a�`2P��DW�+���9q"OB}ғ@ֻ��a��:~��xʔ�����p�X	Ѵ�'�p���K��|:�E�
��DB�tu(9p�+L&9��ء�GC$98lq�j��{(Ļ�-��*w'F!>�ҁz �4�n��H*�ruj ʃ��(��O�8��SmIl�ՑpD6N�]8�'6V��`��'zVI���ڡ���ҮO<٣��渧H�>�8�i_&!�٘5"ي\��
"O�!�4����[�,�y�%Y Y�!�d�:	���c.M5i<��q���!���1���w�U.�dQ��ȓ'VJ!�B��a�䕡h�*��R��;�qOR`�S�U��0<���dG����%'O��#��h<�	X�[���q3B8&*R�qe�(Z�A��j^���?ɕ�X�\��-r�Thv@-�/�g�'�&pڵ��]��1(+iw�O�~���ش m(Q�b� )�(�i	�'�@�wd�#H�j �bD��2:��OD�sB,)��m2*L0Y��s�?�I���pAb%c��(�S�K�v�<B�	?:��m)peݤk2���p�U�28䳣�Y Q�Q�F�J��@�K#C�Q� ��$��It��iɡO�L����<|O�ʄ�U���5�� �k li[�eى9�rիЍ){J�ئ"ַİ?�t�ƐU�vd�T��qت���LQM��Ӓ�1i"�*Ũ)G;����9Q#@ 
�2[Āܗon���"OV�X�+�H�B�1PĆD���C�� �|�D��TD$I�0F�>�I2e��q�Uc ɺ�0>rH��"OH��-�|U��zQ���R`z���4kވ���%ٯb`����ŧd������yAh�9+n�5@�,O�T��{���eB�	��9s�dK�6�L0�6�X�v��M����2%K����Q�,u�0{@J@��lH�JU�O��O\��	�"_��i����)�@Iɰ�5R�&óa��5K��V�.qp]"�ȓ��!��+`X�š���lW�Q�OY�,�ָ
��
:F��&e�%�h��.�H[ػ���6OE�)��]�'!��25�
���
�G&��q5A�f�=c�@�<'��I4��W �Zv�O��FzBR�"�Ő0l��D������=i�����AR���l� ��	J��-��jih�g�$�Pt��'�����	�-�t���&T��t4��"V�c����ѭ�Y&��S)L�,b��O���V�#]3���M�q�h��'��	���Q��d�h���0 (���x�� �F�I��j�J���|��wQ���!�ڃ͂�ˀ(����'" }�@�C�<����Z"^����Q�^ N Q�N�9�u1�%���U�$�B��:��P5��`�a��=�����@[2@����H�<az�H�-چ��@�M�|�����V�V�a}BE�<Q��⑆J�9��H*���'�D��2mJ�z� E1�cM�U|8i�J~�N�l�\�1�Ɔl+�A:��ڢ�y�`X?d�.L!E��szzPA��^�Q��k�M�S�����F�%��s�AIo�p,FY��ɘ�$�:� &�!D�D;U̎T���@��@�MJ*�`�дR��xI���%�|��D��$<�3ړ[�*�R��؋7�ԕ2'�R7y�����&z~���/��`���ֈ��Q2�G�Ig�PЂOp�Ѡ���A��pR�;"��`�I��y�ʦ'�1�&�YC!��*r�e	��TΑ�7"OT0�q�Q��䈣��z+��ID�O4��Ħ�[x�KI��}Z�*\�u3�<�u�������	R�<������X(��'�8x�p�+�OVO���r�JѺ�H߭�0<�1$HG��pI^;Bi�&*o������F�%o6��� �!xֺ�
T/�J��<ʇi��:!��1GH�h��
N����8�Q�c�@
e��P���]���b)�z'�a�a= {!��!� ٙS�X�\ܥ[�+��.����{���n�B~�-�9��~�ug��x*j1�B��^�Zfai�<��i±+��<#�AQ�<�~�Z�&Ue?����	��m�k�~B�Q����H�@k|��A��d��,*����!�,Y��+�-L%#�\m�$i�1$����m`.��'Kw�-�,�Q���v�Q%D�B�x�dP�,d%��=�O�R��H:|�d)� ��)f�[R� ��%(W����wZ�`U�m(��?�D��ƯH*�d�0@.�0��Ez��͞K'v`�'��Y7X8�~�d@K+0	>T���̀A�-9p'�Q�<��kV-&���@�U�&!h�P���6(�b�Br랪�L�(bB�\mG���{W��q���c	��<�vL��}9����d�=1��BL�F���#ω+��i ڑwQ:<�$��OF{"�V(��j�9w��-
�����=y7�"r]P �����-)�����pi&��z��<`0�,9g���1�'>�d�!��/�<�c��/'����}��("��p�F=_�(���ؿj���BB�"~�Q,@�E�D �$�� �\�!+Q~h<�GK�=\��'A� =�.�CGV�y����u'��x�8���#?phՑ�4y��1��|�n����C�KN��������i.D���`$_ H���@�P�b��h2�JF���O8
�9Aƫ��&��� �_"M�����Q���S&��ȷ�� Q����&��$��Gz�ڄ�#4BT��&B�d�Y�`G�m��d;l��kдq�F���O�^ ��ɋHl�qQ$ϓS�x
S�ҝrD>㞌��O�%�Jd*c쉈$v��
� ��Ms��	Og�}k!j�|b6f�
H�1v�6��x��T 2��C*د'kִ�e˷#�V5Bs��=���"FL9M_�d+���"7�٩j�|ʢhށYt� �8T`�X�Ȇ+v�:�K��<D�4��5sv��� ��(��=0e[���_"<PRH�0[��5�S@7v|�����BC�I�w����	�$n�2���l��.-f���[ :n #C�
Z�.�)򭗽:F0���lI�Qq
�@r̜98�t��#dS
Lΐ�%' �0=�&`�I���b%i�8�� w�Kw�+ �Iӂ��(�#�K%G�X�J?�rSŏ�@CDy�EM[$��Ѳe6D�T�A˚�	>��HҸ.��td(ȅ�u�G�1�d 4���O*�a������h*n�5��"O| �pj�(�v�����ow��f�G@?Q�#�n�Xm��$G0���ɒ(�2����Kߘ�C"B�;Fz����AH���ONl��p�@��U�l@��B�2��l��'���P�ۅ7���a��=ר�����o�ܢ����L�kM�Q�d�(St���Oϭ�y�� 1�d�:�k��I.��J����yr�խa�v�����>G}�dY�(��y�O�%.��]�4~z	 '�'�yR"��v�ҁC�Ñg)�h(@Ł��yr"A�M��������]&�8rg�4�yr`�
8���I�8!TC�b���y�\��}�VF�'0~��$5�y2���t,X�!Y�.&��� D��yB�/:�8 r�NRB8��pd;�y�\V t5[����<z�@�y�7<��@�5���d�x/D�����ǚ9��b�"UZ@ ��5D��s��& =�}�`��4!�ir�2D���S��s2����OV�'�<��PE0D�|����%���Do�v�H�7 D�h���Y�t*���D�T9ZL��"��3D���ꘃf
Lg�ZSi˷�;D�H��d�<D8�􀒥�t�̰�H9D����d+�@��C!P $�q�7D�8S'LS)C7��Y�g&�H�j��?D������7v�\��)Hc
��Ȅ;D�$1�B$�hxQ`�0Y�X�'9�C䉵u�L�P#��>a��S�D�4Q^B�I(m��)s�M�섈�
�Y�B�	�fɰ��3U���M6b�C�ɵ �mc%.��B:\Ȁ M�B��C�	��~`;B�ͻ|e�EA2+��L�C�	�E�>p�R�Y�I$���0"o�B�	�i�&�EiZ2,���� '�B䉶c��k0��*~.D��N��6�0B�	�*�-��@F(�8�u+W8�@C�	�P��DV�sn�a��ۖ-�rB�I�P�:$�&<�A:@?8�BB�)� �1@��#!�6a�ǈɜv�B��`"O~���y�������PZ(�(�"Od�&C�mo��S$nl�\�"Ob%rv�˵OU 'hR�[�,4yg"O�T`�A�3v\���R)c��@�"OD����?E�Vc�����t�@"O��	 �����H*%�W�C��qa�"O̽�q��4~L�	�眷m|� b"O8��F�Ly�I�+��?bz)$"O�����s�(�*�i��LP���"O��P����>�S�fƐ&x��PF"O�r�̥7$2���e#b� �@"Ox`cG���k]���DZ�EaFY@�"OzL����:k@<9S�E�Tl�"Oưz�#�0T��$b�CN�EK��J`"OTl	��
~=�wC[=3 v�c�"Oܪq&ʒ]Q�xi���#a 1"O�|��Q�~��X���:G)���"Op܈`OQ}ZB|s�`�;+����"O(�aB�Ӳ[���3w.�,�t��"ONГ���:{h���Q	e�@��`"O�<0��;�A��-�)X��"O����@_�h�L��I�`g )(�"O�!{�b�o�z���j@J�9�"O�|q��,����c��,�F�S5"O��˃�� �(�h���)�Z��$"O�������d��!̀lҡ��"O^9(�� X��0FT?UB���"O�E���<���s�S�p�i(2"O��;��ŉF�����O
���7"Ox=�$mݞ�*���P�;�z�xW"O��HW��tQuAႁ	�
�"ONyh��
<.%��Q�k��"Xa�"OnQH藩{�U�+Wm�r�X�"O�<pD'��]��}BI�)H���&"O����I�R�0��˗}NxI"S"O@����*͸WnH)|V�D*�"OX�䈐9Qy��Rt-g��)"O,͊3J�:��xږ-��Di<q�"O���o��A�f��T��FtA�"OmՄɠ!��=8�]�l�49�f"O�$���Ӳu�ĭ�2�R�|$��"O ��mN�$���%ظ}�"O��1�� +.��@��:~$Ո$"O���d��LD�U�*6��0"OVcW×?�Б��Cʙ?"�{'"O�e��'@@�+����(�:�yB��za�@Eѽ6�xD0d=�y�bD�?��ڣ!��6��,j`��yBo��{�4��D��r�z`d�,�y��y؁pb58���3w'� �y-�!�8��#L<��3��N��y�ܢ^�V�p	N�F'��&��y/�w�����M�RY�.ɠ�y��"֤�;����O��
`&�:�y�+��h���ꉲC���H��"�yb��$uE������(���m��?)��H�N�qώd1p�.� 9JB�$4�Ѓ�9*�@˦D�����-5�X㨌{1 ���Om�Tz �� J*�}3�-Xj�H��'r�`��a��2�B�ˌ#_eXyq�'2����*7��<�O?�����"7�U��/1B��*w�/D��	���C.�`ˡfW[��؁�J-?�փͬ-��сCe5O(�(�B-lz��hFd��\f(ك�'�����D�� *q�6d�P�V�Ge9p�&���DR�Px(�@�J-����:*�cë
��O�Z���c>��B����R	(�S��2�<S7��y2"�
Ʈ��0�Ͼ"N4]Y�C��yBLJ��{��SU���/K(d2�B�	SRX��l�'P��B�	���S�BVؐ��K�Xb�2��q�!���*����W��-Ȑ#�,FW��t�MT�a~��H+m�2�*�+̒F�6��%�#p
�hS���i��(��@��	����Pt���E}Db�$Y�`�ɗ29��ġQ�L'Z,�d�\F!�䑅3��h
�f�P R�]���GQ4=;��铿q`l0�Lׄ)����,��c�B䉝*���{��s��aq�ܤQͶB�	2j�<,C�E�Dh�հ��G�QvnB�	��$P7�H�+p�
����Z�C�I0a'(�T!�<!�L����8>n��Tڧ�6�axo�*.�.!�G�Gz��=g���x/«,�d�z��-����ǂ�E���2��fx����7T�L�u��+2ޝ���;�(O<���C$7V�T�#�3)0��T��ʙ �@��٬dڨ� g"Oh���+�$��BS�ht�p�y�PX�"�#:' ́p�Ǧ#~Γ~ �=���42�P0@����a:إ��8�������Qr�����ԩSj
_=fya嗿ml� �0���?�>Y�k�,H��8�
��&Ҷ#'Y���HBm3z��q�+�/}�6ِ�`��?l ��E��_�.���)R�Ka�(�`��L��)����A�`�
��'��P=s�����R(h�'>uk����x{��:6��+�u��ݯ�yb��$��z5I��}����M�p��e 2��/T����'iY�2�t���O�9B� �*���1�RG���*"O^(��m�FC~<�#'P�r���;Q��2I��1�dƐ=u��+H�0����Q�q�μ���\3V�BԡJ��y=�{���>���ڷѠs�l(h�a��34a!���U���(�aƃ����Z�)c��!Ƅ�T>Q͘>�O�[���4GU�l9�	N�t:$�:J4���+�,)q.�d�XQ���U�<�r�׺'�����@k꤈���*r�Sr_;�?	�&j�bա��9�65)��ڸ=�X�T���d�p"OR����&�^��E.	k��X	S�E8zY��Z�U�X���f�̔3R��ENl�'� h�`j
��Tpwm�*E���H�vӺ��+ˉw�h��偖_�JKT��{j��Bs�	5]H�%�U�G�<����!`YІAY1A ��Yp�,��O���|IԢ�M�3a�{ H����5j{>Y@�F�J��e�R�	s�!�$�<�&ذ���U�|,7`�+uh4�s��� !Q�n�t���R�Ow�ڿ"H��۰"�E}���V�ho!���4��T��V�]�i��#~��`�	H�v���qR0 ���O��HDz򈑎~�f� ��T�1�t��#Ԗ��=	���91VMɰȑ�P���㜏:��=�"㈗Y��B%�m7�٘�I?�O%XXkN\W2�����fV�O��i�,
!g��J8:�>xJ�˛���IH�a�D�a��/-`Re8'�SGX!�o� ��ǈ�D,�z�"JzqРFOnx�\pD�EE�5�T�7��;��(���V�'Q4����X�<�
-(��I`�E��@uVD�WOH~��Ԃ��Z��9$������g�'G�e�m� >'�="�jC�"Z]���6�	�	�P�! �	X���Ș.;�|vԐ !���.�(��f��Li�nX�5Q��b�"��Wq4�H6�	.#n��xЋN'Q�N�8t
¤*�!��P1'1���dۢAd8�ʕ�B�}���M�&�1BcI���)�'"}�q���^~��"DCL�n���=`�0����x*T1���U92l��OP�Zt'ƨtj��^E^ �ӷu9|��F�/q�=��Iu�h=)�L�9{�� n��vUv���JZ1{W䅓wO�`�O��</�9��$�5e3����I g�����ߒ,N1��\���j>��!qb�N�!��"OhTKA!�e�T�� ��i�R��Ў�$ ) $�"}�W�T,"a�)�WO��3��Z�O�!�� hx�2�Чc���F)� ߘ�ڰ�|RiTݜ����Z���4�� �gI	�fz����'$ҀxC�<�n�o���@�')��@�DH�&��X橗)t�<E��'F,���%��U�L�v��'�FUZ j�"[�p��D�i�\Y�'{N�2�!"j6h�ᓞm�X�(�'�,�y&��1+����C��gm^\i�'zr�{k�$H��mX���Q����'�� �P�m7T٩#bM�M#����'�Li�d-U"Mt�	c��410&��=C�
402$����S�I��&ƭ!'&�q^�1�ȓ.�m+%"�!�Xy�"ٗ!�-�>A֥	vβx����ED	���!�\9X� ""�*9Mn	�.V�a��%��'���P*M�pęa�[	J9fq2S��
����L��n��] t�U's:����y�hʡj�,�-	�.����!D�x���F�kd��xTŗ-J��:�ς�[�n,�FF��AZlź�O����M����&>7M�������9}���k!/�\{�zB�_65�B�ѣW�<�1��7 '����.~�HJ@�V}"Ԛr�]��&����<Q�A�\�%}(�`�D#L�@�]���k>��6퇳!�� �J�G=�RQ��"�$�*׭R(�B�O<��!1�(����fN�/{zq�����']���B�5>/ҝ;����ѝw\���� #/C쨛�f e�h�#�',`�b �L�G� � *��['~<�B+��P�.!��'
p��V��F�O

4�o�g\�����|�|a2�'��i�7ß.\��͓z4-�G�N
%�r��ek�+J��-�'H�� K&�0=	ԩӠ�)J�@�P��x-M�*��U���'Ψ�dʂJ�M0νK�@\ Su�DyD"O~@��,�?=<V=K.�u~Y�Ө��(����=a���Oƕ� Y�"`
�ps�W{PI�"O�ya��GR���A"Q�=���"O|���vx$4��ᘹg�(��"O��U��D PU;���;!�@AC�"OZ���X�|��%�3�ʇe�D�"O�B#-�%�\����=nE�4��"O@)��쎉=h�(�&��3��S�"OpP���J�0��`�%�%=0��Е"O`y˧O�?���Ō�֨ɢ"O�y:��M�A�����2,�y"O��K*wv4ؑIR>A�1"O4��c��5bP�$a�#C
8���"O\E���'n�H��OA�^�܉%"O>��拍	 &}*�����* @"OZP��Ċ�
^ݱC�	�y��Q�S"O(0[$L��nd�A��3Ӹ�X0"O���W��6���D�l�&�Q"O�9�a����y�E�Z�jC"O��pMF����C��/|��r0"Oj,��Ό�=��2�*֡u0�S"Ot}a�,���C�
�2S��m�"O�̳1#�Hɰ%��k��b"O4h����U
�|��Ķ<��D"OH����P�OڰYxwϴYm�@�f"O*�Z���p�h�R�R;f�ܤ��"O�):��O�I�Xer�� �=�f�	"Od���fɔ�t�1�ᄑz��m#�"Oc�®-�\J� K�>y,!sV"Ob���ė�@<�֊�@|�TC�"O�D��%E�A(��jI��	Q��h�"OD9J�5�Y���]?�,��"O�d ���(I�Y��ˏ6q~�j�"O�����N�j.�b�_=n���"O���!a�j<����,c>�d"O������@��R�۠A��H��"O� ���$-�+[���;e�M��`J�"O� ��柨@�a�j�i1����"O�`ֈ���pZ�^��I�d"O�] �B��˖��3�7.�	�"O��3wi_	H�j�)s�٥iX(]k�"Ob�B�Ղe�:a��� X�M�T"Oz���e�2j^�LWH��&ѷP�!�$�qH6��Fc�$98�42WE��!��"E��TpD-A<yS�*��!�ӵ�\�!k��d!jx��*�	;�!򤟋aN 8��j�Q- i��FF�[����,ȇ �D���Jģ*���P�+|�tɳe;��=BB��fxTTA�=D�����J7w�����>UV��=D�l������l��%L�B��s@<D�P�ъR�k�
�����cX�m8D��A�â���y�+�]�PX��7D��ZΌ"9��z�bDv�����*4D���C_1-:V��ՃޯwZ�TY"N2D�؃�+��5��Ж�ɱ(�� i@5D�؉u;l�1��Ҿ6'<���"3D�a0�Z >~���or�q��K$D�$���X�t��!�KK�r[�l+��/D�$�` �
x�v�zv懪B>���!h#D��P�.' =�2G�:nr��"�?D�8�!%�8>���k�G��2����:D��ٳ�Х1B���G�O�؄��K.D��S䝏l�l@�Mð|��x3��-D�z'��8�@sG�.����׭�ON��1���M���:?�O�����n<�uJ�*}��x�Ӂ=[�����T�1�6�ڷ͇>
ջ].�����0|Z��"x�kf!ϡd[�}Ð�� u	N%��	1f�J�E����	Z�������n�V]R!B$>4��2v�W�?�-i�U2!E �K# �c�z!����o>Y��M֢H��R֬��yX`agL�[�f)����ę���%��vǶ��	C�T��j�+�� O�l;Rj�`g2PB��/f����$�6#�xf�~����c�8eR5XE�st��cC �-;�CUUuX��!g��87��
�'Vp �#q�ņ)i�� Vk_qQ�����\h�����.MFD{'���P�%�?�x��tdD1��������2���o�1WN����Ц%�!�D@�&�V2U��9���f���!��or"ٲ�o�4W�M���H�&�!��ĵh�t81�	ȧ
@,x�$��V!��O�"�b%���N8l%�Yp�LN�-&!�ϭvt��3B=jY07��4Q~!��hb�����!O��pp��l�!��|}����Ŏ9���SB�.0!�dU�n�^%�7ᑃ��1B
�I !����Z�뤄Ł ��M��gG�m!��;s"��5l�!�q`$Ǟ�4!��*�jmZ֌��X�U�c��R�!�d�>&�2QF��&��zGhVF�!�DՆ�VZ�Z�B,��
��`r%�ȓw|t0��	��͊��!^i���ȓ]L�E�v�Z:_b��,�$!��^Y��h� ��,���K�ImRE�ȓ7�D��
��
��uK���Q%(8�ȓxb�E_�D�E�
A�豅�"�p�˂�^�YCj��bcQ$z H�ȓe��PCV$���҇G_+m�����g���#��!k�<��
��n>N��ȓ$�{��Q�TQ`��֬��t�vU��Z�:����0�"�ʅjG�/�Y��s5�L�3�ay���t���pz��ȓ�@)2�G�RD��)�!��Fʨ�ȓkȤ���#ܿ,7v-a���mT0��ȓ�<���*'���V�	-ɴ���S�? rڦ���Q1H��GGNp1�"O�i05���X��$��G��Z���"O��BG,X��9ڦ&
�/3VI�"O`�;`�(>�\<`e��,=+����"O����e'�3��f��U!�"O&E��W�%���IC	�Xu�Ż�"Of���UHp䈢#��HB 5"O茻��+*8��y��$
��V"O� !D ��0�j�cs�9t!faڦ"ODa�� �'��-bQM��Z�Hv"Oh���ʐ9Z| qgLy|���"O���VH��� ���Y�R�͈@"Od<br���Td��n�s�(�d"Oa	��ɲH��1b��9--�\b�"O����-��p/P���Y<`��"O&�kҏT�I���+�J�u�"Oj���L��E�8�vˀ� Q0ub�"O�r���#Y�Qp��3#6�H�"O
P7nb��Y��j�*���""O����#�d}6y�2��2��)�g"O�D
a�60;�T°��T�@} "O�0�A��#T�j��%�+���;�"O�Ż��[n�xa�dӫZP�D"O���X� ˄�2 !��V%~y!�"ON��u)��7MH�Hp��03��yp"O`�s�gH>�8TS�C\��5�"Ox%+���#*pN d"ŵx�H	 "O΄ ��i��E#"@ڧcf�"O��a��H�p������I2��"O�\b��R
����& �5�����"O�������������WYN��g"OJM���Ɛ{=��s�iM�g@x���"O��Y�	�
pFҵ���ʹ��hrT"O: ����z��8v/H� ��,��"O�-B���9Jt<x0L�	Q��K�"O�P�����b��$����	<<q)C"O�5"�ψՀ��S�ƌg6��W"O���Öz��a�v$U;��HA�"O�33 �x�P"3Q�hl�!"O���6 c����?Ј�z�^%�yr���0�`<�'�	�2��8RT�.�y"�ʛY�`�C�))N����)�yBe�(*�m��jB"1�9R�O�y�Z��U��L�*f��X�KK*�y�D�5~k�e�3�\� ���
L]�y+S�Q�2��c�
�"��J�L�'�y�aD,O�@ъ�lJ){�gɯ�yrB2^��]��ݨ9P68�5k_�y�cZ�K� ʒA�1�����P�y��&�fXˁ���<[Ih�
�/�y�잙��Aǈ��8�%PAC��yrf��s�tek�iޚg��	k�'��y�K�f9ʅ��'.-]�	���7�yb)�#6-Pp0���"�����y!Q`�0xq�.���h�K�$�y�b�����ab��'��8����y"�Y� 7H�:ׇH�zt2�re��y���7�����tn^x ���:�y�B
�T�j�#"�o��p�BɁ�y⇊8f�yz���:�Q���B�y�k�v#��x��+B6 ���K�yrL��*��D	 �&e�azt����y�J��>�*s`�+�������y)��'F,`cT�?y�h�r ��2�y
� �U�a��2&��4�K!�yR�"O0](�g�d�AX�����"O"
a���q��X@��	3Y�0s"Ot����Z$X�Ġ`0bH�J�yI�"O�)�P�۳'�f���t���"O��΁�\�f��u
�A�R�2F"OF,He��!Z�p)�H_5hؘH�"On`��%$$���RrjX�<���i"O>(c���.�� �镐g���s�"O�ir���~�������U3�"Oƥ���>F+I"o�A��H��"O�����ܨJ�MF�߻ �ThP"O�]���" d4�r�զ��E"O�1p�J�\��1�R���'�j���"O^ͺS��.��]� oT�]����"Ov���팗w4�c���	��t��"O�)���E�J���D��,��"OV�1C�6�<�p�̭"�0�0 "OLq�ċA�ܐ4���0��C "O�4I�N��H&�8q$�_(l:�"O �%� p�dhdN/�8��B"O��1k��_�`��AD��qb"O|�G��"@���S�+7�x%kb"O|���߻<�ƌ֙2��p�"O�Di[=��}�0F��fܨ,2�"O }	��׃p�2���]*=�|j6"O�%����[B�1!ՉE�bD��"O�A��JW`DD��?���"O�T�� �l9��+,D��A2"ORm��	ػAr����M9@�]��"O�p� d�8�4qƦG-.\U�"O^m	D�K�iW�0KFE^d����"O�xH�Β̱4&״vm�1P"OH��J��N��Ukae���8�F"O���Ē*�X�C� g;,���"O���K�["(��#6P貗"O�4��E��`�V�s6��+� �d"Ob���3s�����ƊD���u"O�d(C�F& <�#��1;@ܩ�"O�Ie㐽L��	���B�P7��"O��j� �-����d�`���"O4Da/	59�bb]�'����"O.����ߝ@�:�Z�k��]���e"O�X�K� ��ԃa�)[�a�"O�+7��
!c �y�g��n/����"O���
��E0�@r1��)S�\�"O���BH�_��#�l�&��"O-�%ٻ=u`� !|��H�"O�u�t���p^�$H�%����U"O��l��Z)N��K� &����A"O<���#� <�4k�iI?A`E�"Oⴁ�j����)�����@Q"O���d��4��`Rh�P�"���"O�1���h���!F���!F"O����m�A�
`ْ�0�*5)�"O��
�B݊\�EZ�$M-9�<�:�"O.�R�gVc�D��"��z�ڱ�"O�h� 6Ҍ�t"���$��"O����,B�@�~��@�P"O�X�3BWs$�$\(H�4�p�"OH��䃲⤡�r��Z���˦"O�=�
=D4e"��0[��]A�"O �KQҩu�V�e�q��!�"O�l��Ů��I�'�Lu��{6"O� �-��`V��Z��Qߎ|c�1�t"ON}
wM�i��B#[#D<$0�"O2=婅���c'��Oj���"O��)Â��Y�Rt���ـ"KHI{B"O(I�5��#x�	�c�
20�#"Oڬ��,Ba�Z�C�� f���"Oޅr@�B?����`C)) �i��"O:$4͓1Y��T�w��(
hl��"Oy��E&��X�����L��"O�dA���`;���6q�^��"O�}	s'�'68�Z1�%��mT"O���q$�' nb��%
�v��К"O�����B�S
�r��*d�F%�0"O�(�l�h7+
�=��$��gO�<�G��lr��G̙)��	d,Ge�<Ѱ��?`�Kg%]R۴�@!��]�<!��_�\���25k��9Y�IQ��_�<��`��F�0�`%TDY%˓X�<a��#X��\��&M08r�P���W�<5aٖxʜ�i��M�.�U`pI�V�<9��%I�}��؄ZJH�K�� H�<q��/p��v	�*���@B�h�<�c�ѣ)�ٺFQ%x��?H<C�I���{���`������^�.C�I�IϾ@��LK#�-��L
8^ C�ɚ �x�f�d,h��a����B�	�xx�RLۦu*]r�`���B��!V�bp��`�T�^�y�)�dB�I:��tB�]���B%�^�kSXB�	64���ĵg�x��A&%nC��}��;v�ª-�"�y�,�YExC�ɾ_�ltb�"��DE�����U�SQ"B�	:�j�*���7��
T�@�HRC�l�x��ݧej洡��S�A_C�I=P:��tca���wM�)t��C�ɑ����V�6�l�e@C��B�Ɇ���������ʧ�ոfuzB�I l2�%��_�,�{5,ո*3~B�Ƀ*�@7���=�4=��l]#K9�C�	(n(�&��$��Ө�n`�C�I:;� @  �P   b
  t    �   �(  �2  �8  	?  LE  �K  �Q  X  Z^  �d  �j  &q  nw  �}  9�   `� u�	����Zv)C�'ll\�0"Ez+�D��4��M;�(��<1�Y̟H��Y����4gï���b�愙2A��11��A�"�Sb��{mX���c�u���2��t��?U���C�}����B&PVD�S��(*��P�\��h�'�#4�Ibr�λV��݊Wh���ğ��5�^��@[���m&��P���Z�[/�?���F1���۶��j���Ӕ:o�'��'����ʘd�Z��ܼJ���$��'�Rh0w�mӾʓ�?aŮ�����?i$�^cᔽɇG�8m
.2��?!��?����?��C�%�?�p�G~��O���SQ��=J=��w�Ҧh2L`�"O g��3]B���!"�	8�U��S��Fxr�Oh����H����� 
��=�BZ�vz��MU::�';2�'���'��'3�Sμ��H�w?"A��=�"�A��@�ߴr0�v)|��	�'1�7�IҦ�Bߴ���'6�\�č<���ӤI�&	�=���I�-��>m�#T�&�����"4u�!��L�H���k�]��C'Wv�|lm�+�M[�i3��>�ƙid���X�"�5��9M��)R�܈cP���'S�a�ĨKUf�]ñ���JI
��5O˄M��Y�g���nZ,�M�B��6
ظ@mF�EI�Q���É�jU�2��t(F���ix�7�P�2��>&P�� �
,]N|��JH��la#  &Y��aa�e�a����q ��A���M�Ҳi�86mʱ0e@D�� r8p��eU�LL���e�M�4�3���%v��(bcR̦�aT��&<�pE{0�	#`|K��ݟ��?Î�"Y����eڎY�<<`afO�?)���'�R��,�r7m%��������-H�"�W����\�'�r�'�rD	4�\9��,b$�1m�O6��AĐ�e�X:}�F)�7�ù�0<!� �7�TmR7J&yq���4}w��{�5鰑��Ҵ}�؄(r��cԧ�?����N8'M��i�"ϵZҨ�c�
#q��'<b��S�D���bG��T�v-��,ܦR
>����H�A�	h�x!������,�6,�O���k�l)�'�y�*�Č8��ˬ}VM1��W��yB�V4C=,�X� �A��+���y"�YE��E��<_�Ț��y���FY��{�o�'��2@� �y"�µG_����Z�&�����Z=�y�oU�|
|Q �$��L��H��I��?1P��#<E����"R`�����)y�1i���1{�!���uΈ@�N�[L!2�T)!�!��G�L�uȌ�0�2����!�I*a����i�c�fl�a��*x�!��=<�(�ƚ&z��9`���o�!��ɶL6��3U�C!P�(7Ð�=J��=��|��	�&�^ir�K�����O�I��C��� ����(�����t��C�ɹ+Jс��C*a��0PL�%O_fC��lgȀ��b�Ysf��9n`C�Iv0�z���/c"���l�����dI�a.�m`~�^H�Ȍ�`�/t�f��s�ڙ�?	,O��d�Of�$R���	��Һ8�\�堋������*nXl��"��Jb��S�#O���!Ę�*��]k B�Av�6̀�>�T�	�ش(dɋ�gɢ:�I ��p`F�����UP�4�?ya��.���a�%dbI�Zbd�'�哑}���ʳ��{�Du�4	֨V6���\�t"	�M,�AEҴ	�j�����OV�OB���c�8_m1��|ޕ`ea���Z��I�&���q�<�������YW(��<��Y��s�<�@K�
��)���ݟ���Yv�l�<A�@�0��0�vKA���1fO�j�<9#g�8T�P�ye�[��hC/Fi�<��ȍ�0`��I�q�n\I#� ��M�H>��A������?�����dщe���T�i��i��9�Xo�:��3�iu��+�F_)����'p�Q�j��f�b�1c�[�R��5�Y��R-R� 3�����-�O�^!8�+Aq?�U�\�~����!*z����pC��MSt_��W��O�c>�D�O��D���LB(yN~0��J�Vu`��Di�6�X�z3��	:n����P].H�'��6-զ)%����?ɕ'��H� ��'�<�R'� 76�`�0���	��7��O����O����'9��9uHQ���EZ&愥7����ŧ\0�T�Yҫ=U��C�Y�����=x���p'.�:<Δ�2��@�X;�@�fM�A�0��
�+S��(!�e%�c[V�3DH
�<	*F�Y�5x�Xb��џ���4����O����O4���O$�	��٣�0b�V���ٺm^H����͢,�����

���j"C�	5�M����)Lv���OR���OD�	���Ȑ`����Ëc�B�'���
��'T�>������S��=d"��Q��� `��dI�G8�Ps�HW^����B�' ��a�k
�#��)��~r��׌���=�/�4��@�k�$#?!�Q�P�4%	��@��w�Y8XQ��1f�Ԉ�̒O��7LOp �1�cu� ���2�$%���'����P�2]NI��Y%	Q�8�ꁇ�S�lx����MkO~��O���'\������I��g	��Xl.]@&�'�o�@��Y��֗V�xa�;O>�u�F�'�~u��iO�}Ʋ0��+?q��_�{�R�`��U�DI�گ��q ��6�ԏQ`\y�Pc�6qrd]���䆮mcR�hӼ��O&����I����c oE#m���L7a~��O�d�O��$(�b�Ф�%K��	�"��58џ�q��)̊dК�R�H�C��H�dB�<	�ꓑ��� Y�m����I��8�'Ѯ���D$x�����S����Y�����g*.Ip�O{�i�n;����CGϷo	��{�MU��,l��, ,��^(,��c>-�u�>���"UH�Û7�v� ��ϟd��ş�q�m�ݟ��|�'�B�Y�fmLْ�M�qm����	�V�:">a�y��o�� 3��?7�~ة� R���\P}�[j��'�������鈶Sa����\�DP�HK��[�p��a��惡��؟��	]y2��D�)@p�ٲQ��*��		0��-���~�t���V۴E�@'�6 �ɦfͧM����S ѽ"̤"3�ǁ|<���iP3>q�>	��<D���h'� ��F�Y`�d�	˟L&�h��J��<a��ЧU�v][ŋ�7o��(���y�L�,�����	{�Q�ǂ����	gy⇘50��$}9�oܹ!��S0I�&����C�'�����	џ��E���T�#%��$���g�io��#ɽ>�X(Ԍ��(���	�1*
Y�"���U����7�^���Y���t�(���74����F�5?��>q��Rџ��Ia~�P�_q��s���`���A�!��Oj��d� =7L,��ɓ.*M��R�J,�2��OJ�Ӣ$͑|2H����-tRs@�'�	�r�N�A�O�K���'K~� ���G�Rt�+L� H���'��L�?r��
q�~L�E��h�ʦ#|��V%t#�uaV�]+!���0�h�q~��'a.���f�Q���H�=�]�}z�o�Bl�F�T�p�7��p~2���?����h�����G� ��`�	�O���3w̖`�0C�I �P��T+7J����Po�(0�?��퓌��İ����7�t����Mo@��']�	8c���֟p�I��4�'H�����T�$�H�g>�MD�P�
���F��O�M�u�R?P�1�1OX�EB�0v]+cƆ�W� ʰGI�D4�tAЇ{�>�	��Gs9(b>��P�>��� �h�,@�e_�l���
g����'�B]1��?����ڥ'� 9�@&u��lQ�Jܐf%�C�I�V���y�'t�|eI�P
>|�˓\c������9�t��G�C*dB�)r�<O�"2m�O��O8���<�|jm�)i	�#��-֨ڴ�.`8�+`Ƃ�u�@5 3D��z|�yb#�,A?��Ҁ�!=(]#��P�  
P.������S�]SǴixг���
�r� �H�"�&��s��!e2	hP�'�B�h�'@��I�%O ���`%X49k��R�'p�H
�.�%,a�����RHm:\XJ>W�H�?y#Iz���B#Vm�(8�I�U1���	VR�<��Ài���G��X+�=T�B�	�H;���'�/�`P�%�~B�ɰ��12����xȑ-P^NB�I�:ԌIѽ*��d�)K�W8<B�I�oaB)�ЁK�bѲ���>�Ң=��
�g�O�u����E�"�����s
�'<�D�q`��*Y����싺i�4x	�'����K[9U^�Bƭ�*j2�#	�'���"��%On�j%e_ 	٪<;�'^|� �e�[�b��$dI�Ѡ���'q}����<q7�0Tj�>q|���7�F0Dx��)�p�(lZf���Ur�Բ&��?�(C�	' �D�f��/I��gk�*�
�':�-�p��kv�e�ɣd?jEs�'��(Z��r�~@$.a��л
�'h6j���-t�:�cK]�G��
�'��T��*��h��� f�$C���2)O\0�'�,��BG'5`��gƮ7���3��� L�9bJ.��=� IXW��0�"O8�V���r�
4Q4o��Hʬ��"O\Q�mH<�Ak�'��.1"�"O* Y�D�=�D����P�Pm�Ha�'�n���'� ���޹��<���${�&��'�X�k�MUh�K�L�w��ͪ�'�����0�*�$�Z�v�B���'Hz�/�LTԁA$D6�ٳ�'4IÆʌ*54�$�3 ��D+P���''`h��E�!bY� �7-^����d�g�Q?=që�:A����K#pA�@���(D��J3��r��@K���#V�؜لh'D��P���c�|�B���C*�x0�1D�`9���s����"�2#Q��31e$D��! ����JWo�,t��K�� D��oZR��]��Vԕ����OX(�R�)�iv0��Ø�ef��1H�<p��l8�'*|��c�>������ �n�|�
�'f�!�g��e|�����kEv�Q
�'��8R�mʏ|XPj�0f�Q	�'!b`�¬�1/���Y^�X-)
�'��-J`��)o~P�0�Z'�\1c(OZA��'���Gn��ǂK�&�����'{��ʵ�C�h����e��%�Z1��'">�1�U(r�>t�@�d�R5��'NL�Q��w3d�����X�z��'����a)?ky�	i��;i�ma�D�8���56y+1]�H4�劗��/�~�ȓE���h
8c`ѢD9A74��l�F��f������0o�
qi�Շ�b+��V�U�A���� �!�����>=���FOXA$��bB�pn1��%&��cC䈸K�ڍ�᭎��P�F{2�V����X�I� 0~U��	3E���PC"O:��`΀�+�����#�0����"Ol��� �0��Mi��M>G� QU"O�t�2l?"_�0�jQ0`�Pب�"O���f��M��B��Ψ�2A��"O�-��S*�N̸7g��vm����'B�X���S�i+�DXr�E�x[� "[�-#,��ȓ,|��2$RJ(�9��_�5��$�ȓ^M�l"㥆�'/
8��#	_H��ȓhT�M���Ā#� e��EűWt䰆���]Y H8����F�-������������>?�Y�WP�	���'�{	�[L��Q�;�*uztlB$)4ZՄȓf �ٶiʮh{�����ģV�N��d�p�S.�9"���2-47t��ȓb(HP�'��:�����%M-lTT�ȓ�����)��X������,i�pd��	���	9 *�AЦ��tԺ���OI�d�*B�I�)���b��m�Xh�Q�>jB䉓f*�K �@0�Dp�%�3�B�	\�RL3@��w,0���c��C䉖H�6���oT�={@Q36�]�eƔB�I	Kg���n���k�F��:���=��-f�O�%:�����X�ac��*yp�'!�l�#�ƎP��I���.�p��'���7&r	��$���m�P$a�'Ǻ���:7��
%mȋ2�\���'�4)�ձ�h��쒴9�x�1�'��*�(��^�!.�	}�^4a�]t\Ex����Q�,"�-�0r|;2�R�C��9O�Ȥ�nѬ{�`���ێZ6B�)� >��1 ��L�ZU�$K�11}����"OT�;6��q���y|��9�"O*�j>I��JϿ6��v"O`l���O�H(�ۆم�����Y��Z�$�OJ��pƑ��q�p�%5�|�"O�E���L�	K�c�R# ��%"�"OP(@kX�+7�%��1b�L��!"OL��$�_�x,�<��-�~��"O�K ��-@���cD�E6 ���'���:�'��Ac"��nl\��,G�m��;�'~<e6�֥g�Bic�-T;L�'&�����C#����!�Z'K����ȓO2]��!�~9PD����>�� ��VXԹ����+vT�@��9BK4T�ȓ@ʼmBPO	2M�ջԡY�w �pD{2�O�����t#��	ֶ��胦f�\�I�"Oĸ{GAҚP�mj�	�JOv8�"O��O�J���f�i1��2d"O��h�/D(V��`1��ɵR�ܤ��"OHp��C^�4���uA�!]�b$ V"O�Y�d��?MF��9D@^/Pr�tB��'9V(���
���KAh��A�0���&���%(�R��z�VA #���<���ȓ\��9�凚%`FPP�dP�aZ���qFx]�qN�s�I�Q�0s,���[����-�1? ��!K�,��H����8еO��	z�T��eH�s��u�'i�R�tL�!�цF�`!�`ҥ e�ȓ@�6���% MonP��٬2�0��_��3�h��
+R��ֽG���ȓc^�(q%�Äl\�[ģ�Ec4��ȓ��`�E�	!ۊ��$_�2��Ʌ��*M?T�ɐqu�a�f��<��иg�E�C�$bZ�A !�*�<8�I�$�lC䉵
Yb@�Z�I܍�⫔3*�B�I]a���BW�2e�)���6Z�B�ɱw�f�D�!�ę�f@
���C�I�2Z�)�#(�%/Ӝ�"�h��idz�=�FSi�O��a� ��d�S�M��?���9�'�>�H A?2^\������a�x���'k^q���"����w��'��i�'B$1����%��N�TD�3�'�d���a�*�$Qc'`T�F��pI�'��A�@36���Y�Y�
��=K��K���Dx��	������F� ?�հ��?^�C��*g�@�j���O�u�ר݂_ٮC䉍9�l,K��xD���.]|�8C��kd��A�ԿNuz��r�\$tC��R圝���Շ*�l�-�=#�
C�	����J�o�zq)����ʓW@H��	8k+�̚�E^
K��T�b���;JB�	!�� �	�\�d�#f�Y�-�bC�IE�a�m��~1�d�Y;~�$C�IG}l�����P���R'ͧf�B�	':{��#Vj��*H���IV����Ȼ6����v,�=a��];b����e�i�<9E	;~���b��NeΌ��Nb�<��k�l�����*�x��KY]�<��n�=L��wA��b�W��O�<�3撨�v-s�W!D���0j�L�<a�I$%���K3�V�@�Ry`f��S�'������I�~��Y�l�1	x��R!݂A!�$� H�P@�bƯNzx���.[�i=!�D<g�ȩ��Y%rt�Kկ�q9!�� ����[8nhQzWL�+�h�"O$�+V�R�m�d��&$p��"OJPv�����Ct��'T�֘���'��4S���әf��m��F����x0끕sG��ȓǴ�Y7-_&W,��:w�U�k<���&%��fNu�C�W�@�ȓq[�<�1��xx��
��k�2�ȓ������J��0y���0>�5����H�-�zӦ19�.Q�/E��'��`	���5Qʉ��N�,�c�&%D�`�֫��RJ��B�8��HƧ'D�����D�R4���� �8D���rFAj�r�t��TF���T�6D�,@pM	�3ۂ�cT�T��	��5�O4� ��O��q���(l˳*��A��0ӗ"Oj(p� ]�O8�k'hQ��\�3"O�\8�kA�=S�H*�M(j$���"OTq���E�2ے���K�yK�$S�"O�ဎ�edP���	$�&dh�"O�q�燞,F4��Ek�����I�8�~���ѳ	[D3�"�9
��iv�u�<Y1j���Y�E��#��|�&�n�<���� C��h�"̮?�JpQ ,�h�<9pjA3x����*�;܊��� d�<�g�ܕ
��MC�$�'c���� ]�<���W �ʡyk��<r)P\֟(��E#�S�Oux�HDHԷ��e���H�"O�И���&n�]�CCE�XX��"O��҆J+��i���q�>y��"O��NY�3�E� Q=�*���"O��Bd\�@�a�3�p�CO���.�'  9��ٳL�e�4m�O>�'f$�'�5����� _"U)�$B�#�(��
Ů?��I֟ �	��2�Έ;�ظ��A�:T�z��|��Ft��tj�7[#4���?K��L8���k��u���ȾA�l�m�!�����E�0�DqȤ�T,���`�}�'�ȸ��?���癨?Y����η{���բH:��D*�O�q:�T�7���X4�T
-�NEYA�'[�ʓ
��F�X��У�*R���'e��S�b�R���<a*�r���O2��?�}xp��+�p��!��O��r)�0��$�1��/렌�)�l�<Y�͍�E!ni�t(��r���̓	�4l#��R=x�Rm!d�r|7�͐VQ>ay�`ٌq��Ų��Dsp�{ �h�� �*�O��D!?%?��'{p��4&C,e(R ��A��|:ؐy
�'�>M�����&`��o�b�ۉ��N�O�q�/�5;��}Z�.�X����'�剳2�Q��ן��I��|����k�&O2Z(s3dK�Vy�(��Ё�~ȃW�'h�#fဪh�L=!ʟ����J��4�T(Ǉ#8jp*�vC��l���A���}��4�O���=P#�#.�Q��և_(�I�n�s~���?���hO��	I�!	��<�`(1�����(B�I<:D.1x�ox�!�H�;0�˳�'h�#=�'�?�,OND)@"dm���Җp:���X:B���O*�D�O��Şc�����T�SÒ��d��7�*%�B��^o2P*�~'�D	 �'?��{�쐃I�K�Ńy������.R�ȍiG)�+f:�\�d�iE�l��$ܹ1��oЀT�܅��&�P)�=9qS�|���If�'�65�4�1%�#t(�$8O�X�'<E/�� �J�,Q�M���,O��l�T�'ցp��$��(Gudh"KW-Rm�u�� ����'m��'��Ǜ=pDp�$���e������O�B7<F�q�1��a��,S���@�D��@�b] �]m��
�, �Û�H�
��JG#wnܑz��DN�'C~x����?���4�'����慐 :M��3�Ȇ��:�O����CO������Yf��	s��'0.ʓ)�T���(���-��#_�&\ؖ'�&t���nӠ�d�<+���D�O���!Y�#��5�J
a���i���O�uC1��%f#v<��ׅPa"	�)�6����e�J�E٘Y����7��u�B� w�]�. Ls ��M��KK�O��aaH�*��{�'��YA�a؟'�b�8���?	�O�O��)� 5"�k�`�rM�c��px ��"O�s&d�Yz`y��(��$�퉇�ȟ�4 �k��aeoƖZ��Yh���~=�˓�p�2v�i����'>P��I6 ��Ź5�է1 h�	%e�hv8 ���?�1�H�f>��e�Ji����<P�&1zB��Hr��7�r}JV�~����Y_`0d�b�4b*�ɓZX�T�S`U�x�)�$�ʨ�*�e�D��ٟ���R����$`�61�j 2q�A�/�lq�"���y�b�9{
r�Y�$�����G��?IP�i>U��G���W��`�Q���H�.��5���Dՙr{6`�m�/�j�D(E�n�!�$ʔ[�8H[��M/)D`S�G
�m�!�����*�─����,�!����9�f�W
K��Q�-Ѓ2�!��� ����(�_�"�A ,X�C�џsci� ����O���1��̓#vM�eIC,�|�����D�(���OR��;���9G��B,J�` *�'K��jXw۔$Kt�۠�ܤ2���T!v�+��$S	S���*� �d��I@�hOq����%(��r��x>4�Z�̻#�H�D|����?�5�iVГ�nH�햟fO���'J��*3t��3S�\�	o�𰃫��uqt�;��.w����Rj(�Of�'x��J�x�M*S��>O�Z5S)O`�צE��Q�'���O��h�b�(7�����эssj�#0�'jўq �
�����Y�(�@�)��eO�c>��I�?3���(�+M�$PJ≇9�M��X]�y�'@>�����?����?��'L4�zb�B�+�Hő��W"�)"�l�)x�F�'���Jg�'E�B�6����u��#�1g
l,�T��|�8!�v��.~4�}P�@�O���"m&��Iĺ+��?����?y�'DD0 R�õE��KG���S����D��?��S���+���yrf�5�����S�_?a�"Gs���q#	?�$�����Oxx9��'��HR��~�'�?q�����y8@�y J�1T�H�he��
I�lL���'�d���?�ɇ��?q�'�Z����M��T����Qf���'�ܷ`��I:�!�"��&:O����'�bĔ ��I�O6�$�B�鶄̟{�*����&S#���\"k���	�h}N���O^%���?��'�T�x��M+�gǞKtD�cF��j����*ޑ �n�d�i��$֖9-�7�	��]��;r����f�^6�`
�+|��ic��3c3����9`�DO8;oR�'U�$�'W�$�g���ƮO0ɺ��X�W��ciƅU�L6@�^�����<����?�|�' .�'�,~%h���)e���ئ"O̭	g�V�^��u.��Yny��V�0�'��'�'�2�
�G*n�T�ϳ2k�u/�(2�"=��T?�Y%ˇ�1�4d���[ !��,��+D��`�#�=x�����J��2����)D�|�rH�h��pՅI6"b���)D����	%E:8G%e�A)t�"D��r��Y"L�j5h ��2 ʢ p��?D�ȃc�Q~56�`qAS�m1��ɐ&!D���~1\��u@��%`��Ă�U�!��ϯz9�e[ y�2}��/qy!��X�z�<�!O�Q�谫�B �ip!�$�<�3%�&(��SU�RR!�dֲ�V(r�ΰ;}��d#ð2���E{ʟ�)�L�6t� ��� A��"O`�[S�C*X�u���ŌG���c��D�,/�Py�n+
�x��&	' 6�Rҏ�U����b+�5~�Qc�ʍ*C  ��ō�:��S�2H����D���h�P�.�/+X�"̂4x�)+F���
�j1Ȁ�o p��0���B8X�/Q� �$�ZF�D- ��ہdi���s�̴^J�0Ӄ�ԡ")��z�ݳ9֛��?�$%��m�?2�i 5�Y��D�O�Ո�E�O|c��gy©$�U��V��4h�e�R�hO�)��)�S*a^ő$+���Z`��aVOD����'�1O����W�n�ze�F�ɮ��B"O	�@��|g6f�!�V�c��'u�<�"�/y�$D���*O�f*��?�<7��O��$�O0��E�"�����Oj��O����������Q H�������>N�%Kb�"^
^����
��l���;�����N�*���P��a�v@W7~�l�Y�2QtlǮ�H���F�)Z~��ER��J�I�<$�Zؐǃ	�S�0amZ���$F<�O�����R�J�r������d�Jgゝc�!�䘧*�Ҽ�b�B]Rd�&�շ��c{����Od�!;|��N�8 ł�"v�� L�X���*-�z�bH&Д�"�6f?�܆�S�? �e�֮��`p���� ƈ@ʒ4)�"O>�ҩY�Q�੃����W���"O�C%e	�^/�z@�Ǚ^�(aP"OVXB�&�0	U x �=�� ��"O`Q��JA�r]S�n	2}���a"O�`*���@���Ц-�/���"Oڔ�tK�7�"�����.]��"O��#�S!V��5��Ô1�P��`"O�iXŎ�P֪��(^o���ж"Op���g�<��1 a�0Y8�A0�"OJ��K܃(j�YE/ ,�	�"O6�q�$��gM�d)5d�2}L����"Ol���d
���)%S$��}�G"Oj�3q������bmP9:�аr1"OBԨ�D:���S�$X�|W�R�<�N��W�~<@p�2{@ EHO�<9dmH���(	Yl���tE�<1r��
����P��/�t�Ps�E�<����]zLA����+g1�u�2�W�<��ђn���1U�lSv�r�%�z�<������a�$�$@����#N\�<�'	��S�P`��#�M}�)1�N�[�<��e\�8M�ѡGLP/D Je#�/�Y�<�p��b�gX()����E�q�<���>jE�ԯT2��L8T�n�<鑡F6)���#���/B�1�en�c�<)���9G�P�����S���K�CV�<�S�(\�	��牗,P����BY�<ن@D�PWj����Mva����I�<��.P�_��iyp)ѓRlh�$��A�<�V�'R�Z]��߹]WjLڳ��e�<��h�6�Ass�G�K�n�2�k�<�t��+4����F�M�x\� ͝j�<a�MN�@��@1R�u!~�P@�/T���v�X@|��h%���,�����?D������9nM����4X�:�yK:D��* ��J�(�cb��7;C�9�j2D�@�1��6EህB�i�%���L-D����:0_�����_KՓ��)D��d˜���@0,�"}2��j�'D��8��U�V��b�D�5l[���)/D���!�U�V#�-;�� Y0>���0D�����E�xh!.#1� �:�/1D���񏏓$P�D0�*��RGָ�6*0D��կV��q��,�����p�� D�\JFi׋]� ��%��w�\,�I2D��z.ӆ2�͚�#�:@YQH/D�8���X�`7|���h
*s�����*D��s�.�	T�$���F�\6��ƈ)D��rG�r�t�)�C�6�ڼ� ,(D��� ℐ.�@yɴ�S�\t�X��%D��x�
��"x��!��=�U��c$D��i�!J ?����pʓ�N><�� D�`�"�4jc��a�)~ul�d+>D�Xrrd�4/\r��*�	���tk)D�Ti�'�^Xp@G*��Q� ��ӄ<D�<)���R.<A��! �d:��9D���פ�k��M����ll��^<!�$X<W<μӶ�$sP�4�<!�$�9 A������}bh�8�ʚ�|!�D@��$����3dN-�SZi�!���!ܬ�x��^�XN�<��*�3Y!�䆀[�؍A�h��ND�Y��	FR!� A�b��� M�FP�3G�	
3!�� ���s(Glr*��Bh~��B4"OZ��'҉��i2*�2cz�db"ON���5&c��s�Sc�a��"OT����ג��rH�)q�Iۆ"O�	���^az�Ȓ��I��"O�`�C��+F&-��̐'
L�"O&���,Ӊ.�fi��K�]v]3�"Od��G�N
$ ����"�����T"OPT#��^�IbO�H69"�"O.QJ�.��a=-����R6���"O,�J��@*Plz�m�?*��6"O���0��F�����%O:xQa$"Ol�����"Yb��RC�N
�$X2s"O�a2�F\�SF,J-8�"O����Bˆ5I�9ӗ��<Td�"Oΐx�IW�j`Y�#ś3$�� "O}[���0��倝�Y^4y:t"O^5����U� ɹ�&�=N���"O��X�bW,� �����9�x�"OĹ��(݆-T�a��ak.T��"Oj�M�*�t:�$��k9�i�"O�!ԍ�ql�K��I*/�@Ct"O�h�gS� P�H���zl�$"O�	b�ݱ+$�y �;p��"Ot9�b�s4���)��"���Y�"OЙ0�$�{@D�7OA�tNu��"O��cg�ަ$P�ݪ��i�z���"OJg�2Qt< ���%B�����"OZ8H�	��z�(��=p�� �U"O0)x��-ԂMC��,(��"O���4,�V�1�BնJ�>���"O�1[��ߊ-лu�Y�Y�"a(D�\��j�p�hy���ԲX|�d�WK,D� ���
�v3.�ÄU:-�xT���+D�p8`���9)��2% 3W���c'�%D��!��̒S9�uۓ��*=���a�%D���M�Ov���gn�{!L'D�8#�P�ZI�����A�j��8D����fX�w����kF�<�`��F�6D�X�p��7D�ܼ�ED�Wv��C�3D��ч�P�kv(�g� 6XS�/4D�B�Η�w��Uc��(�'"3D�3���D1~��סU�+�� D1D�l�S�� eB$3�B�?��ɱ&*D���	F�.p�q �`>N�%X�'D��آN΁3@�L�i\e��#D�ĺ��6s�������ra0))e�"D�x�K߄bѺ��u��F5�#.D���`#^,;R���E�V�4�B1�ǋ(D��qu�J�~��<��ϳ{f*m��G4D��!R�&��)pLM�/��k��4D�hhU�8�z 	�Oހ˜æ�$D���葩(�4dqBA].�$U#D�1DKݣj�0y��R�dt��� D�d����Z��Zf�Ց�"D����[�oք}�A��.!
mX�&D�P�29�0
��x����'!$D�(���5z�̩O���Y���!D�� `4��|���	�Uc׀+D�,��
�5N~Z���� K *D��J��Z�(Vu@�ʎ�9���*W�'D���$(�M.���
ɿJ:�I�N'D��s�B7S�T�w�0pp�R��(D�x����JBDH��N�QK�98��'D�� �04�T�L���u�+�xY:�"O��1�
��!���3.	s�yc�"O⼉�擛.��i2�_H\TA��"OZt�4j[7b,�٥��D�Ȅ	�"O�,x�.E	�Xh!�N�s�$�r"ObѸsB_>N�䊲L$�`;c"OJtw\n�PY�Ė�f�*La'"Od}p� ��J)@��Z�N��U"OĀ�� iB=��JO��ܙP�"ODJW�o��M9fI�#b�h8�"O@<zc�l��� �� F[� +B"Od�B W�5���"@�]Y�ع�*O�M��ē[��@z���R�(	��'�^��!���tu#@�0F\��y	�';z�����<8+���嗔S��y��'y"��WO�}I���7�v��'J�����E̑��� /PD]8�'�8	KR�Ϸ4�J��!��4#@�x��'�$ufϘ�a3R@��%��iJ i�'5����d]7��I�` �o�Ă�'�N4���"2��Q��x���'3R��9�1���:s,!�'�fa��9a��D�V���6�Q�	�'�<l��^�2wй:�N��b>�	�'}��珝gyΤh���":HS�'$���棝�c8�P�jǪl�d�
�'������}�r(kC�I/8���
�'�0�`B8CT\��V�,Ǩ4	�'�ج��HP�,0��٥ye���'o�䫑J4^� �'$_-c�\��'��qZq/y������W���@�'e�|�m$E�PC��O����'s,��v�	0�F� Ǝ�1�d��',$�2&T"8\j�ce��/@W�� �'�p��%�b�Z`j��2�>0��'q�PC��YL����遵X�ݩ
�'���x+��}i�����Uo���'z <��H،2�Jd�1��H��'뢡�'Y(~����$Q!z�'R�æ���q�lY́� �,D��'ƶH0n� #����A�!t_l9i�'���k�싲}
������re��3�'���(2*J,�f�p�k	5jI9�y�U.�RBfѨm`�
7č��ybi	�%0���	_����F���y��$_��jT�;Z$�T��ŋ�y��JU��+�I-Y���H�y�΃�ƚ�J�M$;p�2MV��y"�Ǌ����օ�(s��13T
��y�l�;K�a����.���	.�y�nΡ` �Q��%e���cJ ��y�&��P�Q�˓�Z�\���(��y"�E�|�9r�nR|��������y4Tu��b�eFM��P�ٖ�y�iWKU�HV�שBH�|j�
P�y�ʎe�QB����= 0$k�ҹ�y2(�<5yfɍ�`.�Q�f��yb \%0������\h���e�0�yRd�,�0��3h�Z�	#����yFJ�S�@�uHQ��Ɋ��yb-�"7c��!��}� ��4�y�8}�(q��O	�U������y�eFsw�e�}�&@���3�y��H�e�B@����r�̜��L�y
� 4�D�$35p�QM
8Z�h�c"O*1�bT	)��pL��7��=�t"O�M��͈K�:���kWG�~�B�"OtS(`Rr<���Z<Nh�`Z�"O�e�$�MM �S.�=.��'�54��*r��a�V��F�
���M,D��ÅKL�FSq�ŉ�!��)�B8D���c�O�F�T�֢4�r!�a%D�<����~���B֊L�2�F�0D�ȺT�ݑi�񋇡W��,`n+D�����[�?,����XT�X���*D�8i4�E;�e�#��!�7D��T��r�Ri)h����Z��8D�+�Ϟ�bL�=��ᎉ(>�*��&D���T��9e}h��聪�]�6N9D���+�1���3����J��� �&D���f�Z BJ�bD��C
�U� /D��P���"�����bL�b�X<P�J*D�� t�FA�� PF�ưT�̃�j)D�pkU!Q����B�%����"D�h�5aR�U��,�V�љ&� R�<D����B`��Y�P�p��@�%D�H[�eK%��p/�޲��R�&D�L�ÎY�,1�L�p�]�X����$D�t2�'I�z.0�q��}	+�%D�tTF�88j��En6�����$D�8a�&i�5Y�F�f����#D�x9��)��SԄ�.✁ J/D�89��D�[�(��"K����U�0D�0��@�'��kf�����*wI1D�(���-��$@Ư@��J���a;D��K����2������=#W��B�3D��z(O,`ZN|����'%A1�	4D�����8Q���3fAE/H�DQ�`�7D�  g��~��l�֮�31Z��1$b;D���5�آ`ࠤ�S�A�J�6�'D� �d�۬,wЍkP�ҋ!�fqJCj1D��0WE�?�<л� �@&��W�>D�Xi@E��n���$
P����w�9T���4Ù�I�Q�c-M�90�[�"O~5I��Ϊ%��)(DK��\�н84"O���l	Q��)����YA3"OH�,���h�A�j��JP	ק�!��ƙ�:�CQ�=���*�a	5*�!��Ġqx�%����x��Ak7 
.m!�d��
�CC�ŉN5�8��H�z6!��G*%2�	��șW�d��I�:R!��� y[����@�0�4�ZsE�)E@!�DGIGd�*ah�n�ɖ��:�!�$V�y��I2��6>r�8ȱ	R0k�!�D��%t�p�Z6:��+��Ŧu�!���=c�ny��Ŝ��=Ywa F!��h���� ��&Jf9CCaƓ:�!�D޴Q1FLIEHEH�0��D95�!�F%��iX�?��	Hv�ܯ|^!�$�
i�X�X�%҇f�����_1|!�ݷkIB��Ҩ���nlcbƚh!�d̟z�x��p�
�v����o�"8h!�D�9Il��D�ԛ*�dxan%:!�	w�B&-��$X��g�qg!���]�0��G�C|�|�dHK$C{!�E
�`m�&J�h��!U�!�Z ,��'��~~��8�
I�!�Ę�T'�-��d�JSN ����$>Q!�� �k�">�r����!��S�"O
��4͂=y�@�0)� sĜ��"O ɢ0�TR]X���nQ�x��Ӧ"Op`�v
V'�@�����g&	 "O	pU(q�,{vM͂��`F"O�Ɋ�"�.Q�1JS�� �m	3"O��S��+7B���H�	�"Oʡ�u���^��v��0q.�k�"O��(�%~�h�[�"\�2m�4"O���O'KS���!�1c���"OR����9rb�JG S2��"O�M)p�Ӻ,�=Z��Y7~,>�z�"Oʜ�t����H��&>��IY"O�!K�@TkiBY�'*�+'��uS�"O�E1�(�C?bdPfhUr�ƨ	W"O���D��RA�0(\#MժĂ�"O~)k�!�	RN�jǯ�;88��C"O�ɲ�a1�d�so�#<H@"O��zDj�[�(8�gK�y�2<�"O�:._s�:��F���t��-C�"O�@p�&�SI����狵{ÚH1�"ONIq�+Y�iN�!j3'��%���1"O|�����4��t���	)�� 6"O ��A�Q�U�LQjd�^/�0"O�x���5VUX5@Wl�-' �ڇ"O,8i��OgTx6�[���j� 5D�l�7	��k�xD�/ET���'5D�����d

sÚ2T�25SĦ D� ��݇~�@�Z�M'�:Q!9D��(" �ag��D����!�#D��X��Ӊ2��f�1q���㒈'D���@��=-��	�P��\q"�&"D��� O�0i"<���۪,e4�Q��/D��Rce\>LD�C� ��bK�\k�D/D�X����1K�&г㏇��� $�,D�`���>S�Ĵ�SG�Fjh+Ɖ*D��`Pl�!R"(�P׏R�5�\9r�<D�p ��3,\J N_�=�\P�:D�d�E�_7��]B�#߂A,yP�#D���'�L@�ʤ2DK� 3g%���!D�0�@l�4���7���2m2D�L� ț5D5R�Cd/c]�Bd�>D��h#��uWH�`��żSjd,çJ=D�p��B��XYfd�$C�}���a5D��'MA�D�xp��Ǡ�o/D�$��˘�T�2-��M�fUx�:��9D�zV��_�|i�d_A�F��Sn#D�\ڃ���p0����W�5�h� 5D�0z�&�d,���!�H�~=� �Ņ D���+���Vk"n��Hb��,D����F�#8Z���L�����P@�,D���S�|s�Ȩ�n
��q�� 
o�<1֌�,
�N("vHӠ_�J�v�a�<�_L(*��]z�εI�/H\��B䉻s�0�C�ڣ;��H,lY�e�)D�d�.&���J��4�V){u�<D����.����P���-��"�9D��:4'�?�J���ָD�@��d�%D��2bg-�(��mp�r�"D������A��p��E�R`�G�%D�H��EA*Y�<iҭV�k��'*/D�̸���bƐ���iDm�׮9D�@ˣD�V���QA�L��T8�#&D���Bf�=mev�����2R:B�*#D��  �G;/x�|�a�� <��"O�y#%�,!GT���-L ��"O�<�G���WG|��v�B%(*ك1"O`��џ_Gء�a�(lr""O���s��y��KV*&��##"OTt0M
�:s������Lf��g"O*��E��r�4�hRI+�([�"O����]�9�T�t���-t�Lk�"O�I��/?F����)}.9Ȃ"OŐ��L��t��hZ�mv��Z�"O��C�#0ؐ�j�e^�L^tp��"O�ez�O&Px�����N�(U�9�"O��1�<<��Aô��Hg"O���BK��Fd�yq���b��c"OF��!M	����!q�SX�6�@"O(\;@�^%(
������LAV"O�`h�j��8Qp<p�-� ���(�"OpI��g�t"J�[�٘}�Ԙ��"Oz�zU�B�A���3W����@�(�"O����T�x�,�ؤmQ�/�&��v"O�!P���h� r#kM!(/�A�""O���`Y���
���b&���"O@!	lڗ&��9����X���"O�${�䅭/!:��d��? \C�"O���Fa�$[�Z��Z6� �#"O@(��iL8�qi����*x@I02"O<@xA摋,�V 8#��.v��X�"O��K3a
"c�|̱W��0���b"OnY����%��B�fŻK���"O\񋇏��I�4���E�i~^��A"O.����AM�����W�Ka �@"O����%փ'd����Ǯ_F2H�'"O y��S1I<�9y��غS܌�y"O���Ɓ�P*���ǡS�:ݡu"O
 r7�����Z�#8`&�Q�"O0I�
�>�\�v	Y(d�I�"Od����?��aq'��p$@��P"O������!��Hl���z�"O|x�.�!D�t�2䏘.I�DX�"O6�PC�g�԰F샾L�6��"Ot�9Ä	�:��As�M)��J�"O�u �ڵ=�F�Q##S*>A��Y�"O~Q�H���:��,T����Z"O��s뎴�����%)��S�"O�ˁ�#�p�z��[�TjZ8��"OX1��T5���eƘ.U�@�"O�}1W�-_�<��$V6yAlH��"O�ڦ������J�8���"O�S�Uq�Ր��ÏO��"O�4k�ϔ%]"l�7�V/3K�K�"O��a0�� �����¿oPL�e"O\,�E�Q�8#¼I��j�r�"O
 ��	��QV.�6Y�&"OE�7M���ّ�L�I
܁��"O�e���%�fp�0zʑ,�!���e�lX�n��)
�H�c��9%!�W�n�j��E�@"uW�Y�F�*S�!�N1lPD8�CM"]Kz)�ag��I�!�$��'R��R��I���$ �!?!�d��DT�딝v����Ə�i!!��׺.�B�KVe
�(�()˰�@�?!�ė]�1�ҩ��}u�f�� f1!�7w
.��F۳0��Aj��A�!!�R�xn��""B��,d�
�.u!�� lȀF`��fU;��Z�/�T�t"OƼ�Њ��j���\�=�>�c�"O��x��O�r����a��G�N)2�"Ob\[�@�g8��Jv��.A(��"O,Ѡ�iO/��D��"_pԤ �"O��fߡM�f1I��ϳf�)�U"Oj�	D9�~Yb�Q�NJ ���"O�q[ŝ�R�ұѶ�� jEbYj�"OD9��EΉ <.���@ā>	X�p�@<4���+�0$K�%�/YB<|;��$D�d�gJ�Z�>!�q�R�&��%M=D���I�f�a��' o`��¥<D��	P��igR`-�&�D���<D�t0%ビV�2�їhХH�&��CD>D��CG��B
69�L��2��r0�=D�l2�k� 0ä�G��r��8D�t��U�#�0�1�@�$(�$ʲb8D��j�Ǆ2WO��P���x��Q�"D�� �>q��� �_+�N�A!.D���6�H�5�c�R'e�4`:��7D�D��\>l�t� !��
�F�D�8D��K狑�IrԠ�)�!����4D���D��A��8��*q� �Zwo4D�:3�?�&� cD�<�� �c�3D�$j�O�k�H�Bw�uA���U�4D��y�o^	bZ����	�vkG�1D�L��=a�X B-�3�^! #D��*a��BcA��$	�b�;5�=D�h�5j�2$�Zi
���t�x4�C�.D�4����n��噲�M�9CRԛ�d.D�8��nS6.���1k�@2t�A�9D����S(rr
�a�fţ.�*�F2D�P�b�i󠈃e�@ ��%ô�<D���g�]7h9h*"&�Y3��;D�����!Z^d�D� m? A��8D��0#;92r�qfk� ��a��4D��S�*�/!��y�B�f���S�'����+붌�.��]��AJ�'\9�h��1��-�0�,'~�b�'6�P�7-��e�8��u�K :ʝ!�'��BC�z=��+�*OJ0{�'w�H��H�w���`���A��'dQ��j޽�B��!J�\`}��'�^��fC�9*b����OU�})�'���8�\�OxX����S~���'5�t�t�C�	H�u��-��N�ɱ�'����%VW�A�K>`M�'�<)҆�HN�}��*X�K�'�&�QPl�b�(4��/Iu-��'����цۀ?�^�Z���~���'�\��gN�xP�hg��;u�*�'��0IVH�6o�F4��M��}=>,I�'��ق�b���$��>>�K�'��v�L1�����0(�\��	�'k��� �6IѢ9�陰%����'����y >p�dEA����'(��i�@P�6�>������
����'��I�։�2qk�9B*�|s:x�'�,���eГ[ ���-Ӳu���'����U�'���8�L_2uf�@�'B-)�'�I �ؖn/C�V��
�'�F����5ph�c��X0��-k�'���"DŢi��r�O�
H���'\B��f�*��ő���#��
��� ���dH�^��H�dS5�2L "Ot@�Q#ʆq����)l<��Y�"O�I�d��{RR���I�qK�97"Of��N.8�y;�(�MHF�K�"O|q����hI+"��5\�逤"OT���D�_�-�e_�&���P"O�I���w-�L���\�l���"OLX���!J�b!�Vm�><T�p"Od=���U��Zhy2�ƀ@:��u"O��!e0����D&:�P�A"O�M�2BV�m$dp�Ȍ#Ar%"OD$�s��>t^�r��^�j�""OΕQ���Q4� ��8�R�7"OH0)4`O�77`���.�>�P�"O��tCϿHی�A�����Y�"O���cfȫN�6��%*X<	z4�R"O ��1M�7xґ87��^]Ԑ�"OԽ9dB�q!���A�AI� т"O2����J �c5�Tr�4�("Ob�!��	�~��<�E�E��p�'"Ot�f%K<�̰��!�>M�z�ۄ"O~0��$��'<\ �� ��aÎ�z�"OP����ìY,�2���'�jTy&"O)1eg�=�N)��ށ,����"O\�"�@=  B��Mۭ_����"O�)�P"�+v�xy�����j�"O�%���<d=x�kǊP}.�"�"O�2G#�� ��*�� �th�"O�s/
.9r-�_(�%�P�l�!�D��p�$��i@�Qrq���%!�dU(�
=Q�{�Ni¢�> �!�Ė(z<��5����1���U!�)[�Xْ#!=����`��?�!�$�=_��p2J^#Fth\��N�)-6!�7k2]
�ɋ#6�-�pmɣw%!��i.�)�.w"�˳ʖ��!�ש�\a�`+��w-�����x�!�D՝#Hݠ4�J$v,��q�G6-a!�dV�c/PiHБg*:�Rg.�!�45�&�jGϺ[���@,�1�!��2xe�"�L}�AqIM�z�!�E8�v��ɭGo�����62�!��i@��u�W2N	J�{�b���!��X@�&��ԏ�T�x�j�U�>�!�dI�vy�,�)�;&���QfAʱ_�!�$�5i��Y�wO�Y������ƕKO!�$��Q�b�SFE��!%�\8��E4?!�D�'H� �PU�ל�$X/	!!��ЀrABI�E�q��t��nH`�!�$N����
<�v8ӭ	�+!�D�%i��M��۰vʹ4YwG�C�!�$L.!ߠ@H��޺%-	�P�H�!�DԾذ���������'�!�D��9D���lQ�I�� i�?<�!�U/^4�G��Z҅�[X�!��8'�,��R:ޜ����j�!�DO8t͠��s(�$>sg��n!�D/.c�|���W��{bF�Q!��,����g�]8�B���$,H!��(.�;���~�����'-!�ۀ? ��@�/t��YBA��,&!��6m�
�UϚ���IS$��y�!�$A$N5��0h����`��(=�!�D��]��̈@$F%��](�K�
;�!�� ��& [EB|�#V�E���S"Oj3�LM�2?�X��%L�8�L'Oh�D�|T^�QfJ	�b��ZD�T��Py��,b�|�+kEt3�5QԦ���y$]
K��'ʻf��q�F!���yRn�&KjQ�PA����	Pb��y��/�ĉF�ԅ[W���p��8�y�?~��r��M+t>���M��y�M��%	�P�W�?:X��MY��y�aZ�b� �hq��1���0E��y�!�/, Z9�F�^�)�$1[Ѕ	�y���T	1
Y�x�!'�;�y2�I�.�>M3�)θF����fb��y��>=�p�IP�t�
F���y���Yp
8���IK�P�v)^�y�	�.�~��׊oU��z����yr)��E�\�h��C1c�Z��O,�y���8< �Aӓ�l��S`
�y2��0�0��� Xq��Q���y���%T��#����
Ӥ���y�B5��=��
P:M>xmP����y�˛���� S�BY$�(���y��	�ȵ�v�9<  `cL�*�yB�b��9�b�C�/u�jw�ԫ�y��G�}������#=Z"e��A-�y"ߵ$f���׼3��遥���y"a$GZ��͊$~N9��	̈�y�k_�N�"Sc�����7���y"�[�d�|ŚЎ�7t�f�ؖ̒��y�%�+/H"� E�v�\Y�a���yb��`�D�:/ղiZ�] ��ё�yb�8��Pw���L�)X��y��N"9�&�q���' Mb Ѝ�y�ŌBv0��$K �����ɽ�y".њJ~�zDK(b8>z��ܧ�y�)�ti$82�ǻ'Vqs7뎻�y�.��qu.I�UQ�UyL��#��yC��h-h�ٱ$��<!�ջ�y/��t�R@ucÛ�� ��&��ybKA��`D��
j�	�S ��y��N�X�
9�fB�4�Z�2��y��^�o`*��d�۽2�F����yR�I�}Si���,g�]�-Ƃ�y"(��.���z%NϢw� i���ʔ�yªJ�|~�<��Λ{�n��G۹�y2$�!�>4B�%�g�tAZFN��yBɟ�o�v�PѬF�T5�yzf�^%�yrg�r\���덊U�,r���>�yr�L$R��d>��*v�A$�yB��+��� �`&��4�~!�'�ژ�vE��(���>2ҞH�'�z5�u��t��)t
E
#��`"
�'Ў���ώb�l�(�B@*p�صz	�'��U���R ��hU!��hcd���'A\���.n��FW6Z]�}:�'w��˷�	�R� Tn��<d���';��C�`9���aVE2K�J�#�'X���@��8]�(�F������'{�8	� �(��DɁ
i28�8�'��-kV��L�䙢�g�s�'`�A��lǷ8��3��2Z�u�'���E�̩�lH����:��Ĳ
�'����HXC�H�rr��3gt�C�'�f�`��K�wwb�;�@�MR��	��� @���e��a/R�� ��!X~��u"O�,��ݝi.<0�'�/�B���"OJ������B�(���Y ��5"O.�x�N�J��(QD]����"O�mr�Ό�,��q�B��R���T"Ozܢ4��R�H�d������P"O�0��*��S@�a���G}�b2"O��Xi��F6 �B�(?ZE�]�&"O �A�A�<Uh&�E�
�8:lL�"O�i�G]�L�ܕ���B9(�9�"O�#S�$g�	�SxP�:�"O��	��C`!10���q��Ja"O&�[��ƣ)�+)\!D��"
L~�<do�"{����U"?��!�FB�<A�d�M��A{��_��%�fJ@�<I�'�R�,�b�����@�2SNS�<I$�e��d �a��ž��r�Dd�<iB׃w|��3�F?ff�Az�[�<A����YX���l��:�d]�<�@��*0p�2���xA�pB�,Xo�<����_~L�A ԣ1]�)�D��g�<92�Z�<3:��QDݟ?�ڴ��H^`�<Q��S�	�^�C��=�2����\T�<���{ 8
!	�4�RD�r��v�<��;,}���Gµ=����u�<��jA �`*4
�]�"��E�V�<�t����I��̣W��@3eM�<���� �-y��!1��u g��R�<y7�)Ad�R���xL}�CaO�<���7J�XR��@�x���ǒI�<�Gf�{l69hd��N�qr��D�<��W����R�Ĭ��)3Q�h�<I��B��{���+B���"Fd|�<1�&QH�%�@�n{��"��x�<1UCZ&�,Y�O<�:��2��z�<�)Ǣ|��Xq�G�Ctf�j�AK�<a5�G�kC���!��S��1�.r�<)�e\���yy�l�-l���U�h�<a�$�=�|�Rf�փK�bq���d�<��mJ����G�n��JeLA]�<	�L�|��� Q)h��L!���g�8���y���܂9T^�ȓC*�g
��.��J®�[�FH��uXV�I3AѣW�����?D�j!�ȓ$,��`�N~��Z֤��H
���!i\����aJ�A��ش��L�ȓz������4P0�$9�ȳ48L<�ȓCJmj���gcjpH5C^����ȓ4�b�\�#��4�)���ȓc��y�BI����0h�+�f�^���[l8Ӧ�X0Y�x���B&Eb���?��,8��
�2�4�qV�5ܢY�ȓ{,\�@C��@���i��
�Ej��ȓYe 眠38-yA%ܑO-RM��@Rf9@�oO�l��(Z]���ȓy� �BaI��O1~�+��쥄ȓ��`�@^#�PcSK�?(�t��ȓ�3�$_(g�\}�d��mc>��[$$�7J,�ܑ��H8Pp��JR�E�r������`�+!����j0	g�Z�ij<Hv�J*,|����B�~5)��.g���g�){,�	�ȓD���&(2��ѐtjΡ!��(�ȓP�ޔ�2�W8T�6�xa��! �ц�S�? �͖�l>&BP�#>��B"O�e�᥆�b�f}�%��'���"O�	�u��)-�yb���<Դi�"O��(��ж|bR�dB�G�
��"O�As֣�el~���J7m���)@"O��1�(S'L� ��$���+��!�"O���D��H�,�QU��n>�5"O�4c䩀%^z�A��0^̼�W"O��Q$OG,��!B��ZE�Tbr"O��!����T� S3E;_Л"Ob�P�1u{��Y�ڿd����A"O��C�Y�1�M�<� �!�"OD��#e^�fw(�职S%��Z&"O�5�D�
���#��1#"O�hN�:�������X(�"O(P�ݍ �a�� �2�"�@d"O��2�k�:R�ع�<j�LѶ"O�����
;z�"���i\'V�hؓe"O�u�-~��lw:�"O�}qQD2�Ν�!�\Ќ��"O�yvcW�ORp��I�^Q>%�a"O SsJ�����iD��'��E�"O>�Y�a	�"�n}p�(�0�Ձ�"O0آ$��5��Y��D2
�����"O���w�َf� ��L�t�Ɲ�b"OT@%N �}0=��	�l� m`��I�Έ�>m
��߳���3,�*Y� "Odp �,Vc�\�K�4$���"OdU)q"��s���3�Ǻ7z�Q"O�$C�^�h-�T뀁.��"O�ɂBN�u�@$1���T�@c"Oh|#6�
@�)X�(	0�J�H1"Oֹ�@��7g(��#�g�H���9%"O�l[%�+~L>Tk�- |�a(f"O�9r�ㄝ -|��҅�=ʉ� "O�A��l�8?�*�`�$�=Y tt��"O���j5XJ�9�-�z!�"O�=�"_yd]���X%�Ũ0"O��Kb�SQPM"���`��0:�"O��2�f� *D��
�*"���"O�ً���
i�ڜ�D���33����"O��k��vN�x��ȃ�R'q��"O��?G>,�7(�*O���%"O6��B��a �PWg�V��P�a"O��hb��0��7L�Ax��"O�=�1HK=30 ��Mdq��"Oޱx�k�3Y������9Q�`��"OZL� ��H
Z(�r ��;h�A"OF	��b�!�v�sD �+ V�d�"O���1e�Xq�\�%oǫ"b}��"O�iHG��(]l�S,߃J��X+�"ObD�D��Q����<�L�x�"OD!06(ٗ7�p�Z�
�L,�"O�� *�Q�$�;0,T;4Q䍰B"O��Q� ��kE�0	A Qd��3"O"a���#f��#����LiU"O�Br��
a{V�5��@Ր�`"O����"Yz��B���fo��""O �ɂ�(O��g�� S� �:S"O-��#�t�˷OV�9���(f"OhY@�ҧ
9��h#/�-�tX�v"O��R-�<�u�% �6D�!"O�0k� ^�D4�S���_�%Zd"OLh̇�w��}�#DʮK�Zչ"O� \�(�)a�GÖ�7���a�"OPy���
N��2�� =�ƥ��"Od�! Kߵj�½�r�
��i��"O
Az�
X2n1��N���`Z�"OT�i�iD�ȅ˱�RG�����"O ����_�4�mT�7��IR�"O�	K�)�"�v��ĭ]�;��P��"O�C�ς�m��{cMM�\� U�3"OT|k�a���P��k�.~�J49c"O��!��o�0���WJ�i�"O��3u6]��HN2lȊ�;r"O���s��?;vx�v��k��A�"Ol��`�$t�@�υ*�ͯ[�<Qu�ۭJ��p@��X"%�݉��x�<Q�˪!�J r��$j��@ �/s�<9�I�?h�T���E#K��S�T�<��I)(><xZ�$Y��h�E�FO�<9C�ߎg^�e���)QҬ�8"ώd�<�A���������D��AHTdEe�<��v�t����D'i�E�PU�<Q���$d�D(�
��hN�u�EP�<YS���P��)�Dټ)��	���RN�<1�`�"tA���!S<Z�u��F�<���bL�p$�� �� ����@�<q�-S�C�*�#��O�!5�F�<�-ͯ7X@�Y��*g���V��\�ȓ!c�X�`�'�2@�����rYN��ȓl3�0��P�P}:}�D��@I�ć����ȶ���8�����.mWҥ����$��M]�c�NUʆ�L� >9�ȓsh�*��V�?fl��$��] Ȇ�Jv&���R ԘY�pˇ�M����ȓfD�)b���N��1��Y�`4���1�\�r#'��}�D0�w��v��ȓG���!��h��a�/�x�h0�ȓC�6${rOƠ���qaO˖�����0�:p$�ՋD��؆�"pd���ܔUNL��`̳��ȓ��t�d�	#��A� +\$�8��褭���=o����"O&�2���p+ �3&��j1�DY�e���ȓp�q�R*C79��ea�� n̈́ȓ,;�l)D��3�Ae�W��]��D�	��d�/U�Ɉd ���,��%�9�G'�9w����s�U��<��qd�+æ��?���X�P\�,�ȓI!�q0C��&�:�gҺ#�ȓG/�Ya�A�NP�7m�8M���ȓ�6�{k�<����/��H��Z�*L8�A[HK����Ó?H�(�ȓL���c�Η9K���*G�&�8܅��z���HſK'� 2���V�ڤ��c20�ƙ٤`i�
�/!4�ц����̜Tt���a?:-�ȓ/e`� A2���H�,������ȓzq�P�`��r�0[(��I_�(�ȓ[|���Y'WX&���� �h��CS��@��44�4��W�?Xt�Q�ȓ{�$�:w�B1�hYU�o�*��ȓyZ�&FJ=Un@��'Q�(�� � 9&�аW��C�<#<��Vt��Q��$o*H�/��8lx��ȓ	� Yi�/)Y��%e�;��ȓD������ٸj��X���͐��d��S�? ɧ�(�f�ZS�ɖ&;���"O��"�(��		0õ'��!�I�"O����+�|���ږ`��!�"O�� b-Q��$�z�����0"O~Q�Q#\%�y���{���"OH�yR��.��ӕn���n���yBk;+\Dx ��p��Q�reB��y�Ɛ�|Yc�I�d��%X�`	�y��<%��Y0%dJ
�*)��$X8�ybMZ� ����W�|�� ��_9�y2�]'4���eS�w���G�'�y2�N�6�ژB���Y�<�	?�y��7�"�f�R2��l�7�I�y�w((��� ��\dK��y�w�y@"!�3}9�Ix�՟�y���8l�4��q�
�e�Y9�yRLK�u2DY`3K ����jtJ��yB�'�a�6�惡��	6C�\PROE�1�^�p�`��v�8AЂ��J1�,X�i6 aÁ��Z�k)�sj��U��\vn��0�� d8;��i���A�m¥Cs&��@"���I�A�'��d����U1Tx0Wn���4H�O��Q#�O��lZ�c���<�������N�Ókŵ�e2�oߩ	�!��˱�欳b��#��v`ѫp���شT��|r�O��_���%F������?(���!��5J�@�:�ƎJx����5l��5;�#@u:��qB?`��p3�DM�C�.M�jڧ$R�`r5.E�T&��P3�/ܡD��1�IF�I����*��4d��QF+ÀK����,��m؈�d�2Z%��\<����0�ٵwְ{�cOKNrQdm�����<�im�O���'z@��C�΁9Z�\�TK�;y�ȓQc�4�E�=x�~�1E�G����Z����ѳi)剉y-,�j^w7�����~	^,� Oi�~P��ʀ��'>rH'K>��K�MPo�R�Eߨw?�|Χ-��P��"�MՎ�EiZ"<�Dz�a`hhX�<Xg�	�g
5�擮c,)(SKF�#�˞�v#J������|���O�'>�l�%z`�!�"�5Y�bǥ۶\���������:��F$�>z���rD����I���O `lڹ�M�ش;���!c���p 醷$3> a�O�!&"���m�	Nyʟ�O��&Ĕ{�8�sgMT��V��=I2��4�J�
��ׇK"^T`xr�����7`[�s[ū
�2	�P�@�.�M��źh��!�����u���Ug�-�~�|�1+	�d�GJ@"hv޴��,v��o�,�����O:ym���<D��4t�n�A�
H�Qs|,ۢf��p<�}���?	���,��,M�����6l����=}��<)��i��6-4�����(��"ڪ��)�D��C�ax,O|�pȂЦ���&I���T�>~���d�бr�����2u�L� ��s#Uf֦�d�$g�M#�L��jTBRQ5yV^�b���m��VQ4�!4]N�4"3h�[efۜD�F#vk�$�Ji8��'l��I��'!67m�.��Y����h}��_�O#
�@�o�jFƘ1q�V��y�N
+4J��O����,WK�|l���M�K>ͧ�
(O��l.dT
�-}^PEx���D���&<OR��!!�Ea��˼q6Q�*#-�>�S/�DpC3֨��!����OPp�s1�����KB�>f1�S+ V8��A\��P�P� ܜ�G~����?���R/IIX�z1�G�a^��9B/!+߆�"D�i+�\���	iyB���/-�@�NL�H�����,�!�8��`I�A������U8?[�����i0�4�䓌?���ēL��H� @�?   X   Ĵ���	��Z��wI
)ʜ�cd�<��k٥���qe�H�4��6X8$<gT��"�ᔩ^�"u�ǣ)z�4�L��M��i�Z7-�Vx�,a�K�[����݉a8�-q��D�Q_��b�iq��a��	�"��6��Xb>:5H8:�UC��Ǯ���Q�Mx�ݴ��	+hf�(r@[�剟R1Qq�#2�HY���:K�De�R�RT�6�[�;����mbm�cΉ>�l�y�t<�FH6���Z�(8C��<k�H��<������l�����U�l�Hu�O�	I���^���Öo���AB�Oꅡ��N6xP1O��t��	��'�^4��-ԒM��1��Z���'"B�Fxb@�W�'r���O�W�Y��@�+g5�&->�9�Z"<�#G�>Q��d�>x�ÎL�^�q v�FM�d�OM،{���P��rg(Eg��W A�M+v�(aŰ#<3L6��
c%���\�Q��Z��Ȝ�>A>�y(��;J�*#e�}���)t��|��'���Ex��A�����l����kR@J�-�,|�!&�P��#<I��O�x�r��g8�̪P��9L����D���Ot��H<q�C�f�H�"�0��,x��^@?)1�8r%�O,�&B�U�M��4y��	�-J���
��IgˎL9@�$OHi�DQ�O�l���(��S��LB���(t,L�/O��9#F30b�'Vp5�� �ēB,�����u���xS�A;+]$�+��/��$GyB%�M�'�����	�`��xH�&�k��X�'R��:@ ������iC�	9�x��ٴ:z�Sϟ������KfJXYcC�ZO�qy )a˛��'j�R��|B[>	��RL�Y+���<�����o"qG�pn��U��m��4�?��?1��qV�'er��v�"��-�@zX��¥��".7���X��d/��|�'
"-�9HI�@�cD�w�DT��/�W#�6-�O��D�O�Q �j�^��埌��r?!����ۮ�8t�ǀp�A�rm�צ�&�prGN�(�ħ�?���?����6*͚���/Fa��/��
B�V�'��L�v�(�I��&�֘�Sv���N n;�L#4C�'*:N�xP]������O��$�OjʓF��a1h	8� �ŀ��j�.�ZHTj��OT��8���OV�%&{��b � �|>P���OT�rN�g3Oʓ�?���?(O��r���|J�D	    �    �  �  $"  d(  �*   Ĵ���	����Zv)Ú'll\�0R�P����=9pn\�Ёba�#������{�<I�d� �t�Z5$��vT�aN�!@ i®�,]Q�����E���I�A���0�2rTƌ�&���L�/xP�A�^�M� maf�E�m�];g�0'h{G��PZ��xv�Ӳ]m^X�S�a���N�y�D�{�e�>;P`���H�F���_<k��ac5���0$���72>���)�-#��d�O����O�e�;�?����$+H1p��Ւ;o|�ԫ[�gS�	`'&��d���A�4L��HR4rP�шw5�	�6����0'("ݑ�<J"��V.�> �ɕ��<\O����(��@*@9����3|r:�"O���$��A}�@85A�.� ���ie�"=�'��+�B(�4��f�D ��,����4R����%+���?���?�������O6���*!���S�F�j�/[�`��p��l�QЊ�0c��_�Zz���[?Q�4�U&�xUXv�վjxƁ�3�:J��X�t�M�W��Q��`�S�'��QJ��gl6�˰iE�|�2���lB�vT��t�i�07�<�I<�H���LH0Yx�P^� �C��y�&��*8�����ɠ��Ƅ����JM}2P�H��G�6��|`���L8�"nӪ(�6�\�g��t����)w�^�"�"O(���ou�J\(^�12"OJ��g�"L�x�&���{pj���"O`s��]�hZǡ�=
TZ���"O08���̹)�y(�B9M����"O~�����q>� �eI��vr4�"O0]��,�a��ə�\2X���"OX�r��4W��Ҧ��;>H��B"OB���#�m���Ah+ [�"O�H��ݎh��8�t�(�(�"O��*d���l�J�qAhU<3�b�Xv"O^ݣp���[�
�ɣ��S�"OZ��N�e���5�va�Ivl!�dV5��@��� 6�bA���<!�dK�XmD�� ��[N�,ru�ߟ !��G.u��ʷ���a�p�ˎ�*!�$Q�8�ZK�d�h���F��1"O��XD@ l�:��P0���)E"OX�Br�]�f�^���@�~ H(��"Od��o��(��smN�s"O�=2RB_�pʾ̈RΏ"QFڨ��"O(���Ǧ^T.���c��_樘`"O�\S��[�+k�D�0�B�PSt��#"O:L(Ҥ�K^d�z�g�\z��s"O@�tH�V_
�qD���9WؕpA"O�}sr���f�B�\PҍZ�"O<-��X8�$��G�8�.���"O�)#7�ғ|+Ar�%J�Y�p�"Oּ"���-��jZ�u���"O�@��eT�l���Q�)�#�=!�"OH!�d,����I�M�cp5��"O&@�Ť����9��3G�F=@�"O^���`�n`��{6 Ʒ<xn��"O���r.�/5ĩ�&6�� �S"O��4��dP w�� n����3"OD}�ag�[U��ҷ.]�(���ir"O��	3�@�0&$쓒��X7"4�"O� I��ء.��q	vlThB�1�"O����_/��#(:�i2"OB��q
ɢf��D����}nb�Pc"O�(ڇ�#e��}`Ҡؼ4Zڵ:�"O&���k.4^���PO�u{Q"OX��.s�a�T����		C�AK�<Ŋ�;����_\:�5�d�K�<�7��n��)ǊR�H�(�B��Q�<�M� bfŹu�Q�Cm�Ty���s�<�&	+!P��d�@b81��ər�<��LH�0i��js�˘4m�YjW�C�<� :�s-rXEa5e�?�f���"O `0ǆ D�����qH앰�"O  
��9����0��\JJ�J"OΠ�&i��`\�9���$i��l"P"O^�
�$� h���7�"O2��aȭ[�`Q��^/#�~�x�"O���7�3,]�̃��t�P�`�"O������8���ԯj�����"OJŚ�bL7������(@ʕ��"OLY�qf�/-���U�!8MH!32"OL�뢏ɲKg���!$S�;����V"Oz`P���'�U�7�y���"O�H�dFEm�b\�g�� k�p�"O�`` ���m��9Y4��[���11"OV�iQԒ{��`s����D8�"O$��k�v����E����q"O4035��T�r�Q�D�5HF�y�"O0���V<oE��(�˝���"O�(�s���^��Մ�=�ht(�"O�|�qm�!.��E�檐�b��t��"O��Bc[�&A�D�1�#?���"O��´m�1e*�A�'[8w�NU8p"O�]�"@D�hP^p�f��P�,E�F"O�$�֫.�2��֏-���r�"O�a������X󮆩^�.���"O:��m�w�9в�Q=+�|!C7"Ob�r$e��f�Q-�N�r�Q"O�-R�̭t-sFX�d��u
#"O4 ӣ�τC��8BP�P���"O����M�)9�Dd{>Qr"O�`� �3���fĕ2q+��@"O�%*q6�1����0�"O�Q���Km�ő��D�	0���"O�0��
ӐU�4qG.7vd��"O\��nI,2�����?�^�Ia"OL��6�ڨh��摜-�=�S"O�6��?�$��EN�	r$Ð"OxH�Ʈ��z\�kT"�4}�ܔ#�"O����a�H�ٶc�F�90"O�L ��J�h�q���?����!"O�(Yq�1Cю(r�$��h)b"Ovi�Ə˕G!f��j	��d�a�"O���I3���G�@��A�"O:bC�+/z�#F��9_��M�S"O 8:$#����QР��woB�@"O"I���իt9�,�N	&4z죒"OV�sB-E-oF�@��B'j$��37"O�Ib���c�l�3�E��w!,��"OZl����Z��	
"Κ�X�� �6"O�q�BL�~1����/H���@"O�4���H��=s0͖�d�J�0"O����	^Ď�s����.���"O(��j�I)��&�._�،s�"O�$X%�ީ:MNm���%j�~Ő�"O��V`�'XY���b�ΨH𠃃"O�ȇ�&*�XmS$�5,��"O ��P P'\Y�\�$��Xll��'� t���'SN��F�J�i��t0Љ�
��qד�u�eO�"����y���Cf�Vbb]�P�>[!�D�>GҐub�kM�(bN�3�E�_��'�N�1�M�7#��q �r@�����>�x�2���C�	8L�0������%	p��,��n�����{�
˓��D9��L��2��->�����bU9V��t!��0���d�� �z\����t���%��1�	�4��O!��I�I	~؞� ���&G�vXtqr��<\��2�'}�Hb���=@o�q�G��'b����n�zESѩ�c�X��eM6�y�A^L��iu�l5�)�K%���lXj�Q ��.
� jăٳ�(�N��݉��T�#� ,�¤�4"Of�p��̶'��8��w_���n�(G��my�F�#yP�x�]�l1�1OVMS��![1��:R曨؎$���'�VLQ��cǢ�`�
��10�C���0(�l2r$
)6/��)�T�az���&/4�3䞮Vfʉ�A�	��O,�JԈް;:Z�+#f�|���R>{ CF���9ˊh�E�Ĭqu�B�	�&�x�y�E(ҬA��!)���- TI�E
P�q@ê^��dӊ��F G8`b��J�v`F�P���!��21���;U��E"c.�.-�M#�=a,�QkOrfr�PԚ��d	 z��	:��'&���$�w�rh :v�(��M��>��	�Eݎ�@I�"|��ejd��8  �q[��'h$��e^<�AK��$�>M�Óls�آ�J�E^�!K�aC��Y[�)�.\ )�M�o����#�M�<)G�R�}��1ah >b.�y3C�M~bZ�x1G�
�2�.$�$!�'^���(vI�7� ����W�̵�ȓN��a��I�-9�J����C�Wg�H���ݐ��>����O�u��aB�=Ȍe�e�i!�`B"O$��`�1)�"� e�ҷE1hd�Ʒi�:"�F$U �P�
�9�$"r��6Y\A͜�&t̬��+a蠘�Ԍ���yrHG�k�d�����W�F]�U����y��g�ȥ{E�=قT�f�.��'�D���C�F�"~�"�=��M��	n��@�3n�B�<��KmR�a�҃@V��#�W�<Q�U�Ԟ|�GX����R4q���pÓ%�z5�3i��XT!��AՐ Vǒ�ܡ�oL)}�RY!"�a~R�@�����[�6���f�ݩ�yB�]�S�~�H��$\x&l4�y��ɡ�ʈ˰I,X|$���y���U�b����i,��q����y�,�?l�nL ����6T�@�ޠ�yPs^0�(��U ,���y��'A�I���H<B���P�ώ��y�A�X"�`�cY	z{�g�
<�y�G�"Wg\Dx��7t�"���/��y"!�4z��$�n4��9�(F�y� �h ��4 ̄l�
e�R�߻�yRϙ3��j�'ϻi�rJ��y��?3<|FiҮn>�U�P��1�y¥�4�"��6m$9�
������yr��?&��QIŢ]6crrt���T��y�&ʼzĚ<F��"��=�Pb�4�y2j�1sԱ�׺P�կ�4)
�'�@]�v��1��-��Eϖ)4����'S���hX0�L��fK-c$�:�'�l�@��f"��D�%N$ ��'p̉�O�?RLT9�U 2��yA�'�+cN (�`�t�F;0��p�
�'�v�X��=j��hC��R.5�����'J��Qю��dE2�z�L^�;��M)�'o�	��L�=rt���I�$�^(Z�'��!j�Ϸ^*(�� ,H)VE�'�VH��ݮ����q��y:����'��Q򋞷[�m2�fB�r�.3�'c(,Q��Q���;��� �n%��'�F�����f��Qz��Lʶ�k�' &Ы��8�2ё6蒣qߎI�'!�-+u,K5��Щ��Y`��0�'Pt�)���e�4���9N Ti��',&pY5��/���W@��@[r���'���'Y��6�P�l���'�I��-�"N�x�!!F����
��� j�Gܠr|���F�	1lP�Ц"O^RD	�d�UY���u
����"O��P�Ë�#JZ���ɻ-���6"O�ӳ@�\(e��"$�A�q"O�ؒ��Ƨ>_���������Q"O*�S�Z�V�P��@�1`rF��2"O��k����󬑙hvը'�;i!��	���-G�{���W��8~!�� �pP� A.�:~��8��-9`!�D'?'�$11�?q�*pk�J]�nI!�D�.hBJ��r�M0�T=;��W��!��%6���&�V�C*dbQm�3�!�E64K:u��c�8=`��#�Ȟ�!�D�=t=���6U i�N��2����.2��y��R�f|�6�O�y���dU���kX��ָ(�n�=�y� ���O�4[m&��PG�5�yF�4A*Νٕ͈�(&�� ,�y9���I�*�#O�j;�hÇ�y¦�1��a�AHԌ�Уϛ��O�Y7Kb�欙���]��HbѾi5M��m�E1�
�3
͊�X�'�Ԩ��;�)s�Ӆ*oL��'���c�Ͳ,�� ��-}(���'�z��'F�_�*<�2��%�A��'��|ZW��Z��偱CC�[pE��'o���Qň9�x�� '��'�<�
��)tz� P��ˆab	�'Rr��Ǆ�,'�+6-��J�B=��' ����.uE��8v�<<�!Q
�'�R��PkɕU+d��5K�-�~�
�'�l����R�|��e�C3J8S�'!*�c��<�B �-k�j8"	�'Z�Q��
J��VBB;n��x��'������y��d��L=O��x�'�v�q��
 GF�zv�B@P�1@�'h��s��J��N|9�������'v4�PC�n����~A�!��'?��6��u�RQ����}��Q��'�J��tj�Q���o�&���'5�xaF�5b�\(��W���X �'�xu�!��U�B9+c��!<�	�'�~�p鋑{�\$�A킎���ʓ�~� �˃2jՀ0&KR���ȓp�	��6,����E�� ��G�L��� �!i������ȓ{���.L{a#�o�P`�ȓ!G�ja	!xNk�O6j��@� �b��B�`�ڄ������=(��u��)��z'��v����)4:�0��ϑqS����=�ȓj�(uy�c�%�Tm��='P��9�f4�#�U�n>@)��\��vY�ȓoOڴҤ�<ȴ�P�
2R��ȓ$W���	�3]洼(G��]*l�ȓP�X�J�AJ��`Ո�DYFA��}�lȣ�B��j�8��Q�8����ȓ8�p{�N�>0��˕ PA�`���R�\I�%M_�/�jh;�,���}�ȓe���b��OB��mb�mSbOb`�ȓU*T�uȅ�g�Ș�2�kA\�ȓ	6� w*�$H�V�����s��8�ȓV;F��P�hRtax�Ǔ*��5�ȓ�Ve��)�M�E�P�4	�����Z���hǷB�5#ײz�<��S�? v��3�B�ɁA'�d�q"O�@�3
A)/��"!S;JI���r"O�iȆ���/R �aMΤ7���$"O:��,�(p�* F=b��H!�"OP�
pB�جx2%�T�h�.��#"O��؃�F4y^��I����&n(��b"O:��4'��*/�J'��.zp�`�"O�8������#ł+ .d�5"O|����N��i����2�Q0�"O��AN�.r�>x���>���"O�(����|�E�'�q�"O:|�b��Bu�H�1΁%�ޥ�U"O�%�#Y~z\jvL�>ڶ�JV"O"��e� W�~�T+E�@��f"OF]�VJi�U*��	,$����"O�}w���IE
���T��`t"O����<�$!I�,�q��"OD��Γ)O�tq�E�^0�i�"O�5��$��4[��:�Ē�F��PS�"O�A
�fA7�R�1wn��t�� A"O܈d�&�%�DQ�ģ�"O��:�)��L?��q` W�2E0�u"O������h)�Yp�N/l%Ta�"OjBF��+
V Bb�je�b"O2M2�ۼG�<����^0�5�"O0M���35��1�É3zp�h"O�����."0�胠Ə2@|a"O��p��߂xH�e���WRX'"O��h��D&r����u�ǯN�B4"O�d��Gɜ\��1��Kn�6�3"O0�@Dm�(r5^�*2�Rz]�%�A"O]z�N	�8�t�g�kW:pQ"OT4��Ǐ=�f ����	J���"O�= � �n��l#�b��V�t�7��h��D_����`E@!6rAb��@)ny!�䊷9�	i�C�
	�Qc#Z��!�$�5c�AZ���k����Q� i�!��5�u�"�W67�.h	ԋ�%�!�Dʪ\q�13�ᕮ��=
�
D4xG!�כY��ɉ��L���� ��;tW!�$�JP�hA�DG�~�i�R�� 0!��1cm6�"7��u}JY8M8Nr!�d�g&a"�*CRRYH�@�)�!��-��JWc��\;�)jvJ�")�!�$�)�|gI��A�y����!�$]Xn�0��_
4�vfo!�䗯,bZ�j6,�?a�F��^�T�!��V3��5�R�A����s���4D�!�C�mf( �@;���X���1OB!�ڞ`u����II6��ń�94!��ݯ�vC�⓺C1>�@�m̤1!�DE�^�J8��!��J/`u	�m�(b�!�0` *���Ė <Y(�͏�A�!��* p����P.4�,*��[z!�
�"L,hڴ��N�4"����.G!���!�� �Y4	^�IEJ��P>!�Ȫqm�:��7B��B�oݣrN!�	-� )�����]����o;!��N��x��T'*�Hp 0�K_;!���5M;n��k��ȸ��KƯ
	!�$�<��}H��&r�B��k�)\!��Š��FA�T`���e�!�^��\A� $6�蜣��O�>�!�U�.��do�7ڀA���V�DF!�� \Y� #�:d����q�N��e"Oڡ3d�æu)*�G7�
T)�"Oxp+�.�<�`�6���>��=r"O���@ Й`��]��@9]{|i�"O���۟��ժ�V-m&�!�"O�XȢ����Dr��( fܰ�&"OH��vc��C����bMF�y�E�"O�y� ���i;�=p\�{J�a�"Or� �cڣ"X������?:<c'"O����{�l�s,�F2�x�b"OV� /	� :��!���&>��L�f"Oܭ���%�u�ː:h�@e�c"Oڥ��`�1�a�#�ؘ/�H�"O���,q��y����%ea���"O.4�#UrK|� �J ����%"O���3h��VP��h��V�n���!�"O|)1�\���|�ӫD�?���"O�`�b�q���f�V�:E �""O�]��E�(Q�Tj���%`h�"O����!y�`�+|�r"O�dCq ц?K:�J�$>��lQ�"O�R�-ƖK\����t�,)$*O<h1��\�j�:DE��ex"�{	�'�{�lO"	� �#�a���'��٩�G!6ot��A2�5��'�r]� O�A�x�1�9 �'���Kһ*Jhad�Y�\>X�*�'��b`��L��=Hs%]�%�V4��'��x"�]�%�
ăR�%r*�-;�'�p#��2W��� RLg.���
�'��gN	"~|1a�׭Yr.(��'�􌩥 ў4���(S'T6���'10X`�C�	��񪶤֜S�B�K�'jڴIF��
WE����AB!%�X��'���$ڂ��Y�H�z1��'��}���M  rf]r'�JE�^-��' N�� �4lL��0&*/-,���'���L�]qDh;�͐�\��'�T��,�<rЗ��-*�����'zH  !t86����&K�!��'��qЅ4$���I7E4�i�'^��i�bK�&H J�Ϙ	Qh,�'+�I˅m��1O��
r��; 2n�P�'�ҽsTf����ؒٹI�� S
�'���`E�!�l��/ےB+
�'��F���a Pc�4w2��	�'Ӥ��@������GO��].���'	,�:�`CH�� � 
��0dq�'؍ʡ+�6"�&�PCn�,q�EQ�'[�-20�\�6C~A�E
l���q�'6,���@2�AQʖ2�|���'���#/��f�R'�b���+�'��zbIˇ2�f��E�D�]�ԋ�'<��Y�A��C%��$7lT��'�����\�j[�U�TB�2@��'��)(���2�����E�}�0} �'�P�����'�0Q1ġ�.L�C
�'}.�����#���S�öP����	�'���+djL�s(9���������'L*ܙs�_s�b��e��2!��' � �1�@O�!qAOJ�
���'8�=�0"џ_���"b@�O�JB�M@�Q�F-�>͠gC�t� B�I�S�8)Z��5�]��,csZC�)� ~�8gM�1ڂ+�Ɗ�7��PCD"O���e��UFQ`��Md�2"O\hg	O�>�(=p�f��	��Yt"ON�cB��[sl���D��9��)K�"O�2��S!|��
D%�����"Or��bE.V�(s��ʿ�eX�"O�āRD�	"� ���t\^!�"OD�[���'$���E�;=����"OB a�R�� d�<���_�yB�B3F�x�Y3�\�&O�u ��y2�M���U���53���*��y"BD�6����Zﲥ)�ʪ�y'�)H��2���L�F%�y�`ܹn6�dqr��G�H�����:�y"�!�AzS �II���5Ɉ�y����F�h�@"m�E:�)��yIΉ�Fy�`a�-�� �C���yb$�7d���)-{P����Ђ�y�o
�u����$�A�i;��`�cy��Ec����bۊ ~ ۶m]'J���ȓ(�r$U�^- T��Ц&U���ȓj&���b"V�|��H J��d��q�ȓYEqЅ��=4�{�B�ì@���DC��޽|x(i���\j@	��[��X� @�?   X   Ĵ���	��Z��wI�*ʜ�cd�<��k٥���qe�H�4m��_;:<u�i��6���K��=�3g��2�R�9AfN/>��m���M���i�����P�O̚�+������ch�i �o	��M����O���4]�B|S&j��.zU�VnR�q_0��'&Z�Q�����݁-O�p6*�p�6h .O�)�e�Α�Zm���
9HfE��$$�4��4M��!���OZ��E�&�s��i��L�6䨰*�3�R4��GT�+��1�nC�
��ɯAhl��j�th�'�����)�~�f3{��T�u�0Pd����k��~�O�PC��J�yb���GBxx�<ID��%��l¤ �P`���<�%� '��"<���E���˖�f��-�!�U�{P�LɅ�I�)F�ɊE�:�q02�*��En@: ш�'���Gx2j�Hܓs�A��&�.+��{v��4B܁oZ��0���8F�޽�(�(W�б��	+2��%�	�L���f���cq��-Y(ȑz���5��d"q"�<�@
*k�⟬
SB�#y���ї-vhV5�6�0��ܠ��	���k�7<a��n��#�|<K��ܘ'|�Dx��Cp��:-"I�����y�j�'�Hm�f��"u���YT�xB"��P��g))��9�'��L�Y'�O�h�'�NxD�̜P��'���fDM����ݾ_Y2���&ͨJU��3c�$��ę:R �Q��D��j`ԭ�M<�����8�L�q��:�p����J}bh�s�'��Ex��a���0�zpH�Wo���y�@4. d  ��D���<��С�'��(=+��:D�X��F!��,��(ə�DJ*7D�İ�����²BSw�LЇ#D�쓱C���^'!WCF��$� D��P DP9�=�ԅm���s��?D�0�4�,m��S�Nl�~���;D����\,Z��:�=(v����:D�,q嫏	m�� aMF!�r��-D�0�R#�cv u�b��8rԂ���)'D�p�J��e� %*�-�5C�D����%lO���AmB� �T��[�6�ˢ�-D�t�d� D@6��D�e�8EO D�x�@D6r��!�i�<P�Q��#�O������$�&��3����ik�	�ȓ(T�{�jB����tj�-�^��H���B��l0� 0Ɓ�+��u��S�? ����NQ�:q�=�&"C�J��Aq��'����{��w�J$?*���-D� �W�,'hQ�0�Ԩf�Ґ Ǫ'D�̛@�-�|C&ћ���p��$D�8ʀ-�#4J�J`!�Z�j0W�>D�� �W�]G"X���X��@��=D��k�cǷ=:��Fb O���3�1D����J�&�R5���18��e<D�\�i�h(>�9��ܲ �1%�8D��{3	μ ��@��)"��:�7D�� �Ņ��l]!�,�F����3D�ʶ���H@��pZ�P�1D�� f��;���M�(	�x�%0D����ir��p Z!SQ�A��3D�,#���3���c��k�na
��.D�`7��=���ae�Z�M[���ň6D��97E��X�y5j̉sVdM�"*D��5K��BN�h%E(NZ`��4D�2T�S�L�ep�G])Y�8yB�1D��!������skU�P��e"D�|p�T�S�B�%�!�B{�?D�ظF��.U���r�x9��2D���Wѩ!9��hd7��p��/D�$�@�̢y����Ԩ�DkP\E,D��#"صI%l�x��JDA-D���/ �^/
	��XD�0�`��8D�P�D��5�2ᱴA�?|�¬��d5D�x�n��^�����K"�X��l1D��A40�"�E��xk��F%D�p��lQ>	O�Ə{�H,�6Ɠ�y�%͵ �HU�B�ۧ��Ǭ)�y�ɑ�7L��tb
#L��Ճ1�y2��#�^U��הE|"�<�y��0�Ba���P�l�
�J���yB��XF`�c�eƢe���q�:�y �T���ן-L���,�y�&�+ O���`+Q-P�bM�q���y�"R�E��ʕ���@���{�M�y�iΨRd��&i:$�nmK`V��y�ֿz-�ܡ�X�{�G޲�y�픅
'V%�Q� ��  a�%�y��¸ I��d� &�7o��yb× 4N5����"Z�x$�� Έ�Py2�E���Qu.Q�i�C�Q�<�R,�nmbcj^�!RHyv��c�<A1�*5��V&�#
��3"A^�<9����|$)fU�5W�!b�Y�<�T��N%t��B��6�ҏ�N�<����?�TaI���)W
D=��DQ�<�GBaz�a���V�0�f8v�ZJ�<a�D˥\Iۖ$�DAn�P�aAC�<Q3	.���5�v �R JH�<9�+_Re���$�!s�&x��n�<�!dȉh4�TdF#�bs��k�<i�m�1�I8e���R�xe򖄓@�<�v�%�,���#�����~�<��!zlm#� ~�n�x"�}�<�T�_�1� ���$�ŋ�Q�<��
���`CQ<p4��A�GL�<3���O�0dfE�L~�ɫ2��|�<� 3�,-�C��t���a�<� �α)�R4�m�z�q����]�<!׫�&,&�XB�=5���'�Y�<��,G��0⥋�
ar�7ɕ��y
� z����l[���aB�8G�Z4��"O��bJFFbU�/I�8N&x�g"ON���O��3���1P�J���f"Or��"#$�H�l:�H9u"O$�-	4>M�Q��
X4*�f�;�"OT@p��!��q�
*]L��B�"O�tx$�]�/r�b��O�
#�<��"O��g�'�<Q��&]ijJ(��"O8���A�jtq1oDK�,Ju"O਒�.:mb8`� ���1��٘�"O�!�#Ej��C�ES"����"O$1Q�,WZ��׃��QvZ��3"O�ř�(Ǻ"h�M0q�ķC��a�""Ot�� �23v�"a�N�i�(���"O�l��M�.�6a�G�ڡP��[�"O�Ш��ŷYֈ�2$�{cN�D"O�$�������É�)y���"O�!�dkO�)�������)hV��e"Ot��v�	j���Eem��Iۇ"O�8QC�E 	�eP��ܜZ[~�u"O���֧]� BV(~HT0sC"O��h"�2��؋��ư5D��;�"O��qj�82mJA���>z��"O��z�է1�(!C�aױs�@A�"O��;r	�
z�h�V"ӔG���"OP`��m�X�*�S'a ���"Or�2ub��HЪƃp.�� %"O���,M|�=�G.�/P��)�"OjH{d'��v�z�	AHӌw�%j�"OzQ$��A>~��p(�|�fmr�"O��:���$]�*XN��j���!�"O�c�;{9V���-_�e��i�"O����ɍ�_t�]�%���OH�ag"Of��Ǒ$ƶ]��eJ�SEZz0"O��1��&@vT�����>s�xH˧"O�E9�/��J�r�k��΁[� ��"O"�j!'Q�
"<c@��@���i�"O�Y�bM�nʩ�R��?Q?��hb"OU���_��+5�D�I\A3"O0\���Y�l�+V���%N��B"Ox�C�n����X�́pf|��"O��#�A�|U�q,ςg]��[�"O̴pr�D�X����$")pX�"O� +��+#�t=P���`?p(�"O^h����(a(�h��
K8�hr�"O�a����'cu�D� ���:E����"ODa;����3d ���T
O'.��A"O����B�4c��6�('$��2'"O\%�� Q@��	1"��Q"O����f�n�Jj��<\x!"O@��j�>���.Јl����Q"O�����3qrDhP���r-�d"Oj�zDX�%�J��&�͙f���2B"Obi1`O�H��K�I%%�� #"O�H����Z���Ti�4��!�"O���$D��Y ��[�Q��P�A"Oh��K�~���Sfܔ�~e��"O��b0`A(kz��@t$Ēn�=�$"Oh�`����z���L�Rn�ٲ*O������q�\��� #Q0My�'˪Y+S�ϋA-J؊f	
n��i �'P�d9Eᄢ�������mn��;�'O��9����L�
!*��g�L��	�'���:f�!^ʼq�NŅz�aq	��� �(���/���h��Y��X�*Oڨ��hF8a��+��	cH)�']b��Z�B�H��g��tRh9!
�'F��PPK�̌��7B=A 6 ��'9̅��ٳZ	(��w�D7JII�'A0�("��7H��0����7�b�s�'��#�	V���рWCC/,�d3�'���)��zF��v&˯x�dQ�'��+��A>X��D)�"��>�j��
�'���Ƅ�MöDܝ.�EKa"O�E�e�:wږ��"#%z��"O���%��X�Z�u�� 7"O>	��c�O%�#gԥ��YB"O���gȬ{������eU��`�"O��a&`ƣA�	�a��Y.���"O��§;���aT获m��� "OV�D�>���R�D�� ��$ B"Op��F��9*	rё�����6"O�A8@*O'/m��jD-ɊBZ��p"O*�D��@���1���=v �)�"O���C��B�:�TEB�ec��"O��`���V��9��Jj�x�"OсQ ˾UC%� 0��"O*��9q�]��ŉ���j�"O�$yD/W6{(M�c˟>�*��w"O����/B,���A!A�x�"O2H%d>���rV�;��$�"Oz�@���&n��
ġ6�4��"OX����ɑ���%H3({����"OfA��K-x5>�Ն5`	4�"O�A�V.2+�XcD���Q�P��"O�����Q�*oؼ���S� �~5Q0"O���%��IAtQ�&N�Mo��i�"O�T3#)H�o Zi���?hp $"O�y3-ܸ

��#B BIvp["O���5GQ���l���Ŧ4=P���"O����n�?g
����!�� :Blr"O\\�p���fe��G�0�+�"O^,p�_�B��c�?��!"Ob�SlL����xW��f+.�I�"O��0HB�@�K�Z�4�N�3"O����]�p"�ԃw"O=׀�D`�����R�̜a�"OrC鈼d�DY{B:6�`�k0"Op��A�*,vVQk�jW�zf0�"O@��B�Z=]�zU���2E��H�5"ONiU%^3'��]af�B&����"OR	ks"��8����Ei�p���"O&i6fH;g��Wg�1q�0X�"O�T��8r�m���f���"O�H��U�'CH��Goe^XXC�"O�0���p�����V�o#���A"O4M�S͉� ��U��Avf���B"O�expa�I�����g�"c"O�(C�͞�@b��2��6AL4��u"OrL��U'-׺a��OHl%�Q"O��ʷ�L�&"~m���Z�|>hV"OJ��R��	/;�@:A����'"O�3���?4���/�����"Ob�àOMߔ9��g
0�X��y"��e@I*^= ��0f��y"�U�5`�
���(dZ�IwD�y�N�;1l����IH�6�bi�5����yBiY �K�d�YTH@';a�Q��S�? \}�2�8DR����IuB	{�"O��1h�,@;^�A��L5^��Ȩ�"Oc�;@�,�B3ǌ2N�2X��"OT=;Q��l
&Y��O����F"O�d��%��,���d� �p�"Oz��`��
,jz��������ɧ"O���`N�u�LE��!�7��p��"O�e�НiƄ[U�	1d��ȋ�"Oּ���?=�*�B^� �&D '"O����z���A7�P�~��$Ӄ"O�3eĝ�hib'��z'>�jf"O�)�󅋦B�>�SR�ŨoT��"O��#E��j(U�u	G(p�T�i�"O��b0Z�C�t�R��,�.���"O ���?Qh�1$(�.ڄ�3�"O�  0b�G-�M��c��(c"O��#�IG���$ T$�)�� �"O,�p�uq�(�u���A��̹"O���4;�4U�f#(8�R���"OH(��%V�wj��኷h��`"Oؔ��b�a���z0ձ���Xc"Ox�1GX��H�AT��4�AH�"OT�8ģK'm�<�0�J+.�F� "O���Sb�':$@Tk�D˛F�MB7"OxM��BJ�t�����!��X�z��"O�-
��|�N���@V:L���g"OzXh�/h%����`�(|���˵"O4t*֡�cۂ��g�М"w���0"O�d
��"�R�ƙnG8,�"O��S��;a�1���3G8��ZA"O����O�T��(�'
�8Y#x1U"O�YRܒ�PX��5? �Ÿ�"Ot�s�J�Eޔ��I�/#���"O� kƍ�$�^�!�o�P�E�b�'��IB~�
n�����,
���g�X��y��'cUe����G�Ķ�y��9Y�ҝ�r�ɴP������.�y���!�Ҹ3�DЅ �8Q�d�1�y"�� ��h0 �/v�t8��/§�y�e�
�����kF�vll�����y芦m�T���/%�n,��@�:�y���ehĂ��Y.8WKA�y��0_F�c� ���$1Ri՟�y"� v�I���nga��nE<�y��6V>�I��";^�DLh�eI��y�)܌_�FE�2��Y�,��M5�y�m�J)J%Z��Q)2�&��*� ��Vd��z��xivj�"CNP�	t��������H�<D|;s�˰h���I��/D� `��׈7�>�J6'��P��(K�-D��3���6B�C�ɂ8h����,D��q�A)\�ؑ�hI;z=����*D��v 0ZR�z*Ǽr��[u�)D��%A�]��]�%�Q?ybf�J#�<A-OX���^�re�l%��X���3��':�!�H8�ܫ!�  �:ڤAE�H�!�$�Tg����Z�ޭ�e!]+,�!�D	�c�~ ��	�$8���?�!�ДY��b&� #�)4o��7�!�Dā~(�أ!kOY�����0�!��Ȁ"
TlC��ը(�(��k�;&�!�d/O�JA�0d]
T��K!ʐB��OJ��j6ʡ!Ɇ�_掼8�ɉq%!��{LqQፘ��x�%��J�!�� �m2�d	*n1����� 9��	7"O2��eKW�+�ř�
@��bŹ"O���qa��L���*���Z��p�"O4 b�IMH�Ȑ�D�m���"O��cč�hS�!c����L�zX��"O���Ф��k}�ia�#��@�Qh�"O��¨P�q��͛ �g�}�a"Of���,F;��x(�)�J�d�"�"O��B�@�;X��`�q�S(����"O����Ja���P�fЪ�!���)�!��&c�]P���
�Μ�HՒ)�!�$Ö/?�4Hg-G�`��ŉ3�<z�O���E*	[��A��*�jɩ�X&S�!�$s�f�d��!���Fk��!�d��W�8DPj�4 �����ꋱex!�dΧ$�2�3�bÒv��ze�ɪR>!���t�q�b��
z�8��f<&���>
�B��������@��y�.�H)<�ʆ
L���b�G�y�ˇB�J �.4��PH�D(�y��Y�xT�j�ag8tæ@/�y��͔{�l�w�7Hό<zV��yhgUb}��+mf��HU)��y��S���p�p��!Xe�J�y��	$��NWmqF�wd��yr��(�!B��Мc��%���S�y��-^�v���k8,��q1gⓏ�y��[�������8�<��&��yb�q�Ȁ�䋅��eb�ك�y2��"hlع6�ק	�
}�\��y�Еjk6��N<����y�H�?���ӍI.x-�"�D��y�"�8:��b2N	#q�
/��?	������(���)��%۷�O�R���f�����L]H�;c�A�h��Ѕȓup���� `�l� ��M�ه�Z��H@0��>���"�H�:Ǫ	�ȓB6�R�`ӱr�߬V��*
�'����5@������CA&=b��(�Il~/��������n�
H�o�7�y��5�>��gbÖ0�1BĘ��yh�"Md���䙴%p�t[��,�y2F]��,�A�*#y�P�����y��C�C:B��Ō�`�i��yj��`K�uB��ԔW5��`���&�y",K	�۱FP�E���"��yRH��H��t+B&&ݮ�����y/�)s��%CZ����ۣ���yba �L���x������R*L+�y1��wo���3��H/�y�d��~���kߟ
�����6�y��ʹLj9�F��4_-�←��yB�R4a�@��H�=V�9�����?9��$8�f��qI�ց6t�� ��#���'V9�f��4s��:���%�H�'�����T*Q/^�L�rM��'���HT�y=J��YN��dgFa�<����O�r�����rI4�z���`�<Q.ӯn�P�1ᇁV�L����Y�<d��(q�/��kZ�{4,�T�<�g̅ ^��t�C�75Ҙ���S�<A��,Ҫ�p �N�}���'e�W�<���M��E�b'��K@E�G�<�a�ٲg���q�9��#��E�<� N��L�_G"	jA�.m����"O�e�Q!K��Y���YM�i��"Oi�6�]e��93g���4<�{���%�S�	@>[�,�*B�&w\K�QR�Ia���b��ުKv�I&h�@
�ꡡ,D��`E^[6��ɏ��5g,D�@ҡ�K2/�h�kG�����3��.D�4��Zx=��+�͘�p�1KTe7D� Y�A�c>��@K���DA��7D���F�7a�����O�,kt\�4²<)�u��,�BO��,@.�ʅ	R�~�,9�?a���~�G#A����kU�~�&���bZj�<�曦#�����9sh���HB�<�5K�#qI�����&%Ι���B�<!$�I,��E	5�E�>��-1A���<ҋ��C0�Ά{��Q�	K~�<��#*2I�PDK9��CQ̊v�<)�AO+N��������afh�W�o�h�?�}Ra�6E­��ƥZupP҇k�<y�Db���6��2 ��D�;�y��8 &�4ؠ.~�&�9+� �y�ω7r�p�ֿ}�|��F���y���w��!�o�'{_�����y�.Xv2@y(c�Ř'��`���y�K��&3zq�gDS7j� �8�y"�Z�XCb�^�
�
@(���y��J&@~�:��T����l�"�y���n���˵-Y	lEh�����?Y�'�!��n]G�f���!�8�H��'�z�B�D]Bȹg��5>�=2�'1^U�ҁV�dz>�n�%���'�^%��,k�j%�fC�s6���'��!㠒+j_e����^����'�1�e�I01Sd��V��QM�!{	�'e I�vIZ���%�'.�At�tZ	�'�d�H+d~���G qWd�!���?�Qn�ػ���;�F4�C@�Ht��ȓ����	��8��mcPk��J�`!�ȓwC�JԂ�tN�Y�u�_ ^��D��R��!"�ڃu�,#���=�>���I��Ӥ���>G��(���;^�5�֯$ܪ�:֮]5J�E{R�OGn�[�l�)���#)�]���
�'�����>g6ؘs 䊸\n@<
�'V�غB��C,����R7T�������3ʄ1��n�2!��̜j^�'�R�|�Z>�'���"�Q��6��BQ���
�'C�4s��S4v.����d��p[	�'L�p��"-�����LF����' �myG�y����GMV#8� Q��'2�xk�Ɵ�R��I闇̕:6%h�'G�X�4|�j�X6K�o�XWL=D�0`��΂F#��Eɚ56��sd=|Oj��#?I�'I�n״QЇf$�P9	�D�t�<�g�e�D�
 �!�%�@�	o�<����.i��|2�BQ�]�:����m�<�W�ϋ[RD1R�M� [�νj'�hy��d�O�#|GC�5[:X���O(F<�*�P�<��V�^�6���ʙ�0���J�a�<Q@�4�p��Dgɮu��]Í�X�<qU-�i����b�%\���W�<yD��,% ����PFj���&�W�<���#,�y����u����aC]�<�DO'm~�)���K4)�Dir	\�<� ~�3��<p#���;g�Y!A"O�P�cMǜ(vD�v	ĎP�'1�	�G�b\��� 2�D�1QC�7XK8B�	w�8:�.��S},��b#Ʃ8 B�I.l�"E;ա�%ig �#я	���C�	�N�f�.���8���_���`�;D��禇�J�4��sj�1 @l��F&��~����[�4�I��ڙ�Ĉr!���B�I�c�81�+!�i#l�^I�C�>�DH�3@�5\���Ir!��| �C���Ur�^")��ש�&e�C�I�@x��F'R�>5�����pg~C�ia�k�a9��
7�Lx �)D���ˑ#c�x�D�T�E`s�1��0|��W�l��|�T��+v:���Fߟ���Ic���ƥ�:�RI(vB�.Vc�]�ȓ9Zm`S]j$hUQ�EDY/`Ї�bu ���](���w\�H*�ȓB~A�P�n�,�Q`K�t
ڨ��,i��8���t,(ҧJ��ȓ��Âg��H'��%F�5�Ƶ�ȓ��`s�6��P�^[����'(a~� G/e�D��>�$��g���y��۳&-tx2%�Q:gН��+���y�=WX~	���>pV0�q��;�y�	:��٨Wa�7�α�F��;�y�5V]��"FJ��<��u��CՃ�y҉$Y���@g��%��!�!�E�yB�ƞcb.8x���	���RT�B!�yBC)o�d0VA���|x%�1�y�H�6g�M�揊��ИB���y2�ު)�Hq+"C0K3��`�9�y��K�N�
Q��쟯u�`c��y�KF��2eW�x��õn�,�y�K�#��爉�P�e��j�<�y�(�'v��e뀕hr�ԤÌ�y�X�J�/ڄ.����Gֹ�y�B93T��Õ��"#S��1��yb�@�� �l#���AHʪ�y�w�%���5n�|B4���y��Ä� ��,�^��C�� ��>	�O�x�'�I�3��:!�w:fث$"O�h*���rhر�N"X*5�a"O�L(���XH��0���<Qp�v"O� �����O�@m��M��?��"O$�*�N33��J��K���P*�"OJMr�J�:��TKV�S���K�"Oڹ�g�!vF`��'KKn�
���"O�IY�e[�I�� ?=�y����#LO��Q�!�;� ���JU��Rukv"Ot��V�X�g�2�3F)�&K)ʌZ�"O�	k6�+e��`���/h�d "O�L8�EC)B��6hBY��i0"O�H�䋯E�>��M�9�4b"O�������1h@CT
~�0ܪ��'���+v�D�p�NC�C�$zG'1���=qç�hA1!Ɠ9����JһS6���0�$�"��<����-ž��ȓ&�h,(���j���)un�3_AT��ȓp2��#΁�uoѱ�)ϗV����ȓ�ؙ�׮�,�Z��b�i��0�ȓp7�$+�&�.A�`���ϋ�q�<��i��թƮN?}&dP`��!vE���i�>��g���b���M�}ܞ}��S�? ��H�EP�DXR9��j�6	�z,��"O�MK�l_�m�T͸�o�+ ؖ!�p"O�M�Մ[�v� �����':�Q�"O��fZt��(�c�69��)iF"O½qdO���hL��V�P�"O��HQk
6$OЉ��7�� @�V�<���9q4Pi/�0O1�xx��;H;
B�I0v)��U~���ԠW=oB�I�D�����Ԙ^=J�k��-Ig�C�Iee*�9Dl�0f���K�j�.B�I|���fC7J�&D�ǺM7LC�	�G+<�g�V�^M��*�أe�pB�	^�
�c�ų�d�i�l�$+SbB�9o5J��j�~l���ȫfNLB�	,�h�ңL��_F��8��A&B�I��h�i�ͅ'?�ʅQpEƺ[�C�	�uL�`������ܢw�� z��C�<���㘻���E�@ �C�8'�Nmi �����/�:v>�C�	�E��H�C?���@�Ć@����$&Kf&q�؉K��h��	tp>���b����Ȓ�
8�0ꃈ9k�ͅ��J����U�&&�HaV'��8��(��U��,��Z(վ��%�
��@��?l��x��ԘOmzܨ�wĄ�ȓ���ԀG9{zDa�G���@%&8�ȓ���3D�\7�m�t��5㞀��\��HO�D���A4��?7��ȓ/;HD�BD�<{N<eq��L^��ȓzӴes�F�a��*5��E�Q�ȓ`0�!GƄ9x=�R ĩxl��ȓE��(���65������4��a��z�6E�&��ni�����a�hY�ȓ-j�hs2���S���(p��$�	U���4-ϩ~_2%i�H�d"�mz�e#D�H�#CA�D��	pR��`��-0�j$D��a�(Zp�0��^�^��p�d!D�x���b< ���b\<؊�x��4D�8��B[	z�j�r�.��9�^�T(D������.P�:��L��D�j�o$D��*���2�Dh@�a�6�ضA-D����2�� 
A.&U
�!�&D�Њ��ͼMb$�$��4�b�/D��Y�J+Ruԁ1�Z-uz@���.D��g/цz+���� ��űr�.D�@���o,҉	�
I&$�81.D����R�9b��$��H@�9�O�I�8 .$K��ݺ4<H����2ش��0?I�*Ӆ1��WnًX��-���]u�<�D#�%9�
�z%��Ƥ*���p�<y�f��5& y��#K���1&�w�<���~���#PM<R8И�U �v�<�l�Y�¥	�#L�l�(Uq �v�<q2D�7I�Ls���m|֐)�J�X�<�V�T�sU���C��ig.0��ML�<�Ӂ <��ѣ*U)60�)�Q+WD�<�3.C�F���0!���j�Z� �hNY�<qGKF�AxH�d�2@�|-���U�<�FmR�j8���&(:eQ�u�4 P�<Q��A<�xB�Ց�D�5D�K�<�WC�<7lp�ը�*g�)��a�R������i���2Z>xق��:��	�<��'�`�f��&[�`]T����b�<�O��1�����M�fѺ�h�/�G�<� tJ��Orah !��Ή"(*�"�"O��r ��-3^t����&y�&D1�"O$�QlP�R蝓)G$0p�̂�"O��٦*�l���f�C�7^ܸiW"O*0
ǭE�r�,�b�?[􎐊!"O�l�5��?a<BYg�t�4L �P� ��ɐEF�ᲄ�?�ؘ�G"��!=.C�I�,,����*s��E��J��H�JC�ɸ8L&���&�k�R怚;S�C�=pl �#b݅�ڰ����I��C䉇/�1js�M�M���bܕg�C�I�N� 8�����a�ԡp�Z��C�ɑE ݙ��ԉ)�X��K,@pC�I;
f<�J�_�90�)dF�iW4C䉎Wҙ6%��O�5xP@L '�C��:��!���2? �B���;CJ�C��,e��(�����P���V��C��9&�Vs�E�/���2�BC���C�Ix6������10ԝ�T'_#;lH��F{J?19V �C$$̠ �Z-���!2D�t�K�(%P�L(�iD�v+�xA��=T�$�`�Z���j��\�$��R"O��K%N��`�(�ʅ�����"O�pU�ʠ ���aC�vrz�J�"O6�:$�|Ϯ�s`F�h��G"O2Xq�Ä�ZE� ��C �R��'iў"~�Q�� �P]KS����Q d�$�y��?26$��E)d:�(��"��y�M�:��U�G�]��X��)�y`|#��DOZV]�&
6�y"��.R��K�F P� 8�v���y���B8X�M 01=����Y�yR`FX3�qel -��k5��!�yb��B;�����|-�ء�Gʢ�y� ��C�LB�@�q������y��v�Y��.Q7uX�0�����y�E?�B�K�g�
�d��-���yr	�\m�����,+=�
Q�A�y9p^�)`!˾N�Ɲ��ƀ#�y��S�C�8kƥ&J66 ��g���x��C���X���F��ݸ���6�!��8Ux ��)�u72m��8i{ў��'�>��$�U2"b4H�'D�
� 1�F�.D�P'@��)�����,�C� D��zg�7|���4��R���R�9D�iwA� #+lDS���)4�H�g);D���R(ZE��`G)���ր9D� �C�*2�r003�
�KƱY&�$D��C"b� @�3E��B�1:�h$D�$r�N��Q3R�#N �OkZ	Ȑ`5D��Z�BH�p�p%-_2[�8-�e�3D�,�GK��n^I��AJ6P�8�;�D/D��:T�Y{����C���#%K.D�k�h]w�f����7C������O��=E����	WC�݀gG��ĠВ�]�[M!�䊁<"���T%��ސ��\5&�!򤃅TR���͸\$e8FK\�!�ě�{j6��'N�;����� ;P�!�$V�@؎���!�4':l�֥��!�!� |_l���'�QV�A��7�!��ͧ7 �)�"ζ_8([v��/,�!�䋟s��\���D9E0�	� ����!��|̸���F< A[�ʕ�|!��&�U���K)%�Pñ�P�|!�� �D	ĮV:�����B��)kv�q"O��Yi�(p�`=WÃ�Q�6"O�5P�n
�1���h	/YB�=:�"O�1��l�m3��+�ǉ_/.�e�	}�O!uI�㝖3�����"����'���蠬�4cxލ1�i�� �� ��'������΄�0�iaW�k�t�'�j�񐄒(;�۠��	�Np
�'�N�:��LJ�^�3f ��`�	
�'�HhWρ�
$�0', (�\,���d�O.�O��S�f�"�Ss�� 	a�IC�P��Ox�O��=��!7*��&b�7 �\0����:�y�@7MԆeq��&:p#4!��yb�܎,�噶�֖NO��# ��y⨉>q����E	R���K��/�y����	�@�!��ϥL����qC��yB��#}W�Z6&�L�.�ADm��y2!����餎Ⱥ9�X���J��䓲0>�Ǔ���NΝ_�<SՋNZ�<A��7��m����bT.͊�gGY��d�<!���
w�L9�\!��"��U�/̬B�	�d�2Q�|MV�xW�׀V�vB䉛7sP�:���*ȲW▧#�:B�	 &��E1�"�t�������>���)N�����A,W�ࢧLҦ!Y6���9�b`�-@$M��H!dH�Z:Їȓ	Иȷ��lv@|`����e�ʙ��`�'b��",�0|�8@���VB���'*p��Gi�W^|̀�/�H���'\DB���M�+aG�%��b*;D����kƗu#�1��Ҩ]�*墒,:����T��"��%�%r
2rz�7i�<����S�
$�P��N\�k�Ƅ�Ɓ�Sg�B�ɴq$�Ӕ��F��p2����<�*B�	;N��i��٣Nvz,���ڔP3 B�I\�H(�F��D��7��+6��C�	�=�\�&	YiDu[��XѲC�2m|�m�X��҂F�XGf����<D�����#�v�C��ɱ(��e,:D�I�l��WX��(ȡEml��
3D�,���t��U��:o�����<a����6�
��^�	'^�#'��0anFC�I#r���9$���Q�	5�C�	�%��XP�ɹs9j���A7�C��*Pl �$��Be�x�⛨dH,B�	+[`��k�6}��I���*=�h�$7ړ��Oz�E�ɖQe���.J��Uu"O�8���Љ ڀ���O b�Ԁ��"Ot� �XL����@ ��P "O 4�Q#�v(qAB@ �K����#"OXm���hbPۇ�)^����"O$��E�Ϳ>~44���!4��D�C"O��r4L�2B\d��؂msPe��"O�R��u������� �mj�"O���snĕ2l��eL� ��0Ւ|B�	d̓cHd�0�̚ ���C�K>
�fI��:���ę� j���k��<�ȓ�lt��G�/B�=�D�����s�2LS�)8,��E��"�r�<|���|�H�� !�n��f 0L� �ȓHĶl �'#��ܰ��$`u�9�ȓ~�H���
	㶭���w��̇ȓ�,�`RƑ��P��.C/%a��?�ӓ�.m����=w���� �;r!�u��S�? ����\GE�V�U�ʤ[C"O��N�`�R�8�j�\݌�
b"O�42�i�&^�BБ�� q�؉����O��d?�'p�z��V�'rlJu���HFp���IX~��C�Q��$����8�:������9�S�O�Mٲ��MJ4x�!�ڪN�Ĝ�
�'9�L���X*i�`�XQ��<b����'2j��霝T�x)���-�6���'!����_-6�x�	��"9� �@�'�0���T�A~z��o
�7_�e��r�)�$A0r���P��-4��r!���y�ɀ�_�P�9�
** Q3�]:��D4���'��#�(�)���	�#�ThR̃3"O��	���2�MY�"�\O�M��"O�{ӏ��T,��Q᜵k9���"O��c��	h]J�#�/Є7�qbV"O���#κI�2Ċ��ж,��������O�d+�( ���d^�vN!ɵ.�d��фȓ�:L(F�$;��9�BYYфȓx�m��>%���h��V�?\�ɄȓkF��a�~��΂N3��$BK�<)5Ȍ:G�`���'bR)⡁I�<!�;*Ͳ�[��P �tM���P�<)s䝼rH�9�e_�!� ��O
M�<IV�׽��-�� 6�|��l�H�<��ʘa:$�U�*�ɒn�E�<q�IRfp�d"b�T�v�D� ���wyB�'R�p�#�
T6��	��(��k�'G�@XЧ�%X�ar�Q�h���1�'vNH�E
�k�ll���˳b<M	�'@��en
6Y.\H V%1��"�'��35MFGrnܪ�a��x�D��'������҇m�^	�d��H�|�����̆)�~�*`�ňH{�;S�*�!�d�>|ıy�΋�)�� ��n�!��cP�M�W/�H��2!��BEF50�ǎM��8a�ƍ9�!��hn��y#�͙
��i��2�!�>�֬�#�F,D�z��FV,{�!�D��jPT��g��w��i#�*�!���Wݤ�xaԝT�4��ĬУS�!�ĉ�,ms)��,(��j��R�!���Q+v�}F�i�)"�!��>}�1!',�eI��e�!�d<m�̄��瞿^@�JJ!���ޤSc�[����j�>oN�O��$��6�ֱ �._�^L*�3��c?!���	^:2$ȲQ	h^�3�����Iiy2�'�����O6�0=��!�<���'�8U�""ގ���A�_y��yr�'���b�+I(�8���
(N b�'�t�*�S&��뇬ֻ�p��
�'1v�s�kĆH��,�G��U��{
��y(��O��c���[�}�-B��y,[�fE�Ls�e���ŉ�C���y�˖&nF�<����D�X�B� �yr �4"O���^{5��S
�y���]��9�+D.|���ѥǬ�y�#�c	�Qy�* �eA��K�H��y��ў$���I#n\\$4����8�y�˟7 ;����*[�N��������yb�	<g�@��L�������y�i�ϜD+�fC$JOR��S@���yB��Aؒ53bFXU�,鸧���y
� ړ���x)s)W	�vs�"O@q�.̨d�X�኎]�`��&"O��q�D2l��d H�x�|p�u�g>}��@	�&�i�&�̋-�����<9�q0�
��e����%�W�~>H@��;�e�2C�e��X�2��8d�Ć�Z,LѷjZ#w�����/����q<���b@f� ���̯�p`�ȓ���y�K�P�i�$B�/~i�E�ȓi�4��f�]�N��6�D�&�هȓW�`r��C!B�X�'�W�`�VT�'�ў�|�
B�מl�`��"Tn!Z��U�<qp-�:/��1P�_�F�6�yb%L�<�ǔ���eh4���#��w͞F�<G��}�B��3d.a�
���E�I�<��K�T�J�s�ʀ2{a<�4�A�<9� �:Y���۠�@/d�mj�'�{�<��+Ə|��\@�+M��4pS�w���0=	�ѡq�b��P�1�P�3��q�<�f��&1��t����G��Pk�o�k�<�b%�~��)�(�\hiG�B�<i%ԥN^�Es�Ɯb�x{�CT~�<�qK��H{��h�����,3B`�<ٳ)�8�4��d�HͲ�:R@N[���hO�|Ǵ-*��^�D�3�(<E�u%�8E{��T�)fnؘ��)�������ρ��y"%ܫ覨�D*�,&�!
r��5�y҇S��0�D��S?�H���=�y� �1!8M�q�L,]nY��W��y2n;j  �z���_��x��jN9�y��R�cǲI�bܻV.������hO@��	C&"u��1���(��� ����O�!򤎚�t���Z�N|�%{Ѯ�o�!�߿jh��cd)V�9�hP�n�!P�!��B�#7\�a'	��Mlq�b�$�!�"1��D�QR
m9�aA�!�$D��9���O.@dS Qw!���8�x�*_1��$��i!���%�|� WB�v!�U�__!�D(Ml�F�'�<�`/KpE!�� �Q���B�L�-ez�R���/1!��Ϲ\��Xw/�96~���f�#g!!��9a�"US3���p�J0Y�!�DB����Ս�:)���悔�M!�� �jp��D��,��ሙt�!��2U�J`�g����JL���C4�!��?	F�qb둌/�����M��C�!�ċ�����l]�j���"� F�!��h
9rѮV.�����N܎a�!�P-D�90��\�q���Em��7�!򄕊
-ؕ"�gJ�{��p�b�V<�!�$�d�@��A��Q��ө�!�$�	A�hD�0�-P}�%�c��n!򤄵'?�}âh5����Ǝ�w�!�d��|΀�A�F�E����� �`!�$C=Xl���2���s��Ҫ]�!�$�@2`��	R&��lb,��|�!�d[?)]�3�\�_�h���Ӂ1�!��1u��:cۺ-ʃ`0N̕��/.�Q� �G<z>�:�(�)���*V4�QiL+C���3�G�tH��ȓh�D)y�� $�k��[�R�D�ȓǌ�s0䓢�����aX�Qq:B�	�l����R�
�WF-y�§TW�C�)� ~�(��� �N���փk�^��#"O��3S!+����o�;Y2��"O $�H�}`�<	� M� �$(""O@�B�@�A/�Q�#o�d (b "OXX�Р���� "��/��b"O\� �Ȝc��I�Ai#��th�"O�H��H��kTftYD猾�N	��"O�y��)�)Y�N5B�
�[�� v"O\$S���+<�jP��%�2c�x�#"O �Q��C�g0�|c���@��̰�"O���VM4?fLӒd�3p�JY�%"OTt����2n�����BL�1#"OaX�c�!M��IR�6lc0�H!"O��8�������͋ZLFԚ"O>�y�ˁ�=� �/�QKH`s�"O�}sVj��Hc��XS-b:Դ��"OR賵͈c��)s��	�PA"O������h䀥���g����"Ol��.���D)Bȓ1�<3�"Orx��*T1�L���� 5��`�V"OQ��N۫;@�"s��;�
%�D"O�I�w��+td�	�@M�	�l�d"O`	�(���u��	�!�X�d"Ot�cU$�� 2՘q�ֺxk<�Q"O΍H3�_�<��Ǝ�*P��u"O���w�7T�k'T.m�`<z�"O.�k� �+D\Ҩ���2J��<0"O,#ä� ]�L"�&��3p�a�D"O���3
H�\��e�?��I�"O<�d ݔv.���B�%)
�e-�!�D]�6C���f�F(�c�"E�!�DP4B}"�Z��"(���&r�!�ڵ?�t��aĠ+\2��^ ?�!��T)
ұ���25F�C��l!��<�X�b���'VA�magjԔ|+!��D�x� �04�d�T��H!�/T[�e�"�I�{��k�Ƌ�!�䙮'�5c�L.1j�!!)T�Z!�D�1at� �S��� �'߃)<!�Yo��c�УN��	P��A�U6!�Dӻ>����C�],�$s��Ѽ{!���&.Ff���Ћ"��{�E)>�!�$�x���"	��a�M#�!�$33�K ��%9�b��b���ux!�d�S��@�_9 ��Y� '�':�!�D��F�,(�ćڳ.��p1G�4I�!�$>-�,��wkH�D~��gg#!�d��������0���Q'�N7!�d�Y�6UY�/��(�(����m!�N� ��3��lPS�e�4�!��ʩRC(��i�)kj�h��?Z�!�u���w&R� Sz%��\��!�ȗ-b��J"��%#B�	2�ޘ:�!�$ �d\ճf!�n-<�r"��-B !�V0i�Z�Q�E$r�RDtF9y!�ڤ8�q{P뚾c��ڠ"]�.!�dؔHb�L�! [�$�Y�Ӧ4�!�XW	�4�M�"� �#��hK!򄒲]��tu�)v�veң��4.!򤒥n��`�W�Mh���a8!��4����r��6��4���&-!�d�#h��s�M�� 8F�7J�!���oĺ�`�*͝J�Ѐ��e��0�!�P�&�Rɝ�F��LJ�dʹg�!�� A���_'N���pQ��/Dh�{�"O���,�?}2�sTL�W?ƹ�g"O�*R�ɓ-�2Ѳk�1
��"O6�h#nO�@��A�Jʹ-=��U"O|� 0�I(:*�������v"O��KP)�L����hC|r!��"O�TWޠ��pnL6\�Е�'"Oxx��L�}BR�ʕM�mel�1"O�([5�S�-�H@G�˛3��Q��"OE��bJ�c�(d1�]�^؝"O"�v��Vf�� *<[2��'"O��P��)�x�x�(�b��"O��� �:%e��Ɯ�N�`��"OB�d�*������?Mo����"O��bghחI�Ҽ�T��'jV�{t"O*�1�L_�U� �,,(���e"O\���oU��1�%��A��m��"O�x�.S�e}���m�3$|F�y�"O��Q�H�\;�`s�b��z?�j�"O�uC��տ|��y���216^�q"O���a��vt��+�˭`/@�"OT����8}��u�����B"O2��T��11�ᓱFǡZ�����"ORQc�eM����eǼVE�w"O�%� �ѡ[A"`ٷ�C�?��p�"O��`��֛�Jк0�	�W��uH�"O�B� Ѡ
cdK��A
N�"���"O�@ir+$��eE[ Itt!��"Od)���I$`�� ��YuZN���"O�ɨ1��-�������j�0"O����i	0 
� ��ǭgՒ��"O$\r�c==�q���^�:p�"Op��!Y�(V,���=T�x`PB"O|�CdP~	Bq:P�ڳB�h}�"On�X�Z�U;Z�O�S|�L3T"O�<��>�2��w�0J{~i�%"O�A���6,��OAi��%"Ob0�(l�|�򌐾/��l�s"O:E۲B�Lf�٦L��L�ĘSt"O�E`��'LBys֪I���"OR��$�T!K��P"�X�I|\�(B"O�|br��&�Ub�W�_�H��"O����K�v�h,��
�>N�k�"O6q�Ȏ'�0�{i��L�\I�"O�!!��p;�����j�����"O8y8��� ��P��K�O l\y�"OF9��͆._L��F�ݳj+8|�"O�����6~�D�3r�Ձ�D��"OJw���{?ha�QNߜ�� Jb"O�h���~��]c4�G����"O���k߆%���qn��z�d��"O�]y#�ӥ"T��:r�Y�M�}� "O����Pfh��WD�3n΁�A"Oj�t�B�E��z�K�;S�x�a"OZz1�
�a!���d���zd��V"O��Cq�f\�hҢ��N#��ѳ"O� �W��9inJmz1�E�,xau"O��� )[?8����,f�Q�"O�����5|t(J1�XA��)��"O��hP���
E��� /^ hɴ�� "O�� ��_)}VH��@炅:�Tpr"O��"��8�� �2L̸k�X�pW"O��qAF�z�hH��kB� �r��b"OF��BeėOa����~hz}Aw"O� �ɰ ��s3n H���!4|uxa"O��Q���+�2H��#�`+�C��!lO&p#@H>�@�����
��5"OR	
��_;|Y�`�
K�bȫ"OZ�	�e�7|˼�8� 2�<��"O��Sf�#B�D-Y�c�$g��l{b"O^A�� ��N��v���"O:!��͓]©
�i�H�:�kr"O�u0w$	����H&	Ǝ}���#"OJ���0 
�ڇ.�rزܸS
Oj6�]��Ph*�̉Č�5!�Ė�WPN�)Eo
���'��:�����k�KϢ,z���Ov�U�`��"�d�ȓQ��܉#F餈���7q߈��'H��(�)ʧ_iv���E�]u,��ٴ �\p��C ��83ʇP�$I@��-O�*�Gy��' dU��tر��Q
O`���'pBy&�.#U�U��/�fn��7O��A��q����x#�� #"O�䳧nC"x�H1�a��.H����P"O� u @�N��T�ghH':�h)0 "O��P�K%����E	F�Zp��"OZ�K$ �:v�ֹ�3�܀|��I�u"O�u���ه/*񰍄?�J��"O��c�HG�OX�E�$-�,Ey�u�P"O�t���K���8��дbK}
�"O��!cF[�w�N ��P�e+���"O�㢃�)Y��P�dO	2t��"O������~
�UB&)�XV��"O���2X(���W�aR(����"4�t���F�bW�1�'$ؾzD��I�"D���Ӂ	6l�`�H�o�H��ؘ !D��zAQ�g�l�rt�>e�li��f>D�|1Wg�j�5Z���T��IxR<D�  NN���X!��ޑj+�-qs�%?!	�]�>��w	�	 �u��&Қ`x���>�˓�M��Ō 1}�� ����e���ƌR?i���l��Y�A����O'knB�c�"O U`B	$G^��"��vV���3"Oy��L�Fޒm�K�����#R��G{��鏠p1�m� �ճ]��B'Y���I�<	�}���ʋ%{
hF�*]�`���Q�H��I�eGx����w����$ޙ+d����*�0���>Oz���5P��h����Y�"OP����
�0K��9��1JĿiʡ�$�L:�S�˒|��q  ����y"D�+
����a�
s
�
��'���'�1Oq� �Z��!�P�#�
����CW�D�O&ʓ1�>i��J-3J
 �jS�<
�`��B[��yȆ�g �i�KV�&d�%3P��
q�������%��O4� Ť =���7Ċ� � ���"O�)��E�K���xfM�C޾��D_��oZ�g1Q���>�+��W:ʭ�`'Ǎ2?�1#rNoX�4�O����(0��@ԋ`�V� ���a�A2�MB%��'�ɪv�؅�d֬�,d�$�ѫ0�C�I>�za�tAصB������<�7m5��:\O���S˪���B@<.x�h.��'�ў����W���Mj�ũSA�>Ĕ���"O�t�_3}(�I��!r���iPT�ĕ'�2�(�3��a"��Dn\��H��h\!!�0��k�矶\��s���:Se�'��O=LOT�c6G��4Kv�-z�\@�O<y�ÏY��n� H�$�$`��n�K�<��UZ)"�D� DV�*��B�'S���"�g�? ��8���No��35I\*,�9��"O�l�a�Ķ�<��ڬ!��Y�@�|�0�S�'+(>�:�,��\ФP+�i�;�nh�ȓ$�.)��ꈵAܔ�G�N�>��=�>�ד'�r͐�f�$�{����y4"��ȓ}��M�S�ڀ�xY+SI'C�t0�'F0��/�9��P.�H:����{�)��J��PTJuÓ,?��=�W�L2	�!�$GU����n��.���(���!��R(��������E�r�3�̋�!�Z�c�ZXuK�3qtЈ(�#���Dx��'��H{�.� ohL��l�)��+�'����V��/?�����Q���
�'O�=�5��0��8s��T�c=*	�
�'�xxIC�D
]��5Y�i��P	"
�'#:� #냠H�T��8s���'M> ����?\����	�p P�"Ú0|�����*�d�+C�܁���zG�����ݍ<�!��z u‭[�;=>�Qs]�!�!��o�8!����`�P(�&�;B�!�[V���f�F�|!҂@г:y!��J�E�Kc�#ⴣ0oT�pg!���,[�=ٴDҁ. ��Ѭ}:�'V�6�'vL�!j�`�~(XPr�4��	�'ۛV@�R�����wlp%HV�)�yR�My��8���C#w]�H��/��x�lӱYd$���37�@��	.k!�*DZ9��
�Ɛ��w������m��(�:�r��E3^� Q6&�K�*aI�"O�ʂ�
�j4(�"���-JU"O⤳�� �g��BG�x�; "OB�"#��{�9�U���`���aD"O�آtK��9�f� ��6	4��م"Of%�.��=����"�V ~�ބsb"O��u)�1P%j�
��B=@~��$"O��X�c��'����4C˺4D��H74��ZPF��Cc�r�AD�bۖY�D+�$�S�',]��� ޚ#�y��ش@��0�ȓ{���w.عp'�8�5�J�gB�5&�,�'��x���-�d���*|\xX��F���?�'�����#]�$�y�v�_,/=쀛�'�n�/V�X�����Iݿ8��ᨍ�$7��]�I��"k�(��kH�^��9��e�?(�!�_����ⴍ�2z�b���E�I��'���z���)�'9Ԁq��
#��'B-�!�Yn��I�$d��PհĀL��	_y�)�mM��h8#P�LFXY�L,��O^@���OΈ
�'�w%�=F��J
0����;O���㍣a�� /P�wu�Pbp�'�'[J9�*�?&=�V&L�+��19���xR)�E.&��զ�(sz���r�����y��)�Tȹ�eIF���b�������<�Zu8�Hۡ�2�l}� ��&�!�Dү*��́�o��t�`Љ	�S[a~R\���i�3 ��ɓ�	�#b��Q�c�)��p<�� Na.1���.W���pqJP�'7�?+��M�c�쁢(<L�*D�<b6&��JH@�Ҟ�]��C����t���iω9"��$���L� J��D(Y!��q���:5�.:[.�)F�y0��$�������b#�����i�!	�F���l��
�Y���ZNڤ@�!\�E�ȓl����#��|���ٶ���'���G|"�ӑ
E��T &�����%�9H" B�)� ���6=,=������4>O��=E��D�$�v쳶�4l<� K���y")S:Ԡ
A��
a7F��e;�y�@�.M ���GH�g�B	ӥ�yr��8��:g��Y�n����\�yӓs'd�r�e��OK�!!�*�y"�A?ct�`��B(�|7$�*�y�_��� ��I�����y�#��Ēd��I8��$��y�H�	a����^�j�:����y�@�Y���3	ͮ�TI��:�y��Ky���L. YCd��y�iߨp�yJŭ�0�d��'j�7�y��C.�ʶd7����N�-�ybo *��)���>:h�ʡʛ��yrgƄ*��|˵��L���� 
K�y��x������<4P�d�pf��y2��c!�`��!�8wR����y�.��q3�/:����bȽ�y�GU�K���T+\�*���2"��yR�ȶj��x�`Ӧ /:9���)�y��m�� ѓBU�Ј-���1�y2$��S�B��Lq4lK��y"��;�~�����&�����-Z��y�&�=�lb1��?`]��̆�y҉��@n0z���5�YBP(ú�yR�
,MN|XRdd
9 ʮ�s���y��1X���j�)��"����t�D��y"C�,�L [&W6�X��W	8�y�3�D|{�J���=�r���y��B(�$��f+V�1�X!D���Py��R>����1*\]�'.�J�<�H9�jLr�6�d�֤�F�<�#Z1��ˣmG�QڤH���|�<�u���O̠�2�8�6� �y�<A�b�0��){�ѳuv���b�t�<	U@\-. D�D�/�"B��<�⃧MK@Ūq أ%��eq���n�'������P�@,�Վ�8V4�:�'~��T�� $(sE�K�>�` 
�'��dk�o�����#��A�6쩂	�'�����eڼH�$�D(/=8�[�'�r�q��?TX4	������9�'�FQ�6��:Yx�L�d�S��PX�'kf�2��Ǡ?{~L9t,���<��'o�a�Lu
D��P�S�f-8E��'�x�l�ec������S��}a�',0���%A�bfɘ���+��'��\ 1����BI�@-ӤQ�!��	x+�iKr��&�P�0k@:�!�䞭C�L���H��;S
Q�~�!�$)�XP�d
U��Q[��Z�#�!���&�LC&GǓU�(��Y�|�!�d��XZ&�c��3T������$W�!�D��%�̤�rK��{)h���e�!�d�:5N���� �07��9�2K\8J!�䘰	�	�i
#Zj����X>!�$<Q��liBcS�r&�-�b�	�5!��*-Q�����UJ9�R��!�S�K�"�yрM*Je<=뵧�c�!�d��ZZ�=���֬s@NA�����!�
)���!� 1o� `�C+�!�$]���8X�k��T,� A^�!�L��FPI'j��)�0�"�4'D!�͢�&�
�`X�0��@r毚q?!�� ���fҷ*���6d\H�:�"O,�˒��B���E�\�"'���"O��#�3I.��[�c��J�a�v�<���ˊV'45�0�!eȵk@K�n�<�P�C=}��hK�OA�,W�o�<� ��|�±��@B�j�*��C�<�T ��Υ`5牻!U�r�GH<�=���
����Y��\��9���+�O�PC�l	�)Gɓ2��!!R�����'��It�ʩO��'X�H��J<K�R�)Ԏ6%�r Y�'�^�����E���:ԯV&��(��OH�,OBqYH�"|��J��L%apK�d P��O]�<�C�
�n
n��g�S�1�"@Rw�C?��'a]�����Ϙ'����H8�\i�jE"�x�8�'��X���4��m���=���r�A΂u��`��\v���z0��g�D0�Al)6}�U�'O�,��dyf\iH��3�nŴ\8(��ƬΗg�=R�!D�D8 -KE��E���*7�4WC5?���H|Yv�Qr�&}���Q�t�ĥ�=&����2Qb!�]�s�(����V$2Gb}�5oX�M1�*O��҄+�3�vb>c� �Mϖx�4y��EÉK���"�!�(1���9��������C� ����QhH��
H;��~���6d�q�Mz���h#h^*�0<���ӌ^g��[o&}"��00\�v�N�i�^����y��1I�V]rK���5�䪁���'>aS�iՃ��)§B���􎓚f�F84�q�H0��8rUx��<�8es��1����3�|©��3����}&��S�G#j,9`�.�<���
p")$���1��KK�	�p�Q�H@��I@�!�@���'T��3uf� %�����n�`�Ă�'Ɣ�� .��BdK�3hm����'�ba)A�I�Ya��	3gߧ7+�m�	�'j2��ؒ?�u�-��(�l��	�'l����3�b�
w'�&ebA��'N��X�B�#%kZx!W/3$_XL������Z q����6i��|{H�3��Y�ݚ`c!��ƀU�<�D$6`����G�G,¨��NAp��|���Q��`K&�ː:��1�!�,��C䉳%p��KXr�v�{�� �:�_� ���c]�&v:��$Q���l��|#�(j��D"Ta}�䑈@4�,c@�A�Oi��x�3�ൣ�bC-ѥ�(4�x��� ���yD�Q�C����W/$ғ{$2́��Q<��6�щB������v$�a͟�ΠPH�N%O�u�"O�쩄E���A��'���ys�i�ڼ8W!7-y�� �ճ<j$X�C�s��Iѧ�fd���,��#D�Lh�._�}xH�KQ���|P	!LAE��������Сk���'=!�$zVA�/���H��DDmN�:\h���Q��u)TLZ�2 �!!�n7�0Z�lb<��嬃��`��c�,��)G�|ܽzq"0[vT���~�v���]�e�(�EgӘ�cp/R�69��o��?��\��!۲�ywJ@�&��=��g	�:�Ҥ1tHU�y��_�Gsv<J�#Ȥ ��1#%�l���[D'F 4�D0��2] �&-�Frr,b��%��s���ywHg�> ���R8"�)��MU'�{b`�A��(aP}�(|�@�[����)�x怱� !
��}x�κ��i�G.�&`�����[�DW|S|��cI$ֆ��+"�I�Z�nmb�=��@S�J:�	�EJv/��*���D���-��l�2P����#�W'�l��VF?�O4��"�*mF��"N�5L�&��q+�Đ���2/�h����:�6������uw��9�>��Ď��[th_#IW����|_�@��j�_�<�6��8*l4�¢�!yR��F/̙jq���B�G�. >-���"k�ܔ��;��"i�ր�]� ��-�@���j��ABНRe ��ə#�I�Fэ����#�i�"@�Q���5. kp@5� ��59��l��d9���b�2.�,{�&�::U�O��b��K>)z���S5`P0IN|
�/�)0N�FX�n�t���o�S�<��ŀ05���8F Ί+����*��?[ kc�`찀R-L�[�lG��'f<����]�z�C`���d��,k	��� ���!���%�A'v��|��!�O2�	@�٬]�`J�
�l�?i�k?"Kvع���:f4����/�f�4�!F=�>-��a�j��-� �è�+��-ԡ��H;���t a�M��{vD��=�ɝQB��P�O�g ��eF���OM6�Ѡ_"HO����I��H���	�'�����O.Y�
�Kc	�0�h�XV@�L���(��2\��ӭ�(�剎w$��A�\F��פ� 2�(C��9K$�0vLT<��(���Xl��t�A�a�H�{q�	�H���xх�y�'�Z��@ǎy}�E�P�Qd����	�>�$A �H�A��� �G6&�(+0m({��U�X)'2��2�ͳ�a"�P:c������
S����䏝Ҙ�5AN<~X!{4�ٲ:���T2��'I��<`�@ٜ<T����m�)��%��O���SӅX�:��$�EPd�����O��0V�����H�wVy���{�'"���H��v���OB�Y`¬Z81�Ɠtc����ՌC
xJ�l�'�zE�U恻_%L���$�$�DQ��(֖[`"?9`�K+>���{eL }W���VBx��c%��y]��� Wl���q���d�+� �']@�@��E�H�`�'���aO�oM�@*����h�:H>!�A���|�Z �I<�` �v��1(�V%�v��x�*�b5
˔51�"Oz�s2O�+�D��H��N�U�åF�"�N�:�/E�����$9[��5��O2Q �6-��JcHèM��x�O޵Z��%t�PYa���	
�~�*!/ث�|y
�l� ���/,���F���F t���̷���YF����<��������-�^��Ĭ��>$v�"�kE�#b�bJ�&< ����*�:���N�~�z}&��%�,�<	+E�&���L�x%���7�S�H�F<��F'0�X�yF�M�0D�B�I"	~*�Dˁ�+@t�A�V�2	0����E��R�u_h�8��!�g~2/)��p���]qN�8���:�y��D�'xF���i_d6Ԁ��lI�V�L�[�ǔ8;���q�Iʔ��dX�Г��Fi��lA�"N4;7�z��$4_��Cm�cmJ���?k�~DЍ����w$U�;|�'��Wdm����$_�~�[�q,�XGi4�IG:�]:U�L&	�zy�ş�&L�	l(Z��ȸ�� vb�& � 9��`������KJ����
�m�T)�P-N�MΤY�Ą*>�$Ӧ�
��6�O	��eGg�ԭ��y�!V�VPH�ED��Q.���#�7�y��R�A:��%�Κc�<� ��
�*��I�XG�a&��	����R�RG�1D�\ 0�P�����6kr� �ጡx/�X&"�Oൈ' �`~��f�F�6��9�T`L��|��O�3u�b8Q����?���A�h�ki&�au�p3!��'�d�g�6D$Gx�!�	f��0�vtG�x��ϙ�ZfL�h��ţ2��2/L*y#��]&_f�� �߾)&���đ`k�x��ҍ�8@��i��}]1�FN�~t*�P���]��u��Oi�d��gӎ�2H��O�NLr7�Hb��=��< �	�2h�a~��4j`ޔ���Y�y�b<ԇ�8M�Ӱ@
3����g�ƱEs`��3$��[���?It��;I����0�y�o/x��y7GSZ��H�v��?�hO�������Co���־.X�m�G,��R�W�%�n�)�++D6�Yꀂ�+pd)b��O@�jcX$/Ơ2' �b�'��A�$G�H�\��tcȆt�h�ڴh���s)��l6m]��4r���w,�"E�ҏ"��� `�8y#�K,2�3M�+�MK�
6F�x񤢓Qx�p�"�aJ.p#�ɱaYv�;��K6.X�q&� 2ʆ,c��8A���0%��!�$X0,���5Ot��daÍ|�C(A8�&�U�'r�Q��*��6�&d����"f�bfP)�b�9����;(~9�Q!�)l ��R�t��Y��)TJ�Y`ġ��',z=i��� WRD�x�BD�^����� ����	A��*�Ms���]�����6��<z�@^�A��ı��9H�b�B��"T��r���hE�ՙF�">��1}�U+Ea�l���}�؀��FA�I�̴z�m׼�S@G͹�h�$��,Y1m��c©۪�8qQ�R�V=K�F-�O�-1a�Hl�� k�P�(�Ը�se�Ď���(�3k���m��'E~��93�gj前f֞�8�͝tl�x 5�%l��DL�/,DĈ�lZ3��W���?j�����"t 8�O�ܠ��\EO�XP��Sm�:���܉�h0��Q!,�=����2��(8���W %���^�T$��	��}7r��q 0}lN�`b?OD�q�%�4kP5�ua���aA8O�E��Aճݸ�h������ܞP,<	��ϭn`�s�$C�=~��)��3�Oܤ����Y ܒ��J X��Ѧ�'j��ce@C�$�\�V�asj��1T�Hp��C�0�!�؎/�Ze��16���l@"bW!�� 0����_�)62i��h$-�L�r"Ot�9��C~�!l@a�"O���UjH#pa��I�"^,�;�"O��ZW@��|eJ�"�/:��piw"Oؔa��L�,N�T����-�p�B"O�W�lx*f��e��B�f�<Y�a�,&�;�Լ.�`]�N�\�<�ū
,�	a��8
H���a�P�<���ϓ
���۸+�nm��N�<�t!��ˡQ�����$E�<ɵ�ƿ3Ј�"S�E�;P����@�<AQi͎S��"� ��F�YP�K~�<� ��gg�y���;o�T��CV�<��&܈jզ���ҽ,u���A�Q�<���PO0Ɉ�K� {`1�b�D�<y��i�R��2�XPe95b�D�<QI!�Z�qk&����]�<���4iԐ����}��d�Y�<y�+A?/�yh��A�����D�~�<���I�a��lQ��RT�����<��,	.6?<�c�Ҭu�,����C�<��&D�r�����c�0$�V�w�<9�a�`Eۄ��2��`�OAX�<�J$vGv铒E˘v�	Kg�|�<Y!�[$���&�+�^�b��`�<���T�g�B](dХ5zn�Hv��w�<�7G������!�Fi��� t�<�����>�(aDZ� p`�@���h�<��
�WDR	�F��"}vEp���<i��:����d�\�va`M�m�<��I���5���A�Iή�96��v�<y�]+UV�H�B^�?��82cd�<�"ˊ�[�BL���ܨ�ޑq�c\`�<	2J �B�t��c@�V�eᤥC]�<!�
�/�-ۇ����Ӣ�^�<��Ȳu�fLRQBݭ$�^R�g�q�<!U����q��[+u3h�2ˋe�<Y��X�q�D��g)R3ktܰ����[�<�E�J�&"R����,eDV��C�^�<���+��p�O�(l�Z���D@�<��C��<|'O�*Td�"bB�A�<	����)����[�qt�Y���}�<� �����Y��ģ! D���#y�<	5MR�6C��1����#%���2'Jl�<p��lyN0�q��j�x=h���W�<14%��{�A�Q@�(-L��;v#�F�<YQ"Έ6D�P���MT��rˍC�<����p�M8č�� ��0�O�k�<)%V_�$\�s��(�4�xE* d�<Q��	Y���*h�xm�W&�y�<��aɝX$l b�O [�X�y���b�<��E.˶E�Ј[�TJ0��c�< ފd���!H5�>�v��P�<)%�U�5�b�q�mR?6ȜI���k�<Q��S�\ɘ"F��W�IH�e�<Qb�3^�.�"&����)`˓o�<)�B�$v�S%+�3:��Y��k�<�� �h� 
G֫l�����f�<��E�&F��mSVg��y��ł�R^�<��w��]r���9M�qil�w�<��K�:ڀ���]L��a��r�<��`�>gP��D��m� D�q�<ѕ��<^@�ئ=�6U`"�t�<�`�F"A5,MR�A�K�|a����<�  �I��B��0��/�@f6a��"OT�ڣ���E�S �/_^�= �"O�x�6˃j*$�s%F@J@��"OL��:��a@���_=��`"O�ز��z>�� �j��"�\�P�"O�x���K?½Jw��JE����"O@���ŽM�sѐ)I��@�"O��r'�W0�ʔ�4���L>�
"ON���Y�/Wj}ī�EK�-��"Ol�8E&�D��������L���"O�I�!c��e��@A�C�0�V�6O~���b_&\�6`b�φ��`x�&�)�m��M*���!Ƌw�|ձ5fZ#��	�+�����X�-��`
��2�؈����(RHB䉝W�D)c#瓓]�������uk"�'��Y#A�z��ҧ�h�S��ȟ6��9C�c�3{61	�"O\��i�rB�4$H��[i�x������	63����)0�3�	'n�N �A�D�� R ��<�C���l�Z��t�^�A��lB�@	���a��*L���1��'k�	�$�\9I��i�N-=bI!�(��Y("��vϔ�'�\�k'�L0,��a+�G�C^�#
�'c�}+���:�*�!a F:L�H8�OjA0�B�r��H�"|b��Q$| zq(6�@"7`�06�\R�<Yp�I�r���; �Y�fX	iѯO2��'ƬBB^���Ϙ'�*4�qgS?:�����nJN�@a	�'� (���a�R�+RL�
�6}�u�	%q�Jƍx����e��`:Y+6iӨGQ(1�1�7O(�0S�۳L�J-�J�$��
�:9���a��=!��,�9D�Ժ�����^�S�B�%@QbX{�2?чB#H��ܘ�d7}��)S<vO%CQE �iL��
�a�!�ď*-ǜq�țE,j�.[���&�(z�.��Y�q��'�4�����%5$�@��8^��'���%LqC�p�d΅�o�<�[P`�9`_���I�@�6���Xw;�|��f�$I�B�I�BE�p{���o��b���+ojB�?V�l`S䌋:<K���R��� �hC�a~��'����ǝ�-��C�	�F Py��	�9X.�Y81ƇB�C�ɮ/D��I$Ć"L���.۽=�b#>����3���|b����rL���պ}b(s��R�<�w�
:`�}35�D�	7l������Q�T�%�"~B'gӷ2#�%+B�B0G�}�%B��y�c֍v&�܉�ц�T�cB�Ӭ���Δj�8�������<)��,d&LCC@1=L�i�m
yX��9��Zw�Y�"�ܕ|q��*�C�?R?�up�
�'@��d�*���1��6R�4 �U�������D�L��X�i�0(�u�Y�t�7G��˳��M�~�h����y2���q�<!�s�D�sH<D����Mca.%BzV�0&N�h�i��撛�h�k�
�#����0`��M�Nd
�`�9�!�d�=X��v�ޛsyh<���:�j��� i�YWG1,���S0Y?A�����<�Љfl��m{v]JR�\e�a}������@D 5� i��7� ��u΍�'��}QD�Q
�"HL0�O��2A��A�d��A�ɜxI�U��LH*��Y����ę��i=��S<o�7mǠ#�A&I��K�cө�XX`��-y�-I@%�T�<y �ZI �iK��\�qat+�)�������Q��}��ៗA��*pIڛI"�AE��6^�eI$�A鼋!b�.R��E	CI7d�j09��Yk��tS�h�`���Q��_��(� G���iV�ߕ`��d@E�v
zd�1	�e��Uv��'X��8� �V�'U0P6�XY%�4Y��!�R�$C�S �Hx ,ѳ"�^ )��#:C>�S�
��x��q�4m�h��c��-�qQf��q>`�Ɖ�8Ta|rH�	�y��a���}�Pm������� j���I]5�r8�g�� �W5	zP
��4L�睶R�(�'ȏ�{�(�9����2�C�	�fex#H�%Y'�<�GCL0O��[�!4�le��� ?�(�4���'>�8�d`��b} �B�yNp�1�ՙ!!̐��:|O^�!�B�
�Mz�dC��X-c'�ŵ	�l�0d��\J��;P)���'����ʙ{��� t�����^�R�U�8�H���d�j�`�B�E�?z96�@"e����' w\%�'#]����4�f��ȓ8Y���	c�r4S��ܰ% �Q��e�ٔ�	�臲��K`]e��~��;Z��Qi�]�)bL�y�����y��T�-��9B7�Y�.C�(� ��{�̞�v&��b��#�TAX��	2A���TCG�|�Xu�3G��~k����N���Y�P h�XP��G#�ha ƃ��TĲ�(�%�x`���|�b���p��g�'��Or�q�J�)�9���%C�~&���>�r�	@G�yRǨH:�ʐ	���b���ҭ�~򩖇I�4��eKLO��S�D_�-q1k�a{|$��K�d"C�2�ȥ!���w���h�(� ��'��0�+�)MV�	���O���6G���mr� �Sg(����'�&�!��۟*m�mu�	)vB�[r��\Y�����Pa��_�}��I�սlF�I o����O���� 	�A�D���!4�)ޚXaX]07C�%��y�ҿ4!���e�6.B5D���!��c(��7s�	�f�^�z�D�S�O�(1n_5"<�	Q�X.����'Kz�����n�vt b���~#�}���7?� d�$.�X�B���}����[�V�a ������C7��?!�!�]����`�uR4�ѬCjϒH "A�H���'qh�:�n^/`���X�	�џ����Ѹjh������ϗ}.�؇�U�ca�$'���y�`57Tpx8���+}0�	ѫ��Đ�dt��YP`Ц��)�'��	�G#O `*�)�phF\�^t��1��{�� /�Б��'-�K>�5K]�/��|�<C�@�+R��1�Ɨ�Z-bm��MF_(<)q`�+c*�k1�#1,60xo��k0�Ġ�"��[ HX�NQ*��⩌�HRڸq��4D��&��L���ȓf�U['6D����.HJ�K�>DX��`�.D��H4�Q��r��#��@Ð�ɔk.D�lⶫ�7,�~p�ẁC�8D���S2\u,��p��,l[�����6D��%�_�b�ze1���~>}���9�>�:Pi��'w^(�@K�9cxQY"�^�*���xb���1�i�+���^�ɢ[b�yEØ����ɼ��ݹ�����(�Y%��*���,�Iı����-P��V�����v�d���1��IS��˧�y�-
� ͈C�X������jW�u*�Γ9P�ZѨ�?�x�Џ��O*��$C�*��T��t"���B�)��|L#	Ϣh���J��n��!hK�$-���S� �R-�`��q(���#	D4W�>�*�ɤJ�f}�񢏞{��a����~#<1�`�.K����Vc�9�D��A�?��$iگ9���Bw�K+��=�G�Q�c� ��k٫v�a�	��4��Y���O�^����B2K��q��$y��@%2l�$0���5��q�pG�"[�ϧ�y��ȭ~����5S��f��0?9"�R!%Dl�3��*?4�iK!N+siN�`M�!f���#��BF���^-��@�N�*qkD�B����<1ЦX8O�|��c��&��r��[�'n���Β ��ɬ�Dpi�f�`zXc���"�b�Be�_��;� �"$���'�������?@Ihb�)ړV��v�Z�
�a�-L���$�r��9 �7�<d�ݴ: a�$��ss���-a�E���S����j� 6$������!��s�z}�%��-n�Jx`�'�u��	I�[�F��n-k%(t+�������+U���ժ"�7������^�xX���?�Γ�.�ř����VGؙ�|%��	01.�*4 �;��9��ׯl�b(�'�\<����#-trݚ�m�~{�x�G%���'���Y"��MA� ��!]��k��ݖ �AvG]$�ў��V���@��i�����s_
�
�@J ?��)���7�ұ��-N�$����B~r���@�{�'���{c�ĭT{��:�酛n��X[�4sj���U�N4^"2�D�iny��:�'X_�4�w�D6j�9�v A1:"���UE� xDp�	�?:��%��8��}��'�_Iv�`��8^�0ܻS�X5|u�@띧�i�W˲�����oy2KI;� ����-(��l��֗��>���,,h1A@�P 5% x9͚}�`<S��[���'���8Fܵ*!JF��L����mbU�O�w�x����hO13q�4z�Z#|J	>]�<=���x�G�G�[�ޝ)sꉾ��I������L<��� ?���LɯY	��2�@��<���π@Ȗ➢}� B Q�
љ[ �L�Pi�={M���f�����'v|L)sg��*t,��a���R]�
ӓ8\�j"}�
�8�� �eI<2�L[��y/��Q+���ʥ0]Rty����y2�V&[�$�C�%��Q*r�Y&�yb�C���b�-_;^&�F���y�(�V���مD7îx��G��yh	���Q(�-��;���g�yR��|T����@��l$��Z�CH��y2��e�U#���!X3�d�ƌ��yRK �c�x�H��W�ZW8�VbŔ�yJ����d�.�5����y�a�� x���̆�z���7Q9�y�iF'n�x�J��C���G���y�F�������U��LDS�5�y�l�iψEb`Þ�K,0Q�� �yB*��UH��đ�(eB���y"�O�YʀJ���3v6=��#J��y���A��̄��B����yr�M�	��y�m�{������y�c��w��E�4qv���@Z
�y��Ґn�b��!ѡZ�n��J��yR,�c�P�K��G� Ξ�����y��U�r�%��(��o�(��$�/�y���4��
���P��m�3`]&�y�ӚU�lpc$D,W`yARP;�y�ψ^�,%PB�P�F*
 �ʨ�y�,�d�&�����-�����&ˠ�y��E9A��1f��s�0�+���y2���W%�a��k�>n�.5!�L=�y2��:Ze�ܠ`I�f4J�
�GԬ�y���)��)���x�� ���y��k�ȁf��4|�8xḘ�y�����r�k��q,ܜcB�$�y�{�JjéG,jn��Q`��yҩ
 5z�ЁY�p<r����V��y�o�*|��d�K'E�~0`W��yR���t���EK\G�j����I��yr�ן����Ý�J��V�?�yRmؙb�-�-�	v�R��G�3�y�fM�hF���ĸkz��J�G �y�g�bh=��UJ���r�䑹�yrmF�PrykRM\0L����$G���y��?yz��Aܧ4Ţ-����y�P�;�a��ϊ:5Y>�"gA�y�إ	�+cR=,}���$��O�i��۴�>�i�*A�X���"O�Y�ƥ�-a���P��]:9/��"O�Q��Ά�q�D�g�k�� �"OD�5ϛ�9�$���f��8VE{3"O:)�����=&�h�2�F��"Oذ���P F�>��\6ʝِ"OHx��R���5Q�-�	{�u�7"O�QW�	37&�:F��*t�����G٦�9�3?���X麣R�?�zq藩Q�t��W�O�hPr�o��lW��z1��D�Fy��)��.�ijvE]�e��!���#km�"!�&fV�Q�ʽ<��S?||�C�H�7��-�G�M�F�����g�T��x+O���T�l�a
&,��Hs�_#[����bmH")�dj���O�1��	ɻ+ׄ �
�'�$eYt��:�!`�Y7��'�r�HQ�C�xd�ecM��� /o�Ќ��B�"ZE���2�'����WQXYT�6sS��S�O�8`�LƔ/�p�PM&u0lh�6�C�P�fH�"/����d�u>¨ò@�]��\�9�^���E0!�8(�O��`��K�'��Sr�p��6�d6�F�f�<�O�`&�f�>����9@Ʉ��t�I�r���%�ށ8��d�p�1��'�qA��0lTAr()=������� �+`@��8������}�@�`u"OzX�D֬A��d���$��"O����!���L�j��u"OfTS'nH+Bu����J�����"O؝�5�PB1r i��^�K�<%j"O:EC T�3vU)a엻3��Q�"OHhP0��@��-�V"�_m�ak�"O��;$h/7l΄Zs"�	, �;"O�=�s�9/<��go�i����"O�0@��]�e��� �٦b�@�"O2��
�x=ڭ�G�-�̒�"Oh-3B'�,/��h�D-T�HҙiU"O�S��cB��so�]� �a"O6@҇/̋p諱,[8 :�	G"OL!@��*�x%A��,x���"O�E��*<�v��X���Ç"O�ap�7-!�iQ��I�w�H�S"O�۰�D�U1���~����"O��R`��o����!C1	z�=+�"O��!�T�l���UWp\��"OH�� #�bT���6Q\�� �"O�`[�$kڦ�xA���
C����yo�=������e
���Q�X*�yC�X�N�)2.Fx3����y����gl�Dge/|�L[#j��y"D�$�����JX�%���C���y���5���Ӣ�E���RӍ�.�y�	נ"}0���Z�n���3�L�y�.݄��+�a��5#^I��-���yr�R������f�*��hI�H��yRn�Ne ����U�a�2�yr� .?$e�D�@�{� ̲� O�y�e=��Y1EJ8+f*l���W��y��ީn(L`C�twL��h,�y��	%��"��Y�oSԁxu�D��y�I��Wa�₣{)�p���� �y2F�O���K�mO<@Jd�$�y�-H<N����2l�"��v(M��y�6}����+[����`�4�yB�$.����$��NΆaI���y�$��O��aș[�44W���y�HL@��wXY��1Ղ:�y���:\2J [�'� Q�p�A5&̸�y"�!9fD��ٲt����i���y�m]�"h|�����].��z�#��y��E)�m���֜XA�}�u�X�y���_�Ȓ��
f���[���yҀ��jT���1�S�\�duj�P�yR�Q[ &Ub��W'X�T�n��y��9�� ��H�*�Ŵ�yB�E|�z�a���!A
�L�@��(�y���>Ko"l���[�6en����4�y���oӄ��$�).a�xb�M��yB�B&�:�z��+τ�B��T��y��U�yc�-R�0(�h#�פ�y�� x�fJdԭ�"��U��y�녉	G�`dgB���IP��L��y��ij2\[%-L����+����yb�ӅAP�!C�%��]�A��y�-��d���s�#��x��&�y"i�8E��~��){r���y�E��m#�ȱ3�M�rͮcB A3�y���/"�n%t
��bdh������ybjh�p�ई�60�p��%Y��y
� *@� /ΧF1�jE��i<q�"O�¤� K�	*�耘[LM�#"O�����>8���qg�
UEd(3�"O
���ܦ3�jEy�%֬}=�Pc"O�<���X���� �b���$"O��w��=D�(��2i,�"Oʜ:C�ƣK��X��I�3���"O��B�,�>�LI	�XT �;�"O숰UטzD�8r���B<�U��"OR#���0�FQ%f�t,�l�b"O���`�|y�;�$�}��!S�"O��` �'BeP(��3�H�#"O��IҾw0��M�E\0
�"O�I:7m�&=������\&�N��a"O���h��YyTM�3�E&��P�"O4�2��>2�I�̖�b����"O6�⋜h'Ҙ�#n�;Z<��"O�t)��6j�鸓,�b'��V"O$���;��9�v˘5?���"O��C&�B@��i��{����"OX�jP�T�,e �X�&R��8���"O4aе
�0ܨ ��8q|RI�"O,��Sϋ�q��	��BcZ�"ON� p�%ir���Ƈ���T�"O�� h8zA�<��EK.A�T"O2��v"�~$>�Q���/�t�;�"OPe�#�Dv`��jD�~֔�@q"O�����N+IR`��bB���"O4�E*W�P�T��Q��#����$"O�Q�;xp!��/�:R��*2"O�!�&�X�Z6�u��͉�@��"O$�y§�Iq���C���R�g"Ob�K�#��Of
�� �6��Y"O�T�4��5Z�+c�:w��*E"O$�c�!ǥ&���JsD��i\x���"O��t�	'[�00�zL���"Oް���ס�t	�q��M(z�y�"O�xUC�	����j�m%���"O�t�t�͛�J��C
M9)�U��"Oly�q�:��͹�	�s#���T"On`�eKA�[�����ԀW4�ї"O�렀��p�r�I7�B:��#�"OP���@��e!A"�-�P|�g"O�Ƀǜa�!j�Nh{�"O�|��"� �̺@�9n�H�sV"O�� ��c�j�H�o� T��D"O�ŉ��?h��(�/L464�}H�"O�ؓ�N�$gV��e�+#*���c"O q 0A�+GŔ���dGd�6�<D���o��V[���g![�)d�L˅a;D�� p6kgj��\@��L@E�9D�4pF�L�}�\��-Ů]���qI-D��`S�W��8����Ĭ=x��V�,D�PZg�M�T�H��O8K���+��-D�����	�(! �	�Y��}{�)*D���AO����� J*|�V���d=D�<8�� �*�t�� �}�(b�:D��' �>u~aHp���I�����j-D���&N�)]������;5��Xj� 'D�p���
��lBN�/&����&�%D��3�!���'+L�t�,��%D���)B<FPX�@*�0�����?D�1��
�B�*��X i~�d��;D����EM=AY�F"�>@��|Sr�:D�� H5�A�<(����i
D�D"O�(G� 4��*R�o���"P"O�� S#i�)_�O�8`�"O�B�O�,z5ܩ
��1
�@
�"O��y��'Q�̄�`H�<h���#"O`)`��խ-\3�# �B��q"O�dy�hń^t�%� A7,�laB�"Ox�[B�"iq�h�!$
����E"O�A5I��y���
�b
�S�����"O@���$_x����`;9��z�"OD0�@a�j���)`o+��r"O�A��,׷}3H\2���kJ���"O��0�N�g����f�� :��"OB�S���0��$B�e�k0��A"O@�#/�3��U(�n��y'qY"O�ғhW!i�"ѳ�A�As���"Ot����٨yx"alN���"O�)�:)NQ�˒	ZRb�(�"O$.�p�	 *�]D�"f���!���,X����J�������!�d���a���c�6�u��;r!��?k&�:��'	�(��u/{d!�\_ ��6'S�v�$q�G�,R!�R9`�����$�����E�P@!�$J�{*(��-'c�>U��A��#R!��f�V�%CI��b�0!�Z;[y�a+���:m��8Q���!����x$i+`a<��E�!b�!�'=��iAQ,n
T�wEExA!���!:p1���#[d mJQO"!�d�@����`�
*\�\s��	�Py"j��F�)b��*`HLs ��yB�s�v�Tj2(�p��� S�y"��.fD0�u.����&�D-�y�.G�d��������}~PXG��,�ybI
~3�x��+8��	B����y�'�+�p%��)2n<�/�y2����2�A/lz!��]��y��q)\HS�")�R�nB��y��E�0��❂	<��*C��	�y�-�+#Č��@�2 �써B˜��y"��q����Bu��Qr�:�y��S��t+rhW����Q���ybeޛiW&�Q����H Uт�;�y"�K�f�m�u	/� F'�yJ��hLX��h[�K�LQ��y�^�o��q����a��]�y�h۩:x|�ie���b��g`\��y�cÿ_����n�~JuG�o�<A0I+
�M���Q�p�3��\�<!#��v�z� C��;cJ����W�<I$�4�����Ș8:>���.S�<��*ZV�<��Z@��bģRR�<�D�a,����K%b�&Ir���P�<�1��
j ٵ���sRA�J�L�<ɕ�&l�Z��ƙ .�llhQ�GG�<12�ӑt"�x���R�"��F�<�#�g���(��0����F�<�P .}	^�[��V�jo2�z%��D�<)c�"���ƌ�*b���:7�\�<ap	��j����گ.C��R/GX�<i���#O�8D@��'%�	K��~�<�f�ٌ,U �)`霣
���*W��A�<��O�K��p�V�;k�j��4B{�<� 4�T�[�zZ��W�]����"O4��WL�uL=��ɔ�A��u�"O�t3��ٷ+�L�i�g�/yX�QA"O֙Xd�W?e� �%�Kqh��"O$Y�e�;e��u�H	Tî���"O(�� 쎑�J�r2�ۛ*��e��"O���&b�u�q�ԉ:�Fu���B�<9�)7;'X8��˂��D�&��<��ݬ^�|�1,��Zl��ӵ��{�<����BMHu��P5@]>	�"l�ȓ� � @�?�   �  Q  �  +  �*  _6  �A  tM  Y  �d  p  �{  Ɔ  �  P�  �  �  b�  ��  ��  >�  ��  ��  ��  t�  ��  :�  ��  ��  �  \ � � � y �% / �8 �> �G nO �V �\ :c ;i  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�|��'����F��a��������yҁ�0��(�A��>@j���S(E��y�M�-o~�C�X#?i&�s�*�0<A����	)���̖7����vW+^!�b,Q���ؐ4l������Py� z�ЩW+�5�)Bc��y" ��g[�䋷�ݘ3OΤ���y�G��@���ף�8Yj�� ���.�y�/A�yz�97O3H�vyh�{#!��J�:x���� ����RN!���8 ��]K��ʙ�2'�<c!���`L*�*V�q������ �P&!�D>�dY�Z�T�DH22��!��!�U# C]�Q׈Ł����!�d�4���{��J���7�I:\�!�d��x.��)�J��W��<[7��]N!�D�r5�	Sv�)~�@H	r�W?!��q5R�B��\�b��
�N��A!�D�+"�@*a&�&7^({�m@.�Ia��(�n$�,Q�+�����xqԠ
�"O��G+�Cΰ%�Ek�
j���"O���[�Ȉ�#��'�`cGB���yB��B:�8��|\nt ���)��d9�O�RRGq��H��D?( 0P�'"��(@4���B�ҶiW8yX��w�NC�	87WX�`�jE��
���(��?q��)�&�b�@ś��%M�cb|���� L���Ȃ/:����#6\@I'6O̢=E�t��,JL�t�� >!��2┇�y�2^��03�1bQ��%���y�,�o��Q��	�zH��������y��bat�ɇ)I�s��9c�����hO��R�h�b� ?Xz������0�"O����oL�P0��s�@��P�� ��Lw�����R5��Ыc./���e���x���N��U@�Ɗb�������Ḧ́��J؟�y��(v��C��8]f�T�f'<Op#<�4�GP/�d�0�,GŠ}�WAI��� rJ�9� B��0�&L�)�bl�Ia�����Xؗ���p�	��o�0��j-5D��"���_XB���.��[���#���fh<u�E	n�ڽ���	#�4�� �h���<17�I�0�Ҙ���g?�$-$�M��K_i� �<��)!f�q����=)����ܒ$��x2��;��)(��ӭ�y��_�xD@A�
h~��(!���y��)�v���睑
?*-����bV�8�ȓE�m;s#�4>��S�'�C7�9�'&�=��w�܋t$]�|��ěg��e8���N~�A��<��*��t�\ңΑ;�y��F:5��2�	7i@�Yc���y�F^�o�0�맡��RpSs��y��Nm�Y��e�2M��k�	���yGx���G�j&�0&�;j�LQ�u�0D��qc@@"��b�%Om����1`�>i�����(E��&~ MY��F{
^0���r̳4�@��<q#������ȓMkx)����; ְ�%$_�1Kv|�ȓVB�p�U����q�#1x�E�ȓW�4y���;� @�� V#�y�ȓ<�D���
/^!Æ�@�8�ޱ��m鮬0 �� �<��p���u �E��!��qg��)@I��Y�66���ȓW�P�!�끅V�l!V��++(L(�ȓX��,Q�B�$_�	�s������ȓ��1zw�Q�5EX8wI80�����j~Y��.�K?�� k:LK�݇ȓT�R�ņ1
bAb��ƫ4�`��(��)���9r� ʗ'�*|�<��oQ��XQ$�*Ì�F�K�aBf���M�ب	�!��O� �1a
	05�8H�ȓ
鶬��+ؖ:�ЅѷJ�/�&L��ZF��5 %IJ8A1`֔d�N��j�Y!�Ԟ!�*�05/�i%`��ȓx	�xk���60w����Hh��ȓ}��J5f��2�!׮�Sk���ȓ��EѲ�A1"��R)=4�0��J�^��gB��<Y��ҕ�޻u��ȇȓz2-X`�+��TzqJ��Fv�5�ȓ*��������>)��3��5��Ѕ���&��@���H-6h��ȓR����� &s�����O��쑅ȓq�fNE�t3��i�R|�e_W�<)Q�V�+xs֏��j�����{�<I6
ͺ_�Ĉ]�>����WGN�<)�����c�!��H� �p&f�<��#�&�|�pb��#7���FΆZ�<QB/I��Zu��&u��� �VV�<����1�>Y�f�	2$�M���T�<�r�E#/�Ҍ�F�~ Ћ��S�<�Ə'M�`�1e@�mq�%�R��T�<�  ���K'P��xC�QRPqR�"O�q��L��(Y�sA�2B�m9�"O.��&������2!��6憱kr*OnP�уu�R�b��^�[�>͙�'�t��"z̰�вfɲUG�U����?���?q���?����?)���?���mfƐ8�撞v��H�O�%\���8��?���?���?����?I��?i�+��8��c�^?�`mN-]�:is��?	��?���
ߴ�?Q���?���?1�@�CQ���	F�V�j�)���?���?Y��?q���?Q��?9���?�D�^ʝ٧��&��
3! �j�$�O,�$�O|��O>�d�O$���Ol�����U(d&J�#�h�"�/R����O����O��D�O����OD���O|�����-�U� ���P�*�V�d�O��d�O���O<���O����OB��j�`j��U�E_|��s�h�d����\�	��Iϟ�	�Iӟ��	{���d�YO,�e�B�֡V�^E�	П���؟��ş�����	ן0�	�&��HB!$�'�r��p�G1]�W�����X�I���	���П@�	���Ϳl���vꐾ*�I��@�ܟp����0�I��	��t��Ɵ����dP!�H��&.)D�Qa��^П������Iԟ��ߟ����x��ҟСE��I��e�a��Hy�$%�ʟ��i�7m�O6���O����O@n�����I�RI�M	�	C`�Ӗ�.l�,e#-O$�d�<�|�'�6펯D]�=�3K4o�D}��J�=?�N8AǕ�,Zڴ�����'g���mYv�Y�I+:��X8`�cN��'M��k�ij�	�|���O�B<�(*��s�n$�efH�6��<�����0ڧ����$&�-���G���"��JҾi�$ḍyB�����q�:4�#T3a%@���J�-�I�`ϓ����N���6-a�l@Ӫ���Zܣ���21�����`��̓�#������'����b�m�uR�lŮwY����'���r��6�M{E��J̓��"#iT�O�6����>f��,�R.�>!���?y�'��Iz� �J�@N���h�'��f����?�Я�%�^=�|����O\=��Mʐ��]�a��y��T�oN��+)O���?E��'c~99b*�;X�xe��&�sQjD�'��6�����MS��O��t����Jj:�0�
A)=� h��'J��'�"ͽ!������Χ��č֒W2$	ХE�	R�T0bØ+�(%�P�����'�b�'H��'��h�(ŐF�����Y��F-��R��s�4)��8��?!���O3�$�7K� ��c��ʲ�`|��>	յi��6�L�)�S=�8O�6~zl;N�"}.L���h�+��`���c��5�'�ľ/�6���+��M&�˓Q���q��.Jes5��E
@����?����?��|�(O��l�ԁ��-J�t���$�vu��
�)����	.�M��ɾ>��ip�6��妍�)͸5z����K��nʜE���\� H|o�D~"��rw.X�S]���Ϻ�;`h�樐�V��L� �]�p��ϓ�?I���?I���?����O�9�E!إI�t����ׁǚz�2�'�b�t��5x@?�"�d��Q$��zf'�k��P����(2��1������/S��d���ىz�6-#?1��E�H���v����?8�%`7!l����i��˓�VX������	�H�&	K�#�L9Q4�خ���3��ޟ���Yy�iӀ�����O����O�˧uJ�å�J9�4$k3/ƐÀ�'/p�U�fi�f�&��B�.Ḇ�ޮ-�f�⦎�>ef�0��5�2�+s�m~x��!��'3hM��yǋ�;yK�Ib���
� �Yq��"�'}��'���]���ݴ(N�I)�&��#�4�{����	9�iJ�g��?1�E��&�d�b}��o�F	�&�� 7>ip�0��\�b��ش�,�{۴���D ><a(�����2e�P�MS#X��`���2�h8[�4���O���O@���O"�d�|��	<�,���H�q�-�A,Ԅ
ʛ�ɓ<^�R�'8���D�'�7=�H�2���0���OԚ2}$x��ԦU9ڴI����O��B!�i5�D=
��鸒숫? \ڔ�ۻ!��ߎɤ���Jy��~:�6U������j�$�\���0���oG�t�	ߟD�IEyi`�P�N�O(�$�Oj"'Έ"�Z�I�j�2�F����6������ ݦ�K�4Pa�'�A�(;Y�2��9yN���	h����,#��4�$��(��ZG�[��?�Ԩ�O�t[�ˇ~zi	T�1B�`q9��O���O��$�O��}
�C���Ae�	=>��
�-��x�Q��vl��	T��'�"7�<�i�݈
]�%<�ݫ��T���ST�n�$Rڴ��&ng���֧n�J�p;����H��\�n�8Nm���"�bx�)d ��$�̦�����'s�'�r�'��<��'C-��-8%B	$��hAwZ����=�f�	����b�韀��ɠ}��ث��8�	4'B�D��ɞ�M���i��O1�T�;�G�/:kz�PC��C�P�$��5a���c����M�j	B�Oy����˓@F�5 f�U�$T���&?^�R��?a��?Q��|z*Olmn��!�j��9��J��T#��kaA��<*j��ɥ�M3��+�>��iJ�6��Ħ�@��ٱ0�*���=�U
@� &�n�<a��I��A���ej$�O?1)V��� �)$�N�HZr�ؒdX*n[���:O����O����O��D�O<�?��e �� �tIT�J6&�:����^ڟT�	ԟ|2�4(����'�?�ӹi��'^Ě��8�@ ���Z�MdR�Ct�%����j��|��ɕ��M��O��3�>����$sS:���I�u����:O�!@�fT�$�	��������#�j��կ�:5��8i$a����Icy"�x��-�Š�O���O�ʧ�� �h�Xi��":%�$��'���e֛�	rӌ4&��'obB�`��w\ Rdc��t(�I�&&T:�Jť��d�غCq��O  Y,O�>;��� �hy���W�Y���#�'���'_����Ow�	0�M�d���<��M@#I
���Z�H	�s�������?0�iN�OR�''7�ãY�����f3L#p�q��	1��1nZ��M�e���M3�O���Ħ׳�Z���<�3�ũ-�\��@��dܸ���'?��U�$�	̟\��ğ����X�OdFl�P%w��G���j��c�"m�Jh����O����O��?����KFI�0���c8vp�B�Č$����sӾ�$�b>a��hM¦�ϓm6�ӤN� t����*��CP(�ϓI�T`q��O��p.O<�o�Jy��'�BZ�U���zQ��}����nvs2�'���'���;�M󐡍��?Y��?!�h^�P����NK=/��"``̳��'-$�0���}Ӹ�&�lBQnݲ3��5��ښ(�8�� g!?I`+�5/�@�Ꮁ����3r-�O���l2B!"'+d����Rgԧw0�̺��?9���?��h���d�$/:�E ���!
��7W�<�d�㦡���U��p��.�M���wv��7W�p他��&�02���<qq�iWT7MCɦ�;3�ϦM�'J0#�J�?���x�h�B���fTɀ�]�/�I��M+.O"���O�d�O\���OJ�"e�M? ��cp��qv�	�C�<�a�iy����'�'x�O�FD�w�QAb�X��$�@�DBl��?�4$ɧ�B��e���X���Y�4F%QF(y�d���=���*OV��Q�?9�ʢ<1e�i�剚~�4x#����M�$�d�!E���	�h��ɟ��i>E�'j�7mZ<-���{VRY��)�(w6 ����f���Ц��?!eU�l#�4 c�ki�ȥ�b�̅���9&'M�Z-T8�ϛ@P6M*?q���>}*���ǧ�������BK����Ř0����ʽ`|��ϓ�?)���?!��?�����O ��SV�P�M}h����^5Θ�F�'B�'�x7� k���M�O>O�1oR��wEQ%&_�a&̰���?	��|���S>�M��O뎗ff����f�Sh�D˸XE4v����'��'���'���'S@	�$%�,���U�u���Sbӟ(�Ivy"/g�A2�)�O��$�Ov�'4L�L���ԅ����0x��',��?A����I�*cPP���dzM�6�̙<5b��%(b�9����-W�o�I�x�H����/g�8ܺG�z�j�����I�<�)�hy�cw� )
sa4=�iK��E�!X���	������O�l�C�=�	�d� ���f@0�/])t����R���c�4m 8���4����+ ���������B�H?d�|�24��P�q`Du��'�'���'���'c��`]�!���8�Ms�.�P�4&�� ���?a����'�?I ��y�Δ&|�y4�L���T2�霤m�H7�Ϧ�:K<�|²�˭�M��'�a���&l]�A�c��� ��'y�MʦGZ��ؐ�|�W���I͟@�!l$&�Ճ�C�*s��ݟ��I��H�	`yB�`�̑�%�O��O4��E�:[�-;����!Ft8e	"�I������J޴/��'"�� G`���2�I[5���j�O��u,�'D�q�-�� �?	j�O.l[�k��.|��;0ĭ���O����O��D�Oh�}��]��P�!m��-!�XA��ʲW=���>���Cć+K��'�67m/�i�)
V�T(P��H<j*��U�g���4%�6�fӠ���{���z7�P�ԋ�����a���\D��*f�_�k���#�������O��O��D�O��$��e�K�[�bP0r���BHp�`Q���۴��Z*O&��4���O`գ��C����r���$��*Sx}��wӌ!l���ŞݰA�(����E�.�,�pJK/b�\�K*O2�� ƨ�?	� ���<��(�)������n�� �����?y���?)��?ͧ��$U���� ��ş��U�"uMhu0��(6T"3�ϟ��ߴ��'���!�V�l�x�nI��)Ƹr�ma�˂������3�֟���SO�K����k���9��G��6�ı��&ۚ�&xp�d���Iş0��ɟ����,�:�!I�-��L�Bb� ���C��9�?���?9��i��2�O^2f��O���$��f��k�3d�Ht8�Np���M#Ʊ���B̴xf����f�	ui4l �"�א��Z	���p�' �I%�̔'S"�'#��'/��ie.��7�T����XgZ�aP�'�BZ�X�ݴVo,����?	����-k��� 7S??t8��΅/
b�I�������ݴ#9���	��4`��%�Z����f�Ұ<�Vi;B��1(��E���bWB��]�~U�8�����t3�D���ה���	ɟ������)�S{yb�v�ZȻuB�f�PӕO�*�B�(�аi�&�$�O�l�h�<�I)�M �R����oA<���R恙s���q��c4(k���W�:������π ���U�6>..t��$gg����6OB˓�?Y��?���?����Ɉ�_&��3�\5W��1֎Q y[@m�e����՟ ��S�S՟�������i��H$��+c㗏E.�y���^{���d���$�b>9��/�Ҧ!�\w����C�2xbrꑉy��̓:� ����O ��O>�(O���Oz������(H.�b1�d�޾"(��OH���O��>A2*��?���?���:k؞��4��:&��Ũ�a\��'�{ٛ�Krӈ�&�, �ūA���7!
�Ʃ��N+?�/�9�X��-�e�'3�V���%�?��ќr�K�W��Q��gRKZ����<���4�IR�OdR�����t���4|yX��rE��=�rg��t��O�O���]Ȧ��?ͻv��(�GJ�8@�Ód��C/t���?q�48H����U��v���A��ɤ=�$D�����̀>��c�����$�ė��T�'*�'m�'�"mB�#�n�����ٖ*�`�ЄY�<ٴX�~P�,Od�1�I�O!B��$
b��-�;|@D8�e�g}�}�ҽo����ŞQhƉ #�X-ttp���R�?��h����A�'|�Q�a�����|�Q�${�CA�m(���K6�n��M����	�,�Iʟ�GyroӲ��5C�O`��kT8�0�C$T� ��@×K�O�o�G��W��	�Do���M+��\�"fB���u�t�kb*��OC@$�ش��ĉ�E��(�'��O`��Z�@}oʕ\樼IGH��D�O�$�O\���OV��?��#|VHp@F	4���T�����-��şd����MS���|���|�֘|rAB�Y��	ا��g�I���� z�'����T@�jW�6���ݐYu�q:�Kܻ���`wDX=C�tIZ�ǜg?�N>�+O����Op�d�Oų�MW���A0F���?��(Щ�O�d�<Դi����'�B�'��S.g�=1u�0m�Fu����*0�O�9�'���'Lɧ��<E�t@��ٽU��!��+L��#����!A 7Sny�O�v���h��	�bɊ>5\m����b� 	���?a��?!�S�'��S����!��g�d�	R�G7��x����&� �	ߟ��ٴ��'�\��?���7�4�����+����_��?Y���dHش�������?ї'Q  ���H<�@�$	�I2�'�Iɟ���ğ��	�\��R�ԉ�8ʲ]�/��zk�@�ь6͒�s����O��2���OD�mzޕ�'�ϹDX
��G�̌r��Y�
B韜��X�)�#�<lZ�<�㛺#�L=S�˕�w� ��S�H�<!B	�30�X��L�IYy2�'����|ui8�jG�xɒe*�O�@�r�'���'��ɂ�Mk�$��?����?�V��fw~$sL����ېJH��'2z��?���I��F
��:�pT[SO��b�
!�'v�Y�֢ϱn��Vl/�	��~"�'�ܸ�	�i���@��E)aTp�1��'���'8�'��>a�ɢT6���5H�a c�c�T���M�2eYt~"�w����)7g怃�E�	N�]���M<�	��M3�i\�7MI�)<�7�7?ٲ�\%� �	�]�n�طc
�DIqk"FT��M>)O��OH���OL���O.i�6�˴/�ĝ��LM!.]%��<qնiތ0x�'�r�'���y�n��cc4�Q'� Z���x�]%d������i� �'�b>����Ш朴󰦋�R�*(�&��+�n0?U�<Z^��� ����dB3 ��ҳ�� �:�K�..$ʌ���O���O��4����Fl���y"�U3a�2Q���Fv ��o��y��q�J�ˬO�9lZ��M��i5����F�"z�x�c�؎uR�yKe�_؛���T1��lb�d�������b_�	m��ă�j�8 �?O����O
��O����O��?-�B�J����RbLEP���	p���	�`Q�4&����'��6-+���&<hڍ �^�'�p\��'�"�>i&��ܴ{��O�:��U�i?�ɤM,�XS��ʎ�R�����'W�x��nտ�R*{��~y�O���'�2$�Y�$�C�L�^���p�Ai�'���
�M��+�,�?��?Y+���r���48��qJ �x{3��б�O8o���Mk5�xʟh�)$a
#?�<��B�/�lLB�FF�F����ճ����|b��O<��H>Y���~\���T$ȻP ���g��?���?	��?�|b/ONoZ'����0JQ�[���I�OM1WW�t��Ο��ɑ�M#��&�>�3�i�@���o�k�DK�K�,T���=����o�x k�j�0�_~��q�d�2T�*O:|ÄB�+-�vղ�,4uJ�I��4O���?���?Q��?������օVO}2�e�7�H��M�umZ�Mɼ@��� ��n��蟔����#��I��I"��-o��;���b�&E|�L=%�b>����Ӧ�� h r�D�b	�=��Ǐ�oq���!�X�נ�O�ؒL>1/O&�$�O�a ���CZ2	QԪ^���" ���'���'�I�MS���?���?�WB^�z�����$i:������'4��j��e|Ӡ�$��1%�o����`
]R ��<?��U:N��9Y��[
��]���$Z��?9M�
.-��q@6�
������?����?Y��?q��9�:���J�kJp�2�C�$-{�&�O2�n�UI^��	����4���y���[���s'��"4V����yr�{Ӯm��MS��*�M��O`��d�Jt� �L��W,�@��B�^ mjU� �d�<!���?I��?!���?���8Q�J��A�~Y*)i�����ͦ5sQnIʟ,�����`Gj�d%� �B�N�Nx�U��b���t�	n�)>�2�rG2�.,�xy1�Nc�d �'�tـd�Q?	L>�-O��b���JC�D�!S S{�g��Of�d�O��D�O�)�<ɴ�i�.I:W�'T���O��$�`13 �Τ<j ��q�'߼72��=��D�O��4�,�ѵ�Ԛ���������U�ʔ7Mk���I<L6d��۟0�����c�Zx�@��10��;�H�=A�v8̓�?Y��?y��?�����O_�K��E���)W��r�R����'���'?|7���mU��O�oZN�I�N� $� J��L���j�BV�3f29%����ԟT�I��=m��<��O� 0����=4�Y���T,��A��[���'�d�<���?��?a��$I���p�Aɭw�6�?�����A��l����������Oj~0*"��r72�7��%K�O<4�'���'1ɧ���'-P��.q��d:2�(�6ju6B5�i�����a���$�L�P)��I��4�͐a^zd:�����	���	�b>I�'��6�M*u�j�b�c@A���	s�dx�d��O������?IQ�H��96���B`��DATU2#d�::���������M����u�fPDC�i�<)��-!yN�:��$,���(�m_�<!*O��D�O�d�OB���O�˧wA�e30��=�&�	���0�����i�����W���Iz�П Y���;�P���)�M��}��q�V�A�F�pӎy'�b>����Ц�̓7��"h:$���7�E(
�.�ϓ#�F�IsB�OT��J>Q+O��d�O�p���]vI �#��y1���OD���O��d�<q��i������'���'�R92�m^.O��jO9>8�U���$Bx}�'~�(n���K�y{�$Š<>�i���@�,.�'||����G
=ZXr��tg�ȟ\r��'�Rո��9h��2u��-.���x�'�R�'��'��>M�	(uzB4" � (�i��(HzlT��I3�M��X��?���D���4�,�5ύ=o� ��a"?%�lEq�3O���O��o�ye~�m�O~��K��$�ӯyϰ�X�S-�q��� �3s�	�|�^���ڟ�I��矘YGg��;d8��CK�0N�p���_y"�r�bAQ�<���'�?Y����[\���˧��i���B0A��I����I���Ş?Y�h��Cʔ=Rѳ��G;M�l��fmO/A9�x�'���3�ߟH�|�\�|�t�K�K��p��ΰ�5ń� E���'"�'U�O�剷�M����"�?!P��� �" �ڜC2�1 �n��?!��i�O�p�'3��i�7�O~偁4:�8/	%-�LՀ����Iϟ|�@Y����7?�����CE�[;[.\�6�׋tTRE���Z�<���^�Z�l�#�&l�P���i�qJ��?Y��)���B���ɍ�Y%��K��3����7�M�9�	��c=�ēnr�&�n��ŰO��6m4?�����|TY�OEڠ�`߶S0	Æ��OJ�HJ>�.O����O
�D�O���t$�8e	 ���T:'�vQ��	�O�D�<��i�D�3��' ��'��S�1| �H��X� i��O�`���5��I��M�iJ�O�� ����CƽbFք���.��R��;~T�(��T{y�O@����S��'�X|�t�6�$M \K��Y���'���'�2���O��	#�M�ԇ��o_�A��(p�0��h�8Qx=����?�i��O�)�'�rdM������&K�6��v���'R�'��AI��i�i�M���Nf�(O�9QC-	��m������廗1O��?���?���?���򉄱�Ɯ��DS!qW��Єl�Ox�0n�
��d�'���Ob�Sܟ����!�i�b���ڕ:5����GA�6�vӼM'���?A�S3aO֑o�<��#O
�%��E~��b��<Ѥ NQjL�dŮ����4���dЌx~��D헤$�!+�/YM�l���O��O��i��&�����'�2���83�4���ى��!�WDZ�FZ�O��'��6-��yRN<e��b A#1gǶ4���r"�o~bΣmFh8�#D��ON@�I9�B�h���#Z7i�ȩZB0&��'cr�'r"�ܟ��2`وB�	kӬ��AT�AK��Eɟ�9�4Q�����?�io�O��P+#�@P��8x ��1D�։��D�O�7M_ݦ��������'��� �j��?	�f�3+:8�c�H�y�%��B�vj�'z�i>��I꟠�I��I�Yd��â��6�(�V�R��y�'��6M.+�d���O~��3���O�,(g�_��n�q�G/|@�e��Gy��'���J/����L�R��e�r	��LS(���!>.��uNY��$C�M}hq��,�,�OnʓPE�XQ��=��9��(S.�����?����?���|�/O�o�	����;��ܠDO߳`P�EC.z�Ҽ���Ms����>9�ix�7�ʦ�c�����:���揝o�h3`M�!�~mt~�̀5�Љ��l�'����"�N=��UV4�hcK�<!���?���?!���?1���H1�p�r�#H�(.�y��B��&���'0��uӰ���4����Bզ�%��� �ʀuh�*m^ �z3����%؛&�m��	R/a�6�??	3�Z�? :�Z����O��Y`��1\��T�P��?YD�:���<ͧ�?����?�`���+
P\��KGi���r�!]��?1���D Ԧ��1�X�������4�O�B(I������`OA#A��A�O�ŕ'�"�iF�O��N��{�O�.���ZÎ(��%{�oؼ�2���*&?ͧt!l�dW�����0��#85X�d�R������?���?��Ş��Ċ���Wd�<���/��]���O*-u� ��O��$�Ц��?�wU���۴Z���h�"��^1vubg[�rI�8��i%V6m�u�r6�;?���#R5b��9����˴L�K��o�=ୂ2�y�\������	���֟��O2#4L�+[�l���I���;jK�7mt��$�O���!�	�O�1oz��+�JX.T�Y�&�qƄ�$ھ�?Q�4�ɧ�9 ��4�y����l���� L�"<�!NU�y�ˆH ��ɖ��'%�i>E��`v�)��/O�,��D�p�b���ʟ��ȟ\�'f��\�K'�'"2����hyE�׵7W~�#�	K��O`�'mB�'T�'�8�YM�:0|�1�H��H����O� �`�U�=��6m�c��(y���O���f�;P|��d	S��y7d�Ox�d�O���Ob�}R�X��С*�I�񨧮I�Iu���8��6ҩ�"�'��7�.�i޹jr�T�G�r9	�.��I�vbh��h�4c���d�%�P o���~%f}[���Ƒ�F�30��ܙ�@{`@�����4���$�O����O�ͼ9�b=0�ݝc��0���)t#��Q=�Ɗ�d�2�'���'L�����D���;���	a?LqJ�B�>���?�I>�|��B�	�V��$� G�6q:D+G?� �4'Y�	!Zg ��O �O�3�1��3�(�f�R�w�f���?���?���|B+O�1o��s܈��	l�@�z��Bp��J5Aݮ>d�����MC�r�>���i;6����vM�� i�@'z���W��n����IЦ���?Qw���m����>�������#YD�p��`����D�t���O����O��$�O~��0��!oƪY� ��0h*�=��I9� �I�<�	0�M�cGS�|��uě6�|r.��!h�-c�ʎb��ۖ �.��O�$mZ2�M�'"���Qٴ��$\-B��9���V��r�P��>]	�d��?�`"��<����?��?Y�@�G�haW��:�r�:��ݑ�?�����d]��]��uy��'��Sf�r�X�㓦[��X�������Y?�� �MK׼i>�O�S�nj��H���6'TY+�E,���&Ϗ�Jqi��Fy�O��ɉ3W�'Ô�����mADH�CD�1M�����'���'���O��#�M��`�-�,(g�A
Z�* �̻+
�����?�a�i�O0�'76�2A�8��Ci��S�\�W���|�0%o��M[C�+�M��O0��S	�3��We�<�� ��?粬XR��2j�J0QD��<�+O��$�OP��O����O �'4������X��jC"ގ�#��i$>\���'���'b�O��Fy�󎂛9���2
�v�P� b��3��m�"�M�r�x��$-�=%���3OJ�F(yʌ���q�L�[�4O<P����9�?i�j-�Ĩ<Q��?��#�P��<CD���wn���7�A��?����?�����DW�uH'��nyR�'���+��Z�$�:T�R.��M0��$[~y��'�֠2�;������� Pi�����X������䳴ω�?�b>���'+�����w���jFBD�me�H���?82��	�p��៸��@�O�@	�J9�	S̔�"d,�T�4#��r�J�@��O��d�צ��?�;i�{��Y=D̪�w��V^R�̓78���y���o��V�80n�B~��4����Sc�N�5!d���O�%�(l���|�_��؟H���@����D�%�~}3���0!��T���D]y2�a�Fq+f��O���O������X>�8�$��*�䑒��{޵�'a6M��q�O<�'��'|�<�W/S��	A���>`)��B�?�1�'|8�_ǟdb@�|�_�<�æѧn�R<�D˚�8�qK�֟�����I����by�$l�������OԬ�@lS p��[�kT��:\o�O|Ul@��K�ɐ�M�W�ic�7�I�V���3��-q����ҏ�`�D�t�g���d��d�R���d�>9��-S�`�rC��u������q��I��x����	ݟ$��{��qi4�
$�	��Lz��LD3�����?�����F@,��D�'Z7m �dٿkb!��ϓZy�ఀB�%���'�@�	��|�ӖpMl�<��d����i�$_7��Cw!A�>��5��&_!w����ϼ����4�X���O|�Ĝ�5��9�0�06O�d	'��?{����O�ʓ0��l�h�b�'A�R>)��-֟u��$�&%!�� {�.,?�\�8�I���QO>�O�,X��b4��ԊV'���Q���304���.��4�LhP��Z�Oh��U�
n�A�#KA'#2*M 1��Of�d�O��d�O1���<���m_�J>5QǃG^�
q��Ԗ[9�����'>�(r�f㟀*�O���}5X�P��
C/К�,$�6�'�
7M�Q�6�|�`�ɩBI��f�OdR����c��n��V�
	-�����D�O���OR���O&��|��	�`&���K:7z�@��	�L����B����'����'�6=�B�pC�q�9#�M@�k�H5��!�ʟ oZ����?��S�?�C�*ͦQ�S�? ��p��3,���;�K,HF�"1O�=��=�?��@$�$�<�'�?I���G�2u�G"D�`�$�ه���?a��?�������;�A��p�	� P��4�rqZ6�Z�r����A��hu�	��M㕼i��O��s@̀
z���a�w�b(q�����gCC�pX��S��@�rQ⤞ӟlJ��Ç"u��I%jU�+��q �g������ɟ|�	՟�F���'�"8�p�_�
p���_��P�e�'�x6풁Y�����O�l�v�ӼS��� 'V,3aE�7h�0�RSA��<q&�i��6MZ��5J�ʦ9�'�rA8�$��?�Tȕ�/�PbrG؛eU ��U'b��'Q�I��	՟P�Iǟ0Γ2L�Djvg�s>�ѡ���j��'SX7�@�2���D�O:��#�	�O�yg@�Qhhx���WT��stU}B�c��}mZ���ŞF�X��h��������{ӎ#?�R��,O�J�I��?1U*:���<YP�X/N!��	U/� {��4"�D��?���?����?ͧ���_�%b�� ���l���p�* � �Js�@��i�4��'P��(�mmӖ�nڼx*9�����qB��2 �P�YQ��r &���'KfeQmA�?U*���t�wm����F�Q1h�BL_�/tp�؜'��'���'Kr�'�eBP�I4�m8�+�RZXQC!�O��D�O��l�kG�Sӟ�{ش��]�±��Yu�ZQ�T-�N� ��x҅zӺlz>��ed�˦e�'�d�k3�_2"-����(T�mb��.u���	1Y��'��	�������	�2c���hR�]�D|J�AĽVf���˟Ж'��6�q|V�$�O$�D�|��kG�L2N�3��ͮ ���`�'VD~��<����M�4�|*�8�%F�/<�����C���,��=bX��gg�xD���|�1��O��H> �F�3��cl����q�I��?y��?y��?�|�*O�`mڕD��0'��Jޑx�³xB���⟼�	��Ms��������M���
`ј��A��4������X2�6	zӨ0�!�u�V���F���S�����fy����Lu)�-�<"���'ޗ�y2Z�0�I˟������Iן��O�d�HI24L�h_@�T�E`��ـ��O
���O2���$�ۦ�]�?蠁q�[�:L�pC��<X[���M�D�|J~*W	��M{�'|b���g�
�`p@�*.���'{�����Pɟ�Bp�|�P���	˟T:1ʍ�|��I�����n�Q����(�I�X�Iaybhv�:��t@�O ���O4��B.T�Odp���O�&0m:��v-"�	��$æ�p�4��'��2Ȗw�q�r��$.6�"�O����=Rcnmr�,8�	ν�?Y��O"�᥋��6�
d�=.o@�ҥ�O����O��D�O�}���P����3F�(uj�aQ-4�i���M<N��'��7�!�i�{���#YE�t�e�Ӌ)�`<�������劣�ڴ9��d��4����m0�x��'*d�p��Ǚ�.����V3�#�e&�Ķ<ͧ�?Q���?����?q�r�Խ����G�)r��[��
ݟ81���<A���䧙?��F�]s��H�ee�ir���Iןl�)��S�",��!U.T�@G���p��8l�0u�B��9R���p�aBfe�OʱAH>I.Oę
p�ɮ[r�Y��ɉ]zPD��O����O����O�<QѶiD@�y�'.<���@�D��y��c�0G��I��'�$6�4��$����Φ��޴���J��%I��G�u*�i���Sd�黑�iQ��0�N��Oq�\�N͕l*YB\�ޚ�rc�֞3���O����O>�$�Oz�d?��{�(�3�E�D�b���4>Uvl�I����	��MS�$��|��&��֜|��4P0�@�Dc�JQ��.f�O����O�i��K6�(?ic��"وH�U�#S(�}�A�K	s�胲m�O�8:M>�*O�i�O��$�O0(����u؊�q��O74��d�O.�$�<QV�iS��CE�'��'�哃iN1�,J�Bs:�J�(ېh�F�F���蟸�	����|��V�R���x&�-��^.em��j�;�qc��a~��Or(��0C]�'�8A�tfG*4�ҤZ$�J\�z��'Ar�'IR���On�I �M#d��p�n00������b�6B�t��?I��i]�O@p�'$�헍$�ղ�a�m�ta��1a{�Nx�z8�ce���t��YP�n䟮�Ob,�@�V�h![SCڊG��mX�'��	͟���џ��I럤�Ih�ԅ (��L��2<�X����
Y\7G�Vۄ���O�d+��	�M�;-If����[�U:��@�*��	��ұ�i�Z6mN�)�8Qh>(oZ�<YSe
8܈q���Z떝h���<��C��M���	�䓛�4���'8���'���]⢆I�����O���O��J��vi�n���'Z�G�9fCҐ���-^�8(�+ϵAw�O$��'�6�禙�H<���U�3�4`zs�++��X���G~��̩V�n���#�>i��O�f��I=i�"�T	5�Ys�N�C��h��̘\��'��'�R����khػf�|,H�ϓ��2�,����:ܴ9͢�a���?Q��i��O�n�|���Z��Õea\��l�0sj�dB����4V��o�12A����� �(c��d�ڢ`�����	(5ք��V%��'���'���'�r�';R�'��I"�ɇ�Z�1����_��	�M[`���?I���?�J~B�3����#��=��pa`�W#;@��z�^���4$�Fg(��Iݱe� ��X�ߓ[V~e��7[n�͢GiN2�b�K�|�Qv��O���O>q.O]��	j��ܰ�ݍV:]`���O6�D�O��d�O�ɥ<�Էi{(i��'��%S�ȓ���0Cj��
�2�1��'�7m#�I ���X����شG��f�2C|���.�|�g(K�3+����iu�	�,U�S�OOp�&?�����FX�S-�'yޮX�'ǀ�A+�����	�	�0�	l��e��()@�5��H�uۨ����'��'s6�͈O����O0�l�]��.:dX���--��p�!J����&����֟�Ӣ{��Dl`~Zw
X�(�PD��!Y��[�'
���1���<a���?���?���+�t�P$G��p�T[���0�?i�������aJSCA��	��0�O��a�=G�Z��)	�s꜅j�O���'���'}ɧ�i[�OG�}X"��5�����'S�>����wĀ�Q�7�my�O�����
�=�c�#a��Kف}���y���?����?��Ş������������]�HL�x�N���m�IџD+ܴ��'�"��?�+�'y�a@Oĸ<��� ���?i� T��޴����@a8�?q�'���i�&�n�(���ox�'j�	���I���	�����P�d�դ`Z��E�c����CK&%*�7-A^����Op�D,���O08mz�y�a,"2N 	��K�]��i���ן ��R�)�Ӽ=�T�lZ�<!.��)�l�
��ɞ>�ԙ��M��<��
۩����n�Cy��'���3����*��׌)�"�'��'���M���I�?����?��&�i|t(5��9HM��������'�x��?)����5��MA��&����*Yǎ=�'Op���B�R`�&D$��Ć�~��'z�1��K�'�x�bE��39�����'+��'d��'H�>��ɪ/m:E��aؕ*�x+��
�2��	��M{�����?��AK���4��ꡆ�.���`+T�m��6�O"�l�R�l�:8��n�i~���lr
%�S
5�:�P��1+�^U�$�c�B�;�|"T�����h�	՟��I�x��@U�A7lp*��`�6��Lyr�`��Z�d�<	����'�?I�O.7
aJ@-��|	�]p��I"�M�T�i)�O1���JD��N��D1C3s�hb���XV�@D���фoQ#$U�cy�i�4���	�� 
�3�W���'���'�O��I��M�#b��?�PD٠7��;e�
9F���scӎ�?Qҽi��O�$�'R�6Kͦ}8ڴƥ��1�d�PA�#k҆����C5/��5l�s~B*�^���x�'ǿv&Y'ld�I$�4���ࢍO�<���?����?��?I��$	EYꢌ:S%�`��y�
&:���'Y�v�\-�V7����OϦM'��X�<7$c�$�$#�U�'���ēiD�V`�� �=R"6�8?ٱ��,YDxP�+R�}&�x��$��!��O
��O>*O�i�O����O��jL�B|J�3�O tc8��dd�O��$�<�V�i� �'��'�哲c4�u�P��
�q��k�O�h�H�	��MST�i.O��,{�D}x@.B4|��W���Ѳ'hT�3*�I#��9?�'ofD��3��)��#C�_�4q�ӏ�0ZK� ��?����?��S�'���C��tn#���2v��/�\�A�䔖/��!J�6�d�W}��kӶ�D٪)L]zꊲX����B`�S�4-��P��4��Ę�Y:�'��S4�9���		�P�a����+D��	cy��'�B�'�R�'{2^>]��@N� jte�d/ΈB(�8!!��&�M/1Lv��ɟ��u�s��������ɔjd>aIw/S�!�v�(5���{��F�l���'�b>I��MŦ��H�Dذ�m��?�ȄGG܌hK�ϓX�>̂���O�̀N>�*O��O:-�q��#~H���.^��x��+�O���O��ĩ<���i�]y�'L�'�
��ת�l2�#'��ha��D�U}��r�dnZ&��jF�թ�i����e�ZF$����������}��Kc�3��!}��S���P�U���A�.S)jv�����۟@��՟ �I˟xE���''`�H�&��*7@�1��l}f����'$�6m9%#���M��w��U���WZXc0Ϥ4D�!P�'�J6��˦!�۴ܞ� �4���I�chҠ�'H43׊�%"tjs�M�:T����$���<�'�?q���?y��?A�%]%l<b�S����Hf�-q��O�����ئ��wJI����	���&?��I�*E�(��
]�&)f�:� E�p@�O*=m���M���x��D#[1 d����*<@�0c�R�{t�����
�;Ƙ����#���O�˓4�riA2lݟt�(l�A$�{Юx���?���?I��|"+O�8lZ0'����@�"���2��x��9Zޚ�����Mk�2.�>!״il7���3g�W�`l�{�^' �D	��"�$zZ�o�^~r ��L�����E�'���cD9K'�!hQ"ۻ]��{Dā�<����?)���?!���?���d����T0��$(^���ֳlr�'2¦|��H��?] �4���|�,��+�@�
2���K���'�"������X�v��h���-^kFe���˸V��[��!>�\���'\��'�������'���'�|D�2�,
N�1/[�XԘ	It�'t�R�`2ܴo��h�+O���|b�?3A,��hP�b|2 �
d~��<��Ms3�|*�� �q�f�M�#zzAb��2V�����6�Zو&`$*��i>ݒ��'@��'���SA�-�r�02Y�?�.��J�����@��ǟb>ɗ'ox6� 
_����$��ŢpB($�x��)�O����Ħ��?�rP�p�ݴ|�"�d��Mᎁ��	��|l"��i�h6M+(�V7�7?�DCڎA��� �T���&	%�'@6^��lW+�y�^���I����I�$��Ɵ`�O���@߬s~���":,���Kb�6���O����O擟��d���]0l�b��uh�#��`H3
E)\/����4����(��Ѿ^:6�b�l P̻k�^H�A�	�@�x�xSGw���v�œ����X�	Sy"�'[�']�I���!�x���#2��'�2�'��I��MC����?��?�W�ZX���.�	%�\������'q>ʓ�?�4!�'�f�kP��5yׄi��F�0
`!��O�	sW×�\If��󉔪�?A�Z�j��Z)8`��É�m8�����	-�2�'|r�'^����аo�6�L���	n�(y���H<9�4#��=����?a�iH�O�.�U���BrÊ*t��9 ���^�$��Cݴu��E�
k����c@�K-���W�iq�A��)�P �TJ�_��$�,�����'���'!"�'Ť|�c�	|�/9�r�mT��ݦ����Ɵt�I̟H$?q�I/.�ɇ@2T&|h#��:�6PR/O4��mӴ�%���R�b��6MYr��S��"
��v��/P�asD�� �s� �]���N�Gy�F�8���ƃ4�.��*��0>�Եiݴ�q��'��y���A[qX���"�>�y�W�'~66�.�ɕ��d�O�7������l��2j\�Oؚp��;�`(S���mq~���E*��ӛ_�O07�Q )h�vK�#a�� ���1�y��'�l���F<�]!�o��U�'���'�7-G"=����M�M>��Y�*2ٻU�""ը1H���.~��'Į7-E���0b)lZQ~�O�1x�*�r �:��̛P�Ny<T�.R蟔#`�|b^�\�?!(ƏR^MB���!�����f�'lf6��>X>��$�O����|��A�1��j���"Z�֜z憚X~Bj�>y�i\6-b�)��i�"Y\\h
*D�X �a*�cBH��(R��ָ�H��/O�	Z"�?	A6���_�~���-��<N��͜�[����Oh��O���<�B�i��؂���$L�����1^�L1BbMH�h���'�27�?������
Ц�xg��A�x�(�"��a)�}���Ǩ�M�i�x���i�	@�zq5�O&�M�'���A�߳|�ɔi)t))+�B:�mK!�� t�9V���d�J��e�ڹ
&@��Κu��)�V��,�#ڔ*��J���P������)I$��I�i��H_D$�t�ޭF�$(���=ғ:��L��*zN�IJ֍E.m���"Ӌ�uܸ�B'���n�pT���!(��H�� nf���W�B q��mbR��5]DmX�>n��k=Qɔ�0�ك�F���`��asT�����48>pA�h3M��Qp���	[-ޘ��@/q��hT��?:��[6� Eڮ�nZ�$��۟|�Ӈ����<�b
>IΈ�X��>����-	���� ��O"�?��I+g;�� ��V�<!��ED�f�<�ݴ�?����?�Q�C��Iuy��'���,<�F(pc��Nh��w�ٴ/ѱO�(�i+���O���O�4��½X����V`��2A0��a�ԦU�I�[�,i�Ot��?AK>�1V�̨H��Y�k��S珐6G�Vi�'�i՗|b�'4��'��~8��!���u��E;���o0Lp�X�����<�����?��8'|,��nW2�:�Ӓ#�(z04(:�dж���?����?)+OX�����|¥���h���U 2<�`� Ԧ!�',ғ|��'-rCޏI�dKq����!� &3(�p�!E�WD�I����ޟ��'i�q��h�~R��q���Q�J	�R�G�<P��"�ik�|R�'j�i��RqO4Ԡ����<�!1��+p9��G�iQ�'%��&)Chp⨟B�$�O���ʇg�����*&�8k󧄆��D'�@�	ɟL����d'� ��y{�< eJԇY��W�P�D�r�n�Yybj�.B[<7��O��d�O��iRg}Zc��52KF ���I{����4�?��>c8}���)Ǳ/�1�!dߝ?\�pѷ��i�vc٢F��6�O����O���P}�_��适�M9D�ŢKt��,A!X��MsW���'G����&6�\)b0�G	j��1$[8Ye@hl�䟰�	�������$�<���~�]>.բ	��Ӌ�i���8��'qr`i`�|��'8b�'����
:����_q_���3,q�����4��?�4����&�$���ҙ4G�qЖ�@�ϹV�|�'����ԟL�'���'O"U�d��@vE�soʣM�̽�G [�����-���O���?��<ID�D���eQ�*��$�V���������$�O����O"�4%�+w;���;�JO��@%�˗����	^���ϟ��p��Oy�$:;��bU p+\퉵��v�R���u$&OX�d�<Q��Y$���+�|����-�@h�1#�4�ʽ2��)*��nZX��?+O4@�őx�1��e�S΃^�Q�ĉ���M������O�-����|����?���K��۶[�*�b��Q8Ha�&&�$�OJ˓$�DxZw�f��Ђ��o@ X�4�S�D� �4����0W/ܕnZ��i�O.�ɀi~
� �I���Ȣ!�&���; C~!cD�i���蟰��)�ħ���ݲ�]4m�N����-g�=#t�tӘ��
�E��ٟ��	�?�:M<�'>�H:�F�:	�y˶$^��H����iD��'�"�|ʟ��O2����^sو�.��q�\*�Üݦ��I�L�I�cH|8�K<ͧ�?i�'����qU�l�l���-ЛX_ȹ��4�?H>]?�?��'���D�ZQβu��@�`h:���4�?	�6��e��D��-�hX'%����a�sٯt��%�8g3?���?1����D�SB�C%������ �,�uY�!Y��ޟ0��򟘔'z�؟�X�7o��W����a��$:���1Ƶi�BX���	��T�'8��ד8��)����Y��+���t$EG���'�r���O,ʓ:��4mE+H�R�))%� �V�� K�O��d�<Q�Q�D-�.���d�:jd�R�F.rW�0��*ŀ%_�Am�|��?�/Of��x�=]���7E�=�������M����?!*O:���CC�̟��s��3"�\� ��Ff�v
�u�&c�Bʓ�?Y��?a�����<��:��us�(��5�ؠ!I۶P��lZ{y2�L�Iu�7C@�4�'��i;?q�$~}Ad�X�R�S�����'�r�'�����g�s�6�����/��4䠁)�MkqK��F8���'�r�'��Tf'�4�:��R>@�Fѱ,bx�9@l��M����Io�)��?����;m;���ޕU��Q��֤G����'��'p���tg�>�(O"����|:��L77k� �+��$��샷�>Q+O�49������P�	���;�W���dW�D�!�8�M��Y"���Z���'��\���i�u��c�@����q�N�3 b���o�z��<��O|�D�O`�d�ORʓi����3+��e�꼺��\�m|$uJ(D�E���_y��'��ߟh�I��憕& $�2/΂���q���ͪ�ICy2�'OR�'剤-8r�Ot�y� <v֨��O^�?��3�4��d�O�ʓ�?���?���<�¡�'_ը��E�49�4�$��'����'���'��T�$0� ����OzU�0�/Go攑���G�dA��(����	Xy2�' r�'g��c�'��C������T"�P��ߗx�tnܟ\�	dy�n6W�b�'�?����"�Ph��񵪝�����$ɰcp�����I���ADkh���	NyBܟ$e ��ؑ=��̃��
�R��ði�I�]��ݴ�?I��?I�'J��i�Q��l���,�KvM��"�Ψ�IzӐ�d�OJ���	uܧ�R}a���]Wh�ic���,|m� TW:U�޴�?!���?���6���Sy"�K�&�P�R�h×h��\c
�#�P7�؏=e�D3�2��,BQfǸ1�lk#��C�f�e���M���?y��I:1Y��i�R�'E"�'�Zw�����D:xsZCra�(e�f���4�?Y/O�7�g���?���?i%eW�~<����(�e<꽂aB�����'Vz}�7�>9(On��<1��#�87��I��Ν <��Mҡ��r} ӭ�y2_�D�	ƟT��|y���c&���fv �:�G:N�ʡ0�>A(O��D�<I���?��[v�1i����X����Ѓ1�ָP',��<�-O��D�Ol�����B@�|���\�,dB��6��7�㤠립�'a�Q���	ȟ��	�+
:�d%���&�48(H�
h�+G
`nҟ �	��	Ay͜�L|�'�?��5�H(C�	f*��B�;>�l�|�'��'�*Ͷ�y�Q>1�p�6%��;Ra�<l�B��aL�<�M{��?�/OD\Hg
FR���'���OȔ�:� ��7� �� ����E�>	��?	�9���Γ��9O��5>��-z�ݴ}P�x�@ݖB�6�<�G����f�'��'
�t@�>��@��%�$g�!J�4����!�6�l�����ɘx��Ig�^�''-��Y��
$A{����X�aj�l%"�����4�?i��?��'.��Iqy�'��-d��A�� �m��t� ��M	J7M�7*��Oʓ��O�$�R�r����A�cټ���
	v6��OT���O ��"�N�	�����y?!qAS�D�.�r�N� I�Ck�Ǧu&�(s�Ø�ħ�?A��?��MQ8P$+2���kݩ%̍�5�f�'mV���#�d�O��'���&�"�N$e���(�O��-i�^��顢ɟ,�'a��'�P���#��ucx�ҕ#[q���`$�!9DD���xr�'�r�|b�'��ѱbT�0B�aZh�Ef-!�xZV�|�'2�'�	�m���#�O��)��G�@:b����bI<����䓓?���rj��'�f�uBȚ0�&a��DT�����O��D�O����<�I�$t�OiDm�Co�uꉑV�H��mCd�s�*��#���O(�DY��5}BdIh��jd���1�J�	���
�M��?�(O�p#���t�Sڟ<�Sh~ |x#$2>��ĥ�0	�<H<����?I�)�<qN>q�O� Z��Ű|�vaذ��ABxYش��ę�/]�l����I�O��I�J~b��?>
Q�Gڋ5bH�;pƟ:�M+���?�JS�?qO>q��T�}{�	��X73TVa�Ga���M���"dB��'Y��'��#(�ɲ}Zޡ��"������D�v���:޴�6@z���䓔�O�bc�X���@�i�>v4��h�>G_7��O6���O`�s��b쓨?�� Z�k�#P�&���T��1/���C��iK�'��s���	�O��D�O��x�%�V�f}���2�2u�t*��u�� �`�iM<���?!K>�1 �M��K͖v4(ʱi1~���'�ȑ���'A�����̟ �'̽P��2w���:"�� P�t� �.͞5fc�8��@����<�	xd>�"�-2'#�����E�S��-�����$�'�R�'��O}���6�~>���'��p��u�c� �($�>Y��?9L>Q���?�
�.�?���ԋ'��u%�1U��/X�]�I�0��Ꟁ�':<�2&$0��ŉ2h�9�aΝ<al�e+GO�QmZ���'�,�	��B��c���Ol���!��ڵ���<���i�2�'��	�95�miK|����S�#$���)Epa�u�� �h.�'�R�'��ِ��'��'��i�u,BȰ +D�6SxAլ��i&���'B��H�2�'�B1O�d�'�Zc���"4�D�K�5�'܍R=�Y�۴�?���3,@xB�EA�S�L\���& ����TjR�~���m��
T���4�?����?���g���d�$�T�o�p������0
C��Ax 7�F,
����Sx�Iܟ4�q��9!w$�����/fu��g�3�M3���� �r�'$�	֟8��~䠥�� � ����U�����DZ�S�T&>u�I��I�T��q���3C��:�A�D�*Ձ۴�y2A��?���8p����&��q$�A 2�l�	U7�)I�դ��$�]&UA֒��������RyiݯC5�m�C68%�ܺ0)�6q�p%3�ϼ>����?���?�r�gx4�@`��.l4��텝�F��s�|��'���'��'�t��ޟ:�a�D�aZр�� =�`(���i4��'{��|��'z�������4B�� ADIHG��D��ɵDE���'r�'|"�'f"�I_��'gBȩ��$�o�+�hYI�٤n!�7-�OO@��O��Х��Tv�'$x����!��EҤ!^�Q
R�`ݴ�?y����J� ��'>����?9�7n�)������N�9�bƇ�M��o�$��8��i�h3(�0?&���iņ6��!ߴ�?��B�ج(���?���y�����L1x���<h���0.X��\��Ĳi��'V&�G����Oni`���<'&�pۘj�ƴ�4Y��qr�i"�'���O�hOX�d�t���V�"�&�ǮW��@m�2x"<E���'�f�#v#(VgЉ	E�^(_f~p��f����O���,�r��>y��~��n���c��*ϔPa����'[(��y"�'��'�� �D�]%�ĉ�o�)#�)�b����U�z��$���	�P$��X'4aH-9v�ȌshT��6��:
�zq���<	���?����$�)j��٥��6�=��b��cYɓ�F]��?�M>����?�E&�%R̮aɠ��&j�[�b)nݒ��<Y��?����dH�_�hxϧV��ƭY�6j��K�l�	~G~]�'���'�'���'G<���OtmA��W7[��A�J�k����Q���I۟��	Oy�t߮��q�#��!	TG*�2T`Vēbg ���IF�����AX�c�Xk�V0t�����Hs�����xӺ�$�O� Ĥ�Ks����'�����8�Ġ�A�Iz�#Ʈ�z��O����O�EQU�~�A=
��p,����rOЦe�'ъ���K`Ӏ�O���OE�4�����a������(i�<nZ�����#<���Ď�� ۼ����.R;y�R�Џ�M�!��7x�&�'���'��o/�ɷ �i;�'˥^�v3F�+�9�ߴP�րDx����O� s�ϐw�}�g�==lY�K����I������"�tɨO<����?�'��=�e���+����%r�}��6Θ'�b�'��xa����5��Y9p�Ķ-f�7��O��B�f�<a�^?��	j�	��T���ؐ0����%ɉu"��O��ؘ'K��'��V�4�TIW V�P$+S�
@x�-2� Y�v%{M<q��?I����<iE-�,1�e"��'�B��g�	�aH2��<	���?������# iV,ͧ7V�k��M:
0թT��#j��'h��'-BS������%�~Z�g�v2 ��� �/,f����J}��'32�'g�	�d�@ꭟ��D����I���+TT�Ւ���9g#vn��|�'-��'�B�_6�y�R>7m��~�~}�C�Ԇxˈ�(B��3Dt�v�'(_�d	RhM��	�O��$���=���H�J#H�~��r��V}2�'K��'%(�'��s�L����"����C�VD9 嗮)2J�n�Wy��L�)r7��O����O����n}Zw~2-�t�] S��%�)�Z{JA��4�?��j��̓�?A.O��>͘u��+��S�E�X銆nyӺ��QB��1��쟤�I�?�y�Or�f]���'��O�����?!��B��i<L[�'��'��b���v!HUF\�q9��	_dQ�!�|���D�O���!E:t��'��ퟤ�{���e��T���`�)it=o��|�' ��R�����O��D�O���Rh�1�����L;���Y�N��	�n�	��O�ʓ�?�(O���ƄP�����! ��;�$R�Z��@�g���	ʟ<�I؟��IMy�S�u�\��Ő�7��U��Ř�"�l�Qǎ�>),O���<!��?��l?� B�ZEkE�A��Y��9x��cCU�<!��?I��?�����C=Q��̧6Ai��b_�rб	�(�."��(m�by��'�����	��U`x��ػm�R@R9%�r���0���?1��?�.Or���Q�t�'��a0-�! �"��©G�o��,��Ak�d���<	��?���
 ���?��'Qv%H��g;�h��h�*p`\ij�☜y-�9��>7�>)5�.�P9���	R� ��L�O�<@˜�(�xT��S��|�$�� ��1)���
B�H5�O�T!*|�������T�[�B�����!Ũ�������/u"@"�#��oY��hV��^� (��K?LI�HYU�V�P�XK%��5AJ��cT&��Cթ���J�p����D�&�֠�奌�w��8QS��*)���a��y&8�(�mA��@��nԌ�?���?��+���)*Ӿp��V�Z-�6倨(�R@'� �e���8b>�O`���@������8d�p� �
iB�Ha� �A�* q��'ޞ�0X�5�*y�wY={����'���'�ѳW�������OV�#p��2JuA�Cұp�8`���74��	E���w�PU��� ����!v%#?Q��)�/O��7�4"��s�G�15�͑d��8�(��&b�O��$�O����ԺS���?I�O�<L��"ё9 ��n��Ht���;CΝ�����d��'Mp#n��c�D����~�^�(��]��z�Ae�E6K�=�d�'�|��(�K>��UbF�J�`d��8�?)���hO㟄������C�"dU�t�t�LB�ɀG�\	#ĂExX���EA�~+�c�lx�4�?�(O�!2��c���'nIS�!!<��4�ݝO��� 7�'U��H�b�'#��:'XDو�i�i�>A!�d}Ӑ�SC`K�a��� t��>�����'-XA+���-u� SԪJ7���OҨ<Lx8K�mH�sk��b���Ɏf	����O�L�! �ߦ;k&�
f�K?�\�<9ߓ3��dSѣHFH,҇��@�^��L@�FA@�<���m�5$a��ȏ�'�[����aգ�M����?a/�R����O:��5-S�Pw@d���'|�&(�b��O����<�4q���9�ˮO�D���B�KÂÂ'+/@"���i���a2HD`+^1)Q�T�O�.� �GM�^��e��3Ps��H��� ��O�b��?QS�C�$��q�dᑪT�-�4 =D�[��^j�������:���CM-O��Dz�j!38�4F�w
6�a^�O�T7-�Od���O�2�Ѫ9<p�$�O��$�O���y�,��E��a9bQ��p�!�6�3lp�$k�%�$-�0a4-7�3���^��$���k"��S��)O� �$�e����U�������|��8i��A�?�L�pE�K>	�1OB�p���Ϙ'��d�Tl�	�Ҝi��٧f�v<���hd�NU c�A�wT+<��1�'9�"=E����^#*�e)ԙ#[�A��f��C�P3W`�"Q���'42�'%(���P�	�|�P�R�3U�x@�FdLdzV��,�DxAĬ2fa}�����J�jc��]������,2��Ka��4 3X���^�i���A�,!C|�ӱ�@C�����'�Z7mϦ9�Iy��')�O�9�ʉ�~��H����fQ4��"O�e:v/T�!P*T�*G/i:��ڇ�ĝP}2T���l[��M����?�A��Fq����	��f��aݖ�?���9�i��?	�O6P��!��!�&����fp��aG�P�!q�G0
,L�O^O8�\`DB	�)��Qe�%O����� h��Q�̋&>~��)�� <0�x2�T2�?�N>���?���E�$��s�.OD�<��#I@���G����Hxp�[B<A3�i���(��,�J�(�ʨe^��x�y��fZ�7��O��d�|r!ك�?���RcT���7��
� ���A���?1�w�����̠X[����d3*�"�'\$��Z��8����3v���O��ɴ%� (Fn�:r�J?n%�#}b��/6VA�G�4I
ڽ��#\[��1h��'��O��O=@���M'E`�����'e��*�yb�'{�y�������2a�c��P� F�
�0<10�	�4��P����|��΀ |�pY��4�?I���?�1�S98�����?1��?�;��58��Z5����� K�L���3�hei�'�� �W������q�BɰQ�mt���#gb�!h�)П+Kl���'\p�S%�J�g�Q�X JM�� �d��Gϫ� -�<��G���>�O|��&�0n�!q�G��k��(7"O�8#0H&X�P�ɿht�	 ��\Z���ӕ@(>|�Wj�AGٰ�G�;x�C�	�:���8Ī�2Bհ��G���C�I��MHbM�m��-�5���{��C�I")?48��X�3]~�R���͜C�)� Dd��&A�Ťm�iF�J%j�I�"O�cdmЯRP����ǟ�:��Y�"On�[�F�F���I�mж�J�� "O������c,����<d����5"O�tbŕ8��ha�לf���(#"O��0�J�BLҥӦ��u���i�"O
�B�خ5� ����x��"O�9yUO�6E����
�T�<y�"O�2TNƚj���)�U$p��L�F"ON�3��](5\L�s�i�9nu��"ODE�f�e&�)"H�>��X�"O�;�&��f��UpP���.|RQ"O֡��A�!��l!����3"OB��ADک5ֆa#�Z>Xp�"O�q3rM��3�(�R�2j�!&"O��XN.fTH�Tf�bV|M�"O�5�TɊ�w�ԼA�O]�7�=:�"O��EIO��H�F虰`P�J�"O��oV��zì�:5� �g���y�(Ϭ}Ͱ%r�@�)Q���y �/~.x8��˯�>��2�y��D9K���4@8���VMć�yª����%��K�0þi�uD�3�y�l��7��uy�瓐%� ����л�yɔ�]���G�. Dxe���y��E�U��� �L�������̸�y�k�E��h�H^,� �6僅�yƃ
 ��)�e�z/Z����ĩ�ya�<b���% �\��ѩͣ�y�	DlN�'��q�
��Fϣ�yEĽ'�dȘ�oM�YT��G�y��B	@5�m��`�Mo�A��U�0=�O��3ϰ�9E��`��K�F�e�N�E"�2scR8�y�nV��PP��Q�O:�s���'G*�Y�s�v���$�'KA�| !*d�x����L����s�d�����LP���L"�pGJ�"vNp�Z�@��!&�g~"o�<d�pXxu�J�w�]�B�Ѕ�yr��7m����K�G !�����]�v�X,{d��:� 1lO��qV-̙?U�ӗ��rx@��'o�ɋ�@;, ��o�J̛��ݾ}�x EF �j�j&"O���kQ�ꈠuEۭt�F�z3�Dگp�V�:��>%���E��`[�\�𭳗 Ӂ#ux�ۑ�ؔ�y�'��-v��m��0�\�$s���=���5��E��O���$m�($� /��6%&�+D"O�Al��U�!; ��% <-�+�
̆I����|}��	%�=��	ݎAH����ݿO����d�"���
T�ޥ|w8�lZ�CI�x+M�I�(-+���22�C��jӶ=���ȃU���Y
3@�c��XX7H���m�!�H����d/Ǚf��UR�gX7!�r�� "O���J�sfڥA��,>�b�)��,+C�dx�\X}�kL3���IG��ʆbǩ!����A�-#C�ɻ������W
2D '��r�P�;�/.Z�n��p B��=9`�.	׸��� ?TP\��^[���0�(,��T�����M�T�E醡��a��Bt��s�]N�<�l��h$␻��]�9r��J�Y�4y򅅈
��Y��R>�SB�D�{*�Yk���e�p81F��C�<y�bV�Ph��*��x�C�'� 8b,�'9~�s@9���I+;���P�,D�p���oX �B�[�W��l�G�	5m�����(�g?����s�D1I�,��7
p7-\"�yljV�h��@�Z��e�!���?��E�$�p��@DX�ԋ�1U�f�#�ߌ��d��;:�qp�O�t�P`�G���Fj@ -��"OK�*p~����1[~}Qԍ����'��1ذ�B����� �!:�Uvq�a#c�3*z�{V"O:�I!���zgZ5�Gҙdg@usE����:I�y��(�7&�-c�$5�N3t0��X�-D����E���^x@�K��NL��ԃ�O)� ���|R��t�����
QXza#��	���=Q�4V��0���AZ4(�St�b"�����ćȓgz:���@!%V����D_&�%�?�c˅�@��TD����&�Zd��/�H�r�0�B;��'Nu(��2�'t/��٣�J�_J=J@g�l�R�wBș92�b��E��'���"�])p�,y���Rr4�#v(Ь)J1O4�a� !�'�yG�1,��4�E|��!a�`ء�?1���NJ��	�$L����L�)׸i����k+�K�,��D$i%��)��L��DRL��}�'��0ۖ�3߈uB��6L�1)
�`�j�(C��l�P�6vܘH�2'�(�#v�¥IU�iaÅ�$a ��dٝgd��	��I3g�P�(D3_��O�(fkа�y(��X��M�6*A�&>�IƁJx�����'���%�;x��ĉ6"��R)_K[MY��$4�Hc�J`����M��E�z�	�˙��OA�n?]Y�����Q�L�<pBF�()!�D71��}Y���1&�:�bwN��Dpwe̵1G
9�6g�]B��O��]w� �ɦ,|�ू��	ވ��CK�>����*[6����'�|qڥ���.������S~� !
��xi��)Q��Y��I�pt���^�|�m��&.[2��$��KG�;�ϝ~���R]6d�+��eO����(�@ �ԩCN�G}r��T���|�2&� �,��f�c��r�'E�-k",��>O�H2"�	7�RE�6.� ��O����?��]AC-R�R��W�:E"�
�'_�p�c�B�S�O�>�Y��|]B���	mh�Y��䃾Q*�S-e��҂����a��xU�O��A��i4�d*cM��20L���'�x���#H�6��i��4�`�#jݲ]�ؐQ6C^_|�]�F�vx6�ɡ9%�����/�a�T�=���	eb��N�.=�������x�d�[D�ӄ�Z1	���\)f�����ˁ'lq�������I��ʧz�xx��L$&	��A��?xK���?��oH��Ѱ�G�����qE
G��pnH<dx��k�f�\��U��(�����<���Z���i)��@���E�D��b�o�ld�bI`w<<\'�`��h����
V���UlȓQ���t�S����b�A̱E�=�m\��:��TW?#=Q�bد�~a�'D-zjf����ܺ�4tuR��'fWL�';b�ր�UCn 31��G���vT��N0�ӁS��Px`"�|�'��x���
����f抴 6�R0�ߕy�ԙ��`��ok��|YwM�(PB(����jL�P�\>��.^$SJ0$т&Q�/�$��M'}"L�W�I�`��:�����JD�OXt���/�U*9B��N?ޱRٴW�����Z�tЫ����?7mG!f!���`�ds� ψ/�$sD$��&��qVD8��L>���Q�/��tz $HL}���`p�y��	 $PH@Q'�'G���Qѭ��^�1q����j���8���֙���b�M��.��@� �OI��1!��w�X��	�XG,	��O��pVe�,δ�1��Ƃp���+��i0�L���d�'�̙�fkѯ��O_Ԉ��Ѡ��5��;i<[K<ɑjWs��D@�| -ʉ��#=�:���V'x���(�-�u^���`����ـxh��z�"~nZ��p
4Ⴘ,5�4 �L�ܒ�I��E�1��DN
�D&� .h���7	�j�C��'��	��O��|�t��~Fz�G�7��[ElS� �FљD�C���ɤx	x���	�D:E
�O�w� �M��t֔�,��C�Z`��ɟ!`[�y��I	H"�s���
O��\Iv�R�L����ʝ?������m��>Ʈ%��	��٥�t�I�㛼.~���ѬZ%lW��(���� 3��bᓵ�j�-ƼV�v��G�J�2�f7�N�^��Ě���z(QUn�+�����5�C�+��ب�"W�C�<���?8��F��&b�z,O��}��Ji�����6LhݫRGb����q "aӄ ּ(q,��ϓ2Zr��8�6�Sæ$���@�i�v6mͦ@�Jaڐ�A�3�Dz�H�)&vт_cʬ,���8V|�Y���4��]"��ڂ���ޚ��O�ư�G�Oe��B���?�m�������7�(��A�G_�'��uȲ�V�\��᛻(�z����?-����N�c�/6��7j̒a���F{Bq�d�и;#���L��6�D�E1�� �B�T���%�Mç��F7�BV�Σjrݡ��}�'�����YgnȲ�hNm�8;�4�~r�.?�Vq���sC����6g�O���6cE��mχd.��
#�?/�V��'�џ�H��-k3򁘢`��tY|�����''���9лi�m1�&��R�pF}��u�z���9�I 3�+%R�Ч�p�"?ٶH���'�H�J/:��%i�֚\M��l�a�'�$���zG�5Uc]�f��Ap�O� qST�A�HYB4�2'J��Y�,����I��Oz�C��)�8�TB���+��92�	��ԧ4�d@��լ�Mc6O!�2����S�L(���1&oyR��V�~�����*�8{��Y��C :��˓$"|�0��G>l�h١ѦO??h�H�ҩ��,HҠ̔���c�ЧD������<���\�oɺ�x%/���(\�wL w<d ��ٷ"�B8hƆڕ<G�r�K6�hM�#�i�d��/B���Qu��`�.���#����x�x��v �|�7�*�1R8T �=
�M�*�V�=Y��c�i+�̓ ��C\�=��㯄�_�,d!�'pD��1+�0����Y���oߜ ��)%�GK�H=	DK̐Y�Xcw��]hd� ���D��<I0�ΰ`�Yas���e���syb+O&�J�{�ڇTE����i��D��ɣ0��)�C,;D%���3+��<��&]�[T��h ���' ʈ��8
��4�A̨F��x��`�\�������(��Ph���D-O�^�ADy2���6�LՄ�I69�����Mj��,�48�jd�W�9��y���ݞon��F�ƀU��,bÍ
v���d+X�T��DeߗN��r�FA�H���1���,=H��:��'�"�PV� 
?3�!�6� 3>ܩ{'B��*�X9�V I	a'j]�Bd�Y�'ӈM:�F�,)��pr�P�RB��E~��z�ڬ27��(O0@0(���I��a�h@pm|!GI�fF�\`�ub����\6���2j֕A���S�(�?�!�aKʏi#f��_�atT,���{��QOc���BO�2;�L�c�o8|O�mi��o����O�6bd��˶v�p�<i��4��˓�J8N+��97܎���O��ɗ	b8��qa��qm@!�VBј  aC<S�<��*���	0"���se�2�	����	P��2a�ʹ{�
�z����d\�"��(���3��A��O(J,�8���;'~�I��-�]��	#�ƒ�S2��1f���J�21���o����3	R0J��<Q���A٠� ʠ;&H�%^�@��%�Z�&@�'�E�r�z�A+WW7R�|��t'h�`n&D��jDcަBj*����۶/��,cЪы��l(�����M�''
��7��~�q`o���ηb�x��厓A��psm�uF!��ޗ"&v4h��(iap����G)5�$�@9O�ВV*	�|�V�["Hf*��)�p��>QTƚ�6q|Y�s��0�0��i������'����l��)N((gE[>K+��b�9<��������屰�ПX���C�ʚ��=Qw�[�1���b/��)���zuC
B~R�N
Q�zta��4Dj�}�7�Ŀ�?Q��FR�nh �k�u2���X�teq��48`��3n>D�p��6U�\�ɒ��.���ï7)A�`Q���lYl�Ѐ$�tt�Q�N~҄$�p|��ݲ�������|�zyz�ON��C�I�S���`�I�9���Nw��zo��ا���D��s��ɥǎ�Ll4�2�=1�!�G�w�䬩��t�EH��Jvy!�d]5X��� J�CT�I��"�5Ik!�[R�tD����f���)�.�B��"t&����ǟ�t?P�ا�Ώ�lB�	<n�~�h����@^,���*�u�4B��<=΁;&� 1T�8���B䉬K4���Q/'$ڝZVaB��B���B�|�ʙ���;-A"O֕`�V�v�n��+ֺ0�"O�i�@3[��墰K&0�t�"OJp8�����v�;�)އ\Kx�"O���Ћ4ֈr�VZ3X�;"O��� �
�H���FT%��q"O8\+�iЎ^|@�Pp��6 �ؼ��"O�L`�h�Y2�h�L+%�X���"O�}kK�  �9��O*I}8�C�"O�q��D0l4L)��H?;|�5�"O|�{eFl�Ȁs�T�*k����"O��:���B� ��[:�4�r�"O�ኵH��JۺeR��tb�*�y�K���@����%3��u!CN�+�yJ����9���}��hqҨ���yb���d���$��%�Lۑ��y�J�(B�H�д�X/T�
�f(��y�%�Td8��/\�{���:#��%�y�%�l�lAS�*ׂ	-�x�ρ��yD��4#�e�eo�2F(���X��y
� ����9:���g>{�(���"O����K�@��4S��W�e5�pB"O���&��n!J�#c���"O��!6N�
�*�K�@�$H$ �g"O2����q�,�8 �R9�:t��"O�\[���$v.�mX$O���b�"O乫Wg��q��yK�*K���å"OR�pd�� �� �s(IR"O���.�
�\���HO�~��s�"O`����|�R��B'¿i���"O�й �c=$��&]�8�s�"O��[K�-l������J3:��"O:�;¥Fjc&��D��'*�:�"Oܴ��M�`A訪��[��p"O��unS����G���6"O$ �j�: 7�Ձ#5H�F�"Ox�u�Œ9�,�H� �
�ts!�$��.�ł��-5$Bűg]�=K!�ә}�(��&�
��+�Ń9m�!�$$�>$�b� ]�ظ*7�FG�!�Ė@��H���&"�)��$�f�!���O벌�s� $�4x�Sd��!�Kq�CDӉ/�T)��6�!�D�G�(����N\h���&�!�&q7�p����;;Q	9pϿ �!��{��� ��xllL�G�\�8z!��K���ؔ�Eq�� )�N#3]!�_.�d�e�'��eȓĊ�]=!��ɛj����T��B����cێZQ!�D�>=���pnſ��Q �b�:xd!�Ĕ�G&lg��D��ໃ`D�OP!�$;Xi��2b�%1���`i¬0V!�dQ�
�<��oX�h`��;ӈ>u!�$I2��T� �$Q�͈ (]�eu!��֍{�pX��L-<F��B�	z�!���*K�P�.K�t���	�O��>�!�d���h��OR�Z��a�M��!��S��eP�")M��E�0 �!�D̀���q%��vNi�,�h!�E�y���9�!��i7�0f�NXa!�$�0Q���g�Ʈs ��%F[�f{!�D׏[zڬ��$�65������sc!�$^#z4��$�@��u��,(E!�_!�镋F�>��10��B��!�$^�k�r8�d�T�
�0�/3H�!�dBRf�%"�O�1{�L�2��8.q!�D��8���!DH�O�xP"n��,g!򄒣i�zđ0,Y��J4A.��7.!�$��6�2 ��? �`�ٗ_�HʱO�=%>	��І`R�|1W�Ҳ~tE .;D���&�DR��ps��  �lI��(8D��9�&��B�0d��<i\Bɐ��0D�@	���':��`��1�"I��d2D��q��T%�@��P�%����1D�@!�j��[�|̡s� rɾ����$D�,���ߏ`jdx�q%��~�~D�F"D�#c�!�2��/ӘE|�(�"D�����U9K��#⏐C�~ ���?D��C#��'�Q��#	�:Shh�h?D�T�B�՝T�ad+�^�J� D<D��8�
�6�7�S�D��=��-=D���n[?�B()�ASN��qL'D�؃"^5��*���"ӆ����"D���@�ʙ-��dZ���=l�j *� .D�� \V	�)Z#�XsR,޹A8��	t"O������
���pѫ֊����"OL�"P��9"6���x�$5"O��"6��l�4!y0�_<'�D�"O��Q���I��ЂG�p���Kr"Oz0*ԥR�TM�x��O�*4-Pf"O���×�,�<A���X�K�JzR"O
iѨک}lP�7F\?~g�!��"O�q�%3G���A�)H����d"O�5YaM�'�b� ��"�e��"Ot@�Rc^)B7�Q)6nܾv.x� q"O�l�!��-M�˧́$o?Xs�"O�b+��Xs,��+=r��""OԌ�0 ��vl� ��͈�-0pʁ"OjH{fC�
�$Ph�L�>�� �t"O*1�#%�1�vȋ6솯�u��"O�jfE��s��K��7E�Z��"O"��(C�G8:��� O�0�Y�"O�qP�
W�QI�՘�`W�R�E"O�H�@�%!v��A�Ƶ@��4�@"O�%h���Z� Gę>��D�$"O8���d��P���3�&�b"Oh��C�I�����$�P>���"O<��J�;����)S!/�̐u"O���ޯQ�`���5$�ٰ�"O��7Yi&q����c�r�"O.]A 푋z-X��i�&|:y��"OJe@����! JSf��`"O�ta�cȰv>�|b�� 3�1��"Ot�q���+g�eRr�O�{{n="OЕZ�J�?n�&�_{^�0�"O��`WN��4K�՚���jH*1 "O2�F��9�rb���!Cl��"O�87*M�b��e�%��i6֥�"OT�0� #���W�^�kU$�XP"Ot0ɣ×�3z6X���ٱH����"ORir���=5}nH�.S�lY�"O|s�n�!^=	�m�l.ū�
O�7�M�#��Ʃ�*+��� �@�<�!���"T��Y� ϭYנ��3�ڂT�!��Q<!���u�IҘ[�.G�Y��'dў�>�"7�1Z{.5z�*�&L�	B5�5D�8҆�M�w>>l����}T�@x��'6�ayҤ���85:���=��ʓ��yR,�<a�n��`E�=O������y���L�H��D�;-�0(��
�yҁ���fH����6&�J���C:�yb��X;b�au�4"�&(��-��y�Ɂ;UBh��ޘH�������y���o��=9`� m	~)�%OG3�yRED*Ǽ�Y�+iasd���y"�	&1�|p(F\xX���a��yB�ҸC��=xb��a�������yrǉ;�l����a�<�f��y2.ϱ��<Q���b ���[�y��;Y�Z,�+E(0l�
�y��+c&Q����yFe���E��yRÞ�s��`��j �I���I_��y�װD��y�2hN����3Qϙ�yRf	-Y��e�U$up
�Ѫ���y���4�$�XH3P�P<Ptz�'��H���}�UJ�lJ�Ds�Ј�'��Uq��Ґar�Y�,Q=kF��
�'{��%A��8]6�S��Z�9�n�y
��� l�C
�g�Hꕁ��r��X'"O8�#�J��5���Ɠqx"�"O�l�]7%�8ʲ�I9Tk�dQ�"O^��d{�mb��ߙa�b���"O-��※-�*�6��-4Ɩ��"Of�Hp(]�Fp�����)2�"O��K"lb�*w�E�eI��:V"O����� 4L�R��`F�e
�x��'r�-0��D���f��#�k�'�L0�%T�LU��{��ޖ^`�R�'x�iҳ�)Y fl���P9�ܣ�'���0��Q<�x��c�"�F$S�'b���)6(�Cd�M�3�
�ۥ�c�<q� ���Z�y�̏�:8��M^c�<a�!�t�|��F9�.��{؞L�=)�$O�3g*�G��$PeD���N�<q�/F�	(��'A����%JK�<��n��3���H%d��H)F�WO�<��D�pc��N<�vԨ`�O�<I2��]��-\�7~���-�L�<y7#ӫ
߄��'��=9��iq�DOQ�<A��ʉr��Xp �8p̀��M��t�'�Pѱ!��"1����A���s�����B،Sv�H�M'��#R-
O>Ԇ�A�̢�(�M��2'�*���ȓ6 �i�*(nE�#Y�^�D{��'�R�걃�l3��:1l�F��Is	�' jT��TOF��#%ո>��E��'��H�&A�,.꜃���'/�����'����w�ڣ������#�)��'Jq*"�	�%G�)��
1總��'�V S�IK+�|����[3x8T���'a�E#���wDd��ǰ�:� ��'۲��2#�806q"�'.�N8��'�. �cƆ/_�����(O6|��'l4	�4,6jր��A۵5r<Z�'���#^�Z��-R%�*�R�'J*�*WBؒ�Ɲ�W P�R)�4B�'8�m8��ה]�<lصśJ3��
�'¼����ХMXn�N6P��%
�'g�U���A�|պi����6y���B	�'��P�q��"���4ʈ u ��	�'
�*��<]�u�G���1�
�'=�I��ڶL�j������Lu*�'��1�D��5uP��Ã�{*�c�'3�a���h�ܱ��	>6�QP�'όԛ���c��4b�%�"4�X��'V|d��#̋j�n�7#�]�� �'����$�蔹
�ͅ[�
X��'�t� ���O�A�6,��S����'�>���h\� q����B�Kbp���'�uhr��#\�)����%@A���'��}� a46��j��B%fv�3�'� ��2e\g�����N�b�
�'6�U+�i�r��p*ἐ�iъ�y�TX����׬A:X|T�����y�E�� ^Q�t��Oٮ� U'��y� ��V&�)���܂7�h0��J��yc $S$���a�,&�l�T���y�$�[P>�:u&���@�bJ� �y��R-6L���S�Ϧx�5A��Pyr�Ĉf���k5��AdDaP�e�<��m�6*� ��!�*M7�8���[�<9�-H48�t�P-�6�\��`CEW�<� aR���].�i2'Gؔu� �"O��c���Z�Jq`V+XKj`�V"O�x�sk #*!�iU��QA���"OL<a�/ü0$Wn�(�@�"O���H);d�K�=l�l3"Od����]�6�R�BՊ3�!�"O��s��-)n�k'�7"��՛1"O�IbWě	`z��p�Ӎ%gZ��s"O��1��M�f@FLKr�fÜq*2"O�Թ��^s�X"d ]��H	�'�.���D-xz�Q�
�<3v�
�'ۚ��L{|��J�)ʺ4d��2�'���f�Ϧk�N�#�.���a
�'[�`���"�z�jg�V/�\*	�'~�Бe%uk8��e&ڊN�n��'�r�2�aK�T�QH��y"F܇ȓy�k�.��Z��L�Ո^�F�.t�ȓ~S�LQ��C*l,p񙵌Z?;kb��ȓ���͚ؖsq�)�U"M�c]^ن�wj��ٌ
�"�	aBEpѸ�B�'D�@�$ز7�@�u�X�aj�a�'�αZ2j�52c,��J�SZT�1�'����Ƙ'`�J�c�(՗����	�'$v����0�޹�&d���	�'<� 15O-�^����Q��'�VC���±�
��r%R
�'����
8y���Ic�"$�	�'G�("$+��#����K����	�'n�1�0OD����զ�w���'�.l;�Հz��#�Y�s/���'Gd�@��\����0e�g�r$��'� �Lk-B�
�E�)G ��'<�i��q�n�ض)� �$���'��I�f�V{����T,N��Q	�'��[�k�]�2�+��EH�^� 	�'��<����
���v@;2|Y�	�'��S�ڰNޔ��/:���a�'�nh�P�M3�S�:f�#�';4��TL[-z�Y2q��5I�2���'��1ä�&v�������Gʞ�Q	�'��ѕo�:>��7���?� m!	�'Bh�w�܆@�R�"��K�9ɞ���'�<P��5'@�4(L�[�0K�'4l�R`��$rXP�:�H;P�A�
�'x4`���
1�%֋KZ6h��' b�i�.T�!�&��Ç�k���y�'ݞX��$�,N��̪sc�V9����'��Q9��,<��5)��F���'����u�ɌE��fL�uo, �'��}�g+��R$E��ޖl ny��'�效�/�wάŉ4���b6�(�'�Z�R��B}�A	��
5
u\UR�'rp����X�X lQ��P��*<*�'��t���F��y�.�s&Z�j�'�$��cD�/l~��48��	�'N̽�!I��*�K�E�(<p�A�'�Ј{�E�FЙ:��;j��'�
������ɀwHݲM��'�z��G�����I],,h,Õ�1D��*.�j����ОT���);D�X���6-���� �� 5��i��,D���M�=l�2�X��"��=y�,(D���w���v�����)�����*4D�h�4J�>Ϩ���I�uR`����$D�� �\�Sˑ�V�������6���@�"Oxͱv@��#`}��1)��-�q"O�����?�����/{�F��"O&4�D>�|�a���/�̉J�"O�Rb��.�a�S'BG�1�3"O ��M]�n�^�R`F�:��at"O�����P�f�����$J3��c�"O� �`lׇ!5�C�8 ��T"O\�{f�?*��*r!��q0�IQ"O��W��`���w�ąX �9�"O��G�	(�����/A&���"O�<	�I�j�Z]�W�;<�n��"OXPpE�FN�ܝ+�%���:�S�"O����ל;�H�ګ
Δ�Ps"OpC� �!# \1b1�db��Q"O6	y��=cX��3��g�4d�V"O&��r+B�#��r� �\�V�<y�<{Ƣ}��MN�F���AP�<a�$�����@Nl(���AL�<A��8[`��䈈�l���b��y��E�K�蘨��3k�8�b�J��yR���vD(�EQ�L��4����y�
�	R�e)��W�>��ۂ.H	�yR�S&|�*���#8���9�"ʱ�y�&N�x)G��/6���[࣋)�y��]�Ynht.�7H$�����1�y�+����\Q�i�WVU*U�M�y�B8T�	�ՅѢse H0��X��y�_H��q�t�ɷU�\E�  �7�y��D09���π�!��P����y��ُxlN��茆/�n	y"�#�ybLH2m�3� �4 �t Z�J�4�yr-Z<Kψؚ�E����b��E��yb����!Ώ��4C��yR�M5"��a�Q	�5�%���y��� ڔ[$M�8*�(h��ڃ�y�kӀJo��1whO� D��y�bԯ�yBeB`����Mш�����+E�yR��b�����
��fÎ�2�A�8�yrg�6o��`nT>�vx��Ã��y��"΍3s��	����冥�yr�b���R�,��p!چ͓�y�f�o(~93�Z�u�$
�\��y�a�U��G�k��ԋ����yB+�
f0I�A���\w"#$���y�MB
�z�Q�j�/G�% ԋu��'ì�p��E�A�&��!^>4���'��.�t�x�r0h�&b��P(�'$��rp�G	V��tP�2Sp��'��3�L�'(�=��f_�7���'W�Q���� Y$ ��,��*��	�
�'�ƨ �V1
*�yƇ�#�z1h
�'W��[DA aT��0��r�	�	�'ְ��	OD����r����'h��`�̛-�(�h��%EED��'Dq�,��L�j���B��H��d�'Ϭ�p�F0�����M vO H�
�'Y@�Z�n��T.�����ٷ9'��
�'��1���v�p��N�3[�Xq�':q8s�ٕ���q���N�t!��'��˃�[�d��30㙹J� ��'�|ъ�%I�s�\��W�6�L��'��T�P#�)�@��$&A�Ps�'�0�	q�G�9�����E%<������ �a��R-���	*�'|/(���"O���u��|ʊ8��	�-���"OD0�U�D?4٢�ЈV�Ac�"Ox����9� KF�G�t���5"O<m�q���r�<9GO�S���"O4TڥeOv6p���'5;��!"O>u*�!`��t�2B+� p"O0�I�)�S.�|�"˓�W!�a�"O����J%�L��#D�"S�=�`"O��3�lT�F
Eb�_��""O b"�?VU�QҤR=d���"Oޜ1���\���skEa(ڔ)�"O�PG�+n�ݢ�	�Y�,5xE"OTt�Ul6��DAbI-br3�'R���i�J�>L�\z`�B�od���=D�l��C%��@T�� z )"S!D�̸��Å�	�ѡuLĬq4a=D�L�gY\غ����2Z�1a�7D���J��z�I�S�Z�t@ڵ�9D�D�##�c*��ҠjҚH�x v�5D�l�� 9 =X��M1N}F-�fK4<Oj˓��䖤q��(�A�*1�!	Ӈe�!�Ć��@����P |L���B�82�!�$�f�0tFA�*(������>!��@�-���@��3pz����ɋf!�dL#w%�iW��W���Q��]�!�(F�bp����&E�pQ�g쐅&!�D�4b�� ���N?"܆m���)��}��d����e!j}1�l�6!���9�i�<	��hOq��Q���U=J~D�C���0%����"O�����O�?�P7��--;h���"O<�y��U�w�C��W5b2��"O4YS����N���Ѝs���Z�"O�HC�o�7&�T��!�m��`1"O[�#��cv���
]��}ж"O�<��h�� 5�R2l��|{S������B�Q�[�	̺,r4�ѪR�RB�/V�.Q���V��n���C䉙^p���2�I;`�(���مC�C�ɸU��x�Q�ʹ)�� �7�U2�C�	�*O��F�?��9q���k �B䉻�䉪vg�fk���7�TO�B�ɴu0�u�$�7��� ��M���$4�\����^�(��c��Z�6�`�I2D�415NL�R�6)a��=F�
	`�f1D�H2�����
}*q��F�b�#+D��IR �2J��3˟
	�3�&�O�C� Y%��7}rNYh��
�$UF���V���SE�]��##��(�؇�H��ݩ�ᖍ��@#� K'F�h��ҟP����*f2�#�'��.r�Q#V<o�vC�Ɂ��у��)���T�|�B�ɘ6&��	#�R;`����B��d�BaAR��y�.���J�FB�	c)*(�tH��G��#�S��vB��1i��H�� t��db'�ѧ)�j�O����?���V� �Gb0�*��?`)��'a~R��1F$&��PO�[���2��y2��
�|�r#�F@nq�rc]�y��[31�&�	�DܬD^ڡ��I��y�.�
,O�|A3	��n$~���d��y�cV2ij
���k2]	�	���y2*M�R�@4RT�G�h�� ������!���'
L���E��r�S�	:$)����?����9�S�? 2��� ��P\��jJS<xp�(�"O&p�$�4��	R�/U! �""O��Sd �$U۰x��]>-��)1&"O�l�0
�?q�kX������
:��'��O��I��Eȹ2�쉸pF�A��p�'@��`K�g��5�"�ǿ� ���x2�S�i�ĘR�$=�A3��V���<���PF�J�-H�]�4Z��a$!�dR�5b���J��;�h/13!��17*�5�׮oӘ��ȅ�!�ݢjj��iÂ�}�:�{Af��Tџ0D��D�z��'��.Qzڜ+�O���y��ȀK��� 'R�6p&��th/�y��/1LɰB�.~����ϔ��O �� §�� �W�8d��H���ܑ~�ܨ�ȓe�"dhfj� �H�	�� �f]�ȓb-(SD��(�$<A��/32=%�XE{��tdZ�,i%�%�K�9<�b�fC�y��I�t�΄��f͜#�|P&-��5�&B�ɔX���צѷx6�y w@�+`&B�ɣ6����I�^t�����s����hO�#<���sԮ�����e������E�<�E�M�M��P��E�B� �a��e�<��KJ -��PP����(Q0�(Jb�<����7Ap�UÓ:3Z��+F�Ne���?Y�'P�;�ꌊX�D�dF=F>�����X-�%��A��kq'US`桅�mP\�d�9�^��g&��Yp%����	�m�Be����|3����ʯo+�B��1�,�c�E�!Y�� s%�ܾ=-bB䉶$���um�w�̄"�+ܟ%����D �;�{����`�"tEۚi���-��<E��GV#v3��829�°sB���!�$Y04Gz)�U$1ܤ��f���q�!���`��N��o��E"�%���	nyr�)�
N�R�x�Ҳ��8�.qr%��yB�ĸ5��`�61�`Yk�L��y҄�Q�D;�m2S0����y�`��j�r��B�T1[�05㡃����hOq��-��J�k�Z�I1�F��25"O>�A�D�QiT��b��s}BT��"O��{��J��(�@���~e{��'!�$��F���9ŁP=~�$;��݅2�!��_���:D��"5y�hY�j9�!�$�
_nݐ�T>+	����J<]�!�DԜU#�(���aXMم��w��Oң=��j���#ߓb��`�q�Pd�E�"O6]� ⃇M�$����4m�e�g"O���wb����rtG�!)B&	��"O��ve�7C1��FQq�d��3"Ob�)�"ŧc���8�$}8��"O����ΒBf��N� ���"O
$!&�j		�m}�-@�"O�$4���F����+{q2�¥ 8D���W"W�1OdA	���MK�����O`��<I+O?�BadΣ�&4���V�7� ����c�<)�՞m�6�G�0p�����a�<A�IJ.O|��2�O\:k*�$�X\�<qj3_I�q� ���|�<�s��FK�'Uax���<�{t����p�!�Û�y�jԧ;H�[�eK�&&L�P	¦��'ў�OZBPrC��=�n%i%�N2je ��hO?�!��kC��c �+Pe��kdb|�<��� p`�f���L���p�<� t������y��W�Xf���"O��R�U7�pQx��ӝ��
����O ��$ �[]6��p�X,D���1.Y!�͒;*Ҭ��ʙ*B�$)�3��NU�O�=�����>ki�U; Oʫ6l0P"O�ȉ�o�J1힎-�b�`��M�<���x`̤��+A. �Hb��K�<y�̠I��IVnÁ��Ӡ��C�<Y�(̰]�"���J?1i�ʘb���?�Ó=>��P_/��S�f�	(J~��ȓx~��#
� �:)QaJM@�Θ�?���~�eK�)��})�,�Wc�X�s��џ�$�l�����d�U��aBva�%�a���Ĥ	�ʓ�?�+�8)C��ȏ	�b@��4Q���!�h���� 2����FR�,]��ȓ8���Y�cX�%A�	� �(������ry2��nE���$	��pC)�5�!�$�*6t�K�㖸{�|-(WJ޺G�ўx��Wt ;v��p��U��Ƒ84P�D{�OB��y��D$C򦕊�����؆�ɰz��l�gE�>6:���ߊ=��C�(Gx��`����W�"��, ��B䉏C�H�s�]����3E*�H�~C��:�"]`��_'�p�8�혩>�
C�ɷ˨e�"A6�d��#��d�&�=açN̩�s���
p�Ӫ�D_����N�����'��'��|����
^S�K��l*��c1Q�T���8p��V(�5[�Dz�!!9�B�	�{2���k��������ý�B��*r�.	{A� vZ�AWoC�EpB�	c��PXc�D2$޴!��eY�C�I�|����!b��0�@#w��C�	 +5Ӣ/K�A��Xp�	�Q���|G{��'���HG](U�����n���)�q�!�$�%p&�Uj�/�o���/�(*i!�dZ'>��X����<�:PQ���0eg!��4R�,T�NZ�b���"�q,!�9g���e, �{�pơ�z��d#�g?Q��!y����g�8|�$X!(��I��?�}���E�F����P7E��#�I]dy�|2�s��A$3z��B̖ �p�X��vy"�'}a|H5c> yyO�6
�@-R,�y�)31|�T�DBI*;��In^.�y�f�pߒ���Ҵn=���sn���yR��(,dQiD�h�$����?������Op�g�'�"��W��u4x���b�5�&y@���'�a�T��I��} aLl��X�
!�hO<��$�(sx �o2m��T0{r�	`�'\�`��I@�,�;k$P��
�'���W�]�3v��R�M�f�`��'V"yk�D#)|!��ŧKV2���'�L�G�ӄ#N}��k #pK����ľ<N~�=�֣��_���Aǆ����;�@�u�<�R%��[��aeꐴ/��+#��g�'a��L��t	\ms���b^�9�A��<����"�z�x��U�s\m��I�	[i!�%kr�4Svc�L�H	�G�
�!򤉺1L�P�j��{ͮ����I$��	O��(��m(��vL�鄌ޠuO҅� "O��b<b>H�R�"I�؀�"O
�z� ݅*aPjsB��(^��Q�"O��i�*��C�R9�p��'E|İ�7"O���#�\�+�,�*��5VHfp)�"O�q��DG4�( 
���4=~��"O� �1ѡ@,E5:`���Ѣ>"x�"O0����yżhbCdK�Q��1�e"OuI�.>h ��!��(��t�"Oh��!ng�K���/(��A��*O����ސyj]Q7읺C���S
ϓ�O�(��B�W2�� �:|��d"O��+�N�n"l@p��O`�D�P"O��
c��>W&�a��l��y�PH�g"OJ,p�@�%�0�lH7?����"OA;G��vVT��*
;B�S�"O���`�"�z�T#߰E*����"O�(�)_&#�����N��Qw�'��|���͌4���ӡ(��d���B7D�x#w��9�r �DEA�q�(9��f3D�`a�+�Z+ �l�)�5�a�/��#�SܧN�̡#*\,g�
�
�Z�B\��+�v���*�>�z)ز���{�H��ȓ@� ��G�S�cH�Y�AJسX�l��0���s�� ��
e�3����ȓ6�(����oV�:�N�%bl��ȓK�6d�c�e=����� s�-��6쒼a0Cíf��;�D8\���ȓx�H-Ґn�]���E�V�z��ȓ>3 ��siG7uEr�"W�T�W�pU�ȓ%�r�auM��|�e��p�:@�ȓa��0'!�:/�т���R�A�IƟ�?E�T�S�C1����5�IAԗ,�!�D }4�k� Ë�0p��fצf�!�ğ�?�<l��MW����A:H�!���|��a�^/b�Xh5�B�!�Nhq*����A.kx
�I�!�պ1�fy*hT�88rc��8�!��P�_���W�[ ٖ���[5��'��O?}�u	�o)|u��@�t���#�/�w�<��# 3È�-Z:A<��uO�q�<��lY0ov�-B-̾MB�a��U�dE{��)�pGd A���!.�|e�P��=G0C�I��� ��mV!�e�הi+bC�	5~����ň0�@� 6n��|��C��"e����	[�:a�7ES�E��C�ɉxS���!��Y��!!1�B�I
V�)Ā��V�:�*�n>GU�B�	K�;�JG1O&
p�&��WXB�	�e��,��ĳa� ��Ȳ��C�	��lѩ��VJA��A�
�_\�C䉉Hpѣ�D!���G�J��C�ɞ'ݦT	EL�#p?�p�ˇ#eN�C��]�tD 5�+T��(ՌG3mjC�(#�,�`o�-�n�`S	5#	:C�IL�(��ƻ��@ �5wI*C�p�h(�"�Ͳ_��	�A��dC�I�\>(�������r��t��C�&b���a�<KբT��`@Ns�B��u�e��̩+cҌ
���9WJB�I�16 �Q�V���٠�j��r�B�I*@@H�4���k�hA���B�	��r����U�6m�H�f��oO��d4��T��~"��>|}�QB�䘼3�P�h�L�
�y�h�%��5�
+FC�
�-�y��[	��R�,V-�0�"�8�y�M_�M�b�C��;0������y�']=����Q�-bL���[��y"�S�{��l2q�>&�&ŉ��2�y��=�|���!~:� I�y
� ���t+��4ʐ�3�!�<#�]��"ODف��!)�hY�`
e.�adS��	ٟ,��KZ~P�p��.c��Ȼb��%6,C�I(J�L	�f���j��P�A�'�T��3�.�@L�g�	�_w�<��!F=���Uz|4;�$�!%,0��	�8"�L���C\��e��G�<��cКHeJ��ȓ�����P	"L�KTBQ0 |؆ȓQ���*B�X�C*����R�+~v�&�0��IC��س�˫Oh$)��q!�&D��  .N�F᪨����62��&�O�#ؐ(�!���T�kݟP�HP��Rk��scA˂2l@L"#�>Nʡ��<��*��κD^l�q5�MEt`���4�\lA�,� L�v�"�Ŗ'/:J%�ȓ%��iP'�E��y3��+y�����s|:S�Qs��5��D�#! ���;�RY3d \f��ٞ��D{�Z�HG��&H� &� �Y�B�9R�y��%X1Jܙ�1QHT�+$S��y�����g%�2B�d�dFV�U!:Єȓ�l �J�;�89��Ls�QK�m�<��M� q����G,���Uf�<A���l؜IE"̟]{��I3�Y�<)%H\2%A3��H�R�E٥�K]�<��/4]��9�d(Ɠ$�Z����TY�<��m� ���b,��;%a�T�<�3��G�A+��18ld��
�M�<��L�) ��"�30���s�R�<	g␪4O�	�`�G�yힵB���s�<Q�#ɫ7$�QP�A5*9�� J[�<���G.[̸�x����@F2��Y�<�7���R�"�³	�+��l�''
M�<Y��K7V �XC#��� �4�bW��^�<�gGS6| �12�����r�Et�<�Se��}HT�Y�JX���iBtțm�<i"EHL�M�g$��
��I"��Q~�<��g��P�P垇0Y��ᓥ�}�<�H��vD҅f\�n�q7�@�<ɇ�	�(4D5S��J�Kt0q)3�Ve�<�.	$�����L�7�����WL�<��Ŏ�H�����тj���)AI�<ѱC��x�@-q��QOZ��'�MG�<Y�,4e�\��G� 4lX��N{�<��E��IS"���L���w�<!fB�a9)k���+bx�H(�lPt�'Na�R�}�� �J�����+�yB���Y�x��_�vu���@
�y�GKf�z��E�{�p4L�y�"�[��bYNZ�a��O��yr���Lx,�c��(�"��y����t�.�\x��5q3�F��y"���0��HH��
.hD�� "K�yr��jZ����H
6�*�p�����y�@� U5n�K5e�d�`���͕:�y"%�I�X��b��V(�`�]��yr���9p��S��R��0�y���p�x�BXE<p·'��y�	�=J@�q�E�q��j��R��yҦV"j�,(2j�h� �U�
�yb�/E�|���\Ud����M�yr��B��=��E�?S�"���K-�yR��?|d�S%JH�s�a���M��yң�� ,#�-Q�B�亠KN��y
� �����q�ؤ"�&�9n٢�"O�]H�d��Y�<�3'ܡr HPq�"O�pe�%.vȐP^5��!@��'e╟8���JY0���
��P�%D�0B3��:rf�q�����Q��=D��
�Bґ"!$D:�L��}��H	8D���CI�TItH��>fς�Sa�4D���&g��*�����ݖ�	�dC.D��P�����p��',�Y��K-D�h�!��=@`��Q��+lp���/<O�#<�m�<f&���L�?�l��cKt�<q�͏l/����û�����j�p�<q����Gc�q��ɑW��T��-Qi�<�qC�Y�I�.Syb��S|�<������я�Z�xաQ-{y�'Ua|R�>0�tqP`Ǐ&^A�#ſ�y� +� J#�?����NB�yB�Z7*@#�����Yr 	5�y"�O�J~�QAa͐v{��[��y2b	 /v�`�AmKh�b�S�ހ�y¥7+o��H�δa^F�����y�%Y�z<q 盒H���Z��&���0>IQm�F���G:Tk8}
���0�y�b�%T���*T�>G�d��/��>�Ogç$L���·O���"O���<b캕.�,	�t�"O2����7P�CM8-ٮ�"O��H�	6-���3r�R�(�<�"O�ITM�7��ز3 J�PBԩc�"O@��jK*=ژ�jRA�/����"O�@�/KXR8�Q����-3 �'�1O���#�&�|!�a`�"u� T*"O�DzRi���Y� 4O�̰�"O5X�n�"0��Yd�C$7�Rؐ�"O�� Ǆ��oG�QS/�
�b�"O�\q2苩F�r@�u�.c�v�"p"Oн�Ч��6�C$�$��@su"O��	a~P�j,e����R"OpE�I�y�ꝲP���z�>8�"Od�#L޷k�^E�����Ub�"O2�D��:�ܴ�g	�|�G"O����G�F��U�V(Ss~]�"O��cWؽ(��ب���,l�à^�Ԇ���ar�<��oР$YD�V�m��C�?!0L�9BHB���!i|�B��1qW�-B�6�J����H�D�nC�	��Lܘ���6 �Bk�6?�C��7Rm���7h@;�a�$s�C�I.+���ȕ���٘�Ă:�C�I�/^�0����;1L�~g���0?!�LH�qL�Y�c��$b�`r��d�<e���,�S��98\�K
|�<)��AˠtbQKʜ7oЩX�DMx�<��DD���xѶ!��!{ܸ0��^|�<y� H8v��ȓ�M�!v����̞|�<�g�h^剒!�7`��$I��{�<�T+�$>�Mb�&���"(��Wm�<9&$5j4Jؒ���$B��i�/�b�<���\ ��{�i�x�v��D�\�<�foǞQ+Ɓ:�G��d�&=�Ō�V�<A"%]<�8��� 1}?xp�AN�{�<��eC�R1���"�6��:V�Eu�<Qt�5Dڢ���ō_,�|*AVE�<ᅮ� ������kM���ǈ\{�<� N+�b\�drRi�Ģ������"O�a�g��<���[,%��\�R"O�Qc�J�U��C��=~,�u"OҬ�s�PM��	����.Sb&���"O�I��ƽ)�� �ó_���"O�a���	P��Hӈ�)H,ֈ��"O Tz"�>H�TH4�#2���"O@ ��ץvM"�f@-z9�"O��8/�l�% �;6�tĉg"O�ИQA�$Y���cƍ$v�)��"O,a�	�G�"�yR�@*jGx���"OX,�w��?�,,��L5D��!a"O�P�*��*��$��B�q@��B�"OFxp$+ծ$�V0yF��fM�"O�=q�V�-�u� ����Y��"O�Mq�'ŽoH�	�7��j�"}��"O�r�dגq�HA�O	�;-jyy"O���b�6��
0(ܨ� �Z"Or�4*SG���uZ�I��"O�-���I�d/���	��p"O�I����3�X����S$<�0"O*�B�΋c�D\(�b˷"V�YS"O�\� N[#3�xH�n�0{R2囶"O,Ȱ���A���Q�G҈%6L�P"O�UHp��4h=���WdB4K�"O$���H3c���#�Ꙥ= �Dj�"O�`���4岦�nc΅P�A!D��d�]�f���{#l}w�ә�y"ަ7Z���"-n`���F��yR��w�2�s�j��'Pu�F'U��y�E� a� 0H&�E�	�bh��)���y�*��uy��W��D��%Gѣ�y[!!�ezC����\ys���y�	ݗA�p���C�$%"0{�-���y˜*cZ
�(߿L��"a�7�y��֮N����b����� ��*
=�yL�~\�x���C�T��b����yF�F��z`@V�J���"���y�!�!R�Q���i��3�aS&�yr.M:LT$��t��f�X�b����yr!
�AB��G�\�(�� X���>�yb��!$�d��BӸ� ��RJʭ�y��1Q���1�Q�CBl�,���y"O����!@�Z8J������y§H��$���.4u֗�����ȓ8< G)�6nE6|q�M��Rh���!���;q�ݗ��pQ#�Ǉ0H�ȓ3|�re�#J
��*_/:�P�ȓ:�4]	̓�A��x���X"i����ȓ~}��,��0��.�0�$@�ȓ|<��c!OH=o�8�u���\����ȓ�JUXd��P^&e�W)�܍X�'�$�A�d�/6T�`Ju`
��`S�'Q:��g��r�r�B�ai�'��h��cB�$�61�D�_�bH@�P�'.�a4hθY�tt7�Ԟ0h����'q��ү�!N�d��fʅ�6�H�k�'�<�@��	)�RfՐ0����'���h�#�!�fl1a���/n�<��'�L�a�%��H,���F�"�����'Qz3+ׇ$�E��E�:f��H9
�'�4)�R�.<lШFhݼJ��R	�' �3�l��M���C�(��p1�	�'Cޤ:�,��`�y��A<������ n����]R�Sꛂ\���T"Ot�j�*J�Z��Xx�h�X��Ke"O����aJ�Zu��#��
P�N�`""O܀�a��.7��������"O��&N FGb�0��VG��Q�"O(���G�-Ţ���0w:�|�t"OL���AA ����R�P;HH
�"O.��� �)����eV/�y�dg��p��يU)H(�� 8�y���Y�<�0LL�#2�����
�y�ߚU��$c�ϝ"���8ģ��ym�7Z<�Z$���c���A�*��yҤ�5l�lbT��'aL,D�I��y���?	�50b�տh|
��v!5�yA�-W����:e���5(��Pyb���b� � �Y'dYt�~�<��hֳ'� �0���6I� ˕.b�<�l��Vp���l@�wi��qr��E�<!���+Z�p ݛ"]��;�
C�<�J�}_p�׏W�"��Iso�@�<q`Z�C��rv얆it,��E�<a���p��GC)TnXⲢSB�<a6�[$(�F��.����	x�<��䘻�@���$@e��!F/L�<!WhҖ�k��O?&#zU�&TF�<�$��<,<c"́�0NFh�wF�W�<��� �!�0hw�,~�T�s`E�Q�<�2挹�h�R�ʤ�����D�<���-�����O�]ܴ���HZ�<�+Ӽ*?h�$�#VaDek�<Qb	G�M�-��B���|�+��h�<��E\<������9�J�<9Ĩ,�^IB1jŝm̾qҦ�C�<y�끐/�PZQ'ۜn)�VC�<Ya���Ktq�
�?$x�9A��}�<A�Kз��M�B�/7��#�a�<)��_*xΈ!�Ȉ�K'����cW^�<T�˳D�Fy��͋}��T��O�<Q���N�:Pu�Q#;bR���H�E�<�w��g��z%�"'�$b5��@�<a@�˯fd�h6���K��G�U�<�#�w��E)f�C�{����&MK�<����r����s���1�sJZ}�<���\9#� Y[��S�w�
q��"_u�<q� ? �ҹ��Fےqk�i� �p�<iS ���:2heJ�%ӣ��h�<������ G �H���Z`Ab�<���Ec�B�qwf�aq�ec��b�<�d� iBY��@<H�����g�`�<�b��Zv"ܚ`+��Ux�dF^�<a��Ԙg�Z���MΤ(^t	�«�c�<��- L"�d�F��.=@
0g[�<�5�٫zcΝ�b핤Dk0��%��~�<I�.к?^αH�!'z�f�i�H
z�<�A �@L4�Z�A�.`�>��pC�y�<1�k�a�E�&o2�=* 	�P�<Acㅕ_�"ų^�E�v��e��B䉃;�z�Cׯ<�Dc���Y*XB���n�0��
�*�#N�1�RB�	�}@2ਂ��8Y�1�@�76�\B䉴6\�]#�`�����m�9jT*������9�E�:jT%���6v��ȓtd����@�c����s�O2洅ȓ&��@��gZ@���y���S�? <�� ��93R��,��,&���v"O�H�`B�@�FmЧl�)j|Fl��"Of,{�+ [K�D�+��,hn�h"O�����V�6�k�KA dSY�S"Oc���+j��Tq���xԨ�Q�"O��bLQ ֠8�h�Z�XPQ�"O"P�W
X�0�f����ܞЋ�"O^0�t�ِ$���*��Tr"O�y3/ɑ��0�UDօZٴ)�&"O`�Zg�Y�A����e����"O�����DU���RA��&�渋P"O�(a%
8[�,h3 ),���ae"O�����'l,E�u���F�B/S=!��H�o��H��o["`r�04�!�D��{Ɉ��'ʎ����U&�?~h!��A�;��,�Ł���(Q��N`!�d]�]Ҁ�c ��MY4��N�!�dҨ;<̉K5��6άQ���9"p!�d>?��h�#�+̮��'ݼC~!��37��1'��]��u��'U!�/��� f�̈GxF����]�!���
M�`����f��5ZƉ�2�!�W�8� ��J*t�$� OV T�!�ċh/~��f��D�re�X�M
!����Tִ�R�A�0;���A�Եb�!���d��@��iZ�d����%Ձ\���B���(ӕc@(൸�n�y��S(�`�sf��L��aT��y"�J��x@̑�ND���y�C�:W��0 �vw�!ݭ�y�.�u�J�bT�V����"��y��[�&2�9��<V�l�AS��y"�E,1Ԅ��E��Ic�Y��y"[[m�s��GC_"H����yb�\�I<ʡ�F��K��XCeIP��yb�	>�D�O�@X�m`�dH��y�Nڡ9j��`�OW.h��#W�y��ڀ`j��p�랪A����ȸ�y�F� sI�ݳBͯ3�:msR�V��yrm�y�=��=(��X��N>�y2� �!�)��� ����'��My�J?!h�p�>�j���'�<DA�ɜ 8@�H�$��m.���'���l�?g��Y#���_��#�'M � �Lv�lT8�H�]@RP�	�'����҇�EVP�5i��j���8�'�ɐCO�X�nl�D恴�ܘ��'0�C�I U�x5b�`��� D��'X��õh0eP\���ۭ	H���
�';<�P�D?m��2c{8�T�	�'�y:2!�D7���I]�,�	�'�0U�C]&�i�
W"Eb��
�'plyBm҉(�V=Y��Cs,�
�'a"�A�F���〒�	�e�ʓa��	CV�R0S�����T�V�,���K��e�����̜Y��]ި��M0���e�� $�t����`����LL]96O��5+T��2���@z4$
%�N��J�2��L T��)�ȓa� �Z���M�}"V�;W4Nԇȓ1�0MU�J$#�
Q��%��=A|��W�~��2�.?i����/��5�ȓj{b����U��A�aT�L��5�ȓiZ4��Oſf��DQ�*�T؇�S�? ��0��ݒt�p9��B�g�\�S�"O@�%�H�?Qd}�v�L�Z�{�"Oډ�T��\���X�D��6���;�"O�Xピ5h�<X���v�,P��"O�}�a��F�>�
���-3�)ӥ"O,}$"�H@	(`(A5G�X�"O��IBo��slDehcf�KL���"O,@˴��%	$L�y5C�-�p�f"O����6rD[pAÖy!���"O�l���	�;)���&F�N-z8 "O�uau��<P�����&n�"OR���֫)(m5��	;�\Bq"O���i�/�Ҁk���,�0�є"O���0�6C�����Jǰ��t"O0�{&�('�`V�$�P-��"O�傐o��j�|x@��:W����"O"m+�T�~a�Q�)K��D� �"O�MV�
p[�esvo@�Tq^<��"OP�#F��A�$N�v�.q�r"O��#fl֦
�cWH�'��}ғ"O,�#���H����+c~�"O�H2��6���@�3Hx�}z4"O}K��B�,V,���1>n�E�P"O���@�*��MY��8�@G"O֌Y�U@���.Y!F�p�"O�Չ5�7���c$O I�8�A"O@�3��� G��R6��(;����"O&��֣ *x eb�)\>1���:�y�KD�nD�D�ʼSvd	�2�yBL�9v?�����Q;d%��K^��yb��y�r�*�Q*j�Ä��y  �J���]AbxղS%�"�y�EL�8��	��Lڼ@`�A�ᓺ�y2ɰ �PIZ%�M2����R��y�)�P�ly�ׂ$/j<Q%�^�y"�F4oWn�g`�.`�k$Å"�y"��L�41�wd�+\oҤKd"�2�y2!IS�`��Œ�h�H��$Y��y"%_�ibD�A��W' ��`[�y�cP�yR6�K��M-LAa�[��yr
�KO��@��ML
zx�T Q�y�'	�Q��#TA]�[QV�q�α�y���?А$�
Ü~����Ad��y2 ��*�q����}K,es��A��y"��=?�*��DV�z��$�E��#�yr@�����#A�P�;"�H��yb���7��(#�ް-@��f���yl�%u�~$�5�)v�(����*�ynDҒLAe�H$ ��y��+���yb�X
t����;tĀ���Q�y"��?
� ��@�yJ���M7�yϔf!,q���7VH��Z��y�a����6�SN�P�p����y�"͞#�`"֏8:��b���y���>[^T�9�d +0k�x�S�y"ˁ������H5`��ˢ*��yR�y�=����XW&q������yB+�/,�D+��[�$�8a���yb͎�l�{ ��7e���p甈�y�h��r�f���,YP	��
�yRA����u@ �0T	A�����y�,ΊL�0�"β)�Qg ��yb�GBނD
W��f����j��yα%d�<���cM�8��ሬ�y
� ���5!�K>rB G2�@U
!"Ol*���U����C���:]vQb"Oʸ[P�C*"��= ��q%�C�"O�� ��#ߠ�q��c��$:w"OHX��м͘���74ݸ���"O ��A�M���1�D��2#~̨�"O�-���i lH��"@*k&��"O,Ms���F�������OW�T�"O�@�f,ڣVsZ�3��'C8�h�"OP����5,�h��o�v6�	"O�)H����z���n�!'D%��"O��⃇�5#���p.Ez""Ot\�P�� ���Г�T��+ "O��S��f2����&DZ�9�"O.QU��+ީ0�-��C�ً"O�J��1ܸ��2����"O�4�&��63P���0�U��"O2L�iGYl���@�< �X|sg"O,�"c��.W�f�I�΂1�̴$"OP�+��d\TͩӮ��|uqE"O�"e�	�L���F�t��H"Ofi#���5ȝJ nL�>�X,��"O(��BC�F���I.ȑc���j"O�JSkE�.�@(���O��	*�"O։;��'fxBM�����xf*O��o�<8����#
�d�Bu�	�'���0���?T6HY��EE�/�(�
�'F�3 ��X�j �²)����'��Mɂ��{��!��_K�d���'V��N݆f����T?�|�(	�'�H	��]>�	��ڏ5��59�'�H�s��\9�t`aL��)�����'�^ ,;V��1xC�7�����'���1���Vر`P`�1+Z���'�XT*ͅ6=	 �@UȒ�'���'>jA�P����5�բͿur���'g-9',P3*�� +�������'٪��1�I(t{L�H��^p���'K4H ���R��t�ٺ0&D��'��xd�Sі�D�)-1�Щ
�'(R<��KQ!5� �Yd�['�ڼ!�'�v�C�^K�Y�#
��J޼u0�'8��@�����B �3YP�\�'�:Q�R Cc)l�s�eR�~��ah�'�> �v����TB��ݬHh>��'��L�W'̔v	�Y�!-H	B�J�
�'rDY�g�'F�F�"��M?Kz�K�':Jܹg�2P�ƴ�`OT76���'��a �+ؕb�H�{��^� �f�S�'�<����Nz���ÁF"88��'O�XF$�,1��3�ȍh|�	�'W& qqeO�[��a�o�;Y"P	�'ŴP��H�0Y�X,ٵ�O��U��'�T=�t��\~�au,��'c����'I�Dʥ�C�Q(����&����'Ӟ�)'D�j{-���,5hl���#�޸��6.5��i�,�=^26�� �i���M1LuvQ�ĥ:@��g[\�8v	�V���W�^�{W����zy�$bW��1˸0��'̦Bܪ�%��D{��D�@wI���V* �W# ���Y��y�e�S����C��V��Y����'jaz�i�i��(�%h�*R�� )CD��yB�� YJ$1a�0H�r������y
� |���.%F��cǒ�
����Gp������*jÏ�P���.Ӕ��2gO$�yr��/��<x�(ݐ'"T�b�N �~��'Z�T�4Jߙ^�f1���@1F#T<;�'�9(�Au�ؕ#f�[�8@y��'�JIx`���|!!��^#0�dI
�'4V�H2��>|����� �~�(�@�'KrXQ��b�����)V6q1��
�'�2�x��gq�!�6ab��B�'��E�lDJw��#�çZ���R�'7��KS�D�~PX�P袘b�'���w��$3����S&JC�y��'�D��^�]�T\�m�7�]��'ۂ0[4f�>o��zu��DāO���I�S�P2���$��i�L߸B8��􄨟�EZ���FB3t���[κ )|)��=D����*K����x�bO78�Ju�O)D��J�ǁIV��A̻R�>]�` <D�S%5m����oL�4r����,D�D���/�ƌБ��/K�4a�c�.�d5�Sܧr�D�FC�m�=�U�.ڒ��x$����U�i^X�BG	�X=jd�ȓ)n@� �2z�0X��W�4�ȓq��X�s��� � 1�,�
����nZ�)� �~�8�h`�/�h��#�^̚5`@�,$�9c�I���ȓ� �z .���aSJ`�~�Iy����P�Y�!�e�H�B�(�5q�H�X�6D����Ó;<\Աh���O�D�pd7D��#I̩Mͦmy�$	9r�4��Ad5�O"O|��� ]�+�> ��Z�[p:D�g"O��a ���'�!Vj��@�"O�T�t���~�.�pw�9w~^�y�Y�$F{��	��{=0�I��B�Qr����]��ў4�ቌ�Q�s�<[�#�]�#�.��hO�>�5���	f0}��I��~w@�a&�O�B���h���@L�L�}���^�@I��uX�4�<�U":W0���0�o���[��l��P�?��a�
.��ebQ��8_�,��� l�<	v��*��RSh6`=@!�m��hO1�����5,�f��Z)4N$�@"O�-�"V� ��!(�iV�����)4�S��y�AD�{�^�W?�:���j���yBL�n$4G�ˑ@�Ⱥ�-���y� �kI�a��_�=jԑ�4�٦�M��'��H�� K;@o|I�%P+7{J!:�'��ꐨX�.Y@�f��6�0y��dL8�h��<��F5VD�z�%��=d@Q1f"O�P����sĂ4Q�N��4/�y�oi�Fo�dr\��^�/�����Ye��3Rl"LHH���9*e}&���6�'\!�a���&�jb��E�r���X��$;�I���M�O�0⭓�+�iA�Tb���'.�I+���7V�2��? *��{�}�X��+�S�g�X�A�ŀ�2Q4i�qhG�{#=���T?)�L��Q�ₐ	=�BP��Ռ.��$%��)�g~�	�">k����K�g�����ē�p>	V��.7�0��kC,6o:�ôc�i؟\�\�� #�J�)8����&��i�ɇ�Idܓ�MF7�jUa��aJl��b^�'�r���)A9ST@겤�3a�>؋��Eo��	Ex�|�"�(!�аa�Up
`g�r��G{��W�,@C��=z����H�$����$D�(��j�9k��`�D?|�ã<�2
+�O� �y��AXj=���Y���u{"OJ2
�b�� ���;Mh�Pf���G{����'��U�R�/odh��� 턄I
�'K� �\?C~U��K�|@ ��y�'�`��ʅ�;b����0���@
�'>�����֫3N��!'�Ux1ts	�'�8+�"ۂ�5�UJA�jO��y�\��E{�O�-��f�6_V����L�q�z!`H>q�'��iRDh��L��'Xԍ��%�¦��t�)�'�a ��"&T}j�@�&�d$��	u�S�(ScM"w��c�e/SƊI��|��X#�JЗ
bJ��D��+T���Gx��)Zc�_��p�wdY2kΤXr��v�<!�E�-m�0I�U~8� UC��hO?牙nh.dB��� �F��D�D|�p����>�� T.U<a$lX�J;���Ä]�>n!��̋G����R����P,Q=azb�FY�sy�☻#h�0`�6Y�dQ�ȓEŬ0f ��*pNIR
�.-M�9��.x*0�JJ1?�!J��F,R�,�lQ�����v��'N�X���ǿ1G�@�j_+�y^3�:�c�i����E��y���P�bRⅹ;����ޒ�(Or��$ӎy}RI;b�	L�Lhdf[";�!��é:��q3#B�o�dm�gkA2w!��+2z. �C�;�E� k�	rƱO��h�}3Ǎw�D���݄��PZ�	�i�<yv�Ȝ�,�#�B�g_�@����h�<iV�F��1i �QS�Lҗ�^�<qEc7$��kT`�;H�d,{���]~b�o�O�����K�?�4Թ��a��!a
�'̈́�I�D�߮	3�F=]�΄H�'%ў"~��
_�L�.�1�J�-6��B&�L�<�7���xl�g ވ*W��A�RJ�<��EܶH�z�sBsǮH��j�<��eٺb�(�Q,T0 ��˳ɂh�<9�GȐ+㤤�g�5b0l�Ѩ�a}R�'cJ\��
χ-26�{�(�3%����'be�@�Q���+e�D<&���'(|Pv�V�{+L�*�d�9k���,�'z08�	#K���1�߯l<�����`�i�-J��Đ��D*n`�aG{��O���R@ ;r��l�![@Vh��'�v���`%I۠kN�W��\*�K�O
��G��o�6i����Po�l�����&��!�Ĕ4�܍������ڡ%���IS��(��(��i��-�����-�E%�"O�n�|�`aP2  C*�Ԩ`�x�G&�O	�0��+O��Ѓ%A�6��A�'��Γ{�!�U-��F)^P`鎧9�����5>����s��q���&"���Gz�i6f�~�Vo�Y�r�3 ��9��4��	�t�<ᱪS�#��؉FMR�h�G-�?yq��s���
�XA��a&�
:Ѯ@ǥ6D�葂ǂ-G�U�E�0 ���!��4D���W�H:@Z���m�1V��a��%D�ljC�Ub�����͡:PT��
%D��
��_U]"8(��ǜ3�,�X�n0D�T��]�͈e8�̅�U��]x�O0D�0��FB�� a�h�4���h�-D�t�E��_����������R$+D�D���!'պ�!��WPV!I#�'D�(y� �4@�x���M|HK��'D�R�+m�Н� ]6��i���3D�� �A�W��&O@r4r��D�R�5��"O��)B(�V���$�|���"O�L�s�(H � ����0�6"O4��W(Ȅ~�z���OB�R��)�"O�{�$H�W�% ��>�>�"�"O�l� ���keNΎyyX�Y%"O�(q
��C�:iۆ̔�Yh�e��"O�,�PΛ.y��*��/N%�3"Of��R`ސ:��Xg��_�H�"O��Cd <o;�K���b,2=�"O��;���W/�h*�%<P��"Ol:vG+H�p�[+�$ ����"O��n��2���7�IA��"O0��(D�~4�m:�@K�A
d��A"O<L�_����#-�@6"O$���X	dZ�3���7��@"O�Y����Ti�	XV'���e�"O<E@�ا&-�g��-^l-r"Op7��56<�%F�QL��Y�3D�d�B�l�"U���qEn��&%&D��q��Dp���@0u���D�%D�4!4�Ԁ�X�h f��,��!y��$D�Xtg_Ҭ����j��YK�� D��q�m�Z�8�g�\���i`�:D�PH$)�0	X)x��#V�ȹ2D��8��;^��;�"�be>ɡEM<D��`-�%��䲆gI		�;�:D����d0 +���(�+q����;D��c�,�.o�lЉ7$̥0�F�"��9D�D��GN0(̌� ��%��:D���f.Z7}��e��ܕ���1M8D�LZGd�p���e�ڄw�a@g�6D�i��+����%�Y�v���"D���P�������q@,��0$5D�t��19�p�q,��@!�y)�<D� s�IݴW�AH'a�c��)�� D�q3i��Mr9���ߌ^��	�e!D��*��/\Z����J������<D� ��j�����^��r$l:D�Ȓ�z%)P��[�N�Fh��拟�yr��&�v�qd�imr���*�y�#���4=���P�\Z�I����yb*�I�d�@�.W/�U�����y��"{�`	D��6Zq���W��y��x��c!ҩ<]9rl�Z�<ɀG�)֬t���6X�H���M�<qR��J@R8�c��2�"i"�e
E�<@�����ǖ�(�|!��	F�<�AT�}B���'À)�J��N�Y�<���_<��X��ƽ2�� �[W�<�cH�
a�1
���A�4�QPIw�<y���2C��Qpč73�^�A���l�<95��:1 \|�R߬R�H��@n�<i�������Q��/�����!�k�<�`KOܭ�"�M�l뺄�g�W`�<���
��Т`P$y��i�̕b�<�a͝w1�UB$��/��Z��@{�<�]36���³'���� BLs�<a��>Q��₍F&54 Y��EBn�<16� |� Q!�m'i,ܒ1��R�<�we@���L�w#O8r������NT�<&\��!c7%�gʖ��'�W�<a6kǘzzla�G�w��܊@�N�<�F*�;�6����Q�J4��!WH�<� ir���:�-�� �4Ql��1"OJ鵠H�����Zl>L�"O4����r�����R$P�qX"O �b��K�,��K��yD���"O�i@�g�O{��C,#I2�k�"ON`@�AM4��z�@�"z8j�7"Oh��#���p�$D�+���B�"OlpbpG��@���f�ξ�<Hz1"O��j��8 @�ZQb�?�L�;�"O
(�`�,u�����ġ=	�`0"O$YA��)H�k��I+N� }�6�'�舉���g.a|2�M< �����ϵg�`Pb�d ��=��W�Hɒ�! @�O �V@Y/W���I���0��Mz�"O��c^#� �5j�J��a7��%K¬�5�׍�"}*W7$��i�)ɩt�Ti���c8��J�)�S}"�E�A�=�b��I:.}���Q<�H�J��ݑ(�ʓF	��|�'Șk��'M���,G?	��#��ޣy�$�!��iN	a\���+P
9��4jV�K�m��8���"n�����c؞h�`$W�N"���J�5�<���N�Ld����~�����3�$��A���M�����+�r�`7h͌C��tS0�`�<I��D�G��8(#I�X�tT!���<Yt�K 7�,7��)n�m�R��
�S�.|y��"FH:xx���gK�	�P���G�:P�QX�'قY�Oڜp,:����.��jm�H���9��<I�j!�gy��J�X?�`�w'á��	���+�O�I�푔�ȟ��h$]���1�E7������4G�iqh�"RZ��$A3������	?-&��7kE�v]<�
I�S�i�(���rAM��D��#OZ�X5��@B�+َy���S�<9���
�T�Q�퇊	ٴ9��!�D��'W<l�@�I�Y��F�T#Y/C�|���q4�,����'<�!l�J�Ş.|���2O�#����P0�Dp�/� ��9?��ŏ�sX�#}�E�݆�0��$3[���jʣ]��i$���ʊb�g�E�GN�p��ɷo�z�rLڰ��ƢȨ��)�F�ԭPC�~r��:��!!
I0I$��qǄ�+}FEz0'����d�><OBQB@�H��lJ��}ڤ�R�ųb�Yp�O���FEV(�m H<ѷM��,D� `�<��K��rTM�Tq�$�[�'��Xa[�́@�+f��˲C$�8	�P P�� ΋g��'&� j�� ��AF����" �j`;Ed�"(��9�#Z2ʸ'���1�٤a0H2��F��蚜7�5S�
'⦜+�b��I���P�>)DE	����'n�=J���y�h�����0��t����"gq�}�1�Η�yiL����I#fWx�0�oP+7T�]��|������R�' %�C�,�J���W'M�pM8sO6:Ղ��Պ=di�D�x"�w6���)�ny򨍙y%���B�%J>:�S#�R���<�S��'O4.�c��ӟD�ֈ���M�"4����*F�bH �h���ēT�����jP�Rp������$��P�5�L-M���q�ɕ/J�q4LK�9Ⱦ�x�*�5��Ob��c�*Z���x�a�	p	Y�&N?t��/
"�B��x2K�;>�4�%���,81釣
��<T��#��\a���=�h��,O<�I4� ��&Q�)
>}�`C�BF�L"��Ű>�D-ȓd�r%C�E������A=ь)��ְ'V��x�)��m5�'N�I��S$��I%MV��eǂ�%ؽ9���'wf,�󄂷-̕id,V%qj4E0r�Պ)@eJ��U�s�R�\�̠J�E@�ɼ@���Q���I�/rnr�ђ�FF�bC]��'~B�#�����Z'�F(^�1�~�Cs�FDs�i^�6�(�P�a^p�<�ۙJ<�)/֡�xA�g޳n����4@қ$�v�����r�����v��h�BU.D��Ȓ7�^X!�D R�e�B��D�J�9��6�1U!ٶ)^T��W��剋'�Ly�5B�+W�@8��co0��Č�i2����	�Q�H�Q�$J�p��7_�b�j�y�a/$��Ƞ��>e������L�H�PUM+�jX@px���0@��?	��7Q�ıu%C+)�9���"D�<ʳ-λh���R`�܉0����h�OഛF�*ʓO?�ᑉ�+[��8�R55P<l*D�q�'�j�
����{��(Z��US���Z�'�L9����c���iÇ�������'^����(�>Yv�V��:��N�a�<N��q$K�g�\2p�׵yHf�cW�;4�� p��3ǁ|�5��lQ9��d��xB�Y w4��mZ4���IP�� `��Sz��̮4_��b��O�
	{Dt؟��Ff^j� *�KʂpYE��
b0�yz�i�rxi��*�@ؤO?���"W�~&0�h�"=p����`�'�du��a�x��4��Ǖ
FS$�Q���y�|�'(Q�Tƀ�>C�5��	���杼YE�P{���2~+��{�S��e�,?qO�c╻qbX�<��- Q#.]\=��~�l�ɠ�=$�`��EJ�Lߨ���G�D,ҡ��%����F/���E�zU�ԫTm(���?j!$R
^�!�O�n��"@#D��$�zU M����7�:��a �O� ��ES��`���<�O��x⤎�*��r$U� �-�q���>�QDZ�XM��za"ZG��*���	8>np�'�9j$��	�%x@��C�>x�ay��(QD��b2f�zJP��F@��(O`ʃ��)S@ȴz&V�y�@'?�+�,d�:��	ӗF�1�ƚG����O�rXI���N|F�����%4���-j�-k'��h��'���
J����yWF[;G/�}8�	��y�h@@`�χ�yR��G����V��qr,���J���n`�H"'�G�{ʢ$�P�	�`�Ը���~�ء���-�&����
P.�U�Bl�d��負�8oG���WO�5F����&��	������&9���\;�-����d���?�LۢJb40�̆3�z�{@g9�I�52Y�`jF"�# Y��KY�+����y5*a�4Ȓ�[�R�qb"(k��H���J�:��UD�$ ����)Nx7.i�����O"���շL��!ցޖ%\x����'����,J�4T�xR��(�����Ѻ&����pCU�%�Z�J�Y��#BH��[����2v%�n�Q��d��K�P��.�,��0C	���� F�e��ם(Hz8̨���lȼȡ�Y�q�I�U�L�YǊ�9��S�0�Y3���T��H���&<r���UL�*���n�6	=i�c'˸Y�P��r��<�`�P�%;~���%�Վ*���S.`��@!�ν*�,'�<+�P<˧O!����P%�^�1�)S#!
D�aѰd�qj���W�*B��)K��Q&�J��i""X�B!�0�~R�6y.�=1�E� �� �?�p<��$GpR,@9[������3�.��U�&9�HZ�&�!)�N9�q�	\�pI��U�g�<��M�2�Q�ī��>�$kS�ޠs�Z]	aA5}�ؼD���bb*z��̳g�fo��$n��/(8���銽_.�� �2�
�SR�D+/�jܻ��[�
`.��$��!�8
U#�?��ɘ�C`钱9BH�U9�#,��>biyVΘ%�B��A�=��7��,/��睬jd�d��k��ziN*4�'8��B�	53CJ<�QL�Q8Bh��B�p��a�&�ǔ!@%�E#p�p7�]VhF �!��P:Ht�A��u���'U(�q�"ĝ�T��P��/��=�
�;����!г_
�;$勧7�D!W�P�i�lxf :��C#�ԦRu����-�	��J@�'��0�t	��0%������f���N>��ʎ�g��˖늒O���#s�jݡ���Y�3��������$����mB#6R��Ȇ�
BҩR��Na���"�⟔�F=���ߓ+'��Y�Bd�LIqʔ\��9�*@�:�b���@1���?�S��h�PjZ�0�$3��HG+PB��.f�`���9�D(�"B=w7.�䋆Y�x-���iP@���I�2�>O�9;ր����hAحb
A��"OL`Zm؝I�`yn/������>)���^7����ĸԞ� �B�Uc��>gF!�$�|�E���	�X�03��<=!��΁b�lE�Ԅr�"�ґ+��7E!�׾-D�E�P$��>��Թ�X)�!�$��(��ㅤ��2,�P�JרO�!�D�Gf�Aa'R�f|4�܉>�!򤈺�x"�Բh�����i�G�!��>��$�G�}�0U6�!�L=g�ڹ�6�B:dT��	 �V��!��ӁI�4���ê~6Ni�Ě�e�!��6 �^(��j�g�� �6��d�!�����tk��:ٴ1+^��!�d�?^�@�J� �����]�!�d�XW0�1�N���!YP��3�!�݀1�\�"��F���U!�$�,��A�j�2 ��W,�F3!��K�(���x7�	'��H�B�~�!��<!@ �9�bZ5Q�%���֛a!�P�V��Ց$�Y�7��qd J�y	!�� ޕq�E����w/҆ 
��W"OP�A*ֆc�|;���G�|�"O�|���S�bC.Su�C"|4�<C�"O��8����]~��7'��R8B��0"O4I��hA1+*l�������"OP����*l�l ����)>D�����
�=X2Ep��i� �Ά��!�D�?��Q�1�T�d4�x���0�!�ʒ%��� �2!l�C��*�!��H�j vbŕ���1�AN2k�!�$��!dXI� �6��� �Ş]�!�_�/�d���^�P���c�@�<s�!��X/�P���̎P�4US7m�VT!�dƃ,�$p��2R�b�+"��
d3!��ġ����I��[h�0"CD	5!�$O�1�� �C�)W�tDHf��:�!����T
p��R��9����m�!�M�8�̈�քD�8�T�̚$_�!���&NV���.��=�.L��MV�l�!�
|w ��!��?��k�M��
f!�dہo X����E�@��P+�I)l!�d��X�����(tٖ�y��W!��/v��؉�)�\k��a�Ǖ-Z!�*�Z�9��N9�Jd�%�9�!���@���� 
3�d���"�(�!��F�"�K��U�rś�>�!�$�"v*|�8�☟x��=�7���!�$��/L���t���A�rYG�U#N�!�$�/_�0Y�=:��%����!��ۯL�y� $Z� D`b�"�!���!�,ˀ�
�dܹ+$.�+�!�D�n$&���� D����-C�!�ۼ0��9�ĈZ�d�lx���+j!��D"j\�ٱͮv��@Ԃ�.%:!��gɤ�QrDpU­�N֝�!�G�ƨ��E�!�&Q3��|�C��*/��� �O�V��LYH��C�ɠ��8g��h_�4�$��X�&B�	w0v<�ra0}����@k�9�,B�Ig�t��iA�vu�����R��C�	?�NQ����xS�B���%t�C�I/x>T���  �~ȃ��s�bC�I N���t�ѩ`^��"_	:B�O�)����V��w�B�Ia��EOR�S�
�(2b�4s0B�ɤ#��hfH B`�)�Gl�m��C�Ɋ{�B��,��V��A�mK�M	�C�	!�(Q�M^.!��M��ƒ���C��;W�"P�A��}�}�ԁ¹<�C��&'���@#�,?H|sQ'��o��B䉝�"���lE�
�Z��7铩B��B�	�\���fI��=��/�~�fB�Ɋlt�q@���[������,^B�=^>p��s�ܛ^|���4IY/}m<B�	����Ӥ�5޺I���5C��C�	�XzF���l}�숕�T�N9�C��4$(�i�ͿuH��m�$v�C�	�T|��H�!"��ᆪ&^��B�)gޠbeg�aS� W�ވ9)�C�IA� 2���U��$��f��\��B䉿IH�li�n,#`��Ş�`�B�	���ا�'`���ދO��B�X9�0��i�!v"\�E��B�I�V��� �)`��p7��3��B�)� �ZW��<� �3$��m��ti"O$\;�fZj?�AkpVcZ�+�"O�<�š�<�����Գzl��"O*݃�L=4�T��� W�PK"O��_EA�p��#�0��p�K�H�<	d)C���A��؏�t �1 �^�<���P�t�Th0%�ʄ��\�Q�U]�<�Ӭ�6�L�a�Ъs�f	���v�<��'�-m�}Bҧء0����C�q�<�W��.y��&!s����4/�l�<���Jp-h�f#ŀ�H�m�<q�#���xЙSJΕ��@Q�n�<����Ҽmx����H�:�Z��Aj�<���`
��q�6E����`�8C�I;8�$(�.d����+d���@���RV�*�O��JG�P<J����s$�5f�n����'~����,��6R���ɦfdƝ�u�@<l*Ļ��ǎ[޼B�I%07"�#u!ǲ-�4츢E��4�X��b��J�$��A�\i�O#�l`T��d۶��O߇s�HiA�'o�E��h+R�zmY1G��k�n)r&�)�"�U�<���(�gy�jFP�Pݓ�'��(@ �����ybGȻ��02SA�jiVuV��v��S�) 5\ؒ�&5lO�����`�����׸#%<���'1z9��I�HHp�"�i��1[Ȅo ݠ�� ��B	�' Jm� L6�I��IN���p�y�E��}X��T���r��i# Ǫك.� X�n�2��<
p!�D[ <���W菋6-~����*RR�-����x����'�@QE�,O����7_�ɢBN�!�Part"OR�� LARJP����
�0��3Q.E,	�(���I�Ą�	�f�옃1��4H�X+E�	
�����@i��$�Aܹ�?�J�%E�<����`������Wn�<1��.n&�Ca�T�&���n��؈�EhN������c%	�;S�x�
_�T �o3��'<P(�$/]s�ŞɊ@�C b��)a��6F�@�D{����#R��D�4`�bd�HC�
�7e� 5m�D�!N>)�S(����I�K���#GDf�)�E���6m]�Z{�"����$������	U�A��ɇ�3B�n���ɳ�F�:PH	�.؍(s��ViF�i��D�<�J�)��xRh	1)r½@3j�~yB��,h�D�B������G��p>!�ǀPlPqSdKZ�ǈ,&"Q�vm��z�A8_��O�0aU��v�Və��)Y3�(0�C��NNP=Bd��[TqO)�gM��)�ʨ��a���,��VbX�z]��H1c�2�h���J��n ��'$��j�/4�3�D�~�U"���6=�8ҋT}:\��_�Uj�A�3OJ-���>���ӂ<�(Z����S����*��i�2�3� F~���D\�)��q��'[O
���@S@�4��r�ݶ\�dY�5$��~	0O�݊뉁]�t�*O,R�*E.OLDe�D����'N\C���@��=���A#�ua���w�B}��F�)����xR�M'V$����%`�O��|�%R"rvpI9�"樌�H>)�nA 갤�@-62](52w��F� ��tp4爆x���2&��?(�~�:�H(}B��{Z�c?O��pa�Jђ�9�0G�ʰŇ�
�d�ɚ`��s�̊Tp�剄
1#$�	Nlt�v�D~���f�ѲA嶅���'��LJ�#�O���l[�!�(v��61��AY�TĢ��p"QH�D�8��Q{w�$?�&	X�y�D�e M.-x<��֤�tx�L� �,(r,ݺ$��h������X�q�*�MٜO]��ZK�n��'��d��UW�S�'�T�7'Q�Z�1�� &��!�KE|2`��z�U�	յ_��T��e�\rݠҡ�;s!�ĉ�/�V�Jt�5H���A=S���(ԭBF �^Ϧm�'� �g~�N�f�ЕZg'�*�R4�g��>�y�eBڊ�&�9B� ׺iܶH�s�@��ܓ�I��R݅�IKD�h��H'=��3�ڨqh��L�h��M�e'��{��1MO c�pCҠ��{B�cŊ>$�(���J��}ڲ��Bv���,0�f� ���nO�r�<�?�z�c�IJ����ƾ&
p���3D��Xa����%i�%�\�vl�Q��O��Q�ޒW^p�O?=� Z�ag-
�rL�(�c͟0@�ݰ�"O
(Y��m��)y%��	�R9aF�>Y�
�<$����j_(Cc�@>*���2oI�9a~�����@���b��E���w�B:\%�}�'��D�E� l����D�a!�8���$R�!b� XV��~����~��A�Ҋhp`p�!g�<��̕=WTM� ˇ*����(����S�AT��d��>E�d�1ZaHլJ�L�2-�6N"@!�A6��lĴ¼���'�:I�I2�8�v�>�ay�A&)cҹY�H�Yp�=8b���>)2�,�H�B$�����DͺH�0xB�A�B�ɂ(���8��:Y�8ɺ׫ŃXyt�=����.k.V�;�6�S�x�<��kS�|��$�`�%D��g���Uۤ��Q.̕G�PXt��O�h5����LiL�"~�2js��!�L�4�h�e�1�C�I�{YL���)a#��I���˓>�����ǕtXJ��䌑d�ܨ�c�O�^׍�u�a~R��;db�4���ٴ5���1�
���f �f�񤟉'ǜ��f�'<Ƒ�W�,�Q��hR��k>0�DԿHl������17��1�n6D�\#�"���/^Bz��, D�HY�̛�(f��c$�`�bH)�l4D� +G
�&h�ѣ� �|�| �47D�h{��ݭ1(l���<��`���0D��b�E�x�TCI=ʒ���N14����ͮG2�"��^�Ж���n���j��'ZDM��F�	���SZ�5!
˓hZ%U��'��I�c�LĨ�&ہ]M���egB<BJ�B�I}��JV�;(��>4�6��A�>���«o,u"��F�}��Zv�-§5T|���գI�Ƚ��$�H�x�ȓ)능3A�`|pJuI�
Q�|���.غC��)��G T���P%�Fi�g��*��XK�T�� cU�U�TC�t{�	�e�08�\᳁ح�V��"���W���U=���.�XX��A��I�w,��8W��5!��Zag0Oڥ@vc��܊d�����DbC��0=r�ב)\}1c�Ү(�B�IY����2���� De��-U��'���J$]�L�Q��<P�m8��	�>�ݪD��~�,0���8{!��ҙ@�
���?=��=Hm�oF>�)$��\�N̓�ك6�扨���!��W'Q��P�NB�y���"��3d1���(^�)�3�_@n�i��Ijld��_#;�����-��hX�&,O6Kf˸jt�(���W/o��'���yv�î_�(�fB�g���j�X�imP����ϵ^�֔�Ag���x2��;��{���.(�n5{C����(�j=kc�%A��3�8U}\b?S��.��$wB��2p��s� %D�<�Y)�b����@�uݸ!#,���yRj���Jǝ|��I�![򵪇�ܧ�2��!�d�FH�#FD�c����ތi�6�z�	�-$LOf���h߳��-��X<F�i{%"O�	h��B(^�~�ˠ�J5�y��X�er�[�f\%���`g�4�y�(×^������Q*H�0e٢�y�jǺ[��d˂���L,�-�uD��y��0/�)��-B�J�%��HB��yB��~7,@���C��T ���y�k��-�xr1`�F��P��yR�١'�\����+�>Lcᛠ�yrJ�&���W�C���0j�/��yb)���*�&�Ye3���ǆ3�y��%��lw�)Z{\�`ץ.�y�F�<;����GWx�AG��1�yb�֗?���M�05��F�9�y���^�ʸZB,� AJ��y��#�y�Q;�,�9���=���K���yrI
�E"��`�]�J4J����y
� 䤠t�ɜj��x3Ѩ"P�@YC"O��0�ݤ ����/)	��'"OZ�0�L?t��ġ��V�Q��Mڐ"O\���H�Z-���e���0"O\�F [%"N��21�a�c"Ob��ǫ[�gQ����U(bM�5"O��ص�G�P��6J�"���R"Oh"u�LtRdz�ɒ-��0�"O�����x��Fj�<�U"O�P��a��t��'D[e��!�"O ����\ �@�7BFнh�"O:IJ�"��F]@X��C�(M\���v"O���n.2E��k`l�Ix�Z�"O$	�/gA����MU?<ȉ�"O��k����Tb�i �h
�%B6"O(�.8.�B��w����Գ�"OFAh�Axړ��6:u��%"O�D���ɉ��� �O�Z���P�"O����% �Q��عF��@)t"O:��fB�!�b�{J�	�
�"�"O��cb��Ÿ]c�@��h����"O&�zV"[y?��z7�>h��1j�"O,�ڒ����NH�2	���ہ"Oz аJ�M�J�z����\�`�p�"Op�sG�	>$�b�X�Y��y�A"O0����:m�@ŭ3� "O�5ZB���6D��Do^6t�0 $"O�-��M�%��&�RC:4�"O�x����2d���@�O�Q��"O�ѩ�-��e��4A�)�-!T�#�"O 8���S���0(H& Rz7"OXh�2�T:/�D�2e)C7P� �"O�lA$�ќd�yj����.L\9�"O�8���F� *L���O�o��5"Ot�
B��5<��h��x�@�"O�,�k@ &[�l1Ġ��r�8�"OnT��<z���dz�A��"O$0[����kk\�2��>N�Z���"O�QPD�V��l��]B�,��"OP`���ַ!z-�PN�6x��"O>�k#�{*!��F��'�x�'��)�3�?a�bL�.�4;���W�X�3�;�\�/(�<�G<��Iƌed!CR)^4�.8
�b�_1�IJ�(d�x�)ҧW0aU�г3�%Q�"^�D��p】V493!�8}���^�|ң��7���Z�hE�t�Y�吼=��q��<��F�C���>%>��c��g�����z��������Q�*��}��/�u> nF�+h����GX^��B��>I��,?3*�2��x�����f@�QHR="�d���~���(1M�W$#����w���� kq�0=+Bݙ��<yεXPmL2��O�����ʎ����K ^5V%�Q苲hzfe�B�M�#�BS�@�##}*��c>ՠ�� ft�K���m�8,����Yy�r��(�b9��1s�Yk1���)ta�u�'��Gy���%T�2V�7�a��牸i6�T�a/c�"On��(�(��@�91����f��Mղ�:�����O�aCe&2�$Q��ݞ3��}�-\>2��}4j2�$8|e���6H��j��G���|B��͘	; 1�F/�&Y�r�7�ɩ`Ў��C!P3i��i���蟾]��@�$��H���C8O��R�̛���C�	τh�8扡���b>1�ƈ��P�4R�Y�R��`�:D��;�K�6�̑��0�B��Ň8D���W�q~����hB�rZɻ�G5D�h�-LM����,#6�#U�?D���Q鑼&������2�%��!D�$:5Ȟ�;�,iQ�p>��� �9D��B"I6d���!HC�P��c:D�� �
P�+7^��Q��]t<�ȓ]�Z����H�U� �	_Ʈ5�ȓm��RBOM�B9XQ#b	ňiyTl�ȓ}���c�Cz�Wټ\ T"OA�e˃�):صSf�F�uؐh��"O�`���(�j�1�ЉP�<K"Ol�Z�L��:|��0@�b��T9b"O��$� �B]d�/ֆQ�|��"OLЧ*K%o`��PpH�*��PH�"On�:t��/�:)8�'�s���"O��4��rX5��'�%y�Fq�@"O%��NG*��E$0F���"O�퐔�D\y�V��=MV�� "OD(X@K׭L�	���^3�P{`"O��"��$lhu���
��a�f"O��%雀5�6LMTB�hD"OڨP�ZwԴC���(\�YQ�"O�H2�#3��uq`O�X
��"O�}"o�M�֬�&n̾�t��"Oܙ��:t
)�p~���f���y��I�j-��#fP�+H$�#�nU�y��ۭ9��)8BP&%�^ɓU�� �yrfB2[V���.� ��kb`��y�d
�5l���˷j��4#qm@��y򬕽EvP�S"�^"^}R {Њ��y��V��f,#��k�8�i����y��҇6��m��O^,b�Ktퟲ�y����9�@�K���h8����ۗ�y�#[�[��<	"�a}6y��d.�y�g�z	��ʰ��RDV�hrjנ�y��ýw�ك�H�?Kϸ!�a���y2���^�q�$iB/��(#!�A>�yR��4�桀��=�"�
�.���y��`�B��q�}�X�P��0�y�ɯU\����r;<�KЩ�;�yRO(8/�Y���vŃ�Ȗ�y�O�KFb���EѴ��\C�f\��y�o�:ٔ(ȶ�@"���y�I�lq��P�A�2�Ľ�anE�yB��<-�����A6_����1��y"��*yH� K��#]�T8�@��y"GU0i����k\"K���p���y��cA������EpĹ�@ʛ�y2䂙=���(G&��y;7l�y�[�z�!�v��vY@ᚅ P��y��h��=��e@�`�(���L�y� Jm`�,�T.áb��k��ک�y�cBu���*�L_ o;�86!�&�y2�@�<4d�xIE�gdh�pƗ��yBHʻ�M
�iP$x��U��y� Na�(eр�X���I�p옕�yR�0!t���ACzdP�����y��_�L`���>�P ��yB.�6�8t��D�9^���(p�o�<��닮7T-��B�z���$E	a�<��^�}2�I���t����}�<���ٯT<��4��:F�2��Z�<�Ɓ	�`e����- L�
��R�<a3lV�n�z��"��*%�y�<!t�HLF�����34�h �hJw�<����>u���D��E�\`�b�x�<��C��A.P	3%�c<����y�<�Ư���ƥ���%>Q��{�<QJ�;OA��`6iw����Lw�<� �Z�(�D1�5���$"}����"OL�KtDI E,*ez���;.QbD��"O�aQ�`�#8�쭈��ϋY/&�#"O�L)e��R�|�bf��p
j)�'"Op��2/9z=�%�#T�#"O|�cRI�/B�YR.E�~O��"O�{Ã\�_V�L���^�����"O���cFS�g
F-9"*��x�T"OvP2򄃀O:��
�l����b�"O�cC�^*78�m0�M�c����"OkT�@09�����ۛ
�ʑ�"OLui�j��g
���6^�,�"O�9�ۮ`Ңq�Ba�7t��ɒ"O�]��s{du��B��B�b�p"O�T��숼i�(��6���v����"Oȸ�,M���I`@D�"�Z�0v"O ���NN�H!��Ӑ`L�h��Ţ�"O
�+�/�6^oz��`\;\�L�e"O�@I5�W�V���u	�%uM�@�w"O�e8�����A0�Y�GB�h�"O�Ds)3,����ԈW�t76Hh5"O�`d�B����Hګk/R�(�"OJD�O26qH���5;�P30"O��ASe͆]������3"O��Q���(Ҁ{�Hӂ!����"O4H$�>%Ԙ�9q�� @4[�"O,Sdn�8/�2t{�gӜ�ti"O�I@çA9�`@1ᜁVL ���"O��RĊP:z-<� ���0i+0�se"O��N	RЬ�`���@�"O�-aB/DU8��ȡ�C���R"O()YŮZ�'�X��A�B,a:�"O�<豇P�Z]��Z�7J릸�1"O��ե��K�U��:	{ �a"O*e�A�TR�&͛M�6.�Lِ"O�}��ne.D�	;����"OD�{Q�̂L֖;�K̗?��"O��
a\4�hi�C�Ğv����"OJ�0�NF�
�40�]9X��	�"O�`����.6-�)�3f�'s��Z�"Od ���=H��s*@�J��"O*a� �в7!L��6��'�0�a�"O���@N�#��]��)_��p���"O�L{bJ�H�tU(�8G�~a2"O�ACZ<dgB��T��W��{�"O���E.���߹�tZD"O�( �CW]���:bʏ��y�"O4hZ��_2F+Q�ܑ)���"O\d��(IY:�C�+\�vYHe"OD�k���oR�)�½M t(�F"O@�@tk[�N��Pq��m�Ɖ��"Oz@�@\4���A�0	����%"OZ�(e���+��!=}*|Y�"O{��J25ex�x��\A"O���Z}�,Y*GZt=!�"ON@ t!:?���s���!2�P�"O��Ā�gH�t��d߫kBPC"O�1�D��5*֒E"��#r��"O(�G��
��A�,�S9J(b`"O�t��
�t HWa[ ��	G"O4��c�̑,a:Y�Ԁ�A����"O�kr�׳Qz�Sr�d����"O� ��T��bfEG?[����D"O�+�Eےq��i�� N�v�ے"O� �58p�Z�	S�J��ԂZ��s�"O�}�#U/Q��!bDt�pU��"O"�!���
! �F�K��8T�`"O@�˃LTD(��C��H�Rzl5ʰ"OLR���7F�6	�O�h�p�"O-��{
蝉&G�n| P�"Oν����[u��P�K��!�"O�E��叝7s �R��R>,��"O0Y�A@�W�	He
�"P��Lh"O��@U(��iI�Z�ƚ=�l\`'"O����W�W�^H�CE׮Ǻ��g"ON��C���`o��8�G���m��"O���&A�#����c�:]�� ��"O�(��/t~���U�Ͱ_6D�*f"O�q�a��s����*c����"O�*'+�;1UԽ;qj'S~r3"O������S�GK�Rd0��"Ol ���o������ �h֕"Oj� ��!@�P�ǮL
V,C�"O�he듅��MHR��\���"O|0��R�lN����M%I����"O����"V�&X���X</�)P0"O
�%��WƖ��V�.�2 "OPA���9*Rą����*6�"O�8ڣ���gȄ�bdC�	���yE"O�}����gx�=05C�&]:�"ON����r��H�t�W
&�.�q�"O���f�V�`S����F?�R���"O��c����Q��	��6]�2���"O��kt_�V�D-{@�H�ID���"O�����;3�E4��%6RёB"O�i2$�GD�f�:��
>$���"OxAbT��3��݊5*	8"��"Ozh�@O�9%g� kT(�� & }�"O\��1N�&$)i��琶*��X��"OJ����`�h������[6"O4��&��)������-j�ʡ#R"O�E�d���yb BG/�Aʔ"OJ�za�[2.�B�!�7c˺��C"ORM2���!>���!X�,�f���"O��TL�3*6�sw�ǥW�n��"Op]���L�,�,���+AX��q��"O��Bq+�)�B0x�J� %����"O��C�ɨfmDћ�	�C��z�"O8���;��A�JP5���R�"O�t��X�J��� ĢTt�"3�"Odu �� ~�l���+��|[�"O�y���\�*gH[1�[m���Z"O&`���
�&�ʆa
�j=@"O �j��Q����5��b��	;�"O���ϔ�Jɒ����f"O�՚1DX+x%8=�seϊ����"O��H��L�W[��[�D��D���"On�K�@�n����/c� ��"OX!����i4�?�0���CS�<	��
�(���F���t�<�1��-e2��̂��Cʗ7�^C�I0�d�cą~���� �2� C�I57ި{Ud?R�q���[��B�I�(ļ���*Ձ$U �"��Z�F�B�2_�}b�hV>"�'�" /&C䉛ZB�    ��   �  3  v  t  �)  5  U@  qK  �V  b  Ok  �q  Xy  �  ۅ  /�  r�  ��  ��  a�  ��  %�  ��  �  G�  ��  /�  p�  ��  �  ��  <�  ��  � �	 � � 0  �& - R3 ]7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6#\���<4�d5h��'�B�'���'	�'/�'�B�'���$��^] ��/U�Z�3��'m�'�r�'���'K��'r�'cظYA��4Z8�xg&�=�nܳ1�'�r�']�'���'l�'���'��41Cl֝wMƩ���0���4�'��'[��'D��'[b�'���'զ@�R��}�[�&���Ģ��'Z2�'�'���'x��'��'T��s�D
����c̚�	P�'V��'��'2�'��'���'X���EAO91�(��@�{�x=���'+R�'6"�'���'���'�R�'%l$�H^�C

��\�o��ص�'���'@��'���'��'��'��12����4��x�Rk��'n��'�2�'>��'r�'�2�'`P��6�.&M��;�	�:�d2R�'��'���'���'[��'���'��u��Ǎ
���z_��BT垲�?���?Q���?q��?����?���?��O�1^�����*J+Q4	zT#�?���?���?y��?a��?)��?i%��=�61Tg�y����ڟ�?)���?!��?Q��?��Px�V�',rl��~
I�"�m���rR"�U����?a/O1���,�MS�"��#5lQ� A��*���;Մ�!ct<�'�47�4�i>�֟Ђ@0TPq���.UM6E�0��P��-H�\nZT~�=����S���NxP1�u�֓��08)O�1O���<I��	�CV������*rAf-�n	0�m�&Z��b�D����yw���P6n5�
N9Cj� C�oK�/�b�'��d�>�|Re-V+�M��'dl$Pd�Q��H��G�w�̉�'L���ğ z��i>����1n���G^;P��"�'A"(~��~y2�|2�m�:Y� 4�
E3`�Ϗ/<*�i�!��A/��T�O����O ��G}�(��<>:5�Ӂ �E�$Q@���$�O�9FA׻-&1��	1�-&��3�����R+)l�麔��t�����O?�I�n�L�!��A�4�w��Q���I��Ms�,[~��{�����&&�ʥ�C�kxnEҔ��**��Iڟ`�	��ۡ���'��)��?�+W�H�%:^	Q���U�L�p�G�(^t�'��i>��	֟��	˟����~���X1e\�� ������r{D��'J6��U�r���Ob�D*������Uk3> ���h��!����OX�d�O�O1�� Ȧ�f�:U�Ӥ�T<�T�#ݧ� �8敟�t�8O��g�yy���_��'@$@ɦXM�C��']"�'�O�剮�M#Ső��?�ƮZ���@Ж�LK���xǊ��<��i��Op�'���'���C�;�pĨCk_4z�B$�wbӬ~�`0h��i����M��=��ݟ������V�TB�X�1
��v�.� `78���O���O���O���2�S������R+���s�
�$loM�������-�MPEơ��$Aͦ�&��uȇ�[����ʘ�2�X�&�O@�ʟL�i>�@���1�'|]�1E�_N
��!�TF\C�I	�nA�	�	,{�'G�i>U�I�@�IA;|�3� PMiT�M�}���	��'ł7͝�?(���O��d�|����-�L	bm��!���0S[~R��>�������I� 3eTlP�!�&2�؈W��N��R�ûi
�F�<ͧ
�t������1z(CS�^�
	�E�$b�//G�0)��?A��?q�S�'���¦�B���$�@����I����Ĉ�B��\��韈�ٴ��'Fv��?ɲ��U����:\�� �����?��~mc�4��d�9�X`��$oT"gp,�Q$���[��0C	��yRW���������ɟ��I�,�O���m-)�)@�R�Z��0�c�v�R�4��O����O������Iۦ�0-�E�"��;W$Dr�$J?1� �I���'�b>��3F�U��x=��^�;P�̳�n+<,�A͓Ij�1媟�$���'02�'Hy{ �̤;y�x'l�Hy����'+��'��R���ڴrd�����?��rsfq�&kƌD3l���[�iC���r�>����?�N>2��Hڰi�A�Qf���!c~�΃�=��� ��iF��v���'C"��()���� ^�29�yp�i��'0��'kr��՟�����6ly����J �0F����ش+ޕ2)O�Hl�[�ӼSSNQ*�-i��Y�M2�4�Si��<����?���:X���ڴ���� 4hs��� u��b��Q�p�#���� a8�H������O.���O����O���k��7�_SԘ��G�ʌw��ʓZ�F�ʳ*SB�'�r��22~:�: ���tу$�*P�,�'���'�ɧ�O�Az�$]�J���a�C�#���{�"\�w��E�<�ED׃����h��Ny���?�D�8QkQ�l��@��F��	��h�I��cy"�v�b���H�OF�b'̟+���`Tl��O�i�6O��n�X�y�����P��ɟ�Y�?,�J��3�L21��	�C�Aʨo�{~R&eb��jܧ��� |�Rѯ�0,��RE ��;KRJe;O8���O��d�O���O��?�A4랧��dAǃ�^�*lr�Aٟ`��ԟ�8ܴ!��;+O��oO�I3Xe�eK2b�z�z$�D1p�%� �Iԟ��#2�o�}~EV}�	PT��W�|)1��.4���b�^@?�J>�+O���O����O^!���a�h�Cb�"��*P��O �d�<���i,��x#�'��'��S'Cڎu�E�W%�j�e��x�p�E�������Iv�)�0�B�_Kl��������J���K@"?!��4����ߟ�i��|£]>T��h
q��ર�]1�'�B�'����X�й޴tjB ��ZVx��[�(6`�7�B�?y��!�����\b}�'�Q��#� ���-.�ieOÉQ��'u�1ص�ig���d��ן|�]����!	���P��r������D�O��d�O��Ol���|�tMX�b��|��+��@D�x���ץo�#POSb�'[��'��7=�ը它Tg���H>r��j�Oz�$!��i "6�l�x���ī]�Y�_�H�t�Z��U�iD�1��M7��OL��?���^�$�j�	_�RZ�ݚ䈇
�0�����?���?1+O��n��k�lm�Iٟ����VQ��!�p5�	bbC�30��?	!S����ş&����
��
H�cl�4Ry���F�5?I�r3�o��b>�;��'�Τ��:X.�|j@��Kr>q� ��8_�T���Iϟ���r�O��d]1�6l���G�G��ܙFW;,Br.d��@.@2���OڡoZx�Ӽ�p�Ϩ.��*�f�v9���IR�<�����$T&;@6--?i�M�i�.�I�(~b���[�{��e�Sf(Y^
Y�K>�+O����O^���O���OD����G"E7 �h������<AB�i�R�1T�'z�'��y�WH� �&"pKص0��9 u���?Y����S�'G-�TZ��%r��9e*�7@�Ȉ�6�;�y�'�$A�M埘�R�|�]���@<G�.���@�-�4`bu�\ޟt���T����ry�l�.P�p��O�EC� ��;�*�J�,��;P���O�o�E��"��I����	����@�s 
���:.�����@:K<%m�S~2K�
=2 �'��'��#&,��|�����'MJ_���W��<����?	���?����?	��������f#˄^�f9��D ���':�*q�*|�4�<�D�֦�&�|C�dI,E�NlÇ�H{��Ѓ���u�I�P�i>�	2�E�1�'��Y���u�`��'K ����V�e�����>|��'��i>y�����&2��Y�H?*z ���8H���ܟ��'��6\�u�����O�d�|RW�˩N6p)k�b��IrVh� AJ�$+�	����If�)*V���e���I�ć3,�����ڮcEH���EJh��W�� t�|⭛�^]n�XbAI�0{��9뗬���')"�'���T�X:�4#qr����!x�N=�2K�#4@-��-P�������?�2[�X��=n��������Y�GЊg;�]�'�s&�iH���Y_
����O~��'1��X6� 98���х�$4��R�'W�	ן���ݟ�	�<��h��J�7��C�OU�;�hbW!J�a�6-�LI����O2�5�9ObImzޕ�`��:ild��� M�Hw�իU�A��,�IJ�)�S� ��n�<)��N�{�u�N�0;J�	�<���[w���U����4���D�6Q��eR'!�/o� �JuO׮D�\�$�OJ���O˓@��)�?1��?�Emڣ6g�Xk@-�$~�yc �ը��'����?i����]�ԝ����OT�)å�[4b���'�� S���d�F5���ԃ�����'pd��!�)`��Q�Ŵi�H�A6`�O����O����O��}����������v~��a���S�����<'����6R>R�'�>6�/�iޥk%闒��h9�'�8f�zQ�cn�(������	�VZ��nZ]~Zw�z�g�O�~}k>v�b�� �L�@�[+:ɱL>�(O.���O��$�O����Oxd�ł.[F8P��K&Fz����<�³iF2t��'p�'��y��^�3�H\+�#��R nЯf����?Y���S�'oqH�3醉t��`f�ЃOC������2�z��'���i�Ο�`��|�S�L�����(�n����{���;g��џl����L����Fy��yӦ`:��O ���C�9x����U�)�B�O^EmZ`��R������⟼��`BKy��	�)A�2���C�bГ-��m�f~�͇A ,1��\�'���0JɘQi�@�(�%�����@�<��?���?���?!���g�&ṔVb�@O��(�Y�1~"�')"�Ӯ�"!��<	�i�'b�u:���8�����>CtP��|��'#�Ow�h3�i��j����
Zxh�`W;uS05 kѸh*R��G�Iyy�O��'�R��3D�������U��=��ߺ7���'��	*�M�^"�?���?I/�*�ac�M	�hs jY $��ظ5���ˮO���&�)�u�z��a@ۈ��ڗ>]����EĠ<���+O󩞔�?і'��
7f���3�
څ|��"���M����O����O���I�<�`�i ��)��M0s�&!ApF^�B��x��GB��ɳ�Mk��F�>A����D�(|����Y�,�)@Q��O$�$ľ}7�8?�D��$=��i*�� ����e�}*�AR��ٍ����1O2˓�?���?I��?�����iDA��as��qK��
�np��Lmډ"	̱������H��Ow��w��27f��ڪ0Z"��q��hh�'���|����X�v4O�t�� ��r�iI�p����7O)x��Ձ�?Yh!���<Q���?���D�V�%�)l8�h� #��?)��?����𦉣B�T�� ����+c�ߔsP��TE�.w2h�"Ǆ���������	n�Ɉu28�c�a#�����o����	�iB,:�&�XK~����O2���|���RI�C�l��7J��&� *���?���?����h���d�r�(t�� ��pW
�R%�|���ɦegˊ��4�ɉ�M��w���qv�Pe��u·q�B�a�'�R�'������F�����G\'Pj�iǎqʺ�9e�Q�M����o�.8gt�O��|R���?����?a��`��)��ɏ�s
y��������/O^�l+qܲ�������y�':��x��bA�1�KA�[���<ZD���'�R�'dɧ�O�}��(P�S�U���%%/���%����i�O\<�A�
�?��f �Ī<�!
��fY
�9� @�vAz���	�?����?a��?ͧ���ަ��ǄΟ|j�!�7?:<�]P$�0U�@�`b۴��'<���?����?��(W�=���2g�6)�)ȧ��	=�S�4���'6 ��'��O�և��q0$�t)(gGW�)��	ϓ�?���?a��?1����OH�I�e�D�`�g	$̎�*u�'<��'4�6X@����O��nL�I� |�0��X�;8q ��@�b����jy�&`����`��ϼTX�F�R���ʒ�U,\��¯����D�|�_�����������b�Ӫp���8OC�9��8�������IZy"�s�FUJé�O����Ol�'w����V-�7	������J/��=�'�n��?q���S��Mɽ=�
��˽U ^��g��0$ٔ��#�2F���<�'HϘ�IH�IP"M@Aú6u�x�aB�<���	T������)��yy҅b��t�SIB�g�B�ră��*H#��,#�,ʓ�&��D}��'�@����/JaK`���v)R�l���ঝ�'��%a�T�?�i1^�l��G��J�LA���ÚD�����b���'j2�'�b�'���'C哛� �‎�;I��iΠA��h�4	�~ua���?A����O' 7=�Zl�u㉜Yg�U���%MT��JĮ�O��D:��i�#7,6�d�x�SեP�����'=DT�ak{�X�����Mm�.��<�'�?��V4���j��^�$� �.8�?��?)����D	禡��ȟ(��֟�;�m@��TYs��1ꦮZ|���	ߟ���U�	��m� C�ۇ�\6�4�Ӏ�W��M�f��� n?��� ����
�kX�욕��^5����?���?Q���h���N�7�e�b �I�jy�0�p���$�����q�Q쟨�	4�M���w��0sE���o.��)uG��p߲P�'$��'u��	'�F����p˶L��1W�9�pg�
���4@P���4���<1��?9��?i���?��E�|ߚ��pa�1/F�����dJ˦��@ɗ��\�	��L�R��S0�9�&�&C��3�g�I����	\�)�S5lL�����$D�,���œC���Qs��̦��.O
�,̚�~"�|"V��zWG'r#�L�V7.K�5kD�쟰��Ο�	���`y��l��5��F�O�P��ː2��1�JCY����!&�O�m��(C����Iҟ$���C�<\���"�04��f�L/��@m�I~��3�����U�'ſ;���2P��f�v�2	g�D�<	��?���?����?���	�4��`�$��UL�H�/�)���'E��cӬ�+$5�������u$���.�?R�Y����)�b�怈_��ɟ��i>5	�KӦ5�'w8qv��i�:�p$k�8{�����B;�a�	G��'8�i>��	ߟ��I+ig����A4����5��P�.��	��'�67+Bv���OT��|v�Z՚��3X�2��FE~rm�>1��?QH>�O��W���" �뗫P
����Q�qf&�.����4��H�@b�O�!2DҼX{P��&':8�)0i�Ob��O����O1��˓Y�v�Q�S��s5*�{th,���:G��3��'���fӴ����O����@�(���yѲ���ݞ+�J���OƵ���pӀ�2J�}'>�,+�`ڷ�N#1C�%�r��F���	gy��'{��'�2�'Q�T>uY֪̿>��#�i,"w"Q��M{�k�'�?i���?�J~Γ盞w�Ɖ�k���6�����U}H�z��'��|��$�@f �V4O�T��H�I�
��f���k�a�6O ���R�?)��<�$�<ͧ�?9P 4)r�2�[�{&(�#Ì�?1��?�������ĦyJ�������֟�`�R1T;�|:����N�I�4j�N�;��Iџ|�	x�I6B0t�R/�N�D�g��v�,���0(�M�R��tAPE?a��8Mĸʣ� g�b(�&�LQ��?���?9��h�����(��yA�Z	%�X��vN�v3<���Ҧ�B���@�I��M���w�d���'�.���cH5��x��'�2�'7����'ӛ&���rA��&��� x���${��i�B
~��\;��7��<ͧ�?����?)��?wO��*�Ԥz�N�����dP�����ei�����<�I֟�%?-�ɂ2���j��F�%r��d�A&���2�O����O6�O1�44Ȗ/����p��[�S<�
'�7m�ky� �6G�(�����DB�^�t�zp�I��
Ւ�/��N�d�O���Oj�4��|��֠D�rr��&���KDQ;'�ԙ�G&�3u�aiӒ��B�O����O��$G$\Β�K7d�xMʜ+��
(��!�e��t@�������>��]6�6pBW�ܞ����Q�y��I矤���8��Ɵ��	Q�'[y�dB`$�u���ևZ�N\����?a�<s�V��+��	��M�K>I�`��E� �*҈I�.���S������?Q��|² V��M{�O1��S?�$x�G�k��(�]����?A�'���<ͧ�?1��?)[�� ��](�A�y�+��?!*Ot�nZ�x���џ���}�4�� n��ȟ�}�����с���D}�'�b�|ʟ\��H\� j��Cd,0]k"��bk���0��i>���' ��%��BCNؙ"͈�T�=CmJ49օ��0�I՟���ٟb>�'��6��3e�d|�
��RH�([�xiCf�<i��ia�O��'<"��)h��u��^Q����dB�5a���'m��Kt�iP��:v�����O��SXP#�#7.��(��!#�����O���O~�$�O��$�|r� I5;iN�� �dX��Ys�60�f�اu��'`���զ�ݠnnV�7n��Q�&DP@�W�
1j�IM�ŞTi���ߴ�y��Ϧ>?��QeS�n`��4�y��%[d�I\"�'_��ȟh��c�U��`�(��a�$�ȳz�^`��ٟ���ڟ��'.6M7L���$�O����*@��-[�>�.�&N�$�t�X��O*�$�O&�Ot��SIITI1 
2�D��G����bE�5؄s��/�S�5�r���4AR�r��9�D��2cL�j�cܟd��������|D���' ���f�dê��D�#��)��'#7m��D��ʓR�F�4�8�HB�T~�|Z�)O�L�jM)�4Od�$�O���ˤ= �6m)?��a�BE�'�XDA��E��C���� ֎�{��,�$�<!���?i���?i��?a�5D�ё�W�7R&A�į� ��D��]��,矠�	��$?牼���xr�_;B��� �3+i�Yq�O��$�O��O1�r��`�*u�z�6	��Ut�A�L�^Nf�����`
X�%��.o�[y�߮AƖ<��A	��\�%��	}�'^r�'��O��ɻ�MK ����?I #��&B.���٤ tDY��?)�i�O��'��'�c�9A[�)3�˒G�����,U{x�j%�il���T��7�O�q�v�.�����-e���X��&lR��Of�d�O��D�O���+��6P}�T��I�jh�v	şU~`�	���ɤ�M������ĦI&��;�ݘ8�h���>L�Z��N|�	Ο�i>��O̦]�'�N-B�@�!if=x2!�b��AW���I�'�'��i>i��̟d��ks�Ӑ����؂�ɾ��I����'�6mO5`����Oh��|RC�/;���6iG 7�4`��bFT~��>���?�K>�OO�xq��z�8��TÍ*K]@8�Ҥ���t.'|S���|�B��O�M�I>�6�� ��:�@O�o�2�(7E���?���?)��?�|�,O,�o}x�(���ͫ&o\� �D�7?`�������I��M����>������D+� �HVM+�,���?����M��O�)��	W��TT�*lB�K^.�$8�	�oM�Ģ<����?����?���?�+�V�Y��D�W@% ^!`7cԦ�Y��T����蟼$?��ɂ�MϻV;�Q(��TE�|`#��h���?�O>�|BTA���Mӟ'�tk�A�=!D&��''Y�3��:�'�Dݟ�8��|�T����T�E#ݭkzA{T
޶i�v��d��������H��Oyb��O���':r�'JlQk���?m�X�(� �P81@����g}��'d��|"��J@p4b0)�=i��b#��.��$R�S�6i�"�G�X01�m���]0��D�}Ԯ$ &���X����E
Rp��O�d�On��#�'�?Y���F��)�b�.L�ǃ9�?aֹiM�q�U�<Cٴ���yF%H�j�$wn����е�yR�'���'K l���i�����z�8Dݟj�kR��n�Z�@�Ҭ4�p(R�&�Ĳ<�'�?���?���?9��ai���˵|-� PԈ���Kئ5H� ��(���t$?牽=�\ Pv��
��
�6y�H��O(���O$�O1�rF��7:z�0��ˢP(�4��1{Z��)��<��c� z����<�����}QR-"�N.a⒩{��DU�&���O���O�4�"��:�$�Z�R�8�J a�t��E��Lܜ*^ u*�S���D D}"�'��I:!����˯1�qS�L�8�!�N��]�'	0�4��?��r����w&&���ƀ�de�uf�+r�UH�'��'0��'q�'��j�Kdg�&rT\�c�̚y8���O��$�O^DmZ�y�����8��4��M茜�Raȃ)��9Bc) �j�L>A��?�'����4��d:4�� 0l"rK@�E�	JA�	0DCP�s!o���~b�|rQ��ݟ��	˟�#�.��<�X\a҄	�����������Qy�hu�d��h�O���O�˧K�H갉��k���b�N�	�"��'����?I����S�g�&�2�c�曟f�l����!r&i��X���9�O�ɟ1�?�s�?�D&�ȶ�+@�T�ڥ��-q2����O~�$�O���<��i��D��7t/b\³�ҽ?��]Z�nY*@&��4�M�r�>I��{��5H�GC�X:v�Cmě�Ι����?!�P��M+�O��QR���JI?�cQD�?���3R�A�	uTS�mb�T�'X��'���'��'��� e� B7͂�{�<٠S��.#�.���4Hh]����?���䧘?�P��yWl�m#�q2R/�H�� l���2�'�ɧ�O0�BR�i��$��}͠�b��I� Y7�;[l�$),�� q��psz�O���|���8�Р�@�@��mS׆#��51���?����?�*OF�l�)0ߴE��֟��I�x�� F���M��Hd#��G^���?��X����h�a������=�h��䇝Q�j��'z���2���:�4�������ߟ�7�'/z�(�B��j��<k���G������'d�'���'g�>��I���"�78�t@ QJ�3�0���?�M��O����̦��?ͻ+1����'
r��I�(@�-4xd��?!���?I2�<�M��O^)���I����қ4�V5"4-x ���CG�(�O��|R��?���?��!�T[�L� F�ɉ�J�S
�(O��lZ)V���������c�S���{�e��
-asH�?�h 0To���d�O��D!��)�(Dʵ��b��O|U�eD�;.�� ��S�X�ʓ)Z���b�Ov��H>�*Op���B�|�XЉ����`@�O����O��$�O�)�<y$�iE�-9��'r��nH6 J�9B�E-$��� �'O�6M%�ɺ����O,��O�����U�B8Rs���1C��Rd�6m&?)n��g-��|2��q�ֵ"f�*dK�Q�V*�M�Iϓ�?����?���?�����Oۊ� ��D8&7�d���
������'���'�D6mA�N���$�M;L>i�OW7^
���c(V�1���ԋ�r̓�?�)ORY�rJa���uc�@�?g\F@�!eF��҈h�.�q���������Od���O�����s2�p�ˍ�~Bf)�Al�J���fT�hi۴:�<�9��?�����)�0e�l(�"�#f4f<J��$l��I�����OR��/��~j@�ȫS�MGM�!�$���$�<H���IB+O�2�~�|�.ȉ&`�ERv�C��f(������'�B�'<���[����4SVL�a�Õx�*�:SF��.]�o�$�?��d&�f��MI}"�'����[,.*<��i��o�P �7X�li����U�'�]�B��?��^��p䟏�����	4���ԋ`��'%B�'���'
B�'�S�o���q2���T�ܨ���Nr*�(ߴbJ�0s���?9���'�?q���y���!Q6�(���?.���L��;�b�'.ɧ�O�8Daһi��$���)�(L�Q$���@jJYS�Ȟ�� �	�4�O�ʓ�?	��8�aC�-o���k$��D�ʁi���?���?i-O28lZ0y6���	럄�I�/�TDh�̓�}](G�֯�P��?��S�D����&���6I�<Sfj5������".?a4�O=Oe�eڀ�n�'Hd��D���?a��o�ZA�Q<3�h���[��?)���?���?���i�O.��Q���j����ӌ�2g�౹���O��m�b$�ݖ'��7�-�iޅ��Ó	*�$5���-Is0� Mo���I�����gԒxnU~�KRL?BL��N.\K��;�x��W
.�e�L>�/O���O`��O��D�OT�IfM�v�Dl5	 �!�)�3��<Q�i :x(��'<��'!��y�%��3tAiC N�C��S�	՟g����?����ŞN�lI���(�h�(�BX%:��@[Ѡ�y�X5�'v�݀��柘j�|�S��"�A��dTb�O�g:�mb���柄�I��������Xy���j<q'�'���D�P�K9Ȕ�0dr�@�'7�'�	���D�O$��O�0"�ЍQ�<�D��-�0�C]?X�6�9?y��ON.���E����c%�6j��@�f�u�f�h��ɟt���4��������J'td�Bw�_�fЈ��^/�?����?Iõi��T�O?f�ڒO�`9�(�>\��zd��!S�ԁЩ)���O��4�4��h�8�Ӻ��Ȍ?	xA$�\vm�=bB�/�����A^�O����'"�t��!)_Le[�	Խ:1����$�ɉ�Yyr�'<��>�x�1�ۇew��QA��v�J�]��	П��	w�)���i�N!�b����BͻCc�$<���H��;m� �+O��6�?a�'�$��Ь����Q(�,��m$n!�$���9��@<<E\�	Ё�$Bִ���Ø�am
ԗ';7m-��'����O����["$r�"!/�]]ԥ���O���Uq��7�2?�;	Z���X]D�;�.P@��V�@2"�f;$<���D(|OB�ѷ3Z,�8 �I���3k	ަy�&`�dy��'���lz��A7�U�n�`�)��"��5�����t�I]�)�S5t�J!n�<� %:'��j�t��e͏�y�>HB8O�q{�jE��?�'�:�ĥ<�.O��ӉT��d��� �~��z��'�6-R@Y���O
����1#de8!�uB
8y� � 8�⟐گO��$�O�O ���P�d�d�����ʬp����噪v��oZ���]:����t��>(�rHXD�jU��k;D�( %�5+�S/p��d2�����ڴZą����?q5�i �O�ӣ5�d�y�����˒��(x��D�O����O��S�c��F�2� #��?]�&W' �k��T0	�D�c
�G��py��ɍU^Z���E����+2E����F�"����z�Za��XU��Q�c1�B�eB��؟���K�)�S�T��+��iڜ[�LF�)b8��$�CԐ�'���`���ӟ$QӞ|�Q��B���[��Y�n��f�l��*���؟�����Ly��~��u��O*(�A�7"ly�V
/'�$a�E��O`|oo�J��	�����ǟ���ό�sG��&S
�� �ޤ7"�<l�d~B�3{��G�$�w1�8��Z�0l���9~q�y�':b�'���'r�'�����%n�Y�gޠ�x���O���Ox�n��b��'��6m7���n�0E㈑ei����ǝg@��O����O�	�U�6m4?��k^� ��0R��^*����^�VC Hx���T%�8���4�'�r�'���3�?0zڴZV�J�4����':�T����4w�������?����iǤX���P�ߥZ��$��9��	���O��$.��?)��".H,� ��+�!B�ϲ8Q���L����D'Hk?	M>ieR|��Q!��~t�-@��X�?q���?��?�|�.OJ�mڸ)E&EY�+'�ҍI�AZ�P���%A�Ty�Le�~㟠I�O���1�����7+�tK�!��:}<�d�O���u�pӢ�E�~lЭ*�S�C\����Ԏ2ܹCש�"c)��IIy��'�r�'
��'��[>����зZK������cf�iaf����M����?i���?aM~z�ϛ�w�B��6Z*E��=�5K2
�k��'s�|����8- �v2O�����"~f� t
G�@�<�>Oh)��W��~��|�[��S֟��S��a8V`�!���gq�1s���<��럤��^yr ��`+�O�O����O�@�1O-|B"@� T�4ܺH[4)�I����O��$5��߰,m.�P���+[S���í��`����W�� �B.�⦱�|r�弟��	�!�b�!
�O�HHCǫ�'���I������D�	P�O�#W�6� P͖'s���5�B�8k�)d�hI��O����˦E�?ͻ������!��)����'-�&���?��?�ԦG�Mk�O"։�*� ��!{J`�U�%,�y�r��(K��&�|�����'���'���'QXI q�?`$}����h�i�PQ�,A�4�A���?a�����< ���H\�7N-8xH�(�Ss��ߟ��IK�)擂3+r}g(ʴ?tx��b�։>�Fp�5��Ӧm�'&��1�X�40�G*A dLB� �d�'��ex��иhT ��A�S��Ts�FJ XU�A� ;h����ׯ3p� 6��5���T�	�8�a3 
�l�ː�w ����D�=\ RU���_4�����@�(�cE�V� #�Ay��G�\X�?!�摋s���Tp�ɂK� ������!�S�J9�v�w��!�qJ���5��DPS��x���$�K���	�V#)������>G�D:��;J�1���R�'j�W��,�A�tcxӴTb���>f�5r%ЯVg�`:F!զ��' "�|��'���w��U�4,����ՙl� �g�%1��	���I����'P|L9�~:�4|�3�&ِ4� ����5;\�Һi��|�'�C��qOv��L��V��@V��+Τ����i|2�'��ɛt��}����$�O^��B08=�bM�.K=��`U`Ұ	�f4&�T����#�΍g����˒{��` �㇀E�!)D���MS*O���W/��m��ӟd���?�)�Ok�O�f���s� ������V���'q��x�җ|����:?xEQ�ΰ!��p���:>�F(ɐ(�l6��Of���O��iFM}bS���ԩ>��$˓�۸7�$���@2�M;��
���'�����Qy��}肫ߵi[X�qA�itT�n����I�P����8����<����~b�H�,U��a�#e
)b!MH,��'�.4
S�|r�'�2�' ��=X8\
��f�BEKB�p�6�<a��'��I���&�֘���豢��W*�@$�(*��(]�J>����?������Ņp.L1��nK�ú����*6�>�����s}�]�x�IS�I�|��e?��ǔI���lLPjf����IH�I��x��ݟܔ'��U�A(~>i��-��f�h97L�N"���$~Ӳ��?	H>q���?ɂ-�~rf�'F߂�c*���d�c����d�O����O�˓q��1�S?��'F�)��jç
�N��$��*�^��ٴ�?�M>��?�DL#��'��=4��<	jLBf�%�����4�?����Ѓ�N�O�R�'���_E�<H)�H%v��O,���O:�r�e+�	g�B��4��aۦN�?/�D�Ģ����'r���Ohӎ�$�O��D�nէ5V䄤8�.���FC�Ͳ�g�M����?�(4��'q�� ��g��5B�N��F�I����@�i`���s�
���O<���*m�'���1c�ޕ�@,E.@��i��猝<�l��ߴ���������O�bmC0x���	P%T�l4X���D.<��7�O����OP8���y}BU�4��G?�#�M�v2�a/nLH,+aFܦ�$��yw��ħ�?���?q�l���L;Q���/j\C��XD���'����u+-�4�>��6�����e#��|�W�L�T��$����R��ǟ �'���)�Q ��xhڹ�^�F���Z�P����Ɵ��?����~��\Nt�B���9y#f�I�C�M{f$VQ~��',��'��ɴaf�k�OV�ٳj_
8�RG� 5-�X��OP�d�O�OR��|��� {^q��M�G�����֪O�p��xR�'#��\JUT���'�xD��Q�~f!��ʙ�r���f�n�b�\�	ly%F�ēy�ڕʱƖ�HQt;��H���m��ؗ'F2nH=u��ȟ,���?��qR��k$ȉ��]6�š]�O �D�<i��\��u�E)Jr�-q�����,�L�h��'d�Ad,B�'�2�'��R�֝��L�����1+mJ��w%}Z�6��O��T�DxJ|�'��c� e��<�����٦�R@̎�M����?a���f�x�OL֤����#�J�R%�=���"k�v��O��5��?�9"L�DY��a��Đ�2�i���'5r&��^�)2I��!O��R��H��p���9N��O<t&>9����h��<�8�[b�.;!4��*�w-�D�ܴ�?��@�rى���'��'� �e��:�|m���Z�+��0�$�O��O��$�<��oAp8Ef�
ں9A'��w�����ǣ��D�O��$'�	�����\�6И��_�g�x��ɂ�m�e�bc����ky��'4� @ܟt�`�Q��ҕ�Y�w3��s�i���~���?�/O:�*6�iz�͓��*��J֫jdX�O<!����D�Oh�@a�|b��{2R�9e��+A
����,/���D�i��O&��<�Ee�S�ɏ7b\�����V���X��&b&6�O���<ٖ�E-�O�2��56É�7>a�a#[rt��3�oӯ�����O�d.�9O�N@�B��)j֣��~ʜ�J!����	�;�dٟ����$�I�?���u�͜�2m�@J�_� ��d�X�M����$�9��ݙ�ɀ;T/�9Б�*vfT9'�i�0�x�e����O��D��0��'T��*LL����#F�M�L$�.�)�b1ݴoh\��?a���?����'�� (�D#��h�)Ձq��隗`t�����O8�d�;@���'��ꟈ�P.��
� Xn�Jɪ��� /��en��� ������7�}��'�?i���?�V��<���")#B�dQh�M�,u����'\"�h��>/Oz��<��s��X�-Ԍ�{GۡAl|5���^}ң_�y��'���'^>�ɯH0�)W�v����0���I�# ��Ĭ<!������OZ���Ob5ibfM.q�P8�ƞw1��lW/@r���Oj���OH�D�O�ʓq���;�� P5������珵9H��r�i���ן��'���'^BM��yj��I���Vl~g-ۦ��%/k7�O����Ol�D�<�EE�G���؟�X �, h���W�L N6-�O"˓�?	��?!t!\�<)(���չx�6�aTO�O�^a{��U��M��?*OH����|���'���O��yc惛�f۶	��͗-�]j�΢>����?	��y �,���9O��3"�9�V��=Q�B��j�*(6ͻ<��)I2��V�'�B�'���i�>��H�)9��C�
�Bmj�'G��p�o���x�I�V#(�N�hܧ{>B�IE
� pW�ɳ�j����l84�J1 ش�?���?��'z��Zy�	?&p�Cd㗗,��u#�P6�I2��$�Oj�D�O��?=�I�x|�(s��R�x�l�)��3&|@�4�?���?�`&��s�IMy2�'����
F.���2iΜP��X�sQ�֘|�Kʚ�yʟ0�D�O���m�ԕ#gB��i�B2$IJtp�6��O|@#��h}�W�|��Sy���5��P�K�Hɐ%a�*4��%�1녷���S�X{���O���Ov���O�˓@�p�W�B�J�2�`�U<P�0�jG���	Qy��'�Iџ���ޟ��dR�,� 1�H�!�}�ФF�D�	ӟL���p�Iޟ4�'� �a�q>=h#k�	 ��A�g4�p�t˓�?9)Ov��O�d�}��	'@ёF��$=(���2����?���?�.O؀�0 ]d��P�ڼ���A"9[��9��͌gv����4�?�L>9���?a����?�I������k�P���+svI �Gq����Ovʓ{��Xq��$�'�����-D�`!��9�NQ�玓��6O���O�Q��(��`B����j�H�zʠr�����������Z���I�~����j����9QƔ�@/����U�!NP�lb�����O�p�t3O��O��>M�%���FDq0�'��i��PX"�~�>�Ũ_��I�X���?M<��ޚℭ��,^��)�e��Xf��!��i�8����'��'��B�$6Y=�i�e����s�"��vD(Pl�џ����ĊS���ē�?����~R�0r>%@s*�t6�*5
���MN>���OU��'"�� PAl��� 8�ڿcJ��ði�N���O���O�Ok1&�6��v���`ێ�j�$ �E�ɋ4*<�{y��' R�'��	+}"�C��Gv(�Xk��9!�rMa���ē�?������?��#W�#���-�Đ�Sc|�X�c�L&�?!)O����O8���<��O�=b��i��w�D�@g�
V#t�vڭZ��I��4��q�	��0�	�����:elʀ�G�2n���S,_j�Y�O����Oh�Ĩ<Q��V#w�O�꼮@ǒ�I��BL�s�!ȟ�f�'��'0r�'Y���'h�=Z:�iSa�]��ا"^k`t�o�� �	vyҎ�-u���������o��f�%���'��]c�KUb��㟐��Ob��	a��j��l϶7nj`���u<(�X5iۦ�'����d�P��O4��O&F�vN�Jȝ�F���G��f �Im�ɟ���a5t���y�	{ܧ_"����j�"�s�küO� m�)c�e�I�@��ן���ҟ���F�t�V�Zlq�U#B�e��
��/�6-�k��dE�EѦ�
����YD�B�Io/�� ��/D���á+R�%����l˰% v-�OvS��O�9f����p���
�'$p/*�YC�T�:�`拙�zJJ��6!��/0	a��l��)Jg%.d�����_�*Eh�#��%S4��L��D����D9xe2�"�'G�P�<H�5dMm$㖤�+kJ��eN��P t5�0�.W�mp�^�\�>9ѕ�\3�|9B�'�"�'��m��#�R�'��	ۀf�1;��ݎQ��8���dZj埅Q����'�#]���G�{�'��\�FƈO�(0�ʃ�����_�!�D����s���8���K� #?Q
 şT�� ��s�R���%A���.0�E{��5O<�)��چgΜÄ�	(F�B�	�K8��卅4^hf�b��Ԯ2ȼ�"���<�SJ�E��I����OF���w� r��DjΒx���9b�Ֆz"�'�R���/�ը�G9MZ���O�ӎ6��:�A%[a���
�J�T�<!6ϋ:X�D�CF�k(`�I|�2Þ*$���HS�I�'@ڶ�E�'�&X���?ي�$N������B�s�^<w���y��'N���T�5L�p{��K�b�n��z��'"��x�m�Nx���3Ǌ#X�:!��'�f�ȔG�>����ɕ�=c2�'B2�><��	$�3#�mp� ps�]b�΃�P,2Pqa�4��T>�|���������S��x�`��X��"�� y��]�	�.<.ٰ�S��?�a�w�@QQ��Ǒ��t[3[�faz��?��O�O(�'�b�k�]$�B�;
���Y��'�����oI�M�E(�����T�����f�����0�"�@H0�$�ip`�#z"���O�ppf
 �z8�$�O����O�կ;�?���79�!����<?������ZHx� P��mFI�`�#��M���|F|rB_*3��Z+� b+��-@�>H8�����/A�&u����R����O����/�x̓(<S�gO�
Nt4�e�G�.h)������@Y�lu�0���O����O��4�<} 0Γ�/؈+��Z#
�
q"��I�HO��0�t
a��0#1T�Yvբw���4o#��|b��~��y�;M����H����Q4�ٜ�R��ȓc- ��rlWhb�As�̱1�fl��Gǖ08Gʗ�R��!�D(IZL��B=���%�L�Y���M��@��<�,���gN������O�&��ȓr��١��D4EI��;:?�,�ȓ3$�(2���x2(Lbfb� 3�P���\�.Mȶ��.�v����y]���?#��q��ר^)�t�� ������A�й�LZ�f�y�"�9(y�ȓ:R�ͫ` K!V��Ƞ�Q*⨅�b�ܸ01.K�^���H%H.���@Rqqa���`vfG����ȓ�P� �
�2�^T�W
Nv��<��k�La�עȫ"fn$�p�L�N����=�Ze[�,�&��I�%
�a�ʀ�ȓ.͌����z�8���N�H�q�ȓa��p$Ν$\�*@y���ҙ�ȓ5����F�ۜ3ThꐁX�Rt8���V����dcD�G�b����	-c�@]�ȓZu����jĶ) �$&0|��ȓ_�:�bR�"m��ͫ��!l�E��O��H�������) �R�J���U��t{p˓&Z�!R��(��!��S�? *a�A�;0�1�,�:q�"Or`��+*�h�6�O�B�,��"O���⇘9D�
5)�3C��p%"O~բ��BVh@�״f)��r"O���dʺfj �Uȃb%�"O|�b'�ъ=QYQ���%����"O&��'/���d��F�YS�"O!�5���	�.i�6�߭�R�:�"O�hp��^;�|�� C		8�5�Q"O��D)�x}r���Y8?TBQ��"OTX�G]ׂ� @<N24Ӂ"Oڑ�+=~�P�Pn�@<�Z�"O8Ա�Μ	��ИE���/4��"O�c�)G�;�Z�� ̒K�t�"O���BM>���ն
�<��"O�PZ�nפ^�y�����`"O<Ѧ�I?\����&\�tCc"O����,�	~�Μ���ҳn_.�0"O Y��"%p�	�,�z2��Z�<I��1y\2H�����:��XcaH�y�<��+,p�`̊��~��R�s�<I��2��Q2��Πz��H��e�<� �J�J��P��~²QQ���a�<i�O��NTݩ�ʟ�~���!7#�d�<�т \� ���dT�$4֑����d�<r��=̩�F��f�P��_�<�%'T7��L[Nɤ|
^!cuJ\�<�o>��},����BǑ&����p� �i��Do��y���U��'���Z� ߺ��Qa�q3t��T�|DS�d��A����~�Ā�ȓTД�[��Ovꊑ���S��	�ȓ
X�C�Յ�^5��aG���ȓX��:��
8��L��%܅ȓd*�աT�ɯJ* 0f�^)j�ȓe�h���-����g�E	����O��XP攟9w(��FX�\�hͅȓAQ������:��K�1sx��ȓߪ��� >b
r)�sC�i����ȓe����U�ʇv�j�
�'�v�T��qCX+��״t+N8$t�"ل�^N �k�l�j�X��
�2!�vh�ȓ,�vD h	�c��0t�-����ȓkfZ}K"N[+	h���^�<�ȓe��	2�S�X�*�3�N���n���`\����/h-d��e�W�q�����s6Ȕ�/��tA4�[�7�(��ȓ��� d��khDq4K��`h��"J��s�#lC�0c�7Enp�ȓV���+��X1����.Ѫ9 }�ȓ	��e��'n���%�Y&c�$������YS�� ���ԡ] ~l���P~�L@��-,`��萨C6cN�D��?�:,�l�،x��2kxF}�ȓc.^)���@�����,՞��ȓGx�8n�=�Q"��"	�����qWk�9K���֠U	�2)�ȓl�0��剎��l���'�K��0�ȓ?G�Pb�J�q��
Ph��o.|݆ʓ�`�deO�i�(�r+�.%� B�I9M��+%kT>xqtp���;(��C�I}�j�k'o�o|kVi�{,C�	�~Q�lA�����#0�ե�C�I,w���wB�;?v9j�K�8R�C�)� Rm�ϝu�"��B6ӠtP"O�Z�,�-���F�Π���Zt�'>�q���­��
�48&�&a\$�v��d^9R�!�:M+V9#�G�ws���ℏ6�qO�`J��FH �?����('GЍZ���1I�H',0D�L#6�(5�ެq���������6f{0��<�;�gy�*U�md�����xYPwm§�y⮓ z�A�&HV1�֬�V�*)ৡN e�}�Oߊh�^4 S�~��SFl
3�p=���ެcτ1�'֞V̖4F�uJ'(��=^=�c!?D�؋g.��3:�<�F(N�y0��C<�ɾ���a��?�'wi�ԉ�jm�>`c�(]	G\Y��&D�>�	;irI���R;&�K&$ K�� �T?T@a5c3�	��II0^��P=#�k-���9��M��|�;2�M�W�B�I�VHB@sa��I�X�;�i" x�'��j��6�@�J�Y((���|��B�;h<����ӍLR١�M�<���ɼN��Zu���HD�`�=Ξ�9��W�,�]ɖ��|�<)�e'A����)�R�:0(rBK<)�i�.͂��P��69T��gJ��Y�ص�T �j}��*K�=&�����f���h@'	�!l�{�
��1�ax��\3Z���gǙ3����Cm�Bm�U�Q&�}�n}ˠ�٭SH���'�|h�!יc���ۇ�ݣGp֔+�Oܴб	�'O`�j�&�=- �8���[vvM�РD�D���PG�A|!�FUz�����ƺx��ёjY�f��E#k�Il��S��(}iTi@��$N���" �V�<SlH�oD	�!�$V�u�4��TB�v�����+D�z�1�J�	+���)1&�;B��ۓ1�Wa��,.�I� ^x����$��jÄdr�P:dq��Q3G�8J
�qr@ž|�ڴ���V�w �A�"O�tZB�@#6�����]8,��u2����;�Ǎ��\��bO���j��S�y��$��GÆSDl����x�>٧ON�NsQ>Y���*wpL�C�`��~4�j$ܡe��p�T4��i�1M�V�Bb>� m�/����l �V����Op\�H�7㸧���0��+��	QDD�&��*���#��qĀ�0��k� 1lOУ���t]<yƪф!��L�f�>9r�T�K���̶5�~���tq��:��
%;�~��O4��¦�v�z�!�1��\�P�~�<����9���.�Y��a�Sz�'�ܩD�-§g9��@gݹa�@M&{�=�ȓ9�RXjVƄ�<}�`#�(����� ��l�rD5~Rt*�)�s@��ȓPp<]�Bk��� ".-����|E��ʦ�A�i| ؐ N��E.L���rfvaH7�(du(����B.�l��ȓV޼���	�n�,ؗ��
3L��ȓiH�
V$�;]�4�j8Ԩ�ȓj�� Q�B	�xduj\�$�-�ȓ(T$d{#��wB�h�.��Ő�ȓ����(E�'�F98c�n�6�ȓ-���C�V�l�"��L�Ao�y��{��2̑���Y�F݄��\��>؆Yy��Vi��Yj�?M�����3�����B�8s���;Zv�ц�#�B����\ ���5�Y����8��8���O�ѐ�FĜ=����ȓn�n��f$|���E��F�֔�� �����8Xx�M�����vR(|��<����-�u��kK!:E�ȓ	Kf�h��%4:֤k�,���ȅȓ=_�}{�U�?m�����J�H^���ȓ_t�1gOJ(:NH:G�W�"�,�ȓ&�A�Z�a4�	ZQ��=NބP��(~`p&�L\�J$	�R] ���W��� X@� 	 ��0��)��L&��p�XHDSУ�6bɄ�S�? �2bm) � �懰pX8�B�"Oڐ�#@�)�h�ȅcH�1���@"O>� ���O4bL)�ʪ/�Yr"O܉���L�+���1�/���Rt"O�)1`Ə����c��ј��L�"OL%��Ӓ%��-B���\�^H%"O&젲�΂Z�HhȠ�B�J���+0"O|���1G^1����/WxD`6"O~�J&E,p��mЀW<����"O��*�әo�P�P�6.!�A�"OX���Z�vD�7'�*f ;�"O��P�)D�ȅ �CM5��*�"OhH؁�¥*7�]�c�:rSbeR"O*}&�ۣr>�a���CJ�ib"O�	�T�p��Å"�\��:�"O��2T�$6���� ��V���4"O�T���\93�poÚv=�l�"O��c��L�kX,�i�Z<��mCa"O8h���8�����N��5�j��@"OBU�� �!W��+�"`֗?�yr$P�wþ9���$)���� !�|��NLRH҇�P{��U�4-�6�x��H�p,�E@� J.�=� �e�r�ȓ.9���F �$Y2�f؃Tk�4�ȓQi��RF�t�l�8 �PV�݅�i����ƌׅ[Ȫ�{�N'V�ȓj~N�K�--*�A���Ů9���ȓJc&%#��BG�{ͤͲ�F�S�<!v�Ǟ_�|)���,E��) �[M�<����U�T�3�P�)a�[S�<�R�\�,�T|�싊�h����e�<�6ˉ�3�����j$�`qb��]�<Q!@��RQ��șo��0�MZ�<�"/�$/��1C ��;o��� 4Ʌ|�<QF�'A<nt'!�5�Xx�1�Gb�<�!�i�~pІ��O�5x���]�<��P�eԊlH`Bm�ȫ�5T���0c�4�� )��"`/����*D��b���_:��Q��7~u�-��m.D�CP�X�-��4Jg�i`t	�0�*D�0R��	3:��y8�Zr�8�C�b-D��B�ލXX�l8!gra(�3F)D��fg]<Ԥ䳒%��VYfL�a�%D���̍�NNހ���@�n�`Hv(.D��a��F�����&�7�r�w�>D�P*$P4l�}�����Rt Ǐ)D�L�Ħ����J���4U��ѡ(D�H��8� m)��ԔQ^��2�2D���D��=.���Ff'{��5<D�P2!J���۴��?j]0?D�(Sf��$�ƭ ��YE<��ڔ
 D��R�L&R`��Z4n��9�|���1D���eh�]��h# �,\4���'0D��d@4j/~i� ��
g� �a�3D��p�,E9�h�X�A�E��	�b�#D��@� �<
L�	�;�ܡ��6D�tɱǎ!��Q�%�Q0E�l�s��5D�ػ�& �?4�$R��9F4쉰n8D��qw�Ɏ|�]�$#M[.`Ao7D�Ȓ��G  ��1֋
1֕6j4D�D�q�Ohw`��$��4a\��X&�0D���ׇ1�T}S`Ȭx���I3d9D���1I�$dy�r冄>.��� ,D���Z-j� 8���z�<�6�6D�� �@�v*�(fK�)�$B]i��4�"O�:;�D!�@ݢY��b"OL kO&�B �t��,��"O��Hdg��[�t�͗�?��R%"O�8У��0U���̦h��H�"O�DQq����Ex�oʪ�M��"O6+&b�v�Fl�3��'}K4"O���ղ*4�j���`L��!g��p�<Iaj@�/2�I!3�$z��)X��A�<�g�.m:���"�s`�5�d��A�<�
�5��\"7`�;6�{�F[b�<BªIE�U
�F�AO(��gG�<Q`���� (��5P޵��'�E�<鶈�  =��P�3g��BӀ@�<i�l�dD�Yb���Ft���T�<����i��k�
�/'�p���e�<�$�B�X��}.c��a�pMX�<1Eb�]�>�xP$�0a��c�n�<�'�M�����@ܒ��pi�gMC�<�&fX� �f�@�5�,�P�[i�<�!� H� �&/�;o��`lN�<9����pH`\�^Ԅ]�G
d�<Y���#ZXBA�c��.$��7�Yi�<U���a4�4�`+�WX ��B�I�<�C��]I XRhι&8��hSN�<�7&<^fF9ba�0o:������u�<�w�i�.����\d�=Q�KXt�<�����'Ӑ�A�?(�1yBb�D�<����<}A���e_�0i��X�Hv�<�S/�&2��ꂫ� ("�X3eY�<�$�D��$�D�.��T`�D�_�<p!]2��A��&ҡFCz��F�d�<��b� ��E�a���[lމ�b-]w�<�g���,��EM�A���ТJIr�<)4�OV]�)��	A5s�|�P��W�<��k,���5�VSD��*�N�<ǫ��mU�u���Q�<�Z��El	V�<���Q� ���+�O���˕+�N�<q�(��C�g�'$O���1�A�<�d�2�x�Y�%Q�|0A���R�<������=�f�}�䰦A^F�<��_�|êp�"*� �`�z�<ѵ�J=N꘴����*��(���w�<��_�qXU&�"Թ�@�s�<E�-D������ 2c̭���_s�<9 B�2��X@@���9h�I�j^p�<!��K�Q �KR�����D�m�<���1l�����8C��h�<���K�f���h���%~�i��}�<1�Ò�V?�����9������Aw�<a�$�:I܈�"Sh8o���jbh z�<��K�#dzA�/�>="H
c��y�<�ù"v�q&��j����wϕA�<@ O�?�|I����-i��{WM-T�*�
�	g�T�1�I�U���X�;D���l�E�p=)1┉�~mp�J;T��S�,
<9��ʤK�����B"O�h6��5t=ؠ��p��8;�"O���cK
*1��(u P\��<�v"O���GF:�h��`��e�16"O&����4 ��Sa�·\x�i�s"O�Z�bN� p�5�H��2Z6�bs"O�����%�F�Y�;$�Iv"Ol��	Na
9r�ƍ2�\�w"O� ~A!J��P� �1�EU��l�%"O��Q6j��v���*�$2K���F"O:����!	�|(h��ğY`N�A"OFxQA�/�8I�Tj[�:4�Uر"O�l ˲
T|h�i͇�$�@���8LOJ]׎ NC��`�*��n��G"O��Hv��4-0�Lq�ʒ��L4�f"O<HHs��G� -I#ʌ�����d"O8h�᠉6~��M��H�<K�ґ��"OvL��,K���`�Ǌ	<��L�E"O�����bt��Ć�X,+�"O��1��ߵE�����I^�
��"Oh5y��Ή4�d,V�ܕS�^i��"O@qFQ{��G�X�pi�Q"O\r�"��8�ށb��jiU"OZuXtKD:F�(�{�*L?iެ�c7"OޤI�煑� A�ڋ'#ص�"O:�t#P62I)��*���	!"O��!�*9
�I�hW�%���"S"O��:� =s:��@'Q�m��t9"O�p�g����Eܯmd�4�5"O"Ĺ�e�Bh�8�s�lM�y�"O� ap�]$_�J��FC�v8��)�"OX���3�t�f�)*�xX����*�S�S����0�pq�r�Ç�B�	:GA
(е�ʑb����凞�~�B�	
���	CÌ&_�f�B���.O]pB䉊)�*�/�)]t����H�)rB�	����7��$k�~��@6O+ B�
HxIr��C(zlTғ�A:�(C�	'R��x3����-�E+�oӒ"C�ɼ_�>�C�D�P���T
�<+"�B�I�-�����/�3hd��.S�,��B�ɫ�dr헐؁�"�ѳV~B��j�Ұ� A~�D�͕INB�	�>E����:j��LM�8�'ў�?my3�A�[�x%��ʃ%N(�|�Ԣ"D�*�	�=KJ�c��BGB�Y@;D����f��p�Fm!��6Hn�)�E�8D�|�C$E�[�����%厁9��:D�8�wlHH��Z�W60m�����9D�$��FC3K��m C�K/8�H-D�tsbi	�<�`��������"$�*D�x�/���j-0g+8Qh���e3D��*�o��H�n���g*
��;��0D��x��ذ#"v$��4���`O/D�p�HO�X��.h�z�32�-D�p3�������5�780>�X��)D�dz�Ϫ-�.mpe�F��p��=D� �!��+o��l�����wPi D���ƅT".U���'��PR��<D��A �3�0z��%i�Px��l-D� ��_�15����
:h�V,8D�t�#gdL�`�S��F[ �Aee1D�#ƄY�D] h����XI���`�.D��YE�ұT� ���� 1���2D�Ġ
!
l��,�#ua�|c�$=D�����X6��{�
�2��<�dj:��q��|;�F�2����5ݢH����"D�,ѳLM-�VEb��f�� ���4D�����B�24�C�,�,E5���E&D�8)��^�t��R�Xz���I D���3�ۃO�p��7�J)b|��k��0D�$#��B1e���Qo�.����� /D�� ��-"�:]�B��X�m�"O�
`�1��=��n<0<� ��"O=*��Q+N�X-���� $x�e"Oܼ�ԍH��4A�"֝4{ĕ:F"O�)���Y�I�R�`Ýr⥳�"O}�Tl�[���bS"I�W����"O`4hVm^� ��ۅA��J�.5�"OxU���#5Tq{G�3b���"Op�r�ΐ�%��I ���L\p�d"Ot� .��_���aP�
�!�:�(R"Od9�o�-)��h:!ϙ���P��"O~9�1k�mb��5�K�`r��i�"OxD�2���R/pd��M�w��Q��"O.𹤩ӓ�.��P- &�0�"O��k���>�JI���Q8�T��""O�C!�R�[T�=����C�tM[�"O(|�`�
'2om�Rϋ�y�L�a"OD4�*�7ո-��'Y7�ȑ�"OD�r�R���n
0&Xɱ1"O�d�6�G3��)amGt �xR*O�X�'C�Z-.U�fB��:�>�b	�'���rӭE+:�\����b�r��'ۮ�QTd��	�U���	Ä�1
�'zxQ�cMY�D���T�.��'�N,���/~Qr=��(u���'g��(FOĮw�.Y�ƍ�k9�t��'�@�!�%]�!�a�,�4��r�'����d1�e���;���	�'qz�3�E�eb�]IQ+P/{N(���'�>|�G)+Ҳ)X�HTnc �A�'%,���(��[i��sbk�r� �'Z�%�W��#a֒����6����'|.�z��E�aЂ	a��X��'��-XE��A����r�ȧ"��=I�'x<���	o�Z��R�������'� �q"
["�$zbIZ'ı�'�0͐�A8�P]�@]0V�}�
�'�(�A�B\O�<�cA�؅#Q6��'+(��W͐P7h���OY�O`�'V��+r�L������ś��0��'pl �DM�8�jܺ�L�aT�`�'�hP�(� ,�g���'�lz�`ċX[n(B"؛��'��B�b'F�h���X�u�����'�`LKv��[���k�r��hY�'������0>gp�sK�i%�%��'�В��z��ia&��X��m��'%v�J@��<Y��1d@�F�B=�'�J����MT���#�.Y.��(�'h��7B��4���g�ߪ��'=\��� X8]��0�d�V��a.D��Y�+�R �:���Gbv����,D����\gVH��Ζ��9��(D��	��[�:�j�G�т9|��o'D����jǪ�\!y�F
���ԋ?D�x��N�4QpA�A�%~öy�o"D�<�DÉ�H����F#C�4��i�B,D���Q�[��ec&#�!C�
$µ->D���'M�&}>T9�G��Z�����/D���;�(�@��c��%�U +D��9�{��4`r�N)}*��3�'D��Q�S�lel��� �-F��:5k$D����,�����b+Ӻ]�~�`�!D�� P�fdܐ���O)��sg�#D�� �tZf��8�|�7��	�yA"O��ĤCq����Iq*IX"OqHA�Ðl�����*e@�=�0"O��q��
U���A��e�4tS�"O�4�#�H�������	s���d"OD��Fe��,l��ֈQ��yq�"Ox���E�%f����%W��,�"OdС�T�B -*`�
�&@W"O��ru�ڥh��<�RB��C��t�@"O@��b��`��HrJS�kqLT9�"O�<X��� ���`�F6LA^)�"On���%�0L�b��/]=*���"O�D���mܥ;�#ģ]/npq"OvM���c��a��b<(a�"O��1��	v��`���3%��"O�i��'*q�0�hݲs/r|�q"O��sσk$�Щ�'U�- = �"Olak�gK�v۸8X�]Y,bC"O�A�׽_� �kH�-��"O�w�?n2�ĢҪD�r�JtP"OX1�V�����/��0"O.�k���?�
):�̢||Fi�"O*4�RK�q:9r%=:����w"O�(���@,~�f8PA������ "O����ܻ��\�!e�|�nX��"O�+���E��9�e�~��"OQ�P�My�I��" �<��"O�q�+Ցb5`�����?t�ś�"O�I#�.�3NJ�勦�уg�Fey�"OB�E��T���X��նx���E"O�}ppJ�P� A;$)ڿ\��"O� ��!�"l=B��Gg�x�y�"O����.o5��bi[:Nj�˕"O�H���%��h�B+�&d���"O�d�&�O	$d�e	��MoT5"R"O*,;bg��w�j����S�`2���"O�I�FE�,a.�W 
2_W.˂"O 1�v�]1Q[��2��<lL�aB"O�H���-!�4!��-/&�µ"OԬꆇ�<\�d[(+ B���"O�`r��ܺ����m�HS"O8�A�>�B �"��0=���hD"O��'�C�ʼKgXzf�ؖ"O���w��*#���t!�OS;2"OH]�dDڊ9&��Q���:^���5"OZ)��ٖ�p�a 8n?`�A�"O�AC1�X�?�b=ڄ�D4�1�"O��� E7!�� �2k��B2"O��!�����p��aP7E@���"Ov��q�OG����-�g�a�"O~Ȩ��_�D~,AcI>Q���8�"O�!�l�z��ETOQ2��|�F"Ot`겏i��m(�.�&���P"O4\���+,�Yb.3:��"O&��F�˲=[�����v��(�"O���6�ʯ�@���[>k�0X�"O�e�RT8��(ar�_�{�"��A"O�t9!�;O�2�ƨ� T���Z"O���Ø�j�v}�P.Z&�H���"OJ�ʓ�/@��i��¥M����"O�4@��E<M�����բ�B���"ONH��nc�|H3�¢6$��3"O�<3 ��V�
c
����*�"O�9��C��!:ƌrUjݪS�as�"O� 2 �S�~�3ꅅO{�l;"O�MK �Ң��I�i=1BL�[�"O�Q�@Ҩj k1(�a4���"O����ō�^k�(��a�1PA�%"O>頰&Y	Z��ara�<[BTS�"O�k�.�	OD)S��Ұ
̌�T"O%!U�̇[Z�y �Ҁ@���"Ov�!eEG�De���'іr�H�3�"OD��B�]V�-[�f� ���"O���1ȝt�<��S;��;�"Od�%��&7��}bg�;��7"O܈A���^* �2�坃?MD���"O�|p'lãVh�ib'�-?Vr�"O"����X� ���_�D^>8R�"O�}hsX���P[G�Z|I"٘f"OZ�2����Ra�)qcdD�*���"O�D��5mPbV䒮o��`�"O9�!�h��"�T d��a"OX���a��^�XT�F'���ɳ"O$�c`Ƅ=�h0D�V2~�=�R"OfA���� zQ�Ҍ�Tȴ��5"Ol]:6MJC�8�W�W3�^��"O�`�df��jY(bd�F�0�x�"Od�!#�;3Ŭ]�b�(M�r�"OR��f&ϽTD(ys���3.xt`S�"Oج2�`�=r�l�` �nod-�p"O���%��b*Dq�b� iRj�¦"O>�zԫ/	@�����5m68�A�"O�`[b�+d����3�@�M,dq�"O�EZ�(`���R���	p�Q��"O �凇4_I��Ȥ\.�t"O��kdI�Bn�P�	\�N�F P�"ODX0�n	�b������ޔ�`��"Ol�G�V�!��\�w��x��+v"O�	����:��Sw皦PoL��7"O�ٚՌZ'�����4l��(�"O��kLB�l�j1"$R2M>В"O6��D*E�M��A�K=����"O��v�K87p���@Ӫ9�S�"O�T�D��\z��ׁ/\"�!�.�K�<!1�_u��[�J\�[2�I�CfVO�<�d��8�ҝ�%A���ܸZ��BQ�<�$��[⨱�Gƈ0L)iaLL�'a��g�2[�lH��.S�5� ����A-�y�@�oTT#��X�*x����$K�yRA����SK1ܪ��֯KY�<����+�ٸ�G�(c~�e���k�<�̏�P[�eن�E/0Gx]���k�<�%	�p���6Ŋ.1�y*� �d�<)C�Q04�p���莪j�4j��^�'0a�dj�=S��#+O�C���3���yb��z�읐�l�.7������^�yB戊1�ظD�E�"%���Z�y��Ƈvi��`	��oR��M��y��1�lh���ӑf[����@ó�yr�Mof�P�ʔk���`f�͝�y�f�9t:��Sgc����"g�y2�N�*I�gΊ�>4��h��y"n
�e'����"�t�X��F�yrK��J��3��Ghn `��펊�yB ё�F0��+D^��9�ϓ��ybFF�&��Q��g\S3� �%Y�y���S~0ܐG���� ��S+�y��R�^m�aY���Z���g���y
� <��ԆL�������
��%��"O��3�ˀx�6E�!U��N��""O����ԢlOfY�Q`F4��;2"Ol����\�����)�M���"O( ��e���Lt+1��VD�D"O��2dm�f�����] UAZq"O��1!↶�VL��E�M��1`���OT��I[$b9\�Y󋀟dv|T�5Üt�!��J84�q`�,39�]���;Q�!�_���cqg؅MG��xa�Ԯ%a!�G8��q�C��|1�����NpH!��>?D2I�0@��1f�%G�!�Dɢ=�T᪐=|�<���bJ<��}җ�h 5OÕ$�pi���Y4a����5�O���`�i�O6j3d�{D�	-B�9�ȓw��d��%~Fqc�
�=vX�ȓo�T��#B�"?�ӳ�� P�ȓ�D�ס��9:��m�8H��p��-�N}CS�U�o6���&�ٻ	�$�ȓ���I!�ςp��E�bCT6dW|��ȓ�h�ȣLB扲�Ț5���E{�O�\�����>@�:c/#x܄���'7�mB�aΝ=�X�h����:m4��	�'�@��rh��v1�D�Q�93L�1�'t� 앆a-���C53�
)	�'r�Q������l���ù���h�'��js�'<e��r
�]K���'tX5�e-�x'�x�j�Q�޹j���hO?�r`
À���LC��I�TX�<�SmB�`�x�r%$0|y�H
P�<aQ	��x�u�N	{�f��@QJ�<)�J�KC�´�� s� d�5�{�<yQK�,��<��Z���<�f��b�<Y��$2T��C$h�#Jp�%�PG�<�s��=Kt���� 1~Q9UB�B�<���A8*�
]9`F����hqb��{�<aDn|z�Q�d�F,����L�<!���A ł4)C�o:�� �L�<��ib�t}
u�)4��=�IG�<�R�ڦ�21�g�Q���%�D�<�Į@#HQ�\p5kI�\�^�*�hXF�<�pg�j�lK�H�qr�B�Ll�<�S٭z��$L\� ���Bi�<Ԋ�*{L�`��*�Q���KT{�<!U ٍ��̚'�ҎmK�0�x�<����r�b1⣀� CN�ȅn�u�<!�I��I���Һ*,��Ɩ|x�Dx�
�$a)�� ��!��u���O��yBoٍ(�vuPs�ف?�Q�!�C���'�O8�+?�D/F50,�|�B���8 ��)W	G`�<%H�)T<a�ɡ'㒕C�jLP�<5��c]2d��w��Y�E�<y��Ŵ8���E�f0�"E�E�<�s��p��	�MK�1ؔ
��<٧�ɴ&|��JVi۝�^�;�!�|�<�v ��Z�0�s�a��(^�p�B�	�iX�42c�P���i�9�B�	&$+��M̯J.J|��!�=�B䉯C�2LQ�	��U
H��׍�NU�B䉌n���1(ٶT��X��U�K�B�,�Q��Ӻh�����`ӑQ�4C�I�/^*%Y�D�`Τ���ǟI������L����:�(�ɝk'���"!��8+=,5J�A�
z���"O� 68سfԟ'!�l6�
%B� �"O~I��YM(��f
�cf��"O
9Ȣ`�7(�8��*>t��V"O�]ş�]I�<Ht
�)A�ּ1�"OH�A��	&��<�S��"3���W"O
X@��~�� Ҧ��/.�)��P�Ȇ�I?p
L��I�x�+�.��C�	�.�)��c�MʂX3d"�
��C�ɿN�F�8��\�9P��ac��R{�C��;�@i2S7�Nܫ��	:6�C�	� �PȠJҢ[� ����I�	�B�	�R�����f� l��@S$���$�WP\Y��P�>M�� ��N ��Q<� N�=�:psb��i�%b��_�<Q�#��F(�A�!z�Z�٥�D�<��+D6�Е�WL�!��<鐅|������:ʉa�Tz�<i�l�)ZQ`Q�H�8�x��'�u�<y�/�?~������d���BIs�<�gm��.|9���@3�%!D��f�'���_���	[�i���g$\]�B�	�Q�f����{���6�J�_l�B��?�	�FJ�_eP����S~�B�'4�4���"�%C�@2� I!�dE<�(�F2�M
'i�e�!�䁴
2|8��٩A�$�*!�ĂlID��*�68���/I�T�{��|2F*G3ְꤢ�~�2���-	!�d�}=�4Ԡ��Eh�d v�;{�!��W;��0:7*��IR��KT�E�!�<#�vX�t�ؐi_�i(��H6n�!�L52.8j���P|v�z`��8W!��Z�`�t�_�`�qVB�FQ!�d%bB<iY��їR~���aMf�!��fW8�"V�۲FNz�`�`��Y�!�϶y���5D�(9Q\Y;E�؟9Y!��D-7,��&��a^�)a�Ǖ4[V!�D�Qn2��瀟 0���i�;'!��7Z|�ᅉ�#qL<��j˗N|!�D]n�X�g܌�L@`4���y�!��,$ ��7nڿ���@�Ub��R=Ob�b��`ȍR�Fߦp`�}�$"OĥږƆ`�jM�k��u~�\�"O��(6��8-o�8��	ė]~!Z�"O�ѫ���<�6 +�IQ���"O�T�U�ޗ19J̱#�WIBС"O�P#3l�z(a���$l�"��'��D��"[����JJ��!@ܱC�!�ė�b�j�@)?�1���6!���<}er�����mHyk"aJ�.!�D�K�TC�i�9Z-�7�ӽ/!�D�Vw�B��ՓT؊�s'o��H�!�0R����1�M�N�|8(��n�!�$�).ٮlj�L]�	��x8���t�!�$��w7V����ƣ"zf�Y���1�!�ާ��q��:j_��릁��!�P9� $��6[�U�b�	!�_p2����ݤfS��`�!��J�!򤊚[�X��%�]'O5>1_|NX��'��Lz`�++�)�����/mĔ	�'�P]�Vi�Bu��jQ E8\B:�H�'n(�r ��2cՒ؂�AV��t�
�'��0{dFF�\��0k�w@D�	�'~��J�l�}h��w!UuJtY
��� �ڔ�ĳS 섡�͆�r�8(J4"O,�����A��$�d��9�B�KA"O ���@0o�*)CA�9�"�z"O�E�B��0hԾ�G��o���'"O\%{�,ϲJ�AHD/�8n�X���|���3�'%��	p��*~Q+����9�:�����)�iS�9�G˺4��e�ȓD�8�cs���<x�QP�a�~���(Lj=�"L-J"-���ܑ㶀�ȓ`�>��q��;?%p���WP�pE{R�O�����E�!�0<b�C��N)H�	�'���J�jK(Vv%�Ú0YbX	�	�'�ijS C
y^Έ�����!�rɩ�'���c��^+T�,u�b/��&���'���BQ��MT^�p�B<. ��'�1Ҁ� 6Ș#l�2�&��'&=r����az(�Mŕ7��%�N>Y���	�6&���"ֽ� Ş�#!�D�4H����wM�uw#��ff�'x�M���4TS��h�䇭$�6� o�y�DT&˜��"c��
Z������yb�Ǳ}����B��P��A͏�y"��U���A�P���K�1�yB�_�����H�+�h�c�y&�^�b�P;X�� ;R��y��ޅ}�����&��B�Z�s��!�y��6J�B�U�M�A�ܴ���Z�yr�T4p�<��fT<nw���v�&�yC�w�
`aF��;gp�9rw�S��y��Cv?z����k~PpY'.��y���l���雏e�\"kE?�y��J/@��ӄ�[��8 2d@��y��D�b��/O���R����0>�� ж/�.ݑ.���ݨ&�y�<I'��N��eSSg��(� ��j�<i��V�#L���V�� �AD��N�<�!����h���������
K�<���ɉzEnd�#
�q�A�[m�'g?m0��py�!�(ř � �+�@9D��� L#7�5���*��K57D� k���-q*�K?Y���3D����+��Gq�]�R� �V��S�.D�Z����Lpهc�� `��b2D���0Ȕ&t���瑈'�%�Bb6D����N�-�D��@珂3\���a'2D����"H�m�R�	�ID}�!�%D����LC��F�1�'U�^�@a�B��O��=E��A�<g*h�t
+�.�؆X�!�$��T�&/
cdH�*7��U�!�$�2V�����C��N[촀�ꇺs�!��Y6{�j����҄	Ft(*���p�!�dL�w����2O��;FYQ�B����'	ў�>u��o�*f5����C�+*2���#D��W%� �ƅ� �C��4��N�<��N�*�B�d �Ol�t�%	]���b����j�IȜ����6���V� Ո�D�<IZ��E�VIp܇�m�0���eEp&@D�2 P6�v��ȓ_�ɚg�!�ڥ#N41����.�f�X�(�pu��4Cӵ�%���xTkw.�S�P���'�j+@Q��d�m�c?8����ƺ2 ~m�ȓ)�vԊ��F��} @�4X�&���hn��"+7^��f灭/��م�S�? :l3�@x���fY�o����"Ox�&oV�VXXa�eS?<{����"O���FBȖ<�7eKY��E�"O60Z�gޏmڌi�C�+���yR	�:H�Q)�g�ҌX�C�@��yb�ɶ>��{�����cŨ�y�X$;}��)�8�"u��l	3�yrA��1�R
ׯ����x�v��yrkW�8�:hi�͖&~C83Ve�1�y��1�*d׈��`�3 ��y�#�;qMN�82!�Q�.P"
�y���IҚ��5.����w����y�dҽ��y�j��9������y� n�`́e��9w~�`��K�y"Iøk�!r2�"k���P��L�y
�$�ޙ���c���lX��y���1H�J ��B�X�������y�ʊ5 ޖ��w���.�"h��y"�;����%�<$a�ή�y���F����DE�$�RB�-_"�y���C�B0!�`R� @�6�ygI*6[h-��4FQ����&Q��y2����<T�޷ifR����Ȳ�y£�r�"ћ�/JZ���a����y�@7:�37lN=%�D����y2��/�بp+�J4�'ꞁ�yB��'j�(	T�G4s�P��GGC�y�aϐC�n� �7������y`B,IrF�� �
 3��� ,J �yS<cF���N�%��J�
W�yң�9R.���`#s�P�+��8�hO������0G`�xʄsՌ�lM�E�	H�O�:�#dkGhb���B�H�H��'ϒ�A�lT
Mz�UKA��;Հ͘�'d����QQT����֜9����
�'����7J�,!8�ˑ6�\�'��l����&�!c mH4�d��	�'�R�A��������#(6��:I>9���,�� �������bK��Cv�L@��B�I�/����󇆓*�r�9�JՇʾB�Ʉ$��	�B�G	`��i�	�^��B�I�uZ$���P<<�h��>�B�ɝ~��� ��'Xx]z�o�<$�nB�I<7��!kׂ�&d(]��!+�jB�I>��ԋ�H�r���$�I#KJ�D{��d bhΦ�@�'� 25���zgH�E�<Aƞ�Dݔ ��N�|���FLj�<����8���SD��|�a�D_j�<a�N99� ��&�_d��7�O^�<i�E�gI��	�oL�$�T!�P�Y�<��!c'4akЊ��r�8\�� T��hO�'|K���#�?x��8��ťT����	}~�O	�6(���Q�s����ݬ�y"&D�a@(-�D)^g%�݊��?�yrǅ�i�aw)V�dA�]ˠ�ǀ�y�gҤgƆ���5W�J��0�I��y��':�49H�SJ�p`�
Z�y�.T�"�(��D�^����y��B��z�(���;?�0�`ĢM.�y�([���;�C�7 "�q���?����=8���]!F��� "^�|�^1��J�`��
"`b,셠���ȓt~���H
�leް0Ѣ]�Y��m�ȓq������r.��t$�>-�8���S�? &�)��פ4�A��W'"~|I�"O~����ԅ_\4xV'�u&ٰ�"O�쨔"�M�����$'C��iQ$"O<q��d�m��c "�\P�@"O���`S�#�轻�CL"d�N��"O���G��?��dM�'wY.�!"O���"]�%�f9�ʒG>�Jt"O���F�W�h�fA����`9�"OL�Q�&�Z�pc��|�$$#1P�t���z����/�+t�!��<TO��ȓl�N5J# ��l���N��Xz8y�ȓ)���,�:W� Pe!M%=�Ƹ�ȓ>���jq�ƴ'���c �&�ҍ��;ql� $�44�d��a�7�x���,K�$���n(^試Y2y�xL�ȓC��1�(��nrz���K��ч�z��\��՛TQ�xy'*�+m���ȓC24�W���
x���j[�T��ȓH�������o42��)H$n-Z��ȓ~- - d�d��ݹ����j��P�ȓl�N�g�M�Q"���[$kv�E��-����7f���[�$�2ؘ��	w��������b[R�䐓c �7�	�O<D�PqpN��}�X@!�B�.@��8�IM���(�Cn�T��/S`�$U��I8D���Sy��4�R�C���D�7D���5�7 ��q�(PW��"�4D���p+^"� �at
P��^�e+6D�h�@ҬGk�q�O3N2m��d3D�0Z�9\��.!��hhfn2D��Ra
M8a�|P��L;5���{f$>D��
Ƈ�+dr,�Í�}D��:af<D��f�h�XPV�*TJh��n,D�XkՌ>L���0��
�xMHR�6D��j§˼*Cl���g� e !"D�L
��5d8�"�<��d�G�,D����.�A���)�"�t�<Ypj+D�����cXt���h�����&(D����NU�q�&9���A%���#%D�$�O
`��d���56���!D�4�3D�O/ޑ�q��y�b���?D���>c�� q�:BBh����<D�h�T/�[���p�`hpT�<����Ӂl�>	z恁1n�����$TJC��d�~�ztG�݆���fZB�ɿkehU� �X-X���ӊ��3��C�	��plZ4����[V6��C䉠:�:(Jk�J��kH��xŐC�1�$\A�!��K����g&k��C�I<ن|3_�,�5��4�>tbш�<q����]�V���kt�`2������?D�`ȣn��I2N��@�H��`�>���r����Id���X�`"O������!�8ᛥ H�3t�p`"O�s�$�z��&Ɠ<3d"ș"O֬!�J�I���7cնX��1$"Ol=�'�� ;F� ��a��)&"O�m{va�J0J:kBLQ�"O2l�re�:S$�Ю�*6v	�"O&d{1�\hEx��fϟ;u�����"OD"�A�BD����Lj�4�bt"Oޕ[��|�+�MŠ_��\8�"O���%U3퀔k��St�H��"OBx�"�]�0�F8��"P:x4`���"O� 8t��"��p ��4|1�"O���#��7W�Dz�
d��y�"O
�xum��)�,4&�|1X��"O��5')���1c�O�} ��r"O�Hv Q NC|���31���Zr"O������>q���uE\�ui��"O�����=�.�a�Q�!S,��R"O���c���P�1�D=�"O:(��;	Gހ�wm����,zp�d;LO���,@�%����� 
�<%x�"OƉjD��;s�� qŽ+���:�"O>�
�D�
/6!��呬j�dz"O ��%�Z�,����N�Q�f��b"O�T�B�j��Q��M�2vT@FO� #�ݞA�������D��0��5D�����2ab���!��2��x�u�9D�P��!�OP@8c%6�P<փ3D�XkI+r��3Ԫ�ac0`�5I4D�x0�M�o�y���ѡ:2�DR�=D��[�i ��
�˗ � 0����BB=D���dͫ}� 1�̰U<x��R�5D�`��$�;9�Ft��D��r�P��(�Is����ʭ}e@U�ƭ��e���� D�(�BmE-�=�'mN>SpC5&9D��ѭF�c� Ds K�1xF��<�Io���i䣋�
E���
ð��@�Q�5D��*Q���a��ឨgm��s�(D��ō�"i&�9T-�7$Ֆ\c��1D�H3@ץL�Fa�&���V!��1D�d��c�7
hl�^-N�<]��O1D�D(��0	H���-��|A`/D�쨧e�-����k��qq���<��(��D*�d
@��!�qF9tʦ(�ȓ9ȐĎ�(�~	�IS2V��9��Za����,	27�Zq�b�����I��0��b�&�/=1(���C2��ȓg�ȅ���-'hE�%�F�w�^͇ȓLK��07NS��EH��!<���?����~Rt�h���i��ǉT1��٦��h�<!�䇪E>V��sa�'�^u�am�h�<1gGL�|9^�c��&w�XI`dJ�<�����-B E�S�@�<�PhY8�|���	�	^�H�ČZb�<��Գh��d�����|�@M2���\yR�'�i��S8i�n�r�-͌o�
��'p��#UT56�D�%.ǝ_O`�
�'f�։
�%!�`�GX*U�>TR�'��iZ#� $<x��E�#_iv,��'�:h27��](�A����k��9
�'��H���9 X��Mĵr-ZL�	�'>j�
�,ɚ(�j�C��8jL��I>)
�{N��CЧ�.r�X0
��I�f�~܄���h"�CC�]�r�駅�7ذ�ȓ"�9 CH؀	H��b�)/^�Є�|�9�G�RI8�!���U�Q�ńȓk�NAȑI�	Pv�����^qq���)�d���sHl dm�;m!82;�y�iE�tР�s�� �\���OF�y��v����W�О\�଒�@;�yrD�w	l@��c�;>j�����F0�y��:OI\�S��ߏ.��-����?�y"�e�4A7CK֨D�Ĉ͢�yR*�"K`��Pū�*o8����yb愑A��h �؜�¥������0>� ��qF�"����k�@=��q`��]�O�"�z��
�WJԨ�e!�"m([�'|P�b��M��������~����xrjV;.M !�%Hmt���#��y2��aݐ�(���2S�!�����yg�8yf	;���*�r�*�-���y�&���yD�r�4%[VÕ��hOX���N�f�34��g1�}�F)�4$��)�|�4�QN���z�e�:U���'%d|s�kϑN�(��1��sʐ��"O\�k��E�yR�3'��1xD"OT�1c���|�$@�/8W�~8*p"O@U�4lǢS��co�k�xع��'~�0�����a���5c�
�3��;D�x�V
�i���[ 	�6���[h8�IT�ИOh�	�G�O�on�󯐊
N���ϓ�OxA��O����牐H�~%��"O�LJaI=,�XTٮ'��#�"O���r$�YǮ�r��ў: ��� "OV*`!�k39�F�l~���"Ox,��׊���cFسvi�C"OTi�2��`�w��k֘S"OH��p4�pR�D�[|�pӖ|��)6Ha$��.Pe9�@�fB�	X�~d+!H
S�B!�g��W@TB�ɒ2�Й"G�T?�����DI�B�IO�x0�e�\�/�� q� �U��C�I�R�0	�b�E�4wjK��K5��C��"/�@b�
O�(%bgc]�d�C�I�e����"KK/bP���#6vC�	�u9�@�A��^f���Ӂ���0?Qֈ�8�@���_ !4UJ�Ʌ~�<�	Ԛ^�
��_�+ɀeX�N�}�<A%H�_�8U��L
�H��\�FA�}�<	B�Q�R֤�1�E&6���w����<�dB�-s�f
A�08ӄC�rx�Gx+�/  1�Ğ_�N)�4�$�y�C8^�F@0p�
�GR��S ��yR��]ޡ��R�r�tT��D�#�yIS:� y��]�0mIt���y@��0��/ӟF��T�y�o�h�Ľ#��M?Ϯ豳kU�y,�fu�9��Y�PL�c�3���0>Ys��G���ab�� e�th9��_�<	)҄V��5"T����g��[�<���% ��- f��;y���C	Z�<y�`4���%�=V�CP��R�<�vi�Lj.�W-�$��<[VdRO�<YsB�=X`}ҧ.��|���2�fCK�<�G��O�8��r�
, ��'��Jx�<Ex�BÞC��#"�$��8����y�o�/ 
�kQ�M�����y�:i�J���X��vI�EhX��y�FƄ$�2�YEbːY����0�y2 c1�`�cbԇZ����?q��d8�c���ʰ�H#L�2��P-4&�neK
�'3���ۣ(.$���I���̨	�'%�#p��2q�:�ca'C�b���	�':J���Y�yb�%���պG����'(�a��L�;8VxX�W:�ܔ��'�μqd	:ܔ�����5g�����'_����i\���ɜ�Q�"0B�'c������5�b(�WNխ/4���'J�]���":�e`��=F�B�B��� ��p��Ȕ����V퉟7x��� "O�)��l��ۅ*���u;T"O�Sb,N�[{%� �e(t�"O��
��GQS�1�'�rPxD0"O $c��L2�yA��B�\N�TZb"O@� ҇r�t(�ÕGD��BF"O5��&ʲ&�x�(D���e$����U>�z1N[	K}hPї�#j钜��%�IޟD{�OfB4z�Gs�JM�w�ֺj�Ju��'PE2Q�S���X�&�\��a�'N(���@�o�(�b��<�����'��ܛ�G�@�����0z�A
�'�h���փ &D����E`b	��O����'�p;:xV"�&r�5Y@�|��)��{�ִn�z�
��nq��ȓ3pJ��Ł#��]� � �b��7�.pѧ�܅_��0���!|X��~�l�!�: H��®L�D���ȓh���f1Y�N|Ss�)6C�IB��<�F�ؑ6�	��2nR�C䉄W���U�<hc"�?%�N��1�S�'����1Ԧ��o��^܈�N�x�ўX�'�>�����Y M8u�ӯ5�V��QO/D��B��y*�b�$!�H@��/D�õ�r.<�E�O"?vD���k)D�(@ h���Ұ䁍
f�[�d5D�$# j��M�:0 �#i.�ȳ#4�Oh�I)�qcp��*7#��aG�R�"C�	f�L��l��,�5%D�'{C䉑 3R��� 7�적锣E��C�I0Y��}h"R8g{d���S( �C�	� dLĨ�8���`��gC�I(W68��e@�RX��#�	��B�Ivۜ��"��3e�L�(3�͜��B�$�b�"�.9���(V�&��B�,U�܋׮S:�@���OR "��B�I/ע$�s��0?P��c���#�!�DU$ڤĲC��4=5��q����"�!��.ZivI�s
�	&-�������N�!�dhA2�`�/�/
�$+5��3I��'a|��</�D� ��0�6��"Ҵ�y"H �M����0��	��\(�y�C¾�d���C�#�� ��/��yR6_U歑֨ �-�j�����y���R/�hx���<���d#�yO��JJ�]��BC t�f�AU ^'�yI�5�<Ęs솚h%�ykg���y�L�?��25o�_i�Y[�K��y҄��O�Җf]�PӀ���^��?Y���S0��Y��J��ɓ�Y�fm���ȓ6��Ȣ�P'c�Y����J��ɇ�o�4< `F�?�4�ɑ��ZN���9��p�)�"<�dD�GY�j�6���d)��	@��X�Bh*��[3U� ��QC�����$%3���ǣhj�l��Ug��Y�Ih�h�D z�~�%� E{���dزqPt<A᎟
��T�y���&�@HQ�C��hIja�ɢ�y%S?q������Si{,�c]��y��˛E^"�YSab�����	O�y�㙬�z�Q�ֶ}x	C��
�y�猞F��\(R���s�q�2L�9�y�
�=y\A7mˠ>Y�@J��y	_#|ix�lF�/GbE"'@C��y
� ]�TI�OF�\�0���@w�e��"O�U
��Kw����G��-o��"O��!�[���!��ÓQ��a�W"O��A#�8�f�C5C�>W� aa"Oɡd�ߝGтq��3s�f�{D"OL1�c۠
���ŶC��ي"O��*ԝ5�`�xg)��<��#f"O��S'&F"L�)ڞsV����"O>Q��L�aM���N߁w<d@�"O:����]��h��kI�C4]X"OL���͆0ڠ,� ꂴy6��"O���������|�D��.+$�D��"O�I���I�`b��*52�0@"O����EBa�S��A&J��P"O�x�Eh��!t��D�!u�9�u"O.;4�T��0��s�M(%՚���"O�5��ƬA��%9�aֶC�A8"O4컀���<�f��%5��0�B"Oya��t����h�L�p@��"O�q����F]���J��o�ą��"O�����YR�@"g�?{��kd"O�� !��1���z��CP�""O(5�sRш�H�A�]�6��"O���⅚����ȣb�R13"O�0��M�6�.Q�BZP�J�"O��0���0D�Hd�v��0D���"O�Äŵ=j�Ep�aJ�0�݃�"Oz�(׊J���KL�&v��K`"Olj�`��	v����:A��Pka"O, G��G���Tċ�{��d1�"O�-Z��X;@���C`#��ho��G*O��
��B���U"��W12Px�
�'Z�s�ON�6�2h����6��{
�'[�@�gL�X�v`ȂcR0r�RH3
�'�*��B(��*��u�2 C�{��IB�'����b ckT<�QM�=w�<e��'��tJb(A�gǆ Q��x�H��'a䑹4�R�{p��0�O�o����
�'SH,��� �|H@!߸8mj�y��@
I�� �. �{�H��ª��y��!&.0}��μ
!\$xb���y�%��L�6�}�<����y�N״}l����n?Y*�`7�y�
��3D܀9鉈q��Ied��y"�I�+ɚt�i9S{���d�B�y�cZL��d� A���ʀ�y�J�*'[� ��P6@��`��y�B�3 ��'_�8���� �y(��&tS3i��[�q�X��y�g~�p)�R���@9n��T�y��Ս�.ek��ۣ<�yZD�G��y�eD:�h�p��6��|�#�y��4�μ��d@0$|�� &�=�y�N���5�Ga�'�:e��/�y����(ڄ}i��3��	�3ȝ5�y�F^��>�:�f��0�gK��31"OP�Ò(]*]v��[��\yB"OЄ�DOZ��ش ��Sk����Q"O���R>���
��-��]��"Oz](6�	V�dX����-"���&"O������F�$���*� ��"O�a֎$�J!��I��Q��	
�"OB̛5�J�4$yӣ�w���"OH����+U޴�ף�E�%��"O� |u��@K��`T��(tGʰP"O��/ %;�~� ��ݺ="1�D"OS�k� �	t��U��I�"O�P�"�j� �aJ"=at���"OXu�`Hњa@��2D f�d�V"O�))��^�ZV�Yk��ٴ"��U�"Obx�c�S� 4����!]��习"O@�RK�o5�0��ֲeJ%C "O����Ù7)�	6M�`J�`��"O�p &MZ�O�>�87+�5	b�"O�d	�*�2��yq�����:6"O08�#.Vo�]��K7Q��`"O<�y�A5��u!�75X���"O`@�t�TI���N�&�@��ףJ��y��ϊ�4M�LÁ$N�'mG��y"F[;q�T��գӥ!��i����y���f��"����T"�ΐ�y��;�P��o�c*Q!����yR �Rq��st��?;�e���N��yb�Ħ`�e��U;5�|��P/�y�.Za��y��C:`It0��a���yB)ӄ*�ju(�NɠV߼I��,��y���$L�&tГ��K�`pw+�yB�_�
R�܃�b�CeҀ�f\��y�(�O������C�Dh���Ӌ�y�j2El6р�蜪Jx:�a"E�ybA�	�x� ��/��dP1�yr�|��h��@O����:��Ѐ�yR�I�lJ�r&H3r���"�O
��yrd��u\�A1�+F8 C~�)��yB���:�F�6J��r�v�p�눥�y¡��&&�tgʰoLZ���U��y���v�@��@�9l��ͨ%f���yR�8"��i$ɐ�`B>�eb���yB��&��0�7g�)I�����y2!� B�ba(6�ח\��Y�$ D*�y�C�D����֞}�h��/���y�B�('�d���نK�Ɖ;3I���yr�M�HHkK�=&d)k�FU��y�΀ ���	����kP���y��Vu��)bÁ�~jX��W�J��y�D�~����4㙙l���1G���y2fO�9��@��D�\jt����y�A�M4��0Ҋ\'�"`�2�Կ�yB�	�La������Ქ��y�+]T��qT-O�����l+�y�Ě�O^���.@�PBхU��y�HM��|k����k�T���y2fM9]�ɨj=cA��Pa"U��yJD1j¡9��.�������y���1(*�����(� ��n��y�� lS� ��m�jp��ВAL'�y���HWLLz .]]��p�"!�?�y��-�>	zQ��Pq�MP�	�y�f�>��Ei�*ɀM��y!#+�y���iV�z�R�N���cCD��y���^�(��g�'=�Na�B����ybI\�2����mZ	ӌ4
ɋ�y�j�� �hu����b�$��!��,wf&���O�1j�����'�!�����p -[K��Ti�)�(8�!�܆Hrqz�҆J�X��TJ�T�!�d�8s\eI�B���dE�;%�!�djzxp�nE�u�nXCQ h�!�� � �'ㄊ*#x��A2D1r�XP"O,sԈCwWr|(u�X�+�G"O�
q��:R3GBn\H�"O8A�`�T�i��HP�%��,��"O�hb�C�@xa ���m�C"O��X�� 1�L�P��ڃS�4`��"O�#�J�
4�����,B|#"OШK�I�|Y�(����5V� *"O>H�+}�x�7��nT�]��"O��:�n�/��8�%C��E"O^��h�`����74��"O$Ԩ��C���[P#H�`��"O&L*�a���j��I�(�uA"On�xr�גa� ٩�h��u�,AK�"O���c��)v}a�&5m�TÆ"O��2"G��̃x|��XU� �Z%!��3�n`j���y�M@�ʏ�s!���@��σ-[ XC�])�!��Q�B�%��i�t���!k�^�!��r��1f�X�;�d�����'���yc�D�|��`'�ؿpv,<�
�'mA��`�'��@:���jd��	�'��)�
EC�lȥ��2�(���'��c�J<�%���'ì��'Β�1k�(}�����b�&����'��I�&c׹���Uȑ�J�Pu��'���i�k9S���Jd@*Z$2�J�'j�m:�R/D^X7�A�!��-q
�'�x�c��͚
fH2�d�1R����'��e�wD�))�t� �!.�^h2�'����GK�@�!�{��TQ�'��0��j��$ u�7g����'��B��C
|�
���D^�j�)�') ���d�})����AR3Y����
�' 5�D���	���`
��QK����'�LzeC� �L��@M�Qt����'��1�߈���F@
�<��'ưa"��9G^�N	�ԈH�'�����D�1�����	[�,��'�
,�:�r�HF	/�"�	��$5<O�}��o�1D�>����*G��l�"O��Q!AȈ3�
d�����"OH���(�,�w�U>o: ����w�O0>XKĢU��8SB ��{6�I�'��Qrς!J�>���UM:�� �'bў�}zЩ��W<A�&��k��b�"H@����>��&�&�ۃ��r�ё��<)��٣q� ��r�� ~⴯a���d0�h��2w��!�Dm�DFH3 �@�ȓI��:�NȢܰ����_u�lE|b��S�D}����3����풊hT�B�I ]�hL*�
�@�liC$�]�.7��(O?7�1S�<٩�9��9Jh��`�!�Z�"D�������B��bE�֣�!���&�ru� B�4?��Q����!�d�RJ�����@ ���� °;!�
"p�#'��U�x򀀞�}ў<���7=|P���:�p��W@]�o.B��9���ɗ��Pƈ�(��@C�C䉋NIΡ9��1�~�s�)��d]��䋔A)�!2���M���	�lR�!�!�ź0|ܼ�P�)s:9�ԫ�&zU!��ڙH�,4!2�$l,�0K� ��O.q���0���A�ܨ=���V"O� V9����4}4�@�f�ߎ5�}K`"O����4��u��ɜ�t�Ԍx "O����R�~e�`OC��	�"OP�+�!��~A`Ar�m޸ؤ��*O"��H��3��8{'��be	��'^V�pgl�6-膁�_[��'�n��2��T�T���&Y�0��'��#�D�)���͗E����
�',�q�aE�98�ڸS��\C�(��	�'��8�#��"q:ٚd�!A�^���'�j DG5j���Nʙ6#���
�'e0��-��2�(Aa�嘖f���+
�'$Q�ŋ=(?�	�2��<�b�k�G$D�쐔� X. 8b�W&c�,e��7D�`�ufG����:Ø	8�!�F�3D��A#�^�gw��&"Y� x�0E�1D��P��@�V�Y��BY(����`0D���c�=��������2�,D��A"!�Z�@�撪'~�:$- D��
Eg�Y�(R�)~�fԚ��>D��W��(���:�&P;p�����.D�T����T�@9��n�][D�@�c"D���A�8{$1�����0x� !D���C�gD8s������y�>D�� �ք|�����.�9��c!D�0�W��0R6�##"PG��
�N-D��ڤh�
j�!��̨X��X�S�&D���]=6���� �T�,�Τ)��'D��	�Sr�	f��B'��@�L%T���۪K"xyK�n�l1�;�U�D�<����O��pD+�#�^8��K�g=N��&�'���	fڐСf�9�P��B��*2�듍?
�Ӫ�lѢf���b���,��$�I��M�����OIF�����1t`�qל-΢�#
�'��]Z��$HD�b��%Q��$��'=ў"~:���;|]H0�$dJ�bZX��R��m�<)p \=P�JQ�H�<¬�z���eyB�'�2Ux��H�\ڰĒ���ZQ(��'tH�a��]S�l��&GR��p�'�x0��_�Ĉ�υ�w��l�
�'�l��,��9�zP�tB�';S���	�'��e��&��+ZM��B�,��Z)OhEz���[zVıR�7�:�9c�A�:"1O����W1}�hx2��4O���ċ<{�ĩ>���'-	 #�κk��haɢ'=��k�'���g/��kQ����ʄk$���'j��[�l�(��2#l4 �9��hO&��ьx��1��"b��H��"Ox��`�<Ꜽ�p�^�=�΁Y��X���)§1������>`�$m�S�Ĩ��lm�D#|O��jS.��h,����o@�i�d��U"O
�hT��]�hx�o�!(�Lx 
O�6Mݽ%Ö��7KE5K��V��)�1O��D3�)�$!bJ��腪<��ԃ2	�P�B��^<��p���|���a4�
��B�	�-'f�	TGR8��4p6Ϟ��BB�I��>Y�J�sU����/@�➨�����<4+R�b��Q�rɏ�w� B��AZL�hAHݿj�R��c
S
��C�^���Z& )aL�a�d�C�	�J�X���%M@&�i�$L�S�zC�I${��܃GM�#��T�B�	�@�$��'��X����7N��tB�I�CP~���IG7k<�$�G��]��b����)� �����1 �$0��� � %�d��'xqOpB�gֵq�R���D /��ī�"ODy�����v$��I_��ṟ��ITx���U�&=����q�R�:��	�1�O�� M�����G�XXiD�i_ꀆ�`+�@��.��pg�[ j֬F}r��
T�(]Ѐ��>CR�b���B�Ip�HJbm�hV���ͮU���D&��O�1���x�OW�A"�01��g� �"O�q&-��u�6dH�-��c�/O:��Φ��S�'��9O��sr��`v̸!�� �]��"O.���şO��)+q/Y�=疘��"O�y�	�7��A��(�T��g"O�y;&-F�l�:u+A-ܐA����0�'X!�ĊU
QٱF��U�j]��jN1O�"=���Tʕ��b9�$' �����kD�y��Ϳ3�|X�q���X"u��O���$�-4�(��DR�Ƥ[��_�!��� y�*�H�oK"+��d�	�N��'0�|�F�(*��Ɛ�}>d� fl �hO�c�����Y�	�1_GB��.�&d��` "OVY)"��Zb��˷-��ai�4��Iw���	=E�4�;���(.�a1��:1s!�$ގwӮ������ $I�`�!k�'���!�S�t�ҩaG�D{�Q}�V��w�X4��?I�'�&�di�;��x�ƚz� ��
�'��0SeS']��: l�0o�Z��
�'�*@���>?�I��!o�@�S
�'�ū�-I�h6F��ņQ�m���L��F{��t
6_��@���-Xt�@��ޠ�yRM�6-GERp�S�d_��ɥ�͟4�4x%����ok�$:d���T��[�*
�)�v���%�INPlX���dq�Hɇ%� B�I5b��l[�e�3�B��5��	x�C�	�B��b�|�:�{G��
B��4YM�|S�j��:<⡯ߤ��C�Ƀ&:��:�%�4�U�جGG�C䉷9����oU#�]ro��x@�C��+Cy���T�9@έ��J�2֎C��'=��ݓR�~˦�q�8\d~C��:L��p�� Y�d:ĉɔ;�vC�	��rp.�K�t4���Ȩ-�~B�	�^���y�O�[6L�i���k�*B�	/.�EX�ܺ?qH�k�|�B�I$����(�&a��+c���l0B�W�����S;x6z�8W/A97��C�I9U��A���;&И�[%"����B�*�.Uò�H9[.�e0��5l�B䉕�L�Xca��S�$���Ā�F1�B�I2����E,x����ߕZ�C�	�e��(�"��4`��D!�J�PB�bq��b �@##���C��D�u{4B�I�j!�ճ��������ʜJ�.B�I��ɂN��s�:q�/ڜe�B䉮K?`p��<'�x���*R�ZC��:�TA��d{�,#ua�;P�&C�	����*ԋv���V<0Z�B䉼1�V��p�L�&h��ѥ[{�Y�ȓ0�z@��҇� kS$S#H�Ňȓ �$e�8��Ua�+ءU��X�ȓ?ߐ԰�+N��L�s��ׄ��M�ȓ*1�]�g&��R����H�>"�V���o��a��[3Vv
��ƒ2PR�@�ȓ.#���.�P8���.Qº���S�? ��	h80���N܄*��)�"O�P
âD�e��������j�nq��"O��ᣪ�#{]朡qB�9֨��6"O�L���myXm�R�̾)iz����'2T}+���o�*��C�#����Aa�4>|�'�dPCE+8!�Q&�إ(�ʨ1�'� ŻTE%l�2�KJ�z$
��'���J�
�����(Dn���E��'���rjΏ[j���z�B���'��=y���2/�t�0��Ӑ'��)��'[�8�G�����@�� nr�9�'P(I�'/�������'���	�|_t�_���'�BGK��h�7.�
\�r�'k��H`	�5n-�@��MZ�:��0	�'(*�:�eɛ�d�
D�$~�y�'��	�!�$nw���0��3Q<(�'Y�̈u��'_?r�*� [�xcU��'7��PD��'H�WM
�j�&U;�'Ә��QĞ�gI�!��k�NQ��'v��$ W��i�HRH�&��'��t��Q)�@H�Å�*I)�Y��'D�$���<�4u�N7T� �+�'�쉣U��zZ���E{�"��'͌I��d��Rt�@�K�'u~tQ��'�����2h�������)n�4(a�'�"y��L
iR�I��I��		�P 
�'���bF-$r|P�!&��%2��l;
�'�t�P�K_$SxT��5�D% �б��'DB�14�,V�:%���
� �'Ax��Q��j*��)!�ܒ�bi��'��|��m�11�|m��C�����:�'#\�S�E�m AH���(1�'V��P���)h ����̫�'@P��r�A�d6jg�\�-}��'(^��s���"o`|�hؖ|��A�'����%꓇S��i�gJ$��i�'��5�S��~�� �HΓ�<��
�'$L�kEm"9 ���F��@�d�'\���:.�~��Ť�+�Vg1D���v�[�W�h�2�
8.,,����-D�Ъ�ĝ�G��	��Ƙ&!(T��D+D�t�� +~��p��ǉ[��2�3D��գ��R	Ti��n|�s@j3D�
q�ы:wl
��]4=f)�5D����M��U��)�'aZq�Z��-'D��iR�ȃ1�LKy:1��J$D����^H��2�$ͭCP��11"D��H KB�FL�%��
%8d(�ա#D�\��
M*�Q��
�F�xso!D��*Ԁw&�hbm��.Ĝ0���(D��Z���B���d�ҍhɨE��m3D�d ��F,i�x��F2���1@a4D���n_�0�r|�r�O��4��"2D� ��%w�P�Ӵ�
(9,�I+�b1D�\y4�¥6!%1(Ϗ)4leXw0D�p�G�l�cG"�n�x+�o4D�������x�̍r�()�6D��ec� >�bQ!�'Ur�j�8D��	db��'�5��S�lRH zg""D��X�Ϙ�gK�u�S�, ���^C� �:���W���"�ݨ"��C�	7D $i��/�#x��Q)M0F��B�	�2������O18�����ɕ"[�B�)� *�J�� *�嚏2�;�"OMi%Ȟ�w���FO_
���P"O��PъL��ҽ���_�"���E"O�II�J�$�e����;$RA;�"O(���`��:�5!Ư�$��l��"ON,z$�ÒL���CdC�Z���"�"O(�д��o!��e��.4zx��"O��ѢH�sOXa(��~Rx}hG"Olpz"�)C�>=���M�B�Je9Q"O�LY���7�0��@��"���)E"O����B��\���i)"O�d3�M Ec$mT�R*�I�g"OV�	��[�mҬl*���e,f�Ї"O̰��B#�X��%0jP���"O$��4I��z5�S�8+C"O4lj3,1�q�w�OYXu)!"O\����#�����$��B�~��"O����K�\a�lY�-Gk���$"O�d�s�ͺ�xB��&OKn0 "OF=9�h�9oȼC�6^ږɚD"O�ᒅ��d[Fq�$%�?bZ�*1"O�ܚ5��)	v�a�fHLf~ �e"Onb�锊�� �%M����z�"O x�(ٴ-��a�$�=��`ٶ"OȷߧpY豙@��:u
�P�
O��ㅕ)$���Q�F�.	�޸1���'_Z�J
�'l�[D�GP*��PEG�5����f��DV8�d��"+�4�b��+;�E���)X��"Y�@�ݏ�x���'���klϹ��!؀�|�̄C�4{��'�_�8s�p)�ď8��%�}g��\�|�k$g���1�ůM���	�GC$v�z�;U3O�dZ�BC-OP�f�r��*q�&D)6�$Š>j�E G(�(��3��*$�^0y����Jt��=ɓBQ �N�W�7��$�R�w$׫O2r���6lN֐-B��*L4~ ᤊ�vx�Ա�G�56�D�� �
�a`P %�Mt,u[4}�ʟ;��|����*PAc�k���;(r 1�EB'�myu��R���ȓ)}g�}P�\�B�wxd+iK�'�{_�|���4qr9��65}�A�weNe�6kB�١!M��%��P��%&pʱ��ɣ<���ڦ��pn��!
z�lJ��@#�l[�h�$|V0���J&u�(�q���@�P`��U?�kW ��'��1҈VO��A�@�-?b-	�{E��,� mQ�ӭ>
h5Ir�%0Z���ݱ$U2��#���1- ��#D3na�cEÙ9�����'>����	0]���8s�ܗ`:l���8/��	�M�p� I�>qQ,�cvkPl���B,@��r�ǅ���4��G��S��"���l��5(��;�㙤<�̱EN g��	��5�tQ�>Y��Q@�]An\�뗀���uW��D��
Ad�	ƥқ���"���xo���D�,���O�䈲�ђ2��h	E՝v�L
q�N+>1q�I�f^J�	��l�K^���/��̽u(VR��D�&�$���&u�a}���O�ҽ��DO���r��7���0K<}�Րd�*a0A���j��˓N��H��2d.}�sʝ�FfRtGz��'_|��vذ�,����0#�E�0��i!���3�]�>��e♕z����'�-C����}y�-� ��ٟ��&�/�z��7�^ �����o�o��j��	�g
�db��O5^���L�5n��B�Im j�3P�S8�"(�����t����V��� ?"�qiB2Y na(WH�|�4�E'
�`O�ثt�n*�hRm?���'���ء^�fo����'��uPf 2vX�<,���Uf��ht�@W�� e��-�B-,O���"�.uq� �$�OP��q�6|V����B�|�X�I�8DzS�����z�j՝4F!I��Lr��a�'fP��UF��,�P�f�J��2�'�NlA��C�B��'K�v�ʔ�7�\|I���;lXp���}��y+&n-n�!��_�f��	@@��+Ey�`��Y�H���z����@�b�獷����������w�I&_�����/B4X�����,�)/(���R'\���2Q%_�k��E�ǎx|z}xR.�-]����ʏP�p����Gx��e�M{p��+P+�'�N���j+}B�֊<L��'n.̳�%��Y,�<d�L�V\n�����=9����U:,�����b�n,�ēE/R��A I���lۂEHdtS,Ov�{��Ĳm5���Q�uh8r������M���� ��q�`B�&�����M�+萹!��'���A���}w@q(Qa\/A�B����ЀV��,�甆��B���O�
x��'rDu�Ol�'��q�HE"'P��6�I�~Y�M���"��h) ک�ħ\oRY[g.6錩�P�\0]И�':ҸcfnC&w�~I��ɮ}W:����G�=2�����˓{�04�6H�0UoF�c�K?�ӫ7&�	�u���x��[��]�X����)$bfF���O�M!�G��f���	a��U��M�%��`~��`�'�b�	��۷IU�Ua�b���O��R���A�No�横�Ib���DˎQ�XЕFفP4d����5}"epv��[c�E�:�P�O�4@�J�/rt$?5k6&���ţ1E�Q���cSB�'�V�J��G%(T]`bf��O�W$-g����\7���1�V7@��ɹj 8��#�mx����:0��e	����d�T���<�����=M�Q�mSn6*���di�4����lM?��RfVt����NCr�<Qa��n��͙2�6:�J�hf�):2��։^�<�c*�4d��|�<Yv������:�iB�v���:�*JS(<�@�S�(:|��GŚD�Va1&�3ip�*�BC�kpL�q�-5�O���K�{�,�+#����̲��'��b�bG)'���ϓF�(�F$����ф�)(�z��ȓh�ly�CS�0�ْ��j�0��=A�b��[�]kF룟�� &˒7�/݊����:]�\�j�D��C�Ig�l�F̝�!#� �&
��86��Yn�'n��$�7SЙ��.ʧ����,^�0�gưI��g V<1�!�dV /,�9C����XX���[�)�h�Z35�ܭ����Ui��֘#=V�B M��ᝮ��\SC�}h<�jQ����҅_Up��Hc%f����k.���.�)h�Ȋ:�4��77��y�hJ;�,�Iq-�w}��@�Q��d`)0�<�UOʸ�y҇@�*;����дEҼѫE`с��Dײ�˵�PJx""���U� ��`�ĝ^/xȈ��L_�<�@�
�dD*�!�&&�H)5M��(��c��>9�>����I��%��0bX����,J^�ݫ4O�DK���#��d3���e����g�K�'��i��N7��>2ɲ��y ����L�ցi�Bex�|� O�ڕyX��!c�Yv+"�:-��H���yҦ%Z8t��g�1 e%��yBf�� ����Ӆk�l)3㍓�&���R��I��B�	�W�PHF�G�OO�=p�1b�hj�*%�� 0`Q>˓x� Q�#�\D�-[�#!��ȓp�H��b�{(|��%�I�~���R��{�(Ą|���+r�|T@�ȓ{�ۧ�yMP��JϤ��]r�'�Fe����_����.�h�'x�Y´���,��Y�A�`��'�<ō��x�u��Z'V�b @	�'�б�0.�a� 1�ݕ4���	�'s�I��KB��ڡ��[A��
�'� U�T�H�V��L�\VC���'tL��� J�"�fWVƩ��'x �cڪe~��;BַHd�T��'�z%
S�TNj��!���K(���'����R�
�@��g9���'��B�I�&4*!cڠ�P�H
�'�pb��S�����-��\EI�'�����ӑP��pq`,^j�x(�'N�}���wIL�W&�#~?le2�'+�@å�{oZ��'&�t���'�*u�@���f��c���A��p�'����r���8�&ʌ M����'�8\X1���N�֌	�+�r�'�ܹP�@4`S����j�'���PoK*p]�8R��&ddax�'	r���G؊=�~Y9�Wcv�ݡ
�';^�(qʑ�]���P�F.S1�+
�'�d}A��ԅo�
	��DGoԳ	��� ~�Ku"�9[���1����1`��z"O^�cI\mO��U��~sJ�q�"O�(�'�X�[���㳮[&eP�y�"O�$)+T=J��US*��7S�EJ"O������L�xұLM U*<�U"Oz��"�ɿ#�l�:��G�sW�i	"O��*&��t���#�]Gt��@"O(�*3�ӒI��Q��)N��w"OPa� 0/@�(�l	g��	�"O����	�r}��#�֒?�,���"O�k �K%$��(��H�c��ɱS"OBP���%��]b�JH�д	�"O��!��$F4!�-[lz|�g"O��:$]�p�lh��L;�*O�
v��F���y�,aa�'�����=Z���7���{�$�Z�'�а���ox,�Waߐw&��
�'�0������-���sg�K<O�\�
�'����P#��{�t�2�*������'�Fi:�\�v�vIa1�K�jj�[�'䊕�� 2A٬D���P�e���''��*��n���r��-,^ܬ{�'��٨3��	�͸�"J�	��
�'ނe�ʚʞ�#�bE�Uf��B
�'����W��)�����'AT�	�
�'3t�i���{"$�p̛��6��
�'��	)F�E�DWt�`�A3��)��'�0c�N_^ظ���6z2���	�'�aC��A��Q��a&[ภ�'&�p�E&D�D���g�d��L��'OV���^�a��QЖ�S�d�r�j�'�x@�f�3F�(�e�W�I�
�'����V�2��E%̓�A����	�'��I��X����4��'(��K�o5�n��M������'��ᨤ`��v<<��
�b��!�'5@�Q�K�E�F�*�O�f��P��'+�%�@�8��y�	@ب:�'*��(Z�9b\`����<q�'�N���9{�
E���b8*�ʓ"��ɵ�Zrԑ����9G1,��H��y� �*of�Kr&1B�Y�ȓJ�+7%�R�|PKG��/J��D��N�2��H ���@3<"L�ȓ|�:����ֿ��p��ۨZx�ф���`���$6|	b���_��P��R��y "lC�_��$*�ft��h�ȓf}��j����;�z)R��L�pNX�ȓh�Kٍ�8ڠmڹ-=r���'4D�8;w��6v@�R� ��{�R����>D��i��C$N@}�k�&M� ��(D���֋ІX�fq
0����+D��Q���=���矃t�xmz�)D��KE�82a�t��?e��ɚ�o3D�d#"�T�R�N7������3D��yC�S�*Q�=y�)Q�T�)���3D���vO�49PAP��Na�r1+�	-D��24C�S/�����[22�ܢ@6D������ �����
$x���5D��p�D�7l
!�Q�0�"W/$D�l�r��'��ڃ..4Zن�#D��@5��G�Ѐ;�Z=0P�m�G<D��XV��}�\���q���p��:D��۰��C�Nh �[ Bv|h04D�� ��Y&/--vAP�B1s.��"O����F��,Q�`�7 b�i1�"O��W��@��,�f�rY��d"O,���D�5:7�E�Fh��"O��p�KBH�WkC�2Ht��"O��s�w����q)G�I(�1�"Or$��R�� �v�G�Y�:�2"O�)�Ќ�>����g�[�l�R�"OV�;4�;+d�a� ��V�9"O�`��/�/j�D��S(�/�]�"O���1#\�<��B�40M�Q"O0 8�@A�e�A	t��<,,C4"O�ٓr]�A�����!_�h��"O�HB�#ҮJ5��G�]/�̐��"OZ�ꃪ�$OC�s��ɸ���"O�<�2���T6f��foU0<z�2�"O�ɓ�3-�	��P/J`PJ4"OV�X��'��03�� �M�%��"O	���Ӯtn�*�L��wI���"O��xa�[L���Z�,�7�0�R"O e���1T�YA�F�"$t�ؐ"OZA��e�	�05�tF��u.0�	�"O⭃AB��ҐB���q�N�y�"O�q�ԧGu ����-3 �H{u"O�E��GҁQ�.)*��ֆJ/����"O�	�����4R8 ��ӹD�8��$"O8�CUƏO4LٱĎˊ"�P��"O���,q�b�#W�	�t�����"O���i��aY��Ц-��B����"O����B�	L��t  l��)��"OB���B�f�"h+Ҏ�5�^<KP`�nI*P�=!���O48(�m2?�ӗ�4��y�"O�����P�D���'ڣb"��ӹi��@JAʘ)S}�|��V-1D��c���ە&ħo����� Y�1�I0�y���8M�*�)rJ��_k���[��y2.�hj��3\U���eR�ٸ'���iG�u_�LG�D�
#U�8���lF�E�x(�C��y�e�a9T�B�ΞF��i $� IRn z6�U-���,C�Q>˓|L	�DH�M9b����@8[MT��ȓd���Ņ��F �V�:WVذ:a&�ZPF�8AτR�@�\!t��B���~��0�0\O"�(�!��v<�(�'�	��CDA���S�Lvd�A�'#� 
��]�S�OQlMCt����,X����W�~!҈{bHW*F�A��b�O=����xzmPBJ�&(�d�'�����$�L�yK9Kd�1C�b  B���Ꙓn�J��$暳��3$��2�Z��ۭ�&�TnN�sd�ئo��E�F!8�c��Ȑx�H�&z��р׌���U3e���M�d������O�9"7��.w9��=}�OR0j%�V�2�'f��#����p`a(b�>�����0i4*
�)��A�a�CN�|iRp(�@��̱�OZ�8���O~l���*߲��L D;�qOl�3f�/��A�ՙ�x�ɕaCP��A�@�N�!�A u�ay�f�7�����Ԃ)i�=�&��p<yS��;P������yz��9#M(~����S��>g�z �4%ٖ A<���'�&��	� +���\�nHH�O�	86l��6��Ű�HP�W֢ib��@���hp��R�z+�]z���G�݅ȓv/R�	v�I�w�չ+D#�d�9��b�������N(±��X����'Z45��H97+^9QO$W$� ���{^8���եn�|��LX�8&Pܪ�-H�z�Da�&���ϊ}蓂D/I݆���=1�6��@G�9Z� ���}�џH��+� ��8U"� x!��ðͥ\���3�מv�X,`C�6�E�O�H�c"D�-�Ƞ,L)�~��R� 
�&	37U�ĻA�D
/T�Xqg
#0j��>{���#�� Ss�Ջu�Ux"O��7l=r���1���'����� ȡ|�b��J�P^0�(�/�	l
�O[4�$��"W \	C �J�̆���1�<�O΍�@=� ��8��_i������22Aĸu'������[�;<3d,<O��@��8�QTLڟj��=�S�>1���>׼�,���P�#`��T��O)LZ8�F��~��!'қ̾8��o�5"bB�W��=!%���6$��LO.��|�'����D��>����<vE\���`�!���ŦqͻEG�S���w�@T�?>�4��	�DB�A�lE�	a��>�h�*�L�Ӷl�6ĘP\>Qȣ�F�#�Π�ImD�n�I����1��'3[.@�r�"!�f�?���*S��L�@�+�)��V
��su��:�)��&<]�I-,��A�m�ayB`Ġ�8vL�/�B3���򤘰� |@p�5ID*�s�����%&�Ѝ�f��JT�M��Q�lm�dD�{m&h�����@'�+t�Y�P�
��X���_9v��	52V%���
�⩣�']*v�铨ywmлpVT)6G��r�d ⦑��?q"�P�T�����D��r'�؆"R���EZ�Ze��Ato +up��'��h+�U��O�6 ��T1&r����M�>"y3�I3PÈ�!#_7]r:��$dM�|���OB��f�0]n(��`�B~lͳc��@V�',��9��WR�}2�#�6jH��/O^A�)Xoݦ@�o��gi��>���υ27F~�iVB�h��Ċ�+٤O��C�"OLT I�"ؤ,�AgAL�@W�E�G���=Op�dO�s�1�1O$'�	�z5�0%�[9QF
O��q@�8d!���-�t���N�@I �b��
�}y��9d	�:eP*,!4��=�`�뉔MeyBD�,Z>��ƛx����lU�"4e�! I�E&!�5�𱠠gI�,��\���H�bqO��@D�0Z�Y�'����SMC�d�̇_r����+A���S�ˁ��y��%/����(���#C�apL�b˛z?Q�F^�0����)�K2o<����ǂU^��0�|C䉱}�r#�&��e�7�֙
"�S�J�63�a��'��@ ��OU�Ez2i��!,<d�6 q�j$.�$��xĈ~��؄���r�Z�ȍ�	���A�I^Rp��	�ąpVoF0p�x!l� ����$�z ���� ���ױE�Ш�`�;w��a���}�!�Ɩq����A+U)@`�q��C�"#��'b�m�%��!&�`dE�T�V4�X�X�O
�)ր���a��ybH��{��"ۇw�N��D�i�p!�g }R)�<���!�D��ț!4���&ӸKJ�Ɠ)yt�%mC�kR�a�D�<`֧A�]�"D��f5�Ob����>N^ŸgB�,+p�\HW�'OZш�-(u�X�'~�q�范j0�`� �`��)�'��[�%V�o8 �퉡�h�Y�y⭉ �b�I#��7nn i�N�	iJ���Êd�B䉈p�]���Ē6�{T�UR7�:�I)�Q>�#�μjq93����̧��U rHЧ� >B��`�_^�̇�K���k�l?(0��8����ȓe�P����!K�X�  �I@d8��7JdmIbɐ88(�L0cJ�4hР�ȓ��*1�'r�����."Nȇȓd4PEZ�H>�m�Q��y�F���f�晫��)Z�咣�E�F�<9��&}H��"�]){%�	��Qr�<��
�c��� �)S�2��!���Hr�<Q���/`�Hd��O�s@�ћ�/U�<�OJ69�ѕ�E��(��Hz�<��A ��Er��8Dz1d�|�<J#e�d�5��>!�x}Z�)LB�<iW��{��=1�����|-Q�ȓ#L����ÅN*�1�Ũѕ!� �ȓ1�t���h�!i��)A��nILU�ȓ^}�lIAk�-_=�|(�fR�>��H�ȓf:V9{'b�9I�rX��@_�7��h��r4��o̊/��u	�����̄ȓv�8A&�,�d�s�� C`��ȓ�j�hׅ�'Q��j��Q�ȓR�X��h�0����,P���S�? ��%DH�6������!��m٣"O�p���"��d8r#��~��<�"OH�B�ʧJ���{b.a���"O���vGѤ"�jW
�����CO�<�w��k{V,�f�Ça��숇�H�<1ׯ3[�(y$�Q>��]�㦕F�<i���� �)��D�kgȍy�`KB�<9t�	:0�Z��s�Ƶ��ѓ�Lu�<��Ӕ/��t2��3m�bĸF�Jp�<���'lT�s3M��7X�E8�n�q�<��.B�-b��m5l��h�<��j�8]�Աsǎ
�up|�c�-k�����f��P$ڝ�f/�i��7(����ec��0D�|RC4\$�����K�u{��9D�p��Jؾ\��	̕��A��@;D��"q���6���ȾcZ���:D�ܑdb̍=&�hrT��63J�iE�7D��B���/	�pjv"��<�z�k��4D��8D@�nBx����
z�n|Q��&D���e��p㾵ئ��=|��H�Bo(D��c��j���"lA�_H"e���$D��`Ȍ�_�(TaO]
�җ)8D��:tKܤc�t�+��&���G,6D����t�Vu
5l�2a�|�B�8D��u���N@	9s	�)!��{��#�$��1�JMG�Č�; �~:��Jq8%���Ǟ,L>��P�N?��	��F>�`i��'}��IS�**@�j�G�K�`��U�G�D�4���"/}ܸ�>E��N(w�H� ��Hb0����ˍ|z��İ���a���Z;"Vؙ'
�r�f��")n���+J��*E�R��L<%?AKp)c�����E����J�+=|O\ &��m�=6���`�"G}�A� D���a�ВX�-��
ߚ^�4#U� D� ���8.���G�0X�6��b�3D��� S8 �ҍJX�8@��Չ}�rB�I(DT�����K��n��դT|��C�I�<*X��j��q.�I�'#��C�)yT�aH�x���HU
��pC�Ij���+������i���u��C�ɦA�vQ����K��`�.<-	hC�	�|���چb�Mm(�IsM] B�I����0DNC��q�(� Pp�C�	&'��q�f@�]�>�4`]�]�C䉙CO�� �G�&&z�C4 X(c�C�I[��8p#.��)��֦gdzC�	�/\`���l���YS��F/�B�I�7�} �U�(�r]�e�]�JB䉟X|A����\/x�7hDq��B�&��KQO�F��ّD �4Y�xC�	�s�`}+��O�Z����p.�)@C�	&(>�M�F��L65)2gJ�B�C�	2)�<� �E�
u�Di�h�C䉏2�%�e�.e���c"ʇ�B�ɟD�6ȸr��^$�C�#ͺe��B�	*�bfB�=����BƦ�B�	��6�r�j�Miv-J�L�)o�@C�	�D��T�QǰS�E�.ٜ��B�IY�����ߠ(�pI��X�6?�B�ɏw�輑C�JQZn[daە3A�B�ɢ`��s%гCA�1q�� LѨC�I �*$�A� -�8��c�ۿZG�C�F�	a���4[��	g��>��B���
u��'�l�pU��=�B�I3N# �hq�<��f�P�-C�ɵX���VB4b6��#����B�)� ణ7��,`���*��ޝI�zE(r"OV��`IW�1��k! �,�U"O�Hr"��
��\�׏�+1�>Iaf"O\��`E����#�J66�V���"O-��@���%�u�ɉ%���;�"O��iC�ʄsA>U�?�A�"O@�2(Y}j����lL�G(��"O�� �&2�]��+>]�| �%"O�A�����'�<��(D�� ���"O05��@9 ���ӓ���[�"O<)"��V����@�T7�X�"OX�%�P�PS��7�ؽ�	�'�.\YD�B|���"�Gl�ZL��'>z� .b�4���E�{ؐ��'���Y��A]���D 1
֠
�'"E�3�8C������uЪ�K	�'�Z�H���>yT%�"��o�JXs�'�lX��<hk�(���ζ/6^�9�'�nuҡ#ΰp���aB�,/7t�z�'��p��I��.+�Ɉ&� 0#�'\�q���/M����K����'�\��dA O �x���Ozp�'�=;���s�6A��M7c�L�ȓ(��Hsg�4���Cq�������C�dX��@K"���S�	u&Յ�=�%� ͂�9��Y6UTo����,��Lإ(Y�q��Xe�������j��"Ĉ�1��1`WC� |(��D�D=���+���z�GB�d]��N��I���)����(PP�ȓ-$�9����'P޼rU
ŷBlvՄȓ*��a���x�`��!ul���
8�1G�/$H��0t�E�#���ȓʦ��
�&�q e%��DNbԇ� ����Ҋ�9q_x�F�<)���<�b�#i�xwV�7*�;!N��t��|ГiEq�be�&
5[�2��^�d�!�L�T�23m�2?�-���F� ��Ⱦ'RŻ��߷E/d���4��-k�M>ny�a�o��'ɺ��ȓ_7~q)t���N���[��O��za����0;��I�v�H��A���>��^��g�'WeP�;��W����c�<i \<t��h��ݶuqK�,��B�ɪ)o� [�ծu�j���S/n��B�I�&�iq�ۑ@�(}HQɏ5QN�B�	�_�$T�� ׍J�R�[�j��wҴB�I�]�lJ��N��R��D�߱
,�B�	/ �
�{2�?Pxh����I4\
�B�I�Z2�Q�B��%���H�u��B�O��=	.ϰ7*�Ţ�b��4m�B�Iz�H�W�S�UDT�� O�>C�	:�xY
1#�Q$��A�¤_�C�ɥ
�H�2ǋ�4ytJ#-�'4JC�	�@֊���.\��������C�I�B�bJ�`C�y��D7,��C�I�W�ƥ���7��ܢ�ʁ�ZlC�I������嘾-�Z|����4e�RC�-#%.0a���3?���m��<(:C�ɑ?��IC������G?M�C�	G�p�� �ݥ�mS�2��C�I�]��L
�@#Y�,(���
]ބC�	�xn�=Ia�$jVq:U��Z�`C�	�
��'������Q#�B�)� ��z�*:xK�k�.ڟV�l���"O޸��%ĻY�� �tnܦaݎX "O�����%.�#�õ-z\�Bf"O8��d��F> *��֏^[6��W"O�`oԪs�ʐ�ᤞ�sV.!��"OpL"'$ƬK�\����͗<"tЛ�"O"X��܅Gqzv�Q�,6Q:�"O^��NM<!�h���A�� �$�r"O��rA�O�0��r� ��"OD�*"l16}$��*�i�����"O��2tM�OvT �F��ur�"O�!���p0��/G*��"O��JUA�xЉ&Lʬ[]��A�"O�d(�၀F�� Eˇ8X(�q"O�p�K������N�tհu"OfA�Q���)�JxB�R�I�p#_Q�<Y5��}��]�\�[����I�<�,<2r:����J�D��q	�F�<"	'O�����B�=�|#v	�A�<���Eg��t���9ZP���E�<�\y`~��@��>^ಬ���F!�čZ�����M�@��c/T��!򤈳rj�P@�L�T�VM���(Y�!�D� �h� �F:u.p�0�Kȵt!�!��#+��
��(���7n!�C�̌AՏ�]��q�v,U.Z!�$�3h_L��f�����ꖽ�!��׵_����ՇJ�C	�u���b>!�dU�Z�$�2� �(u�!��h��N�!�D؅Czr��22&�1Ƈ3=�!��M�S�x�3G�?O~�K2E?eu!��l΁�4-I�Aa�X8d]�xq!��Y4:Z�}��@��lX����B��=�!�$4&�*dV*��!P�⧢�/�!��N����� <N�$�� A=�!�D�$B��ҍ޺N%@��2l!�d�4A���Dl͎d>$��BE�O�!�ҏC5:p"�� ak�����!�=�&0Yb9}6��t�M�!�ݭ0���#я��I�D$'�!�R�(������y�.0��E�,!�0(N	�v/�J�h�V�ԂD!��_	��Aa@�=���2�4;:!��ƈ;�Z�����H��(c@@0!�d�%:hx[�埦\��Dp��-z*!��QUF�}A��3z�L��.�y!�$B�|�t� �<�r!�0M�9A�!�D
/[Rd�x0	D�&��2Q�Ɲ�!򄃗L�>�D�~���R)�3f�!�D�ia���J>!X���F�_;=o!�ޜlyl�$��5<���2p肬2�!��K�6������
)��9JG�1D!��L~�(�P�u
,i�`�g�!�dE���X��F� {G�أ��$�!�dX4�A{`ĊF$�F.�*�!���%�~�x��@0ta���:e]!�D �GY�飢j�g�lk����/6!�DF�J\d�� A� L�dK�O�!�䗒^��Z�ݔU����q�!�U�:�XPI�ÅgB|��
�$�!�d�s�n��ǀYu#Щ�Y���؋v�L��5�5�ܠ+ ����y�˒�wӪ�ziП3u<ݳ���!�y�ɗ�rQ`��� �)0Z
��S�Ƨ�y
� 쬊�朜Z�r�z��ɚ?
6��V"Op0C����LTyv�)2X
��4"O8�P3 зa]\��r�Ǥy�d-K�"O�$�tF�7;h�q����(M�uZ�"O��cIz�"0�W�o4$��E-*D��5➍B��ӂW��(ɛ��;D�p��V�/0�5�6�ʏNo\�Pd�:D�0G���7�xx��S�JN`��"�5D�P�^04���0ݖ�D��M2D�8(�+I8fk���b�,�&��A�!�dU(�6Y�M@�RO���7�%�!���<O8ِ'FоF۹e�:&�!�DN�C��g�$Q�!��B�V�!�$;Wh�.�|��K� M�!�Dױ�$��6�ݰ~���Ak\�$!�����ؠ��ل�J��O!�Ɛ=V�������$���@�#0!��P`FԿ�L)��f�)wN!�R�6:I��Cэ3͊�
��E7�!�]�}Ѽ�ʤ�����LQRH�b�<Q�IG�N�x��̒Z���@��E�<Q��,����r� +`����Az�<y��6@��d[�iÃAsFe@�F�n�<yg�	����fIV��!r�<yT�F� ~�}5�� BLt��g�U�<qTb�
Sr�����f�X���%�M�<��ߌs��Q��.\9I��Q�&@]T�<���[� m V�Է47����bZY�<iaߺqT�񈗪�U�s��S�<qg�m���`��&Ky]�A)�H�<�VN�+X��(KA�1��ʦ�IH�<�
|}:� V�摈"
G�<��f�Di�C��|�a�kx�<����y��{q��A��ՙ���X�<�愊���!w�O�q0e�Z�<qv�_�	�8���;/D��`aG@�<�F.J&�yɠoB	5�H�*�v�<ї-P 3f�rCK��!����Z�<�1�
:�B	��# bd�z���T�<���4a�\*�#]�r)0��dG�Q�<���S�g�@T�e��Y�LX(�� J�<��4 8  ��I��"y�*4j�
=�`d'?㞨zd#ي�(\*�(x�,�:���m���B��3,_�=س�"'�����M�(?�]�����<��)br�'uDY��GE�l0P�	�+§Q:���<(�p�ъπ�� ��y!H�?��Dz��L=�@��ȓ^���Pэ۴]붹�t[�i9�ɥO�ecU��6��O��p�E�!=��$��B.j����'{T�4�@���r��5Y����
�'*���'EŹ+̀qM0H\��
�'����Ʃ�T�|�kU�K���8%�\�n�nԄ��b+U��뜔>�����N�2a��ቷ_��Dƀm�h͘,j�j����#�K�V�B�,>�{C#D�\������v���Dh�bJ5��ӧ(�� ���2`��
)+g
��}Y�!r#"O�iÇ��!:]6XYC �ZM�Y(�jv�� �&��h��J5���S���I!h@�:c�л9���
�V��H�UML_���Ԥ�}8@ �uǍ[�Ό��I d�-Kp��7H����AE,���?a��A�9�8!r��2��_�M��p';�J��A xT!�D�/��lI1��-R�|p�aI�o^�I�,�\E0�'��S�OaN<C��>~te��
�1P�R��
�'N�0XQܭU�D�Sl��¢�,}�'X�8�9r���{�!M��Tqph[�@j�5k4/K��?YӁ͌��XaDXM�b��J���@���D���d^�1[6����Nle !�.�ax�i�>^U�d:p�|r�=M@<����ӷwʄ�P��y2#�i6Pâ���	���j����	'Dj5r1��ɒH00py�LƻFʑå��7!�@��lDS��H;Q�U)���$�!���0&���\�_�Xy����q!��2NZI����YT(���+п*/!�$"F�&��P��yBP���hZm!�ă+=�n�h��ɤg��)���K�!�D��UV�J?��s0��s!�Z����Ε�	m��RTkV�!� r�8��3��+,B.�j���7A�!��+d��5�nY�9F���FK�_!�D�r�Ly"��:m1��!�lO ?l!�D�<j���Qe�.�P:�l:!��F�V��l8��S�ߺpP&ʙL!򤑸���dAw�V�*���/ !�D۲Y~��
�|���q�υg'!�d�+B��Y1A��a�x�(�,!�ĝ� ����#c�*�2tL�3>�!�d�R$���L�lpj I��X��!�DA-�и�o�BwZ$�� �%1�!�,oHUK�ɚ:H0VX��L�Hr!�$Y*1��pq�䗃h'ʭ��g!��`Ԗl�&��$I�����C�*A!�ˑ@��wO�6�X H��=!��+y<]EI�=�Q��D�F!�	�H�4y�r�"B�1�@KT"!�	���e��*�9�@#�-D!��
F���(u��zߦ��C�L�:D!��S�l:�p���k��#5��<!��HL���R>0�ّ�.>!�$P>+2V4�a�C�?����L>$+!�d;Q��`���ݢ/�B ���6i�!�M�SR\=3@�&̀��5&��]�!�֓��I@��$����E��F�!��SW`p*1�ɱB���
:�!��[
C�E�����(��1�ɂ_h!�d�Ő�	�i�`pV8s1d�#]!���Op6��tE��KJDy�'B�-bi!�䗷^��x�+�>6�qQA@9i#!�dE�M�@���)�+��q���d#!�WD��Т��e�����ơ5!�dM*2��l��m�Qu����a"O��+P�,�
��Uf\�J�r��"Op�(�=��#������T"O����4�0<s���t4�Ч"O����Β]츃g��l�F"C"O2B#
j�A�p�5/�����"O2�FZ�(:L;EL��!�r��"O�@��e&,D� ��L/#�б&"O�40�c�U7j9��kR�H��U�"O$i:��
è�	�&S\<J!�� ��xc	Nn��3M�#`��"O,��D$� y�cfćY@"���"O��{%�ӲP��9A3�͇"O�"OZQ%T��4���U�W��]��"Oι
�*	 �ؼ�	��J�Z�8�"OF�١I)�p![�h��
R�u["O���V��.��@���N
3{Ё�"O0!`E�;��c�*ypΝ "O(�
5�Q�f]H��slЏ � ��"O��H$��R��	�K�-K!|�Ss4O �;�L������(�g��H���AJ�!*8��F"Ox���n^3젤
²X�i �_�LX�#ҫ
�f��I�K���3Ñ�i=�c-�~������<�d��	\?!ApqHƃԋ>�bl
��ڻ3�B�
�'�\�ī�7�2�`Ġ�|r:���аl:A��)
��O�8PRDOۡgH� S�����KBh�<�Ӯ�*`bEZD���	�@��GM�䦝�"EM�N�\H�>E��4�� :R����8�AOէ$���~��{0��:In�42B������'e�U"�E�?RT`���
	#��J�8�� k��#����՘;L�!���!{0d:w�Ć!�ܑ�Wa�d-Ԕ��'^����&{6@˲��(5��D#��dZ�,������Ӽ��OY��B%"P�cK\|�1+T#�T��'�X�!F+$?�I ���P�H��۴�.�EdƳ
>ӧ���F��{��X(�A0E28i�\=�yb��O0����ޘgf�p�W����D�S��c�EK���<0(T/Ki�ȫ ��,,U؛��V~X��gi,
��i�Z�]CďF�T�˧*�`��񤏥�4S'"�D���VQ)P�ў@�#I�5�ЍD�D�ĭPƮ)a�"G���t�Ī@�y�⃿, ��%�y9�@��%Ȩ�y�ˁ]�E�=E��S�t*��E�wq@�0�� �yrc�.��� �� dL�E
"��y��	�k6dxQJ��eV�y2a�D��y�'ˤL&�U u��4\�ތ
LK�y�ҏ:wN��&͔P)r ����1�y�PAFQ#@)7J����t��y�bG�m���-D(�'nƹ�y�-X�9 �&�?�
,�G�.�y�N�Z�Pub��AKz�cX��y��Ѻ<�:�
a@�*>��,qCi���y2	�!� ����42벀�gn@&�y��>��ܛ�F��&#�ia�d�%�y2l�J6�-`@�߻�����ߧ�y��C
j������=A��4�5�U-�yr�ͻ_��)'*<�\0��	� �yeΣ�6���%�(�`��C�=�y"@��Z�qrU�=)�LHHSL���y�B�h��<{����`8b���y�I���B�r�f-l�b�5���y�H
L6�0�p��"�1�R�Px2I�&��402H�d���#�O��� ��"q�pI�ъ?кM��Qo�3�	K��� ,�0g\����F&ː��DO bt�-�R��Ox8y֬ϤM�~�Y�F<+%>�ڰ�,F0�����O6ȓBèپ���@v<�6!Z�!�v$E�a�剄idX@�Ț���]"@B�BG�Y����v��q��$ �nS!<9$�@���r ��+�!��U�7I(�i�W'y��3(8T�TAQ���b�d]҇`��:���C5�ԗ3O ��'���I4E��yG��5;Q��a��S��̑�C!�2"�$nz�m�V��	����P���6�f�1�glN��(��+� �;3�V2~�]�&$�����>Q���AyȀ�@*A�2k���zh��|�AG�?i3���h@aB�"`�)��7(�&�1�eʻg68IQ��.#�����RWV����R��a{2!��}ɨ��A!�-���	���V���,
8�M�2��SF6]�+y����Q!7.�ذidS�R�ݸU$�@���I�9	�<!�'��V���;� ��U��T�	�q3h��bĤ �J%�"(Q�I(xz��\$RdZ�/T�)�U��ყt;d��O�EQ4�[&
�� �����Ӎ&N�a���u���|�kS�FƏ�ZH��̹���7@�(���9ZL@'�
� ��yycD��
T���䁀w��pi�1J� � ����'����G�NXځ �hΥS���c/OGu�4�,OJ5��� �i#,ҕp*���U!+������	m��+��K�.N؁� � ����F���Gr�dۢ�]x؞8"��ә&��`űU�tL*a�R�p�.����,	N$;��� �;שR 
�� ��V�z6mP%��DNOU��!%�մ/���[1����<1u
U�)���;�F��y�kM���G�؉-�p)�@��f��`�����<�"��
j^<r�+G��!ܨP�<�1�rA�#������,Ph$qA�|�\(Z|!�$�2.�K�bU�rq$�	>���!NJU���׭Gd0����>���� f�j�(2��i�,Dz�#��b#���ҏ�6���.�%u=�ʓ�~$��O���`s�	b��'��0�
�2R����+�b<K��Z�A��83��'T��_6���J�&�%�ք��	(��B^+��lz�B�ɼ#SVM�Dú��ɼRϐ �N�p��<+������&9���>1��ưkp�b� �GY�u��e�E��:9��x���J�	D�?I�G,�fǜ�h�,�}5xi��?D��FGɐ[{2�9�A
�Lg8=R�!��ks��O�dB�B}�g�	���#��5?��$´�J.+�C��(���P�B�6~�o�!^�{Eh�  �B��'U�8ɴ��BHB��*�KZI˓���r�Հ4��ʓz
h%f�
�r�p�"��Nu��ȓ� ��Qh�e@h8p�A�k�\x$��X�D�)6�&��p���y
�!/�?&���I�c̀CA$B�Ɇt"�]H�B�4��9e�MIi \W�_E���+��p�~&��V��"�����Ͳi��JG�>$��K�G�)a���b��*(���Q���|~ԵB���(T�}��FL�\h:f	Y,+�6E�p�D�<�Tl�3[QTu� ��<�����g��a��
H��dr�v�<�c �'R� �����}1L������I�|5F��㭎>����<v%�����!��Q�P�;D���N^ ���G^-T��#��[�qOr �1�3?���պB���h�KU!J�2�q�l�o�<��(S�S��q�$��!�P�y�`�c�<r��
(c ɰ�l�M4�1�
Rc�<��$��=;д�UhG�qa�Ei�G�c�<�!�ިG����	H�dE���p�<�7���j�´*�k++�P��jGo�<����"�9�B;!��dB�Mh�<�ae6G�v�bG@�P����	�i�<�B(Ry*��6%q�	V�k�<!�����A��6y`|�2`�O�/S��a %�'2']ÁׯE�<���K�9����vH�ik����I�l,0�\+j�RPAׄݷD�OPXE��O^�+��T�|v5�1��f�.�YC
O��&�~L�b����#Aj p��L�	b���W!D�E� q1
� Jl�ඉ�7�p\ӏ�	~ �I�L<�A�#B�{^X�30�d��F�Ȝw;�	2���v�FE%D�8��@F�;⪔��[��BW�<�r.��7b����\�5Dj$���i�|�
xt$X 14ȃ7k@!��+nj����>>��]p��/K���f��=�B�Z3d�P���{�U�?j��P���e���"@J��?��hջ9���{��n�~�*��=/��PpĬ�8t�f0��Ǯ�0>y�᝼3]逑́�33�\��f�T�'��hd�G5�����ÛGP���"��9�����F�R;!�ā.|+dM�M�629��ycΎp>�ɴ���Ȧ���:<��@�K�J�OW.�r�:$�-s ��e�i�'�d�Q�)��i���C.zs.A�H'����y�2�����gܓe���w�>���NE���%��	�d��h0��/�D�i4���.�	[���4T}���Ga}��T�`�����GY���&��0<a�NH�g;J��H>��K�N�1d�(���#V�g�<�$FŧP��|9��P�<|�ƅ[K���{ �z�{��Ti�1|�"� �8}��8h�-M��y"���,P��	4��t� Pҥn���yB.�1����Gm��k(�� E
��Px��	X�? ��C�A���aw�����%	.8�!�D�#��@��̈́J�����S/ax�#6i,DB�|��[����ǡ�)D�Tܺs��7�y�*P�-�NL��_�2�U�������}/�d`6)J
��)�'Q��SR�"k.���V�N�>e�<��W ��	�f��> �	ׅ�U<S%�>Rn�8�X
N~�=�K-D"��f�C��V#�*���B=[�p5�I��r���@ ��,/���pA *�
|;��Z��*ea,Ɇy�tQ��F�'w�����!�a$>�I��m}V�zd/���Mbt��~�<��Z"[�J�r��:9zx�H�i�]yk��{��رՂIg�哠	�Ś6�@�jo�}�F�޳>2C�	D�a�蟔C�nY�/��J0|�'����7.�|��ϸ'th��'�1)��U��-r^����Ovb��t	]2{�
�qu��
�VAB�i�G��=�g� �O� �	�,&ɑ`�C<c�F�rr�'�b��`��'D��j��)#�\*$!B�X�Y��'����0��$2v�s�bŐkZJ��I��
��E� �qO�&0x���u�dlS Ay���"O�$���%)��Q��\�8mr�!�"O��1��ƸP��Dё�b!�A�!�d�U^H�& K>B��T����/*!�D�,���3̔�7�"�t��{
!���-oR�!��9`�L�x�J(k�!��V sC������ Qݜ�ۂ��48�!���=k�^���!�����f�I�!��WG�rTb4��!�
X�祜�!��s�t��7MI;;��R��H�*w!��N(m��ԠT�5}OPuQRk�0o!�Q+�H����~��ì��H!�d:�~h"��G5P��U)���"1!��Dm��;`��/a���!OY�!�ԯ@Äiq쟼3,M�ĩ D�!�D͖8��͛�"ɚv�@	����L�!�D�l3�q��+z�(�W�!{d!�$�WI�H ��6ib�8Z���#|�!��E�k����dC\ b�*��s�!��]nξ=��D��.��gɏJ!��	�Xm���hȘ4�J��g�ب
�!��+��O(f� K�@ �!�d> ��,�c�88��Uڣ�	�eq!��}ހ�`�*B7%D�Uw�ɥ!��1�h����Q�mȭ
�!�܇:Q
��c�^)_iR���BB�]�!�F�%�6i[f���cNT��!�=[p!���^@ā`Az�Pp���@ ��6�(�\X���'�<q⃄�8�̑Po�69��ڴNB~��ֹ+��ȟj��ဇ{Q��ad՚�H��V=q|��;?���)�F����.tF�!��X��kD~�,Ք'`�[�QP>�� 	מ
�����K@�<���"�	���� hz ғ�L>�ǦܮLåa�0��Q��>a�@Z����A�8�~�'�Z��V�L1j�X�E�p�T���=n�� �F΅P�)�'J��c �I��YCv�T1vlq���[��`[�x�ՙ���:��'	�Zmk'*WqU4��጖��y�@��6v�p�͓�j���o1�������Q���g@�{ʨ9�cJ�|�����|�����?a�D���8���:9#J�5��"H��S�`���#�D�^�x-z�'�BA�7޺&fE�j�^��spT4{��3pB4k��	�E��X�RQ��,�<U��j�z5H�1�U����*��s���G�T�B1�����P�����0��F�]�q0���cI��� A)-o���}<��IzO~���.��xd�O�bUŸ#��M�ӵi!F0��А�8:�1��P���	��%��(iR�^�eL@�UJصY=pʚҧ�6ہ+Uo}��M�i�b��;OP1�Ƈ�*AO���N�"~b��ft+td·Vj�c��@�v�x�qfW1BF�ҧ�g�i>��I5l��*�WW�Р��Y_�0YK<Iu�C����h�g�? �`aΔ�(&���ͮd��Ia�J~b+C]
��;�"���SČ-U�D�sO_'�l��]�l��{�h<yu#7?�|��'�|�0�-�6++�d�&��	V�@�*۴��a�vE�,�F�1��WZd��D�d�]+Y��Y�i�0w`d����ڜ)'ر��jޥ���I�M�ɑ
ç!#����ږk� j"�`*T�ȓH@�eڑˉ:F�!E�F}�̆�E.Q*Tk�(�҈Q�n/�����.2�ޝ؀��Z)� B�>�!��ǣ]Hn�a�G�8L�~�
P�R!�HI�M;V( �}o��`!φ�Y�!��N$��Ey�����^-S�Ά#�!�3V-�,�uG߁o�h���f�!���X041d��&|H� K�%T!)�!�ć�^�䂅 )<$�p�i��o/!��0r��$Ж+G�h<x)�*D�} !�#� e获8D��k�6P7!�DJ�U	���-<%��xd+�BQ!��GApUC�(�2MU�7�K*@!���A�$�#��2�q�	ƍw>!�J�)a&�ӥĊw�t���N��!�$�?l���ro8C� D�J4�!�d*Uwr(&�Ӛ/4�0�h�@J!��W�!+Z='�H!�B>!�<AQf�B�LL<X�a�3m!�$�^dF<;��A�s4���UNJ�P�!��3����֯G�%���u뒹E�!�$��n�.QR�ӆ}�b�+S)!��9T��B�߰@�̸��7�!�d	�b��P�]�}�S��ͤ�!�d��Z�(��e� xleT�Y�7�!�Ą�w�H��"jrx�T��T!���	���3%�1$W\�ٴ�&I!�X (��]Ʉe�).�8��8L!�,^�%*�B	 m�(r��#�!�ڮ"Ĳu sBܪC��P ����2!�I�w�ɲ�!����#<d!�$�'���
�s2L}�f?G!��DL�t"p91�:!�Ao�n>!�� #u�]ّFY�S�����֯dF!���j"�� *.$�"��6C�3!�D�4b@}xGb�&o��h�'#ߙ5(!�dT�@|`@��Ӽxg�i��|!�D�V��R0�1�t샲�J8!�d�4��!o�"�8x �ꒈ�!�$����(������"�Is��=�!��!
¸�o�#~��w���Nb!�2���H�E�$i1ׄX9{�!�\zr�Z��H( ��ܩ�CLl�!��@x�qY� �;��@H�ԪaK!��G�:��`i6�����ђ(�:O�!�$�,S��C��ءB�`19fh�:�!��%Z0�m��j��JN�٩���?^�!�d�m�8[Ɔ;��j�&�+.'!��T��k�==����)�8�	�'�am�>0hd`9�^x�'#�8�C��B��C�U	9�L`1�'�X��u���K��h���"� �c�'C�ĸ!L��8���3��]�-��'I����M� ���r��an�H��' ���GL�@s��3M���	�'M,�x����2)��Ҙ3�|:
�'�@]I�Ώ�6C�1c���!
�'	�=�EfֱV�T��T�(���	�'�^t��(?�p[�Iӱ������ x�@���[a��t��'�%څ"O�MbVDP�Y�ӰKGڎ���"O���Rŏ z&�P`s�Q�|�8���"O��`A

����A�D�	��"O&K��H�"N4B��(t�[�"O4�Pđ4#j�� ��$Z�ؓ"O$J���+Ni���ED`v�bU"O�Yd�ɢV��Q9o�6wRu8G"O��7iS���(p2��)PG�5#�"O��3!�89��n;�$8G"Od��qE��Y��`1D�,TM"$"O�lS@jU�Q��qq
y�^��D"O:�;���KX��)a�R�&U�(��"O�� ��և
�.!���1'[  2�"O�aS��H,����םk��M��"O��h䭁7���Pgǁ5%4<Q�q"OB�k�r��S�Hͷ"+�qs�"O`$�u)��k�*a�B���P�*O\帔hԐ]��Ͳ�M�l�0e�'2:Y`#�M��]آm֜R�$m1�'U��#­�V�"U0e�K;J�] �'"�;f�؟ar��G�.67T���'�J�Q�3a?X�Q��V�|���'�>u�%A�����|>H0
�'�I�B�"mۤ�.=pf��Y�'S�is����F̂�ц��	34)�'4��w��oݞLif��\��*�'<�����N�G�Q;sG��Y�Ց
�'ʞ{���<]�b�#����g?T8`
�'B��	�^F��A!���LPA	�'T2�
�6#�ؑkʴy�	�'�B�Y;#��!h㙆P2u�'s�%��'N�
W�K1`ڐgZ�[
�'��EB�%o�2�p1HӴ
$jTS	�'��	�E��(�� F/ғ}�>�b�'a9Xg�K\}�(�t��q��'v��b@֟l���[��A�e���
�'�,@�m Vz���T�nd
�'7�����H�c�f������o����'���4#)X��� ӬГy��r�'���BG�O2,��2��j\H9
�'��Уbˆw�,�I��˃fU���	�'��[��Ҷ.\���
��
�'b���	�1�|m{d�����!
�'����,ƨ�1�$�0z�X�	�'��8%��Z��$zaN�x/��@�'�+cm���t AP摌C��q�'^d�D�4tY�I��ܜ=�� �'j�����?�$ta��-5��]2
�'�f�3���0T�Z��Y�1�*܂	�'8Z(c�Y3T��scפ^�p��'��l�Ê�YZ#b�X4ܬ��'��hPW�Z�~ @��R�J*O���"�'X��$թ&(0���C�"�k�'Q�)a��\�&�����Lq��''�!!'K��m���x�V,��'�.��'�j�
��t`E�o���"�'��tQ��7w�P �*���VY��'�
=R&ㅿ���;��%v� ��'zNy�/��`0t�R�C�~2e9�'ۢx��O(-&}z��
�Ƽ`S"O
|�EoȩF���YH�9!�T
/�!�d�|�D�"�\� e	�f��>!�D5}�\x�Be��r\�� �fN�-2!�� 4`��Ȋ�?�J4�D�Ì>g���"OB�f���{�Ə�hT�h;""O�4a�ҭ T�AKa�Q�nf1#F"O&H���ğ=٠3��K5rI���"O ���Phy�h2��9*f��"O�,��k�%a�&�l'���"O4��4��#mH ��-�P}	�"Ol�+Q�1��$`��@^�LȠ�"OF䈓ℭ[0x��Q44���"O%ǝ�t�AQd���[�*�i'"O޸(Ӆ��%��	6KФU� �#"O�ti��;}�J�qd�R�H$�"O��K��Č!cJѐ2��!4	�4"O�r�L��:�n\��	-�\	�"O�҃GC:rmz� ���\��a"O��ڒ�J�Ќ��JC�"��"O
�
r��[����ANcn��"O�$�vn���2d����Qav�*#"O�U(�,]?|](d��OA#�\H�"O���T��lBD����-���"O.�ڤ�
Sz��E��"v,l�;�"OJ��f	�3A�K���j���j'"O��p�g��$"⅒qeV>�"��c"O@ � �E5iLԡr�d�]Q��� "O� �V��M���<O�a9�"O�px� 	�|�9�PL�U�R"O8[!��[¬x6M�m�Z��q"O����O�T8�X:�ŉ3�8=�A"Ox���Ll���:p�($x���"O�b�Q�V#Ux1�H#8eb�;b"O�CV�_<޼�+�ǟ!]dĈ�"O��*�苄)��hRF�0hj�*4"O�� Y�7�<)���dF�4�"O���o�~�$��`l�/P�"u"O�M��IF.q� @��l*���T"O�ma�e24^$���\�x�"�I"O­�Sf�f�ʅ���;��:U"O� �!��W�qˣ��62���ȡ"O+O�&D��m��I65� 1�N�<q���" I�4g�����Q�<�&�)|3���c�u�`�RAJI�<���Ր;z�X�A�;.^ �� OC�<�v���2Δ�a >?��#�Kd�<�W��<b���AѨ�8c�� "墍\�<y#B�.)r8 +��A�%h.I9u%�[�<	��Fr�mB��ð2�(`�F̋Y�<u�**�걃�+�+v�x�2w'�I�<��b�LXP�Q
S�0�>ڧ�VO�<��Lzܶ8jTLDB��2�L�q�<1A���gS���'��V�<e�bh�y�<���(
����wN�xZ6Kv�<���ߣ:����'
��<�!`�t�<��A ~0�$#CfJN��6&	w�<J�9�&��%O�uw"��GdH�<�&�U+N�(���>	��d�K�<��h͍tR��F�>Ke��8G��~�<��S��`�Q�,��
�*)�G��w�<Q�+�(&�؀��ش�ڜ��q�<��j�^�l�J��O(�%C�D�<���-٬#&T�1��5��D�<������A��C��}��mB}�<1e��ma���5Δ �P�y�<A�3/ń�I��u�K4�LD��C�	Ql�42�$_�h�D��vC�)� �*�/�,?L�⃄�=���"O�$��Ɣ�K���V♚:�:*c"O����C���!^J��i��"O��2vM7i:į�N�P-ð"O�*0��O�j@�n�0S�h�x�"O�\�' �X�i���6_���a"O�S������K��M8b��,҄"O���b�@�z!Yď� ��@��"O��G   ��   �  B  �  �  *  q5  �@  L  �W  �b  n  �x    �  x�  ��  
�  N�  ��  Ӱ  "�  ~�  ��  ]�  ��  "�  ��  �  N�  ��  ��  ��  w �
 � � �# �, -6 �= D HJ �P �P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'��O��P�]�۴$G��d�q%"O����bN�#K��X	0�O�#�yԮ���v+T�4z��s�����yR"?�EP���2.�R	��%z�=E��\Ȭ i��3Qlh׮�	.���<
�<����$�`�(��@�ȓ|�<��TL
!��qC!o2䭄ȓ~��s�X�\]��9�E���F�<I��^�C�}�R��-�h�J�L}�<�A0ho��+��ݐ%�]bUC�^�<���ɸ{�Z\y���6a.�Qe�Oq�<1t
���A�G��J5�-�3�o�<q��w����EQ�*@�p�S�<Qa�,��ms��Q$i�QzREY�<9�����A�Ђ8�3��R�<nM7w�jǁ\ۦ5#�E�N�<yt�g�zQ�EcKU�Z����q�<sK
 1rT�h�$��B�O�l�<!$�x�Z���U�����M�<�V�h1�\� .jV�S �G�<i��8�V�+s"[,hn��UaE�<��_�P�S��$t`�(;���J�<a�C*!�$�r4�KZt��҃�Q�<eب)����.��{3�����P�<A��]D"A�Di;c��%�ЩCM�<�B�<.�j�D�g���RbaDL�<��!İ<0��i�H�k�x�$�Q�<	�mO�
a2�*kC���[3n�H�<q�M&eP�(Q��^� ��%&͛]�<Aԇgގ�Ƞ��$~�$���s�<!�H�E��q�4�
,g�<	�c�q�<#Դ
���(d*�E�VD�9�!��6x<y�&F�(9&P��G�!�D�;(G�̨#`H�4�=�� �!�� 
%���J�]���"����"��,�u��k�O�m2�gӝY��Y�s��A�h�
�'�0	p�ˊ�F��0a¥�;[`�'Y`!��N<�lh!��5dbh0�'�,P	ĩ�$1:�p�0�Y�'����yB�'S:�H�Ļ9f`	:̘�s�0��'j�)⃬?m�F�h��
�|?V9��'��qz�aT<1��:p�A�CO��	�'�+�Ë�~'�$���;�zL"
�'��Ə�|��L9�H�7n�)	�'|RD1WA˞_@jy2�$�+�Ib�'�n�*̇�<����P�R9!%� q�'q��siW�R��´��Fd����'�i��xg\��4�<@�rl�
�'HQ�Rf}�>L�3BǨJ<��	�'{ȕ`7�W]< �;Cl�����B�'A�	��S1[p�i!F+0B���
�'� Თ�ə	�:��5Kڲqp�]b
�' ��A�(�.l�<m2��:o�0̘�'��`��GP	����B����)�'°HA��E����B�P�|p�y
�'�b�(t�b&]q���C����C(D�ph���jz T�V��pe���2D��q��T�Z��)Β��uaw�1D������v�ز��ˊXkĉ��.D��"�%D�wE���0kɊE�¥�!�'D��sfl�6�Z$��n�c����Ո!D�x��(U�!�2q��͵6�b9Z�#D�t��,ǨSY0�C'�L�P��5D�ș������][�᜴|�!
��3D����_\愚g�*}�*��*O���$�wX����F�.m�rA��"O�'ڱWy8��䯓<tf$�"OP�[��A0r����M^((CA"O|�:�%�4/:y�g��*A����"OZy꣪�2���J7@w@u�"O�x�© ��ic�ݴ>5\0�P"On` 쑺l�Ȅ��eގ,{�)��"O�YbW��g�2K"E�9P�"OX�ɠ���?�p#��Z�iA��"O\L�E���7������ݙa�, ��"O�Y�bEچ)a�)
5/� � �ZT"OD�Qt�Y.m��x�c��?HK��Ѷ"Ox��W��KKp,�Ȅ#8;6M�"O�a���2�64J�E��xB�"OH� �c��5�Ҹ5PĤ<9�"O��	''N�E����	����6"O��p�3��!c�枠E����G"O�uf �F�{���w���"O�,8�37�ڵcg�"rx%3�"O�����Ь��o�4-gP1�"Od4x��L�t��hC)�E��!w"O1rnZ?}y.��0���+�"OЀ��F�zCέ������A�g"O.�Q3��%L���ʒ%�NEҵ"O.��K����M.��pa7"O�h0'×8x�kgiE?���8b"O�����Ɏ/H�� �Ֆ$��S"Of�5cI�p�(T�v�؜^��"Omx����scH�q mA6W��H"O^��@'D-lX,�!�ɡ:\NU�6"O��"��;�}5*ӃA+����"OV�
Ԣѹ���1'!
N�"O��`��#��eۇO@� h�`"O� d����Q:W�ޭx�M[�:P`��"O����1�n�P֬�>r1zB�"O��s���یq؇	3{"~���"Ot�{�J�%��A��zB��"OZ9�&k/u��hZ��J�;� ���'���'���'���'�b�'�B�'�:�+�$&�Q���[1@�����'/��'���'ib�'��'B�'!�`���FH�,@��GJ#w��7C2�'�R�'�B�'�b�'H2�'I�.ٶBc� �"0Z�5$퓇���'7�'���'y��'��'�"G[�g��}y�O�}4�ZJO�I���'���'�b�'���'B��'�bϋ:0+� ZA��+�d�穎����'Y��'���'"�'�B�'���B�*��h��^'
J��j�!6�'B��'��'���'!��'@2O��c-f�RK�5��H+v�(�R�'�2�'�B�'PB�'���'���Y��@IY����F�,:�R�'�"�'1��'0r�'_��'��C�@! ٓU팦n\�0�싗8_��'�r�'���';2�'J��'U�٥K��
�c�'_Q��ka�7\?��'��'���'���'g��'5L�Mx|���
z4`�	T�r�r�'s��'�R�'b��'�'��&��ȴi'Ζ�M�ZG��
�B�'��'���'���'��6��O^���FM4\jb���';"�� +�=�T�'?W�b>�7����-���Hf�
t��P�G�x� Y��O��mZY��|��?q��޴.Ԯ� �2?�(��g�8�?A�����4���h>M2�����M)��c-�9[eH �$�5{y�c���uy��ӠD�������x�������*�4ZE���<����f��.�.�j��CE>Ό�i猈[�����O~�Y}��t�3sy��6O�CdF�}t�Đq�ޜn�X��?O��	��?�&�%��|�Lp�Y���ކ@�Y�4��3i��p����3����E���"�6���ċZ)0���.���pl�?�RS���I���͓��\5h&�[�N��ĉ��+R���p�e#�!4Vc>q�u�'W����xo��b���s��Xf(�/r|�|�'r���"~Γ��H+3��" ܊�A�I�	/�*��/�����dH��}�?�'RpЬ��#=Jq.��秊� ��Γ�?���?�s�^��M��O��,�J��&$^"�s�`�% W Q�� ��PܒO(��|z��?Q���?���7�DZ��W���փ�RiN��+O(9o-�2Y��mޟ��	�?�6
�ԟ��I�~�!�� .���Β� llB�Ox��(�i>�����Õ�@̾�ۡ��x6����Q�_����iy�n>Dz%�	�G��'�	�n��Y�T%��x)�lC�b�
i�t�IƟ�����4�i>Ŕ'��6��ttx�D����ѥI�Bk׿0�C�c�Of�m�R��+q��ޟ`�Iԟ����;V�¹iY�����ކ"�`�[b�����'� �e�?u
g��d�w��P1���"uR�@�P�Z.n�쁙'���'=B�'�R�'J����hVy=���o
9&�Ɛ�B��Od���O� oھL�J�'s����|2 �p6��S�c a ����&U�w�'�����D'�3i�&�� � \�7�|@�cI";E =����Hl�r��'1� &�������'�r�'�ֽ�Ȓ��z<-Sz�h��$)�?����dئ9��c���l�I�d�O�0��n�/�0"r,R<m(���O<y�'-��'�ɧ�I�':�Pmp��/�$t��	=A>fx2�C �6q�����@>�%�D�w�:���.T.`�Z �B?n.���Iߟ������)�sy�`x��Ńs%]5n,�,C�X	��!J���ų�^��Sݴ��'�X��?Մ�6RA@q�u�E��B��$	����3wD�Ѧ�u����+���
iy�h
\�,l8�(K>s]�$��i��y2Z�p�	�,�	�0��ڟ`�OG��9c��5a�q��'WI�hԇl�B��V�q@��D�O�ʧ�?����?ͻ'�&QS1k���ǧ��n:�{��?�I>ͧ�?���=ZP�ܴ�yR͂	nW�p9Ao99�x��d.�yb���T������4�<�z�4���	�hNs'��<$�$�O�4�?�.O�pn��E#Ҹ����4��9��ِ�ؙ8 e���>q��?1�W�����$�l{�F		�4����\44�}
��7?)�CK���9�Ā[�'������?a2��e(�
"�d�����?����?a��?�����O���nG�v��K�E:Y�ĄJ%�O tn4|��'	�7- �i�5Y���'�r ku�F�@<���w@z���	ҟ���7��)l\~r#�g��	�5P��(�%}��s��	���h��|�\��S�x�I����ʟ\J���,n`!���oP^���vy"�y�x)��O����O���󄔷07>���
T�)^N�9��Fd��a�'@r��I*Q��b�n�hR��9A��ɯbGެh)O�a��Ĉ��?Q��,�D�<Y��H���m���[��Y�+S��?I��?���?�'����8��ß�HwMƔpX<�-��Z0�U4�T�������?�^�(�	[y�l�L�@髒��/YNRQ��FH�a!4�i���!��e�O��D%?-�=� n�#�T+�m�E�<*�T�I�;OB���O.���O����O �?��h�`H��Q�B�f�T�qu��Iܟ���4rL��*O��o�K�	%S>u���F��IT�Ӿ-�@c���	ȟ��IGh�lZ�<���6J�|
�>D�|9i��GuN "��,W�P�d������Op���O8��X� q�����5��!�a�I�Q�����>ʓ:%����8���'�RT>��� �Zk0l��k��WN�$� Mc����^y��'R�|�OT�`@�R�T�B��;��� ��tE�(E�./�8�O���L��?�q�!�$_;���i'�]8O2Rm��c_�B���d�O����O���	�<V�i����e)R?ht�(�4"�., G�۪X��I%�Mی�>���>�z� V/R3R(�c�e��n�d���?%�?�M��O�nY3X*��)����$��$�V4��jF,g��4�� Jn�$�<���?���?9��?)*���KC�|��{��Ϝ|Ш(�n�>�<x�	ޟ`�	\�Sޟ������5��
C��<PV�C����:�?1���S�'7[j]��4�y"BQ?�h1���U�ΥUW��ϓ�v-ON�D<�Į<��?a�+�n|(gɔ9�p��MH��?I��?a���d�Φ���˟���⟴�wC�aVplP�"�;G�d���j����I�����z��	l�P�mހ~�q0�@�(� ���0���X�|: +�OLS��ݠɛf���4K��
�c	D�Jh����?a���?i����yŸm���?1�iۜ%�d��d������"ݯ�?�3�ig�u��Q��I\�I՟�]?mn�Z&#҃ZG��
���p��	�������x�a@���̓�?���:=����=�ZX�l�N��l�O��"/��'�x�����'b�'�"�'~����#H�B�i�5�/yd�+�S��P޴	)4����?�����)�Ob�$�36�8�� @ȶk��Œ���9N��?����|����?)%(�'[�dԨC[��R��]8f���0�Gy~�F_�p������rt�'��ɪv�.	�$L�r����Z�w�>��	ş0��� �i>q�'��7�ǛGP�M�7Y��ӷD4
i�-;������������?�R^��	ǟ��I�N$�*`LD�o~�8Z���f�0 ш_����'_��z���I�O#G�S.&��&��;�d�$��.�y��'|��'b�'�2�i�?4�,�J�(	�ʹ(�M�<q�\��O@������qUkp>I�	�M�N>�r[iM(6��5%����!����?���|se ��M3�O�\��A/uX�١�/,rqѳk�Cs����'��'��I���	���I�t�M:S�9)E|�Q�T�U��������'�j6�^3)θ�d�O��D�|�7j�v�PG�*+b
4�Ip~"g�>	��?H>�O�VL�#v44:u��S��M�Gb���Q�醊S���|:���O�5�H>Q#��{�|���"{*$[�._&�?����?���?�|2.O2d�Ӆf< �xW!�4p���+Z�!h�1`҃�<��i��O���'�2�WV���@$-�}td]�qگ`�B�'�F<	�i��iݹAdl�?u��\�����`�P�Y�~�Nؠ�$s���'�B�'���'G��'��Y�������P*̰�� �s>9��4�������?�����O^�7=�`�q�ÞC�| �支v*X��R
�O��b>i"�Eަ��F��c�5{�^9i c�b>p Γ��Q�7N�ÖhL>�/O�d�O
L8ckΏ �$$j��M�v�1���O��d�O �$�<�2�iO"`�@�'���'��ݱk޵P�r[��n���b��{}�'d�O�H���&�������V^�1[�����%f�N�@pb��L�S�O���ޟ�)�Dߒ'1�p�g�^�]M@��_֟��	ޟ��Iȟ\E���'��Q)��t����f����>A�w�'��7m�t֊���O�mo�b�Ӽ{��(+\��CUŁ&s.���D��<���?q��=! u��4���g2(q��b�^�#�I�P���af�\�B�5�Ĥ<�'�?���?����?yV���9" ����2/�P��	U'�����Yá��H�	ޟl'?M�	u�\�ЇS�E!��F�/ ���O(�$�O"�O1��@ #�� pY��P̄'�(��T{o.7-1?� gGU\��Iu��ky�F(L����%��alЁ� �8 Q���?���?i��|B,O�oZ�]��	
ZS��R�ݲ@�DU�V(��f^d�1�M{�"J�>���?a��)2,"���ln.!�]sK�T  �ܱ�M�O�-aQ��"��T�w�Dl�F�:x�ki�0u�����6��O�$�Or��O*�?���8 �𰦊S4G�`U�ܟL�I̟��42�ș�'�?��i��'J���!�>;2��dD�&&Q	��|�'F�Ol�e
�ia�iݕ�1+{���m�� Z`l�Ap�V��ɓ/��'��I� ��џ��Io:��2(Љ	8tHS'95~�������'ތ6Mˠ6r��d�O���|��'s�~i "I� nPhR֍�K~�Ƥ>Q���?!O>�OS�ё��Y�J� x����0J��*&�9�k�i'��|*G��(%�(��I�|�\�KG�Բ)Q'%�ԟl��㟠��ݟb>M�'pd6�M6
�P����WOU40��bn�O��d�����?y�_���+:��%��]G� �	�O�,�Ҹ������̦��'ʸ�y���w�*O� n4:s�3q�$5�` �qq09�5O���?Q���?a��?������m@L���ǃ�J���F܆f�ld���'�Ҕ�t�'�:6=�R�	&/�.).-��,D�cr,���$�O���2��IH06�7�s���U�-Ҥ��W��-��
h��q'�@�b��`�I_y2�'���+�Vl1�|�6D��r�'<��'l�I��M���������O�]a�	��z �ᡲi�H�8����'�D��?a����qu�1��a^-���T
��_��A�'%���C��.g�����~"�'��p�)X��z���-�^
��'�b�'���'��>�	'&��M�CA.s>���A.�@�	��MC%�����Ҧ��?�;Y�bd��"٧v���Sv�\�&�z�Γ�?i��?�Cd��MK�O���U/�?�ڑm��GG" qD�SI���6)ܾ(7$�O���|Z���?)���?I�_�03q�L�S� �3�m��p)������I&�Qyy��'��O�R�C�N��k�ʁatH��B�ߟQ2��?����Ş@t���%�H�l��-۵��+��,�>hR���,Oh�ⰄE��?9;�D�<�)؜L�H��pȔ�3���Q�E3�?����?��?ͧ��$Cͦ�s����s�D��T��P��nMa�H�����ٴ��'�r��?��Ӽk�MMZ~"51@Ύ~�bh���&9:�޴��ē�W�2uk��M�Ғ����Y�����O�s�a� [$���O��$�O��$�O��$%���":(&�X�H�+�v��8g�'��'�r7��W���Ob\na�>� D�6�Kk�l��D,qX�Q$���	ğ�Ӑc��<m�Y~Zw� �����7<�l�ue�('2n5�q�Q�^]b#�d�	Dy2�'���'3���:�:Q���H�nΰa5G�C�'=�I�M�u���?���?�+�&�IvKAmaY#�8u�5b���)�O��d�O�O�Ӷ ��P�ag��^䰹1��ˈ{�eRK�~P��!?ͧ������a� ���,̷�4���Z�$,��?���?)��|�7���?+O�!�S^��Ĉ�mF��@�}ƪ8���O�d�O"���<ͧ���O>����
(����!Rvb���O,��� D �6Mp�|��;�" ��' R��hnn@�"֯	�� �OP�T�I��?����?A#�F;�?a���?���?��->0��Fmǆ�n8K��8*�����$5�h��Y<�?��Q�������Q5F��D�&pΙQ�Z�r�뤂9e����OD�_1Հ�4�����O�	��Lh�l�I0thGH#7�����+K̺�Ɂv�� z�'1��&�����'�(��v�܍omT��Akް'G0U��'>��'�rV�@޴jWj�����?���W�b���q�\����F\
�;���>���?�K>A�K��D�$]�C�U����M~B�;B��PQk!�O��@��#r��%Q�$��� �:98�uXs!B@~��'$��'2��S֟h	�
��.!��LJ;�H���՟,@�4 �Lq���?�q�i	�O�n�7��P��F/P�h�d�dq��O.���O(��"�x�t�/L�׃��Ȩ�af_?"��d��nETa�N������4���D�O���O��d��Z���#�������"vhUh�C�<qf�i����'�B�'���y�#r���8VnR�s��t(��ꓢ?i������Ap��Ш��&��`kf/�3i�����e��ɽh��1r��'��1&�<�'S�蘕N�D�F B� �T@c��'���'����Z���ߴ#Ԏ4��>W��̇'c��lKr���M��ϛ��Jr}��'�b�'���P��P4�L���� `�x iF&8���d����<,*��i��9�onĉA�(��P�\HI�>O�$�O���O��$�O��?�Kp&��6����q珑{TV�'$���,�����޴���/O��l_�I:*����*0��g�0$���'��	���� vQ�oi~Zw�����د\{��rA�e�`��d���~]�M��Nyr�'1��'(�#P���xw�̖T�6hQUY�p��'L��7�MK���?i��?	/��Ӧ�2�t{��ܝ2��x9�O\���Op�O�t�j��n��+��X��@7nAl���mK~�O������W��y�)��WѾ��`@T2?����?���?��S�'��R�9�'N]�kqH�-D��*�@k9��*O�8lP�����T ��R��B6	�}��my��Iݟ�I�?0�l�J~��$6��Y�Sc�)\�W���	p�Ol~�X6 WH�D�<���?!���?����?�/����@�
w�\!`1��h���ÏƦ)��������ҟ<'?����Mϻ4�DI�G�:X��0SI�:�,qK���?�M>�|�����Mc�'A(���C������U%{)� B�'�>�:��
J?K>�-O���O�y5G��(�D�@&O4�YbF�O��O����<�E�i`&���'���'�� s6�G頥��`ǩI��ͺ���s}2�'I�OF�k�nԞOM�����@�ˀ��g��`9Ѩ�p��@���z�q��ϔ�$�VEG/q�:PI�Ce�$8�+�����ߟ���ȟ�G���'u$�ck�e$h4`�f�=3a�����'��7+<-���O"lc�Ӽ��]��Ժ�cb_j��<A����D�bL,6-;?9&f����)]B�? d�H��W�Q ���r���c�0 e/���<����?����?)���?�"�_���M�bā�h�$�� ܫ��$�ڦ%�q�����I͟P%?����p�F �`B�"� g�^�W�T99�O����O~�O1��<�4[?Eâ�u@Z'>t�xZW��
�P7mBFy��Ӫr�f@�����$
J�a�HP�FrP�)��	Y��D�O����O��4�&�U����,U�,�	A����"9���8W%9S�"��L⟘ʯO���<�w�	t4����~
Ҝ���I�8@nu�ܴ���B�=)�C�'m9 ����� O�L R	�X�Ti�%�Z.-����O����O$�$�O���3�S�FlˑL��I��HYg�T��'��xӆ��1�?���4��D�T�[�ֈv�,A�e�P�Z��ThL>����?ͧrh���4��d�7}����	z�f���*V݆P˓JC/�?��I6�ģ<�'�?Y���?15I���(0��C�)�䣂�?�����$�Ħ�Xp�I̟0�IH�O,���2��	 ��/f|�+�O6�'����?�S�,E�c�9EN��W�F�h��L?U�R@��mX?P�8���������p�|�+B����l�r���$��1���'���'���tZ���4�~��w,�]�"YS�O����D΍�?�������H��`���؟��P���YP*��AB�V���n�ȟ��I�R]m�h~rn��J�t��}���[(o�5{��-oЅ9����<�.O��D�O��Oj���O��'�0�*�S�u+��౉�(P�ޔ���i] (���':��'
�O8B�z���(U�
���	�.X���*�2?G����O��O1���(��a�.�%;x1ֆ@8L2$aU<I'���cY�9��'V�'�������'*
h
5�H�H`��P>�<*��'�2�'��Q�B۴A�Y����?��$����"mH�2<X�ԏL�wotT��(�>����?�L>���� ))f��ε�D�N�t~2N�k4�b�i1�zT3�'�r��LPM`�F�%1�X��G߁~Cr�'M�'[�sޡ٠f��=8�I�.4��x���Bٟ[ٴ~;8����?aбi��O���لi�0kG�l�����g���D�O����O�H�-}��Ӻ#����M<<��d��̻U��h�ǁ�J�O��?����?���?a��=�J<@����-8@��*G)�1b6nʓ0����J�'d�$�'UV�Ra�+X"$��i@=?ʡ*��>��?�K>�|zVJ	��D���aT��	���ܚ`.D�۴t�I5��,3!ܟ�$�4�i>�ȖJ;*fP�bk=~�fI�WLğ��Iӟ�P��ٟ�3a��uyz��bk��q{���+<�`Ra�^>�9�c��2�C5�(�4�̩oZџl��蟸�	�J���
QcB�����ı� ,dͦ-��?I�  R��i����d��f����\�^�"�2Y�I)�7S����O���O����Oj�d)���wv9kEaW;{�<����7*�0d����	�M���N�|j��D�V�|���O�dm��L���\���R�'������A�~����l���ӑ>�� [�.`����bROQH1��'2P�&� �����',2�'D�e�(�� m� ��M�*�dA:�'��U�4�ܴ<zX����?������H�,�k� w֠IjQ��&��	����O���'A��#�N.c0̽�e�?v�����W1�p�cܯ��4�F���s�,�Op��rț0�`��C�"/�����O����O����O1���A����G�C�ZI�S� A�c�
kL�0��'�B�`�b�@�O���Q�
��)�rc&z�$B0�ĬV"Z���O:�R�fd���Ӻp㝕�0��<��`�W�����	�bw�#+��<Q-O��D�O��$�O����Odʧ]+0�	E�Ⱥ>��܀��	�lZh`�%�	ޟ���o�s��������ˣ^��i�d蓹F��H���'�?����S�'=�t5��4�yR��&�n�B�2e|=r@�%�y�F%Q89�I!��'>�i>��	#��y��DY�yp3�߮mn
a������Ο��'��6�l�|�D�O*�d\�q ����-�xak�ds{��ܲ�O����O|�O>D �@O���Ί����FMi~¦D�!����:W�OU�=���:"��!$�p�N�/!؉�w��:���'���'�����\{CQ����%��RE����hٴW�<%�)Of�m�f�Ӽk��
�&T�5X�BUt�P��'��<i���?a�s��-��4��ĝ�)�����'.��	�H� u���1�OK�!j2����;�$�<ͧ�?��?����?�b�w���x#e�J)(MiV�#��ߦ@��U	u��t�������kkX���ǟ,�B,ލ��H&��1@%��0�MFyb�'�"�|�O�r�'��fһ(� D�e*��<j������8�&��O���A�?y�2�ĸ<iOG,�BX���d
Q���?9���?���?ͧ���\Φ�(�I�2Ѭ��o��i%��r��,�B�z����4��'Ͼ듡?Y��?��%�\qb#���U��݁1��-d���4��D�k����'R�H��&���t�z	z'�\�<����D��r���O��$�O����O��6���
���0E����]�*���Q���˟\�	 �M+�Lް�?a�!5���|b�_%?�(ȸG�/�Zp���L���'��'��@���8O|��ȿQ~� 0E�W��Sʘ u����p'Ҕ�?�1�%�D�<i��?9���?�w *<S�͉4�Z h7B�{���?�Ԧ��'Uh6��_�l��O����|��U;"�$[pE�v��-A"�I~�&�>A��?aJ>�O���%�yZ�i���3#x|�uJ=^(���%����4�B\��?]��O`��k�?C����7'Q�c�QÅ �O��D�OT���O1�*�E��6�=A�0��0C��9*B��R&E�H�l��'12�t��⟜�O6��Z51?V��cAʇgq� ���|k��$�O�m�2~���Ӻ[a�H����<1d �IW*�`�0_�+�����ey��'E��'�"�'�T>AWɖx�̸���u��CM�MSGCԃ�?	���?yJ~Γq}��w��5� A��3�%�ő�'̸, c�'p�|��t��/I�;O�qj�I�|�≪��V�FHf��7O�DH�n�(�?9�D&���<�'�?�+)7�>lZ��6���ͅ��?i��?�������q�G�M�D���A���uD�x�	�[��(SQ�1c����@��`�I U��Z���c�� !��٣f��3Ǌq%+Ƕ�\JN~���O\�x]TD��� �(��ކK2 �����?����?���h����I�-.��9��G�x�F}�'ʡ-t���Ӧ�C���L�	��Mӎ�wm�HمMB�4�F��"D�j�ٚ'�b�'"���꛶���1ke���J�P0 �/4�"��S�̓O��|���?����?���f�1�Q9��Ż&(�q\�hS*O��n��&���ҟ���^��	�����Z�r�n:f��,b�4��_����0'�b>�Q�7�X��E��-/�����$�o_~B�_�Nrj|��䓻�D��*�1�/Z� ]\33�Jd�.���O�$�O �4��ʓ9��ʕ;CX�M�����τt���ӫ��yB(jӬ㟀��O���O���P�9�ep2J�7�ƥ�  -(���x�m���� ���䟈�>���<�hx�"��]<]R�:2�{�|�	�������I����U�ǸFz�X��ۏF���'M=�?q��?�u�i@���O���g�n�Od�#�&���@�u���0&��O�4��� ��{����x�R V6#xlX���+��d�J��h��p�Gy2�'��'7r�E�)avXx�kC&�2�i���/���'���0�M#����$�O�˧��1��[M��MpsmQ�,z�)�'��드?i���S��Ɩf12���-}U�u���wnly`��A�tQ�9P�O���?!��*�D�S��  $EJ�dJ���;��d�O���O���I�<A��i�y��S5'�V�[B�[�/DJ�iC�4G;��'��7�)�	���$�O�����/���uC��%�b��O>��$�7�-?�ċĠ8v��>��Mŋ�
�IdFaD�Y�`�3�y�[��Iӟ\������	���O��
aЕK8�a
�.ր��@c�}��cI�O����O����ئ睶}��<j�K�xJEy��a������'�b>��5����y͓,e��8KH�c�dBŇ�&Le�}ϓb�$����O<i�L>�.O��O(iҶMUj@BqB�1��,�q��On���O,��<it�i��2!�')�'��9����(Qf�*A䙉n��l�q�|��'����?�����j+h����ߟ�@�� *ƤK�bx�'�	��l1��p����Bӟ�pP�'<~��h�2MB4!z��8h`Mu�'���'���'+�>��ɼ�l|�����o�6��K2��ɘ�M��a������Ŧ��?�;[��r�M^O�k#OL�5��P��?A���?!4�@��M�O�ȓ�6�
4kq�dYP�"�$e�g �<�O.��|���?a��?A��/�����u�A'S<g;�q�+Oxdmڐ��1�Iݟ��	C�s��c�ܟz���$q��@���A���$�Od��2���4� 9#�F��d�¹� ���zz\aA��3���y������'|�$��'O��������� eIB�� �'r��'���4S����4x;�@X��h;>�@vKۃA��Ś� 
5m�V����P������m}2�'Z�w�&� � ��⌶o�Z�*�#�S����k�@G����U���9cWH��a'L���#�/E���!.}�|����@��̟h����B���:��Aj��_�B?`Yڲ!K��?���?�5�i�4Q �Os���~�O ��4
��<�Ƚ��GU�-yV���1�D�O��4��Y�@�n�^�@`n����Le��Q�K��D��y��س^���j�	oy�O�"�'�(�(U��+t�͌]v��`�X���'�	��M���*�?���?(��8#���4q��ԏ3*A*`���ӨO��D�Ox�O��:�(��6hW|��	�bA"d�ܽ���R$>��ioK~�O��D����D�VP!C��7*��Hd	<8�����Y�V�R�3ִ�
�J��`$0w��_���03�'��fӆ�`��OZ��*��\Y��[i#��v��c���$�O.�+Á}���$W�[�Ǻ?��'��q��PY �a���b�r��'N��V���3�jOJ�	
��ɤ=��R���2�M��L2����O��?c���k���@|�����O���%ȁ�?����Şa��Mxߴ�y
� F}AJ^�XD�b ��~R�A"�?O��[Gd��?�'E6���<�-O�� *�,�J�o��v:a��'7��,4��˓�yr���/`0���պk:�DH�
Y���'�V��?��������[�-�{��а+CZbU�'����K��+"0�*P���
^���*��'��퀡[/aT1�n��)�a��'��9�Cm$~W�3Vm\�Y:]���'�6��KǠ��O�o�{�Ӽ�g���-%f��+_-�
��׬�<����?!�-L� �4���@�"!�1��O2*0�ŗ'���������"*��|�P�dE�������]%=_qI�G��d𦝚�Qy��'�I;FjZ�-� &@��N��aCu}2�'�R�|��
]>t�TAb�a޻U����M���sC�&nV剞*6����'��}$���'��T�S#4:�X@Vҥm�5�񉼤M�##�?I�FY�z�f�y��Kr%*e���?��ik�O���'�R�'�RK��8�� (U�J�)2�$�i����Ȅ�Rҟ������S5��Iq��P�$@����%,0�.�O�%*�k�-)@49��#<���X B�O���OV�n�3\F�'?@���|����X`�tC�w�&=
���~��'�����T�X�k��擟,�����D|�P��)��	�䴐�J�<}��B��O~�O^��?Q��?A��)9mhȎ%��	ȺPp���?a)Oj�l�P�4���ʟ(��B��,֌H�P\���Q2�3�瓱��dIL}��'/�'����XR��y���.��y�U�d^�%�X�%�.q���'�������K��|��B�;F��p�ZA%0 �(؆	�'���'���TV���ٴ]��$�� ���aۯ3���;�f �?�<���CD}r�'��T�`�ތ��u�#�Z�^�"P�U��z��Ǧ��''�8 �?��՜?Ѹ`�8d�,;��E�~��\0O�˓�?���?����?����i��7�b}���Ay�d2�Ķ>���lZ�/��4��֟���u�S֟�����1��==���Æ\1@..�S��<�?�����Ş	@`��4�y�ݠ�8W�2,��Y:f�O��y"!�sk"!������4�����E��AiE� �6}9�EQY����O���Od˓^*�f��w��'���'J,��C�&sCR�N�90E�O�'l��'K�'8�<���?����v�N٤O|8�-��x��6�(�Ӄ}��$�O�esv��:-�Ԃ���V�&�����Oh���O����O��}��t���҂���U�* $a^�1��͆*J 2�'�t7,�i�m�7�8�,i��N�r�NT1Gr�\���4���E�nv~¨��Z���,�t����lyJ�$�/>=�J>�*O�i�O��O��d�O��r��è>.l�7�N�dT(I�<iq�i-"xR��'�"�'�O�R�_�
�209��$@d��d�>����?����Şh}�|x!B�8�饬��)���j󋉧�Mr[�HQ��_H��?�$�<��Rb� 4�Y��N|��n�!�?���?A���?ͧ��D��ݱE�ǟ�1j�9h��xqa%�ms(Aٟ��޴���?Q]�P��֟���,;�*�k#$TYE"�+cX0��nɦ��'��a�"�O�J~���:���Ғ꟣P���@Y��ϓ�?i���?����?�����O�H08�`�M�pXƅ��69�$h��'r�'e�7-XD��O��l�Y�I6ҕ25�$Z����LPY�l'���I��S"T\�oZF~ZwX��i�m��#/�@���B�l#�2cꖙ'�R�OF�	Xy��'"�'BR�\�m�L�����Ye`�I��T�b�'>��*�M���6�?���?�,�.)�7G�&u_H���M�Y ��8O��$o}��'���|ʟ����
�� ܓ5�G9� ء��΁"~�H�2n�=\����|j�Od��I>��X�@�RAЫ�i�����l��?���?���?�|�/O�oZ	O��l��"�k��tI��S0N����ן��	��MN>	��(��Iǟ�M����ة�b�(�T�x�Ëɟ��ɞ%�Vl�^~R��06b(��'��$؆k<�\Z�fK�؀���oF+7��<	��?���?I��?	+��qi�	9>���`�ɑ�;���ܦ�µ��џ<�	��,'?�I��M�;we u!��z��*q��,Jp�q��?�O>�|�Bł��M��'�ZX����j�p#�%L�	�'�����N	��W-߭��� R�B�9��A1P��<~�ڍ
�h�4Ȫ|�������@�̊)��C-ɀ͔AKj§6� � �>=��q'O(S���:�(�*f>Z��ǤF��ڲ��<KX8��&�&H��T0&
�<�Z�Q�,��ÁY*n���y!�pM� V�W E�� ���<H6[��/+&tra�K�cir�PB�kDx�P��O<!
V��աXĸ�S֔���F�W�Q�ĉ�G��Z�/��t�ѕЬ�����(G�{�j��!�
j��	�2)Q���@k�)�"2.���c~Ӧ���O8%��D� �N}���f)���^6m�O�O8�D�O��������Ex��c
�Q����ʙ�x���'I"Z�<�Ab�����O<���VM�Ff�*\��,���'v�*��NW�I̟��	)g��IL�I]���lZPac�� ���#��Ц%�'?��%I�.���OX���ק5�@Ò^�Q���ȷMr~ �M���MS���?9��U�'�q�� �CB��I�����hԓ&�8���ix�l��z�>�$�O���,Y�'L�I.E
�C➹�l5�#`����Bش\v�����O��0J��`���!�~���b`��e��ߟ`�� ~u��ʬO�ʓ�?��'�����A�j8�\*��LmvT��}b,]�'�R�'Y�G�D=ԝI&ǐ31�( p�#.�7��Od�5��E}�R����W�i�J�`����a���i L����>�P�����?q���?A+O�)�3��\��BFm�������ݵZ��'���۟8&�d��۟�adAZ�]��D���_�N6�3�	Z&�&��	ڟ��	Dyr��&�n��"x�JН�B؀�nW(>�6͠<�����?��[X��h�'�N�u��k�z�c0`G$Z$�i;�O��d�O��d�<yt�������U(Q�pg�Y�V/��1�� ��M����?	�N��{R�UH25".ׂ)��� O��M����?Q(O�`W�Uj���'���OdT)�u ]��;��,�GY`�'�2�'��$S��?�P@Ɵ	S���T#<H�\�$i��ʓbp-�5�ih�'�R�O~�����"`�z�+���ə��
�M��?A3&�1��'�q��1�v!���ʅ�Rf�2�d+�i,��8w�u�����O����^��'+�I��t �J�;�D�CU��~��ش4˨�`���i�OH6)�l���$)�Q�#o�M���?��J8顴Q��'r�O�I8�+�K�5e�A��	*��'����|b�'�r�'fx5�f'߼K��	y)B��X��� g���ć�N�H$��ߟ�%��]�/3V���)&�Ȁ���X�ZOz���<����?�����d��a#���͆D��`�a\Pq#G���ē�?���������<q��T:�\������z�i2X����ʟ���`y҈�Y���S�q�$�)�C�!O����AC�Xo���?q���䓝�4�����QR�� C��v�E��E�-X�'���'	�Z�x)���ħf20�8�ѽ���!C%�2$��	z��ig|�T��ҟ���L��эE�+��AdO�~�z\��ig��'���1S�m�N|�����1�Y���ěU.������c���%��'���'��yZw��2��+|Y�9�%�Tr���4�����qV�i��'�?a�'�	�Q�}�&l��.1��& �6�<	���?)ї����4@��J9f:Ja�3mDЩmړi�:|�I̟��	����Gyʟ��!cF?[t|����R#J{�Be��V}��
�O>�gF��L��MR�b̊V���b!���Ms���?a� n�k(O�SZ�$�!�� ���4o� 
�N=	T�<Gx�n5�Sݟt�"��+��[�x��$M+�l���X�0N]oy��~��2�X
��U���*I�u8��h9�Ol���O��?��L�=-�	� �;!ܦ(�B�J;-�.��+O���O6�d��F?��"�bE����	_��X����yc�C7�ǟ��'�BNf)�)A�1��!K���7����,� %����'�����O\ʓZ[�m��$ !��:���C׶hN:��?I��?y*O�X���g��(����s�_���ç�Q̌���4�?YH>!/O�)�O��O��(��Fs���jS�նNg̕8�4�?�+O���ݲI}˧�?�������(����r���� 倾/��}'�l��Ay����O�.�W�:����#�B�ҷ-�(��Z���G�U�M�_?��	�?e��O����uJ�0G@�}��Ǵi �I��T�	7�ħ���eX!ᄻ|6�u�D��,����VNfӴ-؅��O��D�O��D���S�4��6�d���' 9&--����)��C�6�Fx��I�, B�0XGA�^1��1v�ǅ�eo͟ ��ӟ�ڡ��byʟ��'~À��Y���S';M�x�/h𱟸�䳟����A�Pg��CA;rή��Vcq�p��9~jʓ���k��_�TzE-�Hܺ�@D�Ro�{w�x��^7����O����OH˓;#|���CL;�<�cd�nT"�!`ٍ8#�'�B�'r�'��i�%�EZ
�)@�M�% �<�Z�N�����<1���?�����O�d
�ϧWVA���J6c R)r�N��}�LL�'T��'I�'U�i>)�	 �69AS��10R�ZS�H;t��O���O��D�<q�a�;7h��؟<A�M�V��˦i'/4�@TF���M�������O6�$�Ox�	=Ot��-�����DoD�y��ti�>���O��#3�	J3V?����8�S$0��y1H(u
����)E��	`�O@���OJ���1���OXʓ��d��p\@h(bDĕ
�x3��9�MK*O���dE�)�IПl���?M3�O��@�H�n+��,�h�ڴ���՛�'D��]��y��'��V�'ff�=h$ӊW��]E��;AfR�o��lt��A�4�?i��?���J+��Ayr�9oT��b(ߖl�|��A�X�7�M�_B�d;��-��Ο�Q�K��r�n|��U�Z�R�SG�'�Mk���?a�X��T"S\�|�'�r�O�)*��FL��$��V=f<�D�i�BR���#�i��?������ �P��, Z�>3�$Vr�\��i��(��b� ����O˓�?��b�48� �N��<�0��UG��%�'��'���ȟ��l�:��a���<5X����*�F��`���ġ<������OV�$�O<�KF�F�
Y��ˀ�F�Uf	! ��<����?�����۠MW@�'�p�(�E��:��Q!HiZMo�Ly��'	�̟L��柠�%�f��X�.S3d�e� �<>�������6��$�O����O��tbf���W?I�	3ˊ���Ȋ�m��(3m�.N� ݴ�?	-O2�$�O��D����Of�
�0�̜0�l�#�F�ydߎf�n!nZџ���Hybj�e�H�'�?����s�6팝�B�I=\�q"b�!%��Iԟ���ӟL�	k�L�IMy�ԟ��m��; �²OőQ�X�#��i剎�e��%��(���?]��O��Ǩ?.+�O�\w�4����6B�Hm�ߟ��I� ��I��9O��>��*M"7d���Z�^�ˢ��f뛶��7��7��O����O��)Jt}�U�HJ�-@�.�f�sEN Do8]�u��1�M�����<������8������"kD0.�e�9S2����#�Mk���?9��A�y��[�d�'DR�O��ZE)C;��M��*̒V��(���i��I���a�j���?����?QE)��:��q7�8,Z5Y�ċ;SěF�'���H��>q-O��d�<y���s+����QBk��(�TS�V}".*�y"T�`�	�����Py�`�������LQ�4�(��!���a����D�>�.O��D�<����?���z���l�f�h�cs�	�KU��N�<!��?���?I����d��B�&��'n>�A���7�M��d܈\leo�Ey��'��ş��	����bn�@`E� Iu�J��D;;&YB�Ç���D�O��$�O�ʓA�(PW?M�� Ie� ���S �މ)㧍=�"��ߴ�?�,O����O����y��d�|n��Z3v�dh��M$h_(3w�7��Ob��<1�i�m�������?��e����m��?/��	�Mƥ��D�O����Oj�#�	eB#^���SFGAe���g+�O�˓�}@ �i���'�2�O�f�Ӻ{чUEg�xj�j�1a
rp
���Ϧ���ٟ$�fa�,'� �}��	�
�d@
+�|YC)�%�C��M;���?����X��' H�H
(�j9(q��ެx�W/pӂH��7O����<����'�D([�AO�2|����_-z̘RS�{�b���Or�e��Kw}�W�$��S?��/ ���D<>5�8CpO��I��@yC�yʟ2���O���9>��;T�r�	aW�(Qr�Ql����@�U���D�<����d�Okl�.<c� O�m3hS�B�.1�6�'��!˙'c�''��'�"V�ذ�/�(X��N���J�ht�3$��YʩO�ʓ�?),O����OX�d�"�r%�e�b7
b#FL(Tx��#9O2ʓ�?I���?�(O�hkQ��|�Bˆ�x�8���5��I��M�)O�D�<����?a��V��`��[cI>DMD���X��tl�������Iџ��Iş��'T�H�B�~���T�t�'��v#L�y2�x��с��i��_���Iğx�IU^
b� �!^[�A G�"�tIT�j�Z�d�O��z-�p�'T?���ȟ��� 9�%�q�4!�VE+��Ҥt��`�O���O$���2���ty�ҟ�5�L�w�,|���gql`h��i��	.3tt��۴W:����@������
�*7b}��*,Ue�<�GQ1�F�'�f^0�r�|���ۋUW��F�
�q�+	*Z�f��!8`�6m�O���O��	Y�I퟼�"�
=?< �k�ᐶF�TC��<�M�@*D�?�N>�/��˓�?�G�n�̅K�C��ns��Z��¸ �F�'���'�fU�>��OD���p�ƃ��lV�C�3v/�!Fo�z�O���$��O��D�OkLO+  2��S��*R| 1 ��t�F�'Pz���**�$�Ob��7�������U+U�]i'dB�WЀ�� U��X�G����'&��'��Z�����l<� EK�V4�┪19���}��'��'���'�.4��G.n�3�a�[
I�R%�>�bP�x��ݟ���Ay2��$,���ӋL&L��4삘N���:5N�+�O4�D>�D�O6�L�$�	b��1NJ6Ww��)3��e�B0�'W��'oR�h��N!�ħz��%��:y�ĉ��(�~�h4���i�2�|B�'��b��y���>9�J&*u�0	��9$�U�%A֦��	ޟ��'?8���K3�I�O���H&s�*�!�FΕ8����F�$<N�i%�(��ʟ�§y��%��'G�ޕ{Ԍe��E�F!�z�o�{y2�B�4}�6�]}���'��T�,?Y�g�;l}�ik��Ɇwj� �P���	�I��H����ڟ'�4�}��,�1<a�m��� /���4e�����M���?9���ⷙx"�'^�!xghܚ��ҍ�D�%�R�|�0��^���|r�i�Ob7�^�{-�p+f�#`��S%h�	�Ms���?Q��]����V�x��'���O��U�]�d\��2 �:(��f���;[�1O��$�O2�DW)	���!=S��v�&P0�o�ן`��@
<��'��|Zc��h���O*7����M8jT�®Oz����O�˓�?q���'9�ΘHphۿ<�1J���"Д  ��x��O��<���O��$4&+��{��+��p�F�/K�(��'�O�ʓ�?���?	*O�8W���|� .H����Px�Ċ�� �6��@�x��'P�'"��'�,@b�O��BS�( �بR�2p�	"dX���	����Iay�bϔ�,���"4,<�]ん�	��r��Ŧ�E{�W�$��z�$р{��0q�'I�b`�p��
*�V�'��S���H��ħ�?�����L0vf�����	�*�X�*J���D�O4���=�v�QGd��@0���f��b7-�O��$��F�h���O����OR�ɤ<��r^�x:�f�.b�R]`f�H1���n�ݟ��'��ub���t(�n��0늲7D� m��M�K(�6�'���'����>�.�u�`�"i����I:s���E�ɦm��Y�'p�'�"`Qk�H���M]0��y��0[.26-�O��D�O~�8w��O��d�|���~�k��na��5�Mnm@� ���
xFx#<������'e��'w�Ձ�,R"ަȢ�Jٟ�
�Y�C`Ӛ��_�Jp�$�Ov�O���|�,�,MM2p����,�B}��]24�'��B�O��d�Ot�$�<)��K
�*��;s��W+W����Q���I����	ߟ��?��aș(�	5"�JlM#FK�:����|��'62�'�R�'�,�(uן(�r��V8J�Q�ȝ�i��Y��i���'2�|��'
�	�k�6-��d���$�͖v<%+QT�|����8�	]y��'d�%��^>��I0Jr -�%S�dC��:��>c֌p�4�?iN>����	pȉ'&,D;�n*GYrH���*��)p޴�?�������.9r�&>����?;%k[V�D9+�	�.} �{�� ����?��a|0�#A�+4̌����0��mZfy2��F�7-�_�d�';��;?y�j�)ZӺ}��.�	�A;S�ڦ��	����#�>���OÞ=gmJ�xbШۏ_��Tz�45�:)Zu�i���'�"�OS(O(�dƸO�� �2��$MtM:󄉫6�F5n�7$��#<����'7 ��fJ�=S�5Y ��	<F| ��m�����O����w�������O���g��p���C�2�10oZ"E���$�[����	�@;-��|i�tAѸ�4�X��M�i��,ZaR��:�����O��'h��%K��R9�@�GD,H0Z|PJ<�N>����?�Ħ���ǟ�Ҁ�� ��ݑw ̪���'I/�I�'<��'"�|��'	��΍X�"�hP�  Z�u#�#G�w~��䋻��"�(�?���<9#&ʟ:�*��V�_��y�"O�,����?Tx�[7� 7]���`��ԮBHJ �gP� <��0�� ����%�c.%����Q�<��(��_D���wg�.|a�q�eI�p���Z�I.8cT��e�칡D.��c<80�`�4H	��f��1<,�yf��~�,��g"l��Lc�#^�i}nhKgj�$UH�P��)u�H�cɩK��0�EE7U����G�������5Ș�2s�K*��'L�jD6#i0ٶ$�G�8n�|2(��� w��V���/
LPT!t�>����Z��AJ- ���P�S4��`8t��;.\�!PN��s��'[�\	��?9��i�OX�����`�4*�c̵z|���"O���k�3׎����-b��'��#=A�f�
b��]	�*ѳ!(X��FY��V�'�2�'(���(Z����'#��yg�G�M������V&��6E��?Ȳ���I5��d�6U:
0�r�|��F�{���g�$���3��71���Iܤz����'Ih`p��L>���
Z���h]6B�F���E�?1�O��8���t�,tg(@"�G�0 ~�����M1NC�	1
n�Q���c80���10 �vő��Sßx�'�-�`B45#�M	�C� 0>~�R���=��P3�'��'��`r݉��ß�ͧF���s�O]�!��D�Vm-L�DJH�0��9+�k�\��x�	ϓ�|��'�U �hZ�E�qs���bH0f�ta���"Z�"ϓe��"��=�ڐ�	�Q��p�a�D���	T�'V�O �����5=4`H.�/�d�@"O�qX��!����B�U�N����������yy��S.T)��'�?)d8��YpFGH)2��y���A��?�o�t�����?��O�2����Z���MW����!db	�J0����3K)�ݻ�9O��S
�	^��%8e)Kp?�0O�8<p$��@�떏Qj8��ؑ��O��<I���a�\���nPt1�j	�H�1O\���P�@9|�b񫎁z�-ȵ�"�!�$����!�]�O�Z$���T�cb:as������'�Yɧ�e����OB�'$�N���G�:!�&�Q4����A.�G������?�����/�Ir�Oԕs��i���ɱ|e���X��Mr-����}�$� ��[,�B��e���S�^���"R�A�xڊ����@8��'����Q����7ҧ�*r(�c��ً'��r&B��h��x�#Әl�|$���-c���l��0<)��,m8*	 �^nP­`b'6�,ͪ�O���d_>$�4�#�U4���ďPb�!�� ��Q$�>-����!hC�1)�"Ou��K������OI�Y�Ez�"O<�c�̷%��ɲ �Ψ\K$Z�"Ohx@��zC��Qd���B�"O M�r�0�zp����0[�Ʃ�#"Ona	/F�7,�{�`�Ff A ""O��� �Nv��W@���C"O��س�H���:o��B�d9ʢ"O�LP��ϵD��cD�����s"O���M���`g�4;:�u[�"Oz�����>Y>Ua���q���"O�l����:WFp�r�2�&�a�"O&c(PK"���T�#�,�2�"O4(;��JvɃE�܏l���a�"O����&u�,���&�*��幅"O�`j�I8.04�A �)��iS"O���r�	a���Q�H	�sv���"O�*B�ܺtA�5�P�À_!P"Ox� �-�Z�BFCȝ`�b�k0"O�݋���_#�P�UKߦS�����"O���@�����ũ������"O�<�P��K�@�TfY�s��A"O�L2��A�U��yಃH�C���"O,%�U�J��8�q�֠A�*$�'"On� 5&˿}�)�P$U�h���V"OD�e΃{�����ȫoW ��e"OdAY���1)S�V�&D�zd"O*����+u(d�Me1V���"O���VdV<c��̫�	�F��9�"O�!��;8ZRՉN�-�f@R�"O�e�� ^��B�.β��I�"O*�'O�B! Dr,Z�S�6x�b"O�pX���l����&k��H��k�"O��j��P=�zUؔF�Q����"O��q�W��5i���4�4{B"Of%����+��鰉�0k�ܵ��"O(**5E	x��UI�i���+"O�\�N^�U~�y�6(�'SBR���"O@���gԌ]��s��#&�"��C"Oܕ�A��n�(X�I"i�B���'f�e3�Kaʽ�C��>{>��\�o��� Kn@8s��&ZA��Ac!�wѾ�F}2��7�>�!���2S��Y� (2�ԧ3D��˃*�9;����MʞF��p&n������Vu�S�O�����Ѝwr ���M1����'3�-1B�V,+�z��F���@�O��P�k؞�#�m�U�,D���/;�6�+9�O�
��iӊ���O�=O��Ÿ��˯2	�(�"O�MC\e|~D�a�1�ܛ���K�'� M�C铫b2��G�N<Ll���\9n�rC�I�.�l� �Ȓw�T���C��:�>�LN��Gx��逭\aL4K�-�'(�M*�Fy�!�$Q�.��AI
�B���!�.Sp!�$҃;�\ͨ�ʐ!? �*3喰KB!��,d�� q��U��u2S�kX!�A�*� q�o�7r�T(u��n�!��@�c+�tA)J�bW�(8pO��!�$W�^0�4�@O<`qՎ$�!�D8QJ�[���(2��b��+p!�DO+.�� \�&���1`��g
!�߈uS����0Ts��W	�!���Qt~��i��lkWs�j���'�V�j¦J�$�⩑��A�c�v���'�"��	�$*o��R�D�H:����� H��~�4kE����"O��륨�\�P���Cݜ��*��'���KM�����آ�����"Ĵn����(D�j�T@qL4�PD	�m�t/:�	�	�dI�y�����)ͷ(	
l�j�j���V��4K�!�$�>{ϠH��t�bf�6jr��s�v�r�r�G��N|��ѵl�j��}u\.A�ұ�t  D��r�ϴTc0!1CY;lH��b�,�.-��MI�n��)��m	����b`z��%EG������
��@�Mm?q0�L3\���O�q�4#RC.�]2f+77�p��'�*82a�'��y���+8�L	1n[(ǜ�ʘ'T�y��Oza{b�G��O�j`yf\?I��Z}ۀy1 J^�3�*�`��?D�X��g%�M7!�*	������(q:R��5��+%���LB8yK����HJ(�x�HI�&ިj3>�C�%��:��}��'�� ��X�+����FP�u��n�	hΤ�1 �p�F�@�BA�mg&̒��-�I�io6"=� -��@���ۥ�Y�Ժ�"MU̓]T��&��a�@Y;r��� ���'�l��V;xU���G�-t�~5�ȓ<�H�Y�$��θhT�Hc���ܭU��{7㔻&�5ϓ��O��5�w�p�Q��A�6��p�дq���c�'Mb�Jb"�?4,|[��T�Ė�B۴|	�������븐�֍��:��ʓ�<ړv�b���	�+�̅��ԬY��I��!�+3g��Z��#"�/��웠�R;��
��C)b�!��ߞI�.����B�j�@V$N�g��9q6��=�qO�9��ܮ$�NQ��B�:=H�ę�Yo��"�>�8��=��!��C�,��B�I�"SpmqRꖻpf]!��B0U��(4	�&Ge��k�%R,Qٴ�(����;Q�p遆f@/j��0⣆�����}���ZԊ@��4�l�?r
���'��g@�+  �1�%�,x'��XІ8ғ_L<[$�� )ʦ� 7�-	�DI��4��)�6�47t��#�#oC��9eV�wt�����_����m��s�f�x3H׬�p>i����$�B,��
XY���ly��c�4Q*dm.+3�jv Q�И���Ô$z�q���/�1H��E��y�H	�h�	��"o��I[�lM�\��@�0���<�O^.ؑ��ɺN9�n�1���A��(aZHu s��J&aR�Ըu�LFB���hz��9Zr��BP�<1��I,fh�ۂQ�S������D�'e��16�ؽq�����f�(%� �����0#w��HFjF����z�LZ�<���g��9ER�)�)�,�`�� F0���W,U�B�|���� ��6F�8Cr�s����d�1,�� .�t��dj	�X���	� c�(�B�#��K�r �f�:Gn!��H�z!7D��~Ԧ�@D.�8-��0��02��Y�C�>%?M���L�1�`�]�d��WŜ=z�>=b��Z�B�I�$st�����
�Q�C�Ơ~��Z�X5��ɫ4` y�hX�o��e��T���\�'�ԭ�a$
?r�.a@^. Ҡ�
�c���1�!zpr �M�#j��b3�ح&ܒ�� �<���Pq$�v��h�%Y���>y�I���<z���r�蓰OU~�d{m>��#i�jo �IE��?�W�R;=���LLe��#�]��܋v�܈��C�* �[�+v�|H���M�>���>r1bS��OȄj`��p��ȅhd��QS�!��lcd@��E?B�����'2�PQ�) *R�	zCH�g�P=���NqF�be���wdxr� �<��o��D{"�'$C�\�n� X�K��0<�$(	�e�|rw�
`ނ�ǘ�U�� ��IJ�f!Pe.��-���Z!� Y�Ն�����`���ۖp��	���S'@|d�'aBP$	� ��P2HM<,��t��iC-@F�	&MI�.fp'�U=n�!�D���P}���V��i�Κ�|AdI���,Pj�'V�	�𙟰� ��
V>(5��9s3rx�E�6D��s"�1H��u�c1g�X��T�Tg�Z���J�&q"�' �ˀdE$uf�hT���v�	ӓz3P5��ӥ%�����M�,���`B�N�v��J�����Н��<�&��&KB�0�������	�<���Q���bR*2$�|"�$�9��]�ա�2z��hH��f�<Y����*�e)�^(���V�B��QJD�4L���O��,���	 y,��y"͞25��s1%	,Mh�B�	+ �>upCr՘�!� Ieވ "3�C'g�8�#S��>"��uS�8,O�\��N!+�:�j���h�hz&�'�i脢*dj��P�������LtA�%d]B.L�@�!��$�nhz�
O� �@x�k�=A4�M��&�9�F����>���]{�:�(#�1Ho|L�#�VѦ�>٫ӎ�"�F����F�8��f) D�D@���&2@Z �?���D$$L^m��(�E� �m��?�>�������f���;b�xèE�w��)�	m�(��q�q����a�d����] t�`����~"�ǽm�I�� �?aa	Ր�(O�5đ)2����c$�+-��6�'&��I����`.���cʸC�DbhK
��-�uDL� 5������/a�7M��E1���������a�)]���S�I�6nO�y)�س�l����	��l��'�>���8����E��q[Dm:B9��j�̼Yc+U�Y\^�ŉ���r�"�ݹq>B������|*�۟���u"W j�ܜAb֬����˃P��(c��w��ز��$$� ��Ӷa�>b R1
DF� 戩*O��
A 91$�'��'r�l����b�p��g\+Mڒ�XS��R���c�!=�I+Osꑒ��>IBj]	6JX�ׇ��4�����ϭ^!���+�-lmnJdm_�k����J�^:B݀V旣�0=���Z�l�҄ˎ�`�R�y��H=���)O�H��$f�佰ROU?4��S��S6���T�N%"�D)���P9>C�	�*Ġ �b�$@�>y3��n�:P)$J(t�6i ��C�wc��֧���?qAЉZj���B�J�*��9�J��R,$���'���R �����@�1s�,b�B�@�뎜%����wp0��:��-�\w�0�8g�Ddb�xz@W-I���2C�$���Ï2�IMKġ��2�S�d��Ǉ��w�t�ؔW5G��X��8!rn����IpTq ����S��'LO��9Q���_�i��<^�a�ܝ�Xb��A�ͿSUH��ɸ6p@��g�u���W$jB�c���0��u��ჵq!��P��]3���:G�0�PsO�R���@�G�B>�q`S+uwԱ*A�-����	�?^�>��uML~M��
�e�9��`��I�e��Y�d�<�� �CI �3peIS��"5J;m�r�2��G� �0�#T��Os]��D	b��Q�EW0NΠY�4�T�/Y�O8�p�JQd��L$��M;I����k�RV�H��Κj%^%`���1�Z���׆d����i�b�C'��:.��ؔD�?� ��G�i:\G�E ����|�q���K�!��_�~��#�"�zK ɲ4��$P�^h��cHb�)ڧ!�:}sN�(>���C��[\����O� b��U�K~�CA�v��&���!��mB ��I0v�nk��)p�ver�H�Z/6��dC6Ynu�ȟ�z:�{��T�.�u�EMS�P���uÆ,)��4aj�q*$�۳5�x��0S�O6h�&ɋ�{��lyuD�6�@��"Oց�Ł��:���+��ΔA��u��"O��Hq�֛���B(�\��ؤ"O�]@@�@H����<Tw�L�T"O,`Q�"ȅD�pE���!6�rh�U"OV�[V����MV��Y�v"O�EEC8M!f�@)K��Ȳs"O�q2���:��55 Zm�H�"O�LJ�m�=}TT��3��xB"O�XIC��#W�ޝ�PnW
x�F� t"O� ���"abt�lS�'���ڷ"O�IPǃ��z�4��-V�1��ʗ"O�0�m
$'����t�V���(�"O݀�eێD���0k�����"Od�`.�?8��4�=dm�;"ON�ЮՁB(x�#L�)qE�c�"O&HxAI�d����(Ӎq�*�1�"O蔈�Wl"&`�H� U�.��G"O��j"�G���Y7��h���[7"O��R5oĩ*���MӉ*�ơp�"O�p��	�op^�P���
��ձ�"OR z��	�k�2�4�̸M���P3"O�"�[�1�f	l<N��4#�"O���/-r�)���B%pP� �"O�TfN :��.��tX�T�"Ot �G_�h�0P@5��X^ܨ�7"OFL*Umm0ii�I]�}(����"O���.ab��vb_�`"�[g"O� @ՠ��C<�6\r�gP�%B\)�"O�H��"l޽sa��jͣ "O"�Q��:��J�%��f� R-7D�8� L�,�Z�ʀ�Բ>�)@��2D�l�%c h@d�z�萁0g2D����-J��hوf��6B��PJ2D�|3��)����☛rn�t��0D�Hn�� ����̘�
�J,J#�$D���OR����ee��[]9W�$D��9�d�N@N���#[ ln�-c��$D��E�G1u�i;-��dL D���A!DP�*č[�Hq��aU D��@���+NX��U�Yum�h�s�8D�l��Ls+�qJ���&v�^`2U� D�p��8}a��QKR�z����?D�x��"�#�՘oΘ{�A�Ԯ<D�L['H�"WF��V&�9;N�y�1�0D�����Z�Z���PŊ�%6��A�C1D��х�������ʊN�R��N3D��5��C���z�쉾Z�B��'3D�����Û���C��@̐�.1D��#ŨW�s��t{E�GF��&�)D�H蓢B�\�h)���4΄q�-&D���VC�;'������h�vX�'�����K%�"ؙ��@�U���'�a����#�d����8N1�
�'֜!�ٓL�(�P�
9N��'^�J����T<`���9���'�@���p�.e�w��@g��@�'Eּr�@�g�R� 뜛29&qK�'!��R ş%\���xK	%P0Q�'��S�-=��*b�ק,�R�y
�'�ZpɆ��|�4:�HG�{5B��	�'b���V'��Ȝ�:��M}�s�'��Eq��|����i�{@�'�^�*�QS f�X��Q4q�Ƞ�
�'�����9
���zc��c<8|@	�'\Y'�H�e�&Q��&QE	�'�<�'	٘)��q�Aא4C�)��'�x5�@c��xF����L�$%.@�H
�'�<8#�ˈ-nc��r�l+=8�
�'�����Ί!Q��;cKOK>��	�'}5Jw�O(k��<Qr.Ԧ{�
�	��x"��� �ҡZ��8�̭�"B��yr�˙�`��!�^�<N8�Q7G�&�yҥcM:�jЅ� hmq��Q��y��	�T��A�/O��𩒢ڪ�yr#�,C��QVI��B�D���>�ybC�p�3�e)x�FB�,�y�N�5V �cb��I&�(&��y�R�/�t�`+�i�ݸ`(��y� ��*er�ɔ�_,��+=�y"��35���ò�G=[\S$ǚ7�y�C�|�b���N�$��h�*Ԟ�y� �s!�l9$F�g&yst�]&�y"CX�	��)�Ӈz��, kY��y"&i��t ��X�jw�(��(֜�y2i>ą�{�Tce`ԑ]6���'�hCn�#�����cޕT*J��	�'r:9Zr/
p����Z9�^��
�'��p*�ɚ��yi��V��y�'&���OL�jT��2�o�@$��'qX����M�T3b�ԝ�f��'����&O2F�a�遠j�
���� ��`a��Z$H�0N� 1���Q"O�}��!�f]v�q�MD8*��@"O4�1�V�oj����1a�p�c"O�����=0�� ic)�#�"O��x�O�3��@gj=
��c"Ov�CtgK&&l(����<O_X�"O\�a��?P�T��׌�ll4�bQ"O@L�0�ݥF2��d���SS�t""O�$���ހ�N30{F4	��̼�yR�"��݃G�1$�� �,H��HO��=�OR�p����.�¤i���l�����'_�\&K�uդ��3d���h�'��<�qE�y���"�K�`<H�'�����٨]�d�=03l�8	�'~ؙ'��/�|�C���-���!�'�&ȃ�,ޮaq(� ��.1�8��'�,x��$�0$��0���٩(d��'�B�:��J5/�����G��ys�'��|"6&�$ODB	3@A��h�r�'"pQ�c��O�D��b ��Bm:
�'9�u��HI���k��,:@q�'����O]�L��{�nT0J��Y	�'/���FD�-�A�)3>����![�����'{����E%2`��ȓ99`�q��]�4��,���!EG�}��+F�B�(�, ���q&�Hs� �ȓ1�jm"vd@=T�,* 
,Q�`���K�"�.ǬC�V�$�����"O0y9t�V�pI�yr'��!Z��R"O��w.I2U
�*���^���"O�@*���q��)E���H ��"O��@'&U���q�P�j�f���"O"�B�aM!d��D�i�l�F"O��q�g��Y��C��w� y��"O��YDMH�py���M�����"O�ۤD4��h�周u����"O��!'��9���!m�` 
�"O��Hkɽ �y�f�5uQKr"O����Bm�T� E�3w\	��"O� ��
X;�MȓD�b$���"Ox��#mO3y��p�E�BgG�8�"O�P�"	�4!�tl2��[3I�497"Obl��H_06��q��=͢���"OV�1OP	p��x�VD�4W�4`$"O4�1���4�� 	�;MU�1�d"Or��-͊�t��"2I����@"O"�S�gк�J�y w��XQF"O���GX�y��%��Z!n�I���`�O�^�06
 2H_��k�O1S��<�'��q	0��,vw~H�a�ހ�4��'c��M��-��0����	)x�1���'�!#�GP�z�]�Z�4���B�<� �A�U�Z-↥�3n��w Ju�<�Ε/=���p�$K�|�hUno�<��n��m�����!":҈����v�'Uў�'N> Yեݞ5d��ѴI�V�Є��c��=PJE�!�q��ɸy��5��G�L���Ɣ�I?�1�R%ò�(���[Cn�*�����U��
L/�rĄ�Ub��+q�O=S{؉���]��(�ȓ ~ W�:9)`��a�N�1=@��ȓ"?t�y�I�I908L�86@\�ȓ��yX���I�i� e۔"���j���8anF�,��ۣ̎����S�? THԧ��o4ȡP�$��B�"OB� ףY"cR��[����
��Z�"O�ѻ��
1�>D@&"ϞH�J��b"Oj%�A <Kb���_	vh�=�"O�Ir6�	�IX6���e�\]�"OlQ����<r��@�Зf����"O
�3B�X
E�f�S�2�v�"OZ��@��}g��r�T�+�60�%"O2�x1
Q�^(��р@����V"Oz�Ɗ�x��,J�'�QqU"O��Y�U�U �q�D��./lT�b"Ox��N��p�5c��$��B�"OH�*�@̦p=�ܛ C����(�"O^���͇\�����ǎ4#���!�"Oƙr�#�8�<���T�d����"O�`z���|��12U��7w�u�v"O��x!
��\��D:#SQ"O*liׯI
gFL���țk�&Xi�"O୲CF;1����"��.�
���"Oh��é��Y
t`)��1gtAPs"O�� �7��rV��j�W"Ob�8`��1���B ��kK����"OrT�]"+�� �T�i�~tiF"OrqPe�H�#�^X���w�а+�"O�g��0����+���� P"O6i2q@��5�9H@U�$���)'"O�!��*��,�g�H����b�"O��I�O��^�|����T-{��=B�"O�D�Ƨ�'z��-��6V�\k�"O4��A.
��-��%7b���"OQ1an �8�`
�+1J��"OH��AgĖk6���w�aN��q�"OD�#̄N�4;0j0L��Q&"O��D�%h4��r1h��1��"O��*�a��[q��3��	!+X;�"O�D�fO�jUh��U�, y�$"O줪 ň8����cZ�:�`)�R"O����C'`�h�#�%
����`"O,�1�N�5x�0�!��۾K����"Op�s'(^U�3�
ͬ4�
�;�"O�-�7(�"7u(�& N����"O�᱕��!H>Y
A��3W�U�"O��y�.<�n�LS�h�� yG"O����M8 ��Z2˒�8X��"O4 ��H4E5 Y�@��-C����"O��q&�-|=Za{v/",�x�"O�̱��.K�ŁQ�1 a��"OZ��EM��(� ,�B���W"O�H��fΝM*�"� -b��X2"O����"�%(����p��E"Ov����ۂ�3���\�#2"O �dD@.l���AFm�@`�f"O�`q��	[7~���@��6��Ы"O``J��I�va�Q�M;*�j�ä"O����ٯ^+��j�gB7/Č��"O�9#���
�^�)q�$DЀMs"O(� �!ϒI���r���z� -�"O�1�@�7 +�m�di���y3"O�}T�Mа��RHF�h8C�"O�x�5��)�����b���"OH��oE�w1�a�ǈ�z�Ԝ��"OL����T�i�N�b2��31|��QE"O��q�i�!�����݉#�0�@W"O�4 ���;@QH�G��j��p�"O� �m+uZ��M����oef��"Ol��!��<5Qb�␄�"j[Ÿ�"O Y@㈀I����DM�!P��"O�9Hr���c�'I�N8��a"O��f �H�ܵ+R` #(ȭ�F"O�4Y��s�2��#AI	"���f"O�Թ���=c���Y����"4,�"ON�[1�Z_zT�,�"2�q"�"O�-z0��A�}���:rP"O��6�٢���>�;�"O�� N[LLI�q�T	Ut��Q"O^5e�Nj�����M\�/*Le"c"O��A4m�+�~{�\ɀ"O�l�e�ڤF�8�yw�S&g�P�"O�H����	'��+��͈Q*���"O�m+ �L��r�Y�|�
t�s"O��$��4�"�	�/��=AVY��"O�!	���m-���
�H	L��"O"m�Wފ<:pq"Wi��EтW"O�rV�H��)�JTk��M8 "O^1��Y�v���L	�v��A"O��P��r�z��B:�b�Ru"OF\x�C��HZ*ܠ�)ѬF8D��"O6CI�y���*W(�,:i�p"OJ��	6<�p�a_;��A�"OZqku$�<#Pe��!� z7<Y�"O��Q�H�|��|1��Z�,��"O8A#��Dh�h��/�7\��$"Oj�2*��	ɺ�PƎߢS f��"ON�����T������Q�o���!"O*T3��a�1u/��$�Y�"O�Z�įUV��*D���0]�"O�M"u�5(�� 4��Uո�"O���3��#w��#�n��)�Xl�"O��'�QD�x@mI�8�,��s"O�ybF(�(�
`+ژOȨy��$%D��[�o\�d��ZF�W�[��E�Ќ8D�0@��' "ֈ��'�	Ŋ0� D����_�}�S�p*�
�?D�x;��PCE�M)�G# 3���;D��)4h�F��L;�$�%%���s,:D��!�K�A��i���Gh��p�4D��jB�W=Yds�ȩi��My�2D���E��P������qN�eC�/2D��� � "$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j���e�{�0ʅ/'D���#��`��`��Gx�q�1�#D�� �uѷgA:R�8%��lБ8��(@�"O��z���|N�!�e��24XR�"O��C�dǗd��F�Z�_b�a�"Ohp��L�PȰ� L�G�
�S$"OZ1�hE.?X����"���P�"O4��e-�8�0k�&(�N�KU"O�QIs��g��5��K�~�@��P"Oh�aЎ�{�|�˓�%,f�� "O\HJa�T���I��*A[��(B"O�9y�� /�l�|P��o���y2o��!u�;��ܨO 0�O��y�U�Fݖ���@��Ze�fS3�y2�G�{Z�eˌ.i�1�D��y�!��fp�h�3��2r�Z7���y�k!Oπ�
�E0V�\顶C��y�����i�/
#8����u�ǎ�y��;m��5K���z�����y�iR#|j���`��%z�� S�$�y���/q�0�+��,�ubҭT��y2�^��pk��"���5K^8�yb��;8px�4�O��43c׀�yB���"��G�8}�"�:"٠�y"M�"	1�1 �n��ph�G�2�yr H�H�xi���5��)����&�y�e�v
zD�� ���D���y�-2P�(јg�����A�6�y2�1N�Q+�(�v�T���'�y"��K��1��l��|�%���yr�G7��Y��H�]��C��,V��PJ3mHai��x5�N�d&�C�I&-��is�ѯ1��$����#��C��1p��ZDo\�S�X����֩3}�C�ɡ"��8aK^P�|��٢�zC�I"s�ԓ��U�ED�u����V_bC�I�8�|��`�Ǆ%z��,<`C�	�(���P�!K�T�jS�ˡ�PC�Ia���"â<j�x4g�7"x�C�Ɋ�`RD�^(`	�
թhٲC䉘*הȰ�-J3���h�'S�ke|C�ID��!��A�	c��p�,F7�@C�	�,�(l�,F���s�D�"C�6&��$L>/)fA�񇆬2�B�	�cƬ���.��3�Fd�"B䉝z���9�*�)*W���CD�%��C��+/ڼ@ҋP�q��;�FC�FnB��<#r�쉐�ز���Ia��}�TB�	'R�8pf�'~�A���g vC��/�����%.�#U�x�r�:D���bƜ"���[3��kS���7D�0AF�E8<��d"��<QڱzF-4D���'�R�M��;�`�Y�Ɓs�e.D�T���+s�R��P�65�i�f�&D�DٶA��5x��BckɷZ�d����"D��S%�yj,ݫ�
�4ْL"D� �)�}��-0�'���{� ?D���D��7�,XZeН:���3��2D�d;D���s���ƍ�8)��r��1D�<��),��{��N�Ovx"�0D�Tb�Nǰ|4�	����ewxx��/D�� �1-�QE�ަ^�(�3��;D�#熋S���;�-ЮyC� �i$D����Rvȹ�PmX�l��UF"T�D*3B�9n�2)#���;��1�&"O�)k����zG�j )�F�vkG"O� 6��Յ�,c���$գ3�=
�"O� rS�>?� ��7�2�\$��"OF����ܕ70��#�C!�%["O�����(
��9b��$VD|�a"O|�#s`@$F4TVB��r]�}�"O�<�� ��b6��cZ�D>F�P�"O��sHK	uz)q����[��0�"O�$�&mY-�>��Kͅb5�tH"O�ٓҦ�(ڂ��J�L�|%�s"O�,[AOߘXr�3	�
^���"Oj��d��;�X��Jey��"OF�z���7��8*����԰d�0"O�]9���g^�0�%_�#� �1"O��Q0"X�2%<Ј�M�=��D"O�z��NM	�܀'-JX�i�"Ol1���,�=��"4Oe��9�b���XF�PeB[�.�,�ȓ%��`6� .%c���?+��h��?9�T�K�c��`�f������ȓ �p�e؝3����`�7�%��L��Urg���Z9��*�6���k��cE��:p�������e*D��ɐ4]���tO<P=����-&D��thͬn�d�+]&+��sTG"ړ���*§ �����ԓ�=ے���_Ghh�ȓ�*��RB�;�n����;5L��Z-��Y�Ā����с��8��+I0ȹ`%}��$��86<�ȓv�\���?+����q�˄p����P�
��ƅA���!��S?!����M]0�%���Vg
8���K�y���ȓ5��9{�.ԏa��|Jc&�h���ȓȑX-@�%�d���C4{��ՇȓFPu�U+^�o��@h�-\R�!�ȓ�r`1�K��d�v�ѯڥQl��ȓ5=��@�F^�L��Pd�7h���K�� ��E�X͈��)�4o r܅�(�z�Y�4o���aB<;3xa�?��N"L�f���[\�tA�g�by�ȓF��a1!��V���[ E�T����u�f���NUij�At��$a�怇ȓO�TE���?W$�t�&C:�>�ȓ'��i׈J�R�b��x��T��۠��cʘm��$/X�,Y|��)O���d����m��
_�+�Ԁa`�ڼk)!�P�e+Bu�r-^�� �H0�>�!��M&b�bAڂ@�>X}��z�I�!/�!�D
�A1��s�eۇ�L���^-'�!��@�`�����j�;S���(����6R!�_�v͑ӅG����#xȆʓ)ciSf�^
�Ű��&lB�	D���h����vp��i��`0���0?ٗ�u��M��m�3�*�����o�<Y�Ȕ:U�&43CksJd���`�<قѤc����A>^�`I�r�<�%�H(���K�$ж���5#@m�< m5rZ6�PU�6��Dذ�q�<Y7�5o��[���K���aJo�<a��؈`ZPp�`0\��r���i�<qd�g�c�k�^}�h�o�[�<��W�sT�SB�\����	D!�Z�<��<��8���j$,=%d�Z�<��!P)DV+0�P|P�C���!��@%"p���%��	|.9eݶ!�� ���Ԋ.�<|��8gly*�"OPi��$T�[���O��~��_�����=p� �zC�N���s�f_8�"B�	AF\���Y<�(�%�-D��C�	�OO<	���՛F�F�rq�,�C�	!8e1!˓�D�I�˕�+n�B�I�.!�$bB�N�T�9w/�,e�|B�I��p5¦JY�Ax%���J:C:B��\X��#bL?t��	��=3Q�C��%H�zɒ�_$l�<xe#P	-վB�ɁUi�H@S���#V渠d,#[XB��<|�n�(��|G�hIs% 0FPB�>�΀��� ?�n��ïC`�C䉜C�����"���w�3nC�IG�	�F��R��T҅���K��B�I�E�R�V�}_DY2h4:�C��9?h�4�2�
(���H�nC��:e��i�J��&N�����R1�~B䉟,���QKF)I>�
��2�C�I	#u�kteV�K�Tu ��k�B��!G�5�r�Ĥ6�f��-��PA��� B��sd��%I.����C=_�!�N�s�&�.Y`��e�!T��O���dB1�ְr1Æ64ڴ ��V��!�d$Qbf�2��
s� �R"	˪%G!���7�j�/%(��0�&�o��q�'{�$ë�>E������Y�z�v`	�'��9X�c�*(@Iʤ��"ۮ���'�HH���J)(���S���|YxO>1�r�I>L�<	�Ǆ��zeX@%�iςB��V�D�pE���y�n���n�XB�	r-P��ب�V�U��C30B�I54�çX��2���W"�C��P9�ؒ	Ɂ7p��g�A&�C�	3v0�K����Z�8"c�Ӆ%��B��
|'fD���+~��7 ��+�B�38 ���ݺ�>��c&"��B�ɨ=��\�0��6 �2\���Ԟ
�B�I3iV�Q���8tt�
�ֺHB�I�GI6�3����"��;�DB�	�'�v��S�Ηq(�Ape�b86B�I�y�0�!�H�j��rL�wJ����h�x
䣞�M��=0�� w��败<�	X�'m�Ɉ)�����Y�Y��EI��C�	�^�&X0���^��X��aA��tC�	 ��QBg�t����b%�V��C�	<tvi�E�\�{��ؒ@e]
��C�I7�8��R�$fa���E���[�FC�&d��@u	�/uL)���8C��8����(��4�pB
�Q'C�IK��kvA��Gd�pR�����B�]u�M�� �7:-)���!�C�I>l����-�X�$\6q�C�I5E�R<9��%	�m:����c_�B�I1�8���/ƞ)-�!!�̋��B�|�|t���O��)H�	�Zl�B�ɖ<�n)�a��t�D���]��ʓ�hO>a�)��Bi�Hڄ����R�v���I�θ P�!W!��Ee�<K^���#�f4xV� +(j8�V�B�qֱ��/ ���_4]3H,cZH���t��ɑ���z�d�+d��>	�J=��h�J�[�˟�i;�*$K�fЅ�e����dվd�4�	g勗qc�E+��� "��7AP2|�.e��
�yB�z�U��G{��C�-[��I���:^�ΨU䁘q�!�Ē/��}Q��S�;��B�!O��!��ĉ!Fu�ҦO:_����dOX��!�䁀}��Ӡ/i��m�L��l�!�Z#ưH��U1T=2�3�j>?�!�dI8�`Iʡ��q'j���)DA�!���*.�Fƈ�9K&t ����u��'��O?�"f�!^��B��CK�*���E^U�<�v��PP�A�Rlހ�n��G�H�<�m�2R0��c��X�H.J��QF�A�<Y���F��Xr����}w�r����<QV�_7@`����%���i��}�<���߀G�Rа���af���z�<�R"X1kc���$�
s��9Q�+\�<G'#�^�;� Z�$ �����p�<��ObA�&S4}֬�j�<q����? �tCNƌy�@3�d����<	�W�&��d���Bz�h��[k�<���׵/D�=q�eJ�HƖ	x��D^�<e(�|��1�$�n�\��Y�<�v�X�H��Mi���	k����%�J�<��'��P����ՠ,wc\D[�a�<9��Td�����\���_�<��&
Q��a���M:�����[��8�I��،�c���xy��%��@����t��CQ^L	�u��0����ȓ_�9#L��:�@q�5ǂ��Z���<X�+@�F��PJ���ȓ#z�Y` ��s��ճCL8 �ȓN��-�ҩ�7�8 ź�G�z�<)q�X�6�*| `������)Ym�E���O����́*[Z9q��?�r�'�T��)J�=����>�0�'���HG2/���ρ5ogL����O0uy�jۖ$���hui��f�>�� �'���|\>c�擪lM�@�G^�|bOG%�6��k�P�Y��Ě@A�!"��j=�ȓb����,=Z֘����	->���ȓIz�1Z� D�Z4B�z�E�C.�u����=��苽UbH�V(�(h���ȓR� ���;+�8Hـ��gO�I�ȓ_�(�hU*�7�‐�E,!?�Gb�'w>	�f��!�EH4e��zhI�� !D� �7$�ř�EL�t�bI�* D�,y0�dD�U U��v�PQBe=4��!4oܩr�@A�g�g[Hx
��x��?!����ɢf�$9��[�n�'"Of(��UjX+��ւ$
�m{B"OԜif��E��tP�	!Q"O��7�	Vp�BbG�{�b`�"O�P+GFB(�vՃ�Il�~ ��"O��3B�T!S$}�#��l�֌�r"O>�ʧc�!��U1�
�F����"Oʉy'�:@�1� GՓr�l���"O�E0��V��r�eШ
�@qb�'w��xbOG�t:sB׳>P�����(D�x:C�2���C� ��%�,�E	%D���w����}�eӯi6J�P�=D�4S�E]s�pA 5j�>gB���E&D�����]�0�
��c�z�ڱRǥ<I��哾,P��#��	$�.��D\P~B�	�
�|�sB�^]40c#NJ�FodB�	I�,K���.9wLa �K� �C�)� ִ�QŔ�m�ĵ9A�ǡ!/�y("O�*�@�n6xKb'Q�}v|�u"O���J6O%`��.G��""O<�P@��
u� h�K���p��P�|��)Z�'GD�K�Γ��v��㬚7N��Ax�'�ґ��G4!���nY�K�J}��'nΑ��O�'ؔ����=�a�'��Y�B��ɖ�]>�3	�'�b�IĂ�l�,���2Z�E��'V��s�䍽_��Y�+Y�3�` ��'�z�*
��1j��~����'ebX�6��z߬�Bb	�~`�"Oʀ��7u����F��sϤ��P"OB��cE��jR�7�@q� "O�)�%k���F �Q��o΀�#�"O�����=
Vv��ǡT�Y��i"O��S�&L�r�B!BL���"O	�� ބ{�]�PAI�-%�!�"O6��4��F^��¡��(-��"O�iK��H>y�BJ�ϑ"$t�"O�X�잠jǆ�A�^�}{�"O4l�~a���8>ձ�oǎF!򄎍g�|:�˓I mRb 
3	;!�dD,12�Y�.E%&� X���U(5!�d%�m�K�6��5�7�̓	!�I�W�|�ݴA�R�Z��_�7R!�Q'Q�̡a��ZXP��u��/S:!��E�I,��R(�c~к��^�>�!��>\&I&�N�敱���j�!�D΄ea6y�I׾R��C��5�!�$O!L�9:0j�kM��`#[�y��y���%U~0Z���N�bp���2�B�I�A��`����SJ=QR >
3PB�I)xt�g�_X*� !�P�'�JB�ɜM��H��WUu��2�-H-/!�S�0���#����bQ-�t�!�d	�9�X����D��!�w�� fA!�d�>�Y��GH�d��IԌ	L,!�D�	x� �Ǒ)P�a����E��h�D�.r�<�w�];"�*l�pc2D��ZF�A�,:���"<�����2D���SB"���l�Ct���#�:D��(׀8g�B�p��V7F�V�
:D� q`⊩Q�zU����@%��6D�d�g�ņ1H�8�0
.249�cA"<O"<�C�֌C3~��֩�z��`#�GV�	o���O=lqaСՄ'a�@�@�]�"��	�'Ͱq*f�ʐ'b�si��]�� (�'jr ��萧~�"�C��]ݖu��'O������â�S�'�8�r�'O��z��)>��s�
�h�I�'dwm�����"�b�c�'�$)�GI_�}�� $`��bd��'�%��,���PS��8�8�'��q��+f�ЃglO=kL���O�Z �'¢�ZGG�0��4�@��uפ�r�'��bG������Lܑ`p�uc
�'����.��R�U���Z�\���'���;c�1=�8�k���YkRE
	�''ĭ�'��:p�p���1"���"O¹�� �����(�h��"O>a� (� usr11�08���1���8LO�܉�B�'q��׭O��j�"O��@D��w��Q����"�z�"O� "�S�I�mQ��	���RR�"O�����z���h��Ǚ&z��R"O�`k��ٿX��}�V-ϡʨ�0"O6l��#t�Q��m�8����"O�"��B�r���R18�����"O�-��	R6eZ�ʓ�ˆD.d�C"O��C,ܷ6,��c�ԴN>��#�"O�$k�M9Vtۦ*�\��"O��0Έ�r�;�� k��A�"O�9�tJ�g`�q�#�L����	}>��1��lt������>�Ќ��$9D�@[��ԆO!EŐ��A8?ɶF�j���ҝ!�:��չVL䁓�4D�\��Y$s����P�S'��q��%D�|ۢ���A���y��Ԍ(�r}{t�7D�� G(��2z�SӠ5'� �ӆ1D��`�b�,�FPq`D�m+DqS��0D��(�I�f���sl� %nF�3��"D���Ѧ�> 4ٺ��X3��%� �+��=�Ol(h��0��h��Q�	
��s7"O����^&�L��M�.�ة�w"O��ÃB�<I�IhUGȣB�*%��"O����!ȼ��,��.����"Of���"-yt����"Fj�_� ��ɂ`\}����}�Hy���D@��C�I�p���ؖ �B���f,�:H��C�	Z2���G+Kh�� R��A�Im�C�	#��b��=e����-�FC��&CR�"����6�@���	�d�NB�	Zh�0t��K�9�N�| RB�	�WKh4��̀��<|�%�ЁW:�B�I�b���aM �E����o����C�ɹU$~p��g�-;�}䚟"��C�ɋ5�a�b:"�5��Z�KO�C�	�H\���%U'P,HKZ�G)6B䉪AM�$�"n֥
��p��Y[�nB�	�J~�H�狚<�\z�B��fN&��'�I�@q�����M�@������z�C�	8<K4��&��(���^�W� C䉋<���%�{�B�1�NڍzOC�ɕGpL�
@�*C�\�JP�ׂ^�C�	�Js�u	t�D*
L�!3G��LݤC�	T�@�[������JʜS$�C�	J�H]sqk	�oz��v(G�Vr,C�G#.=����0 �R)��+�(c�&C�ɭr
̩�靂!e$��gC$�C�I.�`��0�82LO�Ae�B�ɛ(I:pDC?y;�M��LG.kw�B䉈w4v�Yա]�3MN�84��<��C�I�@���� �'J�6([ց�3
�xB�	3�Cԍ\'%����B�P�i�(��$+�ɜb�̸�g��F���P�͇sf���%�ɷ$2���ר_,���yKʉ�XB�Ih�0cw͑�y��u��ʮP;rC�I)5��� ̗�<H4Y����Y�HC�	�?��(�CKI�Vp�X��-aXtB�2��lV��n!� �g� �BB�I�MQ��x� Ěd�-ȡ���B�I;�t��r��*T�e@#��YBB�#Z#��� ��MMR0�VJWz7��ȓzB���A\6���IZ>��(�ȓF$��۱���h)e*������i��e d!�
mT�)��t$�y��{���y����K
��͛�Rժ��S�? lHˢD�,�� W&�}T"O�(�g��?**�ԁA��	�Z���"O�M�O��P.<a�$��@�P@��"O"��S�1t�hg.RU�q�"O&=1vHD3il���#�j��i��"O$(���E3�
0���/j�hH��"O��B#@�P�0�����b24j�"ObYqE "Z(t��T+&��("O�1p1�����TA�W(a�CW�HG{�򉄟e�~u+TmY�04���N7I!�E�D���E�P��2a.�}�!��>+��ٓ��E&p�T�A��^�N�!��(�6�0�@	ӘM:��֫(!�D�Ҙy�S��*ULT!��(N�!�E�r >�)n��d�D6�M(�!�D�<&����nɶL���b�"x��O����;��ʭB�� KaM��>�|D��}��K1�Ý<����gD�|�ȓ<2�`Cv�:��)F"�1r� t�ȓ��ihs��B#8��!%��e�p���d,B��3e�� "���)F����ȓ
}���$�A�HQ�U��LRS�>���zR���

�B�����Ćȓ|\� 0V˃�ĉ���'
z���	Y�? nY�+ҁ�:�y��E�I�ҕ�ȓlR(�Q"�2H�z$�"�ܝH��܄�qۺ�S B�2��5��N�:0��ȓYź�ce@��9� �G�D�wq ��ȓ.MkP��<"%��t�� F#���ȓ+��3�!�)<���B��K�����H~��K�5Ia�At�h)a�3�y��	���gG�e2"dȖO�����d2����
�lS4�b�H,Ò�C�"O����S8g��*�ቪsH�D��"O�T f�	}�^��5�G@�`"O$�i�C��t��d��9GA����"OJ�:U�D�>��z�,�H4�S	�'XD�`�E4;�҈Y�C�zQ�QQ	�'�$:&bБ~���s�H'm.��	�'��@�@V�P]9Uܨk�X��	�'Ȍ���Kâp��0�ԯ��Y:���'���S�D�_�: �� (�����'
��c�vr���Îٝ$(M��'c4h!F��]`bec���ND���'�,݂G�Y[~�M��F߾;�>H��'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\���)Ą@/����f[~b!��/8o\��w�x3�)��GE	#U�O���-�D!�3� 6�yG�A'cR�{��Z�cvYS�'��' ў�OW�I�$��=5��e��B�1����O~���
$���Y�`O�n!��F�IL>�S�͉�6YRP��5���3Q�+D���V�J'FpP�)P�s=�8��3D��0rC�W���S0���|@JgE2D�,�P��I�m�@���\��#�2D�pw��B���"�s�p²C�O�C�I0����dD�aZ���D��:;ɂC�ɚ*��bj�.��̲�X�s��?���ɆK#�P����:��u��A�	�!�C,UA�(�+��5Y�,R�@�"~m!��H�eծ���z+�;��!�DIT��陁#nyԐ ��8�ў4��S�'���
B@3���޻V��C�I8Ơ�$��>�fD T'�.f�xC䉚����1�ɭ{MX�����1}�<�=a�'p�`��ρ@�Z�x��	g���w�Z�C���J[��A��J�
�Ї�<��}���W�D�l�@�N@(<������6&pK� ����PB
��'��U�?����~Z�h�#&�V#1�*i�R�*�[�'aax�Ăx�j��B�NY������y�΀:����eͦ\�20Z���y�HUlp� ��]+S<nt�fnH��y��N�3x`�k]!}�����B��y2�ȫtM��"M�!0��S�2�y��*�"��4��Ƣl(�M��yb��.3�`�q��
^>d�mC+�y�
�HoVq�a�� ��IAU�՝�y��G.YiBQ�r'A'w�������y�j�&���8Ďִk��![W��2�y`�M9X�!�ߕd`�;we��yR�/dŋpm�Ms��Cq'	�yr�K^����c�(2��}Cv����?��'&�{u�0Z���ZBHݰ&�.Y)���'U�8E�E5*����ъJ0���@�'s����>�HH�T�
o ���'8���2�K�5�L�� RA^�k�'�bD`�� �ẶK��B<
���'�Z�x�G?�T�����2��!9�'=�hXg�³c~��6A�4U�\]J�'ޙZEo�6ir�� wg�z�2m��'v��[��2Q���qF#P1~�.}��'���1ׂ_�/	���l�y��b��;����� �S�803jϩ(z9��"O�樑,v��,ie(�9Ng��� "O��a@%��f����ć[d0i�"O>
nŨ	w�%�CH�-��U�V"O|��sEz*P�'�(��"OjI�6*J�o�${f�H�y��"O�=�b�@=�-+���-8�py�"OҰ*HȮ$t�C(F@���J�]� ����Ic�h'�[6~��d�a*�j��C䉝Q��I���G�&L�]���H�M��C䉬2 y�|i�i��Ѳ �C�I*2�ĥI��J.�Vb+�)e���?i���S�OHTj�.B�	*��`��A]�UR�'?f�g�,eD Q�E(1!(�'iĜ�҂F+���1W��.)�-�	�'76������sY�H7�
*�J�'d�9h�3�� &��1AIb�'^9�*�<��;��N$��9��'K�	V���1<,c�IXSZ�a+O�=E�� 46��E�E�L;=���kfV��G{��	�:$���aU�/�����)M�'�ў$�<i㫕/]b�`��I��Ȣ�C�<�W���\�*T��?Jǜ-q%(Ue�<Q&M��� +"��FϚQ�Q	�_�<�`��.	��U��5�b\���R�<-M��S&�¾oq�5;�ԜR��ʓ�?����S�O���AJ�)H��{�*�c��y�
�'����'�x��-zd
a��E��'�\R�],O-^P�#ϜiJ�#
�'Hdp!�hˉaJ6%#��G�.���'\r (F�ƨ.���P�D�����!�'!8pS�HA�Ex4�w��x����'6��A�NM�Xþ)�GҿoL���'_����-g��֦�� ���'Bx��u���2�"
��"�I[�O�H�[׭B1u�L`�%���[�"O�y�$���L�RT)S"���b�e"OR�rΘ;<��̐�o
(��p��"O�\*��K�>b ZNʈ>�\!�2"O�#�ꊕ��mA&�Ѧmˌ��"O^�z�21���4Y,m�D$Y&"OR=H#J��^��䡆�ʎ`I�̀v"O>l��Ǝ6N=��Ҷ�
�g��"O��	3���<�N�P�D;�����"Or4���׬`���b��7K�h�x�"O����ͬ$�J 1�d��UX��"O�p3���;=�(}���9_�=�"O�T���ʆ)l��{q�B+�g�!��u�*@�e��k,�xAm�>c!�Z�b�c�
4I\���e�Ǭ_v!�Ā�_��h�D�8�V9sD��<t!��^ oDlYT�j�.�z	�?7�!���-�h�ѥީ/��|!DH�S�!���O��mIb��6E��H�֍�E֡�$�	f���ԫT52��XAV"���d6�O:9huEiGT��WD�&R�|�OrdS0�[:cD����g��G6�`�H�<�ST���T�'.��a�й=�"!��hP^�`�gI�U���6��17H�ل�G8�m�U�@W�����e���j ��:XL�IE��D�1qbˋ+qތp�ȓq�,�q���l�Z��-�^��ȓ�"�{�Ù�a �8tJ(_�dȄȓ6Ϻ4h�kP��Srj��\Q�̄�f����(3;���F�
>�-��C.�"7�Z� F@%)Q&��a:b���4��b�:a�fͨ7F�z5R���<H�@�!2�T�i&-;����=�9�LC*^V(	֥F�5�����LP�5���zN��< �QA��=D��G'	��@@� ��E}9qƌ=D�����T�`�fL�:�9Y��=D�,�+�n�����4r���a'D��
��P�0Od��*y��a��%D��	��'�~5���H��	���6D�TkW�֖KѪeI�I��n��A�0$(�d8�S�'Gn���V*y� ���(@.P��i�ȓN�B@K2��'>�����Im����<�<%�E�q����"�[!�ȓ9���6d�p0BE Z�h֡�ȓnv�+��g�6��B�0�D�ȓhg�$�쒲~���D36�$x�ȓ$���"Ʋ9nZl���/-�����S�? �Eh�ˍ	�L�9%�nQ�$"OL9���V�+a�%cC�E�h�Ly�"O�x�B�9|��� �o��R刬�A"O��pA�����JD�9R��̣U"O�@)�ヂ*�v<pb�v��Dk%"O|���J��0G����M�2�leH�"O>�+FdS�U_(Ȉq��O�t9�e"OB�ɥ�݌)3r���\<3�d1�B"Odu����1is�d����P�����"O��֭��	;ڹ�ŁR,ib��'"Oh�˗͙�K���'�QdT�@�w"O*PT�dw�\��5TL5h�"O�ؘ�� �zNp|a��õG=,L�!"O����.��Cnm� �9pTv�y�X�LD{�򩃼J��!;NŨ%�����cHD�!�ְ%�\��  ))�"5�#��]�!�S ��ͻ���1v�$��ᆮ}�!�'� 	���J=`e&@HѠZ�!�+o. ��0d[�,�u)"J�!�	j�4�c�.A] ϒ'�!��5f��H8���d��+�HBv�'2ў�>`P"�1m �M ���r���d�,D�d�'�"3ΐ���-�2H`�8D���F
,e�	9�Ϻ��õa7D���r-żM*=h�*�-`��=��B4D��Y�#�y#���2�!��Q��4D��RG�G�P���b
�a$)��2D��������kb��ZА4S�0D��a@�V��6�c!��$=Lȼ*6'9D���
�>f���k3*J���&<D�HYtY�1>0��CC�8h{pn=D�t�0L��90�M���P�>�7�<D�81"�%�%hק�15�xPcFM;D����I�k��8�2AѴe2쪁F8D��Y�ט;�]�,9��&BmM!�d:S?���U�N�]��S Eǀ@!�D��/t����|>���.c4!� vp�(�K�P682CN<I�!�DZ�2.�)�O�o28��׍�!]|!���'�0���I�/��Yy!�gئ�R&B~i:u�I�
r!��ڬ�`t���/�R����O$`!�O�X�Ve��c�`���fh�gw!�D�P�t���+T��Qe�66d!�ď:p��) �޹2�D�wbÞM>!�$[+ ^���'�0���Ѧ"\8i#!�$?�n�WE�i���8bY�0!��LlG͉4aޓ?�]����/~�!��M�Y7�֏U�=�*���'w�!�D��E;�Y� MؼF��u�
c!��Z�Qώ	⥈V��D�B��#�!�r��K���]�m��n 0�!�D${�41���v��͇N�!�Y��1�DM�R�����:!�D\G�
�����g4��i��ă
!�Dշ!n��cr��w9�<��N�Y !�$�& @�B#I"' QY"U�!�$T��(��%M�Q����Q-:e�!򤟸p
���䒊<G�P�J�!�B�"�ڱA �d9ʵK�Ol!�d��2Q��A�Ň,9���`'�3AW!�D�4u(#-^4$D�E�ԀOYJ��� g�,dy�& IJ�� k�yR�ϐ':����J�r��J5�	�y
� ̝H�+�?j:ĝ�FAQ"B���ɰ"OH|�chU0V��W-���%�"O�t�v.Z�-�*Q��K4���`!"OZ�y��L�0֌��$�
�����"O�d�Һ'>�C� V�c���!"Ot
��P� �Be9�F�L��!"O�=�u\)
��B����(�"O�
ՈW;v(i��/=��H�"O�eR�7�H�GN 0��,�&"O�MA�Jx)6p2�˳_�A�"O�t�'fq�Z����P�4Д"O���%P�jU���%$ۋ&���"Ojh��Rh���i�bE�YFlH�"O��{��I/�uh� �2::�ԛ�"O���6L��qגLQ��4����1"O��k%��>~qd�РOQX́#"O�M0�	��r�mr� �/݄�¶"O�Qk&��	vըw �;B�Z���"O��'U
����WO��k��(W"O��z��	a����$ǿ�jY{�"Oġ;�����p&��v��8�"O8�
6Er�r�2BS�*:�Q�"O@)!E�8`� �	��ܑ3(����"Or`z�	�*��%P7�`(V��"O�Q�tW�9s2�(2�θT�phd"OD�q��K
:Ȱ�H�<q�.U�7"OT}@� �pn� {�&��)�֐��"OL�sRm1m��K#�̰c">誠"OD���N��|2ŏ�1�Ru�"O�<R����I0v�@��2-�'"Oj���$z����"Q=�6)�"O&�����/K5��V�3muh'"O$�EҊ	��4hF�O��rT"Oȭ�E�M'@�X��\�MH��"O�Y��ъ#d���!� i�����"O�5Fi�(:z�Af��iW*���"O�\9�F�:��t�O�4>thc"O�uK��Z�('�S9D�""O��!Hv�2P9�L٤:j���"O��⧨�);xpK�i���t"Oڅ�E���E�6� �»d���ð"O6��$�� ����QJ����"O�u2�@U*Ĝ�)@+��R#"O
�2a�ƀ|2�5?,x��"O�x8@a8Z�:�`a�]�?v��x�"Or����W�]!�L1d2Ax!"O`�RӃ¶#��suE�8o�����"O���EF0Y}*-2��Ֆu��1��"Oй!S��}Y�#�A�o}�	Z�"O�����\2xYs�+�>lh�-�$"Obi0�L�p�RP�����(ZlST"O:�2���"#�|EI� żY��a{3"O-�¬�h�`a1D�E�ԁ D"OD��MͰ9�4�S�ܺ%��b�"O���+բ&i�@d�7S�p"Of�;뎚&T��`'��]��v"Oh���X�gF����ʕg�*0��"O����Ѐќ����Q�7�<Z�"O��d��qg� Y�� �Wp�3"O�s�N��Y�l���Y�&ؐ�kv"O���c$գ0����@eGR�ެ�a"Ot<2��Ϧ	�4e�D��"O��(��=BuX��ȌS��ĚQ"O�@�r
�/<Fd5h�V��f�hS"O� `��aĚ��`�ڷ�'d�H��"O�A��qS�8Уe϶/QRa"Oh���.�<���`d�[���p��"O|P@	�*-�&���K��(��"O�՛�%�2��e���rtP"O,�C��؅V�P��Œ22�b�"O�Q��j��T.�i�!$Ac����"O�tR�G.w\��
#��i(0l2G"O�a���E<0z t��$O&G&�E��"O谪a�ΝL�D�10dԡd���"O@�rpG�L�CԿ"�qe"O�ՠtd�Sx$"�������g"O<�ڱ$�4J�r�3�%�8#��x��"O~݀�\6*� ��*���M*�"O\�p�
ZW ��(!���@/�Ã"O�Ea�c�S[h!�
�(�`�"O�!�R�3��I�W�K�-�4"O�|r���+����h[�	�=X "O�))�K�� Y!#.U.�`�"O@�'I�+U�x!���ʨU�T��"O�]�&d"_�Г엇1�2̈@"O-�2䋦GN��)ë��I"OX�R��F�z�d�	2� �0�x�"O�s�A^90Xl��J��g0�eA"O2	�fI�?^�zY�r��&z�c4"O^5�3Myc2@��ş@(�0��"O�@��6����<�t]�D"ONda���Μ$�$AEo&�b1"OD��o�7p��t��o�<b���"O8T���"o�ɢ�m��,��g"O 5���%'6�)CoK�?��P�"O`RaN���Z��^�T� x�"OBPku+�W������2oݾ,��"O��y(I���[��T'̺ݫ�"O�����(WR��p���v��X)�"O���ԥ\q�t`��H�r�v�r�"OJ=��%L=Z�@#�!�W�T���"O2���GIq����E�O�^�ṥ"O6��lѱQ�1�͟Yݲ�j�"Ov$��-��<��eB��f!V"O
hRƚw�`�q�[�yG
("O���ʁ�N_|��1�T4��U��"O�p3Ej՝fB���7�*��r"O�����)�� ����"O�T#qeۉr�2D󲢇.��#�"OB�J��� :�.Y � �=I��	�"O��� � �dW�|�S����t�yG"OR�QaNJ{.����N4��b�"O<x�#�
;�Hi��l$�
�"O �z��z .0���P�?��з"O$8h!�CE*�@ڷ ]�]!�G"Ojly��՚r�0�C�U�k�}Y�"OJ)Ip�U���ӡ��?u����'"O"��#�3Ad:CӦ�IO�,�a"Oh�+��]��2ȣү��-9���q"O���5��!�*8b��P�w2
��`�O~���K�S �X������&���!��P�\a���K�V�����A�!�+d(���AO�f�����~�!�d:,�6t�W(�3M��P�BO���!��з9Yt�� *m�L��/�**�!�$�1x�f�5��h�!w�3y�!�a;�)2�J���تV�C�t�!�Ę�Y�t�P�0{�2�bSBS 3g�|�x
� ̙s�O�B���Hw{�[c"O�4 ���F�R����9^�MC���N�O��mJ�=��S��Z,on��
�'r ����R+� ��c�(,M�9��'�qO��}��-x�c;|� ="��@+XK�|�ȓ~���AMS&�$�q����O$����f-b1�UW�e����2c�cWa~�]�|��F�+,�RŠ�o?02<dSbn;D��藃�*���{V�+4�X�[�O9D��@��/B}��+�>���+6D�H�D�K�DD����V-_7�c�j5D�@�C��'��D8��J>ʹt+��3D��ɕ/�?f�5:5(
�:;��ؑ�2D�����א>����V ��Mr<Z�
0D���B���� Ө|zH0(�/D��#` J(	���E��x9Ь� J+D�x`�mޞg&%���ªl� 0I+D���+�=SN�W��,�v��$D��3ҭ�M�-ď?f���xC�!�O�ʓ:x�=b���(6H�J�MS�R�hD��
�R!q`D@8\{(��TM��BN(��ȓ$���L�#l�BZrH_�<��ȓ"����� hd�m�1��YX(�ȓ}�&a[�K^�)���D.�qZ�ȅȓ:%`��.�#'�0�c���r�;�']4��w�^"���*G�*7V��p�O.��<Q�4|��e�PW�Y�Ir� �1����\��O2N6�H�F
"�ĸyQ%�)4]!��p,L8H���<P/R��N�78�!�B�U^�� ��>�-
����ў�ቯ8��0AU� �;�x�	��"kx��"�ɓ�H��I�v��Xu�4!��h�&�&$�(mS�'%џ {�؊A�G�	�+��2"5|O�b��`v�T�Wf�s�F$%�h�"/�O��ɩfbU�b��5&�6 �w�\)��B�I�O{$�0��D�mHI%��3=�̣=�U�8�ddH��b������٨	�`��IW}R��ӌ�IB�<F�~ �P�m+�w�H�Ity�ȯ>%>-Kɟ�ref�/������;8�@̓s"O@1B� oei��@��p���*���'�bn�M�'��9O�4��LLfh�Ja��?��AK�O�0S��Qo�f��ʶ�&���$_UD�Dy��I�����@��+��)TU�\����*�k�n��w��{��M`�ݩ7�z��e̖�H`�֩�R��M�'��`���iR�����O>�����~B�Ϊ(`N�b�>8k��#���8���/�O�	#�,�>��qLŲ.m|���]��G{��)��1��,	bE�e��5�#OX�n�!�D��mv)[�]�K� t�"$ʁ_��	����'4�x��0A	�tÂh��O�]�c��y�ڼiDb�k��ڈK���x�����M3�W�a~rl���
ds��D�B�N�sw����>�5�����ׁk#���
��"�Y8E"D��S��X��𬂯C��!
p�!������
ç^��z�N�$?���`A�0RӔ��� m ����CHڱ��*X e�	�HO?i�L��M{�|`Ƌ�9L|���#D^�<��!���l�i��EbKZ}"�'Ӭ����9}�Ȍk�eY
����	v��1X⩜�e��+���.H!��hʚ��f�_z$��ʅ�F�(�S�O� Tc���m�b�X���c����'����T���D��TmŶR���r�'�4t��o�rӦ��T,6I|������ (H���V�F�T��CW�i�jЦ��4��I [��(�6%G Q�X� B7f�B�	\��֯�I-Vp#$`:I��B�I�dpj8T��!XF���9ijB�I�-�
}�
��� H9��{�8B���-�
��7� ��0�����Ms2�!D�� "�2��=!��)!7>H�� O��=��-��n�@(ӗ�@�b�zQ�g��<y2+|Q��Ɍ�e�Qp 
=T��F���_���#9F"�/:D�D��K�A!�ʔp��c�M8D������/RуM��&�2�x�E"D�4���>O���3r���"]�-�ҡ~� 6�#�O��b�֙~�D��f*?���2�'Չ'���B�j=zO���W+��{�J�
�'�Ԭ+��[
n�YWmY&'~���d�M���cf�6% ���Y=N�!��S��� �rN�\�e��ўd��I';�$�Dj��Q)�hN1'�HC䉰�|��Ɠ[��sW!�)KFC�	%5<���j+��!��0�B��t�8 ��6@X	#�eɿ%�vB�	S� ��F˶ �hZ9R�ԅ! "O.�q��P�;=� �ѧT1���a"O�\�	����
����Ќ:��'剜	|�@y�!Ӱl��|��̳d�C�$?Ґ��0�T�XLh�"�	IT|7�=�S��M�ԃ��Q�bJPIɽb��*�T�<q�,\�O`���7:R`Q˒&�ş��'��|��G�@��ш�E܂.H�t!C���=!�y�
L {	b�a���'Z X�����y�Җ~t�8�� &="�BFB��'^qO��|:񏂚5D5c�+�k���8ሞz�<�t���#�9j����x�'ўb?��ьϲu�:�x�@F�����:4����*U�"q:���=f�tU�s�qy�)�'&cn��`��c��s3��S�T�?���O�~�������,Q�w��5���Te�D��:5BY�Q[�m֏)���!!2OZb��Γ~�� r��dި8I'N�Ն���O9����#�~!g�r������<ى��S�;��L�a눉{4� ٢�ז�dB�1qN�Y�������I�E�E�VB�I0����#���+:X%q�߻O�6��d8��9K�rQ��Â�$�BIF��Y\O����kx\Pѥ!���0`��1O�=�|�U)��CD�!3��<�|���c�<�ᎸJG��@�/�H^r�+��K^~�L/�S�'D� ���Bˤm��B�̍2*�N �ȓt�d$�pĚ�jnPp�ڢj�1���d#lO��G#�L����G`&���D"O(
 L�%p|zǬ�01��"O�ih/�'r�Ƒ0sfԄ��P˖�$�Şqa��Q1@͜h��Iy�@_����ȓ��dhP���hό<�MGx�'�J$cĜ1dL�	��Y��'?�d��2��a�1`f~d�'�"d�@""���(A��n��t`�'��X��V�Ed\qb� �'f7>(�'�%�c)�<O��8ه��U�����'Z&U	����t\.���&��Lp8��
�'����a[;$^�GB��8��B�	^a~����KP�k��ހsضC�
>$t�ŉ[Mp���� ��C�)� L�Rf+�5���0�,��"O�P�D#�nxh-��$#���+0"OjP0$�%j���w$��	�H1!"O��A#��{�)���W�9K�D"Opu���ľ��P▃\=�L"OP9�!����@�V шL\�x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  3  v  u  �)  5  j@  �K  �V  6b  nk  �q  zy  �  ��  N�  ��  Ԙ  �  �  ׫  A�  ��   �  `�  ��  H�  ��  ��  3�  ��  X�  ��  � �	  � Q  �& 1- t3 �7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6#\���<4�d5h��'�B�'���'	�'/�'�B�'���$��^] ��/U�Z�3��'m�'�r�'���'K��'r�'cظYA��4Z8�xg&�=�nܳ1�'�r�']�'���'l�'���'��41Cl֝wMƩ���0���4�'��'[��'D��'[b�'���'զ@�R��}�[�&���Ģ��'Z2�'�'���'x��'��'T��s�D
����c̚�	P�'V��'��'2�'��'���'X���EAO91�(��@�{�x=���'+R�'6"�'���'���'�R�'%l$�H^�C

��\�o��ص�'���'@��'���'��'��'��12����4��x�Rk��'n��'�2�'>��'r�'�2�'`P��6�.&M��;�	�:�d2R�'��'���'���'[��'���'��u��Ǎ
���z_��BT垲�?���?Q���?q��?����?���?��O�1^�����*J+Q4	zT#�?���?���?y��?a��?)��?i%��=�61Tg�y����ڟ�?)���?!��?Q��?��Px�V�',rl��~
I�"�m���rR"�U����?a/O1���,�Mh��#5lQ� A��*���;Մ�!ct<�'"67�4�i>�֟�`��K/.�i�����lm����ޟ��I<J �hn_~B:����[�	�7A��!�6r�.$0�m �9s1O,�D�<���)L@мp�G�'u�$%Ҷ�L�V>R�m�f��b������y7��2������A�J�\��������'z�>�|c�.�M#�'/r @����Yj>px1D�%Ɣ9*�'��CǟlQr�i>���=_%X�PPjlV�cC!H�_(��IJyҟ|f���8��d�
�NtRaÝ�	h����i��㟼`�O����OB�|�Ҩ�t">����('6�b�MKI~��'!�U�tCۖO!�Q���BVr�D4'W�0a6�U�s7�܋T�ž9�@yB������5t�Z,�i�]�\���'�o�L��m0�-6?�Q�ie�O�	�%؈ ��ʱFy䑖g�~M��O*��O�X��a�
���D���d�0v��'Le`���"A�~W��)!�A�����4��d�O����O�����q��P���K�4��J��F'^��˓k��H��6��'L��I
�RZݳ��[�D��A�.�J��'�"�'rɧ�O:\5�`�@�ebp
�g!Y���� BFY�
,X�O`]!�Ō�?	��"���<	Cճ]x���Ǘ�u�$AX�S*�?��?����?�'��S��M&ٟh�A*� ���f-�'n�x)������4��'�4��?���?i7큄�F�Rc��m��Q�]��!�ش��$N.d��I[�O"�O��E�����G��s1� #X��yB�'���'��'32���ln�YȢ	>�U�%`@������O����ۦ����>����MN>)�I� �n�w��2i�|l�e�����?���|��aB��M[�OdR!@J�5�ސ�QJܚ�ܢ�`X><��@r���ƓO���|���?��^���+#�ƚx־0���)%Opy��?-O�mڮJ�ٕ'p"T>-��39M25�q@�`6	�a�'?��S����j�S�ō)r0@ٲC�
b1�,��KQ�@�`�]�)D��$T��Sw`*�B� ?��8Jdv� �1a������	ݟT�Iɟ�)��]y��h��h���L�4�j�%�{��c��Sx���d�O��m�s�|�����brjR!&�PY ʇ���)k7�V��4�	�\o�V~	&TH��}�+�y�C��1nh�c$��<Y)O����Of��ON��O��'�4 �DЫe�B�P�]�IF��0�i|�r��'���'/�O�B�h��NO9#�B�S�`]�''ʔ��g@ ��$�OғO1��|��$z�@�I/�����:qs ��#ϟ�/���	|И�w�ON�O���?���Ŏ0LU������-��Q*������ߟ��IqyKtӼ�����O����ON	jV��/t�$Ӓ���<dp�4�I�����O���&��ƖlʜM3��2O�,���Y�n�I.f%���Y����K~
󩻟���^{�"���h�ֹ)v�č ��5���T��ޟ0��X�Os�$��@�-�0k��8�9PE�F�i@`x�Θ�g�On�D��!�?ͻ@)��n��t td)a-�&g�U��?I���?ѡ
N��M�O�n�&e���۠e�L�J�LJ2��8g-�"V�|�L>/O���OZ���O����O��w&�}ېhB �J��i�ã�< �iN`hHd�'��'B�`� Y�$!��!ƺ\w � �XP}"�'q"�|���'_z�)��7�����0�q㠷i�˓]?�����4'��'�LdcN�y,0�;F�"y��X�Z���	˟��i>��'dP7�_�:j��D�s	�ĺR���M�R��=U6����m�?[���	�|�	��4�6H0ؕ��ߵ"��8���y�'Պ����?��}j�{�? �¤�*~�zI!��{��E
`3O����O���Ov���O�?��d�/uBX���g�L��(�ʟ��I�`�ߴU�!�'�?	�i^�'q���Q*m�^UsS$�Q��Q⒗|R�'��Or�D�i��	ހ)9 K�(���A�KY�ƊF3��'���<ͧ�?Y���?A��=zؽ3���;m���S $Ѕ�?9����Dަ���fOџ����� �O����*�"bl�9s`�\�q�<X�O6|�'}�'�ɧ�)�A��(��T��Pq��
z�Q��`\e�E1Q���<(�¢�^�ɨw ��W��%0c��F�-Z�D�������ӟ��)��Ty��z�����#���0��8c�V=��^")>8�d�O��o�h��Q��	��'G�MP����DK�P���+������8=v�o�X~F2d($����K�^���dK�<�dīu�At�<���?I��?I���?�*��8�D�ɱ2��(:���EB�"����$#ޟd�	��%?i��5�M�;;!�}�C ۬��ؗ'ߐ�%���?yH>�|z5"̗�MK�'[H�ӦM�)/�i"��-���R<O޴�4凾�?�eB>�d�<����?��HM�y��z��`F0'Ӵ�?���?Y���$�������F� �Iޟ @��&D��RƵ<������A��#�����H��t�ɚ>�b�y��
�%�r����[9+߰�K��"4ß0gV���|�$c�O��Q���h�L+U�(p���_-d�y9��?����?���h�p�D��h}
�F�1t:e	�U���^�y0'�NƟ(�I�M��w��YwN�+�((т�^�(�|̢�''�U�D��F���'����2���?MG"ɷ�H��@Ur
={�fAtm�'q�	۟��I����̟p�I�3ژU��D�I�����ć[l��'2P7���&8�d�O��/�)�O�9�P�ׁV����ޅ |xH�%�S}��'vB�|���EW�g0�1�s�_U�D��ژ8����a�1��D�+q���f�̒O���^$i�C_�"�s���,�Z8����?I���?y��|�.OzLn�X����rj2����3�f�c�+�6���I��Mˋ".�>���?9�;>��pQ�K�MV��@jۣi�r�� %I�M��O���N���4��T�w�:��r��
"�A����n�6E(�'F�',R�'���'^�z%�`J�|����3S�0t9E��O�d�O�o8�*�S� ��4��L�H�cQnܖh(����	B���L>����?ͧz.�L��4���4�@*�	�?wV>)�g�Δh��ARdա�?!g�3��<�'�?y���? �T!A��y����K٥X�`���P�'�7�/r�(˓�?�,�� &�0j�P���ę�q�哟̰�O���OƓO���_��䣓��8i��H�q�ϞT��1��M KXI��)=?ͧ!���R���Q�{d-Ĺ@L�aʓ�+�t����?Q��?	�S�'��D�ڦ��d�B';���H��ƅv�*	�4�P��.d��ʟ�y�4��'���?� �9b?@y��ORt�{$g���D� *7M)?)��R��������d�\�T�I�B	��jI���L �ĥ<���?����?a���?	)��	�&JW��"�id�ٌD,M�� Φ�Q����(����X'?-�I��M�;j�@�S[�@�CV?r���0���?M>�|b��8�M+�'�`�p���)F�����@.s"��1�'��c�_��27�|�[���`@���6,j�5i����"�ΰ�7�ɟ0�Iܟ��DyBHl�b9�Aϰ<A�S�*�zp&	#�<5('�d�	����>y��?iI>��К(G��`-ǂ�,H�0��t~r�Z���QbΩ��O���I�92"�Nz-n����N�N3X���.�8r�'���'���͟�B�S�y����t��0�� �	�럀H�4� �;��?���i)�O�.N�[�8�Y"^5�5GB h��U�'R�'q"��E������h��I�S�D 	�*K�j�^t@ɐ�[�%���|2Y�4�I��8����	ǟLP$�
�HU�&ɞU�B�h�(Vy��|�F=j�O����O�����d�\� (���Χ!Iy��e�h�'�"�'�ɧ�O�0�]`�����z���ɀ�+�Z�"Wΐ���$�+
V��:�<r�O�˓;��Q1�D�4� ٻ3�Pk}�]��?a��?���|�+OԤlڌ����ɩocY�&.�LZ)�:nx��I��M���m�>���?q�{ǜe"P�,le�@��Fܪ_ج ��@�:�M��O|a� �1����T�w����t�I�4������IjZ��'�2�'���'��'�񟘰x���A����&n��<2��Of�$�O��nZ1v��S�Ȓܴ���rx�gǀ�L�4I0Č\y����H>1��?ͧUZFxr�4�����~�{�J���1`�uo�Q��ƿ�?�)��<ͧ�?���?ɷ�T�G�H����A91#W�����I���'�"6�]>J�j�D�O����|r�+� ~�np��Y�G��i�(Em~�I�>i�����)
�%�����쒒q@,A�u$�R�����^)1λ<ͧHB�d����Z����N8m��SA�'	�����?����?��S�'��$��uKd!�7*��;pn۽*�(EjfC@uQ�u���0��4��'��ꓚ?9T�ױ"������4oQj����X��?i�(��1:ߴ���I�^�p @����3� lXxǁ�c}�	#a�� Wg�h) ;O��?q��?���?a���*~N&��vi�i�� �+ZY�An�s�,}�I��p�	p�'SW��w���cÞ>)�b�]ή%H��'�"�|���JO�t���8O�:�ę�����B���B��y�N�LN��I�e�'N�	ٟ��	cb<����΅:,m��#/c��m�Iҟ ������'�7�=����O��D��i���gT�"�ny ��ił�H�O���Oj�O��3K��M2R
 +�)><P������`8����mf�Sa?mW���$��o�|p㳒�+�"X=[F��' ��'��ߟ�I7cP!qZ��Jԏ?y�4a�/۟<��4~�@u���?���i��O�,B��ihS���NZb�,V���O����O����xӾ�W����?1TČ�j�8a�4��P!蠫lPS��vy�O��'��'{��IX9R�	�AĨkԥ�*G#剽�M��#�?���?����K[y��ʱhJ\>�� ʖʰ듅?�����Ş�����4`�!��U2\�Q�@�l���Of�B� � �?1%*,�D�<Y���@z �: Ά��w�(�?����?	��?�'��$��)!�M�P0�@�0���;�A�Iv*YЋUş��4��'�꓆?����?	�I�1~n<�᷂��e�ٹd�O�GF�޴��Ē�$��e��'��O��H�>"N���p�A���P��y��'���'�B�'!2�I�@|���8.�p-@G ��U����O���^̦����q>�����M�O>a&m�f�|�j˩(.����[̓�?�*O�PQ�J~��f�z��6Ȋf�#�F�7�t�Z4K�n��d������OH���O$�D�K�mi�n��A1�|"KD?z���O��5Ǜvl@�v���'T�R>��2�ѩ4�,����B�4�TQj�"?QvU�P��ٟ�&��4�؜Sg�_
qI8��u�(r�Aӎ�9Gm>`ݴ��i>qb��O|�O.�h�l�Rrf�k�P�]���K�$�O ���OD�D�O1�|˓��hǍX�R�1d	N�uI�E1�O;g������'�R{���ѮOx�ĕ�s�x��Q �8���%��ʓ,��Aڴ���7iM��'1	�˓x^��I¨�Y�~�R#��Q����d�O���O�d�O�D�|: �J�5 ��	�ڝ�Ӄ��'��6�'bS"�'}R�)�Ϧ�*0�lE �G�Y���0*��oj���I䟤&�b>y��G�y�O-�8;� R7�pUK��2te�s
|u#Aj���%�����D�'/:uYW+F�&�p��^�<�@%�'���'��X�[ش�<���?q�.�z��3�],19 �����C�x�'�>���?�O>C'�!J�x[R,���>8`��]I~��XW��I�i�V�����'bbL��>D8�!!M�M���%�9���'%��'E��S�`�5��!�����eՓ~@�r�M՟��۴M�Z��?y��i��O��p�쭃��J!sN�A��;f5���Oh���Ofm�e$z�.�Ӻ��+���Zw������ό�yh��낵Vú�O��?����?���?	��A�\P�NQ�p�B)+2.q.O�HnڐT6Z��	����K��<�����/��"A&t|�p0Y���	џ�'�b>U�����;;�Bv�3wov0�3��e�B|m	����9��,s�'��'S�Ʌ_�h���Jm���D��!7�8�	���I柸�i>��'�F7͎8m(�������U�
���QulY�L��ʦ��?��R���ҟ��'iFZ�Hԫȳh:u�qē
/�r���'Mۦ��'+���i��?��}���+;�V�8ikfH�3���c�<O����O~�D�O����O�?����~b����{(Tx����� �	Οk�4[6X�Χ�?�i��'|p�jc�� (���O
e~CE�|��'��O�:�x��iX�I\��X�&L� }�,Q�3L #C ��4��n�2�Re�Ify�Ou��'���3Z澸��S�p!6�x�,
�9�2�'u剡�M;�jQ-�?����?.�^u�g	a���t���P��-?!�[����ßL%��'L���a�T[�R�0Դ\���FN��D�Q㈿F#��|*���OR<:L>�$*E�K�ʰgNݡz}���5�؛�?����?����?�|�-O�an�,.<5��E6]�zS�^!"�y3�ß`�	��M���>1���!�3�U1s��ab�8b�]P���?Y�Mӎ�M�O��
T,��O��9m_]K
I�w�31� ;�'��ٟ���Ο0�Iٟ���G��Fн0Y�d��� ��`�rg�$#p7-O6-���D�O���-�i�O mz�A��` Mcq�ŧG��qM�����z�)�S",�m��<ɦ���E�ر��)�NcP��"i��<I��c���D����4����T7pz�ABM�
����Q�����d�Ot�$�O�˓-B�&��Vl��'�R�@'�X�1T��9]e�qH)�D�O���'R�'g�':�kp��a,�D�冗 "Ԑ���OZ��&�O�2>7M�\�`a�d�Ola�+��q^!0U)X�`������O����O��$�ON�}��#�,!lF�q�I�e�,�h��B�i;�m�T�'YcӘ��]+1b AG��9�Fy�� T�&g��	��������r`�T����'�t��	Y� ��xb�� 
�v��ǇB(��a�=�$�<ͧ�?����?1���?�B��\y�@ȄH�|S�oT�����E�%��kyR�'��Oy�jG�2Hn���K�O�"X�����rꓘ?����S�'5Rh�!""\� �*�1s�"y�H�-X��M˖T��$Dҵl�� ���<�#�ُx�ڌ!��L4u�,J�m��?���?����?ͧ���˦5�E��ޟ�p���K�a"bd�}���FLϟ���4��'G,��?����?Yf(�{������$h�Z�B I�^g��ݴ��$�>-�*��ĸO�G�_>�<����ĖB��C�ݸ�y��'O��'���'�"���/5Rh�f�#ZL!に|����O��Lڟ8�9���㦕%�����.0���A����͕y�	⟠�i>-����Ҧ��'��� �a�Zl��d���Ѝ���$��	I��'�i>!�IԟL�	�� =s��R#L�@��_�b�����4�'
7�|�����O����|�F/���M��C<�f��wfT~2��>����?	I>�O�$����R5�f��C�ƌ�ؽaBO�|dc�mƜ��4�$���<�ʒO�qVc�� �Tx�6uXŉa$�O����O����O1��˓"F�fk���T�&),	�P�	����x�Ȑ�'��Ju�0�hC�O��$�1���%,4
r��
� ��D�O��"m�����E)��P�O��܋6�
�b�(	r�Y/���Ӟ'U�	����I�������d��~��k��<(,yS�ʀa�|�ˡ��T�27�	wt���OB��7�S��M�;%�T�p悊33�d|S&f܇05�aR�����Or��2�i8�$��[��'��,F�M9���-&�Pbb�J�Q��Oʓ�?�� P:��'@%5.�,�����|p���?!���?a)O
al=X"���'"2.��Z�tBU��d�P��u�����O��'dR�'��'����*�V��)��E��I��O�����:?��M�t�ɏ��?�t��Oj��6�٨R1�M�sm�L�r���O8���O����OΣ}�����P��S�V��c���,��q������W x��'`�7m%�i��+��,�nxqD�#9��ycRbi����ߟ0�	F�@�nW~ZwЊ)s"�O����S*�=2�h�Ç�T1A�)d��X�Ipy"�'�r�'�"�'x�'�,�vH�wC�FLL`��I�"4���M#��H�?����?�I~��>��� "�6Tv�"2a��W�(X�_���	�&�b>�9FiH+U|�I�
B�<��x�R��=��Se�8?Ქ
p��1������X�I ����Sm>e�r�S�GD����O��D�O��4���q#�V��"�b�[�aZ��q@�(5�=��Ƨ#���u�⟴i�O*�d�O~�d�
Nh����?jU\��v��!dεkv�eӠ�R�a����>��]�qA��qE208nS��A=����韴�	�D��ɟ��`�'_0��ǖGذ�w�O��%�-O��Vצ�8 i>��	��M�M>����~���1��s����B���䓓?���|*1�	�M#�O�p0� ۹�N��'ɝ(���J�S.2,����{�ޓO���|���?��ib���+�+��1s�B�e&�|����?�+Oql�=�,��ޟ���r�.��Zn�qE�߽5N�y��B��dT}��'A|ʟ T���%=`� %/��4|���BB�M+$���d�����P韐��|�+�L���#�-vz[3�A����'s��'$���S��Sٴ:�x�3�ጣ ��"ABX8���1i�=�?�/&���$I}��'�x�bAl�$Q��mk�ۦvD�г��'��oM�!`�֔��2Q��q�S�v�I�5���k�n	�MO�@r/2�(��~y�'�b�'���'�2Y>�:��̄�FJH�d�|�)e-��M3e��?���?aM~������wt�d����0@Zނ��C�'vB�|����RK��V=O�x9Č]=�R��4�4q�p�K�6O����K�/�?Aw(7�Ĥ<�'�?i.��XOj�ɐ���6����&�R��?����?!���Vݦ��e�ɟx��㟠��^"
v�m�4�Z�;�6��c��K��
v�Il�Io�I2u�lm��Ŝb�h�§����8�x�B!�ѦI9^��|�1
�OJ�@�u/����h6���@ \�^̓��?��?���h���W�8�V�2mNI��|�h�#�f���Ц�LVݟ��ɳ�M��wV`TB��Y�W"1�W-]�h~����'�r�'���[�)
����pK�(Z�,��	̌G�$�Sc����X2F��
KrO���|��?���?���,Ynx9���e ���a-ٲU�+Oil��!�j���ݟ(�	p�ݟ�jdMkD�ف�>!q��Z���D�O��D)��I��w�jHk���8z`�) �-���l������ʓm��("��OZ�:H>-O0�ƥ�� �1Q�#�5trd��O"�$�O:�D�O�<�¾i�`M�W�'�Z�i��_�$������*:� �'��7M5�	�����Oʓ4��rc'S�O� cFF�<g��gBN!�M��O�9Rh�����#.�	��r@*�ʔ�Y��-3"I��`RVMx�5ON���O���O����O@�?������H>�)�6Eу��<��,���L�I�0	ٴk� !�'�?���iG�'����Q3�4@AM�����|�'��O���)��i���5;�� `��GP8	�tx���[t-T��'c���~��|�S������	��h8�ƈה���%�X[�� T,`�IlyR�w��e�C�Od�d�OJ�'(�zI��ގG��)����4X�'����?�����S���
�ޕ��F�x4|�S�	+-��1.�u����O�)�?A�&��ƲR/Ja�w'�O@.x��� �^���Ot���O���)�<��i��x;Pd��e,]��ߧA�.��['G��'��7-8�	$����O,r1l�)x����ݳ4h��ց�O~�$�"$S79?�O
Ta��i,��jK�"����GZ ��塵�C��y�X����̟��Iퟜ����\�Oy�x���'-`�`�q�ӼR���cm�,�ʶe�O��$�O�����DX��睬'��I�/Դg]����.�\H�Iğl'�b>-rp�ܦ9�V����U�� Q?��q��'CHT̓X��X��O�q:L>i-O�i�O*��bW+a��4��h�:Vy@��@�O�d�Ox�d�<av�i��Q��'��4����fam��]@DA�9���w�dZa}b�'�O-낫1%S܀�G�-G:�(w���e��K�rh:��r�SJ�R���|9�܌p�TaN"4�n� ֬۟���˟��ǟ\D���'ͬ��#�K�2����&P5��'|�7ˁpS���OtQm�]�Ӽ� d� 2��%;Bb�]�$��&��<!���?��f�d��۴����+ai����h�.�J�Eçf��\��#*bF���2�d�<ͧ�?!��?���?�C*Ť}��4x%,{�/��	��a+O��o�W��]��ڟ��Ij��ڟ8	所�s��z��/`\hP�F���D�O<�#��IQ;xs��p傎�4�$k׌!�	���SR�x���\H �O\9�K>A.Ot�� �?.x���ڤ+Z�����O����O
���O�i�<i��iZ6I��'t�k���;������<d�\JU�'ƺ6�2�I�����O ���O�`#��'��Xqk��Eh�H0:�Q�i'�ɀ ��6����-�Vs��s� ^�z���Hm���I����ǟl��ҟ�����4¸�H��K�Y�@|ʥ��?�?I��?�w�i�V��ϟ<�l�~�	�����[��x2����r\�c����fyb�Č������KZ60�fP����4J���6��8\'X��'�m&�L�'���'���'>h,R�J�3a���(�!�2Nؐp�'�\��ڴ#	H�����?�����ՙ@y�m�Bl�������I����O���;��?�YPi\U�<��s��E��Ȥ�ڟ��"��Y��)O�iR��~�|��8�bm�w+�8���oU�Z��'���'���X��1�4=���y�4��@ 4y�NH������?���W����B}"�'P��c4O�O:��94f߅fZ�j]�<��¦��'��#�?Ih�T�����c�`D)u�ٸ<gxJ3�e��'�r�'�2�'k2�'��	W�T}�G�$V��=	�dU4Y�t��ܴG\L����?�����<1��y�jA�q���{���\)�!�TٙA���'�ɧ�O�s��i#�ܬ%����qB�)��iH��.R��7'j����U�f�Ol��?����&��i�%�hdZ�
�3�&iQ���?a��?�)Oj�n�cs0U�	ϟ��	�T@{�/%e> �#uZ�Tk���?1�Z��	���'�$1�A2AD�`����(^&L��
=?�P��~��)BiŖy���$�?�'
	�������cL��j"L[�?i���?���?Q����OZK��R�yK�F�5
�R����O@5m�>s�$��ʟh�4���y��+L%�ei�� cx� �ƈ=�yR�'m�'�R�{�i8�IF ������޺}�rUb�h�80K���[+��'O�i>���矀����	�5˴(�fA�>����RAK�I8-�'�$6- 0+[���?�O~R��%�zb�N�d{�e�gg��(��<�sR�$�	ߟT%�b>}��H�&Y�v�BD�7M���Oˏ;��ؓUi#?�'�v���ӆ�䓕�$�#V��j&��B_V�����ݚ��'���'����^�|��4|0I ��oK� 1t�J'QA5A	,Af�����~u���D�]}��'���'�VP�%��/VXf��RA� G���(��i|�Ɛ�'G�=��	"�	��T���R�f�n(�T��-t���q3O,�d�O���Ot�D�O�?��BNŔ}������hٜ���͟X�Iڟ�Qߴ
]���)O&Tn�\�I�u�R$ �׮	�(DA`����&�������/�TQom~Zw�R��ԧ�|�i���'3�PCB�ݥ8���H�Iey"���8bk&�R�h�
6%�h`5��+��ةܴj�&����?Y���5x��0�P(�H� �z��ɡ��$�O���,��?�SA�!jtx�g
�W� (�O8N`t�"��}��Q����Jџ��ם|�L�U_���U���o@JurB�ּ�xJkӀIdMeԨİ��M�~-�]o�|���O�(mZo�H�	��jߘ8,��߀ 2-p�+����I��f�m�I~Zw],M˖�O8�'9DyVE15E�6�;�p�'W�t���S�ċ�0ВU�cl��J��Te�U(�M�����?)��?Y��$t��nMֺP���8%�-PC䀃:�����Oh�O1��E{��nӺ�)� �x���=���I� V��%Zu0O�� 1M��?�H9��<Y.OZ��-��5<��bg���5)��'��7�\�ap��OB��PsRX���o�KJp�tE��㟴��O��d�ON�O��	��M�C��d�5�\�J$8��疟��o�'�t�o����'%O��	ڟ��6GN���Xsh�`?��� �8D�|�5/F=&ڌ����4���x5o���۴]d�����?A��i��O󮀅`I�0��`J@X�}�p-]�w���O����O�DpC.n���c��\�h�?A��-��Ɖ�e9����Vf�	my���)r�T������_���ѷ�Y�D���O��V�fB�'�B�	�5�Jt���1�T`i4�E;(m��'���',ɧ�O�X􋈷o1F�{C��!\<��q���aʈP��W���B�M�7���L�	}yΞqP�R!N�QB���r�FP���'!��'��O|�I��M;׀D(�?�@/�#f<�k�*��b�T9 ��?�B�i$�O^��'Ir�'"��hg��{؋B����+��K`���i��I�\�.�I�����$l�F�0U�``A�l2��q�d�	ޟ����0�	����U�� ���J�g�=|h�M�?1��?�a�i��=K�O�o�f�O|1����?)�i� [$�$�P�6��O$�4�܈��tӠ�_L�82g��&3p���U#�R9����_t��l�Izy�O�b�'�B�M #�h���R��d�X�˕&QB�'��=�Mk��ۑ���Oh�'E� )3D�\����AK/8�2��'�0��?A����S�d���GI(`�N�)�^5Ձ[uwJ`y�ѹ/H�6���ӭD��D8���?~�8 ��B��
��)]�^�D�O|��O^��)�<aF�i
�!H�JǊ�t��C � ;�����Zd�"�'xd7�9������O�̫���< "�p�V΂A�ց�b��O���¾	6�#?96ύ�;���>��� 6�dс�H�e����/p�t�'���'"�'or�'�`�u0��*B�R|�v�T�x���Pٴ\���C���?q���'�?�1��y��6J"9�v
9�,�w�C!4HB�'�ɧ�O�F��սi��$ԡf&�pe�*2 ��&N	���DR@Qz�:�'K�'<�i>9�� jUޘXU��$Y)��3�O5dU���I���򟈗'A"7S!:N��$�O|���"B4i��gB��q�鐭�l����O����O��OJ��⌅1R�3Ab��6Mxu�5������Dy��o�X̧;���	��YA	�HEx��� ��J#��9C	՟P���x�Iҟ�D�D�'@t@Q�"Z	vJ
`�H��J�~l`��'k�7͎�#�d�On�l�X�Ӽ��"V:o[t!��`�	/|@����<����?���.��xyߴ��d��&5��O�����O�+�ny1��<4	|�S�|�R���,��0�I��6d�D�"IY�!�?
����.^oy�!fӄ�����O|���O���x���6�|�t�Q$�f*BU�V��H�'2�'�ɧ�O�x��,>)@l$����?[?�\�GaV�i��&������f^-�H� <�l{��X8���`׵g�,��S�ĊbQ��@GO]�[��a�Q�()��Ā�Y�d�7E��3G�i�@�]�'xJ����
s��&^��2r�Tp�xG��*�g�i���!�Ǘ�E/�,q5%
�la~�0楅UD�ǠV�W����_'xr��U��$qRUۅ�
�<"�#d��ay���D�[�k�t���P9L��6LϜH�V���%	>F\�0O�	l�|)��.4A��@#EG97�H�A���×�/�PxA���i�B�n�x��1�vK:7G¹����b8Rߴ����O*�O����OZU�G��pz�gFr�L�8 Ł5��,�ʺ>i��?���򤖊=t5�O��g�&�`E��JrO�6=n��r�iR2�|��'S��^�]OqOr �u�R��Zq�v'NK��q�i�2�'�前6t�H�������O��I�Nz�i�;e'X�iq�.Y�,'���I����O�����)��u�f��Ʈ-.�e�D�Q!�M*O�A����y��џ��	�?���Ok��S��ˢPX�T���-�v�'��[�|���,^���ӡ�
P�l�VD� �FP'�<6��O��D�O��LG}�]�4b0C��Z���q6oS�hJ��$�O8�M�.	���'|���J-`�>p�q��2KJ�%oD$-��Uoџ��	ɟ,�p�����<Q���~�e};l]��LX�� 	�aĜ��'!4 p�|��'�']�Y�*�+F|�TCG	�*�.����w�P���1L`x%�'y�Iş|&�֘</����ԤِgҶQ[p��.I�Z���0�N>���?����Q8E*�Xyt��X�� �f�<!�L�9�"RU}�^����l�ҟ��	/(�vx0$�K�6f�i!��B% �|a�	F�I韴��ӟ �'�ir�a>y�!�P,k���Y�+�W`��$'�Nʓ�?J>���?ـ�0�~�nD�z�­ n�>v=��b�E�+��d�O����O^˓a�Zi��^?��	�z������b����-ɓ$G(���4�?�M>a���?��0��'�l�nB�n�^*v����&-��4�?A����dRT7��O�2�'{�4BH�`��9; �6TJ<QA��D�v�O��d�OPLy�I7�IjZ���wHB	@p!�'�4 g�ߦ9�'Yԭ1��a�t�D�O@�$���4ԧ5f��A����� *�E�"�M����?���5��'�q�� ƨ��Ō0=(j"� %C�4�iE��6�`Ө���O������'K�	.1 0�F�(ޜ����Q��4"A$C������O$�Ks�h����24[�1r�E��p�b6��Ov�D�Od��L}�S���	G?��g��W<0\��h+Tq�m&@Ʀ�%�8��� �ħ�?����?Q!̕4n]��BG�r@��C	�~���'�֗
3������'e�'i܀�Nډul0�d.S$�J����!��O8�O��Ŀ<Q��1�BL�B�
�mu� �H��vj��������O��D0������&�T��@�0 #9R�bP	f�oZ�����?���?�)O��8�`��|��m�\o��2��I�[wl�u�Is}B�'R�|R^���؟�[�V,jҮ���3�~��+	���?�*O`��(Y���'�?E��m �����B�^c���HCF�����O6�!�.$'������ � 3��+Tn�Az��d�<y��L��db.���$�O����L(�98Z��dO$ט�:��x��'I�IY�6"<��!۸ �7kD������S>a�'"�$ԓS��'F"�'��$U���bڌ�8�+*@���gN�V�6�6��[�d(�K*�S�SF�����M�#/�5���U�>��7-,��mZ۟��I�D��;���|��`3m��Y�h�AĐ�A�&!q����'E��'�ɧ���D2�L��:�B��0#��^:}�����M���?A��+T�XJ-O��E�$�92`�e�q���G��Hn�Gx�&2�	�OD�D�O��p�Y2��YaSN}�P�hV*Zߦ=�ɷKȩ8H<ͧ�?II>a���bZ�Y3�>�P��ۅ2��4$�X��|��ϟx�'d���J&�qB�_:{k�)2��N�ojȡtR���	�?���~(80��BW��]��ys&��M{��n��?)-Oj�d�������I26����q�)��7�O\�d6��˟Ȗ'lD�4\S���"�n.��/�~}P]&����my��'9vDzQX>�������'�+Ƃ R�װ�2���4��'��R���4�(��|�XI�������Jp�үz����'2R�ږ����'�?����CF��c�f��"S %|}��OGb�Ify��'N�����u�H��B�	m�*R���g@-���Пp�pK�� �	ǟ4�	�?ɖ�u'@
;p����%�P$F�1�MK�����N7O����U�w��%:r�@򃓝tB����i$�y��+n�����O<�������'�I�+�!As����(�!�C;�6�qڴ4q�p̓�?y���?Y����'kШYe��h�>���R�x�ٶ�d���$�O������'��ݟ���40����`҃��тe�7*0lnZԟH��֟�[�
n��'�?���?��NrZ��J �2�UhG�		 hB�mZ��$��f���$�<A����OkL�>k��0�E�[�m�r��V<�ɞ���	ԟ��Iџl�IJ��'�ꉚD�ן<���qbC�X�(1a�:I�~���$�O�˓�?a��?�G�7|$Hbr��9!�,h`.҂Wق ��?���?����?I*O��ɦ���|ʱCL)O3���Ȇ��X�i�����'WT����ޟX�	=6���	�R��tZ�!ӘYg�1�G�y�Du��4�?����?����dP����OTZc?�M8A�	"ra�g�Ql\H�a�4�?�*O��d�O���	���|n��q�ȑt�4k��e��-؏g��7��O��D�<�Ǜ8)����p���?�zP�*S5x����sz��8�%����$�O����O��s�:Oj��<)�O�� 3@@�#m�gķ ĸ�޴��$�S!$l�ޟ(�I���������(CW�S,6�z�I4��2�i���'��ʝ'V�'�q��4"�������(:��|��i��y)�.u�����O��d�,��'t�)y�#���%_�H�Q����4�l���?���?	����'�HybF����v�A?}�ܴC�ik�h��O���R	�`�'��Iڟ���kUt�U�ےc�tDѳ&�+2F�xnZC�Im� �)��?��O,&Tb�!��J�09;�k�j�Hxb�4�?�S&D��ey��'%����سF�vH��C�=0)��7	���I-V�̓�?���?���?�/Oޔ��!6�<h{���)Q�E�M��e��'���ʟ��'���'*ML�FN�J0�Y�f�tm�Mܽm�v���'�R�'��'b\����K��4F�%&qրӑ��WmRp����M�,O"��<����?����ʍ�':�2�C���(�"AAz�%i�O����O&��<��^*G�O��iŶC}���&E�|0��j$�k����-�d�O��C�H��$&}BoݡT��Ys�
��]�siS��M[��?�(O����j�՟��ӥTt:-`��*#�~����4� �N<I���?!�;��'���@�+�^#���|�!ș�.��fU�ĩ��û�M[�[?��I�?]�O�M�@�oy$��ch�m��ꄺi���'F�-��'��'qq�~��ƂC=0|5����&/[z��$�i��\�W�o�����O8�$����%�d�	4��"�(B7I��Q�0�ʼ�۴W@��������O�B�P�
2�J�6w��a�f�	�6-�O��d�O�8`2�C�ݟ��ID?Y��
h,��d�/IXeYqD^���%�$�oɼ��'�?9���� 98'U�e�ų�-`�����i�2�L,xΚOL�D�O��Ok�ƛ`���p@��M<����&3���<����oyr�'���'��I<|���W�F�"7`�*1�E�T�fN��ē�?!�����?)�cI�Y:#a�2+��}���R��ivjE��?�*OF���O~���<���S���I�1>h��IpE�+<���c��	��	ß���[�Iß��I�BQ"L�	4|v��cR�)�Q.q{le3�O&��O��<)Ň� 18�Od@H�r�ROH��3F�N�~��W�m��$#���O�_�p�d>}RG��S�(��V��?G9�ᠴGˑ�M���?�/O0hz1Hi�SΟ����S�򨠕bQ�r���CnDt��\JJ<!��?9�oY��?aM>��O�黑&���jC��3v��ٴ��$.�
�l�����O����N~�I=t'����K�~ۂ5��&�7�M����?	u��"�?�N>���4�Љ&���tNͧt���$ ��M�����?Q���?Y����/Or�'2M���c蜎{��@q��]�6h:4�iP޴+��.§F�26��Z��y{Ab�z�@}c��� �!�d�<O�QHr�F0L�Z�ޅ��'vHBpo�+q�x|s���n&�R�d�+���7ł:�H���'OrLbP�
1e���򬂁cFv	df�!Yp�2��Q�P CE� �4�`OS�tBVx�Ռ�z4j#΅,�Lūf�
E� �ˆ@B�<�d���MV9[�.� !� n�Qز�42>�S���"Z��p���?���?i7K��?	�����!Bܨ0���Z�i�i1���;�{b%��3'd"�eP%"z>���3{@������p�(		u�.a1��	�=� �7�X��4�M�'IN����?����tR� �7�m���1�>�hOܢ?�%T7Ka�t�^eI�	#O�C��#����$d��gLH �I�d~L���d�<QCA�!����ԖO�6ai����s4) ��h��댫&(�'�!�k� kcd��Wd��I"��O�ӓdx��Ca�I?��!�3.N�<�d�	!
8�@cV'yS< (M|�T!�6\���Y����x߮�J��I�'�����?ɋ�$��3YȂ��"KۣY��*�nP��y��'�n�c��XZ��$��U����~`�'�����լ�����+��̀�'���Qh�>�����C�A	"�'���Q#T"�5o�+�Ġ����}ڼ�����K��A��FA�>�T�T>��|�I�.�`�QCB�:pC��$��Y��dh����J�24�G�~�h���S��?��"�.�m"���&6<��O�;+�����?��O�ON�'�,���b�7�\m�2�T*ud5�	�'�,X� �3��pgӯ�=����L���閧Z6�����^ւ=c�'!)����O��Bn�J~L�D�O��D�O9�;�?y�=uCH�K,b�zT�؛(�4��_0׬���$³t%�m��|F|2j܌�t)�gѻf*;��7-�
M���А[ţR���yn`���O�t\�ҮH̓�b��偣l��E"�7m2���R[8���&�V�f�|���O����O6�4��I"C�d{��qAP)Pqla���HO��%�`[3��[�$8��
q5�ɩ�4@i��|2ū~��y��wr���H�x�G^˄	��d�0��2,4��#ς������U1�U[��V,%�l��Cޒ6m��ȓ���yŌ����%�@9R���ȓ;������t���� �Ts�,u�ȓu��Z4�Pz���bA�߻y�P�ȓ`��A	��P##nͻsN�/_�,���Y��T;VJ&qw�AI�)Z�AC��ȓJ�\, �;J�E�"�)&/܆ȓq�b�r�*�f8�X��,w4��ȓ/�>)BM�+=e,}Z!ǊT�~��ȓ&�"R $�W��l�#�F�vR���i��1qAS D!��3��$K�p�� !���$���+��a$��.󢐅ȓ\�Bh�tIW�CP� �j�G����ȓSz<<�
�-�!b�)p~���ȓ0����4JX�^��Ȼo5NI��\LqcG�0��X��LD/V���ȓ�F-y�I�~�|�;���f�ZI��t�$��,�CZ�-�	�"wt�����H��1�����Z)z����ȓ/⁪D�ܨ&��L����?��$�� � �E �1��!XW�ϵ;��؅�zEJ�2tDԂ[���룅��9?v���S�? ~4
�O���d�3�. "�8��"Ol���՚��8�B�¯#��4"O���Ӣ
�-�r"�I����"O:\�6+^�d?d�%ARR�8Q�r"O��2�'��z�µ`�'P~���"Ofظ��NP�	��O_�8zF�k�"O��ɶ���k�E ���}o��P"O���*�9	P!���Y�ݛ "O@4��$J'mH.1ʇ� Z~<U"O��h� g��e[���b��"O��iůUh��5҅��QR�E�f"O��)%��Mu���@��9?4q�"O��1Lۂ:5\�+@��8L/UY�"O�\6)G�Y�踆��z�fp�"O��Sf+����I� ��L�"O�̲�K�FV�)P��l��""O8-s�0�h�0L''�Ʉ"O�Лdg��Wml���j���t�S"O"��J��W!r����=�0M˄"O��A�͉%!Ty��/~rL���"O���&��=dUH�iv�ڨp�Pp�"ON����9S�B��JU4I��Z�"O=�B�ޒ>�X�!��� THp CT"O�Px'lU����1f��:,�2p"O���Q$?P⌔Cw���Tq5"O�D��ŕ�F�n�Qr\1.�ˠ"Op����M���n�`��"O"\�s���� h�eC�`� �"O�Y2 �]5>b�3���u�JY*5"O¡+D[�b�`�4#��f�
"OP�BL��+"���Q?'��Yg"O.QX�c]�w�,��O=3&t�B"Oक़� Ā[�`
3��0gJT �"O��jU�	�D�$� ���8�8���"O�U������PW`���%H	0�y�ZZ"�b�+g�HђF+ڮ�y�C�����u��gs @�N��yR�P6l<�P'�K��큳���y"@�$o��hU#�.��#D�U/�y�e��L�JlE�g��v'[��y��23x�劆�:� �e��$�yr�̧rs)�$�::�
��d�A��yb$^MX�[�mK.,@dD�L��yR�:P��!1
�`��0BC�y��(B�ib����[x�T8q���y��:8��5��� PX��*ۣ�y"��}���A1��Fٞ8 ���%�y���:8��9�v-�7C8ţ�E���yL݀E� ��BDݲЂ*H;�y҄�����ԍˌz�~�h��U��y��,+ZJ���&͡x����C&ٯ�y"�W	@x�� ۲����+�9�y���C�2䛵&���-�p"�.�y�P�3��%��ż	���5��yr��	�Q���~�yZ��-�y�����G)�F@�Y��,���y"���)�lxk����1��kӍ�"�y��@? ��0e� �)�T�����yBƍUΎ�[�Ƅ8S`6�)��ש�y���.`� ]y��@�,<1�tLƹ�y��^�h�\��.(��0��*���y�d�79.�A�����a�-�y�ꁃg|}�dc��S��أ�)�y�5�D�a��_�����ң�y
� �����Ю8���Q��ɗ4Y����"Oh�[��.rs�M���2W�ɋ��'[>ep'�ޗ��DĮd[�[������.�m�!�LP(t�K�A�B:�A�E-�,|{qO0��@�9h�?�a2c�:_D��g"�����.D���%ìl[�`iэF�<�.X3�i�X"��<qi �gyrmM"&�n ӕA�i�$������yR昗#�Ep	e��=P�oD� e�Yy��_S��}�&B k�<�:�NK'Z��E'��p=�R��(o���'�p�fn�Y+�49��$u�xl��'6"y�j�I��%��G�y��p�{�ݾMn����B$W%tҁL�G�<,h�o;"��3�¡>��iQ��=���٠I��!��$����]0-�-�>9�\?�c�J�}��Li{�*��:H��q b���ܑ�5�[j�<9��K�w��h�rj��]'(\�'�Df���$Ks�q��GT��xk�F�{�O���3�`�f�)j�F�;�u`	�'���
��]�}٪��J�(9�  ��a�P(�ړ�J)1.t�ѵ���Ϙ'f>���a��o^�1�G�S>�b�'����vG�i��h�I!%!�I�/F�g��i��ƕ�nYDPʎt����u� 9�f<8U�֟TZ9�B6O��.=��ԩ�+�$"`�����'��r#Kȳ\6��̅�@ hy�'p<4y$C��`�R +$��i�P��OؤCPDD-:��i���fd)0��	����ɧ���LљfȌM;!�"����1�M�%�N�):�cԬ1pHw�$>�h�����S��jt�M�?n�҄1Qg�,[!��K�|�Li +J���$�w�M2P�Ӥfr��゠� ��0��I5.�s�!G!y��:Q	E�:~�a�ቛm����@Dι*����g��Z��M��CI�|Q�s�艌��L1�)=D�tX��J-'$d�t�3~d�P��<?�����g��)[g��-��i;���$Ґb'�,�r�2�a�Q����"��(� ��j��%�� ����M�ౘ 
p,[�g�=���"�i�1�1O�[wlP�|��iH���Kg�(c��O��c�OB ������8��	YY��1�"����QS�X)W+:���=C��xzU�9lO"uX�Y�r�D-����sPX�2�>t�>s���d�1>� f�"���{�V	sW�~��ݗI'��8U-
�U����%�k�V8��	y�<�5�ĪʼLJ�6<����n�x�'-F-fe+§q��Aq����MG�_'�9�ȓd��WkX�lB�hRe ��L�@�ȓ_�lӧ撾qJ����;n2���6E�����NO�48'.���ȓ�*�����n@��;��O���ՆȓV\���k�"W���sM�";����tu,x g��"�(�Q-#�|��N�@@-���DWc�����b�n�<��),n([0!UF���3���j�<a f�,}�n\�M�m�TggYd�<Y@��<\.��C�A\��tgc�<q���]j^��s�v�A�C{�B���vKM8=
�鉃F�V�"C�I@+�����3"����c�[��B�I�r����B��� �A��B�	X)��f�V��~�s��M;0�B�I%��,��'�%��ڣ�K�B�ɐx�Vh�RE��X��d]�C�	�v��q���iO��G��2N��C�I�.Ԭ��@�-�Pd"d,ȇa��C�I�4D����
پR�x2�h[���C�M��ջ��^/
>|z�AX�	��C�	�9�1��#Z/�ļ��A�zC�IR��DՎ6i��j4	M =��C䉋4h��um�<~��"K�n�B�ɑ<D�2��Z�@�Px D���B�3i���BG�[\@���f��=:tB�)� �\�t�Z(J-R��@�U��؇"O�ɓE��#0�I��4�� ��"Oz�$DD8�|Z#Cދ�`�Q"Ot0��5f�2��%�
������"O��,�P�&���o`�(�s"O�\01�B�2�*=�Fo�Gn�"O��� D+��łB� ά$�"O
5�2���+�P�K��[�D��$��"OS�
�	I����FV�  q"Ov$Q�@v 0����N�V$sA"O�x�ee�� ��ى��$Zv$�c"Oa"6�M�0cj�H�hP#:�^�"O���Ã+K��+$W��""O�8��'Ϧ"�zuz�ɤ6�}�"O�*
��H�󷈎W��8�"O��עO�x��Ç!O�p���"O��@gǋ_`(�#�`�� ȓ"O��y$`�;�x��5@q�uI�"O(u�5ir��;l^+��*�"O.ss`�&h�<)@E�[��[�"O��� �5A2��V �m���"O�e�wo���ڹ;����yVn�("O�MZ㯔xԲ�ѱ�  Z@�"O薦no�A�AW��hq��%� �y��< 
�1�Ӑ���(�!�yb�% H2�g��xΜ�9Pԍ�yBMU�b�Z S`\ݦ�Z4G�?�y��(:��<�G~x��T�y�FT "r�K`��uMEPׁ�yi��F����e_��dѺǏC/�y�!�"�� S��v~���GcΫ�y2�5�BX9�͓�k�|�`�/Q�y����cɏ_��⦀H�y�� -L�ˇ�ˎKfx�I6d6�y�� �jAk֦�!W�V�"�A:�yR�B&M�B��#�-H�8�ae�D��yr]>'~�5覧�Ik\Ac4�U��y2C�=1 ͙1�ܯA��k3����y2぀��$���H�W����6�y$G6R�"4�E%��|�����BI��y���$�u�L �{�^l���ʵ�y§ڙD⦼�o�&v�Xp�J��yBmQ;z}�ȉ��F��<�狃�y�	Is�D�(\��`�L:�y�Ć�+�z@_�R$x�� X�t)�ȓ׾��`>8�&�kjAL@*y��TD�EPs�T�SW��Cs�ՒF��u��@�rѸ����nF0��(��ȓ"e�C������궼B��qB3D�8!s
�/SUD���N?)���7�;D����lM�Ĝ�§��v����L8D�Xkw�Ǚ��2�V.�pK2D�0#c�Q�r�(��h5ұitH/D�H��.˒����-N�<��a��N,D�����w%�X���U�6BN6D���ǎ�h��=��
V*�����2D� �tJ\��r`u�A� Q�i��%1T���%L��8_��A7 ��.�x�"Ov9���|��z5M����q�"Oh�[���mz1d�T��l)�"OnL���R���y�e�X�.�<1""O.Z�*��J����	eIx�d"On����ɼ(x�(cW"W!��r"O��ag+��~�h�!',L	@$�	`5"O� 9�t��8X*����B���"O��cA*�*Q���J�Q1ƅ)'"O"�˧E٪9�r�bvJ
f�p�� "O<�1FP�}`���o�S8��""O�,�aC�Rp�8	#�ʵS��}R"O.�C���Q�JP���,w�l�d"O�(�V��~��(�Qa�8
�j��G"O6��pȓ4wl@{3G�|�d�� "O��!(��v�"��'�ι����T"O̘�,˰\����t�,�x�"O"�b�c��~�
�CCԳR�.�yr�̨Ol ���:��I�# Q��y"���,���(�����Q�d�y�T�J@���
q�܍�B&��y��&~��jd��t"|8Huχ��y"!<T#�`� �(;�>M�a�Z?�yGځ�����N�,����ѭM��y��Z�[we�֋� �L�ڐ���y"��p��𳦈R�k���a�0�yb 	�-�X�0Ʃ;I��Sq�y"��?	ߠ��D8��`�Җ�y�d�wHZ%yw煮21�! T��yr%P!/���0��$��djB���y�̥b��)g�������	���y"�_���%�H
d��s�׿�yb�G�1Pu@���%���A� �y���#��)�k_�W� �L>�y�&�*�U��e ){��ȣ!���y���v�^L�!Øo���� �Ԑ�y�DQH���%�VJy���y��E�e捃�B�Pxܨ��蘇�y�K�YD@�m�C�V�
���y��5<�H����Ǒ�
T��A�y���	���G�n�����&�>�y�eF�{���P��3~Z���֛�y�`�J���C�z�L$zF��'#N�B���5�`aѢ閝"O,i�R
)D�����5�a�
S�}�ֽ���1D��!��SZL�͡��Ԍ@���`1D�|�f �Q:\E �
T��+�-D�"g
��B� Dg	Q�bB�xc�b)D�t`�d��k���33ˑ�g$0Ճ�'D����2r�iQS�:��]�9D��P�J�h�,� b��w��AJ%D�*�Cؙj����A/DA�u��"D��y��ǑH�t�����V�� D���ME.U���W��>I��ª"D�� "HC %�$N�?a�=���%D���4k��t�.�Hr�A^/z9Hw>D��K' FZ������.6T��6�;D���L�v~R�[Ei��aTFO��y"(�6��;v��m�����I:�y�E[itV8rT̓k��A	$�y���[����/ޮ`&PS�F	�y2�� R�<��Y�X<��$�*�y"�:-P�Q���+y��\���.�y�,B�8� �Q�J ��E ��y&G�g�
!��o�"y���(D�E�yR��Q"`x��H$w'��\��y��Q���C�~�jd@��y)��Qw5��X<|���z�h���0�XX��	�X��ǋ	�&�ȓY&mZ��K���S�@9>I�ȓOw� 3�J3f����oƹFUʱ��S�? ��J�M@�]�D��]j��q�"O(��HQ��(#�Aڏ_�D�i�"O���Û�6b�c�ߦX�"O$,��'0z�g`��7Z�r�"O��.��bFA1FM1TT<��0�D%LOb��f��(v<i8�L�7m�@
�"O�ؘ����Z9��f��C��,[�"O=3g֒
v4�i�+�6+�V�
G"O�P)��\cnI�$��t�Ѝ��"O T��J�'s�hu@HD�7�
=і"O�`��L�<�-�"[�R�Z�@"OL)�b��1|��1�D�R�R$��"O
4!��K-1 ͉��K�DL@"Oj����,������ř+����"O^��b	��h�Dȉ5*G^�Xt"OeK�	�
��) ��%C��� "O���0�N�NW���S�|��L"2"O�������S�T'T�\�bP"O� �t�
�!����,��W��Q+�"O�iJp&�_���z��M?l�t8��"O�eJ2��(�ވ �>�QU"O",�cjSY���ݯ�P��"O��(4Ι��@�k��^+>�Z�C"O�@�Fj^�e��3��^��,(���7�S�<[`���(�'WQ@�sv��>1O C�<$^�\rDm���h���b�	s�B�	� �e����ti�U斴@�B��3k�R7�B�%ͼ�B�$Xu'�B�)3�H	���I�ä;��X���B�ɐ�b݃�*�`ʜAa�=?�B�	ڵ� H�����ץ����C�I0"�����EҨQ�|��A>�C��n(�K�"
)W8��R���8�C�I�P�A�#�
�y�fa!�AN>C�4#�U�EQ�dP<��QB��C�7_o������7(��шx��'ў�?1�6K��~�&!c[�r��<� �-D�����R�|�s���4}��C��6D��zB�9n�q����6,*��I5D�����%1�Ub�Н+ET�`&5D���r�ޯ��8 r@��= �EP�(2D�ۄ��p�����)B'?��t��	4D���u��C�(��ĕ�S��zC1D��J��\�m2��ai�W����0D�̊���"�h�S"&/ :����f/D���ѩE
Z�����	p�!�$(D����_=%��z�B�<��Í0D��hf��!���aNUr仦�"D�,2P�جVV�L"�)��p�: !�b-D��a�V�ߞlk���$�i��=D��iFL��,Z"�Y���v��a��9D�����K�/P&���ς*��xQ��<D�\Iny�~��C���FY�,�'�=D�������q� ��5$��e��U�/D�,�t��(u_p|��H1:>���,D�������>lDm�*a�R"�J)D�8�b���P7�	���C�Jx�!��I'T���p��ϴ�{``<�B���?|O��+r!�P��(�b�X&Y����"O$8���\$2�X ꥏ7��,�"O6�@��7w�]d�$�`6"O����1wa�hA`cǨ-��"O<��&��7�QˠS�)���"On���@�".�Rr�*G�
ތQ30"O� B$�Vc�#Hc <��5w�N$�7"O��S�J*!jL����S�V�Iq"O��ѴIZ	@�E��l�=��)�u"O�aA�*�\�t��˟�����W"O"���ĥ�Y�#��
I{Z�A'"O~XX6�1q�e�F�ͣ0���Z�"O$��F:݀��C�sy���"O:��BM���0`��a��vD"�"O�܀��N�L�I�`��
�*C"O�4��3H@���mDb-�a"O0|�w-��H��	�Ab8��*"O}:��G1�u�!�+<"O�]%,�[�=@��=���$"OxhB� Hۦ�:�A�r"Oܵ�0K]0!������ L�a�a"OJ��"c��$Ғ)����7a6�	�"O����?��i�G�]�Ul(�"O�i��́:Sw��?�>)�P"Ov�1��yT!�`A
n���)�"ON��g�^���w� 6k�(0��"O�%�%AO;0z�=�ň�q��5r%"Ob}�P�W�I�RBڷ<�Di�"O�U1 R�<wJ����W�k/��#�"O}�Ꮔ'|��M��/��4{vU+�"O� څ$S*�͛���0v��×"O�)8�� 3Z�t/��-e��RE"O��� j%Jl��.ɕ*��đ5"O`<:')�Tɚ|�!�A1�\PyD"O��"��L�'[Z�A�ּ��ѓ5"O�M�A�M�hua�*ՈI{,p��"O>�x'허g�	@*�+Xz�u�"O�l�Dh	�;�z �]y5"O�� 
�.l��Z�@�Fo2H��"O�i��̵5�N4[5ȌGi���"O���7���6G��1P퇱)]ިB�"O$�
r8�F���6~W�I@"O�l�q�
MV�܊BK�c���5"O��h�#Ѫ�%�qH� �B��"O�AA���z4��CB�t�p��c"O����B
W�2�P@+}��y8"ON��c�@*E����6��Ȳu"Oc��?7%xH �X�.�iu"O0�bc��3)|��7��V�T�zR"O8ɰ"�J�X�V�!�A��l�$�s"O�D����""2�1G2J��D0�"O��YХ�%�Ġ �%�]��""O��ԛ[�<Y�"��'B֕:�')�,℩O�QҴE�$G2k<�i
�'������HV%d'��I
�',�K�@ߡD�$m:6�X _�0��
�'H\-sP�)`�`�r$M�;)}bX�	�'�.`q#J63m:�³`T!A�}	�'���:0+�9A��B1J����'��t�t�ͻt���R2 ��>yʽA
�'zx{�H�!\���I���a_��j	�'u�AP ߟi3�H&׹,�e��'�Fȅ���.<s��"v�B��'���iC���2�&Ğt����'�z�SE��o}=�S,J�x�����'��Pc�'J�*�,�X<j�D��'���p�N��,*`�!ac�\��Ĩ�'����qaB�����Q"��A�'ݢY��cD�%��7h�>].�q�'N�P����rd��"F�Ì��z
��� �c�*�+Kz�l��*˪1����"O"!)�D�]�	�/Z��\�ҡ"O칂`d��A `8�T�/�d�@&"O�h"@�Cs���%L"3c4X�"O����=S0�E��+ZcJR��A"O��i�T1Gv8y��E�d�#�"O�0Ѡ�.-�k�$^���sQ"OXx�G�+X�`P�g$S06���b�"On�+��،�@� �,�p�7"OX�R0ŝO�l��d��d���7"O�T�P�H�6Zux��ecL�#�"O<X�v���	���1��6\���c"O(	�b����`��>֌��Z�y �8>��� 1&R�1�n�B��y2CY4D� ���:'[���(�yB�1*(�my%i�3��)j�0�y����b�r���"�bb'�y�)=)Ȝ���r�\���%�/�yRI&w{�HDHLd�N5�w�ż�yb D�6ЛuB]�[oX�v�ׄ�yb�Q2/T�1z`��<XD�F�Ӆ�y��*p�<��D! 3�z��E�y� �3�:h��nS�-�h35J��y�% $q�5��+���h;�[#�y����i `*��@!�k�&�y�\�M�nlx�-ЏG$�J��(�y2�B(G*��I��\�h=��Y��T��yb�ޚ �q���_7"�Jf��'�yr㇣\�8Yh���0�`���y��9T�����ϵv֬P�;�y���,�8�RA��i��@��A(�y��1x�`QR���2���Y�۳�y��/b6Ra	ы͕v]���AL��y�<լ%�FG��@Z�DJ����y�L�-���7N��u�Υ�y2_��H� �g�O�%0��N1�y��a����J-���N��y�5B�H�F�
G�V���m�"�ya�6$��(h��A!EK�`�u�@��y�hN�H�x ��jA6=����GΎ�yl��6.���5aޯ6��@�Sa���yR��=��4�˔^PyC/�$�y2ƕJ�f�CK�A�̜�Reԝ�y%�-a�T �˚:��%y�mK�y��]�6�T�,�����yrL 2��苠k��-�}+�
�>�y�m�/������'U.�s��y¯����U0#J�! �:a�B�Z��y⭎(+V�$ǌ;�J����.�y"�F�1�v\9��^5H�: �!���y��2�D����<��쇘�y�F�w)���g��6��գ�k̅�y���g����E�9�J�rB&�(�yBg_����@7�J�[L��iW��y�F�� �LԸ�ݯU�|��e��y�)�
K�L���@d�ŉ#�V��y��-�L���$ѳ�����΅��ym��q^<�kpJΐq�� �ybC��W��A#�)�2nj�PÚ��yRd�Q�~���ɗ��H�삾�ybo�� #HD�Dj$>�
!i��yc�1.�pT�� M�J��s	H��y"O� 
�Z�
dYL� #Tb��y����)���z�C�B��i���-�y
� �a� ��|��91�G��\e&��c"O
�d �%Z	��g��",l��"O��J�L$�ܨ�6�ʝ�\��q"OP`�2KZ�\@�q�c�W;���1"Oh1@G��38>�PA"b�'F\��"OԕyÚ�P���R "��?m���"O,�8֪]���T�˭?C��Yp"O�t���?�Dm��	�y/���"O88vh)n�h�1��zr�!�"O���ʚ3�B��H�F�Q"Oti�Ĉָ1���Z�GL!�z�yd"OPРGˌa��A'^(:���e"O���놽T`ݛ��5u>�x��"O6�y��U �5�6�;K'�9��"O^�� �>J(	:�Gl\谔"OXD�DI%[����D�Z�l8�p"O�=�@�ނWj\�p�¾�B�(�"O��sqV� N�UR&l��Ph@"O��r��Z�\�AR
ٌ��]CR"O�9��ҙ6�i��(Vo�j0�B"O��bC���z�MɤƋ��� "Ot *�Ma �i��Ʌw��蓶"O>�J���t�ZI�H;j�R1�D"O����T6$#n��Uh�Q���"O�ؚrL�7��wH$��a��"O؀b��(�����'ކsL�D"O
l�UFT� ���A1�?km�1�"O���U�\���! @�^�ESrX�F"OѢ�
��+����㘩~F&�j�"O� ��!.���zԃ޸8L��"O*l�ˈ.BbX!3���+;E�"Ozt�r�ǀ5�`�R�)�2����"O@uQ&�3T�y"������"O�ia2L[����1��Fy�K"O0L V�����`Q��&l\,3q"OTtJʏ=C�8�L��$���҆"Oz`Q�J:T j#��c����"Or���p!C��Q� =A��>D����aS ��q����T��<El)D������*A�]
dAܛ'R�pq1�(D��$.K  ːЀ�۞ [���%D�tJa��8%n���c���{t�!��#D�x�H�~T�da�oN���!��0|:��y���Wl^�@�H��d�Y�<�C���m����/I�I��9�R��n�<��H	�h<"5j1��3���#�Io�<9����A�l��a%�}*f��T�<9�C ~�����ӥ[�YB�c�R�<I�%�����a�Р~_�8�@�T�<��-M��4i	q����	��D=��ɺ��I��Nm��@@�2�"O
��B�e���Y�/�>��B"OVa05�_�9��C��^��6"O�Y;0极{"��@�I���� �y�Ǖ86��x��I�z_֝�F�I��y��ј.�V���b�kަ!�nÃ�y"-ޙ�6m��D���t�n�y"��*^ʄb���4m�Qԥ���y��=b���+6�0�Z# ���y�$	�8L��B�dܦ9��9���y"hC�K@�!���"!����yj��c1��0���&�ua�B��yb)��w��0�I(Dd�X�-�y�΁����O�*@a8�%[�y
� "�	TRo�='̔iuDy"O�h���I6��E��Z�1�V	��"OtT`�5�f!��
L� XnP��"O��Ů�.1�mSU�Bf���R"ON��3���	 c!9��q"O@�8t+H4]R� ֦�t�r=;�"OT��DHʏA�:����)2�]s����O��i�5�X�#v��&mQ��S�<T!�d�M�r��닭nd �΀ ma!��S�#d4�㉟'B��	k����v�!��'u�*�*�i�A���[����!�3Ȱd;eh�b +��e�!��4z�h��B�`����9~�}ⓟ�Ň�l|"K�Јxk�Z�K,�O��?�$u���:N�(p0F�d�����|�\��2���$%]9k��@��g��5��d����hk׫��R��<�ȓ�2��BE� QrsE�ږ@� ����4�0�L�LU<���@ƜA����aV��%L�80Vy�W� �9|)��m�^cЇ�	�z���P�:�xG{��O����H�`� ���^�N�6�0�'����Nх[I2�0 ��EX��	�'�h�Wo�n69Hw�:0���0	�'�~90�@ A�&�Q��D%z�:���'F�k�g��9ǟr)�US�'#&�f�h|�zU���%'Y�<&�� w�i3�"K�9���q�,�ϟxF{��I�����W�$0B�	�΅��C�	�xW���c �6B��]��ݓ/ǮB�	��t��`��bR�Ceܒ!rtB�^+p� �&�ZM
�!���uyB�ɚ|�vaPFj&)��D�'��2v�C�I��O$r��{�`�!r'pC�5�<M�0��i7��r䫌=:�&C�I=v]#Ԉ��b�"�3'�C��+T]`�w��.G�J�"�c�:-��C�	9�Pq{��x�B�����^.~C�8E�6؈B��,$kSK	�U�TC�Ɉ6J`1R�ߠ�D��O��ULC�ɐ&u1A[�s���j0ϹT0C䉐�-( ���x�W芨m5�C�a􈭨�Ɯ0/0���F�C�Ijb���HT����y&���C����`�Γo�)ʳF�U��C�M;i�##�]}���Bj�P\B�	�]���l���Ȕ�R���&���.�ht�B�ą;��p�C�ɅȓO(�|k��R$6$d�(�- 
��?���'���?�R�J��	\,��ާ1.�B�[�-y�(ϖ#���ɀ!\��B�	=$l��f��G��3���x$&B�ɢ/E�1��D��d6�|��B�&�B�I�=��\؂���V��\�N;�C�I; ���e�ӄo�|��-2B�INO��C�ep�F�PA-��F{B䉑y��-��a�<}2��8G� B䉛w�@yBV铴(hȷ��
.�C䉹q 	�`V�+P� �b��l�C�::�P,�^2�l+w�Z��C�Iw��d����~� ��V�w$C�	�GӒ�s�+�Z'����Q�GW*-��:c���f�S(h�0��@Rp)��C���`�E�)3N�+�bG┄�S�? (�P���.����mO��P�`�"O$xS�/�X\�)�U=r#ؘ��"O>ڲjC�N6^���f�-�a�r"O�8��D�w��5P ŝ
iĩ�"O�0$�G3,�CAY9?N�+�"O��S7���h��*w ��6��CU����	P���q�m����)8�G�-.LC�ɍ>��<ɷN6�\4��L#<C䉨�*9�p�%�t!�dm��B3�C�� �@��G���*�/��xd24�"O�p��$�+��uL"-E�\p"O6��EH�!�4�;��W*����'��X�B��6t�r��4
ʸ]���B��OjB�	�p&DB��t��c'F�nvB䉆��e�&�#�;G^?Q`B䉱EҰ�y���'�p�f SR�B�	�I�y�D�m�����b�"B�	%6��+�4]pe�Wkؐ]DC�	T�@pR2*��<)���>i�C䉒w�"4�B89�3+u��=y�����|ub�l�gl �!h?}F�"O
��P��r�(���A/w��A"O��37�Q=.��p�@�!(�hp�t"O�iR+I�8|<�r��D�U��z�"O�L� ��WVD��v��W; 9""O�e��ĩc��H�7?Dl2"O�-�Go?"����>"V�c��'��'�D���nZ$t�!�j[�z��!�'4@�`Ś;�B��T$�2m!�X)�'��5�% \�O�$D8U1�'�n40�f���X�3��;0"���'B�<�`���Q�b\?*]�(�'ʖ��a
#�HIU&т�����'���
�.�h�lhi���T��'z�A1��sՠr���$��'����9](�8�Δ%�݉�'aP��B�Z=YF$ѵ$B�@dj�'0%Zj�:N�T��^ �@3�'�ıb�_<E0���B�� t�Ը�'��l�&��"b+2#�Dr� ���'�2�J�jڅ?��yY���Rr�<H��y"!� �"�I��D�;�(��t�yR+�vl%9鞕H���D�P��y�#CU"TX�᜹iv>�׭��y�lU����k�|���G��y��^�p��IU�H{�}P!c��yr-V:KϪ�a�!��!Bq ]���?��'�x|�t#�++zP4��j��6&ޠ��'���%Oڱ��Bd�τ�H�'=
��7C�`�{��݁�4H�'[Рj�̐�Z?L�ra@6�6��'�4��g��dQ��i��Z&m�@:�'�@�4L��6�)k�_��c�'c��!�JIԴl�ӥ��6�%a�'��t"�%O�G/��r�ǉ4���+�'{�"��,8� D
�**p4I
�'�j�Je�-T��ծ��pd1
�'oέ�i�!r���!Ł �2��	�'נ���-ح/�0�ϯ׊Q[	�'�P����:Z�D��@�A��':���%fF�e�	  ����'���+3 =�ꬲ&��`9���'��-�ǆL�^H��Ӹ	�0��"O��RN�YT\U��f����Y��"O� Z�C�jF��T�#�eS�s:9�Q"OR$�s ԰]T��DE�
��L�"O�%pe*C$Vx�8!g��d�F�P"O,@D'���2��{z^))"O�j��E.>]v@����Nsj���|B��!�'F� 	�#�%m�42�hѿn��Y�ȓ!����bKљ4ސ�1Ea :"���ȓq2ɂS�]
$]�4�E�W�^i�ȓDP��r��V?I���'σft(I��2���ɆU� ��g�� .!�DG{��O�b�b)f34@r�R&t��m��'�*	c1H�t�F��L�X�vU��'�\K���$ـX��%P�c�TL 
�'��)7͂�Q���+Y���	�'��X2c�!����P/B�RZ&��'��D�#P�����ȯRZ��'��d�Q�Ç� G���<����	�H�b=w�/��!'��!�$�7U���*�b*θ��pcZ� F�'��E����-��)��La���
��=)�LF0�yr%D�(x�����w3t���a�)�y��Z����#I��k�($�J���y�D��L0֜9��Ce���k�E�yr��0|xdbrb�]5z��Rǖ(�yr��#�ui"��M�$a�vb��yB��P���3/�K@�q&�[&�y���-Oa
 f�F�Hj|D��ґ�y2��0Px�[��G��ͳ0��*�y�#<J���b˘C$�y�ȉ#�y�(�5vQti8Q�Y6w��&Ɲ�y,֋/],5�gK�x�y����h`������"?\�흴8��ȓO#r��W���2����	���&���	�R���	� ?8ۧ�Ԓ[vC�ɺa��p%ß�d���M�&�fC�ɿ��¡�8
q�q��"lpC�ɞ|5�q�����DP#��,n&TC�I�>R�򤼙E��U��?i��iL1#ܦcFK�*M��0��]Y�!��,[��(���=9�#L��!�$c�$�c4hX�R-��*�*��!���RTRġ'_�|��g
��S!�dTs��H��'i�(lK.�!�$՗u�rD��A�Dr �	P�Y/!�d[t�,<���N�MP��FۜT>!�;Q��k �B&x5�����)P!�DʔtD�T8�Lϋ^+�kEc!��)�'"4�hzց�=iO�i���!�(��'(��0`��>�H��C#�Z�	�'����r'ɿ2�d���}�	�'ȩ*� �
"{��"[�p��X	�''�H:ÇԢQ���k�T�`H>���i�I������Y>Jx��&�\�!�V�AX�� 2d��=��('�-0��	^������C�q��֥�>!t�!�*D��3�CB'g��!�G�Q(`#T�C��4D�p��^$�@tY�OZ �6(��3D�ī�np���?UT&�Ju`&D� �Uk�=R��"g�6�L�D�)D�TR���%ˎ��H�~א�h�n5D�lf�N\(n)���I��N<�d D� ��i��龈��J�3[��r��>D���d��\)���J��=B�1D�DXQ��#_"��h���,E �%p"-1D�� �	�b�o�&Ib�aD6k��쳕"O�ᡥ�	\���*��"�8)k�"O�iz��G�r:���3�ҡN�.m��"OB�y��A�?��9����l��M��"O&�9)�+A����"o��u�"OƬ��K�JC)H!
9:e�'"O���,���8�$ϙ�L
-��"Oxh�Ƃ�{�F@ ��.>����"O��sP\(J��2�b�"VDt�@"Ob �%(?L�����09_�I9�"O�؛�K�HI�MОM��%"O����	?��lQ1���].�1��"OB;�LՔ��q������2"O*5�2aǿ'�zQ@ m��d�$p"O��#� �:5��ەK	1M�8�k�"O�9�Ā�	^��H�M(w �qr"OD5['F
�����V@o�%X�"O��[Q�}` gZ�H�3��E�<���>l�ũ/�0ew�@�<�����ʝ�f��<���`e�e�<��"ה5�^tQ' �)H<Q0d�X]�<y�G��E��y0���a(~�#aG�@�<9w�)"8�*����qC�)�a�<)�D�n_`�d!�9�]��`�<)G�.Yq�u�@��KȢ�6�_�<��n�.�����F�8*��"j�Y�<i��ܖ?��Iy�╺~8�2��H{�<9ddJ�k�ʙzGh۸4���"Yn�<��.�86����߳$���Yƌ�d�<9��U)mz�\	b��1q_��a��f�<)�G�te��I8��P�"k�`�'��Q�Oإy� Z0'4/�#{�ӊ�d9�%�4�6�T�V�i�,��,E� ��9��)���a22p�d�G��Ri�ȓs"
�zD��&��)b�o��S�*���^���y��H��t�q!N�+Hf|����4Ak4FW))�H�9��#b��m��o�����
���-��J� `�ny'��D{��Dք4�"0�U�5�ll��G��Py�lQ6n��U+�OY���6	V��y��͔!J����>J-x�چ�D��y��m�� r�Ŋ=$>�c��ٱ�yC@d
tQ"`�>�:�:d�֐�y2�Jw�0�R�f�/߀D�3�]��x�,f�p��&~N�8LM�ў�?͟\�T��*	����1dU/K�ʅ!G"O���e��'1=b�V��"t��kg"O��Â��**�X8��
T�n{B"O
���+�U�Ѡ�����"O֍Cu��)/,����I-G��z�"O��PIR hJ�je���/$�qB��d%�S�i�f��ݢ��Ël���H�@	0 �}�������R^档5�&�e`eL<D���� �0?�T踔l�+/��`�`�<D�|SR�  
�31��'R�8��b<D��9v�\l,h�'��7^�
5�4D�H��k�A�&QP)+���H�%D��p��LI� +�1r�fpm�#D�0H�G�1m�x�Ӌ�*r�,��/$D���g�5J�ʘ��͚�A�T�Ռ�Oʣ=E�L��w
v���%X�����E7P!��4=�ѕ��aA�@�+}�!�1N�<Y��끤�(9i�O՝N>!�$�H����	Ȓ�Y�/\�{�!�� �d��w���Zw�@"Y0u@2"O��H�JM,V������ 1���Zd"Oz��1k4�R���.�dl�"Oz��A卓<�B4���M�f;��6"O0A�N%M���ck�B#|PCe"O��YA%�`b)Wk�t8.�Ѳ"O��
A�Ym�����J3��8"O�<!��ª|)�����@!�c��n�<a/�(0y����N��	`�ny�'�dT L�6�LD��Aك!o�=�"O�y��b	I�hm�B!C�zz�5AB"O����F��w�����ϝ�C�1(�"O>u��pW�%�$��nd�P"O��"A�/
�@�9��6u�3�"O�I�p��9����$�N9D��(�"O�MS�D g�j���e�"�^\��"O�)�$�1��5�Ɵ�a&,�2"O:��wo��a�[F�S�ĨC�"O6%3���z�*�8�%�?J��U¦"Ot�� Ƌ����@f=�"Ot�#��Z�A�z��N^Y9�"O�8S��a�����'�(_W�Y��'nў"~��	J.���9�ݒ� �P�A@��y⅞0J�s�lV�y�N�s�L���'Taz���bL,X�'�љcg�dQ�� ��y�U& 6���� QY��,���y���}S@�
��дE�pH�g߷�y2�8����0D��$1��R��y2�W����)ȝi���熔��yB�\���(\�z����HX4�y��f!J "���qE�l11�ɡ�y)qR<y��@�l'J���ϑ�yB#	: G"l(U�J zWXYH�H���y2�V	7V����H�:�R�ϥ�y*��CӤn��GZTd�)��yR�����,�5@.h���̬�y2�S����b�L'a�ؕ�ea���y�Z�f��Z�%2k
H�%+��yb�@�l�:�"9O�4K�Hך�y�ʚ�;.H�R�D5�(����y��ؽ ��(�˕i}J��ᇅ=�y2g�/Ǫ;�HY*`c�$1A ���y��Mj�MBbiݱi%T�c �)��!�S�O�Y$�J�T� h��[� �B
�'YRm�������
D��0u2�'Ǹ�3�e�����L�C�9�	�'��у�.�3J�D}j���$�r�'��z�Ւ%�<|�O*����'���s�D�|�T�wIT+.�4|�'Z����'p�=p� M�;�D�
,O��=E�i_;N��1G��e���)$i�7�y�b���ื��̨�)�9��O�"~j�;tO�P�f�ރ+cP!�0��Q�<�bO�/꽋 ��&���X���L�<	���!XX�#����nf<U�'c�E�<! �X�B������ʑ>���#� L�<�U�.X�\B�З^*��(�H�<��ɇQVu�W��.�F��ȆC�<�&�Е?��xF�ZL���Z�<y��P��С���=jer ZB�<!��U	$�$�a�Ɛ���3e��W�<A�(½(���@��?�L���W�<yե�T�ư��-Ȓr{�th�Hy�<Cg-fZb��E�� I�a�<� J��R�ӄ@n���#�4� �#�"O��ƚXQ�����w�F8�"O8Ū���1*P!�m�7A�ưYR"OnA�"#`0PL�>"6Y"O��aH,4�h�qPK�.{4���"O���1�(k��IU��pm6�p�"O(	2kG�V�80����hNV�c�"O�3'9f6h9!Ţۯ;���I�"OF�w��x$��b�g˛PL����D.LO
���΄4~�PWƕZ��Ա�"O؀�Ӥñ)4�����J%��\Ic"O�h��ːaze���W(�Z���"O�����$40l�GbQ-�`���"OJx�uş�0Yf��B�+�t�EOf<Z���D����-A<Z*V�B�I� ��4��-̵t�$�R?-rB䉒n�t쑷	-S�����LB�	0h���ǉ1"X�X��߹d�B�	�D�(A��a�"�7iR{��B�
wGܰ�wE /�8X1�)�C�	�� �ag���4��Qv��&d�B�I�.$J$�J�4�B��RI�POd����II������C|�R6i�"[�C�	/�����O
���34LB�I�f6�<k�4�v�y�.>��d�鉤zE�)rW!y B�Z��q����ȓ<���wmG2� �"��N.^�e�� �^@
r)��y� �G �VS���	�p�ۗnH�za8*�K���%��T/V�p���s[�;��T��E���*e��d��\�QAja�ȓw�T��jL$AD��.�
>���'+a~��r�����ț2U�nm��N��yr@ Xha�W<Gֈ!P`��&�ybM� u��� T>�8��7���yR�� �"��E��!	�.DCv+A��y��R�0�,9�qÏ��*2w�B7�yba�Q���"�#DlX��&7��'�ў�O����ٗ6,u�@B�'\�J��	�'�z����Z}�QI`&RJ.%a	�'���`��ҵP0���F��J䬒	�'\BA��#���T�.s���	�'��di D�^�٩@�\o� qK	�'�L�dK;:�Ժ ǨJ�9*Op�����fa��A6iL>2�FH�z�!��#"�892����g�vكG�!��-S�0�豢�9���Zq�3!��I)���+݇Jv���W�٠8!�D�*-�`��G� Ǟ���d�#!�D"R�:�1�.׼G�]��C��U !�����cۋ]� �8�CY� �'�a|��+s UzpE-s��<�񪈡�yb�P���I��N�]��tc ھ�y�ɟ�/���Y=�q��o��y��)NB��C�`W�<�����2�yB�� /���8�=;��%�]���'�ў�O�bHɈ�JƝ;`پ�n5�	�'�R��
q�l��&�LZ�Y�'C�m�J�4F�tQ��y��k�'��M ��� [��������0X�'����@�;b����#�����'�x#��rnz��)��UJl�	�'�p����$������K0��ʓb�[��Q�[P��Re��;i���$���)� �H0�@�gz:i�Ì֓1�zm���	G�O�΅�B��?�@�`�ߚm��1��';�lH���W1Y���d�x����xb��/d�l����:H� KT�V+�y�F%	sdt����8�Dx G.�y�.>�b�*V��#.�p�Rь��y����z�lPHu� �Yj�#���hO�������y�@
�(Δ��E;�r�)�'sA��+ŭ�,�xYy�G����$r�'�p��c�٬/�������,jӴ"OJ�
6&>֦�qa�}���
`"OZx1FK�x�n�%@2�pY�"ORx��oF myʹ�O�K=���S�'T��#w]�]1��дKZ)!�rLBB>D�hSP)��B�����X%G�b�8G<��F��O�^��0�H��8�ܐf6�}Rϓ�OFt3�!�u�j�ض횞Pc�xS@"O�y#��C�,$-I �	�b-��bB"O*Q*W�R��$����
w ��"O�ͣ��@�G��|[�	Q�l�]!u"O\0����`��ԇ��)M�0H�"O|������Q} ���t;V���"O6��W��H^41C��1E�1�|r�)�ӻ"9|������lĈVnR�\'�B�� C$��ʤ���^�C��Ԭj�B�	�5����&z0�i��S�o�B�	�7�qqWjB>�@ ��ѝ >B�	7t�H����t\0�DF�3:'.B䉿+K^b�a�$�^M�ʛ�^��C�I�	䱓q��I�Vę~VC�Ɏ,�|PZB�b^`Cu[�#����0?�IPkZE+���<�|p�pe�i�<Y�y�jI�S%Yb�� �N�e�<g џ<:���4~��挞|�<��n�-O,t�j�Y�oբ���ʉ{����<���E ��G�G�F2vMNx�$Ex�J�)̸<�f�+��a���	�y�!�Y(�Sm�������M*�y�c
�RzZa�e�J��a��E�y�T�'b�u Gn� �b��R��yb��~��$@1@��p`�	�y�KZ�+ej�r�%M����c��W��y/B�z�DuyR� (~!��i׋�;���0>����?����̝�l`����^�<@��h)�I`a%Z�q���[`]�<1&i��D�%��^�@Z�Y+"�o�<��҃(�q��L��{�#�j�<�E�L�3<L���\(��I)��R�<��A�3B��� ��2r��P��QO�<��m�4�	���f<�HTÐHx��ExMˌt�y�[��|I���.�y2C�N
`dQ�mL�r�\	r�B �y��-.�~��&r~ި��b���yRɉ�1�f�[b�� ��!�d^��y���M��(8�.��~d��Pm��?����3�M��H��׳R�4{&���E
�\@
�']�<�t�ґ1ϴE��E�&<�����'n�@w$�)� 2,�#9�Z1��'�(��D"�+(J1�boB|4�2�'�k�ő�o��)bG&�(���'�|�����0id� �"��N����'~$�b�D��E�N��&�H�Nt����'�Qx�ECbZҌ��S�H0���'�`9p 
�w!B�2œ�<�Hd
��� ���Dͣh��]��E؍r��;7"On�	��Ɏf϶ҴE�=VFhKV"Of9�DAؐz��U�O)��k�"OL5��c��y�l��rK�2RX�A�"O����� �"W�aڡ)0%ޜ9zA"OV�.��2ξ��҉^
��-��"O��I􍚋n<�y5������V�P>��4j�JR�������!��i<�	��,G{�OAF�����o�t\t	^�B���'�8��C��q��8"s�	9R���'/����%��#�Ρ��n����'p�cȊ;�ș�����w-����'*��j�ɝ�Ax��{wA�ig<A��O ,s�J�G�^�6G$%'�A�|��)%u8�R�
�~U�� T��9m�B�L*��x�'�1;-j��P�ԥ_@�C�*J�8���:p+��u��:rJC�I�f����ö-\A%���6lzC�	�B����'�,�ҍ�4Q6�B�ɸLf�I��N������H�2�hB�	1}Z�dX��YJ�����WI��-�Ş���±:s���bS0S�$�y�b������<Q���̲)��=+$��Es�8��X?z!���lbmR�	ɫ%q����ąa�!�5`HR�R�e��">��+�r�!�$�D�
t�B�ڽj��������4�!��&3�� P"̷H��4�F�	��b>O��A�fψT��X1.�M]L�'"O.ʆ�F* 34�4�4H� 3"O��&��;�x�G���F;�a�"O���A�0B@0�Q�Ս�#L&D��
�B.�zm�&,�[hě�&D��s� �����H@
�T�yB�$D��;�׎k��mˣ )u���#D���/ُq*p��C'
�F��BB�<D���̔$ q����Z�8=��Vh:D�;�bӄ)R�����M3lz��0�7D�c_X�2��ܿT��`���k��C�I�	 ��P�չ-!�M�`ǀ9(�zC�I�Q<kbF��G�0t@�-�L:�O ��$�>	
}��D:� �c�?o�!�Dȝh����T�O�Js#N�!!�ĝ2^�l�c�'��_�D)3ł�	y=!�dӍ^J��ҲGǲz�2l���3J6!��}W�e*�[xSvZ-!��Mkh�����nY�<��䀿X!���^�N�鴍T�2^b�re$�!��K���i�N©Wv*pIN�x�!�D%;$d�����H�1Zdi��b�b�)�'��aљ+��E`q�N�v� 
�'��U��$/�,`��I+L�-D���G��4Y�jP���;��	�g.D��*de��K�Rp
��Z	B��T0�,D����C	X������V$fz� ��*D�l�5k\�MGz�+#��>.�����;D��xf�]�l����C`��e�D
�;�$%�Sܧp�|2�Ծ.� ���n���_y�="�lE���T!�A��*����%���+�f+C����bJ�px���ȓ�6L��ɇǩ/�xXi[W�<���?(�(�"�I/pc`-A�a�{�<�vC��Ztb�f��XoF���b�u�<��
��me�W5{0�$J�oq�<yu통l��ģ&o�7[[�PӦ��C�<�  a��N�R����%l�+�&`Pa"O����#\�t� �ō�,�$I�f"O�&ɜ�<�ZTj��)[�ԙ��"O.�`��߲W�pª�3x�"O��;��L�r�b��U�k�B�J�"O\p��9�\�V
U�a@,��"O��2��X�I"0l�8�"O╛���!��/���ظ"OP@�*V#"pL�V��l��"O��N_	��� ��Z�D�D"O���SN�?I/B@��@�_�(�3"O��a�a�� �_,h�>��d"O�iBCW�\U��"���=��	�d"O� (Am� �@Mj��KtZ�+'"Of� �������P"�ߣ(bjc"O��c�LԬc��}�1l΍��<�Q"Ob�س�E*r`ZuA��؋C��0�"O0�Xa��08�d�2%�;r�p�XG"ObوP�Zp�P����	�$��"O�5�$@q�H��ƀ��!B�"O�ж 	-:d�a ��������"O�=k���: Wf ����"tt$X6"Od,0֯J8�ԍ�#DUU���p"O4Xx$�Jw����M�@��q""O��B�8N��=�mF�M�D%rQ"O�����^	�o$+���`�"O�!��˪�%��XG` 2�"O	%.ˊtt�8MK�+;̼k$"O��ܜh��22a�e�5��"O4�;q��c٢HaiϲM,��P#"O\4�!��3���r�@3u�.|�"O�M�kL!\\Z#�P�X�>H��"O�����+Aڤb�/�O�.AQ�"O�<�2HV�9ĉ�'��/2�(�f"O6B����&��eK՛>�`�ׁ0D���p)�:X����P	�%��$B� D�H��煬1��t��.��p	�03��*D����
�T��٠��K���d��N%D��qRV1�d@��芿eH�P�b D�p��U��)�QG
3FH�=D�����7H�h��0��0�Hp��<D�Xa�`�GI��cBJ�@{��=D�@ԏ̱��Đw��>�Ia
/D��C1 јT<��gA�æ� �!D�Dڦ�O08��j�,A?�f��C�,D�d� ��}�Вe���B����(D�h��"ݑ=X`$���V�n�6�"D�L���$A��RڇD7��b�i D��KD�T9"SDV`���ӬN-V�!��3r�C�g�R4�ǥ�~�!��5K�$5�ٙ7�D�T���Q�!�L�O�����n��fd
�u�!�DO?:��U��K�!�B��t�!�$V���k@��+ .�cR,�5�!��(<��C�-�	���V:P�!�ĉ<$�T�%�G�h~����R��!�dFe NѲU��␙����o�!�W8U,b�JJa���ڶɊ�!�$EGS�p*&��;c��Q�	�3=�!�DO/C� �b%��)T����Q�J�!�����c'�O�d�,)�U��!��	�L����D�w��,�C�Z!��P�fA�e�X&Pl"��dO:�!�$��)��MA�5󰯒#?!�� ��ɠ�@�F�:��Q?�d8� "O�}r4��	�x���A΂r@�"O1J�MU�uļY��p��5"O\���~S���I5���K3"OJY�$��!&ItD�dɖD�ґ��"O���&E�}W�qS�׮w�^	8"O�L�ìɱ>�� z��S9%e~��"O&)*�iOk��H��F�)�m�R�"O�@��ܾl8��b"@�p�x)d"Ov\{��Q����#��]���"O,����8A�N\��Pp&"O���!��#fN죴��!�F�s"OF�z@��n~spFJ�VN!�6"O�K:����M��.Ҙ+�#Z�$�!���%���Z�c�RVirA�S�!���X��뤊
�7Q��q�`ȍD!�ͦ!|.�ySm�2-V���AZ�|�!��/	� �C$6�����U'�!�$O'�f�"s�0V���psoܻr�!�� |ƑkA/��A���n��f�!�D��P{X� �[�E|���6C�%�!�dH�0z�E�d�Ƨ)u��1�ǍYx!�č�pF2�X��?]�q&쎅_X!�ͭc`Z���IH�'@�ͱ�5W!��&���q�)	�q=���g�G�!�D �P��Ö��b�Jpp��*M�!�K�LJ@�"E]�:|���#��K�!��) 5�p"#�	b�t�1M� !�$��.�a�*��bn���V�ùg�!�$�;g�&	+A+��GO@�w	��!�.�PDcDD%E:tR�\�%�!�L�֩���J������-�!��H�8Azh����Q�(�	�V�!�DC-~�x��t��.�<���Y�_�!�DD64���'X>��8`	�!��@�b`dP�-��q����!�B:U�!�Dџ5�´���O�B4�L�!���:N��4�ؖ3E���ˀ�Y�!�Ä+;!
�
��1!>��CO�	�!��2jA��V
ӶZ(���g�?5�!��^7@��EJ�,Et��6l@�!�M�PRր���@lrF�[%j�.m�!��%a�N�`&L��N�X��"��o�!���\z,�#�:��-�O�'�!�ĕ=W���D�*U��͂�'g�!�C�9���P��#z �Y�iC�K�!�DƳ�|49�F�>�6%C2g�*"�!��,��ly4GՐ �(��g��Q�!�DY�*�A�Y�q��d��1B�p��7���#E�K'�y��=D���ȓa0�%�J@�&[���2`^��� ��T0�p��Cݩz�D9���26������ 4჏�}��rg���|,����_!��(���$�q%���!�L��ȓ�:1PV$� ��1����B���7� �� ,��S�D�?f�D����#Kde���G)�&��%�ȓG���)��+��m�,[*v>m�ȓ&}l�rŃ�1����GQ;Rx!�ȓy��-h"-�UT�0�b�K�P� ���
����1$7y�L�	!h��$)�ȓ=�0�BG(#A��ͱ��W�m����P��qO�@@.4�TED91>���ȓn��<�R��)�>�i��:��Ѕ�S�? h�(b-
LNt�C�FҰl^Ԩ�"O���1"��'�֍.h���$"O��*PATA�(�HA�	{ >��"OF�ç#RU�X�ȏ�8z9�W"O<��4
���4K�߷M�� �S"O�u�R`5$��EQ��t8�1�"O�`۠E� g���WLpl�X��"O�����-M�uy��z\"�ʱ"OvQ��(̰{cX��
"LM�-�e"OD����L:>j��֪y��(�"O��a"(�!��5�e
��YP@J�"Ox$���2���XON<#v���"O���S� �o�|�7̆l�xiq�"O�����e���"T;мA�P"OP�
��Ӟ`%�1�4ؙ�����"O�|�s�D�#R�l��b��kBr��'"O�d�>��$��22��	V"OXu��^�
��60
�}�W"O�ܛ�ʇ6fF$��F��C�Y87"OBa�t_4f]8��H���BT��"O�;B@��	T"�P�8jЁ�5"O��� z씐���6kc�u5"O�ɔ��:b��%ʧ���@:���"OD4�l����p֎и L���0"O6yAA)P����O��r?�A "O���(�2"��3��� <F9��"O�4a@�9"^@ܒ��מ��&"O䘉��N�m�����E�'�DXS"O4�`�M�->�z��\�W��L��"Of\SCF��-�]� ���D"O ,H7�ޝ���)�S����P"O*���T7Ow� �h��\ P"O�tp��%T�� Ug�+>�a"O�jQ�+(A�l���
o6q�"O�hX�FE��
���%
}a|$y"O��:�S�WENĚw�MmEj�"O�8��0@�ⱻ��r��a"OK��
�cS$V�`��"�yr�~�TԪT��:�-!5���y�i� ���ⴎ[�ԐS� ��O`���τ%�#P��.U�������R!��Ѭ�To���������!�D�f�֬���Y��p�T�T�v	Q�,F�D�L����� zR�0𱂖&�y���5
�����n4x���q�����~�)ڧ�и#�Y�;
<Q"��
3��ɇ�	`����B��X�X�Q��-F��ȓ\��y�T���%v��U���a�l��=A�O~�~�� L:M��83�!�3��CV)�K�<��$Z�>�tT[Q�S/J`Z�Ѭ�J�'��?������6��.�"P�W�$D�l� �=2���GФyFبt�u�D�����sӐ��R@��1��,c'��|i�Z�"O�[J	�j���c�w��j�"OL���hZ>0�4�8$���5f`�Q�"Oh�U��MkޝP-	8_P�:"O\� 2O"
�rZ�JI%�>���~��� 
�I���ZGHT��}5n/D��c���Gc8!��ܾۄ�kR!/D��s!�'FHh�eO�~VLM�E*D��3��[\����`M�ZR>U�D*D������mL�)F�Z�����4D�l�S�� 0�T9
F��)Z�M�O�B��/5�0�cp�����+rDN)�4C�)� � �NS�SB�	�!X��"O��;ֈ�2��	v��_�9�`"O��bvL���0$aag����|8�"Oz@sV�B'/r��XƦZ%q�<hk�"O�Ś&˗f��\!'&��t�v5`�"O�e��%L(S�(Uz�@�=���"O���R K��Z��Ǣ���"OE�%��ݸ�/,<��i:r"O 12g "�cm �j�z��"O@�qvF�!Y�z�	 �L�_H��3"O�P�ƜiSU�g
��Hc^I�c"OH�)ff�?,���7O�\�eO����V�`�Pl/.����jN�<��i�v5���0	�'h"�{G��M�<Y�*ÂT���C͓�i�<�4a�<���+���[�LЪY�t*�`�<i�L��j��=�N[ pC2GZ�<iǅM�&��(��l�01B&�a$�~�<�#@}#uC�g���|�<1��_"���r�ǈ%´���c�u�<�%�
b�Je�%H�[�j�c��o�<1�זc.��aaGo�U��l�<��Ώ;�0A
���:]� M;��^�<��N�7)�$�E �5P��5�#˝n�<Q&
��d� �˖���y�0n�b�<�F�	S��	��(<��S��i�<�P%�p��@���$!ƛg�<1���8�b1�� *_�A��	Ae�<a5���Hr�:�n�R��g�Ed�<�d�8h!�Yآ�I���yt��M}r�d/�g?�M�`yY��_/j���C��Z��X�'��$x� �+�m��釞v�n��'��'��keE�=�B'	vb@�D}��s�
��)��`S@&[@Ƭ�bgI]�B�B�I,3�jĸ�@U+7j0m@��UR��	T������+5��So4� ��� ^��Ĺ�"O��#�5@Z�����7��͙UP����}:Hً��]�<6H;ǪƟ �
B��3pS@@�&]�!1(4��A.)ߐB�	�Z��ӓ� �>�h�.M��B�I$�U�1c�w(�"b���V�FB�I$
B�5�v̜�*g��Ie��Zm@ʓ\��|��*³?' �����	��H@G���=9SD
9l#0)KE�DO5HE+GfF?��O���퉏%���Wj
3��ɪ�K��Y�nC��2w�@C@Y+pX⥺5l�
	�B��#~v�B������d 27����d4ړu��=��aܱ*̨d�� �,7M��8�H�����+�g��<=L�'V@IFy��i۞MC��[��N4��Xk�ɓ�M�V�>�ߓHh�a���� ���c�*��ȓ,���!r�Sfn�P#! 'W͆����M�E./1�b�pfLv�P��&c�J̓�?1��������>Dk��ÿ������y��_"
��e���o��H�P�Y��yr���<'��ӷ�_$^;05�c�+�yr�ͨJ3d�b�A7YM���mצ��'a{"�e7,�{�A�:Bh��a�%�ybk��.��!�q� '̦d`���y���B/I;O�l��%�mn��'$h� �{���aڇfyh��'E�щ���9J;*��G,��W�b�'��ܲ�@��9=��
A��xe�
�'�DQ�G�ɘ�J��&K��Pvk�y���� �RS�._@P	 ��<i�Bf�'�qOV�C��Ҟ��p�窇�~���r"O2,Z�om�,YHo+f���B��	mx�����l rQ�e#9�Q0�, �O��K�� ����/�
5h�_�lL�����q���01ؕJ3œ�~�D}��S,����A�ʐfL"y0t�)�XB�I�#PUEdˠ.}�<��߃�F����0��O�1���(��ds�kP����G"O`��b��B��p�uEO�jɬ`�6�X?�������Ş��9O>%Re'9�eygd_�SO>i"O�]�梜�S:��)�2j�R�Iw"O�� �B���Q�pg�p����"O,ͳ��Z5&�`���8[��$�'!�dG>1 �Z�J�w]�1�`/�B	1O2"=Y����P*pPsI�2�$����O��y��Ъe�8<��(S�ݡ���O����˵�Tu��O
DG�X�S�² ;!��G�`E.p�� �7K�H��S��䓄p>!ҏ-r�@�z���H�"v�Bn�'�O �O��}qRd�	IxBؒV	^IfhP�'S��pY�H�ī��ʓ%hT����#�S�D�V2�z/�_\��&)�y�˂pk<��2\i�+�9���~��):s��s;���W��r�
�p��GS؟��I�z����
M�諡�X=\3�	��n��<K���xv��"`W�G�4��Vb�� G鑇 ��a��B�h�J1�ȓ;��0�LւA�2��G�lĬ�O��=�r�.�^hԅ�6(�A���|�<aE)�0�P<�uȉ�?uP�ku� ~��O ���]|��ʔ�0��Q�$.�rta{���O��j�zd��nh�9)Ul(rl!�d�0�<8��Q.K���8��J�j�!��H�&H$�f�ߗu��܊�H�;'�!�D��rf�a9ҠEZ�:� u"��!�$ͻ-V�i
�!�%6q�@uo�!������ԪYb��:K
9�!�\>s°5c���Z�pm�@c	��!��5k#�z�ЈM�2}�)\|!�$��Z��C*U��!(���Rn!���-XCH$
T��5��@�(ө !�DǶ&�+�f�f��T0���l!�R�-fT��6�:j��1��	O!�[�V��4�4��7K�ֽ�%�J?h:!��W�'�����)��v0��N�)ǡ��;T���x���@{�\J�i��y2I�F%���D�6^d�2�ꊣ�y"`�	[�ڭj�,2�n�'�"�y��w,���@\�^P�v$]�y��O-�@���F�f��ƈ��y�O�()X܍�w��B/2��j��yR,�&wX�Q#� �I㠝*S/�"�yR&�?"Xv�r��B��T�Wf��y�<�<� ��>^@Ec7���y�/�c�|�@7C��t�m!���y/Ͱ�� ��L��^�r���y��=#�`�!!��!)�0�y2`̑%a��k0[q�v���y�'��y�@�1����X1�)�PC���y�H"@u��&��>��UQp����y"�
$�bQYv��֝B`�[%�y�NM�#N�����}��8��N�y���-՞���I;ntj�Y���y
� Υ[Q�3`bUk�K_�B�%�"OV Yr��({��@{�V K�����"OF1觤\!:�P��j����D��"O\ȇB�*��Q�ňm��k��'x�		� ��J]��"����CFI"|E���	�'g��L�!Ϣ��&�#/�.�	�'V���/]: �
��%F�C�'}��u�\�2M`X�5�؛��xs�'��E��dϤXqR��P�؏,�����'��u�M^'[ar��
�H<8�{�'��q!`[#k��(��U0�$q�	�'*����$�YO��k!%ү6��)+	�'1Nh����&z0ĺ@��\��A	�'\F�V {���s�.�]�j���'�1��F�]v6H�W��]0�\��'�bl#�LE>c� )�� V��0�'"�� H̾A����!��J���+�'Gp̙�k�:DA$Pc��K�L��YC�'W.Q�1�S+hL<p��Õ1�T�q�'��p��N+Dw����(��^��'?��@*�|P����'m��%��'��Ĺ�/uS`,���X�|Q��'���Č	3fM H;���W��%B�'� 0�s霊���A!#۽Md�̺
�'Hx8Rwg��]Q�	ӊ]�r�Ԡ
�'�ZԈ�݃ \�RcNNu��J	�'��r'��<h��LAjF�0=�x��'�(Z��R/�Z�x�P2.�L ��'J �1�	H5������S�( �Y�'TZ,��I��'�DP���h���'�J�1�e���P!�G�C�R�<[�'��j ��>��J�k�%~(�H�'О �bʣW������&v���X�'\� �Ƅ��<(2�ߢ�`xx
�'�츙G�N�]��"�ݝL����'j���'��-i����O�q_�0*�'Ɗ̢�oy4�!�R�t]�
�'d�D;����<>�s1��:u���H�'O8�S��H�`�A��nQ���'�z��b+�g����h�cTP�
�'y� �@Qkܠ6.��g*����"Ojx��Ɉ/d����q�ͦr��X�"O��gM+s&$��X0ت�E"O��Q��LС�+�y�~��A"O�#E��5p8�!C�N��(d3�"OP3��>,v��4H�`�X�+V"O���$�ѣL���4�
	rd��w"O�ɷ�J�<���K4 P`��R`"O!���9VӅ�MHF�0��"O$����M�X�R�;=;$8"Oz�:��e�xIf�@6�¤"OF�I��<J��D��+{ltHq"Obhѵ��[ܩ�£�/[X$��""O (���9SbժFvX�Kp��J!��6L+�L����/m\��bA�{?!�d�)<F���c���E$Ըpg��&�!��£U윪Պ�	�b1E��#�!��	�	�*!r�c�0zA��f�$!�D'Z\�er�)V'�
����	
!�$Â�*U�&o(
��$���[tm!�ė�bnȲDk�>t��ѐ��P[!�D\9��U��k�2 a.�Q�ã0�!�D�r�����M�3r�X˰�D�!�d��yL���)�0!&p��ԬX�!�� �<�� � +���V5A�$s&"O|tP�*:%r��Q��&	+�"O2����.7�� �)B�)�pT�D"O�!�L��O?�� ��(L�x�"O�uCあ@���^�j}�i�"O���%�\�:���� �\�i�$MC�"O�-�g��|��:��L�N�4p��"O�`աQ�1���h4����d��"Oh���j��t�$$끉Q"�"0�"O�0xÄ�S��8p��Q�n����"O"|��O 2A+�ؙ0�'.���"Of@@��!��m��eʞ|M
1"O[�bʒr����˟%��"O����酹l�e:j��IH��5"O�  )��x��h*�v>&4 �"O*��T	��@-`���)�/}4!�C"OA`FN+����G�:�LQr"O$��$ �r�$}��/[4�f�W"O���Wύ�/~�
g��5N^��V"O޼��	� m�lx�
�R�!�"O.!1ģְ�"�BU�\(�Ty�""O�m�a��@�l@�ūR���u"O 1c
��)�|��>��\��"O�9�2�^�r����Օg�&��r"O��H��D�GF��+��J`����
Op�h�
Z������j�Q�s��	��a��'T�-b�ޑ>ܐqs��0đ�c^"w�����S;I�������g�v,�Q���=�ÂҾ��p[�'�h�;5����bs�ۆq���شw�@Bげ9Ch�h� .џ#�$R��	�}�D/\�9�~�Щ�>�#"  C��p:�dO�,Ą�0OĔ��%��!m����C�`,IxSɌ9^Z��DA;<4�pQf�5��3F͜���W�Xd�Y 6%\wpF��=�Rn�9=��Z��'�ӻ9��!Z��w�1��%�? 1,��b@%o��<Cg_�{X$����7�|����m���JEHز?rTS@�H�	8�'},��V���;X M�<Z� K�ǂϼ�nR/u&A�(��*V!�v�K�<����	4���2)˪s��ej�j��?��_�&���jGh]$e��H�,1���SB�Kj��E�Xi@6�$ebx�h MH�x��	�\#ps�Eӿ󄈇
C�
�B8���#D� �d�`d� A�,���_:G� aP?F���ߘ'Ēx��iN=iL(�����nTr�{�F�6>�`�D�d��oL2�lHN[ $�B���pe����+#d϶�p���.>�"�O}��!R��'��a���!#���S�m5Sz$�ipH߇Y�:J�L����C��Qr�-�6ʏ%2�����{L��Ӱ�I׬�JeJZ�[	����-�qg�7V��0������l��⦥P �K��$H(�bV/�5��	�u���T,	
�*��@TG�XD�'��E*����Ŕ~���Q�OH�ID��'|�ѐ!��L����GA�L#��ƛlݨ��ٮi;��:�t�0�&��W�h�ԋɀbu��"���-a}RbS�B]2��Q�X<~8j�iD�~Gx8���2k$tšc�ơr�L ��F08:�=��_?�%�����<�f�/6��Ez�@O/�PA��C`�ufW�~�Ț�Ap���Q��d��T�tL�.X�Ā�'N~y��*�02��Ł�N�q���h�}�J�#��H��\�dJrY�gj�21���>�k�F�V4a�4lÔH�CPLOj�<�%�[|b3��L68m���/{WH���g�2Dq�X�4�Ҥ+�fɖO��Q�SL�	c:�,ҕ�K=��ݰA�^�>3N�����2 �F�9q�*��dFH�S&/�Y���kwAM!B���dE;`�(p��9:cz�R$eN�)y@,B`.\��#>9g�/]���I���@ƍce�"ux���&L�aM2�Q�AшL�:]{�GW�Mj!�d��Ĭ���?!x��1�#�^��7=�!�Ӆy���ZgܜdQÃ?��$E~	ca(�'/��1��ŠJ�@C�eOA%�،h!Ca�C�PL�y�d�RԄ�� `�3&d�%4��V���{T+��,*TD����Tw0H��	$}|��<�Pq��,l3�肈/;^X�3O	E"��@B���<�-\�u?\ⶬ�<`�V�� Fb�Dٕx¤�+O0��� �6fS�	��JL�2�Ѱv���l�T���Č3�my�OJo�!��'��$�K�ls"@��Q�'�D�s_�ș4�يD��:uO�<<�V(�R�۝�u�Q%��6�� �p���QX���E��*Ǽ��V�'t�dⱣ>,<�҈^=�x�,�~��!S1.���3��V��u���'8	�O�'�`ȩE��	��mلj
�_�f}{���� /�
7����'7]��9�]yN��K���s��-�'w�%���Dv��͆�I�̃)\�.��T��āE�˓ql��ړ-ך���`%�	��a+`��`�M��F�xH桱�o�	�T+O����+V�X�l���FB���D(1
�j-��'o.���H�����qkא\�d��OH�]��@L����^��y�#Hj&��$+�X�BBJ��hs*���&�z�`p�C)�,"�xH�&�~l�٢O��`����Ԡ'?��6m��p��y�#FݺD����rKc�'X�}BF�q�}ӣcJ,��ĨNr�(�p@G~6 ��q�uj�Ɏ�f��Fhx�`��C�)�ᑧF�M�bYiJ�<I����8���%+'R�逍��N-�z�"WJ�<y���I��&�D-���V�<)�V"W��z��7��ұ˔3H��*D�ԕ�y�ԓ�F-����y"&ۼefl��"�l���C*	 �Px�-^2S��a:R�P�
i*.ڜo��"��ݧ&�u@�	f���PA�
h���*�K�k C+\Ob��d�C�9����'�����'NbA�i��2+���A	�'�6�"gd�e��(��� A�,c�{bЍ#o�-��Ty?)��ӊ�f�'	��:a
�	�x���*=�d��`tXы��еk)�9pL�W�0�"'U�
��I�b��*��Wp�O�x�d�Fɋ���gqf�#d�`HC�	k��h����z� ��X>A�l����Zx��'���8"�OM0�Dz�!
>��}hw
T#o�Rq�����x�'X�%rRdcU�����桃�9U�m�g�4R�XA��I�j(*DF���\i*q �/Fx���#�DYJ���
����|h0���� M4��b�h[�D!�+Q�t�d��s8�a��Y�U��':�}��	X�P砱F��h�{�^���%�)��E���y����z�Q�`m�'lzQ�#O&@`���;}�
C���R�)IQ�'?T�س2'��1�����$B�P�sDٟ2�tb'� i�l�ed�9M��So!�O�l�T!
j��	B��\��e� �'��rfcK_��a�'��	*P��q��[1,\�Zt����'ؠ\S��?E bVKP#G�r骋yBP�E�x�����~�N�r��?{yja����B�!i��|��n��N�Z���V�N���,�I�I�Q>�*���%!�WU����Η�~Y�� ����SV'lzp(
�
t��c6� 3����dRtٳ��ʳck�-��*���5FE�HG^qC�	�Ʌ�q#r��%�7�!珗�h4��u���F+N������1/�l��1�L}(��	��J&'��	��9�ȓO���s�*p�25䋄x�t�ȓz=���6-9"�h�U�י]��ȓ{�$�2�B�;�)��S ��`�ȓ0t�8��,$��)�m�'^D �ȓmt{�B��ȂY~�H!B�ծ=6!�����S,�L�#F�<O!�$ѓn���[w��o���7
#!�D�I��y�7�"��1pD�!�!�d �f��!{�����#D:�!�	
�26��'x�(�@���!�d�C��t�R"�.K(�I���&A!�
	t�S�!�;MҪ@��@�H�!�� s{ryq+�,��@�o�!��p�B�@��ʘ}��L���!�d�v�B@*�
��*�\L��M��q�!�D��Y'01��W�q�����N�n�!�DX9bd�SoR#T�()�3'�!�$Jr:���Y�"���c���$.	!�d��m�Lm�.���hq#�8!�dJ5+�ar��z�EҴ�U�!�� �����C�!*�\Z �݌&�H�3"O���M�<9�Џ�4t2$3"O �iV���4X��F�	[�"OY�t-� �N� ���.�""ODM�3��0�p�!�N��cN�ʤ"O�x[�����!Ұ�ܴ\��u)�"Ozy8���b�s熓;V�n�!�"O����G�JF*���B�=�
�#"O�IsE��d ���g��u)@"O\嘧+��na����]�A8��S"O�y�3�E�\�zAEH�E�ԉ3W"O��`AϲP)@E��B�����"O6pS�Kr� $���2'ꎑy"O0Ź�f�� �����++���3%"Of9c�3_�&(�u�6�H,��"O=��:�qp�gI��h�"O\�p��X�txjm��B:d�xRG"OL`($���o"dHjj	�wP���"O"a8��.].�E��
?��xP"Ob��e�G�v�ы�;"O�Jf"P1=�&hR��S�Gm���"O��p�C�0�T�!�_f��P"O8m@1�W��q���ɴE^����"O����,@I����J�����H"O��ɁhR.F��@��A�6���"O��� ��v[`	�'��i��@��"Oq�'�0?DR�oT/<�Z�5"OJ$0��T!zZZᒷ-�?`2�53$"O��K���?]nX��Ѩ.Ȩ1�"O"1p�:Y���C!ٕU(T	��"OBa�j�m��4�Wk�L+Դ�r"O�X2w�΅JbՓ�-�a2)�"O��[`�	Dh�j��D ��"OzX�㪆�O��p���ݳ&��	��"O �G�߀X'��Y��%q�py�"Or��2�Ғq�:0����yt��ې"O���D'�*"8�
PG�\��Ĉ�"O�xb�dˀ3�]�H�-pRܐb"OB=��OO�*r�BE�_{�H�S"O@�SO�pւ	�E�*{l�Xg"O��P&W+U�()C��ƌ'X)f"O�I��-��(;�"Z3�0Ik"O�=@'�Z��v�t�% D��"O6$�fmP9N�}�N�/��"O�%��	o l��n�N�Z�*4"Ol2����9O4�q�M�{�RPS�"O��:�ő(M�� C�%�*mz�"O����әo`���,S/{�bEpw"O|���W�&FpJ�!]�3����"O���jS�v��00�c��Ѝ��"OZ)����>�4�A���"�9�"O�,�aH�d�0\��Bu�xh�Q"O���&I�o$QIplskr<���"O�i��!�����,	))S`�X�"O�48�g[35����@��j�ei�"O�4�񉈛B�|��G-N$Z��Z�"OVU��^�E��M
b-F���K"O�|:Q�P�$ �*%�Z'N?��P5"O�HH�9�`HV��))�yq"O���G�Y�e����G�CQ��"O�)p'펕$\�	 �K�)��Ma�"O@`Il�"
�"�R7�� �mq5"ObĲ����R1"^�$�@�pc"O�ؐ+�<@'4A�`��m���"�"O� ��B�kό��3��=|�H;�"O�@�	�J�t�ac��y�V}�C"O�9���>+����M�xf�"Oj�!��V�y�X�!�A/ OJ5ے"O��É�D�q0�G@I�]�W"O\t ,�4 !(jBJ�H%q�"O�Q���0�����&)�J\Ȣ"O<(��㘣w���%���<��"O"��&U�p���Wya�"O�k�AX�w����lD*����"O�$�@M�\A���삙ɼ�1�"O��Q���0m�m������&�G�<!tbў#&��'���H����H�<1�K@�2*���J�?�ܛ#�F�<��I�!;�1y��
0&��"NJ�<y��5"h���S�Gt����ΑA�<���E�P!��:��0��G�<����8�tȳ��ѱP�Q��[�<�2��"x���p��1�Ж�N�<������z���-����H�D�<!��?hU�B���J�9��	I�<��A%�����f�	��m�<	&�% f��	ug��j�`��h�<	��X�\ ������5?��P�l e�<9aR�_�ryb5χ,x�j��\�<ѳ��<��*rF�L�	�X�<17��/l�h*s�ڠ[:�X����U�<���X�(]*%`�%_CnI�Ս�S�<9AdV('�č��M'+�H�ʊv�<	�')
h R/����Jw�@U�<��ʜ=D�Hae�����kΚ8���S��D-�g?��e#��,�΁�jL0�k�[�<��댕/ٴ�r���_^0͢ӡ�ꦙ���ۗP�}���-r�T��(�g���*픸i|����>+�]E�Z��yR(]�/��MjBc�!<5h�C���*�yRƜ�S�����(�"��$����'�pRき�6�l�F���J�I���a�aٶ[�z���>�y��PN��Tc�̍J��\�D M�F�u��k4���Z�Q>�2J Hw�|��y:����>\مȓ,Ʋ~zf$��%%Wؼ�eBO�,ĸ�"g�GHZ(��I�;c��g��5A��`3&Ei����� 6Ҕy��Z>�y��ܙk :t���Fg������~hP�JG`0�=E�T�6����1LK
$VL��5i���'�t�ڔ �n:��D���ސ%k��Sբާ$��BU�����ŽML�=���*<O�� �[�K������̕6�^�pBb�qɼQ�d�>�$$��V%����Cܲ=��Jǆ �.^ k�.�d��P��OH�RΜ$[%��� [�Exp�CǱiBΉ�4D����P���C�i�ɺ�O�	��)�ҙ#���:t^�����-Ea�{¡��{m���'�T�3�gϞ=�C��*[*Xu��n�:"|��9��2����������	+��@��n��֠�`ӌ��P��C�	11e��(2��W�!
b	J�@�1�O ��!Ş�&��i�4N4,O8]�+bqh��R �x���p<� H�~$`t�E�g�Aڰ��i����e���yq1���%3Ԏ���'�l8d�إ%�&0��fՏ#z�q�O�E@"�L�'V�����	��0��DXD�']�& ��jK�hL|�Ǎ�Ek@��Pԁ��}�.Aχ79O�@S����c�:q���pd�3�
w�Ӑ�'��<S�j^�N�|��)��a����]���F�
<,c3b����4�pƃ>;f����!�37&X@(P�ˡ
b8��:7+EA�U��Hc�ʇ@џ�pdQ�6�{R�(5�C��E�
aZ��P���:ed_�>-Mp�O*��w"��Lj�L�d�Gj�����R���Cɓ�=��;c�N�H<���!�;���<E�%�X�)7бɔ��"OB���Q|�`JU����\�D�D�0J��!�GͧW@iK@��&O��ODm'�X�`څ^2ը�$�Z�;�#�O8H��A;� l����]0��d(@)�8�<�Җ�כ��	3�Ɇ ��y���3<O���Čfr�5���>~�8�>a�ɇ�|�(�&d�(�#N���� `GZ|A��:WH +T!� �Ȍ�P�-�B�	�i����,13�]#0 �Cc:�'5�ܸ7m� ������(4��	{l�Y3p�A��}�;r:�����'t�D+�b�:<izɇ��<s?���F�@9xP�i�*��K�p����k����Gԝp�VT��J��	j�	8y�k�	''����+�;���8&K!n��?c/íyA�d�8�I�"��4����}�L�i�ŃGx剈HY�YK�@�ayB휦);����o�ʕIӏ
���ˢf�QJ��>+JY3����!����D�2L�0Q�'X^�S$�ˠI �� ����E!/"�(��(u\X )2K��\���
 �ر*�D"����� - 铧y�`��dN`J1BD�}-ށ�4����?a��A�b�H��T��ma�� �%]Ͳ͚	�)J�}�6�'iR�'�`�Ѝ@ M��O��0x�ҹ8iT��6�З�^���	J����[�FUVp:U���|^x�)Rb�{���rƠS��r�'�i˵,A�S0�y�-F�^��5s���Jz�Ce�Ǚ����hl&U�1�k�Y��7�S�2ü͸�K��
64�� CB�szu� b�t\!��)-�Q׫�\h}rQ�֏A����w��P'``�0����R�S'~L��Ҡr3�	)���Z��G�����]�a��9� 3	:��`�2��%��FM��0>A�e�4t^)cP�.-��ihdP����K
�h
�#4O2�bT��3�<��w�}
����"O��C(Ԋ|�����(_1A�����?"T��3� ��~Z}����?E*���>�9P�[����@�,D��3�"��� ��z�̩2g�?9
<Ґ�Or�0�;;��|��3�1r�D�e�N}���X;1��Pd"O� u ЦX�r0+�H�B��#�MS a��kGs?	�/���2 (3���lap�� l�t�i�&c"��Ɠ,x�5��@"�`��"ޖ"!h�a��\�.�qRO6�Oh�RC��CO ����9l=bT�0�'M*ԓ!�:i:h\�'.�jW�E�9PRb�ܺa�6�h�'�j�JTB,F���[��*]�lԊH>IRm	([�t��0�&�'�L4B��ѹK9��*�)\q��ȓ3
NU��I�4�6��t��-=Zc��O��Z=t�Y��L��R�@��N���g �-6q���t@04� �&�0(+�E�����8��eO�k$�)���a}M�u�!�5^B6�3e�	��<��ޞE8�E��>1&��m�bc���v�c��h�<�g؈~�6=Yf/�V�,���|�V�$���H����^<�¡��~� �O��>\��h"O��Ն^�'.��0��p�� /XlqOr0Î�Y��@�hG5 M�H��"�2c��Q�j5D��)q Y��<� ��Yq쫀�5D�D��ȓa��1�[/m�1"0*5D�|:s�¡[:J�����VV����h<D��eC� s�����*�R R%9D��Eo�6���zC�� ZQ ��dc7D�@۷o	40��y��U�)#~|���0D�8X ��:
���w��"`2(��#D��S�ǝ�I��,8�M�&2l:t"-D��t7E��F!�rv���$D�L�EMӰ`����bU�`8�m�SK)D�0b0��Z�4��h��3tvlX@*D�EW�e�f8S�Ω�X��(D��@�	��8�q쉮�]���0D������� )�7%�������/D�,��AS�@p�{D
'16�x�I-D�l�Vb̀dg$!Y⩃,m�`����*D� �#���>��L�`⏰	x%I  :D���ǿ~$�lVcM1p{J����=D�#a�N"]�ژ'��UV���4�.D�D��	
w��B�����.D�4@bF(��j�i�m=ș)��*D����N@�κ��%��0Y��XE�/D�� :�:��_(e�XȀQ��=ӈ��"O^��E�t�Y;d$�$]h� Br"Ob���Μ]�Fx�V)ʏ{�~�"OX��q"�WhO�!�z�r�"O$̨�!޹2d��
A� �� �e"O�xXS���H��0s�6�F$�"O����"A�`:��K�q�>=�b"O���u�"Tz���a�V��"OxUx�<&lyA��C53�f)�"O,�I׊�m� ,��/��%d�!�yB?B�Up�oԳz3L�*�ۺ�y�+Tp�N� t��s��Aw�)�0?�e՘Y�|�s��?w\zв�`�9\��0S�#MY�<�.�:@@��fa 	NIKu�DT�<)bL3�F�6M ~E�up��{�<qc͌kj��q����oK� r�z�<!�.<\&a��M�b'�����B�<�q����P���:1_ni���}�<! BN�&�:�#��BtdE:�lS�<YuK@�B��͟	��-:p�HM�<!Q`�e�|�§C�AAt��ҏ�I�<�BD�;8C�xH�	�H�J�)�L�<� ��H�;����}ب�z�G�A�<!Peҽ'��m��mŻz30-�P%~�<q���5X�R�.�<;�V�)7a�v�ɼ�M�CN�"��:�u�O5�$j�."̰���/�o}r�����~�퍤~(�|�kW��	���!�=S�H;��� 	c����:C��;��.}��IG.<�e��D�!�	�� �W�u�0	AI�,�O �+0�ة���L�]QrW����O�����&����l��(1|��a�йC�����'��Ot�r�c>m��f��h��Y��"O�e��ȝ	~�F��CH	�X��6"O��J	��k��cC�2I{�AS�"O�`'��??zv	ӦMY�Zz�y�G"O�h !Ǩ;�h���Lعg�U��"O�)a���2���w�60�T!�"O2l�B.Q���Wi�<��"Oؘk6n�@�\���#9$���g"OD��h�	(X���d(Ha"O��c���=Y"Z��D���e"O|���ˬ\5XU)�׋uɚ z�"O0I�Lڎ2>T͙�h��a�j�I�"Oڨ@��)L��3a*��A�~=�"O�\�gfۣN�7��к��"O0��d�O�N(�[&������ �"O9gF��eװ1�!�?a�਋@"O���R��65
%P��[���(�"O4h: ��'� �E�
N��P"O���f��1��SF͎)=R�4�u"O��t���u�X]q��A�F�\H�S"Oh�0 �]�}�F�(B	V���J4"Oz�)Q#�f�t�CA��o���`"OPH���+��Q�V
@�urA�d"O"��f]�o�n���ڦJuP`"O� �g˩3�ډ�����*rqY�"O>,Ctc\�,� �1ׁ_Ez��"O&�)���>iq����nGe�>1�!�$VHB`��� >� IٶD((�!��c�$}�d��=)�)����w�!�D�v�Q9��+Wi|�ȗ��!��=��śq�H@�ɑ2��(C!���J����U�?5b��ӯٴC.!�D�w8N,CeL[��ȟ+S"!���2�����_r,���V�
!�� r ���Q5\ε���%]�ْ"OV	��L�v��v A�%Ex���"O0��jȡ@ �!���B����r"O.˵�ԠHӊ{��Q�I��Q"O
�h�E-�dp�#���bL1�"O���a%��Y��@����%�
��y���%,�&��3KX��@�����y���dX<@�/��lI��qR-�y�̊:l�Q��${夤J�H�y"(��0�JEѥ@ r&�aa�R��y��H�sd�(@��A�B��yrc�	*�T�qb��&�ҙk�d	��y҈�/vlr(�ņZ%X�\�(�̈'�yB��R�fy(u�Lw��j�@O��y2*�1I�ր����!A�`p0r��yR[&���CG�3D���*�ZB�\2��¡�$\8<I1�Mϑ(�C�_�v%X0�Q� >8�ӉX�s=�C�In�d��e�Z�$mȜ	�U>{C䉉jk��(T�@�>���
A'� C䉇䜀1���* ��(��@2H<�B�ɳj��k��
����Ɋ�6�&B��.�j���� :�)曷1B�I�J9����%�U=D��3�A!�C�I�$>�$��d�� ���gK���B�	,F���@���`��HƬ�)��B䉐������60���	�脯0|�B��7��Sv��8*���ǍU�<kpB�I�u��,ABaI-�(�ĆU/u�C�#s�}��ԮC� �A@)Q�t�C�I4=W8 0֨� ����e�%#шC�	��^m1�
�Y�D"A���*?bC�I5-Kh���r���a�N��6C�I�z԰��kZ���8��1i� C�	Yq��b���>7���1�h�BB�<i$�̊r��><RA�'��'��B��"'�mptE�YT2E�ң,	��B�ɀ%I��Y��z�ޭ	�,ep�C�	�^<b8��Ӿu��-���H�m�\C�I$6i�9!g��1�V�`��
��B䉍A%�y�o��Mv8� ��� ͸B��
a[p�ci�4Y6�	����}�B�I'D�F�2�b�9�.x[�#@lXB䉠i��c%��ݚw�]�{�&B�	�.2Ze�E��j!�)���ܶ3�^C�ɕmr�`��\�Cs
y����DC0C�ɑ<�x���Ύ2f�y�4]���C�ɖa �h�a�����+��l�B�	L�\Y�g�K�b)~�`��B֖C��1U���E�ޱ	�LQ(��Fa�B�	�(�X$�GI�(�~ԑv"ɸZ�B�>&�p1�&/�/8�M3�lH�t�B�ɡ'g� z�FI'�Ȁy�D���B�I�}^�k�O�
yN��w�H 2�B�I6f�5J3��
0�	s��h�p"ON�(6�\&�<����/;9���T"O�Yh��� (Ir	�6)��"O�-OO�B��1Rǎ�"����"O�0!��_!m�L���!���"OvQX���Q���gǖ�n��a5"O�Q)7�ىr��3B� �Jy��s"O��R�+� :��h)��������"O��e�*��:!��2T�S"O�z�˄�Lp\b��� ����"O� 0� ��eT  �b�9����"O��Q��[� �i�&�=�!"O"l��eK�"�0�Js�P W�6��"OR�p���%(�\�.	+�@ hw"O�E	#�H9:P|�����E�d
�"O�}�Sb�*Xi�(�J��N��$�B"O���ULWE����D�.�6HP"O�A�D���X)��К/mp�@"O����0={��E̊`a�"O\����� $�4��a	;@���؆"OʍFC_R�f�������m)r"Op�&X�7 P�{R�<.���b"O��aA3+���WK�@�����"OVu�a��@���rV�	������"O��
A)�>fl�����.���@"O<�����p0i�����"OL	q3jF>�t����D�Z�0X�B"OVe)�@�W�\Kr&5y��}�T"O������� BBʘ �fm�H�E�<a�aQ�#���;�KZ�[���1�UG�<Y�)ɜL�9IS$M-����ЫO�<�DG#7z��Ì��^d��U�<q�ü�X�"%��;A��ȂBx�<yF �'צq�a�xȺ�h��r�<р�h�~��ÍE�rM�7�r�<i� ϚA����'��o(1`�"\q�<q�I{����-E-[@<��g�Md�<a�J�42X8=����Z����`�<�3Ҳ=��uڃo�t��4���u�<Q6�P�� ��aKH��`��Ξu�<	!K S�b�CŽ;��d�Pdz�<)&ڕ!Z�� j�e.�,+��`�<i�P�yT���$")�uJRdDp�<�b��W��"@��:��{Q�T�<閦��B�!h6��1������R�<a�"UCZ��2lC{2��c��g�<c!&L'l�X�A�.0��Ĉ[�<A	єK�<������6���ȎZ�<!���-k��ca�C��Q�sDN\�<qŀזG���HGǁ��͛�L�n�<)a�
>s���
#^t���PF��<����#���b�!�9�h�S�Mv�<1�B1WD�%��m̫`>��s�b[t�<	�(b��P2��$.]uZn�<y��'].�S�2G����TQ�<Q�������N�h~���iN�<a`��)}H����r$i� T��y�H�
{ր!��À�n�nD��e1D��{�ƙ�&������2غ'�/D���WCůu�Q�d"mDh4�ů9D��G�W�Y��
c/�/Yw��A&�5D������"Fz@�B>j�� 3D�p�d�)����V�B�R�l�i/D�$ʒBL�
�ժ�k'ɓUg3D�lf��@�Jg��y�� 'L<D���4��3V�T��	��O尕ʳ�/D�xSPo%T�2q�R#At���4I/D���TbDq3���+ո`Ld�	��.D��id�"Վ�`���NPm#�"D���P,�#����`��,BH9g�!D�D2-S�1���RB&�?!+(u��"D��y����╟Pt���BH<D�S�^�\.���$�40���#'�5D�<�/ȯv��`��*�t�E��&D�� D)��רg���!G�z=�"OT�cA��v�}���.l��+�"O:I�
ͱ�j�{�H%�:<�"O��S@CA�u�(����E�.032"O�qJO$d��]Bv�Q����"O��w�R;
JTMX"�T<��S�"O>`��)95�H �R�x�@=i""O>=Sn��x�U醤Ȋ���x�"OV�Ish�*{���У��C����"O(���%�",�h�o�t�����"O������l��D2
�f�C�"O��1�j�7F���b�%ޠ-��E00"O�]���$D`� )�<R�"���"O�Y�r��d�P�v
�"{� ��"O���U�T�!��h�������� "O��*��9<Pi`gK{{"�it"O<a�S�ڡȞ��a�N�Yz�"O�a���%����֍r`��2"O�D��mJ�w����&���9T"O<����A0n���Ǆ�)��-p1"O��	��4|#���ڈ?1"!��"OR��6O}����2�Q`'���"O�M�3��,Ua|�{���k�M�"OP�1�D7c���§Bָ�xk�"OP\����/n-���1a�GD��"O��[���7g=��:�@��2��a��"O2��S��KH�A�&m�$��(
�'����SBR;Ӿ����]�$C	�'p.͂��ƎhB�1�Ȗ�Z���[�'�h(�ƛ]�z�ht�M�H���'K�|PEa��c���<v�^��'���!6��%��$�֏^n`ʄ��',��h��Ģc��,���i`�P�'���ȴ
D+�2Rf,S$���
�'�|2g��G�8%
�'ZB�2d+
�'���6"�>@���	�6��AX
�'BĘ ".~ ��m3|,��'����࡛4����#kR w�$���'����e���_����u��n���'N�±�ۜ��%�5;���'�
@�T���;zd�d���0��M��'{ �S  ���   �  >  �  �  P*  �5  8A  �L  ;X  �c  0o  6z  ]�  �  S�  ��  J�  ��  �  /�  v�  Կ  j�  ��  7�  ��  #�  d�  ��  ��  3�  ��  W  � g 3% �+ �4 �; �B 
I LO �R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr�'��'���'��t�C�	`�J<�3g�@�8����'���'	R�'x��'�B�'�R�'�E���Z�aw�8��T�1���'���':��'~r�'Ar�'�2�'�T��e��]��ĩM #�����'�"�'���'���'�r�'�r�'����E�+��#̆yd��c�'�B�'���'���'m��'A�'��v�s�\���kC�WsԠۡ�'hb�'�b�'-��'���'y�'fzѐ�,ߏwɰMc�� i��p��'�B�'���'nB�'���'�2�'�ʼP&�F���jV�)�ܴ��'��'���'�b�'��'�r�'m�h�6HϣXa&���2^�J��E�'2b�'B�'cr�'���'���'<�6!�93 �r��oX�SC�'��'{��'s��'6b�'e��'	���O	E#� $��[L�h T�'���'I��'�"�'B�'F��'�,�[E+�%�<h �
DL(`�'���'��'���'3b�'N��'��-���z�.�:�O���ـ��'�b�'�2�'�"�'5rdu�l���OJT���ޑ,�P��j����Kuy��'1�)�3?!W�ibdlZC� u�L8;��Ral�8%�0���Y榵�?��<����0a	O�	e�CI�xB��?�BE��M��O0�ӳ��N?1x�C���QAF�g�4�c@3��ş��'�>	�Mʞ*>~9�����W5��"�Ҽ�M[���o̓��O.7=�5�L��8����W�v7P�����O��$a��֧�OP(a��i��G�+��
�W2!��X�?���x��(�y1��=�'�?�d��������e�ܵ0pB�<!(O��Ojto�Db��8PI��t�l`�-�Q>pH���K��D����`���<1�O�3���{��h���3<�P�����ɹ!3@XR��'��9!2��G���� �[�5r�����!�*t� J\y�_�p�)��<Y��"8" p�S@�p2�kC��<��i2m�O��lZP�S�;4����Ysb��2�ʍ� Jq�P��埄��i��mh~�>�&����c4>���	�x��}�l���>�BT�|��'��OO�'���'�/6��R	^�> ��Q Œt���'X����Ѳ Z>�y�4��'I�H����[�l�c�i��=b���g�'�"�e�4 oڻ�M��͘��I��p���4a|T|K�GϰC�9�"b�칇�Ĵ-x���5`\,Re&L�}�@֝��ē3c�I�4��Y�#��]�@L0l�`AT��	֟��Iӟ(�i>��'|�6M
�+����P�⨁���$;z-(eg�S->��٦�?�V�(�I�u2�4
�, @F��	c�l��GLR�����Ɛ�M��O@a�7O���Js+����
�:Ê�/t)���Ƥ��
�� ��<���?a��?���?a�����";fP��A�
-i�6�B�"+�'h�.h�(�rV0���$�֦�'���dع`J��WG٤] N;�ēP��v`���De�7�;?Q�K�0MId�bC��"ݺ%�T3_���1���O(�K>!,O��D�O
�$�O��*���!�P��+��1�6|���Op�D�<QQ�i�4�ɢS��	D��%	�p(�gL�*��-�%�^���d�s}"�~Ӱ�m�1��S�T�H_�I�A��_*�t��F�|3Ы�NT�2RQ��S(Ct�ʈW�	/%D�8�mS�!�yZ7���WnTY�	̟�I���)�ly�b�l�h"���!�� ��Y')>�݋0��H���O�@n��`��IƦ��Ԍ��a��D�M>6͊��.�M�i��d�i"�	�`*�<
��OȊ8�'����Ś:�\�@�"�	���'_��˟�����I���E��oC,e���b!h��)��Г��?ʂ6-�- ���O*�d>���O�n�ߩb�����)��ʄJi&h� �ʦ���4f`���OF4`��im�B6j�T�!ѭ6�I�Ɨ,v���N5<*�R�Fi�O.��?�cH�=�f/�.A'��{�-!#vı!���?���?!+Oh�n���m�'�bgWF�F�+���f����`E�Cr�'��Ȥ>i%�i��7-_a≋d�l`�f��"l����ͬa�(�7	pْ�́f���!K~r�,�O��y�O�}�Al�$��j����`�����?I���?a��h�2�DC:��1���E�q���u��x{,�Ğ����U�Q�����#�M���w̬E�W�P�W�*h��-�:p�$��'e7�Ŧe�4i���iڴ���۠8��Ez�'J��`���G�feJ'ĕ�1��	hBk%���<Q��?���?y���?�tH�S���S�/�_)Ԅ�������d香�@�ş����$?��� 3O}��Zk�yU�(#�Z�O����OD�O1��}��/��_"��KU+��>���y�hY����Ud�<���Ңn3T��W����d������){��h��(rv����O���O0�4���' ��,��;ib�S$y����JL/8zIQ��]�0w��h�F��B�O��nZ��M��i�����P�[������<0�ܱ���>�����rgOT�h����r���� LT���	APX�C��7T���:O��d�O���O>�D�O*�?c�bH=X0D�!�cɒ Ϙh������Iڟ���4!��O�R6M/��I�o�T@��+�0=G���!C�5 2��O8�D�O�iT�4��6$?��B���ˣ.�&��5i $V?H��J�I8�?1Al4�d�<�B�C�>�R�����!�>�۲ 
�O4hm��\�	����I�T�8)b����R�
$KSt4nD�'92��?)����S���	�f؋�(��L=�	x1'�;��H�ы	$1����WW��*'�"�O�)��Iv"�$�#�A��� �'6-�Lf��g�g���P`�=Ru9u��O4���]�?QV\����nT�u��"A'I��@J�7Wà]���� I������ug'A"H���J�eyR�#Q?}[Ǣ��AZ,(Y���;�y�S�l��I�G&�����)^���!w ��4m"4�*��?A���O�7=���q�C\�ec<͹��Z�e�z\�� ܦ	B�4Nq���O�A���iz�$:&/¤����?l+t8s�L���~R&ݱ'u�}�ɢg�'q�	ğ �I8t���9�ͥD�"���Lp�J��	֟��� 74u�'iz6��r����OZ�D �g��J6ᐰ	���v���-��<)����� �����O�H%ɧ0k^5�1_�gV ��0O��_]����`f�<l����v.�O�Y��j���lЊ'�$��fȟh�q����?)��?���h�8���$�R1R�D.�҄c�N�sW��$��������ڟ��I��MÌ�wu:LJb��,�������g�ĥ0�'6X6�ަerܴs���a�4����#��s�'KI�)�0�տq�<��c-�l	�ã7�Ĳ<���?����?����?�!b�����&�F��7��%��@� qk�<�����O�z���wc"��/��V��A��>���?���x���H�:lg��]�<������^�@ �g@��D|����=0��O�˓D��<`D���yq��1ml�I��?���?���|R-O~�m�3c�(��V�*�f��a�|�U/�#������M[�r�>���?yкia�D
�Tu��
3N�4!p,	8���R�֘�̱��X$��$����)�s�̾V;<u)#�K;��б;O��$�O����O��D�Ox�?�
҅ċ%���#�.i�L@rh����<B�4`�)ϧ�?���i��'���4⑇]jPC��]�v���n>�����R��|�T1�M{�O���ש�7%
�$� +>+����/נ`ETqk�MR�OR��|r���?��/g�4r h�8^��@�h>�����?�,O��m�9)]y��矰�Iv�T(?6T�W!�	@���yB�'����?)���S�D�<`�F�+�� {xD,�D�H=P�x���G�s�)�S��?�(R^�[�4T���d�<I�oύXy�I����	ȟ��)��Xyr�}�2�acF�Yw���E/On���)ߵ7g2�D�O6�n�a�G����%�"h/1�>�`��^]b��Q2�M�5�i�����i��ɭ1�>�pq�O��c���� w&4��I�$ؕ����O��$�O���OD��|r�]�YDʜZ���6]q�l2����oʛ6ΝS���'����'s6=朗)׊�6�����
Ɠ
�.a��A�O���KI�)�S+պ!n��<1V ѯ<��=�E�D+?�D���kS�<�sLՓP�B���
����4���DR�"���𣑁*�[���"X�^�d�O`���O��U��������'��W��BX` �ѸC��g���O���'o�'	O61 �f�9-LL����>݈�1ї�����j>�3�B#�Sk9bB��  E+U
.���PE�r���ʴ�ğ��	ܟT�I�E��w	v���DU~ބ�R�ۢp�~��A�'p�7͜�/W��O8�n^�Ӽ[��7T�y٧��(bi8�	fX�<q���?1��L0uPٴ����F����0�I�n]��s1\�2�^�Y��̊������O��D�O����Oj�d^?T�	�rl�E���cZ�x��[�h1�4u���?���?AK~���Dx����M�t�0�X�->U�PW����ݟd%�b>�����5`͓ã] s?ԠۂM0b��pQS��ny�n� Qь��ɟk��'��I��ȺƦǑZ´,�4�ߍ!��i�	��	���i>��'��7͛:O���܁X���"��TX�Iqh�
|���[�5�?YBZ��ڴ*���`Ӝ�0�Q	4��M�V"A3&�h�d�� �^7�=?����!-?��,�������! A����� �	83�o��Iğ��ԟ��Iԟ�r@�ܾ+��a:��P9I,��%G���?����?0�i3���P�H�޴��I.����H���kCBշ<9����|R�'8��OK�3��i��I$��97�/HC&刦�_���S"��p�dN�Vy�O|�'
�&2Vo>���m� �cPe�-R��'��	��MӶeY+�?���?�*�~݋!��'_���"Λ��3��؋�OP���O�|&���x�I����{�������~
�%��N?С����G~�O�z���}�'h�2䣓 ~�Ԁ���C�Zq��'��'4����O�I�Ms������iV?Ǹ��	�OC~Ex���?9��i��O��'>2@��WN����c�$C<�Q��^�b�kӲ ��l��"_��C�����π ��$��I��������4AA'0OX˓�?���?���?)���)��WNH!������D�l�pAo�~˾l�	ޟ<��b�ޟ\(����Q�|���V/*>Ef��?����S�'nGT�!ٴ�yb�S\X��baF1/:��Tb���y⅕(b�	2Il�'�I۟t�I�l�` ���iɘ�15�N9�$���؟���՟�'R�6m�{M����O����5 T�)�U	5�$[G�+O�<㟄	�O���O�O��;#X�V���KF�P�h�N @��X�7�ި?<�=0�`Pg��>;`���
W�
O�pi4��	
��1C��$�	ܟ8�I֟4F��w�Ƥ�k��A��i�*��āv��(e�@�!"��O��D�ۦ�?ͻs:�q(�I�#b��z.X)͓�?���?��Q�M��O��p,V�	N�V���@!z��ur6�]�� �N>a.O����O����O ���Oh�S˞�`�x�֩+0����Ǩ�<�A�i�:� �'���'	�O���F�54�[s�[�H�^�����mr�kޛ��u���&�b>%[�)�++�P��r�Lr�XXfc@�n�X���yy"a�����	�g��'��-I�*�a�	Tx�8���R��FE���<�Iʟ��i>u�'J6��U�h��ķU��{ŤŜnjJ�(�N?u L�$�����?!�_���	�����49�fYb���<QG߉����C��Mk�OV��p�M%����+�	������Āk�\��*��#(�L#�6ON��OF���O��$�O�?E��l�5�R(i��Մ!"<�un�����џ���4J�B�ͧ�?��i"�'u��
�<q��5�Ԣ��pAB��q�1���O@7=� T�B�w���8�V��N��Xc�Ls�P�z,�����p���ʹ�����OJ���Od��~�Y�Ü��~�ȳ�J;k�|�J��'iY�H#�4^��h��?1����I��P��J�bY񥼒:y�'�6ꓤ?���S�d
h/�X񏑴h�P���'�#M�@؀��
!�a��Y��S�.-"�Vu�>o� q�S�Y>U�Hy����"I$��Iڟ���ȟ��)��Dy��pӠH& �N��tB�>^�^�˳�+e3ʓ}��v���~}��'�2�s#� ,W�<	r�6h���2�'�6���d�6�6?IG@��|U���:�Ģͧ:��C���Df��Hq���yR[���Iџ���� �Iџ�OR6Ik�$_?}��S�����3&xӢ1��'�O����O��?yj���+����ԔYSe�d+ !��
��?�����ŞA��P�ݴ�y����yӣ����I���y�A��7+�E�	�T��')��X�	�-��!nՖ�L�D����e�����I�4�'��6MZs����O*�D\���� (ӬR�3W�F#2��㟈,O��DvӶ'�PzƀͲ-P�Xc���H��a�+2?Q��	%|Le���=��'+B�D���?��j/B��1)�͈d%L񺂈H��?)��?A��?Ɋ�)�Or��F�W<^�&L�7G������O�nژ����	���"ٴ���y�M��s�^��@�۾h�@���yR�e�(uo�5�M�i�M�O����ݘ�s��
�KH�tR��aa�
5�(�O�ʓ�?Q��?����?y���j���5'lI��P<p���)O��mZ�]�����Ο��Y��Ο���2�`�h��>����˽��d�����4{��Oql�0�;���C/8/!���@�|� �"\��0$a����nHb�Iqy"���i�!W	&��GDGt%r�'!R�'y�O��	��M��`L:�?�UB˰O֑���okj��æ� �?9�i�O$M�'~��'�2�Z�!���0���)�b��g����i��ɊIp����OB�a%?A�]	׺c�@�p�seoU�V��I����I��T�I؟$�Ie��a\ H�G2���K�JR�/�,<���?I��^�6�
����'�^77��ޑ+H��GE�?Ѝy��&f�O���O�i@8<6M/?��\��\���$R�FLyr�G��?�	8�D�<	���?����?3략��]�u+�'@z���O��?����D�؟h�w�<����=*�~q��O"@	�-	a+I�'�I;��$𦵨ߴ[���i��s|)��g��v����jI����*5' (m��G����7WҎ��ɼV��8Z�%GgRر��� nt�	�|�	ޟ`�)�SQy"�~��8��9^��ꦭ�VP����= (���Ox(mZA��TG�	6�Mkծ��E��S7�ñ'�C��f웖(|Ӷ�y��a�F�F�ͣ��)O�I��mЊh�����/%|qr�7O˓�?)��?����?����)�-gC�T��㖻rw�!����Pr��	�:h��?Y��k~��-e�� mH�~$ ���udp�$�O��&�b>�+�C¦���%b����}#���m�Jq͓9���@��O��N>�(O�I�O���d��v�>PCg��`��G�O:���O^���<aU�idȹ���'B�'�`	���X�P� 5��1u������@y��'���&�D���Ӂ��0��fސ!F�I(�`t2��M�&��K~
T��O����|��H��̨2]��c��=^���?1��?���h�󎒏u[����C0	p,��A�,90�DF���Ο�I��M���w���G{IH�&q��'��<���i	�6��=���צ]�'�]��F��?��� �PKԇ�/6���c��{�%��'�$�<���?����?Y���?��'5���*'�7�����J�8��ʦ}�Ei�eyb�'��O����b��uS񡆡��C�!���'_h6�Ѧ	@K<�|"�E&\6���L�HO�q����_*�����C��d�kSJ�@��E�O@�t~ňee�t�,  v �m���?9���?A��|�,O4`mEѴ��ɿd�^��F���H�F�
�牬�M��r��<���M���i9<�U���M�B��"!��_�����l�1|�Ɵ����V�������(���ɐ 9lx�v%O%y�Z](�8O���O����On���O*�?�(V��-f�4��.T�i�pj5�̟���ߟ�H�4B�Χ�?1�i$�'O��$A�"���eA��^J�bs$>���ަ�Q��|*W�A�M#�O��+5��S���p��K�,�[���#�����0;ʓO���|����?	��PJ�Hґ^hb-J����*��?�,O^(mZ�P�L��	柔��E�t@���u��M�+�Ĩa�+^���d�g}��'�RH:�?��A�G�izBu#E��&p�]㱮���|pK�N8Rۂ��|j�&�O��L>A���`L4y�+���M���G:�?����?���?�|r(O�l�F/�u�!�GS,���R�7�;��WyR�jӨ��ЪOH�Ĕ�~C�c4a��Q��͉Eƣl������%�����M�'�Y���	�?���RU� �@/vn���a�83��c:O��?���?����?Y���i��6��j0��X�kr,G�3�4�lڦ�8�	���Ij�S꟰�����l@"+w`@[�
B�0�A3F͹_ϛf�nӆ�&�b>��va�צΓiD���A�9�  9��}b���~1��O.!�O>1+O��O�CC�J�sJ�+�B�"��1jEM�O����OX��<ٲ�i$��j�Z�8��|���U�OvcT�3�I; ֠�?I�W�X�I��;K<)I�J�8�(U	M����OO~	м��	9v�_���O�����-�©�G���˰'A�zb�X�E`�'*�2�'B��'=r�s�u����5� ,x �OV�~=+pEğ��۴ɥ�Oԟ8�	��M3��w�č2A��U� x�j7.�'2�'��ț��֝!.��S*���1`�X��@�.���h �|�P�������ϟ��I���9@� R���3e�v �x���^WyR�dӈt3���O����O�?��uԵ+4�dB���%N���*��$WҦMY�4"����O����>|�t`�������	B�.`�bS��{�I��	��/H_�	`yB�Di��\S1L�ڀ	RZ�r�'���'��O���>�M��B-�?�CjԞYz-ٖā�a$ѩ@��)�?QE�i��O~d�'�46�N���1�4D�ň�h��L���3��-&7Lp��
�M��O���e����aa:�	�黎�� �'}<`1ئD�!z��$8�<O����O���O����O�?�˶ 'Bq"HZ��N���!'W��l����0޴7h��'�?9`�i=�'{��s��C��cd�h<*��G;��DϦq���|����7�M[�O�`S���0uh	 燚Tm�Ya�������Bp�O�˓�?	���?!��7�p)��I*��ʓ�HyJ��?�-O oZ�bO�(�	�0��N�t+
�~�h���r�8(�%Ԇ���Mdy�'P�� �T>�c�Z~<9�h��(�A��B ?,�83s菂3��!���$���$"6�|B�֗Yd�e��D�Vʾt7ă4Rz"�' "�'e��$^��y�4?Rڵ:vAO[\&��(�
j7I�7f��?�����$b}bKl��+��]�D��x���B�i!���t�I���[ڴ}y|���4��$ݒ	��t��'k!J�'$��� �ꏭk�"Xce@!T���Kyr�'�b�'4��'��[>�k�Şy�\CWm\�k1�@ҷ�^��M[S왐�?����?O~������w�����{ �(h�:��ٖ�'���|��TJҠ���;OJ�cfd�1� ����=9�Ex=O2�����0�?��C5���<Y���?	GC�rZ�l� �F"T.u���^��?����?����D����|,���O��D\1K�d,V?H��o�T|�帥�|��'����?����gz����ԓ(���y��D"Z��'S�j��݅!�D�Xp����ğ�X��'l���CAьj��0�猒O���'��*0��uz��)b�ݷ����B�'��6M��D����O:�o�p�Ӽ{�AҴº�� +�8ظ�@�F|?���M���i��,���i��	m�`�[��O����Sʆa�VH��F�uwL��c�K�	Uy��I�wѠ��r�G�Gm�Ukv�A	9�\�\՛֮_('B�'9"�i��7�2����^/$�x���"�|-�'T�i�b�O�O�*�ȝ-�Դ���$!�(p�.�K���J�\��A�Q==Ab+Ia�I|y�f_�+(zEs�ɏ���P��BT�'�"�'��O��(�MA�!�?9�E�*礜v�A}hX\��@�?Q��i��O���'z�6��lmڞW8ܨ�5���#Jdч�;n~дT�FئM�'��C#F��?o��O��ݻd&�(�ǐ�(|�f	S?�yR�'C��'���'Z���L]��тE�;f�21qU�8W���OB�D�Ŧr��j>����MC�yRe�U��Rj�20h,Z1��~W�'"f6m��iF�Y,6�5?�We	A�? ���c���\NѸ���z��
U�K)�?q��=�$�<y��?����?���L:��HK�$)�mA`�-`4I�����$Ϧ��#��ǟ��П<�S�����޹V\Py�	��i���5-h���	g~��'>�R�ԖO�������ԭ��� %6Q���S�yh��b89�V�\�S <��I�4o�h�6H�|`{W���b,F8���������@�)��wy2�p�2p�`Z>-�-�J��y02��!Ú`����OT,mE��_F�I��xx`��2m�&��1/X�[�B�2c���$��;�mo�Q~Zw�&ɂA�O�B0�'�f$e��,y��a���	f^�@�'���ڟ�����D������	Q�Ԣ>��؀�J�9x� �A�~6m\�$�O.��$�	�O8�lz�����}w. �۩ K����D�����A�)擞k9V�o�<	@���J��7��^�.��f"_�<�wA���:�����O��D�sH*[5��f���W̘)aH0��O��$�O�˓x����"_�	�8�BY�J�M��!�vr�YW��@�	͟�3�ORQn��M��x��{)`�����C(�(�������5���	��8Z�����1�:Z��X�l�ڔs��ҿ5��ɫ�l[_�&���O��D�O��<���k[�x�((H��ٌX�:|��h��?A��i��ēQ�'_��vӀ�O��4�b��BQuI�a��AI0^�fHP�3O��d�O����;]�6m2?�;s�N@h��*���էG�VJ\�11�G 75���9�ħ<y���?���?!���?��E�k���T��M�L�Pi���$���Bf꟨����D&?��I�Pg�Xh���W��� G� �!��b�O��n���M��x��4͌=>ș�FU�f��!��G2x�P]�ƆܨY��ɶS�-[�'�f�&�<�'�z�/
-$w�y0	���(a��'�2�'�����\�t�޴P�:4��U�N R���6����r���0�n�B�:���$�B}��r�B��	�tY2�O݊ٹ�f�7�ŮE{���!��i��ɳ����B�O��5&?����N��B�C�ܠW��-9��	ٟ$�I� ��֟���W��X02dJ���)d��	������?���^<��"R�������&�4ۣGB�k���˔�a�p��ȳ����~����R�\7-8?I^�$����ƕU!�48&
H�R� DH���mkB"�Q��Lyr�'o��'u�/��E�.1q�gә�|�:��߀X���'A���M[F&����d�O�ʧ�$ [����(������;"4��'�"��v��O0O�� xR���s┱"� ���Z�i���M
�2�HM���By�O��(���A�'�Ҹ��K:+�D�3��o��e"��'��'�����O��I��M�ԉ�R����>�[�	���4����?���i��O��'gB 
<�����w�0�)��Odb�'^\鰆�i��i���E��?�)'X��P0*L�
̸�2H��5�Wr��'�r�'��'�2�'��S�6��	4b՛���_�*L���ͦ)QB۟��IƟ$?��	 �Mϻa��z6cabplR���I�|���?Q6�x���a<~��?O*��V��d�`�{.V�~\���q2OLA�.8�?�ǥ(���<�'�?� �D�� )і�Ұ�
�ɢ&Ӆ�?1���?�������-�aI�̟���˟8�p坢7�|�0���7�Ԡs��C��>m��ҟ��ɵ��EQ�-����2 �hY�e_�1����'f ��ҀկD;f-A�����A��'5�3BjV1t�@�q����	��|���'���'R��'�>��I�c�����N(YE�D����9t&��$�M������d�O�)o�d�ӼKK�):�]a1L~�������<���i�6����e2eI����'���qA��?�{����Sq���4���M��nW)�'��i>i������I��	= LR�	�b�K���R�ڂ�<Ӻi�|U���'��'V�O��%ψ7�.���C~�$��P铧l����?�����S�!������K'��ᷧG; ilˡM�l3p�'� �`�G������|"\�T��.��IW.I0a"��5��������Iß �	֟�[y�'f� u�#�O��I"� X��b�m�3S� ��'��O�4n�|��b��ɜ�M�'h�6NV�l���q%��i�py�H��&4hp�i\�I#e����O,v|$?��݉��"�K�:�k�,I�OG
�I��L�	����̟,�Ih��|�B(cO�1w�b�bD/��"T����?�_������d�'{@7�7�dR<t������.��T�	�*�"m%�P�I���S�>���o�}~r)�8:3�i*��Sw2>d��E��c��]矠q��|�R����ן(�	͟Tl�]����n�X�#�P:�?����$
Ʀ�Q�蟈�Iǟ��O�\�)���0۸�PiN�,�,�i�O�D�'��'�^O�S�9��T��(G,#(�1)DI�6�`٘�L�+3O��3rb0?�'_d��Š��Cf`U��Q(D�bzd����?Q���?��Ş���Ϧ����ޑ<���)�ˎ:B܂tUbQ�(|��	ٟ�Iܴ��'�듶?�V V4�B��Yen9ʣiǡ�?qp�i	��վi��I�+Y\zQ�O��"��%l&oABDB�N�!gY���$�O���O<���O���&j�kQ=��b���=��$�6����?�QX�	џ�&?��	7�M�;KiI:��	O�Ȝ{$�W��rD����?�L>�|*���M���� |U�7�5e�>D�bC�TȂ��w<O�X��*�4�?�1�d�<I���?�d�\�X�0�U8:�!NP-�?I���?	������u��ȟ������i�!��N%��ÎS�a��ݘ�#�Y�Q����M�1�i��Oh���K+ze8-!�бU5LM��`Z�K�,�$�0e�_��-�beS͟��^Z�h8c���T�-�͟|�	͟ �	ȟ�D�t�'#�$a�Cڍ}����Y�_,X����'7-��"_��[f���4�ԑd�Z#vt�D%�n�^<Q�5O��D�O�oZ4z�,nZ|~"�ܡV;���#K)�0���p 
B��b�$Hh��|rW������Iϟ ��؟��͑8�@�����;4H!�$�hy�h��y	R��OF���Ox��@�D�\� y�烐
[��HsHA=&�~��'�'ɧ�OQ�@kW���\�\L:ƈ�'���3憶WW(��6_�(�g��bÛn��]y��51��ԋ�h�'����#%�	W%b�'�B�'x�O��I5�M���+�?	���s�ȉ����6JRHi��N��<�3�iY�O�y�'t��')�6�N�r\�%1��+ѐ�

�#h��p���	���O��\�>���o�h�كn�%I�"$��!�p�.��ޟ��I՟��	ʟx��b��?��u����l�B����K������?���(��f��	������M%��`!fb�	�g�	���
����S:��c�O��hܼv�Ɩ��`�n�0]�������%N&�;�D߳6�}��'a�y'�l�'�2�'���'����(@Ȍ\(�m��
�b�B�'�]��Zߴ@�z@��?����IЯ*�$h��<>�����E��I���ĝĦ	�����S��M٘TaX�B��P�B�$R�Zܔ�K5�?2����Q��U�KT�&�4U1���,��𒵧��@R��Iܟ��	���)��|y2�b�X�Av��l�橰d��Q���(���G��D�OX�n�_��\��	��M��i�,\��`×
_<�b1n���y�,	8�jӘ�_��a3����6�2+O�Y�l�d`5��	ӈ2����6O�ʓ�?1��?)��?�����	]�n��q�� !&�&�ŝ���nZ6Nv���埀�	x���������aR�v6�Ꞿ����%�&(��Lc�r�&�b>%в��Ħ��9h��[s@�������#��XΓ7`A�j�O�bH>(O�d�O�$r!	�&�,�C5��g�h��B�Or�$�Ox��<A`�i������'M��'�Ř#�>z��r̉�7�H��S}s�0�nZ1�ē+b^|!iQ�o�=y��ۊX\�'��1yB��:��Ց�������e�'tl�ӗP�$bM\�|qse�'�r�'h��'L�>��	 
������F̤����V�`*1�I�M#�KѴ�?���
�V�4��C�z����7F<>��K�8O��m��M�1�i%%���i���y�
y)��O�����(~��T(�ڬ#!�j�dy��'���'�"�'�R%�>aԜ� ��/[<vE[ӂ�lh�I��M#�蒚�?i���?�O~b��S�c�
*h�b�#kX_!4��Q�@�ܴq���k$���W�>���Y4��b���2/ P�p%+�jGD�ʓ:�t�#�L�O�H>1-O��"ӠJ�jf��S���I��*���O��D�O��D�O�I�<���i2`��'�T���L�������7JL,u£�'��6�>�I����[즱��4\�����2��APbhؖEܵ
ca�=3*r5�i-���Ym�B����9����z�b䄅U\`q0��dN��'6OZ�d�O����O���O�?}5C�9,&B'�C A��T�6�HGy��'6�7�L�G���O"�oL�I�t�Y4�S W[�Pkr,��@���HH>a��M�'��kߴ��$ƂF:��1m�'m���Ɠ*�M�
9�?QҦ(�D�<!���?����?�F)ʬt`�8�0�\?$�|�'���?�����ʦ�)uA�����ܟX�O��!�f��9V��
�ۉz&�=��O��'F�7-ݦ�	H<�Oa�L��)��. �%��/+m� TfJiHF!3���9��i>U��'	��'�X!T<Z�h k���N��mq,�ҟ��I�����ǟb>��'g�7�.`'������*ZQNe�V�2�P<�g"�O��Ŧi�?Q�Q���I�Dp����51�ѺW���H|u��ן��S������u7Ċ06����cy�"�4�p)�&Xnޠm	Ӂ��yb^�|������	����I�l�O���#`�4a�JbC�ʈ6��a)5-z�b7,�O��d�OГ���d����݀`4:P[@e�<E۴�����4�j��	��'�b>i��� ̦I�*��vH]�_.�yD�{ -�j�`Ep�"�O 	�K>Y-O��d�O��� �[� �^�`�!��;������O ���O<���<	��i�.����'�2�'o4�;�,2D� ����3�(T�5��DF}��'}b,#�Ӝq���:��6\G�c�9I��	'l⎀��@�%r�c>�Ғ�'�q���o�����I�5�$T��� MC�	�/������.܌:6��Y+:1����M�͛�?Q��jR�V�4�<���́+@6��һ)Q�d�C8Oܼn�>�M�Ծi����i��ɤvɢ��B�OS���6�y��Ѐ\�N��4�M�	wyr�	"ǒ�qmO��;!�/=��6ěV����'�r�� �X�^Q �_�Z;X�f��R!&E�'�P6������J<�|D�h�? "B$�>�t���o��F@*=3rḵ##V˓[. A�,�O�� O>Y,Oh�q�fS)Q�(��ř'>`����'z6�`��ħol����ӉjJ�h�C�0�N����I�?��[��������I8L��	z cLW���jC"��!(ѺU/W���'8�TO�?���Μ�D�,��6�˃X�f�X�i�:e�`\{gL�:`w�l(��Ӏ3��x����i�|x���̍D�]�k�0q�0�;�I�,L)pщF�Ǡ:Q�QzQ��E�,�!$AP�t��
"�_�ZD0��'�V 9i��N8r��:P���p������2a��`F��� y�V�IT"D��R�K2J�	�ы��dɢ4�eÆ�9d�Ҳ@W���{�F��D�D���ߍL��Q��qC�x�e�� �-�1BR�9�!�wE��P�}A@��/N�K���1����MJ	e��m�dչ�M���?!��h(�z��d�O�I�X��H�?�^=��i�/A�Dc��0��0���X���v��X	�;#�͛,lxq'��M���-��9��x��'�r�|Zc��h��L��hQ�q�'B����h�O���{��'���'�\ʢ��*��yW?-`�BG	Z��ē�?a������Đ%<&v<(�B0!R�H��U�r������O����O"ʓkcv1��3��i�n�8�Di{�Lٞx�E��Y����˟t$�Е'|���O�H�Q�>9�@7 �T^�wY�P������	|yB`� ��l!��>g���&G�S��F���	]�kyr�����'c�}Ӡ S KȽ�Ҡ7b�2|rݴ�?����DR��nd$>u���?��@
��H#W
Ҝ * ��D�����DŤ5K��'�~�0�wV���S��0�2un�oy⅕"�J7�Yg���'��t�4?A�k�<a�"��N]j"'��i�'g�=Z��4��'�����I �'��� MW�D|K
ᦩ�%l@#�M��?���*�xR�':p�+�4{�jxs�� �"\P��nӀ����)�'�?�BN2FK}+�"1�(�c�@�D���'b�'�*p�4�(�d�O��d����P&�(S�B�#䁜��L��+'��;��b��������	�d|(�
�Ŏ�pW4@H�]1z���4�?qE(�lʱO\�?���d����=�Pu�����A�*KuQ���7�>���4�I��'0�T�VɃg�h�1An8��!6�ߠk]:O��d�O��O��~�(p��%�D��j��^�0Ip��A��?����?Y*O��P�$�|�t�UG��|���i`l1�*�k}�'b�|W��
�O�>)D
�3;�Z�ۖ1:.x����i}��'�2�'���'���I��'��'̜����X�2�-*�ȗ� ����2'u�z�D$�D�Ox�$�����xR-R�Y9u�ФHD�q`fG��M{���?���?!k��?9���?���JңC�64�ю�8�����	�0J�'q��'<ܜq��9������-+�.����oy# eɣtHp�yٴ�?���]u�(���?����?����ƺ�ؔ͐��2�J֮ߠC6�Q��i�bR�h�E�3�S�ӣNZ8kꍕ\`����?/]v7�Rd����O��O����<Q(� A���:����@�x1���o}�˛#�O1�x�d� '���0Um�!,
�;u��X�n�n�ݟ\�	�\Zǉ�?��D�<���~R��&h^�}����2i2d��fj���M�O>I �U�E��O�R�'��	��h�'�(%�,�Q$�B�'@7��O�]h�DAE}"R�L�IJ�i����[*af�e�v#α��z���>ч��>�䓘?����?�.OB�ѧ�Ч;�t "cG�-$:��D�͛k��p�'������%�x���� ��X�Q�\�PpD�MfE�� \�=���IRy�'�R�'H�I<x&����O�̅�:tx��!�Ҥ1h��4���O`�O��$�O&8p�뼟L�Iٕy�x)� ��:Z�(���>���?)����Շsa�M�OU�I&eʪ��Ԉ� AsM� �j6m�O\�O��D�Olb�d!�	��9��]$����G/FN6��O�ĵ<�@(����������?�k4�;�8;���5'+5HD. ����O����O2�X�o�|�'�I�2(H4�0�EC��t���zt��R�l�g��M����?�����tV�֘!�&�X�I<L7���t�K76z 7M�O4��J�w�@���}*Enǽ%��t
�͋5+R�᦭�bFR(�M����?i���J�Y� �'
�!�a�F,��"�9r(⇄z�8��gk%��D�'�?9����Y�%jb"Y.���s��^�9ܛF�'I��'N4dC��>a*O����3Qo�R
9 ���"'�&p9�	-�ɪ �t&���I⟸�	������N�*����S���@�ڴ�?Y�c���IEy��'ɧ5&��g���!!��� 7m����^G��O|�$�O��D�<q�f�6���'���8��۠k����f[�,�'Vr�|b�'W")ϮYX����#�m�~Xi6,�=f�aR�'S����D��ٟH�'��m��H|>����D�(P��+R�3�:�tMu�v��?)L>����?A�)C3�~2�U�tȅ��LǏ�R�������d�O���O�ʓ\tn���t"]� �xV��g7�!Q�뇰4��7m�Ol�OB˓Ϊ������D 9"m߮!(����!�=�6��O��$�<��s!�O���5�L�/u̬*u�G�[n�dqcP�����=�&�0�ɯ?� ��SV�Pԛ �*r8c��i��I�^Pe��40X��˟D�S���I�N�ZI�7�Z=��D` T" _��Y��U��˟��J|�K~n�Ld!�f�r�H5_�f�6�Ç ��$�O����O����<�OdPa�P�$Pl�P�Ě^6�I"le�n� ��U��1O?�8�M+[L8y*�&8X�L��/��M���?���e����/O��b�� ��2Ѝ�e���Q��ۧG���<�V�U=8���������/=����0(�<v�J�Ei���DP44� J��p�}YZ��b%i�d��D�p]�$�3T�S�"�Ye�c���	Dy�'���0&�I�T8�w˪�1clb�IџH��a���?1��<��\yw CR�1a�e��m`p�,��	�'�"�')�R����%��t�T�.���Y"O@�p��M�!D5��D�OB�:�d�<AFmZ��?�Ѕ�� ��,��M
�K6�@������	ܟ(�	ҟ��'*����&�i@�c5�t�^H{` h�唘rK�1o��'�T�'�j<���'��'X�d(q���j�S�*�+$ o��t�'����-Y3�SƟ����?�X�MI�,R%EBI��}��k!S	�OZ���O���̖.:U1O���`��$��T$vC����:.d|6�<�`'_R��f§~����b⛟$G˜!J��	�mχ8J�p/p�j�;<x}��m��O���MK���?$h�s�l i�Vp�^ݦ��f��%�M���?������x�Ou�\!щY�H����'�C^�yr�''T�u�'Q�U�x&?�P�X�	7���Xe�3Şpt�i�B�'��]�.��)�K��3g*H$>��5K�b٦G5���%Z���': U��%���O ���ON9#�s��	R��}��|��@��Q�	�V8�J<ͧ�?a����Ě�j��Q� ��e~.t�BE�8%�0Io����a�I�x%�����|�'�6��e�H�!?x��D酵*,~�9��&\ΊO^��O��ħ<q���?���+Aܤ}-e~B��#,5^�ʜ �ś��'���'�2T�T���̳��4'b�[� M�6�Q���M�,Oj���<���?���+�b��HN:��V�����I(���� �i%B�'P��'�I;&�`ʬ�(��
}U���b�D�\���٨c�&�nZ�l�'�"�'��MO��'_F�qDչe�e"ĆD�Q�>�/ F%�I�`�'���~���?i�'<�vq	(7H���Z��LF����]�D��4�	�"(����ħ?-{�D=g[��4� ��%�|�`�paԤ2�i���'f�O� �Ӻ���R�|�aف\sJ,�獌��]�Iџ8ᡪ&�O>�ѴD\NG�I��\#�R�4W"���i_2�'�B�Oz8듥򤈦W�����(	�Y���բy�lZ4u�X�I����'����D�[�B��&!ޗ-�D���◦5���o������|��$��$�<����~�#� s�>��sG
%��`��4�M+L>At��<�O��'�2�܇*% ��:Y"@�&C��v	�7��Ox��� �D}P�t��ly�5���*�Dj�J��7Y��2�습����'���O����O����Oj�J�x5��o��N �Őe�9I����s�3Q���ny��'����L�	ǟ����ʆ6J��5��N���$ƌF���IKy��'v��',�I7'`ls�O ���(��z��� ���R���4���O�˓�?����?AC���<yU��F���G�:p�!:���=O˛��'a��'��Y�`��o������Ok�c��(bL�gO
q��\]��f�'V�̟���韀I��n���I�$3�㙥\ź�y#�&�.��DE��M����?�)O`�1�̏n�T�'��O�r}£m�|�%�4G��*��>���?y���p���?�.O���-b0H	�l�A"��̜WÚ6m�<q�DY�Kf��'k��'N����>��EQ,(��JL�~�,q�/R���)m�ş��I�)j^��2(��A�� �)�� +�-��6M�e�D�l�����	퟈������<4T!��{Ã��C��!��1���ʜ6�y�X���F���?����Fż���hL6>�셺���3:����'���'wYy�(�>�/O,�䳟l[��>T[��D�
L	Fxf�s���$�<��G��<�O���'U��K�̉��^�D:,%B��	��7��O��8�HXe}r^���Ityb��5�ٰc@
�����B׏����Ʒ��D�O��D�O��İ|ΓA��,��/���ua�	��0�T��2|J��oy"�'���������ZBh��(�E�v�هPp�Q��aQV�	֟x�I����Iҟd�'��Q)t>�ɭ7���b7g�u��q�$��?9,O&���O�����3��TrdK���+�h;��G3.�l�����Iğ���ey¥����?�1�d#�ۋL��r�HőL�m�ԟ,�'+��'R"��1�y��>q�K�h2�L�q�\(J ̐�ci�Ǧ���ڟ��'b�Q��~z���?�'Y��M3���pv�T v(��^��@�Q���I���	�q������'��	�)j:ȀEY"x�@���NY�VR�$Z�����M���?����rY��]>nlX��'ҋ{�@�1tP�FЖ6�O��D�����O$���O��>e��D� �>��q�[Gp�Ǣ|�r��@ �a��ӟ��I�?���O��|%���Q�KPx �k%E��o��hp�i_L�x�'��'<�t��MA�? f!�GfW:��@I�*f%�i[B�'��\:d�F���D�OV�P����ak�6e��Pf�,!z7��Oh���O���6O�؟��ן0����[�2�h
XZ �!Ύ�M�6z�L���xr�'Ҟ|Zc���Y�c�輜��m�+�,�p�O���"7OR��?Y���?A-O�]
qmC?s�\�J���x%�A�eB�o����>Y����?Q�{�����]�u��z�Q�1,���%T�<Q/O@���Od��5K��|r���"f,��ha@^Qֹ G�EP�I؟�'���	؟`a��g��Y�g�1F�y�҄dh�C �����d�O����O.�[?d@���4�ѐ$�d$�BÅ Ii ܻ@�IF�7M�OJ�O��d�O*|�=O`�'f�	�Eh[z�5a'�۝g*�i��4�?����䖓L�T�&>����?I���]��!BAE�
&ff�agDի�ē�?���t��t��������y��)4 ŒR]�$K����M�-O�e�&�¦A�������2%�'~�S�D�K��M�$�&����4�?���|��p�������O+>���M�Y��=���6AH��۴A�B�+�i1��'���O�fOL�DE�{CN\�3l�K�Lq�'��	�Ynژ ���Ii�I�'��tG42��E�p�C49|B-h2o@�g�&�'b�'���W�,�d�O������a�l�q��q`�K�+��I��<�ɄvbDb� ��ԟ��I�e) rʜ1*]�3d={�،Bݴ�?q�J�u�O��D%����8Ѓ�`��+]nHU��ظ����"(�H�ĺ<	��?y�����!Ūaa-ռ0���L�27ÚYC��V��矰�	O�矴��̞�p�T*1P\r4�H�R��P8DJ~���'��'�Z��� ?���O0|80l"��N�p�Q)�P����Op��(���Or�DR�C��d>.!HppkG8\�P����Q�]���'=��'�2_�L�"-��'p�27�$���:F�D�5w��hd�i��|��'��.0I�qO�U��#��f����	��PPгõi��'��	�s�(��I|*��2�����ht���H�l�
a��VI�'��',4˜'��'��iX�rt���fи[�*��@̆�3'��_�d��'��M�qR?Q�I�?� �O�)��IN�ɐaJ�J��ic�i�2�'#-r��'i�'3�[?���:'d�a&�7�Y�6!@Ʀ=V�D�M���?���
����:R��1���S�t�ݨ��.g�&�nڼGv �Ir�	���?�`� X�'C7 F�C�C*˛��'��'�J�HE9�4�r�'�n�Zt,����Q[�f�D��-�ݴ��'tz���$�Ox���"op�%s�օ/��Qрg�IVYl����B�����|"���
=��Q�<Wp��Ñ�'	�^����ݟ��'!���:��iZc�_03�8x��:V��	�c�'w�'Y��'��'X��O��$�s����N�;C�Z8XC�i�j�{�O���O��ļ<�L��A��j��][��Kd�ʘ
a�;R��'��|��'�qO�a�D��^θ����,�l�Q�X� �I����jyR#Û7p��N ��[�
�-�������&�ɦ��Ig�	�����I"�c����B���,�k��2@�ӣc�����O`�DJ�*���d�'`��C�-s�@Mz��AO^L���ǞA�O��d�OB<{�t��'�(�kH�5��P٥	�9{�pmp!�ݝ��g�)#��ˣ#�H�HlhQ*�3��Q��~Q�a�+حA�������B��-��Ř�q�����
��g����ߧqqԉy��\$R�Xi�w���Vܦ�zVƟ�`�f�jO�`���� ��3���3�.�jŋZ(��]0qB��T�ֈs�oD�L��u����	|Yp*�<:�L�A �fleJ��H�@8qB� &��@���˼�v�0���?���?YƱ�n�d�O��!��!]el�c#�ݹ=�����"Ux����#��2쓤p.��Zu�'�X���?>"d�R��.kR�Y�H�% � �C���0E6l�4�����2�S���p�֢%�ҽI�a�i*F�� ����Ɵ�G{^� �tG�{�� k�G_�Q9�&�1D���w��m�� 46�$�9�/P��HO��@y���]��6��i��k@��n�֍��)ӄ�>���O:�d�O�8R��O��>͸�C8B������QGa�"���|YrH��v�LIx�P 1o�5?Ri��ܬt�)�r��/��)9�皮>�uC�(]kx�4!��Oj�d�&`D��G0*a8U��>�^�=I��y�B�cD�X�IDi�2	��C��qy��)�G�y�tLB��X��	#��D�<��OPG�������O��Q�ֻz�0(�D���RiV2�'.�,ϊ\���
�&ڳ^�րa��O�Sy/~��T�Xu~��/ʟ-[Ģ<Y@��NA>�"��	h�I�J|�-s�v�jE�{?r�q��[�'�����?���4��	}�I�ޝ��kD�߂�y��'��,��[&Xx$���ĒM��x��Aى'mT�I4@F8ƪ��􅑝H�-p�'\�5@��>����)�HOR�'���3��d�턿,�ڽPנjZ�bb��A��x�`�ѐAc��T>i�|�)� :��%� y���'�,M�:Us���of��ʃ�o�E�wi�0��I&C
;O�q�'$@4%��c')� ��TG�OBHS��'�⒟��>�O�PF��=���IT��-�b���"O���������$KUN��5�6���HO���HL ��,�di��ő�L����px �������	ß`�]w?��'�f,��/�R����kX�ad�y�'�>E#�
�-h����e O��2�I�H0�!��%w�"E�O������_��9���]q8�i�n�+2��qW�S~�@S�����u��Op��<���ɁJ��hu��>8���2�+z�!�ٲ9��#��s^��S!�
i�n�Dzʟ��cB�b��i���r� ��EU����ƃ~���ك�'��'���=�B�'j�(�O,R�'�F��2����X{�$��}�HԨ�IG8�
��"a�h�yV�8 ��&dء=��u0�E=�O���f�'�"�ۚ�<(6�N�a�l+�o؀W>�7��OVʓ�?����S�D!�/[��!�0��ܩ��%���y�"T&S����eBՍE��0�A��y2Mtӄ�nZqy2c�>@�F6m�O���|"��יl��Q�����q��N������?	�GV����i��'�哋Yn�X�L�R�0@C��=r��<�5�(y�!Q@) §{�p�ADf� &�kZ�*D��GyR$��?�T�iaJ6-�O��'m����C/�L��c}�b!��������d�*���D 
�X�8��BS����D��4�?��L�+�L��-��(B��@G�<�1
�a�^�����?I)��%�b��O����O�x�B^A�v���葴|���w$��@ ��ZG�|ҍ���IW���a�����]-w)���D�֤@i��c�|���'���Y���p�x��*�K*�!�!�A��'��'+b�s�(	3�KnCN*�(I�M�r��G3O��$'�Oq"�M>U!楛F��q�!C��	��HO�Sl�<9��T�$�� (֨J 2``��	ğTۤBʮjz� �I����I� ^wr�'̦��0��c�	X�-݈:���!��O�PZ�h�%���������СR��Yh�F=C&h�FMO�i*ց�I!���Cǂ��6쓥ҟў�����Z��taD>6��[r��dH���O~l���/c�u�j0*P*�׻|B�I-8�6��1�7l� �VNV_�(y��4���=�D���,jQ�X�|���Bw�<	��_)0
�yr�F#I(M��q�<yWZ>q�@�q���y�=��l�<I�Ex������@���QWA�g�<�����U	����l	PV�d!��
d�<%L�g��ӄ�0�^5ia�G�<�7aʌ���a&D�!�fQq E�<I� �&j'�+�
����WH�A�<����0����?\�v�Ҡ�B�<�UÂ./��r
[6u䀆o	d�<����G��ӱ������oPZ�<�D����5dZ����ð�	U�<��m$]8�x�Ҁ*��Tː�O�<!w��nn����Z;Wq��:�ɅA�<I�i�:W�l(��D�6csx��Ҁ�F�<a$��BQx|(KY<o���F�@�<gg�B��8M��i�MP���H�<�)�!�>�Q�;t�ҍ���C�<A��i�pib�K�8MQ�3�@H�<i��L�+���G+հ6 �WF�@�<����	
��+t��LHgm�|�<Iפ��/�l��&=f@D�R��u�<��⁑o�$j�!,+��+Fj�<QW��v�\��!��]�}���Q}�<���80�L@��������x�<I�\6��FiϿ[I@�KG#�v�<釂Ƅg�F	�%��t��<���o�<Y5L�\����J�bZa�<�0o x�� ��&߇u�$t"3nO_�<ɐꃾ7��@���,C�@����[W�<	�Nu��c�σN��=���O�<� �l�6��?#:�y�������`�"O�y���DFk��h��K� �R�"O��Q��ɴ�b(BgN�0�8�Q�"Ov���@�P^l��/G�0�kQ"O����e��_�p�O�@9,=;�"Ol������M�BN߂z�0���"O�12�K?-� ]�f�<_�V�X�"ON��fH��h$2��	|�2��"OjX���ޫE?�@s��;ph�	�"O������(O����S�cW�(hC"Ot�[� �'wsxh*��,Fl
�"O�]0��!w��=��T�V8nyb�"O�U@�>xx��W+#rÀ�"O(8��
�R��7�8{-��ذ"O �i6e�:W�j|�3�ˊY<ȲV"O6�+FkS�5��b�±�t"O���b��kҚ5��Og��q�"O8�&�R){n�a��OY�ض2"O���ş� ����F�̣h�(hs"O�`T
A�j@H�@G�c���"O�@:�[�ء�6]�zSv-��"O�y[4aRI��BJE 7_>��G"O荂D�[$4-` �FE��,Cw"O*]�p �9e��y�D�p�B�0"O0�)w�d�������-k���U��ʃ۸h�b��|�#��Qh��{ūƴg�Zq!���k�<��J%lv���/�,*�Vy��*�}�..�FY�5*��4s׎�T�!w,)>��� #8�O�3W���0\@��$"�/7W -�eF3j�*�IC5��Z��&%�,���+��B�:�T�.�>����0�[��O=���0����DT�}$r.-D�;k��-��Q27��hVN�<�7@ňB���zH>E�d��;9t}8ԫK�8ZȘ"p��+�y菘c�F�R�[�/1$y��b���+94Y�gb��0<㫑#Z�`���`J#��SD�a<Qc���5<<%�c톣#4�԰gHβS�ܝC�R`<�G+E�A���pQ���T~�Ժ��T�<��iיswt����W�v�6�z�<�6�	x��A�ǅ�2rйV(�v�<�"A�j�p@ C�:q��Bq�<�����</����^�a����qG�m�<�d��`���8����c�l�<qj[�
b���fT|�����HL�<	��W-(��##!� 0(���B�<T�ԛ:�~�P��X]D�e/�f�<�7n������?H
��@J^�<��S# �����75A,��s�B�<�sMMTY�i�2MX�r,@�<�e})"���O���j�� ]�C�I5n�-�B�)K��e�䋙�}a�C�	�V��iÅ
��&$bC�k������)�rI@`�'#%4C�	�B9���eC�w~���m[�/�C�I�@g6�˅�dB��1Y�DC�	�;�Ց񮓟7��E#B�֦�C䉘7K&�	"oq��0惔�5��B�I.jH-2B�B�L��{B-��5��B�I��\�k��^�yz6��:S!��tP����L�v�Z5#��I�<;!��A�l!�u��n�840-�K!��L�,5Z��#�J1�����D(|!��R�(�S�5(}���&�K�i!�D��nRP���I
�c��;���&!a!�G��"��5
�!%Y��5�to!�� ��!���	v���  :/���I�"OD��ъ�K	򔠡l�#?uvtk�"O��[G��1
�yA	];7X�x�"O��B%��  �<{�2�J��$"O�ؘj�j|�0ځJ\�F=��"O ��s��o�Ɓ�Fʇ)1�@!"O8�؃*G\�E;g��=
���"O`ô��6=��l��9���"O���K�U��h��LP�W�vq��"O��i�M�FĈb�S��<1�"OTc�oI?1'��'.�)'�e�"O�8�k���H��O��LR�"O����+��xŏ�i����"O
��%,D,��:�[�#�D8r�"O��P��P�DP !�#W��@�`"O�I(6��/^X3A �("����D��'.���l�A�c�>��Td��V�uɓ��`�J&��h% 9j��Aw������L�?�x����L���x�ʏA�t�3�֢��[�����o�1�U������]<`��`��S�z��Q��܆>RC�'e�Ɛ����=?�Y���Y�E�N�d\�(��s�N���[��OX�B韽�q$>
��m����/�2Ȍ��'1|O�pi�ٿZp9J�4h��<�s�H�V�`M�9�@E����@���H%+: ��":Fx� �2¥  i�F� �G��0<鐞x�O�+��-��� ���0���y��~�cU	 [�I1"�>���dz�(hI ��&:M8Pk�`�@?�lcF' %m�D��@�'*m�d��af!B��X�Zc��?P,UJ��b2����3�(yG�HbU���[�T�&片1d��"R�aκ�K!`2�Ĭ�3pJ�T�Ou���'��^7@�㐧xx@(�'��xȷhU	F�uB�4'ndi� �g?�t �SҶ3�ci��Y��ú���)����8�4���8GI2u0� H�!�~J��'? ����L�'y*�!���8u8��
�� r{�٪/O��jb#л3��_�J��-c'���O�	`��i�n�3�0�����I�NJ�b��)xn�7�6pM���Os���#��>� �%��+�L{�'������2ؼ�5h�T8��+p(�%-�����	P��7��B�X�f#��?L�bT	(;�0��~&����%QW�)�3��BԸ-��HI�Bቑ�f��C	-'F�	��k �g�O��pf�߰ 0�O��OF}Z0����Y&���rIC�^y$9��'���o��=�Ip��4��������㊨K���Ʈ�����?�D�Z�'�z�{��O|��y�l�)f4tfk�',HI��	��o�X� ���3t����͝�*H|��f�'���0;Z���nxɩ���*�4����2䂆
J��V�	ED�񤏌q�xM Wg@!���^�6���C��&4�6mK���q�	=Z���OW�)@��5^w��A�1)\�M� ���߯d4�i��	t؟�X�2�\�q!��mu�P����-�=�ee�U��i}�p����,_**g��<-'J�m�:"p0��@�i���ɗukX�z���B-��q�Hڋ����3���MI�5J�i��;,����Z�;��� [H�; �ϕR���3�!�i0��>�ᩀ+7 ���V ��p�i��p�- )C��%�`ų�ȓ�_��@ZT�<��b���r%Iθ_2ƨ���WI$����!k��[�x��pH�>�p<�F#ו0�0�ڍw��l�� 	�(��\7,GB��:'��d?���ڪMpR��[��-s�Ń�.[�L�� ���3.��6�/�Ok,� ��t@!�υ1� �Sw ̂��D4�~|YaQ;q����0�A1������ YiL遑f�	wz���㓂1�) ��!OxM���O�__��"�@�B���
7�J�@�B!3�%�<�N1�C��2��IĘ|B��:r���K� c�"��w�������}9�ǅ@��5J�9`6�G�:���g�.y�@m�d-̝k���2$�*=F�%܆i���	�鍲<�}x0+
!Ӹ�3d ֺ �)�'���G3��6���`���߆3T��Q����I�XCխG��|l;EI�(A�X��`ρ7P�z��C�ϦsԴ�Sč����Y��@�Оx�.,°��X���{�� I�a~��w�t�`�b�
���Y�e>0:� J�qOf�*��j���
�G �'�������u��ښbh(��.W>.�xIB��R,'�џx��@�y�m�#E�/y�0���x����Z�=�~)a泼X�D�I���O:Y�@�Y0X+�L�S%߾?�1��>1��(��s�0�B�23��E��(!��ajo�؂�-T���'�аd�?<:rձG��>���z  �.	�@��+G=��G���G��퐄$,O��	#��jd�|F'�s���J����PJ�p��*�' ���:����t�����9���4�Zl>�ٶ&Οz}X\�"O�kq�����'�j8#ԍ�$p��ѻO�07�3���"�I�6������ �S4�P(5n���N̄Tt�g�'���s&�_(�UJB�r �����b�Zgc@�,e��*�H�+=�q��	�z�\�+!��ҥ�u�ͽHZ�"<�E�"`=*��QN�oİ�HW�\�;���k�f8�o�0�~H����7�LB�I�@[�-RDFQ�*��t�+�p����%��!�
�+�lX��W� �Q>��16�*���.X�F�H#���C�B�	��xD�!m�#tͨ�y BZ�c���ĆW4:�=AӀB�g�$$:"$�?�Gz��pZ�[�,̝9�h2pV4�y��$q��б��W2CVJ�:�n��y��˵2�z`(7�·5�6���Dɢ�yBfH��H�E���
L�E�ǻ�y�mF�Ap��?Y\��Dϓ)�yB#�"Ȋ9�A\*ezԸ#�U�y�I�@�U�H�sʜ�S#͉:�yǋ����Ƨ�d��2K]��y����`��C��6�!�T�y�bǹ��y� �[	���f�T��y�[�9!�-���%gv�$z���yr��/.����_��a*ꑕ�y���r�LA�3+��u�i�mI�y�#�#�:-���6d�n���`�%�ybeޜ#C�����J&\� �;"�K��yR���Pqtf"��9C`H��y��8:��12�FD�]��*�yr�A-]� 	���Ý;���s��� �y"S�mT��q6ME� ~�qs1a�yB��a���A#aݣ'��jrCH2�y���1/[d4������]bb�ϵ�y"	j=��O]Z�>��rl���yr�%K0�h��˾OJ�x9�c�7�y�%ϡk�`��G�<Y��Ȑ�ڗ�yB�)�X5�� V��
���yr���AD,��BG�S�|��U�A;�yb� ^��5@&�[�P��m��y�aH7D���Ǩ�AZy9S���yR`�ʀyx��M�<�j�*3�P��y��:Mj�Z� E�:**�J7���y�ކ-#�ɵ��'LhA��ډ�yRn�'*<�G�H+&�z����=�y��3#qİ�7�V+h&�r�+��y��]"g�] ��E�\!@D����y��y
��H� }��������y"�0ڲ�h#+V%z��)!�dݨ�y�c�����lQ�ɩ�K��yr+K�-kr|ؖ�ǥZF�I�Dߦ�y���i�~��ϕ>c�Ȩg)��y���e�Te�׏�x�c����yr�^�Q� ]aV�//�����K6�y2Cې%1*��ܰ� 0R1�O��!��D8�x��w�~T�C�n�!��I�
�d1�	Āp�F�x�.;K!�d=�����̖��qH&X�y�!򄛼T.i�4�S�#�Z�2�AE�!��G�f8J���-�@��D�e6!�o>@ݹ�.T�R���R� O	\�!�dv�}[pH5�!�r�8|�!���RpKU`ݹ�`��S./Y�!�D���pQ��(�d!GgY�B�!��q�$Ä�, �9�t�#F�!�/4Ĝ3򥂀oO�����Ft!�$�+%��c�@G-A*!�U'�9a!�D�D�N �w��A��:�+�3�!�ޫ��£�:A'FYԈW�{�!���P&6�#��ԾX�%��*�%!�� &�#�"ؕ+�$���o��(����"Oƭ��!ɒY(��oZFf88{�"O�Quˋ* Ќ�k�-�8b��L��"O��QGΔ"k����Ӫ|���"O��`�B�Z.�y��X��(\2s"O �y��x�vYI�J(2,<�r"O\)��!^�T����k'�!��"OtU��ɑ�ĝ��Gķ ��*�"O�0!��+(r���)�
Y l�3"O��gɍ�D$��Ȅ|[T��"Oܭ0��IA�h���G	�,Y�"Ofu��N��|P��OX��W"O(1�����}���3&» ��"O�� �I���uR��F>~v��"O�"��<���c_;dh,["O�	��ͼ&�ΐ��Q���%a"OP�*��Q�t����Ѡ��@��]��"OJe�K0D��Q�)߅~�22��y�����杈,��ل���Val|���3�y��39��7��	Yx�@C]��yr��lZ��dJ@5yq@E�X�y�ɞ;>"�`�E5$+� E��y�k��P1��[6�{�l(�y"�Zc� ! gT0���#%��y��M�m4L�����W8$�b���#�y�Ɛ�$c����h�K�6�R蔌�ybƂ�yH��!i�/:�@YAoK#�yA�n�� 9��S�5�p5��� �y�kN�?.U��?b/���ìS��y"�W<#�`��d��_��,j�@���y��
8i,��;r�Q���Kc�2�y�����<�I@M���%+c���y�,ݶz�B=�EB�/�q���=�y���z&��am�{��r6 ��y��M�$5(�a��x��c�e���y� �5M�@�gJ؀p�+%� �|B�	m虪��@U�p�;R��C�	���f�Y4{H�i �-U"^rC䉈BKԁ�uhђG�P����bC��&H��� 0	S$O�`y`�MI��C䉘~f&(p�nJa���C��Y
�B䉌:w��j�*G�c�����˺$��B䉂I����AAPqd�!$�� �\B䉾;�@��&O%H�r%�ͯN�"B�ɘ'�n�Ꮟ''���#��d��B�	�+�^d�ш� �$��f�@C�I�$F��xF������G�C�I�$y���&�����͗D���[�'De&�^�K���ɥiL�hw�}�'@��I�n��q`��(�:b�d	h�'���{Q��o����5o�cg
���'��]�elR���di��r����'kڈ���^�k�h�!� ٍi:�P��'��8{�Ɋ+PE�ӣ��a��}+�'�,�!��qo�AXCʄB~��I
�'��S����A���
cj�,	�'b��� �\`6H�C�p��U�'ʽHe&X<r�JD�$�Z�n7����'�0����t�����Ƨtv6�q��<$�d��O'TԀ}���̓D���9++D��G��t�,)�Q�'�]�q�4D���ag�������X��,2D��hBc�;
�Hh��ģ}޵��#D�\�p�O�S�t���{`M�A# D�� \��b  0�=a7�	#W���I"O�,�T� ��ڳ*O�!X�"O��e�0*�de{u�U%w���ʓ"O
=30`��}J�(D @٨�)�"O,MY�H��E��R�J�B��"OT]��Ƒ�5�B�a`FM�te�b"O2�2���b��� /ӎ}���Z�"O�b�g%2�j�
�$�}���"O.��G�
=	���V����r�"O�h�$O�.�r�fL<x�\ �"O���W鎄y'2)X��Ҁ�3�"O�`�ujU�+$4�ge�kÜ�w"O�J7��A������,_���(t"Oh\3ꈐ�n4�d�R`[@�1�"O�cՍI����%��|X�0��"O~%aF��!���{%�ESL��"O�(p�I��b�@�j�@͵G#2�
'�'��	�WO��! N�*	� �:�)@% ��C�ɗ=xd�� ��+I~,U� 9�tC�I�@��`��ֶh�ڤ�$�P<�<!��T>m�BN8M��h��JK$n��	3�&Ѷ�hO?�$E	m�$!�Gʏq�vIk�-�7!�I�`��၊ZϾ�[Č�20!�G�=����c^3f�N�2+#a!�䈅/��(2�ˁ1��)��	֔{�!�$HBE�t0��N�l�$�X�F.p�!���&10@����(�����1~�!�G�W@���c�)�,�r0��B]��=E��'_\��t��'�@T{��A�BO���'�Dx�d�N��X}�B�/N0@��'
Y�2�T*	c�L�Ώ0/�
Q#�'��	sB��/P|��a�@*+K����'�H��FA����R�߿L�X�'m�U��'f����G�K��h
�'�`�`���(�ې���?�tyr�'���w�	_kT1���\�s��s�'x�K=�<�O�q�mj�'�n��f��(,��$����j_2�j�'2d(����~���#BUY�US�'��س�+e6�8QcIR=CJ�H+�'?�@c1MK�.�X}�CS�<Ɛ�`�'�Iq���U���	s�9]�aq�'��<ZGA�t�@��Ӈy��[�'ˀ퀵mf��և�o�tq�'��\�U-U>I��k�\�bF(=9�'#�`:gl��)ń$R5N
+����'�¸���2 ;�z��W�UR��z�'����&&U�!��oN�?���'>ex��J5��Ё"��'9�b�S�'�p,
�.I�v�d
�]�)X)��'\��ٔ%�� @Rb�N�#����'3&	��Ϗ`�F ѱ�ߦ�p51ܴ�hO?7m��*�83�E�6�����ɯq!��Ԡp��W딱���"��Z!��5_��pg�O
!F\av�]�m!�;Qq
p��ح1
�=�܌6d!�$�6���*Ʊm0�����:t�!�$�O*�h�@�w������x8�p�"O�iG��l	3W�gF*�1G"O�	�dH�\k(��LY6x�K�"O�\H#[�w����D�ҽЬ����J�O�0Ґ#^A���0��-�"ts	�'��\�l&@p�ݳ'rrH��'��Q� ++L����(m��
��� ^��p�;aCp �%����@��"OT�3B������D��t(W"O�|�K��&����8F��9�"Oδ�WjE�wmPI���� y�0I"O,�ۄ7Q,x��1�ʫI��4��"Oj���k�T@�����S� �'"O���M�X@(D��។\|�A
�"O��1���W��� Q�M�)wV, u"O�� ��
#�f�sV��<{{dx�D"OlL�`�>P��bf���9o~�r�"O���֨_���F�|~�!��"O�q $�M8U~�81J��{VQ��"O�]�5�ɠ	��2�h��uqJLI�"O؈�wҾ'�ݠ�͏U��-C�"OR=���؜1V��eb
6$g��F"O�����K��	s��E~T����"O�ds(�0E�*u8���J&�"O�	:�)B@(ڐAІ�� @��:�"Oz�aGI.h�b!��c�5z�bQ"O�M���Y�����0� ;�D��"O��3�H�v���9���Nq��"O��{f�06w֜���݇33��"O����V?�0��F�A1�Q��"O��&E��!�U�r�,��6"OF����5=�$��-�����"O-�T��^��SGC�:	�v8;"O��T���"idQA��&�B�Z�"OT�[��&ex�ZƂ�=�4h�R"Oz�:�Sn��0����"O�����v�2����D�xp�p"OfL�Gm[�W32�Au!S!r��� "O�ӦE@-oJ�z�C�ٔ���"OBDÀ욆�Z�B��D<� 8y�"O�dʑ��G1�ph���-[]�� "O�$�W�Շ*�JT�FMTt�rDQ"O��蔥�j����տd���`"O��D�W/q9���A�l�ȱQ�"O��)�@_�5�� ��^�@A"O$(���U�beP��JӉR���&"Of��`ŉ�זܱE爂&�r!�"O0(�4��?e��p���
�\a� "Of��bH[�D�Y#�DF�	����"O, �Î��;� ��H��=i@l��"O�Ի&dL�[n��"%'��T_HD�"O�(�d�s ��c�)lUnXa�"O�܀s�]�'��qKgcǲx.�H"4"Oby�v�C�E��J1I�58����"O���B��	T������a����"O�dg�7��sKՇi��M��"O����O#&��37�R�H���7"O����ê�9AT�K��m�c"O�u�"d�(V�k$e�2�AU"O(p��I�D ���ڭ@�u��"OP�J��?�(���C�:��i�!"Oj��M�A�I惂x�f��t"O`a) 
B�.Ӻ��F��6��Q�c"O���$�z�X��!�>Z�D��"O@�x���΅���zx)ۑ"OD�R��ץN��w�ɡG��{�"O�l�fo�$_nP� L��E;�T��"O��Y���c�^��sa[!#4ژ��"O��h��M�!b&W̴��A"O��8���;n8����I�9�5"OLQ��Κ
��$�u.Q�$ my�"O� h�N:~�֤��'�3��"Oz�3��_-j*( �&L�7�~ P�"O4(۱66H�Z�)�-`8J7"O�q{g	Ͳ<��JpF�6(��ѣ"O^�ѧPWx��EՂE���%"Oд�6@�d�P�*բ@0�201"O���A�AL;�|���x6��"O½xTϞ#م�C�ଘRT�z���$V�q��84a@� $��Dʅ��y"�ۯu����M ����ˈ�yb���u���I���-�xq"��,�y�b��2�J���F7F6U�q�&�y������  �=,,�A�s�,�y��Z�HTwŋ�)}�!ɦd��y��<M���Gm5s5�C3�y2���Q����*k��]��K$�y�EÈ@�z�|+fFZ$^Mƅ��'� i2�H�">�����l�0ZĀ��'u<��@&u���2Fg�P��m
�'B<�� F�<�
u�uG&;��)�'^�q��	`)^ؐ6&�/<j���'�(-h�I��]�؁��)bB|�r�'\{���=���ɵ��q1���'1N��`��A��`��S�W=$��'��1@e�N8��!��/A�JӂZ�'�b����gdD�b@C�B���"
�'$�y�,_�T��uyS�|�blP�<A[��b� ����	C�C�<G�ӍVؚu[��Fh������\C�<�OܺUN|�!�!W���Ňi�<�&��bYB#�K�h.�Lq7IK�<�KW,4ۤ��u	��w�@�p�R�<鲦��[�8�T䝁C4���b�N�<�R��+V���I�k�j�p#�GN�<5a�.���kDc[_o8<s��o�<���=h�� �,U2`��jk�i�<�&lI�!��s+�т!$Wi�<1W��<#h�Ѓ�疬g�~�R��Sf�<�Dl�4<�DT���F�wM��enb�<���S͊�����)^cZ52��v�<Ѧ&���(2KԺl�0b���W�<��e��肰�:b��#��J�<���!L�,� �8<�ډ{@!�H�<I� Ի_|~�����l��H��Y�<�u� �-��E�G�Q5�����A�n�<qS��L��!�t��)�0�#�F�<i1�\�1h@ږ���r�����_^�<�#9�<�PcZe�:� R�<��oV8��#�f ޲�f��U�<G��=N( )�#	��;��Q�<i3+K�=�6(�W�X���1CuC�I�<Q��|��Yi���&x�Mc�	G�<Aƃͻ9�|��bcM�L��� �A�<�D�ڰr\Ÿw �+ ��qʧON@�<I�mK�M9��a`�<3�q�Sl�{�<�Ǯ��&��a�nڸV?��s��q�<�$Nބ]儽*��A�p�S�i�v�<A�C*젉���]|����UX�<ac"�4^v�� ʃ��8<3�M�<�p&G#���;��Ɏv"[�'�G�<q�f�;1��IHBB����P��,�j�<)f\�mP�m�6DT�RPr}2Q��e�<Ѣ�^m�Ǭ�e�2J �_�<'
�K'`d�� �by���*T�� p�Q�hVͬ�kaO��I�$��"O�8��(r<�����:Z����"O�0�p�ٗ�Q��
>e����"O����)jk���k� j��s"Oh�Hw��2��y��Y�xo 0"On��"�S	��dqpC]�"f��R�"O�<���k�v��+�!ZV��2"O �1o��:e|�Y�jͩaaB�@�"O�\a�I���e[�)
S?>�R�"O�ř��A1!4q�ت^~( �"O�P�K��	j4br�.e$TH3@"O��(��h�����'^�h�"OT52�d&7$�{��Y�[	�1;t"O�e�B��X2"�wʑ�Jn�"O���Qk��<�9
2��9'�&ݒR"O�5���+QF]��>�%�"O�MZ��(I���`��K3K#�i�e"O�MSB$=��Ö�Վeb=
"O�4Ï�]�)1��Y�n�|t��"OT�@I�6�t�0N�u����"Ozq�$�G�H�#�G.Өp��"O�$�8��z��M�l@14"O,��c��P<���
�U�R� &"O��X։L�E�.���� >bX�h�G"OPSą�]v��"׎"=$yU"OH�(PEJ�[Ɯ� BB�o;�;B"O�5��.vQ�ѓ%A�Z�\���"O0�K �Ag�  ��=!~�A�"O�ī��ܓ`K�����bl�"O�!0�BJ��L`���`j�i�"O�������B6��)	�Ds�*O�D��YZ�����؎{�����'���A�	 0��*͞���'`T��f��r�A�\3s�~Ȼ�'���c%�y�x�y&l\�iSf���'\&,J��G�V�b)�)��r�,2�'�2d���L�H��x��i�*"�`�A�'�0=�C(�f�tԫ��$� �'��mz�E0"z C������'��T�RF|�Q�0�ܒ���9�'��c�����ĵ���M ��y�%y����X ,�{��߄�yr���+��q�R'C�t3�xXW��yC�.w�ȜaT���>j�E�6����y£�MeD�pêِ3QmA@���y�o�
�ҝȥŭs���1-"�y�fZ��v�҇ː�8�^'+���y�F�F���T.�3K�uk��޻�y�J�+[�}*�m�5?@ك�.԰�y��I*	M�iQ��پ}i�yhPc��yrʄ�*�eA@٪M
\�� )R!�y���
�i��F�[ͦ��R�J+�y�R?5X�4!�;��՚�՘�y�
pJ@PG�~j�"m��y"f �Ce���q�'~�����A��yZx�ᄄҌJ�q�G��W)n����񳟈դJ@�>$9��]�,qAf�"D��fB����;���g��K��3D�� �?�C���#J�4Z�'5D��	�
�5*�~AP����^�l��e�8D�	����8�P�`H-aL��'"D�\���~�%H��Ȗd01P��%D�T��nA�vc��Rq��E/6����.T�̫ZRdX1��L�x)Z`���y
� x�x� A�,٢���)m�0�"OD\��nհCFf K�`�<K��)�"O�1�Vʂ;	�9SG"[ a=���"O0����_�#x�,ȃ��'38y3r"Or�1��@hTuR��2�*H�7"OnI)�0����l��x��	��"O�L��bڊ̊ [���3���A"O�	�h�9�TsuJ"d�M`"O�ЋJ�)�rK�GC�FU��"Oԙ)�X?8D���eF&V��]c�"O"	3�� $����
P4�>y��"O��kUI�;Z�v�Ӑֱ|�v��%�|�'��Oq�*�듧�!gj
|�Ec\�,�`8Y"O�<xԀ�Y�朰h\4�<u�"OL�d��5S����&&AP�"O\�Ba$JC�ĨVݡ�1س"O��k+:B�e����H��$F"O>��#Q<ltz��̶v��yK'"O��ϓi��|;7c
�n"2�Q�"Ob\����<;^=�� �����"O���ҵ494�2���6��s�"O�8k��!�Dt�t#V�O�X\�W"O��P�7W��ذ��'*z��!�"O��H�B�?OrN���dB]v
��P"O*E�.�?5,�g�N�BZ0y3"O�-���Z.���2$��&XE���"O�ɃC%�!�����xOR�X�"O�@��(hS,(���(%aE"O>�҆�ݟ � p4�õQ�����"O���c�baٰM6cB IHG"O���G��r����rN͓�p"O����7=�~�cь@�Mcv"OZ�Ka��2K��" �d���9�"O��x��כj�>}g���"�qy�"O�,�eO"�v��ꀐ͸��r"O�$�6U�<:`����$�����"O����_M����ªf�vq�"O`9%F�Y�d��Z�m��	�w"O�ʖ��WT>�ҳj'u~&�"O �iA#%ƅ�,����A&�j�!�Λ}M�yPN]�!�����R�.�!��ٺk�K�N
ss�mk����~!��B8.O���0P�)�e�2G�!�D˔Q��m`�g�"(dk���-!��W�`Nf��b��Q  ���!�d�~�b�D�;bo�BCPm!�Ē:6S����as�a[�L��`"!�D�1C��,l�� ɐ \K�����0=�%?s3�LauI�r��%�3�W�<yƠy=�U��[�q�H��}�<��#�U��A��P�b��j*�s�<y���v��;����%�3 8B�ɒk�@�A����-�cR>X�0B�?c]�I�$�4W� 	��S�o�B�I:5L6�"�-�h����/b��O���-�S���; 8P��D-=C�@����%2B!�Z�OS>���ȕ�.�6�Y咏*,!���!!|�%Se+
�]�jE� ϙ6?�!��&<�쵙�T ��%�r�D�gu!�$�;�6E�2�5TkQ �*�Ly!�D�T.f��k�=d�H8�G�):ў ��mg�E �֙Q?��(�K�o֎�OԢ=�}␥:L>��r3fߐ*nB���G�<�0��(VL���t�3�|<�a�[B�<� �����P?L����
�ț�"O~d���	�vg6�1��D)��y�"Ox���'ЄJP\�#���]$v	#"O���ǲF�����N 4x�8�"O���oH�#���y�O�^kI���'�S�	B�0�`��V��i�*���E�(�!����h����N&����Ԛk�!��ځg9��a񫙓)
D��F/�!�d@��T�@�&պo$ �А�B�Q!���S��0�ף�j����h�!dD!�N�X�F4
B�ЊW2����N�p'�O¢=�����f�,V��=�W��5�Ҹӆ�IO>q�cG�`1�Ý����*�,D��Ȗϊ�J�H�A��V�f�xT�.�O��;& Ř �F,ϘA3A���\I$����ϟ���I�BFk2�Y���O=SwZC�I���$�č�<�4��
A
G*NC��#viW+D;|Zh|	!�
�O0��4�)���	<TV0�j�<#�C�Ie��q'Y��:�
V8E�~C�I$5���٦I�PLr�F��P\^C�,"#^���r��dC��5v�6�OD����.t>�J���B,���1�!��.yP*a�G�
����N��ls!���Q�mIvi?)t�x��l��L�}���fn��V�p�aI�I�µڂ+D�(��ܣ[,�ړg��$9N�	�#D� a�WS���FY�0��A''D����lǾC��Y�ք~�p��t�)��O���&O̸P��>>���ǘ�L5:�"O�AgJY��;�*���P
�"O�X���9SV����.�}�P"Ovi��J�R�X��r�=43j����� �S��Z�a T)�[��H�I��RU!�Ĵ7���s�D�qp��S�@ӝ
Aџ�E��N�
��5�3%Ӎ;�^�z�f��y����_p0)���hZ.�fe8�y�%�3Mv��3���'i}�\C�虑�yb��P�j��c�T�4%�A�<ɰN:"V�Q���q��H��'$�'����9X#>�S�#$$b���$C�I�*�,Y
�%߶:� c�V ,��?���	�hFZ�#�
����u�3ꓐq!��@�Q=� d�&-�$M
UOQmX!�{��pyl��J�\hx6@�eX!���E�Vx;D�	!Wp(t�6��F!�G9<����9a~y���A�qџ�F��e���XًT`܎+�<��cd=���hOq�L�Bw�
� }�ƚ�@pH`"O�����[��k�$ɤ ]N��e"OF9�gO�e�i�4΁*��=�2"OH̊dj��$)H�� nE�\�$t��"OD�!gY,Xm���Ш��� B��N�Or���aK��s�ʶ
��7�H�ϓ�?��y�nͦX��I7&��w�t���ϊ��y��!<�DsѠ�w���
RG�y�� =��:Wf�4B3�����\�y��D?�(���A%:2F�9r�G��y"�"~(��]<.IR\���S��y��:j+2QK��#%n&�)�yiӄ,�i�Ǖ�J5�`[d�.�yb���"-����.B ��t����y�H�t5J����e+v,��n���'jў�O��Z�N��A��`���'��Ձ��� �!pǄ�_��uS$Ii��Q)c"O(����U��D+�h٭i��T�"O�-�#�Z�"�@�
S�ry�dR�"O��ê��$�%bW�S�����"O0D��԰8B ��V,r�
�x�"Oj�2���z���0'�ݵ�Ti�"O�T�-�� �L���'�Bu��"Oht�eP:>�t��Ѣ@7�n�r�"O�C���=�U���"4ht`�"O�]ٖ��awFPp$HS���|8U"OFț#B�f�l��X�Y����f�'ў"~���K�F����`� v V���$Zv��`�fTL�����0/�̆�>%
�X�9a���!.:�ȓf�	IG%N'fK~�0�̆2ކͅ�T�| `�n����,,��,��'�n�wm�i�F=��+�*V����Id�v>� ��ˣ\��SdS�H��0G{��'���ə<YU�D�F��:\в�'aHK����j�p&EQ6�r%c�'�����G;;f�)��o�(av1I�'��<%��O �����a 9
�'��P�g����\��������'[J	�kJ�F͜		��^�s�d`�'�L�c�K�������&�>���]�������G݋Fk(=sf�i��D���O`�E�.CB�#A�y�z}��'���ȡ%�=��x� �6A�4�"
�'M<����G�P�N%9u��4x
��'A0���!<dd�`u/̓,�	�'�,�`Q��7
]T����W�FR�P	�'U�p�2��"kt��C�9�N@�'��hc�ȃ1̠��D˂
�L\;�'[�	��L^�?|v1n�+yϖ�"�'f�H�G5[�Z�[æ�ik�D��'-Lm*��ɴ���%i�
��'�L�8�F��y�d�h^2^K�ԫ�'0�L#�E6Y���p��]"T8��X�'Ť�����I�T�7t碰��'�A���ݳ�%�j���+�Ǜz�<9�@ߞ3��|kPov�@���z�<��Eڇ>�����	A�&��gn"T�hR�������0�����Ls(D�T�� �f��,Kp'Z4k��3«:D�l#����F)�s�A�*E¬���A:D�|���ɵL"����̔�{f�<ҁ�2D�tSwF�Y�bDC7�TD~��K�n%D�\2Ձ�{��!�጑�_
VSW�-D���ďG�G�Ld��o�r,�g)!D�<e�Y�3�� �� �xp}ڕC D��#����]1�.S��2e�(D�t��+2D�0q�K_+^� C�1D�@����#o�HҐ�]�s���ۀK"D���� �X�U��$0������|�<�e�[�P�$B�d��D����c�'�?����JԺYHtm�?w��M+D�Lk`eȆ�&1����@��=D�����o�.=���(��ikL1D�X:AA�8�\)1�R�9�fJ +,D����b4N����#!&��.^_!�D��R�fDS5L��7^Q)��Z�0m!�䇸#ۀ�r�$[h)�����7D�!��ǚZdLʾ �肅�XM!��܆gp�4�P�F���Pbf�:~�!�� �̨���3mB�ᅊS3WbR�J"Ob�#ABv�:���r�4W"O�	��Q�^�VآC���;g^!�p"OX�@�J�.����Ff��}6l�8 �'bR�'�Na2���1�&�S�(��F��q 
�'��i[ ��W]�H��H�.����'vHh���X?��`�& J�A�'�>Q�S�[�L!��
;�bU:�'ڈ��׭M�4�(�E�Ε��%��'ff����&X����%���g4�|A	�'�pM��*I���(d���Y��".O���D�!�%�pb��e�!���,e�!�M�p�~�Ғ��/�0"�H
2q�!�]���P���U�z���G7 ]!�V�"�v�{�� :�2HQ�'��M!��<:: ;�5W�DTP���C,!�d�_��p�ǝ%K�@�ag>K!�F�"'ތ a�C<�8�01�R0o!�D�"@,��#�ʒ�_f���BER.c�!���)��]	W$җOZly��,�!�������iI�uP0�B${�!��  ��Aޣ`Eldh��!5@!�$+(�����A $�15��m?!�d�k&�@���.98	b򎓦*?!���i�~����E��;���;'�}b���iV�W,uF:�`ď�2b��葕�#�	_����cAz��0�@�M�-�$�yRE^a�(A�5)���c����y�N\2	>�ta%1��P�d��y��5/E�!�� �Z.rI@�!Z-�y�eؒ���A4��	Zj��٤���y�F�="�䭠0g�%Et~���ʠ�y�aN�]���:�����Ak�
�����!�S�ON�-��a��xV����>�P)��'�|Izg�	�n���Ƣ��(�]�'���( 	�4���"&��+/��j�'<|��b�B�7#�d��,O�0�0�����hO?u�;C���v�ɅRLN��)�i�<��e�0��d�1��%����Ogx��'�.a��Ɋ�,�Ѐ��Ȯu��ݰ�'F���"��2���dəjR�L
�'�b�p�"�_~d	f��1i��I�	�'Yr]�Q�P�)��`z�DO;qK�D��'zҩj������F
k��ز�'J����L�bV���#�PQ�D��'�:����\�Z<bTř0}@~���'1O��ҡ.�2K�A+0�U�-b�)�"O�M���ۏB�$�'n�4K��3�"O����m��p��ՃP�О���"O��A����e�+��<k�!"O�a�\6lT\z�ʕg�n�0"O �SŮFg�ĠA-�p�Bg"O����/B&}�}��C9unU��'�!��W*�p�>V1x��X#w�!��MkE��R4���P�*�!���$����v`�K���4P�!�䘚��!�Оj*����
�]�!�E�Yk��AmB*:GP=PC+�?�BV�P�	xy�O�����"����D�C�[.����$4�)� F��r!F!,\6������Gx����b̓1Ȩ��D?4�PR�i�oJ*<G{��'ھI�6� hXN�(��@% �Q�'�^a��ܫ(�ʙ�b�NZ�$�
�'�T�j���B��Ђ��IJ�` 
��� @hAQ��^�|�cB�m*�S���'��Olb>���N�z��9"iFS֜�Q�2|OTb��D@�I�AB�O�1@�f�
$|O�c�� !�Hm�4��C��7H�)��!"�Or��(7d�U��'�N��b&Z�9@B�	�A��H��`&�: /k�,B�=hF�)���I�j�X*؁1EB�1/8��J���.���Cĩ*�G{Z��F�d�8�z��tȇBB��
.^��yn]�T}pQأ�VAMLU�����yR(��"b�y��E+@8�|2a��yB��gF��%>ր��	��y"oԆ3*��mҮ0�<�H�=�yB�������	R�夔F拤�y���)�Ҍ�5�A�Pa)����y2��b��� .�M��ef�0�yh�eB4$"R�4��Z�a]
�y����E ��&���.� �j]���=�S�O�-�A��nD���d�#@��A��'�b	+dI֭Mg\��7��3��	�'	���%	Nm|��n��^q�E��'D�Ms�*�''�Hsu��#Q�a����*�'���0oK��v ����R�d��ȓxܜ8�r�ZO���
<R�'����	���c����!��0��$5�S�O���E*�;K>�AԃO�Y�x<��"O\�1�)Ѯ� ��Jg�hjd"O�!��D�{�L��r��1kX.�6"O, �&^�ȁ��j
�7Df��p"O���'�L�0g^s�d<˅�'�R=O��V-̇$��Q*d��H�\؛���9LO,�*�/� ��j�O"~Ìi	�"O,��M^���W��zM�#�"O��pSC�5�����،?fd�	u"Ol��6�Q�L5��n�,Y����"O���#�	�*�RA�L�m�C�"O�$� D�T���bJģ��P!��'9�y��$\)�X%��G�r��&8w�!�φ]M���jJ���5E����R;O������:$8}*�ۨ`JR�cd"O�m�I�YR�4q�SF;�!�"O��`��W/h���+���l+hmq�"O��+U�L F%�`���0ذ��O2C�V�}�68z寏"m��`�0D�48$�6si4y��BOg�*د��y���`�8���0-����6��?��M�����H6���7���1�8�'�nl;`�	�4cM��KP�~����'��Q���h���sΚ<[Q��'Y0���E�<�T�^y��K�'P���ǂж �&�y�M�"�)�'젽�@B_����J[��\��'��yŔar@��D	
��:	�����M�(� 0B�,���p��ܟ!��X�N�01c�� o��p��]!�d�9<��)��E�y��Y���,7!�D:+���IBj!O���Ё��S�!�ӑ:T�����lDya�Z8$!�t�TL�4�ΑC�fL�a���!�$׊]f�9�$	�5�XY�̘!�D�0������_iBm���!�!�Ąh�Нh�K�-[��AF^ Dl!�/ڂH�%H\�*���q�û>j!�ՇZ+H)�a\+#�p��t�[< m�}"��� VYSc�07�6]���!.���""O�mj�$VqR���h�%��P�"O@yK%�Ȯ'��1�3��9�*�:��0�S�	J8x�&��Vb�Ih�oG�X!�d�\ߔ�2 =S|)�î�E!��"vTn�w�uK� �,Y%!���k�8�s��P8v��t�2~�B1O�Q��0o�蔫V��Z�1"O���%�LB0xPm�lC�"O^�X6(�H}p�I� ��F�r�'�dq�G�MYiCf ����Y���0D�t�"[uT ��$�>:^�q.!D�����V�nj`p�O����4�2D��E�='�l�T��hiXZS/<O"<0f��?^b�ꗚp,\�����e�<���β�E�3X��駦D��yRoJ�zwN�"q'�0M)nț����O#~:agנ
8��j��#���̌b�<ɧ&͢P	�̹A&��<Bv���
a�<Q K͗[C���\ �t�#F�Y�<)���jkƐQBn�-�����W����<��	bبB�iA�&!r��U��L�<��h����NԎ[�J�qr�QE�<QT��8��X�'�Ow8�)�AA�<y��O/РI���S	����c,�w�<i�׀KӔ���%0��uyS��y�<����f�|�Y��S�Ɏ�2@�p�<�0K�� �x�+N?Qvf�R��q�<�`튲Vf��Sg\%�90��\cy"�)§lPmY�� ].�zl	}�4	Z��d0O��P���$Y&�	p�p��)�"O�PY�#D�B���H�*�06®L�"O�H���AI���Q�ߒ|�X���"O��!n����F�K<B8T�Z�"O�Ї�&�>��t�`)��͒��y�ĕ�^��0A��8�ap�
�y���yH��2w"�2�\����
��y����5d@���4-�<�s4���y���2$H��u�^"'h�];�ǖ��Py�Nv)^��
�n��D�W*Sv�<yVdI�idhc%�Ԓ4,����v�<)& �x��0�E�8Xp��D#�gx���'4L��SM©kPz�yc*�W��ݑ�'� ��ND�Z�~�[���%�̥��'?*TX3+�/m�ؑ� �,���'�V�����H�b��w�R�
�|�@�'I(]8�Tyc`h�9=���'CV��K��(ؠ�����&'����'��U�ʛ�@�����IB��� i��$2�`@��	�:Z�����"̉9��*"O��"dŜ�^��ӢL�@�1yB"O����cQ�Sp( ٠��.9�����"O�(M�@���b�����&"Ob�1e�3��!����+����!"O�L;�i�e/��J�#�W���A"O�<��	^���@mن� u�"Ov�#Pn�-k�-���_���
5"O��ʀ��v-K���c{�cw"O�t�@l�:v�$��C�R"e�j("O֩��J�%m�F��%��<c�"O��7�θc�ip#��[y��@"O�E0�^?�>Y��ō=Y`&m"O�h*�f޾oj�XG��& R,�����D>�� ��>�ء)eDޤH�0`��3D�� ��; a<J3�I�N�C��I�%"O�Q�W(!�p����%Ѫ8��"O�}�gO+ �*YU��>���"O�D�3aƺ�L��L�U�D��1"O|�k���y:���A�0=0�"O|@+7���cf	B��ʫC�~�Z�"O6�!��^.3�T%`I.��ђ�"OB�����C�,�Q�D��"O�l���$H�K�N��!�w"O�5:#ω;9 Z�^�5d����"O�CO��0�j�ޑ~K��h�"O��Y�*ǈcO��
6��J��"O��P�O�0�x1Zc�G�Z<�8Y�"O���%�C�9C�Ӈ4�`}�"O(@�4L��(TBse:p`L�`"O�<���F�R�Rׁ�%,Peja"O�,e-�Ĵ���mT	h|�BD"O吥��#��q�	�I�j!�"ORT�M�>�����^$r�#�"O"�i��.,��ꆂk�D�"O�7�2 �F	5���P"OԽr��=Qi0�q숏_Lx:w"OxhY���[���8b���=���"O<U�#�ţy���*�F:DB�"O���� R�E�w�K �0��"O���E��"����a��.�y6"O�1Dݏ%�����ȯ(,*�"O��
�e�R��8�cY3�ܐC�"O��s�+����'�E���I�"O@4i�M�s%*��Y���֪��y̯�$
�NV����s.Ё�yrH;N�u��oF�5V� ��ơ�y2�
=R����g
�KRx��Y2�y��[$R �	|� �� ��Py��ެx�	�7Q+h$�q��C�<�����F�,�Rp�X����)�}�<���G�\X��(�3p�둣Bc�<uCC-2�{���)g)����J�<��o� ĝ;� �R�^��F%C�<A0���r����W	Ch��a�F�<�옹�z@p4l���L�Q�A�<1���g�h��i��E�V�S�<�!�ljJ�� B�	?A����.ZC�<�TG�!qE�@��;���A�<I��M�����N�g�������~�<��fĳu� ��B~��`u	z�<qD��s�"���/=9Ĝ�G��x�<Y4/^�2��@I�+��b�2��QHZv�<)�KW�*�¥	����X0Ёu�<9�$è":��¬_�^H\ek`�XG�<�gj_#�����  �d���a�W�<���,�tE��c?Gg��]R�<!���	_	�d��|欅Ђ�O�<���4.88�%�BC&��*�VI�<i���9wѾ岕�Y�E�*)I�#�z�<9Ra��}KZ���Ҥ�2�B��k� j@M]��Qh�h�+��B䉮B,����Ï.�\�wȹ���D0r(����Z�1F�X�A)Ub!��6�>��K�N'PL�Z!��<M<P�J�LZ��eȘ	q�!�d�+~d����ډ{6�{���W�!�$��FZ�pz �A�q�0�O�Kj!�D9*�Q��	"L�4�å�$WU!�� ��Y�'��漊��??^�0c"O�A��,C�\p��L�3Y^��2"O0�#�J^'�|���	?}-�yu"O�`��e�I�ժ�
�"O� ��$~�J-)fBP	3g.�Q�"O�=3����n^$�a�JpEvx�U"O��v2�j�3���&Pt��"O�}�ԩ�/]\���,�wL:��C"OLL�v^�/\�I,T%^?�"OJ��H�3��mz4�Ƞ�0���"O�S���4��yx'J�(s�
�0 "O�ɑ�!	�o�[��ڬ7�yi�"O@͐��S��d����)�Z)˲"O��rO�=*ѸQd��}}����"O8�S���ؠ���G~4��"Onq�UlԸF��|��I@��N�<��&_�li
)05EʗK����M�<I�Ŋ7z�K���0i���U�<&A�'a��kEC�<�&u�<���A�r�p��Ū�]Ψ��k J�<�Q&�*\��*�	l���fD�<��O	yn����뉃:�n����~�<Y׋�jJ������Z��u*f�|�<�`N9�$:��K�_�؉���C�<a6θ^U� �F�#C�|����B�<QWL0��)��쇦X>�Y8�J�<1E�;q.����!\�BdIF�X\�<�'(��`<��C�f6�9)&�B�<�C�	5�P�37dA���#�i�<)2n��+H���k�&p~�	��]A�<ٱ�X�b���_ S��B�^z�<��(N�_�Z����]|t� �z�<1�M߰*x���7�B-�8�Z��s�<�/ط!\5C3�Z�I9ڄ���l��1&I+?�q��`�Gˤ:z�hf�<Q!L�5"�&���y��܁U��V�<rfJ�mn.��.�3K�l��oKg�<����xXr�N�X�zLQÄ�y�<�bȉ��%� #:���*V(�TC�I��NQ��'ƶ@Tx�;��#[�!�$E�<���
��H!�4���׾g��}���|�@�(��dT"�25=b�%*D� ɀJ��|��X��)�)8��<r&�'D�p��]�"J���$Q�$D�Z �ª^��d*�K����#D�P(��SRly�1�6a��,��?D����X=��2���D6`��v�=D����Ą/.ٲ �.S'xFF�A:D�,Ɇ�R*���C�۹Z@0�+3l#D����$(K���J��'��icd�-D�8�P�V�#Ƥp�$�֭0Q�8D���I[&���Sa�4&�9�5D��ـ�O�z�����$V�^�I��&D��S$Ŏ,/�I�"�+���S�&D��*0#�6"��룏�A����/D��!K�BTq�閑p��x6�+D�@X�#7���;tI�	wi���A6D��c!�S�5�&I�tNQ��^A���5D� �n����J1��Y�n��P�5D���D69~D�/N� T�3t�1D��r��_�����%3�$��`�0D�d�v��?lh��W�W%Za�,�3�#D�H@1"�V1~5J�������#D��`���IԐth;5/��� D�� ����ȓ�H�0��@�
_(��"OL�óiہ\��1��H��F)��"O�a�ǆ
���7G�#�r1(�"O^�������2�w�ߏqѨ�� "O�a��,/(������F �%�m7D����e��7;�@�!�*u�!� D�0��W>����F�˧W�a2D�*D�4�p��%�<e:%���V�,銇�$D�X�@��5�T�Ơʥw��ZP�/D�L��FVc!~QE��<��P��/D���`O1+
xA��� `���Q�2D��	�hԬJ�ā�N�?n ��2D�������@���^�2`0" ���y��B#2B�@S�Q �]��³�yBi��i��Ĩ�
4N&�x�)L:�y�a��w�b9ۣB��|��P$���y��҉8=�!A7�M�s��ɠ�4�y"�� c��DX�Cȕp�đ��OC��yRK�S����e��eI<�2�З�yb ��R��5�����\5p%@����y��$��d#�o��)��ް�3�'r�\�`D�	u���A����x%4�+�'A��AY R�aEr;�'��X\H�P<�'iϜf�\	��'�\H�䙒yBVi��ZDz�'�d$�L�#t�i����V�"���'�����(�d�� J!�OwTU�
�'�`u��I�O���� !AQ����'F\0r��c�n��捝-���*�'Nl�ƆP�BG�"f#�T��R�'�DA�uڥdXܙ�$�e����'��6LɑBP��K��\V@��ʓ3` x2!.��T�MĒ
���ȓDiP�u��:K�"���eG�sV I�ȓd:R�! �V� ��
����[TNأn�cf�+�H�IP�͆ȓ��	bU$�� ED
d�Z�ȓY1�����x�Z�����
1��)�ȓzl��s�d��]��$��,�p�ȓ�X�Z5o&J�����&}�D�ȓDu0H�O�3ͼ�Y���?Y2�ȓj�^��0��lP�DJT;Qq�х�}"]X��gi4 �5.ޒP�%��q��@g'��Z�p����E�-��I�ȓX"��",�;$ �Iq���K~�L��	�Z�UJ���{�!�p�1�ȓb_��A���\=4#SG�K��9��9'��PѸI����2憚%�~|�ȓ�����ΑS��Y����*�@M��XC�=9�f*: ����O���(�ȓpMfMz!鎲i�qx'��*D��ȓ e��2/�W��و@ �v�0���w�, �H�u�JȘcO�R��P��tR8� �"ͶF"�<3A@H�E*���ȓe�^Dӣ�8-mf�t�̈J��(���X�8ªM�h
V�zp,��'x���ȓU��*���;R�2]s+ ;�.��ȓaR���� ;G��Q��3T�24��OO�!��K�ri��D�o�T4�ȓA���T-��|��T2~���	n<���<
��"�GϠc�T���]�F�h�Ѕ{� �7�	�[�����FӪ%կN�-��4QC�?�\���2�VC��Q_5�Y��a�K���S�? a��LR$eJc��4��x�V"O z@G'��h�Af�k��d� "O.͂���$N5��Xu��;%"O:<x.Z��t cc�|���A�"OX���#;Tl����tt���"O�E���C 6��᦬X�S\� +�"O0(cA(Æ`K����)���P�"O��`Y?S=�"�Sf�����"O��E�0~�utl�*S���E"O�E@�kP%"x��KS;kĶ�2�"O�ā���7�� �q�2�|��"O�����;~�C�d����U0w"O��:�$��gdYb�_�j��X��"Oy[��G�l)e-E4x��&"O\<y�l�9-+�)��fB,�sG"O�E�"�:D�4Q�d.wn=9�"O�8r �I�Rp)�%/�����"O�ɢ����k@xa�	�
���P�"O��@U�M52�� �U'T#
UR3"O0�per-�Ix��P��x�1"O���Dw)q��M�_Dl�W"O�-���<��Y��oL�?�ԍ�A"O�嘗���7�(��+dI�5�3"O���'BA�r�|�dNZ�8V½@�"O|������P��`s�u�Q"O�RP��S"m���X�[�t"O�U����B���={XhA�"OĢ��t�#dӼ;���"O}�I
5�F5����v'�Q0"O�1)�N$�����

�/�
$��"O�pËƊx�8	b�G�1��<
#"O�L鑍�(n�:ѡ�拁{�
�"OZ��eF��r��9�$��o�m��"O�Չ��Q'6`B�CZ6'%\�S�"O�xP@�)e|�q�,��3:���"O4��E�G>�X���+V���2A"Ol1 G(�3��5�f*C��<���"Oʨk5c��E �qcS)��L�v"O��0�\:$>Ai��=I����s"O4���O^7H	� ��nջ8����U"O�욥E`��X�@��-sy����"O\i�1n
�J7dP��&��L���`�"O�Q��A΂J�|���D�O�ZH�1"O���Q�@'J|�B�a�,���"O�D��f�JV|�����ꑃ�"O�L�əp�M��E,n�z�"O:hzR�~���rfG (��e"O��y�OۓQ���T! �cb"O:�@~�{�*B{�`�0q"O�Y0SL�R�2t���1I���"O��8@�3Cx�du�B�4-r�"O�A�A�Ƌn��a�'�A1e�XH��"O�|�"��%z���*Ъ$d�Y*�"O���ôj��(r���+WURaa2"O���l��0�tq�NY@� #b"ON-1�ī}�`!��cJ�u5�YD"Ob�&�ŵ��c$�D��"O��Z��%,�p�P�(u�xr�"OT�9��?A^�A@�߈4\e"O�(��1`�,�'�ˍFZÆ"O ��B�Kq�]J��پ���ӑ"O��Q��H�_������ R�^]s"Od�+�����B�,>ò��f"O�DPp(H/b+V���A\�Pd٠"O� X��a�ڥ?��� �!B.7�Xx"O����kGR�
l���:pIU"OL���:S{�Ř!�,�̜�!"O
�	�֞xD���Pz8L2W�yBi�	����f��~�������y��� 5�{���v4�X��yRd_&O@0FC<u,�V��h��'�z6oFI���(�"QIr!��'b9�E���@�'�EB���'�v�J㈎�4~�Sь�
@����
�'z8	 &�NM`	jPKP�7�|�
�'բq�cBP��ѡ�i��)n�x
�'%�(�G�2%�8ĨT�"���	�'��;�g0}"�04��E�Դ�	�'�J=YcI׶E�j��t������'}X!A�����aP�j_�颹K�'�Ԣ�M�p�$��2�ך\]Ld	�'2lyx3�Xin��+�&���0�')<��f��{,
�:�BC' �le`�'*F,AUfH�	�����,U!�'m�0G�ٶF��� ��)A�'݀�(�!�77�l�FL�`�`�+�'������
�r�����&
>����'�xڇ`]�+����U�řUl�)�'!���f���j)^�U�
�xLR�p
�'Z^�I�-J:W 
t�(ǔ}W�Q 
�'�~�U�hphГ�. 1Ti[�'HșC�i̧ �Ը��)Y�V��`�'"��q�����S-�926!#�'��-	����D0�C�h��w�4��'�4Pk�$�� �	�X��T;�'
���%`��8�
r�+@b֤P�'�2�p��ҕG�@(��E�6	����'7ў"~����� �x9��Jp�a�i�<9�O�mx��D\�^��i�oHj�<p�y���׋�Y�0���j�O�'nax"oE�I-�r��LāEl�s�<�"_-R�b@�D���b��PR%�X�<i�H�l���Q�RW�D�'�_�<�U�7E\f���ȉ(�`�6��E�'raxRJV���K̀�.F� ��
�'�V��" B��Lp����M���
�'p*  p� rb���ԉoRP�'tў"~��J�F0	2aP�(���@k�p�<�1�L�pA�D3���6��2��q�<����='��a ˥J85���V��`�?)f �H�H��@V�W�c��L�'s���ǄJ�<st

"y@�gk��Q1O��'�Q?��kO}P�a 0�Ό7�T��Op0��������s��ϵv���i�N<"�H��d'���	��J�
ĄE:����c߄.�2B�Ƀr��5�k��Xi��<&j���$aӖ�sWE�c��= $S��e���y�@��QQd�+��ةC��# @&�yB��-���8E��>�]�G�I��y�L�>b��(�#�/l�=�tߴ���O���O����/j��L�b�.P���s�'�ў"~RB̠!����� �����ԤE�<!��E�K�!��
�*������	H�	O��
�mޛ"<q�EA�h�}Z�g#�O��ɗ4Dd �d�V�_7J|෇� {!��qڐ��a��.�`�&�iX!��J�3Ĉ0q0OK(s'� ?!� �J\;A�qJ�!Qm�7>��g�� PDH�L�b�<yY�e��` V"Otp`/J� (�cM��7��y�U�$��	/L�4���
]B��;T%�3D6|��d�v}R�)��su���$pr�ST#�y�4���o������?~��>ь��Ӣ<��!���l�U���/W'!��&_\����
0��TYWMь
#�!�S�O[�`8p��@�4=(׆܂f��-`�'�0�	�.�r. �PG�Ӿ_�u

�'�a""@���i�#�lL�h�	�'K��+�7SuJ�j�H_2��䘉�D4<O0PR��)�����"}����"O|D����E\�8��HY�f�>)0"ODd�g̎�6�xth#�H�L��1�P�O;*4QaL٩e��CdA^H����'�a�!��D��#kM�:,x�'Lبe�&dp`Rc��6 ��#���~2H̝K<�郦��_6``�ӯ 7�y�@�/<�J&_�F
����<�hO7M%�~A9���81N�Pq'�c3Z�ȓ|$��P2n�b!�q�g	�/}r�=��U����|��5h�#��0XW.̟+@L�G�0D�D��c��I�0QbKN-wK��pJ.�d(�O�T�W�;wXH�X�#��G�e�!"O�|�Wm��|uP�w�K�n�r�#��$S7�0=9��Swc�8���Q;��g�@t(<��	��T����S'���'��xŖC�ɬQ�F�d��T�ʥ����O~�#>aO>�O~zw�[/;r8���Y֥Qw(m�<)�EZ�/7���@+��ya-Vi�If�'	�	�L�Ԙ������dk�l��f�n8D� ��L�� �K�g�wʴy&�3��*�hO�Ӽ>�l��.]�N�b�����v C�I7u��Pрo�Hi��߅JB�I�*J���V�;��y�4���Fb����ɝT�աB�u4�a�C��E�B�	�E	4UB6�tN�0�B�h�"<9���?�۲�M��p�gcZ�]��(H�,�O�OT4���A�:�}���K��pĨ��(�	}��9O�U1��ĖMSՎ�|wpEr1"OD��fV;(0T-ku+�,J���U"O^�H�뛋���iZlB�q���<����Ap��� �KJ2<��5!�B(I�JpBԁB�G���h���0�!�dȄ^�(m��*	5f�p�Űf��~�Y�$:g�V�t)|p�Udפ�(�jP�9�Is�����F��%`�`yi�NݞB�I)d�\�qV��
�(1�FM�Q9�B䉧S=��x�jԄP���Aj�.�hB��E�4qţO�Y��A਋�}y�B��a�!ѡ�YK�	tBdC�� �A�*��rɊtx��Ɏ+*xB�	,W�f4���'9Œ��e�]�L<:B�7F̠���osz1kT�]��B䉕]bnP2&�y��|r�Z .8B�ɳ!L��cU��,G��1�=gF��/?ɤF�35�T��׎�._>B	I4$F�<��S�Q�j���������B�<A%@U�Z��\a2	��-����%K~�<q����ám��z�r�Q�z�<�M����0Q26 &�8��wX�EyRoӡL�l�uX�$$�?�y�[/q���	a��U_9(e��yR� �)�B���b�
W���T*��y
� �K5
ګ`�2�)P�
*c�x��"O����ۨ+$U�V%K*Y�l�c�"O�hHa� 2C�\�\�\h�"��E��0=ɂ�[��1�E��횡aq�(<	�4cR^��W�
�x#j'�1c B����y��)e���y ��xlIp�-�� Ф�H�'����'��x~X�R�&"]���I��*B�%�8lZ^؞d���wl�d�KA�n�J`.�$IKy���>�I~�OY&�A���2�vTUG���6š�'�^�ea��=�ő�-��#�*��N��At����+��.<2��2��*�v�C c��h��MӰ-�y���X���#SBM�DR����y�aM1ay"�Y:G�|H�T�aҰ�8b/[��(O�������}���{�@͊Ĥτfz��P2g���H�Ɠe@p���C��A�X�Ҧ�Ѳ�hO�r�'P� �׀Dɤ�hS�#T�!�'k�����U1��	2���<	��~���%z��g�Ǿh����fM:��$��B�h1$�-~� ą<_6&����I�I��0�ݓ�hيc4�B�>�E��n��*�&Y���B�	(m���`��0��x�p�8
\�B�I�z�MZ�ˌ�:���B@fJ#�rB�ɭ�섁��N20\t�n�tgF�d<�S�Ov�41�bU
���s�R��P0Z�"O ���O	�Y�� ڪy޽��Q����	�,��Ty�:r�x"��3
B�I)nx���c�� :fQռA�B䉆T����#W
�>({��TW�C�	4!8�Ka�@�|��]��NT�E��C䉎O�lk �ڢb�`�*$Å�H�C�	3ag"�ċ
�x��V�{��B�I�0�tŸ3c�8�Jacd,Ԯqo�B�	d����aj��(�z��#�Әsk~B�ɣM<L�Al̍��P����6+pB���1��i޴��#��̵uzNB�I(c�~\����k�4`p�%V�NB䉪���	tN��T�,�ФEF�B�I
2̾�H��(.��e�dB�"-�B�	��8��F�R61���Q��ř�zB���AElìt�����RB䉴a[����,H�j�j�ˡ�T�9��C�2lQ��u��9�~�җj.^ĶC�	� �0i8MM�f���B%?o�C䉝1(�d�C��3Ub͈�A�"u��B�I�{��0���*-��d�#j�_�B��9w�R��� �RfpX�Zq����	�'^0�!�C\���yrC
5��0�	�'�Q�%<_|v��aC�)�1*	�'f�D��eQ�'��A�kg&U:�'�6���)"E�bp�7u����'����a@�\箌�FW�.��A�'s���$��G� xyf�ֲ�<]�	�'2�h"��ŐF�9@��ņex�		�'�Y:`eB�1Y (�Q�_�����'�fp���cI���W!�Qeh,��'LBH�%�����*7�Ca4��'��`�D�[���e��o�e��'.8J�� ��ɋ��5PU�M��'����7"�8M|H����_:<P�'�<��o,x�c�F�7G�湀�F�B|�)\;eM�}i�F�4�%��W*u�
�'_`���n�Lyp,��C�:�!�'Τ��a��
_^��k�L�1�	��� �Yå�
6t�����{���"O�$��eR=  hY�	�
{E�qJD"O���um��W��Rp�9Wd�"OH���/�2�����(Cj4���"OlX��e�,TD4Q�1���i{�u[4"O�0`��Nw�DI
�eU�Az���"O���tu�`�Dv}n�q�"O�ES�AZW(lš��Mg����"O�U��Ƅ�r��Y`�OY�m�l�"O���� ǕZ�\Y*1�>9����a"O��K��D:E��� R�\�K�0�y�m�+S��`R�h�R�B��V��y�c�&C$��͢b5�]�J��y�'A-�R�/��d���a��W��y2�6xd�J�%H3��v�Q7�yb�Х9v,�;W�S�V׮�jF,ȱ�y� �NHlq�b�/T�6))����y���  �qZ%AK{�pӄ�	��y�	��<V"�x4	�O\ja ��7�yB��6��<x���3n1�dS�ű�y�ʵ0p!��t�|�#�M�y�eE�~["��mA�kF�l�R��+�y�%�,���-�6ԅ�Ha���
�'T�A����%7��04+�+2��,�
�'����wl݄T	�q	
��g	<9
�'���B��˓[9��#6`��	�'=j\�3F�Y�mH4śr��-��'����Po��������t�Y��'��z�`O>8Q<A�`��
��݇ʓ%��:r�	ESl�z�NȀ~oL���U>`�Dfê�88�u'հ�� �ȓ1���↋�$^��(�^�Ą5�ȓyTtt4[�?�8�M�7`u��~�& 	��T�S�h��#ݲkU��ȓ��Qd�V-*g�́D�Cy���ȓO^� �g_�.��M����v�ȩ�ȓ!w�ɳ�d[��V��v��'~�.��ȓ 8��`'D"x�6�I���?)\ą�6����݃)�Z���I,3������yj�g�U�ʘap�T-($���%�֑�F�)3��9�`�p_�-��&�6٢���w?�� c� &��y�ȓ!Z�E8!�qBQpe��Qz%�ȓh���Vl �Z�����]l��ȓ��`E���5c��G4@�Q�ȓB�-�ʈ�n��*�ɋ�M��m�ȓq�M��͢;��٪�H %����1�L��K5-����C�?D
�$��[�gX�{~�y�c�$5��J�i�:D.rX��+�p?�&��<\X0�)`�Ȩ���1n�Kb_��xBG�03%��I�E=,T��vnѲ܈O� ;Fĕ4�`����͎*5��U�$�T9bFCE0�y��Ԭ~��x��ϝ�d�	5a��yB+�n�ȡ���\���";���-'�~P���U��C�4Z���jߚ~���aD$P=[�,�4�$̓�"y����˃-�%@��B�>�(S�@�aa~r�
�5Q \� ��*]� ��*ɜu�x<���W�/�P��{��VnT����4:$�ybT��E�'�6�Y�-ݫ���}�� ��FJ|��@��c����B�<9�E�2m�h݉�$�v1ڡ ��<�fK֟=�:�p�+7}���G5t�J'CC�A$-����`!�7:od�ʂ�a�$�"�l��S���z��U�5����xrF����=�ԩ�o���v��p?��"��;7v�Ha�P6Y b1�2�M+=���)@j�
��x
� ��q��$>�p9�Ĝ2(E\@ ��+q� ����)\4Dzd�q���j(��;@��.�!��Tk�B���.��R��&`�!���b�<�2a�&1
ܲD���!�R�GNP4��S;V2��0�g�!�5-� D
��,�$��t��f �O�h9��&븧�O�^�"N�$c r���^k0�-��'�Uz�l��ޜ$*RK6�m*v�|B��}:���yRh��4m�2�@Р�#|�B�!
�~�����!g܀hPL��u�4AQ�G�(�e��,�	���Q��Wns�:=�p�c���~���Dx¯�7�4�(��,qp��� 5�iO)n��P��tA�$(UF�-�!�d�B����B��T[�|مC�|k2�th

+���u�ɔX?n(˧��  dȜHK��.�t�PW	*D����37�8��c�yN8�sE�	(� C#��2SNK=+����ϨO&=��A���x ��NݎBLq���'���x�A�,!�&�ۈdI�-�1	%:�v�4`�/���^R؟�!�#P<bI@�Y=p��ԘK5��4v��`�!(~��]�x�O�Ҳ��,�")�Mϊ0�qb�<�Hx�8�p�����Zb�^� ��7�en�, �/ܮ$gyD��' :�	ҫ��f�u肯ޅ.�y[�'��հ�l�(}���� *�97��ǹiԔuY�Hm bGF�:�?�q�"�JѹǬ��;ɪ��G�y��,��l�x�愓a���-8��
G�O�� gȔ=Y(Eˢ�ܯq��0��Ɏs���EeS"�IS�b�+<��#<q��U:�����"�L|���E���&�ҥ��۶n�
x) (E�!�� ��ZPcV;3ޝ�P!��
$A@�ϯ0b�3������� �@S�O��.�[� �٦ ����/�.A�!��k+��C�½��!V���j���❐>><�+�b��%A��O)�Ez�%�+$PP��s���,1��8��=��/�6�С+�e�+%1���%�X�>��6�<__��GC�]�����3�ON��q.�%K�,}x6&�.Z���D*����3J��M�P�%*W�Z����cvj�3tEXY�c_S��	"O�����Va��-��cv�����t�A��]2z$���V_���D��;�tla�qبe��|f܂�"O����^���qp���=b�8*��H�}�����c��у ��6A��G�`�'��\�OW	nY�3GA1Ox�	ߓcs�)�� ���T��",D}C�5(4�y��
�FB:0���Tc3���z�h8*RC��to4�󐆓��tBcS���X�0��|��aMg�$C��* �Y(�I�N�
�aU�y��2kfh���k�y��� : �$��!�<-r��m�*�>����'Ԁ��ŏ�S�N�0fG�,h�̕��'��M#�ϳ[�&�#PW�k�b�PH�D'���k���ҁ�'�\)rrWt�Z�`@��_�L�0�3eHHOV� �(1b��;�h_*H���4e/�8����5b�RTe�7ʪ��T(�2�;Ӧ^�FP�c>YH�Aʁ �8-CpgW�n���"D�lXQ��3��)cD��I�d��ﮟ���O%���`ҕ>E������I�I�!�0i�ViD�B��$�v�{�+�n�L�@C$l�'߰�p"� N,Є�	�:�M���x�\\� ^4�p��d��f�,�6��at��*��{�*�aVC�:B&$�'���Z����@�ʥ�&+�&XhN�����T���t-�S���Y�F��|��P�Q��owB�IT�����xk�D�@�λ49�˓6�2�"�)�'~#X���BZ�:�n��L�1��ȓ?�d!��E<a�i�$�3^N��ȓ �� ��1cbH��@�B��a$D��( I�]:� F�X03oJ�#3a"D��s�N�7���* T�e�~Yqp�/D�X�UL���N!�P�X.4�X5"+D��!dMEJM�go�/"%��I,D���V�5Yl��ʜ8��1�-D�h;���2'ߠ���I&Sw���u�)D�� ��SG�U�-#0�C�S�Dt @"O����c�u�Z\@���M;~����'<iIw�EX��H�RqE�#�7⑋��1lO���=p����+2���cfg�M��MݽXSʓlO��Ie��t��y���)ђ@�/K>uJ�,Yrg)��'E�8�Cj�?k�I%>7n���Hs���`S�)ՠ�	U"`����IIf��'�a��ϣjX�:Ac�$�4���s@�,�I�P�C7%��!ԣ�K~��g�=B@���Rˮ���G�/z3Eb�1D�(�T	ܗ {̸ӧ��g������L��y��;{`<�[�O ����r��T$>7�w�HZ.�*Lij" �0𑞌���;s�$C�,	q���	��4 I�^�(С��
���qӎ����΄u4xP��uay�h�i؄��@T,�
,
��ЪA����^Ub`, �i9���#AT�@'>%"���D������ף�Vy�ցH�{���A��84�~C�5&�4�p��.+d���*f�x3�.��e\�@����Ol:İ"�ȴ%�8�P���D�	���������Rf=�j�	 � ��zR [u��b`�� ��*@(��v��<�*��$���VU�A��k��<�q�j��<�q-ԅ6�x!�5.Y�".��r�g��e��G�h�"����I-q�&� �\�Z~�	KZ�&�zpmߞ
�ڸA� S�o�!�#<�d�eH�5U���m�>8�J)���@�[�D{ I�ې�KTc�'%����;׈}�"�Q�y���c��U�-В<��5��!�\�%�8�3��֫{��IPa#��5�	���8'�`���<O�}��ڡ^p��B��Z{�Bt�v�'q�j�NZ��TX��ܥo@y�I��x��*��>��1��T�[�!��!�n9�4�@��}ZUC!i��'�mr5CR#l�V(B���M%d�P�A�,[p��2�Tyc�mN�Z�!�D-[�X��C�C�+���Z�����,T(<B��ADK1s/\��e��%?�Kǫt:"�����%V��k�!�eh<q��R	'`x��p鍙V�r�w��8, �H�Ɔ����	h��|�r]�Ó����A�:�VtRR/�"�Ʌ�I��\h�OK�y���p��;2��Q+�9.�vY �o���|Ӫ]e<	e��?1��`���(B�|�"�Z�C�v�H����V*P�C�h�k\���|�w���ą[�bҦ��}J��z�<q��[�r�y4D�n���ȏ�D���ICK��6�^�p��P���O�)����ɕ�Id0�`�"Oxy:�)�F_Vh��eQ�=?x}��W�a�Nl)d%�jV���p<�R��G��`(��˩5z���`�_���K�e��^|)0��{xl�mX�p��sH��,���S9ѡ��D�7P�a��F���0��Q"YqOHA����/ ��9��}��b?��MH�:�����4�9��(D�`9q�=\h��p&0��9���˖���Նe!�(	����|�'[�4�H�3|���S�W%[�|a�'��T��.7�R$�"T����4��ʥ�Z�Ph���1<OVxP� �8MD�cʓW'���#�'Q��"A��P)8,@��׫g����%L�^5���ʻ�y�X�~��i��>G�Z�ÀM���HO.@T?�h�V���6	r��D�D;�����"O^��\:0 ��s׀��1�	rt"O\�(�\73:��� �B��J��"O�x�7숦^{�U8cMޫItJ��"O�i�e�<z�B=�`���X�n|C"O���!��iε0�B
	�=�A"O��r��Ŏ^�2��a�#;�T��"O��*�E_#�؄�gɜm-6�"u"O����A��9�!^(�ڱ"O��@E�΀Vs�������-qB"Oȅ�cB�{A�}q*������V"O�`�'$�Cs� !7I��z@hI�$"OF9�E�0�~� ��#,L0�W"O�$�  �tL�!�V���yR&"Ob���7S~�x�Aϖl���"Of�ң�\��H<�O�����&"O<� )�(=���UN�;{�xY"On�`&W�p�԰�4�4
��q)"O�)C��+l�Āq���I�ja G"O� ڜ�O2BxVQ;��S�d���"O��Z�'��4��\K��B+v��Kd"OB�I��3ԍzr�R�Y1�HJ�)D�@��>Z�T�c	�h�iBN3D���3�?P����V�s|�c1D�l�]"hɘF,ݝ1~P�Ũ1D��Y��������C �kZ��pe1D�������;P��gZmJ�)D��R-�U�޽��!C2t� e;'&D����R�t)������{v&$D�8��ᐷD��4kw�*B�(��
&D�L��e�pAJ�J��;C�����2D������n c�Ή(#$9a��2D�l����y��y�&�V�Lբ��0D��ۑ	���Y9��_P�j,D�<�&.�#�ڈ딧UD*��K+D�����ݐ$P��Y��
e�p	1TB&D��pJ�q�V���BS�
�X���$D���JR�V�Q��!E��XQ M.D�� 1hS-f�:��G��(Nq̜�W�,D���%��E�^(��Ѵ7<@��#O&D�Tx� Z�4��)���"P��;D�܁ơ]$`2l��3	ɡ"����Uc7D��	��H�x4s�EGl��h� 4D��0�-O�E��}pdH�*:1��5D�ǈ�U�N�A���(�����7D� An�#_C^X�犅CL���p�2D��	D)L�?W2�x�(à<��P���$D��#1a�[8a0A��AՀh �h?D���J^W��L��枔s-vr;D��Z%��,<k�� �\�Ht��SG*D�<ң'�,.���Ђ^�$�&���,/D�0`n�V�u�ٶg��XXW�.D���3jÛg|!�� c�|ps/D�\�`�U�GW  �kB3:@��p�)D��5� ��@ ��|%���`i'D�4�5N�	�&tk3�Y��X@�&D��i�,�:�bL�)�h��|�&D�|3Є�| ��#���]|���,1D�|� ��9Hr���
	+� ����#D�Pp��>VS�t!�d��c|Z�Q�:D�̘�d�1D�$ bVl֏�n-҃@*D�$���͛B����o��s�B혷,=D�x��EO�9�N�8��v���b�%/D�����Yf���>B�2���!D����_&6<�L*�##z��aȆ�3D�t�����|`g"΍,ن�PR
-D�0��H���x�HU�[o\A�cB(D����Z2!�z��T#D~Jc�#D���P�ݫ�⠪�o�9k�"�`�!D���a,�3�xt�2�R+=�x�"��?D�$ Sf�-I��li�h§iK*�Y�8�Q�Nђ\�ϓx�IR I�Pk��#�A;X�����$��g����(��M=A�PY�ʚ 1�>���/�v�+� �[�=)���r�X�F|�咏u���2KTcܧgYh�2֍֯Y�N1��c���6��ȓNF6Ei&.� F�sœ�oB�5ϓg�.-0 !�>tT8ӧ���zg�A&c����B������"O$���C�B��ђ�mȲ:���k�����Uړcy6����'{��X��BV�LU�o� F��`z�JW>�[���;z�8ೡ�^�%$��!I 8ɡ��z��9�,\!�Fd�6���ZW���3O߀4�����iY�x0���A��p�^�`E!nN!�D��q�����"\��pX&W�d �d���(	������)�g�? JM�1�1~�����������"O<��BM�\(|�`#$	�@)Ó��� ����%ҕB��'P�����O��Tqa
B+iˮ� �+6�U�'�ڍL���ʞ�rA���z�Հ	�'���9&�<��L��L*QA��O1(������i �d��5A"7�����#�y�ʞ1؀�R�i�_��B"��y2e��x���)�F��g�p	����y��P.4,�@^+ ��3�ʅ8�y� �xA4�K8[�QbԄӱ��q�����i�"r.�M���
`�s���_!���rb��9�@�9�|�5% �@:n�O�t�e�@�B81�1O4U�taΦb�p�y��D�_�����'lt	��
L�8A�ȎSC(��mB�(2JdR&	�<-���!%�'�T����SѦ$Z#A�+;�B�@������U8+��e	��j�S�X�0!hr�J3�ʠRIY�0rjB�	�訵C��ل�\�"D���Z��n����Y�p�Ȗ*H��+p�%�g?�@$~آ��A��r���4IV\�<qG�\:7ƙ�%�W�������_�u�̭S�a;Yxn� �M�
���3���������G����*(|Oz0Y���]���X�䊀%E����'�t��E�Ж88�a���?ᕩ� ��l�w儖]n�٥$�v�6���6�ҥ8��p��.��������\hѪ�z�䄯���"O�;��)-v� �EF�Y^p��ϺF����'�	A]j����N�>�I��Q�Gɰ
+�d:��"�VB�	�R�N������v����	�j�$nZ)R�j4(pn�{4 ����O�di��]�� Dk�-ݠM٘H6�'����mI�g��`y��:9��1��[�^�����>�D���i�r�a~�,%��R�1X��w�f������LPՖ���c�O���COJ2�ʧa�na+���c�d$��ꝿb�J��ȓȰ� ���V�nP��y��-(�̋�a��qE� tPm��ڃ�Q>)̻9� �1���<3m��� ̛R�p��%�z�� �1!H�u��Ǖ ��R��	��8C"��&{\a!@`��?��`�	�^��!�W�"¤IY�懶Ǵ���&afX�ѬK�_��]9�$�1m Z�����Uk\��@�@FZ)��B��ΰ>i���{1�A�7�sn��E��g��q��Q�$@��.�f@�V��D�� 0�˾~zA��[��sB!_(�ƙ;C#�E�<!��٬�0 *���2�䙺V
��pȈ��1N�! -�#��m���	��ټ�Q`J�B���
��?X܀тE
y�<q7�U�dX&�����%&��1�
r)H�I�e�l��DB�����`��ӛf^��H���3��P A�S	r�c�*|O8�!� 9��@����,+gE��*=S�@ ��\���f��>�(4��3Zdh��2�)e�ѰD�"Ex�(\% c���b�P�Qa�j��`���9b�j�T� A���#nԎs�@B�I�&C�����Y��nq$a� gZ�`䉮[�Mc�	V�EBbF�%����VgXh�e#�
���/!D�����܆r�F��CC�_�:d�E�!}b���]� 
C�����Nՠq�!�,i�:�O^ԋ�bC?Mb� q��ӯpӖ�"'LJ�-�����H�x���j�s�ǅ;%W��{�oW4��O�$����8avR�C��di�ɴu�N���X��!cD��y�bK ?"����վb\hy�#[��~2��&2��@��KS��EAr,��Eoe�AJ"��,NC�ɼ5��`�`�
^��Bv��l�'�|q%�65*І�ɒ@�peâ�W�gz���d+d#��$YDMu�����LRpiC��ǆlp���MЍ!�`���'�4U
 `�g�� ZF��E><����� J)��'0��{7�3�F�l����T!LB�	�%h��� bF"a�r����K�L����ڥ*$�)�'2u�}��������w�˼A�Э��m�FL�g�٘Z�~0r�nA?�n��ȓ�4����چ��IŅ#��C�Ɇ3Ä��K��
�6� N�;��B�U��H8p���E�:%�#r��B�)� ��@0G�}^ ڱnY��(H�"O*%Xf���h�A�n��8��M��"O�	Fʀ&%��$�M�c#�I�4"Oz1�BB��5ꈹ+c�ժ,yD��"O�����8&&��p�,{V���"O(ywMO.?lX	wlL;A�%jg�'������QX������Pp1��%U�� 9��#lO4���&E�	�DB�-��&Q'j����Dۮ�e�L��!"F�f�yrGZ�~Ȕ�p���;�,)z�Z���'��0͚�8�6�'>7�hӨȩ�I�� ��4���12J����oC�cf |�'�`�l�<Sr8��"o	x1��J�"�j�#M�,1da�.E'���Ǫ�g~R(b��
���!d,r!,I�p����=D����$ϞjT�y��|�|����+ZN��6E��Kh���O����8J0��$>7���3�|�uʐ�!��{�FI!��zB�H,� �"(��<�A��`���J;`�Y�P�l}� �Y�-뗍��<����;7�4pt`�;x$ℳv�d�t�qۀ�Sn��搋�ᝦ<���K�6+? 9Fj�1z��r�'K�!�$NJ����@��M)~��0>|���~	�ax�Y���3� $���;����@Oφ<��t��B��j�� ��[���(��/9� �[�n�[!�!�emN�zv�c.�|̓y~�#NB|�'�`�����$x���[�B��7`���<~O\�Y1�FL?�q�28����	
=N=N�y��]f�<�!Z�;����%�9u�|}!�Y�/^3�"���u�A�Ӱ$�Q�$���]�6qY"h�	�����o!2=�ȓ[vpj�ᔏ|ݜ�0͒z;xQ�ȓ�(Ԫ1͎Fz@��\)F�^͇ȓI~`m��D[��h=bD�ˢ@��=��;jj��D@Դӎ����#zBЕ��y-��d֞U�JC`טxl$���R;�l���� t��)c��?	AD5�ȓ?(`�1�(­y��:�E�4x�p��ȓK�>�	�#��i�Lh��gD35_Du�ȓ-0� Z0M!T�L��0���T>�ʓ��Qb�ݞi�T����l*�B�*3�LA���QƬ`��S&sj@B�ɓI���-�
y��٥ �<a4B�	�?ת<�2bݺ#0�ͺ6�$a��C�IlKD�@�K'޵kt�>x��B�,g=�iBv��X����Ɵ0-�`B�I�W)�RL��Y�J�E]
c@B�I
	�>q�'�J�n:"]K'.۫2�ZB�	�x�r�X'/��9DV�8B��T�s���~A4 p�hT�	52C�Ik6P�5KR��%n�:N�C�
V*)Hro�f� �e�VVB�	/��m�mО7�#)�(t�PC�2y��� d2"�� iGEMcj@B�I1r��Ju�ޒLhz�q�I�M�C�#uS��e�B�u| @��x��B�IU���Z��ծ2�$��Ү-.�B�	�j,9*�M��T�p�KC�tR�B�9" Ze�̬zRLt��ˣ^bBC�Ƀk�xM"��8�X�,D��I�a7D�;ٲ!7�Tز��=P՞	�J2D�(��L�j�J���K�|�D���2D�l�ql(�6���o�/G[^��S�7D�l!-ɽ{I����J�>�P�J3D�́�"!G�*S�˦R��z��.D��S��T�5S��p%�6 �"�2�e)D�ԣG���,1��1��Y*ͻ�'D��r'D���p�ʄO^3CRd��.D���1��9&D��0
\�r)n(��G,D���fIL'�U�e�]�yE��B6I-D�� �l����z	Kr��wPZ|zP"O�X׫�!��D�֋��:��}�"OP�
Qʉ�H޺�񇉛&�&p�@"Oμ�!g�(X5���QF��F�Y �"O�l
�'؊;�.@�b CZ���'"�M����8C`,���oj�qv&��G��q2�'&* sL�*J�DJu�
�b`���'�\�+�`��!	Dr���!%�r��'�Lu1gX<�	�0���&D���'ǖ�b�)-2a30�B�Y�؀�'p2|X��N���ht��Dg����'�X����H*n�ṃ�խmn���'�p�x�ӇZ2A[��ݓ��`��'!Pp�A�Ro�|�AA� X6�!�'��e�2��mЁ��ں�zMH�'��5����-�\DHb���^�p@�'�\ӴdͯN���A�eH�]@���'�M�j�O't�{�͓2U��9��'~����I��޼`�f�� 9w�ِ�'�b�Q�o�_��@F�1\�.��yR�_�\�,��=�|b�.�~|�Q�-�iɔ��"�l~���Ґ-�I>��ɐ=KL���@�G��� [2���D�[�usT[�D:t/�O>7-H�B 8��nފ�U87I�*Lw��`H�'���S1C@<
�$Z����@̧ngJ�Y�K�3��2-I�\��f��%�=3�oӤ��+��O҉OL�U�m,<C�V�61\là��a�\�l`��0�O��Ŋ��PW0(�QÇ�a���b/<?���O�^ª	`��/��ͣ�@3#��9hLi�ԋ���əy��IsjS$^��S�O��%�����<ո�)c�Q�i~j<�4$Tqۇ�Z�8d.8�ȟ䍰�ň�t2�%�r%�#�9�Ac��K_�̗'����FM>�"UIؗ��4*�%D^�4�iЪ���� lz��Ї+�0|r���=W�L@T��W7�p��H�<�1�Z�V"���@X�:�6�
�\O�<����g���d*�Kd����I�<yw�`�i�r`��B{�z�F�_�<����$nT681�^�bWl9��R�<�5�S�W�t�[B-˹x��qJG�_Q�<鲫�I�4�WJְF��{���r�<�q,�T�p��EF�,@ ��@�Rc�<�ț&a�0�Hv��5�=i�Z�<YOV-C��ň3K��B�˔[�<�T,G�WDɺ�K�@��iFZ�<Ia탇vD��"��5�ƕ��W�<y��-ê���OB#��Yx�m�U�<Q�C�*+d��1��!-��A��M�<i���Wk^��0F�}�%�k�H�<q��A�L�����푨��6�A�<a�C��n ����-�A��y�<ѡJ�%����D��`�0�Ф�y�<�r��c�i��B+n��А0��<�����F���k�㏧L���	S`�<y��Z�$M�={!�����D�_�<�ů̳.|��r��!.ξæÐX�<	A�C5Y��  ��q�v�˓L*D�D�#h7c� (h�䉈v(ݓ�d3D���ՁL��)�+�a�  Q�,D����@�a�S$&����&D���N87�l#��#S�$[�:D�`�s�٘���@��,7�����;D�DaQJÅygZj��&��qGk:D�0A�U.2���N30o4uE�3D�0��V�����I�bi�S-1D���-�86�V<�sD�6�0���*D�Pp��؍n��䆃��@�q�(D�<��+�F�x�S��4/�l��&D�� �x�Q%����J��mb֘ʰ"Onѓ1�?��A��)
%�ܲ�"O��a�M��QK	� *�d4�`"O�y;R+�ic،�j�#��U	D"O�(�#F�� ���K'	B��ۡ"OԀ����#i�D�6-D *.��6"O�Q��DN����I0��*��"O�{&��8Y�d����_@�|G"Ox�CR�
�%Z���'>�5�"O�� ���O��03����٦"O8IS����E�$0����6�ڹ��"O	���0;
��vI�9GFF���"O�5�,^�2W�Y�3��*.�"O�x�2�=���I	!�́c"O��y�C�>�򠺆�9����"O���ք3$�JQAf����"O��Iek�>.���%&	�`�F��"OX�� h�&�ֆ�+'�vEZF"Od����&�>��a�l�d=�"OxM���ҙAt����S��)�V"OP��!�M)3�6��!ć!h��Z�"O\Ara(�/`,h��Xs�(t�"O�Axc#����41�E�r�yp�"O��H�`�#uT4�%�s`8 V"O�9�����P0�Y�r�I�@G���e"O2ppԣPG0�Z(Ɠ0?\ �"O&y�S�z���5$\52(�9�"Opx�r剿p'��
sB�WC��"6"O�����_G,˵�O#>Ej��v"O��0K^4x�B�2� ��c��P!"O����ч���˒A  c�2Ԡu"ON��i�:s)&��&���yP"ON��T.ޮ]�z�y�e4b����5"O|	ңG!W|��Ę#=�.]c"O@ey�ǂ~H@��Ӣ�'�!C�'��h�a)�L8���5��lZ�'P$S$I�#�����!�9e�XP#�'�l����r���dά��	�'�ly����档��J�U���2�'�6q�r��}|ꐈ5�B(dJ��q�'�&(�S!BS>�s�7�B�'�p�1p�z���/R3y���0�'[�%�DkЬ#x��$�n�*š�'C�(�6��o���ALW��y��'<�d�P��2�%`�#.�'d\LG�>�A��A�)&=*h)�'Z�S�� gy�������h�
�'(^D27���DP�E+!���	�'9ZP�dm\�Y�����"�	E8݆�&z�	j��\()C �M3fU��Ud�(�SLp ��T-�(m_�Ԇ�jh��ʐ*��4� E��F&N삕��v��i3�*�z���[�%�LE"��ȓFG�����/�����h�
����K����.nf�<;T�I�i0 �ȓk��B� *�}��_*LJ8Ņ�_�H�̒�O)ab�A��.�0��ȓ	�x���͆,}��0"�aF�<ˌ��&]�0���2ҮѱsdP+sڞ`�ȓQ�Y!L�<P�����Ѫjz���ȓa����o�7��Q9���3_�d��<���'_��-a`�D
k�j��<�^;��_L ؠT�G�CJ1��Hu�Xp��*n�:pxs��)Tx��S�? �x�!\0\A:ƪB&���""O�$����X��I/��.h��H�"Ob0r��5?��pz�m΍:Vɧ*O����UG�Y�!
<B�E��'��Y���^.]� (%�#�N���'<�p���*H��е�=t~x�'�b�hRFL,hu�� �,ʜ��'����F��U�M���Ny�����'�x�qOGX%��ŭ��i ��8�'D�x*A�wB���4��]���'"0�ұ��9���@�n��e�l	�'���ʰk�q�ހ3�MB��<��'o�%�7Z�?�(�fE w�`��'��q�e(!3�D���쐩a�$#	�'$���6~��[f�
�J�XL��'
^�hё*I&�C��E
t��'z�
��3t��Q&��)f]X�'�:-��O?Š`{��V�3��%k�'��5bG��)�@i���%!HN� �'����NmT��DCM' ׼)�
�'��܋���)2|:I�u�e�

�'[���Di$�|2�h� p��	�'0��$b�M�L��S�b��'(�u�˞m��Q����J�b(x�'2�S��ހ-)���Ё�����'V钤�֎]^+cLH�:�и
�'�0��!h�F�6�5��?����
�'��˗�&����d��5"��x
�'o����T4_и������t��'Ȇ��v��&;ܜE:��Dm�����'�ؚ�	�%wg���`�3_S�l�'�����l�?)�4���oљ $>=*	�'�P�ВeUp��_��qO���y��T�_�@�s�Ԉ!�t�!ԃ�3�y�d��D�`@1b�){�M�TGV��y�m����@Hg�nr�Q����yB�U��y�ːG<���Į�yB��	ZB�2�)F��N�h�	H �yB�՞F@���Եs�`I;�y"+�"�����aK�nb$0���y�"����u���Ղ�+C��yrHE;�l�͝=�(��ER��y���@�2�� ���>㴨�y���^H���l��q$n�2�y�.6����n֘b�T��� Ì�y�O]�i���Цͻ\�4Zr)���y"�E)JH,1�P-�ZG^	"�	?�y�k�2��p�d&=��)�&π�y��P>R�B���&�8C	`��m]�yr/6=ߊQaog�B��f��yW�Z�>ys��>p�� ��H�yR/��|����Bl���;�΂�y",�*�N���"Vhk��Be���y2�X�� Y5�+^��Q�f��y��p%"�ـL�0]�@�C�'�y�Q������3'8�i��B��y`��Y�ȋ�/T�$[*��y2�Z&Q��k��4F8���Ώ�y2i�#S��q�g
�˅L.�
�{�'LNY��
s~H�!�_�,��)��'h�$F�(�X0��H,�f+�'�Jaj�N^�P2��[�hA 
�Y
�'F�Q˵M�d��פ�MnD��'�J��$�'yJ�J7�D>��QA��� ����)*��l;���#!���"O�d�å�_PhS��� z8 3"Ov��$��o'Z��w�Dt9��k&"OfI�*F3s�����y �a��"O�3!Nǩ�Π�����X�b|c"Oqxt�=��!Ӧ�?\m���"O>5KE���S���7��`e���7"ON��0j�*S���
 �ݝ\4�+�"O�̙�D��|�Xȑ%9K�tK"O�񊄮�%���sDN�D9I��"O������^�k��<7^�j�"O:U� ��� �bhC�	"Nx"�"O��b�G��%���  �q�}�"Oz�鳍�[����nŎbT�҆"O�ۄm�R�Ƥ�D�U>t�"O(�H��ظAZ�Ks����a�0 D�p�#ަDe�q#7��u�0L@��#D��00��%��lڤ� ����!D���u�T!0��a���|��U`�O?D�$Qo�@�ʍ�vپtoZ`���<D�@� �	~����'�X�8(���A=D�8�r$J�.e(Y�!�x�21K�<D�<9�)��+M*�TPC���8D�80�!ν,&��g�tϘ�B��4D�@���>~܂9�v�:p]Vp�4D���f�ݠ5@nD��)!'$��-3D���C� r�Z���#~����<D�\P�%L�ryN��mN�) b��1�7D���6Ȉ�Dt�d���*4v"M��;D�<	E�#*x�=ї�V�^E���,D�H�� ��|��D�  ��g�8(��%>D�@	��D?Cv��#�
�\Y���&D�����A2/>Å$[10#�I�dn&D�$��]�;��7�ć_�p�!D�l[��   ��   �  N  �  �  *  H5  �@  L  �W  �b  on  �y  ?�  ɉ  ,�  [�  ��  �  0�  t�  ź  L�  ��   �  ��  �  u�  ��  �  H�  ��  , � 8 2 � �% �, 4 4< �C �I >P JT  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(՘xb�'��O��(⃯"T�����Y3s��eX@"O�-Q3�&&���PFi�&��{W"Oݪo�����XsmF%b�N1��"O�����?l-�pp����k�j�w�"4�L���%U�\�5�Շ<`u!r�!D�����7D=b}�����z@Bm���:D�878B�lq�ɣ%�6o�!��޴%��q���T�D��=��@خ�!�ā%"�na���̥a�A�Ve#�!�X%0��I�3bZ�8u [�6V��}B��ȹ�V��T�S�&����pb:D��1�)\��j�;�lֱx�v���A$�B��?���ӽmTm����X�P���!D�Rl��A�65I�`^0�P,�bƪ>�������B��a�B 	�+��B�	�x���s��q�i�5@T%,BB�)� �}�Q/nI��x2�ݡ ��B��'��'��P��:Ar ��b�-7�\P
�'+(qh���NEV���럢^ti�'?�<�̚
<��$��+F��l	�'� ���J/&���*Ł�1�T�i a%�S��?�«D�5`L�����+Z�d�{�<� �׷,0��0��i ��#�AN�<���׵Y0$�o�a4:�Gtx��Fx�#���I2
�+�`��c�щ�y� :8�8� $ݧ
�z�2#��1�y�n�5"�T�e�ʄ�ba2أ�y�'�BH]��M�>/� ���yr�&^}�M�4�$m��{F���yr+��9=�㭍;kw�rJ�s�!�Ĕ�>Hr���FЉKg��*�DK�!������	*8�r��`+ �!�$��U�@ᆖ�<ڰ�um�r|!��� �4�r�I88�N�-^4F�!��Wdf�H�/ƶ����l��#!�$�*�L%��dԁzh2�¥�t!�ߺW�Y  %�ox(���=2Q!�dϞMj'螁(n�|8��):!��]���l�7�ӏ4��WM߰!��ٛD�6���V� ��*��
�!�ÁOn�X��U�v�����B\)g�!����)�"��i���V�!�d�>H�0XQ#��j��9��OU%I�!�GX�b����ڬm����W�/x�!�^a�@plTR��6ޞ�� "O ��0�	��D�a��Ա>r��W"O�t�3'P,s겱�aIA"��]�""O��A�`�7 R(iUOL5p��!�P"OF���H�<p�1�ED(G��q�2"O"p0"��I�B� C$���3c"O�<I׮�f������9#L�6"OlŢ4e�!"�`K0MS
K0�Y�"O^ Ct�Wk�LۧkS�Jwl�xF"OF0���S5C=�(��oO���"O�����U�L����?>8��"O�����p�<	
%��i6�X�"OxxVD��xt4ahƈ��qs"O64�ǆ�JW*<2Ӧ��]ߚ��"O�m���)Gp�P���o򠹘g"O:4Zg�&<�����
)l���"O��h��O0(|�1aԎR�P1
P"O,�%���r�jƟEY����"Ot@��@� �XR��6K��b�"O<���cU
�^ �1o�?q3���"O�Q$��
W�Q��n۷
�8�`�"O�TD�� ��U�r�3ŚhX�"Oh4�c	 l�Ƽ�k�!��ѐD"Oyx�3���;G`�F@8�;�"O2�q4��7�nb������1"O�	���8~�Ȁ9&-��4��L� "O�����9G0:PA%:��(�"O���Մ_�x�Z� DA��b����g"O�Z�k	a�l���ӼF���*6"O�J���;hfB�!/ݯ6%J�A"O&M)v�1X����͐;��"Od�b@���?@����R��@�'"O����(p�hF�V�6��g"O����)B�a�F擌���"O"��C�čC��}ل�ע_�,��t"O�q�aaW�{�������$���"O� �EQ��šV4���ɪ�l�SU"O�Dr%�8�*ȫE�7%��Ȳ�"O� Yg
W���H��L�8 "O�k��=YYxDC͜&�4���"O���/_���쩀�!$����'zr�'Y�'F��'�B�'���'t*�y��Ջ6��Y	A��{Ĕ����'Z��'��'(��'"��'�R�'T�A���I�6|p\q�+� Q���E�'��'�B�'���'J��'[��'�l�0ҡM3���y ���Vڨ���'��'I2�';r�'�B�'\b�'����ܮcM��:�eQ~�)���'��'%��'�r�';��'t�'��%�T.W/Al�Z֢�&��¶�'���'6��'���'W��'�'�� ��g���Pd���h%�d:��'E2�'��'��'��'/B�'Kؠ����Z=�U��V�R<�a�'�'���'��'+��'CB�'�X,W��������Z=p��)�?���?y���?1���?����?!���?3�ۡW�A�%R:S�TqZI� ���O��$�O����Of���O���O�׀(�x��Ӆ�2@'���6/�z�H�d�Ob�d�O8�d�O�D�O��d�O\���ư���޿?g����D!^;����O��D�O>�$�O��D�O���O��$Y8�H�ŝ�.����8'�d�O&�d�O����O���O�mǟ�I�.��Q���T:]+�,��k�N��*Ov�D�<�|�'l�7���pm����lʉg�f]#PC����Ŗ�L�޴�����'��aԘa�z��4̀�U��P����$O\��'t��K�i��I�|*0�OU�'N�"\�g��:�����F�(+5���<������>ڧ���hWC:o8�d��@"m�y#�i�2A�yB�I���]7r��-ٌ���h͡xlhu�I؟�̓���I{C*7m~�ȹG�ׯ`�6�8G�U�U/f`���a���s��bFf���4�'�a�d16�@m���-h�
�'w�	B��MK��d�n����G|T	Zc�F!R���m�>����?�')�I�O� �,aRҤJ��!0��?�7ɞ�J> |�|�'��O"|���%�@�N@�0��y�Dρ0�R*O���?E��'�����*X���,� j��es�'��6�&?���Mی�O,L!���
i������*^%ز�'���'��P�8�&��Χ��������8h���dh:��_�r��&�����'���'��'V�qQ�@0Z0Je�7��0&Ҩ��R�'9��9S��j�'`R�'δ�T>�I�[�Q� �4x-{`
۶V�fd�-O��`Ӻc��I���$�U�T���_�A����h,=X<Q���q����
?���R�e�'9���]���,��	+������A e�3ʔ?+��I����Iڟ$�i>5�'XV6-� # ����N�S6��4�@���IW�V��dI����?Y�^����4}�&�'�\�+�ǆ�(yB�����F��=�����n�f��<�6K�W��d�~zT��2�*ft���ЙOfJ��@&�/g�d�Ol�d�O0���O�$6���Hpj F�`�tq����Yͪ��I某���?���Ky� d�ؒO�`���B�(��$sH���Wb)�妵���|j�0�Mk�O�``��+��Bo���s��
�J�V$��+�t�)ћ�R����	Ɵ0Vjj0:��R�i`�	��ޟ`��oy�e�O� ���'���'o��7 �A�C�O�D����&>`�R��	��Mc��i�ɧ�	��~��0�/��zNer7Mݕeh	r�R���X	��>^w��d�I�/��i��Z�P�p+�Y!�f�25�fɺm矨�IޟH�I�b>��'��6-��%�-�s,R���e`�y�m1!��<y'�i-�O��'a�6m˵tB�Ó�șn�P��o��]�Mo�ɟ�X�BP���'#�ˢ�L�?ݦ���q嬂4�P�R���H�&Qs�o�ۦY�'���'���'��'���gb��s��#�U����:�$��2Қ��	ğ`��\�s�������$��C��Pa	�|�z�"բɉN�i,1O�O*����i`�d�=p5y�a�++��,I *ƳJ"��!s�Zy�IQ0�I"�M[-O�I�O :��}�B��k�R�,�{"��O����O��<9�i.�����'���'8p��í�*~X�麦���3�LP���K}�i�0YoG�I	Rۈ����$�>��w	ӛM�B�K |��̊1:�@��O�]�e^B�ɟ��E��2!Z1�a� � �w�������(��̟hF�D�'�޽y`�Y�l��=`%$����_�?qC�i��iT�x)ߴ���yg���pDaϪ{F��{'��~��'~��'k��(��iH�	�m@��A�OP�6Jƞ}�H��[Vj�	��Leybn����|R��?���?)��EI`��2f�?cO��+G*r�tɃ-O�Ul��TP����@�Is�s���v��*��1o�8���W��$�̦��ٴ��ŞN=b4���U�O_\u�0O�e�80�Z�&�pI�Oh�r�#������Y�8��4���	>

�8V�O41_���f���	La|��e��Ԉ�D�O��AW�<��$X��z��5=O�=l�F�� �I�t��������@;q]>9넁I01=�%�Wצ�mv~��\��5�'��ܿ� �U�ē�;/<���A����@:O>��D�	 یhqB."(�V�2R��ʓ�?i�'u�M�O(d7�4���2�IfNñkp���WI(t�%'������S�K��9n�M~oY�cV&a�,�nR�CK�&}vLI3���T�Q�|RW����䟔��ԟ�[t��58i"�"��ҍb�'����	cy"�j�8�27O�D�OV˧~	��X��$e�k�@�9x���'���iy��a�@e%��d*����k]�0��� ��s��s�"P9ZM���'kA~�O��L�	;�'�.�ك&�3'O���GY�.:8a�'Sb�'|B�OG剿�M#G%��%��F�UF�ڼ��ܨ�K*O�n�M�@��	��Mf��!q@�.�؀1vŊ-u����4p��:A���h�É��M��4�~¤eԈC*�	��J/O��@���<�/O>�D�O~��O����O�˧j��I3�H���j�'	5HmИ#��i��9�1�'n��'���y�l����<t�S`�˸y��� b+�>w�%m���M��x�����|3��8O�1Z�
7�L@�g��b�إ�U>OڠЦJ� �?��=��<ͧ�?� o�o��pF*V�
�H�8���?����?������u�w�LMy��'�)�Ǉ�^�pi82Eތ������'|�'g���?�ݴ-��'r@h�@@��5J<xn�+��(Q�'+2�Į�\��P	�����쟒�x�%m��DZ�|R@���A���Y��Q�{f�$�OP�$�OT��!�'�?�b)��tl��f(۟G�,��	^�?�i��}��X����4���y�%K�s�k@ˠr� {w��
�V�	��Mu�i��7��e,�64?Q�n���)�9*Q2iX#���p�#���75d�ūJ>,O�I�O�$�O����O=�P��)���E�@�Y�����@�<��i��ŻV_�p�IS��xqU��oDv�� C�z�6T��/��$�O���:����F�>Ia� �
�ՉB���Jw�L��'GX��-�e?II>�.O���P��.?��y�"�Q�[�聚U��Of���O��d�O�)�<���i���#��'���{���w^���&片9CЈh��'�7�+�	<��D�O����OزeZ�y�H
$l۱.`@�$���7�'?������L���)@ J++4ʌ�+��@�����w������@�	Пp�I����z�o_�2	�8��K��=6!7l���?1��?B�i$*�Z�Og��vӔ�O��
�����I(_16D��D�=�$�O�4���-tӎ�Ӻ{���!j���i`h:�q�qMY=%��'��'�����|�I��D��(M�6x��K�a���P��8n��@�I���'�7�AL���OJ�D�|z+Z1 -E��b߷'�(�A�ŗU~�>A���?H>�O�.1Ac�(H�K�,�*1�8 ��(�L��i���|"u"��4'�� v�z�:A,�^�W���S_@���ݟ,�	�x�)�Smy�As�TY��`D�xDH���vTR��]0yN���O�XmO��P\��۟Ċ�adU�Ux��6y��i���R̟l�I*3�o�a~Zw;�ip�՟$˓Cgt�ڗaХh�ℊƁ���͓���O�d�O����O��|Rrc��Z͚�`R��$|�(qX3��=m��e�H��'b2����'��6=P��͊��ˇ(:m�d9��O��0��i/v�6-c�<�ヌ.q^�p�P4^��
ak�4��ᕋG��<�D�<	���?9�e^4���*�憢b!d��U��9�?Q��?����d�����Ug�����ޟ��0d��Ak.�3�"N�`�bb�D�{�2���ɟ(��J�ɴK��űC��2��#w�Q�6�0��'�� ��GQLF�6f3�)΢�~"�'פ�hvC�8"���)݇AjЉ1��'"�'�r�'��>��:2���e?�����D٢
�P,����M�Mѓ���ߦ��?ͻS-��2�'"oV������\�q̓�?!���?)���M#�O�}0alB�7,�<Rfѱ��Ş��P��^7��O���|"���?����?��8;��������R	S&S�8 S+O�nc�0��'B����'<�!j�M��<М��á��=p8�Jŭ�<i��M��|J~�2[�xs,��A���YNޑ!#�G��1�6G j~F8�.9��T<�'��ɓE;:��I��'K���&N�
��Ğ�����ҟ� J��v�@�� /uм:��n�8ߴ��'����?9���'��n��K�J,|ݸW)� //P�Rs�i��ɥhF���ҟN����� [�b�6��*0����	?\��O��O����O���9�|�&���(/� u���X���!�'��byӲY��=�����mK��S�,��+(>u �ؠ!�T� M>1���Mϧ�N�ܴ�����7
� �P/ё)ĀQ�Ǚ?qK.1�`�?�Bl1���<Q���?)���?IfƋ�?dL@$�Fqq���׾�?a���HѦj��˟h����ȕO& �ӷ'��g�d�rwOG�T����O��'�b�'ɧ��Z:T�u"�0m�>�%�Ok���!AeΚ&�~�Ɲ��5H���g�I�	��z��:��J�~�J�з�'���'�"���O��	��M+���2��C�~$$��U�^u�ux���?���i<�O��'=���34�8���p���U#�6�h7��ަ� VA����'0���k�?9��W�� f<R0V0	VY�#J9m��	��>Oh��?����?I���?i����iE�18(3�'0(~5 ��/<94�m5	�`��'l����'�j7=����PՐ�
�V��$�O�d9��ӽ/�v6�n�p�]�+嶨��@�/C"��ݕE[�u��'��'��I� �	�~��g/�+6�ؐ���D�$���쟠��ʟX�'�@7E :}\���O��ѱG���")(Ʋe�2�ֻ\�X)�O��O��O�\���E�F�Bػak�a��"������֤~� mZ���'L����ޟ(�p�N
	�5�îճX���ө�埈�	���IޟG���'���� *�}6`��熠
.$i ��'�7�3v����O��o�d�Ӽ��삌?u,E���- ��ʄ�<���?�'v�9ߴ����:���N�?�9��]�PP���u����T�@M�]yB�'���'j��'(��1a���q� �(z�(���e��	��M;6_�?���?!H~Γ`B�+��5+	~D�V-ЀH_��
�T�X�	�H&�b>��Ǥ�\cv�3���9z�+�⟴B�R�l��D_� ����'��'��ɸ����Q _$��$A�D߱$*��	ٟ��	՟4�i>��'e�7��'4����XH���'��˲�Hw`�Dq���@⦹�?!7X�d��ҟ��:��,ѡ��}�����B; �rH��oOߦI�'�A��{�K~B�;��ۇ�
<�a ���7�2,��?���?����?!����O8­�	=o>��0��D"����S���I��Mk�$�_��M�֓O�̒�$C2�V���!�#)):���l�	㟴lz>�е�e�'@f9{H̱+���0BKŁ�@,�����<�	
#��'��i>��Iן����e��9���-��)1��gA���I��<�'*7��L���O��$�|*S�Ce�L��ǫT$�r1��R~���>��i�H6-j�)�5�j�xSs��0\��RI2 p�	�,Q�׊�����(,��Q�I |�@kfmӏ�"�	WI�b������4�Iڟ��)�Wyo�ܼ(1P�<2����J�: �R 
��I�M;��O�>�&�i2ļ1�gʟ��#3�p9�)�''l��HmZ�)�hl�i~G�
6���T���>��Y��ZK���Eb��o���<y���?���?����?�-������9�4͠`���K�^i�r��Ϧ��3$u�X���%?���M�;b�Q�mV<-Vd�
�7:�ҩ ��i��7mK�)�ӽ>��9mZ�<q5*It�$[�A�'}��B^�<yG�20���ϰ����4���� �Z\�RdՋ#�~̀�!X���D�O$��O�ʓ�f��y��'eBaęV<f$�0A:u��l:R)ޜ9�O���'�d6m����K<y�qS��s�a��Y��@��F~�bçm^��1ŉ&��Ou�%�I%.n2,�6ag�Ѹ��lc�p�qV����'>��'����L�FH�S����J�@��)uk�֟��ߴu�8��'��7�/�i��aãYYdLD�� �"rO�����h�ԛݴw��|�BI� i��C�6���C�f4���1 �����@
)S`8�6c�	����4���D�O ���O���Z�JW�Q�p�@7���^�˓_c�F�@6�yB�'�����'[�����Fp�I�f
<���+�>�r�iA�7m�g�)�Ө{V�CE� s���@u�N$U�T�Q6�24^j�K�����l�O��L>�*Oաև�"D+�����&W&�8�a��O��d�O(�$�O�i�<)�ii2����'F@��J��4xS�u,	�G�'Y�65�I.���Oj���O��T��9���q���B9�r6>?A�J�t0��q�����j�c�t�V�`5b�^f�a�|�,��ǟ`��ԟ��	ڟ���b��t���V\۪�FeM��?i���?a�i����O�b�v��Op��*Ҫg:.�����DK|���b7���O��4��%��u���Ӻ/*3R��&�35�I�C�j[)��{?�K>�)O����O���ORa@V�@�����҆`�A�O,��<���i�"9 Y����q������$�WB�/CA�#�<���x}��'�r�|ʟ��ː�уZ�,�H��D�h�,ZFbL�;�|����z�^����T�TM?1I>ѣ�ζ~p�p�	�0 򮒃�?9���?����?�|*O�@o�>�J=�����*j���GՃ]T�P��ry"�z�⟈��O��d��8���3��4���:G��e�f���O�FbӦ�ӺC�MS���R������9Ҩ�t�ڲB(��щq�̕'���'r�'���'`哗=�v*�[�{�4l�a�!"&8�	ٴ5��pk��?y���'�?1��yGjWRBR���@�[-T�	1�N�~�"�'�ɧ�O��9�i���O^R��"ɘ+-�X�要�!��D������'�'��	Ey���e��Б�U�MU�6���axBeqӲ��)�<��x���t�ك ��&.^=>��E��ɽ>����?�6�x2���kl�23��<������$
	Py��	UM~�hm%?��C�O$�ء0����ņqu��+�p�����O&�D�O��;�'�?��J@�`pD�&��,\A�� ���?�iʾ)�U��0�4���yW "���c�b�;.����L
��y��'�2�j��S�&h���`W����?� ��RO��,��DY0�41�%�7�d�<����?I��?���?1&�H-�CW$3�:�w���$�ǟ��̿<����O�� yc��h��P� ���c����'�>��iR�6�UU�)�S�����na�3R#m�p�&�#��'J���%NΟ���|2^�p�c�ؿBp@0���dLjaA�"N��(�	ҟ�	ǟ�ry2Cr���)�Op%֥�u���Q3��?6ˠ��%�O��m[�L|�I��M�3�i��6M҄-xf�!�cM����t�M�j5��hD�n���4�Јu!Ꟗ�I~��;O6� �&�9���s�:\�4͓�?	��?Q��?�����O��m�	�-Q�*m�@@�6?(�6�'���'3�6��%֮˓)��V�|��F�#V�Y�� �4��g�hO�Xm��Mϧ*/�ߴ���t�C1kW 7�|W�4J��ӢD<�?yp�$���<)��?���?��g�]�I"F�P��$8���?q����Ċɦ51�*�ʟ0�	럸�O����2GV�o{��j�D�i�*�p�O6��'�,6M�֦ŁM<�Oas"L´
�fLhV��y����waP�'s4��!iE��i>I��'�'���'��1Ή��lQ��x-0������	ܟ��	ʟb>}�'��6m����X(b��"uD勷*({f��@#��O|�������?q�_���ɵ09�ͪ��^�D� ���'��I,�Mk��F��M��OfQ�r����d]��A��KD��c��,�rpY�m��'yR�'m��'��'H�Ӎv�(yu�TpϤ��`��G
b��49%��Z���?A�����<!R��y�v�:HZ!)#R찪���@x��c�(�%�����g�zӴ�I�+����^�e�Z���EɈ�F�	
J7�iPV�'N��$�l����',��VhV���"veY�g ( Rq�'�r�'sQ�@J��6�ݕ'*�]/&�l0���11D�����O�8�'u�6M����@H<Q��C ���#GQ'�83��n~C,$b�9@�b~j�O@���~!���#Xl��*sc$T��yj��S.���'��'8��S�h��^`���NXEZX�qnȟ�9ߴY�(Щ��?iv�is�O�N�/�ne�Ǎ7����!�j����Q۴Aj��&�MV�v��R�%����T �p��(�d'lk���g^:Rh��%��'z��'���'���'���Iץ 5�8Y�j����Y���شP���?������?!��M�<�r���
�Ie��2��Iꟼo�*��S�Sz�l���- )4PC����������;��'�
 ْ,R՟��v�|�\�t:�J;;�U��37F� ���T�	֟��	ǟ�~y��g�Ȩy��OF��t)X�I�x�E!޺	J��p1OZ\o�T��f��Iԟ�������4hJ�0�����E�����f��pn�A~b 8���Pܧؿ{��[72ʨB��Lw���I��<)���?Y���?���?я�dH�&x-ʳ�Y���>�b�'w�z� Pstð<�$�i3�'�N�bc�� Sb5�w�+&ӈ�A�|r�'S�O�HIq��i��	�S���z� ���da� �	d ���(�OVf��iy�O{��'�BA� �����կ	4�ݠW���$r�'~�	)�M㓎@��?���?�,�P�0'Ìe+��4A�Dz�P;`���;�O"��O:�O�S!?Сɲ���P�ʽ:aȑ�6}L����L4?ͧ2%�Ę(��Z���y��£e�jXR � S�,����?)���?��Ş��P�Yh�i�0[z���tF�xA$��$�'��7�+�	���	���2��&jCj�P'�K�<�E!�CP5�M�d�iU�e��i��I%k�j�p��O(�;>����ºj@v�� � +���͓���O���Or�D�Od�$�|rcI��U�ʠ�c�L�t�q鎥/̛���p��'?R���'�:7=�9) �Cw<);��Յ$�X�{�6-�ѦiZN<�|2��6�M��'�x�(Y1K�0�4g�;T�h�+�'��屄� ��C5�|�Y��̟�ӁNz¼	҄+Ӏ7�D��u�Y��������Hy��u�4M����OB���OZ �df�-\x�+��1]��ps#�$��,��dB�q��4Ɖ'�����M2x�$I��iG.xd��O^Irs�����h4�	H��?�4��Or
��V�竃M�<q���O���OF���O�}��EHD�bØ7�y�2��8b����7l��lϮOY剿�Mk��wc��SKW�W�����_&o��s�'uv7��Ѧ��ߴ#AdĻٴ��$޿���{��K|M��kB�%Z��fɃ�@�n�P�1���<�'�?���?A���?��M�;.朱��H(wjԀ�M_,����yw ����	ԟD%?�	�N$b-j��4_���uI9[��O`�l��Mw�x��Tm� r/:�gC	;�8hhw�8��k������d%|p 8)��n�O&ʓ%Gnڳ��5A#��S!��US|\���?���?���|*OJ��I�)֒�� T��KQ̊=�U&�<����˦A�?1QR�p޴\��6�b���v
�L��B�D֔O[r���*m�|6�5?鑊K�=|���1���q���ثkH�0b�G�2��8��c�����$�	��@�	� �Z�GF
	�H��!ʊg�t�Y%���d�O�n�=�2�kh��|�#�.zit��h�q�`�' ;0OX�lڋ�Mϧ  Y�4��dG�0� (ҤoEo���� �F�"�3�A!�?Q�)9�D�<�'�?����?1a��8�,XsTf��J ��ӈP9�?	����d���)�C\����I�ܕOs(x0
�X�� B�h�5DL�tz�O�(�'�2�'��O�)�Ob����As�}B��Ym,��tC,,ح��-{�z]�'x�t]M?�N>q� M)u�	Q���^Y�%b�E��?���?����?�|�,O�\m�<b�Ԉ��Ȇ+-b�As��?1Z�J�m�IyrHl��㟜A�O��D� F���R�EX�d����7����brC�֦m�'}v�r�Gm2.O E���KQ���5*K�s��	��2O���?��?i���?A���Ɋ	3���u��>|?�M������m��f�L��I�(�	T��������d���(Y�d"�a�-T��I�K�$�?��C���OL)�1�i��7: �`z�e�x��V�{��D�]p,��'��':�	����0�ipC�Y]?�cY�l�����ʟ�����ؕ'h6��4 ����O���87y.� �d�>X���i �����X1�O��d�O��%�h`o��5:�L��h�M�!�2?�v�ٴj�^8�ܴkI�OΆ���?�㳲XE[�RǄ�"�l�.Ґ���O.�D�O�+ڧ�?ٖ�+ ��σ�0]V)cS.ũ�?�!�i$$�PV��ߴ���y��(k������={��T�I��y��'���nӞ�JD�k�"�=v~Q���?� E�G1ndJU&Cr��Q��_�	Gy��'�b�'R��'1�5�*�#��Lj�E8" �I��M�Qo��$�Oz���D�X��A�`�ž6��
�S�$I�'��7���QzM<�|"%e�*l���R�j>����(5��*4�S@~"�	?Qt���iA�|2W����iٹDb�91��7kl`��Qş��Iӟ��	ʟ�tyҍq�p��Ԩ�O*t�g�57����ԡȊqt���9OvqoZw��-��I����Iğ �a���&�=:R �
Lx�];� ̽[�QmZk~R�@0�hL�Kܧÿ[#F*tlL �!ꉍVh>��ej��<I��?��?1��?����h՞|֑�^^��3�˺���'��v�@��Dc�<��io�'�Z�HQ��D^~_�25��	a��'�2���4a�<?����d{0��6N�.8�7�G���%�pjR�{D�%��'�zp$�8�����'S��'$�m����Hf�4Ut�a9��'�2Y���4%>�S��?�����յO���de�0�b�+I�6�����D�O���0��?Q
#��)�h;"���m��Сo��0b���䌅�#�V��|:�i�O$��H>y ěA�>�q��%h�B=�ը��?����?����?�|J.O|`l������
 �XmY #|02'�Myr+`ӂ�\Y�OX�D3=�Z�IG��&g��[o?Qd�$�O$ЊU�v�n�nr�"�韂�O�����Tx~�cB�vPT��'���ɟ��I���Iӟ��IQ���"7
Q9#,h�آn$a�7��;c�B�d�O���>�9O�oz��J�Q=���k�k�b�Ȣ4��ܟ��I{�)�#I�@o��<�aDV�S�J`mٝ1������X�<)uj�!ל�$I��䓎�4�B�d�=�\@�*�{��Ir@F�:j���Of���O�˓(M���@��I����˜�Xr��Z�-�93, �����j��5���8��x��
[وl�ȃ] �����������;'.� :��|�7��O��R�eA�<B�H* "��gč�l%�Lr��?!��?���h��\��p]S��D?k�nɡƏݸ+���DP㟸�Č�O����Ҧ%�?ͻ'���r��&`"���&єUj��w[�dӶ�m� 6p�lZ~��)�K����ƋEɚ�+�69�p�c�>�䓛�4�`���O�$�O���.s�=2p��"[$����K;1�����_8�?��?����e�W�򩘐$����hC6�/e�2�D��k�v&�b>u���h� ���2,ЩQ�։o�f��An.?�S#�-�j������d&G����v�*��d��c\ �P˓�?���?ͧ��$���R����R�� c�8HW`��@�AA�|��c�4��'��e��He��DmZ�$4��M����0�C#|Кݱ�j�˦��'��b�e��?��~��*oB��D�H�-�N4�w^1_і����4�Iڟ���㟜���Oa$�Sţ	:.�^qJ�m�>�P�O��$��݈�a9?!P�i��'�V�X�U��<�)Y/u\x8�L5�$�����|"�i���M��O����n�>-�@i�J�sF| �n�{�`����f�Ol��|2���?���[��)R�o��:�H��ql]�$��1����?�*O� o�h��Iԟ��IP����>rR����7X�\��h����d�g}�@`�r�oZ���S��ܓ{���٥+K,�xw癡EU�m�&ײM��ł�O�)	��?�A)���B^�p��ڔZ��q)e�A�x���O���O6���<��i���'fa	<�@E	3�8�ȵ��qa�	;�Ms��@�>�W�i�аRpC�w��J���3T����@m�~`ne+�nZH~��w����Z���((�X���͙8���1�TN��D�<���?I��?��?Q,�v0B�/4N�j�'|\�m��N���K���ȟ������$?�����Mϻ}c"Y�3
ͻxvཙ�i��
!���?�O>�|�E ��M{��� ���al�M1�܀�e�"f��'8O� ���~b�|2V���џ��c�d�&���"I�v�n�y �՟���ҟ���Sy�ir�N-p���O����O4x���W��5��j51H"�ɛ����O��d6��D�b�f�:�&��QD���K�V8��mU�"��Lͦ�qK~JT�������L�7��;�|�#��#ڴ��ğ��	� �	V�Ou��ݜ|V�5��һD3���R&�
0��u��i���O��D�����?ͻfp���&͕8e<YZR�޸��̓�?���?����M�O�n�8��S�"�h�	���!mT�P�L�LNl�$�̔'5b�'���'��'<�ԈR%��$D�M8�S��̸uQ����4<V������?�����O*�ȓ��G-pp���S�{����>i��?�N>�|Z��b좬�����a�p�Ы�5�<�B�4V��I�^�=���O��O�t�ġ�m�F0,9��Pj����?9��?Q��|/O֬o�^=����w14����/Cd���H��gF]���MÍb�>���?���-r�H�5ћ=$t5J[�vռ�� A��MC�O�U�a����4����w��E�2m�?"O0�Ex��'���'���'�B�'a��ܰH��?5֥GI�|�0p��o�O����O�lon:���'F6-/���a�`�"�T�H�D���K�AG�)'���4J��O��|���i���:dJ��6.�i�݋#%`�P���ũj�!o�iy��'���'�Ң�o��ucv�`�d	U���'��	��M[SK���?���?I,�^���PSZ	�1+ؐ �`�[�4A�O�o��M�Вxʟ�EhȽ#�:p rN�%<t�H�УѾ�܅I���%�P��|bVf�O��K>����X`���W�K+�^r�!��?����?	���?�|Z(O̔l��W@e �!�0g���w�N(S��H˦!TGyR	~�D��ѯO�lo�*A��$�8"t)�O�7:8�Pk�4	U�&d��
,�֒�P�Rآ2�$OMey�A9]>I��Ŋ�x���%_��y�U����ڟ���ڟ��	�ĕOK
A+�d@�h�2mC�/�Ř��{�x����Ox���O����d����s�����y�b=H��
'w�¸)���M�|J~����M3�'��m�婜�&j ���[`�'��=`�� ϟl��|�T�D�I�\yӭP�j���c��zj��'�şX��џD�Imyr�q�n��"h�Od�D�O\8��G�K�Ub笏,&�*�%���������ܴ<_�'�*D��E�r�:��ǻ1h���O�u�C�ó464��逳�?Y��O�=i��g?dQ�G��%pX˖l�O����O����O�}λ6f21�v�ϛV�����V�{^�
��tMR ,�?!��Fl��4��H����|�H�d�M�z$��8O��m��M33�i�R����i��ɘ!AH`�A�O��-)�aǓb�R�3C��20@�av�R�IKy�O��'m2�'���a�$�	1�_�x����ߨN � �Ms5@܀����Ol��B��аL{��BP)޾� fOJ�)��$�'��7͉��i�J<�|�@+��%%<��N� mFZ�dC�4G��QBQ@~bȆ@u���� ��'p�	�Cf$�5��uRJa���H����	ܟ��	֟<�i>-�'i 6�ǰmR���R�,;�d<(p6a1�e�-jl�$\��?	�\���ڴ����i��ٚ�@R� 	|ȓ�'Բ^DY{��6x�7�)?9emG"�2��*��ߙ(��EҸ�y��� Hsތ�V�p�t��ȟ���ȟp�	��`�z�&�L ��c�I��,A!�7�?����?�!�i���O�R�s�d�O~t��`-_X(q�` �)8�)q��g���M������cI�������4��0�����x�\Y��R=i�B�Ǫ��0:�|�Z��ǟ��	����q���k�ᘩ0�^��#Zǟ���ty��t�j����O��D�O�ʧ_&	� **JH�t���]n�@�'�*ʓ�?�ش�ɧ�i�O���hI�	���h� �,�P1`G��f�8P���S�72�s�	�c:�0��>�<�5�ĳE
���͟���`�)�Soy�s�L��C�k(�3�	l��	��t�Q>���DM}��'��ԃM[��h��Xx�"X��mT��,�I5ކam�U~�`ӂ'-�l��g���uP1g�@�{�>�K@�$���<����?I��?����?�-�4��Q'�fH8`qԪϘS���@�hEͦŲ�+�ǟ��IПl$?�I+�M�;q`��2ǁ�p�b�`�;e�XL���?)O>�|"!��<�M��'I,բ�F��L���#�-e���'m4H���Hߟ�R֑|�Q���ߟԛD�חɖ��Ƌ�3�|aQ�����������	Uy��o������O����O����_�MvʬX����b%��� ��OD}�'�R�'��'�NI땈%Hz��f 8La���O��ґM�5�4,���)���?鑍�O.M�Ҍ�--4Ѐ�`ؼ]��u F�O����O����OZ�}���:J�	IB�R:�ؤrfD��m��9��f$�T��I%�MË�w��*�D�Wؼ���+p�DÛ'���'��G�.��&���+e�
�2��t�Ъ v��t�_�z��H�Ĝ�1��&�蔧�T�'���'Y��'0�����?->ɂB�1��J�P�<��40��ؘ���?�����<�B��� �^�A�@"�wh_>�	����y�)��'��� &U�v�G%[��M����9 Eqr�]k�	�sj,L���'� �$�P�'�xxH��H8 C���-T�֠��'Q��'-"����V�p`�4}�<����v!�hX�Æo�r��dn�)���ΓS2����N}��'3��'!.�y�O�i��qB�ʞ�:�T��oj��V���jPdRm�T����4H�+V�`Ğ1���]0<I9O`���O�d�OB��*�F�I�]�T���}ϲ!QP,P��O�d�ƦaӢ��Jy��g�ГORh��)YZQXe�T�#��)7�%���Od�4�Rt:aAz�����gQ�A9֔�щ��:�I��Y|�$L)����4�"���O.�Ѷ��@�� �T�*�YƌL�G�>���O�˓*��6���y��'�V>9;V �"����B��A�\�!w�5?�U��0�4Gś�(�?m����1�����Y:][0YF�\�}�Սo���|����O�%BO>A$$��ժU.�H�(�3���?Q��?��?�|�-OralZ={�,]��V1*�9�(X6dT�F�2?1Ծi��O̜�'�7���k��h0��@�{��ٴ%�M4��l��MK�
�M��O�l��B���L?���GV(�������g瘝f�n���'��{���D��`γsr䱔V"�J6-S�	���?���Bw��Ε�gb��1�E^{�Q{�IP���D�OZ�O1��)��z� �	�@l�@���q\�@p���%X�z�ɴ�*���O��O�˓�?���}����%�h��)��;cO�%���?I��?�.OPlZ�3� ������I��bu�e*��:�R��	�3r� ��?q�^�t��֟�'��s`�1v\@ � v � +9?��.
z��PBA�c�'s����#�?ATd�z���iD(-J.�}YE��?���?���?)��I�O6���n��#t��:��-�Z�H�O6o�H���==�&�4�AxՃ�>}����qD&]�t��g5O��o��MK��iP�Z�iz���L�4]��O�z� w7�b@�BLS�sŸ���H��Qy�O_��'db�' ����|�� i��'A���q7 ��'�?�M��%��<1��?AN~Γs"@���t��| �K�3t\h8�R���4 ��6�+��:rTp5���d�vPHc�'9�X�PD�	=O&�����'��|%���'�z`�����1� �Z�[�A�b�'7��'iR����W�`aܴ��m�S�2�򰭂?#�V�ӥI!�F�Γ{ћv���v}�gsӔ9nZ+�M�egV6k�.#��1qR�(F�,�I��4�����2�<���'̸O����3A�����3܎�S�oI=�y��'�2�'�b�'����FN����+D�r�1a�B����?	�'��x�O�H71�_�w�zL�A��{��:b(���$� �ݴX8��O�x`1��i����f��"B�?ı� �ܪK�hu�!p�BA�Y��`yb�'�"�'�R�O�0� ���S4p:hc��Ϝz���'�剖�M;r���?I��?	+����&�%]��0�N�#{�f��束�2�O����O��O���my<ɀ��75ݪf����ۖ<d��r�9?ͧq�j��F3��\�<����P$!ꑨ�a�&Xv�y���?i���?I�Ş��Q�Q���*_��щ��/N����u�.,�Iϟh��4��'�j�����;��@y��M6B�ݓ�8�6��Ѧ!�h��U�'���{"l��?����eҳ�'��0H���H��V�d�<���?1���?q��?,�.l�0����]Zc\{ܦ��P�DЦ�3�'R�������T$?��Ɍ�Mϻ^IZ}�AB�^���*7�/����'&�F�4�����1ԛ<O�xj#*�b���@�/��b1Oȝ������?�Q@;�d�<�'�?�u���J�=�D)���4�C�ɂ�?����?�����$P��;��AǟL��蟬���ϸG�Hrw��6H��y��KK�_(�	㟴o�4�ē"��زK1<9HH:�E>-���'}r@���� ]Ѳ�1��Ta⟌1B�'���h� $x �(u��U��A�'���'���'��>���613j�;p�W�P8�!WA�#%�8Y�I��MK��B��?q�h�f�4��p$UW���(OU����Of��f��lmZ�m�vHm@~Bg��*��M�Ӏ#��h���&<�*A������=��|�\����I���	�������?F�]�����\��
ec@Kyb�l��1�P��OV���O���R�Ĝ�� LS�H�^���I�Λ8=�0�'�2�'�ɧ�O�ƥ��G�I�ش��(K,U0֌	�A��]=�F�<���A�"�Ip�IEyr�J:�*�R�@�+I�*X*֍�7:��'r�'��O�剩�MC �ӿ�?A�B��]�*�h�m�$ߢ��0���<���i/�Od��'(��'+���d�ȅ��L-J"�c��8oz�a���i6�I�+��ݸ�۟N��x��Q�j�ɋ��"�^R'اWc�$�O��$�O��$�O��$*�Ӄq�tE��I�)뚽��(ͼ'�,��՟��Ɇ�M�	�|��&Y��|�6i���F��^�*��Q).�'�R�����P˛���֝-iY��I4��(n�0��u+���F[?!M>�*OJ㟤�T��(��}*ă�)!�|�D3�7I��,��h��x�O8��f�(�\�Ï�/o4�X��O��'���'o�O�3� |)qkמ`R���5e�K�����l�6&w�1���Sv?)N>�B�F�0d|@�� �d�.qag�OZ<Y�ib�͈����:@QlJ�%�8�%�Xo�I��MC��l�>��,��)X�iN�X�q�`��##z)���4����՝?������M�[)��<T�݀@a�A��Gu6Te�"
�<,O����ۅB>�ӓ@V�{T��FG�(�5�	�l˓�?���$u��Ŵi���id*�l�!GY�Do���M[��x���KT�%X��4O"�:�Ǎ� ����GFe �A"?O��@�[!Q��<�סŃ��P��� �r�fE����srlH!�	>] @=Z�d�9q�.�b)��  ӋפQɳ�o���o�"��U�R��[���9`�&��J�$TH��!�O����	r8�	xU:9�#��9g,�������! $�$6>2�ӆc�:���! �\�f��A���|��֧���E�V�2Pr9`t��'^��a��Q�Z���C��H�")BU�� �F%��T�"�V��n*a3�����_�t%��΅H��`���6���0�,X� ����������џ �*N�z�.1�K�{@@�`��O$�MC�����O �$�O��T`�O��'&��7�R:@Y�#��~)p`�4�?1����D�&4�
��O���'���D#N�+��̽"_ʁ�g�cO��D�OBS��#�ID�t
ӄN�ԩ�ګ7�0�Pe���e�'�0-H�*f�����O�����ԧ5v��g*�!�@PyD�� D�2�M���?QC��:��'6q�"Y�ѴG��X���C55	��2�i�ް�f�tӜ���O���<��'k�I$,d*�!^��+c�S*(d�Q�4��s������OP��+�Bt�w��L�RKF-47��O����O��V�c}b\����w?A$#�D��e� �� 1Fq5�g�ϖq�L>y���?1�SP�ٴ�[B�TcTXR�Xu�i�r&G�[l�����O�Ok��#%��i�M�2� ���c���+���IPyb�'�R�'@�	�DS�m�3��J`�Σ씬J��N���D�<Q����?Y��B�p�с ��eC"�I�,��a#l��F˕���?y���?Q.O&Q�ƦZ�|�t�Z�^��u�+�:uh1�ӦI�'8"�|��'9��6;��$ʼ��3'&	
YӪ� ��['m�����\�I�l�'���H��~����}s#I��7��U���$F!	W�i�|�'�r�_�h�qO�[��L>@��L�uK
�uh���i���'��I/[b��驟h�D�O��i��O��ZD
ޡL� (2�иJʘ%��	�P�S�T���4'�.�����8�U��a��M�+O(���O|�$�O���������2qs@Q0�F�P�)��
���E�I����`�S�']A���lШKE�L!5e�)�-o?e4�-ݴ�?���?a��Q����Ĥ ��(���k�)�0M��aF�b7�$j!*���O0���<��Y��	�`�&+��Ӣ�ڧ�
3G�i0r�'[RMĘc�O��O��A�%{�H�=�i��}�6��O˓`��1W?��?i�'��1A�*�`�(#���l�d��4�?��	�����X����	�LL�Yj@�'p��V[c�Np��W�t�%@�!��c���	myr�')��{��$2d�1�ĈZv��x���L.�����IO���?��'��� �Cl0&�9�Ʉ2�4垈�'r"�'2�P� +�jH���t	��J�����+��1�ǎV���O����Oʓ�?y/�F�D�5�d��sh{�p�����ZW*��'r�'VBY���I4��'��Y�3��9X� ��]�w�z({��i22�|�X��s��ß�� |8 �[�N�jD��o���G�iHB�'�剓]f<�J|����1A�~t	�(9�DM�q��LJ�m�Oy2�'��kء^R��t��5FEL��#�M�`��i��J��d�O�h�Wh�O��D�O��$��d�Ӻs��ZGf��e�֩V�@����٦5���@شF�a b�b?U�Q� Kx�YЃ�Q�)h���p��1yv��O��O���Ꟍ�S�D�<����n�6u=#���b�6�:2$p+1��z�`MaeШ]������ϚU��iش�?���?o����?	�OP���
���MH�G�a�J-�e��C̓0�<=����O2�ɞC}���	F?t������D�7��Oh�����<�GX?��?�#OE)v������X<8�X�)3�	-�	^�="23?���?Q����(~�\q�f�>l-���`��d��Q@�gU}�W�,�	fy��'-��'5��K1X��H���5	��"��y��'���'���'��	*\��؜O���C@�/��h��ӌ^�b̹�4��d�O@ʓ�?���?�7JB�<!�G�F:lXpE	r�ة���R�@���̟����� �'��!�@�~B��F�$k3@R:-q���DJ�# �q�i�T���ӟ4���X���IP�D��1h��#��F�&�B���p����'d�X�@���Ǣ����O�����Qs�ĸj_0l��MLb6&�"�q}��'c"�'x1�'�s���'X�ր���:�j�Y�#�ɊEm�Zy���b66��O����O��IF}Zw2�)�\/A��ȡ�N��	+�-�ش�?��W�����?I(O��>�ѧ�oD�U%��|�
أ`�m������� �	�?=I�O�˓"=��x���.�h ����f�ib$��'�Q���:��� �5Y�M�x"�%".()����iz�'���ʓs#�ꓔ�$�O`��t���Xc��7����έ,��6��O`�eH$X�S��'��ߟ��B�ԣ1L����y+̑��i	��ɗP@�����O���?�1T�X`���I�@hҭ�ҝY�.��'2�'�R�'B�'�"Y��+s�<�j-P�ӅL&|��&�)
B�ЫO>��?�)O<���OF��29��[�`j�QK �n�X ��n�)��O���O����O��ru��v3� ;�MM�MX~���ʷ{����%�i��ȟ��'���'#��yb�ۤ0�\5	�	��=CF�/�J6M�O����O��$�<�T#�#��S������ݤE{eqq*�pĪh�T�5�M����d�O��d�O�Eh�1O&���O�,��@	g���� ��6j:�)e������8�'w��H j�~2��?��'-h�Y���m@��T�gY����������}���J��'��i��5ܴ��s�ػj�܍Ro4{���V���5J�#�M[��?����S_�֝�&�zzA@ߗ,sz-z�C-07m�O
�d�|����}�u��t"��s�O.Nڬ���ަ�yEj�M���?����bV_�X�'��7
�Mc�[��0U��$b�B���e��j���	_y��i�O���A*])G:q���Ih2�������D�	�7 �<(�Oʓ�?��'x�J�)̌g�P��$L�;=���ݴ�?�)O��Q29O��˟4�IៈJa	�LU@5��b\��ZЬS��M{���t�cg\�H�'D�_�L�i�Ղ�n
e*N�Q���p���>i��<1��?���?)����䄥D�v�擧vJ5#��em��􋘬a��Iky��'��	럼�	������30���q�յ[}~�`�L�<f�Z�I˟X�����Iܟ��'l�՚��y>)R��!m��3��ʈA��wemӪ��?�*O����O����3��d8pRш&�'�p�Jܾ=��5m���	ߟ��xyB$\q����?�1z9ڝ�U�����Q�C<q�<�l�\�'C��'��%Ւ�y��'���D<g�Q�
XDP�G،C^7��O
�$�<y���3}��S֟����?	@�&E����q�J�EG�KUė��$�O����Ot8I0OʒO��ӳ0
I��^�n��ѓ��?CeJ7m�<qR�����f��~"��:F��4zSD��e����C��F�g�hӈ���O�P!s��OJ�Oxʧ�~ \����O��(�����MK�oT�:<�V�'���'a���'�$�O �Ь��4�1����1c���Y�J��}����'������O ��ţH�0�RI3��Y�$����A�צ��	� �	�!��x�J<i���?y�'�L�B�9R}��yԌ�l�&�S�4��M8D���D�'���'��P�b�҄q�����*��}S��eӤ��G v`&�\�	ן�&��X,j_����:5�q	��,�¦x����Dk>��O&˓{ڈ�Tlz9�(g��e��\)�@��5ƱO��D/�d�O��Y�':����<��kvb's,x�2O^˓�?����'5��9�6|�e�~D�Ip�VTP��W���	ڟ�$���Iڟ��"f�ן��2@J�=��к0��l�D ��R���D�O����O@�N��S���hO�S	��1��*���#+�=566�O^�O2�$�OP0R�6Oj�'#:�`�I� -*��֫ыg`d��4�?�������$���'>��	�?�`�@+�ni�M]�`��c3�L����?�e
��`��ܟ
�� DS:Ɋ��Bo�'�i ��?}�H�4]��ş���?��D�%W�T�[RjȢS��YcH��l����'Jb���a��|b��Q2YN525EF�tp�P"^�U��F@\3Fk�6�O����O��i�T�ꟴ��!o��I���(�u�U@�M[�e�(�?)O>),����?��MۻwҶ�!D@�LIġk�(��:����'=��'uD�X��>��O(����0�m ��\H�N٣*vB� }Ӷ�ORIj�`z������Fj�`�$�����6��Ց�����	4 ���M<ͧ�(O��1�h)h�`v��8pX���V��[d�����ş��	����|yb�<(�V� ��8�d
�zݖ�i�o!���O8�=���8`�{7̖$\؁I���"Tr( %Ю�?i-O`���O����<���R��C�]�R��F��8{�v���m�jT�I���F{b�'�6�:��'�Ĺ2@ծ{�$��W��I+jL�aDg� �D�O���O�ʓc~�kМ�\c�|[f"���
\��$��4�hO>�d4O���D+}BNU>�����)��e�&`�q�О�M���?�)O:�(���_��4�s�)T�ߔh��$�W[����$?����;�"���$��'8�r���$5eA@	�?i���n���4j�(�������I���^yZc�<ɂӄ\�i���K~���ݴ�?��QQz16 ]H�S�'Dp<8���ޒq���-�7%<$o��{�4�@�4�?Y���?��zK�	p�$�0�La�QA
'�6LsӇ)#W^7�OQ����}�ןL3�c�T��s� �ߘ�����M����?����V ���?�/������h@O�4A��jU@,�Aa�M1��'��8�m2���Od���O�0T�ȱ �ލ#��8�;3��1�ɷ.f�hڴ�?���?���M��y?��C*"|b���@J$\i́!L�b}����yrX���	����O���:� �x�&��;�d�І�po�����[n�f�'���'=rʭ~�(Ox��L~�鱊Y�,��:u��9&�� C2O���?i���?Y��?a�d��1�&��N!8B��ӾE�����I�@Br7��Ol�$�O�d�OV��?��`��|b�iy0少%QT(�5,�I��6�'��'�"Y��#�.����I�Ok�R��͑@�Q1R+�B�hk8�nZ՟�'��'T��M��y��'ҭ�D��P��U"}�$���+S�Q�$7�OV���O~�d�T�`o�����	�,��m��meR��@t�U�$���4�?Y/O���T*����On��|n�>�u��76�L����v��7��O��� /��]l�䟸��џ���?I�	E�0C���4y'��#&r�����|}2�'��"��'���'Y�b�	�-M?�ݑ�/UW\�"#�	�T�/�&;�&6M�O��D�O��i���D�OP�$�!��ˠ��*9��,ʴ=�l�lڄN��\�IҟL���t����'��] V�O�8�D��MJ�FA�6�fӈ�D�O�����N�V��'��	ӟ��mi} �Z Ŵ`�J��v�tl��T�'�I�����9G�&��'@��HަR#V�A��Z�j��X9�'�f�QF�F�>�)���jU( 8ד{�$i D�	��e�X�yʕ3��:S4 �)�.�N$:�#Z4}B]��D��A�nF�m#�5sg��0C�y�g,����{u%W�I����'�('�h��t!\!o:U;ЧO%D�}� �^;����'Q�b�$�%�$���j��61��aCP���q-
Dô @���t6���	�<�SCKƟ����|"��D�[��q��_DZ4�8�9P�a��$ ;c���DԴn�j5z��	���dh ��5�l�*�m*6��A�U�#�T;@
ݫ �����׏��O���'��S�:��?C�|	�Ђ��N�8���3�Iz��P���x�Ɉ�"�_���0��p�4u%4yv�b|a��h�",�T̓��D]4
�6��'��X>�������|h��J�[B��!�ހiCL��u��ßT�I$3� ������k�p����.�?�O$�S�o<&l��bUUI�!�{���'�LTb��O�=�,Q��˄Z��>�ᶧ'Q�I���5H|��-7}R��?i��h����tUu�ġ%*��`"���I�ȓf40d
�̈́{���GZ:�,���HOD5�s�������
�)7tu�@,Ts}��'kr�ܨFJ�5:��'�r�'W�wy�;Ѭ�
8~��9�����s��65��-���O(��#���(x1��'�ʐ��%���@Q��_ ��$R�o �X<n%���O^�C�H�9����	���!��ř3��ȉ��K,X�� ���dK�X��Obў|2�͜�;Ĵ��fJ%c�f�Rr�1D�x�!φ�D��i$�ɜ+C"��@2?�$�)�-OX��!\mT��f�w��Z���-T]z�f�O����Op�D����?��Oe�!�bώE���8��Nı�у�`(*l '�kA�"�<��<y��(v?~Q(H�_���u$�&`d�cݞa�ԕ����iG�� �A1vQ>�<YW���B��[?Vf(|#K��5�����o���x�+/+��� e�.ȉPm;D��eAщI���"����_g�64�I"��=�T&IR�&9��aɩc�8!x��|�<Y�J�CC9I7	ȡg����CFw�<�Ī�/Θ97n������%�Cp�<)�,�G�n 3��C���iv��s�<�WO��I͒D���9iJ�s�FV�<S,K�>����� HR���V�<q��7qpZ�v�!%Ǣ�7o�I�<���T0Y~�Ɓ!&@B1"G��H�<agAD"_I@uCU�O�'�r鉤
BC�<�Ç�+&�a�̊�+e8�q�$�{�<P��$*<@H�Ќ2}^����{�<�� ס0L\���^ ����'�r�<�7DR/(T�J%��T�1у��b�<��'F�8%2�0O� J̀���C�<	�`�%�:d�u�j�~��U���<�g�)n9��i��H�����)�z�<9�� �Mk��P�A�s�<Q�O��s2�T����J���!p�<B^=�n�a���r!������V�<�M�"�e��T�&pS���O�<���ۤ)�
����@�f&���kJd�<9���7�ʨ�$
ͱ�.X�LR\�<��#X�j�Tj���)S4�����p�<�T� C8�	2ڤ=<J1I�Nn�<� <Kg��6���`D�ǜin��"O\}��K&@���	کh�J��"O�$Iw)L�^�ꩁ�Zk����r"OH�#1���D��&��5�$"O���� @�� ���L�N\�@z�"O4�c�N��[�z�[g�/p>�� "O�A�h]=g�]�@��\X�
�"O�D��� �}��9���2/r(��"OvpWȄ�TXa��ѕU��r2"Ot�y���mzx�m_�Rfp`0�$I�;(� ���e��H�0< z��Q�@�*�B�I
O����rMX Q�t� ,�.Q�ޅ��o
��U�Σ|�'�	8l�V���+�Nؙ~x^PP�'�nyPG
��5�B���P�zԖ���q��Ic.5�O�@@���I.��	�A[$ۜ!;��'nQ��I�4c��ɒ#q�hrǡY�B�D=#���~W�C䉃:���BG�"�Hy�J��ɚ��I�LS�`��E��	%W�򙱗l[${�I�0���y뀙���)$���p�Ĝ2@���t��ip󤄧�(��	�w��D��ݗM.�}��&ާXk�C�I;1q�@�5�ʶ%����f�]&N�C�I?[޶��S ��BA!M��B䉉IG~tٷEÄ9㒱A�핗�ZC䉛@��uq��˺7��9�@�++8C�ɣ"�:d�a.�<R���/>^��C䉶I��܃t�@3^x��A��q}~B�ɺf)0x��怶taēD�n/LB�Ɋz�4*�ދE�2U�w)OZ�B�I�I��AYPO[�>)�1��;-�C�I.17�8�b���Q-�-���!�'������C�m6��q�	)V^$1��'�8��	����JC�@P�'���W�D&uΩ��ν�J�{�'dBJ;2��k��
�] | �'�����E`tK3)�I�'T�d��ˊ�Z��n��sl��"�'�����(��L�L�*U�r���'H��6�V=y&cQ��'d��*�'/Ɣcu��5u��)�h�2��	��'���0��[�����&���XQ��'�´x��К0ּ�����=\���'%�A�玘�%	�1ՁW�3��t��'�j,)��:7�q�F��!#�"
�'d5B!�*�2�4��Y
�'v��B��U�V1�Y��.40���j�'���`"X�>��H���Q��a��'}zf`R��Zci�Z<|80�'>ͪ�.C4 � �� ~~����'�X�k֬�1��YY��b#����'�bM)��L r�Z��A���q��+�'��t{wOȎ8�1��		�lV��R�'Fr(Sܨ;�<p�h�1����'?�`{vGխbʤ�u%L,`��D@�'�$ݣqk�:�L�!F⋌T�Hu{
�'d$P���Kޜp�GS�6�y�'mRA0Ӫ\�HĚ��X=KO�t)
�'���DU&��U@ �ĄF7ƕI�')23C���A�P)zg��;7b��'J�h�ÒH�\�1&jJ�f�(Ik�'j��x@L�"����F͇5����'�0-�n�;n"�ي��_.3Cd��'J��s'­u��aB��2rp�'�u0�C��#� X2SL�u�x�q�' �(�r�M2q����bJ&r��pX��� ��R��ť��(�j�t���N5.^]l�aWRm䧈�rB�(J�8��QP4R��b쏰�y����0ՠ�`(�
K��]�f�թ�yRڀH������',��y��'yE�e��h�9�h�rł�0>��HC�k�\1�Y,nU��E�!U��8J���ʂX���F�{ݤ����#:f�H���+&
�0�G?X.#<���I�t�B�H���c$���+>׾���k��ud�i�pI�2k�!�H�A�VE	� E(��L���{]���`E�@�B��6�ؤ�0�,x�#}�w�Hu aL\}X$�s�&\�@Pb���'brqq�$N�O�6����[}4�4�$.�O����bS+	�4�Ck]��u�͝r�'�X̂�)�x�����Mݕ:��%�ۓt���V��d_Z���Y{V��a�2@�{P�4^���oU�y����Ā�_�QS(T�h$�qc�ڸ(��OXy�2&�	C�}��N]���������:)iC�,Z�@�3����m!��F�e��9!�R&j����%n�l�XƎ32� d�bgO�Q�"��)ʧ.y��[_�� �_�4��EȈ1d!�DZ�Z0��
����Hk��P�,R3�D�I� ����A<LEZ� 1��j�ʊ�����D�f�[�z=:ab��@��{2�ǃS�		@�
�L-px�6*��!�g�V	^%�=A%��.#���%�/�O��B��LA|Т��"O����I�X u�� l��
�ME�<�O��p��" �oٲ�J�mL1�'�B��wG�
�N����|���OK3�����4VN����
Q��hk��9O���Ed�5,�>��g.@8hy*�cG"O� ��Ӕ\�� w�\z��e Ta�|(0L�1C�O�d�EM$���I�n�����@�:^�J�"��8�X����`��7-Fu����ƴ���	b�l%�(׮��+�pmy��'�ؐԏ��YD(J3����	�Ó>T4Ԋ�J@�]V�'B�С.��B�z�P�oɝ~��+�'�rH+���:���PcԆ&1<	*� ��rݠ����.!�VL*�˂��h�J牋|�8
�����f�30�C�I o�T��!�|�~`�P��
�8��Q�(�ry��OE�@���c�9 ���S�	�L@�$�Ʉ;�,5���-/axb
j��{`��Wlx��!�$)�:=3E@Ʈ�$L��]�#Q���d��I#P�p���[5�Z@���)k��H^�ϓ&�`M[7�(8d��� ���|Rw̜/E���Ib��	��B�\U�<���
vW*�:*E�0�n�C�K/8���bs��I}r#
�?�O�@�j.k>I�w#�U���=r����A,�L�8���Q8��2�O�9�ՠ ��S�l�p��ЋY�hu�A��O�9q��+�����F�uW��\�'��L9���Y��݋�:ެ 3���%���q��H�E��)/��I�,��q1�"G7\
���C C��& 7c�r���[-"̭2�ȝ(���$!�CZ��P$��
#�(�f I��R0�=�O��ݎ4*T�AʥZ^$ `Q��h�C䉻;Gx�I�O�'�	ei�[�F��ec�7���J�����6�"}��X�!4���U�YV���4L ��<���L3�)��a� n�\�2l6vK���Q�&D	x�p�Ņaa�l��Yuza@��W+�\���w����*كLab�H�dN�҈��'����ټ&�q���V$y��Q�6�v�1��X>q�%Z ��>L4kGODX�d��/�a��'ɠ7^�:CL��a�V(�vi�L�ў�I6`ӭW'�ͻ}��	�2��9#:�ѳ��o4����ɔ_{@bÌ���{sc�1j��}�.����'�d�I&(�)L�N݁R�ݭ	F��K<�QO�#��p3���sl޹��
�L�'��Ǘ�!�l�a����f��۴,D�q�mH
n��E˵�E���%��J�;gZ����!O�;Z���
c-@���jX���A����R����CJ�b!�}���r��V �	9�P�'-���fصg��� �.��U.B�;�"O֥� ���)�v�2�/!��(��gE�I�<x�fdg�����l=֤�Ӻ+lH->��@R��wށ��]F-��Jr:1��*�O�ig	�.Hf4	�ïWL����d	I�m���BcK� ����f�'�U��`]t6��ţO*,v����{2��t~����S��Ms$HB ��OFT �	Z����v�A�	NH
��'iR��%=mΒM���ξY~ZY!�8�����$�4\y��	�'|��aI��P��-��d�2t ��ZV�
#��"|���"EH*G�|��eA��2�,Ål�<r� �s�ϗ?R��d� �� ���kp*����z�T@a��J�#{pő���0[�� ��E$F^�U9�_y�h	�W�:TAc��Z�c��Ē��� ;UZ�;E�dA��%M�7r�����P�FV"��IKQ�(!"�)$a��)���G�PD0���%I�C�Q�2�,}q�
U$s��Z�L�D��*���7'+qO� :����=�x{"#[�_]�¦�I0#\��_ ��e(��ӣ#�DɧN�4�2a�:�&�E툼v@�}�A�c���'`«T�z��Z�Ȑ$�F����F�	�~�L�1��仵L>Vb�Yb!��?Q�@����b'�V�nނ)�h���G�ɋdk60h!�$�"4�x�r+B.vc�9XAEY��ұ*D�Lw"�`3n��5���g�i����=A錘����R?��*�J��|�\B��!)�C�A��ZҨ@3��[5`�x8�$�
0�$��#�S>T�b����x�H�+r8��ݝ�}Bg���0<�ť��$~�˓�
K5�` ��@|Ta��b�.<��TC�Jqh�O%�����+K=����!�OT��G7?A��[_��a�-��9�^�ya�W6�8�>m+�9��-c�ç}�գ5�4D�`ٓ��y�����ë#�k	�]9\]��勚l�0��Ce� r{c>��G�>y�o�~9��k���~��£��e(<�hW�.t�� ��!����5d���F�R>2za�ߎ ��JެA�7��/t�4M�D��FG�|�ȓsV,c�hGu�j�/.�nȇȓ[^�-�S#M�az��._#-SV��k`�)R4Y�58I3��q?����:�c(�+�����KE�"����܉��X �͐dL�X'>��ȓ"�9a�cB�a�r�k�D�g�h�ȓ@����!�`�
!�� �/P4ۇȓ�pQ2�|�a�!T�ZE��I2D�������*Ia�ǁs/"�2ë0D�h�%�]���(�ǚ�r�U� �;D���U�ۤw�d��/T�P�
�P�9D�h�`�*�0���Ѽ�����M6D��"2�d� �r!��-T�!���2D��B��sf��!B �#f�TH+�n3D��3r�+vm��pi˄�*��/D�@�G��,Yn�A��&hk�,�%�:D��p"��=0!������.�\��c3D��#��\D���B�.J�B�AA$$D���e�ʲa��	0R��
x>�`��4D�@1���:Z3���c�?M���+��6T��"*Q�}v��!��
d�x �"O
�j��:@�<܁�(/6��Qg"O��BcF���p��D���"O�X	��/��+���&X�H�f"O`�'�&b��%��\�p	�� "Ot�1U�'=�(����*'JJĚA"O�${$-Ryz��E�5꼠q"OH1���hn'�0#(�9D"O����ct,�d��F~Iw"O
@ �׃%K�����٥j��mb"O֍S �X�Hq��O >]2��"O@=�.@0?��I ��Ԑ,R��A�"O�!)G�A &"Lzd́9rL�V"OX鋱n�f��2�#Mmy\�Y""OtM��d� v�]#sY:K�ܝ��"OV$��D�5YE�d8�P�lYh*g"OP\HwȄ:Pؔ���Þ�	��� �"O�0ځcǻp���1��u���`w"O�4�$j*x[��eJ_'^��93"OJ�+C�5�&%*Ҩ�N��x�"Op�;��vRਔ&��:�4�"OL�
vcEf�����'����"O���&N�` �8ab�u,	"O�l`��fQ� [� \��"O���9a�!�Վ�9l"Bpk "O�]cG
<���B8cy�"O��ĢT$i���������w"O.��2AG�q8�@Q��S=���9�"O��� 
E�6id$�q`�.��E�P"O� �[���&UD���Dj���It"O��QJ�j�x�V�*r�5�"O�p�&�r�XйP���'k�	�"O��p�ƀ==V|�󠎪Ph�S&"O�5�0�����x��7N
e�A"O�l�R+֣t� HxL"���"OV8Kt��3ɔ)	1@S/S:�4�t"O�i00��+K`1���5��XC�"Ol�A���6�G�N<(���"O��j�԰(��D�B�7Z 0G"O��{3�T�(�P1$�w�D=C�"O����ԸUStA���!�"O�#@fѣz��AV"�U�U��"O�[�JI@�DD,J�1�N2�"O�]1�d\
p�vœ5��8*@�թ�"O�i"AQ�j���,V6\*�Rq"O�x1��3Q�%�F0G20�2"O�A�J����亲��0�m�p"O�-b�i�� ���;7�ݺ.
,��"O��&�����5��͕
8�E"O�J��`9�4�W��:0��I�<�5j��JE�;� ��5��\)� �B�<���ء����'?,@ds4 �W�<1�o��n
�D��&p�F��b��P�<i���r|���ʶL����#D�<��-���,a#fg�j� ��	�j�<�D�j��`AFI�=W�ɢ��d�<yC
����e�4����$����`�<1� ��Ye�PR"ҟ[#j܊�!d�<)'A��bY0��doG�*��G+c�<�� �	���L����`&Jb�<qa��B��X�q�Wp09����]�<�����2�4��)�a�B]�<94gӎ"1v	����(�SPMQ�<�랳i�f���Ϛ�:��*3��d�<�r�C�16`�J����]4��\�<�T�=#"H���¼n����u��X�<1�P'T�1��9Hoॺ�'�N�<�FOů~N؜{�Ѯ�P�5&�L�<�K=��SS�[gXl ���F�<Q�˕�F� �����5y��*�@�<���މ6D�i�Qغ�t���BU�<9�B��|�X�� 8��k �F�<��D�4V
�!`Sh�4�qw#SI�<�'ވB׶	
�D�)���A�<QE�ٕ��L �AʫS244�#'R�<�d#	7l L�a%���@����F��w�<�BDiO�8I'�ۡU�"ف&��Z�<1�CR�[h@h֯9p�v�Y��IU�<�� ѝ.,�-8�O�R���.@x�<a���	3 -�"����T�g,�u�<�G�G�%z2Pq��_)9�f�B$z�<)���0���b��$n]С��k�x�<Q��(q@�pyN�w#�As�p�<Ʉ,ߺ U^|�!�� 墥 VC�P�<���0
�?Qb�*C+�.8�ȓ+)\�[S���E�������J7���ȓ+l���c�H�[m6j�ÀU&���ȓ0Tm�E��{y�@�GSD� ��ȓ=dV������l?f���h�~l�`��N�%��o�Cה�Sv	A�5���ȓA�pF*�z���C���-�lنȓxkN%�AÃ~��K�cOq������� A��d��};0�Ӆ*"���S�? ����uV�Pǋ�?�	2"O丸�Ȃ0�6y��=N���b"O^8
��� ,�A�B"~�3w"O��q�	{�58�HQ�#^pD�"O���w%ά~Cشj�SO��3�"O݉��A�M�F�(ċB�>A�W"O�P1�h�B%���־]�	��"O��r`�ęR���Z�Iʎ=Mp�(v"Oʜ %I.�N��IK�VDK&"O�����
 ��a��B��Р"O`a姈5)r<r*�� ��S"ODl1ҍ�o�R�+��X�N:U��"O��J�g�]�2.:�w"O�T{`��i�V@��N�"�Tb�"On���A��>W����[���,�f"O�!�'���y7���oH�trR"O�T2%�
7ζ �UJ[�1lI1�"O��+�D�FE�w�|#"��"O��`�Ǖ�cF�HbtHA#-c"OV�!A�ˀw�����?Wx�Dʡ"O�!��D?g�x`�"d��w}�i�d"O,y1���u!�}I���lݲ��P�'_���!��Fm\�aT-�`*.D���!�\$A�6V�J���>D�\��]�r�����:�pd1p�;D�Dk�A��LU8��R�ѳ�D	ѡ;D�\���f	��h��M`T���9D��gC/z� ��5$�1s��#1D=D�DR�@Cy$��Cc"g��y{`a D�����b�Nm�����K��݁��O2C��#"	��t��Fm����B�<K�|��ǣ��A�ъ@�0��B�	����H�*�zd�Q�R�n��B�ɚ|J�0���$�B�� `]�!5C�I�Z�8miQ	��HHshَF��C䉟43��V �)��Q"0$Kl(�C�ɜoόUA��A
 h�z�%ʔ2��C�	x��De,Uh��h"jL�I|VC�	r���ȵc(��#'Х,hC�ɺmي%�sJ]�)�Դ�a)F�8C�	�{ V;�ß�,���[Hy�B䉯C��X`Vh�:q���b�B�:,�B�I�L]�lH�dQ"��8�
5�B�I�nV�3��B�~b� R6�	�P��C��!�,:��[=
�XmP��Ϳ+{�C�	5iX�@�� ��Eᴉ�4�����7�I&E��P���\-Y�S%��o��C�ɑ� |Y!�\�8�!���b/XC�I(u�h���*��=~`�-� �fC��iݴ��fV�C�
5�F�����C�	 B�Q�k�P��ȢmA�ʈC�Y��I"��*YJ)*��w�NC�Ʉ6��$*� $~�0yۑ�]<[�<C�	8jU���Ճ=�mbA� �TB<C�	dԐ<P&L�L7�����_EC�=gp�`�F�[�q�ڼ���;��B�	�*g��S�\���cB�^�B�	%&�����ɸAf�KQ����C�R-B<�E�-Ƃ�S�	��x��B䉇"�@Y��H�q�Z�	�B�	�l��C�x*|۲l����ꓞp?�*�[7Tq����
'Z�
�M�<��ز,�2��pmV�>�y�UK�<��G> ��D�%ޒh���#7&]�<� <��@�Z��u��c�I��Pz�"O	#��m�E��Y�x28"O^���!ƺ{(���T�=�����"O�i���.VO~ipuN
�
��"O0�8��?C��cu�Ԛv��� �"OX���&�5#���E�;\���"Ol��&�3U�0�F�#Q�����'L��j��T-uU�%��$��_p�{
�'nu��ک&	>�j��]
 n>q*
�'1"(Yb�-E���p��;}�#�'.:��Lo�h�,�/	���
�']2�qQ�S,7>��R��B#>v5��'-  r�Y�2�����b=��'��T�ER( �c�g�E�����'�8�pG�]$�H�/ډ9���c�'�@ydjրc�5(� 
�6ژ�9�'�����&��{
(1�K�7*p��'�����jx���Ø�!R�I�'A��0e���1�cJܴ^�k
�'�bq���?o��A�/D�	��'#�82�բu��j[��rE��'n���R%�%-8P�S#4��M��'I:肵��`�A���Q����'aЍ�#�J�f�*z��{Ip�j�'������U�a'�89���'�J�pU�ۇ"��͒����Py�'扛�B����0��a��O��k	�'�`����/)8Nu���F�]r�'�x`����&5��8�wi	i��x�'\�IU��,<��
Ga��p�
�'�40��(�欈���-Y�n���"O>� #���\�Z� a�U�N�b�Ѐ"OLA����;<��@U��"���"O�Ex@OۯS���2�	Æ7�p�PQ"Ob!+ Ň�dƼy�7��6v�B&"O��0�͋3E��R��S�?Z.Eq"OT���j�.Q�p�! M�<CF��c"O�$���OV!��-A8VC���"O�ܛU�
h��ׁ܁"�yy�"O������'iی�B�JB�|���"O���JsE:��`ҵb��	�"OVQa!/V3Y���snؐ��D"O�!z2�^�@iA�8�EW"O0��\W���N֣�|�p"O\4�2͊I�PH�͑�2$�y�w"O����kIN�f�K���1"����"O��h��կH�摪�L�"
Z �"Of�0jB�H�BD��1L��"O�ġ5�K�k(|�5�ǯE��"O<�V�ۀ�BL�vhΧ
.�q"O�4XD�Q'F��]�GE>�(<��"O�!:�ER�[k0h��%�h�"O�P؂��}��(�e ��@��"O��ӨD�F�0�;B�!\k\�4"Ob�����g$�ɀ��ƳwbP��"O2��FR�`	��M/ICBp
6"O>�p'��jf<�0����U�v"O���Q��h`������9����"O��bG�Y/R����s�~���"Oz �w)�/�t|� ѣo=�|Q�"OX����Ro��tQp�� 5x ��"O���H܄?���"�܂F�� �"O��Q�kj�4�!ljni��"O>	��Ǘ�$Gd4)!��9�� �"O� xLSv��$m�$`�̌sDmjR"O�Q�ІPA$.U��`�A�� a"O��
ԅY9��I�E��5�F��U"O���p�Ή�$�JG)O 7����"O,��l���@� 7�ڟps��zS"O�m)���i4�٨C��3Pa���w"O@���H
8O`�0����wV|��A"O�!AL�b�2� �#P��"Ol�Ɂ����YeR �����"O ���@�)v�2WŁM�F�b�"O2��j�=$S* �%D�~��p��"Oj�����2��(r`�Q+&|z���"O���nH�}�r�b,>'_f���"O����m��l�Ҹ�0m��cA��I�"O�yآ$�:r���"A�T�W)6Q"O�]�6b�?C�irtj�{��"O�ܓ�g1@Z����;z��	"O�Yp�K]�Al.Xf�Ͷ_l�"O`D�d�A+�X��H�K���F"O2A��@�c����ŝ�G��C "O�mc0����RT9��?�X�W"O�L�� _wP����V�Y��u��"O~���cG��(А>�̨��"O�p"ՋU������E:>���A�"O������~�r��ՌƜ+I�l��"O��B�&Fq�*��K�(�t�s"O����&�:���R��B0@薍�"O��2R
:(��!f\_{B��"O��ZQ�W�5�H�{T��R�F���"O�1��'�(	w*�f^3]��lɔ"ON�	A����\jr(�"w@�8�"OJ��F��7k�6�gE۽\md�J�"OZ�)ićC�� �n�K�"O>�Eh�6����GVN,��"Ot;+ۏm��0�f�mATUR�"O*�	1ћ	��ԉ$D�(~3<2�"OD@�r�V�`P�H ���
}B^A۲"O�ez�Aۆ"��+aD>T�Ա�"O*u��(/r���_;|�,�d"OTdC��	�D۴@�YЊ�G"OL`�l>�����CZŲ�KA"O�lc7�	y���K�!�!HP!�"Oy*�S�{|*u���?)�5�W"O����� �Qs'OA�P���g"Ov,��͚� :�t�1/�T�hq"O��FS1RR���-W����y#"ON��Q�ݹ'��p�;,]�@�B"O�ѵ$��0���b�1��NB��y���*>��P�Mٝ`a��Y#J�?�y�F�9q�K?	:-�b/��y"m�:,�\$B�	�Ȳh�S"�y��Ůk�V8c��-��B��Ұ�y�`V9
��`g�{P�t��?�y⍎���s�M޹pI`@2@X��y��G�0^b��'u0eAp�Ծ�y��E$!���y��I�nC�|`�H_5�y"O���<sEK^"yp�UJ�����y��5K�1�DE*$��܏�y�%����l����D-�y�G�2	�,)S)Z52��M��e���y�nڇe��ԙ�	�&{�y�썷�y�ƅ�r�^X����#ED���N
��y���	c�
����c.��e�H��ybn�2K��(�R�# )*�fB�y
� JT�aC�'��]�$�M��\�"O��Pצ��k.h�'��6�D�"O�@���K���bD�Q�]�4A�"O�*4D�S�P;pe��57��04"OQ0r"۳;�jȺ�Œn8��$"Of@�RDG�  �c�$
;.���#"O��ړe���SR��T#"��c"O�R��M�T+B�۷���v�x�G"O�h3�Ά�< Ό��C	v���a"O�q8У�m���4�ӹ�p�w"O������>m��i�-E2���"OfQ(��H�/
��h��7b
9X4"OJ�ȷn�>����h�*GjFA�!"O@\�p`ۯ'�4L����& �|�K"O�����l\�X"�Q'��A$"O ���i��	>�1sRn@r��3�"O�<�1Zvr$�&�ob$���"Op`"���1?�� ��N�=K2�t"O���"ԓ0����F�U�ڜ7"O���1ŉg��ya+��d�Ρ
4"OQ`�L�$OZeZ��?u�!G"O8�X�j�pit�
���*Z��"O m���"Z����s#�wG^�u"Ofd�A�R�	�����
�& p�0"O^�).�
:s���(A�j. 4�"O�)
�"�V��4��&��t["Oޕ[�@-ztk���X� +Q"O���5E[�B����a���:Yb���"O��B�w����&���4I^H[�"O�({�"EJ��b��ŭ'���3f"ODŒ�o�ʴ
a�	h��ճ5"O�!+Ad�&Tj��BoߗTτMP�"O���[V�l1��ӡF�ȴ�"O0  � �1'f�s�V��&��V"O�}25)-r0b�x���)ax�b�"Oa��B�Tk`��$]���e"Oi�p�34\*�r6�P��L��"O��P)�-`J�y���]�
�I; "Oj�H��9S�i�(]���I�"O~�C$g�?�.�bB�<c�5�"O@���\�e0P����*r��!�"O��
��V>'��E��"3e0z�"O ؉fI56�L�EhB�0Xi:"OL��5 \�"#U�VG�B���"O�)C�D�dh��D�N�v�"Om�3�-4�0
Ձ�2�����"O�l���� w`�3��~��C�"O���'ר]M�X��`Mb<d����U�Oi�5˳M�<*�F0��hY$�� 	�':*(��DW"[`�Ҧ�X��+�'��5R5�"xt <+���m���)�'��$�C��9_��u��I&;ߴ]�^�<���.GĜ�����|�qa	�oS�C�Icl���&�nfn�PW \�C�	&9�!���t�hm1���)tWzC��>�.Qbc${���r��0���O��$؁Uh�h��>��iG�L7&8!���$2�ͩ��F{�	�T��!!�d�j�<9�fIA*LٰV�ʔL!�b�|pX�`�!����-	�W!��q�q(�D�6XAzFB�Y�!�̸u�t�t��/)_��(s��!��n8��$_%ANv !"BO�b�!�B?����g�>Om����C�)��y�)� b���i�
 �l��Ņ�]0�9z"O$��6L �w4X� 7 MA��'�ў"~ւL�Z(�ㆈoM��a"��y2aD~̌aS���3~e������yҏ͆/I4�ɡi�1	�L��8�y2&L�F��hs%�@>~�P��$�9�y"�T���Up��
Ǵ�aL��hO^��-�A���#aQ��8�J��h����Qa��R:Q��A�pm�%��d�'�a~�*S�/Y<��#@�f�pe*�#�yI,A(�qB��@12;���� �5�y�ׄ`,��ţ��M�����y��W��t�֪�"��� #j�y�q�lq4�R&�t��"����䓓��䓧���7��lCS+Mxb��<�!�D�]�^�oQ�[g��)��39!�X�Cx���tEҵ����,P7!�99�:��
4]^j��G!Xw!!��[>Cئ)�D曦L9�h���K�.�28O�L�OD���a��M>d�xP;�Q���ɉ@�
�`���n���c0$�9+m.�O.�d9ړ���\��{�;=��p�G��h���b�"O��9d�u�.xR"�2%�~x�"Of  ��΋j��%B,�Pљ'"O֡�#��S}�p�i�Ao�CE"OT�k��y�d�T� \QB�"OƸ�M�>�ȠZ"/҃PD�"O`����vN�4�_0O�NYI��'�1O>iIԏ)&���R�� h�P�!"O�<�N�5�\��3���2�Z�ju"O��7ȏV`�R)^�}��Љw"O�}Q��#�Z�)ι7����"O��(�FDoK�9�%i��2�rl�d"Oh� Fː�M�	�d�RhH��0^�(�	c�K���0�CV�D VJ���g:�O��9����t�-�WL����Ij�O���v
"?:���n���0���'�z-�ዋ @`�@e��{��A�'�@�"���!s�A:'�:�e��'�"���h� 9��Aʜ���'*T�Z�OЛ]z�M褮'�(%y���?Q���0>���I�&��ۦ�����C��o�<	�L��h}tX�'���#h�<!�H:'��:��."$<����c�<�s�Ƥ��� ��ȫ.�����f�<����k@�ڵ��K?���Ad�<���N�p�5��x��fh<��痳�0lH�B���^ ����"�?	��0?a$B�%p��|I��{?��$�^�<1�AE:w� %����]dyZ���U�<�+\o�D�6�F�S%J*sOƟ�$�h��	b�ܩD���>�䁻�F�2�C�	��>:MZ��p�b���(�C�	�Lɠ�BSN�,��,�G�:��B��BhyڄE[�LZ��c�޿`Z�=��lM6I��\R�����*~��C�I$��U�b_�d>�e��#�:uՠ��5����G��Vi�ь6\�E�&�7D��k��	�1^�Z���l���\C䉿=�@Y��c
8eLq�Pc��h;C�	P2|m�⡇�u����#_,<p�B�I�1�FH"AI�pw��1�����C�	)d���3KC?Z�Pr�/�C�	;Ь\H���
�|K��X
�<B�)� ��2e��T�<QpFI�`��Pj`"O`XK�'G	fA@�R藃�r�ڦ"O��s'mO*+�&tk�[(���E"OZ�� �O�v��zbgDiN�e*g"O�����-���f�?|$n0�"O@�z���:y�x�#�C�Q�LC�"Ov}����"�c�M	"4��f"OX���ڏ7a2�+ ��s"OB���V��\�Bl��#�P�"O��jq���	|�`{�� �r�����"O���Q�85�0���7(�v�����f�O�~U��dO��8���nD+G;>��-OR��^$V�ty���<Y�4:f��#H�!��Р/�����HއXWb���ݢ xџdG��ꗡ0��!�2�)���¶���y�A�I+�5c����x�D�r	�ȓӠQQ�t���7D�e�Rńȓq��q�@-�(1�i�I/��r̔*���o�p�XQ/e�م�	_�en�� �.R��0�Z*t�6y���u��DҒ~eP�P�J?X��̅ȓG��u ��ѢƤ@GB:{	r���gJp��O?�hz��J6n����n�jY ��F"Ph���J9K\���3 �4*���R�Š��M�;�4���3�,��3��>|/԰(S�6p�&����Y̓����AB�r�$�oΜm%\�ȓ,�l4 ��]fJ 3Q/@rZĆȓ'"�1։!DjPyć�=�č�ȓu����ѣ:l>	E^8{�Jx��S�Ĺ��"u!�� Pĉ	.	�E���MP���C�
�pq���2��ȓi]()Ё��M%.�I"O�(6�~���	M̓g�&M�t�D!�Xq)�
v6'���	)�J��V̊<	^ڠ��l��`*�C�Ʉ��)��7�`$�gǧ:G�C�I�^ �m��G��B�G�.�bC�R֜�1rC١Z|L�� L�/]q�C�	� �"�C'A^�aR��9�n <{NC�ɱ;�P
Ї�<4���#�_*P?.���n�'/�D�׍H�V���S�-	�J�XTb�'9��)0�޶*(�lGB�����y�%S�x��	2�m�p4�ks� �y��P�'upq;R,`p�-�"B�yҁD�N^�x��BkX���h��yR�4ma�IQ�'y��Q � @ �yR�P�}�8ip�K��v���YW��?�?a��hO<"<����`J�8Av`�%oL��B�q�<���P$��CH9��]cSY�<��K�= ����w���!m�<��J���˙�;�Xј1��g�<�2/̇a�6�a�? �8���A�g�<Y��BHҽz�;C[��k��Z�<�OT`Y����0����fT�<�78
&����'�:�M�S�<	�H�>n� ���
���2���d�<V�#j"R [��_�y�#jh�<)�����H����]�|��0n�i�<�2�� ��1��䝦3�֥0��N�<�DHD�i,h+�	��"4����Hh<Q��k�tU{���fq����y��5q��M�8Z^���V*��yr?+�x��� V�C�
�W ��y����!���RCY%�8�1�A*�y
� �I� ��;5f`h ܴF��u��"O�帅����Q�2�K"wd��s�"O��{� ��gp`�1��Ή(B(�� �	K�����ڤYyPϞb㖱��V?�?9�'r��B�$تkj�@
�KǇ	�"
�'ݸu�9!EP񒂦ލ}��'��{u��8��$��AƖ�	��'ۦx�n�b�<�����R�d8�'�b�R&1�Jt���Ӟ[��y�'�&���������ᗺU��Q�'��3�n_�q�I
���$Ƞ�8�'� 8r
Ԕ#F��q�ŕ���Y�'j����%�-~���[�ʹc�
�'�VH��)��DTJFeخ	$�2�''r8��jO8WH���B	b`%�	�'�>T!(ty���ۇ`RR<X�'�By1Ɓ�k�� ���Dך�a�'v��!��)+���`@�I���'q| z�G	�6����Gx����'8}C��ȼ8�h��g)D95��y��'��cDJ�JM�I�hD7����'Hm�S@�X��)�� ~��{�'����V&ԉ5�&�W+�/my<\y�']1H��f�T�\�gs� 0�'\ ���<S�5�&`bi恫�'�L;uH�l�$�(sEF�Xo�UC�'	D�����*$:�̀�&N38�h@�'��e���Qro�ec�3���O�<A���+)���dN-�-��Vg�<	��XP=��{aKӑm{ڝC��CO�<��$ֵ�]!�G!��mK6�HM�'k��'
>��E
� pJf�)u����2V�#D��2�D�"X"6�+e*�1�f�""�#D��hb��%�`�#L�'p_��Ct�"D���d암8ԌPP�k�zW|Ce.D����75lD�{p��,+�f�
�,D� Df]*AZ`c3
DB�j��?D��قm��dN=Q��YN�"��?���?��ɍ6]��	#Ouk:��"	X!�$ػq�θa�(�6NV`��Ǐr�!�	�<p��GD'PJXՠ�gǞ_�!��ڱ<P$庖�Q�,2h$:��M�r!��o�<Eɧ�ɉHC� q����!�
�T0i�&�;H��jE��I�!�G��P�ᔨe?4��b&�i!��۱B�� ���!HB|ɒ�'b�}b�',�$�0a�V��h��W��L�N�&�x��D��\@',O�mTT!��n�!
	S� 3D�h!m�.J�H��'��	��%D��;&�Q�#�AY����0#-#D�����G�;Z�����'������-D������2!���%m;cî\��*D�xQ����e:����2�t�;�,(�O"�I�"�.D#��� l�r��A'�/�D�O��$%LO�T�wM̚Y�ar%I�$��"OT�hC�ܷR~U���谡�"OB��g�5k�.�"���4�f���"O�}��� N�����L
:&��t�"O*�C�I�c���l��#�F�	���:<OJ-����>p0�7��;Z���#��)D��X�$�`�����քΜ*�E(D�p�����U�`�H���f���y�o���P�RH�9�&�óg���Py2�&v��\YA��]�~�9/�x�<� ��Ç�f/�(�FYK�9�"O�05n�2����Ǥ/RPj�*@�"LO�-�j%P\Q��M--l �Bc�'�!𤁳����HJ �$���X�!��R�:rb��7�;+�v����ؼ,�!���Թ1�BӰA�����<X
!�$Ɛ+k �q1��=q��d��'K�:�!�d��mp� �Q
M}P�����Ae!�$�<ywr��tcH5���&�IG!��۰����cb��x[���t��_�O�� �b�آ��?'�)�A"O����*@%V������4Iq�)5"Oƴ�J����ׁ�J�6���"OD�K�Fدn��yk���<���`�"OT �&�/�C�j^eB9�$"OP���
^6^|����g�܂A��<���U&w���"BO�Mn�����i8�B䉝E2h��\4� �D�� @B�	�;34�q"!eFpq��ڒ4-�C䉚0l��dH��w�"к��Z�4��C䉓&�n��$V>;^& hq뗊%B�I�LC�=	�c
 �ʋ�mC�C�	>sӞ]1�����B&���>���O"�O:��9�'.c�˅,��iM�)B��8H����J�.�3E�,>�h�a@$�H�%����ɤP0hl*��JNB��g��>R}�B䉯9lt0��m_%�@CUMم+�BC�3/�(��I��`�ħ�3bNC�	�a����Pʐ���%A�n��B�	
�)�Q�K�3��	���R$M_���?���)��6`^P�q��B��L�!�$�"S0��hR+@�/��(
��ɫH�!�D�l>��7��J�v���M�9�!��@�ش����R���:iH(�x�'�2aZ L߸[s�`�l�P���'���ZE�� \jbgݔF;F0*�'2�@x%!ǨuMdb�`��¨�,O�=E�Θ�*X�S�j�b}�@�2�yra̎*�Xk"b�x�����yN�	!#��0��q*������yb�'�����_�lɻ��
��y՜e�� ؐ柸I�8���A��y�M�`4����'W�<�.��dE�yba�=M������D����T�U8�y����ĭ���	97ft��3��<���?�+OrP���j�V��u�JhX0|��8D�`˧$%P(��l�x�@��6�6D����
�.ߦ�c�.�Ȁ`m8D��[���f�^���g��w��c6D��C�(��q(�̅+�5��4D�!A�D 32�H�#`^�MZ�7D�����������&�����p%�(<O��d�O���m��(3$�	���Ǯ,I�ܠ��3D�|�jH�/eRl�'dءb���ئ�5D�, g�Tur�x��#�<j��.D�(	s&�t�~�1�Mx�� �$�'D� Yr��q��5�2.ʲ2�j��s&D��"�K��|�hԊ$EL�D���!#D��Kڍ6�¼����&B hWn4��?i*OX��u>�k�.\��T�J�gir݉�B8|O�c�d�.�;X	FTrgL�8�Q�7D��!H�')���p���P�0D�Ē�+�.|!��E2�q��:D� �U���4�̺u��G<�`9Q#8D�� �4e�J� ��!#R@�	E�t��"O�%�a�6V��#��n�()�p�',��dE�.�B��ד4,�+��C�s��y��'J1Ox���a��Κ�Q�!�G����"O0tE�b�F�H�ש#���u"O^(�S�Z�3�:����4�i�"Olj�L?A�X���/nu���q"O���Аq94��u��+w���	>�r��>+f��a��Q����%�<Q�P9=��K�V��I�Ԣ�-B~)��	]~ra ���TM���c���!�y�#�fmD�@�c;���@�-���y����hW%�`H����B�y�'ɞM���'�|Pqv�I�y��f�H ���X�6���f�+��x2
� ��@P6	�>V^��&������R��'Mm
-I7��I��0�O|�=E���#���S�G���n��6p!�D	8X�q2w��}O�����!�d���8�x�+�;T�j���D�!�$B�f	Z�!���vB�4���ھ.�!�$Cr̀�^QH�T����l�d��ȓi����M�;=�v���^�����b<i&n6U@2�Y�TH-\�b�A�Px��'K�\�(O�\��H˕�4Rծ$K	�'�0���
�O�,,b��	{���"�'~����_�#�\�xQ�ųk��[�'!�Ӧ�4K�VE��%�)1�����'ܠ�D�%���G��V�`��'֎�WMB}�4,���Ք8bh���'�Dq�E�0�\�˗bQ�E���*�'\����R4Y~�
'%P�I��@��'!f��T�
���mӆ�	TZ@�p
�'�ܵb3K�S�tY������'��,�we�%q@��2-Άءr�'�D7a]*mS�K������Mg�<��捭�"��nΣM�(�*�B�dx��FxbeP�Q�*�p�d�C�4��Ь�y���-A暵@�h�K(4���NѠ�y2F���J��t��6B.�qe���y�!t�Tpqu�;���#��R�y�0�J��3d=�''���y򁕾>���6�N�/�"$�Ħ��y��)9\.( �bЦ(���є�J��hO�&�u����¥j�И����(2B}���t��p��K�������N�*!��>�z�0䯇q\,xr��	k�>|��)�65���-5����Q�<��(�ȓf�P7��a�r���_a����C�P�S��U��ń� ���ȓ\��;�"#O"t�8��9]K����s�'~�Tʱ��M���Á9v2	�'��@[���c��P�˞�1�����'=duJ�N�?�d��%�Ȓ(�fԻ�'������
H&�\�6�T�'�
E!C1��M��!ѳ3�~���'�ƀv��j�l�U�2����'��%��~Z�q��Aǐ��'t���p��1F��ܸ�
�p�ԝZ�"�'��l0Wo�	K��R�*�	@U�j�'�TI33 ,���/=� ��'����ը�$8¶H�aS2Q��'�l}�(��A{����F�+)R���'���s�
ѰL�&Ab��7�4!��� Zd���H>��$9�"�8|/�yX'"O�m��O�44@��eb75 2�#"O `�I�<%�B�!�,0�
�R`"O e��+>m-�T8�۰VB���"O�bނ(�~e�1���hD�E:B"O�aq�ᕺ*L c��!L���ac"O��٧�Y>t.HI���d�I�"O�!��F-0�A`v�J�/�d���"O�	�SE�WF $��@ ]ϔlC�"OX�t�:~"^�	���zR�xX�"O�		�Ȕf�I�ą�TD�$"O(ر��'N���h0G�m�V"O&�����3�ތ��'��5��	a"O�-զ�3~���d[>�=��"Orm@0MPT����Ɛ[�8�q��'���'��C�<Q V<���՗.�.�"O&�B4.�"d��]�N5E�\���"O����f-��ԡD�S��<�q"OQ@���-f\���}�=[A"O�ГF�ۃ-�V-1���zv�(�"OHP�E���d�	�}�LP�7"O�j$��9V��	�"������D�'���&3�|Tr��	>g��ŉ5B$k�RB�ɥ5KjarF��7�0��7�ƋME:B��(v��X��ǬUx�	
ʼ/޼B�	
e��]qA��D�l�;��M%2bB�	*JȔ��OܤD[���V�-/�C�	$9�c�a��tU˃�Z��C�I%i��l%�66��t
�c�C�I7P�(�x��1���i�e�(lC�	(z��DA�PY�M+F��s�
C䉳N8� ׏�ID^��4�L<��B��=�(`���!`	�b� c8B�	2ML�X���n��p��˛B�(��� �m�q��I�O\ĲB�I�<����$j��:p)τ&�RB�	�X{@��q���l;����D�JB�	�W%p�p��OW&!�wj��8~C��;/X����V�" ��x�&ݲ)�NC�2Z��Hʤ�29�X��� �>�dB䉄f粍��i_1|@�1��%M�JB�I2@ĈpR�x�`��N���C䉌	��C�㙎_��pG��:�O�!� ,��IZգ�*a�@!�"O,L1��H�L���j������q0"O(-�!� y�t+saU�?�`�"OBT 7A�3�9!ņ��Id���6"O� ې�Z&F�|���j|�c�"O0�+�k ��ؖmC&ji(9�"O�9�t	�%?F޸�wJY�W����"OH�!/��#�����9<�x�
�"O%kѾ�Ҁ�L_�'�B�҆"OP����~1�]rb��6d���c"O<�8�M�frP$b�7��e"1"O���2+)[Iְ�e��F�h�ic"O� ��L[�_o��v�$��y9��O.��)^.�<!��f۬4
��雑G-�'|ў�>MS �,!�<�G��G�ġ��"D�0��U�wg��inȅEx�1�W�"D���F�.5�J�Z���KoF��7 D�
�#�qvҔpAO�0��2Cm1D��a��R�N�0d��d��e:D�\ E 
�2&�ܣAe՜�Ԡ膈9��0|�S,�.p���v��*-��A1��p�<� |a��.� Y�P(m#��_,$QH�"O�e�w��~��A��	��\�X5�"O���OҀzѺ�s�I���|��E"Ou�e��J��AӶg�"�F�v"O�����^<�)�%��Pb�"O����N
�i(�R�f�� g���OȢ}
�'����fV�>v�"c��,F�V��	�'�I�e�%p�\�ڷ��R�NP	�'�`�)�6|D3mZ�S ���'F��D�X�??�$�anS� F�{�'¤Px�օe-���G6��\��'+��#ER���c�]+hh����'clL��N��at�$!�Jh�$�N>����	��}�����R/QT�����]�C�ɠ6e8�u��*'O&�oM1#uC�ɰ�:��隃Z����Ţ�'	,C�I
��$�Ԉåy6ف�1�.B�.����K�����+��� B�	�5�ޝHI8��𺧊���C䉟{/�qp	�� ���.��: C�	�g;rP)GT�<^���C�"��C�I�vH���܀V����.�:�C�	:������ ��u	�G!=��C�I1�F$��A�	\��yITA�	>�pC�		 /y�\8�BAͲ � I�"Ot$;A�Y�(�Ri��� )R�Z4(�"O�8����s��jD��S����"O�j��C��Upc��F�T�¶"Ob$@ņZ�+{���7���s�"O�p8���/�"a��a�~���f"O^ ���Yh����A1�X��"Oz�33�@	?�̨֠Πq���0"O��xe�Ӣ=����[��dH��"O�P�& K6!�f�C���'���"O���RhơD�0�%�Z{�v�r"O&�`���DE�ݐR�W����i5"O��sc��m��`��k�|�a0"O|���oH�#²6�k�V�P4"O��5��,�(Hс��![��jG"O�;�G84[jp#3�(X�Lpx�"Ox:sK[��y�Ҭ˴/���PW"O��ۖ�+He��H&aşB�HI��"O��F��
K��Ja@��-fQI�"O��ɦ��y��m!�	Tj��X�"O��Y�ϋ�7����� 5wm���4"O��J!k�5dP<��6�Ҙ o~X�'"O�����X	l����X�RWּ	e"OV�F(�	l):�yp��o8��"O4��#i� L�!I�R7���"OTܻӌ�o����R�j�"Oθ����O�Tl0E�O3M��$��"OB4y��D�@a��⓭H2]}�5��"O�l{�E�:N��T�
�Ht�"O:p�ᄮz�ֱY��ցzm����"Or|{/0C��Q�`eF�V^��"O�<i&OH�F��l��dM�Zm����"O��S��:VlN(hA�]dy*��B"O$���'?w���7c���S�"O���G��J�{�C9G��pw"O��C�l_�pQ�!E�V8P"O|�4D��1[�m0��>G�l\�"OHL�D�2I0N��e(Z<6����"O"@�I֨0c�0�G�5�2͛�"Oj�Ó�S(_��|�g薌}�j��b"O� ̼ہC��@�����P���5"O�erc+��H,�h��nuf�;"Ob�(G*Z�B�!SG�;v��H�&"O4RB�B�v?xT+wa�)N��E9�"O~]�u��<B �@�B�����e��"O��%�K�J��5�@��s���"OR�ò�ͺ�V#�$ٙ'��T�"O�1p5([F�Q3R���!�bh5"O�8f���v����^�2�fL3B"O�a�$E�u��H��P0c{�9�"OB;�B�I�^ ���A�|n!�`"O�]*&�&W���!�F7|���T"Ot���ڗlT]yJ�	_���"O���`����sv��g~ʈ	!"O,�ꡧX3���`�5fdi!"O��ӡ�<
������0�"OHp�7��,m,��KDa�
2���"OF��%)r� �bn�_!��r"O�Ea2��/���pHѵV<�k�"O��ggĥR�y��T00�8ل"OR��!��uK�aR�2� ��"OLPiG�K/>��1�v��h{1"OZ�+c��(.�x� r ��-��yc"O���׆��tq�H/%i܉B"O,}��O�0��Aݸ:b��"O��&ˇ.**��X�Nx��8
P"O����bP�R��$���9R�[T"O��:$��8�`��nRE&�B�"O���V'��C�vY�6LY/Yjir�"O4p�2�� ���&Ő>�rM��"Oʁ	B��)��f؛�����"O����m�*4%��Qr��D"O`�%��>;�(�)��q|MQC"O�t[��pe�lZ�Bap�b"O��qI)A L�bR�A�5YNpI"O�	�@�Ψ[���p�		�`P�<3"O�4k܄�(�(�M�:$s�"O$�P*ˆ\��#6�;g"�Z7"O��Cb�f�4��)���"Oh]:�bB�u���@��4)z�\��"O�E�iH=(XHXD$�w���"O �Q��ԥ`�d�Z�BWor�3'"O���A9e�(Q��Ã[Eę*�"Or �AJ��xIk2b�>���1"O� K��܊dvFUS���Z�
�Q�"O��{A�G�
�R7 6aXݓc"O�@I�'V�fn8|��h�fCh�Y&"O�i
��̨<��!���'���8E"O.(��ƙ�q	͓t�ZM25mV�<��)Wg�
��'Iy �i*Q�KG�<Y��dۂ�H'̖�`� j�CJ�<	A`ѕ�L��0�{� A!ƌ�I�<	׎�	<�p�Y`J�h���pR�WP�<��j%'F�a���6<�p$�A�c�<��ެ5Ta���ư*Or����^�<���2*�<#��Іq�0���]�<-4D�x������E��>��݅� .�� U��=3��K �=l� }�ȓ9C���p�v ^�'	=*`~���z&���ꀠI�8���T��5��`����F&������1>I�ȓf۬�I�Ý8S�YX�M��3�l̆�4Y5��g�Q�@�U
��P�ȓ^(e��l�>A��K!��|v����S�? H%j�_12��Ǯ=g8<�!"Ova�%.M&QHdm�&~�`�"Of9��$̹n[�[���5&�\4��"O�,!�,��x�\�r��Ou����"Oh���C�+�(1����-Ga��"OĜ�(�3@r\��f!1?,Q��"O�)��S
���B�.k�y� �H>�y� [�i|�@�#�ɳ1 �1(��B��y�-׆"Jv-��&�%#��a�g�$�y��H�9E���=�@�2e ���y��Y�j	��r���&4ZD�4�y��Υ*48���̷M8ӆ����y�� -s��r�Rx����fl*�y�h[@�"��?f=}1�͘��PyҬX��"�/��+v����}�<QcC��v�.}��W �|�7e�<�P�.�LH�aԙ4s��X�z�<�b��@(�5Ca�`�ؼ�0�s�<QFA�f�����4���T�l�<�sc�]�
,�7e�6@Le;"�D�<aר�o�t���/G{����x�<	C�r�0�S�A�)ɨ��o�N�<�-Όa��dإ`�	!^)�w��L�<Ad�U.6C"`r iO,zL��͡"O��K�)��X�T���\�{���;3"O���.8JM�a�QA����4"O@t#6M���e���y㴅3�"O$P qb��d���&g��3�"Ox�"�NXq����c� 8N�`��"O�ع�O�f�V�Iv��:s0N��"OQ�����_� ���4&��@2�"OBb�L��ʎ��s%�y�ДA�"O�AW�K=��$1��V���#u"O~��2�W�$^���*�F])�"O����C&+���x3&�Q���2"O&tBJ�@�\�����d�� "OAc�DS�vD�a�����zYj��"OR����2W,�r6i�6}tŘ�"O��H���;�������/Q��|�6"O�@�e��/d <9PN��W�^%pf"O<{���25�Pa!��+���"O�m��ބQ ݛ���	;@"Oɛ�e�"z��nȳ;$�
.D�L!Rh^�
���J�I���"� *D����N�$V����i�8Y}��R,D�P���?^�$yA�L�YK��i�h/D��q�� ;|P%cPJ�"A|1Bƃ!D��S�"�7ό����
�~䙲!!D���G�R��X��o@�_��P�M2D��)��3bB��:�X�'
��s�<D�4��	��`�=J�.�F����҇0D�h��
�9���0%��f$�jP�:D�l 7i�fY��D'}�"��
8D�x�w
[�9�d�#��V�X��B�2D���%�,.R�9x3���BD�%D��A!F�e8Lm;�ܳNJ�P�*7D��[W��*V]��	?$y�f4D��c����
�h�ԇz�BHS�0D���L�nf��C�)g>0�9D�xI4M�(�ZQ%!4�4Ԡ�);D�L�u�>l=^9�T��<:��=D��ფ��`����參#OV�B��;D���yz��G�+m�P��Z!=�!�AT�n�bA�H�F�`�G�k�!�� l��$8�؀H�I�u
x��G"O�yزl�L�b�2cbŨ\�lXZ�"O�	ڂǐ/5���K�NU�����"ORㆉ
�\�#��9�Zq��"OP�i�Z�N���{fၜ2��8�"O� �reW5d��`�2 ��ə""O�8@���7_����:/n�IQ"O�����I4)s>T��D�Up�"OT�Pb)��p��`s%��).���b�"OZ���^�^A @â��]>µ`�"O��-A7���sdj^�;>.L�#"OZ�x&%ֿ"(�UH�Ց!�u��"O�� r"܋,w�!�b:a2""O���;z��AhC@�+'hHy��"O�	Ñ@H&C���YGl� (7"O��	>Xx�ݩ�
,V�!�"O��@%�}�l�2ǩ�H����%"O2iѓ
�QdrHo� y���"Ohتk���`�Sad�xcB"O�� !��C��=����)y$����"O�1�v��"TO�X�EƟ8���"O��x�O�=P+�-��d�NS��#�"O�K�I�U�Yb��6W�XPA"O�yC�m��}�Y9�C0f�̐�"OP�Mu�.������D�!�O$A��	��=�n�R�=0�!�ćŶl�(=��Lz���c+!�dO�|��0Y��A�\�$�U�ڮ7!�DP�Yf~HYB��L�����*|�!���-ͮ���ڹ5��C7韷4�!�$�#Vޔʶ	@�������q�!�d�9����NE���GXy���ȓk�çG�k���sUF�3~v0��^@� �Қp@��2��N���by����L˽eh���b�t�h�ȓ,2X-���K4�F�t���@W�=�ȓ�x�f%�in�1D1��1�H ��C�MXz0gb����ȓs�����T��s�_:Q�漆ȓ��Q:"�GE&�JSL�Wl�	����9�aBH;�v�j D3uGJl��(3�U���Q(	*ʄ���j'�,�ȓ6�T:�P�v6L�aAD؉�����ma��1��ĥ�L� �⓯k���ȓ3��UYT�E�jr���l"aI�ȓHu�����b�r�@Ճ� An6�ȓ�tC���&��,�6��%����iJ����p����#@�8�ȓ*�{q%�
(�X�Y�,Ҋg��ȓDؔ�fG��9o��	�I�w���ȓ2�L��#"Ҩ]���#� (��1��q�I�b�
�6NZ�]Q��y�H�j�4e
BIX�@��i�%���y��M.bI���IΑ6��l;�MU��y�B�?8��E0��0Y0��_��Py���& ̌�U��!<82d��k�<����t�R\�v���h��H�H�@�<�.��yM(�	$H�f	ԍ����<QD��7d����7](=��MxG��<a�9P���a ��3�XM���<��@�bZ��ڶ�~:� 8�Ib�<��7�f5y"�ʆ�``�w��C�<ك��z���UF_)f�����B�<��OI�S?Ftz�$�����( �<� �2���7"{���-5��ɘD"O�5�%M��yk�Ey�픱}����"Op�XQw���0��7�P�зCK�<� �63&F��+��F�X�+^F�<����6+KP��%ʱv��j��SC�<A���`�ܨP0��-B�Q���x�<yu`ǵ65�8;�k�7ozpr�s�<��բ.�^h:@"��x�z%��F	p�<�N�8#�
�a���qK>P)C�Pl�<qQ
S�&�>���
*(�F(AT��e�<a�䔬h�N,ӲKN�k��5j���x�<YQ◈TvL#vO�0�t���J�<y�hY�0f�0E+?ɰ��s�_�<��":�~y�6jT�9�1c��B�<y�ћ5�����?{�:CD�RI�<Q`�זs09h��ۻc�Z�cJ�<	�)jG(��Ĥ�[`��M�E�<A��^�r%��j�$`̦��
Cx�<�$�P�7�űwGCJ@�	:��t�<qe �>2l�����/j�1!��q�<�b���=�L���F�	æ�I^G�<a��I)pr7j�2C���;"�Hz�<A��� �P!���{@|���y�<Y�/�$ ��Q�((6�p��
Ns�<��`� (����2X؊z�<���ѻ>��� V����A.q�<)�nۚ$�@�#���:3�=�2"Ml�<��J M �K�
�1]j�C%�j�<���04BD��qՑ`��t�w��d8�,Dz��P9S��|:����HMr�Z�D9����]ןlhbH>u�X��Gğ�gL�d�0D���rb	!V��"$H\=+��I�#"����Ԉ�qfVn�8U"7Y���)��d$�S�4m�4�+��м��x��N�Q�&c��:��)�ɞ�T��lK��G�\�\A��Q���	�,�F����������G�18~��=a	ç2kR��Wk�9S�捹��ʖth���In�j\��3���q�u	��N7��X	�'2�-P%bB��Y��/�:�

�'�,%Iu�ݻN �L�pI�,W����'�XC�d��@rXq�w�D5q���'a`,�Q���F�$���D!f�'z�b�6+�����((b��Ó�hO��ە�T�b��z��C����"O�Ԑv���?^��k@�.��䁰�'��O�q�5cW�4�ha���lk'"O���DD�"A��@-��(��L���d#�S�'Or����AŊ+�F����H��@��t�	�v��)��M�=nL�ѪIkQTC�	C�٪j� +���bh�:v�0�Ў}�9O?��@�4<$a: �P0��!���'��|B [�O�$��-]�q��,A�� �M��""�O��ɮu(���q�P%����q�B���B�	�0�VXXbFH�n<����*oK�"<�ϓ|���*�� �A�2�ߓ/tJ�?����~��.0�Z��`��'���ŦJ�<q��a��p҇%�Q,�)C��H�'xa��ۓRt�ؚ�ѧ<��L�%�H��yr���z���g�9��r%㊔����i2�g?ٴLǮ	xP�𓭞�Qr��Lb�<ף�.Z���!U�W�xQ{iߟ���a:
����Qv�`� a�=E�
܅��*Oje����#�%K��(5��"O�����x`f�V�;��h�p��P���� JTa� «A�*h��._T��$��"O8�)Bn�k��4 3��)/��ps"O
%��2E��ё"�H����B"O�I hä{|�k�G�/~Ɯk�"O*��f^j#%�%M�jaV� 4"O���!Ē�A�b�H�!Z�J`~�Cd"O�AC�.���Ph��6cHm�!Z����	�H`��%dM:��E+N3<C�1*�l@Z�c&^��Ȣ��O( C�ɪ%9֙Bs`�f_�l3�D(>��B�I4h�vm3��9,�9Hÿ9T�B�I�d��k�<I����
���B�I!�p9zs%�P��8�C��iТB��3
>>dh��g�֥A�EL�>q,C�	�/��B�L��Y�A�%a�B�I?m�Xӕ��(K�>�1ҍ1�B�Ik0xs����< 0��"�*�B�I�@0���ҫ�vɸU2DJ =+"B�	�I%���W�dӔ���+Ӻ"WVB�ɯT����6���R,4�2B�I:#p�[Ǥ�>T	P'-�F#=q��T?MYЎ�6�`�3�G��j�脋�-3D���B �V>�;eg�2����b0D�� v��I�&iX�)\�%�����-D�l�C�S>
�HVC�#mZճ��,��G�� ����54
5��H�P}���$�p���Do~P�Œ�Y�	H��Q�C�VB�	=k�3�	^2$jr�䏣��B�	+E�� ��% �Lp��K�!e B䉚2�$EK�C]�$��S��h�B�	&FU8,"4���Ph�W	�"��C�Iu ��k����[�f�l���'�b�9 ��L�"=Iq�͐z@�k�'e�Z�����,�`g�M6zAJ0:��d!O�8��Aӕ|Y҅�vh�21�Ri;��'���I-.�� 
�;}<�CЭۃX7�*��T+�'pU��Aa�4v��Ij�,*��m��>��]�jh��I�l�)��#D�8���-{�d�sD�H�c�K�
!�DH9 X$�1�I�C�U ��[Z��p��H�J����N	=a��i�g�-R~MHv"O�Q�ƾ��{�@ç6\�!#�x2�i�'��)��@>C(���'t�9����;�!��ɦ�X�Z��޲�t�L+�Q�Ѕ�I2c����`���Cd�� �nC��#2������Q�vACtc^�Q�6�F{J?p㟅-d�T;��Y5.�pu0D���ɢ ��	�YlY0��*�I�P��}���j�݊��9��D۾vN�㟨���5C��)!�͘5�niY��5N)�O�3eO�R��z�I�&�
����'�
�1�y�b��o���W�̏K�Ȉӥ���y�G18b�K��ՐAxU�t�����hOq�:u��ܽ	�b�q�߾E�Bds�1OX�	X�S�O��s4gHG���7��:d�	�'���SL��e�Ec��+R4]r�y���żE��aR�CA�3Y���g���g�!�D �3�Rܨ�E��iMȭ�vE�&���	�O��?e�vΌ�Y%z ��Ƿk`J�['�+�O Onq�1!�#/z`: ㈅e*�@���LE{���ʵL���`e)�51��c�
�!�D1��|�0��>�ɔB�,[�!�"8���^	5!"h�s G�Q�xD{���'� ���� ��;�`N�0ؐ��� ��ϟ�ٰ΋8�p���OD��d�:U��у5L >b,0������!�Fc�"���
�hd�y$gM�/r!��N�#���gc�el89"�F�$b!��P�Z��w�
Y�DRpD^�8Q!�$P�-����G]�t,�Cs�R.,�!�D��d�xx�%��d��9��`8A"OHm9�&^&|��0!%1w��#�"O�Y�GZ�%V�<��cҡ �-��"OJ`5�,WuF��c��rwĔ���d<|O�T2@��n#��D���ZrL��'|�O�I�q����U挓?tz<��"Oƀ����CJv��*~bD�1A"O�Dj�;{ŸE"OU6�U��"O�A2�ܠ8���dҖ���e�O���$�[����"π�hp6�]�i�!�GCh�RG���H��4�^&Gl�O���d_*N���Zv�7C�n��򩀏Pf�zb�$�~<�*��\����.$k!�$]�8Y���1�&�a!.�h^�'���)�S}C��h��C��>9�W�L�g4ZC�
qc� )ۢ-�(�f�I�NB�u͂4��]fi.0�c'F�U��B�I)N����)J3R�d[IrB�I�dIb����
p����B�Ɋ��}����v�zKJB� SB)r���+1�\��a�8?�C�I�V���⇆Ғ/p�1�>6M�B�I�4���V�@5Y���.B��6�2�S��M����Dհ,��a�# ��rS�l�<��%��G�r�:ѣ؆5�Z�{�FR}"�O ��DQ)E}�$�&��zZ`9d�	B!�nq�A�G��+)���(��L5b$!��}�E�/�@E2�eƁ!�ҖwI�T��E�2��:p��#v!��U�O���XV͑8�
i���0t!�]o��ЄMV�37�$�a�Z(�!�$F=~�]�p+��I�L���
B��!�	7�r@D�͑&��i�ə�!�� 	$�(Y��愪l��@�U)XF�!�C9-�DL���N�Pp�M�#o�|[!�DO�*�I83�6hl���5T�!��S���	C�.M`<����,�!�l����/K"D+�4S�g�B�!��B2u��x�wŃ�I�~�# ݼ!���,J������$k��N�)!�$�M� ��`�޵o�V����f4!�-7IС�F˛�s��\1r$]�^�!�C-�tXk4#�o߼���"�!�$�Ht$�{��C�1k M0 �V�z!�ӕ��5���B�Q�d`�4��=#�!�dҝ(���bۚX�H�1�"O �y��^L
 �2w�M���S"Ot:AN�Z<&�:��ȑx�J�W"OX�A$�M�cBd���%
96�� �"OH�L�=	�|@�d��3�M�d"O�4`#�N�W��\����(Ft��"O`��˪G���wɋ�QZrIX�"O�}R@��[|D�ZD��K��A�"O�Ert%ÜQ����	�&?4�c`"O�j
�Q�<�����X,�"O��ړ�D)J��]��'A&Jx��b�"O4u��D��t�%�p�ƽ\j�ت"O�5 Q��+p��6����0��"O� �h�CBҚ( �Fƞ�A�%�4"O�]�@f8y���ǯ5�D�p"O��Ӎ޼V�P5he�Ѝg�JP�"O@�e��1&,%"  �P6��87�'��y����On�c��Ʈl��2'H�#=[NK������'7a�é� x�m��c��f�!�'�)���;&y80L�a2(�'�\�a��e`d GDƢ��ȡ�'��-b�)F�cfp�v'Z�Elmb
�'�	0�O�f����g�"����'�����IzQA���f��1�'�8a@ ²>�\��%�K�I���'v�Ag͔Z��[P!�:���'����Ed4��ǣa�� ��'�� P�#R���z�*�\�l��'�"I��-�"P�e�V�|Y��'�:�³8U_�Ȑ̍�L�D���')H��<'u�5R��
m���UD>D�@{��p��yk�dB9ʍ0$;D�T�%&Y0��, r��/m��H��
$D��%��
$U=�ue�"f�l0*W�(D�x������&�@WB�=ʈE���'D�z�G8l�����*t�����0D��
%E�X�4�I4(D�J��h1e,D�Hj�HǉfwzTɂ!f�n�0�/D��� �ě��d��C�VFpE���*D�W�,v�2=�p͓�2 H%b�@)D�����
�Y�dU��Q�t�� ��&D���MEa�	I@#et��Ȓ�%<O�Y" �#dv��]�6��O.�pd�'c�:�t���y�y!TT�8
b5y���A�*�$��z��E��(E�1�S�����Cᙃ5<(�B"�^�8�C�I�'2�΂�`#D��k-�����>���������L>Q�NK8_���l���A{�
�(<q��&+S&�;���ZL����h�t�I�%�� \��{%n����\(=H�D�@nA�Y�B��>p������ �l�'߾e��on�P��ׄ"H��r�'�X]p��C�?E�l�7"�U�"��K����/E��,uu�k�OC.�#�!�!�����aˁG�*�'���&��"@����` /'�[���*l':˓ �� C��8�3�S*�H�h=RP|Q  �R��d��Uq�]H���N`D���:�.m��X��
��D$�O��@t�U(a���#0��¥q��'���K�o ,>h�V���o�R�HCP�ϰ?oH���.D�����K[U��c�G<Z��]U#�䐏z��Q�V*����$yaD˓�n4���^<A�D�U"O��`��6c<L��/��y��X��	��'x��H���>1��I�~\��� �:�<����Z�<��՗?� 	�g�N���W��~�<	B�^KD|8֭�DziPK�~�<91�]b�$����E(1�u�<���ݦ��y傄���"�n�<����%��D�D �6d	��n�<�4�ŷV����)R�W��J'��M�<�Z�Q��ZqNH� Mn�
��s�<�EeZ�4g6ѺkߵD[HҡLJp�<��ǵr�\�IvE$R%hرvm�<q��WI���`L�qt�����j�<��ӑ=�!�3"� �2��ЫR}�<���@
��S����wm�[�Hv�<��閜dV��*�L�:��U��[�<�ۂ C������|g��RK�m�<	 �ՉM<� �5�^�@IޜH�
B�<�U�C!#7���4#Y� #�R�<� ŋ����K�� c��D�4f"O�MbPo�5#�8ٙw���&�\��W"O숹u�Ǝ)�D\A�ӎX��e��"O�Q���n,�� �!�:��"O6Y[QHE=󴉱���|r\{�"OƁ��B��P�Bn��TR�"O�ݪ�A�DXh���{�4�"O�I!d*J:O�L��Up��W"O����+I���˓lD�"dh(�"O�DK&��(zhT���ƻ��)v"O�PPk4R�� "J��h3"O-���SqӺ '��"��K��!�DP	P��5(h�b������8�!�DG��h�`5���QةkgFW qs!�M0w-xyr&��w�\Ѫ�e2k!�DY>�8|s�d��\�JE։Olb�{��Ԅa��p�'yJ��F�җ]w�����;�
�B�'%�4C��9�h&�	>=�<Tc�}���҄ ��pR�ؑv��?q��Q���0(��C��
P�j��*U͗U"Dy��$]�S�,�fɀ�S�x1X�Oأ|�'���ǡ>c��2P�ϲP7:���'\t�u!�2
�\� 	̰_XH�ҀE�]f�q# Ȕ	����ŔP8��hv	%b�>�� �M�Rn���f(\O2TR�*�]m�1RB�?[�0��%F{l���� ~���%���x�%(_A���� �NM,�!K�)��' ���%��*vJ�J�Ƶ,�|�|R�c�g�R�ڧ�G!01����ZX�<�� _f��<�F!S�S��ac1CȚ- �16��h*uj�o�61��E�,O8�ACT�p'�����1��C�"O4P.�$1ǈ�0�jT�������2`BӌI��R�R�l�J�axR�E-v�	b&��:�JY�����p<�Y�c�v��R�Z���������'�K�bM.��s��!�����-�P���@�A�����"~i���;?!���G��(���6hpH���67XHT�|Rp�H72�֤��Q�X��E��r�<�1��3r��5��$oj�\xv
H�q�53wk2=�n\چ�J�b����|���
G~,��,���e�Cˀ�2�6�xB�R8+b��g�
|Njt�C��m���Ф��my���5�q�s�'؂v�H"}�:�3L�e�Xm��b@�㥩-?��-i�Z���$H�q��	s&�;KJM�&�%$���Gh�0$��k���SQ��xQ�=?	�Dч���"|ڂI�??����g�DK��\�<iw �8Ze#�n�1ǘٚ��Cܓb�d�j
˓ּ���`u���S�A���0�ȓ:+��h"+�?An�K���1�HŅȓ>n���aP3r2���F�vNɅȓ=5rMB�kw�DIk���>�Z��ȓy%������ ������� 	.h�ȓF���҆�8������T�ҥ��-ƨKd�ܠ�B�7�U�_2�ȓs	����H��@i?
4T���-2N ˑmZ�{��))2h9Jtƈ�ȓ[6�a�C��/�p��)_:��݆�*i"���g�#L���!'�;1�-��(�Q+�Oތ%��Ed�+�T�ȓQ��8 �z�i+Я�c*�Y�ȓeN�H�N:DRx�zC�Ȅ���G}R���%퀥G���ط6ۊ���=/��m �&Է�yr�^�� ��J  	���cT�y���/����|��IΠW�\cĉ¤=�T�F��A�!�d��ɡ���]�޵��ʔ���$�R���S����<�L�}]x����L#�L�bEHqx��BwE�3���1��SӎiPlE����TQ!��~�f�1Q�S�#����Ɇ9[�ўl�2�޸rXȴ��&N ^��P?z���[Q�T�#�!�K-nv`r@fB%v����iټXB���'h8� �^��F�? �qS��&Ͷ˥̟�x����"Ol�A/A<3�����+N���R�l#t�F�y�,I
��'��C�d�9&�V�I%E��:{��a	M�c�wΠ9�t"J�*����W�bИ8��SH<���ɲ���RF��m�&Y�� �|�'�=Y<4����~r�,�91���z�旕@^�p7��W�<)F)�=zV�Zpf_����<у�/b.��M>E�����$����ռ2�b� N
��Py�&B��:���m'|�FAm�d��*�J���,�����vک8Q)K=#n�� ZZ�����J�*ɑB���c���ȓ�ztI�t{��1!);8���'p��a��d�S�O(
`z�DM-�^����̇ct���'���8{=
��N�5��D�O<1VKݧRn\a���=:v#[i�TtRa
6��TG�X�mo�ɖ'��@�Am"�9�D:t�j�͖����Љ�s<�0)G��HW���3�I��_}�9��0n�<�TɃ!Dk0�	0�vڒIi����Q\�P���3a�B䉋?�J�#H0�j���o>����i�zY�f�10����� Q�)�)Xin���O�=���7D#���4��Mbe8��'Fi�VH	= ���@�`�	g[� �e��g* �A�ȉ%B�x���UP�(֢R^���+A��%���B0o�\�*��#�Q��8`ڀZ+$���E�c�6�au��58\b�եY �����6q��e&�l���ɚ����'�S4z2��L����u��6�����aߑeְ�q�d̋^�z�3��)�^��m�g�*)�La���'(�!�����)Z� %"C�R%V�����i�TE�\R�"5�8u"Ř?��RD��Gh0�?fX�"$.L�r��dF�'$�x)���P��ac�U�x�<�����j�ƇDNx��'�By����`kyBD��'�\ѐ�\"l DU�&��&Zd=R��d��'R8xbHڊT^�m��I×[�-X��r�&QD�������7m�4)�'y��R�g^�k?x�A@K���i��%zv��>���Ti�e|��2'_�h;|�>)i�&��.�
Pir�Z�9ޝ*1�@j�<�q��]�\!y���N@��Rh�~P�5�TPu��P`dU�/�|��OIX�Q��Q�	�v��� ��F�J<�Ѫ�$�v���$�x�:'�2r�v�б`�p� RB���@[����8�##�.-(	�c'z�'%�*QV �ǟ1��4G{¬�F�aQp*�Rك�ǌ76����a�O��$a#VY6z�b�3я� ����ē�:�2D�f+�M���c�2��	�RD��+&�6!�=h�.�+}�*�b�D��d)q�r�3�U� ZR1C(�	|<�	P�3D�4a)��6�\\��ƁE�H�v�!��MB3	��[mnt�An||˧U`��`0��*8Z��ċ�,�\�O_	�a~�ψTR�p�B��Pf( ����x����q*�A�f�����P(׊/�y�Y&}��#���[KbY)�߬�O�)��OלPj��2��ɭ)����u��M���5"X�|b��sM�#Q��BU"O,�:�ҥ7���碅'�pe[�O,�Y'��>*�$��*�N#"�P� ��q��6U��S�(�R�<��hő~��"�M�4@�sSBA
H�P���'�QC���5 ����On���3%ʵ�d��;�����'�0��N� )�X��A��|�=�p횱8�4�*�"H)v���	5E��2�4"�t�K�E��-���D��1���"��I/��p�OI<v�zHc���6ZF�C��%S
�I��Qv2���C�<V�DOf83էN�����OV`�8��[�����Y8s݀���'� PQ���;:�\E{W���c�,���'��� %��K���P��!�i
�'!|�A���õl�!v�d�
�'�
5.�V�D����s�`P��G�L@)JA���;s��0���l=�2fnR�5�F<���oG��ȓZv.Q�h
B�,=���V� �ތ�ȓ@J��̛a��q�'�F�S|t��"����gD�Jz���U�RU��ȅȓR�]81+��C(��e�r�݅ȓ.�X�#���e��B�c^�A��S�? "�&ζH��42�*ٽs�`�S"O^�K�ꖋ@ծ@׈	'���Z�"O�����(e��1C&���Je���"Oʼ9��7B|.2g�C�k��)V"O�����8Ya:��KB�+�Ju"O$�Z���3�R,��Q7�n��`"O�2Ɯ�,;P)��?n����"O��8I<?n�DC��@(N:r]*�"O`�b��<�}֊@`�B"O\��B��$�0[�wz2}�%"O^�ae /�R��2g�7We�	�"O~���/Z z~0�f���� �"O�̳Bٜ|ْ02$�2]�F��"O��Y���c��9��AY�U��H�R"Oa:c̀=�����VP�.ě�"O�cC��n\�� ����d"Oީ(�.N�*�8�EI1�;�"O��"p�־Uru*�M	!�T �w"Or`p�K��S�r�����,��0"O�yJ����1E�E��&�u�T��"OU�1�H!~`�M�n��\�A�"OJܚ��
|������7��2'"O��Hah�0j�n˽s���R�"O� 1R"���m���"O��G�:�D�AՎ�:��`Sq"Ol԰-1�^�!��Sac<��"O^���L��l! b�G��0�"O� *��ؤ��^�N��-�p"OF�	۬bZ����3�L�i"O(�r��9s��)%*���a�"O֭rY?\�(��1�l���"O���
��  �'u(��r6"OL� S �0%��0.r��'�  C�1/�I�`r�p�T �:t�R��
V�q�C�0Q�Ц���j:��B�)[�O�|haH�)Q�����*B&@Q�F�*]-�X!���nW!�DY��ȉ �M=6`0��iG,\�9���Hy�쟦�Vl�}&��"��̝����F�,��0T,-��k��GѮ���l�~e5i��ɒY�)��[�+��)��ɚ<"%v�OY����ڀUI�����<|�$�ʊiR�J%<m��Z�8ZM�G�2sG��ȓ#Fܸ�`�̴a� u$E,��<�O6,��j��^=xAA"�(�'a���!�&:^�)ڗ�~<V��P���/G�u�$hۡ��y�v�bu
_�m��		q�i����|���=;�����͗�`�6m��`��PxBg�4���
�+��X��.�7_T�	S�
�;ʼ���'�
 F����|�D�)=�����kl(3�Aד
�����O,L{���3V�D����"(R�0�"O�HƎ�Gx6@j�➡t���xżA&(���GW�OI��bPc�d��)�p�\�,hԅ��'�  k���yn,-[�U"_T�!pH�0��"]P�1��L����K�M<je����g��5�@5D����+')~���`A�{�e)��)D�����S%6��ȱjC+x,��"� &D����߄q���cd�@�T��Q�2D�\�A.� T�po_��=��A.D���� ��q�l��u��	�ѩ/D������-��$��!��-�q/ D�x�h� v?��$��0��S�!D��(�,��N�&�q��4X�I{q<D�t�� �!Dx�ڷ(^)I�f����.D��yV�
)Ł��|.��`)-D��a���)3�L�jE�П7�8��(D���FhS���X�5�+ٴ����&D�� �T�Q�ĝbǄ���'E>K[�U�"OⰘ ��-w(@`:C �h��kb"O敹�ŏ�
��Y��7�zIQ"O.�����'�8����83��8P�"O2�ɐ��f_i�bغ{�@��q"OtIk�͜9�.5Zs�߄��yI#"OF�Ҳ�ǙhI�Q� ��0JтY�"O�@)�D���YX��U }�5SR"O���E����^�Ha�y"OX؁� �Z�IP�j�>]F����"O�pv�H������g[Y�l�"Or�h��'ZD)�a�Q*�	 q"O��Q�W�,b06,H�g��;"O�Qi5+�l�Y��Ał[���j$"Oj��D�
n$.L�1ƒr:�kQ"Ob<�tΜ%��U�҃ rcFh�"O��q��PE" �8,ϳJd
p�7"O!h��]�-pHi�e,E��^���"O<P�B�]�d&L@��Q�c8.<`�"O�P$.��[�LH����o6X����'���F�M}���5^�b�'��Ea�<�y���N~��zRAB��-y�.��'JZ�i�k
NQ?�W�L�� ���Q�-KP��!�He8 2Ԥ_|ڹ�GnX�W��d�$FC#BL�����۟�j��<y�,687�H��.�W�tp���o�<�B��f9��C �SO�QI�m ),Fb� 6c�>@Ȉ��\�v���D�M�~�@��:����=8��z"cC�`r�3��'B89��_3;ת���)|3�� �C]�?�1��g�D������/7�]�G�?̪4�=1i`Z�+u�<9Ϡ\�q�2�Ӯd�>P�g�G�/�䐠P�A�s��B�I�q%������9n�P�W�\,2�mx��j�T�s!F��~���2q�:�gyeN#T����f��;6��
�y��F��A"�kȹO_6���	�U!lQd
�&7����T��V6��J���a��#Y�\&&Ź�n��,uj؅�ɉHt"���q|�[F%Ҿ�zX��B�RB�i�ΟR�6��0O��J3��m�H1c3&��mc����>x�mb�Md���EL�'U���Kr%٠!i�5* 2V��ȓAG�{�F\����s�Ѭy8.�	T��Vj���聙?R��	Z��~r�Y��ic�5f�y���:�y��I�X�,��A�)��ڃ-�8�ē2Q����$�p<)a(R<�R�t�ԕw�胦'R��$9Ah�Qx��ɡ+��Q�&�%/U;�4�O��D�O!"�t5r �&\��0��"O`� ��] ~�`��t�t��"OT� �1c ����̡�"O�,Q��B�n��7�WZ�(d��"OBX�R,T� P�	�b!
��� �"O��2bb�/)H�c�]:�4� "O���@!J� ���:h��!��"O�H%B��j�D8�DBÂya�1%"O:Qs��:7օZBh]*HVvUr"Ob�r��@�PyقJ� Li�@"O^�֫�0���J�B�ձF"O��2�$��I��)BC:���a"OPH�I�*q���υ��5��"O>]r�_�e�t Ë9���if"O���i6FZ$��OL?��X�"O�Th@��l� e�VΖ)\��"O�HYDi��Hx��J(p� t�ɔD�r�P��$}d���� �b��􆕅oZ�B�I"P
-'��0�����ҸRqP�2pv`d!s�a�)�s_�-x��ڑp1��
�`5Jq�ȓR���j�ϔ�7�S���ɗ'Mr(c��L�2���	�?^l��K;�� �f'�v0��d�u8٪w#%� ���f*�4K�M���E+C
�!@YZH<1�e8�DhÏY�ΦQ�JG|�'�Fx��O"����~�t�V!Ӭ��_=�((R�<yѣG9�h ���P�Jކ	؀&����+���I���ĝ>E�Tn@�n�űb��i;�U��FY�G!�ވ��E�C��8;��]��I�_#�2"�I�uWay�J�0a�ZX`�A^*<�lY�ϱ��>IRFϳ}��(#֬ũ6�xt��h�bOҗ*�^B�ɧV-Z�K1��
<���$�Ң=A�	�
�\Tۗ"/�ӳ1~� ��' �c��!�% �N��B��a�\�(���g��- �6 '�扈)jLSJ�b�)�u���d��@-��K�<i9R���GoB-�f��S�܂�%�<~80�O<�%�ˢ�0=	Q�ڄG����?>�k���a�<��mN�{����Z� jR��N�X�<)P�̣$(�Mq*O�B+��r�h�By"���=���=E����4��mҐ�O:Y���	5mM��y�G�xf��c�B�T�J�+T�����4����(��p<��!X�e�3���5:ޱ�r��|�'�y3P�fyb��=�I�g4}�ЁJ6o�$JQ�@a�1BzRE��W�Й�dG	<��2Ӡ�7a�*��'9N���f��L��'v *��N&6�1����(A�m�YaGW �P�"O�C�$7\Zr eL*�j1��O���2㑃,o�X�4+Q��� U�x���� r���2r��PbJJZ�8�P�K/�O��⃈ı6� ���)�,{.�H��Os֥8����~��Җ{.f����EA�$�"E[|� �Kd��9`�����?�,W�}�7�?G�N�IV�X�b-�zČ����1=���e �*4�݀gO���p.�l�Q�aY@"S�Ot�KA�B�a�T��'~���'C	+L4�|�U��s� -�D�֑.����r�~�<��6tȸ�"%��7y��H u�~?I�E�����+V�+P���Oba��G~BH�9J�!���m�21�`�p?�G#p�<e;�O�"���Ȁ�'k��5)fX� ���	���e��I]�c7�x�C�;:�<��B
�R�(�GJ�٨O���((���R~������8z^�1�`�$hb0� �֚T��aÅ�%$��K�jQ���ѯ]�I.���3�>d/�	|��Ez�'zƽhڊE�B��~�h�,� )�u�FN-E�^�<�0�޴A��)�Gf�&\äx���۟D34L�1hbq�5
'@Y��?m��xrdC`�>LR#ǀ�7Ӡ8��g���y�@ϋ`h!�A \%Y�3@2���F�j� ĥ���<�!�]�s�!�c�-�ш¯�}x�ؠ��>n���`�D>N�㥋�BX�@A�G�	�!�&�������;�M2��
6�ў��扆�=�v�HE��ү,���q҂��U�ID�.J�ȓ��)&aǨE�(pOޥ_ ���ɲ`z�b!d����S�O�d* �K75ι�3B��(��l�@"O�IC�"	5>��If��<vR�ݓe��8�l�{�l��	=E�l�K�j��G ����˥
x��������e�,?$�,c��ʑsޮ�S%����y�lG�|���+7�k�y�P��y��e�B�L�l}�3��PyR��R�
��؛k��E����D�<�� պ`EP`�MH{�����DD�<�A��0@X��{�I�b=.�rx�<Q$���1�ؙ*q�҈tMDh���\�<1s)��3f�J�2jP٣�Z�<��AO�x�-A���6�#� �]�<�&�+H�"I�sJTz]4r��LY�<�A�ѱ{`� q�юK-��a���P�<A �ԲR��Ua�ۃ�h�E�Q�<)�OI�?|4����̼\W���@$NS�<ᔣ��Là�;�c�`�@� 1C�N�<�p��{󖉙O�z4
ui�D�<�f��cc���3eC��t�7�I@�<A��1��ƃU�>�~�B���Y�<� �AQ'+�L���k[��T3�"O�c#-��Y��"Ej2X�'"O�"�	�4-U�,�'i�'�ݣ�"O>+�n��+�A��O� ���"O�� �dD6��I�ë�	r�D�)�"O��BK#�9	��5�H��"O�q��'��r�Œ'�$w�J��5"O���qkx�d��T�H!U���!�"O�(cRF�rޢ�ڷC�%%0u"O|Q������\1A#?<,�"O�l6�]�ui�C>#��A"O��1���k������դ]�"0���'���* ��tu�f-O�3�����'Q�
����>J��2�'��J��X�6�N(6`ٝª=�'�h���q-x$"d���"ș�'���Mǟw.*`���>��'9B�- D $k����(��'J�@*Ԍ�������kت��'3z��B��򪃫pH�]a�'���8���>��=�a�Pf���
�'�d��F(z���U.�K#���
�'�4,�����gz��T&� 9�����'T$�ۂ+�!�h܁�FR<
��O:հk�$����)ςq8�$��N2`�dʃ:�K�/N�?.�D@�%RБ� ~p�)�'4
؈s�Ԕsҕ,�>*6:A@���1�LI1�������i8#�uN����$ t��30�5�'ID��ӥ7�ԣcǤ.c�%���Z�es�Yr#!}~EI5r��ć��%�����*GŔ8���5j��'?�-`jk�,�'D�O�� �\<$y{
K1g��Hb�I������ ��سDE	��H�� ��\��x�r�P����)v�ʤWOH���Oͧ)A�0L�bF�Hr�ԋ��OF�ONB�KS��{�� S�_�`�	���84tI���M�U_�a�Nа��i*ʧ)��tO�3���� m�:_:a�B�A�A�&<k�ɏ)�d���S�)��>�x���[1y��$�uUh獓X��k�g�K�<�X��v�:��I_�x�e�4=�T�f�(~�F�����PW.D��h�`Ԍ��O��X��i�}�"��pO�0Xt�̅(�E�G���v�����0|6�f��!Ipbr�Ƙ��C�u?��-	"�K%�����S�}1�d��%ˢ5h ���ٝq�v�#6_�(R��@�����O⡱ �"~,R�A���#T���"OD���! �G�`t�R�F���k�"O�E) JX�_Ye���U7�0A"Oz&фL�UY�H�P	*��W"O^|r�샃-�E��g�b���d"O�� k�%u�^e�c��	�B�S�"O��ʲn�&JL�7�F�FT�"O��k%%�>d������r��X
Q"O��@�8��U���#	w�%��"Ob�8#$1p6��� ��#v8�� "OdA���S�KfTp����:�h"Od=Y�G���:f��|���"�"O��s���T֠�fnE�@`,؃"OX�,�
,����-E��"�"O�kA��j�(3C��9k���
�"O(������tq5��.R���"O �����R�Jyc&g�=�$�s�"O�\Ჩ(_]Jh1aE���P0"O�ѫPcY�]2*y���U�B<�q"O��	���N�:�0cb�\��]C�"O�����zҘ�UÐ'n���d"O�	�	�2j/�(P@c�-���*"OMʒ�8[`�*Qc�Ms�QT"O� @���e�H�0�`�v�T�"O�Hې��8�rT�c���\q��:�"O�Pc�V�C�|���å]��"�"O*�B��*N����=MK��R"O� ԩHG�����	P��l���"O`4��G�>IL�) .C
��g"O�8���UQ&��#	X�8���;�"O�,#�GS1N�9	CG�o~Ԍ��"O�<x#�C�}����%�(s�޼ۄ"Ol�aH]�Ex�5)x>5{�"O���G������CS�~��A�"O4�A7�ř-U��Y���I���a"Od�`�f%K�ĩ�l�K�Z�r�"O$��@ĝl�����)��Ĺ�"O L����nX$�FŔ5H����G"O�L���|��<~�UX�aO�8��[}��*��^�<��r��W����|�����.=������ �s�>����B��U.F>�Ԓ��["�*�ȓ������.��@�h�A.�ȓ� ���g�e!��+�vj���Z�*�j�,L'!b	0��I�Z�@�ȓ��%	k��f��K7훻@�A��R$��p�#'��{���W���5�l����ƒ,��K�]�9S���ȓ`hJ� �+&�p`suR�[
����~k`��E�V���	�CǶa*�ȓC 0JB!_������Z�I¶|�ȓx;�<�3h�  Y	vD7G3���u�|D��F\��z���6^F��ȓ$@��;'N�R�\)q��4e����j�+��-/��9�Ð�v&P݄�n��T�QL�	���ĭ�:4pp�ȓ\�%�p�S&�@�:��TVMFنȓ7E��z7�qF�������A 
�+�����ME�K�^���1ƙ�c	T�T�0�EE�$Jp������0
+1�`����'h��D� �[dhJ�Ff�q�'	�;>�0��{Fh��,T�a'�# [�c�$��7S��ö�O�.�l �� 5g"Q��*SP[�&x괌��Fu� ��m���cHQ5<�^i�D"�y���ȓU�0��Ji�ęP��'��D�ȓ~�W�I�s/PD��L]�\ņȓkQZl#��V2}��4±I߇cu�	�ȓ�Hȁ��9��L�W )U#|�ȓ#)\�K@ܷ:�z,�"���#p|���J��
��2o��	��.b.H4�ȓW��Q�&�F0D�x� �+Pm�1���FѫO��P1��<;�D��W|��h)��P��i�B� �ȓ)�����Gc��u Ȱ�J�ȓ[�F�I2��@	�*v���ȓY&,��޷�
m����${SM�ȓ_E0�H�@��]�����ɦW��p��K��4R��S�P�Z�k�"J�t�ȓ*�2,X��(d��3Co��*C�-I�l��ÆM۬�)�hN+��B�	�_�H-�qiL�l6��!��N�=�B�03���!/R�a�f��`��.bC�I �l��F=/ij�$C]|�>C�	�M�x�g@F�LC�_2��C䉦��kf�M �:��d&I�C�C��$}�,�YVj�Xx�ք5}�C�I�����0�� ^�څ��惦
ȈC䉷+�ڍ��d�V_�堶'T	SZC�ɳW��M珕�sc�����Q�^�.C�)� �`��F�O8�y�vKB;W�^ (2"O�ِ%�O�%�r�ꊬ@⼹��"O&�CB�$`z�"����ji�"O���rL��,���y��D��͋�"O���1��imڧ��%�HI�f"O�Ȋ� R?xBnT(pb����z�"O���9<B0��JF#b��!0"O"���#��0� ��C�<\��*�"OxL�4L��]�LE#���4+E`Q�"Ov���ҷ	���I;"C�R�"O��c��T�Vq�ƧLH���2"O<�v�	�����2k�$;P"O॒��1l�$�)A�<���"O�(��E�	w­;"bés�"O��B �I@�`���٘��"O*��f�)���DNJʀ`��"O���DV?�@��ѭA��c2"O,�k��7~0:���	i���Z�"Ox b��H�yp�x��� 5�fl�C"O�`#�
-rxq��d׌�"O��vS�y �����O�HHV"O~�{$D�h��A�C���"$1s"O�Yh����ap�B+{��t8�"O�}��+�J��ē�;W���"Oy�#ы��l���%E ��R"OQF��Y���-Q�!�U�S"O6��5ۏD��lx��2�0��"O����A�XL��!ơǨ[�0=�U"O�ɐ���0���9��K�Z�bC"O�ղ��T�a|,��!E��<0"O֕1� 1sO�h!�`]�i����"O>-����m��Cp��,��ب�"O:ʥ�F�k��Dk��%n�~���"O|ٲ�A�9:7���%�]�"OV�2g�L:U�&���M�5�Z|
"O>�0����8�Tă�ֈM�����"OĈ1!�/�:1����S���9�"O:]8����J���h�	�";��( P"O��:B�Հf���6�_�Siv`�t"O�����
)2:���E�1pd4E�"O(�#@�F!aC|�QQe5oa�yjB"O6�A��ܪy�~��dCJ�t]�y��"O��K�q
��.=I�*V"O���lDL�t��W��VG���g"O6	�`!�u�.��7φ{%�P�#"O�!1�+W#]�N�$ϐy�,�C"O\���+���8��H�F~�)�w"O�p�v��i��LRb�̖Au��"a"O���H�b�d�!�4ia Ȓ�"OجڠIC�^lv� �9�f��@�!��%�����C�yH�B�E�:�!��G	`�N�h�I]*3�x8E�[!�D�8fȺ�ѧD�>�����n!�Ě	c^j-��'K)v�&����]�oB!�d���}�7��E��a�!�-f)!��ǜ�����aǾz!p�BȀR!��
�w�����������xE�?e�!��-~��bE�֬&�VTY�W�&�!�({\Y���E��	�fD�	J!�ͩPW6y��-�<h!�dB�ě1"!�d�o�d	� �<>Z��tN�!��!m*��b�_�tF�2!��$'�N19���2���Q�E!��U�N�!�g��bݚ�itL���!�� �\��EG$�9�M����Mt"O�D���������.�h���"OLɚ��Z>�y �
�G�2��"O�L�#
�FO�$)�*V� P1"O 5���+m7@m�'�5e�*Y�D"O��k��"��蔌ۜZ�:� "O y�"��Y#Sm�1Iw}r����<!T�;��V(rp���ᇝ�<ޜB�I�r�jh�WɤMV�i�dAl	�B��q��Q���\�qV�����=bB��U�h�B懐�q3.����ݢ�JB�	,��Á��>�^9�7&I7� C�I ��!�[n`E �G�qS�B�$2�t��8&�6�	שƷ�B�	�v��8';B���I�`.|&nC䉾E1j�KC`�4�e�'�<�NC�ɇ_f�{o��Y��� rANC�I*z4�SE*�!:9����$U
PC�IIx���a@xq�ͫ���
&x,C�ɀ.ϖi��P�EQ$A ����(C��2g��a;�)OzZZ����V"Q)�B�	0�*p�d��m�z��h���$B�I 2Tv93�\�b^%c��R�BR$B�	�el���HZ�~���!�iM;�y�$Z1�>�NѶ4��D��y�ǟ�^��X�e�dcD��ဒ�y��پ������4���8�
P�yr� �L�j��p+V*bf�!t�Ȏ�yҌ�}I�`ʜ/��Q�Td���y��Ѽ`l�!��O����#���y)Y�U՞���"MB�lIT�Q��yri?C�*��']-E��:���.�yR@�gDM �G� Tf�p��߫�yr��,�����C�����yr�/�I��H�AN&�9�k��y��
DP\t��k�*O���i����yR��.GDrE�K5N�*��KY��y��G�&��\��"�F�����oF7�yDيlb�I��S5�D8�f��y2��"}r5`��n
Hv��yB�L	(��G� ך]�E�K��y�a�22 `  ��     k  �  �  n*  6  �A  !M  �X  Kd  �o  �z  ��  �  ��  �  ��  W�  ��  J�  ��  ��  2�  v�  ��  �  ��  ! � > �  r! �' . G4 ; B �H �O �Z =b 'i �q :z d� �� � ͐  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�O4����C|���D�4B�nX�lWCh<!�ER��x��ĕ20����,i�'Jayr���<�r�h�7Q�r`�rOF�yR+J?@˸�s����MQȬ���-�O�Y�㝍`x��$l��}AP�$"OPl�`h]�b�t"�!��r�!:��d�U����RA�]�>`S3��5"�B���9�O����J�0�IL�Mg��СϏ�=GxC䉵{��pP�k�2F'��i㇎A,B��ug�`��Hn!AIW�7vJ�prH3D��h��fGF�c���_Z��Z�)�>ٴ�O�>�9�H�h
��WH�Yu�q3D��QB��M�~͸n�&F��@�
#}2�i�V��� �YC nJ�l�X�|q���v"O�h��ɰ>�茹�.�^^���b"O",�P!�ys��I4��RT2ix�"O�p� ��
��eR��9-$�Q�"O� RUe�
��"��	�E8��C"O�c�O�q+���AB�.62(r�"O>���"�E.�Y�3/!(}��"OP�XѬP-"[|:�A����Sc"O:p#d@�*!V�11��r�hv"O�-����(R��6.6��rZ�Gx��S�R��B�$g����脡1�,C�	Up8���J��0��)�W²����H������ VC\ѸX���J��'����P�]�:0�A`�63�	���n��I����?�ƻD�B�8!��4v����K}X�GyB�
�Ax��S�J�mV�8�mT��yr�"i�L��b'�iq�|�Rjз�yB��""ǜ�����0J�ɲ�!�y�盫1L��!�3"� 8��Ƅ*�y�ͯGL��f'�	��-�
�	�y�*�h�H���g\�T�yQS��(�y�bkΰڥdP~�e��k�"�yR�#Nq����E��9!�Aܓ�y��
;��@�` �HtV�+���ybǘ"M��Ub&閬t�ބ�w�T �yRb��l<j\��h2W]fR��)�y�,[�k�N}`�K�G��Kl �y��W�JN����7?3�4cw���y�b�3>tX�`��09��w�Ё�y�g^-4���f-.�� ���N��yB�E&&|5C���Rd��!G@�?�y2iԙ{.NP�rGQwf�5���H��yBɀ�v60���^?!�R�A5ω�y��3}�BYِ	Ϝj���Z��y� �"@p��� M>[�`��J\��y�/ �#�\k%-IW�2���=�y�l�U�Z��ЋX�A� �2��Û�y��6$�Q��H�+ь��7�R�y�	{�\03`E�9��]�eW9�yC����R�^�-�dJ����y�g�Z;�4˧��-(��8�׊G/�y�PCE��!oé	�A��e	�y�S� $��w�C�ⵢ�Gۻ�y�(�sИ�x�T,]���W��yR)��k��3'�&u�C%LE-�y�J�"���%I�#�L�$�V��yBaT� ����N$Ԕ��Z7�y�ģ&Aj0S2i�q�������y�B�!aZ(xSB�g��e���Ӆ�y�aJp�Q;t�e.X�*k���y�n\	L3^�����W��h ���B�#O�x�)�W?l��P�J�'F�C�I�79<��X�L!�G�,ܲC��'^ކ�J"؏h�ț`� >#m�C�-h�ܬ
���-al�c���-3��B�I�v�D��C��Z14�x\�"OH$�E�ި_�ND)ҭK�u��A%"O��Z�挏[K�ȨǏ	�R�:eӔ"Op�� `��<�l��퉹~�z]1�"O�P2q�	Z�͡������"O2Xh�d $N�e�@�u�,��2"Ov)	kIw2�DP�yu"O:հ�C�[$JT2���\��9�"O|��������1NS�"�.���"O� x4i�T*E+.��p��44����@"Oq4o�)�ҥ:&L�V���2�"O���4ĀmhP��J.U�:�3"O8��͜U|$(�dʓ�@�^�q'"O��"�I;a�9��NW��V��F�'�R�'���'�b�'���'���'���%�	�:�3��EN����'E��'f��'��'���'Dr�'K2���[W��H4G�`lp{��'���'�B�'��'�R�'j2�'�P��(���&�a�G�0RR � �'��'`��'���'���'��'.�b!�<9C$�T��+l�rE�'���'��'���'�2�'f��'���e�ԣ;�Z�KF�[c�P�T�'y��'zb�'�r�'�r�'i��'wR�όYu��#d�� e�����'o��'z�'���'Cr�'o��'��ǌ�+
��:e�wK�Iu�'ar�'�'�b�'"�'�r�'�dTZ�BU�'𴹡%I��ti��S��'���'i��'Y�'B�'cB�'۾�Iˎ�y!LQ�&$�/PA�lҲ�'���'YB�'L��'7B�'K�'����  ��"F�����K�@mZ��F�'?��'���'c��'p��'g��'1hH�eE�N�A{��Cn�Ѩ4�'���'&��'���'r��'���'��=�*VQ>�1D$�2|��̡r�'qr�'|��'��'!�gӖ���O�y
g�N�DgҠ�dlC�O�@#A��gy��'��)�3?1��i7� ��]43G�P��M�,Lq.�;s�$��dƦ��?��<9��{���9�0IIB��2���3��?q�\�M��O,�ӡ��N?�p��˙*`�WG�w|��0�>�	ğ�'f�>�KD�7.�>�Y j��Ш��ݶ�McA�G���O��7=��9CEW�	�b�!��K/hO������O���t��֧�O�<0ᒶi󤁾9�t�a"���\xC$�6���v�l��7Dp�=�'�?هm�%bB�$c�m��M2����<).O4�O��m�KP�c�HQ�5-v4�m�'1��p;Df�T��8��	�4���<��OV}۵�Si�>�C��O撈*���L���aF�E�+�aGR��꟠�u�Ɯ5�J ��H�i����aFzy�\���)��<�s�W�A��e�E�S8����#��<ѥ�i��O�Un�n��|����&�,y�׉�o^���
��<1���?��Yh�8�ش���f>����z�0��q捽x*&I+�H�x��� 3��|r+OF��d��'L/�$Us�퀠9CH���1Od��
�H �8C!��ʦc>%���*�C��׊�Bh+�O9��d�O���y��'>i�	���s&���r
LK����Lu2��5#�X�*�@�>�@(��ae���Ҍӧ�'�1��J����fz꽢W	�4	2T��'�'C�7��D%���>{��m���\�݈U�7"[$�$I⦝�?��<!��?�4e
�#�S	O���ZQM)7���G�\7�M��O����ʌ���l��{�J��L��D�$�J"QnV�Z҂c��	DyB[�"~R��q'��a6]�+�Xp��UL�7)��T=��$LȦ�%�X:Gۤ_=!+rB�#���2Q���<�O��d�O�)O'o��7�6?�����@"#���U>����ù��$K ��O�P��4�.��?���,:��*.̋p��)[D��<�K>���iC�y�X>�Y���;�بiKE	y���t�1?9�Q���Iʟ�ϓ��O��E�h�%�(I硔��nEb��'fV�qÏ҄��4�¨��	>�O���mL$V_jĢ��.a3Ԁ#�O���O�d�O1�|˓vB��
@�
����$���Dt��D�5o�a�0�'1uӎ�0ѭO)o�<Xѓ��۵n�l,�`�H�I�MXش�?s���M��O�I�pۘ�).�Dk�6Z�Rq�
�4;��y"Z���I˟���0�I�� �O�XA �GPܼ�"��,BglucfIb�2-����O����OL����D��#4�"�ЁgJ�*�έ01�N:s}@��4k2���|��$�śF=O(�`v��@�M����Oj��3O쭙"^��?I��!��<ͧ�?��b7k��b���,������?	��?q���$�㦹�Qi�ҟ,�	��p��X"%[�Y��d����v�eL�	om�	�k�>�{�Խv(�l[��Q�#�L�~�T��>\G�I�|jbM�O�I���6��[K~�m����,����bK�Oo��?���?���	�O��u-�o��H��K�|<��fc�O�)m�&uD�i�	矘�ߴ���y�FK�%k�MJ�)Q�r^|����ç�y��y�vn�ן�B�o�Ц��'U|M����?�YÇJ!L\�uƉ5�p�u���Z0�'��i>���ԟ���̟��I?bA`<�a&6q˴  ���k3Z)�'�7����O��;�)�O�u�r��9Pr��a��կv��j���C}B�mӚ�n�v�)��#��|��O�������x-�!<1Z����U.�O�(�K>�-OP[��R.`�@��E�J!ڲ-�O����O��D�O�<qV��e����?�sFBX$qj��6����)�<)��i��Oa�'�"7m���޴`2�	'�uli�����:4��d��M۟'�RD� _�T�����?%�=� ft�g��
���eۀB�r}sC;O��$�O����O�$�O��?%�����5h^S.��Ɩ�h���$�ܴ���J.O�nZQ�	5,���CVH�xf�Z&��
6Rbq�J<!��i�6��4��Q)���ҟLÂ)�'u5��0�-�'��Q��w�2!r��'�\$� �'��'k��'c�4 @�_
�Q�B�6fo�aD�'�S�\q�4"@�(OL��쟪�)A�D���*C��vh��D�It�	�����Ob6m�q�韈��6:0��݆8����E#��%��aӱ�W+(��m@S��<A��U���$N���qm�	h��Z21ɞ����Y'����?����?)�S�'��d�Ԧ}��$M6g�-(b�����a[��۔ch��C ���d�D}�j�~�fa�Ξ8  cN!_3бC�KΦ�K�4uJ`� ڴ���\Ϣ(`��S3P˓L�����	S:|u�1�B z���͓���O����OD���O��d�|�#G�k�$$�S-�1�X����*$L�椗'$w��'�����'�7=����X��*�J�	�H���^ȦiشA����O����i���P9#D��B2n��xR�ެ]l�@�{4���-�l�Oʓ�?9��'�S;�X�#�j�����ϟ���Ɵ��	Syi�����O��D�O6��*��<0g^De��@s.�O0�O���'8�6͇Ѧ�3K<ѥΞ@��&KQ�H
@x���<y�K�$q����m�(�/O"��܆�?A�l�O��� �Z��i�P"^}Xj!��O���O���O�}B�'��p��ϛ|'8��T���[�d���� ?��	�����I�MK��wϺXr�E=1��0��ЫJ� Q��'�"7�O٦�ܴ'*�X��4��֠[�p���G�d]�֢MYrZ=�a
%v�N�C�c>��<���?����?����?i���W�p����˾r�D��G� �����Ѧ�;�JDy2�'�>��'�7B*03��5m�"A@u}�OxӺLo�#��Ş��}P0o0]���с�B0-���� B���C�򤋿t�����14v�O�M��l1��-�ѡU"`���2��?9��?���|�.O$�l4q�\e�ɟ�`�" %��b"�Q����~��	�M�ҋ�>� �it6��Φ%���I4E�6����n�E���)�*�o�[~bm� fW8���M<�OA��[<O~��i o�:Lq^���n���y��'���'��'b��i�N�T������&�t���݈i����O�$�ئ�)�%�ry�`Ӏ�Of��^u�d��1@�W膁7,��+�'��7m�����ld~BE3+:R �]�x�mSk�L(ƢL� ���|BR����Ꟁ��Ο�ir��������
3.DHc�֟T�	fy��jӄ)�q��O:��O.�'dLi��)7��rg��)�x��'�J����l�
�&��'@���5�[	NȄDi�H���I$�<JNH�1�lK���4�)A�!���O4l@F� 3�`��N�~;��E��O|���O��d�O1���%����8� �$5F7&��B�թV�m��'Lb)p��올O,�oZ�U��yC��#d�L��>:�dA�4k˛�A\&�F��D[��V$f� �nyb�CKu`H	��(H��ʄF�5�y�W�$�	ҟ��Iן\�Iڟ@�O��txr��:��u��!FA�ư�'�h�N�T��O6�D�Of���dAܦ�ݍ�p�-EN�b���� ���H���M��|J~J�L�M�'�.�:����eK��-v꜓�'�H�q,^��<�r�|�\�����d!RO�yVz�Җ�U�Y��<*lQ؟T���0�IlyҢy��u+���Oj���O&�:CN�]x���h?i�t{�"�I����ަU0ش�'{��H�G)F6��jV�͇c����Ob�	�L�,7�N�)�f'���-�?��F�ON\�B(gFDeٷi�$.�yw��O��$�O��d�O<�}�;w ��P�N�e����DȈ%m��C�뛶m2��I��M��w�҉P�JOXP^X��IH#4���'��6˦]
ڴ7��J�4��R�Ji�%������I ×�Y1j��@�� S�X�A"5���<A��?a��?���?iLܶMV��S�Z!���wb��D���	S6(���P�I͟�%?�	�4�����*�H�@䇈4��eګO�Dm��MS��x��D�űM߸���O�/v��SAB6'����&����V�8W�'#��'��'�h���� $�@ʖ B���5�'���'����dY�BܴZ�����}�*���7%�E��I��T��?�ſi��|���>�b�i��6-���!���
k�ժ��5Ua�1sHڇ,�|�l��<���f>M�����ȫ/OL�I�a���(\f8�!##ੂv;O����O@���O���O�?aJv.T�)�c�5_����$����Iߟ�ܴke�AΧ�?�v�i��'����s��KY( ��9r�5(�	.��KߦI���|f7�M��O"�y��߂z����7c��|��\����`��=��p3��O�˓�?��?����a��ʘ�9����UY6VԂ�K���?I*O(�oZ,ks���	ҟ���i��C�zà�A���l.�Öc���D�p}�i�4Dmڲ��S��LA���3��!w�����.by�����!��y� \�� �rH�`�4Y�}�3�܄F���`��kڔ(��ɟ��	ٟt�)�SVy"qz	�=�h+���(]��-q�K�<D���׫�<9��i��O�-�'��6F�+�C�j[��$ѷ��%��oڃ�M�R�E=�M{�O����X�����<� 2Y1�*(�B,���
�\�92O�ʓ�?y��?q��?�����IF �P���G�+:�x�#�d`k�l�Z7�d�Iϟ��IN�s�X�������H�L�!�2b� )Y��T���Ar�rM$�b>ef�ۦ��w��Q����%Ϩ�
�$q�r0̓+j<���O�A"M>�*OD���O$��@+I��|i�*HG�0����O����O��d�<i��i>M[��'&R�'|�3t	�TSF�*rč0=�p�����j}rabӦ�l���/�R@h�ʕ14�2,`���,͓d�D�霂HV���n�/�?ɮ�0��KOݺ���'�t�7%D�=i��T4<ƴ���'��'���'*�>u��Z$��B�T�>�h0��[�Xy�I��M�Cb�G~��tӰ��*�i�����Ź�e��>���6�M�ǲ�Ųi�B��i6�ɜ:������O?��Z&�M��a�!� %y��`�D'�I`yR�'��'��'��.��~r��S�L"6c�e����I��M� ���<����?�O~��x�̓ ^	�ŀS#�G�x�^�pj�4(1�V(�O�#}��"�+^�X��Vz����rhOw�V�H�%�7���!C0X);�Ÿ'��I�WN�#�A:Kp�]�Í��}p$��I�����P�i>=�'��6�M3t��D�5W�A�-
�Q�0@��!šd�$[Ԧi�?�3T���ܴd���n��q�"/�US��ؤVҵ�w �:U/N6<?y׮�l����������e��/�D00���M�����,�<���?����?���?Y���K�'g�u�\�_d�A�f��'U�q�����<���$����$�H�%c�����c"��M����[4����v�~��	��s;T7�)?���&1�]zCH����f�{�z # c���%��'f��'���'˰u�0��7ÈT{���n>�����'�bX�P�4Br�M����?	���Y4#��0(���
�B�K�B��ɜ���˦1����S�@�$��xs��?e��*�e��^$PIR�ʑGHZ�R��
)H�hY�ɞc��W	�$U�(يhEHQ���I�����h�)�hy2$��8Re��:P1���S&XYY2m��*9��?�e�i��O.Е'���)�>6�ƨ��� ?G4��;	״]��6��ئ�3S�����'����e� ~�.O�b5�30�
A��;���9O�˓�?���?q���?����)ܝU��A���8@z�s�B��%m�
���	�d��z����r����Uk��,zJ܊�G�h�� o^�·i�����<%?�h��	ۦ1Γ%�`dp�h� *�h�P�C4��S�� �� �O< J>�+O����O�آ4*�J7�g����B���?���?�����ę�1@��n����؟�0�*<�NybV,��Lo�y�#�x�����
�M�i6�d�>9���	,X���-�:s�L9��Um~"�)uJ�H(�!� f�O�x��k?ᓉ��6zm�#�OF���SE�?y��?����?����O�h#Da�2�ZH�A����ĩ!�O��lZok��vț6�4���C�	3��x2�jʿ9���v?O.�l�	�M�ҿi��p7�i��I�~�
5�'�OA�x"wo'K�t;t&ҝ!��hs��:�	]y��'���'A��'��Į���#��/�:���i�剢�M�I��<����?�M~�.��]Q0�טF]��3��SH���^����43ܛ�i�O�#}j��V#P�
@ܗ';x�ȗ�>{�x�7b��^�j���Ը'��E+W7
�dY�@�*a�v��d�'r��'<����TS�ܴ'�~T���i�y��չu�ltY��#D�ɒ��l�����_}�ld�����¦QCQ$�*k�vI��]:�Z�X�`T�Ed��m�S~�c��Q�Z(��]��O�� T�X(d����^nR�HvlƘ�y��'J�'��'xB��^;s�x�1��L�RKʲ!����O���N˦y�m`>9�	�M�K>A #Q�k�~�g���*PR���2�'=�7M���ά.�V7-?a #@�!x�YvC�)r�I@������G�O*�K>�*O��D�Op�D�O�-	�� �(|��0肢N�2���n�ON�$�<	�iS��[1�'���'�哉��\�q
�
����F<�Z�j�	'�M3��'4���I�;L�ahr�
@VU���;%̹�P�ܼ/k�y�o�<ͧ|����>��
Ҫ(b�����kT���Ȼ���?���?i�S�'����at���m-�x%$\(Î�ط������Iǟڴ��'*��G$�F�P�Bv��S1LYSprA��L�k�̑1�`Ӵ�9X���VF���(O:�
A ��=KpH��I?���R9O�ʓ�?���?A���?�����۝u�ԌH2��(-�02��5e��%m�2E�����Ɵ��	u�')ƛ�wҪ��-*>�cj�d��yp&�jӜ���u�)��O���n��<iv'�C�6D�U�[�/�+A��<�jRR���Dl-�OB˓�?A���*i��˛PX�4�eN�X�t����?���?!,O��nڧyޘX�I��P��(�~p��4~i�E��DV*<Fm�?!�V���4�2�x�M���5�H
`Ö�{��Y�L&~�͓�?Q4l���Xbf� ����p���_�����zNn,(�ᒴ%?��Fi����O����O��3ڧ�?�P,�??B�S�ޕvP�����S��?�i� ����'���zӌ���T�t)��$	�_5����̋�>����MC�i8�7mT�>I�6�)?�OؗPy��)�n�? ��`� 5�$���-TU�%���'��<����?���?����?�f�9��ԒŪB7h
L䠕b���D���ۡ�`��ޟ��:$a}���c�
ާ"�
���� : �	;�M+��i�VO1�����L fB�X2�*�|"�L��R�o�`6�VMy�e��@�Pm�������,����D����Y���p�<��Or���O6�4�ʓO��^T���<p�h�g�� \[s�S�Tib�k����i�O�	l�)�?y�4'��)�%�ź0��[D
�'��|R F��M��O��:�銿��.%�i�� hR��48�Vh�'�`cq37OJ���O����O6�D�O`�?�ؠԹ����P*<o����	�̟���ٟߴ\�$̧�?�i��' `�"F�а'�~Q3���f���CB6�d���y���?�U���Q�'$`� �I�!i��PX�g��-���G��k�n �Ɇ0�'��I̟l��ڟ4��3]���F�˻AU�X�c���Yv�Q��۟ԗ'7�	�����O:�d�|�C�L5=�RjJ�h��(��Jk~r@�>)��i���'�?����8�$�ipg܄<�Ta���oȚAQŉ�x.l������ܹ֟ �|BN�,l�U�ԃ�	��Ȃ0���j���'q"�'���^�p�ܴf�pQºX,�xT ]�U��ks*[�?������PA}Ҭt�.M�K�1p,�@܈ ��pv�F���l)M:��n~�"�!������I'?͠�k��]�^
�*&�� j���}y�'�b�'�b�'��Y>�i�T�8ȹ�F�G���f�[��M�bQ�?���?�K~
��jɛ�w��5Q�aD.O�r�7H�z7���������n�)����mZ�<1׬0QD��* FSM��Ы�^�<1E��-e*�D=�����OV�$�
\�&e�ԉ(;��PΖ'2Ͷ���O���O�s'�f撻{B�'W�*C��q �	x��ǢQYA�O}�'}6ML�ŻN<��G[�SE(d�i�-n���t�[~BҢvѾx�c�M��O��\��M�b�.O�ΑZŝ6g%���d��D���'B�'r����0���6Y�����۸|�z���ܟp�ڴ\.�|��?���i�O󎝺\k��Nŉ{�4����?G�����)ٴ+N��,�R�����Dq�Y�}��dkM07π1���J�x���Ŗ,ň1&���'�r�'4��'b�'<�Y�)��w_D��FŘ; �(�P����4r��4���?���䧆?	�.�w,j�RU��'>`�u�A�	?f�����M�"�i1O1�*��w�3���R7F�3F��(�<N 8+�Ġ<�G����D�������:q���tC];LZ$��2�K���O����OJ�4���Oݛ�R$%�"��M9~�Ѳ�D�s�4�b�'q��e������O�alچ�?��4/��҆�ŋ[��C�#D`h��#�8�M��O����Ȁ�
��?����,C1�ߋj9��ufI3x)"��6<O���O����OF�d�OD�?�QR���E��˒H�D���Ev���	Ɵ�yݴq��'��7m.���,D�Љp*�'U9F�����`��E쟌�''����4���|p�֜���U�Ѻd+pd[c�'pB�C�*u&<�jv�'EqOZ˓�?����?��M�i
!��/7o�Ъ 	-]|�C��?9*O\�m<c�6�Iџp��D����'n���$�0UT��Ř.��D�f}��xӺ�lZ�?ь�T��5
B��c0K^<:<ѸP͙/,ڭ�@��&��`�S��SU���ĉ�?l�YS��'vW
�;3�Q4-��D�O����O@��I�<�C�iň�T��6���� 6��ŃU扛��������?�D\��[�4@�ƔJ�� Π����2����ib&6M�*��77?Y3A\�#˸�������F����@S�y���S�Q)s��ĭ<���?���?����?-���G#��G��0��)�62�&m�Ϧ5��mt� �	䟈'?�	����w[t5��ͅ.C�|h$���ЍӴ��OT6�ӟ8���'Y���4�y�L�\���_=�)9���y� ��y*��IZ���$�OJ��Q�4�e�sa��Hb�:GD�hl��d�O^�D�O�ʓu'��iG�?!���?i�OB�*�&��&��7Lk�MK��K���'D���?�ٴMj�'O�}I�oK�k=����D>���Op4��B;J��6-�A�v����O����	�d�K� U<�uN��f���'5B�'���s�����W��HC��\�Wp�#�@�����49!�����?��i��O�n��L����g��B�����V�_��ă٦����M����M��O���7��tJL�9�JL�с�!_X�0��5U�V�O��?q��?)��?	��c�|D�� ��$c��w���.Or�nڰF ���?���h�t��Ne)`�v��!iS��ot���f���_�Oc��K�+�~�ġYr�3Z#���E�g�2�@�]��X��9���<i�h8s������b�P�&��?y��?����?�'��H���G'u��!&���2F��?�F�lv�|ٴ��'2`�?z���d�J�l�<C����7��>.x�
�I��'l�hñ������'DJRk��?Ah����p��z �S�n�L���Oٞ~��⇤g����ꟸ�I���	�����I�a�~<�VKX�TI[/��<	��?��is���O��nB�I�X��ʢ�׏z˔�C�k�T�{����!���|��j�4�M��O�5(� TAK��
.v�[u�ǥ
��P�����?��{�^�@�Iܟ�	��
�'mn��	D��h����C����YyBqӢ�Z�=O����O��'p��)x��K�+'�yJ��H�N���'�j�>�� q�H��	M��?���������1e��(`�R�HP��K$28P	�<i�����D,�ɋ0��ɘ!����TB���MmZ���ٟH������)��byr�k�6�H�l�v6����lr�*=�bW$˾��O*Xl�g�\����
�dG�N��d��JU2�Y{!���?�� `�Ul�K~R�Ӏ;�$��Ӹm��	�'���&�V^@�#+�'�2�	@y��'��'D"�'�W>�X�F¾K��s��D6��6$��M�e��!�?����?�I~���`қ�w��<0�"=L��d��"W2�HU���Of6M_^�)���W�7Mt�`�c-E>�p�2`ıM~*����l�@���,�=���<I��?iU�8F�a���T�q�\r3��?����?����D����A~y2�'�䉒f�ˋE�N c���:��M��Āuy��'$�x�鞇b6��WK	 M��
�����$�D�Aӓ�N����� U���6�D*8%��攬��s1JWwi(��Or�d�OH��)�'�?I��&/R�Sq!@�1���։X�?öi�za�q�'�Bhe�����p��C΃u9�i��*ȃ�D���Ms��'����W�X$�Ɯ�x�G"����G;S�8��BDF?s*T9%�<Ɛ&�@�'�2�'���'���'��ىufG,r��A��	���;�^�Ӧ�3W/D矠�	۟'?��	~D�J�`Ҫ��a85'�K�4r�O��l��?�L<�|ʣ��%u?��PP.�)��+7_E���+�C5��$�48,�{��*��O&�g8T͒se�\'�]�1�_�:a������?���?���|j+O(4mZ�e�r(�	�m�dI��%R��[Ct��ǟ�!ܴ��'�,�J���,�O6��&7�5�vi	6!6�����-U���g(���d�Dd"�)쟼]H~���]5	 ��Ndn4��j	1@�,�ϓ�?����?q��?Y���O����dشF��82��T�J9��'K��'2�6�
%Y��)�O4�m�M�I1�ܫUN�p��S�(�ʹiH<�"�i�6=�@$�&Im���4�y��/4Cag��(�TB�ɘ5h�t�IX�uy�'B�'�"��&B���aG0JlXS��2���?)(O��n��gO�$�	��d�	R��� �V�L ��B��;�������P}�'h�l���S�4�
?hK�0��SǣYIf�
t���Cr�lӐ����	S?aN>��CΧi@�A��K	�+Kԅ22v���O�q�����O1���f���K<rJy�ei)n.��fB��Zfڤ�c�'���p�H⟜�,O�6-fB����(@7VH�d�]]��m�?�M��j��M��O��0�7��dZ��9B�^/q�a�U'L+J�nm1^�y2T���Iş��Iß�����Ou���HOhT�h'Nܠh�t���Do�R!I�O����O�����Dʦ�]2F��y��7��Y�S��2�$s���M���|J~�`�(�Mk�'�4�:�MϰQԔ�����-Kz�Y��'��D�l	x?�I>i.Od�$�ON��$?��zeNb�,(9Am�Ov���O��<�i�V�;�'
"�'�͉��U<:v:r�T*��"���P}�u��yn�?	�O@��rჲE� L)f��i�2�㕟d����qg�pEUh�S�skB�O�I�Sg��R��,Y�� _�F܃*�O��$�O&��O��}
�^��y8�$�&
]<!k��JI�9��[v�#ڲ��$���?�;koȈ��B��8��f<�<��F�{�XLoZ'>���n�u~Rb�h��)��Y�yQ���M!*���(̍���ȍy�X�`�I������|�	ݟܣV�� ��a#��R�.43D�VzyNs�ԡ0f1O��$�O����$ͯpU���)ň]�=�c`��ш��'�@6��!���H��+�f�0,���
S9Gu��Cd�\�G�8	+`�<Y�εQ���$�	hy2JI<v����3z���2�� @�R�'��'+�O\�I��M;w�Z�<it�H�F�L�4����9�!�<�D�i��O|�'Z�7��Ʀ�ڴ@���V%;�*���]�"��8�'�5�M�O��Ӄ�!��T�.�Ip�!4j�&o��4��I%([W���y��'_"�'9B�'BB�)��[� I�ݡf/ޥ�UD�9��D�O��d���.��I��M�N>u��6(���F�I�y3 � T�"P�������S�w�l�z~���@��vN�?,p�ИQ(�ͪ�����t�=�-O��$�O��d�O�0xs�L�<��b����xDe�Op���<9��i�Jٳ�[�@��v��/W���	��mruBS����$�Xyr�'R�|*���+�gL0'*��h��]��=��"K�{0�ɓ�R����|���OZ��H>�4Jԋ>!�|"�=z{��B6cۇ�?!���?����?�|B/O@un�wɔ퉋f��kW����C,?)�i��Oе�'4�6�u�R���.��X�T�����#\�1m��Mk��Ը�M[�OV�2���������<�$��t���� %�'g�]��*��<Y/OZ�$�O���O�$�O��'Y�b��g����j9�1@]��2 Q\/᪴������m�'P���w亜{D$�
{�D�r/M��|�F&kӈ�o�4�?A�O1���Eu�@�)� �e�r�?s��pe;:r��2O"\$���?��{�Q���������&�N�)�g.�L����W����I��4��lyht��3Oh��Ol]�h�,�8�$K
"5~9@� 6������O7-�ڟt�'K�\R��A�v� �ʚ1o,Ts�O��V*J0
���2�I)��B1�?)�'����&�;4sP�B��T�%��	�T�'{��'���'��>���.�@䡷D�1!Ԅ1eMɓpw���I�M[��Z~bAaӂ��ݶ-h�ȣ��T(z`"U�f#�扑�M���i�6M�RlJ7� ?�d�O��^�i�<s������Y�"���'^|�.��<�)O��D�O^�D�O���O���`hĨ������#2��dk�<�7�i<���'���'��O�BmPf]̹�D��d.�| �V>y"�j���hm����	d�Oe���d%ԛE��SI\�*�0��A��R���<��i�/���������Ĺ�&Iq@��3uE���tS|v���O���O�4��0˛�@K' bb�$�����!Y,%xc�9
%""b��<�OrIn��M;�i�j�q�P�uH�9��£��x2�,Z9-g������#�\���tgA��>�5�&G��uC��Bv�%� ��0�y��':��'.��'�����u*���Γ��h�W-��As����O&�$��gNn>=���MKJ>�wi� H�L�᫛��6M��C�z��T�$�	����j��n�y~���9�2�p�J��1MJx �@�'M��`0��̟d�|"_��Iş������H��~R��I�b�1]�"q���ɟ�	_yBFe��(I��O��D�O��'f0�҅ν��l#ր,H� ��'�
�8��Ƃf�p-�	a����&�%8�؅0�#Z�c0�@
�,Nqp���O^5��4�lѱ�vՎ�Oz���hA�K3��@"!̌���#�O$�D�O���O1�4��ܴ<�N0iH'��$�C-�y��NH��?a�� �v��L}�}�V����!R�ƅ�w�9�2�9�aUϦ�#ܴX�ܴ���!|Ԗ���'���	�t���&,���7�V�A���	fy��'f�'���'��R>c��Q�`=�	LI�D��
[?�M#��K��?Q���?qN~J��
I��w�-�u(x�1C�	ރL�t�;��O���1����F��m'�63O�)`dmYH��2���o���0O�u����9�?�&H(�$�<���?Y��.#qhuD�-q֠<�W��;�?���?a���DIǦ����������@�1L4C�b�1�LT	[8\�rď�t�
��I,�M�@�i'jO$@0�L
JD��	sI�@�R-av�����R$��=Y2l�W�S,��l�ğD�l̢ 4q�������{6��'��'�r��ğ QA��'r;�5#��3Cjy�e�Zҟ��޴O��'�p6�4�iީSG�T��@]j�bO�b�vm狺��I¦�8�4���s�4���Ǳ��������hk���#! ^dY��T>0�
���<i���?����?���?�3l��N�0�d��	%h ��׾����ܦ�r&(?�����O�� �f���ܑ/
!ؤ
���>�0�iQd7M�۟E��IU�U��e�Q�L���V=~�:&��#��I�Z���e�'yqO���Q���S�i����	��R��?���?Y��|2*O$�m�{�|����:��Js�G[���`�u\f��ɇ�M�"+�>�1�i�7�ݦ��3:��?�8��!R�
�M��O|����!�b��7�I����B�q�4Y��/�:oVLc�H��<���?a���?!���?	���@B6m��ypɀ)�z .f��i���?���E��@_�����':(6m0���4\� =Z���t����ž��@��c}R�`Ӛ�oz>	��L�妁�'��k����c�)��LQ��F����'T"�&�ܕ'���'�R�'�&�q@�5D �d���@���r��'U�S���ݴ|@Ո��?9���)�(L�d<h'Ǆ/%�"�_6D��"��d�OJ7ß��~�F�Ld�����;�p�{v�Jodv<�D�^Z��)O��]�?��.�$B�mT�xC��5휑0`Mԛ
!����O����O ��i�<I�i�v���,$ob`J�� \���q��Q�
]��'�n7�3�I����q�ıB��}J̽@��N�2���B�릵��4���ߴ��dUyK�������j~r��#	Z@��Q�F�N%����d�O����OR�$�Op���|�2+@���j�	֗F�V����7��VmR��y��'����'v>7=�`���ݷ7�.@"�FݼR;��b���֦9��4�"_�b>Ic�AҦ�ΓL��LI�I�Q�H��U��a� HjQ1���O㞔�'	��' �iy�hJ�K�Ny3�\����"�'���'BX��k�4L+��?��Z9�iӑ���kw��`�N�7N�
d����>ѧ�i�6�D����'�&Ap3�МA�`��!X�Y"�� �Of(��V�^�^!�@e;�i^��?��'�tY5�Z�Jt���@\%P�\�t�'Ar�'���'&�>]�ɨA���j��]�O���X7aP- ��	��M�5!�~� r�&��)�|���1j�$u�O;$��ɯ�M3�i�F7�%O�T6m7?Y6J�UM,�	ړ��@Z��
.i�=�Ƭ֘N�"p�<�.O�$�O���O^��OQ#�č=L�� �ď{Z(yC�B�<���i�܍ښ'�r�'���y�J�;]i�@�eM��~] �E����o��jwӦ`�I~�O3|0�� ��6��!|<���A�'o�������|��˓�F R�o�O�㞤�'d�q�ŏ*,�Pd�cE�>*ʉ���';r�'����P��`޴$i��ϓQ��!���&SA|92��/{���ϓK*�&�DN}b�w�l�n��MF���l9��Ä���Z���1C]�9ݴ��D��H���>[��� ��y��X*�-�/`����T(T8�����?���?i���?����O3��2����yʶM����2$�z���'*b�'4�7�ڂ6�	�O�$o�L�	.r���F�Q�mlv��!?pD�B�y�	��M������U������"Wm� ��F�H�N���$
(kvP�6�'`��$��'6��'���'�f�8�N^Lj	@Q��#���"��'�U�0c�47@���?q���iX�P��m:�B̼k&���b#̈́M�ɳ��$QĦ������S�d�οa�¤0�$u�H�zA�=y�����&`�q�p_���&h`2Ƀo�xƠ���ퟪD��1Kr�Ϟwb��	��	쟸�)��yyb�yӎ�Ѳ�F�mzx�R�N	y�j1����I��M��§�>�u�i����Q��q/�|B�k .������Ul60��lmj~r�Bqi�L��.�I� ���bo9{d�����J�9����my2�'�"�'�2�'h�Z>�#���_zȡ�*
W�@Y1��2�M�@a\9�?����?�O~���}��w�F���ѹB��BB럜����t��0���)�S�5���lZ�<�6O��T�E;Ӯ�8[�X��஄�<�G%L�>��d�9����d�O�����~Ea���p�ы��F�CG����Of�D�O�ʓJo��DӒ�y�'�r(��}7p�W�V�4r(8��闔��On��'�6�P������K�ol>���/ѣ[�$�D F)E��	�GڴX�0 ��R�"t%?U���'��� �9�г��9�n����_C��$�O����On��&ڧ�?��]'']J,h��9!���Co*�?�3�iUDu)g�'j��a�����2Go<�q1�Q:j������I�X�-�MK!�'����˩]��������4K���ÒN���8�F�@|0!݃,�f	$�d�'�'���'r�'�v�;� �[�Ɣ"�� i��lP_����4g�~M#��?���'�?�'m��6�V�����
%�ebGh%+��I֟�nڻ��S�6�f1@���gB�J�$�
i=���N��-�-O\H{��ǽ�~�|�S�$E�O,��P�+�O��В�hXwy2�'c����R�l�4z f	k��Fh��@�B�+Z���(1�Bmc�&=���$�K}�Eq�D$nڣ�M��?Y�\#̗:YG01t��e��4Sٴ��d�3FAc�O*�O��
��8q$�ba�u�~p����y�'���'���'c�)擥��<��@щz<Zt��fB�C��I����I(�M�Uk��|B�E�V�|�Bռ|���ɕAC��
��'�m+VOpn���M�'K�4ܴ�������	��東!�r�{s��E��j�L� �~�|^���	�����쟄�b���R���'��r�A�N����	dy��n�@@�?O&���O��'6�.y�'j܀f�����O,R�0�'`�����n{�����y�]3��ؕ�Lqݔe���ӧ9�U�5��'����-];��4�<���'V�\#ՊU��x$��n�Hz��U�'���'�r���O�剛�M�#�'�� F��+Cc��y"A'V���Q��?�iM�O��'�t7MβB��X�r���eJ�a�t����1���VԦ��']@���?1�Q�(�SA7,�P���>��Qy�/d�d�'�b�'���'���'y��)5s�����I�|� �®@�k�|��4Sw�<����?�����'�?�S��y��1WF������6��/���S�i����?�󉘷H��7`�a�ύ#�fqH�B�8�hՉQH{�(�` v "�O�IAy��'��Q�iI V�,rmX<sU	�#jd2�'x��'����M��nE9�?����?�7��>_,�1�w�F�&)�����'���O/�ƍ�OHOۇ��5n�b��&j�7a)�����1E�,�|����R�.�Rƕ�� ����I��0)��v`{G� Ɵ���ɟ0�	⟘E��wܲ�h�R�X�˓kZ�B��4q�'�\7֩<xz���O�,mZm�Ӽ��L8%ݔ�HP(��Gǰ��#��B?����?)޴l�0� ݴ��dQ1hy���'4� S�B�	�	p2D�;js
p�N#��<����?9��?Y��?Y���T����NmK����M ��d����	w������H'?�	�M ֔���R!^kr,�_���I�ON�n��?�M<�|nV+*}�FJ8X��%�bҊ�[W�$�前/�%��'�D�&�,�'�,���".�Dadf�2����'���'/���d[�\�۴x�|���cZP�y6��RN��%i���!+��71�f�D�H}��r�F]nڱ�M#¡�t�4��O=l:�%+6�,>��6�'??i6/�,6v��J��'!k���y�d������X�[+�P��'���'�2�'��'C�&,ۢ�W�;���qmW�~�&PY@��Ov��Omoڻ27*�SPߴ���4��Ѥ�Ec���w��8��ub��x��hӴ�oz>��ʦe�'
�!���`�d����ЄWy��[V��o�~a�������Oj���O��Gq�ʍ�uf���Ve0K^~��$�Of�e�Ƃ��~�"�'�_>�s�F���#hǳzYH)`�7?�&W�(kߴWa�6�1�?� ^�ZWiL�*���K"(��h�E��F�z��f�^P�����b?�J>�b@է%B��ǂK�1�V9z"'ά�?a���?9��?�|r)O��l�&-/&�#ED4K� �A`�$o���B3AB�H�	0�M����>���i�h�b���0 �� k̺2�Y��v���nڏ~�tDlZd~�斐09������dC�q22-Bq'�<�v�#p�x2��<����?����?���?�.��M��g�"U�.��3큥*C@��O\���e��ğ �I�x'?%�I�M�;/�`i��#S��!�D�
]�����'9�FA8���D�A�(��1O��d�@��`�q��ԫ6����3O�֮�~�|�R�@��՟��M��=Bu���ԹC?l�9V�����Iݟ�ITy��h��	�PJ�<���`��|��Y=[����x���%�>��i�7M�P�	.@�`E3�J��\�{.oaM:?�qC۫[�� ���	��'_���9�"�?oH����#|]`�N��x��'���'�R�՟|�B��=��ԁ�H\�k�x����ş�+ڴ.bd�k��?���i��O󎕃��H0
�H�aREM��&o��Ħ���4E���#
�Ƒ�<ʄ�ڶ]I����vY�d(�],e��4�6�ɪ#Y��O���?a��?����?���iP"�7�<rv�	7�6nM�t2.O0mZi��a�'�r��T�'ll�� �S�HXCic�욑��<1���Mc��|J~�t�@�!"�)�����+N`)�ܖ �1#�4Y�	�2�xpP�O �O0ʓE::�y�l,x��$�tfU(-�����?9��?I��|",O ��p�V��O���HDNW�|�#G�0(w�a���O}m�\��M����M��i~d6M�1x�9�g�J�ص;������`W�i�
�h��eL�?m%?���&b@�3j��Ex� �p,Nx��Iğh��ן��	���	i�'<^�z�.1WJ���Ь%����+ON��G��p�t>5�� �M�I>�7�5i���Ǌ�Y�UE��2�'�6m\Ŧ瓳<�Im�v~�oF3 ~�bV�ȍe�e
�A��D�0@9���h?AJ>�(O��$�O���OƥȄ�Y�à|Zc�Z|X\*p��O��Ĩ<���i�0��1�'D��')��;_�������cȤ:��Kwd����I��M{��i�lO�ӸF�<�FWN�b�;��}0�@���`���oZ��4��c�'��'wj����Nc$2a��A~j�s��'j��'x����Oh�ɓ�M�wA�z����!(�"_s����������?��i2�Of��'}"6+g2����瑴Q���O�x�Хn�M�h9�MK�O��电��Ӂ&�ȝYU��xW  �R����c�Е'�2�'R��'
��'��'=M^Q��܉]�^å+_���"�48��ϓ�?�����<����y7ˉ02i&<��EI�b�Xi;�΂�r�6-ĦYA������݃f�6-b�,
���n�E�� �K�}�v���o�I����<����?��J®U}|�� F�@�(}�����?Y��?	���d�Ц�Á��蟼���,1�,�3��Y8"�M/n?��2��Nӟ8'�d��O�l�5�M���x2�O�ٰ��S�R4{B�@�V�y��'R*e�*�0%�j	 �_�P�ӡ�Ҁ���I1�� p7h��Q���"�>����؟D�	̟p��֟�D���')<�=�h|�v��*���t�O��?I��ih�Z��'�B�aӆ�杪�̥JsĜ6(��i����!Z���I��MS&�ie�6�;�6Mb�h��:ސ���O���E�T�&�X����
H�(!S�C�Ky��' r�'��',b���O!�Xd^�J���э,T��I��M�a��?����?iJ~���9PjI�	L�����vO�6	t��&T�|��4=���F!�4��i�h`����Cڈ$c�@ՐD���揎�U���@��<���?*�D�䐋�䓫�D�=}����k��W۶�X@�A�N�R�d�Oz��O��4���`�� ��y���*2yʥz��I�f�T�/_��͓n����Ny}R%u��pm���M{'j���\�Q�GW6=���ٶ
�#g>T�4��Dڪn�R�z��`V��֍�1%ZE"�#�m�֐�Q����͓�?Q���?Y���?�����OL�	@���zd"k�Ț�Uz��'���'��6퍸�)�O�lZv��=D��]ʢ\ ?�Y��g�`��[L>����Mϧi�.e��4��$"A�x�q�K��x�:$P�i�� �X0aA ���?�
*��<���G����FV'I (�{0,���O��lZ���	۟$��r���İ��AZ�q�*X9!�A���py��'��n,�T>u��<)��c�<?g�@�PG�Q�(�a���Ѧ��-O�L��~2�|�n�
)0�Z��~'
Õ�G��x2�q�����%V�:aφ�CW�K&��"[����O.�nb���㦙�5�C�>��B���
G�h4S ��)�M���is(�Ã�i��I6�qba�O�h�'$P1B��?����Ł��D40�'��IW��\;��R����*%s�`��-ӻ�M�q
�?����?ю��q���bZ򸐂��v�j% `bƩE��lZ��Mk�'�)�S�f��nZ�<���)<݊�l�T�m0clM�<��AX�=����ӆ�䓼�D�<A�ψ�,Y��9 gI?QWI�T(y��9۴+q\�3���?)��q��i7���B�E�o$ h�I�8��'��&��&�fӺ��c}
� z���i���l���l�h7�Q`����H�fي);� �[|�S +5��@��=�1#��V�-5��S8D�D@��ˢu���ᖼ`���Ҡ�ǟ���4>}�ز���?ᥱi��O�.R=z9`-ǆK�r�ۦ�
7-�¦e�ش]�V�� '�f���Bw�lT��BB�U����j�ug��q#���%��'Eџ� �E�b@����D��ɂAa;?A��i�p��g�'4�'��}h���
*48۱�@�<� ���MC}B�yӈ�l����Ş]���VF�^��Άf�`%r�"\��McR_� &&Ѥ���7��<y��K^,P@�
[�dt
���o�8rߴ\_(�b�Z�p�Dm]�o�"��������ƛV��u}"�wӶ4l-�Mkf(�WG�9��'GP��c/�D�:0��4�����LC�	��'o������$X	�)�Q���T�J�؟Ia�?�OP�I�Ƅ�=}v�0��2_Mą�ON�D�O�o�*1���'KS�v�|�����D:�k�e����b*�'���O��dx��	�$B*6�'?�ŭ�ae�)�cњT���P'�99Ui�F���'�h�'��O�|���)_���dX�z�ph���	 �M[�摒�?!���?�)�d�k�A�.c��@�8F��\i������OnTm�<�M��xʟ[�g�y���!��q�j��A�P�{�V��&���|J!��O@��H>���<�|������dE�k^~<)�i���j�[53Ԕ��d��(v�����O#&�R�'�\7M8������ߦ�Ro
	u��Cn��u��)� "Ƅ�M;��i�� #��i���uI�ޟʓ0�Ar�J�.��0r�G�o������=|OX��mU�%\:,:B�N-T�rب&��Ҧ-"s�KƟ��	̟���D��y�-ϳ,����1��+>�� ���6��Ԧ��I<�|�4%�M��'j|t�I^��V!j�NH�b���'��}�Hc?�M>I,Or�f\�@��NZ&#8��B�#=.p=��ɫ�M��P�?���?��%�Q�b�E�نY��!"�eV��'i��ΛV�~�bY&��[ƅY�Z���Qe���Zt:?ٓ��:YIrԩ����KM`��	�?��'�m��I�6%V:V,�q�JH�<)�e�$��� hѶ9��Xa�L��?��i8f��v�'M��i����]�~�LL���� g�ܥ�! �"ea\���M��i�`6���Q7M:?y�I���#�D�S�V�]����¢&�$�$��' џ4�U�ҜZ��Ճ�OQL4"' ?i�i]B�p��'���'������D�wr���dƁ$�D�F�k}&|�\]nZ�?q��[/i$�a�B�C�0�H!��K�?��E��o�%P�ʓ+1F�;F	�O�@�H>.O��b�Ώ�@�M�B�O=Q���'D�7�L<<����۟�����!M0>�,�b/L�P���]٦��?rW�X�ߴ�ƍo���i�ŋ7�vA�(�<����B U�(��7-/?��K/gH�	L��䧽�+��©IO���p���:��M�<���?���?����?1���hH#̌L�s��16]T4�p�܆o���'��b��P;�=���DG���%���5mߋ2��P�(�9pJ&�����ēc�F!{���cn*7�??3+�>8��(S�-4Iz���eO��{#I��L$���'��'���'�T�!&��p�u+U�B�W�<t��'�P�\ٴN�����?����I����y0n(h��@�����	���O6�Q\�|�4nP#*�lCFNѸd��ChO$H�4:掅!�M��T���w(�� ���� �tx����!�r8���Q���D�O����O���i�<��iLJՓF&G�*�޽ gP2;�!A�R�i`r�'�"7M&�ɞ��r����m��M��j� e:� � �4��m��4���̰$��J�O�	
b��	��^>&��*Ҫ�=���	Ay��'���'F��'�b]>5{�i�8b���rEj��0��Z�%H��M�T�P4�?I���?)N~B�����w	��`��S�s�N���H��
	:�hz��}n�$��S�'$4��۴�yҊX��T٩p���b��� ����yRI�
hh	�������O��DI��j�`�K��W����ىn�����OR���O��f�E[+���'`�EKb���pc�(k���!A�4V�O~A�'�B�ih�O�(9d*�	S�E�"� ob��a𚟄��(7��lږ��
o���ݟ��B: �܈�A�_Ev��f���$�	��ꟌG��'kҽ Q��0��=��/�<�iq�'^r7���~��c����4��KǸ�;a(�5Z��b��Wy��� ڴp���n�)*������E̍16��d�Q�+O����\�/k䤠��K ��@$���'B�'W�'w��'P�-�7,��%0�n߼-�ta�RW�0��4f��h���?y����'�?�����C2��K,(�"ƆR���	:�M�Ѳi��O1�:$�BDJ��&�P$��{U~�j&�8^�*Q��<�q��-�j�� ����D�y�T����a0*%�b��<LȀ���O����Ol�4��ʓ[7�f��d�B�L&d��Q�/�
�ZL��!_�\���j���:�Oڼl���M�e�� Ҩ� +n��r��Lj��!󊟱m@7M3?Q�`�+%�R�邛�䧶��SO#xKDa+ӆ��!�����<����?��?����?1��4�Ɯ{\Ĉ���&#��(!5!D�20��'��Io�fX@f�<�`�i��'�މ�C���zCrQr�/�%?��t2"�=�D�������|zD,�M��O,�S���U=���C�N
^��T1$�����Tv�Isy��'�b�'�b�K"T��e{��ӫ6�hܙrl0Er�'��ɿ�M�CB����O��'>�4#G,ԙ3�氹e��#���'�>�C�f��O�O��
� עV�{(�Qo_����`�e��D��=�@�Hy�O���0k�'5P�ڡ��?�:H���н|�����'���'�r���O��I�Mc'ʙ�
P6�g�\�B�8`�.�N�|���?1�i��O��'6M		?�����B���@=���	Ȧu� �@Ħ��'�@L{�gE�?�Z�[�\{E��o-��IЀXY��5Kcw��'r�'���'=b�'���p�|�:$ ��u�b}�s	�1ws^��޴-6!���?i���'�?Yÿ�y�G�:Kf�	�(F�P�ұ�d�H@|��Of�O�O#�@��id�L ��xcd>�zd�4(U�[�s&Dm9�0A��ON˓�?	�w�.= Q�PI'�Ȋc\���f��?	���?1���$����A�M���T��䟤#���Iv����%XY��q�Fx��-2�	0�Ms��'��'�Z���� '�Dt��ٵ(d���O��į�T9R�Q��=�)^4�?)���O�tj5�]'qL���Ќ�c=��6��OP���O ���O<�}��R@LI�*ޜk�eɰc��^y��z��Q��v�T,��'	�6-4�i�A{��/��h6Iͷ@�08qF#v� ��4�2�i��m��i
�ɶAJ0\Y��O��-�\;Θ���G�j^�#�G�`��]y2�'�"�'^��'���	�y����B�Ǧ'���^�Ā�4N�8���?�����'�?�`�cҽ۰�œo�.�۵Ã����M��'9���O-����Jך*gJ�� G1�~���Rbt�	�R�L�����N��&�Y��Hy����NAD�Q�ҤD����!�G�b�'��'W�Oa�<�M���#�?itC�ܲ��YV�4�P�ێY��<�	��M����>i��i�b��f�N�)�e�*�r��#�29]�H�I5?f6�,?	#Q'_tT�IK���'ѿ�R�2�2�i@�[�d��r�c��<!���?y��?1��?Y���*L@#b�!�h�6\6dd-�G��'��d��M0�8�@���M#K>15��0����a?I��P2ǋ�S��'�>7͘��)��
6!?5�!U�$ڕ�-O�"���㞝%"�! ��O�ѺN>	(O����O���OF9ؗ T�Yi��K߬:F�2��O�$�<�U�i�H�A �'��'�哷:�|`�+X	,'��e��&�DJ����M�A�'!����2y�&�X@�.wت���D��!�cZ�L�.�
Ǣ�<�'f�,����T����!��q�$H�C�"<B���?����?�S�'��$�˦U��f�+�(�HGGðm�}�Q)�t��I͟���4��'���FϤh1ٸ���6/��IF�ĥ>t���pӤ�KAam�z��|]+%����$c.O�ty�g�Zr��?�l B�`���B�+K�[s��4,�a��D������4�T� r9��[ %G�mJ,1����X!r�O��NJ�x�E��@��	/Ŭ��'B�qr\�Q���je��z��qm�q]Ω��\�/@�ĸ�,��� ��d��(�%XC�J��*Y��o�me�I)r[�;h�dXQ�@�p��	 슩P�Ή��_�#	���ת�<ܖȪ%h�#}��ӣK�d���`Z�y���&i��y"H|
�S2� $-�q��ߛGX�*D��
BnMn�����I������']���)�70��B��,
�)[�Jr�����C�O���O^��3����KU�EH<9pA�yQj� ��D��Mk��?i��/�p����?q*�|�d����Fцk�&Usb���dn�6��'���+��,���O����OJ "".M=`h����c[��´`Ц��	N��������R�D.�MK|:��LG=`Ϙ��햿'����'fF�25+���D�O~��Ol���O
�a�@VSD>=��ל$~�p�do�=@˓�?���?�M>����?���7yO**��]�<�np�&'j��k K�^~��'���'���'6P�dݟ�YӡL3z����2�1T\<4i�i>�'<��|�'=��	!R�H�4��pi �	M�:uK��@q�'*2�'6�'TRFx]��\��V���E� �v�≙D��M���䓪?��JH"u!A�C�I�.��T��b� 
��R�і_ְ7�O2���O�$��]��'�?	���b�&^;�H챕��"�*�Ӧ�	��'D��'�tL��H�6��I��n��$'�x1k��GY���Q��C��&�M�Y?����?���O��P���M��ܡ�g�B��i�5�i+��'D���2�ӕQ%��R�!�.� d�Q��7�\�FKB)n�˟�	��T�S����<��eK�`Y,�*���Ih��T���Oś���[��O��?��ɥ,�DU8E�X�-Â�R�����J⦉�I埨��2\��aR�O ��?��'���GI�?��0��	�:	�~���4��C�f�������'�r�'��Á�����&���R�p�aU�{Ӛ��ӗ���?I��?	M>�1q4��EP�f�]0��D^��'����|��'���'��:oz�P%��3xX4�5I�.	�a�����<�����?��p� $+��,1���*��%�!�Td�$�䓽?���?y(Ov�P���|�3���܈�T` �(E"�;0�@̦�'�"�|��'�%V�T�$�Otę�()��Ǩ]�+�	���	��X�'Pj(�~��Ot��zwk��E2ą�ׅ��;��ǰin�Z���	������iO����y�d�a'�(RÂ۲|s�9"�[���'w�_��ᡢ�
����O�����Ɲ��_o��b��C�2H~�(��d�	ǟ���ck����y�IC25+G*?4!�M��������'��R�+e�>���O���ԧ5��];r��&�Z�#��N��Mc��?���S�'�q��A�b 5��ы��q5V 
u�i[:��,t�.���O@�d���'��*?�Lq��\-����0��%b6�h:ش]�Ve��I�Oظ;�j`R��[Ə+y���a���Q������	#cΐ��O�˓�?9�'��+�Α-R0���fʇ��([�4��C�����D�'���'�
tK�g+e`�IY�<Y~��wf}���¿5*��'b�I䟨$�֘�otIY��
l�*�FZ����P�e�N>���?1������!v�,�p�.��k�	�d��A� ��V̛M}_�D�I�	��@�I�H�
�F�+qp��3E����	�g����' ��'��S� �a��#��Td'QD����93���I��M�,O���"���O��d��+�	�
ʒ!����K����#��y���?����?�(OF$�tiE_�Ӳd��I�]�5�P�Pm�;@�p)�ٴ�?�M>Y.ON`� �O��O¼p�G���Ĵr�)�/Րy[�4�?1�����^��'>����?��a�n�(`1P6yۑg0��O��.*|�b������D�C9����5��YV�����M#*Ot�xEHTԦMث�f�D䟔H�'��az��ʜA�J�{�$�JbLJ޴��dF�^)�w�p%'>�'?7�׸L��D[6�S�qz@��GL>^Y�6솠h8�7m�O����O��	�p�i>m���	(d�ٖ��
I` j�ȋ��ܙ���֟�Iby����'��a�O� *����]'@�"� H.27��O���O$��ɘf�i>I�Iq?�k �g�٦k�*ƬzH˦���Wy_Z�X��<Q��?������o�J�@��ek��iUZ��
"�x�O�"�|Zw���YՉ�,me�$�����KN��ɯO��r&��M�K>������O����uBB�pU(� �v���i��?��˓�?����'���'�.�3���/f�P[�揋5h�h3�+����y��'���ڟ���@oj�+4|��b
;u�u�������D�?���?92Ə�y3$9nZ3}� �wj�����0v�LOV���<Q��_f�ٰ/��$��p�� ���d��G75��mZ^���?���T7B��d��O≥-E~���ךW�t��#D��6��OZ��<�v�͖V<�O9"��5Ƨ�!����v�������䐿�V�=��?-���N�ke68�*��-b�� *gӾ˓}f�� '�i�r꧳?�'1��3oxr�ȆA��lC���.s�6-�<�j�!�?Y�����4Eh� UJ�8s^�9�����>�
1m�&�HE��矸����tyʟ�P�@�R����*܂b7B�##XϦQb�J!��b�"~2ڴ5r�
�1���1�-�5&46-�O���Oq��$�<�O��*�"h�k��0�˲�,K�T P���Y�
Ī�'>i�I��d�	Mh�L��BEzM�py&舝y��Jߴ�?)���Z̉��D�'�rW�H��&�r�ҵI�c�&F`'D�&�M{���������?������,F|�#���b���`��0���	e�Zy�����Iu��AyB�T�|0P���a�p1w�
�QD���d�'.��0�Iꟼ�'����jx>��� �Y����"� 3�N�q�M�>����?q����$�O��DQ�	J���D [#d�(�#�]�U���	o�z��'���'���̟����}�t�'!j(!��9����2�Ǉ ��	�j�P���Iʟ ($�a�|OP��J�5���c!C�1U��ói���'-�I�Y���HM|
����1���a�K�. �6��!T, o�_yb�'�"� �R���D��5��Z�s���٦!Nv@6D��e�%�M(O��ɵ����s�����럘@�'b|C�d��!���q#��9^n�Tܴ���B�O���$�`��^�D�Od�	k�5��5� �O<^����`�i�|h�v{Ӝ���O8�d��>l'��ӨX������	 u���[�G�%�2x�ڴ^N�p���?�(Oh����O6|{���!�fz0cL$'� ��P�\צ���̟��	�5�J<�'�?q�'V��(u�[�6�h�W�ɤk���4�?�*O�ex`*�Ob�O��䳟H��v"���
_��2��6%c��DX�V˓$��N��@��U"#�Ԍm��*vj{n$H0Q���Q��,\N��?���?�/O�I��J�v����I�g[��ٗ���`�t��'D�	����'E��'����:��A`i��d�DI@� 9`�@ژ'���'�b�'��s�p��g "��T̒V��Qq�}������Q��Ms+OZ�$�<y���?a�� ���Γ6�t�k��G?Z�&��ᖐ/�pPBֺi���'hR�'��	�3�P\������٢~2L0R�☖3>P�ᗮm�4l�џP�'���'F"E���yb[>Ic� ~͙�bO��pa�?`?���i�"�' �	q%�lX���$�O��i
p�8�(\?AyP��R!���Fi�'���'���Y�yR^>�	h�s���o�PG �Q (�`U��ƦQ�'�p��dӈ���O���$�ԧuG���V��@*�c��-0 Fյ�M��?Q'N��<�VP?��b�'02D��
�
�p��"<t^J�ov�Z�Hش�?���?��o
�Ify"«�����f
�
�JI���O�4��6��?$��2�$5�S�芲B��lT�d��6F��Yw�[��M����?��1�tk�S�T�'��O��)�$�* �� �#� t�V�i��'�����i�O>�d�O1g�)��;���5�������I�ɇO����O��?�/O���<(�Q)��kN��v�+�[��S|���'��'��R�A���8�j�d��f�2���SF�i��O���?I(O��$�O���3����D�	YԼ��
���q?O&��?����?�(O )��J��|:� W�h�a�e�X+tcz$�t-
ܦ͖'��R���	��IU��Z��D`��n)�x
ԫ�,����'��'rW�	qŬ��)�O�DI�U1���M�j�l� �֦%��fyr�'���'K���'?�I�b��pɕ�*eEZ\)�G��,ڴ�?����$|Ph��O]��'��$וyޭr�F�2K"0�`��>i�<듴?���?Ag��<	+��D�?��4�:����ۊ5L��Ԋq��������i���'���ON�Ӻ�=E�I#�C��l�
�ɴ���������0�9��O��㑉�&a�b�x�N�~7��P�4Y�4�i��'2��O��듳�d�|}�=z���.Ƽ�	�ΰ6��o�\�����ܕ'��z���#,� ��"DԃaX���&�B��Tn�ϟ���ߟ$x�!��D�<A���~��Þ7�<$ ��\�@�T��"eG3�M�����$>�?���柌��C(�q�3lm���r(ɤIː�oZ� �!�����<I����$�Ok�%*�l�CeM�{�̩D�H��ɺ%�t��?i���?����E>�2!���HKrUkb��(,Af�3�*�r}[�H��\y�'�2�'�>h5�R�tF�t��I� v��LQSh��y�T�8���L��Sy�W�5mp擌P�A�pM۴F*�q��Eҥ\�7m�<Y����D�O��D�O�� =O(=����PN�1��O]Q�( ��Ҧ�I矘��ɟ��'8D�UI�~"��d��@HI�5�@����'o2 ��i�W�8�	�����t�|�	ҟx����ɸ�Ʉ��M��_�}<�lZ�����py�Z�Q
b��?�����'CC2� 11���gX6ט%{�HT�''��'�bl�7�yB�'���I4 ��E����%�
�BDP�A�cC��'�|(��oӨ��O����H�էu׎؛~��E��żJH0�J��8�Ms��?� 	�R�'�q���rĢI�Zrx��c_w�,��øiϢ]#$n�T���O�����r��'��-ƚ(�F*k8��Xdk�[��A��4Ò�ϓ���O�?��	%be"sO�%l��8��P<(_�(b�4�?����?IתX9/��ey��'a�D��
�9x#�d3�/G<���'���3G? �)J���?��x��&*Q-�*՚���8 {^t���?��5��Ly2�'x�L��"(Z�k��d��zf���c	Hz}R$��y2�'A��'p��'R�I*6T����ĲNT��Ƨ�5V�X<a�L���d�<q����D�O����O�|i�H�Qہ��0�N��D+h��<����?�����۱M����'VkHxFC�SJ�'f�	\e��nKyB�'x�I˟��Iџ( R�g�����=��*�f7b^��Ё�����O��D�Ov�o���#�V?���=��P���$�z�sw����Bش�?�(O>���Oh�DNLZ��o?�	�#i�,�u�ξr�Z�DH��������ܕ'kN���~���?��'d��Ͳ' äs>1�S΂0S��S�Y����ݟ���3 ��������ϟ$�'j\�|b�)�(��d��$er}n]y��F#&E"7��O��$�OL���d}Zw���yS��_��1�G2V�@��4�?���^�N��'d��CܧzyL8Yamχ�N�s�iH�5�l%nڙY�����4�?Y���?��'.��Py��I,o�0����
�,�z�6���`_�d�O����O���4="9 �eߑ$�:��L��7��O��$�O���)�~�	�d�	D?Q��($d�p��ĤjMpl�����$�x�c�����'#2�'�Zc��\��%�0V`�
�ϋ�p.��4�?Y �Ӵ=��O��D-���ly�c̛h "䢤��^�xPjs]����Ir��'9��'��[�P*��2=�*�ql�:n7�aAC�eψ��K<����?I>���?�F��cO����a�ɒ�GK/�Z�����O��d�O&˓%H�=�e;�B������u֊�kaLI��F� #[���	ӟp$���Iӟ$[w�Fٟ�����i�n�Cd���XrL��c�;��$�O2��O��"t�&��TiZ�}	���/�:�2��0_��6�OV�O��$�O��)34OF�'�X��H$��P�ꘗQ� L��4�?�����G�+�&�$>}���?��ѧ��l��A�↏kf�Pq�����O~�D�O��zb�O��O��	#���'M�?��5�#
��@�h7��<9��\���掶~����:����QȄJz ���v��c5�x��d�O�ѸG��Oj�O�>� L�� �6 �-��_�hq��iv��l`����O���b �>mj�ⱨ
�y����Qi��hQh7-�,wH�2��2��՟8R$��{�4�H�ǩX���s�I�Ms��?1�:�z<I���O0�I�Fe$�rW�U*	�T�@DW�p�7�,�$���?=�I˟d��q"��܈+����q�d4m����F���'�"�|Zc(6F,{�1�N��+Z"��O^�u��O0��?����?�,O��:�DT'5�L!���Ӫ9� %�D�$H�x�>�����?�uG�-���
Al�RTK��,v()�"�<�(Ol�D�Oh��<��ΒF(�i��N�)�smf�f!�7��.e'�'���|R�'�b�Z��d�+yI$`j�@]�5��H���6Z������ԟԖ'E��3h3�i^bJL��a��g�jH"e�ȉx���l�џ$'�@��џb͟�O^D�Ej��>ej<�&Ƈ�"^uԷi���'��	 b T9M|B��jEʇ�)�BEȆf�,��!�� M'Y��'	N!i �'��'��� +BǤp���+��".
)��VX�������M+�Z?M���?��OZM[Ƥ�%�!��X&�N�;�Z���'e�'�ɧ�'�p``����pH%h���l�A�I�޴�?Y��?��'Љ����(�-�7���GY<�c [7L��?����Ş�?E���;(80'���՞g���'���'�|��s�"�4�T�'d�� ��I:d��F5Z�N���4�?QM>i՟���'�r�'<�d�g: Po_�[�6	*�r���D�'c:�'���Z�'�0|rb��)N����ݹ>Yd8sO<����?y���?A��?�-O�E�
e�,�E��\n���v	J!�|%�\�ID�'�Ę'��Lr5nM�X��k��W��'��ٟ`��ߟ�''���j>�D�K?#�$$D�R���PnjӘ˓�?A/O��D�O@�$�kq�dٗJd�D�R�86z��] t���n�П�������IRy�ʺU�ꧠ?��&� pJ犟l�e��I:��lnZܟ�'N��'p"�O/��' ~�20F�ۂ:3HWoԸ���4�?������ϔ+>��O���'����@z��k$��$Q���Z��L�H$@��?����?����<	�����?	Y d����xC��OqVe� bӆ�P�P}���i��'���O'V�Ӻ��CU e����FE����馭�����*!
c��:���d'�ӄ?�X� ��X�R �T㓥G�7�?���l����I� ��)����<I�bJCRj�2Q�v�T
0"���փ��y��'�Ia���?!&e��+��\�(ްl�g�'_қv�'�R�'u"��d$�>/O(�����Y��.O��=AѡW)�~ȓfIm���<���]�<�O'��'���;w��)�s�BM���r��oL���'���"&�>�.O��$�<���[ք��.�(�W�.�L��/Ȧy�ɴ9���Cy��'�b�'�	�}�� �C@�
�N��Q%�0 ��`����d�<�����D�O��D�O�iB�,�Q�T(�ů�~Y\Ԙ'���$�O(���O���OP�+����;�������x�Cg�@1"Y�iR�IƟL�'S��'��yZc���ӧ#!>�yʲB za�ԙܴ�?i���?����䖈4��h�Ob�1Z���cJ��.*��	��&1Kf6��Oj��?Q��?i���<���~2g  W�H"f-�jXv���M��?�(O$�!! �M���'�"�Oh�3eF��@�����@8� �0D��>��?��H��Γ��9O.�ӜW�R���'�����Tz7-�<���-2�f�'���'���ɢ>�;F�P�Cr"�k���� �5hr�5oZ�����0<���{�	cܧ}J��J��)U���*T�H.���nZ-�P�8�4�?a���?���e��	QyB�T�5LJ�P���'v���BƖ�dkB7�\�J^��O�ʓ��ORҠ�_{40v�WD�y�`	��c�67�O����Obe	f}rU����V?�r+ +4|�E	:4�T�H��M���Fyr/1�yʟ��d�O�� A��c�H�FӞ9ۀ*>2��1m�؟(��Mڍ��ļ<Y�����Ok,���
��Ƒ�-Қi� %�5�v�'��Q�'R�'��'x�Q�ѩԉ3A$�n��l�� a�G&H}#�Otʓ�?a.Ov�$�O(��_5D��0nށV�z�*�h�;m!y�8O����O��$�O��d�<1���7K�H-6s�<X���>B�xQ�`�2�FV����JyR�'JB�'�,�K�O����τ[�Lm�wC-w�
}��R�4�	�4��WyrAZ<��'�?�� H	 Db	BE��lh,�Pǖ�4��'��Ɵ��	ȟ`��.`�x�O�[��/Lr�0��?Nh�ъf�i���'���'��b��'�b�'���O�����i
�]�ɒ�œ:(�y�?��ORʓ1�fExZw1��(�m�%T�M8&�I+{��ߴ��䃏1O��lӟ���埼�%����n=2��1ˠ"A,�l*ȅ�3�xr�'�ўd�O���R4Bj
3���#e�"�kR�i������'f�\�d��㟜��ry���Z�$"����'�V!I�΀�Q��J�Fx����'2�piq�O	+�!��hԌr~|��buӤ�D�O���`�С�>1��?��GW��і�՘ ���� ,��'[�9ҍy�'H��'*� �w�ҙg�pX�T��P�5J�W�ܢ�̚ay�R�X��e�	�:�dQ�[��(��fn@�e��hK<qd"~r�'z2�'��I�L�|�s�`G�JK�Ps0���g� �؇�G��ē�?I��?����3}���B$@É �L{ �Xw
�،y2�'��'"�'j lr�П�]3�h��r� �//�,�ѾiB�'a|�'`�0	3P6�0���qZ�
>�2U�G$.��ß�������I؟X1e"�E���'b:����	�*X���TE0NX+�c��)���O�U�~'�@Z�O�z�Q!��;�
����bӊ�D�O�˓_�(�����T�'��N�a��xv&����T��.J26�8�ɀ7:#|J���#΅�R'�$�A��!2N���&a�����OL�C��OZ���<��'��ƨ� ����������!K=�UP��iE�S��vC=�S�<N�дa�@	nؐx�F#��-�87M��-^l������h�ӕ�ē�?م& �0�%ٞ*}���
�\��F�Н�O>��	�L	
v$�,�,@�gIӪKzܴ�?���?�/
�<��'��'i��G$ZhL=h�"�N���Rq��	u�O�l#���O��d�Oj�i��-{�d�
��M`�!�E"����I�_�P�I�}B�'kɧ5&�Wa�7��")��*=v�	l�Pb����ߟ��	dyB T+�Dx�&�
0��]����3�,H5/�D�O�d8�d�O��ŦM, 1�嗰O�}�Q���Q������Ol�d�O|����3>���c���5G����-U�> y0Ӝx�'n�'��'7�lèO�uf���'5��"PN�"Pu��U�<��ϟ���Gy�c��\������,5���936|��� #PզA��}�	��D�ɥT־c��!\�A��H���^�tq�Em�4��O��4J�P6����'x�$\�t��ar!߰�>��`@�� ��O~���O:���~�@��n����%T7#6�R�"�$;z�Q;րA&J���g�5�%	t���0Kx�CF�T|,���,/�8��KWDk�%H���gg ��2 -�Vm�� Y�.����6��#�����ӋW0���s_pP[�	�i�X8��H$����&��	[�tz���U�V�s3i-cw
)x��I�]��X9��C2-�N �7$��cƔ�$�H�m ��'� ]��oe8>��GS�AL�4��]�]��`����?����y������O�eI���	?xd�a5Aަn\���g��d=�`��`�a3:���d\��ND�'>��b��'a�B�li^��j%*l���Ё@4���Ѵ�2����*�vt�V$�If���qB��4���!"P��	��`E{�U� c'�EX�Ĥ�a!��+ P��,D�,��jÛBM�Y��>g���p�	�HO��Sy��2�"6MΦr�>m�A<6�0qr��4p�����O��q����m�ON�db>1`1�<�:�+Vk>Zv�r��K�^R����7�,e�3��qx���B� ���Ӳ�A+dDd@�CĤS�A���X��0#�"�_x�\���O���kߦ��'%=S�vh"���0r���=9���R� �XX���(�
<��O�!D�!�dX�U:F���������Q�P�Mv�v}�_��!#`6����O��'fwz����D��������Ь!����?I��?Y����&�\s�P$*"������K- �G_�3�"��bF%�Q�d)q��6�܀�*���$>mk I��N��T�	�2mV���*4ʓy�B��	����D�����2�Bۤu톘���Z�<�	����肊Z.C<��2関�0X��I��ēDz8Ub'�|���:�A����#֎P��R����m�A-Pw��'�"���iޠ�����*Ⱦm��*	��;u�W +�@,ړ*��_Q��T>��|���>����"�܌XP�0�2h�yh�ȓ&��\ph�p���[xŉ�IY,�"�>���?kp���V���*`
,0���M�W���\��M~J~H>����q�	r�,�!���&0�ц����Ju��7��ъRhÞ4� Dxb)(�S�$'�7Q��JDM�Z<���R�&$��'����Ʉ/u��'�B�'8��ٟ��ɛ!i���#��j���N�"���#(�.�
I�e:@�HǓW��-��S��b�"e������X�z�9�E�{,���'����F£H���R T-{W��c�'E���?����<�3m��j�Z5�N]ݘH�O�H�<�ܓRS<LR��O;O��y�ń^%�����d��v�loڗ/� ��� v���h0��/�@L�������̟�vd>��I�|z��ǈ�M���x��#EHϾ:����k�8��ɸ%�8�BM��A3E
B^���Sh�5M�pK��'�V4��`ћh���h�hތM�X�" Š0��6��O˓�?1�ʟz4:�^%��䪐��
4A�"Ovq�U�O�E&�U���E
a[]�B5O6���'X�	l�vZ��*�d�|��P,�@#��+.��Q9a��H��z��?�������B� c�X
�i��8� ո)�� ���BBP-I��m+�DW;dT�"��I�8J|�A��4Y�z�J��#8���>��ZŒ���*�V���N?�����O>:�:���Ę���H&K���'
�"k�-\5����+[]&��$K]��0>Şx���b��k�	Ls�Z�<�y,F���?*�<�����O���O$`S�� �Aݬ�)ȅ�'��РN��$��x��bь���,]՟ʧ��?Y��;49v�LuP�*1�P�&m���8W�bI!�`K����OB��a �[��P�S��',�XB�'D���D�OP�S�Sݟ�'�vA$.S*}�T c�S(mx0��'���o���n��Ab���q���Hi�'���wwz��@�e,��Q��9��m����?��n[ 
9.����?��?a�������OJ�;�C[��^h9 jEoJ��!E�O��ѵD�	qD\���-jb� q$H-���Z�J@�Pt����%��9�8lO�J刞�k���P`LK�?�n-��OM���'s�{�	�?4aQ`N�]���ǅ��yb*Q1A��3&cәXaV�+�O�6~Y�"=E����
z�7���&��|��M�(���"�,J��$�O����O�ӎ�Ox��b>�	"ŝ��D kC̓&O�K��e���;�4��l�q�'��9��}>���$VQHIM"fP25P���l�.����MV��E�U��8�E"Cm�5����`Ə8�M#�B4��<!�hB�idt�*z�<�7K�C�<�dK�U��dƟ��h�]�<�2_���'���%�|�p���O��'���T��d�
ؙf�W�^Sd�#T��:�?���?iE��!�?Y�y*��a��b�{N �y'G��R�FX"G�I�E��
A���R!v�@ҭQ�X�k��x�'W��+��h�r�@�d�{NPe�,�"�����"Od�[�n��OC౐T($c�E:��'_�O`�����^v���3�@4O��"O�9�e�o����@1o�HH�"O�
�i��	�p���]�n��}��"O�u�����܁�o4q��A#g"O�ۣg��)�r-`SȈ1H��A)�"O��� Br�;���7	b�9D"OH�ڠ.Y?؈�{vIƙb�\�5"OѲ�f�SP�bhQ0A�����"OJ���f��=Bs���t<�ۃ"O�tH��S�2qd�w��x�uk"O\lJ�l�Ԇ�����yj� aF"O�$)��#?���'�
�b � "O��zG��=&V��d�\a^`�`"Ov�sV���;�R0$�<KJR@ "O���T��Hr��
�B�3� �"O�
& �5�[B���Y"�2"O.qegj5��G�9|�����"O�u�Ѫ %E���`�-�:Jٔ��a"O:�wF	��Zy����i�����"O�����-^��|��Ȗ.��Xq�"O���f@ШYWF<qA�rkF6"O̒�gµ.���WF1ax�4"OY�Bj%܈8[��O=3��`��"OЀ�t�R g��(s��B�W����"O��;d�K4-{j��$���MH|P"O[�R,�H`�Վ#=�4�"Ox�X�톻<*lXp+���ș@d"O����H�6Yur�Y��V�E�d��"O�Ż��P�]+�����6�P"O����O�4J�CP�U�j�c"O
��qDCr�J�+��/�%"O�l�E�ƠL����䏚o����"O�i���q�5�Ӂ[l�XzD"Ox�Ei�h^ jr�K-v��E �"ON���k;7� Ʌ�׷�$��"O(��V�H�У�),�%�b"O�e�E�mbej g��>�`Y�"O� �`�BᎧj����7��0C�4��"O&Р��x�Q�0M#:T�R"OVYK��ʊ,�T ����~�TP�"O���Q�&WV��R⋴<��5��"OT�Bv-ߕ
�>��tg� ��a�"OH��U��08�$ժ���T�nIPt"O|iAr�@�d�(�Z�C����W"O`�q#�'�� ��A| ��"O�Hsaɐ2�k��ȇ"f����"O��`5��&0`{e��1fF�؃"O�t��aWv�@x�A�0s6�� "Ob`���1,�]q��mJ��	V"OPy3ÊЊ�V��5�E�R"�%
c"O��B�	�SД&�èT^T "O$-��A1KwbP���F=-ԸeQS"O�ВgG�$R�L�"�D$ǜ��"O��#���3WpXHP��K�Y�!"O,������2F �6�@�#"Oh�Ye(�"V�fQ��K�K����	�Q�	"eo7��Z�#ł]�Q���3#b־��B�I��4��`mٞV⠩Sq�՗1Ӧ��o��R�M<�)ڧgk����A�'[��k�d�H�^)%��+Wd�L�N	9��i�2q�0�u�	�d�;���w�8��Z�ZCx� �U�D;1&Dkc�ر\]���JXX�%�d;�%�j��˧>��M�SK=6��{Ƣ��I2Ԫ�'[�p�d��>8Rd�EAL�m_�2�G�J�#$�)��G[��I��i'V�Ū�o��݅�	�m/F��E��	��D��O�,�ԩt!r��.�ȁ$�O�]�ԊE�g.1O?���pv@K��ǅal�i�"O*����D�D�n��q	�+Cؠ8��x�&S�:�	˓ai;��τ>�|`����8�ZɄȓ ��y�����}Pn� �ַ r����D$�$��e/�e(s�óR�<��ȓ{2�$�� E��w���F���ȓN�l0��/ 6,Q���p�j3K8D� ��
�lVdT��K��Q��p�0�9D��R�.ݹ*p��yʒ#W�z�a�+D��Ӗɋ�&�ܡ鰏�@�f��֥*D�l�r��H�u��1FWH� �,D����у1�� ��� ��$5D���@��`^%W��2�2�pT�6D��	Bm��
��}�e �6��['/:D��!�Kȇ!$�z�g˜Y����8D�(�!�Ec\񵦌9kǔ��S	,D��Gk�� Cw�˕]�px��6D�dY����P�4�y�%˜=�x���?D�(��F2
 ��"n���� 2D� �w
C��X�E�?8�^�1O�8:��[�,j��u*�*;��$�"6!@���}�=�2	��,'!�$�4��Z�l	�f�Z1[�B 4��*Ť�"6N�D`*3 �=� ��$��$)w�.i���fD�! .҅2���*׃|I�X Ƥ@�2}��b�D�G�g̓CN*`���8=�:4[E��L��u���GF:,� A̗oV�)�B��1�j�SE�A�\�� �f"�Ɇ�	�R����1�z�޼j�(���ቹ����3�� ��$�9",�ɁDꕒW���o���"%�G!���)��Yk%n!N�6%+"c�'��*F�2M
�DǸ3F.x���7�9�!���Z�_U,�&��j`�(��FҶ5�q���%7��!T��@���"�mZ��F�(�HD�J�����a�L<��y�B(��_�p9P�H�*A$����}�R�R*3P*�*4�M=���k]0+�R���&��h�>�D��|Z4�*sdƎ�~2$:�nd�u��<h��2�Z��0<��#ڭ_ ���㍕M�*U̓��x����,Q��\�E�a�:�'b�$����)2B6t*�ˋ?�'���o{�Qr�%`��mIC (x�N�b���8T�$8cm�x�'0�p{�a�Z�? �y�CT;�a1�(�� Ⲅ�'��\�:C�K6��$��(��Ɂk+S"�]��`���ٷ��=�6��2!���	$��];��ر�P$�-�iލ�q�@�s�f�;5��$�`���ֈX7�;Cg�S�H���'+r�p��QMn��A�U�Y���A%�'&��d&�{|Ȅۉ}���vp����윙2�N'khl!ق��4�<�b�vHU�#� S���&�%G��� T�<��U �&萢̌�a ��qg�U�AZ����o�5=�P$Ve�.����f���@܂��3�%)�P(uO��)�X�NZf�h��2U[����Zr�O��ZE�ɮ'����`�BV�t��S	�q,��x�ȟI�.%bKןyP���>���?'U"��+� �|����lV��3�%C�<���-Kɰ	���'�2%�'� P9�Dxމ)���/5^n����R�7���9����r��P�햚],�{��X���OԵ�${�ޙ3a�-W�±yG��1�"��s��Wn��p�#������ιs�i&�a����#~�D�_wv��Sc[�bv�l�8)��̞7�Px�Վr��YǢ�v���g[4
�����0���Se�*L1&e�Ů2e���*[OT`�5!���rm$)E6�#�j�')��1�c+�YX��ad�Fs�.l����^ a*�GTx�i@�m�����R�Dd��O�Ʀ�Ҥ�u}�A�J|�'�hm��o�P��5� �� a(�0��(lhlc�06~4�&���|�]��H5+�3o�� G�B�$]-�J1#�/���W���<A�!��&@ e�&K�&̺A��5@��(҅b$0N@�ba۞L^}�{}���l����/�����*!^\�@�W<��D{��T`�a~�*2J�F��6�+{]�sF�\�e|<<��Cܶ�����O�,�����>�6E�֌��|�C��^���'bC�-MH=Ӥ��7 R��8Db�x5(�sD%?�I��\C��[�G,&��S��r<Т��qQIA��^K�N	Q$Ʌ*~����$Y�4��\�p��?��HB��O$N'��q�Y�`�L�N3"��Eꯟ$ۀf"0x�1��������� Z�i�& A���ΓN���/BIttJ����"�:l�f,M"5�`IW�k
�*&�3<O��ӱ�ζ%?������n`M��]�mY�KGO���f
�&��^��)�MأU���l�	��NpC���`�I4�V,Q�f�:�0?9�d�Dxj�A�H�6/�l�7`D^̕�t��> '��j�Z�x0UB��<a�3����'���i��)&�����?nzD���+��P�ۓL��Y�'(����@І0�&�h���O/���Y,��MC�<��&�W�&1T9�)�	���5���$���uȃ#�n=R�Jؿ�axbn����Rq�B?q��s'D0Ja
�~֮���Y�D4:sJ�T&@�c�J�1*iFR��+U"�Sã� ʺq�e���L̰2��t�%�2I�.��e�O:�	�T��OB\,��ƜM��E�rL͡6�*�����wFQ>��t����l�B*
R��0�5�����d�5�P���O$R�c0c��TAtC[��xi�	���y�SH�<�%Af���O����j�1��[��:_J�s"����摔'��}+Eƙ�2�D}�D���F`JϛX�m������\�M$�`�޹uL����Ǘ��sU;h�vt��F(dS\�	���!	GP���`W�	�l��D�e��8u�Z!I��Rt	��|���³�!��&/q���o#Q'�]) � ;"
.@��L?�y�'x����S%�<UѤ��H��QD"���(�~��qᇞI��h'�F<8c�$���_�~雰恫6��Ł�fO�h�~�)�oݾ@Q(�}QжB�W�d-���'o�jt� �����,�S�'-��- Uj�"A��dcǈ�zL�g� V���d^6؀㵥הa��b�b�]���U�Ѽ-;4�#r&��{�����;,OvI���]Ow�D��!]>*<HCJҲ[�X!80"P���`�HˋT$$,�a��C���I!x߶a���߁tɀ�X$O@l�FO� y5@��zXt�* ����9�&	�S����|��EezB)HoN�x�h���F�M�<A`.ǽ|7�9QuZ ?F�vK7@fr��s+�3����kԂi��QC�t�ӈES~H��w�T`
@I�3��qS�T)E�� ��"�@W�����c0���&���M�'�P��-P%P��q���5s�yET%P��TjpQ��X�y�������1eP���,���ه�Z<RNqZ��|���I�=H�����y'KB-hT�w�ڎ+���!-μ�y�$T�:$D��,�^�P��	GRu��J���M�6 a���>,T�V�pS�>q'��+���0��&%�ذ AUF��P(��DE0���4倅��GŪD"�[���#��m�T�H����P>0푟H���To�h��(����>�y[*��F��2֐�Fm�;/X.�o�~
4��&$<�I@��G�I�:A�� �D��MB�'������|Z��.~���'(���"/> J�� �'�D��)&b�~=#'IS5b�䨒�'�](A�*����"��a0��C�'mV��Dh��A�����QH.���'�lm��CϏ3s�%:��J�D%��'�l�{�m�+2@xӑ���5o���
��� 8p2��;?b��B0�Hm]�T3�"OJ�x!��+�n��E�;KB�Ͳw"OV��N3����˶`l�p&"Ot�P�ś��(	���[�Z���s�"O<�`��0^l\��[�N96 � "O(��#M��=�x㠌�R�.��B"OH)CGғ:��<0"J��Vpb"O�LS�p��2��'I���"O�8`d��W~���"�,<��"O����!Ҹd�h�b#����26"O���	�x�aj#T 4��<�"O�I�'I�b����5ȟ��x
�'�p��!��w`�� ��Ts��
�'Q����'�����2�t^���'�z!�+b7���$cd���'2~��d�8r!�"�^?���'�:�2��B+C��y�!�+%�.�*	�'~�q�����~�8�Q�k���'0�̓���L�а���&g�j�	�'%�-���U�4 r��f�����'U\�d 7�Th��`�"���')b�z �.PG��9d.I�$�*�;�'0h48^H�[w55�*�a�n���y�͈�6�z=��jC�1��-(錤�y�XT�A�rOҭ���K4��y�d�1���J2/| r#��y"eϡ?�*��pI"L��C���ybP�Z"��[�c��\\�s�P��ybA�8��5�"kP�����#Y��y�ɕ�A�񐲤�=yجV�Q��yҬ_�	�81����pr�z�T��y���K���q��l�����	_��ybʺNH���-�Q��U��P��yb�J)~dz��ӤPxBk��y�ه	0b��-P~����$�y҃ �&������F�@�x���[��y'A�.����<s���;��#�y�*��m`z�k���+o�
|���y��<r� ��FjL���)b�ߢ�y��oД;A�ňfr�d�֠
��yr,Z�McD`�cA�b���a���0�y� >K* ��O[�d@�j���yba±p���aC��e50dr�m2�ya�8��YJ���Z��e#�bӺ�y��%��Y+ ?�z�ȏ1�yrFQ�F�$SE��,=1 |ђ�Ϩ�yr ��+��@����7k��:w��y� H�*d�D����6��͈��y�ʛ��6��un_�{�2������y�I��24 ��2��'^NQK5�V��y��ȦnS*q���ncB}Q�W�}N!�� c8tA�Wd�r�:��Ƅ�md!�$��Ɛ�sj�4i\�ysC�z!��:<�S Ԣa�q�b��}!��B/��T��m�L�4�)�i	�.k!�dv<-P'���.Ǡ��S�U$-U!�d�LM�A�#�I�\X$kX�z�!��W;{�nR��џt�zQR��K6G!�d��O|.�s"���xċ@g��!�: T�1�fд� ��%a#�!�V�KrĠ<G�TY��7!�b�J�Y�IY _j2�r�j��!�dA&IM�����<RXl2H�<n�!�D*�DP���ݳ����4.�!�� ���W�J3R���a�B�2\����"O�|h��C�4��P��-�4	92"O���W���(�u�@4��YC�"O*d8ň�K�y	���
et�u"OTY���U��tSA���iI���"O�I3�dU#$8�RD�,B5�l��"O� u��h$�L�}2V	f"O2 ��+�ܐ4 �`-��8�"O���G�{�QZ��� $~t��"Ob�`eY6*M�p�΃�t��k�"Ov�`�㝿=�*��4hJ�r�&d"O��;���$�6i�6 �ND4�4"OT�K�-0!�E�E�R�2Ʊ��"OZ}��8g)��A�-�=�ژ9�"O���+P;-0〯ı<e��J"O��P���9.fL\���.4HAq"O�I�W�tJ捈����e�l�;v"OP�q��H<U(pL��J4ւ�a�"O4����q̔&@�F4�""O�i ���2�f���aݳe���"O�9c�MF]Q��F�	����"O�]�5i�~^�S�O׫^8Mh�"O�a��^�X�>X���h ����8�ŞBbx��
�:T�J��)	$ ӌ��h.�`���&:VF���LoaD�ȓ*Wr�Z�#�[�2���K�$n�L��
6������<���yڱ��Y�Lx��2����V�2 f���-��m�g}����R�AE�̅�(8��PU�dl�AC�(T&��ȓST,��N�;��a���J�mӦ͆ȓ���[��1l7��k�D�X݆�L��Q�` ?'*8��FWp�����+����@D?֠����n��ȓ<�����C�AI�Y23b_�RNVA�ȓYJ�)&Dsh 5DEY�a� L�ȓ9�r]���S/J
b�!�	uk`��W�CEc�kc����O�BE��+�؍Ȓ,Y�8~8����T�.��a3,�V�+콐�o�[؂L��,$HA!�Q�Hb`<�ӈI�S"���8�p�����@A�ĺ.� ؄�eV�ѩ��W��ڢiR�A�8���	�b`A�j�q��i�HW0ц�E~�[��I�8X{��K�W¦}�ȓ*��)c�B�9�-���X|��ȓ+�n�2Ȉbzh��B��pՆȓk>tC��s�p�be��tht�ȓ|�бuI����Jf��0c�Ň�|1duC��j9.����W��ȓ&"X��Vj�n^Z��@�G�B��T��F-&��"h�N���)1�
�8���ȓk�l��7�U?P&�8H�^=F�Y��&d&����FX�}Qk6T
�C�I�V���/j�97��24��C䉸b
q�@���G��B Á�)LB�I�.'6�Pc�m��a��O�%C�	!��\iwl�O��B�+||C�I'=~�鳭Θu�E��~�B�	M;U�A7&}X�:F�H�@xC�I1d�.pӱ
G'%�*���%9�4C����4���B>1k�MtB�	g��qk�oC	�(=˔j�@1\B��X�J���ցe!�͢*'�<B�)� V��q�%�8x�(+i!ذa��']��W?����럩*}��b�i��_�C䉄`� p�3#�":�h�������d3��Y
6p�3�C�-2���*�!�d�	W�`ܲ @Ϻ\�� j$o!���)� �j7E�]պM�T��|�!�7=׌�+��Q�N�8��ƀ�z�!�Wh�xK �<w�F41`��6!�$�|��;����EJ5��!�!��9.nr����?Y��Y�C�
�!�đ�=�����ľg�x�!	��X|!�	�r�:���I����{v( c�!�$L3;�%Y��Y5+��X���=�!�
{7څs��P�?������5NT�����	�c��Ԡ!S�$��I�P��<��B�IA��J�D�Y��E�F<4�C�ɽ����>8F�E��FG�}&ܣ=�ç9�̠�w�%V���##�	U���H�>$��ʍ�<��PO�	&��_�сH�_��P�	�x���QP�Pp��R���32l�W�0D�\c���g#�u�/�{�8L���>�'Z�O�O�剤D骱�v�� 24�]�Y��B䉣���ۄ���[�
L��\� b�B��1|Ǽh"�a�?���2��D��.B�0���j�Ǉ�c���[���9v[�B�ɥyՐ�cQB�J���Q�C��rB��b�pK��w��v	�&IlxC䉡�H��eˑ>)��l� @]Vv:C�I�V=R����ؐx�z���$+�@B�ɒ^hl���f�8Q �W��&B�ɪ
1���'�@��j�hǆ�6B�	)$��T@����Ъ�m�h�"Or,�5�/�F �t������"O``D���AB�$�C'�<���R"Or��#N��2�;F 0j�Z-�"O�A���.�R��RN<�*4"O%)�K֤������X�'N�S�"Od��U��7���:�ፃ>�����"OJ}!�)F�����[~p��V"Ot�J8��P@uJ? g܁�p�'nPy�<��"�0|x�lG(ɝk����у�A�<����]KB5�b�Vs�N��� B}����>��`��bl6��S�Ε4���;���o�<��FDsK^���ݘ0ޤ0C��Wf�<i$�K���v�	jS��#\m�<qv�	�	y���w�ƛ!Cz�S��p�<i� B�S]��uL��-��3���p�<Q���?{���Ded`;��h�<�Td@�jl�mC򂎘� �����O�<��;@��D���Γ(�(�z4N`�<s�Cz��
��ؕG ��!�D�$"��8���;C$]��G�e�!���R�E�d�S�3> PuOO3�!�d9��훢n�z72�ӱ-�_!�
g�R����]_0����f�!0�!��#H�x*�N�%�d#�]�x!�$��O��KŎQ/������x>!�D�G�n�k�!�A�)Ƒ�'=!�d��0�p�% �t"@�1ꑦ,!��=�,�U@:P�ԧE!��=}��t��'�p�H֏�I�!�d\g;�e`��4]��݉�W~�!��{2�9���|� (�� 8{�bY��S�? ���5J�>a�$֯V+"�\��p"OP�G-:	P[�#O8Q����&"O��ᚈ(9F�ҧc[^�(��"O���b} H������"O0��	��tO�r�N" i:�C�"OH�K5 	>y&���D6aN�u�"O� ���2+��
E�G�UG^��1"Od�+b	�<UЖiz�gL�50X�rF"O��ӳ�#@h֥P$Y.�hs&"OlO�<���	�%�;z`�I�"OBh���)8�� �JRR��+�"O�r堐��lD���K@��"O��C�\�6�#`�".3E��"O�<��E�Ip<�SDȬm%��""O*9JG��m̈�C�H�}��&"O�-@��[9�it�ʾz	�uQ�"O�I��M̥l��E�g��,� �P"O`��i�1O��#�l#ZѸ��"O*�pjT1pd���d�~���7"O�]�S�6rR�٩U�K��T:�"O*ᒏ��"ulċt�
u`��P"O��o;`��"ǩWx��"O8)��K�b�J��J�(m��!�"Or������z�*�Fi6t�"O�mZ�!˻_=�-+��	c�(�JA"OLc�(�F���SF��% vt@Ye"O�I����A��8AM%B[�� "O��p���"�6��
��\����&"O�\y6��z�6P�P�>P�pT�"OB,�҇
0hI�Uc؀k�t�H"O0Pb��_�ԼRġ��r�BL�3"O�P�@.ڳA��G�M3��A�""O�AAă��L`Bo%	�T8 r"OPВ$ټ&̶d�3��.�R��p"O����l$@Ƞ�^F��H#�"O����ֿa�P��"X7LܼHR"O��c�ުM�2������~�N�0�"O�����ؼi� ���C��F�D%�g"O��a̩X���8�BE6�h3p"O�8�A���%�0��aD��0��q"O����8p�\ �̟7N�yT`7D���D��:�����&$��w�6D��`�.����K�?4^<�
2D�иGf��E��D����a!B�.D�4����
�2(kYF	(=���-D���viH0�<!ѐ�L��Z��N+D�@�*Еzt@�J9�LX2�)D���*H'cЬx#4�C/(B,�E�$D����'̺
v�� �j������C"D�8��ͨvz�
č�* ��i�h5D����?,<&���9#��!@q3D����×,f�p�y�F���	#D����[�L<AH$�@%�!D� �AcH�*�(hˇiĀ:�����:D�TR3'[�"_���T��
s(�	�$D�l��	�/c@�:�B�~a�Y�&D�ؙA��1�p��� p�]�E�!D�PR�+��D��X��=Xth١)?D��:��Ʃa!���%`�S`����=D����ݺ+�q��cB�j!�5D�����h�M�BC��\0�td4D�|(���0c@)���lOȡ�l0D��D��<o�T�Õ�[���A+D�<�t��&\\��Q�9$��d�&D�� ����E�x���;�Aڰ����c"Oݳ���"-YF �$!�&
�l(�"Ohpٓ�7��J%EQ���A3"O�<0��L?,њ4#��S%Ww���"OF����:%�,EzCkׁm� a�u"Or]�A_�Y���+��2i����"O���#-�0B���"#��8V���C"O*����W��D3�٠2h��&"O�%�v�:p���Q�+�]�y�"O0!��#�*Kt ��Y��:p�e"O�٢b͑lc��yw

~��0�V"ON@sG�� X�
W��#�Vdc�"O�)Y"FҰ�;�L�T݄���"O꠲���9pf��똤��XH�"OV9�aţKKF�!A�	���	��"O��a���L�rD�'X�jq�"O���3�.`u�EKăE�x�|A�"O�zv#pg`%80� ����c"O��*��X�"+�=�F&����"Op��6D�Z2r�9���8�½�V"O<P���0bĦ!3�'�>y�"O��p�;z�\{R`�r�R�e"O��+5/�$^�U�g��9-p#a*O���
�W:�@�%�,͎͚�'���ڡ(��F��P�6.ԑG;D���'����r�i��X��lS=DpZ�'���YD
�l�&8��Ǹ7f0<�
�'xĨPWFC,)�I��	6*�*�#
�'d��Æ�pH�ׇ[>$��� �'U���e���p6��H����'���b�̍|��𢦄�h�<�'S�MS���+I��T�F-f����'�z�����uw�ܨ��\d!K�'��!1"Iք_�@!�#e��Y�p�2�' !�3�1�T�COƆ R�q�'�n��t�F#|!�Xbf$G6t<�8��'�<!��Wd�:r�`ݩ����'��8�A��#�ʩq ʃ�u�&qY�'���Y#ā0.�������X�$I9�'�6$0���6~�H�*bвKF��'�@p0��O2�e���8:dŃ�'�L�@��s�6tAh--�bT��'�l� e� �d��`��?��'�Єh�A%R�I0�k��ȕ��'o)���,jE`K������(�'V*���S}W��y�EW'|P��'I>LA)K� b ����ǻo�\!��'Sd�q�_#S����A�7�����'�}��˕�j�m\�D	�	�4"O�2E�*�����R�F�#"O�t�PĂFB>�)WJ�%Aլd��"O��A�_�T��I�#9ú��q"O@�����c'x��ŋZ�`�"O긩u�K�A"j0j@mյo38�"Oj�:�$�0h�Ԫa%�72 �[�"O$��Lۿ1�H Q��m���"O6=�Ũ+b�X�[&��4 �Ѓ�"O�h�J�� @�0an�E�eI�"OB�����]���I4G�U���"O�=!7��*e
(�&%hJ��1�"Ol�I6�ɩc�Le ��>o?�8��"O@�d&w6�2u/��Rݼ{2"O��Gi��jB�R�G�!h�t���"OBi�"HB�]|�D�fԳ}� ��"O� �1`0߮/�X�{�R0y�&A�!"OB��E�]�-G�[6�E}����"O@Lb�)ќ@Y.���[�b�@�"O�(�%�&IT�u��Y��� "OV�T"�!(�����d�PlÁ"O0�r��%� �4![�k�J��"O*48TⓄ\�flJ'���f4ČIt"O�
gkN4:Z�7��B���"O�\��'^�RG �w	̥���{#"O*�AYX�R�K��kh����ݲgY!�N$0�����g:�
��HLM!���*�J(J��U�m��3ӥ��oK!�F�.c 8;pFQh5�gE�J�!�DN���*`��t��A�s@�Zv!�Ā�2V|3�BL�{��y��M\�W`!�Dս%��O��6#E&T/aT!��=w�Ȁu�V  �f��U��>@!��[���#��%a���@�'qO!���A߰Trҏ�f��=����2G!�K�wa��Ӥ�J~���
� C'!�D�2��@��R�e^N�{��l�!�0E֞P�v��Q�(�Pb.�!�=2����M��S�;��_�e�!��i|d�b�ȭ>,H�r��M�!��Q�z��]�'�d=��0ņ�	\!�$ɓdv	P�-N�d�~x�$ĳ!�ĉ)@XB��7�Z�<������Yw�!�$�7!�L���@�[��!م9#{!�ˆ
�h@�"~�r��WC�3w!�D��]�6��hϦ<��+�C]!򤞜yx��`�G�%��8�+� %!���(Z���q ��P}�]���i!� x���Ht�d¥��	�O�!�D�:�x�:uă&]G����H0>�!�#	4�H0�E4!-h�S�xS!�d�4��C��R �h��܎G!�$�u��D��X�__�س�E6!џ(G�$�>\n�iPF��)�Tb2,
���d(�OR����\�L3L)B��S�29<TZ�"O���� �d;��w/A!r���e"O�h�3�ƥ\�6I��+F�y���r"O��ȱ�4ց��kD.s�����ݟxD�l4��|˕��'K�iۢÚ��y��Ň*襃����q3�^�yr/�3gIRY��-�/�x�h"��yb�B�Z\�Ѩ %�"�Z%ѡ�Ϥ�y�H�n� H�(M���!d���ybA.~��@xEG���]! MU��y�D����c' �[]��
j>��O�"~�f�?hI4	�.�'��\I5b�^�<i��C&-P�sJW5'c��NQ�<�B�\)%��M�"b�8B0���O�L�<���/[
^P S��)o���B@�s�{�h��d̜a��+��З�.08.4D�(��N��Kp����H�8i8U�?D��j�G.9�x���?j�H�I��8D�Py��
�.����
9P8H�e1D��I�YRᘑ�ԮhJ���ë1D�L���P>2�t����_2;7r���/D�\rpL�2�xK��R[�R|� )�O(˓��<q�'�tlY�aG�)H@�vJ9��а�'�V<��! ��%�f"�-�D���'O�M���a�8���� �$�	�'�� �f�A>H!6)���gb�U����?�
� ���b����H;d�73���t�'�!��8Z
,ۖ�A�!�4hwk!!��6k&���]� ��W��:��	]��\��*pq�9�k�g}>�#�L8D���3�S�m׮a ��؇2�:ɓ@`4D�$����~mL�)�,I50�1F�>D�l��$�b�R�I+Q\��H��&���O��$� ��H�.Ày�����B�F���O���2�O֡b�L��M+0-�иhc��w"O��X5*K�O{ �[�	;VVX��"O�Bf��T��P��wcڈ� k.D���B�Q�˚����t�>D�8�q�V/?u����X�j��iR
;D�T��j�մ��W��
5Ǟ���9��4�O��`�&_I?��jb�@�u�0Y����d��	f�ޗ|F<�CcmM�%��[�b1D���g)W'(%��捪U����2&.�d�OH˓��S�ɔ�f�θ"ԉ-sD��)"�q!���`\j�1�)�s7�`
c]�Qb!��:�H��È�U5�p!S /!�J�Psq*X�`�4ۀ�àG�����I�|̄m�&Ř.�(2�ТZB��;l���`�����p�#�"�j�*B䉡p��s6E4K��i��Ɩ&���=9ç_s*�D��:14 �U���+�� ��L�TQ�s��V�(��`̇s`��ȓ���Ei�~�� )���6��ȓ��[")�|���м:x-��n�R���?�Ó$v4��@��:l4K�Oȫ\�p��?f���O]��08�ڥw�N��S��B�/�O��9�5�A	9�`���o���	��;'��QևMUf$��_�t����:%�%	7l�\y����@�e�I89�r����~uN��D��M�$�G�
y(���Lb�%�Is����&��8,�Ry�m���T��%D��J� 	+u�.�ؒi��u@xDqr�5D�0��]ڼ�nN�F�>�H7"�OD��<9�����	\�l��_�H0��$+
�B�I�p�t@�cK�W�С�eߓG�C䉍谢4��;V��90c��*Lu��?9����$ �x�*A�z�tĳb	/E���)�' �z�ǃ�-.ZD������<� q��'�=9�P�ue���^9�$ak�'m� �62�l�XU�,���O�����1��DU�&|�� ǯ] b@8�D���!�҉��1�g����Z��{!�d���y��ܮ2B�Cժ��Q�!��'��5 �XA �F�zM!��҅t��QᶂL"$��RG�'�!�� �'�Ru�"iW�~(�葧P�!��P��A���޶H0����'"|"�d&�g?9&J1ey���"փ������]�<I���$�ࠁ�	tN΅�4�D�<���C�8�ѣ�fD�2m�!CD~�<��Ok!2�`䄎|$�Fa�p�<Q��&�@� �&�{.H�w��U�<Q��H��6�rr�a�X�{ebXy�<�����E��|膉^?I*@�{�E@L�<QNQG�4x��ȸ||�T��r�<�qE�tlB��t�*+�����Ke�<��4b�Dqr�C{��}ȲΌc�<9e�0J�hMR��B�f���04�S`�<�ïG!a8�D���]�)в��6�I^�<� j���Dݖ�`�����;2D�������G��N�9pZ�{t�ǼT���{Q��
�y¦کP������^5F�L�	�Gg�y��R/�D�C�EE�)3�/X��y�@S�-��e��@�-)6�%!�;�yB$�)�в @��EX���y�Kޗ����%iT;RA�0"&�y2KEO��)�פ�%y�.q�7����>�*O��Aw�P�Y�,4���޶u��I�3+$D�|Ȓe6�UWcX2s�4x1�dɡ�y�+�S�4`תɔr���k %�4�y�$A�,��j�ꔪ�p|�G*�2�yBE�
I��d	��٣��
�hO������Q;��e	�jl�RS-�f��y��I�K6T��5X�D��U��jձ�h�$D{J?%  �D�y,h̓��]�k��8��3D��CdKP�yO� {�F@�~R9ŀ1D��qЬ�3!d�V'	��Dȉ' 1D� ��jF�C,���%Fi��$���4D�d��dE+${B�q!C�sx\,	��?��7�O�$�V� A����J@�(�X���'�1OV�0��X?)̢� t G&��sp"O�4k�@�t�%Π@�&�³"O2�㖭�7Ed] �"U$m�� "O&�&��5(w�� ��c� ��"OFՀgC2_���� �:aZ���"OD�@Q�&NV
��/�(*��4�'��Oh��Ұi��y&`�P�N�!Ѡ֛?F�}b����'�6.��ŇG��Ӓ�&��#�Sܧ%vQ"�n�(6��0��"6�V��T��9CQk�1l�.ib#�Wb�ꅅȓ]Z\��2Më1���[+pŇ�(�@���H�C�N�Q�!K�-�xU�ȓ�`e�t�Ȼ<�J�� ��#v���ȓ6���$$Ǫ$����EMW}�(��A�@���'�L{lD�BdݕF��ȓTv��Q-'/��,�'oުh����ȓj��NF,��"m�(�,��ȓ)�������;>۰c"�!G��ȓ�H��@�&����I� &���ȓn�dҤ���9����ċ�*PH�ȓ<&4����K�HieE[6&����zs԰b }\]�F2�\	��6�����ϫ ��txW���e���F{R�O�l�>p�0���4��y3�[e�<I��s������&�(p�
LV�<�R��>���b揞1�PQ2t�T�<��9 8~I��eT�>O|�k�"�i�<a��G<N�|��/�6(
p����<9'�C3Th���Aj��N�a�Ew�<1R�A�����sdh`���Nt�<9@-��A���$̪a��鰐��v�<�!d��9w �B�T3�~����Mo�<)��"p�J$ ��6Ze��b��U�<�ab͏R���3�_�d���:�W�<a��6�@�E�N�Mq�鰳c�V�<Q��
�81�]%?��|�F/IU�<��A�p���B3B@�OZ&���LU�<�Ŋ�>=zXJ�X8'f0aAG@�x�<��ǚ,�u@���2n�%��w�<ɥǘ%>+��*�ک"0�p�r�<1&��$�2��$f#.�@�%Tk��L�<a���>L>�!_�cG}P"�4T���GJ �X��-���-6��<�4�.D�� �=P͚)#��4Ð�k�"OzY8��S2'�l����OM��bu"O @&��J�V�I�;О�QG"O$�J"G��p��%���s"Oi�q �7+��7O�Ay���"Oz͚T�D�e�G��Nt���"ON$�D23k�K�Ύ}nB�"O�Y��	�1m�(�`��΂uS���"O�9�q!��0�phĎAu�Ę�"O��'�C)���!�mC���,� "OL$ 4���5yÍ J�dA'"OL��R���^%����j��8S�"O.8��H8�DX�����a�"O�0�c�ύ钀����(�FG"Op��%����#7�n�D"O�1׌Y�Ox	Z����|y��"O��0W�\�z�F!�A�=���g"O�����ܚf��-J���[�"OF�9+ݭy�B�gL�	U��8�T"O�	@�[�|<��*��1���"O�������+Y��cWUy(X#"O�4"�\�4�65����[Y0$3e�'�ў"~�IQJlT���/�	n��F�y2��]<
X�WKN1��5w�Ź�y��	��,�H�JH�u��ac�$�yM�$s:"�		J3g�&��a��#�y�gkG�E�5j
�`��i94aR,�y�d�6`n�8��_�Q�h9#�@��y2�����K$e	-F��5)c�]��?y���4�P����0�d0� `Q%��-�ȓ
0�P�H�a���郃�G'���x�h�yЪέ>����Q+\�T��U�L8�$D@�v.8�+vCϽd����ȓ..�yz�.L�{���K0 ĻV�
�ȓB%�����ET�1��bD
|(e�ȓ:������#KH8A��uX�	@y��'���S�<1G!��^�}buo��Y5v�"��Ur�<��ےr�j��/эhBQ�F�u�<�TA�$A�|Y��2����L�<��dC�Рd3�Z�c��Zӂ�T�<�P#�G�08)�FV4 9v�8�H�R�< %D0$�l��gAI���]yw��g�<Q"lT�9ڂ��4쀩�*|�ߟ|��ԟl�?E�������H{A&U�I7�}��Cѧ��4�Ob�(��_���٣��"��y�)��wEN)6I�D>��ɑ%��y�nL/F�ÍD�C�nh�M����D�OP��0|Ԩ�uR���F�����R�%[�<A�		)Z�J%D�^kv��@Ka�<�]-��	�g�L�Ïxg�	D���JT��9U��|!���'^��q�rJ-D����S����i�3s-n��$�,D�tV�S�k�z�Y�ϟ�g�4�� �5D�d���g~d��*�>F�����4T� Z&̖Q*��Vo	&���$"O�%A �R���!8D��	���"Ol�@V́*��&�Ho�JÙ|"�'&��E�֩?؂�Z�OQ1oC^�a�'�l�S�T����a�_�^?�1�'^n!�«I��	�)�x���OpX�(P�g���V�'?��j��|�|2�I�l����v��<Hn1�4m�9pk:5��0
麰!Ҟk��0@�J5ry�<�ȓ~�գ1�H,.}�Ƨ˳,t�'82^�HE{�π 䰻��I�pU��X��͆wc\$�"OpLYqk'/��p����bXRR"O��3��޳^�ԥ �̃��~)8��'��	<<J/^~c�+e
�K�T�D2��|��$�p�dH���T�������@�!�ưƴ�r�E���@؁$�y2�䕳5E��x�gS�=�lh���y�6ʓ����O��$�d?�` t�6�4m� hr�Ub{�<�`���� ��!�9B�t��0@_�<�pix�)���d<9Kq�J�j!�ć&U�n�"7��Z6��R�^�K!�D[:ߠ̢FoFL*0m�NȮ|I!��ɢ�y���9��vm��G�!��8���4f��oMJ���&��'ў�>-Yg���|S&��k�����1D��2�b4ot�9��"�<Չ֤:D� ���>�)7�W2��k��8D��q͒�S�"%����>J^΀��3��Z����g׼G��uX��	.�fQ;��7D���AEM�3@s� 4�J�rv#D���d#�fDQ��_�V��T;�%=D�T#A
�+B�t�a�	3pě�&/D��jF
��DH��]0�$��i)D�X�rIM40o�h&$�+|��}�)D�<4gs0�䈦c�$1�}z�M'D�����ϙ0\`����b���p0D�����ιl���˶�C�bJ}b�#D�$�uK��/���1U"��4B��G�R��ҎZ�%����8d�lB�1E�$ ��gsʅC���5�(C�.o⠨q�B�|���`w
�(4�B䉧!�|���B^;J��hC�"$��B�ɥ@"�S����0�R\�P�Ф/zB�I�yJ�00aȞ�vt��K�PʰC�	�
��S�H �g@�|�lU� ��C�Ɉ�:Ձ� _�dm8�#�v�C�I�a'��9��Q�/�H)��ιC*TC䉰"*���	^�.�t��2 C��B�ɮx	�� ����l�S�È9>����O����O��D�|R��ܘ'���#�W�!ˮl�Ejи!�t�h�'<�)I+Q�~�Ib(��T���'?~�i�JC>������.1�
�'^8ؒ�B�|��ؚ"	�N�N�	�'�h#���DRu�R��B�pdp�'�xX�d@660��>�B\��'�(�1�lY�R�̤���G6Kd40P���?Q���?	���	�O\b�|�7�׶[T��P5_�ᒅ�-D�<�O�=B��`��
�E<���bo+D���F��%X� ���މ�Ip��*D���aZ���8A���'=�8X[uD&D����ƞ=$qP[1PH��H��yr�F>xb+S�����f��y�a�{c����0�����?���?1���?9*���� �ɿ JT��s�Q92ݒ�:�?erB��)䕂��Ɲkj(����TB�Iz�dxC��#l4�E@5cG�C䉒�xJ����?�b�ˁ��Z��C䉜[`��Ӈ��-Y�N��b#C�C��g���sW����xb��dC��3G�����@�Z��P�1�5M��B�I�M�8�jg��T�.��3��#�6C䉎U_J��`Y�`�!�U5JL�B�I�hǾ��5o�$�dz�E�2NzC�ɿX�U3�G�0����F�Mg�B�)� |)�����#B��(���"O�����Y���c�5.��A2"OPL
0��4=��"�)u�@�"OT�! A�<�D��~�Ci��yB"B�8 �V�Y��¨����y��	�� ��Rl���B-�y��LUy��{���g��b��y�gYz������~ "�����yf�-e�@�����)̍;�yb�D�y76h�a&�M�&�A�Б���0>a���SSh�{�aԑd�*�3%H�<a4!QmF$a���1n�s憗|�<��FŴWS����*s���Ũ�M�<9�.�"^�b���)qJ�����`�<�'[0!=��j��R�u��P�p�<y��M�L�t��vL_��4h:��l�<��]�k�x8B.�*u"D�hBh�<YV��y4�x��33���_�<�dPepU:�g�hŠd`կ�[�'.?-��\!��0�@��Fs�B�	bx���3ڵ^�F	AF�a��B�I�F��e�E`ƫlP}#hB�vB�	}#D)����g-N���LAxdB�ɤY��ej#Ɂ�)C*u1��_�4B�I� ��#��DN~�24��J�LB�I�Vú��#� e��=Q�B��Җ�kn߫%�G)�~�B�*��`fw�\�����B�	��xU(�,G�����ؠ `�B�I�T=>��v�L2E#D ђ�dK�B�	�@1đ�T�i&��Z1�H��B�I@
��A�F�b�%Y��s�VB�In��@a�=|���)�+�3(B��Q�J|Z0!@"�����Q��C�I9z-8��@B�,zy���(1�C�	�YE�����O�B����d����C�I$��5A#�@�HXt��/k�C�ɒEhL�b�W�$;"��$cA�MiRC�Ɂ{6V$�5�('%�-��QAC�I9^���{d䞤��q0�+H�	��B䉖AmIi �î'e��S"ى$J�B�Ɍw,"����-�nl N��`۔�4���$#������ǋXb�Ra�mu.B�ɌUS����Ѓ+����#J�B�I�T��)�������������$'�S�O|���]�LҒ��b
R;{���t"Ov�@/C����C��#�NP�f"O�S�O��Q@"-B�˂�.�8x�"O6���4A�]�-��p����"O�9� �+U@���k#]X�a�"Od��7�ڂ%AV���*��Y���[w"ONyȦ��",K�H#<�(W"O���hX�"OܕqDh몤I�"O�4�Bo�!<@�DǍ�n`�"O\ۗ#�?@�����M7�ܨ["OFɛ�bO�\u�X p�]-c~Ȩc0"O���b�Ź}.luE�Ow�*�"Oz �E
@�F0�⣋8H���"O���f��/)w6MBw�ǘL�\�V���<y��I�=u��)� ��//z-
'c$
{�Ofk�	!&-�I�� ݴ�ux�"ON�U�޺n�Z@� /��z���"O��5��CT��ۏr ��d"Ox�i�����R���R�Ng6 K�"O� ֠0�NLt��(��MnD|-r�"O\�"D)F�G-f��$�U�gs�����|��'="�|�|�#��G�(�0�ƽB�l��t�M�yp!����qz��/����m�"j!��7+����EaF"N(ށ(b-��!��AvNt���XJ�
E�%.ͩ5�!򄀌v���I�DV)K��ԧ��.#!��"b���kuo�C�܅K5!�K�~�*�q@�Y��)�3�_)�O��D,O�K1$� @J�gGO1O(	i�"O\Њ��57rS���Z���"O��P����S-����BQ�m���Y5"Oʔ�P����BDh�jQ0Jڶ�`�"O���ݾ?�(%[����k���Q�"Oz�rA�ʕ#A��������6"O8)!Tgm���6,��}�ŗ|2�|�R�t�|�#k��Vā��
P윒T �]�<I6��),��uH-/����bGZ�<�!�53h�jp��4iLd���(A�<���k�h�s�ԥ.=��A�<�G�П|��5��gȟ5֔x��e�<	F���0��g.����)@C�d�<���I�6����@�(��Ѐ�j�	{���	�O�zfK�Z�H�C�J#Oܠ����4D�(�2�]��V��2�$I�aa��y%�\0@BE+��)��(K$�y2���z��
��]���Y�u�F��y�"���ؓ�(ÑO��͠$H%�y�]�\m!i�Q�"��+�1�y�+$Bj�*�^%�1�F�y�m	+6.� S�Z�4�"������y2�On����".X��*UN�<�y��¤qK��`@���y���<%�̪1d�wl,A���yb#]�J��bb�	Ԧ�@$��$�y�W�WK��"��՛2��pbk�=�y�� ���Å/K�]^����O��y��1M� �fB�d��x���yr`#~��dт�ށE�p�dI��yB��,<��i�O����?�y�v��E�?G�|ذ�����y��[=$�:�9B���}����+�yr��>@읓SC5q�Չ%ʌ��ym�#��ˡ�nBh�{E��yW JQf�{���-U�(iSe����ybf
�j��0V�a�P�Q�fG!�ybIA�|��ȑ�Q�,����]��y.�1%@�AS�ӥu�ąxb��y�Zq�t��IV�p��(1%\�y"d��m��(�FѵjJ�e��ʓ�hO���i�wi����2�H(�5CܢuW!�d6[��r�+	�*�)��1)!�d �m�j@z��i��pJw
ݚ$�!�䚗G�ICʌ�D�K@�A�!�D9iJ�p6o*[���`a�,!�$D�(����u��(a�	>�!�����4�*����c�Iߏ/�!�$���g�?l�zǢ��*��O���r,��g�"�ʂ���n$ ĪQ�&D�,2qG6*$ `d�*k�6졂`1D��� ��d;֌aQ��c�N��0D��Y��Y'nD��A�B�=2�.D�����C�L @���mz����H'D�҆�ڂi�P���('c8��F@2����� 0�h7�L 3���	".��{�*x�U"O ,+�	O�Zo���c�Y�(�z�J�"O�1��I�J�s��#�u"v"O����Q
SF�����I:0�,R�"O<u�dGB"]�:ݘ�f�)�h-1$"O������lh�%�J�� �0"O	�ؖ=_�>Ͳ��5��r�"O��H�-�
h�A������;f"O��{�
J�@U�Y�u�1S����"O��$��%%p�;k_0�❐�"O��Ϟ�7^ �"��į;��X�"O\1A�?� r� !�\c�"OBi�ѫ��22���&Z�q"O�@��&	����+�x�d�[V"O`����ǸN�`��3�A=�<�g"O�iw�\3c6 uk��
�h��l:�_��F{�򩚟4�(�F˃�*FE�@�X1;�!�D��3����E=y�&u��㔯/�!� U<J�b��G�?��IPPb��4O!��ld�c�Hȥ5����o�B�!�D��N���	&,�(����-�� �!������C��)z*!��K�-'a�Ip��x��Ɣ'u� (	q�~n� ��'D�P��	
�~�a@�̙tJ��c �)D��٤#�9?n�R�K-�v�`"2D��x�I���$D�RM�� *2��B�=D����*�7�P�Svp�9wD=D�0�U���.��F��?`}N�H�	=D�4�7��/vNȘshO',0y��'�b���T���ǭN�lX@AM
��O���� ZHȈabi�h�����!�X,C�VdR��toXQ�9\�!�A{��LR(	�bH�`6��U�!����&hѶ#�nĤe>�!�䓅�,Y�%�k$=���$	!��-q�xu�L)h��IX3�G!j�"�)�'w 2�k���LWj%"4��10Q��'�~����1�mht/H�V�r�j�'��y�CѾ;�����N�!C���d�?I����&�ǮM$�8R�H��W�!��U�A�J,���h�4�!��Y�%W��P1��:5�(��&�ɨ�!�
?�D4��ÀwԢ���K��$}!�W���85e?_��`BA��g!�ܻ$p�!��Mº��
Y!�d2�)bEa��_�8���N^Lh!�$�/vT�$Ó}=��C��d[!�Ē�/���9d�ȧQ�b,7,�F!�ʿ*B����ݯ˾IcTM	4!��L�+Bn�8%�(�&0�왶G!�d�|{�0�J�]�J'!��SS!�Ҁ< �e��'?�u�  	�s�!�d��Cx`�r�L�~$��xuH�B�!��*4 �٤�I�<:Z!���b!��Q�v^̘�gEP�aS�a4V�u�!�dR>�:)��V�W4Li�!�E�!���)[��S�N #�*��/�ў�Er*�)h�tá�ڍn4����i(�ў���I�2��D(�DؕM0 တ-"�C�I�s!$I�'�1fF�eb3k�5��C�	�(��U�%��`V.�)$B�B��!) �g�XV�`�y�fB�I�-`R��R�H>MD��
2\edB�ɡ��(c����|}2!��
6���'�	m��ߟ��O�� ��Sc�Ss���W���~hH�d7LO����Z=%"�p�ю�2
���+�"OҰ�OΊ��s�#]eH�#�"O��  ��s� \;��ٺ	H@	��"Oa�V�h*EHR��6B�8�A"OA�Fㇰ%�.U@�(W�`��"O��[D��4#��ZA��Ne�$ۀV�|�I�l�'�ўЁ����bb��m��i��[��E�yb.H�xz�T�,L2���%���y�`��w쀱�)Ђ� �B��y�(]��m��kɏg^�9����yB+�7���P��e��� �I�y�W2~���X�o�[�����yC�;���eG�Ya�L���@	�y��1,�e��(4<�����ԙ�y"#�%
쨬؃	Y�
��� �È�yr�_ e"D0x��ͯ.,mp�ܳ�y���C����5'��&�&�y"%S= ��P[ �ؓlu�t�g�yr�V�[x��i�h��Z�Ŋ��y�䑧.Gl��Ն�5g���FG˾�yB0
y3��Z.X�
9F�y"��D�Ń%͓�O�8�#F�E��y"�% �bR�U�XN��E ��y�g
k�v���N��z�aF!ƶ�y��A5lú�����E&p���E8�y�o2���s�g�9yx�B�bN;�y��J�2�[�	���kӀװ�yBOW�HO�0�t$T#lX�����@�y��҄tCޥQ�Ĥ�vi����<�y�*��D�Y�ga�%�bd�%H:�yR��3\����'��`e�%�!�ݘ�y���V�yt�[�.b��|c�'U�		��Љ*��Es0j@�=�ڵ��'�8�D��[B�
� X���Z�'��P���:�h��W̜�
 ��:�'*b�K`�݌/������}�I �',��I0NmН�"���u�����'G�������u�+��p�)�'�~|���A�4c����cŲ	��'ܾ��0���dm�\l����'<Иe��\���ħD�^�ٙ	�'ٴPҲ�F�h9�	���.E�X��'�T�a낉|�z5��ŏ�=��H�'b���"�32O��a3�K84jԸ�'�D�s�A�]E&� v��.�L��
�'�.)��'�'�D�`��/+p��'Td���e</
8 H�l�B@���ȓ2D�xT>'"�<��������ȓѸm:"�P!/-�( ���Z����v�.\0-w��%'�'�Z�ȓ%[����U8���0F�tP����1j`��!�|�NP���ԧe�d�ȓh��E�5�V@u��s��-��RR�M�2-�x��|𲠐.H���y�`+(�p��� S��ͅȓ9���ue:ghV8c5�F�v�0���q�$8�Ug��M�[�a݊�$�ȓs������6c��Jj�=c0
!�ȓ��Qk�#T�z�bG�_�%��@�ȓB�(�`��X�N!V1"��G41N)��aK@U�� "H *]�����'D�\���dS\m��N�G��@�68D��&��$h)Rᙐ`@3�2#��6D�� ����mŴs$���Z4_��`�"O���aI�13f�;��Y����ʦ"O�ٻ��
k�ڵٷ*�0)J���"Od4�\(J��R�ˍ'?^`�V"O|���LP��|%C�2M���8�"O@aj��T8�}h�K�`M��"O�mz`�X��j����$7 ����"O��áb��:�[u�D(d
�K�"O����\���Q�G�.]߈\{�"OL�9b&�%:H�Qp���k�4�`Q"OXe����m��2ͅF��H	�"O|iҢ��sJ��P���q�ܭc"OV�JR��{*�ii�	�+d�����"O���sJC��N8�vhT��ۡ"O����� �1YF��C)���L˳"O⥺siT�G2�9��Y���U"O��BC��f�JlҶ��'C�$�D"O�����[|lys��*���&"OU��	Q':��r$� �����"OB�����#�*�� d�%�H� �"O��hE��47]�ĩ�ɆE�qE"O�l2��gq�Mb�L�b"^���"O^���
��q}��R�)k��9G"O8y�_�`�9���J!+X�Uu*O`��NތqX�1�ƇK:J(���'Dby���m�r�B�HĎ0$����'��x)�!U��Ѭ�%6(��'E8��G���(���$����Q��'�L-pDKZ��[Azj��k�'�������:�as��p�0k�'7|q��q$6M�ǯ�dJ�z�'.�L�C/Y�+#� +��� k�&��	�'���z�K�$�@�0�)ػg�f�`	�'��l@A#)���4c "\��'�d�� ��1Xolģ�F�W�64��'��(�a�"d��Egk�#:�Lh�'�
�X�&��i[��֥':f����'��� �R6wP��V�K�+��'9|���®��q+�#(	<x��'��A	G%�޸�y K�m��	�'�V4�N����[�+Or���	�'D��$N�;a9Ԭ�@$����b	�'��x�O�$[4E
�K�a�P 	�'Dr�i��"{l��������'��SтG�f���UV�*�p�'�]����� {���>�z�Q�'��`0��[!��}�Ňӟ1[Ԅ0�'��$��	�}�Pѳ���0G�Q��'�>�C`kK�.��S�O)��l 
�'F0���R�p��s���F ��	�'�i3���y���(�HD��p���'$���.��"�b��3�3:�4�r�'��M
�^�i�i��
��;.� J�'ۂ���`Y<M!Z���`�0L��	�'��a��EX/RT����s� �Z
�'���Ŭ�-?5JIp��ϸw���J
�'����bF��j�K�'H:sa�	�'T����6H�L�%+��v/��
�'��c�A�9�IB� �%6���	�'���8 �	~pL��
����Z
�'3ܠ)ѫU�F��1QC,�cth��'{:��r�J.[Vܡ��LS.f\a	�'I���Q�~�>5��F�+���
�'=>��t�ߘe�|a�2D����U���� ����iJ=�b�S�DD�N)�l��"OމaB'T"A:�Y�b��F��[�"O �t�x��-rQBφ*>� "On���C�7��Qu8{"D Ñ"O$���5 ��)��
�Cs�� "Oh8óF�6݉�B��:8h1�"O��S��N&j�3���>��d"O���%��*-�<�����Ck:|��"ONq���
�(�V}�AoT�8f&� �"OD�y����eF�I�c��#"`��"O��mҲf`X|X��O�n6���"O��4jD#'/:�t���9�8+�"O*�*d�ѧ5�`�h��I�Y����"O:�3��X
�
� �����"O��x2E��<�vI�uhބt1�� �"On9U��E6\`�S͜4V�CU"O���2��_I��Ct뎔`&�q7"O���AɝJ]���j�<L
�,w"O����H�"��xP��>*���"O�鳓JȄcޤ|2��l
�1Ӳ"O�)K��E�W �=bчL<�<�K�"Ot��ҁO�#q���U�@�jS4�r"O��i4��y/��h��">d��7"O^q�)�n��IaA��0�m��"O��!�)Ik+H����S�VW���*O�����M5j�`���+�Y��'o~Ee�)��I"}�Q��'��а`.g�F�#��j<��
�'�V@\5.�����	�@�� :
�'7`�H�d�Y�a�@�a*�d�
�'6. �c�ڧ �e�e$��\I����'d(�:1�S=y6J�&g^�`)��'���<p��K���>_�a��'�Px;@˜�gENL�Sǌ;�v@P�'�^��D_T�2A!�%/(��j�'|L1b[��z�tjR�&H��A�'/�S�O�b̔� ���)-���
�'�BQ�#Ħ;���b��J(tb�iK�'�й�e�/~�F����K�q�$3�'�~)0U�<���a�8Y�����'� �����KL��g�D�M�,�y�'���`c+ӓA��1w
ֺy����'B��S�ɬ־��V�T�r�J�A�'7r��թ�-@���ؿe>�x�'�4����O�8Й�#٤�F=�'[�鰂�;�B��n\#J�D��'�� 5
�U���S3�C4~����'h�p����B!*M0��X+@r�z�'����v��)�6QYE�'ER�Pa�'G�;���h�����#ɧ>�r���']�xx0��3.E��""ҵ!HJ��'��C9�h`[d�@��]��'&(c'!��2y�ݢC�Q��>E�'�f���铵
�������=Y�'�.W&U��0qb��|���'ET��,t`.+��7�Z�!�'4
�
h�5Q,J9�!��z��i[�'�m;�L8Y��<q��E 1B�',� J�f (4͐�Bb%��%���'�4t�b�ˏ:䡃닎,� ���'���ˏ/��$�5�m��'�y���8Z~���� 9|�r�'�$ܚ����z��Й1	{�4i��'e"X�e#GY�(��j�/$�j����� ���q�:aXJE��B-n%�g"O������@���kF�*�0:�"O���
�#
��`�l�%v�y"O�0Z�@�5��MٲꚒ	xt���"O�Yp��Ys���h$��i�"O(e�c.:��ʄ�r
Q���(D�����(93.�E�ڨx"#4D�`����9hx��/A�Z^��H�3D�`i�aQ4eY2�3�j�St���u�=D���Z�N:Ѐ.u����h=D��p�"=�
�s�K���t$zC�<D��+���ab��)�~0�c=D��	���q�h(��N7�~�8�f<D�� �b���.�h��C�Ƥ1�C�=D���rO�d��!V��V�8��c�<D��{�K2ŀ���O.��%&D�؀Qf��!S�p�a�$3��*PE(D�X�E�E]ھ*󫐞!3���@:D�P����z=0��̆+8��w(<D�� �`.ݶ�J�+��a��ks)$D�X��X�w09�֝>ڠ�N&D�,[Qj��1�J�+3��k۬�ʒ�9}�1�S��bB�Ȁ�
)KRI�j�\0��ȓ6�Q�U�
!;-l n-cH��=�6�1LO�3F^�t�d`0eV��tm�#O�l���F�:���Y�G��y� L�$4�S�'e�@8�-Ҿ2�Ҙ:�hʕ=|�-�ȓ~�$�3�F�6]'h�S�Maٜ��V����!�R��G��y�yr�i�'��{y2�NHJ��/J*9��8����<���I�@n�Y�FoӅ=G������,q5H�=Q
Ón��x��[�X�&)@�|��m$��E{���CZC�N���*r�X���
��B�	\�����鐝8/2LS��8�Zc��C�<,O��c�]m"���x\.8 6"O�zta�j�dt*OP[�L�@���'��y�lāp*��6O�U�(A�Q���=��y�KH&�~��UP J$xq�X�Cў4o�H�'�yò��*n؅r�II6	�qjv��,�S�)Ŕ�ấ"B4Jx<����=�d6�O�P@�B8�,��+A�.ڎ�"O�	u�_8O��H2�*���9O����ْX}�����C�h��G����I`̓7��V�X��?;r�Z�'t�e�Z�����&|O~��y��vH
�!���?\ܦ�˖�Ԉ�~��IY�O�Z�ٲ턊@��u�ؕUgP-�yR��Q���O.rHSʔ�J�P����F6Nݘ+O��$��l�O*#<��
�3��U�*�+z}<i�tIrX�Ll#a�7��*w�ip�0%p"5�"�λN|C䉖G���A�kڹ(�AHu�̾Iǰ���I�I���x4��.��#|�S�ʬ�I�Ưw0]ѕ`@x�<AF��3�Pљ0o�_D"	wLt�<�կ� T�q��]"	���a��l�< ��}.4zV�Ȝ7�����BR�<�#�
|����.I�tl�t��WP�<Q�W�ik��U�ԅ.���ҵ��I�<�4@�w��1��zPh�!�XB<���3O��;��0�愓5�!%�TD��N������s�Z���;cTd���H�'��@��(�
`��� �=7:laB�'����B-�PX �CRoާ!�z�	�'�� �©:����U��F���' ��jRlՖ���'�\k�u�'�Jtp��:9|���E���
X[��� Da1���i�V�i�("~Oj� �'��'�Z�K��ہ����Ɨ�r��b��hO���%X	3x�E�2'���*E�t"O��[#oQ�����&Ŧ�@s6"OT5	���X%^E���.������x��'����a� �fR�N�h�9�I<ϓE~�E&k��������F�D�3�RH!�H�]Ep\P�`L�B����R�S������� �~�A��!��5#��_�3��z����9�DIț� ��ؐV���jp�$#�S�O�=��X#Ǩ�RF�1�4<)�'�Ԥ�� Ș`�B����)r䲊��!�S��E�#�XӳE�"� E�Al���y��2t&Z���dq�a���'���2�Ol�QhB!6��B�`�*���b���!�d?>�U����]#(	5К!az2G��v�'d h�g$V�E��!��U�$�3D�D�`ab��ؚ���.�L��&�,�Iɟ\�?�|��M��@&�˩|��0*�f�R��%��Ё�̳6"�����l�옐O'�IT؞������Sv��Ќ�6�Ƒ��?�hO��`�Fl�fI��^^�B�,��G<8@�"O��.td��͋�:HI�m��W�!��>0�f�(mΕP�2ti���q�!�4,mJ�a�δ�:��(р�!�?����e�-<����V�I�!�$)t��D	� ��|�&,�1T�D�=E��'���3��,8gf٥�4Fn��
�'L^ �R`H0q�Ȍ��܁;�*t	�'#���' � �X8�E/X�\(�����$�:3NQ�)�!�f����B�d��'}ў"}�����x>z=	')�^0bbXc�<�e�خe-X=� S?�TX� ��a�<����5� 3U�S>**49�^؟8��'@��)?�̜�g�Ҝ���S�'�X�xf�\���v�4m��u���(O��Y��I�7r!h��R�z�,��-��{�$��W <�p AL �J[v�C�B��	P���O��d��A�����߾Z�=��J�0@O!�D-k�d�#A�E���! Y� �!�49��)� �;
 	�C���!�D��hR0buK�@���M�*:!��ٺd[6H �$WHA�M��-�f5!�D�b�(��ϝK!V���,�<!�䝘J��1�Q#؁�.%ax��>��OD�ɱ ɡ)�	��
5��	�ʬ>���S�&���2���|-�ȈР�9��"=��ĵ����ÃJ���T'`	�����*D�Ĉ��V29at��|�8����2?a	�y��T����&"�����.Z�9�q��M�G�
9y�Ha�
[�\1�-+�+IH�'4Q?!෨��,�ĝ��J��l:� #D�`�RΚ�RmZ����	���$`�>D��5��13JbD-&(Р�ێ�(O��'���?�s��H��q �$@>r��٣b�H�<y�\v6Y�h�W�	�5
�9����ȓ8�bS@kʻ�l	ځΞ3 [@�F��~K�X�7/��)K�Lң=��x�,� ���[+t% ��z�(`�'��	G�)ʧI�yF�ɞ�Xe������p@ ���O&���@˧M_�����L�Y��T�t�|"^����/l�m�pl��l8�80�BY")N�I[���Ȇ/N�7~ �@vmZ�,���8�A��y��WF?�Ĭ&��b�'B�xE-Ý���r2�׈O����C�)� ���#D?+����a
�C=��]�4���/
h��馮��~̀��&�f�C��\,�g/��)3f�� M�( ��б�ET���Y��0͒C��/�T8�dn D� �"cyb���X����ɥB=D�țSF��r���{�O�:�3��;��;Q�b>Y�+%UP� k�
Ң=�L � �:�OD�I�<���R�+������Qg��Îxy"�'�A
g&(�)�qA�8Y�xx�'y���&��A�$�0�B+�4���O*�Q �玑�nJ"tT�i��'�qOv�0�P�\^Ug�Ap:(a��"O�탢+c��rs���m(j�x!"Ov5��+c���WlW�-%&�{"O
,j'@�y���1I��@6�D"O���� S���JE.�1 �"O���ҎU�W�:h�PlP�*ErQ�"O�h�s�M�9�@;��D&��p�"O�y���P�A����N#Zĭ3�"O�]�s�?Nt���G�k���R"Oj��#o�
�6]ˡ½Q�x�p�"O$�����ga�A	��.{�P8iC"O�"��H7N�!h3E��"���"O��P�J�%U>]�� �٩q"O<,�M�&JT�Zg�X4I�ZQ��"O�DI���tmB��ţ�ut�$�"OX��C�T�^����bΰ\ZA�#"O&р�/ضk�E2cBG*C���"O���E��a&��G� :g�n;�"O�![�ƙM������j����"OP�zF��e�丐7�
���1"O��QW�ǑD�9�M��$���"O � ��B9�&�r0JK�@�4��C"O,qk0뜏c�Z]����$pvf)�"O���F��N���0o���"O||r!�;�a����=i
�"O�@�$+MR�H�Ɨ=�ZQ�"O�$;Sa
b�NE[Ə�es�"Of�3��SdM�����#o�N��"O��D��^�Fe+�V�A��I#6"Oj�Jq�h���v(�);�b���"O֑2���#u�e�$�V���a"O������@�PRp��7s�H��"O� �a�>s�m����,g� ���"O>�H\��w&��z)&���"OD�x`�w���!�D�J�4R�"OPu��n�-E����G$�;�t�Hs"O8�y��T�cK��������"O�ᓡˀ2�
���ˆ�&�r�1�"OI��SM�`�pƬ�<����p"O6�hu�ƭ(�x]���԰rޖ(��"O̼c���8K�0�ѿ%�"$��"O&���O͒o� �åGA/D�j�%"Ov�2�
��^U�aR3a���X�"O�ɠe_	Rn�Hԭ�zє��"O:u˖b�`^�P�攟\,��0O�|sЊbfPű!S�X$I�f�[7�+���$O�B )�
����C�	8��A�e��k���
0��,RGC�	 >J\���ȇm����6�tU�B�	rdV\�b�	�A�<�b�*(r�B�5kE�왂�,i��q�t�LpR�C�	�l�${������uW�N��C���I�"�#�́��Ƒ*i!�Z����Y�T�d�W#�W!�� *���G��"� �R)�K�j�"O�T	�G�GLزDG�	���U"Oxh��@�+#�J-p�D6;����"O�Tr��C;e����Ck@��ƥ"%"O�tٵΖ�I���kޅs�����"O�@�fO
~PB@"̔�XƦ�S"O��
���<������:�h�B�"OL�
����MR �(L&�%X"O���2��a�m��s**�{�"OX)���u�6����>A�8�sB"O���b^��@}Y0��mp���"O�=Y6�@�Q���H���x0�a"ON0��n�0*ݲ�A�HԵt6]xU"O6܀�J��j<UYp�Ҕ����"O4���_�{� @�A�F�tƺ���"O�8��N��ʁ"�s�P ��"O:�&�L5RN�i�ք4j��0�"O�A�U۰6�X\�q�O�"_��@"O!g҇d�x+���9?RHy�"Or����<8-b� ��W#+D�{�"O�$�v%�7!�*U��9,4��"O�`��ОZ���x@��Hڌ�H�"O<��U�V\j1�߄^�lܩ�"O
y*�J��7(4yC헓s�V�j�"OZe�W��Ddy�-�<c��%��"O�<�F��z�+ʲxV��9P*[r�<Q0��$�f�2��[�^�F$y�F�w�<�P�K�MH� ���l,�͘�)o�<���֝|��0�*���\�)P�<S�S�0=����M_�T�B��i�<q���{tȤ�&P+-�����_�<�������րQ�T�e�/B~�<kP�yLy��A�-���B��R�<�v�;&�Rx��,�6�y�E�<iGk�.�D�A'�ޮ2u�e����C�<�c��Mtnh����Q��PVDx�<Q0A"�TQF�'���&��y�<yФ�����!��S^�(&
r�<Y�̂�Lκ�z�ˌ�O.Q��BNp�<	�A��[
��1#�V"�Ho�<�s�S����*
=:�d�S�N�e8�lrRjè)��&����B k����o�!MЎ��Ԉ7D� Q���B4�{��S�F��d�6?!�,�&|8�ʳ�4}��	�9E鰸����4@s�5�U�ؿX�!�d�2gDvi:k��[rZe0�&5P�9cVT��y�Ĺ��\%?�L#��րO��J�/̰	�c4o(�O�\�ד�,e:b��]h���	{oJ�p�S� "^��āZ>(ȋu��_r���L:R|џ��Po�hSd���O�p�����:��H�!m�A1�EB&gQ��yR��=�6U���90��pak����ď:|�� 6B/z����銳r8���BB�7{V	��J%!P!�ɵ�8�����7j2�(G)�?d�@�PX�����j��%?�H"@eR�xY�ӧCH2����+�O�X�%�`2�,�EQ% D��"�V�_���Q�#� zU��$QZ����bJ�5����'t(џ��K�n�@jKc��B�H�@!�F:[��2���yb���@M(��/�4=�y��HS���d߄k.1� I&��)�'g�ȵ��nl�I@��p���"ڠ����s���і���D��0�|�����@��}&��{�I���<�Kr%��4�1��4D�X�]%�x$)3���IaB�&�p?1�I�Z7��A�ͦQ�\�1 K��ZM��$D�0r�c�;?#��B��-J?P���.?�F�p8[��5��O�6�3�$N�J� ���˟8N\-���� Vy��;^C����ܳ(��*��'�d��Ed�X��9�O?r��ǐh�cAm�=�X5��AF�<Q��]�<#�+��Y���	@}��^��2&Xϰ<����8~iic��.�4<kp*�A8�xàl�Q
4M�V���"d�_H��0	�����ē�Ԩ���zyp�����>}Gy�iS��������.x{��LՐG�Uf���¥BJ68r��
�"O"��fȷ]� )�k�(:{��R![g�L�E���w�|������ P�җ�G�����b�ʽ�y�D(Y��(y�"
�ͦɚr���~r�	
]��8�MW�Iay����qQ~�9��O�mR�S�K֘�p>Y���-_o��D�\�"��uv�Y�/��p� 
�'�R�Q.�3�nhV�)wP%���DU��F�Q���2�fd2f�0�i5�
d)&k�E�(�Q�gB��!�"�l�a�_#z�d!�CvsXM�pB	�a�!�'��56pp7��OZDɗf��E��9��&3z,�a��"O���`i
����p���$$��Q-ڨ��&��&a�;6��g�'[��!N/�<��j��@��1�B��!�E���-a�+ȸaǞ��bl��q�x�U��a���� ��p�LK��b�ܵg�>�=�@Κ�G �ɒ3Vf ���q��	0&=�"�!��,�B� A��?\�����0'>��P�.��<�g�r��'j��D�f ��zQ&L�Q�٢y��ҧ�O��=��ڧr�J}��J��W��5Ӊ�䟃�m
�,Ԧ�Pr͟��څ�^vܠ�5�5��;�
)^{��k7�a��&�3��|�-;P����@���Z�6�Y2����D,CM���A�=�'��I�	����Q�J;�i�tĄ'V��X�L;��>�v��'�vT�	ŜxyM�1�h-s��H�Xܡ�g4 ��O9�T�D���:��ذ�O�I�⬒
B<]ё@ƼRZ��0���T�'1⟔ڒ$� ~�*I1v$�uaI��q�ッ۳sO¼i0E9�Q���284��d,}��C"v�Q��g?a��٨�Da6*9�{$�1�����:��)S%oF%B��;D(�h�[K?6�yA.AۄQ8D�H���/�!È�L�x�D^wѶ����@��a�ȗ'?F�	�-eʼSdJЛE�vu�c�rְb?��C�wh|��$�S"p�Z�H{�>GFVK�8�=����;��`���g2Z��pr��%z�}��1{|�,����#���1b�Zu��&��t4��'�����4J��<�r+O� 0
]r\�tiqO(�Z�n�;��O�����.�!l�`��g ����IJbώ���@�����ɝLl�{�LH*��)��tJn��Ӆ}���R�T>�q��&�	��k�cT�(���[HOa����9��p����F�<���1m�(�%O�z��O �u�3?)�g](z��S@g�	=AXZ�o����o'� �9������5-Ht��I���N9;&�-{�`	K($�G��/4�N��C�\�V
4����=uq��É�#�̱�i.<�J��G�>��
�!L�>��њ#^?}Dybk��U�x�C	M)�q�e��İ>	�j��|���[)��EP%®\�4�e�X�nr���B.��P$��r�>�p%%K�ȝk���:-\dqG{��2*Ri���v�!��.�W�4��10�*e.B�jzR�*�
�p�<�ē�a%�Q
�t����1�L��
v����׫I+vĨ��i�8dV�ɱ�(\����#$�Ir���� ��B�	wº��%'�0�#�8���Qg��t���O?d~�K��uǰ���|��k޵���+Qm�l#�ɀn�x
e�4�O>�*g*ݬR�6l��%	��ə�/�h��p��X��A���ݝh1�D��R<�j��R�v���<)���:H�pH`̐�KxHԂ��g�'�H�����D�Š��m���˙
�~ �.Ƞ�ZH��)��(���PJ��$�!m�߈O:#4�1Љ��Y�:�����P��4h�Z�� C&|F�Ð|r�C$xL� �(qe��ȳ���>�H��F��|� ء׭Ed�'���C2O4)>yCgˏh�{fG^�B���e����	� ��Q��&j��\�a��m"�Z�8��\��H��;oj�qyW�
7|�7���/x�@��M���)�'��d�G�DF�a����d����e8d�;��LC�P1�	�]	��9F�FD��g�dEM��+fe#ZFč�AP��1)�����Q!l.��7��U�6(ׄ�e�'�~�
u�`�\��уU9e'NI@�DG�U�`Q6�D(7H�sV�	3�0�bc+wg$�E�G����"�2���I��3p�2�#L0zǬ�p�i�;���*����3F��O�\��T՘8bQRw·/�(�bN�&A� $` 2ғ�&�[�q��?�J1'ؿw>*�!6C�'��Iy����B �>u; �1&Cҧ��QI�R)w��C�3O mj����Q$ט�a�Vđ�*^��)S!ʌ�/�Z�r���y���<S��� M��'{�^�
SK*�:�c���-��� #k��偔�^Ohe!��WP�Z���Mp?qb���m�,����̭��>� �!1� (!ۦ%9��FJ���\� �Fm�*z8�\��H_c�x@�i؞��'��%j��2��-i��Z*>��Zb"�%Vx.,s`o�k����		Z�L��p�@<{h�����R�ܢ�	�]����f��Ot�1�H�/���e�K�?j�S�Z6	a�˕�0}�d��0
�Xb)܏LЅ��I@e�� PL� �n4�4�Iצ
����A���(,�#��Җ3xq���|%��"�;�"q�AW&����g�ѤV�Ĭ2���D�pc� u�.=���\V���*H��'bov9��$��uT��'	Q�u�,�b��PMx��̊	}As�o�+'(�~b��6��&�����;�ņ����<>��{6���yp���-!���[wយ3ʟ�*D��v�TRsm[I��!��'���6o!"숡��&�(��xz7l��	�*#�n؛9jh����'uŸ���-R0�(�(�'�Ф:�i��f�fD�&��T���0�'���2��R%^�2%�#OS��+ǧ(c[ A������MY�iK���q�'���we\���|��ό*k�.���[�Ƞ����O
���f["G��'סP���R��ve�%A��Q��0?"�V)UBt��+��%{<��k^{8� ��N/s����0��41�`H�D�X�m��=LvxyD#8D��h�/̫0f�y�C.3^�jYX/%}'�c�J�����J>=�/D�����Ԁ�4m�� ��&D�Ty��čV�@i���(��x8�CD�t|J�'R�ٱЂJ�g�Ɂ
���ɷk��`���ʊ[1lB�	}�,R�/�q���'�܊��[����nW�'��Xee��T잵XdF$9���˓?��)C�H���	�Ei��W��tQ�JL,p�
B�	4c�"	Hg�Ki��b�+�3�
�O��r�kI�����O�X�h ��"`�7�;y����'B��SA� �W�#y�����'a��S��Ԃ&$�9GrH����'0\4�e�׶`B �1-,�'v*Uj׋I�>lR竍�"�M)�'�ᓆ�� ��[�^7*��X �'��H`��'$�<ӳŞ�1A����'�j���^p4�"��]�X��'� �j��	�2i��Ѣ�N�p���''���a�E��-8��8���K�'��k1�I�{ �y�f:��'�N���I�Q��5)+p��`�� �콉+�>M6nD��KX+X �ȓ���6��g�Z�9 G¼��	�'����+�=�hr�$�2rW Eq�'�R(��G�d |ԫ���d1�,��'�
���jA3`��M���ҿ!�\�c
�'����Б3��qc�� #�4`
�'jࣔe��e���"R�Y�vn����'p����+y���&ѐn�؍��'3L�BU�el���T�@,R
�'T��ׯ߱4�>UH�!��V�Jd)�',�3ҊD;:��&�Q�LS��'��庑H��NbL-:�1��'l��,7?��� �K�1,�i��'���¢P�)5��G���*50��'<�=��	:Y�Jʿ)&)P�'�ԈXGHڷ"G��qC)�)"�����'�1�g�H%<��a�������'ֲ�RcA��z�
��-H
=��'ޞ�4�[��l%K�Þ1=����'�����iD8���3d�	�'v�={�i��$�mHc��9nD`�'���)Qc��L ��'Pd�'� f��:��I�ŒhU�z�'4M���ޛ������	jw���
�'�H�#	)SD0��Κ�0un��	�'s$�ʇJE�%C�W�7!�,��'�F%� ᚙ4>ڔG�4/�B�p�'Is&폵���b��$�"��
��� �����8-�T�2'ց."&�	7"ODa�Ò�tO�ZF�;�f"O��Q�W�8 ��pf^�pG�w"O�A`�a]-"�&��/H89E"O�1�'NR�H(�f'�^�� P"O41�M�
Q�x�;��P7p�&�k&"O�h`A�ύ���t�\�4��8�"O��q�SK�cV �;K��"O��	�@A�.�RU��i�!"O4H:7���:l^�س��4t(8�"OD ���ֳa�(ABG%O�y<Y�"O.@�6n�*TU�E����_�J|u"O�l8gG�8[�6\�'>����"On��dh��$u����'����0�"Oԩp.�<�P9�/�����2"O�ؙ�.ћ��zW�A��q�7"O�d�EK�3ܖuH�0Q�조�"O��E!I�4}��2�f�b���r�"O���G��A����C�U�)�d�3"OD���)x�0�� ������%"O�,��Xx	��Ӭ��5����g"O4x2�/�!8,�h� ���;"O%K"��I���3o]�&���G"Oj�I�䀟 ���q|"1��"O�a)�LF�"�Di��"ߝ'j"O�ؐ�Y�F ��a�W#O���""O|�RaY$
��(D"�7g
x��"OM�v��Ov< �P�}j��X�"O��j�a;0��Q1,��#JtYa"Ob��Q�!x�l�7At١7"O��۷��J�έ��+>�y�"O�T��@�S��p���	;�5i`"O6��oR)\�t	�F�D\ `"O�Y��-�H�`)Ǭ1�l!0�"O��w$ڨSw���h�6�H$�'"O�l8hT6��1�/���"O�hю��V�N�S�k�l� t"O�I�D)�5��}y�jO[@��T"Ov� �(0B���F��T1""Of8��eع'^D)���j�s"O<� ��n@6��a�6�,��&"O�I�ł\:��C挺kpdu�""OL���ծ.5�)�a�V�fnvp�"Op���BC�P���2�BBx�Ж"OT,��Gί|�B��AfV(A5�(��'���e���X��'� ��k����*C#�����'V�I� hn0T��>`����O$� 0N-�0�K�"|zL��E��prGl�`_���u��[�<�W� v�<�Ƌ�?4g�Tj���{��D�'�Ԉ)#II�h]�ϸ'{�F��3R�B��g��CKj��	��8AF�?7�I�1@˝%���s�F�&>��##Θ��0?���Ǒ=44�ǝL((P&��O�'E�̀��I�{&a���?!��!�^Î���(ͭX�����E%D�!C��N��aɏUwN�g�<�c�9L�Y�Hߠ�0|r���7jʜ�c�mΟH8�@�"�}�<A� -޶��Ӊ#5" ��ʒ7A	z��'B���@$�)M��ϸ'�D�d+��Z�U�����M�2`���}�H�Sd�@mO�ͪPO 9�,ȣC��}�́v�ح�0?��(P�V�,u��|2�d�F�'|^т��G>@��(��?	����#L���eӹ�D��Gl;D�H���Tp��@B�.qN�!"K7?�7�Y��cd6}���?	���6mB�HZ��R�+]�+�!��lN*�S���g��1i���<\�'�4y�腌>q��'��I���$I�N�+'�ʆM������ hd�qD��Lʩ�P�Q�H�Z����'�x�����&� 4���;��ώ�)����ȓ7j�׈�8�a�A�E�l�D|¡F�B���S�	-W�$��6(��|���(�ϢZ-!�2(��	���QHh�9X�IL9?"��
8�����C��ӬbJ,�y��iIv��f(ݜت(���R�'�))h^5v�2f�n��p@�>I�*A�Ą��GX�Q7�»W��d�f�f�p��5�O��3��L<PI����&O��(�Q,g�4�G �z�C�	�L������{���j� ݮY�`�<����I���EbA���Or1
f��2K�m���<`҈	�'�VUsd�_7/y
���.F7b���if,�D,�E�R'���f�S��?���ޢ �^z��]5WHx��s�<y�|E����;I<֬3�d�!��d��-��u�&��%o
����,�8�M��e� �؆��|��CfF0���T��قa���2�"
�D��4[�Oԑ{d��'����`ե|�l��I=�Ĺ+ć&��Ѓ oUe�S<ߜ�Y�A��\	��S�A�}PC�;4��k�MO05������y�Ki�<e��{�k�yn0Mh��!������
 �a�T%K�z���.0D��*Y�fu��ZiR�m����fڲX��7��]�*Y*���d2�`��HO>%k�@$�`9А�@�k�1z��'j�9j�2e��R2o�W0�hR�b�>:<���ʮ � YC5�'"��╉G����	��'8�
���z`���F�2���wr�0@����Q)�ɟJ$L0��0�:#�@զiS����ߘoB|h�O� ��T>4В���'1�P 4�2�\L�qL˘
�^مȓ ��8�U�����wm.��S��L���=-	H����L>і��B��ҁ�Y��D}ɀ�}(<Y�!��z���BK�{&1 �c[�L�����9-�����gRP���'8��<���˛D��L��=NtB�)�4�L�<�ܔ`�j�C�D*$Cu��͆ȓ SA)p$L�*~��Y�,�Ĵ&��`�X�*�Ш"�ӭD2` ��a��)
Y(QAH; 7C��
�v��+p�� *nU%�ALP���ɦV۾��O��!��[�T���8A&��6����ROry�t��(C� : �͏�\�5kȶL��Rt`O���>��dD 	��Q
�/�� Z���fx��1
*��8z�R��Y���X���eIZ�t"�l,D��sv/һO��3.�%b_�X�+4�E�`Y�D"ƋT��ȟ���a�7F¶u��4Y���"OJ�!N3)����`^�8�D��CT����OFɂ�3?ـ��$5�.�S �X>cT"5��S�<�$fۯw����:~�0OЌJc��j��x���S'̖�6�֕��'��J֪%D��	`"��=�ʹsRjMz�����,D�@"Q�\- ��0 �GL5g���)D�)�b��V8Tӡ��F��%j�K&D�X���ݶJXH��j� ,�`�	��:D��iG�F�}�����N�W�J9���5�OH1����M�vJ�p �a.Ŋ9!!�	i�<	�b�!e�����A$�H"��N�'�pTf9���#jN�TrqJ.k<����1�RB�I�8�\`�˥E�Z�0/Qj ���k��w�Dr����@#�<A��șY�eb���5�z�)��d�<Y��S�S����ƃ�&�0�"6��ȉ�?c( ���RM�'Gr�P���&|pHƀ&R�^؉g&��!|�ϓR�T���/+d%��g�!aaT�acƊ�>���竁9FE����d�WqҌ�B�/�'PF���oW�a��Q��T(�u�>�㊑�X>�Y�J�!2�����O�L]�R�˼p��$
�v�CF��7JE��cb+���q��q����V�>E��V&K��(�!|G8���ѷ~�����/H\�ԡ�dS��?�w*
.�<�aEK^�L�D"�,nrV�I�X�J#�4e�>��M b�Vu*�m�>A�'�jk�
�	��d�t�~��d��Ry�pq3e5H��Us�m�N� �q5g
4W�#=�Bl�&Y䲑�f�ݸV���J��UV��ʂ5�ޅ{5@A��Lq�e��5�<�q#��~ru�K(-��9!N�s�̽� |�ፉS�"�#r�Ζ�iP��	�o9���0�(W�8���9	N@ZC�Րy�b�(4��JM����`�$5�\	��@y0	���K8�ybI�|�z�H��� =1� X�Z�����;��[���Φ	�"K'�*J��>�O�c�+N�6J��@Yo���A�w	XA�}c֥	0j��Gs�  ��E�~�n�Rܢ!��G��],�3}�n�!ŤPP�b�_���:�����+��rf�1m*tu1�n ���a�@x�S
�t�$jA/ �J�c KG]E2�!V ���*p?��xr'��I�z��@40��ɰ�(�)M*I�Ӭ� �rdc���8����d��=�~)P���t����%(s�����<I���+s0u+ɾU�*�ZFA�A�'�� @�Y�=�D����w�D$�����]�t��V��}!תE�-�0�5�G-n&<�'�Q�'���"q�].>)��B��Ib����4^&����cZ�ҧ�ʱ/N8���(���
1#�q��u�o�.�:��E�Ṯ����_ĸ����L���Y5�͈|@�#g*�0b�剈7'�I3L\�|ȜQ3V�S7{zR�X#���;w�?ac@�}%���a��\�Q��:�O� �@M��
���c��<�R4�Ǖ+�� �%É�%GT�q��C/D�v@���
�[6Q>%�u3O�z���$+���x5C�#�t8�"O��wb^����SCH��H4ѕ���'�!��
�M1��#�f�ݾ��OR��KN{8T�D����x�'/N�+��H̟��dǋ
������)��l;�
�dv�����Ѽ�a~��u����&
��<q3`G��p<�W�*.tʔI,?y��MM(U��$�X綈A���^�<�%!\�C�E�h�
i�qI�MC�d��ب�2L��0|�V�k��h������Ԉ�Q��<�d W����z�@�0��P@ �P�J z]�O
�� @ӣ����0�RT�1b4�ՂR�M��z���
�C�L�N�Dn �(��ɹ�@�G&¬���$�O�%0P�m��Rw�(&�N�"��'+�t��N�&PM��ò�8S{J��r`si3��!D���*ހ=C�s��&(;Ud!���纉��4�)��=U��[�b��5�|Y��h�2C䉎1I����F�i�xl0`$�>^
�C�	7"����l-�l�q� <A��C�.�F {�#B�K�8����TrC�I?u	
 ��V��eY#�y���'���T�ɦ*q�Q��*|���'�p-�3F�;���.�vv���'�����3QO|l��jR�dp�'ShYx��y�tK���z��e��'�J��Tf52��E�hl`�"�'S��8a ƔyU����Kݜ���#�'���eg�|O��yVe� ���
�'-�q�B\J�a��k����y
�'G�ȋ���?c���Ç��©$D��`�
ԨG$.@b�덭��iy��(D�TS�h�9z;�椟�Kp���'D����) V�:/ݠn
z����#D�t���nrH����X�\z �H�h!D��r*��pY��2�A��>D�`ا��P���
K?"Uc�J?D�بD�jyZY@$�O�j|TASF<D�`�A)JMD��2qj�?*2���?D�3��4O�8A9$����ۄ`:D��	@M� *w��v��Q�$D����E�82g<"&�1_)jP���%D�DaC&^'{��8!�%߇��	�S�1D��2��Y�,Ҕ���s��L�:[��B�	�6��=���-J�ERA ���PB�	��<	�,�9����v���m�C������7W޶I��~K�B�	�fp�Z �g����PBG�8C�Ʉ:��mZFB�yrY�%X�K��B��<���*�Ɲ}4q��*��y0dB�Ɇ�&����0�QY�A�@�^B��Wͺ�XčT=�,����9|�B�	SM�Շ�)&L1��/J�=\r���"��4N�ԈAŐTB#>� r������}�o�S=�i��"O��8����&�uC�^!5�"O��sŠ�Rp�E"�5�Ģ�"O�%pa��=2=��*4!�?�:�"O�!�1J�wy�U�a�j��x�3"O��ЎM�u�ЙRE#�(
~�tj�"O��ѵ�P�U����"��<W�`�"O�y;P�� EH�bdV��P"OER�	/M?:0�p��]��i�"O�г�2�tR��۫o��d�"O���r	�-sT�q2��E�R���d"O2���n��$�Pe�ˬ��hi�D��ē�&��~��m��~�7hњUOnq�p��3k�4X(���q��Q-O1����|�!��o��A�ƫ	��󤥃�����l�����ߧ-f#nZ�Gd��R�����F]`�<Rpp6�L�[k����(M:��������O���[O�9$.l(Ah�;f���QP��<u0�S����Y��0|
gWlŠ��	�A�L=��p�r!�6��
?ꔣ n���өg�x5W�9W�qSB��]��r&��<�c�[�%e�lӵ�?����|�.��i⦡B���U���0K-´@�Gܦn(@� �
����$y��t�O�`���"�L�,�!䍄���c�4V�^ 
��Х3���8�!�8bla��
�.S(P{&ݻ:F�`�נP�)��%�"�B5gsҹ�s�n�P�
�'bu(�-��O�]ig�n���a� X�eCw�S�<�'an��T!�@�(���@'dؘc�>p�5�x�n�01��z�)8(�m�1)̛B�镇���y��N�W��Pℼ@�>}	�F��yR SL`���R6�R��f��yB��"/��*Aњ�~��ѣ�y�J�~�8q���]�b�囡�M��yK��a-p1jQ
�JD񱇧�+�y��6, ��S�=�r��g����y�:� ٵ(1�`���^�y��/���!�D̛6�ĳG����y��M�C2�5����3�8�:��Ӧ�y��C�������T�,vN��"U��y�ZǾH���ԟPFN��P�L5�ya�.TXR9�H^�W�p������yrϙ7���`ǅ�TRj4���yR�H�9�����D3#$\�e���y�W8i)���C��=���T���yR� t�Uq�m��3��2��yB�T�<Rf 3��!��r����y� �*	:�9�B��#\��7N@-�yBjU�^�L��f���Ԡ�wN�/�y� �=!Y�i��1��i:�4�yr�U7f����QR�/6P�GLS��yR�F�E�f���z�t$C�*©�y�,���Tu��°sp�a�f*���y�n^=@DE�&c�o��y��Z��y���G���QdbںNFѻ`��y�M*bЮ�"�ɝ]ڌ��ġم�y���-����DI��VdL��Siɚ�y���8?xx�T�U6H@ޠ#c��9�yr�+'^|�7-�7s�v����=�y2��7��mЄ��f���1ǁˋ�yR�/-ɀ��0F��[ڑ��ُ�yB��'.�恉 eH:K�ҍ�U�ӧ�yr�C�!爸�ek92&Ґ�!�>�yb�Z5�8�7�Ɨ>@(�fH��yB�[���ex�+Z\�P[���yba�KhL��`E�V|Vb�ʳ�yB�oC��� R��aO�+�y�Ɯ�X���-�6Bx�qrp(��yҠJ'#�x�+3��)7�ڰ��(���y�&4]܁�U���欘�o60!�� �q��.Ҍ$B85���gƶI��"Oq!�#�w�>���DE!؄ˢ"O�!��A�����&��h M0`"OdѨׯ�d�z}�t�X�Y���"O���[0?����刮!���"O�:��}���1j�*j�A"O^��PeտK��bp(�&b[��p"O�-	����;�����A�8vnѐ"Od��b[~��zR!��
v\�"O��G�8������4e�Ř�"O~��&Ħ⪱��#D!z_P:�"O���f#2RzPٸt"�'5�Z�q�"O �E�:���s��̶5��#�"O�l*g�W�Y���RAؐf0TI�"O�M�הZ��`sPB�'0����"OX-a�m	�`L|z+A�:	 ��3"O�9JGOOpZ��Ý�)���"O��r�DB�����/�䥱�"OX���҄G'��Z�3a�Tԙ�"O6�hR�s���0eQ(b�Fq�"O���� 6h��;�d��8c�"OxPFI�"�!��߉	��m��"O�9AF�î(�jH�#.��I�"O�xx&,�U�X(3+M)��T��"Ol�&Cõb�� �e�ũe?
1�w"O�1)��@[��Ѧ'�;Z>ف "O� )��H$SC=x6Ŝ�!��s�"O�QJS`Si�IR��f��"O<K�.�&q;�}���B�[D"Oԉ�է;���MR�or�!"Of�4,</��M�	�Y5"O� ��K Gg4kD뛽-ʒ24"O m{�!J-�m�D
�)�\\��"O���K�u b,���(@��	�4"OB!�G'V
�Z��p��m�3W"O�H0�\q �i�׋s�XI�w"Oh��&	����� �2���x�"O\��J�7+ǈ�s��ҩ'�@�z�"O"i"�N;o����#��7-�,{R"O`y���1����_�}��c "O�)���=���8sf�n%�a"On1�E���g�]�P�U$|�"O����/*~���r���+0�H��"O�	##�īu�#d!X�=�F���"O�[񂍹�1���T�R���"O$�q��	Py���F�T"C"O~9��!��A�l�b�Zf��N�<���M ������zV`�I�<��"8\��G���+]���`M[�<��-Cˈ�B���+���pk�V�<3�i2���G@�?��	�-LT�<i0,��rY q�E 4D�f1�Q`G�<A�`R�j�j��ݭq����U�IA�<Ye�
�X���n��zz�-p�T�<Y��ҩ$��R�+�����vH�O�<IV�؞)cJ�
g�� 5�!�W#Iq�<y���9�0�3� �/����Qn�<�b�>Q��<��	>u���,IA�<a��ˈ��"G���� l�<���;�����eN����Go^|�<k��~2�ȷ�Z�&�1����v�<i`J��| C��P
b����Q��J�<1šV.i�$�p�Ø�ceD��ŊL�<Q����
A��;S�MR�4�P�Lr�<� ���&My�6��%,�?:5TZ�"O���JG�B�@l��%���"O�]E$D:!0Ȕ�X�d��d"O09�v�M�5d]À��r��"O�� 0��*z��ʎ[�0��"O��H�$1'M�Q����Dq�"O$�ۂ�R�nyV$�f��06���"O� ��^>q�Lq�ǘT�`	��"O�5��Hd���Zׇ��;"O�m����j��)8G�΢y�j��B"OM;qlU$_��8E�7N���V"O��:灌!_S�����`�n!X�"O��'W�nl�ly���x��ȓ�"O��8��QF,��P��� ��h�"O�]i2�]*=� ���3Tt����"OƠK�V$WmHPk3Ө\�$h�"O���J�F��*�(P3Ix	�G"O*E���۔���A�"�`3XG"OĹaN� �*�Q�=[0T1(�"O�X)�M�8p!ܡU��!B�p�"O�����P M��8;E�SS��%��"O�����|���&?��
"O�hJbK�'A������r�!"�"Ot;�+��JKn��n��XsV"O }�W�>�t� �Ѩ)l�8iE"O%��H͋b��j���N(jV"O��	��ڻT��Q�ļ�1�C���y���0{�6�[�[�X��!�u�0�yB��9Za~쪵G>X�٨�jZ	�y�'�L#X� �󊆧�y!p�H�f�;%�R1xӦȧ�yriS�l�J�A�&�j�Y�
�yRJ� U*��"Hn��1��A�y��ݸJ,�̻��P%7PX�Ҡ�0�y�a�_=��+�B�A4 �!�.�y�/D�����4����5ͅ$�y�8K�yJԡ$P,������y�C�9���3I

f���$
�)�y2G�"9�0���	Ι9�,]:����yr�N�x.�չ�n�%h ���`��y�/�	�$43��[��@��D*�y"�L!y$�7@X�N���_��yR�F3����ǭ�8y-��Kȏ��y�l��:̺a �g�q��(�R����y��_r��J�gT"p��u��e!�yR�DX1
s�i+n��u�a��y�ĳ�����O��k]� Y�DU�yb�[&� ]�$�HeKX\���y�M�t"�����\a!��Ɛ�y2��ba=��ț`�ޔhPC)�y"х2k��@I��#L&���ƞ��ybI���ʴ񐁛��:D�S�L��yb
�2W5������z�����_��y�D�q5|)�C	�4;"Xe�n��y�C��H,<�$-�2,0�ô�8�y�ʛ�s�DP������`M�y2�U ^�x1�iI�e�6�@$�[�y��6bp�L����K����2����y��[�b��i��)Z"r�Z��q"�y�'	�0�Ա�A�ޡ=��T�`�F>�y��s�$�K�	@�98����G�y"I��y�n404�2>�����㑶�yb��xD�͸� �'63��Q7́&�y��@�=�vD��L����%V>�y
� ���$�V�����!J]�h �"O�m��3^� {D���D"�"O���қZ�2S�X�%Ҵ@PT"O�œ�GO�o���1�n� $Pd� "O4��6���`+AȢB��څ"O�ya6��|/�|�Ȕ!�.q�S"O`k�N%�Ze���$"�8j�"O�I��:�Q@ �ΒX�P�k�"Ob	� +��_�n�	 �,Yň�C�"OШ�s��L̠�CG܌u�Rps1"O� 0�]���E	p�x�Ρ{�"O�[LG�Kl<���ٞxx��J�"O�g�E!e�)FF5do�L�"O$ ����^�����b �L� 2"O�����.l�.�Aǡ�T��@�7"O��01cD�Q����$���=���k"O�@ d��!P���ұ1kX�8�"O�@rs��7]xL� �U�/U"�"Ov��6�(��ҊW<mi$�y�"O>���hA�'$֑X��[�%L�,��"O��0v"ζt������/[;���s"O�T��<*�lp�@��$��W"O�aْ�?�6]�u����U��"OVb�(�31��ئ��/�F��"O�0���G2K(�q�t(��H�s�"O��ca�4F�"p#s�9���� "O��bOCH��xb�?X����C"OK�6!,|i�#Ye�DK��ƹ�y��0,.�3�A��z�4e��ܒ�y��
� 0  ��   �  N  �  �  1*  ~5  �@  8L  �W  fc  �n  }z  a�  ��  �  '�  j�  ��  ��  :�  ��   �  ��  �  ��  ��  @�  ��  ��  
�  M�  ��  � 
 R � K% 4, �3 �; C ]I �O R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(՘xb�'��O��(⃯"T�����Y3s��eX@"O�-Q3�&&���PFi�&��{W"Oݪo�����XsmF%b�N1��"O�����?l-�pp����k�j�w�"4�L���%U�\�5�Շ<`u!r�!D�����7D=b}�����z@Bm���:D�878B�lq�ɣ%�6o�!��޴%��q���T�D��=��@خ�!�ā%"�na���̥a�A�Ve#�!�X%0��I�3bZ�8u [�6V��}B��ȹ�V��T�S�&����pb:D��1�)\��j�;�lֱx�v���A$�B��?���ӽmTm����X�P���!D�Rl��A�65I�`^0�P,�bƪ>�������B��a�B 	�+��B�	�x���s��q�i�5@T%,BB�)� �}�Q/nI��x2�ݡ ��B��j���'4�UAW5= �@प
U�=��;�~�D.M�]<�2Bˑ5� ��ȓ�r}���X3O�Z	3fj�h�ȓM���d��a�0�"F��SBB�j��)����V�o�Nur�,��=��5D�X��5{�,�Y��M)%)D� ��N�^$��Nߒi����V�&<O�#<)�F( ����� �+���2�Tq�<A��A<0�s'Γ�N�6Ѻ�
l�'�ў�'X�
 ˑ�I�G?bb̓q7����}�`�S�.'w�h��M�s�dFx"�'L&��ħ�E?�hbl�v��'�\�ehʲ$|Ra���l"�'���K@�`o�T[�*�']a� B
���DB�Y��As��0Zt����l�!�dL�d-j��F��_�~3�iU�vZ!��8�T���	3�MK7뜝xM!�ޛ�	���4t�p��A6!�>Ю̊ �I��R�r��/9!��0K9�E�P!�,Vzډ�sG:�!�
#r]0��)�.=�%���B䉱RR~��E�A/^S�ɇ\��B䉰-dXӌ�<Wy,�x��ɌB䉚��#�]���-��,�>E`B�I�$wD���!ż��9�e�ͣ6�PB��V��`����I�����U{�:B�	�Z�փո;�M[�dA& ��B��,|��1B�	=C!$ccM��B�I�5���̝~�:5c�c!h�`C�ɤ�)*�%�7C�`TI�-�D��C�ɯn�l��3
��2,*к�$8:�XC�I�LP���E�3ZY��q��ϩRd6C�I�U��{��9Eֈx�N�X�$C�ɚa�4d@E�Phu����ό6,#�B�	$Rl�@�d�I�H�j�ba�GhC�	��N�brD�!t�XT��UT�,C�ɖ7>�Y�#Ó�y� ����HB��9?�B�P���?5�q�񥅻b�B�.zY@S@ �*l!�(�1"�B�I�s�X8��`��9�L���J�f`�B�	)PN5c���,[|�jE`D{�B�ɻ}c�PbC�
4 �[ o_� ��B䉀�82�CD���5�W�A�RS�B�IS3JU[FK˫W��M�*L$idC�	����PM��U(�ꊹ'�\C�����'��yM�U ��!>C�I.{��8JF�Z4mq(�@�C7 �|B��z�\$��m�|�J]�5G~C�I{|6<�f��6S4��h�<��B�	����ha΋=�~��`	O�>��C䉂E�4`�R7T� $�L�y��C�	(���F�F(C:<�C��:oF�C��x��Dq���u��g��C�I:sb����;g�} !%�>@BB�� =����
�1!оY^B�ɜJ���"&R�/�d���L�k�&B�
^#�%���H7�vQq�		l%�C�Ig.(���0o�XM ��G(n�~B�I( �Z����IczDq#�#5�|B�	�5��5s�O�{ˎ�	$�UBlB䉮qDؘQ�dqN͙�C���B�I/ôX#U����#p�E���B�	�+aF�r���f"!��=1J&B�)� �q!O��<����*;2Yh�"O���UA^	4 h{���+ �*u"O� ����T�!�kPp����"O���#�Y�9p�0��o� X)Q"O�|���^�w��4p����
��'dR�']r�'��'��'��'j%{p�S!)<]�쇵^�:u���'���'Y��'�B�'�B�'�r�'߀�/	�����%�1�HK��'V"�'c��'2�'���'�"�'X~�8��UxZv ٖQb��R�' r�'���'���'�'h��'�lT�0*� '(x�:�aɨrZ�@���'�R�'a��'k��'^��'Pb�'Ҥ��� �dԼ#0�&u� IYq�'^��'H��'`��'rR�'���'PV�����C�t9��Ň�?��J��'���'d��'Jr�'���'�r�'ܲ�#a�?����Ĭ��@52����'"�'?��'F��'�"�'���' ����H=8�<đB鞡7���r��'���'�2�'%2�'�"�'b�'qrMw�N�M�H�3��y�	SF��?���?���?1���?9���?Y���?���q��e���M�,��UK��5�?���?��?	��?9���?��?�V�K�@6���,ۘ
{i2�G��?����?q��?����?q���?9���?�ԩ�lQt����r��1���?9��?���?1��?I�-��V�'`R��fh�d���jBt�����Y�`��'�U�b>�l��D(1���A?9n p� H�I<\���O��lZC��|��?�)O�F*�YP�T�0��$v&@%�?��VX&�M#�O(瓉�:J?5���[�,�V�b�u�0�Iןؗ'K�>�w��2f)4J�:Q��T�����Ms���l̓��O��7=�^�a�'ˁ3���k�윶w��!r��O2�Dl�`ק�O�nI��i����
�2���ґ}j6Uuk�4+$�b����P���=�'�?A�h�c
�����T	a"���<i)Op�O�\m"��b�����Y��Uʁ*
 ,SX�B�n�Q�s��	ßT�I�<��Onȋc��;�@�%#Ω=|������	�~�.L 7�"�~�"�͟�qeA�g�(��*Q2^�R1�W`YyBV�4�)��< IO8n����C�����o��<ɣ�i$脹�O�n^��|�7�X�`���J�옠b���OR�<	���?���#{���4���{>���c	j�xT·�?k���&�Y�,\��;4�&���<ͧ�?a��?Q��?�gBR���ZJ�2]v�}��eC��?q��,jZ���O�'�?9��?�������Od) ��
o����t���b�2X��jFy�'����O�4�'�n�1�Μ����3EX0Pdn|�@L*̜���'K�)%�Ƌx�\1 ��䬧ON��(O\!��$���	�,�"�����O<�d�O����O�I�<qq�i6�X���'�����J
-U��z�0{T�庀�'��6-7��)��$�֦Q8�4�?�Q�[!D�[ f8`2�;���y��ٴ��d�7�\�����Ӱ�u7�w�x���� (HY��A
Xv�}p�'{��'Vr�'���'�lCbaL�ȼ`"�H��t�5�g��O��D�Od��ɡNg���O(nm�ɊC�Y[Uޯ<����ދH�Ĵ$���ٴw���Oβ���i��ɋ��]�e���QsF�B��$I��I���Z.rf�ny�a���|���?���s��<`�j�$j�&m����2q|n����?9/OX!�I<�d�O>�Ľ|zV��^(P��`,ظ��#Dv~���>���iO�6M7��?�;D��9ur���Sa�.IxWmT�C�YPT�W�M���'��n���?�'�<ͻ�ؙ8VÁ1��Xsb��[L|1��?a��?�Ş��d����r�,P2oad�S@��aL�ś!iU#� -�����޴��'��nB���>s��x� f��bZ���Q�7`�6-�O<��q/mӰ�z^�M�#�����O|�5!%�υU��=���@�!s-*�'|�˓�?���?y��?9����	��sQ�8��&@n�Rpsp#A/h���	!l���O
��5���O��nz�+E��J��H���x��� �1�?�ٴ����{�:�B�4�ymR�C}�Aʀ�6p�����<�~��E��u�7�\ʓ<ɛfR�����	�BJ{�ˀLT�_;�C"+�ԟ��	� �Iuy"t��M*5J�O����O4PY�I�\a24;���g�xa #����DT�eC�4��H��H0������	�q��,�'�,�y�E� ׀1I�\�;R)��D�	�?��
�S�1��Bx ]	��ݭ�?���?����?����O �J ��^;�9Ȗ��c8F�¦��O�`n�3B�����ȟd��4���y�O�=;�,�S���,yN��L���~2�'
���'C�Ur׼i�ɞS@P��O��Ћ�����2Bf$�aU��W}y(y����|���?����?)�\]C��D��ge�9Ѷhz(O�1oZ�o6���Iß���c�ß�h=��p�E�Q����.^������
ݴ��Ş V�6�Q�b�@��:��a�%NQ:z#4!�OR��j���8BD\��Aݴ��$D�� @�N�H�fD��N�a|�t�� �w��O@���k�g�"����В+�4�K�-�O�HoE���	�����蟬 �Ǎyo0����(b�F�{3k��r�`nZ]~��M�]� ����'տ� P�K�
T�ى��K�:����<O���m�`\�A@-sϬLb��K�%� �$�O������7�r�i�'/�TH��4�����M38a@���B)���OD7=��4��b���H8��s&�&��$���O%/sԨɠ���.c���H��䓭��O��D�O��$� i���@
��
tL �����O �z4�fcؓ�yR�'F�[>ɨC�=F��@�@<#�0]��i1?��[�ܚ�4It�֯1�?1Vf'}`41�S�F���-�2a1�qj��?sP���|�� �O���K>��m�o����+�9W�&DAU��>�?)���?a���?�|�,O�o�r�vp��V/-��p�	L��cL�ǟ �I;�M��B��>�Ӷi~�m��x��I��ȉ�(�+��wӨ)l�V�l�V~M��x��i��L�IS�:�>��gʓ3�Z$+��-I��D�<a���?���?���?�)��Q����������C��M��.Ȧ!p0���T�I�� '?]�	��Mϻ(&���A&�;isr����|h(�D�i��6M[\�)擏l�`o��<9�� ?��$r)�iXL���E�<��X"y�v�D������4���D_!i\� ǎ�:#i�W�#_�����O����O$ʓ!��T74,2�'�b�(��uXQ�S�3FX�3D��<�R�|��<����Ms�xҤ�e[ba��@')���릧̳�yB�'���bʍ�LG�l#�O~�I��?yF��OV�ք[]쪩
"�Q��Au��O��$�O~���O�}J��B;����
K��Y��^'tk|K��\���( �3���'�R66�i޵kP,R6�.����o�0�(U"v��ٴۛ&�{Ө�z`kz���ܺ`��埢E�A���X+X�r4g@抴raN������4�����O����O���L>�*ǖ>�Y`P`ŐW'��|N�F�/��'����'|DQ��k�/]\ %��y�Z��S�>y���?qN>�|���<L�ƨP�	ړ>��J�f >�r�9ݴ#b剢6� ݱ��OV�O�ʓ'�°%�v�x�A�ǟYNV0q��?���?!��|�*Op�n:QO�,�I�Va���4 ܛ%A�$#i�g����	�Mc��>I���?ͻC�ٱ��(k0��b�B:ZE�_�M��O��>�����4�w~	�$IR<)츬�K��Φ���'���'���'h"�'���y�!OX1p*����`O.Z�H�嫿<	����搱���'�6�&�� �J�i��b�&L �ʔ�Q��O&���O�	&9��7�2?�;2��h���	��0ж#e���"���&�~�|2V������0�	ޟ{@�իI��<s�f�<r��c�������~yR�hӦ��
�O��d�Op˧8�]� e�{�XY�B]�o�L��'���?����S�dk��t�v����(F�	t��P��pJ�Ɖ$r��š<�'0O ��Q�I�YE�V�j�SuCN';jI��ԟX����)�}yr g�2��Ԋ�+J`P8k���:z�t����ʓ{���D�OH�o�l��~��I��@�gE@"	nR��)(l�Lԟ(�	�8��lZ^~Zwgn,Z�ݟ�˓n� }3�����X!-�e������D�O��$�O��$�O`��|�ƣ�v�@]3���,f4e����*L��� 1k�����\'?i��+�M�;ecp�g����h�akk!6�?�����S�'j�Ep۴�yrEȝR��AE�O1��9�N��y�O�/P���������O��$U7�V\���-���%��S�8�$�O ���O�ʓ?���� ��'�"c̖Q\hTI�˼ e^\���(G5�OBI�'<�'f�'���<mqӢ#H�K&�r�O�0����a��6mg�ӫN����O���f���HB:as6�M�]$��%��ON��O����O�}�;[4��N�$���ht�Q�)������$��N���D�OޙlN�ӼC�m����8h���4M�v��$�\�<����?���~*�qߴ����u*���.(]��/^,=5H�R�ր<�Z(।2��<�'�?����?����?I��=.o�9	��*E@<���׊�����iK���ƟH�	ԟ�%?�I1u���G!UƆ}R ���-�q�/OR�$a�ld$���$�s�H��@��}`tbd�&!�j! �8��OH�B�ty�kR5=���{�
܀���0��T��0>���i�,�ʖ�'ꜰy'�C'	��e�P�>c����'w6-5�������O��$�ӦM)P��0�@�"�	�1�B��qjBf�J�mZs~2oǸ	J�����'����dԖJ��3��9��t��<����?I��?Q���?����) 4�(�I��ֺbȘK�G�g�b�'�Bj�6�s�<�
��R�]%���s�� Dp���׉n������(���?���|��Ɂ��M��ON�q�k�F���&F+��-,VOfaA�ʌ�0��|�Z���	�t���� ��εn��r,�:F�B���J�ş�	dyr�d��Y;d��O.���OT�'؝���0*����%>Y�ִ�'9p��?A����S�ċ��7�^��L�z*D9�
L;a���{S&K5*�d���O�	�?9�� ���r���3a�43��1�f�+a����O��$�O���)�<�3�if� �� �^�H�0$�E{a�Tx��'D7M$����Ā�m��O�^�,�Aj *����s.�&�M�i|.
3�i"�I�_.����O������ |���݀g=.0��g1<��0O�˓�?��?����?����iR@o��@�@�M��=�r��,z��UlڦcL��I�����e����	���s�e��dF�x/������'�?����S�'mq6hq޴�y�he>0���Q�Z�p�A��yb惘b���������Ox�$Z~ZVu�D��;|9Q7�ǹzS:���O����O�ʓ|)�f Ȅ>�2�'����WS^��g�47����A ��Ox�'��'��'u.EI�c�-2�"4��k�);B:���O�E�e�Ea6�BO������O�p��DG�0��RoͺLPdU��f�O����O@���O
�}R��V�N�P#�J%7t�1�cN�
� ��6����fFr�'��7�$�i��[5 #u<0����Y h�D�S�ee�0����ɌLz��nZS~Zw�D�[�՟Jt�QA�&��:!K� o�0(�-�Ī<i��?i��?�����1)L �{g.�Wq�iP2^�$�'.67ҳ|�����V�'a�O���/ � ���1>kL��	\�k���?Y���Şd�V,a%-A5[d�9#.^ߪ���Bл�M��_����c����6�ī<�'�fb�u-A�^$��-�?���?i���?�'��d�S��V�h�b$כ0k�T� T��$�jR����۴��'f���?!���?!5`ֶz�(���(a��|YQ�۰n�JU+�4��EX�V	��O�O�'.ȒGQ�+�{A�qju ��y��'�b�'R�'���	ѽ'��7�'0�dR�G��1���O���C��3[���/�M�H>A�B6��gl�4/߼�����$��'������A�h��曟0�*ۧ;v�ZW&ߪ٢=c���1
O����'q�&������'�"�'���[e�5u��Q�F^�8�z s �'��^��J�4_بΓ�?����	X�k��@ZF�J�O�H�#�/��Ƀ��$�Ŧ@ܴ?�����^�."�-;֋��q�xl��H��!��H0� Z�|�`�����&�2WO��!{�(C7 B*tn>�hT�<_���I��l�IΟ�)�Cy��aӬ�s���T�H��PC�G�֑K�ˆ�Y�����MK�2m�>���i�p!+�K�h��c����%kw�l�o�%dƎplT~k	h,���\��qAk��{<��cgZ� v:O���?���?����?�����ߦ+(�Au�#<r�1�T�Ƨ-0`�n�V5l������	~�s��i�����nZ�1nL �S%{s !�� 	�6�m��P%�b>�c��͓b߸���.4�2�	De�ER�I̓?��TR)�OQL>)*O�I�O���AIԘ;�����K�yb�O�$�O��$�<v�iEl�A�'���'�Ber������X D!�2kѐ ��O�e�'86�	ͦ�M<	rU�m�V���%ɥ)�VԁH�Q~"�KK��DRS
P��O��d��@��Y�6�z��I������Q
^�r�'���' ���c��nx.�(#m#_�n�����ҟ�K�4����'�6�=�i�i�3<pa���<��(v�X:�4n��oӼ�JG�y�z�x��/���J`-��x�a	v���2`b�,��A%�Ȗ��t�'��'B��'T��TGF�:�IQ
	'Arj�@vT� IٴH���?������<���ԧP	h�P�A���=!�-/gI����M��i/�O1���YQ��5���`VK�-O�E���U�����Zs;�{��5�O �L�ޭ�F�~d�8I�Lx`���?1��?��|�(O�nڨ|X�q��(j���;��M�w(D���.��ގ��I��M���>���?�;r.��Tl�7�B��#ˉ�{�(� �T�M��O�M�h݋��t���w7�=�FNR8 c�=�%Dou��B�'��'�b�'+b�'�N��NCH1�(v��<�Ju�wn�O>�D�O�AoZ�X���ǟh�ٴ����C@�Ь)4��㠣ٯ`xɫH>����?ͧ)�bSش�����chϦMx�ͣW�$��R�HY�3���Io��Xy��'l�'G�T�\�i�G1N�����-cR�'��	��M��eB��?����?�(��-J6+͗l$�ib�9a�h3@��,��OF�D�OԒO�S�rG�Q To��b�	J��	S�Y+�B�	wְo�)��4�Z���'��'DM�1���9���󉞼�D��'iB�'�r���O�剂�M��J$���J�Ä�%�| ���<"`@��?�0�i��O�D�'8���;�*!�U�EQ�t��Af�%	��'VN$��iR�iݙ����Xb)O�i�Rd�ܠM*f��5,�
�3ON��?���?��?������e��
�F�٪��!#�oڜ ���'qB����'!Z6=�d��P�T�}ux�E��+�f�A�O���7����-��7�n�$
�!�>Z�x�raڏ-BR=a�Kb��S@�̈́/�� �$�<9(O0�8�f�hB5J��<Z���#�'��6-̯�&���O(��ʗ�n��vQ/k������m����On��O�%��2!��<5�NA�p�0[$2!*��,?�Da�h��h+�4��Oʜ����?a2H f$ "�CP>mL��ʵԶ�?����?)��?�����Oy��/֜�! ���)�@�ë�O� n��-� ���`cܴ���y����R͘�R�OڠH���h4����y��'<"NiӜq!�jӐ�pJ�4��n�?� h��Xn���D���q,���?���<��D� a� x(�7s`^	 p�(+���:�M;,��?����?	��$
�N�H@P#�;%�Y���R�T�1ݛ�q��I'�b>a����|�Ȁ�bn���	h)�0���\>v	��_x���� �O�%I>�*O6�)�"��SqV-�2��b!;���O2���O����O�)�<�D�i�H����'N��ʵ��:5n=���I?\��`i��'��7m&��0���O����O�E� BD 
4�� 4�B]b�/��>Z7�.?uI�?v�8�SS�S��Z��0Ri��Z�K!:��L+�Nj���I;I��B]=5�h-��}h�����������MÒ�P��
o�
�O�hb�M2w4����/��1�"� I��韌�i>-�^Fb7m>?)P"�1}�x!Y���� F�I�oY#Zr��)�� %���'I�OY�A�F%<�X,3q�b ��F�I�M{B���?i���?a(����G�9$\Ī�fĎӘd������O��D�O��'��[��-��HF�a[��yV���m�H����עfm^LJ�4 ��i>Ys��O��O�����D�&#θˢ	�8c��b��O���O"�d�O1�l�Eݛ��Ob6 ��4�&@����L� &�|"&�'@�yӞ����OP���Sֈ`ȑ�ǀV�P嘒� _Gx��HƦ��E���Q�'D2�IF jz)Oise�ւs�"U�HB�=
��3Oh˓�?a��?i���?Q���򉂚P� ,���5Fx܅��M�>.x�xm�`���I�����D����I�������j��x�f�?i�Cq.�|��i�ڒO�O�މ�Ǵi�$� 5vL*E*�8.����k/U��Ǥ�\����v�D�O^��|����`��-X�����'�ב@?6����?��?�-On�o��#ZA�I���	�-
\��K�,-xCi�=TVh�?��V�ܛ�4����-�DU�b�����J�]�.a�CC�px�ɔd2�]�2�H�*�'?թ��'�*����:����ʙy�z-!E;���I�����Ο ��o�O�R�sY�uᘤW�.U�1k�!��v�����O`�������?�;i)*D�-N\�|
S�Ӎd�(ϓ���k��\l�b�j�no~R���E���h�p�rL�&ÜH��#
��țp�|Z���	���������Iៜ����Q�N(a$�M����!cyB�b�P�c��O�d�O�����>s���%Y
����ʬ"���'+��iVb�O�O�<��EGFx��3�ʇ�i���㮒�pd�)#S��k�$��H��L^�Isy"�J�a��kg�
��X�	ŋx���')B�'��Ot剮�M�� <�?W���ʌ"s��0a�C���?�ûio�OX��'���'�2�	�aT�x�����|,"bK{���ųi��	-q@��`�O�q�H�N�Ƽ��, ���J�g��D�O����O���O��d*�S�N?��e]#��L��!_5eL���'�rex�l!�=�V��Ϧu%�d+�C٢+4����ʳhQ�ٺ'�Uw��ӟ��i>u i@æ��'ۊ�Q�9�l�3ǆZ���͒�G��Sȅ��8sm�'�i>���ӟ�	(,��ܱ3�Q����b��V(/�:A�	؟��'��6��Xh���O~�d�|��
�}�Vp�MH��`�H}~�f�>����?�O>�OӠp���Ĝf�Z�@��6M�
�[����Ԩ��4�fm��!r��O�y��E�+07�#��nm�M��O�D�O �d�O1��\j�AM�T��l�C�-�A�`P+]A@�@E�'&R$c��pX�OB�l� 4Q�u��[�1z(�DN8O�>�S۴*��a�!����@�D��3�T�~���҉&����A�6Ge�T�7�X�<q*O���O��O�$�O��'!�֝�lD�mh��&o�=H8M` �i��8���'�b�'E�O�2Bk��.Ѧ[��5�b�!':�`��=hnZ�M#w�x��D)IM3�V6OVb%f��^G�ա�/4bɆXad5On�p�?��L(�d�<�'�?�QޛM�v���tm��raJ�?���?9���D���i�,B�<�	ߟ(kvl�pF]��@>:��a��s�l,���M�#�i��O\�ꀣ�#D�
#˵.��1@V��P	�M^&r[�1b�%��rS���8" oQ�T�|(����"	|(��B���I���I���F���'��@PlǬ�*��p� ��2a��'�6��l���ORAm�c�Ӽ˗b�]Z�<P�lԼQ�LPR���<ѳ�iʘ7�TĦ��%����'�"�@���?]��$�HO���'� w�6|r*X�bN�'��i>��Iן<��矈�����Ik��^ 2�k�@.pjy�'�6��12�t��O��D)�)�O�yU�W�Z�9�VMF<;v0-�֌�T}��iӤ�o'��ŞD~�����/�����B���01G��,,�l�'-\�`���P��|�_�0zv��3l�K�;z�P��A��B9d���O&���O��4���l�/�?�#�_�o0��z�˂�߲-�����?Q$�i+�O���'ü7^��ܴ���WC�'��]:"/�L����B�MC�O:���"?�b����w�~8���T���K1@�)<ԸS�'���'O��'�2�'��*�(W��y?���"��p����Oj�$�Ob�lZ *���'B��v�|�d]gޘb�U�z��D��K$O�$n��M�'�x�	�4��d�$N�� 
-�� ����Eo��brf��a!���?I1N;�d�<�'�?���?ys��=v��pyS��_���	lN��?������������(��쟈�O�$�HS�F� I�\H�,��'��XX�O @�'\��'�hO�i�O�}3�T�:L�i`��q4V4�4A�7?����u�ݖ'����i?�O>��V�n����.� �D}���W�?���?��?�|)Ob�l��:B|i$�E=��T�T듯{��@,�֟ �	0�Mۍ�	�>��~� ����� xY�)!Y�5�������%.x����`h���N�I�<�&�	�<i�nf�q�NV�<�(Oj���O��$�O����O�˧Bb*X)��Ѣ�P���#�*�Zf�i�RŰ��'��'��O�R�}��N' d��mG�u�H��Q����D�Or@$�b>�Q�K���ϓk栵��mR�o��P��U����xخ5 f���H%��'Sr�'��	g��'s����ǫ^�9���I3�'V��'��^�`޴E~�C��?y��sD@�Q� �AT�KQ�њ_]XEY�b�>Q���?YA�x2�A04h��a��hߪ��u�;��DoѰ<21Kd�x�%?a4�Od�V�-	�0c�e.OX�k�
��\6 ���Ov�d�O��2ڧ�?��n̺$@�x CM;&���W���?!@�i�Pj��'��h��杓>h�A0��2 <��͚~�,�I⟬���M�!S�M��OX �dm�?��4��.#�z��d�@/4�ʰ�4˯/Z�'���֟T�Iʟ��	�T�	�:wXlSH�5l@H�O7\נ��''F6�0���d�O���-�9O*�u$�4}!6(�%�0-��ԱÄ�N}�qӘ	o����S�'}���a��]'@�<�B�$k54��V
P�]i���'�j�P�,�⟼��|�\�`���F-6�@V�( "B) �ʟ����H��ڟ��{yfӄXBB�O,��(^�	?v��g�M�܍a��OHnN��~���ҟ8��䟈��±@��H� �6K.p�3]�|qx�nD~��tv���Sgܧ��S�lT j;p��4��8��G7���O@���O����O���7�S��U��!N~�Z�i2X���I䟨�I��MceN�|���P�V�|��љ�y*��S3�����F)�'�����iQ�u!�V���xt�D���L�L^a$R�)3 b����'���$�ĕ����'.2�'����#��(I�2����l2��'0rZ��hٴ,�,đ)Od�$�|�Տֆuxjћ�� Ojl���
y~�h�>���?yO>�OM�Ms �-)�n�c��8YH����d� �p�!�V���4�����qa�OJi�aK�"r\i�C�$]�N�@�O����O����O1��˓u��'B�i�e�$��2�aX~�U���'IBjq�6��ˬOZ�kظ�a����h-x�!4Z����O�0k��x���-f�) t����O�( ��$�
%y��+�L	����'H�I�L�I�X��ҟ\��o�d����� �_�7:��W�
,XP6�ڱu����O2��"���O�mz���Ԭlj�Q8E��RIʹ��П��	D�)�S�yL�Il�<i�A>Ô9хd�m?���ӪC�<�3L��TI|�D�����4�f��W&*���qnl��'�d�O��$�O�ʓb2�v�2?��'��+�f��J0�P�K�ćO��O@��'��'��'�\MSU �7qZ��gcE�f�D�r�O��KA�EH���@5����?5H�Or)&��?�t-@�.�6D��-R!��O����O
�d�OJ�}�;[�)B�@�v���4'z)���3<�f�����;�M3��wC�� ��2sL�s<�@��'�7��¦���4
n���ٴ����v�J���'d�-��H~�D��`�^�.แf;�ģ<ͧ�?���?!��?�I�9ܒH��м���be
����Dڦ����ky��'���c�Oڵ8g�;EM[0{~���d��{}��}�4o����Ş��!��\�<}��'��2+�@�ٶ+XS����'S�QbC��򟜣��|"\�X���ͽ!��=�h��!8�X��L}y��'R���]�,�۴���͓$�|�X�\�T���f�;��H͓S���DLP}RIl�,=n��M���? [��8`a�"�ql<��@޴��$A�Y�<��'��Ͽ�&b���v-�Aƀ*3j5XM��<��?����?�����ɀ%���Q�(��a1*�g'�Iʟ�ڴƦ��'y47m(���=`�\�cvd�6s���A��/
��'�T�ٴ���O�	�#�i�	�{�����-�+��q�$�L���O�"��Yw�Icy�OJ��'��#�9�޴��Ç+8<�+bN�L��'�	*�M�C��<����?/��4��Ɔ�-��Ÿ%�^9C��җ�0�O�o5�M�q�xʟ*ɠ�S�(<"g��-'�\�6M�\��ңu��i>�� �'��U'�4�ì7ybq�(_�{�z��V֟��	�x�	�b>�'C�6�M) �e�4�D����$F�i�Z�ۖ��O��D����?Z�4i�47x��!kVQm��j�J���@r��i6`7�B'�\6�*?��@�]i���<����BO1K��)J�&p�-���y�T�@����I՟����ėO�BB��S}�#��V�k����4�b���`b*�Ov���O���r���Ԧ�L ",Y���&ۖ�����j�@��d&�b>�*�f���S�? �h#7��u��5(��� �°�0O��!Ĉ��~��|]���	ԟ��pd��Ny�m�`��W�ʁb��]�����<��cy2/uӆ��j�O���O�e�PiԜM�Ts��� ��׃=�����d�OT��3�Dx�z�Q��:�pT���֪@D���ub2a2e�̦�PN~�t������i�ޡ�����0Dy���Б~=�!�����I��d�Io�O�"M��M�*A8C+,\t���� J��.tӐ@��OD�d榉�?�;zA�A���:v�(ᄏߒB����?q���?ar���Mk�O�N�C��S�g�0�7#[��T�H��S.l�� &���'�2�'b"�'�b�'�ʄ3"K�Hh��Ч[�w�z�õ^���ٴ6�����?����O���{%�έp��I�p�>C}�LS��>���?�K>�|�2�F�|��Œ0�Z&u[&(V�V�2��4nZ剰"ۚ�h��O&�OP�IV�����O9� ����2*��z��?���?	��|r-O��oZ�`3`Y�ɱ+�����Nֈ��t+<[��I�Mی��>���?1��S���˥e_2a&6٢1A�,
�|ծӸ�M#�O�(��������d�w{�����D<w8�:n�c���p�'�r�'�B�'U��'?�@}Ht�%(+�<q��(uȠ��s��O��d�O\\n1sw���ޟ�ڴ����%�q��|�9;����i �xrbb�>ulz>� ��Kܦ��'	��A����]��Ix��[,g�5��`�	,~��I�g��'�I�@�Iȟ �I�}�z�k@9v"���(/_�����͟4�'�7�������8�Im����Np
9�r#GX��E������J}�	qӲ�l����S��Lli$���lMD���ߌ�,d�T
t�8$�uP���!Rb�S�ɨ+�03�`�Z���X:�2T�I����	ɟ�)�Cy�nlӺ����58a�l�.PX(�� ʊLo����O��nZH�G��I��M�Qc�(~?�8�$nد��[Vj
8_7��g��i��q��|=�=�e.����,O:(§�޹��!�󫄻Z��['?O���?���?��?�����)�lX�(W�o�dAz-��n�lZ�w䨠������^�ퟠ����3ШD] �5@�&�~H��J ��i��O�OV����il�O��~Y`B�yJ���̡R�$GA'J-���i�Z�OB��?)��G� 2�J�A ���eԪS� �����?����?�-On\o��e  ���L�	(p�8�Y7�Y�e����2�� (�|��?�"T�d�Iɟ�'������H�PmJ�gK�w쭃��.?��l�"˪��4��ON�]���?�V�K�_.�9 @�#0i���?����?���h����PWȕ�bO(GL�!��E=t��T���Y��HIy��i�T��^�贂`,۝(Y�U���1��I3�M�0�i]�7-��r�h7-#?�"��Pg��I�G9L1�� �>�2k�*��/��XsL>A-O��O���O����O ���(��9+��Rg*��J$(Sg%�<�5�i��8��'�R�'���yb��1W�&	8e�!B4�`'Ծ7�,�
�& s���&�b>�[w��Fid����l�B�����<k��;?��	$�$�7�䓟򄊁}nq�QÃ�=-�|��e3(���ON���O��4��˓(�f�HWb㟴gA�"�D�A0�q��F4BAcӶ�4A�O�in��M�ѿif��f�@�f^��b�@X�kBz�C���g�����a��[����	��99'h�;h�0��6�"w�V�p4O�$�O�D�Ov�d�OD�?)��lT�r"��>T$+1�_3@^���OR�����9��By�}Ӹ�O���P���O0X�`m����V�L���M�ĳ����3��������@1l0�Q����A�����o��q�Ld��'\5'�p�����'B��'Eb�����IV�J�☪c����'o�V���ݴ\{�Ub��?	���i[�?$�<���ւX.-IBmJ�r�����D�O�6mKc�|�%�2-/|�J��	
ɘ��FAMP�)S �,�-��D�ן [R�|rFҶ0#���MҤlXhz�
�!yQB�'���'����U��0ݴ�,����(�"�طC2F����G(�?��W)�����N}��'�V�qvI�e�����A��N�+&�'�,���f��DGdY�#��d�~BFJ*���;F�ؒ7��'k�<�*O����O����O��$�O�˧d�8e	�[��\�HeJ+~�:��i1��#��'��'��O�R'g���
�r2�1g�����"ȎS,���O�O1��4��z���"J�p=�֏�R� �P��B���I�h�x�)��'?��%�������'윈EM�1� "gC_̞��6�'���' �]����4�@����?y��{e��"sn��@'�ds����B<�F�>!���?QL>��������B#31x<S��t~��F<f6��G���ߘO%���	�_UB��
$�@�p�]����Q�ZQr�'���'���ݟYƉ93�ˡ`@9H�ժ�ARҟ��ڴh�D8��?ᐽi��O�N�wu���SM�"辸x����<I��?���0�
)c�4��$��_���R��ru
��D�o)�:7�
J�X��Ɖ0�$�<ͧ�?i��?���?�G�Zt�P@@ �<�\]CA���̦��bȚ؟��IΟ4$?���8fkvA���"Ep9qc�2����O��d�O�O1���2� ���c׍v���"ō/)g���ǎ�U�	_�(c�'���&�4�'�t�Ői�����E�i�F�'I��'�����tW�D�ݴ4L�l���#�����͐��������2�Uț��d�v}��'�"�'(Y�7+�7���6�݇	=�xt��g+�6���8P��F�������A��Dֳ@��ؔ�Z�E�mQe5Of��O��$�O���O��?��C@̏1UL=pu��>6
�9�*�ܟ��������4@��ͧ�?�»i��'�V���͒�r���$˕u��Y��|"�'��O�^ݑ��i��I�U�d#���o4r�r��:����#�Բb?�#�o�Isy�OJ�'��&2L��� T�;�\��	�B2�'�I�Mۄ�J�<���?�)�l�!!H�.@�#w�|(@ ��X	�O�l���M�g�xʟ�d�ߜ(�R\Q�ex ��&�L�K��Qjӕ2�i>�Z��'
d�'���t��	� m0�_���a���I�����ϟ|���b>!�'�P7��:Qy�Djv�
�sʼ��S�J������8p�4��'W��N)�V�@����Z+Z��a��`ӧI6��h��Цe�'�M�4�Z�?]����qV  �/�~e��ʀ�4�*)؂7Oʓ��=��X3l��CF��3)~-R�
�vn�f�tb�'�r�i����@]�H�6ʞ�0�i�6LP����%�b>u�̦-͓8D켒�^G��q�فj��͓x 4e0�ﾟ%��'E�'��I��hS�Q�|EZ�l��d*&�'�b�'�B[�z�4O-r�`��?����X	!Ԯ�9[�Y�AA<Y��Y+����>!��?)J>��ǒ7a:d�@-�V���F	n~Z0ۺ��V���Oɸ����j�b⛒R�X���h�z�D���ɺh=��'���' ��ɟ�ZЩ��v*���T�_#������t��4GP��'�26;�i�}����&�h���k��>MмH%,h�l�ش��օoӊ1��'h���-|2��J�����3U����HD��ũSFK�h��O���|B���?1���?���/�v�1ԈJ�C��CwC�?���(O��n7{���ğ<�	a�s�\�D18^LS��F��Y������dRʦ�xܴW���O�:A�Q`Q-�>P�ņ=~�����C(�	��O$�y�m ��?ipc7���<���_jҥ�C�C�=���$ؓ�?����?���?ͧ��������i��S��]ƽ���V}�����f��Iݴ��'1v�Z��f�f��-oگ]�9b��DZ,�sA�L�w�,�g���I�'���$I��?e�}��;e�ʽ�����7��Z�g� R�Γ�?���?����?i���O�A�����f�Ed��f�����'X�'�F7픐s��S��M�N>��b�!��"�fS���ӱE�=*�'��7M_֦�7a.�oD~B��+xbqkw.å[bi�ӥS�Z�2h�ƥ���`��|�U�D�	���ß���l�>�܃g@ˏE �,H��۟8��yyR�w�H ���O��d�O��Rt�'� g���rCG�`��	��8�Iv�)JVˍ5�N��6�T�g��Fe��e�|X��%��;X!��t��B�|�j�/m >d����Y�!�.�2���'�R�'����W��;ش}`��5�Ш~PB����&��iY5e՛��d���=�?�Q�,�ڴ y^�Z Kр@��*��C�
x��i`7M:9�7�+?1 �� T��.��+G��DPꥤ��y�´�(���y�X�X��韘�	�L�	��d�O޴��0��!g;�v�r)ae� k��7m���p�D�O��D;�9O�lz�!TD^ز�VJFIl�A��"�?ٴE�ɧ�'+��9i�4�y�Z�l媜)3��X�Lܭ�y�ʴ2ψ��I���'��i>e�	G~Z�j  1p[(�;���)K6}���|������'�r6�*`�˓�?�t�R)~4�`	�m���	�ʚ&��'�~˓�?�޴�'G̐H���^���pb���U��i�Ox��Q!�N1I�R �?���Od�[�c^iݱ@$A�q��!
���O��$�O&�d�OP�}���	�y�ćS�\�� #�/cX\@��jH��Gc剘�M���wt:6E]�c�yQa��i2����'��i>n7�O<7R7M5?�qٴ�P��ұD_�$&��ژ�� �af.�AL>1-O���Oz�$�O����O쉸C`
RR}�r��=6��m`�μ<9��i�4 x��'�"�'��O�R�,7�FeK��HB0���B�?}�$��?���S�'>���!p�ړ1�v�*�D�?TE@``Ʈ�M�R���@,<L�a��J~΢�P%�8���i�e����a"+"GU8]�f�	�t}�t�*0�:q�Ѣ`�����J�(�:�p1-�5h�1;��º_(.8y/�ǟ,Ζ�>R��j_?u���g�.�I0]�*�qTꜯSj�h���:l̼s�.�I����!�}1r!gD�pt��S�J=�	q_'^�)�� G$�\�@>$e����$�21`1eC#\�U�"�ON$�F����A�5s* ���4gx��q�:���2���i.�����,��YR�+�v ��E�(��a���l��CV�L�B6��<�����OB���O�Ģ`l�O�[`��#��Y���;W�}j�,B]}��'%2�'��0r��[��(�$��Br`���� '�:E	���$%�rYm�8$���I��J���gܓJ��
3@����j�+=u��n��4�Iay�L�Ib���?Q��RU�ަJ4d�[����\��\@è���'���'z�P�G�Ĥ?� PY2W(H�I�hʦ��m�����i��I
�J�s۴�?��y�'m�i�-��N�/������%?���)�
q���d�O��Cd�O^�O��>%y��ك#�NE� I]�l��4b�nӞ@�bD 馱���@��?);�O|�g��%1��2t��%ˑ�8a��h��i��T8���$�SǟLH�IОFK�=�2b#[߀�	B˛��M���?i�'_�}�a^�8�'��O�CEN1�N�p�J@(����i��'Ȇ��G	<���O0���O�Pa�S�kO����nޫ[!bT@ek\�q�^���`�O���?�H>��J��0�J��*��C7�� �J��'@�#��|2�'\"�'<��8ϴm�R�ńXŠp�A�_�u�8�diۤ��$�<9����?1����R��J� H���R�O�Z�< vhֹ���?	��?(Oj|���|���	�.����ː�Sf�1�c	��!�'��|��'�֢^��T�d�����ȅo��mRNJ�E���ğ���ן(�'��|�p��~r�d�X!iq��F��q��}�����i�|b�'�ҌX:qO���fd��,xl8 B&����M+���?�*ON=�q�|����y�'Jk T�@�	n��U.Ѿ~�1{��x��'����:.�O�S�`�T�@�i��_���:S�5&�6��<�����c�6��~������X#�ϕ�zw00S���2 <�V��M�/O���O:8'>��O6��;t��$:0j��L%����!ݛ���i�R�'C��O'FO�)�n^�A��ėdS2E�@�Yo�ƁmZ
n��-���8�'�����ڑ4ۘ@�-;.׬��$��2�o���I��w� Cyʟ��'a���B]!>���`�3`&��I"�I$r��9����'<��Ց�0HN�hb$-RV*���'!B�kfP��R���⟠��F�-�	צJ4L&	�����g��'�B�'2T��z�Z&T�~DѲeÙbX�4 .4~���YM<I���?�����O ��2K�b<@si�.y�:��4�����7-�Ot��?����?�-OTaÇ��|2A���7܈�0MޤB1�Px���x}��'���|�V�|R�IܟD�%iI @�xv��T0t�I0�U>��$�O"�d�O�˓"Ѱ���T�,_,�h�F�[s6����Q�b6��O��D�<���?�ˍ��?�I?9���7��$J��C!=�tGw�F���<���?{zUq+�����On��Ƹ��樏U�(��e�t� �xR�'b��'��y��X�C���Y:��Pe���T	0�( ]�������X��՟Ȕ'��tY���P��h8r��2�X�p�^�T�d7��O,�d�$0%f��)��j�<P;nR�yM��𤃓3����K�jHr�'��'���T��'j�*lq� �6a|3v!G���MAйi�<���c������d$���e�b��S��āY�nC˦���Ꞔ���P8�i���i=}"�P&З`�lD̉R1+N,q=�b��ȴ���'�?����?a��յe�L8[��	)Ά bch�~���'���I���>�/O4�$�<���cF�ŬpH��SC�ǭl羉�E������2;�����8��ş�IޟX�'� |B��̡�jś�TT��+�%�ꓤ�$�Ol��?���?9�'	xx�׮�2/� �"TC�^����$�O��D�O��(��qp�<�΁��	��6@�E��(΀}�R1鵱i��	Ɵ��'���'r*��y򭓭^0��RC�=\y�Yi-
�5\���?���?�*O�EJ�+�w�T�'_0�x�� @ s���Gh H��}���d�<1���?��[p\�ϓ��i2����I�ـ��[�:�Y�4�?	����d�����O<B�'3�4B�N"�i�A��%Hu�k�R�<����?����?�i��<1���?���]���`�ٗL���$q� ʓ} `�r�i[��'���O��Ӻ;�h�=
G�|�uM֬@,����Ԧ��	ޟ��A�m��	jy�I/��
A�K��;F,�'6�v��C�&6��O����ON��	D}r\���aO3>��(H4��S |m�Enޢ�M�"��<Q����9�S��S$����R��X�-sR���M����?!��m���6^���'�R�OxLj�Ň<#�,#te�z��ҡ�ih�W��R�@w���?q���?a�L�i�>�	b��#8��c�%��1_�&�'��h��k�>Y+O ���<Q����֌71�U���P6`���Ċh}Ҁ��yr�'���'A��'f�	@���a���Z�(,�󦗆 �������d�<)����D�O6���O�0�eڏ3�r�i�R�h�����_�$�O$�$�OV��O`��1A5�X�2�n�:I�x�����0��)�i����ȕ'�B�'��nZ1�yr.��8T�P�B�j�p�F�#$��7M�O0�$�O����<�CJ�AK�S���P��.[��l��`W�o��C���M����d�O���Od�i48O��禍r�7O*@a��X�ȀU"%�{�F�D�O�ʓ5o�ygR?��I�l�Ӆ?�"@E�.YWҩ��&Q��X�Ov�d�O2��4&����'�f �gӟ#�(�W�V� �fem�Ly�+O*"|,7��Ot�D�O��Pe}Zw\��&��;g���E�شGR$��4�?�C�B���?1,O��>����O9t���Y)���Gք�M+�LW� x���'�"�'���k�>�-Oh�yPA�^�L͂:7����������{���	Uy���O�8� ���!I��+vPc�4v������i��'����>�V듫��O����`��j` *~��u8ӈ�"6o�6-�O�-�D�S���'��'����J5��!��Bk�0l��`l���dÒK2l]�'�ޟ��'Zc�����NM�C��÷�۫|�Ұ3�OF�6OT���O����O��d�<14��/m���Ҁ����+�H����V�ؔ'h�^���Iϟ����T!0��gC
;6eh7�mXi���w���	Ɵ\��۟0��Ny�+́E�~��y��sG���Rz��*V�ץ!8"6-�<�����O*�D�O8�h63O�$�c@�����MR�3�H���æ���ߟ��Iܟ�'��=٦G�~z�x<Y଎�73���7�C�O��[��ij�W�������	���A�D�c��$�~�3&�H&(�n��|�	xyZW��� L|
���vͦ%��E:��^�<�Ͳ��R�
l��џ���͟��.�ҟ%�P�����g��9~���a�hQ o�\pm�|y�e)F^6MW��'��d* ?i"j��vꞍKS�ô9�
��aC�ɦI�����"B�&�t�����,m�ʄڱ�Si�$��6.�4k�v\P�07-�O����O~���f��ȟx��h�,%^%@�I�6Yj�P��J;�M���];�?�N>ً���'G��B5ׄdDH	%m��xxn�b��tӶ���O��*Y�$�&�L�I����eJ.�Pb�"c���n8��oZE�Qg�HqO|R��?1�'��L"*vP����.���c�iV���, ��b����`�i�-�qn!�z4XB�Ń~WI��J�>qb@�<�*O���Ox��R�f�8K�<�;��^L���VH[*l&�'� ���&�$���\1F)9�|��V�v��$dđ)Z���Wy"�'���DJ�P�S�;pP�:�A�
I a��ɋ�Z�듅?A����?I��Df�%Γ;(��AV��Cg��(t��W���Iӟ|��Vy������i"a��1p����ޡl?�Mx��Gͦ}�IJ�	ϟx��
����=Y�j5�����苞H�
�{Q��Ȧi���x�'��b5�:�)�O��i�+V�����{HQc!L�mլa$���	؟\�T(Bꟼ'�\�'O��,�Q�
��Α �!�/BIl�_y �Dp6�D��'���k'?�E��?g0%��G�i��)S�ڦU���4s�,��'���O��D�1:܌�����(�D�Q GEV���&9$�7��O�D�O&�����͟���"ޢ6�t�dH�i,,�2�!	��M��m̀�?�N>Q����'��,���hv ���%00A��p� �$�O���M���&��K�P'�
��4&C�Y$A���%*����'��	�>��L|���?����ԩSP��qr,21%�1*|~,��i�j�EΠO�i=�T#�2�M�!��<1$ ��R7���'�|�[�'��I�l�	ԟ��'� (����<$'NP�d	�=
��)%�B�XdHO�d*��?�6]�����Ǡv���Tm�J �y���?i��?i���?.O"�a���|$)T.~�zE��.Q��H�u}��'�ў����5�Q���\��У�h@�v�Z\xm��*	2ٰ�O&�D�O��<i�%��O��5��'^�h��)V[�\@8�5�d�z�=���V�݃����OxT,�FF��#S����BB�$H6M�O��D�OX��I,D�����O����O��	�
����55P��J��K{�E$�8�I�����n��dc��'R��]��/�(��2m֘E`�aoyyR"�hx�6��O���O��	�X}ZcMx��Ț$Q^�|:c)S�4�u�M<�������'����>�B�m�:A9!�;��B��]�QIƢ��0�	ҟ��	�?��'L�S.Z��Ӧ�*
&��ϟ�E�b�ܴpH���.[\�S�O\BK�e�n�hu�Ȼ	�a���Gؤ6m�O��D�O6X)�DԦi�IΟ ��ޟ��i����YW8�$:4hˠ0�֥ `A}���O ��3O����IJ
b�0g�TؒP	���B��A�Ɍ{�h�@�4�?a���?��H��t?���%;���1G�X<?���Cn}�b��y�T����ٟ��ҟt�I�>��8bu�	�o&X��l�)�t������MK���?���?1�Z?1�'}�Q�|.�hS����n���ؑA4�D��'��' ��'n�Q�$��G�����شBP����/G*.�&�
P�Ŵ�M�.O��$�<���?I��)�����-ՒO�&�C�.9ul�������	ȟH��ݟ��꟨)�*���M����?	�ě�?��l����b�Z�[V�UU���'B�'4��ǟT��c>���j?�L[�b(`S4Ş>c~�6&��)�I՟���ϟ�9.��M����?���RB�Mt�I���A(� �2ě��'��	ٟ�h�dk>y�����Mk
��B&@)4.�Ur ��q�����ğL�hN�M���?����
�'�?����\�A��,�!9���2.]=��	�� �������ny�O��'O�Ȱ2%��i1�6��'�h�n�@	��"�4�?1���?��'%��{yCF
fhMk�c��!� ���b�'v`7�,�$�OPʓ���Q!ӡb%�bQ��[ 퐢㗆g�.�Ɠ��-I�����a�*^RI���	Tp4���9��`��b8�oE�hH�sP+YM���P��<���.���T.�,��5H����i�݁�g��v���jdJ�4��Š��C��hQ``�]�L���-_p�Fdj���!mX�Z�4�C����n4�!�$�f�;� ��� u�I��Z�u���2���Ol���O��I8)����O
�SB�Z�� C�	��tlX�fD�M$^�T��R硇�{�Z�k���Oj�GJ!R�\3�$
K �D�ĦY�7	�0��D�
)P���F$rDmG~�ќ�?��U��i��#�"o$*l����W�N،�3��]6�^�M�f�:2S'�Hp�ȓw�rlx���8^,Q
�Nm�\�H��Ify��9.� ��?�,�^"����)t��T������똇\N���i5���d��\s��Y2˖�����O�S�^����H�� Y�-ʡ'���<�p�i�Pi���Y�<� �`M|�cI�CV<�;D�6BR����q�'̪���?���t��F#.��E.�<������
�yR�'���df]Y��5pV�
O�DHk���'i|\��_���E���DD~X�'����I�>����I�V����O�d�(�64XC��z�CBh�_r��H��T���ˢ�Jt��|:���v��y�VC�@@T�ⰣOq�$a(�*YZX�sgBѾ>U8tad����"�֬G�Ps�gC�%�Xy���qbb�z��'Mr����&�O��� b��Peܵ�`�������"O�����N1	���U-gN�c�	��HO�SZ�t��d�}�Rܻ�fעo�~m������R�O�3�v)��П�����Գ[w���'�jMsꁟ����� �81��J�O�D��486��b�������::r�=3��&?M��PcG%4\0���9x���!�%>^�s�՟%��l���'��j��Ae�"��@�F���'
�(�����=�f�T(^0�
E��Z����S�<�B���4;���r�<m�P	Inґ�"~Γ��kc��� ��q�&�8 �ȓ�88��)K�B��J96�������d�Ԭ;��d��2�z$�ȓF�3"��!I�4�`R�b�=��dk��1�CC,1O�|��E�
���P܎�h�h�j^Mb��ͷf�*��ȓ+�,�҅D8'��l����&��1�ȓ���Yc�F�Nz(qq�U|���}V��{���6XzQ r�JM6	��#�����HI �Z`gS���ȓ!#.T���e��@��?H����DCԹ�S&#�` ��>o�8\��N�}x�	�$R ��S��"{T���J����7B�l��U3PB�7o����_X��rǫ��Y3��jF�@h���h��L��%V����$�U&����2TgW�8����L��f�ȓ��Y!�BJ/�lj⠞*x��ȓ���B���$��{�Ĕ>n�dt�ȓ`�8�`�\�U58�3�⛞T)⩄� >xR����Np��p%�0+���/���Z/r��«�T/�m�ȓ�Ń!�FV$N�`3o�r�$��3<�Pjw�\?v��pD�E�<���A�+�vP��X�V��%�O~�<tA_��АېN�T�p�2�z�<QmISj�iE�����!���A�<)V��A��}r$Z�`o<���z�<�`���Y�̑
FH�?l�I;��Ey�<�TI�Y7���%�Ua�ʖ��o�<��VxD��T(�?�q�t��n�<aK�i���\>ODL�9�g�<��˙�#>D��	����G�a�<!���ݸa�EG�8R�8i��_�'�H �Q�4��OP,yspΔ�6��i�W����UZ�'w�����#�vLS�kH��f���'��<�5c��YKɧh���OH�%���	6�C����"O����D5D*�{�M��/b��4�>1w��.;W�˓l�R��aA�a��e��? Hه�	
V���
�^3�8HP�Y�Ԥ�=v��e�ē����v-֢r���aTbԱ?�D(F}rl�i�rj'�� 
-�JPy��P�Q�g��iQ�"O��S�ДNٲ��ɧI�J��O�T�M\�d@1O�>�rpJ
;%˖�طm�����fH-D������Ai\,)1T�Yt��A��7D����֍3*8�ҹo�حu�*D����8(BP��Q���I)`�5D��H�C�|X��/q���ȴc>D������#U��r���	{Ѻq��E>D�$
DgB�F�kw��]���x�K:D�$��(\{Wb9����bC�ԙv�;D��Jv��3[���s��aѪ|{a";D��ڄ��2q�P�Y�F�P^p��$�;D�4ÉSKZY)���)z�6X�CH9D� �%���'Ϭ����w�����a8D�x� E]�`J �B���:.T��"8D�P ���.I�l ���_; �q⦯(D�����|1a$nʚ)r��U�$D���c���J��aG�@�l8�?D�T8S/͹l^�j&�E�/ʜD1�<D�,�6M�K���c��ǎp(��&D�ps�Ě!@�:���8r���):D���!�MCl�(ӣk5C-J��Q,+D�l�E��nL놌��f�[��>D��h���[��� �/��m��ۀA;D�вKЊ6Bfls���/y�VU�!�8D������m8@	�&@�]O��Ib##D�d�S���Q�$A m��!t#D��qTBBEn�񶀞(�4��$ D�|��'��"��qj�엄��f�(D�t�poC:3�`��I"�:���1D����
V+_yt��	@���F(1D��*P��]��;�(�.[�0��-D��Q��LXs�	�a�u��H��H*D�8x%i���̚�(H2*Rx��,D��q��k�$�!�N�QS<�� +D�HP�͘
V�\JƊ��oE�ڶ,,D��8q�;]
��B��!�̹�!O(D�l�'J��7�x�XW N�-�ܸ+#�#D�Pj���'G��D8��͇B����i>D�83h�8$��E$˳,B��r4=D�\�������8פ�6�6D����` <-�\m��O=�pi�N/D�`rg@�y r,��GO��IR�//D�$�A
�A�:9�t���$���- D�t[f��}hi��m�!'sP���2D������2K5�(p�UWSpEɷ�5D�����7�N�"5H�QO$�Ȗf2D��Af��>�a��
�����*}�"5X��6�8.��?�` �B>`������Ҭ$�6#D�,�c��KZe�GK�${��0:�
�n�&�'촐��\��Ϙ'�������{18,����vGȡ;�' ���^#4������0pc�p�B P@ �4@��N)<F�3.��0=	��#V>����L�}��j\���ޏp��E�s䚥7�`����� y��ȁ�f
V��h)��ܙ���Ɠ4�B�RA�^�_�����U8��H�'Q~X���[/7!��0�)T�p�Q��t��P��@���f1��x�%\�lb�q��X�x�bf��4��� $N�J)������MPv��R���� ��B�S�Y$�'HHiWo«r\���N�o6p��N���fUS���G�
%L�[֪��wuV2�S4���VΌ�m�󄗰���yD��"Q�@X���_�8Y���
�f�*���J�G<����G@� _h�)�!%e��J�$ߖRZ���Oƀ���Q��тΛe�d!x]�� phH�v�^-�#��@	�҉�ئ�?��λ� hѠI�6#���I�8D�8�� ̹!#"�4|��o���@�4n��?A��P8F�x@N>� ��H��ΗfK������ ��C�'��J��ºm��:@L= *
�Z ��:Pߨ��@R�c� ��ȉE�����C�� I�I+��X"�l��m�ax�X27�zXJ��
���lH�)@�:>�#�O�&��K�*ТOpJ���O�92OÝJ*4�zr��9"��0���hj��B��P̔�UÎ��t��j�O�R�Y��Ȋ!�d��C�8����')ҭ�B� �s��*sAO<�<d;P�F,ay3)�v������S��?�F���y�CܭB6.�Qr���b����!Ƥ��O
غ�N�b��'bnxG%��o�D �CS�yJ��ԏ7ԛ���*D�x@�GX0�0=!Ṙy^�YB )Ȯs�~��fkUM?�6��:�q��/2Yl�S�t��-6Q|��Ŭ�-3hA�Uaʻ���#����U�"O,I�C��;3��0�C��?�vH`dɂ�y�@ ?�@ȓ��09�N��]�zi���.I,�"+�L2tE4w�ԁc�?%�����RxX�$�/&8�C��. ��]p6��<kb�I,n; �s��0Ks����Y'v��	I�P�5��/�����$˪o��D|��!J9��Z��<�e���yB�P7�Sg��*}ܼ��n��;t��qKP5l��c��[��0�bK��&cRز�Ks3���SFi��j6.�m[��33+�}�bC#��2FқVR�]@���S�F�X.�������D�;&z�#DlK�~�r�3L�f�$�a�D�O�!��v}r�b3n�,Mf�ݿ�FD��lϦJܘ��WEF��^����#5��<�2ʐ�,n�¶���)?��#�V^��ɞN��@4�xT0 .��?��i�/��/�왳ᒽ.���jSl�:FȢMDy�$�$ob�훷邝n��hWd�H��	/8ՐM�V�� �RrVgʢ��W�,�X�U#� '����$͇e.�B�M�<T����j�Uk�}Zr��
_�A��\,1.6�R��'R�4{�E��Q7j8�c�ƄM�"O���ʍ5/8p��#[�>�nl�@��q*�x�-��,M��������%��!}	>4q�䝄n�Pт�x�t�̐�V��ȐG�06d ����9%v��%�O������/�̈́�#�4l��(�G�%�ݩ<���R��߂E���i�A�
��(;D���PH����E$h��h3?1F�?|B-��$��G��h*A��c�A��/Ăk�{�'����<!�Kα)��-��e�3N��S2>��V�͒zڦ9�3�ԉ� 1���be"l��-Cr�0CTC!��Ɠ2Tx�	uC�_�����m*�}��FG`	pg�U|����+� �ص�lS;m�h!1����������4��MB,�S�&�jr�K@i�:%�a� Kѧ�"�ؑDvP�W��M2|E&���O!jpD�\m l2$��(*(�`�j�)�d� �F�t����"1O��&��N 88P0g�,X� ���.������jT�����M"Q\Ua���-����B�Z�X�%��E5z��G{�f��hn���7������V����+[T!�dM�>���e�m�����}�ў�ANC�O碅�aN�[���ah���s2! �7R��G�~���7�1LO΁!��Bqd���`��I��e��`�e5�5�2�G�VPL����'���RR+M�h|j��N��d���$0>,���&W�^�D��1O^�@�>R?b QT�ӂ|1�lp��$#|�8��d)"x��)h�˅)-[�0�c��:�p?�ҫg�l�+&�&}1��B�3a_(�x��Ɯ�i���p�'B����4��`b�M')�F���="1��s�"O�M�IԵh�6i�1��.�n����ɿ0S�iq%���d�#e�[�[�&��()������Dw��LjE�H�U���$��&��t��
$�DH���D�,�f��IH��͂���?>�f�{��	�f�;����T��O<ɉ6�[F� ��%�Jʘ��s��W%L���bA_�uF@�0��=m1��򢌻"k
+#�Z`˦��6hXJ�z��k2��06�'P��R��I�5�4Y UԠp�M	w��7G�5 ���SA�?E��w�
�QW�&� �`�3H�}j�'��%���J�ך|�V��Y=�?!���u�p���eU���$��e�'Y(�[�Ƌ��r���� ;�L��(��$�lۍl�άb�#]�l1�$rL��>��X�f$�6�Ҕ�Y`G������r�Ї+V1��I�G������4i���P�G�~���@)�O�IN���!BV㍡1�p�ե��>!�բ�f��&+�i��I�F$Z,h�dF�+2����T�២|λ�/ 2n8�Bf+ޝw݈�������˱.��s��]Ք|�e!�.���d�gA��QE�wb���ƄX���j'�S2������7�!��j���;M#p7D��ϋ�'�!��O�X�aJ'�	�z,欨V�E+/!�� �P��|��u�@��h���"O +t��3H�E� �
]#"O(P� �WkZ�2��0�l���"O�e86��$�ST���|M��1 "O��I]�*5<!���x2A[�"O~���h����,*�&I�ލ��)D�8��S�Y�&]:�	�^���T�&D�aCC�&<��aNۡP��%�5E%D�`���W���b�V#"{޽�D�"D��Kd�K=�6�Y�j�m}r��d+D����BD;Bo��J��<w">�K��*D�HPskӾ9�=���φ _"EE#D�\!��2GA��2�BK~��#5�3D�x$Z�R��R��L�U���4D����"M�zr�<��ȋF���d�,D�l��Έ1_�ӕ�ɉJ!��ӂ�=D�L�o�*:��ˣ �.њ�C�(D���g	��Z}�,��.��%(D��Ð���ε�$!�(4��]�*OEOC-[�|Sf_�<5@�"OF�F�9J�6mr����t�"O.y�!�H�`��JT����x u"O�Th�F�1��� �BׅW�F��"OH����u�ʈ��*��%�<1v"Ofp⫉)�6��3O�$Ȋ���"O���!�Oܜ�H
7h���#"O
=�1�1tI�غpgw��xS�'D���pɉ�`?d����+F���`�B D��B�˾ ���ɸiC�Ҷm0D��B�I�6J��ZP��D鰨���.D� x7�5@옔���P�z�+D���Ӯ�gm@)Z�(�*�n0��'D���cK�-;-x��U.�Sml���	1D�e� %�B*��D"53����0D�Dc�X,�гS
Ɵ6�����8D�ܛV6y���p �!J,�8� *6D�,���T-]��3�!Q�/�D��Ն2D��r�* � (p����4z��<D����,B[��UB�I�� �ѭ'D�(�e��L��{DC	���3 �%D���׃C0f�t��f&�d&t0���#D�88���8][N��C��e
��ai,D��[��Ьy$���!k���2d8D�����
5"��X�DT�V��:��2D�px���6b� �rS�n ���0D�Dh� ��*�Q@L�}��o0D�4�V���J�kӏ�r�\}���:D��ر���u�xB��3^�2�7D�h��`��!���M�<�$��%5D�4�*�0�As�)�8a���3D�� ��
�/�Dm�dn�`�ّ�J&D�`qv�9�9"�A�7�I�W!0D�8qAd���}�hU	x�}��,D���',�#�l���@�{����)D�8#�/%�r���D_�ay&1s!�<D��B��E*l�� HcB©F��Kc<D�tq�-�0,VY�6��P�h�S�=D���"i�q*6]�2�%�~���<D��DM��S�`'�аk�F���'.D���%����JŁA�YB.��ю7D�\um\�'�N�J�����5D��{���)�nĚ֣�k��RV�&D�|k�� >���ťO��(�Q6!&D�D�3� �t �kN$������1D�� �����ޯ�Nx�P�^�Hj��"O(q���8z�rz��ܛ!N���"Or0!�*�/,��HԌ�^�v���"O��	+j�@rPP
r�&)��"O�I����g>P��91xlXC"OꀍN[~Z�JT C���u��"O^���í0�h�Q�^�fN���!"Oh���O�4_K�l˜e��'"O��XE�D t,�%�C-��r�"O@ ���Z�t� n�=`oF�[3"O�
����Iܚ�,KV�
�z�"O�� A��4�u�*q$�y�"O�q�D�<r�Zu�FT~DYw"O2bc`B<v�X$;�IcȌ��"O�!���M/#Y�xi�f�5�Ȅ��"O���3���S��4�P&S�p����t"O�hإ��U�F�6�
�{Y"X`�"O(�pH3,�R@ZD��A�xű�"Ot}j�k���l�V�<rz�4f"Or�����z�-k�B����P�$"O %�Z��(р+�5Y�Ĥ��M\�y��_���|��O	�O��`ϐ�y�FT4O�����V�}Nj�c�����y"�� 2~q��jF�rN�B����yrm�`��%�D� ��m��M�
�y���5N������z4akSO���y��?N\|��IM�
�EXSbџ�y�BфM�v�*�����9����y����ig��O���r"+�y2�Y1s���KQ���M���y�m�;K��,�ⅣD�S:/��1+�'tq����!7ݬ�{F�!P�,�'=�̡�*:x����^!����'�t�ç3;W��$�"PF��'l��pQ�$Qw�Q�f��K��i��'�(a�$��B2)v�ԯC[�h��'+x{7��F�4�+�a��&��Y��'&6XC�gɄ�Rt�P4$mHMA�'�y[�)oe�8�Z1���@�'b����J�Z<�]A�����R���'E��K^��4ev�ӯH����'I� ��"� �E����
���'Ǝ]�Wd��*[���Wx4Mi�'��H�cnB*i��Qcʀ^����
�'-&$�BJ�/ �Ԁ,�Hc��
�'�r�#2�R�d�@X�A�<?�}�	�'���RiÈ�Ԭ1�:��:�'�Rp"
 >g�*Ax%�4����
�'�L+�)X3>v��*� Z<.��U3
�'����T��;����3��z�>x�'^�I֡]�w�ҭ�RKֺ^�����'-�e���S&l|>=eD�*p���'zҵ����%^\�a@W8'T 8	�'��U[�-�*��b4���N!q�'� ��&�L)/`$@�#B˦e/���'p8eiƀ��?t�m
�fCW�v�	�':�P�@�G�
�'i� x�� H	�'0|d�� �=�.���������'���;폣x���Rį\��`���' ��#6G�;0j
��C�BҒ9��'ް�P0�̲!A���"	����
�'�Z`��&I(4&]@@	V��	�'�ĩ�B��e��Y��%.N͚�'E\�u
�F��� A�< ���� l�k�CA�<�c5ό���)�"O,Q:!�͜~fn����_0j��Z�"O"�H1,$e�#�Λ]�T�r0"O )C�B�)��))�L�_����"OP}��\$Qd���-υoth��'z��HV*�Z�ț9,��tQ���Pu�C�I<Y��|;�n�1A��ɺ�
)��C�	3|:`��'χ�H�So��C�ɒ�p��@I'a�`��Cµ:��C�ɡ7/���@N&rMP�8F�ñ	R�B�I����l� �Ϣ�X��'�<,�V$�,%�*E  b'#7Ni�
�'��4���/.�@x����) ]J>a�4,�HѫP0<�k6'V%�,���v�i��
c�ݺ��`��M��KLbp��3`'�L�UhK�����������'E�u�`ڱzpL���
�,0I�N��lJ�5@�dQ,�J��'�i!�׈>F^������]�ȓX� i�UM��b9�@��D��K,�����a���K?��b�f�&hR��ȓ �NHkrS	v��,` �λI�NB�	�sPD���W�T�5(��7#t,B�Ʌ*R)��i�%u,��� ��B�	�&��R%ŗ .8̨�M0�B��x�2�k�C�30iޱ��' �c��B�I6S�2�z6I��eqdU�n�=*�B�I�1��|+P)�	,S~d��JT��B�I�4�*	����<rQD@�Ǌ����d�`P�-:D�fY8� �ML��sJ7D���riF�;��AI`�.���J�n5D�@#&) �ԝ����X��@���3D��3��T;N��BDՙ�&p��3D�Ly�K4C�a����"1D���A���X�;�4h��٠�#D���Rd�t�0T�W�l���'>D���0%ܖ>X�
�	\�Nu��E<D�t b��P�^,K���5d��8D��sP��J�q�I�f�8 Z�(�y҃�:��c�M��8F���y���Yfc�o,{@n	�y��w�<�e)O�mo^�����y��I�P��s���]� �A)ݻ�y2�88l��O/&���)4 D���'y�z���qa`E�5��id����?ѐy�E�xYVT*�1E��|Bp+6D���D�>)8��pS&X�=��<*d"6D� r�N]�7��Q��J&���&4D����U�)��j�!E�%լ`q�(1D�l��`ՖF��J�E	a݄�E+D�L�R-�#<R�L�B�Į ]��Sbc=D�j���<*�r�xb�h9���W�9D�0IW���(�04Z0�B�Uc|X�2D�`���Y|� r�F�	C�!�$	1D��&��-��4J�Ćq��cm.D��`��ի)��<���)^��U�H,D�@�E������K/f���(k%D�<J�n؉)!D��Cb[;i����b�!D��c#!<bo�Y3���N��At�?D�l��R�<��=I�GF2"zy��'D�$8׫��A?0͊�i�	l�@�Ǭ$D��B�(=A�wB@����	5D��*�Q�y6�K�K�ĘP)-D���E
*rH�a���O -�H��@%D�� LzE�N;(�T�3投o��͢�"O�s� � (�Z��ɫm�$Y��"O�%Z�G��$���2�	8q�R9��"O8�� π�2��E�1et��"O"q���1�:iɢC_��� �"OB�i�Jزs�p�uț>HR��"Oְ��Ɋ8[>�Ӥ�7s�^iS�"O���Fi=J��X#��Y���(�"O�h`#��6V<a��rV���"O��s��]�M4.X+�@�G�E�c"O���F��RA*1���W�!��"OT��1ϒ 6�zUa# �u�"O�y�4�0	 ������k���W"O2����$le� �7�D��PT"OPJ$�P((�paal�;I�xT��"O��a���ZC�#�$�)S���I "O�1�*>7�jU�2��)Cy�@�B"O�3Eݳ^�~I����!�X��"O`��ڻOZ�X��HV�o����"O�p�"��Vhy#'�A�O�d���"O�A¦��F�X�zB�Ŀ�|�c"O$�8�`ڲ`Zv@s�Q�YR*Hu"Oh-��{lx�3�ͨq"~\BB"O\h�JH�wA�p	�e��c����""O� eo��M�X�r�Ԃ>P�"O�|����j�땉�P(z�"O�E��=��`K&Ґ��"OB� V��g5R!�匓dZ�ĳ"OP�j�B�0�2\�cڅS�%��"Oܸ�s���|y�C�RJ<�"O��s�1�j'X66�`�1D�Ԃ�(-[RtD�W�p&��U�9D� �ؑ2�cG�5#F�Q�g";D�t;��
yf͹�`�+l>�Ѫg�6D�`Q!���e)��K�C�U ��9�K4D�L9QO�v�44�tC�,mV�	Ơ$D��Ip��
����#V��h��v=D��1��%���a�^f�+t	:D��Kq�W�#a��Հ��>慒e%7D��`�ԯJ6��P��d���F�4D��PĤ��6|$ZM[�I�Y��'D��q���&lo~��:a\(���)D����NޏV���@�	��Vر�4D��c!Ս}x�+�D�~)�.D��2PK��]��(�c��O�ލ-D�9��O�hv���v��]X�3P�&D�4�5\<A�p�{�J��G��p�P1D��ZF�ǬRp�e���*6�zUK/D��ba�U(	��m�Wj�!R<�q�K-D������0{����`%�3w��1�5�-D�5��e!x\�����ax��-D�h�3�H)�0�v�Æ`�"V*,D��(Q���V9�  D>L&=Q�c&D���U�àeP	i����,�D[0F#D��"�j)^�$�@��.<}f��, D��YU�٣0�ʅ��̓N(�2�>D��hr�Q�Q�DI�@"0Rn����:D��Y@�B'�s�09	��8D��A� ������3_1F�Vu:�(3D�0sE�P�V �	"&Ș���I�D2D��Q@K�<e���C;[w�};P�0D�DK��)4����L�s�*)�b0D�ذV��/nȽ��Q�T�"ъ(+D��çb���G�P#T��U�C�&D�� �P�c����G� �:أ�"OJ��މm��d���]v�Hi��"OV�E�	J`�h��ON�{�����"Op�� �D)���sS�Ԑ(�&Ļ�"Oh��%V?E��P;de�Q��C"Oृ�H \��P�q&5�:�ʓ"O$����/VM�D��c��h�S"O6iC&$T�NID�i0�ԏQ��X�	�'���b�]�J�Qb��W�_��
�'9��A�gO;:8��ދ��Y�'����c��+�m�b"��~�$Z�'���Mԋq���' L���
�'��h&E8��M�'J; �K
�'P��G�_�c��-�fJ��`@�L����=�J�.4DI��^ ��Ʌ�F����3s�B�ؗ�X[��8��'�lt2�!B�Sb��L} ���96�0c&ҧuP��!��QmK"D�,`��)w��F�H��(L8D�\�3�E�>8b���@ߐ"�Hڗ!!D�D@�Ǆ�B�X����V���d�)D��⦢�m�J�8P��Q�%�&�$D��Y�eA$f��t� �M�kO����4D��
!�ɵr��)	���,�b�)�-D�T����l��5cް!N��2�(D�$1#��-e>µ`'�F� D�g3D����h��Z�P�tŐ�kz�� &*0D���gωe>*�BCȍ�Qa�e�� D��@(W�C��L��+9v �q���>D�\�B�0v��d���D�P`Z�0D�xp�F�*T�8Qą֔>�e�-D�\�6C��C1����,I�� ��&d8D�lp����M��5��L�c��XY0A3D�����n�d��e�ʪhR����E;D� 0�`
���1	jܥ�X\i%�3D��Q���3a/ �h��]�B@aK<D�����A6�����Y8 CD�j��;D���d��`.����Y4
�b��6D���AНa0��IE�	(l-J�фf)D�x����h�@$ ң�	s�R =D�@YF��3\* �[�hE=Bb��b&�;D�<B�JV�,����n�H�d��I&D����8!��8"T�*����"D�x"�֑Mֆ�{�L����.D��'(f�P��B�&b`��,D���H��
P#jN_�v8�)D�<&��_�����	S�A��(#D� Ʉ#r���0��L�t:PX�&/D�����?�$Ջbˈ\���j2D��9�o	�_�Z(�^��� �N/D�l�@O�$Lz�XզݠMn����.D��ԁ�*<�])cb�1x�x��S�+D��h+�v���0�^;>���f7D������BÚ�Ca�]�<:��:á3D�4
�LH�G��8���-���ڡ�/D�\@�狴&��}[EA��8
� � �.D�� !�=(���{�C�$h
d@`�j)D������Pm�I��F�n���c�%D�(P�FQ�K@b�TA����Qc�#D�@�j���Ͱ�e�|���x�>D��bC�Ǔ@��I��I+��ؠ��;D�4�!dFɣ�G	._��49n:D�$����,���7fF?3+�(UL-D� �O# ����dQ�<b!�� ,|����c�"�� �[�<![�"O�<�b%��/ĆY�Ь��P�Q"O��	�'���� Ǧ��|���"O>��Aq �P�O��J�z�"O�X��>�uH5� |����"OU�`�Q���Q� ŤaeX���"OV� ���>�Js�ƁU]m�s"O�����4u�l�RwNK�qK�9�"O:���A�5S�����OJ�ɗ"O���Wk��7�b��UM�=|��"O&���@!N?
�"��R�)��K�"O�0�\�Uz`��@*/p���"O�I�5���-Xz=yP+03���#"Ox4�ǯӂhz�#����*̨�*OT�Q�@�B|y��K�����'﮹WN΂(\�m���O)AP��S�'&谱�M�z�z͢��J5�H8s�'�t ��*ً5+a�f �c�!!D��9!���W@JQ�š����;�O=D� kse�B��*���aF�qr3!D�r�\��4m�s�ط]8ty3�,D��3H�)Q��8�,ՠۜ]�H+D�D�A��*|�2'd,�@��B@)D��;�i�M�MI!(�D�x�"D��[F��T��Q�ԯ�Vu�m���+D�xk� ��	<ɓ$*��9����,*D�x"���&13��x�e^�r�l�s�*D����V!�d��6[	˔tK�D&D���R�f�P�$:/����o"D��RBo�,0^DArO�z�����;D����$'^��˕�>�x{��'|Oc���k^<t�i��b�k�tp)g
2D�����W
�~�S��(#�Z8p�5D����̍3ƆPbt�I���
��>D�����i��j�W�ve�v��<�.O����,V�I��͇g �:U"$!�������l�le`dX�kN;k!�d5l�¡d$��kDd���N�!��.W\K�"Ó*Bv�g�%oў��ቄtƪ��o�L�|��4���C��	t�rB���<� �HC"W�f�C�:`�H�7��j����k�P �C�I�FLn��UDKb��ly#ʉ�O�pC�	lNhpq��O:���*�AFS@lC�	r��*��u�D|��C#[�B䉆Q�t)y!���s�@�J����DB��q}���lȽ[�Pt����9�b��D/?�&h3*���0�	c�ȁ@��^H�<�I ���fɟ�����,A�IQ���OuTT�a`�6Px�� BQvCR���'f��:ՠ^�M/�8`H&pZ���'oHy�V�҄[�����a���'5�cW�T,���ǋV�����'ּC��V;� ��J��9l��h��?��yҮ�sk<B���:��@3
��yBb� أ�,�u�4]�S`��'gaz�!��(&�]z6.Ui��`�u	��y�-Ӌ!�v]�4� e�BL{���yDF0�X\HǇ2����(0�y��ޟ=��T�ń�/C~�s�Q!�yB�.4�DcjҎX�}���ޅ�hO��O��O���7�G�w�Ҽ��*_�W
���8D���H�"���

@��SRJ!D����ʈ�xTz���)�-�p;_�y
� 6Q&"�$6���f�QxI���"O����$UN���7*E ]ո�"O"���k�E�08{7G�.2K��'5�'�az��I;9q.%�"��+�BIX�LM�?��R�s��y��F�|p#F �U�X���HG�<idD��d��&�Y��A��I]k�<	�LO5|�H:��A�t�Q��K�e�<2��2+�pK�4#�]
��_�<�p�J/1x���Eѹ
*�`��DUu�<�vO�:�CB!�Q�6 ��Z�!�D^&M��lЎ���%�S��Z���=O6rCJ���8u	��M��5�"O$��!�)
�(ܒ4�\����r�"O�1CE�5�n|���:.8��"O�� ��	a�q��Ę�SB -�"O<�	U��.Yq��#�c�>F�flQ�"On9�c�ܱ7g��p�$'.�S�d�Ot��͎h�,ɹ�(�m�b����=~���U��\5�%��ɛ��J	�����1�^���c��B�,�@�D�}
�B�Iz��
��]�H�)�0ԗQT�C�I86hp�J�&K�e��(���C�IG�4c��"i!�� 1͑%~�,B�-��9�GlJ.c8��@���0�O����O��𤟬S�re�n�>~�Y@��<�!���]n�eȂ�Z� ��xR�~�!�$
�NӒL=&3z\@�%��G!�ül ���I7H풥��H/!���]b�DY�`C�R�x@�L��l%!�dϒ~�	j�*�>1���1����!���lt�Xv��5h��ĂG��IꟐ��c��S�e��b�*�F+],�ѣ�.=D�x#EȣY#V��`�+3���"gi<D�4Y��\�J�b����
5Pj^���O����S��{r&�W�xq)U�JXR��ۤ�y��:"*��0�+�A����W!�y��2}vIkCC�'5ٶ�y',���y�A^$-hV|r��8*ƌ(�fƔ*��-�O�$"qL�A �a�+d����"O:�� /�vʖ�a�\�)�ȴs��|��'6D��$ڋ	���Ӂ�޷ ax��'��p�7��VO��p� �E����ʓI��ȳqJT%u��T��C�"'`�Ն�>�q�r�$�������z��
/�dұ��1��q)v=dx��v�p�ME6M1�=�d��?�䄅ȓ�
%ab�L�b��:��O ��)��dl�Q��,T" �H�����ȓlҤe2�K�qP��Yul<`L�������Y���&��C�4����"C����*�u����4(�ȓh�P�Ԧ�y��MP�Z2���	O��ea�8)fdH�Mډ3/�����8�5�ђ;36��@+7����l{�bʣ7q��+GJ�'M��i�� �L��"p���ۓn=%�@���GȨ0򪁀L���{E��0"؞���_�E����s:*(�5.	,a�m��Io̓����࣐�[��dS�"�*g��E�?�ӓI��!�d�L��ʨs"N�;DB�ȓM��)�ԃ�?1��x������	\�m�,9u�ä()>z��P_�8��ȓ��Lf�O�N7@<�(K>�Q�ȓ{|:|j��D���)��.F���S�? ) �N�%\:�j�K�8MN(�V"O��  F���D�����>4�����'��d����I��C
m����g�;7!��rj��cȝ�l�> �'�30!�$��]�Z����ڜy��x&J��%L!��<w6$E�w35�|���"1�!�䞾l�p�1U�r�e�� �SV!��!�&��� ytp�1�Ј!�D�_0���� A�O�f9`�]*"��6O�!c���4i��h���\�����"O�������m��y
��$J��!c"O�c��)mx,@+%ڦ։�'"O�PR��Ih�(����-y.�"`"O��j��W4z�VX�D��.2���"O�)t��.�`Pig�ѪB�"OΡ�w���l����NƦ�q�'���6a��=�׬G�����k[�7�ў��ɓqĮ�6�Y8�\uaԮ3��B�71���xF/µd���QҮTel�B��:��|q�,֤B��ku-H�d�C䉄&~܀�1LV�,��=s��I�C��4(��y��5u��E��	�,}�B�	�ro�8[j� 'n�<"D��;�˓��<��O��p�jJ�]X~�r&u�@�"O��j��H+/�r=�D�_�&p�"O>���F�9+v �i�Ɲt�^T�E�'U!�U�+ttiH� �L�"��!���KFZl{�kLu6ȉ��,�+t!��Կ%��x�&�5Q��ܻ2쒳a	!��5F��a�˫zJ�����}��'2��~~���g��@#��*��#���y��ǧW�^��1���̴@8���yB�������b>x8���l�8�yrDѪc���d�ن9���)&���yR�G�U���W�#-v(H��G�;�y� l��đ�Q7#��A�d�B�yRd�	[�P�[���.�)�d��(�y�Q�2b�JB�ѯ9P�M��y��r�$�#���X�UC�BY�y��)e�n)h�ەg���&��y�Q;F����Ə�8Sȁ<�yr��`+��"S-L�|��\2S��yBBɾiJx�5�F4f@���2�§�y�E�e$�oK=P�F�s2�M$��.�O�l�u�P��2��T�44.�K1"O`���&V7�8�&���L����"O��0��ɾw�>PaS�Z�8^H�T"O
B��n��q�V-W�W*J�"O�ZF�ϧW|�����LV
`�`"O�T1�M�]J`�j��6��ђ�'�1Of�K#aAlyV88B��s�z��t�' �	M�hy%(�-W��͐r��O�<��h-D��A���+Q��]�poً~�"=Avo&D�x���
!K����U�¦Y�D�e�"D��C# �;�flPrg LI����'!D�$�lּk�2�qa,^�%Q�u`o=D�P�3!�:��(���]2a�ΩZ�a=D�$(%��y��%[!�H�@k;D��r�AΜ~�5 NسEW��2GJ;D�胂��CMva�����m%|�rg7D�,�Ӡ�!QRܡ���B�\�Y�rC�I�<�"lᑄ�8t���S�H�M�JC��,e�H�1�F�"	�0x�&D�%B9C䉵r�P̢���6-��m�TĦ;�B�)� ��fd�he�艵�\�Avp-r�"Ox%�f��Cd"���L�-� L�F"O���ïҩe�`r���4�N��p"O�10�I��2���}l�أ!"O�Ѣ�K��@~���BO�+Z
�`�"O�� ��;|�Եyb�:e0:��"Omy��C!`�P��CPJ���"O�y9��%�z0�b`J'��l�B"O��s�Öc\<8��Y��9��"OD��w�D�=,P��V�;-��Ac�"O@����ˆ�x1.��O{��"Oڼ��dJ�d����m	�pzyA�"O�X�%� 5��0�*}�G/xY�ȓO��Y���0�L�ɤ��nI�i��	��IR~�Fj����$K&4�6�[�S�y�1h��Ԑ�,G8�����y�lҜ$a~���x�|�@=�y�cIH���(�%��t�l]S �9�y�ː
Q����S�@�8�����y��]�^~>psTk��38ш�aO4�y�Ҏ�0��J�*$�X��5�9��=����D��rc<����/3�)p��'Pp!�d��бD�=T��6��^V!�����z����{�& � 	p8!�D�]�X5	�d�������7�!�Z�Y�����Q&�H����9X!�d1_0!�P���WA����HMU!�bF���(��4�t�tGŉ6\!��Q�ȉW���ۆF�"O@���C$Ѽ��N�g��iˢ�� R'��D>�	ϟ@F|BB[����`	�0}�^�)&3�y�S�%����y��lZBg��y��R�Yq���:X.-���%�yR�S�G���rFI&|D��� �y�Z���F��VTM��g���y⬆�,�� o�+���P�I��y�i\�j 4��Q�U����?)�r�'��y©G����dҷX�Q��<D�l�c�� }�2������r���3��<D����a��.��T��0aV�D0�:D�l�!�DoP=�Ex؈� �7D�h�H�^��e�!1�����(�O�=E�$+].M|�b&��r򼼐�n��%�������4� }�����I�@w���d�-D�4˴�"���;C�F�IXmP�,D���s������oF6i��1���'D�4�����v�R�b�-h��YcH1D��B��Q9v�
��!��
`#�m[��,D��a��moh�-�s�u9���O^�=E��n��D���"�;��-0E�'�a|2���#��]�	.������y���!Ar%�2mI�yfN ����y��/ pi�S�Rs�6��� ć�y�&��T�&�Pa�؀pJ�L��%V.�y�`���=bA��Z��� F���y�ic�|�rd�>f�.� ϝ0�y҄@/�� `v	�B����
���0>�6�[�Y�~E�C`K�4��=�$��o�<aD-]�X���(y4�b�ǐh�<���W"}�r@��D6�,�K�a�<qa�٘ptD����ɇ ����T�<	��{����Gˎ?���2+Wg�<q�nO�[b�H�*���d�#����F{ʟ�b��S���Ls,d�� y��!%?D�� ���3�E��"�9�`� ��RT"O� ���۬VP��B���R��A�"O��kb̀7/9�ܐ��VR�TxJ�"OT�`���#Z�ژ;��ۮ����"O�����R*�T���`��[k�p��"O������.�*0�ѯQ��@Q�Ic�Iܟ@�O�Lrt-K$:I@��Zgʶ�;�'9FI;�bL�NT�
���W*8�ҍ��=O�x�-^�6T$!��
̈+uT9B�"O��H�ԉnR~u{o]�B���"OV}�ª'8FD���(�2�xT3�"OF��uP�
�݋E�T�>��l�B"OD���"C��a4ɇ�-P,00��D�O ��)��7U 2$+��u��2��9!���Wd� p5o־tX���9^$!��f��,��n�|M,���N;S!�dO i
�- ��%LR-�fC�+!�dd���㘸(]|9c !�D�2���gf��Vw�A@ >Lh!�D_g��Q��{c�0�aǓ��O�=��
,Y�J�C�P`4Yp0l)�"O�$Bf!D�Yb���S��5mI��"O��p4�N�z	ČI4E�AO"u��"O|�U�N!������e@TI��"O���F�P�$�c@ɓK�,�ɂ"OX)0�D*fg,��^��!�"�!�S�~�z�Cq���<�6Y��N֩lS!�D\ D=�p����j�dD���/45�}��'=�C�:602�X1(X)krN��|%��j��<�2.���؆�f� ,�d�$D�$Kw�%���T	/V��� �!0D��Wh@4m;������d�v��/D���'�Μn�����>0yl�R�,D��Be�]7`��yb��W�33lѤ6D��qBկ:�`���F�T�2�OT�d�OB��g
.8��DC����G2x)J��O�B�ɔ A��`��:�<�ӌU�=� C�	AhhI���Z@�XA�_�X� C�Ɉ~+V���DI��(�����B�	%a� 3��̀'M�;����B䉬�&��	D��0���({�TC�	#���"�L3&�8�G 2<���O&�-��\���@�,F��`N,�������>��'L����n�w'��;�k\;Hn���'^n	�w��"m����⎎ED�l��'bн�w�kN|԰p���A4>\K�'K̽�rc^�!�Z	�gl��:�l��'� , !�
���\B��H]oȅ�'T^�z���@]���P��x���?ɞ'�P�KB�E}���s���W�t�����ϓq��DX��D�&ڈd�գ��RQ�ȓh�8V�0M�PD�B��LLI�G"O~��%R�$$�,K�ƅ <���"O��
��6X%P����/ �1�b"O�����y�01s�B��N#��'��ɦcO�k4��B ��P
�ds�M:��M��� �L>w疱P@��{y���Ā84�tPB���\͢A$*6�ҷEBq�<��0�6uJ@̀e�ldr&��j�<1���*��%�a&� ��x�%�k�<���U�y
%�a�֔\�����`�<��JM�m	r�kS�*a����T�<Ia�+��Xr�;O��H�i�Py�U�����RM�FL=P�����33<�O��=�}� V0C��^�+�t��lȁ2P!1"O٪�Lݲ,f(X�L�8�b"O��j� �Dw:9��$]��x�@�"O
�0�?����#����#"Oz���Ȩ�
dc��hN�4"O&��UG��چR�'ߊy�pyi�|"�'MJ�PQ���o��Y��j��x	�'B
d����[C��6d��!"Ol(`Q�L	"��	�UB�`#P�""On��g,1z��ª� � u"O
)�N�����1C҂ :<(a"OD]9f�Y5w����S,(��a"O<�`�(C.+\R4���t!�j�"O=Q��� V;�H����IAp�@U"O��1hXQqPtɲ �5nͰ��C"O��9���F��@A%�"�҈��"O������/�@�D��H'��[D"OLM�Sn]4����b� �Er�"O��8���$T�"�p�m��Q)�"O�Dkt;,i�'$(��"W�'��	�<�N���Y��e B瞷O��C�I�N�
E�]�:�j�c@��V��C�	,3qD���j3��T�Uk��<B�	"cx�8Kc��QFB����"+#B�	ql���'�&:�>E8�	Z�y%B��{O��!&k۷WVЕ����>cB�I�K����.QA�Uk7���Jyϓ�?��yJ�;1��ie�á%Td�#4�A��y2��K
���H*,�P1�H���yrɅx	��E � E2rA��y,�?_��mBe��aAh��y���/w�4ВԁV�M4`���O���yBIָ2�N�Ju&ŗC`r-��ڑ�yRlM��J�i��@���d!�&��>�O8uaq�L��r��F��N|J-��"O�����H�����9`X<�%"O���H�)�r�*`8("�-B�"O�9�W�Q-
(̱��G�KplA[�"O���G�&+rP�q+ R�p��"O������b8�6K�4C>�+""O�Ȼo��t���K�)�i?-��"OV WF93*�y���W"�*�@�"OМ���(r���[!OxJ��$"OHy�Ĝ"H����!.q���p"O�5xn�)yL\h�2m�3n���"O���㗢l��1�ҩ�TFt� "O!�!�N�L�X�'	UE�0�R"O2�k�B�I�DXWFW76�hH�'X�����8B -
ӏ^���ͺ�'���h"T'�zlc�i_�5.#�'Ő݋�c�7F��T�Q#͡3���'�(�풺;�ႁ�@3�va�'*XZP+�e3f���ͧ+6̚�'���v�֗G��h�M�8�<ؐ�'�\�֌ �r�b����4\�e)�'
�b�L֑a��*�˕-��)�'&�)ce�������C�('+��j	�'l0�Q��
�zJJi�4�^$�`-`	�'c���Ԍ�,HR��8qA�}q���'4D|@R�K]��ī��C�x���j�'����L��M�X�I�āC�<I��'�J�S%P�/{<�[uI9q����'��bn�.��a�M�2�4pR�':���敋yWDi��D�W�#��� � ������m�-\�9�A"O.Y�Ў�pqZ$Z���w� ]�"O2���ɏ�bk�E{�H�&�.ɘ"O���G$�m���aW��vخ�p�"O�z�M�cH>��(K+44@��"O�����G�Q� �1�Ҡ*y� ��"O8�Q���i�����t��"O��)��\�L+h�Z Z9!����"O�������t \�1#�ԝ4}��Z�"O~i	���@x�3Ų[
��"O�` �f�U��e�߼+�iW"OIz���-4[ �00�|M
5"O��R�@A0AOj1{'��rk�՛�"O���G��"���������8b"Ov! V�ɉj��magd#}<y��"O�l#\1
()GML-V@E��"O����"�Z��0�4�i�"O&�ٖL6�����M�4v�Q��"O�[!e�wD	(���	��|�S"O�rU��)�������4�b5�B"OhT�&��H�F)R�;���8u"O��5@FT���@���]_���"O��2�Ǖ7E�8���}3S"OLm�s!Ɩp����QHae`]�#"O�@Z�GQ�5���%�a�H���"O����M���(���K]�zT"OJi��I�V�4��	�.�(�QC"O�d��GB�C���@�:y�\�Q"O���`o�:qcl��n	IM�L�"OTEK��'r|��x�,Wt]C�"O�y�AIT�}�Ҋў��� t"O���4j�{M�=�	�E�u�v"O���pǒ=��%�TǕ;S'ּS"O�l�1j��x���VeF
ڭ+F"O@��c,N7>��0����S�$���"O��1,M�p�I�B�ڹ�Ƙ��"O�Y�Fn�9j�lH��2�~���"O��Xf*�"$�J$xR��	I����u���1+ٟ1�J�C��܇;�¬G��'Y>�S2G�;g�"@\�|PY{�e!ړ�0|�A��X�09J@ X�A���Z��~�<�,��_.�(Dl�;)&PʂDX}�<	�ߖai&��@�?#�lqPfͅy�<Q��
�N��y�L�:W�0(A�Tt�<iU(ͥ\J�A_9��Y+'�r�<�.�02�z� �)ʊMJMc�^Wx� Dx��B��)��cިA�|8�RI(�yr�M��L�At�K�;C�0�a%���y��[��4��ֆY�8��T1��ˡ�y�ԿAǒ]Af�=+�������y�"�bj$�W	ˁ.Nb��6�y��Pk��q�VS��8���y�;9�༛#��7ER�`�G\���O��$*§J��
.Ϝp��+��U�?��I<�i�����Dl���JgG�ȓ ��R��4K���Ǽ �t���t!2�JR���~�%ꏐsS�,�ȓ[��)�A�$1�\��N��qq�ԅȓ$Z08@v)QE�
n����ȓI�Pp8�Ő�#��)��&Ȕ�E{��O]�eϺJ��P�T�C&�@{*O���B�2�\�O��,r���`惕Ei!��r��'�Z�&-�#��L!�=c�LS�	�3�\�'�Lk`!�� *d�g�R�86ڹa��M�9)|)�"OH B��J%D��9��c�(l�r�"O��C��L1s�
i�����R<Q"O��G%�z�í>$y�"Ov�y3@Ř,&xxq�I�f��(�5"OF���ݑC�TI�c�)��	�P"Ov�zR��=t�h�F�3L�T��c"ON�c�B�g�漉�c� p�J0��"OT-PI_T"����I�T�M�A"O�E�OK�U�&e�v�0oʅ["O��ȵ��C�Hpv'ɮ~�>Y�R"O��	�A�o� �� ���p@�G"OD�hPA�>��fQQL��E"O8y��ôs
��[�#�	(�61J`"Oh�pf��/�tx�R��>��ժ�"O�,:�	��NЪ��Q�^mz��E"O��
�  �<C�����M�2F$�"O���C�^+`W��D�w뎴)�"OniR�S�������85�`�"O�\@�"<�e0�"���N��"O:�!�$LL!&!W5���hB"O� �*h�X��
E��IRr"O�����D1|�H�/��|����"O��;Q��xj��B� S�"OX]kg���Q��;V����"O�`��G�t�(r��	\�d�k�"O��F	rip�h
[<���"O�|Iq�
�$>��[0nM�^���"O�ؒ��K�I4lM���΍��!"O^�c�Mqm",���G�\��\�S"O*`! ��:G�+㌇�`�a�5"O"��R�� �AE⍸-	~�aV"Or�f�[)E��P�Q;,��(�"Oh���$J�rp�y� �F�l�Flp#"OJ�넃C�{Ͼ�8�ʐ1�&u�""O*�� D�	X�0�*�u���1"O�r��@:Go�ːjL�Nu�I�w"O<4���I 5#sf�ӡ2s��s�"O�Ŭ�=��1!)�*\(-�5"O��1ׅاN�b��0�B��!@"O��x�'�]�L8�Gx�Ti�"O&YG<N�Q��,yq���0"O(DY��2��I�D�]v ��	�'�>����N;7!LZk3�ٜ�y)�n�p�d聂�$@$+_�y��ͷ+fp�;�(Td�93�Q��y�Ö��4P��	�FBL�bh���y҈�8?�:�i���@NЙӆȎ*�y"�,%x���>�F4у)�yB�[@�{s�#l�m�s%��y��gx�MB�*1��P����yb��B|�yyQF�!�P,�E&�4�y��ٔcV$tzP��;~ɢ���y�oįK8Ų#�X��*V<�yBΘ�#��W
�@��BF�y2�Z:"ٸU��$2�,���G��yb�H=�Z�ccc�>����)4�|k��,.rf�Y����;>b}ˤm;D����V1p��e�ЁZ�_6$ R�8D�<;e��
���ue�+����,7D���v�m�R5���	����h3D�����V�^�"L��b�J��5��*%D��Ir��]qCj��?�ʥ��/D�l��	6�*�`��iL�r�j)D�� ���"�R�?�I�d��2 ���B�"Oʅ"� ����0cD�$ii\���"O8���A�aў5Ó�:�ᱲ"O�(0��.�ɆC��+L�1j2"O|�2�ʈ(y떅[���<s�N�R""O���ub�~H �������Y��"O�Lٓ#Z;z�)�3���B�(ʔ"O��'�Q�.(a����i͈1�E"O<%��a��!H�����K�bD�"O!ˢ탇~����4
:B���"OH��R��Q�&���xs"O��j��]&[v���M.x�N��f"O�	�r�?�b�	�,Ƒj�(��"O�؃Γ�T܌���Ꚋl�
�U"O(����F@���*��S�F��"O�HS�!�kH2);�H���� �2"O>D�l
�BP|��$.�z�Rp�v"O�"si��sPXA��lP�8�{�"O�)�	C�E����ާǤ=��"O0e���6g��gK��Q"On�;A�$k:n(Hƣ��%1l��"O�X���HC,�TZ0��3	5�)w"OF4c��"G.4 cM��z�xd"Ol���L�m�ꄠc�A33{��"O*�ڡ�ؘ	$\@92�J���Bs"O.$�JZ<7�\���k[7��bV"O0�( A3� �8a͏r��3"O8 �m�<Y�ݻ�@�%!�����"O���Ê� r�	��mX�rQV"O��򷃑<+Z:$��	uA�=�S"O�ᢡ�X�f(*sH�5)$��f"O��X�D�#;��Qe)�8���"O�AR3��F�u��-�>m��M��"O@ #!Q7ꠁP����w5>ҥ"Or�0sgU�Tڐ�S�)cTX}P6"O�%�����@L��ѐ�>y8��1�"O��s�!!�ԛ��G9DL2٨�"O֭��M,{��Ec�(?Jv��"Ox}�s�� !N�<����;E|��"O�ت"�ǰh�JA"�.Y'	A|�!R"O�� qeJLq���E;���"O���噓��!C/�Q0��c"O��Q�f�>j�ibGZ�`ߘɢc"O�E*�ĕH��3��ޠ.����"O�� �	Rt��a��*�&��a�"O��i�!	f�f ��,����"OZ�Q"Z�Sv
15�8'x�"�"OX8�H8L�N��㥆�3*��V"O��z�d[0&����Ą~��8"O�U*`�E��8X��E���`"OT�$IZ w�ε1���Pq!"O&0�u"��C[T�s��-C�v��P"O\��0�ͱ>��rC�<#Pn���"O>�����@u�1;�G��N�����"O��T�y��i⧨D�����"O���F�$5����UH �({�5��"O6�+5�i�"�k��G�[p;�"O��x/؛;�T�b���l���"O�r��F_�:D�S�O�Fh3"O�	Ɇ3쪍�SM\"8�>�"O����ĕ/�����)�	�ؼ�"OR�B�ʙ R��<	��G(/~r��@"O� aA$t�\�s��y$D�"O��3eS4 �yf�,q�%k�"O� 8kACE'3���X�@ :X���"OH�{��й`�~�p�ɖ"��}��"O���R W�q��/����p�"O�;��K����ܒHb�q��"Ot1W�%��X�Ώ/>\��i�"O��i�NR�@d���,g�L}�P"O�5�gM��!�)�o��V�~��G"OʩR3��EȨl��g�"Z`^� �"O�	�]RX	�ܝM����b]��yr�΢E7~�d��;V���1�P��yMǖ9��)�%|�����V��yB��8ym��%.t��$�y��[2d�Ȁ�μ$��a��?�y��%O�X�W�(e�x����y�D/o��@QJ&Np� R���yR��z�Bܻ��MJ=��)T���y�,W�a���@@���V�T'K��yR�"y
p�h� E�[�PtY"ٸ�yBL[�sP0�%O�8O��`�᠔�yA��ez���f��F�B�@�'�y��Q5V�J��*D����ތ�y2�H
kh���Wb:5|����#�yeT'rȉ����3R�1`���y�#ǡse�\B��Z�,Ϥ���B��y���5;@LtѲS�&y�јV�G��y2P�M(���H-g=�����PyR)7%���l�SE�� x�<�Â����$��<2����!XO�<Q�΍~����l�����b�Q�<yĦ�0qn�"7%�s�\��3F�O�<��!T�9W��іCX"�l�EE�a�<�a	�^�1�%�[RZT�h�'H[�<�A��'�N`2��U�TN(=��V�<aA��
�~q�$��##����mP�<9E�:wD�ks�_8x�B]���GP�<YE ]%
�F�����7z�JL��Kc�<��B	�.�btYR�D6r=��YF�b�<�TdE:Հ�`ԣ2 c|*���U�<!��U�Ip�R�A(�d
'@Jj�<�EB�L(B)J%k�`�`�l�<��� �MSt5�W�!Cg|����i�<1�\<Aؽ!	B5`{� �c��<q �ļq1!�		�Y�XK�a�u�<�o�/$Ej1���R�X�� KԎYW�<�	+GR�)�wM�Q�<�w�ݠ��y��C���b)�K�<�w��N�����������lNI�<�hLX����Գ7��QRD	�F�<!V��B�*y����/Z����kP@�<�p��%d}��	�t�\ �Vl@r�<���W�k�zPCGS�=K��aJb�<�r��-(�;������W�<����%1n`(�J�������V�<i◀]K
�*�k\�J3����^P�<1de S�I2��,rS��a�Yv�<9�W�W��X1�H�'b�=���y�<)�$�BBPǉ�n1���I�v�<QdJ�95P�sn��]�tI�h�<Ad��x�y2���=e��1���@c�<Y@�/p�z��%�F�tlĝB���F�<����>.�x�.�n0���U�<ᑦ�]���V�|�lk�G}�<q��#Kq,`:���u���T�LS�<�P��0��p�ЇCv�}�u@DO�<� �dy�B��i�>d�7ӠF�hIS"O���1�|��-2���"OJ]��`�	)�6 ��L�?X�TkF"OKѾ&Xma��2o傰�O��y��!R�I��`���A	�y�&�w����D͖g	�lń�y2��S��yK�J��0��F�y����t�֑��'!�eq�)�*�yB��,�b���0qh�=r�ȩ�yRe�$2!y%&�,m�����y��J%� S���8QX�����y�3if2��!W�*��i$N��ynViK��ban�)"Q��TG�"�y��
�!}�t� ���"��
�yR�7 �(��h��H<SH	>�y"J �ƨ��*�~�x���,�y�F[ ]��}�d��E��܋����yR�X=^H ��!ƚ89����2 5�yB�����%�aE�m(�	��y�cK��z����R��8�����y���<AN�*���K`R��siF�y"ϭn��P���'Js�i ��E�y��X�h�`k�����'��5�y"�ݝP$�Ŝ���*,�yr�	lMޅI��"/����J��y��NN��z���*tw\��`���y"��OvxX�*�s9�Х�;�y*�f���BE�zp~�"N���y�,_��Y�7��H�������y�b�4#~B���k�$U/|]c���y�e�v��[����S�8��QkL��y"�׃G��hEl��T�4-�e���y7?�p��� уL�8���	��y"�[��z`�S�>B���m�yg��KR�I;r�=%�ر������y��Sz2�@�%�"W: �d��y�͑!�rp�`�+�e��Ǔ7�yb�A�aF8�i#+ߘ'�Z�Q!W+�y���uCnh�rɥ!�x40 gJ�y�l���)9��
!� e��N̳�y�855x`���*����I��y��'k'�M�E� ���Dl�y���h�p�*�X��
E��iG��y.�&Q!vɅ�t�a���yB�Ea%raQ!S���Q�ҭ�yҡؖ&�b���3G�hp@�1�y�b:�� B��6NP\p�A�3�yBh�Y��5�r�|������y�ω(f�t����dX�p���H��yB+շO86h��DſUD�1�AP��y�^� �A`C�]N��X��D��y"%��)u0@��IU	:u�P�@��y�kމH=��f/��1���"H��yҮ�1<����R���-{��z���"�y�X<E�=!e 9�
��q�ת�y�X�w������dm�� ��B��Ts�IО �A(��C��B�	�]�����d�!G��)&w��B�I+$���P�3�c��6pB�ɔg�a"�D�#�l�� ��-4��C�I l�H��!鑥hF��UO�~'PC��L�yBA�>]����5� ,�LC�I�c|X�����0�8���	�JC�I� ��i0t:g(ȫ����P10C�)� Lݢ��
�_$ ��N�1U��y�!"O HRKԈ#�`y��u��ň�"O���j�*��=��mc� ��"Oy��! B��� �-�<9Ǵe�a"Ou��j��m����S�u��"O����
Z�V�8���E�0�!)�"O��9!o�+z8r�����Y��Z"O܅3�n�3���U�o���c�"O�}�4Ԉ;D�2T�!����"O x�m�F�M�b�!֦�"O|�S˚�h�]ї	F�:��h�"O40z"k�?tj,���&���e�'щ'��T��w1f �r%M0im�x�M����I�v�,*v�����e�V�a����{��A�ب0� )���ַ�8Q v.-|O�c� ��!�~�A�#ԇ1[(�9e�(��ȟ4 [#� �B�	��F�&����b�I�:}�>m��D0��¤i�<]��L)�F���E{��)6b��9���9����ѦեC'�y��1M`1�#�=-��p���3jb������@�X$V�J����n��1?A�C\6�qS�L�-XAT)"&����B1@tK�ڗ��-	��x�n�ȓ='������<9���P'�kz^������a!���H��e�V�U��ՇȓWD�i�HCʼ����
".7�O�O*0��
k�ȁB ���rGx "O�i���k^�j�A�1O%��G�'E��-�ĀfJX-6��0�DH*{!�C��	D�P)�R��V��P�n��d0,#>���ƻl����fE�6H�]���T�!��O���#)J)n	�A�u�>dƄ���"O� ����" �R98��GM����'�>���.��n�P���6�y��,<��p<�$L�u�p`fJ�	�2��#��r�ɕL�{҂�3p[r����ԧ���#"¡�M��'��;��%T�8�Cʉ2��1�'�ў"~��"��2aׄ\N���"�Li�'�?�P��{v��R�fS������0D�|���2J�J$[ԃ��M=���m9<O�"<��!�,�Pq�1F�\�����l�<�"�"U���4�2�� g�*p��	v��M�?i����<�N�{�,^�� �sf�*P�!��j�J:�R�u����H�~�'�a|�.#A�a�5N� @�ҕ���Px��i��ɗ�(B��Io�k����'C���iC<&����sd�.W�-��(O<�s�����q3'�R�!	�� "O�	q���V�(ysR'�; P`s�"OvG��:Fe��5&�
���W"O���&�Y40X��&@6ۀ;"Oy{�֢Q:����P�tQ"O8�+'��u0�j���B��}KQ"O\Yjw�M
-S��5mB�D�6�R��;\O� �n�p�����i��q��"O�ej0J�V��y��,'w�I0�"Oz=���)�A;A�޳bl�(j"O��q� N?�,H۵(���"O����g26�(����2�$<��"O차�\?o��|2W�E.;ٱ�"O9���]�{���� ^/Q$>�S"O��0Q�Q�<mh���]�ʰ�"O@���>��ԪW�֞}�2}��"O�9�SJ
����mG�^���"O� b��g
��J1���Yv.1�"O��3f�Ӛ0t��b��O�<o�K"O��`$���g�pP�Q��J�$��"O�m��H�p���G�����w�'�Q��u��u^b�1�O
�*>�(	ׂ8D� 1����|���G���Aq�)D��Ye��_U�\B �+/����f,D� #�	�����Ó�'Rw�Ik7cn�ڣ=E�ܴP"p;���aÊ��K_;mb"`��e�j�#G��0q\XakCI��8(:1���?!��6#�r-9��4+ zm1SM[e�<��'��poba� ��g��`p�
K�<Aw�]��A��.�ZY��lI�<Q`��!�|�"�)AJ����F�<��;5�^��â�?L��9�G@�<�샐L(�u�'/.�%b�o�C�<�n�V�u��	;#vy����c}�)�'*G��`�+�Pa,����L��ȓb;a�&���3����EƗ丐l�;��$!�O��Q�0DXM�#�C��\��' ��O:-B�"�tR��+���#����e"O&x!t����yQ#�\�\�*d"Oq�PAV�@h�"������$7�S���}���Qz&`�uET��B䉒Qg"�;@H�y��q�Q��:a*#=��4�䓱��O��t��F��JD����|�<�
�'K�H�	�(���ȿ-2���'1ў�}��'E�l\̀*t'�e�ȃ�Q�<��/N�|GD�K���:EHalVv�'�?��@*�;x�nat��N�N�7D�2�J�,�F83�B�>2,]����O*�$,�)�'+����Z�]�TTƌ���pH���hO?�*� �0Tq�Er�?,(xx�c�n}�(ZTx�PUMӘr�(��t�	�a��1�9�O��?O��I��'UT ,Pv��x]~���"O�x"�if���K�a@"���I|>a�W-	5(�ب ��W�g�~<)T�;�IA?�{����9BĚ����7PI�1�1��9�yR�֍x*F�q@�+F�,YaI�y��6�r�j�D�D9l�1�V\ �X�L���&˩'f��	ވ-���I	��d�<���Nvd@����<�r�k(<q޴R��5�R6L��< ��� C�*�Ex��)Z�Ѳ0��Y8u�9jE�O�W�<�7��J j$��i檀�s��i�<s
U�8�]
�$S�$U`�[%	}�$8�S�'*�:���Q�&��3���?�<��~66��wBW��Z�[ ��-=��=�	�s�QDE�(%�r)۳RB���ȓ�nő��
|L���]�V� ��e�yc"L�Pzؕ�'N���1��aM�t26'�}����(���ɇȓ=����`/���K0�ȩp=$��ȓK| �B��&D�� {R�N 2�P�ȓ[n�O'��z#���F�؆�>B-��kU"B���։��}"px�ȓ�Pzqb�K� ���Ɇ1�2@"���s���A�=I����$��L.�O(�i	r�&�N_^|U��.X�o�༅�g��E�`&���$a`S��>5W�Մ� G�a�$m�/ X�H����=����i�$�E�_�̔�1��2U��H�=qۓ+|dj��1�ԙIEL�$cr�4��)����*��	ڤ�_�v��EnZD������ L� �g��cܺ���G�;!d杺��'-����Ha�c'ڟ,Z.�Z���eC�ɣ^�B<��[1����*Z�q'�#=Yڴ�ȟd49Bc\$֖�HfC��0�)p"Oh��͓ a�����\3X�D�!&"O����+�	ǠaA%�?\�h�@�"OR������aE�v�z��F"O���� ������Ôo��8�"O�<(�%�"�S��Q;���0"O�ۆ�D�ĭ��		4p�q�E"O��k�GY�X���(IOzf��"O�u���  yDXB�%z��a3�x��)�S�sl�������&�Jq� �&(o�B�ɟ��Lh��wp�H��k
`FQ�=	����~�q�FS^"4��ɜ�.\�ȓaw�x �L�s&�a笎3m���ȓ$@��S���C�¤P�@��$�ȓ$�ƭ��N�Q,���@]�;鰐��[Yn x� ��Z�p�X����P��i��P򷃑�D�@����B�� �ȓ ����6������ �k:fE�ȓt�De�Jܿ=�2]PSQ�U~
��ȓI��(��g�+!����F�@Ϯi��*��h*�R}� �!%��91����ȓHz�]��T����WA+bgnU�ȓ'�.��.�F� $��R�p ��ȓ欙���=��X(�h�L��|�ȓc�*�s�QҀ��5�S�Ax,����ė�kh�ӗ�U�K�|�ȓu�0�D�]��(�T#Z��]�ȓ R�xq��A)�u��H"1_���ȓ<���0�������Z5B��h��Dp�;3Cb��VTnm�v%?D�p���ε8���a,D)RN��)D���a��o!�L���\�PF6�`�B5D�Py��ȐU�B����[�zLU��d0D�t!T�;�Q8���5��L���2D����R.�(8 [;ene��I1D��gE^$�r0��EAb�k�:D��ࣄS�j���R�B�S�(��;D�V��U�q�aE�|��"C�\$�y��ٶ-�����M�oD��R _�y���:Y$��%k:g��uR��$�y�X�\�D<h!G�))��2����y�_&����0]�!��k��	>�yD�/�4��Z��E��y�X� ���  ,5z��U�yO�#���c���Jq�,�$C�y )r2��� �N��!�⅔�y��LvUr�L�#9��Q���L�yr#ۉQ2c�N�;93@��M���0?�֥�P�*��
��u0��R _�D�eOQ�<�Nv"� ![0Q��lQԫXy�<��XK[���g��&m�>Ѣ�O{�<�R脪EA���
mP.�#c�r�<6�
O:���fZ�c.�)�fo�<�ǾV\� ����^���I�d�l�<	�c��3��vF�"X
���f�B�<Q��Ɖ:�I�LÊ�AW��v�<#�A�*'ƔHÁ�n�ހ����w�<IV����(RJ����[$L�s�<qU��?p���N�+�|;���f�<�4CFe�faR�i�9^��=���`�<1'mX�a:("�[�,�e��x�<� �)QAR���(
6ʤ����s"O������ 5��X���G"O,�����$�ҕ��<��K�"ObՓa՟D�H@Yj̕K�̱(w"OԠB4 :]�l��ǃ'�Z��5"O�|��)+�.X��4a{`��"O��@wf؁Z�� hP��q{6H$"O�#ՌM�SB5�2)�nj�a"�"Ol`�f�
*6�d�y��V	<\��"O��qGƶBb����"S	�`�"OVdzC�S�HQ`a��9Y<)�s"Oj�RDCO#$hlx!��H�!H�uv�'I�}V��)D5:�R��ANgʭ�� �#(�T"Of9��ɟ�o^F�1�a�1:�>���ɵ9�lʴ��6.���p��c�1i�0}b�B "O\i[T�i�M!@H(V �9�նD�0�����������F�)�й��/Nb������yB���4I����H�1#�yJ�I�<�~"�C2�I���#Oay��U�H2%�B��,ɶ�2c(���p>�+�Vʊ�uȒ!�DaH���+eD�;�ͅ!�2M
�'װEj��^p>K2�-!��yp��߆Dݨy
� X�]u:b?�&D�x��#���#�4T�S0D�T9��F�~�ݢqP�=<�ڶbU�r?d�����.��j)O?�D]�/q�h)PGS�u��1�4`�w)!�؝(���?J�hx"I�"��Ĉ)��y�� �JF��W�d��}K�����tC���w�|�M�#A�u���Y�$p��~�s��R0zT�0X2O�`0�M,UCǋ�mW��Jc�	j�B$�6AI�'���s� ��M�ϓFa�E��"O�)V�Ä}���Ƀ-�%Y ����'�>D�JY�=�ɧ���5�
�%y	"��s���eG���2D�Lb6��	QPe1�̭�� ��c4D���R���L��hJ�^��c!D�|�򪈥7i�� sn��C��%A�0D��QUȕ~6dD��k"�)��n/D���Ҥ�*�Xl�P���ZeH5�-D�
R�* �Dٕ&#-,eY,4D��ӳM��SpiS$�F�!2A?D�8qe�00_�\z0�О/|^��w�:D���CK<Y��͏�B�F� ¦,D��
��M8@�Vy��G�@~28��Mt���gx��kC
�%Z<��A��&`�Ť4|O`����B���$  ^���2,��7#�b!��K/lv���3�!"���ee�O�0�s�M�ȟD`9����1�����\��p��*O��Y���	}�`Y��K�l�S�!�`- ➸G��'A���+_x�r�ۗ_@��	�'Z��W�Z�kA���&WJ�9��2�)�f� �O��AmF�Y�RMK����|�4�a�'����@}򬈢J�(|0��݆w
 ����O��y��Ut+���+_e<\�[�hҀ�OA:�F)��3d�L�N�$��T�A���ȓ5{
@����@+B�zr��pޤЄʓ^��D��-�T�"�xtj�B�B䉵(p�J1�G$&���g�B��
q~�ւ�10��Ha�@�FB�I�(x���b%5/��Б*P�όC�	Q����� 2nT���ĕ0�zC�	n�f@BE�֭E�J�K�ă<zB��|�
2��S���#�.`��C��+P� ����-"�%�.�[ C䉢W�m��đ%���	�呾s�8�g.��E��?E�5�̒l�
 ࣈ͆\��3T�(�O�L��L�L�f�����ۦk�qP ��`�'����Y�� Te*6�<SNa� 	�6Y�p�w�	�h3��2J�D�'i�z@�O�: �Z��!B�=xPHyu�Ǵ|�\�#�Ʌ�#����ٴ~wj%2��2$	��=H,��n
�� @��D��Ir�Lz>��`����h4(�͢�#�>��������M�X�J�dB�I19���(�C6s�b	�B{���]�.�FN�'lq�r�Ԣat���a2O��X�`��.�B1�;_a��	WL]8���N�j$��	>Nh�����\H⑰6j�{���Ab^�uH8��U��k�����;'�1i���9^MF�[�z�1O\Q���!0�<|j�)�pV �p�I�g�(zC�&t�b�Y�`�ś��Øq��C��S�����E耥$���)�j�2f(q���)[�
���N 6K8�qs	�1GZn�:� ��>��Hʖ	��K��ԅ���P�$�d��)�|1��]�p�I"��?���"�J��?K��������$�n,u�S�6iTY����D&���B�Se:�h���Z�F��B�j$2E�ӊ4oDq�eF!�NDQ�D9Ĭ��rtvl"���_�~2��JJQ��`��wk>�2��ĚF� ��U�O�/ !I�&S�ULN�i�P�_�(���S�rg&�b�dD��d�𸳎��+� 5�W�L�>��Gx��O����.ο)�(-���͎:��KpfJk��d���@B��uB�W���F莤,@4hY�gt��xϓk�b�(#
�,�6h§#�.��O�mɖ��mj2 9IX�`�z�	E���i"ѻf&��E��AV��;IRPC��:eU(W���,4��u�j|��J�.��|hD+H�	��q���j����B뉆E��lÐk��p�x\��������y�ƍUP8�A`}�.����T��Ig�I�zj�pe,J�^ʰ����;a����T̨4ɕL��*i�+&h��xEl��uw�|�7D�0�M��Y�D-p���&�O��=�'KԐQ�\�K3R�7�Hm��BV�N��a%�0T,�YC�4LO<!�B�`��}
�&ڲe�|@�'�����X�lÆ�s��@$M��s7��o: (�-͞}�E��mAe�<��#�7��)ɇ�XC�<04-Z��19�mPf���7�x�2�Fz�O�@�CEi
:aHC	Lo3���
�'�����_44'��0r(�v�F�	�Jٞ2�U[C��͟\p�
�����{V0��.��=��`�T�V0z�d��Ɠ�^��/H�.�<�a��O����ǭՀ9��$��/ ������m`���a"U$�(�A�JʫO�z�Ĥiֵ��*��<q���RZ�̓�K]'r^���K�w�<Y�	9E .�K�Q�dϪ��t�t� %��)�'���a �vg8��f�?SJA��$��,9!	�'Y��YF��0�ȓk�,p�Aǣa��E��C?�\Ąȓ���r���~�
����ϙ�����`t��*}P\�[ ��+E֙��I�H�U��P�b�%�䵈a�>A����7k0D�L�נ_#��%�*��$�4(��*�0�tF�T�O�Ι��ɟ���Gh
kӚ=
�'/�1��̕y���a�K�^�^TY��/b��'�L�����>a �
��p`F�� �rLBLh<!p��un��ր[x;Fx�<Ӷ 
W�h	����-��`6k�I>�2��؋@��y�E&�b�-XK}Bm�;'�X= DhW �Μ� ��y2A�'{~���F�"y���e��;��#|���-A�u�#җ38��	�5Dȏ#����gA@x�<a�Fo��L�d�8R�XrP��-@�|x�v�>��@�#����=�:��q$�%,B�x�̖\zC�ɧj4R<k��M�U���4R�,�&#D�!��ye�'�\�� �%;b!ꆫŒ  t�i
ϓ;h9��KE"v�uhY�#ꅠ>�� 3�]�16ԭ�ȓv����#
�p��t(�!�>����<!�������b����.;��1�s�BH�ӒH�5$�!�d�K�����]�mB��D��%F��x���Ē#�(���&'F��rV�H"Hy�a;��J8]��B�ɬDDm�B\�{}��F����B�	��XK&� =E��Y�C�1&����)���],�?%�e�Æ ɔ�HRO��wa���R�+D�,��V;�$04�Vk%�%k��`U��|��&�g}rK��p���vk
no`���A����=��F�XF��ZU"�&�)9<L����بS�����$1h섢��o���(�
�]�T&�14� e��<�I$A�<�Wțc}b)̥gb4)�ԡ��|� ��t��!9�2,�éN� �H!B�"O���p�ŌN���(#E߯8�DpP��8P����Oz�Q�"�SR�a�������Fc��U�~�ӣ��.$���7I�^�<�d�؇ ���C!j�B��,iGLD�M�U��?�>��c'�D" ,CLr�#<�G)Y�$i� ��+Ӽ��D�x������7)(:�$>OV��5B�0Y�T�p!+")�PmU�Y$PPhSE��a|���G�4�i2�B�z�!�N_4��'ɚ�*g�B�"5�Q:�	&�9~�\�S��d�W��I��8�@�-0�ZB�	 ��\h�ᚒ_<�kã���6(��JM�%�O���C�@��n�:���Ǽs��F�{	N�󓃖j�u�A
�C�<Q�◒)Q�%����m��\����w)|%���ܰ-n�͓:���S�b�-[ʣ<��61+֝���Ö?���;R�t�����%�u����#�'ِ�C�>����db�6�R�KY <S��� �X����?c�d�Ǎ�/j���ʧ�:�I�~��}�6���<�e5c���ˇj�~´͋��J!�7ҳT��sA	�s�<Q!�̚?e�U!J]�&%S�	1P̤�s�O6����K�����x�EZ5�
�|˰�c��A�s/0����7D��IDKؘ�\���ؤ�
�2'IX�B��^C�䀪p���?�'�&Aa`�_:��0�â{p�a�'��V)Z,o��crf�F�����ݽd����F�P|X�@c�G^�N�8��N���B��+<O<�+0
��N���O�lS���!?(F���D��Eg"O�|�,�0ZK�q�F�Y��[r�|R��Z��k"	�g�Ow���D{᦬_b�R��
�'�4��4)J@u�ٴ�F*4t\�"�әM��'uX�:���rb��Hȓ�i�.g�����m&D���E��s(�a0F� �~��q!8_�T ��-�O$�@p�K?=�P�-�z��("OV� ���_2h�ڐ,I�
`䘳"O�hС��	��b7KP1���
�'�@���PI�Z�d��a�D�q�'=���fN	V�]P�b�b&\�y�' ä��6B�t���'X��"OD����މ�H�۵C��2@�lr "O$����͗2����#��|`�)F"O�U�F�� %o�4�� w"O:1���SY�QA��	%���b"O��*�OE���t�f�+Z�K�"OȽ,��x^�0*]�?��a�S"O҅±�R
\��Q)֠�:�@�Ғ"OB\��Q�_>�ز!���c�4�p�"O�L��F(d̴(Em<65dH�q"O*]�v��$�eӁM�{+P܂"Oĝ�ŝY�ĸ��P�|���$"O(0K��Щc4���kH9:��"O�' W�s9��k�JK��dғ"OT����	|Zȸ��o�&y��"O"Ԉ�
�+NclP���77��"OFD�M���R5h�ÕZp��yR"OT�S��'� 8s��ÓD(��"O|8�vf��XTʑ��[�/>!b"Oܽ�6�^<>�l�D�Y�X�Nk�"OZݑ�D�X�M0�	Tk�x�P�"Oz��##�[c�	
pΊ�g�v�S�"O:1��J��PQM��OG08`D"O�@��L4+��u@���W��Jq"O��xQB�
�����31��D"Oz	�gjZV>���8/���S�"O�9 ��H�	%~���v"Ob�s��f�Z�YV�J�m{$ᒗ"O��2"�� Ҁ1p��MG�P�+�"O(IRu�m�~;���xCV�+c"O�[@	�V��z����PB�"O�A;fJSM��Q,��I�"O� ���OĬ��M��,�H*0c "O ���L�BX���T�=j�2)`�"O11`��,����FO�\���"O��YAQ\l,����V݈T��"O&���FK-�-YoU'&��j""O��,6��S�,���$y��"O0����r������9_H9��"O�t��eF�أ�	�W\T��"O�%z���L��� ��R�i0�("D"O"�u���p�'�_EF�j�"O��jƓ5c����7���Y7x "O���$�ܾ9�1��
D�I�F"O$��`e�>[� ��P�y#��-�!�9�$�)R��ZA<�P��9�!��D3A�X����
i3X�נ�>s!�D0��aւK����OY�`�}�ىb@	��*>F�,�K��	�(j�@�h�Nd!�D�8/��\���Ē)j� 	VJ���Bb��XE���w���dTʭa6�L�]S��9!oY9�!�d�>0_���Eg��YL�{�l.>�F����(^s�t���py���'r�\qU�Қ7u4�����(z�'�>̪�n�d�:�)B(�s��K�'�f8�u	�G���K��'}l)U�U��
A��;_�h�o9�T�c"LQ�/$|[7�X�YH�0&DL�c#~�:�'��t�Ə�)�ڰ#��� #�H��d�g��H�6_�*��b?�(ǫ�=6Ac΃XY��b��;D����Y�z(:x�c�
w��$�7��I���G"�4:�Ҵ`/O?�DB j�0��Q�3Cr��V�y�!�DؤH�^%�,R.Z0m����"+c�d�c�f���(J&���d�\ڥHiϙ�q˳JZ��|�m�+j2^��-E�~���
�r� �+̡D����7O*���N�X d� �%v$e{��+?����RX-3�n�� j�&r��τ(�a��"OD���A"`����oB 
`���'�,�A�B�|���&!^��M��&��ق��\+0�xC�	�\~�\KT��'���Yu�čz�LC�I `a�Ү]c����Q��D��B�ɏg�<�ː�,(&L�򁖗k<�B�I7b����/S6�:4��W���C�I7{�%r��O&�P����(wsnC� M���EOύENi(���B�It�<	z�iŴq�:�Ə��r��B�I�v�� �q%M'e`���@[;O�dB�I������ƽP��L��ݠTVB�I'p&���7��X{c���B䉾ZG�50��"F�2yB�b
$��B�)@0M�fb@�k���˵7�*B䉇?_:��S�)u�����4h�C�	/Hc�x{�J%>P����=��C�	�f��҅i/Q�� ��� ��C��Z���9_.E������C�	��Z�Qv��by���GG�|}�C��;l�J�D��	7��l���L3X$C�I�{��Uf%���Ƚ�C�	/ ����5�ں�(21�K%�B䉞4(5ic�ܑ"ܜXR��ˍ��B��,]	H�)� U�j��p��I�B�	�LjNXX!$D8�@�:4M-
�B�	�\�\X"�˅:j�~Q�� i�B�I�%�l���M�I��0�bRm�HB�I:������\(�xP����7Mb\B�	��FUɧDS�g[l�"`d�i�8B��)L!*��nV�8�hm(�MO�m��C�!2A�	W�_,N�� �X]\�B�)� �QP�$�01X$���ӃY�t�
�"O �
�/��)�t�T�H�;��Pr"O���3`�=�tX�aE�%�z�p��'�����Q�)&¬�ԫ&9Ā��Q57B1��-`Us�P���!@�MB0x(( E~뚢m�H�kF�韚i�^�)&@�,D��SC�.D!�D�/�!Ѝ��7rڝӵ��O!�$ l�
���N.]�\t�-�'I�4�;3)N�Pnn����H�(��1��c�&8�4��9äq!��ӏF�=��¢O,6-�5-ljP�Q���3�ɣ����ݑ0�(�R��>������"p�H�d��[���e���v��n�CĀ��"k r�`��'ބT�2�Q�g�4�P �u�ܬэ�)�	���
4�	����de� (x��i'l�.�J�S1̇�y"�\�d���Ï})��y�FP�~��H&r���M�3��B�r�O*�uZp	�9 ��MG蛶
�LX3�'�r<�.�����	-*�ɣ�(����΀j���PbR��3�I��<@s�KQ�]I���	BA�����)kt���(x��Dy%{�9�݅X�����ԽNt�����Q�x��l�(kf$���ڒJr�@�"�f�LMs	8TІ|��Y�)ʽn:�6ᙖM���O/!��K�_��z���8 `�Ǝɯ�剪�
���[:%���«�F�O4�)���#n�<��mJ�� �#�'Hȵɲ�B����Mȿ=��$.�:�$�而�Y�0Ɂ��!�$B#�SY�4`P$1D�Tr*��s�,��ズ)i���Ҍ�O`�+���!ΰ>I�ńh��@B�L��b~��&�v�<!� ��(�R��mзak���	i�<���L�LQ�-��ws�EʓM��<9��ƺQ P	ǡJ�H�R���Wa�<1��A4`�$����ސ���[�+Cz�<�5$��K|Y
�x�h��"�R�<���	�bJ���R^�;�I�<9D��T�(̡2���]���D�J�<�C %F=m['&N�M�R(@
_�<�D�X8`7��y�,�6�1���Y�<�'ہ|��@	�MMMZ��O�<Yև��Z���ZFҽ� �@�<ad�ڮB�Լ°OD�Pc1�	�~�<����.<�4��L{���I��u�<�f�ɆH�8QhsCӫD�t�)7/Al�<��L�&Tb�k
�&RʈS�bBi�<Y��Q1F�p����݂c$��A`��hx��A���=�sHG!=�"�Xt���B��B�I+zjU�d��\�5:����b�0*V(X ���F�4�I�1�����ɵ?{�q��)���y��XB�����]#!L�Xi��-��M89}¦W',]��O�n,w.3r���ʝ����ƓD6�`��7? �j���D��`� ��SDDX�C �O�!`�U�pl��V�	�dp��a�'rf肖�aw��'g��Q�?�4��h.6A�@�'�� Q%�%g+�$��T��R8�O>��DԤ�J��+�'���!B?z����鞾1���ȓ �n�Y���S>|q�Qm���>�kЮg��~ dUb��L����肨G;����_�<�r�`�':4�TXˀ1?���uEW�2[� �'����0�#o�^Ua}�Ȕ��S��L�c��@8A
��<Y�g�?`��Xa*�>��l�<-�P��1�6�z�;�e�<鵪��?���q���&h%˄�g�&`1�Ԅ'��걛#E�h��s����l
a"O������>'�()���%^��t���ʩ)qO�P���Y���F �R�	J��Ц�P�C�&D�tX$fwF�X��Q<<Z��kf�$D�tJ���BS�H3r��	��Á�.���p:�����/5��%YS&P�=�89B���#r�C�)� �A���.��'��!j�9�B�^%_�t�H>�b�>�¯�9�J1��3��m9���v���)3	]�R�I���k��7r����Ɉ�@���ѪL8^ndg�(�OȀ�"��cyx,�P$G�D=�T����5&�#n�>I�aH��n�� Iu>)�d���n�����.Ɠk�W�2D���M��ANZ���D� �Y���Q*]ܺ11Ą��T(��S�p�J���)_��y�'3!�6(�Q���x������y`�?kr�X	՘�~l���]F
��㶁։q�\�i�'�8,l��D�Gx҈F	$e|�x�Ip�P�X��S��p=A��-+N����m��r��&�h�� �a�N�CS(v�&�rG����D\��ްz�Փ`<�)���BRqO؀2tN�"/�L���'M��p@�բrHA�'��୕*y8!b@��T��ȓ~lK~����J�f%��%`�=0}V�w��0;G�) k���c�	��yW��9Eq�}�ե�?Q��A��R��y"�J�)ޔ�H%��,U�jĉ�J�#G���"MH�Q�4�B�'� 	"�J�*ր�Dy�eS�B� ��Q�ZA2����p=�"��*UW��	���Om0tJP�`�J*ғe�l�#)I�A�
�2��Z �>�r+�6,����N�
�ꬸ��L�:)&5QT�J-�y⣔<�>���b�R���8IN`��h�K�Dy���Ƣ�y2��&�������.@|2���T��Yy�￟��a"�>�0G�ʼoV�(D����
0�M��y�ǅQ^@�u�M�<�,=֍��bt ��!}"ۦ ��l$܄����)z�(��Nƭ�2�Ɠq��H)���aq*���Eh�8p����B�"F�2�Oe����i�ף�*�XђR�'�q�w�T(�P��'t@I�+Z�nl�Q1��^bdԍ	�'if�1o��"��̠q
	�]�� @N>�Q��.^��8h�F&�'m!�M��FA7L*�8RTGL)���r�`�0+�+w1��I��N�
�J8M�q$��W
*�g~���t��D(�I9&��P��&΋�yb�� �h�@"��{�d�c�R�-F��p���0?�cȟ+L��3��h�,�	��M�<a!/O�i} �*cR�I��a�m�|�<Y'.I.��ҥ@y�%���Q�<Yפ�Q
���9�L����N�<16L�.� X�K�M�<-��·q�<���[dtI�lխ?\��!o�<1� �iጰh��Y�K�k�j�<��&���+�t�HD
�ȓPs����Tg?��$ꙉ>ܩ�ȓa������!R�*a� O�qT$��pP�|/�--2�kҵ*�����
Xi��Ħ�:T�I��v�t0�ȓ��@���׸ tN�*S�­SM�������#`��Zq�&HMA4���E��2&%�:!�Q!��e����2l����̐�{����߼|h��ȓuj�Y�-�aV�놡�7U���ȓ<=��;F��mG�	cn(,�Fh��u��R�LD:-���;WjB|M�ȓt��e ��H>dFTk�'��x�L���$U
�U#w&�-�+Kt��,1�)��$J(N�Vh������9�V�a���A�}z�J�R(:���o�(����uV�����*L��ȓ(��h$��.H����c�b���RI�	�N.D)��@]�?�B��ȓ 1�gkS�s4���恕Y���ȓY8��I�`�.4�@H���'tNم�	�=����M�p��|����8R��)#���6b�B�%z}v��s��D*ve���Z,O�B�	���uB�K,(V$�(V@�B�	*ct��!&ƌ'_�r%��/~B䉼!��=��Ġ0��1$���I`B�)� T`pqbU����B�InЉsG"O^���ċyS�a*�/JFh�]��"O�m�pƚH`��j�m=J]0�"O��
sn�d�
�aE'�Qc"O�P@��+�����I�M	�yz�"O�p)T�
��  ���#�2�
�/OB�qO^��ç�`|����2�6Q�C�u`��(�����En�<�2�'k$ܠ�4�ۓQ�&��oضT���'��IR�	�0m��ᓪC�J=��Oَ\N�4B ��z��I�|�t�zR�Q�@���S�O�"�yt*M�wn��NGKO@����G����a���tP��4O�?)!n]?s����C�{����v*����;GJN�z>v����i�L��Or����J�L���P�'%�U�&H�� �ܴ�V�����8j�� a��>��)���2q�D����.�����*��-j��(��˩�?E��DT��dʕtquQ��>I��IU��0N�^�IG�O��	�'0wH<�'.�R6�QYH�Te�0vJ8�7�[?ys�&*����)EZx��	؅�F��!R�^h�B��7*��Y�LT�a ����O���iF`�)o�����W�}���r-f$�����+^�~1�'̎��0|��&O��$��KG.�V�����Zo@t�4�"{�v�:�I:[޲���S3E)h���U	z)H9c�i]>(�x1[�����Q'u����çz12t���M~>��Bn9F�v�S��x@BJ9I�����OA>A�DD6ސ�2gi!j�+�'�Zp`����7�$�ǅ�f(fh
�'Ǌ���C��p�Ҧ����8K
�'I��!%G&z�0�E�.3=s�'�\����4?ld"Cc��#r����'_B������lh8"ʜ=K�Y��'b�]����'N����镎EW6�c�'����Ū�;&�ˆ��?Bq�(H�'��в�Fr�E3�Ǻ5t��'���*@�$ϾX8��4s����'Î=�I͎10�d	U��ʐ�'�=��\+u�q��ڶj<ة�'���y0�	�_j��2T�Ӥ�`�k�'�d���A�5�t�#"F-0�ܣ
�'r��r�OÀ}�<�#È}3�t��'��Ġ爋�RB�<�aM2t3��[	�'r�D��H\�� ��.�n[0}x�'��]АbZ	R8n�
��˷Y#�=��'��P8�̀>g�2 ����6Mn-�'�l��k�OU�L� F�x7���'@p(�W!?� ��g�@ l����'�0
��S+�h�*�L�&8g�j�'븘��EͻN�;viҶ[��Q�	�'����& �+܎E�UnH[H����'�Fd'����@22�ȶZ*��
�'��@y3K�9�8h�1 ֽB�<���'OR���R���HR&˗<N  ��'I�H���V�%�a��9C4P��'�p��reɉocD�ɑ��=�@5��'����! f��Q�!I��*�j�X�'����gV"m�t����Q$(-�� �'� ��2*Ϋy	~�X!gH�1/T��'vF���b�8#��ː��6)��y�'׆� V%X�o�D	����12�QY�'DsĦʖ}9\BG�As�����'r���&޷|��yS��Q1cp���'G���q�M�r>��Z"+&&�����'?�x�5EZ�Av�Y�d!��2�'���JF�S4xC2��lf�S�'K"��D�Ѽ*���(�,(lČa�'`���g�S�}$�
�i[��Q�'�d4�e��(b�� �a�5MOJY)�'�TT�D� 'Ɋ�CI�<L*���	�'��W	H2/�& QcM�U}j
��� ���]�$]ֹ��g 7*�hy0"Ob�C#�=�Ɛ�fZ�0����2"O\�����(p��Q�BE�?|���p"Op����_ϐ)�ecJ*'2��3�"O���V�Q��	#Bl�@!ʃ"O^]KW���4�H@Rq���"B"Ot��$-IR(b@��ꓠo�b5�G"O0��҅5}�h0�O����7"O)����|Yq0o�	��Mx"On���(ګ&����'P����"O��2e�ܡ�P�Q�n�q�*��U"O �^y�(m0bm� ����"Oơ�㄁5  n|sT�N�U�~�pP"O��+�bةJr@	pN ��d�9 "Od����2
&�E0��G�4� HH�"O"�Q1��B4�-h��&E�pd3%"OL�"#���`?d��A���f��t�!"O�kg�a��IB��9�RdS�"O���0/�#a�����V�_]���"O2��e�H�>�a�G�ʂ}J�� "OleH��@^��܁§�./xh��"O`��ɸ86�Hq�'��4���F"Olv�N�
�q	Y�35J�"O����IH
d�G)�(���"O2 ���V�Y �g �U����"O��JT��bFq %h۷E ��"O�t�'GH�&��0���Ч7F���"O�I�I�y��l�L���I�"O�l��J� �*}:a _TNI�"O����=`���3 N41G`cf"O��d*��9��؆�(*L�+0"O�������F`N�y��"O:uP�ʆp��t���5ɶ�"O��k��_!�!��Nc[�廖"Of�BEf�M�� ��g�<I�)��*O�
P���gj�C(ĬP���'�ޭS�̖+<7��*E�T�h�Ԝ
�'@B`1Q
�����$.��e>ly
�'�&���j�P �7J��(�r�2�'A�<gk�yH-8��� (����'v2i�5C6�{vk:+�Ű
�'#�ЋT�ݮ�V��$H:<�B�ɕ)Ύ$CMQ�
,�DȊ ��B䉅t�S�O�7� "��)G�pC�	��L���.��3�]�(JC�I�^2
��&e�x��o;1xC�"O,�Y:!��dH��e�7�B�	�Ed�l���P�#-����*6>B��O<���ㄓr�6�p�N3	�B�I8�~=�j�+G���C�	�-�Q*%c��4����LwzC�"H�`a[�9�&AnN��zC䉞`�̝
��еK�V��g��>sNC䉿n�P8�-[."�іK6&�(C�ɼ&��  e�F�\c@�"�Aw5C�	�d��(��C�|A�b��^�,A�B�I9m����J�#Zf�p�g! ~��B䉯j}�` nB�����&R(ԦB�396��c5��\Yd)%焐uX^B�I�R%6�[&���G�@i!�aX�n�vB�ɦ+��ʢ�	W�@��$��jb<B�	���r'ҡiD2U��FU!4�HC䉤e��̨���O_���E��	t^C�I�y��&m�01�h��Gg|C�)� ���0�ϴ[��T�7��j�<c"OVq�C�J�[XZq$لܨ��"O�1��_^7��y�I�\�
��"O���,@l�8�"�?7�p�4"O�S"*5^Z�0����t��Q�"O��)��Q�v�|h��"_�K�h�v"O�9���b=:�����v��9��"O�$�RʈB���BH�z�R i�"O����FD�1�Z� `x�"O�*V�̔W���B�e�Ջ�"O���Ta��l��$�Aפ+�Ȉ�"O�<a1�W�5� ��E@V c|P�"�"O���2�_8H�p��mRdal-W"O.�q'��50:š0�ƎvU�-K'"O�⒍C6
�^M��.͘3M����"O�1�R�k���K*Q��X�"O���L_�$���s�P57"h ��"O�9tG�C�>� �'F�\�&��0"O202��.��X��gCu�h�`�"O~�pg���ж�G�
-x ��"O�Lh����j_���s L�w6\�q"OB��RAY�E�4���P8��yA"OͲ!^�,ZqIc�Ĺh��"O�� �F��9PI
2�����"OT\�BU
�u*Diß*�6��"Ol���EhL�S��G�t�[�"O.��'�r�V,b�O���ˢ"O�Հ�P`�XyQBo�*�"O
x�Ed �1��ajg �=%!n���"O�H
S�0U|V���Ů{K܂�y2D��a`)!��6�D�8 ���y��ż%&�8�Vb�0��I�c�L��yb�
��X}�(��)L��hf��?�y��Wb
F�����+�b�9V%^)�y�̟�a���MЖY4� a����y��;��@&°O�5Z �V��yRm>O�h2�	�p�.e"%�y2�
1Q4L���CS!��yċu��\r�IT�A�@Lړ���yb�FY�B��wnK�$�
Q� �1�y�iM�g*Ȱ��ϕ�M� Șv�_��yRI�p�m��E�F�ha���y�I�"&�^A���Fc��[T��y������>�P�y�I�y2N�u�>ܱ �.f�Ȉ�2��yRќ/4���ǗR�0�� �ӿ�y��݈1��(Rs	�)@��]�:�y2M�(�	6 �?(~���U$� �yb�ɗl��Bc�ȞL$�bg^��y2�	10�L)ɣ��K����D��y�	 :x���6K���[��yBiTAy�nB��*��.�<�yR֕4�"x���%{�d,[G�>�y�יTI����Ĺ�F�[:�y҂�e�H���X�MQ�l	�g!�ʘ��iy� C.tdn$�7��f�!���oDųvKt]�YJ"��C�!�d��|�p�%�W�mP��gG9e'!��P7�$�cO#{��h��DS9M!�d�@��ٳǏ6��\; �?!�١c���qA�W ����%r!�$�&r�pr��)|���ҍL �!�D��Ǩx�@Ia��M��B�-�!����Z��$����,QƌD4I!�� �x��~�Nx�
O��2=b�"O@��ffO�ji�`���������"Ob��7L�!� 	�jH	m�t���"O�� sߝX���2�P�<�Y:�"O����R$wپ�
�IT�j��;2"O��[�+�0��ٛ @�2��"�"Ov%b�/l'$4�r�p�"�R�"OBá%�(�թ��@�d��0І"O���d)���Y����#"O�E��윧Y�
��6g� Խ�3"O�t곣��>�����,H�L��"O�J���֙�tj��`�n`��"O4��u-�@N͓fi�=t�P6"O��i�ʩe�d� SG�1rp�@�"O a�G���;n�0"Ve�?T�#�"O<�5������� 4��Ȩ�"O��B2,V$1�Rl�4^�B�	�"OB�y#oP1N5�Ě���U��`	�'�>�"4���k�r٘�	�	;;��q�'��5��!���=җN� ��s�'�<���I�����4@�L��
�'(�����H�����A�����'����i�*Q6����@Y�'�}��'��4S'�GT��ض��wa���'_
�"  ���   �  >  �  �  M*  �5  :A  �L  6X  �c  o  z  �  |�  �  w�    �  ]�  ��  �  J�  ��  +�  ��  &�  ��  ��  �  W�  ��  "�  � p E � $ �* �3 �: �A �G <N Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr_>����,�	!K\j��s(ԛb�SL�D��Iʟ����	ӟ �	ҟ�	ß�ɉr"���bM8����R8,�I埨�	���	�@�I؟�	Ο�ɦX�\`x�aZ!�p}��$Et���IҟX��ӟX�������$�I柨�I�lT �(�P�`뤈�ƆC :�Iޟx��۟����,��ٟ���ß��	�m�R,���1v�\9C�rq���	��d�	ӟ�����D������ʟ����^wp�I"���i=*�:4DZB�p��I՟�	������@�	ҟT��ϟ���IP�]����X�|E�A�	�-~�����I����ٟ����,�	ޟ��	���|�/�̑җo�>8�)���|��ן\�I㟬�	��H�	Ɵ �	��n�`�#÷_8"�����9H����˟�I���	ޟ��I���Iß��I���`ūR�5�v��ՂH�zq���I`���P�	ޟ0��ԟ,�����Ɂ+h��A��'(���DT�Yn��I��	��`�	ޟ��	�������ɨl�49��+]�Y1<�C F: CR��Iܟ`������	ܟ�������۴�?���Y}f�å��/;z<"�b�g^HJ�W���	Jy���Ov�o���,���,`Ԅm���
��N�Y��"?!r�i��O�9OD��H�:D
��Q�^b��P�^���OlM�Q�e�D���d��*�O�^�blG�\m��BR�ӟ�t�yB�'���q�Oi���3N�#�`ґhW#:���b�&��E�-���M�;y����DKӡ �N̨`��D�8���?��'�)擾�IlZ�<��b?*����?%{P��F��<��'{��$U��hO��OHi!�ؚ�
���N�5����v5O�˓��A%�V�\
��'��P#΄82K��ʋ�u^d�b��$o}"�'�;O|�2B<CEfW�Wl>� G�4�~��'�b��` @����d�Zӟ����'��<�&��1Q���dc��d�����Y�@�'���9O6��A�Rv������B��I�:O��&;V i�O5m�S��|z�>���"B��uz5�@"�<����?1��c� �ٴ��De>�@��\���H�B��.&H��2�0�&�>���O2�4�V���O��D�Oh�d� J'(Pz"V;� $�,R2�t���OK�̜&��H����O����A�3?Y�B��~�a G�|���!���?��0���a�f�m�k��D�O���fn�hҢҘS[d59w�ź<�lt��Ǜ�L��Ă�OL��sF7Lx��J�tݱ�M<��^��±D�r,ݐ���`x�@��N�@�Iß���ʟ�Ky"�q���b7��O2M[W�fT`�E�i=F����Oimh��T�	럤o���Mk7	T5 `P�J`I*6@\�5 ��"�Y�ٴ��D� A:�A:���������A9Y�P�Z�����gΈ���$�O:���O����Oh�$7��h��qJ�=Y25���چ4\\A�	ϟP���M[ת��|���Cu���|��D�7(���g҆BcLE"6N�4R(JOƝnژ�Mϧ�Zyc�4���ŉ�� Iʵ>=�p!d���e��P�H�?�?�Ӄ"��<����?����?id�V�*�pQ��:;>Z�R���?����٦Y��.�ly��'���aF@����g�����ڶrm �@����M#$�i�bO��`�5��Ȟ:��};p�Y�1������>�ec��Tey�O3�����S��'�j��?}�t�4̋�[V�8�'���'�"���O��	��M[2a�k�ʕ2G%�,s�J��ʕ��$�����?�3�i��OԵ�'֛��2&�|\�tj�TX�Lq� �.vql7�Ϧ�j�ۦe�'�x4����?YqsT��Ps� �3{� Sn�\%�PRB|�H�'g��')��'��'���B �mZ2�͈�s�ʍ��[޴5��	��?������?)ǰ�y�ˆ�4T�:�i�ҁ�'i�_�n6�ʦuJL<�|B����MK�'R���:t&z��aO
1n[�}��'. �A�×����|�S�D��ҟ8�QN h�NqI��Ą�ȴ�5˟(��ߟ��cy��s�,(Cs�<��yX�d��(D�h �KZDO��O>y�A����M�Q�i�xO"��d&I�4_�� V0��T���*�@���Q�b��v�&�2��D�RiĂ>�x8Ȁȋ�~�� C̟,��˟h�IßDE�d�'�VP���I����SRŤ��7�'�@7-�%VQ����O �nb�Ӽ���o��3��ِW� �i��<�7�i�t6�����Ō���'�&ih3I��?������F�.`�!��ڌ��'c�I����ӟ��������A�ܔ2�O�h�z:�HMn��=�'�>7͝� k���?YM~"�|�����4_6 �h�A���5C_���I��$�b>� ƫ��RKPi�CE�W]B�p�&�(N])�Ty���$�\�ɒo�'��	(u��)��l�Q3W�Y�9�*���ڟl����(�i>A�'�P7M٭@����$�R�`M�/��eBAZ2�h�D�ϦM�?)S���4Y�f#r�҅QP#��H2��K�
Lն�0��V�Zn6�(?����{b������'��� ��{���_4F�
�;<��PW0O���O��d�O���O4�?A���F1W��M3TΒ�L�$}p��ş������޴;��x�OL7�6�D���`M��$V��
#���9���O����O�)��>��6�3?��;���i�%�������|2�i�%ǜ��?�A�6���<��R�D(;���#V΅�_�����U�O��oZ�D*�(�����I@���ѥq��ÇB�P�B!i�c�����S}��'�b�|ʟ�%� @�bΤy��M�)3H:db"�X""fy���]����|"Ł�Ob�L>9�kGQ�|T����	SuC�l�~<	�i�xUj���X�`�����ݒp.�v���'�7m2�I�����OqD�ϸ"Q��� �-t��a��O����R�>7m ?��+
Y���(t�A<ڔr6�ܥ#��Q�ah�\΅���&|Ox�R�L�Tw�ŪP�p~pec�@���)�����<�	���:q��yW��3=�\���l��?:�MS��6S��6-��-�M<�|�	��M��'B<a�#g����03$��&G~$'vֈ��Oɟ|j|�Z�4��ܟdX�*O�A5�@˰�p��#`�ן0�I�q�J0f��zy�$o��X��������Oz�# N�9KjUb��]5;F��/�O�ʓ�?y&_�ě޴�r�xB,B�(Y ���,ߓ��J��9�yb�'���Q,	!�����X�h��7&�B.C���t �F����ĨrVr��n�ܟ��	��\�I��4D���'��p��@2s�x�&�T�Z²@���'��6m��`�d�O(m�}�ӼK�\�Ta��MR/g��R�eI�<I��i��7����A8҉�ݦ��'�<iE��?���FP8�:bR�UKB�kT,"$�'N�Iɟ �I�D������
n���8D
�0œ� �	W4T��'N�6-[.�J�d�OR��!��9d��hW��\����6!��1�O�$�O��$�b>}����r��Ձ�.Q+�]�6��!z��+��3?�&-]3K���'�����Р{Er��f_%$=؀�*��4�L���O~���OZ�4�>�.�VMW�l�o�p{2@�F�gT��D0�y��b����ɨO��d�O��oڐo��щƯyZ�-��� ���	������'�F,�v��?I�}2�;5��9Bǉ�R9�	��A�B��?Q���?���?�����OV"JC�(Ht�`Lq�S�'���'��7m����'�60�$/
�CG�<S.Lba�0LB�&����4'���OX.Y���iY��
^@$@�&&P�Ub�`M¶g��x!�FǑhe�%L�	Qy�O���'���:~��m�:+�|�hT�[����'���<�M����$�O~˧B)�Y��	�48-�R��]H���?��S�l�I���'��K|P�k� ��萰i�W�����G?G̦���JI��4�>9�� M&�OB� ��)E�*��4n) "�OR���O��O1��ʓsf�vJ���)�'#��5b�1?�pI�T���4��'/�˓�M�����)2��p5`Ns�|��!�;���ef���K�At�"�,3>����b�O#\T�w!޾{ Xѡ�C�1���A�'�	ϟ��Iş��ş���f�� Eצ�Q��(�Lԋ� �dO�6��6L��OF��!�9O`9lz�aq!i[�B"	��N�/+6L��d�����Ş7�ڴ�y�@��L��X�D_*|iC�Ї�y�@ț%_���I5D��'Z�i>Q��e�~�SW �c�9�æN�X�>��I��$��ğȗ'�H7-�,�"���O����z��L�Ң��|n�Zш �& �lR�O:���O~�&����.+o�(����K(/�Xg�&?�ס�\|�� .�P̧W~���Đ�?Q��ȯM��9	G�?z��Q��MK��?���?���?��9�0T�F��XG��ܬ*���&��OvTlZ"���'�67-&�i�ը��D޸��١EY� �|���I֟������m�B~ZwN	�p�O{�d�T��'��Eh�!�1!��d�t�D�	qy�'\��'�R�'
�%N8B�z�A�+�(E4��Q�H�^�ɾ�M��D��?����?�M~��L�j�c�:���`s�9�%]�����'�b>%�e��:HN(��� m��#�T�p�� �py2��"~1TA�	(��'4�	��e����$k��y�K9l�\�����H�	̟��i>U�'v�7�ΎJ�v�$�	r6|���M�*+�d��eeV`�f���ڦY�?�EV�HݴId���d�R�ƎW�s5���X�Q�h;CGQ���7M(?ᣭ�^���	=��߱p�$�
��5F(dzdhZ�Ol����ퟀ�����ڟ���v�W0�R���;�����ˋ��?Q��?�Q�i�(ؚO�R�p�`�O����W9a�q�g㗻b �uĈX�����mz>%��$
��'M�,�q�'��eR�!}x��"��KV�}�	,,X�'S�i>���ğ�	�x� d���M�I�.1;��c=�Iҟ�'@7�_u���O��d�|�&�K.p]�r�&a�r0��.H[~�,�>���?1�xʟ<�yS�"�@�� X	
�2�����Ud�0�o�y{�i>�r�'�� '�T�F�B��A	��
5 ?|Q��k����П���˟b>�'�*7�
5eB�����(^n�B+�(q�0�AF�<!źi@�Ov��'���)e6�)�AL�`�P%
A�3�BAs����eӪ��f�y F��π ~p;�H�$L�@䃕.��"��5OR��?!���?)��?����I���YP�K4u��@�'KuNX�m
t�hd��ܟP��[�s�����w�(�<d�%	�R�0`qP)ّ�?�����Ş�z��4�y���2��vM̉0�!��K��y.�7j����� +��'���� ���j\��Hso�*�(@��	~�:H�	ş����ܕ'RN6�ľ9~���O>��X+4 0�8��^
G�U��m����+�Op���O��O٪/ӗ!c�5���I�&�ra��PkB���)������s�S�(�R����W �8��IV�ȓP�Y�������IןxG��w��S�"R07:Zec�G�C�9B'�'f�7M
 )-��(���4��С��K7B��	�ǃ�q��� =O��d�O8�d�H6�7?��\ޡ��'˺�ʑ� p����/l���U�"�Ļ<���?����?a��?)��;+�`�d(_[!�\��)�;����+�ǒߟ��֟x&?��+0�y� �"�^�K���3�r�p�OfmZ5�MCR�x��D���p�X$� AH	+@-��X46cld���7Z�I9bK�����'	�D$���'w�=�WC��G����C$4ڔ��';��'cb��DQ��8�4G�Ha���k���׬Ҫ�bP'��;�Ԭ���4Û6��^syB�'�F�~��q��EvB8����V"K�|QJ�^���6�&?�EiN�t���)�����stk߶Co0*���G�\�% ��<1���?!���?!��?y���aš�%B C��2X�W�X_��'>��jӊ	 �;�8���-%� x �N~A!&���'���t������?���|�7�U:�M��O<�cg�}� ���h׳z�<Q��R>�,�������O*ʓ�?���?)�l�RѪ�j��/oҖ/x_,	��
�����	YyB�bӌ�Q+�<���IJ�&]�Mǻ�B]�C�?n��I�����Ot�$2��?5*F�P8RZI�g	ɟ/���֦Σb9�gD\�z�~ܔ����^ПX��|b����=��F80�C�Ծ8���'iR�'���TW��R�4> ��P��$���BR
V�1���A���?���m�����Hi}��'N�S���c" #f�')"`���'��6M''j6�$?��O�;��	2��fI�~����B#n- H鑭��y[�������������ß�O�.� V%�2M`�(�٬�xٳ,{�zp+W&�O����O �?�y������ȠPc��3��vCp��0A��?	����ŞS��ڴ�yc�;�&��g��;^ɀ���D݉�y"k�}ڡ�ɝl�'�	����	.aGp��Ƀ
6�90��A��d�	ȟ,�	ş�'f66m�+�,���O*�$&l� ���&LȤVE=�㟼�)O��ds�D$��꒦�Y.�(�,�Y�hy%�'?�Q�J>x��d`��Z���'v���DZ�?q�fN.��kC'Z ��֋�?���?���?y����O�}�f��L��څO�nh�Ը�K�O�umڹ:����	ן�ܴ���y��� n�s�n Anp�?�y��v�inڐ�M�r.�2�M��O��0��X����E�-4I6
Z��Q��%�29�̒O˓�?��?����?���>��B� �����FF4U�*O��n�0.��8�	ן���I�Sן8��*��V�\]a׋�G3��kq*S����Z���q�4z/���O�t�J�G_g��d+�(s��e�%���3%�Aɕ[���7L��R%�|�	_yB ��tp(��MB�c�ME��$C��'��'�O6剹�Mkc�?	qB�)ErM����Tۀ͂��Y�?	��i��O��'	�'"�$;��e)֣�V��M�EE��j��1�i���!�)���OS��%?u�]'2����n9�n�H�S	,���I̟���ğ��I���	v�'P3��t��`��9�̓�o7` ���?a��`��6� �剗�M3N>qУ_)�H��Z*_ܴ��'��;���?���|jDHT��M��O��T)T2�H��+j���bSE� k����c�O���L>�-O8���O����O�X ABFWd�O �S�
�	�/�O�D�<b�iI���'�'0��'�ӖM���|��E����m{���OT�'[�6m�榉`O<�Oq�U� ��Z�%��%\_�D4�&��	�d�뚡��4�2����D%��OʠG�6�B�+��_
1�d���k�O����O���O1��˓���̢qyP#\�t�ٳ��
�
�"�x��'4b�x�T�$@�O"AnZ�m9��B�"��6�����%/����4_��v�Z�v���R4+7���wy�I�!p��a�� KDu�ЎU��yRW�(����@��۟ �Iԟ̗O�vݛ���2&@�;!h��u��z&�~�����d�O �$�Ol�?)8������/'	�Ѣ2���a�ʄc�h��?q�.����O*m��i_��3�}Ĵ%8�J�T�D�$��<YFP�X���dN�����4����*d$��*tH��ˁ�D�::���O��$�O��G�&�Q�$R�'��f�!R
��# 9�ysF�S�=h�OvA�'���i;�O��0�ݕ( ���%�0	z���`��f���OF� x�ԟ�YCL̝.j�d��O�|H��'LΟ��	��0����D��w�D�.�9w��k��,H 5�'�>6-�w��$�Of�n�i�Ӽ�P��U\،�T	_+�H��A�<Yֵi�(7��妵j�*N�}�'P.���h��?C� B�P��}IB|�6�˥+-�`��B-���<Y���?!��?Q���?�Pc��u���\,���g�>x�'��6MU>)�˓�?�L~���!4xƎB�W��U!E�
�|��S���ܴp�v�0���4[��k `����"U�_¤u�e�>w�˓V�JK��OܑL>a.O�X�ÊY/2Ά���@ŮY�Tt����O����O ���O�)�<1R�i�����'W����lVb�����N��t�T�']z7m1�������Ov6����*�([�(�l�)�h�iT�x!
�t� 1mZp~�>��<�Sp�'ڿs@�E�$*������}�$s�K�<A���?����?i��?���)ۼE���y#i0�
�����,���'�bji����%�<iP�i��'�8t���3b�(��
W�\�0�#�$��{��|Z�ɜ��M��O�q8���]Zm��ݗ�h��)Ɖ.^�����ؓO���|����?��7��)Q�g������qI��R��?a/OJl����%������Ix�$�P�w�Tqy ���;g�Ѳ�Ρ����V}��'�k5�?9�6?k�i�OC`��8P�^#k9Tc	Wp����|"���O���K>���i@F��qH_�p��v��?I��?����?�|:,Otxl��F.B�j�+3q"�s��J�E�XK���8���MK��Ͻ>��
f&�1�	�Y��W�j�������G�f��6����$�ϩT���~�w֩1��|طn�51\�S�hC�<1+O����O��d�O����O��'�p�{-�R\�O
;Sz�M�C�i�jI��'���'5��y��n��� �*�� b��Ђ!ԈD�1�����H�4{���O��A��i$��#`iA���;]�bJ�eF!>�d�i�����s\d�O���|J�F�t�`�IH�.�Ȉ�V!�Q�@1���?!���?�,O�Uo=0F������I�g�J!&�	l�|�ʡEȄw��	�?a^���	���I<	�N�8�c�-��YRi~ǌ(J�R�Т֩�O�V�	�i��ڋ'��0S%U�Nu9@g�?h��'l��'MB�sޡs��ݫL6዆&2����W����4H|�a���?��i��O��K�x� U�)8D���i�F�2���O����Ol�Gg�"�Ӻ��Ƙ.��g��a��gJZ�W���ե̖jS�O�ʓ�?���?����?)���2�p�T�Q���0��;^D�)O�)o��e����	̟�Ij�'qu����
�%��Y�%��B?�	�W�ؐ�4N��f�'���,�p ���rN��.Q7�!��Z�R�ʓFe�!� �O@q`H>/O�-��g��H�lś��אg�����O���O&��O�	�<�ְi(�ۅ�'�܅���f�h���B���4��'`7�>�� �����5[۴u��̅�@tuJ�Œ�L�P�0��"U��P�4��D@�z�:1K��_�����N�	h:�������#�a��~b�'���'�R�'h2��o��Q��04�� 1@ �M���d�O��Ąæe���w>i����M+I>��(��m���K��H���-=��'�67��˦瓫/��n�q~��nI 	�����z��ژ5�U%�џ�Ё�|rU�d�	�L��ޟ�r���D,Q�ƅ�x��(�c���X�	Zy�fy��d��O��D�O^ʧ�^CfC��f�<��Q:#��D�'RJ��?)�4e4ɧ�)�9�T���R�g�X�x����)m�a���!\^�P�ʼ<�'l�~�䙫��}��"E�H�y>�b��Ԟq�(|���?���?)�S�'��򦹱�H�"�~���V�_H i26!�5I��%��ٟ��4��'�~�K���A��?��
bC�QB.�A�D-_�7-�ݦ��E��˦}�'����?�AsW�X��	I  ]����p�T�k��'���'m��'���'|�+�vTQ���4L;] @��S�ġ3۴Z' P���?Q���䧊?����y���G�(媔��7؈�y��S�^���'�ɧ�O�zH�V�i��dR�>�,i�աGȼ��g�A�󄒖sTlY��y���OR��?)�������I�O���� B`�T���?����?�)O��m�51�j%�'2�-{-<X
�l�>bVp�@�M��'≬>i��?�H>��D@./Ʀ�[7�K�*�5b�!�s~�n��&��5���Þ\P�O��)�I�\�+՟|;H�X�̓%1�D�i�2�y�,�="��@��ھ�X�
.�REu�8����O�����e�?�;a� �t�дAG�,�qG\�����?1ڴu�V�M_����Ĩ�'̊J��	�#�p��uA̖!��� �O�t��m%���'Zџx��mT Ux�$��Ǝo�& �!=?y�iS8�� �'_��'��d���<��p�Ù3/!MS�Ryr�'ϛ�(:���t�J�VP4-F���t���ɬ"�)؅հz��'&)
���'��I'��'J�Xp��<t�h-��KQ���E�'���'���4X�#޴ � �r��W����U�@:D�ѰHK����`��˛F��Vq}�)q������������v�ӓ'A;��Rei��j��xm�@~2J����I�S�:��O��!�0�,�VD�*25�bB��y��'z2�'y��'�2�I��*.��!��K k5���� }s�$�O��d��A��On>!����M�M>Qe$�k���N0����T�UD�'@�7-�ş��Ƅ@|�7�'?qe$�G�? ĩY�KF0,��q��	�|�"��s���?���3�d�<���?����?�EZ�$���"�%
n�jT �7�ZX�����d�Ҧ�@�ޟH��ǟ(�S��M��%�ip���P#h�6���id���I���d�O,�%��O�����#1���g�œ=���L���}�X a0T��S�\?�B��&Uf�����GK>���@�[�I��H������)��yҍ|Ә,�P�
-@D���+Ռ)μ JЏS	J��ʓ=�����L}��'U�AI2Ŋ�P�;%N�>n��.��'��D�e�i��i�KQ@��?��U�D��h�;oB4���������z���'��'���'�'f��=D�h�䐽��]�sH�/;��%��4%���/Od�� ���O^�mzޡK��P̺�H��N%~⪡y��ʟ\��O�)��-oZ�<Q2�%��hÔ�D��J�D��<A"��6G�@�D
,����$�O>�d_�i��X	0.Hp���CߢS޲��O��D�O��?�&cO�8�I����5�� +��9��ʞ�D�p�CTz�	ܟ��O\m<�M���xrC-!�����L8!��ק^���$ߙGp��x,[=B������@��@�l�D��`a�=+�q����=V��$�O��d�OV�d%��S�.DK�(t��D�f>����m���?�&�i*�b��'��+|Ӡ�O�9�*��ł@�[�Uf܌s�B 20O����O��D,Obn6m+?��^�j#�'[,:��%�˨G�NU���%x�H���*�D�<���?���?����?���ȕM����2��B\��C��[���B��1�Ԭ�ҟ����@%?����g���ɗ ^֜B�A4_�,�
�ODlڹ�M�ƛx��$l�nh �$�FCX���� �*�҄�c�F�t��Iڋ��?�n<�d�<1K��.ѷ-˓���$R��?���?a��?�'��D��I�#	�ПH�3�D�x����
;H�Z��Ukk����4��'n��V���J�O�6T����j#C�d?�!
D� KNQy�vӊ�I�L-��N���ȐN~��Fݴ�B+�"`��P�� & ��?���?���?i����O�f|C,[�0����I��C2�'��'�7�(pI���M�L>�ը#{)��MO�,��!r�I^]��'�l7͑��S�+$,<l�y~«�Fy0ɗ�<l�ԵQ@f�A7���<�q�|rV���	֟��Iȟ�p�Q< �,���:�j��ß��	`y�ohӨ���h�O���Ov�'v)^=4j�U���E$\�t-�'4�'��j�OBO��W����i��@�ִ�a�˄s"�xe�O�3r��
��Cyy�O�����1��'�z�Rq�*Qt #k�� ��p��'x��'����O�剭�M;S�Z&>."��m9W_�ݰ����`����?��i~�OF}�'o�*�;qgr�z5�A�g�i��I��R�'�.{t�6����W�8��剏3��u"�s�wB� �N�	fy��'�B�'���'p�[>]b����[��I�۝{^�d{��C4�M�5EP��?����?�L~�#���w��d�4 :R�ر�v��C��'���=��)�<<|6�r��c4���)�԰'��#�.�vh�ěB�	zE��a�IHy�O�Bl��^"9�"�����T�g�!���'���'��I��M�rF�?����?��m�jq ��� D�ˆ��O\��'��'�O���J� @���f"��g�<�#W���Qu��?�΁{�N,�>�BN�ٟ��!&��j�Us���m	�I���I��|F�D�'�l����h\ɳ��YG�$%�Q�' �7�RS���8�f�4���H6�c�U��Uf� �'��<�ѽi|�7M�٦��E����'��x@�$��?�G�*BQ��k�� ��lCSg�S~�'��i>��I����I՟P�	� ���kW��z6�Ջ��K?6pD�'9t7�VT^����O��d/���O�T�pB�rd��흯NC��N&g[�Ɵ��	W�)�iHY��CQt�a�mZ�d���ZW"^�7K�˓k����V��O�,M>�.O������|��xb̒.D��)#W`�O����Ox���O�I�<�G�i^�#��'{йz1h���dz��4t'p���'z6�=�	���ě�����M���,R��)��I�Ą|�c�ɧ*i�H*ٴ�����b��4��'p@�����[��U�ȃ:L��e��k�����Op��Oj�$�O\�D!��� =��`�'��D���A���� ��4�Ms���|Z��MA�v�|bK�����/�3sx-��&Q����Oz�q��)6v��6"?�%�?MvVdTTbU�e)��2M0�
T��OJ�yL>!,O���O���O6�W`W�b�lz�$b�n�׊ß���Fy£w�(�E �O2���O�ʧn3�����N�E<�8���$����'d��?��m;����P`�P�҆V�t#J��蚇[E�TJZ�In3G���Ӱ3���
i�	�E
z��N�*��Lі,N �����՟��ןX�)�Ry�xӾ���fC�H�<�'jķvYP�a�⁕&l0�Xћ����w}��'!D�+a�'3��Hs�(��p���i�'�7��q�6�2?��ȘKF��)=�T��!T�Se8��L�U�
�yrU���I����ݟ�	�ܖOT��R��{aD)s����P��2��|�ʡ�d��O����O4���č��ݡn:!�����E�q�0�	�%�b>��e�⦽�S�? �ih�C�*��!��9�$Y�6OP��CmO��?�S�)�$�<y���?�
�$XRy�'B˹kJ�ygې�?���?1����ċŦ	0��៸������E�	����'́Ih����)KR��?��I�M��i"Ox�`j
�i����U�_oh��T��TQ�ʝe����wI�}�d�"IJ�H����0H� Z�,G':J�Sj�����I�������G�d�'�"�"��+�L���𩅢�2��+�l��L���'>7�.�i��dIH��|a�'ƢBL���a������"�4n�@M0ܴ��!l����LB��3����<���atȚ�u�����,���<ͧ�?����?1���?��¥ ��d���r"�8y�C���P�x����	ß'?�	#&N�� M�mȚ)г�"nM�O��D�O�O1���1��I`|�8)e�C6`�S��ό�Q��<��bG�8�t������1x� �x�h��
c$�u�_�d���OR���O��4��%�FK�w��E�.�bls5�>-�i � �tY�gӞ㟼��O����O�Ll�B��QY�M�3MY6Hy@�S��Wc^����' @$0����?Q�}��;|S��`T"y�
��! ޴$�����?����?a��?)���O�t\�R&�H� z��[�\�Z�s��'dR�'l&7-�y�S��M{K>apĜs�,AR��8fy����*5�'�t6�[����¨>�@6-!?Ap՜F@>\9 �&6�1Y'��cֈD�T�O�`*I>�,OH���O���O����E�i=���c�Y2���b�O,�D�<yҺiq�"�'mr�'�sU�'��.|�6��d`Ƞ]|�d �OZT�'<�6-���'���H�ET'(���"�(B܂��������F����4�D�;��x~�O:��U�W	y[�<�M ��� �O4�D�O���O1�Fʓmk�FMχmB���&>��a��Q�x�|y���'mr!}��� :�O�n���،I��\$|(�1kY�L¤9�ش0+��oʕw�ƛ��Y!�ܣ}/�dk�Zy���h�a���>,���sF�"�y�^���ʟd��蟬�I��O�R��%C-ngR�!c͚:" �x1�lӾu�խ�O����Oܓ����S٦�]�mŞ�����2<hV��b�łq~�t��4F���L/��7-b�0$ڵ	�8��$�zt:�`�&o�L���S�aH�CZ��oy��'���?����	��,Hh��� <��'���'���MGf��?���?���ٮ\l��(t,��o�t�ˆ�ۯ��'FL�m�V�xӺq'�����c�r1K�JiSP�#�<?A��-����CD�$��'#���䕤�?���ܨv���U'�)2(�7�� �?���?Y���?Q��)�ON��]7�6(�$I�*�Z�bQg�OTMn�G�&��	��Zݴ���y���!U��@q� ';'�8ʁ*�'�yBDj�.lZ	�MkV�[5�M��OBࡐÖ���*�Ӳ��O-/�P:#�^�%�<��|_�,���l�I����ޟDk�K_;��!��LQ������	{y2Ba�z�����O����OΒ���<
�U�޾2b`8�g�ˈO��)�'t�7��q	I<�|C��z̚�d�J@fhI����V�>X"�I6����b����&�F�Of�B!�H�L�X�B	i�GQ�*ޞE����?���?!��|
*O��l9� �Ʌ 洸���J/P,��� E�Y�I/�M��"�>	v�i 7����y��o��S������q]�TxDN��a9V,lZN~�1@����'��O\w'�<G<�ÑD�9:��S"��y"�'z��'R�'1��I�?'�|s���rNv�1c�&r�`˓�?ѳ�i���+�OZ��f���O�8c�gշQH@�s&3���Э	s�Iןoz>�r��]�'K�Y�Ce��4��|YU��?��"��V�`H�����U��'J��럈�I����	lþD�#�!p�$�G,�.s������Ė'�P7-a^����O��D�|Z'-L�a��k-��4�^��	�o~"�>��i��7-�n�)��l��n�A�U#n�8���̲L�w�LX�V	a(O�	�?q%�(�d��e��ha�/�6 9F�8�	yT��d�O��d�O���ɷ<�Ŷi[����� ,H`�� 4e2C΋k���'�f6-#�ɞ��d�O�1&�F;e@�BCb��#<�å��On�$7.6m)?�;eh�z��&<z�R��� �8�:� �I�6K~L���$�O�D�O����O>��|�tp��q��̈����7�A3l���N�2�'�"���'i�6=�0�*�n��nx�@�j�#����O��d)�󉏑i�07�w�D"u�� �>��CK^�vX�7mv� �1�<=���UX��}y�'�RHk Ȑ�l��mh����!	���'�r�'k�I��M�tD�6�?i���?�@�Z�fr�����/<X(����'��듖?��8Y�'���k7���>�\D����,9<Uq�O�XR)M^yҒ�醞�?����O�=c�	ð�\�(��@ Hjp(J�"O,А���.kL�Q5i�:l�̹FC�OZ�oڇS�$%��џ$�ٴ���y���g�湠U�^*;�l���@��y2�X�*f�i�h6MX�^<�77?�F�͖	yp�)�3)�l)�)�>R��$��㘓O���H>�+O0�?yf�O\.)�G��37U\I2�`~�Kw�Xz5-�O\�D�O��?�zs䖻U������W���� ������̦�xݴ���O9�B� �A�2A߃�(��P,p�j���i	�,d`˓n� BѮ�O���O>Y)O��*�jJ	!t�%3�ꂿ'r�����'Q`7-�������4ڜ��2���"�qB敥5�~���ۦ��?V�D��۟��I�<[�1�G��2 3RT��cL�}ߖ��R'Sզ�'�Zk�?��%��TꀉT~�z��;d�j!y4M��ar�%x$�ߦy�f��V,�Q��Y���Y�YV��:&�5x����O��uZ��8��԰UmC���B 1���_)\/dL�e�8(-,�uCV�s�!�D #�ͭ��B΅ �>��4�F.x��`�eV ]�dx��j�-^_2T"6
	+@��r�̀
�NlB��A l�����	S*q��q�(�&������<LΔ iFH��o�z�)�<�Dpc���x���[W*�:��iac�2X�Ā)�J[�C�Ψ!�@����q�R^@�us�۶�Mc��?���^��t�����Of�I�@��С�vm�}XSF�o�c�x�&D;��ҟ����QS��2 g`���6a[�`�b�
�MK��Jؑ�x��'�"�|Zc�4��ː |+
�I��)��O��B�{��'�b�'�u=�QJ�� ���T�V�A@\�RfM#���?9������DL:an�(�7[
 ����Ԥ=s�?��'���'y�P��3BN!��t�N�w�LQP�lO��ԧ�>��$�Op��2��<���a}"(�(.�К��+Ae}��M����O:�d�O��
�l91��t��J``Q��L��xz����.чR�6�OؓO�ʓ7�T)�?QcZ�䥘�����)kӤ���O���t�q4��$�'|�d�p�M�� �=`��9#  ����Or˓Io�Gx�����,۔7�5(�!*Az��i�ɮ�jLٴM;�S��ӆ����-����g`�����/V���U��p��p��|&��#��,���1%TX�ԅAFnӂ�Ñ����q���I�?Y@O<�� on�q��(��#n+�$�� �iV�����Ο�pQ��k����EѨ]N̔2��
�M3���?9��r��5ןx"�'e"�O�,q�(4YMXup�d�	&KFTcS���: �1O^�D�O~��#b�$�� 
.�E*@l�T�Ul�՟��d� ��',�|Zc��ic��}b6����)y�۬ON�J��O$�d�O��9��,B��@�	�I*���h�k�F�"P�''��'��'&�I�c�4ڢ "~0�k�0�`L��"�	ß��	���'�1���j>�9�*Ю\�m��� (���>q���?AH>y(O~��'Q� �"O�\+b	����1����7)�>����?q��?��AL |���?��'����Ց`n�u(�nC�TW{ߴ�?�J>��?�e�9q.�'�x���i��E(��\�D���If���$�O6�d�O�<cB�O��ĳ<y�'�lu����?1 ��Q�ϟ�: �C�x��'� �*l�y���a;Po��]@���UG��%�iB�'w
h���'�2P���SzyZc-�����OP2�:��,�ƽ�ߴ�?�+O�����)�ݦg_6d:"�4���2$�Y��CT"L��'C�	�?	�'G�I�/F�FO�f@"�	�n�����O`����)��`�BQ"r\�����D/.� ����\��M����?��@�Μˁ[���'��O���a���6��$�}zm���iS�'X��#!�	�Od��Or؉"��N��P��"%H`��%�֦���;AVĺ�O�ʓ�?�L>�1[��	��b71��"��";W�Q�'�̜Aї|�'���'��	 ���+̍?��,1#�iz�t�`&���ĩ<������?��y�Ĥ��d.zf�%��J��|��T�?�,OH���O��$�<!.ҧ/�	̏+��eZ'P�,+�-H3@���&U�`��R��d�I:Wbx�� .�ͣPJX4�d�@���3Z�.��'���'�bY��8ɔ��I�O���i &t\٣#�PC"�J'�ܦ	��I�	���! @��=I$��<tYft�be\6Ț�Dʎ��	ڟ��'� ��D�~2��?1�'n����j����"C [o>آuZ�P��ş��I	
�@����?����>*S��sӬ��\q�|�pr�ʓ����%�i���'R��Or����᪂3w20dL�pZ����I���Q�	��dA'^����O�,,��H�b���6A��A�ߴ%}�(!t�iTB�'���OL�듸�D�֐l jBv�h�´H�?Xj�lZ�a�4Q�?Y��T�'~6ٱ �'9���/B��(iB`aӸ���O��$��YM�!�'8�	ޟ��QU�\�5Ŋ�U��@���Q�l�,�>�LM��䓪?���?�s��j�@S�B��lR�퓬mP�V�'�Ku��>�.O2��:�����$^�	,�A�)��ԅ�>i�����?	��?/O���1��?������S5m)�B�g�J��'��I�$�(�	⟌�Wj�*�D�Z�Љ� W,j�x=1�h�Ox��?Y��?�-O�Lj�
�|�V~�0�!Wb:�LI�d���Ŗ'
R�|��'�DR��$�W��qxq���t>����(ʺi��I˟H����H�'g��'�U�K�p���lD^�A�  \'��m���'��'՞$��')�'W�6�H�_+L�L�� ���@mZҟd��iy`2j�`����k�WM�E#I�C.��J5��f>�'��3e����C��s� .�� �[�N��cf��?X�� �i剡*����4R���8����D2-,� ��(Rh&,3QB�(|>�VV�p�S�T�I|:M~n�Y�h��5��g����%ć[L6^>?�����O���k��i�<�O�h�����D*}P�����< ��tӶtk�i�p�1O?)�s%L�7���Y�ں	o��Y3e��M�����Tc�)zI� �s��;.(���`B!XH�Ԯ�ǘ'�<��'A0������p�Ud*�F� ��-�"oE�Yo��<	uMCy�ͺ~����
�Nb�Ec'�X�g�L�rύ�rWh�j��ړj��?*O��D� �f���#�nDq�*ðZ��)�2N�<i��?y���'��"��U1
]�e�C~9+��.X,����3=(���?I���?�,O�Q2���|�¥ܸ;᱒c��\l ��Ԣ_G}R�'�2�|BX�,@��H��8w�I>K0�}ai__��!�Š����O���O˓?�������}B���L��*�5J�� 6�OV�O(˓K\T�����7U_ҙ�F�[�]��9�g�D��6-�O�˓�?I6��*��)�O���kܹe9`	�H�.���;�!�>�']b�'���E�ؓޘ���	�J�ђᓪ ��YP�F�FY�,���0�MC^?a���?�(�O�`6AOl|$d	�
�
#���D�i���u�dP�I,��'��禁��0|L�M���Ӧ)���!��Fɗ�|�7m�OP�$�O8���w�i>qk�E5<�B��B"�"t�������M{�)
��?9�����:����Ã� �Xj���j�pTcD���M����?��'A4��(O�e�d�����B�	�c�r8慯Z��d�<A�c8%S�O�"�'���;���[�m��K^���c���7�O��a��_�i>Y�	��'���S��,q�:���0
�n��r�w��d�	C��d$�$�OT�D�<Ab&�'HkzY�&KC&s�n%*��C~}�xb�'���'���ɟ�I���(�J�\I���(�'xl(�b�g ǟ��'�r�'5�R��p�����$�;�p�b`.� ^S
�����)�M3/O��ļ<9��?�f��q�}���[>i ��1(Z.lΕ�a�i���'"�'>�th��l�$җ~ǆ(Sh<|�����ն!�No�ȟ��'�b�'#�C��'�U:�i�#�ڍȗ*�)�����4�?Q����}!��i���'�b�O�NU���N�]Cy�U�[3H
PL�>��?I��u�'f�qs� ����³M������Ŧ%�'��5#0�|�>�$�O��$韖�קuW��
嬄1�nW�N�l���<�MS��?ye�\�'*q�D�0�8?�&JF�%��8yP�i��dרwӢ���O�����'�I�9��`P��A����`��eְ,rڴ�t���?i,O6�?��	�(��%$��0c�J>XB\�Kݴ�?����?	�����ey�'�$�r踨Ck��T����ڪ|ÛƓ|RD��yʟD�d�OV�D�5���e�L`ҹ��ʗ�+F�Ilޟ,��,L���d�<Q���D�OklA��4���<��e4��& �ɭX���4��ɟ���ʟ�'�$Ű�V�$�irÇ�.~��!�&�����O~ʓ�?�(O|���O���[���1��Zְ�q͘�4�l)57O���?���?�/O�����K�|
�+�Z��(L*9��#I�Rʛ&X�L�	Ay2�'Y"�'�@Iۘ'�H����)��G]�4���'oy�B��Or���O�˓H�x���^?��i��L�[�=9�� "�z�Su�B���<1���?�y����?��g�����V���Y3t`�4�`1��i��'�剎�������O��IY�V4`���օ4U���v����:��'�B�'��N���yR�'F�GR��^���a��6E� =a��@�՗'��q{�iӨ���O��$䟌=էu��׃X4�� /�a���9r4�Ms��?y��Bn~�P���}ōM�
Ѱ��oY���A�禽����M����?�����FS��'V��#P"��B&�<o�v�Rdʚ*pQ7�c��$�<����Oh&!7D
A��/9Q�D�@�'Q��6��O����O��S6J�P}�_���IZ?��Ƽ��dQG�̇aVb�s�IK̦���Pyb��8�yʟ��$�O�$�<��Q �/ƈ����`�`�xl����� ��d�<A���D�Ok�R�v�<���;XY2�{0���Q��0 ��ß��	����	y��'U��3�AJ�X�l��K�B�@��&ªs�����O���?1���?Ye�#q!\d��D��dV�C�)|��\Γ�?A��?����?�/O�� d
��|re�!^�����W���$��Ϧ}�'eRT�x�	����I�oe��ICeP]Y��>��(!A������՟X�	�����{yBJ�<7�N�'�~��0:+�cЬ�<IZ]; eN��M������O���O�y�T1O��'�kԲ��b"3���Ǎ�M{��?I,O�����c��'���O�A��nL�D"$�c�H�Mr������>���?����Y�<!����D�?U�5�ڸ]fY���J*1z� y��8CJ�hg�i��'\��O*�Ӻ�Ԧ�= `���"��@�2���EAǦ��I�����~���ϟ0�	a�'j���ǧ��"XDb�@T&ߠel�!��T	ڴ�?Q���?���VB��hy⃆�o#b����;�Dq(kU�&6m��4�$��Οĉ� zAH�l�|$�s�I�  |aſi��'|�·/T�����O���6[ �SCnO��j�{��͐H�6m�O����ORTC�0O��蟤�IƟh���G�o�;�i �W���'� ��M�� 	�ÚxB�'e�|Zcnr�3�IĊ�
E�cs�M��O�`N�<))O��D�O���<��%cX�����&
A��c�D��0��!��O^�O��$�O�]��)ثv�:�)D��2zʦ������<���?IO~��KQ���)��d&bE��B�옊*�g��'��|��'�"b\�y�, 3|���T!N�{�2m���݆up8��?����?�+O:��`o�f�8C�U��i���D'B�qE�D8�4�?I>����?��!��<�I�,��2PMl�[3�޶FAhy�Cm�0�D�ODʓ^u�����'U���]�M( Ă$T����=?�O���O��@�*�OP�O|�SA=��X$%�|���ը)�6��<�jɬa����~��������u�!.�	XF��#lr`4���t���D�O|�	Gi�Op�O*�>� K�,r���R�\�!�N����~��eZ٦-�	�8���?�0K<Y�[Z|h n,l'��W�l��xsv�i�nM9�'��'���S�?E�!W#ƒ��dFv+��o�������HyCNE���?���~2��c��[Q�NG ݺ����'����y��'���'��%��+A�ya@��
��|ZΉ���z�p�$�/Y�,�>A�����a,񰴑p�>V�ڜ(A��q}RbE�/��V��������[y�-¯ r�:����I߼���ÞR���O7�D�O�d=�d�O��:�	�h�rt"�1D�P`��a2OJ��?����?!-OȠ�Ta�|���"F���ڐ =���\}b�'�"�|r�'�R���y"M�5F�y��O���P�����9����?���?�-O8<���J⓼d^�Iud�>=#�Ya$`���Q�M3����?9��bHۍ{R�I2}����ԢT5@�ҥ�׏E��MK���?�.O���$D~�S˟��S6}>R�
��\6|X��g5vW�K<����?qQj�<1J>q�O*8A���<W޹"E��	k��`�ش��I0a��Uo������O��)�u~B�עp�f�YQ�v|%�֏G��MS���?!��9�?�M>�/�p��t��9[�m��4>����K�I�p7�[(H
( o���	�����'��Y+U�W�
��WW9����iv�V� 6O�OH�?��Ɇ^fE3�_q�}yi�`t�$xڴ�?����?�g�pL�����>9�e��B��`��* xq�M���?�����'/��'*<�`�E�qh�qA����brӺ�$G�:5��&��^�'�� F'�z<!�F�5�h9L<������O����<��C���'�Y�$�~��Z�KP5q3n�:�?A���?Y���?�O>Q��~B�F�b�;�@�/�|Z� �M���s~2�'��'��ɝQo��O=��V��(��y���Ҳ
��pcO<����䓑?�{��P�b���;�!!�������O����O�ʓy�x��W���!�),��#��]9#t���+E�,7��O^�O���O݁1�$WIp�v�)K�ԠRH�E_���'�rY���⩋��'�?��'_I�	��U?Y��#�)��rz�ɠ�xR�'����O4��"ऍ��)Y�z7����Æ�]Ubd�I��0���D%?㞄Y'�*C�� ��[vX��9D��sц�Z�WQ�,����U�D�Q��TpV%hb_� <�x���cC"Š&�W�8��������I�4`�Ƃ֒ld�H2�)]'=񸱂��-hP��h��?e��%rS,�Ќ"F�݄@< (�g,X-)����#tc�����i�VD������3�ٰZS(�Ie�
 ���rA�=���'��'��֝��x�ɍiX�Q����=��,i�y\I��ǋ*
�����9b���;���?� ���֌b7���<3th�"$��(`��Y)6��:�uB@e�2R?4�ٟ�hDy"���Z܀��]�	�)�	��~���?���hOP˓:� g�#W�D=A�F�
[����#[^t@A;GE����o�:���E�)�,O2��U�����!��U#�J�Ȁ�8X�L���Mݟ0��ڟ���1^ܐ�	��,�'p򤸚�ǉA?�}qC��Xj���+��f�d)r˘ �L(�ϓN���P��\3���݈��"��j�"5��\��X`�M�rx�:5o�O���84px��(<5^���n����=ъ��M�O�|������d,r&I�]�!�đ�o�t{RL��TOZ��@�w���H}B[�蓁H%���O2�'F�\5i�ٹ!���	� ?g>�-`�K�?����?��ԟr3l����+�|$x����i�t�~�꣬�1O�	�P��}�Q�x�dHCŠ	�"�&>�&>��!NJ���R  ˷y8�`��>ʓU;���(����_�O����X�O�����<���;<���F%g�z�І	�t��	$�����~��a[����SR�����<u��X��П��O$6����?1�a�hm�"�a��|� M�8�ȓvo۫JG� k���9������I8��O� $:��ӻH\H�u�W�0;Z��p�@6�ڂ&=N��i e�#�֔���,<q�w�Q:G�1�J	�_J1����f��s��'�Җ�����OL���$eB̸���©D��)��"OX4Rg^7-/���r���`�Hu�����HO�ӷZ?��Ca`� \�DۥC�k^(8�����k�%�S�0������I��L�Yw�r�'s2�q�J<=�ȑ�nC���5
�'<9xT��,C}2��׊=O����nK�`yxc�ĽDn����O¹
3.N #I"��be}X��8&�8� �����(0��Oȥu�'=�Yy�'�Qq8Q	�h�kׂ��y2������@v6��gZbr���@.�S��V�����:X���(]�]P�(F�'?&9��$ѓzA2�'���'�d���'��'>���V�'L��^+X[��jr)�*&,��0U.L��p>�e%� ��Y�䬚02���+�����-�<E�2��$�P���'���bB4_ ]#7�Q;MF��pp��B�D�<����?�I>�O��h��O/�&`!��Dʆ�
�'К��T�8[��C�O�C��q)�'�7�W����'��M�5i�x�D�O�˧ ��!0���V*x �w�ϕ`z������?��?���Ǖnx���|]>sGS�$��hqU���P�:y�v%�B��ZDF[�>"|jc�СQ���t�1�D�G�' �p���P��Lp����|�r�Q';r���(�6m��L��̚��?A���9O��*"�P)F�6����l��!��.-|O� oZ��M[��,�`}��`�-y��=����:�luϓO2*\B7�݃�?�����iݖ����Or�$���G�	7a  {a�h�m�"�Bn�F�&��'���?���\b<��,�:�Y!7�Q+�9�e�*f�ɧ��R�B� b��X�Ov\���+a* 
r�'���'��OL���IG(@Ud�WYd}�4 c9Oh��%�O $�T	��b�R�qaZ2)iٲ��ɞ�HO���V������h����I�Sot���Q	�(R�)����%JQ��B!��+�t�ѡ"�<[��[e��z"�ц�X&�
�*��͑S�ْ+���r�@��fй<x��) 6Z���ȓ��%H���63�}y�X�Z�<�ȓ�a��i��^��Р�) : y��[��H�T6꩙f�Ġ_bd�ȓ~>��7�� �@�9��	�����
�L�R�ȋP!��95/��8H��r��Zc�ߐ4��t�G�.�j�ȓfn�@��!Y�(���t�X��ȓj׼@!�Kߘ"�r�i�`YLF`��,��� �N� q6��P1H�f�����2C֍��+G�g�n�pӄJ����C�F5+A��b�!�҈һJ��ч�9Y�=��$		%�5�ׅF�<Δ�ȓªX��&0�����^5[��ȓ~�b�R�g�/uz��C�A��4��B,��;�O�l x����S�:�lh���8P���R���� ��'�`H�ȓ;�d	3c���;~�DYE�]�XX�نȓ|D��]�W��`q�oj��m�ȓ����\�
���SS���u��4�ȓ�M�� �uvv����x�'/0D������)r�h4�1j�0?�� 0!g*D��� �8 ]��%��RaR�J��&D����L�-]G���e�O��M2g!$D�(�늦y� �����)p�ps��!D�����
[~>�āݎ���5`4D����O���h �Z>pVr3a�0D��:š&LV"�Y`��\�.��@�:D�D�D/C�%�� ��W�� 8D���D�0$|�
Ԧ�5U�$AX �(D����c�*�L���<Hg��!D��%O�XH���q�84+��1�"D��)ЂΑB�|�����\$�a%%?D�� ~dZ�F�0N�&��j߇I@܋"OHH�%��֌��b�S�|a$"O��Q���>rhy��ǐu��˃"O.�$U�6P�:׏�/,$
`"O��
2�G�#b���V!9+�^x2"O����*Lp����%t��}
`"O��P��81��Ǎ@�L �"O̝RD�!���d��<h�8�6"ORh��$�%;L�ꎕCn�ͻ�"O0��74sF�8��CXiv�y"OP�Qt��>�F�+�
��\ �h�"O�zuIH-����^�r�l��"O�L�f� �:�n�s�?�	�"OD����EN�6�pg܂<�q{'"O���Q�,��@��ݷ�r!��"OR�0��
Q���ے�܋w�d92"O��y��\/w�,�0�Z)G!�9�e"O$�0!�� �M�FH%N$�sF"O�B��ÝW��b3m�O�*ԋ��		|AB�,��2~�Z�������59W4B�	�OE8I�"F�U|�(D`\�{�˓�Fѡ"@���S�O"�=;wLE�j��P�fR3["
x��'�0�أ,�%RS����,]�FP*M>��.Y�VpjÓ?2�M��Đ�Mp i��fI�U8E��I�;:�m�t�D�_�"���)�~�"{��W�H�^D���)[��.�y��8揟'�B�E�Ź$��}:���؆5����� ��
�K!�$F�&*�Q1�,�=	�*�	�	�7�ɱ,�4���'�e�)�'SI�<��*E����fJ�n�l��ȓ=f"a��7'���&Q�^�ܸ�<��P�Z�̘��	�~o���!�֓���V��}��B�I' �i���T:9m��c#�]x	�B�IN��q�i &?�L�X�ZG!��$�����D�.$<b�O�!�$��#��lQ������3w!�d�ji��+��,�X�`�o�,Q!�dۜ�z�A����E���^&HI!�ē ��\�e�0X5z9`'/Db�!��yĆ���iڵ- ���4~!�DH>�q[���G�J�1RMط%f!�DM�[$Z�)���>�>ј��&eB!���|HDr�&V#,�h��E�Q�!��L\���p)�)h���g�4�!�:N<�qH�Zoh0�3�Gr!�+I�bdXr�X�n�F!��@.�!�dۚf{�4�P�D�.�j����!�Dן5m<U�@"�L�feX#KS&*�!�D�@�p�Q/�2c|�h�B	�rz!�Ѫg
���B�3uy���G�:(w!����r�F�zs.�w��7F׭	`!��cJ�!���*+�� E�3]!���@��%�I-��t���T�d&!�dH	p\�2�@�*!��1���t!���']��J��N�4�cƒ�Y9!�d�C���".���aTFI�H!�ݼ&�>��&��=S�B�;Pl���!�$�%�*�#�>~^Dˡ��F�!��Ɉ)rdQ3�Y2l�����Y�e�!��&Jв��Ή\j��&��&7�!�d
88遀��0¤@��U��!�d�2�������3QH��"�n)n�!�Ė#D�!ʵ)?��r̓8`h!�Dt�zy:��ˌY3H`81L�vt!�$A �n`���Q�` vJʴNG!�� ��B��7nD��� 	{����"O����J�d�����N$��5"O�lIS�Z�i��'�[�Z�,�"O��rv��+-|Q&'9D���"O"��E��\&\�FEռ@A�`�F"O
�X��)=$f��U�%E:-�"O6i[��-#yh�Z� ��nԠ]��"O����	�YO�)�d/@)��SA"OP9���62��;s��
`�ִ�R"O��b͗1`��8kQ�%�@�'���т]|��
"�Ly�W��m�F����Y}����<���&�����O�u���U<2���)v�F'v�X�t�d	T�����ة��'V ܻ�%,�>	�% �N20z��aH����������c�Ȑ:�ʘ+T'v��f�Ƀ5X��p���G����O�yed9Pq��ԮR[�4�*Dqb���|���aݸ0:��@c"O�d0�*�Bm���d/f�r#�'�:���"�4�^MB�j��~҉�W����b"���f�N|���(�yaH�� !��	ܦ`G)R}�>p�H�o�,�uG 6��S�8��\��)L�/����|�b)M��~冀N��<Z3�]�8��`����0?�a�Uh�u�듃.��v!V�k�f�aA�":3.J�1��A|v|p��$ �#�uI-/Z��sXY�\4D|��1Lp������H��8��UE@k�n<�pFE�6`:�&Q�U���v�'[�}1I�Y�y��߆f��k�'䁛�Q�7*�ljbDA���S�&�Dٙ�'Ͷ��f@��9U� �1Ȗc��q��cd��a� F�+q�%Fⴵ�ட�Z��[.h��˓� ������@���y�g�1�l{f��i��� T�J �p>A�@�j���L܂S�d�QĄ�
��i���,ry:O�Y׮��,:AA�9̈q�L|Γ_�̱�$�!�fX� N˦Z�R$FxR�M���!�gAY>u´̲"	���?�'E1`8�f�c�9Q�턅�,d�/�� 2�3YNYڤ�2Od4S�
��st�&���tA�BVe.pX8C� �,B\��F�{�J?�O\��kI�%�ҭ:SO�7��O� :!�dYI��O�;����F�_f����,�O��1�A@�-l���֟���sRZ�L8���2�.P���ç�߳LGaybX ���G�#����*���"����E�� �]SZp� B��RXx5nL�w@�	7K����1�m�O��J�B�5��� D[�0 �"�$XA��dHZ�aF�����BӒ��'V��Θ�)���ǌ�_T0�C�����Y9��7�z��a��3O�k��&(k���̋�H[9� A_�_�M�6��U@�Y�4�x�i����x'?��R�v�1x��#;�1���1IjaZc���� ��`*\zr
L&MіeS����#���hR2�"(8?1���+t$eM@�)��1z�h���496�B�'������a8�����ȠJ�i��O�B�X��ŦN�Tth1�G�#\*��V`��M�F_���dY#2��sbR:�:���!Nϖ4�O��q�&Y�\x	��-Ռ5 b"�>��K�Y�jA:�L��v��iCE��F,�r�j���b�W,ڪJ+�� �ʈ��6��V&N�����-@.��J�7
Vtx�!�x��-�rOz.�s��r�M����$����O����h[$c0lX�N�d�<�D�S�d�&C���c�,Q�@�����D��dZ�x/��굨MH�ܭc�K�>y3�^�a%�`�djx��Z��U�0��b04��`�&z�x�p�)U�D��$e��Ӻ����;)z$  G� i˼��RM�$4�}�mH�-)Le���'T}I��֕Y����,����S*Tw.��2,ݶT&����{���)Oٮ�YnۄY��3C΋b��	�-�f4q$�o���0��B�/����iGQ}B`��3^2�ZA��rD�`�I܋�b�Bnțu��8(#H�(&ļ*�!F.hd�x��^0�(A�o�c�2x)�K�\����0`r��s�)�����_0D��X`ːt�S8h_�P�aU�ƬB�K{������'@�l�z䪰 Ih�Z@�[�u[�T�TY &ye���d�� ��)Hl2Jaʇ�H�����C�Q�b��@9p"��R!^��0ǒ�#��x�ЩH�J�z�G�>Ҟ�p��H�4*�-;�L�)`��?h�8I��!�/H_�H��Q:U�-@�ĸB�h��H<)/�H˦�)W�&}�&��"�d�'�R���&O*A�L�W�z�L0�S�R���~�l��s��y�=xІU�<Q���Qfb �q�_���[;E��S�.�\��xt	��%`0��)��R��H�T��j@��E3Qb
}�<���D. X��@�R������P����I�10�*q�m-<�'� �<1ǌ8�.9��+����t'�t���3�͆1��aB.&�L����c���!�ڋ#�l�`6��1j�j�3��'T@J��N7P�;2�M4f�*���DM�BT��8� �_n�Zsl��(L�O���w'S�8�΃VTp �
��� ��;c�B�M��rT��ԉ����s&.5؀b���Q��A��
ٰ�E���BZ��EO%_Fl�g���z�Մ�=z=������Y����Xe��\�U@��v�4B���|����ȓ)�� �Q�C*2�q'�6W�r4��VBHql�®�2��3tHJ���*~8�s�E��~���QҬ]F��i���[w��
�Q
��ݱe���ȓ*x�Lk��}�a�M� 1���ȓ^k�� �G�A�X���D4hȰt�ȓ��y�������X��۷
\d���$���ѕ\q�,u�v�^r�� �ȓTn�8�`��P�n05��m0�=�ȓp�j�1�腴��t�OZ<+�tH�ȓ�@��% �*E�:I�c�� ].��ȓX*,PG�V�2p�S�298@��p�����	ހ6������@��ͅ��`��dA�1(<`8�II)gfI��&�����AN��J	�p�B��ȓ*#F��tOÊW>0�3c��#(# Ɇȓd�H�t���:��n��j% 9��g���D��2���ϛ�R���p�Vmӑ���Q���P�jd�ȓ+��	r�ܺ�@�cኺ;pb���i��L@R&�����"ߤ���kTىgN�G�<��#K�6"�ȅ�n
@JQ׌A��Q;р�(	�d�ȓw�up5�G�:�Qۡ��lXb=��Eb�չ!�ƴwE��ʓk��} l�ȓ8�쥙��#	����.vذ�����9�-=T��bG 	LLh��ȓŎ�I'��5�"!H�"ЇU��чȓ"�e	�]��}9���h��	����Hd2!�(��o��>T$�ȓq��%�̖#������z+d�ȓck0�Sen�;j�Rү�9����ȓ[6(p;��-�D�� 4g�谄ȓT�����c�� � ���X0��p��{rn�@ ԭS����'U�!zхȓ|�̙r�V)|n|�Dj�)k����ȓ ��y�7L�H.�9B�g�A@�Y�ȓVHJ�z���˜�+�)A$ډ�ȓ�a���_���1��<C
�ȓJIJmZ�L

o@2�:P�-�ȓ&���b�:3��(S��h�:P�ȓ@��|��
��Ik2�c۞rb��ȓ}�Y8���8@,F	����w#R��ȓd��c��/OhHY�cO=5ΰ�ȓCO����*0��286 �ȓ4�a؅`B���pjC�[k$��ȓ5� ��,�&L�4ҶY�6#�Q�ȓ>L�T!���9Vr!�βxl��	�Dr�"��	��("�fY�S��	���J�h��\,7n��X�J6�RC��8�0!q�� ���Hم`U�D�C�	sI��{"a��-"P��d�7y�C���I@��~�l�X��Ӷ	dJB�ɋUn����dK`5t5(f��48B�	�=C� �q��7m`h���%>�B�	5P��YxG�R�^L���P)En�B��>�*�m]&�N�x�`ϴt%TB�	
 ƌ h���,%>��F�˥chB�	�'�L2a/%��4��I�I�&C�ɠ,���Q�	
������B�)� �p��޹T�R��2HO0n܄d�%"O�����;�*iȈ	�h�j�"O6咑F�
�c��+i��4B"O�lY��A�C>��@͍c����"O�4[P X/9��bg/��QV��"O X��"P) )Ҭ{#0�x�P'"OX��um�A�W,��H��ݳQ"O�9���>��F�-���"O�Y�f��8e�m��#c�6x;�"Ont����0�H�2��+Zz\�"OL}{b�G�t��"QGG��"O:���+���H;wa�Z8*�j���r����^�"uV-���7 D��%�I�!�ă^P���p����0`�1|!�X�~Xl�K��W N��r��S_!򤃠P�����&\=��`[�r!�)�^�H�M1)v�Ɇ`�:M�!���S;Xt���,&97F��6�!���o���XT����z���04�!��B.r���J8V�zŚ6AV!�d1
�,I&mU�8�ys���H�!�C�#F@��c �":�6�3b)J4v�!򤞋�Nd!�����`�
V�1�!�щI8�aHa��:��dz�*M�!�䖆Tۆ���̐+~� z���'J!򤑬ܬY�O�p4�2�H��J'!�ыu�BIP�ų1���&�F#!���z���)�p�\(p!��g|j��F�.��B�G!��?x)����:>����%X��!���t��2K����r�#Q]}!�R�X(��&�B�9�� �T�	�(A!��\�A�Qq7͚�W�~ ��n�-E=!�$W=d��e;o��S��e��mܘI>!�$э>I6%�$MtFA���G !���	zH\�*֔|�Y2�
G�2!�DQ�Yu��"�`�� i
pP��C!�D�<"f� �q!T�Y�A9���mE!�z@�;��H?k�� �5��A!�C+o|X��TEϯ���R�Mټ(�!��]	 ���kg'O:��TP ��(�!�$�]@��GG҉H̖-���>^�!�dV h �`&�X��`�pѢE9Q�!�Xw�MH� щ+�N�aW!A��!�$ߎ@
$%���]�y�V`c���<s!�dgS@��K�1l�1��iИm)�B�I'K�aiF��3��}cS$ӥ:�fC�	�y3d�S���Fz�i:�QnAC�I�6`1#4Ǘ�x);2aʥ1 C�I�+����� ?[���i�Ǌ0x�B�	�[)��R�G�@}�G��Qu�B�	�-�9x�gD�;�D��+�W~vC�8r�V�i='l-���4N:�<��a[0�C
x���d�T�C�̜�ȓ!�aca�C5�̴�T�\�2�܄�x���j��J$%04�ޏ�谄ȓE�h&���E�`��6'�B�ȓ`����\�|�*�"����Y��8��y��ԧ�b�h�j. ���}߮D���*.N�����7�@��ȓR��U��� ��q�`�Z*g�%��AE���G��u-8dY����x6p͇�Q���OG0?,6��P�8H���ȓb"���%�2��+ܽ�.���S�? �5�����[k@	Y�N�-��X��"O�1Q�o�#e��$ÍU9.��\�3"O��;B�ĀPQ�Pv���v�~,�"O�h�c�8g� ;��T.��i�"O��)�\9z+�G�3]���b�"O��A"d\�O���	�fŐ.�̨��"O6�v,�a�����,7�^@2"O*( fmU�8��
�jT��R݁w"O��FE�Hcn�����L�<H�3"O����F'~���"e	DN���z�"O<p�A�Q�b�`�7�@�ސ(�"O�)8��L'8���6�¹�`��>���Ҷ�G���	���.,Td�� �4A���Ċ#PD�ER
� ��I� Mfx�4
�:i��8��?R��<���T>� %KIC,;4�_
o:���$D��y�ȃ�lȨc�Ɍo'����!D�X�3A�,�c�Bc7�)`�L%D�ء��W�xLl��QN��N�)b`5D�샖kJZ_4��F�g&zdrƆ2D�����-hU�5��E�0���"D�"]�`y���/�y��m6��hO�ӨxA�Yr��-<V8�ȧ�A��B�
7��(�a	=BJ J�ƛXi�B�ɫ<�������~?�U�&KŮN�B�9Qu��at��4�ؙY��<7��C��<`�1Y&��X�ڨ���&�XC�		("�#7�Q�]�� � ��/�BC�	�6_4��0-�6UV%8saWX�LB�I�S�����E��QHԻIBB��b^F���'��y����?,'$B䉎r��"g�գiD��)EГ/L�C�I5l�xRe�i�P�����s�C�	�y����ӋJ�E�8��Bƒ�[mdB�I&� �0�)65�����P&ku�C�	�jY��W�[n��Q�L%<�8C�	�G�4���B�u���@��ֿ5QC�	|f4$���Q�D��wo�B�	!s�\��s��P�kBbֹ|MnB��� !�#�a���#'VS#�B�	�$bT웁�¦uV���'�FB䉛c���h��:^��a��X^B�	�s��*�I�rW�qP.�%S@(B䉬s��{��̻n�^����$�dC��!����VV�%sfQ�`,�*G�2C��B��d�ʲ|�,�'�7>R#=��T?�狞�9Y,4�$��fe5D�<[C��;��Թ��7&�� �ҧ0D��k�O��H��o
0(�P����<D��ca
�0v�4c�ϒ�
Xpk8D����O�!�^����O&^3���5D�tC�� �Hլ����&M��jqi2D�x�@O,C�*bJ�xր�A�C�I�t�^���)K�G�x�a�Á/B�	�R�#o�;rL��ת��G�R��ĵ<��G�1a�qB��ÿa����D�F�<) �:�6�K�gH�\9Υ+��H@�<�2U���sQ`J���@R�<��.Y# @A���z�i"�Ph�<9Ab5Μ� �G
?M@��w�P�<Q�m�'�raj��u?�t��e�<���T�B�B��&D�iq��I]�<aǠ�k����B�e���d�@�<I7�S"=�0�!Ì�:��@B�A�<� �@���>������dC��`U"O8 �D�G��nu�����=6.(q�"OjASFC��Y�0��F!�F��5��"OnTb�M�
I���{ �	0�N��"O$M�g�T>bzmK3�Ñb�� ��"O��9�ašPͨt��fu��P"OHD[6N�>�%i@��;
\r�
�"O�y+%"H!$�x(%A�z{0)Q�"O��h���\�.�hQ*�A�B���"OB��L�*�ڵYgU8l�Qٳ"O������2 |�b�F�%R��٠"OB��WI_�I�I��̩>����"Ob�ۢʑ8mB��M$?�B�i�"O�D� &�B1�"�mK|Q�"O��	G"_~�� go^
R��pV"O�xq���Z(�p�̌=� �c�"O��S����M��lR�I�#�����"OP��Ɉ n��%k%h�
��� �"O8ш��Q�p�^|1�Gݚ~z �y�"O�)r+�cjlX��G9v�8��"O��ٔ��j	C�fH�#p܍�'"O$�":_���E��F��|��"O�H"s�G����OĆZ�f��1"O~��h�1Mh�b�Մ�Jd�G"O� �T�¦)�&�.d$�:p(��!��7`Tc�\T�5!�F_�9�!�J�X���C�m��&�,����5R�!�������ϛ�y�2�1 �BQ!�ںZ6$101
�m� 3�K�r�!���D(��K�]4f�B�1.��!���-�6<&��J�V	���R�?l!�D�� H #U�O������eZ!�$Mf�F�[f�ɧ/�Fl�� -eA!�dř<c�,x��H�]��IUo4~�!�$؄
��uR$�?R�l���GUd!�$�ps�h���ܛ�r4+�L�kS!��0�t�h	d^y�!��,#!�D� ,�  �"�+%bT1��83!�D]�b�l]��hQ�� ��$a�!�B�RUAK������n��ITb�H�'�y���R��,����Cn��:�'[���Sḷt��%z�<a��"aK��^5�h�SJ�s�<iqaB&ֈ�u�;J`��� �d�<�u�T�^dQ�M�:-%�uӃGc�<�M1(E���%��ta	e�b�<a4κ���
�Y�O�b�<���ˈq�Z�����z�Jህ�c�<Qv��V�����T��IPӠ�G�<)"�yC�����^�0�H��N�<��ڃk��mxRg�d8DB�p�<a"�Ųi�Bt�1nԏ^ʂ�����c�<�%L�_���k��KA!�w�<� �F�F�mS��W:X��Bp�<G.ʮ6T��g¨fW�ґ-Fh�<Q&��?s9��j��Z"0�q�?T�x(2�:b�&��--?��c��?D�T���Z�.�r��]��H
�C+D�\Z��ĿMl��1'ѵ+|�)�#D�|IuĐ�h�^[W��d��'"D�D2���-*�"� #D}gb�;��4D�Ӧ��$oT��V�&�DlSa�.D��ib�6��I@�Œ�7�RI�ǈ*D�hG-[d�hQ�&�Q3-~���N#D�� N�b!��=T���Z�%Uu�F� �"O*p;À�4'ܐ쉆�L%b�,��"O�X��G]61��[�/y	��"O��#Vj�g�}�tn��J���
�'�"�;U�,�>Pk�R�"�'�V$r7l\�W:��p2��J����'����� �r���KR�I�=f���'�����8 �$%��g��	�'���H��$v�D�C'b��D1�'�HԒ�^&r���.�e��c
�'�������;rI���\u]�ɩ�'�r!Ru�\"@&�,	��Ա�f�<a��ۯ$�4�
u�ѽ9xz=�6�Bz�<	E �/װ]H�Ը�n�+���{�<��I̲nji�1B��[%ǖx�<a2	R�(3��C�J41ve[�@V@�<�у�Y��J�/	�Lc0�a�<�D�;��� ��'D}�UT+�D�<	� \�v�� �6�RQ�qi�t�<�T��Nnh�#���f�v P���p�<���11�}xG	�Zӎ@Q&�G�<	W�D�Y
�Rp*M���i�<QC$A&1JP,bB@�icb9�!c�z�<��kK "�H�C#�I	'VT"a�x�<�+���"���܍0-H�%��M�<�4��<=�Ƶ B�e�|P���Q�<q��#��dhV�>$����[P�<9�jU�ǀd ƩW�y�踰dHI�<	Я�2�ƀ���4{��@RL	M�<@�>-Ѭ�0	&q��T�pJGL�<	 �ҍ{:�}��̐#& ��RS�D�<	%��`E�y�'O�8\A�S-�w�<A'�[9Q��1gɟi��x�e��X�<�3�ݠC�$��W]�~*ĤBe�V�<a��j,�8����=+H��VLI�<�ƚ#Q�]ydO�>;o c0��F�<��*��MQ�����i���F��\�<)��8n�^q	�����ɐ�[�<y�d��]ú| s�5�	�d`FU�<Q��.N�QíP�n\`��[w�<Y�dh����[M��+T��p�<��̊�Iw��(2cԋv�a�#cT�<��bׂ;�J=IS��� 7�Ԣ)j!�?��X��#�1l����ч�%=;!���2�0��@��U�� {�&�>!�d�E��E8P��A�Rp��T/!�_N�489���7[wHLK��Z�!�$�7 �]�֫cZ"�˔��M�!�D��0(��ቜXv搻B瘸*k!���$R𘱦+�c_�����L!�Ć���R�`��J�>E�֤I4�!�$��p"<�f�� ,Dl�QrCυuq!���D�y�g*Ӱ2���VI1a!���	U���C�mE�O��Y�`C]%!�D@�$0��S�I�ܜ��^�F!��F���s&���p̂w,E/!�d��	S�P�uǕ�N�v`ʔE�6A!���;�@˲�� ���iQ��!��P�Yh«5k��9�e/Ǣ�!��/{���a̵�R�Kc��!��)9��@��-��r�J5��N	!�C�ASx���{��ኧ
�T!��<p62�Cdʣ4����QC�&cC!�����I�L%��j�a@>o*!�� ��4N�:`����U�<����"O�\{Ġ%���R�Ǒ�S��#�"O*-��N�-Sz*憊%w�� "O�5�"���Lvjy��h�4|d�i��"O&�����٬�y����0e�$�C"O�UpcY5Y�4ٚ��:u��9�"O�Q3�F�hL��S����=k�"OZ%�R ��w��g��i$t�F"OdM����=1Z��kA4Pz�4�"O�9KP�X�b.H=e�H$Td���"O�iء�߷�\� E�ӫoL�9��"O��J��ׄi��� $�6/�i�T"Om�����0��\hr�K�V�� b"ON8��,B�a��dh��\�Q"O~`B��#~\͘�G�=�ҡ� "O�\�FI@� �D�[�X@@�"OE�R@ �c�c�7����"O����i��W�Z	���Y�r��G"O>�7�E�/4N�2�=x�Z��s"O�U	A�X�6�z��� �}a9c"O�4��^�\����̬I4(�"O �z#Hү{�<m�b�L<Ұj7D���Ќ�j��$J4�T�pP��2D��ٔ��)
 yGяԜe�U�:D��
%��4��(���2�<��c�+D�3�J��-Ba�9��%Y��-D�ؙ'�L*'�H%斓9���N*D�T&L�7CQ�����V^�p��)D� �>�,x !�� U��:g.'D�Tc�+'[������H���1D�t��,�v�s�6S֙�Wd"D����
����&^$At�� wf!D��� ��!xh�2bN1U�l��f.5D��"Se�:/��I1���b�k��4D�bc�f�z\KqI�`VM
0D�8�u�c�, 	d�W�{� ��1�-��<�O��KS<��ň��K4oq`HX"O��JEh]0"	ș� �+>p�`0�"O:h�/�S~�١��� p�a�b"O@�3s��#j�F	���G*;��"OV��q��$�HQR�O�\6�9�"O��S%Ɣs�Z�a9�^���"O���7�E)	Ml��G��%J���"O�4�
+N�B89�Ä�sq6!�W"O�@afT>�>5Cc�Vfp2"O�	r������5$�薤%ar!��V����h��\xqq1n�e!�Q� .�g�7k��XІJ#U!��C�/����G�ep�EpV&��L!��X�Q�X��)bm|0Z�$/{��O>�=��P��G��*#����k۔Ө-�"O�bG=o�2d����ϴ�"O�A㤚�1Ѝ��gҖ�T"O4�hte�7e��6Aѳ�@�@�"O��B�tRbDˑ��>ZA4l��"O��8� �]�	R3ԜR"�$�q"O|����p&E�rN/�HbB"O0 ɔbX�_�W�%F�$4��"Oh( �9ռ�JS 4�9��"O�$��O�'X�Ī�N�!���	s"O�d�EY�H�����R�S�L�xS"O�| � �>x|}��k�?+�"�0�"O�8q��),�P$r ���9�"O���S*ؖ-���p�`�:ie�Mˆ"O� Z1�d��O.LD 2 Y/eB��"O�!�C�˯.(���@/m�hDAp"O�M2q����M�7��-�y��"OU��M��:�0`�s%�^���"O��f OF�)�j�[�
q"OZ��GL&B�F*�(�pa#�'��Ă�6�N���"N��zA��j�m�!��p�����ϡ+�P�u�ı�!�$2��P K�Sx���ÿ*�!�D؆-�*<�D�X�s�N��!��-�$B'ׄ>�*���/��q�!�$���I��(֧?��Y�aO_'Z.!�䑊U|�����%e����" C!��	xP��F�LGes�J1PG!��,Fe��S�
i������!�$<�А�DdRs��U�+@d�!�� ��m����O�EؠKJ�Q4!���0�Ubf��=	��3�Ō4!�d�'B���+���ę���X�W)!��� �xYS�dQ(������<(!�d�9b8�7�ɿi�\�:7ʂE:!� 	`x��)W
ޞA���,!򤘛L��	��+C5=����͝�	+!�
���$
rN^)L��QY���D
!�dS&&�X�c "KJ\(1�g��[
!��[�E@��?_�,�v(�,!��BiXRU��"������@�/ !�$�1����A@N{L܃wM��%�!��� N���4�Zxph�l�2!��?A	�l���r19�,�!򤖻J�X���g%��Ê¶
!�D}�.�H�Dͽ2��*6�^�b!��.�B;q���<� 窎�N!�d� �Nh2p��tĳvʔ�dd!�ҕ;�����@).�,P���ѕE�!�Dg2 �P�}��7�)C�!���9Y�1"Ħ�a)�;�Zt�!�D��_��Y���+|�����!�����y���]3Q�P+aE[�!��*}M^i"�gR�x`�Y�'�!�ϡF�Es �@	� ��Ϲx!�ě)8Z��g	�P�DUZ�:08�'��D��~b��J�����`q��G$�y��#��Mq!��]�:e`@hH2�yBbR�|*8��u+�&~��D+�bS��y��2,��|zG��)�La `���y�/Njj8�$��'�����iج�y�ꒈ+��x��'�&�f�yr��/A���i��T#6&��F�����!��|
�y�Ò�~��\8��M�lTr#�]��y�k�
Tnu3teH�����G��y�i�%;�h|�%#�BW,��y2Ǌq���+�
Ě z��c�K��y���)$`"��ΜM.>��E]��y���y|��QQ%�!=�R$�G����>�O��Z�mF�C�}{��6k{F���'I�X�����w8��쌝0��L��l$D���'�����"��5U:���P&$D�h�Ă�0+%���e�n���R�� D�h��Hñ`*L"�(LA���:!�#D���A��4�"I�Ӄ֕=��i�CH<D�$�*�"�������0i�1ʐ�8D�L�U��_@�)s���>V�u��5|O�c�������o�"sR��9�(1�3D�� �h*b�ڦv����U*,{�T��"Oti@��SJ�Y��J� UjL;�*Ol��5��Zhz�s���x�'pF�I���8t�eRc��1$%�q��'�F�CW�ϣN���	C�޿ �`�@���'H����M�u��` �i�	Pڡ����$ ;D�)^��mXä%��/�!򄍬n�-k��q'6l�#G�u�!�D��;R����G�k"p"I�l��I䟴��U�Iy�O�,�I��Yx���0eƳ>�����'��`[�(!I�g�P�0іx��'��Ex�Y(y.L	�@�߲��
��?A�yҀ��d�Pa�Y�	Ҕ�K��?�y"���k��U�b����y���yR��k`�����3j�d�sdJL��y"��	=��R���[��	��@J6��3�S�OG�0�`*X�U+�96,T�6[��P�'��d#���5u��IEE��+ڊ�)�'�t9��LT)�#��e4|�
�'e��c�dT�a_Z���aɚO^(`Q)O���䙼{T��Cg��6|�,�h���,
6!�_�|F�Qx���l��M؀�Ey!��*\�|q��¥���8k�	�4��H�)ʧ.���
2��hI��ɱ�^���t���M����A��|����	 �2X�ȓ{Y
�"�B�
u4,с�͇Z;&���)��asOG�JV`�д�	/�����B̓E��Y���� 0�h@���S�Lp��E x�Ð;y*(�3�lčm��Q����<��FZ�0l�+ 2G"��˴��U�<�b��3-�R��ת%9N<P�k�S�<�
2{�<�[�%V$<hǴ��ȓ�����_3c�8y W�[ �n���=��8����v}� �B�!.�>����������$��"uk�.T&P:���8�}�ȓ ��53���=�*�3třk�Tń�	�<�!U��dx(��M;�z��q �q�<�� ��DAX`�OL]La�l�k�<Po��n��`ؘB��i�VAE~�<�JW�,)�i���tLt�P�T�<���p����.".��BIP����F��9j$(\<M��A��p]���	u�'i8�p�fP{2z$nڟyp�Ń
�'�根%#�7A"�t�ւk��X0
�'���qD���)�"@a��Zx�Rd�	�'�����F�m�z� d̕?kS�@r	�'{�lqR&�aD��(�-�8�hp�	���y�N�"*� aC�<�>dR�h���xBa)I.�)�Tŝ�{Nl���燰Y��O8r��۵ ��kT�wk6��P"O*lb�ɃG�Y[Bb��,���x""O�'E�kTH�pNޑy����"On���m;rlP��U�V�%�8�+%"O�]ʁO�u��]�D���H��"O�i���Ψ좥�C �.���(�"O���B��`��3�ݑ\c��Б"O�%z�X��6���ݚ2mR$xD�'�1O��rOݿm_��aoQ�D3$ @�"O�Rvm����yr�rOp=y�"O>��A`4_�x�0�K�*(QR�
#"Ox���ظ]�^1aqj��|5�m��"O����6 ,1ŉ͙J�>���"O�����]�J��T�$�^��"OF|S ǎN�h��g�#'�P$0P"O� (��ń�,�PM	�^�-�����"Oh�R��� P�����!f�:�jf"O�X�c*ƿ�Ƥ��)�B�	�"O�9 %��,, �R �Ic��]��"O����< b�����+[��q��A>��ۦI)0A��"!N�h����"D��@��S,%�0]��)��y4\`2� #D�P��h���AP0o�hӐݚF� D�0��;N؄[�.��%;�� D��rq'ڗ�MQ&	N*C|��l=D��� ,y���
.eɜ���@;D������/����ĝ&nyr��O��O �=��`A��K�'z��J�O�t�����"O�#S�N<�2���c��d�R"OVX 2�
FՊa����<�����"O�m f�w[<���=F�a��"O�x�OG
 ���;$��'VX0�"O]�1	���z�!_�rRHI�0"On�3��14L;vR}+HA"O��%��%V��c���	}@0�T�'���������`V�H�� 9��9D�����e���Q��U�i�v��F<D�0r�� H|̜a�شwb4�#W7D����&�T$�e!$$�K��5D�ࣗm�B,�b �ة:�|�`/D�$����hI˕CY�3��� t�-D��� �/5�p��nˉ���6D�<��,��A����2|~����*D�ıF�=�(0Wㅘ|E��@ӈ)D��yc��?�=K��6k�rh��*O���"A3pN�� �/1���"O��b��c}�����-8k M3�"O�T(S�^�,r�Z4	R��f�#�"O�|T�Gg��r�H�$�i`"Ov���
�㓨���Ib"O
8��I�jM�萀7	
�	w"OL�Y���q|������0�"O*4um�^'��Q�?P��1�"O0lC'���V>,�m��$�dy9T"O�y�N�%8b�ԙDL)٪}x�"Oı��J�kW����?�4��"Of���3R����壕�w�x���"O�X�t�]�n���,�Д�"O���Ԧ�#d�`MyRcU�F�@���"O 8Jլ]����u�G=_�p�@c"O���ʙ%U ��O��M�e�1D��ZC
�-\�te��(8��ׅ%D�d�b�\����� ��YQ4��t�!D�X`�Uw��[Rk�1M\@�&�=�O~�	��xh`�D�x��M*1 �^��C�I# l���@����y�Aߩd��C�/�\ur�dY�nj�5X�I��C�	�N&|���N�2j�x���-ȱ4�tB�ɑX�I��� �	cr���"�XB�	-4���C�Z+V�J�Xǋ��#2,B�?F�0�y��V�*ٰ˙\�B�I%f�tz��Z2��HjP!G2��C䉗;+�h��&��ox��S��	|C�	�j��]��X�a��Z��R�w<C�I�������%gF8�2#/a�B��&����`���S�N�Q~�B�	4F`z�����_-"0���
!h���:�IX��~R��v;�혧B��`P��P��y�jڰ;u��2�Kdx�0�l�y
� ���B��5Q�J q�1v;Ŋ�"O̙�2%Y7z��� FR�6�V�*�"O�x1�gE���poM�
��L��"O@	��s�Yx�Hޜe�0�"O�t�RX�Q�	3��=*� j��'rў"~�����K�xcRmeGZ��Q:�y�L&@�t�S��LC�lJ&i��y��v����I%���c���y�!]��0���B_�ņ�Y�Aи�y�$�QG(� ��}i"�V��y�)_p��y�3A�{�.)��M�y���5c�t[@�zJ2Tpch��y�z4j��0C�t�>}R�,׏�y�	HT;�e#��=��E���y"B��Y�D�PcޅO��,��-��y�FF�s&���]0�ș֪Ȥ�y�)FR%!�cǪ�ceA^	�y��87���e	4b��!J��y�aY�<��Q
1KJ7$
2ՙ��̚�y�"A7.ZX$R�k\�3U�,�s����0����'��HB��<WA��H�HI.�����',R4Id��;1�Rh�7	hd���'��(�Ԍ�/���*��-{"\��'�<mâь����i�|�.xK�'�ހ�p$Ջw��ㆎ�
��pz�'�`�����1��%(s�΢v�䀚	�'m�I�RSN| � �7�x$S��$2�k`�@�C�_���q4)�3W���AD,�H��*6ZiS���V��ȓW����$�Z���]k���{U�5��kL���ܿp���O+w�!D{"�O�T<q���{>j	���@�'v!���M�;y,)��y��T{�' ��B��!��c�B�(le�x�.O�����X��@Gʈ-8�,B�L�!�ęH¬� D$�&�,�'N�%`!�$Q���Ы��n@�[�?2~!�d^I�(����WQ��ɳ��4sf!�D\�s �Չ�NR�|�X+$�+Q!�ښ'Vu@�G��D��Iy����^J�O���$͔Z�ܠ$o�}�V A����>CO�)��<BPjh�b�;"����"Od�"�:py�YYW�]($��"O���l�5e�y���̄e����&"O2�mU�/�`��♲&���yP"Oz%I�� �_�܄�����f��Ȓ"O�t�$�D�, D�(0-�'5������j�@&و �4_^��e3D�j���<@^�@: ��11!�.D��+�GG�p��h�ĕ=b���di1D����ãT��8c��Ba��ۆC0D���.�8����fH�pd~�t�:�����O.��,IɃ�A�w\�e��h�0��q.D��8�g^�I��1A�������-��Fx�$+RE#(�l����[@�h�'fFԟ�&�LE{J?�b�Hmp�L�q&�nf���5D���E�GJ�DA$#9�#��3D����Y�{�Z�Y ��[�f �D1D���e�9{8��hс��"
M�7��O��=�O�1O���ꂅ0���c/�c~���0�'�!�$�<}��(���,M�ш��btBOT0Ӆ��B��Q&9Ip����'�!�$��wwb�b7M�Da�e9�	�'�'Ia|��P�]^n�"&�kXʴR�jʪ�y
� �Q
��� ��@��#%���zD"Oн�efӗA:�D����=�dȃ���2ړ��č�Wd�sb��1�0�[d�/�B䉶z�$�!�F�k,麃�2B�I�[G>PRR(��P� ��eb]�0S.B��<���� {�]�ʙ8b�B��+Ly�(�ȄD�BK�he�C���(i�CKO�8��$ʎ<XB�(`����F��&K�H8U�	�ZB䉼�B07lLw �IyPN�mTB��7��J��]�d��{a�D3�
C�I�~& 	�d�K%b=��� [�Ң?����ɟ/[�u��<`8Cq⇌%�!��M�����̈́�7fr`�W���u�!��.X,�:�Y� ��1��`Q�lk!�d'�x� b�P�z�ָ �aǌpN�R5O
��#�׋J@IyGH�&$sj�"O����(�s�D��M�xo(:AS��D{��	���rbd�?&J�����4�ўP�ᓾlhP�����tct�6�%	grC�	�m�4̑!��:�Ht(��Q��nC�ɩ>�l���A-j���a1o���DC�	[�IK D�V��P��X�pB䉡8H�iB�ϫQ���`���#Q�$B�I�xy"ܚ�n:I��P�gXʓ�?q��D6�I6 ]
�	�É�	�0��b�'^�C�	=�
=�0��!6:�;N�C�C�6K���PE��Ԅ(d!S�"O�m���t���1X�y:��G"O(�ą3p�ڔ�%�̀:�!'"Om!q�h�$Ÿs�S�hj���X��D���7�]"F��Fh@s��O�C�ɣ\H���݁h�N���ĉI��B䉖Tx���m�$ dZ�I�(�p�O@��ē�N��0��,>;U��[2!��A�unlb���X@�J�I�,#!��Gl*��A��Z�Ƚs�.D�l!�D�XسFg������[�1W�O��􄄁9D���̕
k�D����Ψ+-!�d�5_�U���47�-FB�G"O��:�L\�27�5���O�)_�y�|R�'az �;/� �CN<+T(H��I��yB�d�Z�&R��0��$I0,�ȓ2�ꔈ���o�n��F�^h��ȓ(�j��F�H�e���1�h� pR>��ȓ25~�@픬`���V��2]8BI��P�a��,
�L�Ӎ�_`��ȓ�r�K��TZG��Ge&��'~a~b�>]2����_�@������yBOW�$�x�@V�9�\�@�A��yڧ�T~�|a��@;F�r���<D� ����	������@�r�6�Y2�-D�lp��Nn;�0�b�߃^�Z�l'D� �B�փS�\h�D�:2���(�%D�d9`h��	�͈U)�4*Xy$D�,�1'�u�� ���V��A���$D��z4 Æ}(� j$+�'����l D���
-w�X���	Є9Qx\	��2D�!p�O�W(p]�!�a::�[�g�<i�D�R���H�=݀��@��<\`���ȓ5��ؗ�Yu�]�p��y�����J̓l����)F�ĹX�G@>*E�$��\��Y��LٿahƐ��&ɷ�(��ȓa��I�D���ab�շ)4���S�? �qz#,]�����MY?�&��"O ���6����?v�|{e�|r�'
Nl� �;+��BӇ �-Pd q
�'�$(X7̑�1@z�K��Ha
�'�N��dJ/$����wɦ-k�"O��Q%���m�M0��B O�Y%"O0����ȵ
�"��n�Y�G�`�<9t�΄�j\����Ps�P��f�`h<��"��i9�DY��E�ǆŘ�y�\�m�d�IfiM�yd���Q�Ҽ�y��\�X� pš��"8IH�
>��?y�'��H@���+��%y\���'�P��w��\_���q&�
Vui�'>.�b��H�H�{��W:T�\D��'�yB��HԨ��Z֜9H�'T����*_9f~�0�gS����x�@�o�ƌpw�'%¢�zV&L��y�E�Q�����+ �"�����y��D.h��9;��}��8#D3�yR,Ɛ@�h�Ǫΰ7Z�U!�)�y�ϏDH�S'�V(S��DQ��y�dУ�6m��.���\��	�
�y���!�L�3�Y���)����O�"~ʑ պw�ЕA�?j݂U�5�~��hO�L����)5`Dx�(�<\�؇ȓMF��]	t���g虾2D��ȓ1}`��#e�.@6��η!L����}0Q7dіD���@�ʹY����ȓG�dbeִf<��B%PVu�ȓ<�D�!f/��`e"�"V ό	��q��]���)E�}9z���N�l;���ȓ��S�	E+]���26D�[�݄ȓ$�dM0I6��
��ߨB_P�ȓ�Ɯ�0[63J�r���=✔�ȓ(Hlx��ƴJ��b��C3�E�ȓ{���P��I�b�E\~�@}�ȓK���)]�r D���Ǜ�H�'.a~���a5�X�����8� e��y"/�f��2���Ж��d�T��y��U!x|0��Ҿc�A1C	W?�y��D�_�*,�PG�VT�S�"�y�A]���PVbހX@��Sh�9�y��Cc��A��ƈK�@1c�H9��>��O.�ʶǊ���ш�8'j��"O�l�b_'�]� �R/3h����"O�q�E�A�ɸ�-�O0��@ "O�-�'GG�~�=e�Ƀd!�t�B"O�}e� � �
�̃�s0�#"O:Y�%I*"�����*�s��s"O@��d_�dBFM����+px�$�!"O�僧�]rW��M��pI\�z�"Ony$�!��-Q2�z���!�yr�	�:|�uJ�T�� U�С̭�yR'�c;B�����?`���)1�y� �p���AV�ڍ�\)�'%��yB�J@/p�jrO2N�q�E�7�yB'�'G*��mu�f�,Κ��>�O��%j�	������D�}��Lr�"Ov��`ז+�T�s���n�Jt��"OZ�1@$X b}���M�Q6�y��"Oniad�2�rUa$\(#���6"O��x�J��o"�!C�[�eU�}"Oԥb�.�:P0$вۦwI��Q�"O�-b�FZ(�HXV-S�=�\zF"O� �p:�`<!�0��g�I<����"O���uL�	 u��C��K(��"O0P�)��um�(Z�i\�ȳ"OZ�#�lG��L��d�_	T��L�b"O��#���BDT�D�?J�tɣg"O<�&AI1xNh�j���B'T�Xw"O��`�aPEz�����"g>�)� "Oz�"��ǒj��� �T�f�@4"O�D���e���C  x�Ĉ �"O:X#��+�\��s�&i�6tpB"O��� �?A�@ {�H\51�V)��"OJ���&QsI�gσZ��y2"O��'I�&,�ȉ�׆�IJ�Q�"O����)U� t�9}3� �r"O�E�q��:3�p,9���$.�"O��{�eøl�n����4]��X�"O���X�����Դ\�� bV"ON��D%���ٰ�# e�[�"O��1�\>N���'��-�X
�"O�\#,�N*�(B�K�~��z�"O2Q��O�>6��M�aS�J����F"O�$�U�]>[��d�ĝ�u�"OV9(�c�2$v=0��\Q�\ȳ0"O��!`�ڛ'�	
4P�.;�e@�"O�q2ccL7s�V���'�:+$V"O��c��h�  rm>7���"O��Yq)˥����թF�{���;�"O �cc�5$=Zxa��\�sF���!"O���A
�;� 1��Ď79~�F"O\$3�ɪd%"��s�P�(�"ON!�P)�%Z��V��B�Ш#7"O�ɩ�C�G�!������ �"O�Xbpm
�+�xab��#xf$AD"O49����&2 8�K����村�"OH� �mނ<_B��ȜQ̙��"O^	��*�����E��W�*�"OhmBt.F 3��ЂZ4d��#�"O2R��]�/��+�����N��"O���!δ4�b�RãX�zT9�"O�ͪ�락(-$��I�T}2��t"O0�3����3a�ɺ��Q]�p��"O�}��L!g�T�b�O�)�Q "Of�õ��b�~��5�W��"O:eȖ,�.J��7N!H*t�"O��AQ�n[t��N0�2����$��l*�z��#��uh]�&�^�{A��V�<)��Y�F"L�q4R�M�Zqc@XS�<�`�'Ğ�;3��M��k4�IN�<���hi��Ei��3~R�ⷍ�I�<�`�D*a޲���&�e��	٦�k�<A���hh� Te�5���v��f�<9�&��K��	�"Ӿ}�b$��K��0=���7k���CK9	�"���N�H�<a�<�pyCmɫv����f�A�<9���05�<s�)ԿF� Г��I�<9A�F�lƂ�C�:o]xx3���F�<��ē/��9�N�ҁ�6��D�<�v�K�g���q�^1Ew���o}�<	r��&>���GV�	��
��_�<���	�n��T ���W��m-Y�<���-4VjE�rh��v���Q�CW�<YăQ��E��C�N+@d9�O�Q�<��\B�2QSC���&I)�%QM�<�t$��t�tU���� �Xi�6��E�<� yÇ�2'c�=�7�<�ܵX�"Oz�Ԧ�Db�#񧄎/dՙ@"O�lxj�F F�I�~ld �"O��!2�R+�R�s�M�"_��Y�"O�,�F�,�PhA��#5J�I(�"O|-�Q�.I�]
�
/�؄��"O��ӷ�<]1�,�4%G�vp>ͣ"O$�(r!G�OϚa���+4U��Kp"O���*$Q[��_�wb,u�R"O����9�X���nǯNK��)E"OLPP���GQ:�ZŇ�J@B}�"O�H�+D�pg0Ԩ��˞Uf�H "OV�+���z��6f��%^�Q��"OԄ��d��D��Ъm�8	b"O�Y���M7��h�SRFq�"O��[��p���Z�	���p�"O��H��,��x`�޴6Ī �"O��	WϜ��X�c�`Q

$@ݡ2"O:tIG[�X����"-:y0"��2"O�a�$d&�H�a�,#��"O���cERc(�)�2��`�t1��"O��R�|授�M��^����"Ob7H��@���	
 ^6��"O�AA��j�)&�P0^L@ (�"O�͘�"�1't�L,3O>�m�"O�%��
D�V�Bu���ڰe=B(��"O�(k�#ʏ3�h��'�"6#.1+�"O�(�g�0	纀{�'J�F���J�"O���aƀK0Hu�F&�6T�>3�"O��S	����C�%f��5d"O��BÌM��0Q�&p��"O -�U(��wm�|�s
֊id��@"O�x�-��a��d�T��+�)c`"O����l�I�����A���@ �"O@%�֦�C0M 	��Q�.��"ONձ1��LXL�q(�`�֑s"O��c��.Q$�Hbj�/ ��ʲ"O�R����'0�X� ��^y�s�"Oh��*дA��0vϜ o�fU�"O�h��.҄�>��B��e���"O�3�MՕ}�lM '��2v��QW"O�d*�'�r1Ѥj��*fu��"O��z��_'K�H���݀�R�`C"Ov�!riې$�V0�T~
=�"O�9"E,����e3W�U:�"O�X���ѐ\���m	�O�,�g"O� � �8�f��&n'2��}b"O�Ъ�C���a��у_Es�"O�aX���GR,Y�V,؆bpv��"O�`��ۛm8*�p�)ָE�0���"O��k�U�uH�a�7h���c"O��!#��� @2 	<��"O�X`e��Y��a���:��u!t"Od�
�+�%;����$��jВA�A"O
�l�6+�̰E�߶P�"Ot���#i�yP�> y�"O�z�(ɮo@:�0�l�h��h�"Oz����L�g�6�²��CJ��Xg"O���$�Fg��
� ݌4��C"OJ����W��4�1.̖j���g"O��sʗ^r�6)����tH�D�ȓ2��rv�C�.Ve'�6X��T���
�Q

:z��aaA�W��!�ȓ>��
��:�4����y�i��S�? �Q(�CƄ^G�@��D�S~(�(�"O�@h4I	GDL}1�c�Fq�)��"O��K�,L���=��\�eeXEj�"O�� �AXT
X�@W�^�jy2e"OX	�#K�LB��ҨK%ote�"O ��ݯNMt�󆚿+z�s"O��X�&Ѡ`�~A����>g��(%"O�u��"��VLx+5iف$yC�"O�D�(�v�9���ފEp��"O���('!~�S2jW><6��"O ��b�:XDd�!�I̕�4D��"O�Xr��Cz9��.˽U��ŲC"O,��P� vJ��g��w���yS"O\C�*H02x���(hԙ��"O(�ks��2eP�B�hߚRN�a "Ox�c��Э7|�����*pʴ"O$݉�l������@8���"O>�� �5��ɚ&�'F(]�"Ol�-nX�����@FI��"Or��Fw$Hh5���s)�h�"O(��ኼ;��M*��X$���"O���_���ᡥT
�❈g"O��RF�de�f�\r�J""Op��o�11���;��¹ d��0"O@�0Ϝb��T�������"O�E��	V�9t�Q�G��p|z`"O��`WH[�v���cHo�j���"O:�k��L@�Lp���H��"O�u�3dG�������>_��AG"O�A��F�@&�/��+T\ɳ�"O"}Ѝ�;b�Jy�O[8u> y��"Of	jV/�Q�ޜ�7�FV:�
 "O<�(�iR-AΩi��8:Y��"O�d� �S&
���ǒÀ���"O~�on�<�Bs.Vr�� ֆ,D�����wj|9%�{� ��7D�H����t��Ё3��&��27/*D�([�c J��r�'S���(#b(D�h����p!�p !��J�f�&D�T����5>X�U�2� w�/D�0c�I���#��2Y �!QL-D�(x'�	�T�6U� �T:��s��0D�,h��4S+�$yw��;� 
!D�H�1`�
O�����La��Rp`!D��vT�~��]� �L�$����#D�����|n��!j
? ,��a"�5D�,��l�4*�vh�˕�^T��1D���1k�HT�s"Td{کs��/D�h:���{���cH.e�0�:D��Q�J7^ș"1��}(�� 7D��3�	�Cl��9'/�K���F� D�@��*&v�q������A�*>D��S�ж?M�@!�đŜQ�т!D������ I"t�J7(D�y��C!#D�4z�拶U���h0�T �t� 4� D�|�BF�B-H�SR�R�b�����(D�b��k�� ǎҲÆ I�1D���u�	m0pA�T��%R^d�w*<D�#R@թBo�y��DQ�F1J�+��&D��9�(G���rR�Ɋ|&V(��8D���OӼ{16D9�#�
L �1H7D��HB*C`XzmH�JD�0�A�:D���S㍷#J)"vg���Li+��6D��cǌ�� ���ѵa�b�R��3D�� ��W�Җ-y�tr��/�f�0a"O�Ġ�h�ft-@AAV[�ʭ�S"OPu�#K�d�����OĒj[�"O� ��DZ�}
 ;>�|"O��c'*z���Rt.����f"O&|��o��1	�<K"-�}f���"O�(��M�< ��0+O��`�P(""O���sC��0�IE.�e��z�"O�pذnL�q_-���UR�p�"O��!�'�v�l�"Ƙ�`%�I�"O�%��2<ʼ�p��(v.l�a"O<PmӀ_n�S$V�.=�A"OH�x��יmv���*I�b�b�"O��3��ж@�c�m�� 6"O��*ĥ��P i�U����� "O�� �$e�0����[Vu �X�"O�P��:E��Jڠ���q�"O���'&&N6��U���;�&�0"O�Ř�gۇ{m�<�A��!mFV]{�"O,%��Euz`�ұ �,d1����"OF�Fŝ�aҊYY�@��x*�"O��(X�jW�<
A-��,�q�<�&�5�D[��:���+��F�<�D� rz"��S� ;/������x�g�5gf0�*%�Q�#ϔ��$e�͸aB��
��ub���A�T5��p�������'O�,�g9v����ȓHኴ�� L'Rdt1*B�4u �݅�"tHct��4`� @����4L���N:"Ӗ.�/,NtX#A�|����ȓ|� �`��M(}���e��%����ȓ/X�e�r�Ǘ3I>���ū����w�μ�Í�"�2�`�l�,P���ȓoH�S"�V����r&���J��К��cm o��q�H�zR�1�ȓ?�6҅͐�D��$	��CO�2�ȓb:L	!`���a�0�,U�;�$��ȓT �,�v�H0W�~�Є�Ċ?����&����{�X<x2��s�-��mE��c�!
t`��fRr��c �%�`8�,�X�@� �jt��s�XM tEBf�a@����eu��ȓ
h,T��ǌY, D�ʵa6D$�ȓJ�tya�R�N�y�@�43�x���j�@�!/C`F�k���?�����K��m(�FШ/z8���Q-F�y�ȓ�2uWFLb`%+�V-l0�L�ȓ��"j�o�h��� )�$��=0J�:vk�p�D�J�L&N�$\��)�����I�#�Q��#��?�,�ȓ{z�����ӊ@_���R&W�-��Մ����SC��N��c%�O�̙�ȓj�RH3��IN��!B,�<q�ȓ%^*Is��+69�9!������[�N��V��-C!��Hdi��$V؇ȓ!8��TÀ�lD��H��ƥ+�����7��u�������<���"6D��� �B�Y���reZ�m��tKCN1D��0���J��a�Y !:�!SM;D��8��Š`���P�ء_î8!#<D����Qn2IP�*V*qƌ�R�6D�l�P��e�n��6��U�����c(D�ԡd�,v�p���xX�v�3D���2�
>���Z�/�
,�8�0D�<D�� $��!fJ m�-"� �z2}#�"O�Mq5%�p�b��M�2Oa�PH"OPmZ�M�{?�Xs�͗�vH�8�t"O�5���1��pDmͭsF��"OR����y˄�4�ʙ[���Re"O�AB"`)����J�^��1�E"Op<��"U6T��P��4�H���"OPj�1KM�|�#�O�4���"Ot=�B^���L��/�y@�"O� �b�D�}�4fљ%����"OtA�@ꊺLx"��!f�D���"O���J�J�!�o~cƼ�u"O*ܰ�k��8��H�;Zp��a�"O$Hu�  U5D������T�1�"O�1��.K:,Ȳ]�����"O�d������
�QI�j9�"O�MzQ(�	"ԩ�\�Dz��0"O���!�%[�x=0Q��7FuH�"O@#�>=�D0Ps�U,W�e
F"Or|XiJ0K�$����M8?����"O�,�S����H�P��V,8!�Ǖg�J��4�s��Mpt+�?.!�$�1���е���f���jF�!�DЖy�6Q�O��Z��t"�)[�!�Vl�f��V/�2f��"�l�!��Z�i$���s#A�/K�|BAE�)'�!�M$=��	�	::��;e�(5��HE�D��?��t�W �p�a���E'�y��J7O<.�S��T�Rta�D��y2%2:n�8WG��F�n�x����'>ў�O3�{S�ʹ�8m
�o��,8��p�'~8ģ�.%#v��K�!����'�0i#F�� ^��������'�0��By�~5 5�����0Ӎ��)�t��J�(q�bH��c���yU�g`pEMB�E9�8�h���yb�ϤM�"p*�62�X�X�ޥ��O�
 Ǌ�:������"@�`#'�D�<�1�R$O]�A#D�_�h�C��@�<�w��}�DL��F�-x�!'I�u�<9a⬻��8kА��
��p>aa��x)��647>hHb�Y�=U6���	8LO��'���Q9 �X�.�Cʠ�cI�N�ў��e�'�>!�7�/����U�����T�0D�@6E���@1�#LR ��0@h0�	E��$�3���`l� qlܠ�G��qh!򤖻
�9��R�h���i<|��'����!\O����(-,���_3�u��"ObT�#�M�VB~d��Ή�ڨq�"O(���/BȂ�j¨�ɱ�'���[g�P>�p���E'~�Z�%����U!c�J� +h�
Qd�r6�I�<Q��_�{�(Uҷa��M���Q�(D{��鄪]�|���?k�T&fQ�V!��9K�x��%R�%�DY�t�҂!��'�a|b�ɭ<	D4i��D�M���@��y�N \��VhL�[Un��۰�y*҅Y�����P=X��h �T��y�D��f��� �ɾ��ˊ�ָ'ba{��1	6t(�-o�(:2a���?9���>O6��fcX�Le��q���L���ȓz��k �����	��/v��-�'O^����;4Մ���Ϗ� ����\;*��~�[�Ęb�S�Քy���/P�T���<D�� ����--I���ڤY: �#B��B�O6$�y�@-l���
�}�V-q	�')�k�FA�H0��V�H)n/�I�	�']1��/H �=��̫5�V��'�xacQh�KI�\T��=KD��yB�)��DV^���Y�A�p�DMZ��<B��$�H���V(��x�7��XG>B䉜�D��Iٜ2����ۿ\R
���<��/�R� �	�JX���u�<Q�%}	���Q�蕓go�G�<�g
�����yDdӔ	>6�p���i�<	Pi�#�"!ps�K�D���b1Uk��q8�Pi炘')'��S!oƘ��U���>A�4�~�ޤ��a�B¢(�f�#0����yb�֞T������h�Fj���hO���I�K����eމJA1E-A�!�$<����'C�;�Tzu�̸n���@��(��X+	�Y�J�!p醷:T	��"O�Q�kA*%�Ii��ӠcXI�>Q��"�S�'�!�6.��o	%��"(&�1�ȓOp�l�&*63���eg��{j,�=�0�0LO||�!ɓ}9�!`B+�2:G9��'��	9jl��§�Y0H��q�F�E�l�	|���s�H��m��KC�O�X�����n"<O�"<1u/
s+���f�%@�!����<᳂;�O����&l�4�"�� K�fMȗ�|"퉰��"�4�H��Q�.��qX�Y&-��U��Kp�鵀YH
�y�N��&�X�ȓq��dS��l�����'�ў"|�rJX�
�,�㶃N9WOj��R�<A�F�"����-�6@kJm*% |�D$�<q#+�!޺�{w�^���<D�(@���y
�q��D��M����`����&�X�<	��,�3�0��0�	P���Հ�y"IXB��<�v`�9Ř�б�P��ybގl۬���`T�0D��ِE��ېx&[�k���D�b3�8�A��(��B�ɍQ�������Ԣ�#+o�DB�	�uR�a�vkGA��i�.��D��C��?+
�-;�o�`S��Ṙ�JG��'�Q�P�<yU	����ɪFdՅ"Ɋ�(�NYu�<���~��`e�s�X��V�Eu�<qU�%�t�y���]!���@u�<	5��"��� /Q�r��t�<�e'��G���� ����RG�<�o[ <5��FޜC �y�I�B�<i�N�w;,M��.^�_�|٦,�g�<��ҽ[�~�����){�(����J�<��aJ� *8zS��y*̠��H�<�K6q��	ZW�*@�r*�lA�<) P36��A&6|��zy��'ܐ9r�V�6Y�cn%+ĩ	�'st�Q�O)�K�$hPi#p"R�<Q�E�!hz��W�Z;�%���hB�]�� @�@�vL�af�>��C�ɚ5}�A�CװNP�!��P� U��'4��JN�,�r���dU>H��
�'�
�ؠ�S
:lz'ě�8)>(b�'�VYru%�,&yBW�3�$��'۲�9�dvނ��'إ'mb�I
�'Ö�R�� ���E���4j�2��I�̊��)�S�7�~����U:P�
�c�%�3r\B�I�l׌�p%�Vv�)���?u6��'��$2����yuB[�����V�	4�)��'��I1�� ������ri.�#׍^���R�<o�b�'�Q>5*W`L#��H�b���ۤ./��Y�ɺ���>�K�<��U��#@x�[I�'�y�F�)�<@M]�{��ڃdA����j�'ט ��r�a>�S`L*k�|`S�%�~��4�ȓY�&���C��{6�͛s+�����y���9E�DBx�'���b="��h�4���~��h��If?1��ze�\�s*�0?�̃Ǝ9�Jh#�{��N��<�p_���k�m_�V���NYP�'�ў�B
����8U�����Ҿ&�<S	�'1DXd�;�T�95��
H<�0�����XD��[�q�P5X'I��D5��x%f՟�yR�@/=^T!P'	2CԁC��H��d"�S�O��Th@dX^kc�U�R0���
�'��|��J��'��0�IK�D	��'8�PvÃ�\�l�P�1P�*@��'�(��� �^��Ń����P�R�'S�1���z+(=P���#�ny���>�H8�D��TtA`��Y2:\���"O�1���
9H�����P�3��h+��'�ў"~��h�  �#N,�y����y"B�jo4���'��U�7�yrN
�$���ꣀ�<g���׊���y��Y�X�h����W$@�U�L��y�@=��)�⁯M�P�x�lɃ�yr��%J�+�+C� ��!�P
�y� Ś-�����? y�F�?�yr�Ҩ?�>h��CI�14�!�yBLZ�n��0����F]h�h�yr�Z0C� ��M�?/�n��.��y�אd �hW�	8,lv}�b�K��y�m�/���b��2��W�+�y�P"/�������b��(����y���C��(E�Q�l�.��受�y҆Q8Snrk2�!:���9����y�Ҳ��(S��˛,�\����,�yr��*s��Y[�, R�^<�$N��yR�/:��j%JO�:����m��y�
K�w�b����,��h5A��y�[<J6���@ ;,snI�q�(�y�,G9&����C�(_t��>�⤇���" �ЍT)H$i��Y�pم�`(�e�Tk���ȁIO�2��<�ȓu�b��w��4r4�R���v����g�qP6�"`:��@���
;�h�ȓ"�*E+Ո�%g�FABQl�7Q�vy��zQ�u�āԙ5M�ui��B�et��g��*�D�n�F�ag.)�.�ȓm܈RțQ�>����Ndq�܆ȓ�҄�!�̩Mæ]r7#Ă*��؆ȓ �<�y�.�0zs;Sت��&��Բ��T��Q����~�T�ȓ8;�H�c���N��	- �X�ȓt�`#���#���ˋ�C��ȓ0��OJ�*+�ͺ{���)�"O.�!�A�9���C����@X��e��[��'�Ȕ��X�
�Q+<m����'f��!���� .)�mKP�d�<A��E�N�kv`˰D��|S�L�`�<9��ǉ.Hp�q�3m���d�_�<I�`��xM ��m�1>�������V�<Qr��~.F-)�I� JT\	���u�<!򨇇8 �P`VMW�"�Ƭ�&��v�<)�"�6,>œ�H
�6��E�n�<� �m�Ꜽ"����[�y"Op2��V��c[�7�ZT��"O���pB�F"��3b]9�"O YȄ�F�e�2���_,���P"O�@6٢^?`�n�0U��-�"OnQ0����-E�*Ha�A"O��f]NC�PC�j�Q�w"O|D(��<�f�0�»D�"�y�"OHa��K�%%��ԀXn���""O�i�/38$Q�e�آ��"OI�1��2c��2��(�P]��"OL��BO���$Y@��R34$P"O�Piĩ��H;0�KY�����N��y�m��<R�׈	 5��2�yR�.:�9 �f@~֬�؆JK��y�$bq�]�EA���3g�L��y��k���ؕo�
E���v_��y�mW�
|�)���#"�xs��%�yB
��{e�B��<��D����y�/Ƨ]3r��QȄ�B:���k��yr,���z����5�����	l?D��K�+T���'��l����9D����Oĵ�����䎐;�v�"ԅ7D�p� �ۿHA~�I�>X�bQ(��+D��k �U�3v0��T�?�D�0� )D��b���E\���� ��%w
�Sh(D�����"/�b�"!�36�VuHу<D���d��<����a�J�.���&=D��9E������0m����M8D��k����V�Y�]�ܩ�Q�8D�ls7�ܓx��;�)�*	���Z"(D�xr��ƅno0d�"*�4F�@!*D�4��(n��
0g�:�L��m?D���5��T��P!��aj:X[!�Ō88<�TJ��@p~pa��U�x!��R�T�󆁡moDP�F_�r�!�O'HW�����U�`��1S��EE�!�^?A'
x�$�а^����c�/:}!�D� �ʬ�r��:9봉� ���h!����ع*��_׾=�3BK�w8!�ߌp�D%�!m��7�8r'ؐ!��d�4�����-6D�	׍S��	$)Hd�1��Q��H�Ӄ��<2���S&�ZB��<`�J�!R〨 4��Ga��7�J�'@l#a.�'hnay�Y�[߮p# #Nf��L4�	��0?��$�'ʤ�Z���<8�󤉁-=d\`f
�'��B�Ib�
�@� $�,m��d���R#>�L_��40��3�ӡ4��Sr/��L�>%j����N�C�	�+;T4r��Z�g8�0A&Z-(>�ɣE|�5��ƒ�f�S�O�\��0�a��Mpd͉�V89��'�����.�8��ǇAy
�@�O
�I@	N�� �	�^\(;�	I(6wH�r���)��	�z���� X&���  ��PsKM��Py:
O�d�5A �A����EV�Z�`���I�n�6 p��~�q��4#2)a���ί$v��2H��y�ϓ�
�%��[օ)uV+�yr@�nF�\��!X��S!�ީ��Y._{\'-��1�C�	��I��G�%�>y��Զ,���'J�mn��Qٰ��$����\""���+� $4da��̮ �	�+>w���4�0+�p���Qh<y�ܔ��Ԙ���<R̨c��U�<)R�@��EyS"S"98����h�<	7C�'U�P��&aNP0���_�<���Ȼd�T�
��Z����M8��id��*a1O� �u�7I�[�x�@�� �$TF�+�"Oh�3 \P�����fJ8u釚��ӡQȐt&�"|�aǫg�T��&/�5L�h2cGg�<�����S|�@L�)�`*�"�ҁWU�@U����'/>��g�'�K��@Kivt���)<+��I;^���p� �F�*�_������OV"L��� �.��G���
	��C�ĸ�Nޑ1����wW]�a�?��K�O�^�Yg��%oUc�<���.A��%P�RJt�t0�
�0q�!�$�* �R��m�&o�4�)ROB�*�ʴB�j�zݼu�֫��'�.���� ���I�]��9T�W�=����3D���Bɶ:� �)��:z���nۏo(�x�S��$�bd�'�X���	Q.B�8��04��C�HӥIs����ۿw�,a���]R&V�B@hA՜�S%	���q��X+�d�4�¸z ��>c&��Q"�0GT�(0����*d.�Y����~�@(������?t���l܉.�<�3 dI��y��ߚbq�$��G%0���p �U~���y��M�#�zD*��#�������� �hXWbPz�t�2 8D��!�N�B���:��e��eP��Bc��	t�
,P�$Y�h�t�,�i+�>�X��L�J�Аǝ� ?�����9��q�Uߟ��:w���i�h�V( 1���I?KkB�[�h
Yx�<3$���y~������1\�r��)��Q+r$A��&��l��cE�n��R?�
��G3=`0)�&^'^ز�`&D�t S�5d	r����P�C4�3E.K1�Nx�ǩ_=5
�Á=V�d0��ik�����	:hh1Ӑ�ҥ=�)"m4D��k��CryӠ'�pE 
�$��T�ᑤ�4p|9WD�!CFZ��U�HO��XuĚ 7w���H�)Mk�I��'�n��tƘ���XU$�0����b٠SM��"���-JvH��	�J.�����~���#W�7,`8HƏ4h���x�v�[�$�{u��.2hL�P�ޖj��S?
�&�Q���
��1+��� �
�'��}cu�

�n99��U��r}xb��5Sm�@�p���RZRU:mօ%��|j�w��<g��	$��'mY��F8C
�'�4��X�w�h���Q#z���Zb�S��Bl
:m�L���葽d�L1��,&ő��B��Q�Ze�9�M?O����f'�O�q�T͝�79n5k��_K�,�7��u�tH5���
�͑�h��z����=K6�(@hƬP���YEa��UXQ��K�E�<N:�0���Q���IU�?�Y'[,LnP�Cf��1_��(D�0��D��#_������;Wj���"��ٲ�ŷ+m�	�r�>E�d��M���2 JX*/m:-SR��#�y�ę�^��%���n�ZT.M���	�:8��u�P5ax�!h�4��d��o�akdK˒�p?��D�E��%h`��;Jr�m�eb��|8W�� c:C��l��"7���k+B[�I.db:�>�� *t4��b4��^��M�� �36���CE�c��C�?�0�ŭ�3Y�-Y�
 :'@���(l���J�hH3U�S�Os��au���t+��)�@ !,��'����d�o��b�)��u/p�yO�$�����V�R�"��'z.m����9���	D-[�u�Н��3��H�c;���;�a�Ow��h2��{��{�O�l{�D���<qs��&�jD�clU=o~�ʅ%�h�'�<P�1��qy�e�6�|e" '@�c�t�aC>���EK��p ��L��$l�:���p���K~XG{r,S�@"{�mC�k�"&>5K�C�jՉ��Q�Z��H�s*O]�E�R$�4���AX�5U� D�i�lY���v�8���
!�H"nZ,	88�s�*�La���T�s@NB��7R�L͸2�]�ͪen��^�\l;��'�V��Q-Y�a�UM�~Fz"��>X`�@R��j� 
���=�p>1�H�e�.h�0�
����vm٘UFR�h�^z������lՔ��d��t,����0	��5*�j���Q��,?&��#�,�P��UU/����)G�Jx����9h����ׁl�!�ğ%,�@�!Q��.� ��\�u���I���I����B�?ҧ�yG�:$+�q+��:o� 	� gD>�y"�@�	�xI�ஓ:9���OFK�������,�� c��p��\w�"`�ui�J� �$����E�6St8��� O�&���+,\O� �W S2J���R�oJ�_�t�j�⁌A�i�f�
A�4<2�-�*� aDY�i���(�#,O� 4�J�*��\�h�ŬY���!�č�@�n�@"AְQ-ආk*b2���Ȗ�"`	�]�O+�9���F�Q墌���wY�C≙O>-Iƈ�-]�杢��>!�ΰ�1dR�`�N�u�ߪ���+��LD*6�,��	�*�y�皁EƸ,3�"$J���I2�A��y�kZ� ���;�ˆ9_L�+��*���m��| t� "gJ
{)���EW4>(e��"��'x��$��`E�J>�B"<v=�eJ"\O�D/OH`�*��Ն�~L1&镇A�:�"�LB�F���F4f�Ne(�ïq�2�ׄO��ay2	U��&�@�<4���\�k�48ێ{b�T4s�E��Mv�L-�eA��~�DU[�!7J�� 8�A	R����d�ZK�A	q����xr��0U�Hթ�#�%��
A���k%m�i0�a�J* !�P���T�@ٹN?9R 1��`W�ͫAQ�c	���"O�[�h��V�"6"��{���ё���}C���g$~�j��M�N!��D�)��2/(�$�G	�("�4A��	�}��b�N��N�YgN�-1��$U�(��tҶ�w�<�
�a0�O�
��T5L��Ɉu'I�!p|!8��I�=���� e1d�A�����,����pݭ,��BD�L �y"�Q�|����P唹$�Z��ЏZ�yB�Y�VH�SR�9���0wgf�x�a��n�d@�CA/'�bC�ɻm��DӲ#%hHCܿlH�Ol@c�?��<9ń�24^ΑJe&�Fpv�G˚e�<9i�B�zm���� 
�T���b�a�<�PB�.$z(1c���!ZT�cNG�<	��g&1��� W�T#��I|�<)ajG$?��l��$��$h����{�<I6B�%��Hx�NW5�ZӯM^�<!�
�"H�v5"%�
��Y���Y�<� �f��Ss��	$�� �@2T�,����)�]b�='�Vh:�(,D���$\�\�r�U�wY�0�,D��E��n�� A<_E�铴�*D�� ��G�7rfe��&Y��-E`"D��ѣϻf>�\a��+g���&�#D�Dv�oO4��`+��S�.ah�%D�$"H�Xm��&J�0wkD)�F D�`�b�B����6lm:��$D��x%=	��<��j��69�B�$D��:C��f-��9���q�A��9D�CG����(%L�<"���� 6D�4�%�[�j)�I��&qI�4(!D��sQn�,a3ĀP@�\�H�Z��l5D�����5-���+ �I+�o0D�A��O�pnŃa�ٔ/�f�r1�+D��H"fZ�'�%���>�:���k'D�P�ra �I�`tA"��]��m���.D���D.S���G�D+m�t���/D�X��ቁa< ��@VN)���!D��:�H�G�L��S���q�X�S�H"D�0(d#�e�郡��a�����L#D��#щ��~ċdMߢ��I�C�!D���mZ�A@��<��-��<D�le�S�A�3A��`��l�`o;D��He�.P��E;c�V���B�;D�ఇN� �̉Ai�
k��p�9D��І��("��{�m�=w}�@�6D�p �
T�Lu��)Q7e���7�7D��[ �mF2�`��(w�e��6D��;��]м{�Q�I��G�2D�`x���qO��4��&Vv�)�0M"D���h��?��E�e"�)FL~�sT�!D��G�6ޥc�I��;�N%s��-D�LS��1C�\��*j�����<D�ӥ� �Qj�@�Ɯ�Τ��A1D���H��aU� S\�h1�i,D�Pa�V/ R��)�/�ؒ1c�L!�� h�rC��B�hU�$,W�l`$&"O�尃0%�ݨ�̗��$()�"Ol�)v�-k�Fh�u+�T�|�` "O:���K'T�8�@D�5�hY�$"O�I��Z�iԦ)#�כC�r��""OZ��Ĩ)�~����:�R��q"Ob�q+�)�Պ��ʤ`�^��"OHp ��\��1���'.���"�"ON��##�o�^ �����.1!�"OK��NXR0��œ|g����D��y��ez|��$�$!�"\Q1��y"��/jl%*0/��r��V��yBW=�&��@��. ����yb�˄G���a(<i��yWl���yrJ)%G��+d ����#f̍��y�!�5�<ㄩJ��Y26%�	�y2��0�H�J!��.�}!���=�y2�=��0o��W5�qz�)��y����k�����_	G4ب$���y2��S���D�AiJ�iE:�y�(�;>|����8C�t�����yR�ް;�u�7bV?
�L��w����y��U/z6iɧ`�} iS��L=�yB��}����� �~K2<a���=�y2kˮd|";�ԇv��!�Ť�y�%F�N��Ȅ�X?Ѱ�Kd,މ�y­�>JR�XW�+h�K�G�:�yR�Z�j�Dyj�E�1K���EBý�yR��5�1)�"_&�S5N�y�j�6�T�3 Ă�T�p�ā�yrfQ7`�v����Z�p��T��y�oW�-��@���>1`siƗ�yB�X�um>ݑQ�\�A�fۓCЇ�ymJ=o1��{P���	U�u��5�yrʂ�M�$�%: �2�_o�<�0�Т[��Y�Tj�g}���C��q�<��!�9=��`�N
?��,zg�e�<��C�y �`�g9'�J�Ȧbg�<�mG�vF���94F 6bGb�< (ls`c3�ˢ$�Jh�`�e�<Yd�?r4\�G�X�O�X��+Sd�<	�aϭ`�h�ƙ�SB`�5��K�<��jT)w\A�fÊ,*YT/�K�<�a�܋�2i��h*
�59���D�<���S"�Nᑅ,%v���H�A�A�<��o���3����
����V}�/5.T �=E�T�đWzF�{��<����J�y�j��AZ��JuKѳ����F[���ɢf4$+Ao�vX����fث}]�c�Ѯ1���X�$�O`��"_<7�ސ�;�"q�ݠ�sfB���PxrC9q��k�a�x�-rQl���Oj���4xE<����k�84����Th�$�K�LE��y��!%���"Z�~
�ɇä�yr	�E$�U��@Z���9-G\���-\6'd<�Q�ڰ��C�	�DK,D��Wc6(C"�D ����D0v�׷%�D����
P�@t2���m� pfl�+�a~�lE�H�N������]��H��ҹqB��ҦT4T����xl0A�S�ʃU*��a !�+d">F|"�',~~}9���|ܧdɦ]IFFK,H_�!CE��\��u��}��4K�o�cin �d ~�t���,a���K$�ӧ��м�Q�J#xԤ��F�E�^��"O(%�s��3h���i�ESD�p��%�>Q��'6���˓:j����b��2vL>����I!pp�2 @C*����f�H�aA�mH;��� l�C��3)$�M�u'
�Hڦ�	Q"O��rQ�r�`����`��h*2"O��Z��W�zBХ�P���6�ֹ2�"O|;U��C(t�Dp�ƍ�'m
���KPy̓F@|$�3��<k��5�#��p�ȓ ��)�TH�JT���r�ã<.0��'�����E��Fxɧ�4�6�� *,Q1�M:;m@q�"O��1Q$�=j4�2 �E2:#�E�r�ߟس� �(�^0�C"�%)B��I%�:Ց��R�M��Y�i��`����B�M���P$� W�~�3�쁡:Y�8	����N��pe��?7����7w�>�A�BնF��"��(H�TH���(l�Li����k��9�e���EJ�+>��/��y�F�1���y�/�29�P �d-X�K��J�EЃs��	�H"Nӌ]ۄm +[ =(���O�|�� !P��e�#�U\iaV"Od�����4���N���e(��V�>������4�����\�G����������kb�G�N�.5�6s��{BO��T��Pc�
���	+7+�Z��q����}|�)��v��D��	�v�p����g�$RWGG;X����@wk�-���4-ǯ:�4Y���4�F� {��ߠi�Q��!�6�y��	0�������!dK�=�Pd���ԸP��ʪ\�j���
D���*%!7@|Q3���	j<B,'D����I
oǨ��(�%h��S���+o���lڭ-�H�Y�:dɈ�i1����	�ɗbV��4��6�B���ɤH��V"�̟8��[&-R�Y��"S�����ɁRߴq�b��ux��r��:��X��G���:��x�\#t%^�"u(��G�1�h��Q?�Ȅ���qM� �����f;D��Hq�v����v��"jà(9bN��/��0'̿l��8��L�&�L�X��	d�%�O��v�+e�6,� ��G���y�NP�R��2$mc�m��	����Ġ�,S�D�q�6'ظ1���O	^"=16���@����G�V�P��
ZC��̈��}��)��E�*�"t��
-Rx�CͶ
�H!s���E{����'�R�QR
/0���S��8�RJ��r� �tA¢�v��0�J�@���κ�{5��X�I�Ο�y2iLFZD�𨖱�p`bunQ�V�ʤ���D�	�n���$S�Ju),ʧ�y��fF驵��ch�S$����y2�;G "Wʁ�y��[�kȟԆi�s���q�@a��ٹd���!��;E
#=y����P��D�&MΠ2��PK�0y2�ՈN�^,q��δA]b���U�k��bƭ�/8�\��#KZ����^��MS�D'Fdā��IAB�<i0dD_��Uk��ĦDf���'�)j�NG0:���!ÂAʷÜE�<I��]�6�$� �[zl����F?��a�"4��� 3}��I�$N����Ʉ�\�E #j�'6�!����`�I�3i�RXY ����f�&��r��#(���F+~�q�䍎1�DZ� F9��~r�N"�^��@c�'>a�f�'L�Np�֊��	3l���r4� �����~�iҫ_�I��aE}���	gvR��J�Z�'9�T%�w���"�p�� N
�B6��$����2\5Wt��wf�;Zּh��䦙�㌌�0w�ӧh��A�p�P8#��Y3Ã�P�<�`0"Ona�%X�][���Pb��g�*P+��>��D� �fM�v=O��
T��;�a��(�|^��!�'!�YIEʆ5�JI���6E۔q���&�6|H�
O�Rf�Ǻ�X8hd�:
������=�z$s��	�v+��gH;"�T�P���!�d��w�j����N,���L��!�fݸ��I�8"
-X���5~�!�� B�����:@pr�K�?V�!��s-�LZ��N6$�P�H-b!�Ɍ Z69 ��D4̽H��H,h!�D�)s����i��(��	%��<W�!�$���I1֡�V5�}I5��!�0��%�� �s��s��!!��	�:C��!���cw�$����*w�!�d:8��6ȗ�_m�p�%I��z.r����Pܓ�h��� ZD1�Řa=�t*����	z"OX�Y�"�_���i�N�����iJ^X(��\:8r�&���JW�usb>���mTK�A9!f����B1��K���Iu�6?�\��2O��2!�@Obt:d�G6s�!q�W�RbC�a8���PO),O��P�o�s]��s�Ŝ�0�;���X����&���'$�k��ˈ �*`ܠR���0Q��u+�5�B���͐x⧔�O����dhۛ���q'��tR�������37$�*QiUu�}�'jF�g>M3qiM�d�
e�6LظmEBC��95����'�`_Z�Y�!�,�C�i��	�,J�9H�	�f��5�䘖��禑�B�Q�	r`�Ҩ�h�|u*`d3\O� Rg�["Y�ɜ'	E��^0R���v��6Rr(<1�O��zFG�^N���c�'g*)Z�"�g�D�+2O��Hv�{F�%1��y3�QR�Ӥ<��#���+(��s�O�&!F �e$S!l��ĩ
�'�X|�QE���	�U�I����nS��I���'݋>��R�4�*��t�T�e9�I���W�nl�E8�"O452��y_hA�F�g�2=���i@�	cO#�a}��(蜱�O�K��2��}�����A/2<�	���P�QE �Ty2G�B�,B�ɯ+��XS�$/����`�j�B䉿C ��ѣY/ml�u���򄆕2��b����"&t�qC���>v!�C��4��%N(6@�^�dz!��j> ��IN�W(�Qr�cZ'F!�$�8�\=�Q�ʉ*���C�	�!���.l��T��]%���sKO�R�!�W$L��8 ��P�u-*�Q�T'�!�ė�DpN1#��
C���H�f�!�$ѓ=��,���RN���GI<`�!�ʯE�~���T�,&�!SA㞊x!�
�	QFmB���#�l��B�=FI!�$�La�\�6-N!\)N���0b%!�$�|��#��٪D�ؽ�7��<�!�D��#-x� ��r�*�Äb�-@�!�J^*!�\$s�Z��oް\�!�d�5n�M ���"@�Rl�#�R�w�!�ć�Q�,R��>v�u�n[�2|!�$G�h&N"�Ȁ 5{䐃���~f!��[N+�X0C�������ˑ�{!���o�X �A�Z��$�Ѫ��gS!�d͋��@�h�T��I(PC^8YV!���i���a�+�[���@3!��z��8CH��H\�1��3c�!�D�{50A�rMԏ]Vh �`Ȓ|u!�$D�KT��h��_�?��B��[i!���|��("C�7(z`1���
+$!�dX6Q�B��sր&����C�!!�ֻT�~y������c'�(sc!�d�Ǌ���A�:U�.<c��L<mg!�Ę�T*7N�7}������x!�$յP��gH��#~(tC%��Xk!�$	$;���4D�
!,��!dܫ3!!��2�Mr� �LA�͚�!�$�a깩S�b
�h�BK�!�$^�>B�R-�����@K�@g!�.,�����m��ht+��Q��!��"�铧��_b��j��ݜv}!����x�;�f�D��-��,v!�d :���u�X�olJ|�1�A?R!�dć��-�CX����� ~V!�1Wfy����0NF�j�Q�;B!�[D@�������7-��I�!�;bi!�dϻ6=��`Ā�`	ʴ�L9R!�D���nDa�(«-oH��a���Y!�d0ֽʒ\K�0��9S���x�8f�a~
� PQ��*՝4ąV�]�a��Ex�"O��ӕ�լ�wJ@!U�@ �B"O%��O)B�j�t
�-�,�"O�)����>f�`9���t���"OjxN�2d��Y��3\���*�"Oj%"
�(�x��&êK�H�`"O��z��#RV����%��$F�(3"OTE)E�OL��@�J	�� ��"OF�B�\7w'f�X�Q�D���x5"O$IB��ǦkV|3eG��<{|Ēf"OF	�Ϣ&�(;7�)zy�x��"O�)���֖��R��L	S��p�"O̸��GX���n�2[��s"O�L5�U$d�Є�&��)��ZB�'i�A�֩�@�$ӵk���I_��}�U�Ը|X�A�a����S3i����вS�}a7�ʆ,�.�6�K�)'� �Ҁe�ş�ݶB�D�ƸLWRh� �9�vh#4�xb��d��y�L'�Z٘bj2U;N4R'�Ǥq4����͟$[�4�y"��� ^~ם�ӈ����O�	V�@�H���2
�D#!�Џ��Ղ:~�,x�����Ob�q ^*,QY�`�8��eK�OPe�p���:�E�ş�"}jcФ�"ѱ�d�$	
�:Q����:w���4�>E�d��/s�M[w�2���qd���>����"��4u��Q|���OW�D���B¾. ��$IV�@�!�2����'pL�{yA���O�������N����M����'.�p��$�<i�0�_��}��h-[TI!���6���{2 �|�<���D�>l���b�=YĶ��ȓ.)�0rF,O0�Y
'�ٝ!1�u�ȓ�$0p#�G�J��D�$Ohm����0�چ�jخ����J�Τ��`춨��@��f��� 0AK�y�ЅȓD�b��#���5���F�����ȓ
��˄>u�N�`k�*C����ȓ-V��x�n㕓��A��e"O�u�T-W&Y��5o;�h8"O�!Kk�0��0	��0"/�i�*O��I>�t;�c������'g2��Um�}#ZXぇV�ssJHc�'�čaR`Ѱ�FY`���4< �[�'��@yCω�p�a��6.T���'�t�ئ�H�/�RT+&_8-�~Q�'0�$�Z�_E��kU'�	�X8
�'s$���p��1��Lu��
�'�U��R�S�4�6��.l
�'_�����!'�{S�;M|�y�
�'Ě�83(��L\R��"s��0�' qˠ��gB�yC���j����'�hx�f^�w(B����1c�԰��'G�U"�@ڰ&.`;�E�S����'C� ���őg`9ȐK��E��'�h9�^�X` ��J�rp���Qc�<ɷ%ho��s�j��EW�<�Mʼ^V0 Ӷ���pt��O�<Aw�(��(�ܨ;��u��[G�<ٕ��S!}��"�-�D��,�C�<1�m-7�5�!A$��w��@�<1�dX�mJ@����"=�Z�W.Yy�<���#k��k�v�4Ǩ�J�<�a˕v∅��[ �F�*�n�G�<91ʅY��X �i �>H	�� �o�<��� �z�b �eE�$j��u)"I��<���R��Ep��#	� �cs�c�<�5!W�DԮ�7eƥU��p#G�Wa�<1��G� �!U���K^�@��[Y�<I@پ�<��em%%���ZqZ!�� X��b�V!���52P��S�"O�SR�^�7.�8��Gw'vY��"O�Q��ƈf�
����;
");�"O���E�*`���4FD.�윩�"O4M``KәO'P�!&��3c����"Ol`qf�����9���d\I
�"O�)��'XƦ	q�3Pn�}j`"O��q�ߞ3o ��Aa�\Apu�W"OeIh���<I���m]�9��"O��+&nG"G���y�F�T��"OVXi��u���pd�D=�b��e"O�\)e匂g�4��D|�L]�3"OH0[�dЄX+��:P��4���U"OR�9�X[�Xhrd� G����"OrH�hT)zLm�u�S$T�B�"Oز�n?J�F	 ' �\�b�"O����"�A�4�Z�!=~���"OBL1���4����Đ
/2=�'"Oi;`��	l�Ҳ�I�H��"OZt2�J�W�t'���z���!�"O��Wcʊk-�-�F��vZd ˓"O�aK�B�p�|�#%5YG���T"O��A�'7���:B	и6��A�"OԚGh��^���#�� <��	��*O��Kp�h�6��Ƭ��m}���'(iIw �&Qt�j��eB�`��'�f@�%��-�p�u��S>H��TW����yI�Ă�W�1�܄ȓB�dC���h[ԑ��͚;L�x������[)���^8<�f���`��HynH"�r��X1�<�e"O���􂓋D�e�@�{n�!�"O^����+�vQ����8X��1T"O*�֦Ȇ|����$�;�@˰"OT��e�ѡ?|0���^:%4Ҽ�"O�M�`�|Vٻ#�	 ��9Q"O����D�!mj*�d�#qR�*�"O���@�ӛ%�!���
^�D�#"O���jN�mN�"Sd����\�"O���cC!�0y��b�y��1�"O�-�@�n���!���R��"O~i"�'��M(A�����^0Y"O���C�R=I��\a� �g���!"OT��4D�+/
���iZ3g["O�q4Jʐ!�\�1�κ�X��c"OD����A�! �@���"O�Ia@yj@�� ��f.�L�s"O�m�"m��gw��e@6BD�s"O"�:凘�%��/�6/��k"O��`�h�(k�vI��J�,��`"O�|�n�	|��Ǥ�3ks��f"O�Q�%OA)pf1K��$����"O�����0�����4}S�1r�"O���Q@��7NHHgDoL��0"O� �N3S"�L�#�.-x̸�"Or��W-�.c��*dC�<2(X܋�"ODyc�/R!7vTz���'z&���t"OP���D)_@2�c�@\�S� T�"Ox@Qa�4%���Ʉ���8t�G"O�y�� ��ψ��t Y1V�(93"O�h��.d'}r0O^�P:ʥp�"O�,p�ψ!V����Ӕ+�R�E"O��פ��Z�jQɑ��%,��"O�q�� 8�v�8��4#H)��"O� �YSW�Pw�v	�AX;5�8�`"O��;��O�:jE�d.�~��$��"O�t���>P���L��L�\�r"O<`�X"iY�X��J�=ip�"O��x��&l�� ۧ	�|:���"Op�O�9��]��F�:�ҵ"O���V�2E��0CK�x#ơ �"O~� �+�� ��x!u�D�JE��"O����B~�lB4�,=��Z4"O��DZ�+F���A�ųv�~��2"O����&AL�8c@I�!&��9I1"OX��4��6i������7�����"O�p�m	����AjK�Q��"OJ��coD�#�f����)+>nMF"Ony�`�b��h��ɹz+hA+�"O�(�c�H��Y�C��!b\��"O��)+ɤQ�� �	R$�����"Od�挏�dB�`�X�q��8�"OZCO��K�d���n�f���+5"O�k�*�H�R5��c�Ȱ�E"O
��C����ɐp�3z��a"O4��4`��$]����+�!_żA"O�9��)N�f�r J�[�q��"Ol �d�P[V ��Ɨ8sZ����"Od���'N;2�i��Ȃ�4�d]3�"O�Z�%ƍN1`H�v��V� ���"O6��n>K������=Ȁ�C"O�J�BY*W��K��3E��#4"O�I'�	'l���E9[� ��"O�mѶ*�jfUS���B�"O�����)�ۦi	
ead� 5"O� �+�ּ�+�57_*�I�"O��S��^�:���@�	%#\B9:"Od8�v쌵0�z� �&eIRq�"O\��eч�\�p�Ň
P���"O($�b��B�F|�dg$su"OF=��DK�1���# �Z�6�Ұ�U"Or1����23�d�{�D-����R"O~�ѓ�t��� ��d|�U�6"O�,��&�K�`e/�Bl���o�!���5V���d�Z ]Jj(y�f΋ !�7n���@1#7	C��R�C�K!!��O�$(z�H��-/������'�!��9l�\$���8~B�cD��y�!򄈯E8v-yÅ�$8��P$�ݺ$v!�D_bqAba�j�� �O�"!�N�,M��s �=�����2�!�$�j9���P�K�H'�E�e���H�!�d|���Z�f?��S*U�j�!�$N:n̪dy��	;�uH�X/_!��a���0��Z\�+6�G� `!��QdRR�&BR�`�P=�%���w�!�D�9�(`���\�d��OZ5�!�D��C���Y���a�Q�G$ՈSy!��S����
AjP�pȴB\� ;!�4%�,����Ɔ�5���ˉX!�d9�^��Tň�{��xVϕI
!��M��P�0�M�[���i����!�A-2I�	�݃,�R���(˙�!��oY��#E !z�A)CHL�w�!�
��2�[7�[�4zdȐg ,�!� Rfb=x��|� ���hL�p�!��(mfI;�N�Z �p�bGW!�D�Q�C �Շ,=�Ց�$�6B�!�� ~���h�GJ$<�Wb�4V<��{"Of�0�旤r��hXt`��'���"O���'#�-Y���ZQ��,yzݳ"O*��VoPbVF%qeU�<�B ��"O,x�`��;Z���U���\$�yP"O�dZBAY>�tH�ry�6"O���ƕJ����T���_�5!"O���q\R��9�ț�g:P�"O����Q+	�tbČȲ1MLH�"O��FI@/}	p���'zX�� "O���Ac� qHh��+��$W��"O&�YE����f抧%�QyD�k�<�T)�2R������@�E��A�<q�aE?&>� m%)�4do�f�<	d ǭ��ʔ.ϫ,B�;��Xc�<yf��y+�c���vlM˰^�<q"#M���0z��$z�$aYA��W�<y+	�Q�J��@�і;�-IQJ�I�<��%�an(�)a
f?���$�\�<b�!�
�z���=����SY�<Q�]�1[F,��M������T�<iV*�e���c1M�Ue,P��NN�<��o�@�¬Y��>����o�<)tH�?E?� �㋒�|�<ͫ� �o�<�r�á
q��'���1rs��R�<��`�R��q�X8 ���%'�Q�<	ƭ�7=�|�g.{�.�ءN�I�<��h�*]R�m�'��!4gHC�<�4�
�����U[N�����W�<�Ʀ�7   �