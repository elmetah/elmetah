MPQ    Am    h�  h                                                                                 ��C=����.���e�u̐��=��.׫�lVҏ�c�8����IDq����NN?n�z�Ƌ9<��=�紲�K!�c�����q��[��Adr4���ݍO�=��p��~C�/ e���_��X졗V����e��W&��j	Y�,���6����k���z㫏8�������/��a�J >���1��8���?���%ebC	If"j��8���u��*������{h�_���U�A��8�j�l� ���󳯊���};drF�ce������d�elé�-_��>�6t����rwJ�@��~d�g���J ����V�O	�(�$�_o �A���
2�/�i`��S�&�A�;u��,��ђ�bd�6��� e����
�Zm���2:EՎec�����u�9JMܰ�{$ՈYM%-Q�(s�
F�<7�1�#�ϣ?L�i��Y�a4mx��
gTdL�z�b=xC��9^r2].�n ����;2�{s�,զ�8�hA&䢑�S��|1*S�)�Kt ��ڥ7�	(5���_��wA;��1�@P�ML?z��[��tG����
� HF�YC���UG�K��ӭߪ���i�q*�+p��	[���#����;��6֮�ӥn��7��?�>�	��(\���/�uDЪ�w2?�/-���YB���L��f�#"��� @��M��H."�������D�q=XΘ�4�Ϫʹ�Wj0�x��� 7�0��t.M5��Ń��g��%�j����(l��M�ò�)��9�]i:p|�Rl'���q���X5�������~ڕbpMH�C7/O8��ٛ����\�%��9�o>%.�����?E|���΃��}�d��C�E �5���H�t�D5Ƴ��q��~7�D�a��*~l�,:V�i"$�2��9��%$�4������a�\�..}u�M]ܯ�jF�k�0`�Uo�s0�����;1 \�&���gf�i��^a�u�*��Vb���\�A��3�Ԅ=�y(y�G��@���z�w��B�7�(M���z�B��~�-\�K{;���E�sA_��x��c9��A�<9���[͇�.`������2�#3fo?�fQ�ľ�jl`���O��H��%��!'BvV��/��#��-[72(��$��[Ɂ���;���<��3x|Ff��C�D�Uz��Gq:�)T4����8��S'cJ��aB��6�*�К���	.g�@�0A�(��3��F�MF���~��X8��(�0K���
F+��s�x�U��f�wgٗ��n�-Ɣ��` v�ȵ]�=�r�w����]�a4��{��Ӌq���Jm�=$�{��|���[�U����G����!��/4r�C��RȾ?@~!�쟋�EIyl�zw��]�6f5��ح�G.OF�p��;c�������P��p�%EG�XXBT�{��Gܡ���{����_���&J�(�yFHf����6����D�-EZ�����
M'�gz��;����ec��iT�>���0���,>L֛�܄y�!�qK�(�s��f͞�"���QB��%�ҧ�ib�WF)0'�P��*��g]V���۹�RC�`���w=�+Z[�S)�*��`�g-Ee��s̲Q��fI#xkF��>��@�4R)F�}Ǥ!��a�W��_^Op{M2_�a�Ug5���ײ́*���f�N�k.�3g�7k��f��W��`^ܓ�!K�a7)9H�!��C!u1"��p�>R��+�WDW89��̗e/H�;7>�_�����0������>�����{��C�ެ��e¸�!��_#�4�jN��V^��n'��i8�eN�w���/���.������ ��ԫTm��s�i(�xE��p�l��Œ�b��AƔ�}C�e��
��	����c�ڶb�������ƴy"�j�h��IhOQ%� )����X|M�+���qr�EHl���N�_gٌ�:����2X>�
��.U�J}hf��dP"i�#ur�7�J������+���Zs�7���'�ߙ�&���pTo�Y�vΐ�����q7^��]ƺ6u�ۓ�˹��-�R%@:��<��1�MxV��-���:ϣ�@0vXe2�3�aѬ����۷���L.�,� ���<T�����cfm�m]��b�ݴ�ϽGM��$km=>��D@n�������LMa	��Y���{���N�.�
�(Q9E[�E�M��:q4�'���$��o{��͂�E�97�c�:��ov�F`%B-NC ��{����6����T��[���9~l�1�US꾃&���k�A�N���g7y�I�K�܎�;X��G9�2��Q�ؿr�o�0DNj����� �S�u�����姇Ļ�s3����r�	,]+�W|��`ܺ�_�:7��6�?�g�!�����f0�7��}|"k���	���꣧/&>��ɯx�T+B]��-���9�*qoE�B�3 �!�`M�����</����_�m�sw��O�vLe����ӋU���Ts�o��q�w�r�g���H�h�'�Ee�xՌ5t�J�㖧��F��IaN�:6��}�jP��$,�7Q\��@��t�"d��U���	Ϣ,-�m7� z_G�eȚ�(�֯_�q^��;��T9�=��P��L ���xU��B��y�e�(�!B�dnq��(����Y�a?|<~4ٸb����ܸ/^}�w[�Dr�b����]QB {8�������(��$��R��q>�ii�B܋�D�^��{��I�ٶ����\΁V��[���f�C�ϐHUp��4>�J�l�A��59�fS��ϋȤ��� �$�5�k��aI�Y&A��+cә#6'�k�*��!PS���h,wJ��YS���H�h��WT�&�xo�-4�+�sj"��~^�N)�+�+dc$Ŕ�����p�C.�X!���9��;C�Ůlʃ������'O}1X�F�E?�@K�/J��)L� +���6����6��� @$��5;\D.��{p�8�T�k"��x4�D9M�.a��j�O��D�?��oӖ{'��(	eӻ��H��kH��e⾄���V	;�� �kXl׽  ��ѯs�$u�%�d䷄���)�����	A��۾1/zMw��i�G�M��a;�yE!t���h���Mj�=�_̵���W`b�Ry�ı��(�����NMǅ�`�G�\�]	˳�Ơ�@�'R��lR�n�OOx��ס�¹���LU�c��ٷ[/�l�f���y/�K1���/�9� m8��߃U�uY@%�3�8Թ@4xO�E����y�o�q�n�'�*7<�Y����󻯋�t��Ǉ$�U����q���<�HeL�&��ZΕ]��rEP��c�Ǿ����ȏ�]7Y{߈�YhPZQ��s�E/FR
��w�1w��҇}�Ni�����x��g����F�=sb�ߔ\W2�n;p�;hsY�%�A�W�c+(���$S�#�1E?O)��qKO_ R\�@��	#�y��@_ww�A�Ԭ^�PdWY?�Li���o��a{
j��F�E����0�
K�ۤ�z���Zϼ�Ա++w�	*�g#��+����јi�λ�D�B7yc�Z~��RD(7���cu��_�r���-V����]��w��Zc#]��ؚ��ʔ�>!�.�C{ٗ��L�W��p �j�%����Ws�Z�(����d�] ����M�*��~�lgZ��%����l���Í`M���3]�&pw��l��%ۖ����۱'����ܦ�wPb�V�>�/�S�^����T\L����m�V�%ɭ ���P?�~⒏[Ξ��}?��`8Ӏ�~5U��H��Dib��X�ʑo����S�j�B~�Ci:�ۈi[��f>���E�@�r4<�����%��_u�Q}73�j���K&(U��s�ګ�k�_[ W^�XL�"��i�3a_�߃WV�le#�AΘ��/^w��}�y���4`x�҉{w������M�)r��1B{(~ �!-�n;KV�2��������Ҩ5�N��c��A�9@�[��0.��#���-�~��o���Q"��3k�`��6O@����*�%����|�L�D�V��/]#���[rH��w\�VZ��M��;��1/���?3S�.�5�����}���Ռ�G,�p)oR��;�8��E'�v�����1�+���ϟ.��ݎ\���g3(4���d���
7�T�����K?+�n��|�ޮ����3�a��g4��fԮ��K�9�g�0]��mL6w�y�KO�_��?�f.��T	ma���vR6|c���Y��p8
�.����Qy�Ēxrx��M�?�[O��(u�`�lc�����qԧ5F,��0�O��g��O;�#i��f���k�BE�CiX�fTz7Ë����cD��0�����tJQ4yAǐ
[3��ٱ�uD����YB��rw�L��S'h�zTu� C'eޫ�D��y��k�T0��,� ����y�X�q��W�N�fD"2�AQ=�cl�C48�rh����+��e����]QN��6�9R�SG���(=^�,[�R�O����:%b���2�s��XQ��I��k!+�>6����)A����M�8a;��ڤ1pVc]_����_S5����Y�*���f��:3Bhk-��͔���7���<�K���)T4!~��C��8l	*�ZbM�����pW�c�9����sH�R�7y�K�9�J(��ՠj��>�L��u���h�C��5
���YD�%��#�����`�eҷ��+�/z�H��`Q�w)�/i�I���R�[ ����Qm�L�|7�����+6���� N�_����}޾7����d9���n|����U�L�ɀW���$��|��O�Q�w����|�.���符�E�'i��}�_��Q���c��*؝��»�͝���U�qHha�+d�[���و�R�-�ME ˼���=��Z�!��P7'K��TsG����T��u�Q�%�R��DQ�l��7��ي�L���euU,득b���a-H��@5i<����~����ցM��;v�І2Xa��=��ׁ��/��g�V,B���Wӗ U#���m�F���b�����PDMw�kH����f	1�[�Q�6�:��a$�YU$�{�Z�N�
8<�9 ̴נ�׏`Eq,���K����|o�K��nQE|��羦d:���v��%�OC�G�{���m*��0M�r�[t�9��a1ex�S�0z&WR��X�6<��W�g�K3I�u�	>�Xb"�Gtw����w���m�[N,��|m9���S9D��E��%��3���s�	}/�+�����.S��*������t?��B!���y�0ͭf:p!}#����7�䀭�^�2&Y�~�DI6�x�+<&�{�E���͜�/ )J����q��'�:�������q�_�V(.�m������{�@,�ΔU�:��O��o���Xg���u��0Q�C� b We\��x�̜t��-�Q���'�ǹ�&���ٮ��j�^�77��5���(я\�dq������(�-1�,��OG*�(�Zi�ʷ���ݣ�ۏ_-=E�RPԮ�L{�t��D�a���̳@!ن>R�B,�q{kp��ǉ�2�|m<�%%�=������3}���Y0�rdD���]�~w{����K6 A(�6$/��qYņi,ʙ�s�L^�2�u��Iߦ��a.P�CT��q���z�ȳ��5a�j�Uk�~����Jv��\5�SԘ΋��.Y� ����kw�YI� AlX^c��6bP���!K�p�HV
wy�YnE�� ��h[��W���R-/���΂�"��^��,��+��UcI�O�/������'�PC�AL!�*^��];� C��ƞ���\�7�xO϶�1s<���Ӓ@�n�/�VW���������
���96ul����m;��_�8mװ3�����c�V�_����#<R楢9�e�:s�o.�%'��	���h�T�����>e}���ίdU��
ts�콛�b۬D��uIXb�_j��m���������[��l��Scz�����G-���zݕ�8�tT�C��߈K�=>h ���gW��ڪ�ߏ����4���P�JĥMb��`�.�\$)�n�2��i������S�		�RYM5�J�4���\�¹�m�L�,���隷�1���j�/h��Gtr�T �m�3���UQðf�%���8�o4�^F� B���-iy#=ɛL�jn�?�*�[�Y�ޠ�BfF�F�M��<x$��T��菬����Tez*�%�Z�މ��ҼE�5<c͚L�N����|j�!�{�\�Y���Q�e�s���F�C1S�P1z�P�Y��8+3i>�W/xtg���Ű2=n����z�2��`nV?t�2�;�;�s������^5��XDS<��1`Kf)jK*�%[����Z�	�ӧxN�_2w�A8	b�'9xP?�v?�+���+jgٷf �
%UF����óѵKL��zm����'�!+�:	E���
#�t��0��l{����p��74nu6����(���uzK�m��M��~x���B~�5�#���V����$������*�1��Q#�'���Ҹ�}�W�6E>j&�]m��� ����S��Mk���y@�gl����qs��إz���h7a�%~�]��pr��l�\��Q��&�	��Ӳuۦ�4b����9Ԁ/%�OA ��\� ���<�Ǒ��%d}#����?����J��ι�}��؛�8}ӻ�^5�)�H�p'Dį����#�:�1�E�~�!:O�Ui���D�ʿi!a�[��4�N���H��h��d/Yu�u���aj��q�f�U�es捣�Y�OI۽ RMN���y�i(aPa�ߖ����V�kR 
�A�R]ߊW�����y��D������Xw%�T�mgyMͮ��04pB6�K~M�-R�	K1�҃�g婚�������5Ac��LA5u9�R[�q.֪��(��H���o�\�Q��䮋D`�$�O{�V�~��%��
��Q���\V�o��s�#��Q[�~�� �Q�̨�u;��J3N2�N3.h��vi�yu��x-c�0�RG���)�����{8�$�'��х�ɓ�,VG��ǫ�A��.�)�	�/��u�3c�����"��L����kZ��fS�����^��g�B�W�\�-g�pj!���ȔƔ��Ph�>pW]�#��h��w=-&����j�ӵq10�A�!��m��qŧ|����Twoɋ���$�� ��r�*�H$o?�X��b���{��l��@��@T׬b�5�cw��9�O�ߢm���>��F������|E}�X��T�a��F�á����q�;�^�&��J�_Fy<f�e�mϬ_c� ID�)>����"21"���?'�(�zJ���eY�f��û�Ot�w0�;K,�ԩ�@|�y�qA�)��fC	v"�T.Q8���ۉ&��2����&����v�J��]L���R��q� $�=٬�[��ʓ��c��}U]9��sB�Q*�jI'�k��<>q~���o�)<o��ZZX��a">��U p1�_&���x�5��\�hs*k��f�
�aq�3I�kh��/?'�.��IaKL�h)o�!���C�l"�EҦH�Hf���ڢW��89�S�̍�#Hd��7��+��@-��G�%TU>��������J�CN�����1�̱@��N#^���~����W���Wu��w�[t�wp��/$s�d�{���� �5�J�m%��w%"�.�����ߎnňs%�:�]<�I}y���\����wR�M���H��T�*쪂����w1�OG��b�e9|;��5�����E~�����_ײ����[b�(ᒻձx�1F�U*�kh\Ʒd��ә^��m�x����˗)%�xe�Z�7���5�'��?��l�ŐvTe��,"˿�p�-,�gC�7\����bu�a��xG�/� -�A�@0��<U��ã(���Ɓ�ڣ�@�v�[T2���a���L݇��ཙ���,�w<��;���G��m� ��b\5�IM��Nk#驣5g!���7��;���Fa?��YЅ�{�� N,g
�ow9�rJ��}"���qG&�����	o�͸�Ew���X:>dv"5%8��C�.�{Cc��lw���m�
O�[/9c9�
T1�S�&�n��4)7�4��Zg�>�I�܄��X=_uG�O�1�Yqҿ(>�(�NG����Ek��]SYN�=S������qb3q�K1�L	�R+�]���>����z���q'�?Go !����}0��%ui�}�C_����?4>���&t�	տ �S�+w*%�%D��Н��O����Y����T%�u���M	;��;�_8`2����ŉJ�l�p\��B�U;�X�J}�o^���'���,�������(�%|e��zx�,�tW���Bj��?T��?O��Fj�H��b�7Q���Ѫ�'d�'���H6�d�-̒���E�G�������/��g5���ʥ�=�
�P�o1L֌V�f0���<�o]���y�%B�5�qv��ޑ�D'򩗻�<t7��I;��t�e�A}���f�rFP�*-P]G�:{��� CX�N�(�1�$]��Ȥ�qt�i�qËNR�^��i6Iړ�缺���kV�����%����ܲ���rUfT��J13�w��5/TIS����>�����t �
��닿k2�I�A��\c��r6���`z0!F�$��cHw�1�Y���Ϧh6�wWʵY��-*ʗ�)�
"K)7^�u8g+���c�4��po�
�2Ԃ|C��!���/C$;�T&;��ʹ|��Aᗒ$�O�21����;�|@Ѳ/���_y��էp��l��6)�����;Ҹ���~��.b[�!˾8}�z��~0�����w7���5��o���'\�	�W*��SJt��j�enf�Ɋn���Җ����ɽ��ۇoe(�Mu�~�Z)��>B� o�7����@��i����
z��a��+�G�N0�5yt�K}t����@l��L�=ِ���YWf��15���ҕV	��Ž�аM��D`�5�\w
	�)b��R��6j��>%�D �R�K݁E�k��o�3���ALK����0L��S��y+���/u��<��o��m.ָ��G]��@%��8�i94.�]��������y�*-�'*Lnx�*m�lY������fj���0$ ��]��K�r�7eu(j��(ZDG��RZEF��c��J�Y���F�#Es�	�{UPY��Q4�s�a(FȜ	�X41u�ϴ���i���� �xO^g1��K��=i ��J�a2��mnq�"f�W;�/�sρ��wg��Y_@�mCS�,�1{w�)���K} �&�v�	�����i_��AS mԢ3�Pˣ?+7�,��e'f����
��F��@��F�ŐKM�㭰���Pм���+���	`�ih�#���k��~g��G<��N7��f���z�(�;�Y�u���h5D�@�D�9_��iͽ����^#�Cv��i��	���Y��S���L�ٍ�T��f�I�����x��W)����#����Z�� �H�j�Mh��t�)gǼۺ�^(�/U+��{�C.e�`PE]:ipm_l8I9�yG�AF��hӍ�/bA{;�4�/`�
D5�!qW\B�ت�e����%�l���f?V�L�W���Z�}5�p�~0����5��_H�%D���ɨ�>�K����� ��~ ?:�Fi�,H�w׿$� �v�42�ʰ���rs��_ku����jw�ꦁ>U}k�s�������vX M\<	���3�iCR�aU����*RV�l��A�,|��p��F�3y�{**�N��&w`����M�S��x�B�s~6�-ͣdKɂ�:D�DwX��h<���cjN�APǍ9�
�[^.�s�Sp���۷4��opB�Q8<��)�b`�t�O��pr%����2�sfV��%��#_��[��7����L����;D�me���̜3	�؆��X�s�]����G�n�)��V�1�	8�u:'/n�2���'����!���.�U	݄��q�3�����N��
M^&��5�d� ����$���Q��W�Bg��;+�A����y�y��]SX|�c�Aw���ʎ�&����~��\e"m���lX�|�w��Mɦ��$���v��:��r���C�?Qv���tٖ��lYŇ裓w��O5|ٺ��bPOWc֢(�w�Y�i�\ӊ���n�!��E��X�T0Ս��-�ӯg����9-�X�,J���y7%��wh�gɱ��dDy�������]���ͅ�G�'�z�>9�6;XeԪD���c��)�0��J,Oɓ����y'�q�aZ�E f~��"h�Q3��6� ��)P��������!2��f[���Q]G���8�Rt_��q�=T�6[u�ŻL�1�]X��v��s��(QE �I�b#k�`	>��
�P=R)7�~ǵ��S�a=a�Бp�c_a�ƽ&�+5�/�����*&�*f|�B�3�I�k�������E�ܤ	�KG�)��!t��C���74�AW�CH�<��Wuݎ9�7��<@H?�>7����o��b���N_�+>����k3�L�C�6-�k�M��)ٴۅ�#J��8~�[�������:�/�V�w�MN/�`R(�HA� z�1�EHm����r3i��M	ڡ� �����wO@}�Ð�5�
��2V:�+��K'"����eU͂;%o�r�8Ob/�Qu��+��|�9t�����"o)E���;;_xd�k�}���4��U����#�l��U��hW �da.��Tb��,�C���rؗ���gZD	]��:�'9��ʲ����T�Q�|���uzj��b�7o+#�=�]�	uK��SL��j0�-~��@+"&<���~�����~�C���m�Bv	v2U.a�~����L�虝�x,8c^�Z�!�v�D��{bm�Q�n:�b�̞ �UM���k��7�p(p?��3������9aZb�YK{p�XNg3A
n�^9�9�V$-��qb��ĵ��zeo,���S˾Er���t)�:�`8v=�;%��C�5�{~E"������M�eK�[���9ω�1[�S{t�&�[�ɳ2�6�ghQ�I/*���x�X�!G�G>���d鿃���VNb	#�r>il�S���ؽ��ց����}3,�Lӄ	s�Y+��:+����9�uuU��ύ?#�!/@�o0�Iu��}M����g藚o��%&����:�5�.{+�N���z��臭;�v�������
x��ְ&)��E��%�_������ud��:�����}"�U�q�E2�o�&/������
����`�j�e�q�xƬ?t�h,�Ǉ��],���Y�����.�hj!�r���7b���M�D�ŖVdgx��p���S�>-gU���[�G��
��J0� �0���.�̘�� ={8�P�P�L1���!<���k ��Ch��lꆴBbΦqq�e9�����U��)�<�hA��e�1�� Ç}�|���r�gЮE��]�WJ{���;�8l��(�s$���Q�q�-�i"9Y�)	�^B7�BIՠ��g���� ��Ʈ�\�~W�P�ݠ�kUa,&�EdeJ��憒ּ5��<S��\�y=)�d�� ���F�?k�_I4	lAb�'cda�6ؖ����!A=�����w{
�Y����chI�Wt!�I��-%Hτ�"��^�P�v1+u��c��b�ea<����ݚGC_�!ᖩ��;�jvˀ�T]�������mOE�b1�~-Ķ\�@��/��|��?�񘇧�b��'�U6D��>�h��;���n��)ǘ�|Ϩ�ǧ��n*������mI��3n�0�o���'�L	��]�^	�OXd�j�e�u��ą���Q6Q�#o���8�b�c��us�U֫�#��ZQ��R(��Q���D���'z� ����G�����4���~7ta������mY=t���afWqA���x	��/��7
�e�����oM�@�`�\�\����3��\@��8�ß�ƖW{R�j݁@�o���ҏo��5�L��Ȭ����=��</� O��#���m��\�pYy�&��%��48��4�M��v$��.y8=��]n=��*��Y�d������cˑ��$�q��gŜ�"{���epF�7�Z�����E�\�c�����
��b	.xHu{d�Y��Q�"�sm�Fv��/1p3�M$��H�i9
k�MZ�x*��g@�!���=d]ߥ�2I?n���;�C�s

����T�V��"S��f1���)��K�;��G��6	���.��_��AnW �N�P�4�?f���`����
���F";�n��ڛK��Q�K�����j�ݓ�+\�	{υ�z#[�6��h沢��´�U!�7���������(Ȧ���u�FP�cv����{�����L��8�m����#���b��,������gM��T��݀v΄��;y��s�[W��Z�M����ն� ��a��Q}M�6��odg"�غVk��J��p+��EY��B�]�A�ph�[l�U����\������h��j�b��/$;/�U)��f��<��\�[G؅�)��M%�|���i�?�E�� ���}��ԛYH��1�5&��H���Dz�ӳ�.�Y�w�0D���ut~X>�:�,�i�š�/d�߈$��P/4�k�p��M������u��H}�j2/��8U�T�s��E���32+ H�fi/�S�i^cba�(郖�VN�Z67�A�&��@�e�LUy�wx�~\�cv�w�K7գj�M�2����B���~Q��-HnKK��B�u����s����)�_4`c%�KAk�N9x \[9�Y.LKj��ת��귏\�o+HQS�X�,M`^��O�x��B%���Ǎ�.��V�=���#:�5[#K%�H[H�G�(�^�9;��Q�9(��3��HRY8¯�:�n�t��ގG]�)�l����8a�<'O������"DT�<tV��.Ӿ1���N����3ٙx����Ӡ��e���v����ߨ��p��_�>�x;�R��gE���K�5jꔼ�l�����]���^�1w����Ic��ﳵg���$~�}m2|��g�|t����p�����i��QI`�u|>rI.�> �?���؂�ٱ�Tl�Ⱥ�~�"�P5o�����O��M��J��t�\��!۫b��\n$E��+X�}T�h)ü�;��5�g� ������AJ"qy2y6#�"Sı6c�D�ҩ��Tۯ��*H����'y�zz�S��Q�eOڎ����*$�<U&0��,��}���y#�{q7�-��cf��"��Q.W�����tT��ÎVp������w���]BN�G��R/��6��=ϭm[P�� ׉��b>S��ђ�s���Q`XI�4k�+F>����*�)2�w�c���aX�W�K8!p�d?_�
��	�5��w���*�'Qf#GmW4�3�j�k���e�p�|Z���K�(�)��x!���C��e��܅�>J���=�W0J�9�;l̃��HW�7*Cȕ
TZ/߯��>�#�>�F��^n�Cēե�����6�#��E������p��Z��6 �Q�w&�/�nU��|�é� U���Am[|�ma���:��\���y�~����9�ͪ}�/~��.�u"6��y��FcX��%��Z��Ơރ�����m��O�r$��FQ�|�����]E�q����_��!�&61�O����ٞ�d�U`��hRZ�d��f��$��uG���p�M����$Z�����_s'\�h߅�����T[����E���Ǫ�]>7�x��|P�&?Wu�,$�.q3˥��-��@&�<��9O�����|�H�>vD��2�=]a���H���w����,�nl�5h�w�}�mᢹɪgb�2�;�jMv�k�V��	S��-O�bR��k��au@oYƨ�{Km@N�#
	7~9� *ױ�����/q}�������ogѵ���EmAi��:�}CvXW�%.K�C�\�{�G�ݢ�u��G��g[�h�9�(�1֟0SVF�&\�)~�-L��h}~g#��IJ��zF>X�8�G%`��g�w�����g:N}~~��V3G�'S�B^�sH���_~�'}A3�*Vg3�	���+i��uYp�R�r�p��'��?��g!z����0^�T��}�����j���?�b&�חյ�w�	8�+풽�L���.�*/1�������Om�ܐ��u���V���/w_���_������bʋ�9���|hUq��@to�n���_������e-~�x�L{t��B�x�57
ۦ�ʮi�j��7����׸��cMd����K(�ώ:�-8��G;{�������ą]�9�����@��=�3P�QyL�����gՙ�eJȳ�BK�賂B���qlo
��Ǻt]�ͷ�<j���*@�l�*��}��j3r���`��]=��{�'�vq�L(�Փ$��>�q��Ni� [��8^}�)F<^I��
�r3�t���H���Y�R2�;c�U\$���[�J����U5%/�Se�담���g� �p�����k���IO.�A�Q�c?96j���!<�!�Y��w6�Y����h�˞W@R]��E�- \��ߋ�"� ^L��+P#�c��J� r!� �$�8>�C !�|�%v5;��]������������H�O $W1�O��1Q4@���/6�M��&��R��&\����6_I��~�C�;H���	ݰ$LR����w���/�t%L�J�V�o�P�V�+o?�'���	�[9���9*�l4��eN�(ݿ�vud���%Ġܽ�U�=�����u�?�P�
�~iY��k�m�i�������J�z�����mrG>�I�������t�	��+#�9�m=B���ݏW�<�>߁�0괕97�@���H�M3�`��]\-7	˟%�2�C�,���z�8���(R*�5�;��EjT׍�JLA��ȇ�G�GجЍ� /+}��x+S����m${��K���aN�%T�48���4���1�p���y�e���ßnxHm*�zY�ס�S}f�w�p�'\�$��BMo�]�=�u�ek����:Z�xg�"�ME< �c^Ӗ�Ϙ��|^�7y�:�{˗cY�<`Q1�sH�aF>�v$�C1k��j�*�i�iT�S�ȳ�xP*g{YYŁ4=_� �l2_�n�bW\�(;yw�sE�SխtE�O��i��Sm�1�/)|�K��{~ڬ�D	�ɧ�k�_c6;A��Ԙ�fPо.?���b��[T�w�N
Vv�F4d����n��K�\��������8��+�	��i���#6����C�=���Sg�v�7e�����p �(�1C�n�uK���^�ޏ�n3�Vv�O8ͳQ'��3�#I<�'{6���ڔ,/ɶ��;�ك<��a6ο�׊��¹n�W�Y�o�j�
�B�P�h ~@v�Y#M<%�j&Wg}����>�e���r��{=��T']p��pc�l�Mۂ��w�űm��C�7��,bw䀑*|�/�[瀩�W��\89 �`��B��%5�ܝ~��?ȷ�{҅�
E7}+��4�,�l��5��LH�ڴD�WG�D[�to����T��Xe~�|�: 2�i�~�Uq��l̡���4(*�K�ڟ���5!�u����dj�ɦ�~�Us^isw��
A46 C���E_�-iy�WaK}��qҍV�)�}�A�@�ߛ ���Zy	�. ֈ>�wֵ��>�M���Aa.Bg��~l�-�X�K�����z�L�������c�cA���9�U�[��.�˔�_%�Y���6o�m�Qnֳ��`9tpO,d�O5n%�8o����G�V)hEv�#�O[^ᆽ���B�H̹�[;�	�����\3��q��}�Jo4�ia��A:G��)�
T�'o�8<w�'�gÅh���4���K�rV�.�G��zN��o�c3Q�T{������-����O��Z�$rW2ޚNR�E��M��g���R��P�G�7�G����wF]�!��Y��wN���V^�9 ��y��a%��m�[�b�d|���념���L2�B��,1���_�r�x6�9��?�����̩lO���Y��]��5�$*���OTE����ޏ�W�R�7�=F��gVEN�X��T�e�w��	|+��Vջ������
J��Zy-�v������QDtDo���t����e㥯���'��/z@��l�)e�)E��t�e>0׶�0���,h�q[Oy>u�q�v�����f�J"�Z�Q)����G�/����0��U!��+C�Q���=�]=:���-�R�ꉎQk�=J�p[+S�;�g�N��,H;ssV�Q{�=I�92k��>"�*��8�)-Rl�kC��
�as����3p���_�[�\�d5�'/�yƍ*��f>���E>3���k{�� �i��o�ZVaK}*q)�% !j7_ChпX��w�b9l���yW���9`\��j�H��a7e��������XGV;�>3�:�a�x9�!C�����M��y޴�Ԥ#�o$<�Q�K�r��pƈ�L��w���/U���ҩ�>2� 0���K�m�v�h���?H{�Y�0�����4���O�k�}J�0��G��Z����a��AD(�5x��ۇ΂q���h}PO����^�a��|��j�r��瘷�EOV9��y�_.a�Ꮸ�4�����̻f���#hU�K�hMԄd��ʬ˱��ʩ9�c�(�M�)d�Zzy���'����@r��f�T�1^н��>�r�CN�XQ7%*튳wg�A�MuA��	����-���@!��<f�A���b�#G�9]e�#��v��2��da����]�ڷ²j�Ӷ:,.�f�1��m6�׍m��$;_b���V݇M�hk�Z��
�u�������&�a�>YAj1{&^�N�+�
���9�'t�т�LLq��z����k��o��E͉��Eh\�*,X:o�2vs+�%���Cg��{�i��=T���>��[`0L9�[1QBS18�&CGq��R�(�����@g�֗Ie^��3mX��
G`�J�P'��K�9�:YEbN���h��"(�S
�d��n��]"Ă:e3������	i}�+D�����������k� ����?x��!:刴e�z09e�&6}�e���o	�P��J�&�-��0����-+(��燐���v��h?��9�ሳ�_���&孒�a��Y|_I<����Ќ�y���!���AU�
�;��oo/��D&I��e� Z�˯ENUdeȪhx�Sthǫ�=�	��˹�|gہ�Ю���jW�g��B7� ��q��Pd]yk�&������-�:t���5G��l�F���6X@��g0����{8�=���P�rL�������(����p4��8<�*W�B�_�qg[��s��uK	��e�<�+���ʧ�I	6*�}��{��nrP�{��]��M{]s���8v���(�Wk$nt͓�
aq�i(ɋ��g^��7�U&I����#�/s��݄iu)o�4{K�����&UW<>��rJb�B��j�5��'S@����F�W� �S>����kc[�Ijs�AX:!c1�6N]��1*�!7yj��KCw��Y�ED�
�h�n�W{P�A-՜�:$�"|��^g��S�++q�c5��ś�����ԓ�C�<�!���?�;]���ʊtd��ؗ��cO��1�@�Ĭe@b>F/q�0-��,���u^��.6z%?��:�;�ׯ��s$��28}OG	��ܻ���q�y%摷������&s�o��'�P	���T�3��o�:e��ݺ���)���>�=��?����;u�b�K�E��.����ш�G�����s�?��zT�&��>�G���f)� E�t�!��V�t=��a��y�W'X���e��KHb��Z��X%�6�
M��`
\�})�Z7>�MΎ����U�z��%�R��6	��ۖ�H���~�L�J �b� ��z�svW�z��/��3S����gm�}H�&��Ü�W%���8�aA4?�d��L���y�a���n��*>�Y�j��o�2�Y�BQ$|�J��������C��ef����ZuA$�=��E��c9&�
G�����_v��9{��NY��Q_�s#�VFyh��o1f�G��ч$�-ioVd�C-�x��@g�E��r=Z���[42��-n��ׄ�;T�}s��q�H+�J����i�S(��1̻�)���K��GU��G!�	
S��_(_�nA�%���xP�h�?܆���YV'��ҽ�
� FO�'���wdBK�Lɭ��l���Լ�b+�#�	�Iw�#���?z��E��	��17 ǩ�V\��;�(~�:
u{u��s�YX&�Qk�j��r��.��롉#�}�³���4��j�B���I�������b����G�q�6�i��W:Pp*���%�Ą��) Y�Z�?��M�3��e�g��r��������f��������]�p^��lI���=����S�����v��i#bɇ�%�e/q$��;��r?�\�6��;0C�}@�%��ߝy�?gj͒6�O�%�>}�7�رӧ3'5\T�H��FD0%���d�����&K㫱[�~��f:�W9i�WI� ��Up���&�4�Z�&@���M��б2u�E����j�,/���U�msR1��E���	y >Io�O�� 'i��a��k�L�cVĨ�l�A�z��|��wuDy$�L�ݻ��.w@����M�t�nB"�~�)s->c�K�v�룜�ͪ��x����c��A���9n�[��e.�k��$X��=�E1�o���Q����M�`$GOg���G�%���C'���VDP5�a�#�?�[��\�~6i�=e��;ue�����3��*ȻW��WF�d]����KG���)�����8(R'�3|�X���Q���-�
.	�Z����J%�3O(����H�ɤ9�aeW�����Q�շ�M^Y��0Z��n��HMjg��=;,kH-��^�"X�*e�]$��T��w�
ʿh0֣4�]'�ӭ����mh[&�]��|* ��@.����0��:�9��b�r�?�4\!?b���N�����l�/��4L�ט۰5M�U���OOh���Y�1ު [�����-�ҀE�F&X�,�TA�@�2�C�$�I�]0������	�JXN|y("���Ϙ�5�lEhD��E�O���/u~����v'/�z��;����eE�g��m仠x�r8�0�O1,`fR�,;�yYL�q-1y��f/^"9G�Q$7��G�O��	����][�r����t嶔�]8�����TR��ĎlX=�.@[�ϓvm �ȇI�U�s.��Q�hTI�kh!>]W��!f)(3]��C�Dpa����A�Rp���_�a��%5������*W5�fY�Mw�3��kT��͛����I�ܵ��K8L�)�~!�9CC���m��C?4��M ,W���9+���y2HФ�7�G5�@�g�(�����s�>N����
{fC:�b�<!2��QK�쫬#J2'('���e�&����8k�v��G@�w��/�'�מ���N U!6�0m����cg��u���1(K�%�t���[�(*�}�ې|��+�z�c!��|�Ѽ������Q���N�c�OsY`���|��|v(�MY.�Ӌ�E�9��H�_�m��	��O`\�sͻA���U�jhHn�drZ�Ӆ�V�ٍ���������dNzZ>���	'���*�1��TQ�6ИI�y�K���SC 7�Y��n���\�u�wQ��
�ч-O��@�D<�9ҫ�z��>|W��]����&v���2&Da�p���2a�}�����w,��L����'�����mפH��bHd��q�Ml'4k��B�!,�\���T����a�\�Y�K�{o NX
?~e9�N��g�͏�q���	ꆀFN[o���$�wEc��]�:*v��%$�CB
V{/�Q��� �ۡ��v [�9 �n1��SJ<&~���_G�#<R�l#g�I�I�(��pAHX��GG�����������G�C�N�ȍ���+��2SE龵����{����3]��S�	� �+���s�����f�P�݈�?3��!Up9���<0#�a�-}i��#ė�A����&��ի(���+c{&���o��7�L�����!�.�8<:�<�at���#t����_������1�"�XIW��7�.�U�b��62o�����e�Ic�{t�ˊ�i���ec��x���tæ�������20�+�p�\���G�j�fv�N(7s���~bm�^�d�)���P��F-8]���](G�ŭ��;�QP��Sc�]y	۶�r=L�LP���LBN߻R��C���[����N��e(<B3X�qbg�J�>�0BY�4�<`�6�����%�э�}��6 ��r�鮖Q]3�A{8�����=ɰ(���$�Uu��q�1i�O����^�9|�fIƇ�(,X��
����J�=���!�q��URt4�V�<J�����}5�Sy��*�#�5g �V~�WU@k	0I�غA�BPc�H�6�p��̤�!2G���w�TwY����]#h�1�W�n1���-nAϕ��"7x�^8����+߀cp��6�3��b����jC���!2��)�;8�U'��%0"��=M���~Ov��1�Q��'�@=�/�Rl��S��&ŧܮ��X�.6�!��]����;�!��?��9���g
7@�����j�#����������!�o�Y'H˵	������F�+�e�L�ݵ6o+��҂����c���n
��uP5a�F�\�4���ѣ����.��ղH�z4z����/TG��c�!(�ؖt�F���߯�R=Es.��57W�����_�f�7�
����R�qA�Mi(`z� \��	�i+�h7"�"~��00��R`��1[��l��f!�8��L7"��=�r���`V�u�\/��m������m���O.�׈2%�O�8�I|4�����v�5��y� v��ݳn�*�َY�O�	������]f�$�:F�����d��ު7ea`gH�Z0*E�X��E2�c���EQ��i���oY�[{A_�Y
�Q���s��F�A4Z��1a� ����Fi�,����x��g��ŷ�=U�&߶�w2zRKn�ĬRi*;/?s�~c��M�EG��SS�11�g�)r��Kq8l�O���b�	�ڧ?t�_�U�A���Ԏ]P�2�?�%���`Qg��-�x
̫mFjH�y^HR��K9]ӭ��������r+��E	̶���#���WZB�sȄ��f��7�3���f��(Y��E��u����T�i���"�%�Q���ͩ~��|�#�HR�]��������?D��wJ�y���n���5�k�d�d�W�f���@���F7 4��z��Mrb��`
�g3��Q�������a@ïI��L��]���pY�9l�:b������B�	����Ŧ�Vb��&� ��/̻ ���rɍ>\.T����Ǹ�|%kk��t2C?�,#���]�@�}!�ɛ�O��⦫5�.�H��D�O��l���m���]��~�~	Y\:V��i�P�������44��ڟ�� �kb�u�	�Y�jc�8��jKUiѝs-�ᫀIQP%� 9�Mz ��Z�i�VaA���'�	V�Gk�A�Ԑ�Q5�2:y?,����wL�1�t��M�'O��ɭB�<~�p�-��HKx��&Y��)���h��p��cV��A�ρ9� �[��3.�+���B�����KAo\�Q�����`��mO�z��z�%�$TǞlR_	uV_Xm�#˺�[�m�����8`}�o� ;0�Ѳ|�fM3u�s��`p�_ya��PG�ɞ)����8��d'  酞˖����Mgw��Y9.$�[�p��%�B3�ѕ��n��V�vR}���+�P��(�p�3V�I��C�ogV�����皔-���)`�erJ]�j"�O�wRg�z�&�-����ӈ;H�m{ �X��|��x���o���S��`�&��rn!�/:4?�+E�	�$�J>lE���f��	5��y��F�O�Ĵ�f"��Kf�H���!8��vE���X���T����>>�?ȏ��)û���D.�J��y#a~,1��S����f�De@�*půI~X��߯j'�W:z�QZ����e�(��f�D����00�$!,��<��:�ytC�q��p,�fj��"�S�Q�e�f����1�����m�M���g��Q']3�B�X�R`�C���=@��[�2ٓ��9����D��3s�wzQ� SI���kCL�>������)#4J�!d�A�a�-C���}px�2_M^h����5����/=�*�ft�1��H3d��k����6����N�#"K�K)��F!`P`C��:ҭ�s/ӟ���WaP�9Fu���H�{E7��ٕ���U9�����j>iG��W=	CukG�ׅ���IT�G��#NCa��G� ���k��E��B�w7z/�W���[�4�� �,�q�&m,̊�^����mڍ*�f�W��0���c�}��}�w�
��+]���ٗ�e�7�^�보�Q: ����^��O��v=�闣(||�(2M���E�-r��7�_�ݲ�W���j1O��g���XLU1�EhC(�d�S�@�ű�I
�/����Þ�XZ��u���'m
(߶�c�L�ST�&��s#������]�N�K7ۨ7�)��w�2u7Mj���=�V�+-��#@�q<���j@މY�/�/~i���v��E2���a�VS��G�84}�	g�,$Q�Ƙ �b���N��m�U
ڻ�b@{��c�M��kjF�\mt��{�b�s�샜{naƚ�Y7M�{ܟNS�
�Q-9╼���؏�3qγ�6��!*�ow�Ϳ�E^V�ஒ:哽v�3g%��2C�{j��s����~ ��|'[��9;�	1G�|S�{�&����[�䟯y&gT�"I����n�X�o�G�h'�8/��o�����`~NΝA�^`Z�0S�lm�D���¹��8�3�T�w	_�+���&���#L��aٜ�8��?�12!p�[�
0� T�'�}��g������s��>�&�9�&�F�r�+�������3��E�b��<��~�K֜#��T�����_�n�����Lf݌�8_bv=�iK�UBd��1FKo%�-ºŹ�/�����e9�Ŀce�cUx���t���r��t=��g&�7m��j�>=��7���9ح�1��dS���g�?l�-ӟ�����GLO����lh���~�8����v=�.�P�HL��A��`�^����1�b�Ά�tB�p�q]����]��XM�"r<�n��_m�"�l�}��-{VZr�.z��*�]���{k<�''ط(».$$W��oD�q�}�i�鋕$�^.�/�I���X����r��Dk.������QBUM����J�@/��~5�g�S���e5�ЖR �yz����k���I�]eANkKcЀ26ģW�g?C!-5��j� wg�kY[�ѐh}�W�ɵ���-'���"�[�^S����+�l�c�b{��ca���b�I�CK�x!M�!�2�;1Zb\u�������Y�YO1��1��Ģ�@��/籹�f�y�@�7I�?6�=�}�%�7o;����ڶ��g�� R�F{��m��a^���Z�!����oP��'fv	"Ҽ�J,�+��qe�0ݰ������==�ս}�u����O2vu�'��A.P��M�FT�Ѿ�	�=�t�퍾�� z�f-��@�GO 1��c��6�qt��w�e}n��2#=�;���W��Ъo���d5���Ƴ�Y0��uMO�`u8,\>j��кܩ�����*��*o�kt)R�$O�,�V�׾Bz�SF<L���sԷ��G�i͍p��/<�͂�Y��zpm��d�����V!%%��8�QS4����b/�P
�y�6�n�n)q*t��Y��?�d�ǯ����x��$r�ӤǏH��y�Se\��u&Z�2ʖs�E�*�c�+қ�R�M�e�s�{��Y%�yQu�s�V�F�:���1\C��{Z���i�"��9��x��~g,9�Rw�=P���ѝ25�,n����m;
�Ts��)�~���@I�z\bS���14{)�KLw�i��}�?	 ]���R_��A�s��	�APax?R�`�3� L�K��\>
���F����C7-n�Kt�������.�I�+H�G	�C�m�#�����^�k(���6�7�h '���a(4�z��u�w�O����Z�ๅ4�$E��W��#���������,�� �J������������IĖ�pVD��Gƹ_EtW�����[Ԡ��h� ���.M�]�[,Ng�c��B�����\	 Ê����K!]Ah�pTy&l���۳�j��QJ������ %�VD�bH�]�D/'s��1\ɨ\\��������0�%��o�(?������[��}�(^����:�5�)�H�d�D��u%,��:��īg��~D��:�|i�i�fQ����ܡ�|�4�%������9���30u��p�Jj���U�:�sC˫��m�`� 4�hՐp�?�gi���a�:�>�V:]��A�N|߬Ϗ���yZ����ˈ�q:w��m��M�l��R��B��x~��-4�_KS��a.��K�/��x��˱c��A�!�9d��[�.2.8M�Z�������<o�Q�-u���`���O�ef� ͼ%�ʐ���#sVz����b#�U?[dd���j�3ё���;�|����3P+M>������Z��R�GI��),����Sf8��'';,
�9_���?��M��,.?����� =j3�6�%�쨿(Y��cu���lm��FU�w�KUF��!�>g�g������������z������]Z?��J�
w_���5�@�U�S���c�;�>�m����S�|�$��ɢ�-�����u㽨��aɊr�ۡ*8#?���e��ʱl������X�5�����O�,��Y���y�Û��ο��HeE(�X�4{T���è�ܡZ��SC���Y����J�hy�M�o�������(D��d^����I���ٺ'���zq�\����e;���A���M���$0��,o'��Z�y�Z�q#��Kvf�H�"o�3Q����%%�`?�/�ƕ�(�E�����h].{���� R,����=�/C[��2����8�1?]<=(�s�8�Q��9I�k�k��>Ӄ��W!
)U3�|�'��Va���7�pS|N_��-��5���׊�I*��Sf�?�C:3?.�k�O�������k�"K��^)��!��C�S�	�M�H� *����1W=�9a���o!$H�r�7�r�v�U�O�i���BH>��G�ҏ#�5C�H@�r
ø�a����#��^�E�7�D��F鞪A5s�=�w�Y%/��
B᤯�� �$���pm�&�YY��P0w�HC2��q�jȐ�\�3��}��rR���ÿ��H�ٲ�Ѳ_��ƌC'�B��Y��O)�-� 鲩�|��'�+�I��E ���Fv_?̸�]��"��
|������!|U��yh>�d(mf���&Ʃ�A�˹"�ڂ�ZK��}3�'�N��q���g[KTGы�N���υ�yɕI376��'�ƒG!u�B/��D�ˑ1-�@	[<wN��%&�t�Ё����?Ov0?2\H�a�\��n���󤜙$�,��ݨ���������m�&�5�Fb�;��Mb��kE�o��ΧFM��Y����W�a���Y�n{���N��
uE-9����D��}!gq�����9��%eoS���ZdVEYI]�; �:�0Yv�gv%i(C�7�{����Ql��{��,2[�GZ9V�,1��S���&�)═R�����Hg��I���f�X_lQGd���m�b�J��rN钽���T��}S�p�߲�Ƚ7ē23Ӎ��7	��p+�n�aRF����\凓�?��(!�沴���0��s���}T�~��덗a��{;&�ա�8�u�+��_��
֠�jl���m��W�����;�k)���+��p�����_Z8�K�2�g���NH�=u3��%�U݅��,��o��m�uE��J��q	��@�j��e��x��ty���n}9����!��]�UDj(6���(7)/���m2�L��d��	�g>�zg�-n��ة�G��P�w�7և�$�I������,��=��EP���L�n$��V��y��Q���=�o��*@Bi�<qX߶ vǦ��90<V@�:n��X>��/}��`�L�r��ή�#�])�{�L�bN	sƬ(��$xe�*��qb�i����p{�^i��bOI�� �ޤ`�Q�.���ॐ� Y>Bbݧ54UHD��yJ��ۆ9G5eSѲ	��fz�k�@ Ѽ2�z�k�ĕI��Aɳc���6����h!(Cm��S�w"&�Y+���}d�hX.W,ֵP!- �K��"�_�^nx&��+��c�˳�l����ZԤ�C��!hU�\i;��д�[F���뗴�O���10ԥ�c5@���/"1ۍ��ze�����μ36�y�������7;4o�u�˰��C�<�v����`�+9'�BѢ�"���4o��N'� [	=�8��t*�0p L[e�{NݫLX����R"0�c����۩���ݭu�:�<���>	�%��pdɸ�,�HC��b�z%䤩�q&G�P~�����Q^Ttu1��@�R�%�={$��OW8j��*���"[� ���
��繹M��j`p��\�ˋ,R��i!�����!��K'R���'_����y?��n�L-1	��y&�3��D���kU�/��-�d�����mEŋ����MC$%�X&8�y�4PҌ�%�kty�[��Iw�ndil*��Y������c8�����$�����ڏIK�`HeW�����Z�[����E(n�c��p������"�V!{��)Y@)�Q�'s���F*TB���1W����-��UBei�8���YCxq��gg*A��"�=K�.�lσ2���n�"H�\;�xs1�����;�+�Յ�SYI�1 k)h}	K'ֲ����F.	�ܧ���_O�!A�J�Ԅ��P<&?�����s8GG����#
BatF����oI�#�K�݃�R?y��2v���3+��	���j�#�s����β�-���v7Q�q2�(�\�(���G�u����J��b���=5��͟+��2K�#5���T��ج�{?�Q��3{�o�$%Ϋ�ЊBK�Z�WK�[�*�v-��<�5 ����M�%�Vng�����������+�e�/���\]�ArpO��lZsw�n�J��1����ӯ������b�6-��/�Jf�l�i��-"\$�<�����.��%��:�jX�?x��gIF�v�}Ѿ���"�X�5-DHH��%DAM׳0����o��B$�~��:��iڢ'�����;��X�4dV��	�tI@��#�u��q�)j٘8�#�BU_Ăs��d���>��� /V�0?���-�i��a7�ݡ�Vu�o=�cA�����ʗ�#ZyuD������w�ժ"�M��yﭲ-BS�~�^�-�BK.D���#���BV�����&�_c�AA��9�k�[��`.sH���@z�=�V�wo�D�Qڊ����`��Oq��?�%֐��TWU�J�V��u�#�[Jz��Oo��.b��%��;�8����sn3+��y�]¶��U����G7�)G�/�5�8���'vX߅�T�	��T��^��.Z�5�f@����a3 nە��¨��,�M�C��#`�F�=�2oކ�*��t�9$�gW]>�B���#F��-4���]�3�Ew�@b��`'�b����>����Pm9݀NjU|;���q��Ha����y��,prP�l�%V�?s�B����8jl;����$~�I�'5;����+Oy�$��m���A��>�"��}�ヌ�E��RX��TR)��c\�u����|a�[�
��8J)2y?Y��
��㞱��D[)k��wǯ�|�O����#g'@J�z,�C��#�e��W�JֻQ��C}�0�.u,q#�]�;y��8q� ��&�f���"
�HQwG�X��
��J���+j����=�c�[b])&���fRց����=6�v[��ܓ'?����J:�y�]�s_�Q��Ivgak�>J���})����u��a����X�p.��_��1�Ȥ�5��&��3s*���f�}��3�k,�lX~��n��o�Kiq6),J�!V�CԿHD�5��N�%4t�^d�W�IK9|0.��H�Ha��7Q���4���ĸ�B�)>�E\�M����C�EM��o���:���#{:y5��=>��������D��8�Iw�/A�b!�.�*�� �<���mb�s�T'"�����|��t����7D
�$�}�k��m��<|������JB�-���o���l�(�TM�O����mS���:|r�i��C����E�����u6_��~��6/�3������l8��`�Ug&h9��d���ӶP�*"�%�h˔����!Z�R�x��'#�R�,q���B�T�)7�*%_v͕D��7�����,ƭ�u-X��u	5�̑- w�@d <���+j��S9�%�����vk�&2��a��;�ɂ5��5 �?��,���|���؆����m����>byW��iMMݪ�k �^��Oo����);Ճ�aa�v Y-�i{�aNɜ
Ye9؃��x�/�8S_qf�z/��A�o������IET��疱M:[��v߻�%�@�C��[{�2ݩ:V�̘���<[L��9q$�1=S�?r&/<��0�m��/g�a>I�F���)�X:�GL�ԥn���ῥ�E��N��T���S��Ƶz�ȸ�K��o�3�vH���	U�9+����� ^�YW�WK)��a�?d��!��{�Q�0�$��}吝���������6_&1�9��W�P��+Ȋ�Sv]��I�]����r}�t������⨒�G���A*_�!���������w����1Ux���'�o����0�:�e����I��:��e4��x�L�t�,�)����XP��ҕ���ɮ��j�M��B7���#��gE�dI������ϵ�C-	�=��(G&��2��֢�@��E��yq�g�=�P�6iLS/���"R�� ��J^�P��\�B�qSK�[a{�a�!�T^�<�1���֧�z��x�}���1cFr<���<�]���{��+������(��b$ڹ����Iq1fi���K�^�D�M��I����9���4�I�@a�%��B�y� �B:�UCܿ�g5JN&��4(5��S�������V� ���h<�kOҮI��AD�c�P�6:j"��f!#q&� A~wݾ�YFF��0h3:*Wg�V��a�-�ϦŐ"h�~^�F|��+��(c!U�����Nn��N/C�7�!��N��d;�s�d���"������PO��1KE�Ę�3@��/]�Ѝ��t��?������6�Փ�s�����;o�A�z��7���';���79@�۹��2�}�[�W��sAo��'y�c	X]�@��qUi[yeUC$ݦ�<�Aҳ�KK�sD�ۄ~Ũ9u!m�7˄E�%����x��3���f�h�+9Vz����G�K�R;��lQ?t�������`Հ=-%��)W�$���y� ��{ ������"��M:``k�7\��+�F����2����m�����B�R1��"�a�4\ع��]L�h��Πh�n�a��#�f��/�ʍ�2�,��m�Ǳ��dtÈP;%[8���4����W���Ay�(��$��n���*�صY��U�y������e $h$���=��n���eR��Y��Za� ��SE��{c����?����1�CDj��{rz%Y[t^QkYgs�2�Fe�'+]1R�1!���ji�n8�/SxL�|g�n�ň�4=F���)2��<n.�����;�Zlsl2մE��6k�0��S�18,�)�cKU>3��ڳ�	���Pq}_
�eAB����;PP�?�[�i�B�R�>{)
��-F�����n���K�M*������y��q�+��	��c��#}��l��D��!�wM7�'Mw���i�(��z�͸uR8\�E����J�V�yP?��2|�!�#p�J�.�����d�p%�	�O��\����G��n��n6�US�W�i���񑦝���' ���+]�MC�D�Q�gD�(��W��qХR���@n�����]w;�pJ�tl�?�)?/��Ϡ�z)�ӊ�̞ib~���/�A9�'כ��g�\�lrا#��i��%<z�e(?�3��"� Α�.}���{w�ӓ�15�~�H�`(D��+���������V���~���:'.�i��i"3�A�ѡ3S�4��°�7��2>�<4�u��jq�j��.�>��U�m7s�Ԯ�1��!8� *ER����Ǹi j[a���%�V��Vؾ*A��g�b��cH�y� ������w����Et�M�V���mB��~��-*�2K	��8�������0�c�I�A&�9ZA�[[�.�,w��Su����Z�o�
�Q�4��`�#�OS��V�)%�v�ǯ�����V�0�O�#\�d[��<��lL�)�̀��;a�"L-
*3�� ��Q:�P�K��FG��])b���6�8�+�'��h�o���^zY��].u�������)3;Ş�[�,餇�C���>t)��U���V����UY�4igg����ׄ��(z�_��Zg]�H��@��w�ʫ��B��I��r;��mԙ߀Iݧ|����,���c6���\��s���ׯ�r��֡ ��?����:�D�S*Ql�}K�W�ׄT�5������O�ݜ�E��������[��%�EU�<X弢T�|����*S�I��6Kǎ���J�<4yޠ=LFτ-J�؉	D����� ��+��V�Ѝo'���z�o���e1�*��(���&�~t0�c�,������y��)q[��jFf��"�9�Qw��{����e;N�����7�xx�"3]$���i��R��Y���=��v[rr֓b��n<5i���s�Q	�I��kԌ�>I0l��\�)���2��0�Ma��w�-�Gp	�6_����c�5��j�@�<*CЭf��^9}#3��k@(��܏��e`�!FdK$�)G#�!��C�K����~=" �N��e�W�v�9��&�e��H<�#7�Ѐ���$���}��>����Ȕ���C&cn��s�����XI#6}��ϔ��i�>���wt��3�wH></�`�<,D���� wtm"m�;��On�k�ھ����^�`��'Qc�}Qq6�h�ٌ�T�O��襼Ѩ���|�|���x��O��Oߦ{n�*�� |�����|���EV`l���2_���0{�d؝ ʻ�P�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4Hy^�gАPi�1E�{�p%��������Y�]㾗�1���~uµS�	"&���P,t�������]��x"]��/]$
.i��7�7+����O��������qD�}ei�%7��<��w�g/���'�Ҭ}9D`���kS"�D�2�E��7S����o1V��W�)bu4r�\���qt��$.�
밶�������i��}hpv�p=��H���V�l�M<4_�N�D�/^�+S�����S�ھ'%L����ʠ�y4�������e�X&`�^fI�덜�j�*�@�:�X����
1��x��d� ��-v��cbx\@�EGrU��y͑���� ���%�rv���
��Z^K�;yͬǒI������1�ާ���(�[*Z�E���Y�lx��쓿��7�ա����4���03��l_8���<�[\{c�'��[� �BH�Oˋl��ZO~�.fcMk$�U�w�m:��^�jy����1Pa����l�0�}��w�^�H�T���O"j�t2����2V��hͥ���jR\^w��vЀg�- MA�2���D���Lx��$�[��	�ǳ%�����f�+��Y���2���V1c�4%X��.1l�I}�Gi��Y�g���+�#��4m�3:�4�׬�m@s�-���B7�k@F����`�3&�����B<4D��1]�:N��@$Z�e������1Xk����@{��h���Ҽ��߲k��t���K��h�q/�1I�gAe�Ô�K����[%1f���W� �I9z�Hx'��Q;,�l���g��Y�&@e]�NE3i����� ��<+��W��ě��0��cVNQON3~�`���������I5�E��+ ����1b_u��!���c�cq����:�|{�>�`M�S����u��e:��G��^F���O�Ɯ�y>ͧ)gp�V����a"\Ӕ}!��Oj��T����.M��h)Ol[�S�\-'�+��p��������I�)�on�g���z]|H�+�>���=�>���m�u�ݞe�P��o9��\��UI�n����W��6Pz��5x�������jpkhK`6~݂yp��x�q	?�����-8���j����V�|^Zw�z��R�卺��c�G��L0	� Hx�w��FR1K�t(fi�#Vy<\5
�Y��c��[K���cG�}��kk�l!*h�Ho�]0��OwM�x�"xӄk�J�:����so|���E}�"���x2C��s�
t
i[-���ĳ`<mE�?@
��@y�l��c�f���S#�7����SkQ�6��,B`Mj\k�`$t�FqT��HK[��ښ����,LY����^�� ����J���� *�>C�8�ZJFo��J~�ԇ�U���5k��Xe���?�C����o�v�X���%LP�z�ϭ��Jw���׿-�r}��ё73:Ppѭ���r�x��A~fo��q���-4:?U�)Z�L��Y�HQ���赶���Ҍz#�'gK� .a�W�"��۔�_}9	�!&��w\J�lOӠ�aV2��%ڴ36E�b�T;���<^�)�>��v� v`��CH[�����;�c�G����8Ls�n�V���H���m�m���98�Ģz�0��*Y����`T�����:���ңup{2��T��DP��	S�v�p/sz���?���wAk1�9��ɤ.�� `��J�B�������0mՉ�V��m�k�3���x�+��n臘�iQ���VRS�;�rh�{��	d��j�Q$1���(vO���d���/}�m��|��0w��I��B�)��N:�
^���SK}X*�Bk��O/F�N��W���H�
f�/o*K ��﻽�`d�cG��6<W���\����_�Y-�1��'��50drlb	�W��^vyգ�Y�t��1? v:~ �kւ���'[���rI��*p� �;��%����=i�<�]�v�Y��r��&��)��=λ�9��	�r�r���S��s�%��7��Z@�3����z�@�4r�;S�������# S��_���;�.��$7�-B�]Pꤌ�oh�ZE���	��qFq^p��=�#&e%n��.;�����lSUkd���W��s���t�hg&���Ev8n*W�L �A !T+	s�Z�"���2ۄ�b�M��y��^��_�֥R��f�q���tz���%�Mc[}�$!.�X_�'�p��^��Lc�?�)�쮍����4<�UH)'lɏ,�S�y��q���&}����#4O��:���{d���i���y�����qFF �S(sR4N�������,j�s�ߠKˆ�%	��Tm�4 �B.R`�S�-)�`촇����[�&���o���z<�8�1r�B���#�����z*9�Մ��󞏸�S���Bh�קsB�TD���4t��!K�ğ��uה*[���� [�ui���**�ל���A�N�.�HD�9C�˕�W-��i�<�!$�;����M�o( ����&r֢)��ZV�����jX���;�}�!-�f���R�r�~/�*}��l��%䈓�ŝ���
~'�e��v�������MB�2��n@n,�>ȇ?-��(���
��G�b�f�C��l�O秞ď��,��I�0b�b���l�te1�z2ټ�������&�����R�z@�{P�;!6J����΂a���N��:-�he�ow�ll�R�%Φ�[�CU�͓sc�3�d3	K�������(]&G��gp��8�eSc����sV���t�>�=d@~Ω1p�Z����
^a]!��Ds��8=����"
v���!֘ౢ�e$/�c��*��{츑$���E~��`w�f��i��U��8���q����$9 ��`d�����N~����rW���Q6鶁�k�~BJ���͋�ib�~�&�cO[̐����2Q� �My��s�P�0��sJ�2��ɉ���V��E��R�j����c�Q2]	�<4Xj�Ww�Y v�e�\F� �n2ȿ���D`�g�Ζ܌�E��� 	[F�<
�(g� �Y\��9��P�V1e.,g!x��"���GkݨY�𞛜�+kVª6��3G%�4+��/��/�N�����8�@pC��͹3h�q�����D��!��.Nc�@��e�J�9�1ڂ��[�{������>���t���v�O��"h-늚���i#����K!l\��'D��"@_삡?9<��x)Ԯ��_���W��#}����h�e��N!��Ӟ��b��Y�ڷV����0��&GN�R3��`�Q���_^�I7��9�� p����=Y�3��u�x��U�}�%�g�ݕV:�w��JTɳ��G5u'�	:;9G��&F�,uO/�������gr,6�����s\��}#�pO�ƹT9�꡿F��)�|C�k�\�UT�l���*��}Zf�r��;
)H(}nP���~2ъ�T|��F�����U^pY��׭wj;=���
!�D�J���΋������Y��
 5�<��+����xf��E��� ��[3���� ��%6�גV΍�m�Z�EA;�Wr�v��SM��!鞻���j��(���Z ꭿ�clB���Kb�����+lȧ�h���&���8��U��(�B��7��UY�<F���%ԣ��D{o�3�*���[S�S���{[M��\ې�`#)�d�E _��?�_sh{�	|9m[�?��?4��b�lؒD5!�v*�Wh���⠼���Y�)i�ێd�6��5$%��&`�"+PP������=�D''�$����s8m��:=���S@�)Ca�n��#���P��hr|���B��hH��S�v��Pe�鄆+.%���&_�:d��&K���^v3 K[�����^��ȗ�Sgq��O�חtH������ ���V�F=��~���9b9Z6��uw*U<GbϝA"�bx��o��nTM�w4��>�*���]]<�5����+���z��6�wB�
|��R��u�b�Q���H᪄c�2)�
{�����i��y|?QZ������#�o0� C�+p�,X�t�vZ;�U��i�E�z8��T�+	��1_`}�k2<�����F_��8a�F]�Z�R�
)�ڒ�9s����Xʲ�f�g���MZ�-z`�-Ȓ�`�����R7�C��������+��䪰�1c�dp/Mx�XXzR�c�B��c~� �]�>F�h�Q�h������l��5&�
M�)�)8�>�BF*r�+v�X��ow��ޠ2�Ai�y��[� .h�^4��t,m/��!n��p��Ň4�2��r��;F���۷�gm�h�2]�K?_�>���G�M��{\��c�_�!�8����TT�w�u�ΕG�{L1+י�����O!&��H�T�����fg�*g�� ݮ�dW�]L!U�f�{n��!r�2��R�������Ma�Nz�45��2�F�����V���\�>��Mj���ZՖu�T���=-����F���+b	ڀCx��9�^�w�5�Ƌ�����q�0�jsb�2��t����\��=��W�N��'��z��@ ��cNNJ�w ���Za���N�^u-���Ow=9�zV��΂[���7�c�\Yd[W��c�S�(B�G���p��iⱱc=e��ix���Kt_;=�e}~�s2p�i���2?�8a����l�l�� =�;���[?ƣ��B�����4p�/��l�Rt�{��$�[E�4V�@H��Hi��$��P/�����$aOɈP(�����\~�Aߚj���6!�Ói�Brp����Ȓ��~�)�cwì��X�E��HKyF4��.4�Pf���Z�H��8��T�>��7�jAɋ8�2@p�)�ĥd�j�z�w� �v��,�W� ���2𺔗�u$D�[y�����D���1V�d��P
��(-Y.i��뽌xަ1�
{����بh�3�SG���Y�6���+����^|_3o.%48Y��W�i�W?���P��:�@0����K3������Ņ,=@D#����JN�W�@�Ae�r�a |1v��G{ٔ�"�{�f��ߜ�ޞc���GhUP��}��s,�-�KIf��U�Ohn�J�f�o<9d��xQ���|�q���
������1e��N/\n��>B�����`�G;���X�/�N!+N;º3�f`
b>�w����eI_� �a�` ��i���e�[��unq}���`�d�Jd0��S#tb[����gEv�l��b��@|�;5zA����t�	�,��W�ѣ��IDY/f*�AE����Q]�9�e��Sˏ�����\ﳒT��D�F��(b�Bɉ���J&�b�m��,�,����6��(�i\M�����3oP��{4c�R���&���T�Ǟp��|���>�P�u��Ѫ��b����83��������N���Nԫ�"!�.?`,Ӛ��^�jK�?��Z^�"n|z*Mp��6����>F��*���{<���1:2���O��L6)tSVzHG�g��i�)�1>����&����Mޤ�n|�]|0\���W�i�L9�"?�e������\��tXg]'�}" 2/6)8.b$�7���,��܌�O}����[��H� D���ebM7Ȃ<�8��uyȌ|�a4��eLD9A��d�[�]���~xc����������V��㋉/bn���u�>�o��ȴ��CF�O��ϫ���`4{�b���@Yp��y=��v��'�š>��o��v�KY
���{��O��R�[\3u)��4� ��3�=�[�V�C�d�� �IRX�L�e��dx�G�Z���ޑ�>֟1äh����|0]ъy>#�:��'�]PQ)\T>������7Mg?��yE���T�KKE�8^S�a�T|�o ���#���f�72`�K�?�S�����j��d�c-7��n��2`�������,Q��#��v��eA-�����,����0���V�>���&�C�*�v�� k��y�R�5��ao|Y��Ę�q��˓��XN��]vv�ph��J�n�΍�g�O�zB{&��۳z�27ԓ�X��R	}nêIS4`w��)������i��Ȼ��@���G���<7?ֱ{.�i)���NZ[��,e�"�0ƭ�����Z��g���f��!o��-���"����Զ4��W�־|��o�G�qoT@�t�u���� N�II�U
U�|�=!���ZI�I����7 �;I ?��,������#r�$�M5��w
���Q��QV0�=��oOV#��K�꡺u��4p����a3>���0u�U2�D�7!C����G�k�g��:��f����$׈�^�*���	�Y ڽ>C�RP�)���V��_0N�g3��Z`l�{^7h�iIEI����ú� :p��ٝ�}-jun���N�/	T�'��:}7E���a�w�Sru�-�:�@�G��tF��zO����š�Q�g��F�?鳭�\�D>}m5O6Z!T�D����cR})���bž\���a�c���G���|�<�D�)�Zn���{`z���uw��p���T��9h��g�1��tN�i4��>E9���9D�Ƃ���8���L��ݎߒFm7ÎV`P=�M���Z��U�w|�����/ ��cV�:�;��h%�7�8f���S�Q� ����(� �8�紽iW}����|���*�+yB�4��9C
 ���㲛}z�=BͲ�O�2�Naa_WƳ!�s�`
/�om;�4o���dR���y�W� T\9�Щ����;T1�^��\�@d]	�\c����ܭ���?V?813�kv�$��ޢ�̓t�#���G�wfr�r���"p���|┹�92▐v�k]�Z���c��&���=�<�[^�	7��rS�\S���G~��G���Sg��ǿ$�@��rC��״�؄�7�#���X)��\���ď+����P�뙑�#Z�æ̫��q(�^�m�=D�B&�w��`t���+�΅�kf��9�[s���t���&k�u�9,8��yW��"��Q!6@zs����ݝ�����M�Z���/�4l�%9q-��~�ԝBM���2���=:�p'�%f��93����?�c{����TR�4!�DU*��'���,V��yw ���#��v�aTO4�We���5�����P�ﶽ^��aFq�����UR��ϔ�y7��uDs��ˠmG��	��`����-�d�`��-�{���˵�"��Շ�����fz^��ٓ7BJ��#u��2�z��_�w���F��X���B
jX�U^Tf9��:������������m�z�� =�i�*��<�*�A���."���m+�W�qi/ܮ�nZ;Uen�b�C���D�����$��*���{'�9gP�$�.�C&
������P�T�5��Z^k�P�nu��(�sAj����󋅶wP���V%�����Ҝ��k]�x�go��؇NH{�kx�[IZo��0%�\R�f��2��I�Q��d��	(�&,2(��U� �f��u�y@^��%�ש���[)6M�$�"�s�>�����T^��C���pxm��𴸹4)Y�(X�W��0Pb����j�W�:���pƽ����݉��J!R���j9�<�$��RJ��W�VG$�_m�x������:w�Í$�`�kQl���屢_��+dI���ѦX�mU�9g)$�0��li���}�7tݝ��Ɣ�'y�9.�~���dz��K��*~��KƘ9����sإ&���ύ ����'�����x eM��$`����.��� ��tE�;���ҋg�{z���[����;�;˕�Y�+O6��Z�H��z��ߎ�ƒ�+����������S�`��Xs%��X.���4�5b�!��0��yN�fyAdEEb.��������6�Z�s��瓞{!7G|3x6.��0E
H@Cy_vt�x^�)l�{
O� ]�,�X_����U%  ���,�/��o���zy��B�w�x�V�UH�CVI�'u��&���/��R��h����G��<���� F,<N,�]��/�F4�i���o�^��	r,�ʕ<h���r��*�x��y�{�'���+		��N-Y`�2�1Z���D6��8�O�{EL�P��˃��#�`�>�sHhBO5ԩ����(���T7�������8��#�J���+'q�%��T�L��D���'=xJ#Y����\�R��r�0�Ťv�V�|�,j�ր(�mqT2�4ȤJ�I�;6L09����_Y�zq����o��C²k�p�WK��)L0�p�Rf�㵍Z�jr/��5X�ݾ����K}�-�)6۝�!\.�%��fgdiXmh�}����\�I*�貮�ؓgL�%sP-�ڻ���]��x��ҙa�1����n��@�!cUq=Ij-�ͻ���`�xQ�`^�M��<����'��*K�ݑv}���f"i�QH�٣�"[ث��*]r\�=������f�Z�K�x�I���U���-Va�F$�ސ�8�	�g
��͍U!G��3�<=���ATR0�����l�ި��:�� ����<Q(��d����[ا�N����z��8@iZ���}B�=�v	YP�#F��a%Z��o�>o����DJ�S9��ɴ[?t�\Y���b��� QҰ?��@h~25	.��[<���N�l��5Iv\�th3��؎��0Y'��M��臩5���۽;~?�~��"�� 'Iw��Ɇ�sj45��=ZC��% :ha~�5��`��D7��A(��[���Ү���$vNv�`���g�vӎ.W�a���[:�G���A1v�ڄ[W���=���m�Ŧ�qbܙ��� H6
�Բ�;�H��>U�3t��W�b+t�����*���ϝ3��b��oR$�n��w
f��/*<P�AP<����Ȅ�B��F��w4>�|�a��������Q�K'z&��li)�d�
B��q��L�??��AQL���%#h����.�+b/t,�x�� }�{�[�@"a8}�[���+���c�}5d$<K�&���F�	w8Ӳ�]=j��D�)D�6���sya\���\�����z�X�M`��������D�C?���bc��,��8�ܘz1�ړp�	��Jl�z�R��,�ͼ~�|A]���F���)����(��/9��O%
�E�_��p��F�+(�JX��ow�ݠ��hA႓�{
2LR���a�S�m�ɮSU��vg�9�N2����k��� �i�*m��2���?�>_��G�Rȭ����[_���*��y���m}�i-�iB���ɣ�x�
����~�pm�5�#�
��6lZ�N�`B���pP��l��~��cq��IW�rU��*Wya�D˩*	P��&����uR��Zw�ck��8��7�j����f�2{�f��N�_xWjW�>w�2�v[}��� ���2+R����iD��n�Q2��ɢ֭�X���I�?�ы�=liY)�a7���3&1�Ix
�G����n��G.�FY�N��+N�<�y�K3ꛖ4vr撯����z���M7@���5�3mO�tk5�g �D��>�?�N�!@ɨe�m��#�1�s1��6{t*�Q��P��W�X޹N��0L�h0/ҚV�C�,t��( "K����hT1j>d�ł�8 9�o�x�7���[�q/����3�����5e�fNjK������?�A�]��[�֧���ȡ�)@�Nv�v3C�F`�����B5�Iz:	�� \ sy��2�)��h�u�ܶ��z���� ��:�����-Xr4���uJa�:��GF��O�������-g5��>���fX�\x��}fW�OO��T<��"����Ȍ)�
����\��hl��|T̀6L��,�o$�)k)�nӳ���T!z���-w���ƶ�fɛ����c�瑲

+7�.�$��ᦖUn�1���ݼEH;ZY��5�����J�w�j���K%����k	��E/�)ޮR ��P8=ʅj��jϭ�|���������@��Cf�H5Z�b;�	ΆH=e֑!3yR6�����iU�V^�5�Cw��5������Z���c�R��ބ7k�F�l����N�4}M0J�O|`�xA��S�_kϜ��ν2g|�I�E���_x�X����j
Y�i��b�(��%��E���
�R�YG>e-b��6��x��7�W,�p}�;\�,�	�M�����$�Wqy����(��t��q�,� E��ᾯE۝й�����oT��Yg>H�J˫�mJ����/���;p���k�����)���5��y��P����YX��%51�?�ǭwq��O���f<FH�rbw��8�:,aI��}�r�er����~��q�V�
�:d�;�LI��MA��F�������m��{�L"�N@�aLp<"��Ҕ8%Y9N)v&qy�{��!LO���a���*4o3�����;�ʙ<���cVw��Z ۢp���H M+��I�;��q��+���˵L8�}E^VR/Hf	Em2����w9��Т�Ńvo`d~�eMC�| s�Mﷺ�p�nC�����-l��
�S�=/���=���k��uCrA�؀����	��%� ��d������>�mZ�V��b�0r��`/D}xz��4RC�򾃤)�Vw��;e�}hhU ��ր���qQ`F�����(����ܴ���}��\�$~��չ�ՎQ�Bũ��ӶC
������}��Bp	WO�]�N��?W��ؖy�
�#�o��h9VM���mdUP��TW�+\\���ClZ��17����Wd.~	N<�C5��(���~u9*!1v�qv?T��X�0(�|Ti�@����O�U�B�e�^��Y��D��%��A�]'�Jy��׉d&�!����=[#���j	Z-7r���S�6[�~�ꬕ��p�xX��ʍ6@�rƛPחq\��ʰ#%�?���%׿�L�Ĳ@�g}�P������ZJ��̮r|q�%^U�-=g|c&�/���}י����qg@k	|���su+�t�&�N!��C8��zW��M��o�!�ɬs�sq��K���g����M-:��ܓ��:������kqP�]ڙ��SKM�A��������'|����q��?�L��	����G4$%U�&�'Qo{,y��y��޸��)�@��K4��� ���6v�沎������FRp���@Ry�����aܜ���Qǩs�۠��*��轻�]�!�'`&�Y-N�Z�y~$��s��+O��ë6D�z!�Zٶ�*B��U#X��u��z/*^�z��1:�����2׬B�4s�8#�T����9�蜳ҽ	[�Z3���������  li_�*/?N�-�AA�~m.ȁ�4�����W�viV��&��;X_ֺ�C��D�1>�$�/���#��e'%r�P�[���C��~ӕ	g	T��(�^�P�u`M���A��Ϫpţ�h�$�T���C-���5���.Cx�����1����a�[�kD��%�b���8*�U�iIq�e� ��L�j��0��u��@&�)~�u��^L6ӿ�\B�+k��-ߣ'	�"�b�yx���^h0�Cw��p�ҏ�ۉ��s�Y6H�Ɔ0s�W�4��:��E�`������`J�p<��a@��"��o�� �J4űW��V��8_0$���yw�B�$$���>l"�֍R޺_�Bdlt~�T(�P�9����i0lli络L�B8�"���`BX\�h�ͱ^����G'j���G�����c��9ӸM� �j�� n�����brx��E]n_l��'��c ��%�lo�"##��[�Zt�~;�g�B�s���ߟ�ە�.ǧ6�(��Z̭ܻS�p��C��B����)&�{�_� Į�͟���5SU,�������HG���(+<y��d�z��}/�UO�V=�!'<�&'ǆ/G�5�x���2G�q��"�}�簮<�Z]���/��'4-��/���v�	ymZ�|y�</ ���Gα��Qw5�����	�N���Z�NG�AH�`�����9{l@l�Wt�ǲ�~�Fp/��%�hr-�5��Ƚ!}��;~��Լ4v�Ă�i!�p�J"�(+N	F�,�2��L��P��bǗ����Jj_ݯ���\�}�Y�������K���!���>�b3�(&t�q&�2�`i����I���6�&���m�ݯ�_��q����V��C�2�XRKK�sL����q�����cE/ݲgX�44�k)�K�SА�ŝ�I\@��%�'�fNu�X4��}¹��m1I��ɲ�rߓ�.�%zw���î�ZbM��o�Y�5�|���%ۡߜ��_Oc<�%�-h"����j�Q�$�6�3�Cj}��3�z���5Ȟd�}^3�fi�)�x�j٪5�	H靖o�*5�����=��fp�K��rx�̒�w9b���a@�y�e?�8�}b����\�}�Ѓ=�u�~r@R����'9{��>?�7�CR,¯_.n^�ĩg�����Q�Q'w��,À�ˎm�t�E���V^g��Tl���z����A��	�%PtuX�'ăfo��0��dh"/��wA ���+�F�qݒ`��WT���k��GB�OQ���(��Ʉ:�7���m-�:,Aj���%6�I�(C�=M�~��pzk�P��`:c_ێ�d����E�9����`�,LPP�.b��z��5;��h3Q[�ܲ�����)��f�!��i`����L�j�C��l+W��4n�ݙM+mK6�8����~���;|{����,�z�5���2}6DO�
(H��g��V�Ă198��x�o��^�hZ��{�]WȞ%gԐ��G~"�m��D�v��+�]xl"Q��/ѥ4.]4?7>����
�����O���]�����uD2��e]�z7#�<������3�] <$ҠODԓ[}�;
�I`:���}e��cަ)����1��Qv���^�u��G�Y׻E�œ�+�2n��a�31��4:�m�N���n����$@r��A�3R참��ƅnmgD����
�N���@PA+e[ȋ�#��1��řx{[/��E�h+��޾�� o��wy�hWe�]'1�pN���KK�������^�e�E�9�!�x�*��}�b�x��A�����Q�R�Je	MNq��}���Lf��Q�DPI=-���P��N}�O3*�;`��r�BC����I�6#�4 �+��9�I��@�u΂ֶ9�����͇O�:�f����y��{�u�:C,G�sF5�`OU�%�8Pg�O�4\��.}͸O�I�Tc�6�),��ÅS){d���P�\9�hD�����ͧ����kV��)2Z�nz���#�Sz	Dt���~��Е��GHșk�8�z�@�����e����Uu*/�M�݃$���?�5$ʕ�5A�1j�=K��ݮ!%������l�����*�8d4mj8?ϔ�|�n�@�~�S�9oԷ�͍���?	�H$쩑薽R��xĠc�i�4�V��5�$��}�,=��7�|��cs[D�E�Ek=��l͑��B'�0�[�O#��x�5Y�K�k:����\� =�|���E��H���bx^��0�4
��im��/40�?E�oM
H���s2����x���;���7}�u���˨,nn�M���2�$ �Kq���������z�g��,x�р���>��4�^�_�V���L��>��r�2��J�8�v(�3��Ǒ�k�'��E��}���o@��N�~�7�X5pi%<�]�&��>d@��HU���)�^r�u��=�K:3�}�9��rr��p&~Hj��p�1�:k~�ը�L�����]���b�k���&�M�S��5[a�@"bGf���Z9�_�&�|z#�?�O�}a�.b��[�3b�q�]'; %�<
&�j^�ˈ� ���H��H� }�Rn%;ɯ���͍��3L'DB�V���H�S9m�.\�"(�9� #��CY�]�'8��������G�� p������g���SwA����ǖ�"�����A�<������F>��}�v�*�Y�x��KZm��V�s#�N��'�$���U���ܣ9#L�P��V~H!;L�Bh/�_���Ű\Q�4��D�(";���'��R�}��6��]�\�O���9B�6���
�w���s}��B�O[ɨN+�7W�ؽ�
��^o֩6 һi?�d�R��KzW���\�ü�JZ�x�1��a�۝d�Ǆ	n��L��O����"� �1=K=v��3���i���&x��!�<MX�,(�,U�!�����<�����].��`hO垚&^Kn<.c=�R��eѱ	��ar�HrSn���Qfg���L�"f������]@,�r����~������#̔̋Tm��B ��T��S�n�P�w����YZ� ��5�?q�*^�H=���&��Ї����:�muk�6��݅s��t-x&�����8�**WGR�m�e! L&sC��|�	����M�T�`PU���*���}/�qw�nڠW!���TM�3|�Zx�X�'�~��
���x��?��(������4�;�U�T'�C,�"y�*��B����«�44=����^!�b�<z���z�F���F�����8R����%f}�Ç2�X��sm?��wS�і�D�}���8�n�`M�u-U���`�I���T����J�D�zh ����B�C�#?��<�z֞�����tk��-�YG�B����9 Tp������:�B�p���͔֢g�$" y�i&�A*�!�����AK�$.�[m���>PW�z`iM���M�;�-m�,��C��vD�FT�+�ۭ��5U'��qP�B����C0���;�#�8cT�@�^� !Pz�pu��~�Z A�p��w���O�cZZ���}���U�u��x�H���uz�u>�[���::_%]�N�!V�|�Ix�,��A�>O�p]?��V�3�p��u�?�^Sc���*����\P���a<"�k>�H�@U,^ot�C^_)p�q�6v��Cc�Y�(Y�a��0�|��;6��!�ꅔ<�,��$�S�J+���.��4H��"W���fJ��=W���Vx�_w���E�Xw��Q$�Uõ�l��P��#k_�d��U�[���7��9q�k�z��l�f�d���A���.���'���98(�~B���:�m:6^'S-�"/�~paد�U�Q� k�`��#|,�h��eׁ>$*�����.�ΐ )�EPa��������zy�[��u��f`���e���߾��P��:H�}�z����X?��P�+H?OԈN��|��]���m#�6WX�ೡ>&b�J�Ժ hy�df�^�EV�.Z����|P�탋�^�s�YF�a�{+�I|}��.Fg��@Mu�_[�v��+)6��{@` ��`��:���U/�ۖ��T��?������-y׹a�o� �ZURS��'��M&J	v/�X�����a$G���%��J��<�L]�/'�4z.�r���(�	|�L��<�<�O�<�D�49��44����^�	��Nw(�ۼ]�Z�����G��C�4�ټ�{�c�Z}���%�	ƻ�*�<��hUP�5^���/�$����Z��%�5�z�m�1Je�@+�c`�/Y��*ܛ�ևݎW�_eq�J�y�Y��\������x��n���`m��vv��k�(ɴ!q)t.2:V����IфF6VE����� {J_#<�q�7����CL��:��K�r�Lz)�����(#�^N/@�X��g���oK����s@��Iu�\��u%�u
f��aX�p�}��c��It��8�Y�1;�%}��$�o�P&�B(f��V�_�4�h����(� Sc����%�-�;7�	$JM�QIr-�ُQ�F�Y�7���ʱ����"s}ATMf�����٭Ϙl"��K��*'4��Gߚ� %�fP@K`��xŹ����w�h�Fac2(���Y8��6yī��_���3į�����WDR:r��ꍹ|q������:1#R���_Ս~^��g�_�>d���,�f����tf�v�"Vg#�El����\���Y6`A�'=?�t8�eJ�q �o��Χ/�ivA#o�?�p��`��n�#��Iu����� �����_�{��u,����v��m���%L�:;����W:S���uo�J:a��G�-FӪVOw+�C�O�Vzg���c�5�+�\\ݸ�}k1�O��!T��T�H��aX)��1��Gx\��{<�!���H���!�-])�c.n�2���z� ��;����>��[���e�V&�o��3b`���&u�US@�$���)A �n�r5�:��d�K_�8jz,&K���������{?��Wh���>8��j�Iu�2�|�o�^A]�\����[V��MM��h�	���H��l�F�R�;-�~2 iZ��V�5��4�Ƨ<����4�֚.RcQ(^���k�	�l뙙rN��y�05�OA��x� iXr�kt4�� J��FT|<�RE�����x<X�μ�
�|�i%�4�<����E�'
f'�:�L_
o��0�}�]�^7s0���� m,L3>M��W��$>��q^�(��}��#Vd��w�,V��'F�T1ѝR0m��`�������>��J1J�`��Ԙ��Q����kY#f���%}�M����E ӕz4XS*�%����p��Qa���˛;Kr�r�[�[�M:	��L��	r��!�*~�^Y��Z[O�:IxݟsބLC���7��8� �އ0�ߌD%��1���NgaqO'"����ax9S�|&c�A����Oyva�q���3@�ϲ��;;~��<(��HR��i��  ,�f�He�8��|W;'�r�4����)L�E��#V��fH�qm7��ڀ��9m���3��� ���4�*��ᰂ愡N�\��p�` ���W<�N���S���zC��V�y~C����Au(瀃B�.�Y��D��TY����͎G&Pm���V�]���s-ɅaB����/9����{-�nK�V\0�;��h��ч�B����Qe��(d(@�������%�L}�������:3�Փ��Bjɡ�`
h[U�K%	}�EYB5_zO9l�N�ǏW.�^��)D
p��otǈ^�g��<�d��օ�ǽW3<�\��(:��S�1\����0d|f^	�#��\�mLU�c ��i}1�Vv����5��!�%P���£ڤЊfo�J���I�)������v]��}@��c&&|@�ǎ=``��'	�&�r� [S��寭媯��� �Ѷ}q��o�K@J�r�Қ���Od#�d�i��s �\[Z��#�L�(P4Ƿ��ӆZ�i�)�q��(^��=���&o���6�`� ٫�6Zkn��ꡉ_s�&tK�&�į;��8�i~We}��KP�!���s{�썔��q�F��MR׎~���i`$��ʨ�D�q���~#��<��M�n��8��>`'!9>�(��Vv�?5���8�����X4��GU��H'�{�,�W�y�u�4���ɰ�4Agل�G�{�Z�>����ȒCF���]��R~�ۃ�w��Gs�6�s��Ն���5��"1�b�\�̞`k�-3�L���W�J"���s�(�I�z�0���gB�!#��I��)�z�����+�6��B�tw�Brg\����T�0����%4�%���=��Z1���" ���i��`*�����N�A�}�.ma�yc�����Wwp�i{�f��">;��Ⱥ�RSC]ғD�z�	O�K�3#]k'��LPj���C}C�-Q�Y<o���T'�0M�^�q�PX#�ue�j�o~�A� ԪUa.����}�⾑����+�:���P�x5����E�b����8[�����%�j��xA����-IV����f��q]���h/z�G��}>��[�u��^1a�?���P�)nZT��Υ"�tի�+Z�^��^M ���U��Z�H@�=4.!Km��2����c�!�������n8hJj��Ϙ=�|�D����#�=y�����w�	��jH(X2�l�SR�M��$��i��V)��5�z6<���\c�h�ր�?c����I0Lk�_�lѴ��~�O0[�O'��xL����k�Pr������|�m�E-H톸��x�x��4�
$_+iҳ?���VE@lT
LQ�)�����0�Z��@7��:�H_���,��WM;\}$$"�q������IgR�k��,���фn۾ze�8�q��6��Zd4��f�>�q˶�kJ��Q���]�7O�K�Mk����R8��g���}��R�ӻ:�X9��%����*i+�´n���M�q`.���r-h�AB�:��S�$ҭ�+Brv ��5F~���!��5��:�e��ـ{Li±���_�Q�2�f��V�9�*|d��'�9�ta��"f�2�C��9�]T&<;�'w��B�(O�'Aa����̻3����;�'<y���E�Ϭ� &m�L�~H�1�V�t;M�>���K�L# �*(V��5Hqmm�x�ڦ��9�ۄ�*��a���d��W�_���$J��dp�U
�J����N�#��V܈PoKD5Y��T���N��M����ݷb�o8�*lj<�����|�Y�xf�Ķ[��q/q�ǔ¼��	U	�H\�� :�R�b�ش�i��V�q�5������ đ��oִGZc�di�}�ku�[l���'�S~[0o�O[%5x ���3�kN)����Xڂ|��SE�Z����x���hx
ثYi?��g�z�D�E��
���ݤ�����W�J1[ҷ��7�e�B2�n�,�W�MN�g1J�$X�q����,j���������,��KѸл�.��l��;�>��"��I�>'�g�j�(J*�Ӯ���k0���[k�͘��3����Qǁ���o�!Xm�S%t���^���v��.���%���	�r�l��u�4:k���\��qj\r��T��~J��siw�:�����-Lu��,�M��ᵚ6!�
�s�^��ً"m�aK+�"��`����9�w�&�[�t����O�;a�)�	��3��[�F-F;X��<B�)����� �{c��HH�a8��L;?�+|���'�LW��|��V�[H%m�m�n��Zo9/���8����_[)�D$M�;ӷ�(�6 p�������o����S�����Ww(�S�b��`�AϡH�������x����\��B�!�!m���V"���O��_��\�^�9N���w�qJK����V��;�1chg����i��FǙQ�ۣ$h(Ze��R˴���}���K�����-G�BDSM�2�m
¼��屵}�e�BOz|O���Nc�Wd���A�
��%oN�86M���id,z���W��\�������=�?16���%)d�Xy	�М���ՇX���uX�/1u�WvMI|������9?֛�9B�t}�dn��d*>"B��Ǝt�����]f�����֥�&��It�=�2B���N	���r��S����)�ɷ��Z�϶�@�I�)@dfrJR׶瓄��#w-��}���
�6n������&P�#|����Z)���mw�q*^�-=Ƽ&�{��Q���s�P��k��	�;��s�j�te&9&-j���8��VW\���H!8�RsU���j��A�Z���*M,�Z�������6��g?�q� ���<ϻ�4�M�F��|��9<@�'�m�B�yڰI�?�ܗ��Y��4�;U,��'��;,ء�y9���>��>���w�4u�
��`�U�=�t�k�D���� ��KF�C�ӷ�+R��]}����ǎ���s��S��F��	���|8�����ۦ�1`��a-�dY�����CK�
��wk���z����P�Byx#w���t]�zi��9���Ь=�m��m�B̖�W�#T��c�HM�rq̽��b������<�] ?Ōi^��*\v��TmA�O.Gf��c�/��W�iUذ�@�;g�d�C7OD�9�c���啅�x�'mCP�3��0	vCh�b�sЯ�HpT���'�^�5P�Wu��4�I1�A�.��2h���v���Y�P�B��|��=zxOPʪW�?PY2���C[˳.rS�%�N�Rh=����I���W��Kaw���k�S�W+����Bu!&^���~U�*�0�SC���s"!g��� �x�A^�٫C�kp�ӏnp��{��YՐj��"�0����sSE�Y�e�̇��?�ǸQ�݋$�Jc���2='�	�������J8EW�`�VIPt_���}�lS�2w� ~$#^����l�����_<��d�-���"�o��9�H����3l+�����ydc��E�V��'�{9pS~z]&ǊMm:=�_AS�Z�櫶̻����H�� �*��ۙ;� ��4e�?$b����w�.�� ah�E�� ��(��zF��[�ñ����Zſ��6�-Ǉ� �VH�9z���ߐÁ�\�+������\�Ǖk��Q;���X0��v�b-u��JyP-�f�� E���.��=��p�%�{��@�sՂB��{c�|��.~l�GY�@��&_��q�:fy)n��{LO� ߕ�x���O�Ugq�4�������Q��Pyh��9�`�X�zU���$�'7��&��9/�?�*5C�Q�G��w�]C:����<�]���/_OM4H�Ǩ�`�7	�����<*��t���l(��l
U�=~��Ңd	Kt$N�Z�����Z������t�{+��{G�&�� ��M��A���b<��?�h��f5�����5g�\$��������E�O&C��J��+)�D�gL
�b6L�)��F4�S.��U\J���[\#�������шŦh����C����ݠ�(�qa��2r ӤѥbI	��6��m���Xh�_[��q�R����C��L�r�XKjAL�w�u��t�2�/xH[X�}��Ƒ�K�ApЫ�p���Q\�%� f�u�X/�}MG�(�I��O�p �i�)%�[��\/�UA��z@��v ������5���XNnc����A-���A�0��HQ��&��{�~dɚ<Q����Jj��y}y�%f�?��S�e��:D��ë��*_t��&��XS&f�5K�C�x��ɗQ{����a�*7� �G8:�>�����3֍��r�k���J���Rr)K�",&����
�r��Rǯ_�^�ngFO����̪�Ra�,����)��t�� �OBg[3l�ˋ��k�����A+[w��tp���;!Q}�I��ߤ�"{R|��U��U��
\��t�T(F�L^+E X�w7aF�a��Ax���=�M��.�0�8m�p'�p���Ŗ��2�L������3��F	�m;��2�-?�	�>��G-�J:y����__�C������T�N}ű/Gt|LL hԙe�'�~/�!�EK�U�T�or��¸�E�ż����z��)�!�ыfKg��w�r�-6�A��c���[㓕8G��q�߁z���ݩ�l����]�VM>������e�.$z�-}�ġ����0b��C���ը,:��x��B�U�����uL����(�Imi��|k��H:�E�����4&Ԗ%u>Lw^H�6�6��'%@ڣ#k�"��k��I�X��1����S��6���`3+a��g"M�h�
�9`U�&�'���u
O��hag�����3��粹�M;+��<um��5�4��V� -\p3��HҢ���Y�;�r�^�����LJ���0�V��QH8�mD���-dE9O�g�q�5�����������N�����	1rp*������;�EZ}Sbw���C�#��&���'Ab��^��[F���n����
��Z��wm��V����B�ɲ��ƛL~_FţD�>��� VI^;weh�:-�mfJ�YZmQr!���l(����7����}D�z��ް���ՠ�B֡e1
U����kD}^�B}�O�C�N֌�W�M}�(f/
]�GoK4�у�T�sd'�ą�IjW���\�X���h�0�1��
�.kd�w�	҃��;�պ���P �Kg�1��v�\�#�B�Ό#r����hy�gߞз�@��QO�VN8G�m�+�]�������)ͣ&I�%�/=m}i�pQ_	�S�r��S�I����|��m�2�����\�@�<Wr�Fjשv��@r�#��d�֋��cf�	M^�DK 9��P��`�&�UZܵ̀�Zq�U�^�/�=��&\>���f�M�Z�ݩkۣ���sǏ*t��&�M�d�8%$�W2}T��I�!��s(
��9���Yh��h�M��K6���v�����:��q��*�k�Y���M�g�9�64��0'��"�uҊ�C�?���e�a��=4�QU�|'��),mUy�4ɸ��e4!���4���ّ�J�(�l��u��	�﫡�CN�F�sX��-R��D�0t��.W	�#�_s��N�o翼#K����oPF�y�;`��- ?Q���D���T.�c$V3�zsĕ�H'�B�6#jg���z��؇L ��Cވ���z���B_7��J��T����˃✅#	��5����A^	��L� 2��i�G*����ixA�~.�c��W�gi�/�����;*ߞ�ט�C
��D5x�������Ps�'���P�H�FRC;��Ȧ6���1~T�A�z��^���Pŕ�ur���@@A��BBW�z�G�Mp�gr�c��G@���o�x�����BC��� ��[~��Wk%���%���羮IC�L��Zў猒[82纤��t4�{4�uT�%^ɮ��I��}��;�\����"�($�Sa���s^:uC�y�p�؏!�h���WYH`Z�l��0K�ҕ�L�Ņ�X��7��d����� J6�ݩe8VkH��2^�r	PJƔIW�SBV��_��-�P����w��O$vàV-l�P��d̀_��d�.x�&5D�b�@9��,�e�l>A��L���RLc����'�
9�N�~-�790��*�A�H��ѓ��l�:(���U ����\=I`��Ӿ e���$U�L�4��.�<3 tJ�E������L(^z�Q�[��+�o�Բp�`��@�������HO$�zQ%߃,p�[�;+3#.�ӯ��0��hd�̄NXzE(X#ɦ��Vb�� ��iyÚ�f�E�h.%>B��_��x�	揸;s��x�\�{6T|�7r.��:�r@��_FC�M7z)�}�{�$ 2�ͭ�ߌ��HU��7��x0��k�g��;,yB�)�̕0�K�KUݬ���z'J}�&���/��]��,:OG��.���Г5Z<#q]m��/2F4{��=���S�g	�7��=<<=n�����?N������,3��#�	��Nb���NZiL����V�V?���U{:u��B� tu�T����E�s)h�DP5)��<u�������Z���D�"}�����J0�t+���F���!��*��&���	JJx������\v�!���Ӥ��7�k�\����p��(�`q���2%�ݤ�T�I|N�6aD�����h�_N�qq3�ٶ��
C��%���SK�L�L�D���X��ʐcFp/+��X���9��K�G)�ޖJ��c\�L%��f�TXB�}�'K��?vI�����\ӫ%�Q�Ԁ�h|a���������[ٲ3L0�/2īK>c��}m-6l��j��	;Qgb�%��������𲱀m	��C�}��fw�d�F>��8~W�Z��u*�Z��R�����fkrK�+�xPÃ��r��`�aԜ���b8mȴp���^	��_���u��Lt�RE$ޱU�G���x���;Rzf�_ \�^���gm��(m	_�bE�,Q�����t�� ��Vy�����tƂ�p��YPӌ��V�0�)�<�±�3{����U������Ԑ�!��`Q�Q��<Yj�0��ֽځ��*n��KMU�76:�	�cTP��W���I{A6F��҂��S��/&6��x� H��g&��.��1�+!�br�h��ҥA��4�]A�H�O�n�\�x��{�"� =�nW�y�˙e�]�)"{�S/;`�.<�7(������a�{O����G/���D�;�e�7�<��t��_�ȱ39&�5��1�D>�)�	�^֢���c7�J�����E��V��_�b&�����B�q������`��70�e?����!�p���=~�p����f�"C��{'�J��2�4�R23�4}��>O�5{/�B�������N �\,R�k㷊DId=�7PX����.����vJ2�M�s�]�0��Ky}�:Uz�<eQ�>��n��agd��y
^��\|AKP.7ʿ̒S��TaF����H�ª�7k��`����S5Tf��7)��Zd4�W-��nd+�`��zM/�&#�Qk\9�;�
o�-w�~�_P����_1���߈�Sغ�F�|�̢?�kb��:�50�)P�T�Y1
���$��P�ݢO��]k#�4����u���n�]ό#�?O�&?���B�2�fH��h+�7٠nHw�SY�΀ߎl�5?t�$L�i�-$��X�@��x%�X�,��.��K��
%9�u�^��c���ῐޠ_��3j�^wz,�v/� Y�� l�2�H��&VD�"���R{��ֻ��?~K�ٛ��e=���
Y��8��W��{1�r�d�z�M�N�HbGHxYj�����-+(p���Iv3D�4�G��l�F������[�@���O,�3e-4�7��A?�D����N���@���e���6�;1w9%����{���w��[S��1���_\犀�h�0?��F�����vK>���B�����q����9y\�x����C�&���^�6�=�e{�e|��NDr���߄-�}֓�_l�&n�-+	���6NP@3]$<`_ֆ�vרs�I�33�6� !a�iK�_.uagжr���5��:O�:�\6�]�wL�G�gLu��:6ƗGY�VF��O,v�И���"�gO�i�)k� 1F\Rw�}��9O��T�6��8���,)�w교~\�|M������@���/�.)��nm�K�v��z�.�5�JC���#�����,���+yy��~�H�_x���{*�UH��}P�[6�
��x5�ێ�}0���jo�JK?<��A;��� |��6®l�~�==28�A�j�����ˬ|k3���/���(���d����	�r�HW�ؑ{v�RТ:��s�ioOV�c�5)������hߑ���o��c�����@kPa.l@�gg�N��0j�O�x�mlSk)q��Y�r��|���E<���|�x������"
��HizI����?�-EO�
;����a�Z�u����D�RR7��#�Vi���	,��M����$�QjqS�z�'�E�XպZ�,����35�	0�����2?��-�߲>�k�˅YJ���ӉN�Ԧ|�����k���=9�p����h�����J@X�;%�d�Ymq��>u��u%�@��`O�r�a]Ѱm:JC�紭�T}reK o��~ŀa���g�h:>ޕ�JLx�P��ה ���������}�&�h8~a�k"U=��_�9h�h&ˑB��
4O�'�a���Ĕ3�SȲ��H;3�2<}���='���kK 5;-�H������;܊|�fC��֔LR~��n+V���H@�mLv8�5f9W0�yR�����G$�����VB�a}���p2z���7чY�M�PSj����y"�z�.&��I�Aj�T��\�cŊ�q��4��+\����m��V��f�J�Lɺ@��T~�N�L�L����VQ�|;�h� �u'�a��Qz�ã�q`(�
g������T}LHľ��U���6ըBL��m�
]X�����}T�B
4�O���N�%YW�T�0a�
e��o	(M�O��\8d/��j:W�A�\����U�8y{1������d�L	!{�����ԾXl<ST�1�UHv�lKd.�J����
zo��\}�oT!п���Y���^~Ojj�3�]^x����1k&Q.��o�=u�;�x�y	��%r���S��"��������uJඒm_�$F#@�g�r��Lױ�߄H �#�����ۥ횴i����L�;A�PɊ5�.
�Z�f̈�gq�.X^�)$=4&d�ۇ˃_�Ut{�\�k���T�s�t��u&�3V�	8-j|W:���1F!��s0��A����9�ە�M�w��Sů���ӥ�IB<3q��s�����=M"9"o�a�._�غ'��}-w�KT�?�:��m�����E4���U���'�=P,PPy�x ��g�<�(�A4���ٙ�u�0����y����+��K<�F�"��Ҟ�R�ML�8&��6J9�+�s�jG�
����Z���N�wi2ہ�`�\-(w�TеL�����i^ԁz{���P*IB��D#rL��Qz�跇T({�KV����R�Bg#ΧR�T����R����\�#����]�Iq���7 :��i��1*��u��_A�?L."f���\����W5;i�Mͮ�`o;2�!��Y�C�D=����yk���X�'��P�Vn�ACC��Ȯ�v��=T�ζ��f^��HP�e�uz|��$2�A'K�J�!���d�0��(�k�
�O�����$x�wʪ��DK;ټ��[� �7�%�;�-�����IKf���Ѧ�ǒc���"����Ŗ��Gu\c�^&�7���>хHIC�j���"��[s��;�^B)�C���p���)^���I�YP�l�tz30&��ƼT���'U���V��l�1��_J>��m�.^/��x�z��J�;�W�ۤV�.�_�-R�;��)�w��0$~�è�ul�`��lݐ_�d�б.	��j�9���mԳlF�Y_��Th��ZGb��X�'Դ9��z~5��AP+��,�F��,����� �B.�˜ �Q�d�*���Ʉe�+�$]u��<G�.��5 |zE'Z��-e$��z�En[�^?�w�V�x�%��՟��g����HW?lzY�ߋ)�c�W+;�����C�8H��p�>̌��I�X+Nӡ�9b�Ђ�ey�cf��E�J�.-ʕ��lW��zp�'xs�@C�d3!{>�|���.��B �@�N�_N�a�Ux)�V�{'�� m͵6����VU�B	���9��l��oi*��=yJJk�Թ��SQ
U����v'Re&���/݉G�e"A�4�G�	���j-�=�P<+�9]ufr/:��4��8�E��[��	6f��T5<Ef��p�G0H��Ė����`�	���Nj���Zq���ס��9����{B:Ө� ����\"Ց�ʁ㨝�hȯ�51�����������;���$Lۂ*/��� J8++$�J� m�)*ӎ�C��.�L��J��M���\~����aQ��S�!�ӗsSz����x"'(�E�q�+�2- ���|yI�w�6i���/���Tz_VP�q;Ң��v�C�rj��.K��L�W���̚㲿�k�J/3>X�*z�A��K�����1ܝ�(\�%֨f���XJBv}��6�"�I�6��:�d� %\g�;K�p�x��&��+��;X<���ĳy}c���=�->=��\L�<�Q���3��ٺ��rI)���J���i}�Qf���N���@��_�L���*�;��Z�8���\f#%K�P�xX�o�͈����}a=?��VR8u��x(��I��@�&�^�ec�Te�RM6��]�wO�H��a����R��_(�Y^�-
g!&�0H�g�M�t,Y�����t�����5�g6fl�d�/����Ag��2M�t�j����^����z�/��uA�OU����:��6PoD}/��'�OC�㌥�O��=(���Z{��]�st�mC)�,&��7�6Sf(Y-\M�5ں�Da>���c5���*�\��O�����J��R���F��X��%��䝵̭��9�-�s�<�{r�t���ب:���3歐)�r���3�R~	O'�tV���:6V�LSL<��+���*��Y�߇�������Zf���ajHo"��`��|�9�t�&�0��[�U�O�a��:��3y���yN;���<�t�#�B�| �����H� ��I�H;�1����D�^>�L�ހ��rV�'�H��m�X�����9����=>҃�b"~4��C!��p���G���ifpv<�]���Դ9S����+��7��Xc�S��A.�g�\���'d�����j�Pr��i{m8v^V�c��0x�~��[Fٛ8��E�(���jV��;��h�凹���% �Q��գ�0�(١��Y���B@}��H �s�4��
�B�,��?4
!\��$=�}�X�BN��Or!]N"$wW��1�t t
)�oM�W�㻠��d��A�Bm�W��=\:�ጝ�|��1U�:�ݚ�d�m|	e��a��5������m1��Tv�( ����1�����pL����Ѓ��c�����A��w��]���ׂ���&�ߔSI\=��ݪ<^	8��rt!S�bL�6��h��9���փ��$@�rdr���k���#��̢�����Ͽ�!�Đ���P'��.�Z(j��L&)q�LF^s�=E�&(���$����O�k����v$s�|�t�k�&�_�^8��W~IÀ��!��^s�h���`Š�>�>�MK(Ɏ��������Ig�q.db�7��t/M�mI��oq�&�q'�h���q��?�v�1s�խ�4�U���'o��,W#�y����O ���)4T4�������q��P���������ZF���Ӗ��Rׇb�����z%ǎ�K�s�&���)��8��[_\�����E1`<L-����L�֤�	�G�ar��z?�ٔBk�#�*����z΃��Æ�M���%�:�B+�o���fTǎ�<�Q�(�g�M�x�6��\� ~|�i}2�*�K��7�AB�R.�|j�/���WP�it&��R�;����#�MC�V�D�������$��v`'�P��\���C����'���T ��F��^�kP��u�ֶ���WAkFȪ:���ؖ�h����B�/}d��i�Lx�vi�����5�̳�[��Qa!%T�U��i>�3I�J�^��jN�����}�D0�G��u�jR^��u��:�I9�������"��p�&W��FD^��C՚p�^�mk��Z�ZY�Gë8�W0Q5F��Ӽ�����M��>h�0��J*RJ�]����"�2�Fl��>l�JQ�W���V�_Nl���Ri�)�w���$B�����l�����W_��dJ�α�l��s9�����l
��[����-ݞfYƵ`\'Q��9��6~y�	���ٶ��   �  �  1  �  ++  �6  �B  �M  �Y  �d  �n  v   �  ��  ܑ  9�  ��  ޤ  "�  ��   �  _�  ��  ��  P�  ��  ��  6�  y�  ��  v�  K�  �  . � M" R* �1 �8 �> 0E �F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<���C����P��1�ޜ�F�Ai�K���3bH-D�x��U�Y@�L �2�3��??�
�"�^��"D�*N��UOB?U�E�ȓ0�v���,[�� ��T�Y����ȓp�s�MӶs��yU��9�z`�ȓaZ`�;׎R<g�����;UU
)��X��qaE��?F�d�$��]�ц�rBj���H?�dg�A�5潆�%�:��(�j�  ��I��ȓs��Iȟ&�������~_����@J�<�%��"@+'I�WưH#�'�����˗0oءh�hY-O�xm�
�'�x bi~����N	�/>��	��� �5	1�#!�����:(D�D"O��B� 0X����IR+9^���"Ol����yӂ(��'<x	Z����	�j��[�M�e5根b��O<C��K�����'�a��`���(
C�	Jmry;�	('�u�!�B��B�IR�����a� J݂ �F����B�"'ޖ�V��
yH�q'$ʷC����hO�>�R��L�%����)��x%��Z�a=D� j��K\L�B"�35T��:D��qc�gN�x�&+
�E�U"��6D�ػQE�2��B
-m���颭'D���c�57.E��\�Ĳ����'D�����G�:��#%�$rR��V,%D�0%!X�Zք�EL�~4J,�@�.���<q�.uR������0G�y���X�<�bJ�?c'hA���	�$������]�<��2m�~i�FHͧ_�\Y���p(<A޴Pd��J��?�0�_^�y�ȓI�i+AI>0�L��'�ƛl�����6�X�9���&[^2��� -��T��~t&���\�(4��C��?�N5��Sj�pZ���k����FG�\��@�ȓ{��؂4�J-$,فW"L���ȓl�8E��3zAA���2h�م��zy���w�r�.������R����y�b����9���p:)��%���O��G�4�03Nx�A2f� ��xPŎ��ybJA|��|3���p�ˣ����4�S�OVxDG^R�H���ʨ$R��	�'B�T���X�T4�qk�W��
�'a,Ƃ��j�	��C	���yR��G�4�8��
R�Ip��8�y��sV*�򢫜��*����!�yAW)W�pl�4�y@��(l����	�'8�MI�,�1�6)��l��X��'^��N]b}j�����/����'a��Z��°O��Y�F��`�N�І���2����g�%;Z̀!$C�h�b��F{"�'���%ph�bE��6'�:�ˆ�	�U�ȓ!JA����T�ai�7L<��>��'Uў�M`�jC�Ԏ\%���AÈL��C��:!��M���C
b���ۥ���(:vC䉸 �Xe)�ꔹov����^;wF#?Q��iD4?��|�&�·��S�Nե4���
O�)��6D+��B��Ԩ��6Z�8D{��)Q�
F)PEn��z��V�o!�D	�5~����L�at�����w�!���^�)��ԫQ�p��U5yQ!�DV.E�̬P�#��w����2�W8gN!��I ��W [�>�n؛A)��BA!�DJn�T Vm�^��i�h�&^!��*I�h���G
ky@x[�%
B!�$C9:�lu@w��'sX��;���d8!�D�:8���(T��*��S� �����<y������3���E��h�\J4�~2�O�=�}J5mF&Vy�Z��12l�U���Hg�'u�yR
�=ͨ����Dcz��$J���'az�+�g�����C�*=R��,ޏ�y�`�_G�Ѣ�o.T���7o�7��z�C9�� m4��a�����xC��ۋR�t��dh��d�� ��G
�@���N4#K<�ȓ,�2l	S��{pz��VJ��h��Yp"�e�I(�:��a��?���S�? �=pS�޶9�TQ�S��)V�,Y��$�OZ5Gz�O�@ek��4�v�	bi�o�u��'[ζuI�7^(#�[�nm&1�'-ў�}�W	�W�T]��h�
��avŚ|��<�>q�F-~�P)�WHǢmx
%��CK{�pɦ�=�O�$�g-�p��Q!��(,�x�y�)�S�INX�J�-�!p�DqpK�1r����(�(O?���ɉ6����C��^���ɔ�UE�'��y�LȾ,e�8!"�o͌�;T$���yR�R4�3����aR�}�c��yҏG�=�P͸3�G�S�V������yT�M����1D�`u�Ը����y�'H�f�Q���^���&bW!�y"l�6H�gS��X�M޾�y�J�?<����쓻G�%�%nA��(OZ��d�F��4�ۗ?�$,����,Q��D���֨����-�]P��OX� �ZQnMr��}�TD��'�<�����=*��$`04NE�Gj��SF����iN�n��P�#���TԠ;�b�Gy���)G~��YP�%gՌ��U�Q풲�0>ќx� P�Q2�KքH�.�
�(��y��;�f��u��s�DA?�M�}4O�>n�r��I���˺�"T��""O� �#(M7_��s�+��;��dq�"OQ�B��Y��
�jY��9��"O�����޳l�.H�+F<�L�Ǔx��'8��z�`UDSQbi!o|�P�	�'��5R���3YZP��)�8>��';b���i��q���s���qyL��Ҋ��)�)*T�����M�pPM��D`�!�d�zk%X DM!MwhT���ɹG}!�D���19`�h`�1�%�:{{!�D�d�B��i(E�$�4E�<!�>6G��{P��#r1H�+A�$+�!��M�5kA��7��R�΁�
z!�D:�����-��u,���j*M\!��ni���$_�P�>���Ӱ@!��C�G �$j��I0yv~��U�ի#!!����J��67l��+B(	�!�d�-D� �q��v*½k�ɦH�!�d^�G�j��QM��&
N��bG8|�!򄕐9��I�bX�Ic�(��.\�!򤅐oӘ�@��U<XЀ:��܁�!���$���C�	�;^U��9�A�W�!���>�PU�v��M]Zt�T�A�'!��Z��E �K=LLd��Y�v�!�$UR��!�$EM�k2�hbAԭ�!�D�6jX2�rM�[_�)���HH!�d׌g����E�kN�ԂN�F!�Ϧ'N�@�5���<�x3��AB!�T�B`��Y%�K��FAje�^X=!��lCV�["�H����Kˏ8E!�$U�>k~�X�D q�թ�"V2!�
���	1/S�t.Dh�N3;!�A�@,�Ma# @0%�a��8C�!�D����k�e�	 �3��!�ćU�S�퓘~ �0jU�ݙ$�!��C�A����>E|�p��/%�!�}��=����\.nYy���!�$C�}�8Q0��'�y�ɐQf!�D�a ��^�sh��HA/DJ!򤇤��X���	U�8[��8�'o ��W N�N"x$���=�|}��'���
P�k
�5�&씶j����� ��H�h��X)JWǑ9(k,�a"Oy��	�&q�c��X�9b�"O`Xrrg�+|�*P�E�D��z*O�d��	�1$��9�%�9hn���'M yb�D�uv4� ���J ����?���?!��?A���?����?����;�M>�P�����]P��?����?����?���?���?��{"H� thN&NC
9��K��Ckb����?���?����?1���?����?Q�ܸ����62��eS���Ng�X
��?	��?Y��?i��?���?��n�@�X90�{6�^�`�����?i��?)��?����?����?I��9��0Y��Wj��Җ���p��b��?����?a���?���?��?���	�<�Z!�Ӏm����s�T�\. Ai���?���?���?9��?	��?����D�&X�Q����VꝂdY|3���?a���?����?����?���?9�(��Ipl�hꘂ2���y�$E���?���?I��?��?���?���&��	�r��`+:�D"L0t�T�����?���?i��?��?���?���$V`��t���+f*�ӫ�`kڝ����?Q���?!��?1���?a���?���VJ�*A�\�p>�Ea�
صx�B@���?����?����?����?����?��ϦY��<=xD'w���p���?���?Y���?���?�Q�i.��'?�� �U`Bt�kE�¶y9��Y�'�<������8!ش�,���#Ɗ?�4ЂcF�02(v�����{~r�i����s�����'M�
#��:!j-..*1q"C�Oz�d�:�87�1?��Ow@��9�$�����鐬Z�0�Hw����'�bV�0F�D�\�`;nh��e�V>�U�%�
l�7m߸`^1OJ�?0����u�ٲ:�v�WH��J��쌮�?���y�P�b>�`�Ц�̓d�A��i&%���FA��R=�̓�yR��Of8"��4����G*^�"�h�.A2�l����Œ|��<�I>���iɚ� �y��*D�2=)�"�:VH���� ��O8��'���'C�d�>	$ Ոh�$�9��!���A��X~��'=�Z#�J��O=��	z��@BaHIBGeS7��e80eƶh~�IUy"�����d�aB�Bt��4a�<��'�
�����18��<?!W�ig�O�I��N��a�u"�9d�,��n���$�O�d�OpK~����tJ�8�d�::�  �-ܼ�j�b*Z��䓖�4���$�Oh��O�� |���%,�lI�ޑ�˓$��vC��b�'����t�'�jX+�](O�(��V �v�#e��>a�iMNc�b>1��޶6�$9�I^+�b8dF�-�4+S/�ӟа�)�C
���RM𺋄�x���<���	,f��禕v~���6�?���?����?ͧ��Ҧ�XM�����X�|�|�'�7Zv|���D���D�޴��'6��>���`w��	o�$i"�� ��q�ʲ@^Z�#�
����3:�QyHF+L <�
����W��I�.nH�9�+��F5���T�7�y��'���'%�'_��ϯ`�`l�2.\4cl��A#NVn@����O��$�Ҧ��V%�_yb�"�O,�5L��$��\��#	�x�Xp�V��q�I��Mcձ����J@A����\ �h~�,���$��JٱL^5D_�X�ağ��,	%^�h	�4��d�O����O���Xl7y��K[33>m˷��>JҶ��O�˓}��)��?!��?�-�L�Y�NF�v��H�0ӣh� r���X�+O �l�`�&��'qn�D�3OL�T�D���#&(���O�}�8��������ۺ��'�OD��)O�.�V�Y���d����(L��n���Or�d�O���)�<�B�i�Ȅ�U"נ
��L�ԏ�9�&,	�
Z!��'�J72��=��$��Ǎ�oI�hc�M/6p�1�i��M�нi��Q{�i��	�n�@sD�O3p��'R�rCXt�2� #�S����` eӀ˓�?!���?i���?����)L*b�*��$�U�O�bY{v�Z9:�NTnZ�����x��X���b���k�N��d":�i�FQ�IS���p�V�蛖`dӞ�%�b>����ͦI�I㲐�b�P�SH���7�J-̓+�buKE �O*x{*O�nZky��'�r�L�"���gj�]{�GGy��'�B�'l剹�MK$/�.�?y���?it,�:�Ĵ�6��)&�8�#���'��Y���E~Ӝ�&�t��'��(�� 5�Q1꼽+�(?9@��
���rV�V���d@��`��O`E������l
�е��)����R��?���?����h�B��N��QS�lڨ�6$M+�����Ѧ=y��Mڟ��ɧ�M+��wW��qTˉ+:������?�i��'u�6-Ӧ}h�4Y����۴���C:j,���:����)Ȥ��3 /-��
�Ȳ<�v�i,��埼����	����I�.t��Av���\�0.�"�����3�Fy��'��@Q�`�G=`�TLC��V����XO}�Fz��oھ��Ş'�z�re�2��;qJ��#DY	*��⎗�����~U8����\��ʓ=B��Q�� mQC����p�T0*z�U��+�ʟ@��ޟ��I�By�
mӲU��D�O ����X<`�v��@�R3F6
8�4OPao�l��g���5�M+�i��6_��ޙ�E*�/=���R����S7��Ѓiy�f��"ݐw��d��*O����� ] REߠj�A�Pʌ�(�1O����O��$�OR�d�O��?qIb�����/O�T���֟T����ݴ�p�O�p7?���(ɮ�	���%; U�!$em&���I�<�|�X�ok~�HӚd�j)
��� l�X��@��X�Cr����R�|2X����ş��� ��K(����D���o,��������{y2�iӾ�1֥�O��$�O˧?��4 %��i�N����0d�'���?��ʟ��i�Iڒ3}x�z���x_X����M������E�.%8���|����O��pI>࠙�c��ӥ��!3��$��Eހ�?A���?���?ͧ�=�R��̦�D�.J�ɡrJB�U��ꗫ�GΦM�'�\7�0�d�Or��'���&��M����O����4R���!�i��7-β�@7�h���ɾhɞʰ�O�����XS �q�pJ�G>�4ϓ����O��D�O<���O���|z�T?/�d�2h�#=N@p(���4�Ƌ/P��Ѐ��')��Ou���'wrk��ܻp\��je��r�����͏�s������Q�K>�S�?e��.8JʁoZ�<��D�h͌���f�"+`6��L��<��L�fn���������4�N�$F1q+ `��tn��J��F�%� ���O����O,�i=�v��7yB�'�֎E�nq���u��b���r��Ox�'�B�'�'l&���J� 2���� Q[ �0�O`H�3�=0��@��$�	�=�?���Ox9��Js���m�#X��q�Oh���O��OT�}��RO��zr��)riF4��ؿC�l!y�ۛF�*f�B�'��6-!�i�%hq��m�PE� Kh/xa"�f���ILyiQ55#����t��A '��$��,��`#A��88(<��pF\�.ph�$���'&��'���'�'��"+�]����Y(a��}x�Z�l1�46������?�����'�?��DȰSBؐ+�n�<<�,�j�H��_e�I��`Γ��S�'[ �GkM2er�yR%)L#R�@"� ��8��x,OL�k���?Y�e9�ĵ<�Vl��T¤-Z/2=��D��?1���?1���?�'���æ�������`ؕ&	W�V��c` �L����m�<9�4��'(\�
��~� �n��L}��@�A�n\�ٰfb�.mi���&�G�a�'�����o��?��}Z�;t�PA���f.U�`l��K~�̓�?����?a��?����O/~�{V�?w�����ى&*H�#��'�R�'	�7M�\��)�OrAo�C�I(Yr�)�#T�-(鈒'�	D4��M>����?�S��nAl�@~2J�.\	� :e
�3�k�6H!IT�(�Ò|BR����韤��ϟia&L�z�C��C�<"l`��ٟ\�	wy�zӌHYf�O��D�O:ʧD�F%��&G�dp�:5��>kڨ@�'����?I�'m���i2D���w�D�)�5zf/�a� �%���qq����<�'��d�'��'j���6*�┬ݵq�P(����?y��?��S�'���զ�+��
�F-a&��m���;�I�}���'H�7�>�ɋ�������/@=A���� A����a�(E��?ܴU�|��ߴ���� F}�e��'x`r�����$E`S�S#)��ϓ��d�O����O����Oz�D�|ڔiL�Q��Q�A۩k��B���n�B�U��?����?�L~��]��w(��Hu��hﮀ"�B��r�Tu���}�nyl�:��Ş2;�u;޴�y�'�k"JQb�J�Y3h�U�T��yb�
�I���]��'��i>����L3Pe`d��L#�����G���I��$��ǟ�'C`7-ɪn�8���O��\&#���f� z�>�2�CF�;��TA�O��n��M���xr��!p@�2���Q��	�BΎ��$)C�Z�ٴ@�<1�z����<����x08irhͽH��af�/8*����OV���OX�$%ڧ�?	���
�5�(���D��b�=�?�»i����2P���ٴ���ygo�	oy�Lk��> 6�}c��8�y��'����nZR~r#X:6����o#��J�	�r��*d���2��|Q���I���Iß��ݟ���C.SH���4�&�P]�uk]y+t�D z�j�O��d�O蓟��D��i_���I�F�X���<=j��'�6�Y��'�b>q�C�CMkp��*�,2"��pPgN�&��)�&Uy"���9���ɚH�'��	�b�lQɃHG�t����J�'���Iן(�IƟX�i>5�'_T6M5F`���- ��(+�m�&k:pBGe\�u�����i�?y�\�8�ܴQ�b�i#�R�KnR:` _�'���$�����4�V�R
r���ƒI���i3 ��e^���޳F�bd���p����ş ��ӟT�I��8$?1����?j��c����m[�+��\X�`��� �I��M#���ĉΦu&�T@���K2 �S��%b�l�ȴ�D��ƛ�osӬ�	TD6mk���	toX)cEO�;>��P�iGD�R$B4T��� I��ty�Okb�'�2�̒-�Jh����.� �beΌ�S>��'��	(�M3d���?!��?i/����cҝs��t���,I�
�����O����O6�%������ueM�<�V�[���g�@�WIG;9�b�(1��Z~�Og ��Ɋ5J�'t�-k�J�>X!Э#6o�;�B��'���'���O�剌�M;��̾3UL����Va�MB`[�T����?	��i�OL��'�N7m�&��S�&t��bp�%o���I�5C�˦��'Mr1��l��?8�Z�� ���E���Y^V@�C�]���j�>Obʓ�?���?����?y����	T���\�����\�ATK6yr̵l;����'y�����'�7=� ��&�	�m��"e��w� I���OZ�b>���/����!T�[�a��bϾ��E&ϖU���u�S�L�O�l�J>y.O����Of�ce%�Y%�T�s-�/����f��O���O���<Y�i"ѳ��'�'0��
���j���F�V�Qd��耓|b�'B��=���"o���&��'�A3��A�V$|<�(@cd�l��	D�`A֌�� h��bp��Oh�2���}�A/�-�*����
@�<T���?I��?������?����?��9��BEn�V�r����Շ�?�S�'>��y��?iV�iv�'��w�f�A�Ӭ;ؘD �"+LZ�k�'�87�Ӧ�:�42&���ش�y��'��R%��?�!�a��9ctm�tS�U��H�z#�'Q�i>�������\�	3P��q�n،1��k�#Ǖ-޺y�'u�6-/`9����O��D'�9O�U���խC��q����2ѷ#O}B�{�N�m����S�'L �H�$gZ�3J|�aюהcv��؅��qr���'��lX�J��L�a�|�Z�XIa�&�ޅ�`I�
v1#�MQӟP�I��0�	����ay� e��X���O8*w����(�Ór�,�j4��OXDm�Z��%x��ߟ��	��MKV�X8�^��dc	N�@� Rk�h�x��4���H�z�v.��@�>1��6Yh��"2C6`р
>r���Ɵ���؟t��ܟ���l�'6\L�B� "k��$��`I�0z��?��3��������'�7m#�$G��m� �ͱ7���ä.��o{b\%��BߴXD��Ow6TAT�i|�	�*�\UB��� VI#W�;B�5*���#Vd`�t�	cy�O���'�����X	{Ì�3��q �I,c�R�'��	7�M�AA\�?���?�,��t���\'5�L���ΐ4k���ƕ�	�O.���O�q&��X�
�p��\�����g�Τ_:r��U훎^~�����Kx~�O����	�p��'�(�RQBX�
��`'� Fx��p"�'0r�'�����O��I9�M{��Z�bvH{�غx�(upGkϨ%��P���?�Ժi��O��'�Рq	����n��m���#�E��	�!y�oZ{~� �'	�b���=��IFYt��T��g�IB��{���oy2�'2b�'���'�S>�QS�I&.[NH�cY,����7���MK&	�?���?�K~��ћ�w�$��O�T�FA����/��:%jb����h�)擼=Hl�<Q �jr��FC. ��(� ��<�&�97c �$�	�䓵��O<�$�'.��)q�e
�w�l4�����\�T���O��D�OFʓXv��UA!r�'���;df�Tjj8*���2�*Q�Oh��'�6X���J<Q�H]1k�B\���U�<5bqh��C~"�ņ4��$w�d�|�%/�O�dZ�?��Y���a�pY�Ο�\�e��?���?����h���Ӿ1<�H0�.7<
p2$�9x ���Ŧ��u���� ��:�M��w�T����Q�KRE�tD��)'�(�'���iC�7-�(x]�6!?9��Ĕc��էM��`���Z���刀�ouPT�L>�-O�I�OL���O����O��x�ꈤ9pE+0+�4 �b])���<�׾i�8�$�'���'��O�ҫ*#�C$�3 �65"��N�Iژ��?��4	vɧ�p�B��!k�%[r�1
@dK Co��!FL	U�� �'�ބ��П,p�|�]����n��/L~Ipr�� aR�<� bݟ��Iɟ`�	Ο�`y��Ӡ-c���O�X�Ïn� m�`̈́F������O�Xlb�?��)�MkC�i�Z6-\�MMRL��D�G���F��|��1P�m�,�z��4�*���>����0���w/L�0�r$��*��/
 �����������I؟���a�'m�~���)f��X�� XX�5����?��d�"��$�'�x6�9����};>�A�Ŝ*P0�i�����&�`�۴#v��O��D@3�i��	_Ov\��< Θ$〙A�E(��S#C�B��y�cy�O#�'��M]� �H�qDe] ����ËGS���'t�>�M�?����?�-� �9f'��,pP�w��4o~u�⒟|�+O<��mӺ�'��',��p�`7-־0!�i���ҡ]	)J(��`m�F~�OO�p�ɗ!�'@��f̓�_� �NT�)��P�'�"�'�����O�剁�M�~T`A�`V'g(n��H�=9*e����?)�i�O���'�P6��\_��"Q�'N���X5&��@� %l���Mk��W%�M��O���TNN'��M?�#�?.c�Q;P@�)n%xV�|���'���'^��'���'��nX��+#� dk�K%a�	ߴGa��a��?�����O�6=��rՄɑ>�Pp��2����u���IE�)��Û�F6~���&I�,�]@��]�I�7J}������eRo�F�IGy��'�b�զdG|`�b�=^C(�{��۫k?�'�R�'����M�2.W��?���?�ܿ>A\�q�FE�s��[Q�.��'LX��?q�'��'��]����F^N���tl� ��O�� �!$�J Q�:�I�!�?��OT�ĦʤQ���˜�{4�3�h�O
���Ol���O��?my���˟�3����i׆��QG�?	�Rq�����{�4|�������?�6�i��_��s�}A�(ӽ\|���ԫ&�&@�Oh�\��4l�&�i�r�2����㟈z�gB�b���)3� �TSPKζU���0��UC���` )�$�<ͧ�?I��?���?��b�$J�$K�kI�C�P�;P/�9�����]�
�����矰&?�I��tI�L�K0��FF)D��3�O��d,�)��6>���fH+V��e�Bf/gB\p��%B<Jj���'���qA��֟��ƚ|bQ���d�]�[+=��M�U��Ar�Cޟd�	˟�	ӟ�yB�rӘ�I�!�O���ҥ^�~��5�2��?nm�Qh��O<Am�w��|y�����	�M�r$�+]�|pu�W>З��	+�����]�'��-�פ��?��}���=_H};a��bb>)��ڮ+X��?����?��?�����O^��(�ꎿqF@�z�k��E��:��'���'�6M�&�	�OB$l�~�	�8yx��g�x�ٖ����2p�I<Y��y�'0�ڍش�����f�C�� 2B� ��jZx��A��	�;�?q#%�$�<I��?y��?qc��"j_~���)�5>���☡�?i����OŦ�Z dQ�@�I؟ДO����K}fp!�F�?!��,P�OD�'��6���l&��UX�L�!�#�����
@�K���E��A �Z��4�=;�oeO~y�ҊD�Hn1�#FW�Mntp0���Ol���O"��O1�˓|b���<�x��ջ<�(�	@mqD�s�'��d�2�dj�O��$>�|0ՠ��*_"ԒVN?����txm�p~�I�wP@�ӵ*8�I�D�~�j2JT�fH��s�ʿh�(�Iky2�'�R�'���'rZ>�KQ@��p���7�	x�����hV��M���"�?9���?���P�(Χ�?釸�y���풙k���v�� SAY)O���4�����Oν*�Em���.I���`U/�[Ҷ���*�4�.��VÂ��u�'�2�&�Е'��']���ն_2JP�c���|��'BR�'L�]��ܴ&�:�A��?	��+̄ ��$���q���ё�r�>����'.9ڶ��8++�������A`3?Q� �5Q*!p�`̃��U(����?i3N�?"�R�$��0�FIR����?y���?Q���?1��I�O,�%��N��J�	˹+�R̢n�O�il��FP0i�	ʟ�ߴ���y�mU�a��\BJ1LA�B�E��yr%k���lZ��Mk2�G��M��Ob�bWE����6���3�T��5�M:y����$E�"�8�O���|z���?���?���2~�7���XP#Dγr�*�U�d�4>U|e�g��<����6�?���j���,�> ���q�F<:���SZ��Iۦ��M>���?��Ӥ ��1܅(z���'��Di��yfY����)���;�b�O�ݱH>)+O�58w��im
`�g� �t�$��O����O�D�O�i�<Qƺi5�'| ��h�a|��r"�!�u��u��ݴ��'������x�,�l���rfW�R�,��G�-Z�:�$�����'~� H jE�?��}��;M+������LB�19��Yi$�(��?)��?y���?I����O�<(h��ڿmj!�֢N�@r����'�b�'i�6M�'pSD˓����|��� !�fF�_�艑C��50WΒO���b����2�j7%?�Rf�MD�}����=Cl��Zp@����u	d�OD�;L>,O��O���Ovt�Rkv#>���.^�v��9bE�O����<q@�i�ر�u�'.��'O��O�M�qi�E���7���@�*���˟�l���S��k�!܍c&J.o,j֠��J�&��'ϷL���J�O���?���#��}-�� 5�e4>`��+�	�X���O����O���	�<q��i�h���߶� ]����)�p�I��
n���'q*6M1����g�`��"IoܘZP��."M
�2F����Iܴ�5�4��M"o���'��3hE<��EE�"w��و���.HV��I^yr�'���'n��' �_>�f	J�ڑ��`D�}�9��?�M�p�;�?���?�M~�.��w��bs�Y�c4$�w&�qݺ*��'�d#��	8��6Mr��B��M3����_3Jo�ic�b~��є`Y	�R��d�Iy"�'�b`_�M�H�cD{w2��aעdR��'`N�K`�'L��'�M�4��=�?A��?�'��0!c�:���˔ ���䓕?9�P�0��4��j���Za�YrJ�5�>��v�C�- �͓�?ѣlD�u�T�"ӂ|~��O��}��JD�.�+`�N��Y��)m�\`��K@o��$��K��Sti2I��\4���I����5��#y�� 
sNKC�f��"�[p�\p���.C� E�ڲE1��F@z7
LrU9ʓE4�	 f�A8���N�)D��؉p�U�skb�"� �:͜)�U
���&���� T%*S�M�'P��x-a�Z�����(�dY*eJ�d�m��
6.l<J��H6`޴
���+�Đ� A��|��#�dH�\�͢0�<l\�#!I�*>4���2o����������5��7:���'�u����?�.O.��8��v��a�aC�ɐ�c'�4w�D4�'B�!Qv�����O0���O��d�O45sQU�	ʉxg��K�L��¯Ul�t����OT�ON���O�q�vDw'6钑��<-�t�����f:������	����������-���	�cxLa � &�)�D�.J���ݴ�?���?AM>��?�g��jG�o�b�  Af7C5QF�ϻB*�ꓘ?���?Y��?1P@������O>��U�$��B�ל/��]WĘڦ5�ID���0��<t�La
!����dk�DBL�Y�|d���'N������q���'���Oߊ�X�+.8�0m���h6(����<���On��3�p���g�? "[4D[:|��(E�Y�:qf�x3�i��I/l|�mϟ8�I��T������Ɣ��ȟVk�t�֌O�<_~9�B�iy��'Ш˥��;�S�u�����L�7�Z�i�f\d��d_�7��O����O<��t}�V�|����<a��f�L� �^@SFE��M�����?q�� t~�	�O��`�%��(�b���)Z#vT�D��Hզ��I͟@�I:XB=��O`��?a�'�0�0 Fa�xIt��܈	�}�+Մ"c�'nb�'/�(�;�x��lٚ�ڬS�i&	��7��O���g��[}bY���	I�i�)�F�!~����!����ɸ>i@������?���?�O�A��䙀g����� L$f�lģ�ɰ�����d�O@�O@�D�O<�X���4ͩ����	��ٛB�F3�2�O��d�Ob�d3?��7���I�`Dy'ܒ(nl���P��MC(O��?���O����Z���䞸Fy��f��4x��`!�l��c8O�$�O���6?��&���i�O��ӭ�	H����4�AA���3�D�q��u�Iɟt�	u��b�$�g�Z h�ˇ������CrӐ�$�Ox�Y��L«�p�D�O�i˞?� �
F��@�p"_
Q{2l$���	����eƔ|���Ԩ�2��ؕ�����X��P�MS�O|�a�N���Ob��쟌,ԧ5�%�BB�4	��}���a$�G+�M3��?Q�ʋ��'uq��(�Lү����z�`	F�'��bv�i��'��Oh���$P0p�&��.W�	�D���PnZ�5j�A�	�^b����O|"@�kf���,X_$q�oE�X�7M�O����O�(Pcz}�\� ��l?I�o��c�"�3 �5T������8�T��I>���?q�M:�)�#��I��#j�8]�"(�F�iz2�${�B���D�O �Ok,����������8h���1��I�G�h$�X��p�	Kyr"�g��1��49�UQ�P	43d}s�//��O��$�<I,���*�xC"�~��A�(��au��ǹiCr]�����x��uy2�ݧ>�S�B�	riY
+�8!c@k��n���?	������4����14j@ڗ̯]v�k�̬`fZ�'a�'}�R�@!���'�����$�F�<-�d�8#�)�S�iX�|bW��쟴������a��s�����HF�*Ű��B�i���'��	�g%|��H|����1V;,9)E��m��	�p�$b��$���'^��'%��yZwA�Y��(B�yRd)�s�^�=����ٴ���9>���mZ����O�I�^~"kΌT����_&�@�x����M�)O��d�O>�$>�%?7M	{�Z�2�+�<7�@ا&�w�FL�=P)p7�O����Oh�)�n�i>�K���hB���,�V��y�/��M���?�����S��O2Ek'��(C�Pu{�mt�p�����������	�x��d���)-}�ŅV1@쉑��}�z|ӆ�U��#<�����O�	0=T� #jM"��5�P��$&"�d\�,Oxʓ��'U�̣��2|��U����)70�D�*p�1O�ī<�&�h�Ü�/b��p��"�f���fB���d�O���&��՟���f�D�ڱ�;=6�zQ ��#иnZ�&�hb�@��Zy2�'���֟�ro��ndॐw�	u��b�iX��'��O��D�<�dDަ���k}Z,�pf��yr^p���>����?y����-(�&>��H2,��m�
��M��@�@N;�MK�����4���d/��ۮKM�hK5��&/"�R�Nگ�M����?�,O��m
e����s��8���:E�
B?=������5�<���?�I~�Ӻ��*Ό8������<T������'�΍���j����O�B�OC��|\"��S��."=�s�h��($Z<m����۟��	����<�*���
 �
�d�ǌE�\����L���M����u����'s�'��$�>�4�TU����w�d���d�!l� ���U�	ǟ���m�)Γ�?a���))�DA��L�8(�NB��WO����'�"�'xL��b�4�4�p�����0֯##\(R�aըBB|y�5�tӠ�D�<�R�^�~��s�p��ܟ��	�.���sN�>8���)���% ��Q۴�?Q��:L�����'�bY��3�$��T�G�2L~����\��M���jm������4��$�<���!�rG%@-w݂��E�5C���C����O��>�I؟����n�������Oq8qSm����Q���>d���?���?9-Oȕq�R�|
A ��\��t#V��PE��OOŦ)�'��[�,���D��9!p��IT���I�l��8��Hq��l�2�4�?���?�����D�]lt5�O�Zc������(��o;Z(q�4�?Y)O��d�O�$�~z�|£�Y
d֦Q��$�|�Ӓ�D%�`XK��?A*OZ(�sDu��'[R�Oج9"b�=6�z2k����EϨ>���?9�;���'���}z�I�j��	w� ���lNʦ5�'���2uon�f���O������էu���G����t4�Ȩ3�M���?	v���<�H>I���g�T�M���BB  0�Q�M��d�4r���'B�'#��a�>!(O���E��t���@��4ޱ�/���q�w��'��<���	럈 � ԈP�Ö�e��G	�DJ��i~2�'b�$�H���d�O�I�?N^ �DJQ��()0�[1#��6-�O��3,tM�S�T�'_��'O^��遆#�v��vL��0�p-�Mk�"��]�~�'��I㟰�'�Zc��Up��(M�V���i��B*B�z�4uQ��#���<����?a�'�?����2<��YD�1�����B�%��Q`�^}BU�T�	`yR�'B�'�d� A	
H��(Y�B#��H֧��y��'���'D�'�副��U��OI���MőJtq'&�&c���ٴ���O��?1���?ɷ�W�<Y7������D$�x�Ssd¿i?���'�"�'?"]�@��
���)�Ok�["x��@/���F&�	�zT�ٴ�?�*ON���O ��̎��D�O,�I;&B	�2��!��!����פ6��O���<��#L{���|�I�?9u�R���l��,-��eR��˹��D�Ob��O���=O2��<!�O3�Ij���2: ��&G� lW�޴���G�{tlo�l��Ο���0����D1iA!�2Aa�ɋ7�F%4��L���i,2�'6�i1�'~p��<�����	/ذ�3$�h�[��M �Mk�J�)����'��'}��ʰ>.O8xٲ��K��ct�_��؄���R���d����۟�QB��_���b!b��E��0��f�s��T�XS�&�'���'�,����>1,O>�D��p�F���^����/>Tl��-{� ��<q�L�<�OH��'�R�^�&����֣ӄ,j͂�-��v�t7m�O����m}B_��	yR��5�`��3���r�X��I�2@����A�N�d�O����O��Į|�j��UL�8^��aK	-V�yQ�I�#��ILy��'T�	̟l��ҟpѦaM�JЍJE
��!f���d\7L����jy⊍-���'���+�:�؜O�P�$k�36�c1�;�#�4����Oʓ�?y���?y����<� 	��q�M�ŮOT��s�f���'�"�'j�\��cwF�����O�8�'�`Ɗ�q�K�yϖ�H���ߦ���Uy��'���'�2�'��s�>��g���7.��hŮ�
_%  �i���'��I��Td(��H���O��)�	~� HD�ɾJ�$�{T���a��9�'M2�'��Έ��yR�'��4����5=��*�#��
�N��HK��W�!H��M+���?!���z�^��ݗ9_�f�8:�9rEߘ`a�6��O��d��NJ�$�O����z��>�z��V�k��� �P�B0M�#nj�Db��Ӧ���ҟ��	�?b�O�ʓ�n`#�k�{����;s���ճi�i'��Ia�N�z��r���;�I�S�����S�XS��i���'���b2V�����OB�	&0%t!S��ײ�6�*� �c986m$��W�R��?��	���		]p0��3tb�$p����kC<�)ش�?���xm�I^yr�'��	ޟ�X�(��|0�	u&�Q�i��U6���
�Γ���O����O0�J+��bp��C�v�1 �6;�����*z���Cy�'���ß��	ȟc��>C�a1�T.6����@� ��Iwyr�'Z��'�剱OO��+�Or>����/�dB� �tg:�K�4����Ozʓ�?���?���_x}R���T�xm34�ډU)F<���M���?����?1+OƁ�e�j����56l+���[���'HM�2 ���M����d�O����O�ѻ6ON�'pf$�B�L�t�Js�S�|��ܴ�?�����о2�m�O��'����b8Q�ߞ$�b����*����?!��?�PG��<	/���?a�Rjݮ-_���e٫Cxb�B��h�H˓(��J&�i���'^��O1b�Ӻ���N�e�xݺQ
֦f`j��˦��I�dsP�i��I]y2�i�k�0AZD%���3��`�v-ӵH9�6m�O���O�)U}b^���'��lW�}g��\{����,�M�T��<�����,������": �;& �}�Rр���M���?Q�6�%�U���'��Ore�҆�Q�JݡE��+�f9*3�iR�'TA	�����O��d�O����"�!h22�i�v���P`�ئ��Iri8mc�O���?A.O���ƌ��p�7v졖�@�Q���V���F-`���	ȟx�	��y���5�<B֥М����qˁ����P3�3�D�O��D*�d�O���\�%.�m�e���_  K��O�EI�� �5Oʓ�?����?Q(O��0����|��T*�hh�*Z!�U��BKk}�'��|�'��["�78�a�1�(b�U T�꓊?)���?�(O@d�!f�C�G��a�T*��I�M7Hr�� �4�?�M>����?I����?�N����H
��`P����j����RhӤ��O0�("f`2��t�' ��I��m!TH���5J�J�VO���Od�ِ�O\�O�����1m�<��A��@(]-�6�<	�C$aɛ�`�~����ҡ�� AW.
ErVHwB^�Ln9�2*���d�O䜠r�IܧPH$-�t X9��!�CM�L�mک4���ش�?Y���?���`�'�bi���.�� ��=r�U#� mK$6-�%PC�$.��5�Sӟx�ԨE�-,�I�E���f�L;�Mk��?��~r��0�$�O�I�aE^qs�	�9eW$P!�nG�.�@6-(�� ~@�$>E��Οh�	�WU���Q&H0?�P9�/�Fk�T��4�?�$��V�O���7��Ƭ@	�d
�$����N�0/��e8�]�x:"�ܟt�'G��'j�U��� $(	�Fٟ8��Djq�M�[oJ�r�˒<o�'���'h�'���'��y���L?�$�J�n�'ָ	�]��	ӟ&?�X4K&��d 	�HtιI Ј\"�����ʍ���?II>y���?�p��?�i@3������* (�a�ߑc���ݟ��	��'�FP%n �Ќ2"P(����5� EB��'=���	S��쟨��=zE��	~����:$b��BF�����#�ȩL3�V�'IrP��XgGY��ħ�?a��#g��Y�`X�#nj^��ɥ�M��?�cK��?YI>�O��wAӈ\R�f�"&^�iܴ��D��
r��l����I�O��I�O~��7|#�i�v`[p�`{�+�'��d�<���ea��bU�|�СҥZ� �,!��M��d��GW���'C��'h�t��>Y*O����g��= �K�}��� ß��1K�|��I[y����O�б���5C�1Y��C���&�M����	��|�Ia��X2�O���?)�'ڒ������d
Q��,]��ش��Č7e��4@`3O���?I�	ğ���v�|��"��)��  ��F��M���>:���Q�ؖ'�T���i��A3�W,LӖE�F�A�_���p�B�>�m\�<���?���?�����d�f�N��$*��>���bC��:����Ky}�T� �	Sy��'��'��bX�Xs��!�m�EЦ��f[��y�W�T`�Yߟ,��^y�iؽd��瓅dȴ�2GU> V,]�����L6��<�����O����O���72O�Ira��G���B�+X!tT� ��
ܦ	�	ПH�	ן\�'A���°~�����)˫^���X0A9FM��a'�զ��	qyr�'`��'�4�қ'�"�O�H�ǥ��`r���2-�.�B�Aױi���'[�9�&u�������Od��sf*�HD?���u��7����'���'������<��O��#�� ���5��?u����ش��>?^�oZ��I�P�S>�����0�.S�;y���ũ�b~f��W�igb�'ta�'��'�q�nL#� O�O�@� r*]�lu��R�iB�\�V�|� ��OV�D��ڕ�>ѳ���.�4��E�2kwR���ďs��gT<a��O��$�O`0��C6��`֨ .�����Ҧ1�����I�dL2]XJ<!���?���&�f��)Q�\��a ���>�����dF	31O|���O���ʦ7* ] �~�>�`�G�MUL�l���X ���ē�?����?�)OkB�0Y�E�#MV��$���b
�I�hSc���	ߟ(��fy��őĶ5��#����a��)"�ܥP� ;�d�O����O~���D�1�v���E`<؉�A��,Y���{��p�� ԄV8w]D���T�S�r)p@�3D��s��:g��<g<:C�	�i��I��NF�B ��/�W�p���aŪW��l+�.�q<,�P6c� t~ܚ%jȳh�� ẗ́$�BDH`�?T��F�J�d8b�G�Rf9�3Ř\�J�ˉ>,Ē����7G�)��@�~��L���M�%K�cP�\��.�)[��Jݺ����|�Z�s1'�`R��
Tta����l�9�?�Ǝ�L��`�!Kλx��y���3�?���:l�$F� �N:�J�K�jҍ�?��O��|	T�Ҥ7�Vt�ʃ&Ik.�L��! Yz��+����vɛ���v��qO?]��
?=�)�צI����4}��M�?a���h�(���]P@xa��qP`���F�7<�!�䍯"�X �qEK)B.���!a�ax2�/�K�5J���^O��Pj�o�.	���i���'r,	�2~��i��'���'��w��`�BI�a��m`!���ꖌ��gIH �� 2�E[3�D��1��'9��5h]�~f;rč9�!"eEA	x�
��W�ڰG|$Ç�9¸��2״����_
�ν�������$ߜ{<�O�ў���;h��P�g��E��a�֭*D���v# -� �D�%��o{���I��HO�)�O�˓P�⩹0
���P
�T�A��ӂ�~�����?)���?�0��L���O��S�	��i`G��C8�-Q��7DR<(�g��1Vz :U�P�%���	"&�җ#��y���5NǱx {�S�zk�!�@#P�j㨀���r1����ɱK^`��e�1W��Q��L�T�4�O���=���'.jI#-�Q�H��5j��z,`x	���U�\A�p�؎K�|������R�
��<�i�"[�pV'��i�O�p(�W;C�j]p"��:���O\����~'����O��S�t�h��t�����]�'H��2c�V�
�����Oڌd�ɣ
�rR����A$Z��4�O�h ��$�{@'�[�1�'KR(����?�/O�8���̪�EW�����7|O��S�D�8R� ��%q�Fi gOPLl+zA�z��ƈR����aK���Ioy�iVSb�6-�O�ģ|�#M֒�?����yr�e(.�F�!���?������H�����DaD�FW�$BR$���4y`%#}���Ac����NZ��\���iW�R��rU��.\�0�I*��]"��	ԟ�bM|zI~�$�S+I�M��B=~�z�I�Kc��?�ϓh��1BQ�0�������ufj<�'�l4�yrms�R�d>�� d�i�#Я:�&$����vbzIʳ��)��ǟ��	8Q��H`�+��x�	П��i�Y��I$��D%���܁�U+��
�p�h��?�rI�Z�R\�|&���1�eX�y�e�c�8Pi$cR0(�șaգ�?��F^f�>�O�ES$T���&��Xd�Q�)9�ɼ}Xl���|�lE&{���FM�d� e2J���y��ނF�*\00����ŉ�������]b����|�ǅ(8]��Pb	�<JrC�+8������5)��'M��'Y��]ɟ��I�|��i�<V��nZN~2������u� �bS�y��Ý{Waz��F,�*�����a|B��5 QO�y	��P	n��9 �e�hd����#��]Ey��ܕ3�ά��J��LP|�(�c�!��(��?i��?!*O��g̓0���h1('֞H�GI�=gKP]��	i�	2/1堦�^�T�������'Vlb��ش�?y*OL�����e�I�L�����{���R&�=S�d˶'_���	�`������$�'X���	�	�-`�M��� { M��GD<a����dS9g�O�AZ'&��g�~Պp�w�L`y7d8O:-s��'��'<)�󯟲mQ�0��LB6')S�'b$K�,A H��!3�BR��Z�'��7��h�[��Ʋ]r�daٌTÂ�O�$���-������O�fy��'"���B%��1nA�%�O��q)��'4�l��T>�5���34 F�R¬�a�D�`��O
咀�)��@�1r�ʨW��$���ܿw
�'�B�i������O�M{���-�6��2�55�i��'C,x0_,~���r.O4-�p�@	�n��((E��:���+���12��p����M����?��g��9PQb��?y���?��Ӽ�� ����#ׯa�tYaJ�5n�'��@J�����
���#��uH6$J�\4H�d+sl݇;�<Z�� ����@~ܧ�� ��x����$p�
�LM+I�<��y��M+�?�}&�|�@�Jy�R�F�>�>]��:D�("dƟp�J|�$f��t[�Ⱥck.?3�)§u��e����]c,Ԑĩ&}�(�9u�� {�x����?1���?���b���O���unz1ʴ�	iy�qH�\)f6�p(e/;�,�w�^ �X����:D�vmY���"C�� �!����$�D�3 �)/Də���O*��$]2rpa���T8� ��U=(�!�$�&|����ڦ;�Bh����;h�1O���>A6j�0m��v�'b"���^]�4�6�/z�Њ���n>��'�>%��'U�5�F��u�'�'-�XRJ�>�2G $?�ܕs	Ǔv"l�?�A�6�F<��E8b�:�7OE8��;�d�O��Oxi�C@E�����L��
����"Or��҄�SX̚LD2*R���O�l�R��=ɐ�<nX%j��U�&8�c�;beY�M���?�)��4{�O�O�a�b�Qp�	�ʄ�/��Y�M�O
�Ě ���9�|�'涰	V.v���"ŎĿ�"�hN�҆1�S�'�Fm�ӯ�o��=�e�'|�j��O��{��'�1O��iOw,����m��1����"O�4�D��+b 	�qL�	`�ZE���'
�"=��jѢ4������t�b�i1N+���'@"�'&p�{��K�Ed��'�b�yw�WLY�Ê]�-�6���?c�Q��O�![��M欒�1O*�0�Np4tRʜ�ǔ-2P�֒Y���q�@���Q!ժ4�q�2L�O��Mɂh-f\Cc�@+C�Qji�O�$l̟`uH���>��?6$^�7�&�`nE"\�{G O#��=�M>9���Y|>���=���"�a~��bӲ�$+��|�.O*Ɂ�F��8i�ai�e�,�a�����O-�(B���O��$�O��$�ĺ[���?ɝO��Qh10�H� �Mn���J̊��y!c�_f�̅�	+"�P@��D�� |��D�UN:t���Kqh"�ђ�.�On�C3��,�J��BGB�M�e!5��c��t�TLl��X�'�"���D�Yy�(��d��`ˉ�bO!�k���0��=b0LPK[�EL1O��'w�	=��k]w���'��]�B��y���b�_Y�FU�D�'�¦�.���'��i�I r��0Sz��ů��c�8{Tõ":��&�"7@��`@j�'Kt�q�X�
|�J0!f��{��94��Xq� �7�r����WG�#?wǊǟ��I۟��I��@��.a�ڱ��@>$�t�'�B��S-a����"|�ԙ�#�V#<	��4��Lo�7~N�[W�O�;�f�1�U)w�dx�Igyn�~��7��O��d�|j����?� ���3�'?�ðo%i���u"�O��.6��ɣ``æ{HzM�<�M�O}�S*/�65��CN��ak��J�+�'i����5Ƅ)v�V6��|"�L,��	�7yh�(��!{�So�2�c�J���O̒�f�䆜%�E[����)z�*D��@�P��O��$�O*��D0V.� v`��~Q������ax��;�l���Y���%њU�dC[�pBH�f�i�R�'�r�V�(H�s�'���'7��~�5�T$��
7��J��Ȕ#5�qc��*_,�as��R?�F!#]*�-a��L>�3�I���X�`F�X��`���Ȁ�/"a�6�Y=&���ˉ�L>�%�Ԙ?���X��
:X�I�UO�$+���'iG�2I��OhB�'6��'�¦E,̒d�Q�)F�T�c���Mu��d�#>��]�G��5C �eO(^��I��HO�in؟��'	�TbN� �U���3t�@}ۆ/DV�!�'2�'�Bnnݹ��ğLϧyu~��'��h����!�HF�U�'D�0L��ܨ����aɚO �R�g�01��b�KG4s�N�� �rx����H�=�M!��7�J��%^�n���O����O���?������3��ORV=�A,��y��aF2��5B /�9�ݨ��'�J��hO��S ����e�ݓ�@�XI!���PL���/zRH��m��L1!�ݠs��t��=Zh����!��Ç<o�kvj��&S�u`e��>::!�МWB^�8S��+�bbCl	'w !�ʻq�� fb(��Bb^-!�Y#K�l���AD'l����Rn1c�!�D�(f����C<P�e��fΒ,�!�d�t̰%h�58�*ɢwhL�*�!�D�x��Q�֮ΌP��D��U�!��X�E%��$�9d�H��ɗ6U�!�	 A�����J�DH�Y�X3�!��3Ԥ��A���)+������c�!��֝0B�huO^�Y*������!�d̀D����՚]!�m*ѯX<�!�d�)b�be�J�fp@�ѳ�݊B3!򤐴�Jh�bD֚L�0�+$h�	%�!�$y�PD���C3_�A�F�ב5�!�	'�dP��H���K��#~!��[x���CX%�ցJ��� T!�䃊R� 	A�A#S��X�b��]!�d�W~.6�Q= ����	l�!�D�y]�A"���W�쀳t�[�!�dD�'^���,�F���a"l!�$� �RGM�i�d`�-CS!�D�{`tU,ٝT�2)�bmėJ�!���\BB(Yp+H�
���j�L��W�!�\0ـiKf I����	P�!�ҡX�9��j�� ��t�� �S#!�S(T����'`�Q!�Q5�!��1IwD�JwD
^����F�+H�!�$�J�dbWcA�;��Y��� �!�DZ!_��XAE�؞f�xM��-�!�R�Sy����ˏB�F����y�!�$�,�l]���>x�nT��R�T�!򄇚0X$h7΀��ГF٠!�!�$A����B߃A�d���I�W�!�$��2&����`:n�qE��5�!�$�N�YZ�ď�_L�ա�LD�%�!��L:V����2g�b������!��^�1��E�ED��C������D�u�!��_$�a픾�(�)�e�*�!�̹\�f�z�o-T�<�a2'�4B�!�֡8�4���IɆC�DpI�D!s�D��6���=�Lݘ���
0��@R��a4џr�c����� P<C�)�4���B��W�A�p��B�!!�$D�l��*b�D�:��%[	副!�l�|�\%
`0�g�? ��4bPH]r��5A�x� "Ot0
PǊ �x�{��ɈP��R�N�@��	b�'7��H%:O�ϸ'���h�̙j�xPC�I����]���(����n���ł/{b�($�@��y"�V.�,���	O�z]�0ŖE�Ųǡ��x�?�����y��z.B���U���bL8B�$�v&�-׸�ȓlM����̒̔�e� �;��y�'C^�7O�e��%K3����YٳA�:ފE���H�o,]�"OP0��<.�HA�_Y��yR
#Z�Z���'�>؊���Ϙ'���cH�i9��k�h�"D>���'>pEk)@:�X$c��V���P��'�A5�UR8���S��I�}�T�Y�)xhdrq�6�OL�G+���~�4P� D�&�`�U۰'N��y�ˢk

��0-�6h������)���	`������?�� U�t�6a���B��٠D)�O,}�m�&e���dAdr3$H�!%�@��G�rF��Q��������I(�����.K��ke�O�O�@ۅ�Û[�&�ʦ�;�'��P"�o��rҼH2��Q}�e�	r}6�)#śD�{U$�H9JAK�+"����G獑�ґ����T?��z�O?!pDc�|����11�ҿ,��g�%ynB��0.Rm`�̖�Y��鷃�&V�&m�&fIl8*�M��>;�aydj�?�'��25=���=RH�3�(ֻ~�摄��>i$ИK�M�/sH�����%r�>)y��
4��튱�_�&] �惲�n��OTLD��O�����Li���Rþ��C�
�C���G�ܰ*;JQ#��Ɇ�(�~����H�y����D�P�KlH��GO�����YY�'���Ċ�<�Eʘ 00\��N�6ze�B)�/$�(���'j���6
	|�I>�d�K=2�'E���vL tp�v�=LiR�S�)L�z"~O��a������5���#vަeN��cIM�GpYwfO"7�lX��'��z�X>��!��'R��`q�fD�.Ҹ��d!R��`E���F��9��~�)�i϶ !��(,�a�Q��>&�	+
%w�Up�K�^���d*��R ����o�""|�'���YD���Yh
@�� ��X���ߟ��������4�;!��������O�7�G���Ա�n@qY�˙[�~�x�F]=+��!�r��(OPPe��[}�Z�j�`)0�ܡCJ�lP oMy��Ԫ���F��8�Er�Փ�O�@i�'�6�ԟ�q:��V�]3��A�+���4���0�p8����|;����lO�/�X<�$N^ *�3+�:hL�e������:��Y��'O4���O�B��&�qfϖ���b7�
�ax2��w�r1G�Y/Pa�)R$,4���=%h@cs��1Y�	{B��M��l-�~���g�����O\MQD%�-w4��K�`�	ư����p��`ЪW�,�c1/��i
�����Oq����v�QCG��*֌�%��[�H:.�d2p���"M�0�ד���Z����Q���O�!�����.�)�f�ȟ�� � `�,OD]�W��\e35��mR&ԉ����8|t(/�d11��s�}���5�
p��M������>1_n�:C�T���d�{���O8�������8������Z�P��1�.�p4���/o� �BޯQ�6qۂ�I<:���b��Y6jmR���@��Np�K�O�d��.�|������t����O��gR"{Tx�"�d��`1�B�����ʶ��,�:ŀ�4}ء�S�'-�N�9r�'"����&�t����f��c� x�$
N�o���D�5J��X��]!T�)RˎJ��Y�`�ߨ���E�'e��`�?�S�d�K2z�&�##��������w�!�[:D����0-����S�T �h�.���%A  I�IB��'��
hj�.D=s�y*dΖ�4����@]��g�C36T��p����5p��KA�D=2�&dZ��+��$ $���!��O\�z$T����� M�2m� C�p2e���X�Dx�I�zad-�2E��|	���M�Mt ����ln�Z��C!�8L��o,DGN�����588�F��$�p=�lI������� �J��T��-!N��dc����������?�I2 ^9j���6��
}X��c�@�P�Е��Aqʌ@�@)��)�1����6K�*`9�`d�Xs�����Ofi�D���F!�Ah%ez�=�7��x�}KB����4X�4��%T,&|��I�f���'(Hm����}G\4��D'Lh�$ɶ&ơV�h���-xZU��Zr?Q�H��c��l�ע�򙟨����%=|�hpi�-n���w*�*n0|]R����*�l|S���8�bb�]y�K�^�:��䙳�fٚע�">T)で��AϞ8yef�M�ϻ.K�9� ']
EV>�y�@�?pRA�<aB	�vA����C��b��'g\n��fI$h���ȳ��T�,����e���f+�.f�@e�2�
�4�Ur7o�5�#����ذ�1�P7S���#�Q3���4��Ir��'���C2ر�5�H7s�̘4OF(jJ��ٖ��y���BV�!?�%8Es�T9������HEE�~�I5G�&̑� @�l Da �"Hr�x��i�!�,4"���Db"X ��g�0RHBA�?�p�W�(����BR5q?.�s��ЙL�l��"<�$T�O���wU<�\I� �ϵQn;�톟Za��	AH�1%��]�	%�d��PtQFAȥa��y�w1�8Cf��t`<	��2J��q�'�(�A��X� <Q��+��8!�E��<�Oۜ i�b�$+&:�Z#��q�K�l�X3�a�:Q��O�L�b��!(���4'E)[n�b�L�Ɗ����*`3�ʓ��	ϕ5 �
'm�-�씪�@!^�i�F�2w���5�Aʲ�X�O���c�)d�">�fk��$�������.�<(���N�z.��A�J��J����p͋��l���J?T(��]
>":]���ª<:���Ko�$I�U,�9Iў$��"�p���Ki����kF��?9roI%W����L{E���IX�cw�Up��xO@�S��yǥ۱^��C�V1g�,�?�!(܈H0u���q3F̓ǡ�a~��#C��S�ڢ@�I+A7r�Y��b(� E͏M,���iD�L֤-`CE�Y�HEHߡu�T�fI2���M�O���хD��ZiT�V|MH�cU��*��fgפ$7J��^���P��{;&$�U�>�{��(7>&%�Af��F.@ �*�����ҷ+�6�}����
_�ם��@Ο���#|��0����f80L��Q$vd��'M�'��qeGEMp�IDy��ƐE,�|������oѕT�j[���'N:����iJM�'�R��p��ܘA-](D����=t����,*iB 0�'� С���$�h��g)I�Pʴ�	%��!�A�~��	 �M�)ʀ'2LH�v�\�$b��b�D�gx�H�r�L�d���`�L��/�z'���)"�+�(BN��V��C}�H���q��G�Py2M4��ʻGod���/T��r�2���_�$��T�C��g$��P�S!{B4��$�	SK�y�=�#f]����#^Hi%ځDR$���o�5�v}Bg�	'wB(�6�F-hV$����7"�Qrv/��/�nՀbM��{`џ�Z�w�DI��!_	R��ֹ/��m�'��d@�B���Pq	 %X>V�s����t�+f��Z�' Q��kU���kDP���ɬ,��y�!ҩB�� J��/=����$�H��
}_����J��P�ٖ!D#>��@!�Ǳj�h�	�-�BU2��,T�|���	!:8(�.$�a���ҙ$HX�tE�g�2�"��}�8�Kƈ��@u: �d*`���"�I�(r( ����].���QAT O��U�&� YȨ����������A[j�W��Y.]K��Z�ب[0�W":m����)ۅ+)=�d�&=Ph�3
ƭ#d�!��-+\O����	�r �A�r,�q���"�@��?��a �O�'�&}3��D�d���oCL$��z�Ä/F�dS�0z�,��Ќaj����'PXqO|�0�*(����Sg$f�T�V.g�8����[8}�je{b/�!F 9�M�&g�:�"�'vr Fh�X�lpҢr7jވOT @�U��F�b��� N�y�pE"$�P4�d���=�-�If�,�+M�<
�s�C���!a6��R&M>�0?)�-ܻ	_����� _#ne��/رR\¼���'q�9�w5DP玾z>~E�s- )d�����$:���PKg�bJy8%���;E�h������LB(�)�D;8r� p�ğ�+��=e��M1z��v��'Bcў��c���y�Cb�(��γ��BU��������R%�`��d;/K
�Z E<؂����b���ΩAL�M�r��yYvy�4�i����i�p��m�
S����F�I8�DQ4	�qU"9��RLnu�'pqO&�*M�ğT��@V~"Ț%7�)�J]i��Y���hSv�!�O���Rb��YK��J�$� �B�Ȫh�m���)҆�i$�O0�i���v��,cd�+ƉX�eT%�$>���rƌ"}�ؼy����&�ЇA��<��(�S��{̓|�ɓ%O��j1�L��˓�8��a�P|:��GMV O�=��ɕH@���)�*2xh���-Z�XU�ѷqe��ģ��E}ȈˤOP�űO2�Ór����2��7�DZÏ��|�'�n͋�"�?g��<�PF�S�f��S�'B6&��+��v��U�Ԧ˖I��n�d(<���og&\��f�0wOZ	� CR	{A
�rnҵK�v	��L�$��|r�%}"i>>��B�!�*�x��Y�Px��#D�X�T�=���3�	�7)�U@����ž��+��~S��x��'���ҨI琀�ph������'��$3���?T:	�jݒ{��)b�'b�{�Ɉ�J)"�8�b	c��r�'N^-c��_Ƕ�0de��k��K
�'1���(���C�;2��s
�'�L��R�*��X`�0��I��'����6�XǯW�.?�-��'چ8����<*DD�3&Ȓ����C�'���b-�O��[%�+��p��� ,����:*��Xs k	�IV,��"O@Hz��B�}v�%
'��q�X��"O��a쀾yXr��T��:6���0s"O�]¡A�%ߎ(��.\����%"O��	7�g�0�pG#?'kz��"O�x!d�[Y<~�(e��7U~�xF*O��1�"��O��%�W�۪-}&P	�'���K7��=A0�;�,��T�T�K�'��p���L�7`r�c֢ݗH�0�[
�'Y^��N�)y�Dp�Ē&=�d$Z
�'�lm��
�,r�HmX7b^D[�!
�'�j0����3s�E��e5:�:�j�'���"��V>4?ZEKg�*�2��'`�=bH�!t�|$H�.��c�'rT�bŪF1v��l�� *����'��U3ՃќIr��P���
T��'��L�S��&w(�@�]]<� ��'|`����36��p`�[�)�~��ȓF�t1S��ƉW�0@��F�
���d$Q�KD4	�x��ؐD�� ����H��� O��KP傊E<5�ȓ1�HC&�C�;�B��H��
0Jh�ȓh�f0J�'ɺQJ�k�L_8jC"ņ�[Τ%�L�)\��Q72�q��]d:(86ϟG�$��d*^� �Δ�ȓ[I�!�3BR�c� c�M�0O��U��&�ֵ��BX/D%@A�[�r(�ȓ"`� Cƀ�F����Ў�K�bT�ȓ7����%I��fPk�`K�z�j,�ȓoZ6��$ɸ^u*��b� �^�<Q�@�%u����`m+2�V�*�LY�<1��Æ��MY`���
DY�&�S�<$�A���k#��c��H��.VP�<�a�Mf ��bH �U.r�`��L�<!��		U(T��ODM�%h�G�n�<��VnM��N@t0�����f�<I��LK$ �i��3���Be�<�7��+t+怃�N�:�~�*�f�]�<q���i���C�J���FV�<�։��Q�tp��اv`$�P���Q�<�@f��=�5 �B1����cIM�<i� Ѻ7kʝ��#�%���(��Q�<#d͔n����k�UF���q�AQ�<��FF�/Hꔢd��A�j���\f�<�00�fӁI^��P�B�el��@70]�� ��b��l��J--?n���5���P��:�XP�D�,-XzL�ȓrz�z�E��21�1�0`+d��W�F�c�3���+0f�<�xh�ȓ����CM�2��A�L5�1�ȓ9�r!*uk.T.ekԏa	�i��l�D� K���Q3��	`�E�ȓ4���P��F�i���(�)��T�~����8n����Yq��ȓ=�⡚F�շ�� �\�|Lj8��cҴq�c�8t�(�xC������ȓ4��E뷪�5sE���э]�
��؇ȓz%�Bq���|ք1��TEN���N`*���獙z��X�c�G$��Q�ȓ:�FtR���yT��5��G���ȓ>��c����a�d(�rn|�ȓ?�� �ũ� e�(ĭ~�c4�(D�Z�bL.[R���n3=���� 3D� ����gB�2�*��Y���¯.D�� ����I�e��M ���g��a�"O�TbR��6JN�0��*i��d����O�O�&�A��,"�l���Q w��Y	�'�ĩz��hD� ��ω�X���O|Dz��)ߏ=(��2����Qse�&q�!�$�{�<��%	KP�D?��'ea|��
[� HF��$,��pid����?���w�2�CV����d1q% �|.Ei�"O��r��U�=�A��$b2I��'�ў�		S'h�� �PA��/�]�RC:D����V"-����"��oGx�@�g*D��!"����R��F�jr�j'D��j OG�+��,� o�,�D���'D�tt)��������Z�<�Y��8D��Se�,���뢂7x�2�9��5D���V��Q JIK��)j��m D����Y��xD��ۻ''�xc�9D��Zw��&p�aX�P�
�`e9D��{�J��li�Tm\��j��4D����QKb�C [o�6�3D����H<ޔJ�[!Y v�z�/D�4��Ѧb8@6&	�Q�x��]]�<iP�&E�@��+��4X\�B'o]�<�����}@V���dU>YqY�<���s�Vla7�@&8,�@3�o�<���	*������N!"!B�)�l�<9�mD�P�`8�e�S�U��DAU��h�<�p*G�j\T3�=�΍�a	b�<!��D�Q��t��;n\na���Wc�<���ța
����G�8_gZ!!Q%]`�<�S蟲%6
��w�ɿ9�	y��^��0�<!�b��$$B$�@H� �0X���[�<���<,9~��DQ-p@��U�<3dƌ/�JU�P����XBEP�<���N&lPrΒ�a�≰�`�I�<�"'�.&��#���eI�����A�<d �'K9�Ǟ ���z�<a�QVn�5%�m�=0QKb�<	��L�QZ^a����2��d�P`�<y�䋎^�Y��ʈ�;E&�(�iQ\�<�Q�֦"u�(�6b�g���g�V�<A�*�O�������d ��N�<����u�����Ϸ�1�#`�<iB
 @:��"�ƵTtڷ�Z�<ӃM�֘�&��0}Wh�7�P�<���( r�Y�%��79vU)d�XK�<�6cT�\���2���>��� ä�n�<AQF�Z���S��.Rc��a�Dj�<��bؼw�)���\(�tM#% Z��4�?����&�p@��Y�,��F��z�<����'�������:���j�J�<��cӂ�Z�K�*�]�4��pBG�<a�N@v�`���VJ���3�E�<q�`I-&Z�@�c��a:6EVX�<����L�iY5AW�E(��Db�P�<gIG8zD��C��=��Q3�PT�<DJ�1-ʤ�M�.G"1�Dx�<��aʳTJb��f'��D@�l�<�,J�5a���@.Y�u�� �ǉb�<	D#��B8����c�"
��,PBn�Z�<��ȊH@.T��d@,���P�<��/���!�8C�U���f�<ɀ���w�m�Am�3J6�	��e�<�2��5	�l�$M�x�Aa�<� �"¤
+*~��g�`����x��'�r|Y�L�*M_l@�%�)r�x!��'� ]`�
ܦ_F>;�LT��I�	�'<����*~� �	ԧB?������y"[*�"<*��U� V�a�ѹ�y�+�ϾqB����&�(������6�O���U�:J(�Vh�,�zА7"OT�XD섛%��+������ �"Ol���^!%�$�c�*��yp�"OJ�ʤ�
��n����_F�В�"O��R�d>Y��@�xS^��"O��%�ݠURT��#%P��Pp"Oh(Z!��)�D���dF:2<p$�u"O���F���ЛVCe/�$!�"O�̊S�Ehzx�U"�={$N}H�"O�eɢ)�7h�$�S���.�!�"O�b�&��y%�՝z���"O�`E%�?�`y��$�4А)��"O<͡Dlձ:���7�̔]�~�w"OB�q�	�����Ǭ́@y�0F"O���C*w�b-�qN�	�r��"Ot�[�` �;���C8I�,��T���D{���� H�&����n�5Z$�R7X�!�d�e��g�:OV�����9���<ߓ;�l�g %����
֐fr��>������*��!�"c]�ܶ|�脜�yB&�2�!���I!Q�Ġ���	�y��S�~h�+�fT���y�d*�}J� ��Z�!	��y�J]c��B�-a��Z5l�'�yZZj��RJL�":pi�R���K%���ȓ����t��wFFum����wV8��E��J�d������C6H���y�"5�a��5d��y3@�^�w6�9�ȓ2�pRꍞ&)~	�7���u��3����?�������8\�8��ipnE��%B;x��`@��Hm�ȓYHr��NM����ᖥ^)iR�8���Bq5��;_
!�`§qf,���$Y����ÿ/����7Kۋ|�h��>5&	;�N�/m���i@�����ȓ6��(�Ս	�t(QcS�ɄȓJӊ��ցF��yy׃� ��D�ȓV$�(�ܚ6uH�hf�
�ͦx�ȓ[�liRG@s�xX��˜'f2��ȓ��!�ѩ�]�DHT㓞 �6m�ȓM�^���KF��E14$ii�x���n�2r�t�<A�R���H>bp��f���(s��Ȧ��5`0��ȓ'��uri�UX�PA�H������M���+M�a�  $"p��$M�<��Ǒ��lyr��T"Mj81��MQT�<���9|m�@�*M�%Z�<	r�� ]�	�{�|i��Qy��)ʧ5B�=�ҥ��x5b6��u��M����F�yl�@�A/k4Bp	�L�<��*�����J>c�2�A�a�<�䅛�t��=����/ �4����R�<	��X�xXhA犑�W���vN�J�<quc�.g���֡�\Ij�F�<��G�v5��;��ҝ�<U��"�j�<�*N�-�*��rĪ$�L@�<�0�[o��ܒ�W!�1膊�x�<as�H�&���S"�L�[�b�{�<� ��+BOJ���+g �tJ�"O���[�<��-"�̸dt�t"O�ke�ߦ\P�k�%��gLȠrP"O�A-E��Y�m��{4f$yG"O�ѨF��7Q��l�$LR�vL Ț@"O^��m�5 Id��J]8;�h��q"OziUD=h�x؁g
�hά��"O��9C��1cg�੠	�.�P&"O  @�fʘ:�Ne�KD�C�L�T"Oz�C-`��1���R.�ҍ�b"O�Y ��$U ,ء��4Du��`"O���&��$@��P��ω�xgt} c"OIB! P%��4Yr3 �j3"O�hIĎf�p�I��7@�PC�"OpLP�'� A�p��k��,�.%��"O
ذ�?`�듨8���s0"O��9���J�\!�
�Ql�as"O��������!��p�P��"�!򄗛Q�V��cgɅ w��G�b�!��2&�r�cB%˙Z�L�l	*Q�!�6l���'hƹc��t��W�!�D����-��W�T��fd�!&!��� =��(�&Y�d�¨;��Ҙs!�d� A4�#2��8ÐIQ�k�+	!�d�"�`�Э��1	Qk2~�!��W^���BϗmH�qª�h�!�D�56\�ҳf� bM�����B�!�D�mg1�D-I�C1��'J��!Z!��-��YæN�w�RlYň�?.�!���F��\��煆\��aҌ�i�!�#2�|����Y�m�J���]9@T!��)"Ҟ��* (3����QOM;]7!�DM< 3��pS ��J�ٷ�M
)!��Ā�<��,3T�̱�l��!�$yB��a�C?��P�P���!�D�u�x�%��i~Z�tJU�c�!��w�������Mt^݃6)7O�!��ʪX�N���͑��Td!&I�}5!�DO& E�tt)O�~����M�J.!�M�gwyR�ՠmX��AG��Z�!򤛕A�,��A�1n;�DZPFg�!�DѼ����T��h\)y��v�!��ʲV<�1�B�K���i��ʺ[�!�$��'4�@�  �>Y�4�(��*8�!�DђI��(���?��8+�R�!��_z�ZbB��G���s�ҵM�!�D��`i�C�G�omҍ�C��b�!�dD -��H`��F�vg:]�E%D�v�!�$��,�3�@@�&��qb���Z�!�Y���p�*�� w����(0�!���*�QI��y���h��:n�!�D��y��I:���t���8rkV�V�!�^8�4a�I�<Zjf�"�D5�!�d��d����B��F�̴�a���v!�D�]l%��lx�I�	�R�!��Ş`��81�S&W���'�ÞVq!�P\��$�8dD�p��%gR!��"Nlj�g�/ZN8���Q�DC!�U�t:�������t!�$B!�ă�i��8�$��Y�搣A!��"=I.OX��f�ӵ!��	m`���S����v�$!�V#-��e���W%)�4P�$�P2t�!�$�"a��1Ҕ&�#.���C$��E�!�� bXY��;M�-��F�B�iE"O�i�r(��-`����T�ī�"O�-�e��'��AS��4!C�1"O����gS��2��BXa�A"Ov�&�R�6>�U���ƇEŤ��"O ��dK�JN��腠�F��"Op4(@�O
?�9Ȅ�W5oH"���"Ob��i(|x�"��G�~8��2"O�A���8&`%��MF+'Xx�"O��Cp�/�@�� �ؘ����!"O����c��v��[��!f���[�"O��J�"�Q�@����(R�"O��ȑ���3'6D��O��w����6"O(��r,��Gp�u��wɂ�`4"O:m���IA}��z j��1#��J�"O��؁��P��A��I�
7�h1�"O�=9G'֟)R�p ��V�.�0p�G"O�裑��M]b��F@	�gX Ö"O�� �!T�1��O����"O腒ԂG��e���\ -�D��5"O}�cO�֠�A� ���"O|0&��Pj ��c�ķ��
1"O�5�`����h�'�ܼF�0��"O�QcT�J'?�Mr��*
�h��"O��(���1:`�l�r�R�i�Z��"O���&�A=)k�P�+��g�\E�"OP�D#��]vq��j�'lBMv"O�xg�/ugĈ)E�3!C�t��"O(1cUDȳZo�i0�^��ґ"O��1� o<r��$B؟;�Ni��"Otx1v ԝ"�n���k�͠�r�"O��*��
�`BLZ��t���"O ����'&��D�r¿2����"O~�X�*�P3���E��T��"O
����$_�hԱ"�Wo����"O���� ���{Sa,q�:`0�"O��Zub��U�����͕ݒ�!B"Ojѣp�H����!@�>,��X�"O�("�C5mE�w X�B)N��p"O����-�|�b�O�n-B���"O����ȅT*�bC�D9�d"OB����[�z.p`���;�P Y�"O����bK�_ے@sb�<+�H��"O��É��u3��� �="x:�"O���g-�n�8�I��l\}�!"Of�fF�,'�0�8�����Q�"O��C5�	'5��z��1u�0]�e"O8��L��*��<#�K���u"On�jJ�CdbHv��� ٲ�"O�9���	1q2o�s&\��"O���� ���k֮W�E&�`A�"O�\zT�1v�d(ۤ�	mh0��"O�I�v'K�:�� K�&��ah"OJ(��,N�?�#3J�����"O0�Yf�	nLD9y�
�3
��]1�"O� V��)f�jI�N��d"O�*wĖZ��!�da?�0�b""Ohi���K6�l�5f�S�@q �"O[�mX�{[��i�L��"O@H�d��
7�ڴ���|C�"O` �mTk�h�$��3GӺȊ"O��A���u,�� �S�)Y��J�"Ox�Jq!T�.��D?|��IV"O���A��b�CS̍/7��Ճs"O� �q��Ö�zCZ�:w���ӂ�J�"O.Ph�F�?v&p���M=# <�s"O�M���_�QV�|#)�-]l��"O���� �4����B��j�F��"OP#®ނj<�	"��[!b�T�c"O��W��!.�ؤ�I=2]*qi"O��5W�^��d�� H�h��"O�$��@7��L;�nB�.��ѣ�"Ox��E�U��Ǝ#��,)G�	��y�C�/%e���(%������y�F��4{�p3�]�%���A�$�y"�ӬkB%�AQ)�Ùo��C�I'|bБ#��m�*1��Õb�nC䉝� �b��f�Z8�7kA�f�.C�	X�aȡ���N���CXB�I?|����yf�ɓ�oYJ��Q�ȓ�$tC�/�������+� w� L�� <���W
� ;�b5��b��0���_@J�	�,�py�V�.x�H\�ȓ �qz�/D�PX�8�$��D^��'&a~RBg�!�WN� [�ԉq�5�yr�+��۵�;NԄ�3�Ŋ�yb�د+R�Ặ�AM������y�S�P��i���D���ӥҽ�y2Ĭ ~eA񥀽F�:�y��yB��[�>u�B9�rE�r�^��yҥ�^�p(��[6 hR�� ��9�?)���;�'�x�I�㐬bH�Pc�z]v@�ȓp��S�g̑s DĀA!���u�<�$兏1;���V��.��$��\t�<����E����	�y9����s�<��@J|���R3�T�8�(��q�<y���B��t3�\�h�Hl(%��k�<IeE�y_Ԅ!r'@�y�ȱ# bXf�<���X�UL<����$a/eC䉁j��8!3�§Cǈd�v��<C��l�����ל_�,U2����|dVC��+1��\z"ؚa, �5�>C�I�T~9)'���3�<��"GϺ8ғO��=�}rG^;f��I�*+���y� \@�<�I3s��ɢ��_��
�R�g�{���<A �
�e!���󇀊5�px���H]�<�p�8�@��ҊY�|2��F\�<�G�)o�"��AĒDp�I���b�<��C��7�^�Au�@62��yE�F�<�!&R�)f\HC!�ؘ
<���x���hO�'}�&Y���-���@�mY ��ȓ,)<<�D�_�Y*����dےۖ���ɟ\�'�mZu�	:�� �3ت
��� �'&�ȱ��%	$͚��q.u;�'�$M��C�T*4�#�He�f�i�'[�AiS$��7t�[�a��d��<c	�'�4���z��d+����[��Gx2�)��F��>�@���Ψ/Qt��D��y��5vxL*��7!'��pt 
�y�+�F�*q�3��7.�������y���<Nj9ضY^��@hЦ�
�y��*��	W(�?��L�N��y��Qv�$H1͙ �XلE��yҤ�7<�:q�s��5!�z@�2K��)��Y�O^f�zw`G�*�t"�kM�%��j�'cN�XF*�)D��5a'�)6"�rV"O��rC�̍z�!;p�N�h�t���"OL�X��؎D�(�aN|С��"O� N�PfՃo)P����Wa��"OD�����*�$u{�,�,O��Kg"O═�f�-���b�oE����Iu>�)��¼qBDM��"�0Np��3�$D�|9�d_����+@g	� F�r'?D� ���>c��Q(�jCA3r��);D��[�-nI8;�M@��&�r��8D��8� �2�~�c&nڲ��i7D�\І�Ӛ{�l ٔ�Y6m���g�?D��劝$*�:QV�5k�"�I��)D�x�%^	b�Ѕ��  �V*s'D���/�!r*�U����.$�4�#D�(��CȹIS�,�S王mw�)C@�<���<9��ԟRE%�L����A�M4a�d�07"O$E.I8N>ūE�Ҡ|�~q�"Oڸ��_!<�y��9`[��!6"O ��M��~^v��-�?Jtb���"O20ص!��2M��R?t�X��T"O���#�"r��tc@�o��l�6"O^���Y	:�E �����z�Z� ��I&D�$�)�P�qZ"Eq�M+�*C��&%`���}��� n��R"C䉧IJBi�p��#e�H���9�C��~tH)��*=���F���=y�w[�� ��կTq�3���*����	ퟤ�<� ܁���Aef@�8q:�!��j�<����,>��A*�c��|�B��d�Ta�<	S�\9y�	�2�7?���	s#�Y�<�QAśXY��釺"%Ɣ��\�<�LG\��
@�`=�I0�A`�<1U�N�S�`8 6�L�yf%ɂ_X�<Qse��-�!��݈-��y�2��R�'E��'�B�)�MB�9�íin���Y<<!�ͷ����%���[ ���	Y07!�h��6L�>�@i�(D&!򤘦5��AIև��%
1�j�!�DǠ& ����i<y�XLڅ��?{�!�ě�g�l�Z# N�z ����!��]�}����4�t�!d��[��|B�'�"�'ɧ����(A���P�C�z6��Q�4�yª޹~�j��DœfK�XiF���y���ީ�5��<qYj�0F���y���	*�,I�C�
:r��8G��y�J�=y�glԢo*�{�MN-�y�aY��a�$0zK���Ѕ� \�ËF�(�M��E1+J���W�".66��2{�x��E�%�F�և)V�!N/ ��P�ȓvU�IE
C�� ��B�+	8��'0(x���5N����+v�����n�譳���Q��`(҂�"'����ȓd�s���}	��+��T�c�A%����b���'�`���N��HM
=���V�9T�0	�'�Z�J���?�d�c�F_�Ļ�'�4A!��@���#۳U����'\{3-��>�����Sa�e��'[(����ǒb�`$0$�A�D���#�'Q����L�Ѐ
�ӏ/<Z!��'g�Xٕ᙮.�*a�S��+����'x�h"��-Z�2ĚcM����'��eJ��B�W�	0���H����'+�m
��Q	�M� O6�)y.Ol��$�>{�٪�ω�%�V��J�� �!�$�u����+�3O�x)7I���!�� �a��I%g�ʠd+��(�E"Ot���>,��{1] @}<�i��'�R\�������I>=����Ά��-��F��L�rC�	,b�L��&{�ɂH�?s`C�	����Ā]��YS���RA>C�I�J���
��U�9��T�F��|:C�I$r�@&���ڰx�D�"C�	_�tdq%���$YDLU�u�B�	
�B) �F�hHz� ��ҿ���OT�=�}R���%��qH4��	�\�'5a�!�?qH ��F�u��=y#c��yR�7gJ��-, vpP�r��$�y"O�.z;�B�����T�Jc�y��Y��L*�O���i�b)��yJ�?��/.�d�Ql���x�d�#��:PC0�|e3���:"!�$YjǞL褃ۍ*ߒՑ���!�d��K!	#�ʀO�KV�]�!����s���^��u��݋O|!�$�1�N�4΅�;�<���A΢Q�!��EE��q��ƃz����/U�_v!��Q7U�<°m֣9�r�����G�!�$�T� [��Ȫ��IC$ ��G�ў|�቉@�X�H `�^r�铠4�B�ɰt���6�T7�IEЏLh�B�
zyB�i���}rlV��B䉆����2m��#d��@�X�*C䉡\�@��G�� ��vk=iF�B�I�Z5���/�3b[���M��+~�B�I�a�pX����r$���ï�J��B�'���?Z`y	�m*�B�I%s��4)�
 F�z�D)�CfB�I�Is�X�C��/\:�k�`��2�nC�ɿ'�R��瑲j{ظ7�V		n�B�ɩo�8�ѭ�=���faUzfB�W{�	agX5@�hDY �*��B�I\8�3`�5e`�Y5��n3�B䉝IN���=���;���c��C�I�r$��K
utHх�"=!�C�ɏ2���z��ȡMcj�@�g#qy�C�ɂ���v��s�L���GR�Y�.B�ɀT�h�"��&�XuʲIN.c"�C�ɇn��,0���,a"�$�(ki�B�pn�EbM!���5	�<�&⟘D{J?�ƍQ�zFPE)��0A6 J�!D�r��]*s�BY �O�h�0�ql3D��� mB�p���0��j����;D��r��3N�I��
mm����
9D��2]&��� 7��?>f�8"gh,D�J$kD.5���Zի��XW��r@?D�� �S�xq8,��$�%k">@f#?D�̒�ː�3��i�Vmʵ�̪(<D�X��!�6�R��U��-;DZ�b8D�`*ԫ��$�fӠ&�)w���/4D�HSO֛x�YjǮo~��;6-D�Y�� �n|���d�6U�r��!�/D��12cN(��}�`)�������)D����6F�^��d@;��P�7+D�8��ͻq��=)@ʘ39�xԨb�(D��{�݆>��
@��
6�T^�B�ɧ�xJi�'F/��M��'D��cQ��
Iw�K�l�M�R].)D�|R�b®@R�Õ'_d'��1l%D��+'FU�Gҍ������U >D�� �P�uo�#tZ`ܚ �-���p�"O��Æ%җ]�4�aAРQ�L�"Oby��DF<W$���V�- ��4��"Ov����:mwv�Y�M]�=���d"O�E�#��bL� ��ًc�x��"O0y�ŧȆ&������D�J�nUH�"O68�$A�7<U��
T��ĪI��"O���ă���a��ЩT�t`�O~qr'��,�
(k�O�jq��%O�<	�<� d 3옣>�B\��ؖ*���ȓt.m�e$I.r�z9�@�Ʒ5
�ȇ�_� |��J[�
=c/ͫFV�P�ȓ �B6"�:�,ej@�S�O�d��+�A��gY����z�%bX�<�!Wf��(�T��a�Tp9СWU�<�"*��������+nd�r��T�<�sC�6$�zQ�,E Oq���+AV�<!��8��zwIL� �f<2`��N�<ir�^*@j!Ȱ���Ncذ��
�G�<���*��P��)&Bj1�A�<	��u���s&Րvʹ񕏉c�<� L�F><��p&�:�P���l�c�<�G$޵��J�CK%Z:N�q�?T��%��k����Q�v;��`W�?D�L���Z۔������Dx��j<D��p�	�7h(L��T�lt6$��8D������cȱA��].8��`�2D��:���>j�`�k�z�Bh��4D�4�����#��M@���%m,�%1D�4c`oG�	��P	�f1[��q��a,D�$�FGשlDJ<�c�ץy��e[	(D�̒%KŦ<��T35hI�	��� P�'D����ē [�.�9F �u�֤QI'D��R�j�먬p��*�� ��&D�l[W,��t�3'��n *`�%D�Q�O�S��|����md�k4�#D�t�'
�x�%	E��	6�w%%D�T�mX�rK�Y�a��;�TĚ�-7D�RCǅnD��I��F�b�Di�D4D���g���+�$ĸ��� �
��0b1D��
7�6LHp@e�5{�b!D�0��)φc�%P�@˾�C�- D��Cرa��p�� :|�6���>�Iu��X�E�9Ź���u��̨��!D��! 'Ϩ+>X�!�PR����%L-D�t�H�5���AD���D�֬,D���S�2nޠ����Z�:�"!�(D��c���9��ذ� �4dr�!;D��A�`FgT;�N�PNb���E&D�\����6�h󨗰����,��ǟ���ɇCQ��+�L�p�R�E �/NB䉕 �Ԭ� �*S���A/��A�C��zIԭR�g�X��A�}C�IB/����<s�ir��37��B䉥5�v��b��)W���B�I�:�T)��O�b�(p�^�WS�C�	��:�Q������cw��W��C�Ɇ �*L�$艟P?P����Ƈ0YfC�I6K��bE��Q?@Y��&�&�*C�ɺea�}���J/
�X"�J!�C�	3p����O���0�QU��C�I#[�$|QE���rhtq�CQ.
(�B�	!N>8��S�>G�(�f
���B�?bK�i��F�
U*�)�t� XԊ�D1�� ��!�	�d�M�R(-F�0�!"O��k�)��F|�s�[�R��ep�"OȈ�÷2Ԍ3qƆ4�$��#"O*�3爒k��j���l��͚6"O��CdO�wb�D��E
�Wm�U��"OJ�Ƅ[�i�u�N_Uz)@"O �� ��u�d!��ȼTwz]��"OY۷�^�lˬ�� �6v��ň%"Om�0&�fOv|YM���l��"O�T��J�'Q<<{��B!	� ��"O&���	$}�X��	��i�L���"O�%z�.a�ѱǋ�,Df��e"OБ(T��*z1�8�P .�p0"O6�S#�\?�E���� �$�;"OΑ�o'#~>�3�Yy�
�"O�c�%#����C��l�θ��"OzI�L	7HBL- ㅬeBpd�Q"Or�[�F؂P�BX��5D��a"O��16l�шt�t)K�|T�D"Op�K�G@�	�̕�FjT�+Q�`�"O*�C� U49���Qt	�=P4�I�"O.!���!qIƜ��^�*׊)"O�`��d�
dũv呀j�r��"O@��$\4Zzd���^�+����"O$���l/e���GCW3^�4zq"O��"ۑK�a���B�o/>�@T"O�-����^Q�h0���wI����"OҀ�3G�>�&1��$=f��6\���	|�S�O ��p��"e��B��[ ��K
�'#�G�_�@Ȋ�G�>��(
�'o@	R�	D9f�a2����Qc�'F
�K�7~�x ���4�"��'��a���c�!2�V��!*�'](d�0��Qj�82���T����ȓb~)�g�4;�V4�v�Z�hC��	�,�!iӎ��bl��*�B䉵�f	B'@)���bۻN��B�	�"<Z�0"X;f��&D�
R,B�	1)�B�X�)��9KN�SmG<-RbB�I�)�LTzgc;=�.�KE����<B�	��h��ғY�q94jDa�<B�I�r^����0$�P�𕭁U/XC�	�S*4)"ƯC�&��Iiդ�67�C�I�Lb��+L;�"P��-�-�:C�ɳo`0J���;z�h�UH^'4+^B�	�fdT�b�j�Q��p0�%$B�	�"�T=:Ai�B��CC�G�B��-	<Ja;ec�$H���AND0�2C�I�"Fe�䅔�oY���Z�\�@�;D�,�K�4H�P��(��[0��2"8D�0:��;Z���3�J/5�H��J#D�hB5�&1��9c�*|hPQ+>D� y�AX8�4����j]*mr�j0D�ҐOj��;s�̪-����c!D�t�Я��I���5��G�tX��>D�HЦ���w�yZ#��@�f��5�1D�p��6>;�X!��E��R���<)���0>	uI� G��cs��t|~��n�<�B��:Df��&�O�/&l*��O�<��I�=O��9���kZB��P{�C��9l�$�҄f]�.���m�Q9nC䉵dZ�mR�mR�J�*��C��7M>C�	� ���X�(�N�S�g�'l�C�	�E ��'%�7.�Kb�=x�C�)� �I -�2o�DQ�5v��q�"Oh��E��jQ��KL�J����"O�sqc� 0�<�@cF);���9�"O6$�N�3[l�&�� {�5�"O6�3 �w���y�A� hq"T;�"O���#ҩYb���V+-m�L�s"O\@�4#2{�\�EL�, =~�"OH<��W�d�Z���[4G�1��"O"�3Ġ�q��X���Ok�h��"O0��!�AQI	'�%~
"�K�"O4��p(�0t~��@�^�,	�eR"Ot�;��U�q�fR>eΕ��"O���o�,l_��e^[<2Yi�"O�0˲��
 -^x3n��p:�U�"O��y��A�q�):���<@	�X�"O|R&k��2@`��L�
S�"O���jA���Ep��	��@p"O��K1
��R'���d�٦~ΖH�E"OV���@��a���*|(�"O�)��h�$M�Ҝ��	�#��T"O4��]�"�
p�0�X@u�f^�0���+i],��%�+�
��.B�� C�I�i��3��Q+Q؈:�b@#"s�B�	3X�rY�ʞ &��D��=7q�B䉵?Q�e���:��,P5�!F_�B��g\H��6�,�YA�(�&]�zB�	'.�"Y��-��Tކ�TK\2$�(C��=�V��ph��}#ry�G[=u�
C��9�ƴ����0wǤ�r�_�AyC�I/��D{�/&�P) ,�}��B��0�$+2��m_��cKڻ$�lB�ɍ\Һ
�E�'*&I�'>szC䉲.�D 㑯_�y�ToߟR*pC�Ɇa�0YK��Q�e`�yb�O�G̞���ɐ�$���*�#	�~�r��ܘm��C䉤l����AD�V�}�P!>!tRC�	<9�(h� %HH"��D�U�FC䉯$��%qܮ{Z��Pi�$�C�	�01�t�)εU �R�(W8p�PC�ɭT4���ۗl���e+T�fC�I�$�l��/_Q<X��' ��O�����I_�"��� ��mz�GC�C�!��@�׼��3��c����\�F�!�D�;3�V9�6�M4%Ĥx1�cS:�!�D�<(
�ich�|�Fz��G�}�!��Z$x6��r��<;l���ɳE{!�M�s���7�|@���!�dD��z"P*س� �8����!e��)�'f,����j�
e�fg��F�e
�'��)EI 4P�I:q���Q^č�
�'�
œ�&	�W�AQK 4i� 
�'��@�(�}���� /0c���	�'��� �".О�� I<#��aY	�'�� ȝ hY��Ĥ	L�I��'ۀ�iA�Ɨ FשތtblD��'@n����ۊ�^�����'2~A���S���2�_h���'� Ѐ�L�&H�����v��MJ
�'�:�YV���ZkY�~���'��<����+{px��-��K/�NC�X��8n7����ET���C�	�u\@�c/I6~J�X6m^�kn�B�I*lb�P�r��* �Ȑg]چB䉊l�jɉ@J��	C��Y�@�^B�)� ���:�q���m���"O|��Dg�J8P�Y!����J=*7"O����N*t2��s�Ś:B&�8C"OH��󅝭?8���N��,-�5(�"OҜx�M�;)����o��Y&8Ds�"OR�P�I�_&@C%�W&u+�"OJ}*�Ǔ�����Κ��@���"O�mk0E�~i8Z0l�t��%"O��#`j����+@�A#X�U�"O�lpR`J&����J�ͫ�"O�̓��V�~$���ʖ~�`���"O�9愇69Bl�v���"O �%eX�Z��Caؗ^L��Q�"O��E,��-wn���OK�_g���"Ol<�⌁BL2n��[�H�"OZ@���  >��3o�SW����"O��ql�$ �V�3ŲyG"O,�!���-4(j8��nG}H8I�"Od؉�%s ��KWm�C-)�"O�Xrq�w��P�hҔ��b"O`%j�쏕dY������7@�
 ѐ"O�� �B($M�Q�!9��J""O�L���'4��|�X"�T��
�y��X+)�(͒��b�J����yb���f�(�T��8i�m��I�$�y�A_* �N��p��dքMs��ސ�yRn�2.<� �%�Б\��ɊDN��y���;
���pÏ' 5�HC���y����Y%<�r�oմg��e[B˜�y���.�}`1U3gHl�P@��y"A: �ʀC<y�a����y��G�����$�91�<ң���yb�5J�x��� �5}�씻҄���y��B�$�
�����
*"�yC�`�y��1$c��ئ� �!X�+���y� �@U�i��jҌaz��9!
��yė�*S�Ʉh�e�z�2����yB@��R^����lu<�(t&L�y�ڸ.T2u����j%�=�&�C�y��,���P$�Po@�{v,��y�D%���'�^�sr$�26��%�y���_��RwL�hDh��ec��yB'�����A1h�Nm�%�Ӊ�y��ڐO�i#$��6��Uɷ�·�yr���`�gL	V��x�,�<�y�mZ�aH���sEEL�p��֌�yL�>���j��J�8)P�I���y�HM�;e�bf 8C�r�1猃	�yR��\�T53���SG$̡� �y�������a���	E2�<�셹�y�ǓDV��z�(��*���է��yB	�

���1�$�5"��hAP�T��y2�&$qX��.�P�E�4�y�#�+NzMC��է ��h2`LØ�y���(�J�2Ӌ��(Sp���y�.NF��`��͘0bRI��y"�Ԃf[�HA��4��T��씼�yr/V�j�Y��T{�Tu�R`� �y��q�2��Ŗ��h(g�I+�yR�]�J�l��M؀t��(�V��?�y2B�'6J�}�Ќo�"��5�ݯ�y��Ԟqn�J�*J�`��l���<�y2�F���Q�dۀT`���%��y��#a=bdem��D� 1�G��y
� ��yT-D1@�����\.+?HqF"O���B���G}v�AI��[/P0c"OB)p&)��0��7DL)��"O���H�h���W���[��P"�"OFC�$�*>`U*�'��p�"O��sP��(t2�Ia��^�N�(�"O�� cDGE�:�L^��8�Q��'<�I.?ڭ�`��g8X�@�'>�n��I���IG��ra)XxbJ�NH8M*C	$D�D���ٔtb�&h�.-z�%ʶ. D� ����&q8���'O�< �����1D�๷�L�K]�� C�A������1D�L�G%� +;�0)�ۜ����TH"D����!�Hb�:��Fƌ�pP�"�O��6�19G�;݌;tn��^�^��ȓUp��(�ö[\�+c��=8�
y�ȓ9.��Q��;x츒Q�_�z.�e��a���Ї@-�LD��EM	;���ȓo���(���H��Ic���5��ԆȓM��Ͱ1o
�%hz��5 ��Oza���r�RD¥d�P� 	�<����5�c�V�Tc�xؐ͌?�
��ZF$A`����i��<h�8���:�J�K5� �/�r45�f�2H��Tr�Q+vn�<M���&���~�	�ȓr� �"g�nu��@�S�4��P*��K�_�m4��nփnB�ن�+��5��
^����q����ȓ\�(��뜿5 � ��R�8�Նȓ����B U�z��F��7,hޅ��4��a�倛�h؈ؤm�i)�Ї�6/fՈ㩘4��-�t��L4��!��mk���EY�5(�AVs�-��K��Р�,���0�ZՇ��!��8����$�c��T�4=R򦉰]h�ȓr���ᆓ,Z�l	�p�˦A��,D{b�O\Ƚ�A�:�ʽ��D0{��Q"�'���:'�Ή_3(	�Q�/x�.�H�'4��oD�\�E� �k�NЩ�'�8�x�Iڔ[xx�@�/P�n;����'ӈX�% �,1H����D��Z/pQ
�'RD�yq �5"�`�ۦ��U
�+����G�86TH��&c��5���Һjs�'�a|"�l͹�#�$�TQ�kՐD�B�I�\x@�C�O^�(UjG�%	�B��K��I0�� }�����Ȃf4(C�	#P�-`@�c<�� O�)`C��472`@I,,a�pH���#��B�I:k���RÆܬ��f�=	��B�I�o��q��W�MS|��Un�7��B��3z�a��5�.���	��B��9���k4cjzZ��eĆ4+b�B䉿N� E��g�	J��b�±B`B䉌6gb�X2�%����ҳM�DB�=(����%�
�
9r��]�@�VC�&6up�[��O<�����(�@C䉭1u�`��M� g�V �`��(s�B��7=Kѩ�([�i�t�U ^�t> B�ɚ|/@�8��C�����֗i5B�I�W1h�G��o��ѪP�T�E��C����a+`�><XP�kr�$2i�C�	H����V�N'b ꖋ-�B�I+*�
�!T>�&8���G�`�PC�	
;e<0��Ǐ4�2Y;1"���C�)� ���͐3�f���(�54�lL��"O�<�E�A�r�^mHF�=2�	JW"O�i����I��H�F�Lyi>�!V"O�c�/3�H��``دj[8��w��s>�+����Y�B���ވL��� �?D���wƍ�y�.���h�}��h;�j D��AȠ3�j%�a�rH�M?D�@�cę'-��#��C=0-�f� D�4s�N�~��!a+L	��kԫ>D�"�(g<q����?l�ؔ�R�>D��2@N��M'x���C�����'?D�ؙA�/P�T��t�娇%9D�D{w(1��Q�� �l�h���2D�`���.�dE��l�=}��IW�4D���,X�V��(��Z�M*��[�a&D��
a��O�nmsS��X["�*1d6D�4�O�x���JԭNw� jv&1D�P
�	N6(�򥠤��[�N�zub3D����GȄ2a~@	��o�*u��2D�H�"c1E>~ؙ��m�u��N/D�hP	�:'�x xU�̪qF�!�/D�0A@eL"4YK#�P!� e�,D�,%��/_��`�@
,]��,D���1��jW�8I�	_7��5�%D��3D��t�DDy�,����"T����(�,6�Y��ƈv n�r"OT �W͛�LG>�3�j� �@h�"ObE�𦔥J��9p�I>x���r�	v�T� E[� z��Њ+�����)9D�\��!0جP� M*�,���5D�4e�d��Yk�ao�ei�G5D�8�񪓯ܒ���˅�(�� C�I D����ԵI�#�J �@�dI=D���a��^_�bq)�I�Db�<D�DR��)N��ȶ�0L�!�g:D�� ׫M0��;f3
�Q�I9D�\jRk�
&��\yd�,x�>��FK"D�8��!М4:�`[��:��Q��m<D�x1҅Q�HY7�L4 �~����;D���â����%P�(�n%D��*4j+g@.9{�L�	k%��u&#D��C�c�Yz�����P�~�+�!D��0gi����	BESgB��ad>D�ぐ��( ?=o*y���KWfB�I�s�8�Jfh�v\F��O�U��C�I*%- ��/'��#�.�}�C�	 ]���7��*%�]����<4�(C�I'|��U*�I��#�h�c�]8)��C�	Fs�]��P�^�"�{b��3(�C�	0�%o�}�|��� �m�F�y�"Ox���� 2�`���$?6�X8@"Ob��#��~��h��ThO*H!�"O���CJ���YX���1k���[�"OĘ�r����$�+q#�= ���"Oܸ�����T��Q#W&i/�ك"O�((�$��q�qa�?�<�"ON��L¦p��5挻���Qt"O��qg3O;�XR��H.a����`"O|���}R�rUF�%tn���R"O��u��1x��E@�:�����"O��''W6Z�z����0�2�@"O�4qVED�;0�	��'�.�8E"O����뛷xDZq�Ҥ�O�6Q�C"Oh�k�Cn1�2CH8�+"O�  dzaE*4Z�9 V�%abv���"O8p�B`V�~[��t)�7���(�"ON%���О��\����?�F�2""O"�G	�M&=�� xƜ�6"Ot]�SNL 8�tXa&�.Y1F�*`"O:�Q����B�<If�Z�/�e��"O��ȶ�I0T�)9��/E�Б�D"O�8�l�,i�U��	{�@��u"O�l�#�I�[~L)�S�Z8&<��c�"O� �B��8DQ��"c�(*5�t��"O� ٵ�V =h���'߶^!8�"O<6��lx@���m7�v���"O�����!A.�;r�8��"O2aT�^�L�r@�-
7mmJ�YR"O
�:#L(����c�>F�H��"O��7�#�j�K`i�>�*�"O�-( �G>U2�*�(�^���I%"O>H��.�7Vkp���R�r��I��"O��A�JT7��苧���R��$!�"Odr��/�Je��ݫi$J #"O�uQEb�Q���S�̻
7�mK�"Oi�s#)cS�)#��tJX�Ɂ"O�x�*��yd���v��ސ��"O������F@�)�;K��]�"O�QzR�^�@Dd r�<��y�"O2��pBYW�n��'M]#܈�u"O��8�`S-IX��d'Տ/���"O`�z/�
ӔK�
�E�H�p&"O��G�Yx6V��aAZŴ��"O��փ�2,�������X���f"O���ǥ�Nd�d�>o���c"O01J��)$���4�4D�>���"O"�;�!˥OR��E
�4Sx���"OJ-"W+�E��}��+�7`_��(F"O8�Kr�aW�!��!4yF!s"O�٠"�$���r����B
����"O���f����"d�4�伺�"OP�0f�c�2��ÁH��m�"O��4�9���� �Ã.�IY"O�(@E�Q�n{�XB�b66i�"O2̩�.[8d'�Y	�aבQ��Z1"OZt�UCОwB r��9���D"O�xkI�w��}�5h:U}�E�`"O��s#��'7m0�J��ؽAy<�"O���"��zCP`���Y��p"Oހ &�/^x�eB�*��;�"O5�$��C.T�u��)��<��"O@]��ɚ m���U!Z(v�\Q"O�1x�)�.B��%�ȪtN(�`"O��0�&�l!����G3V%"O��a�Y�\(�2�G#�R���"O�ɉ.6N�s���<I	���*O�����^5d|=�f�.J��
�'#r�z��N,D��
�2�]s
�'���2 M�D�i8p�H!*�x��	�'��0V�Z>�f�B�Z�%J|8��'{h5(��Y����v �&n˂�#�'.�Lz�-=�>i�%G(T�\�B�'5�)� P+q�#š�|�\A�'��śV-M>h�-�5^�'�-c�'zР�т�=�܄�t�� &Z1!�'�6��_�o\$+4Iï�.��'R�s$
1%إc��86H��'BJK�eؖ{qR x2M,X	���� �l[�	Ti�����cE�K��$"O\�:6�	�-�`I�� �nJ��"O:m��F�V��q�tB\ͨ"O�řa���6���b&�6 $��"O(`g�V�kbt�S�D��M��L�p"O.�J4D��@$0���w��1Z�"O��`hE4��{ �	�7��D�d"Ox���������͗�L�1z�"O��C�c��c��K�Jڹ�"O~逑��6+ܤ�c��K��8�"O���D�1k��t�U�Y����"ON<�7L��N�ِ��s=BD��"O��YV���;��u+B<��"Ol��w@M�1U�� �TR"��C"O���]�$����i͏A@��"O�1�N�  �Dxh��e@J�k�"OT�0�iF+Fiܡ���Ę(vqy "O�%��a����Eq��ڮ�u"�"Odp���$Z�1� �+ n��C�"O�-���'1����nX�]J�1C�"OL�P jK(�J���&_0`�"ORECW��0y�V��Dk -}=8�B�"O�)z�*ۋ�2P�b��o%DĐ�"OL	��·w}P!�����t"O,E`����~��4�k��\jd�y�"O
��(:R4(cs*��'�Dl��"O|Y�s,H?!� �j��u��L��"O��+N%e��������`�"OXTI4$[�%��<;qɎ�B�v=��"O���m�#=�j8a�WVN��t"O��qDZ�h�(���{Dʅ�W"O^��E�ڇ���ô�_�<¤��"O�����	6�0�#���+8$�0b"O��8uG��	V��eP�[���"On�˵$�N���"��V$!���A"ON�%�A�æ��7��q"O�D�g!K
W�d��#d֡���ȷ"O��v�����a)�>O��5"O�22�++�����C�fѪ�"O�T���:�88��Z	EɶMY�"Ov�y�A� c���A&����`h�D"O�p��N8G�A��J���jYE"O؀Xq��P1�ECWdZ�b�D"�"OX�j&�Ӹ=0rX���/3J-Y�"O@��g����t���ǰ_%�p�G"O8���� u+Z�A���v��"O�)gf.o�(jCG�M	�"O�x9�G,�0X�1o���0�"O����'��&]zܢ��/��@r%"O��a�ܳ |<4P6��=+���`�"ObHC�׌n�QC�BD�rU��e"O����-��>*p�2K����"OаR��+��|R�n��.�!""OZ��c�+S#�(�N��+�5Ȗ"O.yx�`	-H\B�C��WI�t"O�yC�V�!_Ҩ9�'�
i
@ h�"O��2f��2.���tǁ�&Q��f"O�pY�a�	j�%�sA�W;,%�"Oڸ�t�ݖ v�$8�o���B��"O�x��F�5b���J� �0D��b�"O��Iq��� p���#�I��8�)"O�	�O�c!B��ծ�f�R�u"OFŒU"�1)�,��� c���"OJ�[Dj��Yu� �EE�F�X$"O�  �#��:*��V�\5�m��"OT�@�.R��b���,fEZ؉`"O�C�Üe�椊��1n/�h)g"O�}�q�CԠ�)a��4��|""O�h����n����G��-�R�h�"O�y3�-�!:؂7K�F���j�"OF�i:).����^#b�& ��"O���v+J 
�FU���y@�
�"O��%�^��b���N\h5PA"O
e��jSi~��B'`ϐ��h�"O½��a��e�q1v��<���R"O�m�$�)}4ؤK���}���y̎y�<A��6��� �o[+�N]�aN�sX��Fy�`Y�?҄*ª��LנY�r�H��y�"�U��X1KP�m�Z�ۆ�3��s���O!�0#bg�;7��c�N� 0i���ʓN�*�bGB	R�����o-���=9
ۓ3fP@9AJ��x3� M�D����ȓH'9�eG�5���jp�@�4�ɄȓmH�ۧ����+16�~Q��tV�}�gK^�)�D�)P���M��M��*x@��2	�a1�D�L�XDz��'�(��qNs1J�BbL��;Q�ـ�'�.`��	@�
���BH�f���j�'��|��I6a(�z��ڭ;�H ���I�c��Dy���,�z.O�EK��_��H	�B;,����sӼC�	�H\Uh�b��G������*_"�b�P�'��$$�'g�����#9�"d�A�=9��q�ȓ5hFL	��p�~�r�mݹW��+���)�b��I��-�7���R
�
d&����_�'U�5��*[&ID�Ը2��(>�L}:�'�
�0fC�qߪY+��5�8k�'��I��f]4�)�Q�J9,��!��'���['��KVEa0c&,�5�
�' 0� f�+!��;Х����-D�hp��O)LW� �%OJ,<�hQBT�,��p<�k�eBB��J6MLܣVDL�<�Ѯ�q6�tEW�n�X%k�ɀ¦��=I�d����̈́�nF YDg�+_%:�ȓ����CmZ�6��s3DE''2���'�V90���'��T��C["O(ԔJ�{2�)�I[{� �낅��%�`��V)��k�!�$�|� �8g`[�Q���9�eԛ2�!�ޣ1�*�raS�Z�>��r΁(;�a{���� $]�=��m�|���j�!�$P"(A@����X O�L�#&�Pm�}���xH�$�v}�uK��q�r5�`�,D��`�f��N*�5ٲ�N�~Z|�#`�O���1���|�<ͧ�&%������[�Y�y�B���4O�����6���4�&傉X�'�@�{B+[�I� >b��� �.����MN�s�f� �u�RG>�����r}���'	�5Y{]�*��hO�S�%�0z���2V����/_) �m�I���h��$I=[~���P��"d��P�K0F'!�D��:A��se��U�D�	uA	�!�dY�P���R6h	�g�^x�g��&{k!��ߔ4�����8qHp���]!�d?�X�с�=p0F���n޹,O!��
̀�(�j��"߼B6!��S���!�"Hx� ��	F�a�	�'���0p6����S�5�iH����y2�[�k!Ҕ�A�'h��1(�ՈOt���"��%��q�c^�5��|�@nP�<a�Hݒ֬5�/��{߄����J8�x��~
� ��AE
Q�)<i�摫 dZ��"O����ꕘl�X��7�WD�>�5�	��ED��\���]j�OC9,��3@��HO��d\�x�V| �,�*GJ
�Z�ܴR!���4H�p�U:5�����̠\���>��{��ӲD���� @�=X�RXK � ��B˓��a��	�rzV�8��ͦ3�2$��l��d��\}*��v�aA��6nY㕣P9��'�ў�O���kQARM(@�IH3m¼�Z�OƒO|�=ͧJ�-0n�H/��Y�/:���ȓq�m�¢��Z� �4B�5\�, �ȓm�l�Pw+	�MRؔ;���,o�ȓ1�l<c�5�����ٯh<Ȅ�4Q�T�����@�6�p��6DY@��^&����I���P���$5otT�ȓ#�(��O��fܤ�Ȁ9Eޞ�;"�x��'����"!ЛL!��V�,��m����'b��ɵ�C@"�A����N]�'Rxt�P`d��|��h�1[r]#�'�] �CC61C
i���X��y
���~�E^���x!v�UMQ�geӌ�y��'��OD��"aK"_89�6H� in �@"OK��"w�9��`�%-Np�N���'�ў��0i��̵2���S�f2��J|��Iv̓!vA�eB�vV9b#�1OP���j�v!ai��i;��
�U�(��O����6?�U���3sVP'�D#6j�:!Jm�<��]?L��97)̡&L �i6��%*-!�IMx�DPKʕFsB�8���a{2�DX4f֒I����|�DY���ޮh��'�ў�>�
�U8K-�mi�̔ ;Tb�8bN-D��IFfE��IT�B�D�)��B�ɄAK�u�$ �0��7 ��m=NC�*M���w&،)w��;"�C�IcG��;C�Q<6�б�iDX�C�	�E:�%�C�
V�z4Q��(seZC䉃T�dbwŠL�P�����SNB�	�#R� ';k��9sd^��6��F{J?��Ot �q�]����+-D��֨>���*��Xꦩ!ғiJqO�OH�遉>��T���Y=*D4�Q�'�P蓠mG7/4L�y����u���'�HB �p�|��A	Z�N���'��ce��#i�8��a�p�왍�D%�'� q%��b�@Ap�i�
r��P��+�("�N�;5��ɋӋ,T���?�	�P_����Q�f��d���1�=�Ɠ#�@Z&�[�* Y���i_���u"O橩��Y�[��� ��$!��A�"O.9d�M;+t�X�Ši��"OP26l�H�����kнE؁k���x�O��`'	$)3�����_bl9�'����&u#������)lt ��'�&P)���g�L�p�f��feh��'O��J�
B���gDG�0aشL	p9�4ð>�%I�y�>��a�#
ֺ��Ҏ�X�'ў�'bN���R%ڷ\֘�ɢ����܅���c�9���Ҏ=�r����"�Hnm�������Z�0_�P��&�
Z"�awCG���'�ў�Od!{��Fze4�@�*�dEnU:�'��!��*�:D���z�b�`��h�'������i��1Q��s1�@L�pI lUa~S���L�tz,����#(:-{b�f����i�iDy"HԎ> <p9���=i�Y!Ӊ�3�y
� HݨWjʀ��k��6YNu��"OD�'�1�.�!�j�,�0!��"Op�&�<_rr4�3�Z�p�`�u"O���]�T�����׳BZN8��"O^Y	�*H#P%����;=f�2G���Ip�����hC���0���b�`��q�2D����ߓ[��st&
4�4�C%j-D�����
K�����N���;QM�>���_^�U�7�K7,�� bA�$����?t
10�c7U6��"��]�+����5����ۃD�HI�fAO9`΁��O9:� ���:!S3��4o�R���?_l�ؔI��[�ΰ2�"�+�H��o�xXZ��=Sƺ�q ���oZ@�ȓgB P*.��KnЭ��%`|�P��ZP�A��!�
`)UU9�x݆�nr^B���L����/Y7?}�Նȓ2G�I*�I�,�|�(�#31�ν�ȓ���b�O"xq�bG�D6e�ȓc�2��^�
���E�ԉIϘ����Lpg��� @�܁\�<���E�ZH��5f��T�_�I�@����xf\�D^���#�UsF]��e�����ύ����`���;a�!�ȓq�
�"�JȐ5m�{�Ѝ�ȓ+L��x���H��13�%մ��D��tx4
��^m�,4;5Gȕ��D�ȓx_dm	�+��?�<��Ŗ&�@!��b{f�`�b��p��V�r��h��̄���[+�ة� A?��x�ȓ�f����M8+ɤq@�ΐ��؆��V�1��,��dj� �!`B��w���#��йW�������p�4��ȓ!!b���Ԑj�8��ggX�3lҽ��a�����2�RM)��[;��%����l��+(��I��?*����NH���l �	���k6`���q��``ZDS�<�2D�?x[$��ȓe�2�0�K�+�4����Q�2`�ȓ� j�CX+*�蝐�Ê�G_�D�ȓ;x"��A�\*g~t�16�;����lfH�#a�G�Ј�J.��i�ȓz^�KC���pD�lHG�ό rx��ȓv���#�<��V'� ;����3b��D�߇Cq^9�KY���0��	"?���UL�SM�i��&S((D!�,q����HVxK\B䉦`f��ݦ| F"��U$"B�I>	*Yy%`Ϛ�(@!�קP:�C�I>BF0�rU�>AٔtK��W$&�C��A"�!���Q>#k6	[��	86��B�	�[�0��� '_2���Ʉ1|�B�I�&I��'J"ަL[��'*�pB�ɘ9���X�a@�݆���*�.�LB�	���H@%��Pb��kցV$B�lC�	������hP�\+FlB1M[�L�$C䉼#�~Pu��i�X�H'Ȃ�"C�	[�$i��E�sz1��&Z��B�	T2�[W��f�\������B��?S�l p Ag"\4����B䉄+W�5�$5&d^�X�c�91��B�	��r7��-�ĸ�Ue_�UR8B�	q��2 �ˀP̆�z�9<�FB䉏;��KeE
�B+ܽ`���-E�VB�I�a�u�D�[ juV��$1�
B�)� @��+P�@ tq��*	.�@<ZS"O\�F/��}��ى�ʑ���Ĳ�"OF���柽$�u��H<M�(��#"OzYr���!8"58 � [��w"O�;�DhZ�M� \�Di��{w"OFY�AI'VaT9��VVB�a�P"ONe��҅(I��/��C3�%�"O�iz��]��8IO)u$.H9w"OR�*�L
�u',�Z�"O���#܀F�"��U��0x��"O�dy���B^��z��DAB���"OtMk��O�s&Б�@�CY?�%B�"O���! O�P��!��*G�Gt�p�"OPat)<[�Z](�.	���""O|Y��ݓ.^0 ���<Ij6�"O@y�d
d����L�nl�� �"O	"d., ��l��C%Z��r�"O���#a4h|�����6vF��"O�HG#�\tX�4�����Hf"OU�ī�"8z��Sn+&|J���ɥO�� F�tW&g�ّ�������(C"P��y2��h��<�6��P�F�r��Ƕ�yr��m$���=E�$'N|��苇P����d@�y�I�}� ���/�E���������70#�(��"ēs����@ĳR�+�Oum�U���;5��I�ň�q�ɀ
:��]J�ϙẘ�,���O�d�axҀ�b���gk���x�AR�ۈO,�M��OO��x���C�:P@�A�+}mF���H�=2'p���|���ɔ�q�Y�g/�G�\�m�B�#w�8�	6M��K7L2�	�n�; i�v� ���N�'XtPB��'���b��3 /��r�ʕz�<�'AV����U�!,��J|RU�A���o�<qb�ꄃQB�<�*F	7椌P�*ܭKB:���lP� ��I�H(O&lPP �_����/Z��ϫ��x��  G���3�Ü�I��G?Iؤj�
O�y �E?)Nr�s��WL:0l(3"O��Yt�ڥ{�d��v$��H��Us�"O�q�D��)n��(�3��C��0�"O�9�jK�8��̪cCS�c���e"O��;FK�UƬ�2��/ �`�g"Oz��7=ߴ٩�C*rxz�"O.�y,K'O?�Ux�V-o�T���"O`l�@`�2E��R �
�R�b��gZ� R��B�S�O�baa��^�_��۶���~�Bx�'���*#"ۦ)^��sv�!v,6��O����"�0=�@��������?x�N��p�Kv���2�p a��,�=ג`	�ߢ;�$*�"O��k��%Uz��p�ϓ-�����	<t}j���0r�!����{Y���f�TW�"<9��
�Jb�~"S�ѧ<��t��%�7%�^)��[s?A�ڎ*��㞢}JUÝ%>#���J�f
\��&�{�<����ME�
�*�x�&��G��J���]��YRӓy�haEOF5<?��fZm恆�I�Q�.!�2H�5��|A�(�w��h�H���y2�	K<L��p��Y�`9eC���y"I)_����6 ��X�I�yR�"�ܡ8E�DQz�LKI�T��3,; �+@9O��!nJ I�n���M�Nu�s"O։��H�g��bL	�����I�:8�;e�P�O��%�&�F:m�H�	؏~�z��'8�)�d��$Ģu�� �p`N����kG�@cb:}�`�3�gS�25�ԿA�p]p�	(D�|Ӯ 6��q��Y�n4:Uk�!�O�P�j�Ԝe�F�sYɰ�˘tdO�c;tb�����j�A['4�L���'7tb���
�h��h�BMX\�� ,
����
�����7p�D���A#S��� �P~B�����I�[֞H��B�(H���㓤:���VS���EG�Kr@���K<vAH5%)�S�l�1L�J�<�EK'�7��:����"Hd�a{r���~|�@C�q��s!X
�ԁ����2�p �N�=�-�H|�@�484#�^��ف��͗+l$�A��[��v�=�O�ɱ3�̋ �2��g-PvH݀�,��F�PB�Ӽ��U~D���K��T� �R���Dؖ5.n�(���',�ƣU�M|�5Y���)\iD�ڎS).��ĕ�aD�l9�Aʜv/��AS���L5�f�C�zv8q�M3��QT3hW�I	j洹��q��c��S J$ji<(sU#K�rd6`8�m�<��,Տ*�ҹ��!�D� �*�	�	�R���(��l�na�)�w�	�wwl�3�d�1z�]y4��O�dC'��`KK3|O�Rw���b��G�~��=Q�(pkB �oׂw�dd�'(��2��rGƅ���MG�y���=�,@@&��$?�Y@ǟj��s��'�$X ��I'~����?���ڤo�3M̀@�@�K@���(�H�& ����%z�ْDD���')꒧�[�m���+}�Jq����<YbY�I��Q���K�$ً���{�`�!KsB�p �.|����c�9	�9�'Ŋ���G�:LOT�ˈ+�F`�f̾$�� ���� �.�Mh1�J�|	�1��	 �Ȩ�7��\� J�
|�@� "&
%E�Y#Ɇ)Nq^C�	x��8I�Ο5��ѐA	�J�	�G�J'���@�(��6 �䈐�|�� a����|�aI��K�睢gP�"�/UDQz1);D*C��-�(L�F����E���8�"	C[DrXn�!W�����|���IH�zM>1_9Q^��wgO�r�J��AAW��|�#�\S4D:�m��oA�>�%�)gް��f�
��
p�W�L"R�f�zϓ	�fl����m��,����y(̄�۲q[��?a�D�+�Dແ�I*O�*l�և�*D�4�z4���y^�B��$L�lX��	�&o�h��^�Vt�M�|�:�ƾru(��4����2�ٌ��J���� �F�,+�+ր��y2��.*� ����R�! ��U聟�r�¢JA�&5!b@]�ܹ���|RGG�<_�<j����}�d�F��xB�>A��;2 I<yX�i��h;r~��+uDL>'	���'��+�L�3��'�4�`q@}+���#P��$�Ig��1��	�W�TY�ℌ�)N��4�ճ�|-rg��dkJ�Z2o-D�P�ԄF��J�6���GdR-��o4}",�3I�ĸ�M�*N��ĈAAi�OH�`�Ȃ:8��u��*�����'����Q	�7�,
%j[rj�q�ۍ��Xc��� ha'V����Kb&��Q��,@��2Uf��*���I>꽙�)��EK��[2k���	A��K�8�P��v��-�דd���xab*7��(��F����I�7�+����D��C��i��I[�C��P�\��B���[���'�����:E�na!�c���֭s�{"��N�е2�%M�O���xk���	ّ�:�ؘ�'g~ap��#V�X�Q/�ưd�W�w���F��'w���I�Y��<�6�<(y+�'S��+͍,C�v :VIԨ. �b	�'��!�k̋,�0Ui��V�$�<E��'�.��Ë��.O^,z�������	�'�&���ĊKO`hy3Ō�'ߞ��'�N��E/ʞ+茵���og �1�' �i6�U���P
s��bn$�h�'��	��ܳ0w�]��d����S	�'��u��@�I/�e��7R�,�'�:<c��SZ�Zu��,�	��x��'��$kIwU^QAD�t���J�'�.�Z3$/��h���d(%��'�j�iڴČ��L���e��"O��h�.���K&��8x�4mq�"ON�t����N4#"��fl�R"OX���ڂ��h�&��Y���)%"O��Ң�&U�Xlѐ��)I^���"O���Ĥ� �ā��\�bM�"Oza7�޸ 4ܩY�G�H*�[&"O%�0=R��I�y�ڀ�A)I(w�!�D��LI�f�53}���V��!��K4H&�BrY"e	C*D!�R�(�LS�OȠXi�lÄ���)5 ����D1�qO?�� NDjjʰnD��E.�<��a�"O���ǃ��u�)#�	�^d"%f1O
�� 'ۃ3����E�?�^�3	�Yƨ|��C�) #�{r̊�:*�2bBئE�dD@.�|�� �V ���PE"D�`Jc<O�h�qHF>��!�C/=��6p���4$Gz��>Ar��GbL�")��iPs�/D���.N�Y��Y�����1�x�a�-;k��$�(޴���Z��~2JX�^<s�ȮXq�d�X��y�BP+Dv�s킑 ���I$ʈ��?���=Q�6012(;lOR@#�U�+���Jv�X�	��Q�v�'E�	�0�&k�XlZ�9���;�ҡOp`�r%��fC��Q� ���rf��9@M,:E�⟠�%�I�&�tYxu��6k��Y��^ �z-gMD�\�C��2U�����Q;P�"!��+@U3��2�M�F��'x��`g��=���#a��6&�~�
�'%(�9҃O�>T�9���@ȡ��'<�D�c�U�H�{�NV],(:�g��\�L��&%M��p>9�j�5W$�I�B���A`��h�(Y��<@�RC�IR/�\x)̳&�<��R#�$Y�XC��%�0M��oӾW��#���|xNB�ɩ'a�+ D�,t��ŐW�WT=B�I�S���q�bܛ42q�u�T�!��C䉬�\�%`� �8�%=^�C�I� ������
;c9)`�.)L�C�	d�*�ReY
s��<SV`�5}׶C�("�:�s6����)x4�AlގC��'3,uR�ѳP ��RWnS7:HC�	/��;���hxk�l�C�I<,�֑cWC�	w�"	�pC��+�~tq�閦
��K��N�M|!��IFʽ��I����=���ӪJ�!�$�����͇y@����hLd�!��ȭAN�`�&Z�K ���}q!��3	rb�����^8H� �Ɯ�g@!��Y�o��]�C͹x�"I��Qc[!�r��Y4��$� �A���DM!�䈪9\9j�.��B�>=��[<!��$CxWcIKnD�捃5�!�$�j�h<vP1���`�@�7!�Ⱥ6�|=J��깢U�T�-(!��ҷ�"�̞9'�Zܻ5��$,�!�d�V�(H�$Ѫ���r,J'3�!��k������o5R@k���!��/O�ܼ`'�G8� �����i!�Ʒb+�@D	��`�P��D'!�DY�1��!��I��`C��#b!�X�(!�D:f�@=扄�fX!��'T@�qC�5��(�@�!��G1hؠ��bM�pLpC(�'�!��^��H�4`E�EuP��i{�'���Yb�ɺ7��% �[9V��	�'�����$���0P*I��=��'�ޥ;����$@xP�O�'A(�DS�'
���c��D����v�ҟ;���y
�'9ޥ��n�?BsL�Qư�k7 !�
�'K��CA�޺|��Y��+���	�'��x#7Jg9(�`M��,8���	�'��}�@�+=��<���M�2��y	�'��ZQy�Zt��O�Ajp:�'v���vh��a������ �ꅑ�'C
=(�n]�.�8��5'	IL,�C�'�I{r�!.9iФ@(Cpu{�'e��Bb�	�\j�T�S��y�!��C�Ht��O�wP�jD獂�y
� �aC�­:l]@EmȬ�����"O��	���+0����6%��B���"O2���m��P�]����<~���"O��U��)h��saW�Kߺ8��"O"���C�k�fT3j�!� �a�"O�YkdT�E�d᪑iR?��Er"Oh=���6ix�Hz�(�S�����"O���B�{/:\Y�iG :�h�"O5�@(�Uo��'gLEp�;�"O���j���.��Ѐ���R"Op!jp(ʷ�����`R* p�ҵ"O�T��b���!#�-I�%� � �"O��)%E(S�В�,F�rRA�S"O�C���\���J�^'��R"OD@6)R�S�Z��s��:��(r"O��P���w��y' �6�y��"O"�����m�X=���N�	RE+"O�%8䋇7Q�^1��W�`(��"O>U&�>=&��@n]/A����"O�x���Z�3�Ґ;��i���P�"O4@ir��G;�������! "�"O�����ݪM=ι��,�
	��x��"O�	�.�~�H9�����*�H�q"OV�3�_�!���,���A��=X�!� �	���N[�ED `�'iU�h�!�&a)*	���&Ԝ��I�q,!�O�p�;�m�w��%��ӡQj!� * ���D��� ��SQ!�d�8Є�;uc@9Q�l�Cg�J*�!�$.`�e0 ǉ6�`�r��͔%J!�$�t�Ĉ'��Y�����B�W!���Y)�ؙQ�޹ZH���&۫S"!򄂆2��#��ŬlN�x�q%P�1!�$�d�i���Tg7���"	�(,!�dN�-�jȠ�e�9HQcł �$!�dϳE�
=)���i'�Y�3a�Q�!�$�[�^����( � �p�!�P1_J� �4a
4H.� Wn�t�!�|����ť��$��9�M׎"�!�I�h,|���k�?>����"�!�$..+���q�ˋ6�v��hI��!�ЧGvm�ꘈ������b�!���$�Mh�+��*�\�"���n*!�DW� iL�!����J�d�����]!��2]�8�6�Q��@h�"�!#�!���(lՐ!�j�]�C#�a�!���J���"� �B5b� Iu,!���H�V����O��<Us��Đf,!�ޝ3�^� �)�}���2�&'+!�$��6��I��K3tZ���C�h<!��)~T���GF��b�0U��*=!�J"%3�9P���B�A�!�2l!�����uLv<�����K�z4!�$FqL��J�\�Z��P"�Y��!�&jY��5/�C�͸��ٖSj!��քwj�[��7���B�X!�77Z����ڄ	��Ƭ�w\!�$D�EΌУ�G,.�|�" 2!�d74��0�׌�	A���T�V.c#!��ȩ"�\h1 �޽S�DŲB���Y.!�DN�z�b5�v,��\�0�H$EF�"��|rb'���dS�DR���,p���3U,�K�%��o��(�H�:=��05,E�
��ExB�:"ۊ�@�8s��I	Do�8R9�apA⎷~hxB�)� ��*�NS9}H�!T��(>aƅ"�����:���DXB�$/�g?���*����+Kj	۶ �Z�<Y!�Q�JM�Qh���F������$��c[X�@���@m��K#���S��S�F�����	�6��f�H�56�x��[&|`l�૚�$�����ѥ �r�9P���K�`�z��%#����^�)����c6�7�g}�#ԎXZp�@X9�
h �������� wZ�`���h��a�ˀ,� #��$䊠Z�������6E�F�D �=�M$k]�RЁ�H؞��E����2�N�gr͑���=�H��!�,D�Dxf��
}
����P�O!?�8`��i�B���P�!K0�3�F�7�(U��~�N���'U(�`#gE���[���Ysf� E�3x��a�ȉ;#��Ӆ��V"�vAh�;�zYx�B�%&t��`� �@ҝ�R�I�
F���AcC�Nqꋨ[F�G��R��-ђ��G4�4��(ޡxIV8q���/;��<A��� ���O|]�Y0>M�bʌ�m	j5bQX���De��4��9����#Z�u�d�JT���|J���  �zhGKȧE (&
�(�H� u��hJ�r�HS7|y�큒�Q�;��[Q͂2YTm�Wg]�/ ��S�L|�S�+�����<q�LهT��H�C����e�~���S�LXypp`��ɛ'K����$$7A|dç�7��I�d�KHVY�pD�v�XX��$�4`��%1�����4��7��`�)`e�� ç�(Q1K�,~Ͱi���f�j��)ܲU����'�p��/�;��2�
�B� H�O��#4��(�5 0��
��1
#�Z���O>�Q��gR��!�M9JV�+�'�x���뎹C>~�������f1�(�}���ģ	x�1-�3��O��'�9KS��%��%��hE0���I
�'�!Ñ���}�f=2�&G�dɒ�'�~i�7��"Rm�{���0 ��ě�B��p5�9х�/�p>����牲a�����;c<܍�̃�M�C�IF�`��\�B�����j3Iq�B�	�-�dk��O&`�"7`�A�rB�3&Z�ݐ��Oo`��CaA�</@B�;9�J|�6a� 

v]ۑ'E�`� B�I�0�٢7]`���V�DB��<Jr�3�F�E�Da:> �B�ɟ�:��tH��	R@A7��C�ɫ+v��P B�rٙe��>A-�C�%I�n8�`�5:�("àݥ�FC䉋^y�u���<���A��A�0C�	�7ݼE�q��HB�����E �C�	�|�Ei�j^3_�����Ϙ5{�C�~<1��&�>7����7既rC�	:*R��(�~�daڴD��rC�ɱ�RD@�+�21��q�ᐿ(r�B��L�li0�$S)`�Đ��HB�ɟ]4
�[wOP�D)ذc5M�"fB�ɣ\<2�C�'w�z�0��^��B��'O^���S�ЍZ�8��+_3��C�	1B��p�F�'	D�$�,_�h�C�Ʌ��	���rƞ|�Q�"B�P�'�p2Aos��bl�"`���'~l!��Z�]R�h	u/�e�(|��'l��ZEb�n�+�垍^V�M�'p��Cc�6Dq����K>V�:���'@�X�A�/d�������!M��AR�'���A�E�f��K#M8˦�Q�'��aȷH�/y�XK��9�pQ��'X�7��C�8��K�y����'<49�N<8Z��p*�p\R	q�'g�
C,'�N1{b�sx��8�'�*��a)��m�ᅕ�b�v�r�'wD5�ac� ~�sP��b�̀��'h�0��g�����r(�aP�У�'��\: ��;t��E����qE���'�6IU$X2n@�$W,�❚s"Ob���J���0�'͒^�,���"O�aN8�.���Lڲs�4=F"O� |��@�!MEF�W�D0!1$1�c"O���p�U�@���`�8]!.�8�"O��r�=Jin���Ga��٧"O^��iU7�����H�H��[b�1J�R�a����O��C��G?-m`�ҳ�	3���`"O��ғ��U�"Yi4l�'-��-�:O(�xe�ҔD����Ks�|E�QHU�c��{�	P��{��P�4��,1ՊӦ�z���#A�4���=\,�UC1D�$��	Y�^tN��!�(��sem5��{���"c����>	�L+"ళ�����t�2D�,	�'�+l���� �<��:#l�3r��`ޜ��IN��~���b�6�#ƤC��0���y�kH�tI�'�L�3�	�t	@��?�Ī6x]�L�@;lO���v,�hi�I�!�˱K��+T�'p� ���@�GℕoZ�q��D#hւZk��p$��C�I*S��@WNۘO˄�(gύM�㟰��)�Q�}��?8���WW2&��%�a�2n�C�02�X�8�g��z<Rlc�$F��ck� }���O�4G��'�r�����7T&�hA�P6'M��'�z*ׄ�0-�h� MU�EE��'L��b(>��{2m�cpx{��L=Q �W����p>���r\4�	"BÄ�R�-����%Z'T�|C�`ir��!j���!�;X�NC��25�P�`O�)q���dCZ�mcNC�I�2���(�"U��nM3��?	pB�&� ���l�=.xDe[ň۶B�ɰ
 ��IOy$���V j��B䉲Mp����#@8ऺ��0a[FB�m�xC�A!=R���>�.B�IO�E9��8����Q�9�&B��/I��a�Ń�� D�̠M��C�	�t[
-��N :C�
�:ޒB�I"6M�YJcBʶ��Q�0	W�{�RB�I	�JH G�^d�g�֜#�2B��0:����E-{pX�C��0��B�ɚg�Lݘм�ns��&,�x��'���KT��4x�����)�P���
�'g�4xŮѦI���s��H�f,�	�'=⁉���8Wء��%2UL�8	�'`�=1B�q���"M��5�����'h�=�$ń�|Yv �F�p���'!���6��R�"��Um�G	��'��#UE/��$��/�*5��[�'�D��f��t�*㜒+�Nt��'ư��7�Z�B��m{S(��$��݄�0� �Y�[�t�����c̻'�B��A����2�))@cI1����ȓ	o^��3@:w��	��%��i����ȓk�f}�ң��]�hpPDb�zCph��M1F���+Q�|x�cCNŉ:X&�����)7�I5g!�l��H�6�:���N(�J�!���"��g4�U��Xn�9��\ ��|��#Q�y�����ak t�aȋ;�`�
À�e��98R��@���Í	5U�C�F���b֥ATz��!I�9�@C�I;�4��ǟ�nP�ҦD;�>�'&4ب���IÏx��u��gK�;�L�U &���K�<Z ⟢}R���%�6�	Ѥ'"�DC�$EH�R2��S���Ab���	AE#�Y0�!��KƺS�,R;��IHR��ֹ�6@p (�|�F��EM�Fn�3������O,�?U�O�z�˄-J�4�3c�]���B/O���OV�k��O�hez��>$������T:Z��1��WO�	�S�j���jp�w�ŐO�TrAb `������<Yu�E	y�d9�f�A��^����`�_�TqJ�;O���寞_?�Z�"~� ��P��J2n=-��%�4P`aH�%� ��$��)��P���C�\�#CM��4+R���y"d�<1Ì����S�\�zY�Q��VKlM�jX�f�"l�K4(�a��!b�OQ?�r�B��h��,�ҥJ2w)9�����D.T��S�O\h��ȍj�py�R�IO@�K�gԒHNҪ@'*"�>��@r����6\�`��A�՗gجlR��f"�l�(�<��ij?�}�����	�hR��+2OҔRn�L	���|ylI�0|�S�V�32�x�wd�U�n4�%�� 1+OV}�I�"~��P"A#�d��HPz<�Y[�n~bK�`�����k%�O&6��+����e�&�(;O�`j����<T
 I�S.پB[���ֳn7p,K� 2�	79���ȋf[��FϘ?]��d�IĄ{�������	�?U�Oʈ�`��>�xa �P@���8[´��C`� (��Q�(��dy�X•�46! :���F���q��')�Lk"B!C:H�i,O:�}��3H���k��.��B	�caNB�I'd�����G�6D؅P!�Ȅȓ<�@ �Oܪ[-�ͫ �[�BN�ȓ3�l�2�ə��*��_0����ȓU�tJ�*�T\
Bp,d4����H������D��E�U!���'�F$���٭/�HC� H�����'d�u�5�k����b!�<F�����'��5��O�>�B����'�0A*�F���UjGNN)"H48�' ��Ct��#ng t��$_�0�'|�P�
˜�nȕ�*���'q�h����fS�q���	��P|�	�'���(��F�H����!)׳;*-b
�'?�!*V�fU��	,#��p	�'`�t�'uJ��� �|��&"OT��1.��T��DJB��#� $�C"O�5I�V�0\5(��^�b�Cb"O�Ms4τ={E�A�S'�K�V%I0"O�]���f�Z�S��T�(ڲ�P`"O�;�����X��P�O��U9"O��H��"M6����+3c,�
"O~��T�ų�xth�4gZZ��p"OjŨ�K�kKXu��U$lb��"OJ�CEֽ]n��a2�ըw�P҇"O�<B�&��$e@4�Ѕ�@"Ot(X��Ŀ:hJYJ��y��0B�"O��Y͌(Aj�Ő���5�Z���"O@��(_�m*qBv`�8\9�@"O�`:r��Ky� ���΅$'RU"OdPR�8���S4S��3�"O ���K.^BP%E����=(�"O|h�C4�.��֣�Z��pa"O��8���
g40�X6CN&�ؚa"On*F�(,6	�4'�|�`�"O��h�jP�t"zY��n�����U"O8���
�!!z�`Q��Ԉ\|L�P�"O>\����5ZOrQA�������"Oq�EZ�;N���gH�)]<h*3"O<�2��W�x-����)���0"O����䔅baD��� |N� ��"O.0���-g��H�fG�v��0�"OT�rf�J�ܵk��&���8U"O�D�ԉ[�7BP���E���"O~l�B�Q���Ux�͂)�"OT`c'+��p ���p��|����7"O��j�,�A`0E1W�O*����b"O��0@�,V����f
����S"OT���|u2qB���KWި��"O�`{oC�oV��qH�:Q�y""O� J���ŀ&#���!g�6&M^9�"O����^�,x��<�e�'"O��ذ��s/�=(�e��q��y"O��,�/8=��1B�I-9O*��5"O��b��ך ٶ��U,R[>���"O0u�J�Z��$ �� _��"O��Ab˨��=�U���<Q�"O��,/`D����A�.��"O��a����x{��.z�r���"O�y�↭6����F�1�F�s"O���S�ȫ?%���5�Q�f�(�"O�l9` �|2�H���-�����"O���Ď02��A���=�.<�'"O�P�ˢSk�E2୏�l� �"O��K�ҵcn�P�JE�$q@EX�"O�PJ��/X���K�iϗi�jMc�"O�1��K�T�P�۠iA3�|m��"O��kg�ٰ <�+uʙ���ѩ"OH��C(&T�M���I�?�^���"Oސ���
�b)��:����"O���`�P��P�a(��p��4"O���P��k�\<��F<w���g"Ox���Ӆo���@�j�����"O(d�֨�:n��I�ܽ S��q�"Oȵb���j�Rș���3`�R9b"O^5���L0$eaPȏ�Y�NA�&"OD� a�I�$ ��u�?�1��"OV9�s![m`؉�̠Zi<��"O
�G�H�wm�dW/
�uP~�3"O�l��o�d��J1耮mN��K1"O&�Jè�2h5 m �hJ�&5��@q"O��piN�,�pPA�ǀ��0��"O鰔��Qd�V燠s�UST"O@��ޠ/�6i��H18sZC�"O�A1�ă�u��L!%��Mh'"O���Jσ7M�nO� ��E��"O�kaH��)"���SQ�1P"O�$� U�e*<XP-V�;G~(��"O"y���V�d�d�b��;��L�"Of�07&�a���ln�Hs�"O�T���NF��u�*	D1&��"Ohx�t)��"f���P���`��("O"}�3	��%��\3P��H�"O�aEM�
_.zQjT�����2f"OX�ط'_��D�$B���av"ODE��K����4�#nմ��"OB���H�I�68�p,Ҩ�ȣ�"O�jU�^#r����r	�n��(�"ORX�qM�I���zTc\")�"P!�"O%YdÆ3�81��ۡf��홥"Oj요���ns�����bV��yD��<���M�$,��Y���yB	�!O�� ��BX�b�35�S��y����M����E��r���yrD^�m2f/�8�T�c��\�y2���e����*�0�l�aADѢ�yr��L��\Ќ�	��}��ϧ�yB �Rw��H��9E�*0�P���yr�ݿ ��Q�"	,F-P���D��y�;{�֡2�膿.2�oK��y��t��SFƆB�x�"*�yR�&}�`H���!/���RjD'�y�
�s@t*!�'l�`n��y�Hٗ3R��I��Г1|f��倡�y
� ���ԨA�hE�����J
2ش�"Oh�p*_<������>W��y�"OD|�wF_�+W�(��ŝ�/p�	0"O�E��m�X�t�b���+TD5+�"O� db[�}�� ĢPKp9'"Ov��&��������p���i0"O��J!@�=oy�%�2b��w��=��"O��pB]�x��3���� d��"O�ٱ� єh���vb��H��=�"O���"�	@AB��`Aɍ:xЁ�u"O����'8�����c_"�81"O�d��JS3Lp��G,�"OL���C((��}p�
D"~�@2"O�) ឰS�zub��_�I^���"O
1A��ٺY�:�hR˝;u�Qp"O^���A��Ywj�A�
�'���J�"O~��`���s`@��6�;{ʘ��3"O��G�=2�𸑯�g�2Mp�"O���"�O�T���#���"O�ě$��>Ԫ�B([�h
d�3f"ON��6ϓ�R�9�%T�^�X��B"O\[E�/*E��! �R�B����"O��˶D̶X�@��Jρ��x�#"O���J�Oi�����
hq�U`r"O�Q�iHt��pU�:ma!"O� A�$.�0y�N��.���7"OhL��I�a���1DIHX���"O�c7J���P�B���<�H 0W"O���M	m��L0En_�i�.��"Oz�b�(N����X���A"O����'Iv{d�	닺s<�"O�j��GF������wvD=#"Ob s�T�1>���I�%(m�E"O�t��!R+��z#��a�"O�%#�"Ģi��3
��J�h��p"O ;""QSv����	o�|��"O8�ڗ�K�-��|@����G��	��"Ov���F&�  �1�	G���`�"O�DQ�z��� snʈ:�:�&�R�<�S�"��)�,�v�P؇��G�<��ǅS(����i�I�*�s"LVF�<y���#�H�T�e�l5��w�<�� �zQ� K���n�P	㣔^�<A�(�7h��놐dv��k�b�<12�25��=�%��y/frf��H�<���D	�5X�CT J��w��@�<��7@�xЖ&�T����2.X{�<)�)�B!P\���-|�l���u�<Iq�0R"x���=@o�����j�<	d��K�  �M=eelEȖ��p�<�S���(.]:P���Wp�<� �ʸ0�*u���ּ��j�<)��ڮD&6X�v�J/6�8����b�<�qG>'b؉�g�N'�8��J��y⦎3,�����D�ys�usb��*�y��W"���FP�r	<5������ybC�	�����JKi�l�2�/��yraǃg�}C��\�c�dl�JO%�y" I�s�8�C�H��>�`��J��yb��:
E�U�!�G�n� cA�8�yb��!6]r�iv��<Qҳ+ع�y"��w�\m7@Y�6@�c`Q��ybLƚ#�0]�&n�8+�^�y��A&�y���7�DmUE�W4Ri��f���y
� b(����s�0�P�u�J5`�"O�U[�ϖ�T��9���2hgݱ�"O�K�(�9FD�2���d=���"O��k�BÈB%Z�k(�^"��["O�5{��K'|M��)�œ H���'f�+a�ؽV���*ʁ,<4��'b�K+�,�3+�`
�'N�e�Ȳ>��и��J��
�'�6m�!P�2y sfiҽE���	�'�ތ1���0N^���4*�	.2ui�'fP�qr����v0W��M��ؑ�'X���ǔ�0�Z�X5��0W�q��'Ȫp�&e��VtqG�[-b �'�&8i��\�Y�P���ꅴ1Ȥ��'� �1	ĵO;�(�CƊ'�����'n>��g�˵Xy"� O;u�H��'Jp������`�A� �;8�3�'�V�aďǖ@��`eLс4%�\@�'�DQ   ��(e��0+��9�"OR|P,ȟ{{��9��Ǡ���Y�"O�1Y5�\P�|;�A�g��u��"ORX�#BR�RJm3�`C��"O|I��gX#)�B,)ԮԚz,���"OP�ҥ   �����	�`$�E"O~P���$�(\
7�k�u�"O�����cx0��G�$n �}��"O�D�BW�
�0u���[�����"O���ō��i� �3�\��"O�P���!J�q���`��y�"OX��T���+�0�4()%�Lpq�"O���+=E�PIW%H�l-�DS"Od�0���V�f��IY�G+h!��"O>����� I��  �jֱrp��"O�Kj�;sO�!��o@*-���"OHA�֭ӭP�4c��!8,Z}Z�"O�;�͝0$��ع5�8&���"O�h��M7K�vQq���@��17"OL}�� �-F�+�✢?����"O��"��}�%{V��G�ΐ��"O\���.f$d(�ЏC�,Ţ� "O�}Ӈ,X�L5����Z� ��Di�"O���"�	�݋p ��2�6"O��P@�B  d����X���h!"O� ��ۉa�����Z��dyل"O����[�,�@emM�	"��"O�d��m�L��Qx��˼-���"O6	�s�єQ�b��bD�1Tw�M�"OV��b�"���9#c٥=n�Z2"OD�;#a�"lȥӒ��#*�iI�"Oh����<2�`� ���0xT��D"O0�ÇJi��=�DD۝cl��Ic"O��2g�Y?���@!>T"��"O6��d�ɵ%�J��!-���(&"O�P��K�c �� ,98�*�("O�D�`��Kz�$s��3l�hي�"O
iq�G�V$|Ļ�.�z�n���"O��	p�,fl"��V�0Yy��2"O�4[ss��Ȩ" a�x"OH ;�,=X��ـlGH�9;�"O �Rn�%kiB�C��GA�dW"ONX;�KLv���B��d;&T�B"OlDhF��(^����Q�2"Bx�"Oh�D #L�4!�e���\z��"O�����{� i�^,U`2�P�"O��Cm�>{��Sg`�3W�i��"O�5x6	��hh��Y��O���"O�K�eU�c&ظ�F�ʦI(�\�"O6��A�w~n��P暷x< �U"O� ���
ܗuAh�ѶB��z?F1A�"O�!6���r���ӧZ|�0q�u"O�� t�Ă�	'�W�>��p�"O�`�%�+7�ѩ&J��q"O���k�?'z��.��$K�"O`���46h`A���X�C�"O,��@��(����ьM� �Y�"O�%�#K�CX�	$L�9Q��챀"Ox�c��D��bPHF3B[v���"OI0���v8��ZI���9��T�<�'�_���:��  ���J
R�<с��D�q1ȏm���R�K�<IУH1,� �I����0�	P��a�<��@-[�T��1���&u)3�`�<93 ������'�V|!�g^�<i5�M %ڌA*	3��XAh�S�<�c�\�NoT��@,[#�����Z�<q���$=[�����Ћ.�l��T�<��D�Jώ� ��C���񣤚E�<!�A Z�h���ۅ_i�(!�m�\�<q4�@"KY`�`�lo� �e�M�<!�^>9�z0��<T�TRQ�<ن�ˌ6�l���ϊy���q�@J�<I�hV�*;�e�v�τS5��j�mo�<ULG#WĂ�� �x�FD��n�<IǬؼ~`J�C��K�App�@LTm�<9G��<H�bk
"ttra`���R�<I�)��=�Le��mךh}�Ț��N�<Q�HZ�6#n��e�g���F�b�<�aiH�+NpѸ��Q����᫈[�<aqo"R:����,!Z�� ��	a�<1��y��`1'O!S���k�Y�<9c���$@<$�C��!Pd!���R�<���H$�@#���_�݊��K�<�D��,ֺ���(�$�}��O�<��%șM����Kь"+ܽ�wK��<���_)kv��$'��c �����s�<2!�/qް�cvLHr)ьHu�<���VE�j�;�l�xk\���mBo�<�%�R���E��E<M�$ʕ(�R�<���׉}M�jr���x����GJQ�<9��ׄc�R�sB/�X�jd&f�<�˟�?���9�	խI��p�!Ub�<�U(�0J0�%�(T\b�DS�<���K!
{���	??u:4"�"�z�<��OW�C$�Zt;w<�=1Bn�v�<	�� ;�@�ꦆM;UQ�����Yr�<Q�A��$ٰ�9qc@��t��pAB�I�}a����.C�I�]����Yj�C��2w80h��`T�ڕ��{��p�',X$j`L�E5�@�U햗o�N �	�'�ڬ:f	L�͊�Q�Вmz�	�'�t1�RkU�d�����.;`����'�@ ��eT%g+�)*�O�"]�����'�*�j�ł�l@@���	`���
�'Ԕ��d�qb(9AD�ӒS0����'#�Bf/N+4[\@J3���ș��'�0��dДH�����	\�ܔ9��'PR����ǯh�,���������0�y�K�5��$� A��eL԰�y��%q� ��lC�g��5b�<�y" ��D&t�{ �b}�$����y�@βk�bB��DmJ!ى�y҉�3Eap��aȜ������_>�y
� �XHv+G� DJe �*N�ŋ�"O���q�=Ok�Ё��]�fc^�rS"O��9C�_������
�gVP�w"O�Ii G�Z/dl�`��39Z��"Od�0�GR%�%��?_��4�F"Op�n^"(���+AE��A��!�"O�� r���4��1���զ�+%�y��'\5c׫�'bj�p���y"�5d�ÏN�	SV�)����yr��@ @  � ������4�Ms�:(�Fs&�MG�O�=Ғ�_��E{�,@�v��Pi�"x��b1�4W� 0cG.MF(Q?9ڂ��i��_qYp(��m��'2.��,Oaɱ�7	+�̰�s�0�t"R&�$�y���kTr�;D�T�¥�'4�`ic!ӣ��0���4D�T(U �;ҪX���>Ā�#��4D��Z2��z�ԉR�o����{tL1D���℆z0i�!���*��tq�	;D�HC�H��
ѲxI�.�f�LxS>D�Dx��Q.��-[����C?D���p�W� ��'�Aey�����=D�P{2��k{>|�`Ք�X��=D�@{OG~d�d�2�� ���:D��Qd���^�@z��6X���p�-D���Gω8�Mc�T�Nj�Pd�7D��X���%3����nT�d���t�1D��x��� �}�@��O}�L�F�4D���G�k�0�hrJ��C�N�;��$D���'�\#�6Z0��'"D�|��!ˎz(F@֍A,t��k�!�y2�O�R��Vy�����M�8�y�m\���|bǂЏhRR��/��yb��	7gh���H[]��
�J2�y�`���P-�TX%㗆�y���5���R����xL�H�3�ׅ�y2+L�}��Q����j�p�������y���.&	�IX�
\h}N�R�,�yrF	�j��u`4C���y�`��䮴9B���C>!Y2C�:�y�C�]���Y�.G��98�e�0�y��8M���HWP�t}{�
��y"d\�s���2����]�� 1eA��y�Ȉ�*����P�T��e�  �y���z���HJ�y��Ņ�y��[X��O
	) y�E#�y�Ǖ� *��Ug�Y����B��y¢3����P��Q��H��y
� ��P��N�R<��P��Y�ltm�R"OB���A+=�e[G�T=n´�"O ثaJE		�L����@b��q�"O^��p�ٛ�H�[B��#k�7�$D����T$'Ѽ�p��Y7L���-D�����T&X�ҥV'/���!�*D�l ��*	�Ȅ����\F�!;tc)D���� ,P�a��� G�b��(D� �h��,��l�Vjԁ{�dg,D�\GNɗ)A��@�F�<�ҹh3�)D�TP�@��@��ŕ�b����3D�`�bLH�|&vx`�f�P�R�CE0D�HK�Ý�GĽ�1�ؚdB��AL.D�
���!a�
�k��sJ��B�ɭG�����@�+䰭��`ʄ|i(B�I	V0ب[0�[6��xr	�n��C䉓,�0"0�]H���H��	��C䉍B���ݮH�d���y��B��V�8Li�N�$_q�%B� D�J�B�	'H���#���h��1y�]\"�B�I�jp��R�����"�ڭ5g�B�	8q&;��^�������Q�$B�ɄJ
<�H��L��$3���C�I�\:��/�18�<�r�Ĳ!l C�I-?�ndx�(Q,-ltX��BB�,B��D�vp�#f�4Ԋ,p��C��KT�0�� 7ۆ�sR�-mg�C�	/Ft�Rg��4��jPf0@l�C��)_����!��|aI� �#2��B�I�)
��C���`��c�6�B�I#>|@�p��_c��#F �4\�B���JG�ӵbv���bP�z��x�
�'?Nl�G�نh� �J4�#���	�'O����8���SO G>*���'��s�h�yJ��sS�1;i�}"�'H>d��C��?�p�
�} ��'�	Sr��\�6���*e>��	�'�������Q��ʤ&��m��'`D`:a�M�Z�,CA�C P=J���'3b�KF�M8A(�Q���0I�fu��'�Ԅ
��4#�D
Ǝάl_:��'��$B���=o�T��+ aR�i�'jR�1AI�#�\���X�Y�'��uC�!�[d�-���@�V�Z���'�t80eBW<�@��S�M��M#�'�m	��?,���6C֥Bs�x��'u:4sңA�/t���M�>�j���'N�sAK+1�ix5$�(��$�
�'���i�J:*����E[���݁�'�٫#���d�@�b�4m0,��'��9���	�0���1A㕑vt`��'�ty6��]a��2gDߟj�A
�'~��*�Յ\�[���aw�!��&��Sc�8?%ܰ��m�PV���r��h��M师uʜ�X� a��st` À雼"�t*��/T&���Z�fd�#kB)}v��)�g �DZ�q��lRv r e�|���Q���ȓ�^����+1}���"cN6CwzŇ�&&@8��c�j�P��.g�I��|�<��n�Dp��T�����ȓ}�p�2�S�Y+bqP��$�ȓvj�E���_�Q���"��1�ȓ~d,	��T�12=�C���#p`���S�? ��	T�ե �vh��� P��r"O�l�t�/��Qbjٔ�(xU"O��s@.� 0�H�1�(��g��J"O��3"�7�]X6ϱB�F�3F"O@l�jY"5˲1#�Asy��"Otۡ.4T�s�J}���"O�����(���k�6��"O,P�Ձ8@_�� �\�f���D"O�m�� �&�� �3Q8#e���"ODh���&�hՁC 1����"O��J����[!V-�� \#��+B"O��k��L�M@�Y`.�&E�Pe"O���RmS��Г���,�c"O]���%|V�<��b�N�8�"O~0��/L)�t�pp�ŗu�d`�"O��S퉧{����f�^<-��+�"O0�B�J�x=���JV�B����"O���JhP����5v��1�"O� �5BF�2=��H��k���"O~Iڡ�s����-�3tߦ��"OF�;G���.�l��w�_";����"Oi�14z`f݁�DU�D���:�"OH�BG�T�/\��W�F���w"O,�CZ�j9 �8�˃�l,H�"O��@}���� ޴P�(�7"O�}���4Q�8v��o��U	C"O���&@�#]x rh@��8�H"O�1�D�m,�@1� ���]@V"Oj$PEB�1��p���<{�eS`"OP@���b��!pÈK8x��5;�'y� ��0�+�τJ.��'��t�R�ɼCb�(I���;<�v���'�t0R�)"ul�Z����4� �R�'�4��c���.�`�^9�j`�	�'��[!o������6!#�'�Z@R�M,5���beHˇT��R�'�T�0g%IE��Бt���V؎��	�'Ԋ�S�ƀ{lV�@t�G;N�*�'z�)��fڋl���@朚7	����'K�Tz��_�T�$)	�X>6�TH��'�����o�*T9�	j&����5��'q���Cͦ<+Α!}���b�'�ja�Tϗ�Y�bԆB v �qK�'�Τ pc
����R�w�b�9�'�:%�֮�Rs$(�a�qP晇�_��TK�E��|�@B�]|�$�ȓb�ЩhR! =e��b��5bC�8@��,�ЮO?2�$=�v��5(��C�;h�8�f��<I��,%)�>_�C��9Waxlz��R�HΕ�v��"O�=	v� �i�r���-��'�p��"O�1R����X�6�R(�"O U�e�0E��QJ���'���"O����嗎t��LᑊȖ7�8�)"O�]� ʛ��c�鉍tsN<�E"O��A��zO�S�ǃAX���f"O���p*�"q�j��B��6AF��"O��*�E��m���EO1*5:�!"Ot56m���Q�.  x�yt"O������ `V\[@,�"O@�����UR�hc��@jա�"O����e�0B�v����E�5���5"O�PH#-M�)�<��*���B,��"O����Ye��a�&��Lq:s"O� ���h��z� ��"��9wR�i["O��:�J¶������!t7hp��"O���	�<�v bd�Ȃk���"O^�˃��yt䈦d̓O���0�"O���Sk�0m�4�n�U�4�� "O��Yѡ޸@{.��g��1(�@a�"O
�����>W`����Y���0"O^��q��Yh�����8�ŀO�<��b�4ʰH�j�*O�����]P�<	D!J�2"��aMϤj�����`JI�<1F�ܮ�D��fQ#d�����}�<! �)QiV��dZ�`�@(��gP}�<٤�O���I���!���@0�_�<�&o˚X�b��rYC�ƨ `�<�#l��n��O5??hp�BY�<��L,gļ`��N1`��U���L�<Q�;6��<��ٸ�6��n[E�<�	F�x�z2ٛ:���`E�<!�Kұ���a��1;���ȜG�<qr��Y?�U�����i��\@�<qE���uPG�ǥ&�)��dTF�<� = o� 3#QI^J<�ȓ1�nyx��v�B��N�:^`��L����v ��g�Ή�3�F�,�%��W�P�3'g���J�D��>MjȆȓW%.[�l��`9<��u�M耆ȓn�A��aŞ�9���y#r�ȓK^�	��˶u�����JJ�ZE���ȓM˪��&��.�������lzn�ȓst�0{�	T�c��a�I!��%�ȓjm�Ĳ2`��k�x���Z�[j,8�ȓL��H�d�ߚ6������ۙL�nȇ�Iy�FK�1Szh�q%�2ڬ�ȓQ"i@�J�
�2�x��ʖJ����ȓ����s��..��2#�_�{Ld���/Y���	C�PЪ�m�"�4 ��8�\�� @�?+��d�dBG�"9H�z�;D��1��P�c��U�E=%<�1�9D�����E�+��X&��L:D�pX�n����a���9���q�*D�,��A�0����Ԯm���#)D�y���
6���H�w�`4��O%D��* �N���Ҥ-|�6��ҥ!D�h�1��?��H1��
�N�$�8u3D�T��̒NzƸQ_�$�T4W��C�I=[�x-5�։j"�=z���p"O�8R�ͼ
J��L7(��"Op�*�F	T��u��悖$:��"�"O�;�E�N4ά��/�O�F�G"O�!�#�V�&9vL����&m�hb�"O`��@&E=*Q҂c�b���Z&"O� \%�c��*"�%�a4>�@e+�"O�I���p����p�jL�g"O�0��._�;���礐�$.�y�"O��7˘J�m�D��J6��""O�L�h΁���7�7?|�"�"O�b&�wP����� 8�DY�"OV<Ɇ�\5`����P���r1"O��THݵj����Ј3�N��"O^-;�G�&�<��û&��!��"Oac�oG�J���&�
|�:�k�"O�mÁNY)Q �H�\ 3�2e�"OP%ipg
q���2$ڕW��=A"O�@A���8Ed	VC�f�}J�"O�AQp���#�СT%qH<S�"OrS�T��6����TZb	;�"O����֙_���y��1I����"O�|��5�6�h&	�,3�a)P"O�(r�@As��`��Q)�Y��"OJ��BdZ�7Z�L��o��>��0�"O�l�%�:t��9���ƀ`�f�#"O���ƣԍB�0��Եa�:��v"Ot,@w�O�L�$I	��
$�dL�@"O�zԫK�[f�����B�_�~��"O����i9L��0z&��,���Kq"OP}�+	�` ]`�O�&H�t��"O4)ɱ�֓*^�	����j+>�au"O�x�ՎTBT�s4�޺o8`q"O���Β�d�����#48"�z"OT#b]1L�^�����/d2@���"O�!�!� ���k��QRn�B�"Or�
�Nʖ>���o�&�Q�"O�%B�!S@��A��a)+�a �"O�� ��9��l���T�OR-��"O�%!�!��T�*幕���oZ��SS"O�Pᦩ�|"Hi�A�.�`D�W"O��q3�V����U���r�=�5"O��RN�m������'mEP�S�"O��`�W�S�A���R,�吳"O$���G0.�n� 1f�4v���"O�i�wE�>��b;<����V"O��;��ˊt��W�#~b�:w"O�2�(T�s�P s�E�5z:Ĺ6"O�� ®�L|�,WG��Փ�"O���G   ��     �  B  �  m*  �5  yA  	M  �X  ~d  7n  �w  ��  ͋  g�  ��  �  o�  ��  ��  b�  ��  '�  ��  ��  '�  k�  ��   �  B�  ��    �
 � � �" �* z1 (: B J OP �V oZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��	��M�#�?q������¦Fr��,/`,4��'�6m0�i>�	��p�v��.E����w��`Ǐ�����-��5$���';��đ>�R�ӂdY��N��Tf̓�?�*Oj�}�0�^.8�����֘{78�R7m̋H��$�'��'�Hnz�5�Т_v�x�ĉe�n����Bӟ��I�<A�O1�����<1.� ��Y���ؑ���<��'^��D��hO���O֡� Aհ_���xZ9��2uʑ�<Y-OX�O.aoZ�,2b�4A�DZָ�b�뜂&S^Bo S��Z �Iݟ����<�O�4c@o��d�lS�_�W�d\ ��	�6�>��P�>�'Tl������dTC���i��
����]
�,i!Z���'��9O��Ђ/�?X�ań�.�Xh�:O��m?Ϛ�3|�V�4�8B�` �j���H aDc��R�9O���Ol���2�6�Ot���J� Ҹ;��I�&˔n!Z�(�B��}�"�OX�S�g̓W�� S�
*��r]
,n(�'h�7͟Z(��D�O��D*�Sxê�q`l�8#�jyxG&�	 �H��ODm���MC0�x��d.Ёx
z�h˕��\�f!P�:�p�B)A�7�剄@��R�u��|BR�T�e�O�m��}K�/D�
jK	�*Da|�a�}V$�O�t���^�l}v�k���9|�Tu�p��O��lZN�u���pnZ�M�It�4���Wt�L](��H9XZ�K>��R�1��^�S�ߙxr�	g�V�"P`#	�0��Oe�����3g^���W�=F��peC�TRj(��ϟp�	�M��AM�dBg�t�O4����՛@2DmJ�+�
'
�:�!#�$�O��4���3�''���4=b�G	�Y�����k�iM�A�"�P#|��IO��Py��d�/Rʦ�:�A��pd	%�� N��,�ܴ9	X,���?�����	T l�
l(#�
$1n����l�62������d�O��� ��?p͚���-Z�͊'+vi[����YP*�ş�����D�i?QI>!g�S\:�\��FU�C"�L�1�?I���?����?�|J.O�5mZ�[��DC.0A�IGA��@$ND_܆�$�Oڍn�F�/��I�M�N9M�ea@AE�S�d�	O�i�Ȅ��%3��œ@X^\0�'w���B�N�2�c��H-HјV��	ܼ����D�Ol���O��$�O��D�|�D(��r#.���̕c���u�ˎT��V�G P�I�t&?5�	�Mϻt3�E�ǋ�^x���Y�1��H"�i��6-�g�)�}���'������ wP ��ֆK���ٙ'L�A��&C?�N>q+O��C���Щl�6�i �O@�̄�I1�MK�d�?����?!Sb�"7��+�蘔)�.��@?��'� ��?)���J<�s��[�x�0�ȇm��)�'6������1C�t�E?���v��ْd�E1=�����������?���?���h�����|��ֆ�+��`�'eŦ]���d��e��۟��	��Mc���4���Y�Zφ�j��� AV��g��q�d�5�4A�����?X�Iퟴ���\�P	��B>9�,�W#T�x���ȓl�)a��O����O��xcaE�7�|K�-�JiP��0&i�n�r�'""�I[�p�P�����l	�@Ґ�'%�6�Ц��I<�|b��<ک:� 1wڄEJ�>,������/{��@��'&�'A�	<��T���*7.����N�f��ݟ��	ϟ�i>��' V7���F2v���C�pc�$F�&h��
E�g2��d_���?A�]���	�0sشp��U�7$��]����Ŋ�Q����d�,��Q0��w�����>��=� 4�y��^�d��Rd�T�{�2�+`4O���ć�K���+�gT 9@C+-�t��O,�DU��)�a�3B��i��'3�Ы��wP`���ܨB�Jt�(�d���� ��|�G�)��Ax�s�l�2T�:��,�z���O:I��ӟ�����O����O�dКk7���T�`i���w�W�\��O˓)��AC"C��'��V>uQ4HC<uhe��bݪ(3 �-?Q7^�����CO>��?M+��Ohf��wb	,k�v�x�eL�b�̓0���"��*��O�.6�D"Zz2��@�},��SC�Z�P���O����O��I�<q0�iC�pbQ�x�U�e	O,-�m�5vR�'.r6�$�I'���b�P���l��=޲C �0o�� F+�ڦ��ݴC��1�(OP��ޚk����	�0{�b7�=����r��O���	hy2�'92�'���'n�U>�Q���%f�8)�N�)*f�œd�ې�?�� ӟ��I���%?�����M�;rߌ�bgd�fL��צBTD#��'u��1���tꖎ{��I�1&��F�΃q����աbgt�� j�� �'X'���'�r�'��l�!�T�4⣣K��Mˆ��O����O�$�<���i ���'���'4.��k�=+h�{���;S�D ��F}��'�"�|r�\/D�*%�qZ�
��DT"0
8��f?�4�H<��'��NײO�a��L	�V�����l�"�'���'t��S�����'�0s 6@�&�6/|Xزg	�ޟ���4hb�����?��i��O�� ]Yܙ���Y<I�2�@ڄW����O�7-�A��ÝF�@���O���խ�.T>��q�)YO��!�Z͟��'C�i>�Iȟ���ϟ8�I23�(B��8~�bM`����Q�ba�'��7m�'z�"���O���<���OD��d��YЄ�tO���D�*Bx}��'B�g2��!j�����e�Z6���n���(�1�J]���	4-[��3��u��|P�P���="���'\�0lni� Hɟ��ɟ �	���pyBKo������O,��W�#Nm�'mD	O
����O~<o�A�F��������ğL��g�&"�ht�S�ը��̚$�*>O��'�bo�<k&��`���� ��/ N9���-%�9��;>����O��d�O*���O
��,��@�R�	�p؄Z aH�#q ��	џ���&�M��C�|*��!z�֙|"A�_������^�&��1
g2@O�o/�M[�����,O �����$��ԭYA��x�v*üZi:��5E�+�?�h'�$�<����?!���?��I͸�	���J'�@����)�?����d����#v@\Ο��ßt�S�?�V��QI��H ��<@��1?�#]�<b�4cܛ64�4���ɒW�v@��	(4��Z2#@�,���V�L�M#���ch�<Y�'"�.����O��C�ǝ@r��[�l�&a�(�ON���O���O1�(�*]���U�l��Pa����v5B�B�:0��f�'��E�X⟤ۭO��oږ�B� 6+_%��U`�gE?:��ts�48ƛV��\$��柌0F��$��dfEoy�Nٜy�Y�s!�nQ��x���&�y�]�@��şp�	���ӟ�OO4T��+�&a��}�f� fy��1'`�,U86L�On���O����D�Ц�*2��(!O.g�j��$C�K\b�)۴{$���9�4���i�����d�<A6f�'BK���� �I� \�0�	�%"l����']$'���'�b�'Զ����Y�]`�T5i�~4V�@�'#B�'�rQ�|��4C����?�����)��/�4*&�I�4����H>y��Z��I�M�i�FO����F�N%�ƨ�8����8O�Q��4Aa���O˓���<�I�q9��rC�¸i��(p�@�,[��\�����ʟP�It��y�&�=Oն�1�ɓ8�,��d��`�h���O�$즥'��s����]�o8��w�J
oT�*vOf����43����{ӆ�y@4���7N�0��'T�}�c��FG�q�"�M5<�TRd�9�d�<q���?y��?����?D�Mo��(�I�t�}�Q	J���$�঱�'ŃLyr�'���^>q��H��IR��K����+"����OXn#�M[��x�O���O��a�g��1�&�[���1;SNöm�RU�<"��L����#���<YAZ�{��piEzH�!)��=�?����?	��?ͧ���ԦA�C����s��I��P��Ô|J`Ѝ��H�޴�?�J>	3Y�H�	֟���15({P���0�����:I��D� y��'�$�[�l�E�+O��I�Ԣ�%P$,��qH��+�(p�78O��$�O��d�O��d�O�?tm]�R��J-+���������ٟ(j�4ydyϧ�?���i��'����S�m܄��h��ƞ|��'���'���X�^�0�'40��b�O&[�n,Hf�&h%�Ɋ'"�-�~�|�\����������� ����?�;Q�/N��ek�����	~yreu���!p%�O����O��'+M�=�c�
��ل{�(9�'����?������|���_���A&�f�@����q\1���4���O���M��D$��S񆁠s?���b�Σy�Ib�A��D�Iԟ��I��b>��'�b6-հyT|H�4��[
�/A�>����SE�<�զ�?a�[���I"0�4��B�6$�
0۾e��t��ȟB��ny�П������?͖�� �J+��R�M�싽;vL�x17O���?A���?Q��?����	A�ߒT�$,�a���JgfW)?^h�nZ'�U�I՟��I@�՟  ����3�"Z5�|�B�(�CJ�?������|���?��&��
�(C��b�Ꭺ&��$y�b&.�d�*��z�'��'x�����I(��h��DU�|c2=0Q���T\ @�Iݟ0�	ȟt�'IN7��D�D�O��$H���0���!��<��� 
�xH�O���O��O���&^�e���[ÇQ�~$�-PĞ��鷃O;�tZ �>ͧw:�����Č�~�JDy��gyt-��?v����O �d�O ��.�'�?�'��:�t��-g�8��2�G0�?Y�i�� h��'_�dhӒ���q�:@P�a��LH��L+�~�	��`��ş�p��D�I�t����O�:�`-���N�[�h�`�ny�O�R�'���'�RJ��y�~�a�Ԧ<0�T��.l�剆�M#����?���?QI~�� @�T �Ϟ
g�"���[�5�tq�P�������%��Sޟ��	��nXP�J/BN��We�3�ZM�PJ�
��Yg��
��O�7��<1�ΕT?��q1��/|@����ׄ�?����?���?ͧ��$�֦��qLȟ �iP�5�Pё�Q�����Sҟ�P�4��'��ꓦ?1���?)DJ��h��p���2.��CG?+%�M�(O���Y�"�z�'���?�]"L(,	�ًkV�b�䍈#H�ҟ$�I���柰�IO�')ҩ�"���`�RЈ�U]X����?�����& ޜ��I��$��:F�<^ ���S�p�xb��h�I՟��I���Lny��'�����ӳp׆(�U/Y�F�(@��kʄ7n2)�	�[��'l�i>��	��\�ɰy9,}�oX<}�8�4%	U��l�	�T�'b7mP�3�N��O��d�|rs��<Y�T�g*��!�4�H�a�O~��>I��?��xʟ�(��A�0R�2�8�.[9x����"1�dP�����i>m����u��|�M�~l|�!�Y^�����U�1��'��',��Z��۴j�X��s/�7@��:p��-5*�+SHΊ�?)��_�����i}R�'��9H@Z�����A��^N�"7�'?�7��%g���?Y -C�|}T��,}r�ӱo��y�s���L�
�P�yb[�H��ȟ��	���	ȟ �O�te�V�:�^E�!��?I3I�/tӲ�"Q��<�����?T��y�%w���ibm�
0T�ك�G�R���'ޒO�I�O���ʀQM��2�>��U�)t�l5��ĕG�ϓ^�����o�OV�yL>�/O��O6E�F�Xp˶�$I�Z{�1�J�O��D�O��Ŀ<A��i. q���'��'��㳧ߙ3w�2�Z.�����ĆC}��'�b�:��σ7�hal�2tp�gx���Ox(�'D>�p�O���Ӎ9Zw2�AK~��Ʈذ,���ä,�7I���'���'�"�S����a�T rjP�E�(|c^)��OʟԪ�4Z����?��i��O��;/���ȇ�
h9P*�z\�o��l�1�M[恏����O�R��:�����E�`��[dIsQ(���UK>Q,O��Op���O��d�O",����x��X6��_� ;q(�<�g�i,�4�'8"�'��@�"b�}�Q�C.˜.!�{e�\D}��'�2�|�Ou��'���ÈؗEے��%jRj1�A���V8*��U�Of�d�-�?�;�䓶�d5a��6�W�o�t�(Ѝِh>D���O(�d�O��4��ʓO0�v&ƣ�R
A�3�B�h%HƵg)~��b��� l���
)O|�Dt�^)lڒ[B6Nq�}8�Č� ��J�m�S�I� ��}) �O$q���.�i'���ᣏ�:MP �bV�r����O`���O���O��)��?qT�7��D����ԏ՟y��e��ԟ�	2�M��*�|���<ț�|��&)8�a����%����l̢Y��O��o��Mϧ"��!M>�u��0��S�nZ����Պ�#h\Q2���O�%�J>*O�⟨��\4c,E#q �lgF�x5`>����U
r�"�'�2S>	`�EO2��惀 5b$ 5�=?1$X� ����('��'��A�"E�����6,j*�낺�dq�����4�FԂ�' �'5XL��S�D� ���c`�q:�'*�'����O��I��Mۗ�Q�;�.yU��-�*u:�n	�U ���?��i�ɧ�4�>Y��*Tf
`�z��1�
 @F� Y���y2��
��Ӻ3��ٹ���\���D��~���(�֫@v ��os�T�'���'Ub�'��'�������N�i�$�*O�b4R��Wf60������o�S�8"������Ir��Q��,�h`��@��?�����|���?1������$��\`=K�l�0C ]�"��:L0�dֳC�b�'e�'��	ٟ���r�x؁"��q0<l��� `���ԟ�����Ȕ'n�6-\��d�O����<i��[��$�U��j�5|LN�`��O����O�O^�� ��A�Pr�M�
���P����L]�.�����y�1.����O���B�#�6�J�Ĕ�LF$�p��Ob�d�O��D�O,�}���0���Td�ȡc���J�h��[ʛ$�;��Ŷi��O��X�B$�'(���yRA��$5��$�O��D�O��!H�<I�k���H$��v�� ��@��T9�^E�Ď� GD���.�$�<ͧ�?����?����?�"�Z/|�y�4E��tp��k����$Ҧ�B�@џ��I��l&?���9'�̨�*�.�\��V�I�y<T��O����O�O���O��䙐4���)E��D+�"�xd����/�O��P>���K���$�ԕ'�(���C8������4���ar�'Z"�'Br���tW���۴m�p4��`:�{ Ϛ<eVX`"GcO�~�+��ܚݴ��'���?��e8��\57�ءx��ՍR���`b�����|Rb�
�A�SK�'��{#h�f~�P���I#?ӄ�i�j��<i���?a��?���?����ٝ)���J�֣�e�r�ݎ/�"�'��#~�>d���<Y�i?�'�b�Hq�[�"��`E���`����|B�'R�'D�*�^�8�'&)|]�pΐ�J�lsԣП,D0RR��%�~ґ|[�p�I�D�I埀��Rx�<�`@A\?�9�M��t�	my"x�v�d)�On��O��''�N �Gџ@���`�� �J�`�'2�듊?q�����|��\��A��R�6�`҄T3~|P���Ñ.��L�����������'M�'c(I��)����� Oh *!z��'��'B�O$�ɗ�M�(KDȔ�ՎM�l�dY�M	�Q1܅����?AW�i�ɧ�D��>�ir��R�P�?�VTi��O:"�|�)��p�zn	Sح�'�2�І?�TD�'��̕���[`NC:O���⃋/[L�D�<q��?���?A��?q(���1��(<fb9j��]�0 U��\ަ���l���I�H'?���M�; A$5w��¯�I*�����?	K>�|
��E���ĉ�nMj`LP�U�D u��>7.�֤5�@�j�'G�'��i>��I�O��S+]�;�1p1`^4]x��	���ʟ̗'��7m
�@�\��?V��"g욐hՠ�`�+���.���?	�T��hߴ&��� ��*:���`'��(9N(8��D�W�IQ�r�*�噠j�0�%?�2r��u��'e�R\tZ 5(���)���y��'�"�'���'I�>��I�~x�qJ�#�2qoD`��&��y�I(�M�)ƈ�?I�3���4���S'�/'O�US��Ҕ��<J�5O����OpEm>K<0�'$�)JX^1��:���b�#֭?�r���	�O�D+�|�W��ǟ��Iן(���x�I	d��82�߁7n
̓W�cy"�oӞ<�G��O���O���d������ƾ �� q�'T9Mi ��'�7�JЦ�"O<�'�*�'"(8dSte�[�I��Ǩ�W,D��?�/OphؖC��~b�|�^�8!�ǘ#"G4X2�Ӫ���w�ڟ��	ş<�I���jy2�b����N�O��Fgӻ8�*�pf(?bƴ3=OB�n�D�I��I��MŲi� 6�ߕQ��!@vC�		���qƈ� u%�P�*�<1�Lp� g�?�'����wj�Hq�P�l�{DJߩZ�}�'��'���'2�'���䁤��1~F���-Nd̑p���O8�D�Oʽn������'�\7�<�$
��(�d���2���a��P�T'��mZ)�M��'(1���*O���
�jϨlY3��$j�����Y����/���~R�|�T����ܟ��Iڟ`C�$��-�� �0gÌd�����Dy��hӤ�҆C�O,�D�O�' �q���� nQrܫ���(_G�y�'o ��?	�4�ɧ���|0p���mS��ɞ�&�FQ�8u���[���p�>�Č<	gDe��\k_Ft31�
�+����O����O���i�<ђ�i��a򉞤tǾ�c�͒&���i� ��&�B�'�R6M>�����Ħ��s/=*����E�
�TARRk�2�M�W�iw���0�|"���4ڬd�'���@4Pak�.��7.������t��<����?)���?����?a(�.� �K��	�F9� b/W�����lE˦	�Q��iy��'�O�R�w��n�Rtɸ���dn�P�Q��xͦdn���M+`�x����*I��	�x�F pG�G[�)�����I��ps��O��O���?��AB<��⏬c�ԁ��_x�a���?1��?�.O��l�E0�@�':�-ϝ*(�xFEM�I^����"��'�$�>Qc�i�6�K�pФ�EF�
 I6�(�ȑ7 b.�@mh�J
8>@�\2I~��j�O���O���F׾R�9���J�a���8��O2���O��D�OҢ}λ}���+^Z�9��5,Ҙ`Jwa������4�������?���i�ɧ��w�Z���iKL��K�m��X�5�'x�6M���eܴ"f�HK>�&�U#ʈ�i&A��a��`�����4J���^�YN>�,O���Ol��OL��O���V$S�q�X�X��<� �i�l�OB���"��T� ��s����̙q^�U�#l}��'���|�O1��' �	k�Ô� ��,��`	�.bv�U�6Q�'avm5&w?9M>1+O���H�P~biK�Ŗ�!.t��PJ�O�d�O$��O�ɤ<qջi�M"%�'|�i���&C8H��)�#%����t�'�,7&�4��\�'���'Bn�$�r���<��eQ�x�X�0�|�eј딹����'r�"��0E�:
.���q$�8e�е�I	�O|���k�<��[A�찙�G�0�	!�'�6q���K�/̸:��!#0�Af��@d������-�l���rzf�r��S�<aX��C�ί82Z=�G�5?��ǘ�]w�HsG�=[��ژAN�eٱf�3}p� X�D�O��]�%�]�_����f�4�ߒUf��3c�%р ��Su�@�,��A{W�-.Ş��B
=["4h���a��B�o�57`� ��G�0͠����':��	�� ��oO�TkvcH�Cd��C�9����i���'aB�>T�����O��Ɉ*,2H)7��z�D�p��LNxc��1ӦS�	���	�ȰN�|x���HW�<VP�!���M���%5 슥W�<�'�"�|ZcDX��'����O]$	4���O^�8%��O�˓�?���?y/O��!�ǎU�u��o��r�@E8D \3���'�	�P'���I��@v��:/���F�@��5q�-�(�$�����x�IKy��4KF�S�>Q��ҵ-�W;6���A8)&6��<�����?���?���'!��W��E�&�!Т̙�@�"�O�d�O����<��Č�E�� �G-�5�P�@GDˎ|��dP���Ms�����?y�
� 5Љ{B� %�>�S �ڙC�<1�W��M���?1+O1q�]R�$�'���O �Hl�l2l�!��ͼkq�qq�&-���O��H�
�㟨��3p���%=A.L��خ}>�nZAyr��p7-�O���ON���n}Zc
�}
Q�]��V���]S�LE��4�?��y��(������:;��T/M&}ؖ}�E��//țf�\�7-�Ov���O���R}}�[��%I�u�Q�e!�?u�rH�j�M��K'��'T��������bdW
h�&�L&c�>�l���I͟��$���D�<1��~�c��y�	k�g

v�T!�0	Y���'�D�Xd�|��'�b�'��u��hԹPT4�h%d[�z?v��(l����U�a�'��I���&��؇#6��PAK9���ZPh�=Ȭ�A�yq����d�Ox�d�OʓA]����1F �
� B%
$�1�&gJ/U�	ay��'��'��'ި��F�r#�Q  �F0L�x��J�sh�' �'9"R�@�ˉ����C�!�
��'�
u|�z!���M�/OR��4�D�OP�Ē�8��0�޸s�BN��ҡH�����ꓖ?����?�-On=B"��z�S�7�����SX�س��0G��ٴ�?�I>*O��S��O��O6rl�F�'F�
�IRM�}���4�?���dó+8�@'>����?�؆p}����b2|Ollq�^CRH6��<q���?�qk	��?	H~����aπ	��!@WMD�=G��{@�����'��i0r�}���O��O���gޤ�ɱʣm-��H��E1Pp�l�Ty�͋�&Rb'�i<��iy�Ȃjԕo��$_�V3�5I�4S���2ǽi�B�'I��O�O��G�9�0�6��91/��	c���t���nZ>3v���ٟ���ߟ��S��R>Ya���N�� �#�����hۛ�M#��?y�Lبis+O�Sv��ma(�e�̆:
j0�C��H��m�<)Em�7C�Ow"�'\�-�a@��V&F���E�� 8��7��OH-��(N@�i>���ܟ��'�)���%�v�`f$єpm:-���t�<�$_�k����<ͧ�?�*O���8�d�b��=�Di��.��b�o�<���?Ɉ�'b�i��(��ˌ	`uѕ$�=D ؠ��P��d�O����OTʓh�,%B�6��Ly׏\n�}��@'PRF0PtS���	�����by��'��! �" ��s޼,�U�N�$x%eH0IN���?9�����O�s҉�|���h^L*u-�&Q6��C��bU�БB�i��O����O�rB��9��'m.��EC�A�>��B�
-X���4�?�����D��&>����?��	xqv�# N�0ia�-v��#X7�<��?I�E���?IN~���C6[��^Muf�o%�hJ��Qަe�'�B�"(sӒ��O���Oh4�A9��gB��`A�S&@':7UoZ��I�t@T��ɫ��'�(����>v��1���X�m�>4cT 
9�M!�9?����'�r�'��d�2�4�k��YP�!1�ω�e�|12G�H�DK��'k�'��X������N�2�A�����RQ4��yo��8���@���Ҍ���|����?�vLU����4��Ri��!B��Wś��'�B�'I�	3��~�'��'�*J I�pk��	)^�"��A�i�F�$N�S��5%��̟���{yJ��,����$�F]�W��%t6��O��9]��|��'��\�XX�(�	`�\�{#"��Ԁ�?~� �I<���?Q������O~��QBv�� ���I������ӡR�E�G'�ONʓ�?����?1)O
�!v��|�e�]�K�FX��+��s�9Y�fBD}r�'(�'�ɟ����9 "��ie\H��G�l����B0Z�؜��*�>i��?Q.Op��:ns��'�?�ҐM�i�D�E$1-I"fJ������O~�@6"�:I�xR�[8�NP�p������C�M����?�+O���-�D�S�� �s�	[a╕zzݰ,C�N���17�!�$�<�C%	�?�J~��O����B
I�0�ֱ0)^0��O2�DO����D�O����O��)�<�;l�
<3�ʑwRtJ��lRTIo��D���N�D�u�5�)��|G�d�A�F� �̠x�I)U�7��%\<��l�h�����S����|*��+�s"�	aa����,D)r̛&O[*{`��'��IN�4\�x����tC��8�b0k��K Q0"��ݴ�?I���?IT
n���xy��'�����eJ�h�A�5(�rU�wn�&Uۛ&�'��'׆���)�O���O�)��cת��2��N�%|q��o����	w�<r�O�˓�?�,O����� DQÊ����p{#f^�-���a�i����y2�'!2�'F��'R� x�.����>Af��A�ԅl��E���°���<������O,�$�O]i6i�)���aj����lP*6���OB���O0�D�O�ʓ^��[�:�v�b��&+k���ab
Ѻ �iU�֟��'Tr�'[�'��yb��1�Y(e�8.�����W�V��7��O�D�Ot�d�<�6�Cc������<�:�I��1X��%5����7��O���?����?IwF@�<!���~⁘����!ȒO���r�A��MC��?Q*O��2T̑D��'y2�Ov"� �aš@˪���4�v��!"�>Q���?��v����Om�IH�QjK�V�J�mǉag� S�i̦i�'j�P2�oy�(�D�OT�D� קu��P&a�ƠCf�ӚW�,y���M����?�F���<	���-�ӟbr�� HW�V�y�rE�5QX6��<J�n���p�	ԟ��S7���<ɒI��8��ńL��i����֏C�y��'l��O���?��Гr����a�Ǚ}ۨ�CFbR�9 ���'8��'��#�h�>�)OB���4pg�Np�,�����yd�2�`����<���<�O��'�r��9j>��s�]�B4֭jc�v��7��O~��D�z}�[�x��wy���5��E
1�~�����gc�K��,����T,���@�Iٟ��	|y�k�hdr���O�0Y
�I��E���F�>�.O ��<����?	��S�!�����Q���ly�H�<)��?A��?i���$˪pF�1�'F�œ6g���ة��B�6v���lZ{y��'��	��(�	��@CM{���WÁ?RӨTã��211�Q'X��M���?���?!+Oz�hrjDX���'�H}٤�C��Ai��N�^���O`��d�<a���?Q��&S�@̓��i���j��B%��t:���+x�^�r�4�?A���L�в8�O���'���ɁD�R�RuGS� ����4�~��?����?�����<�K>Q�O�	HU.ř9��G*��o)0ݴ��č�y�HqoƟ,��ٟ�������Z@B�k�v��l0&_6v�z��i���'l�@ �'��'q�X�k��)����g$)�v�j��i3����Os���D�O��d��I�OX���O��"WMV!��;���>�h$��n�˦�A����p��͟ s�������^�]�^IӐ �8-~Ъ�4T�n�����ϟ�pT�
 ��$�<1���~����ov�y��. �@i����Ms���dɢ:�?	��؟���o�D�������3�D'CzX�"�4�?���A��ky�'��֘)f}�)�5��I��iЁ~���F�����?����?!��?�,OԼ{!���֤��R���	���b��>�,O����<���?���2��"`%ܰRn�)����QX�dꄦ��<!-O4���O`��������|���ʛ�j��?
	�౱�Aئ}�'>bV�x��ٟ��I�`~��I�76�-j5�<�p�g�4��0[�4�?I���?�����W
���O�Zc���$�
�3�~uv���@���hٴ�?9)ON�D�O��d�b����Op�Ċ������.��r�pcw���dZ*�n���|�ICyBl�K�h꧂?���"r�J(�H�ʰ�
T!�iـ$	*6�	Ɵ���Ɵ(���z�@�'��֟\�cUR)�@2�NW3zARb3�i��Ʌ[�=ڴ�?)���?���[A�i�A{�A9O�$rp&\�>)(��Gu����O�0OΠ��yB�	�t���	���%���
�j�����%2��6��OR���Ob�i^}R�@S��L�1S��C��E鹄�	��M�ah�@~�W���R��vc ����#�� b#O�C�^����i���'M�ҭ�������Op�I�	�����H ��6��S�$�6��O˓w��S���'ur�'�� 0W��4H�r��7�a4jx����(\~��'���۟��'�Zc��a(�'�
N�x�k��?ɲ��ON5:O��d�OB���Ox��<��	ǐZ @dE�Z��@��Vo�iBQ���'��U�����4���6O��@�1`�j�nQb�:�
`�c��I����	���	qy��2NR����p"�Fr��)Ë&?�7M�<Q����d�O��d�O�ыR7Obi��V�F�\��B �d(\Ij7����	ԟ�������'�S�n�~2��+��m��L�1U��p�7a��9�	QyB�'��'AD�'G�s���P�'����@ ��&z[�9�@�i#r�'	��d7n�����O��IC�p�K7#�;�����F.syR��' ��'cr�������#�0�y4��+A�$Z&7��(nZFy2h67�O"���O��)f}Zw�B,�K��vü!X��Y6=S��i�4�?���S���ϓ�䓅�O��0���p`�g�N�4���۴&|��Xưi���'���O3b�� �!(T���Ͻz��}+�'��MKD�<�O>)����'ц�Eē�\}�1�f�	�Iz\x��m~����On�DM:�H��>Y���~B-_�[X6��֛7��cI8�M�J>q���?�*O��d�O����TmZ��D�D,Lh�C.:h��io�I	5xO���OH�Okl�?��e�'+�-���2��?��I�4�i�	ay��'���'���r��HZ�m�/�luva� <��Z&�����?����䓟?��=6Fd���)/1����q�*�2�䓊?����?�*O���@��|
���%(��`��5ne��L�h}b�'�|r�'��h��$� ZuX��ՍO��Z��%i�x�qY�d��ҟ4�INyr�S���t���ЁF����a�}�Bm�Wn�ߦ��	t��	�����i�$A<���2�ݷI�x4���qu�f�'"Y�������'�?)�'�d[� �	,�����Px+���f�xR�'���߮�y�|�ݟ�,K��7"P�B��M%j2��i(�8�v�0ٴXJ�П8�����ÑzdJ}���B�@����&�G,(7�F�'��%��yb�|�iV�J��pI�CR9i� �F�(8��( �.jp6�O���O��I�N�I���B�n�z$�[%"�d�XŴi.\<��'��'�Z�$E�֮5��oW:-����E�8m����	�����-��'�R�Ov�ꖤG\�  & 9eX��ӳi��'���b5�'�i�O��D�O��'&U�8Ј����G�F#"�Ǧ��	#q�:���}��'�ɧ5F�Z�J�q��/{��,٦�Ǯ��$�2+��ĩ<����?�����$� P��J�>Am:�a�50���1��j�I����Iy�	�����<ruC�%���w�99���r�v�@�'�"�'�Y�0�1�$��$��5U��"/\����C�����?�O>����?�ъٯ�?���B$9<IC�л_��Pr%�+�I�\�Iß\�'`�,sw% �i��F��P��$̠|��@�bJ�?A�doD�'�g)m�B�'N�$ْLЙ��F�e�*՚��$13���'�\��fHI��ħ�?���ö���`rDE�k�5�\0bǧE쓗?)C�ߔ�?����T?�%y����h:�>e!G��>���rA���ʟ��I�?���u�]�Bm]�MIq)G-� �4�?��Lݸ�Q��l�S�q$�M�LմN����B��M|�o������4�?���?���OӉ'��m
�j"���/�#���6Ɂij�7��������	�9�v�ݍ{�04q�f�ZP� RG�i�b�'JR'��DnO����O��;��M�fg�	�i�^]0c�ЊFJ0����ܟ�ۆa�A�T�I$*Z�v�&]��P��M���X�D�,O��O��|�iP�N�T�!�NYe-X��.q2�:q���v/�z~��'#��'��I�V���*�ڶYF*Lywd�$J��m�4+�����O>�d�O��D;�ɹ
�6dy���VT������@�D5@���S����T�	؟��I蟈` F�C��O+y�F�q)�e��}��'Wݦ��'��|"�'��E`
6�=\ Z��f
ܞ]L���&��$n����|�I�� �'����3�~��\ ؐ0r`�3N�x���9*k0u�s�i'RW�T��ܟ��I3D��Iן��I�� ��!z1�i�`N��]X��M#���?�(Od)���H��'{��OB�A�*iT���OA�a�	�%�>A��?���V����9O��ӵ9{,9߻D��}�%W�6M�<��-W����'r�'��d�>�;jP&xC�L�}�d�!�"^}��o�ğ���u���	|�Il�'G�������E�,�AR�2g��n|Az#�4�?���?���g��dyR��!I�P��$fʜрӫC�xl7m�%���9��3�SП�Bd�v����_�a��iB���MK��?��i池�_���'�r�O��	Q���
�����HA�Sp�"&�i'�'ϸ��S�T�'�2�' 
%�B��]i!�/t:H�b�
b���D��g��i�'���ڟ�'�Zc������w�H���47ڒ�!�O��h>O���?����� �e	$��+u7���iT%!� !��<��Ify�'j�	��	П�ap��-f:���ڗHrƜ���
e5��	Yy��'��'e��'϶�1�ҟ�y�wi��*�&�X���7-���E�i�r�'���|b�'���\��ݴ���3�i�P�z���&H{8��'�R�'U�Y���/0����O����	�Tt"1�Ye$��`��@��?����'��x�&�$]�d_�����Dku8L�t���Ax�F�'�r�'�"��l���'��'�����(Ⱥ��W����@
���(��Ob���OҬ
�(a1O��;�Є���LaK:tH��	�Q�6-�<ɤ�*XO�f�'���'����>��u�f̩PhÑ(p���皍m�To�̟h�I�nט�ԟ�����0�}
���� �ڜ w��>r��8AU�y�`��/�M���?I��:rR�X�'7�������@z ���
%eh|�tӢ�<Ov���<y����'�4f녺K�H�G���r�2���&u���d�O��_v.��'K�I���;��Qi��XA�ă���rc�4n����'�x�����)�O����O�Q��#Ρ?WVx*�
4r�Lh�&JEަ���a򐠚�OD��?�-OF��Ƅ	�n]�Mu>�B���5hXpek4V���oy�\�	���	ß���uy����^��d33(��Z�~p15A
>��%g�>�.O��$�<���?��"8L��[2.j���Պa_��٥�L�<�OB�8 F�
I̠��ooj	;����BlV�:��x�	�;�U���+9|(��O�-���"]͂��U���������K
K��q��n��@4��l��k7T��l0�.���H�_�(J�+ؓH��:��י��	�D��j��m)NQ�5ŔMx3M�?7|�e-׍t�<���ڃ9�<�Q����4��� � 8�4�
#"�].���SJ�X2�P"�j��1N2i@��� �PY&�E:��{�N;dM'�"��A�E��p���m�X`R�'N��q��
����W �j�r�X�.�� `ts�L�-%Z3�� �z}Y��>����n�I˱D^^�D����T	*�CC�~2��ƚE�P��Q�Ӷ.��p�t�D��m}R�'4�>��>	|k�$�J:�"�F��=��C�	�]t��Af�	�����R�r�h��$p�'�V@��`:�6�X;�*��ei�>���?I�BS�>��pQ��?����?ͻ �����H�} e��ѿ�@z��:X�F����&P�g��83� ��Aj�7HC<Ds$̀v�1��.����:���|�� �~�%fX3=�BH��Z8}�����O�	=ړR���vbZ�<��	tEW:7?���ȓ*K�Ĳ2��4Rc�NQ�;����'��#=�On�ɶ�*�zs�۬2�Q.SZ�Y!w�*Q���Iڟ ��џ�z_w���' ��b��C[�[��Q'�]"{6|�8��K%JQxe�׏݄A,��ā>p�D���C�-��
�cD� XJ�g�{��t� K�24W���{}֍Is�]6�V�8�]�=`(���'�r�	}���Y��bT?d�5�WN	'�8�ȓ�� ��=)�b��ë��h���<)4T�Ԕ'd�x�HhӮ���O�<��t_����AN��Da�`%�O��d�����O��B0�m�_�"6	BW�n�4�;��B����$T�'�lc������8Y:��1��9�E?O 0�4�'�rT��" ��oDP�`��,�k��~���	ş��?E��a�[�*I� \1�qrwJE�xR�~Ӣ,h��_6�@x�$��*%�AJQ9O��?T��Q�|�IO�4gŷJA�(қo�@�DH�V0��I��I���'P$ȖEV�D��٦� [���T>��OH�@!���",U���T[R�r��H�b�í��}s��F��/�Myt#Q A�"h{%�����ɛA�P��O��}���X��p��ؕ��]�%�O�S��d�ȓ@
T��"F�����oֺ8� 0����HO�<S��&0��� �<8�@�Ӧ��I�|��.~�yR�
����	ğl�i��C�LX�
B�K'` �]dFc`7>�\c2�	 Mk���I(����|&��1"g�=D"���Q@�.V�de�O		>I��� l��Z�[?{�X�>�O�)H�� �`��oǬ?�"�#�?�	�=�*���|��ī9�,`�Z�q&��`�`���y"���e��	@%�,�9�V�������8�t��cM�Y�JVW��\�^7Af��$�O��D�O��dB޺S���?Q�O�������=2�:i��j'	@9���O}�|��Щ:[˸�3�}Ѵ���I��m�L���X�*���qB�X����p�M	�$E�q�A�@A�p�'%��6�"ؘ���-%�����m�e���$!�O�!�X+y�6DhCJ������"OF�Z�ĵd���(ЭQ������R�*�PÓ�i���'���e^2~^����.�#0d�����'NbڑM���'<�	*O�j7M<��V|"<��'�1a��}p"j �_i�x���Y��O�A�W�Ǎ^��a����F���"u�'6x�����?���?iwkʱUD�p@�,��I["�W����Ob�"|z��T9T�q���A�p��B�n<�`�i:p���F�a����Д
�-c�'��+kP�ش�?�����[ �`�$�#D��+��F4� @�O�&ky����ONX:��O�b��g~�r!���c �j(f�������	�C��"<�*tnW��@* ���dF(��'�S��@.c������~ԉxu��b��T���ɯB!�$.l�~8C�^�b #̘6.axd?ғ��%��ףiʐy
0ş�j�YгiX2�'1bA"-x�H��'��'�w�J���âS��a#�
c�-��
U��yV�en`��%"&X��ǝ���'Tr��ϓ8?�`��(S65[������5��yr$���?�}&���1B�w�LE@v�#	�hX�0�<D��&U?,V	Ѓ�@�^�[#�4?���i>}$�T���@�r�P���o8$s��/.k0� �@����I柼���u��'�?�6��B��8D�����՜y �xk㄁TN4���'�O���r�*s�p��'.ؕ����QcL$�'�pA̡�A'QTX��hF)б�B��&?]8'��u�
��,�O�iSPOB��15��	�����'w�'B4�BO��n����l��]~���yB�p���OꄹaJFA���'��P��DO+>���I�,Ȏe<��3P�'_2��D��'��)�3�r�K��ĆMYNz��`�p� � ��m�(�	AD4N�jP��'p�7�Y�&�x��Rk%kV�� ��������wB����#$�'C����?�)O^���C�;�� ����m�|[6��O����68ƅ;l�*)��qr��+H��G{�O�7�D�#��Уu�ݵv#V(2��"0N��<�f�Ʈ}@�&�'	�]>u�1�ʟxX��=5�"caD��ȩk��ğX���w����z�S��Oڐy�%])*OpAi���[~�)3�>��ȍN���O�� R/[���eNoo�٫N� �j�ON��O��� �ӓ��1���&�h���p�c�X��ex�hK�Ď�Y�,Hu,�}����<O�1Ez"Iӧ]���Fcý+rp�w��^�66��O��D�O.�K�4�����O$���O�N�y����˹e9�L�*�2$��@����v�h��4
�uSF"�F�g�I�0 ���B���f��s-9`?�: �=D-���i9p�l�h�g�I4n'���E,��Oǘ��UhV�i���<�hV̟�>�OȜ�Ѩ�+q�bU@�d�<|��t"Olp� ��dG$�K'Cˌ�F�w���Y����~?^� �l\ �N,�f�+sH��A��Ň 8�a������ݟ�^wS�'���]�!"LQ�Cn1:��l�r.���aO�퉐��M��� Y�)��(���!�d�M�N��B���jS�,+ᡎa��y�'���-��C�Y��suB�y�o0E�����ѡ8p :V�[���'ǎc���!�O0�Ms��?--4*\[R&�:;&�)�a�A"�����,��\����|b���+{����b�ȹ6sb�HѤW��#G�Xr���"���9 l��d�"T-+�4q	h���F��<.��hi*9��@�-ڕ=u�m@�%5OF���'@�'*IC��	@�bSń*tq���'>,+тL61�kbLǰ�|��'��7�+|<�,�cݤ-�aj�"��u�1OV4�t��ʦQ�I˟h�OQTp T�'L8�S��l3�Q�w�ݪ�����'�2"�.MCb�T>�9iX���̏�2����"oF 7zrȥO8Q��)���Q(�)�N�=E����#�_#.t�'�����Θ��O�.��cZ	��Ҷ,͡q$�'�Ƶ��nI?1R�%�Q�@|��A
�
����KUA�k��X���٘/ΈtK���?�MS��?��e�q˖B��?����?��Ӽb�Y�S��[f匤y2 @Ǐ)��'>� ϓi� �ӶT�܉`�	�Tm�=��	^x������+�f���d�p��m:S �G�s��}�)�3����c=�(��/�(�  �ߥZ!�$8k��DA+ׇ)�D�ؒnY&2
���HO>qj��À;�� ƃ��a���^.Y|x��Ο|�	Ο4��q�$�'X��C�/\R@�e��!1��Ų�A�:u�x�Ɇ�)�O�&h�#!��3Sh[\:�T;7��i�<��r�ݡ�l���'�^}!��!��=bh��3� ��	1�?�2�id7��Oʓ�?ы� ,�0���QU<�a�Z��Oʣ=�O۾�P�F]�e���_�T8�����|�i،T�7��<���	�A���O��7i����0+T��͘w�R��z�D�Or@��	�O6���O���C�K�C��O���0䘘t)f88)�K~\h"s�'&9���V,sal98������'ǊPv9P�C6j�d��Q8�D�� �O���W˦Q�I.aE�l���Y�F6��En��_�<��'����SJ�����Y8?T�x��]�-�T����O$�n�:" d�Z�L�4��`A��G�j8ڴ��d'@,8n������b�D�R�[�t�k�oD
0�l3iͳZ(��'�� 9R�'�1O�3?FթZBR�g雁E�Z}�CmZg�d��2���?59�� �
�h4��:w��I3n/}�Ĺ�?a���?�����OT�qi�OV�Nt:)H���.(,�ˈy2�';�y�h��\1�^΢�E�՛�J��ቆ�HO��I<%[��ht�+�����Z�e����@���I�h�)� �՟�����8�����r5L�a��F!� ,L���k���)D�0�)�l�g�	�Y��M�톫"��5(�*yV=!N>�B̒Cv��>�O����lԍS���j_���'7�����,O<��=��F�N�uŶ�ʴ-�-aTC�W+jq�Kϲ^V�����������?I�'���c���>( J��$�[$K6dr�@�G����'��'�x�	�I��<���D�� �奇;T.�Hk�b��1��XQɓ�e~���ũ@A�3 m�/'� ���S�]���1�C�7캵SF��f��X��h��p��"u�N�HH�a�D#<a3�7� �����W�t�ʳ���z�D��Dg�O��DW릱��iy��'�����Q<�Y�'J4 @ׇ��8�)
��H�h��h+�'w��#]�,�&��_��H�y��;�,X0ņb�P�dTL}"[>�2��)�M����?)$+��.�n1���Lui��c��H��?i�P851���?i�.춵aS�i��'⢱�ק���ڤK#*Еm]J�zǓO��4B�� �P-|���O��X&
�%� \X���jʌ-'�'�Z������f)pӚ�DL�!zh�U���s$3��!>�ʓ�?����4�'+��ED�P�j�Ȳ�Yޮ��	�'Ԯ68i48�E B9���qs*�	520�o�[y"�]�{eNБ!�'ARS>!(&HF� z��� 6�
�F;�\����^㟰�	%I�)�,ؤO8����0t|૭���'I!f%�$|1���KJ���O��rRL�3B�A�2o
5v���B�(��Md��gdK6V�����<V�'����l#���'w����'>�z1�u��if�H�eت��'���'p��'&� @��ҽ�Vg=R��a�=O��FzR��%UН��&�3o�@���C�p�z6��OR���O�=��I�SJ��d�O�D�O��;|Ϟea�Z�1e�P	�� �l%�s�yrB�_�ʏ�D��<
J\R��	6&��g��.!�Zc���J�& �q��'*�Xj��ÎG�*�
�!�ͅ�:G��'��aZ�:�)�<1��7�;�)�,-@bJS��b
�'�U��.��}��Y ��2��p�O$�GzB�AZ?�*O�4ш�D6��"��Ҽ��J�ݢ9F��O����Od�$�պ����?)���̒B#(Ť%��B5)'*pC�'���<��+p�1PÌ�N
�0��R�~��A�4S�8{���g��uR/�E���b�=(�l�cڂ5ڊ,�Lɭj�,�$�O�	lџ0�'���D���|�tjW�L�n	ī'd��*�ODyХ/�z5���������6,4��^��j�l�Ky"�M�1�םퟬ�ɶ;V�2���>lg8��*T�n�����	������|�b&����z�*]^�Ԥ�4J�d����Rr �C�#*h�	��6\�����؁o�b$�F�����Q�I)	,4�P���]p�4���:O ���'���'��ҳj�Ё�A`DR�&�8��T5L��ß �?E���O�LM#s�_�G���-�xR/p������()��1�᪖�Fk�s<O,�R�Ցb�i��'��S:/W���	�@��� W8E��!_R�
T�I؟��wgިB:v=��)ML~*�@ʧ3tހ����PYb&k��(�bQ�O~����*V>�ŢA���r�"}�U��� �|LXC�$]���2g�Jl�Ĉ;H�"�'��'o�Dly�bI���Tԡ��o������O&��8B�$CG�U�}�h�j`ߦ�ax��&ғiq�Qp��Un(�%"3�F�-@�\�'V�}R,]	g�2,�WF]�/�ثMN�y�m�dL�f�� 8Ā	ǎ_�yBKBJ��%�3���[���3�C0�yb��}&��zO��|�d��R��y��Ғ^�(��"��� ����y �)>�I�5-Cy�qF�=�y2���]��uB�oW�Nf~������y�d�b��ҝK�r8��k�<�e��(A�ਇ�!� i2F^u�<IT��L��u�R'w���cǞu�<�@�N�ꕁ��H:���P�Yi�<��  B���9tA��J�~�<i��ڪg|�ӆ�����a�x�<�SA=w ���s�߁~��s k�<�udJ�Gt��1SA��P�$��r�M�<1!]�&����`J_	"`�-
��F�<iP�ӟh6��.���x���@�<�c��	��M����%0�(QI�o�F�<qKοyDUi�-آ-8�@���w�<��պA�H`�r!�a<]����r�<Y"��4V�} �L��8�*ݠF�X�<�"G 0{+�P�$%B�Z�������N�<)D=Q�\�Go�
{N  K��u�<�"�\�q$J�䔂^՜�Z�L�<Qp��=�^��d�N����W��M�<iGN�9=���(T�0L���I�<� N��E!A�6T��/Ir�y�"O�lÇ�D&�xi�Q�ǙX�T	�"O"}�����r�D$�J�'�x� 7-�j:9�'>�����O�Ϙ'*�@4�U�3<~��e�M�/L=Q��g�T��@ҊH�.�rբ�7��"��1'g$����zxs�&[ʠq.�6/m�t86�Ś#��G~R��0a�xk��Ñy����ן~ ��؆�H��L�h��
�"O�8�B瓔M�r ��cI�(1N�!1�O�m���_��E�q��Y�]G��%P%��f��ՎlI�*1�yb���"�`���G�x�<�kT��".�Hh�8`��S��u�-�媘�&�p�э���Lyp�:�㝑2 ƀ��v�azr�Ɍ� #��Q���dȥ��4���� ��u`�K1�V:�L�5}�RiKU�'�2]H&�_i"�	5n ��x���y�n��hỗ/҇`j�*Z�caɴ��?q�$�K%<؉P]�R�d�I�H�)�y2�6�� s�F�.�S2/V	2{ � í2�h2�.B e{r�b7�-vT�O�r�`�w��Lan�k����F�.�
�'�20�I[=l��hjw
��'D �X#!;��r��r/�{D��U�"�7IZ?h��b�����M�����ewV�#��0LO�UI@��?��税� hP�� � "Ϣt�փۖH�.��s�0j��!�$Z�*��l�דT����&hA��"F�ǡ|^���<aƆƣxV��i������`������عBԸ��u�Й��=JF/T)��ywA�U�<g�>�ژaӠl�H,�5xF`����+R���0��"zAo�~��O�����wFp���Ev�M����O�DY0
�'b��B�έn�`Xاj�6+�U�J�>h����� ��"Fh�D-D%/j�ϯj�px�=�qB�{D��ՂȈl��9z!kAO���*�dE4`���5���w��M�@O�k�\([R0�43Kє!�t�pǕ�eՀP��'��l��j� ^�f��42 (H�y��0:�I�x#��
䩙�ֺ�J'�����;�x4���{����Φ=�C�I��l��vy��eOB�D��S$�A?���R0 ��M�f9�#2�Z�8	����'b*����n����(�%ޜ�s���t���+9܌��AK�?���|皕h�q8���!��1;�`<���X�R4�Qc�8b���38o��*A15����'��{���3M�8��@�[nP1�%�G ��'�4�H�@b��7�F�~�Ad�Z	���D�>zm����F[���k���-D��2O���q ���:!�I�������ɩӮ���MоYW�tsm�~M
����K�(�͛u�]'qW�i�Ӭ��_S����E��9�qOz�i��E�#�:��`�X�B\J`�Ǧ��F�^;ƦӉ�p>arfԽl!��p�� w5ԈpOf�F���*��L��,2QO%�3������m�Nĳ{����ҡ 3>��2|Os`#�<�:M�FT�&o�X� ���J
�"�H�1�ax�Κ$ ŜUP�� �R��� "A�w�r���?$�h�k�m�&�$�G��� ��Q	(�6�b�D�d�P(J$�P.U����]��@�g�H�Oq:hiv�<)m�b->�뤭�= j5�1OD�'��qħ^6�xH��U\|���]Ct�E��')X����^�<���s��NE��yH�y2�D�NUPa��Ό0N�& �wJsN��P6Om�	��	;&���! `��kd:)������aF?F���®��MS6j�ߺ�O*C����Zc}ܰ��eB�w��,#t�9&p>�;�'��c ƵG
XA�AY�T�T���b���~b֕�X@�II�|��.q�|��ʒ�r�����H2uMVAS�y��h{e,��f+�(	�#� xAcЅO����!;Q�8� tY���"�  4lD\�@��x@aԍ_���'(�P�@D)I��PX��3��y��sB���R(E�D��	���'����,��:Q���v�ɐ^(ljSg��~M�9�M�/'�{"oK%,?�I��ݗQ�r��FOY<9r�U��+�@�|��9��'#`䔧��c�� DY�!�#��c���C(<�T���sR��p�aK�&��EЅ˚*2�#<QA^����-A3_"��a���0PuF�t� �ƍ�4�U���%�)��.$���t�Z,(h�-C3EQF� x�e*$ @�H��zt\ݲ��!}���}u蹸a��#���@��$��'dTX�]�h��u�*[�1F#�O���v%E�"�b�0B`��J+8���'_Bdi򘟼*Ճ��(8�Hr��W��D٘#BӋ�X���7�|���V�my@�f��/#Dq�"��-aj�ے��!F�Y�6�'���0��OqP�Z挍++TQښ�y��GeB��@V�ytt�ڷ�V�*�!��7�l=wl�j��pY�O�7Chh(5�Ǳ5O6X�Rf�Qt4�9����V��t�'m�q[�G�w�hi*�O�B$�O�u��1�C�T�U����I������P?'�h�d�'IH �ELh��E
穑���g[R�T��N柨QЭ�Ey�1�M<�=�Rd����v�ԻJv�]�6��U~"��3���DeZ	k܊�0��
��M#���=5��Z�n�eS�������G�ŚO����6�M!�zx�D��==�a|�J�e���#ŗ�
���r�.-�(R2�^�|�|��ϓ�y� U��Q 0�
�H1"����HQOT��Z�9a�4hcZl�Z��v��H��2�'�5jkJ5,Z��r��`!�Rb^8^#2��[��Г��2U(f�Er�ؘ
�n��H_:bJT��1�����c$ұ7|z��邟h�(rT��	}���X��E��M��jN�]�#���Dy2m3<�p!fiB�����õ�����tr���t��4�2�� ���}���K�i�J�&�VX�$3oo���i�&*$m���:<8���r�@��b	�shJ�G��`�SFq�O�����>H����D�z⚯o�8�����������t�.}���V�yv=�=��F�^�v<�0OlPK���7K����8�% �E3���Pk��WZҠ�%��U�'D���NS�=�^hK��x��$=6��e���;"~Ͳ��W�]˲�a'�Mv?�`��?���|�<�Q���h��)�Dٳ\ff�tn�L���'9�d�l�3}��3�vU+�K�no��	F�D�D�Z�@�dG�?$����M~���]�BVz�f< \���R��69��7�:���<��H��v�� ���Tw?�ӥ`�u@ᢕ,1[hё���M2�$3��,Od���H��ܸ'�ȅ��!z98�C�MP<�ez�)H�H�����tX��g)���?ex�w�2%!'g�X���s�P;4x�J�O�L��������T�ߩJ��&䇡Hr���у|?ϐa�E����u��Q��Z�;yx�ܪ1n׉��@��a;�ɩWF�A���|2f�|�rcY�[�t����Cj��ap��f���DǏ�x�;�N=lO�N˰gf����e
�����$솃��yJ>� 䖣B'�d�I;hۦ�)u"�Ο�'o4����(X'E�����E��R J3�	697�^h7�� �(���o��%rV��흋P�.��gU�yz�Y&oE,\޸
�ү>�V��S��y�h�5~��Qcs�>+
���j ^vXᓄ6�n�㷪�;)(F ���e�D3y�,0b�ݳcMp���#
�?����"c�<9���<��ם�SMў�9���&��01���<)��y�@�q�{�虼�?i6f3���Ӽ#BG�.qK�u�ӎ˿)��$㊜b�D��,J��hO���gZy��� c=��Ѹ� �C��,�ݖN�����'F1x��ڲ�l�O�1`��#��*H*6�n	d"V��J�cE�U2�؀У	Rh�r ؁ҧB� �b+4�D^dc��J~��}$pB��_\��0��"��$�+IB&]s�r��"�T?	��� l�UZ 9O�չ"L�IB��5l��`�H�kB�p�  DzhQ��f�"r�O�-�ED��Q;�b\�r�8�(Ѓ��e��?Y��jL�28�*ԋ�B����s& hT���e� Dvr<�5��	=o��T�I���yc��!Q��Z�`P<�B�)E�?8��(���e�"=��8�Ȅ�W�.?��nѰU{�M�UDޝ~�̍pbϓ�2�'����ۦ�9�iʂ!+����$'h��kנ�*c*��#)�	�j�*��+��1jMp��Y�6ZA궦#?A�i\�DT0ūҀ���4F�k~�V�qODUrA�âF����0N�4�z���V�!r��Q#*���iX����ja�G�4��c�8{���?˟����C[}�< qd�R�#O&�p��|b�B�c�&�r�+����Dӣ�2��'�Ƥ�!
D��Fx��֗/x��� e\
��'��>�I�՘Ł��E� d� ۥb���xT�I<Z\u
D���qO�Ӑq�2qϻ���$+w쉷M
�F�h�����O���{��}��6b>(4��E�YfH�ӌ��y�1OH�ׄ��9�a!�R��t8����\oA,}��jӕ2�^(��΅�Q��y�bõrS^)��ƕ�u���,G� ��EpjU�gLؽ#/�$U�rU��O$'!V�{�b��IP���?���`	�x�D�$,h4Li'Kݡ^<��螧T�I��FӴ62����$ˍEQ �p��F�7��t�al�+���Z�DWAj��>�Ą���&�u�'bJĊG�N9-�\����0xj�#�T�8���&�U)/�.��=�O��� P?��YK���-6�䋃M��O�^�"a���d���`w�L�xXy���Rf���O��PS�k�*\_Ȳ� G#(����/�I-c�����u8f���M�+�rc�<�E��l@&�pB���q�z4 b`ΓQ��l�<ӣW#`����9#P�;��F�`��(��Oߒĭ�9���+R�n�
�A�"*z�,K 薼S~�xR#��>dV�Y�GQ�}��(���0d(���5����/�)�'(rpd 'jV*�=i��Ζ&�:e�㉊��e��zۚ��	�O�8�(�Ν���Y/;�ڙ;qI^����e�̉]����{*�j�1s�b�����]4��p�@��F�\pȷ�!}�=x���gQ#�޹E��F6�l�ÅD�*=�މB��zi1OވF��:��aa��V�t��w�ĜN� J3,C�Pɦ��	F�y���� ��tC�$�'���A(��dJ"ɔx,�h��bX��E([
R*���gy&�B.��z�Z���(U�"��ys��'��` o:_�1�I�)���GS2Bx��a���1S�@�Ƃ��4$!����y2AK�v�V�9$��+E]X3W i�铗�' F�{���+�X1S
6�y�ρ�`IV�+C�����97)�UV�$e��6��H�'g��]*i$,�ƅ��1*�kW:g�d�DàjT�A���F:v�qRGF�?-�&��'j�$�3u"���tt "��|$���#����%EW'��	'�?� ���J��� 䲀O�H]�͸v!�p*QOp$L��Mʬ+��I��A��� O�T�S+r2"���	G,	���sF�ޝ!���I�=pŐ� X'$�S�?Kd�)žith�R7�+!q�9Qt�8)F}"G�5CN�/�3E��郗j���Ϙ'αؑJC�;J�1U�ì' ưX�O�Aa$�Ƨ�@�c5��;3BI�=Y���]qΡC��l]&%�,�v���Z���@��mBH"qF}R��yg%�B$���kX�6���&)	ֲ�"4AC;��c�l�T���!��-�'D�$�-{b���dS��|�y����#>�aG�Au�m�j#�S�u�������Ov�p ��ϔ�'��H"��(+�f����|�uH�~]�"R��<���<���5>�"d{��3}��I�<>c��c��)YH�k#ɉ\��ϡvn�{����	Ь����-��鉠!�4��g�L��IS��<)��
r����b�#۬e*B"�b�������Ğ�,��٢�	�4{��CvW!�D<M����p �+x��T��F!�$I8|ڄ�[=&�|`:�%R9K=!�d^�%M@lkW�A&L�y@1CL�E�!�č�3�֕�K[�0�+�G� %%!�H�F-hD���y�8bU�B5);!�dI/lX��X��ıyjt xI �!�D͊њ�ҧ%�sc���! �!��
 �Iz�MN����i���MY!�0sY �ф� �z�@�b�ƞd7!��d��X�(�!U%���R�Bg�!���0����� �.\""�ԁr��C䉠>���3%�W�F���e�?VFC��(_ƹҧ���v�t�#Q�˧��B�ɯH�zY�'�ץFVJ�b֝��B�I2jݦ5!pJ	%&I�H��һ��B�@�NVR�@ L0㣞$��=��'u��M�;P�'fG;�H�'r�k���|�1	�Z�2�yr����$y4L��afe���>�y�ϚWS��7#& �:��1�yo�$:�R|�Z-!� ����yN?i�<��(\�D�nH�f(X�y�'�2��i{`"�9�� �T��yB�͜e�,Y#Ç�$�pq�b��yb(�Q4�Ԉ^��Xly1���y2)�(K�fG���D��s-�y��
�]y\e��!��h��T=�y�`�*j7����l�j��e��y ���Ȩ����^�dA���y���0P4uC#�� VIЃ�D5�yB^�N�F���@�p���iC��y�$��O�L��E�Μc�y�s	�yүD�dļ!�dj��X���S��L�y��=�����|��$�B 	��y�dN/f摸e��:{�q�򭑭�y2DT�,�R蛺)'��� L��y��YR�*�H�"�v8���4�yr��	�F���K�o� Us�̖�y���U�h��O��|�\��R@���y��	�&v����\�r4����Z=�y2I��o(杀��"m�ƙH�چ�y��
�`��q��bܘQ8��	�y�Q��1"O��H�%�����y2(L�X|��JBC9N�����mė�yR"���V���_[��$̎�ybO�eޔ�5j�&(sR���S��y2�Y�R��:BM� �d�Kt���yba�V� �"p�ˬGҰ�j��J��y"�M2B� ��@��iA�H����/�y��Ɉ0����3���54`Q��P#�y�%*��t��Y$��)��͈�y
� D���B�Kz����p�T;r"O�Z&�0-���P鞗o�,��"O }���}��� ��Q����W"O�\�q��(D�����w��E"Oʠ�䯗�� �#7!DV���"O�Y�s�W�Nfh�����>*&"O%����q{��S���$D8h�6"O�ա�����e ʕ8#B`R�"O`���#2)�}k�,v��cA"O$q��*li2�K'lh�\����y�n�2f����%@m�9@�П�y"��d�����$�pTcB ���y�@V�.$xh�Y�s�J����yRH�;��e0!�;3�}C����y�J�'
	Н�!G�@r���D��y��o�ڳ��"1��1��(���y��=qL�c0�_%�>��@$��yr�Ɣ�^�hdȜ#����e�&�y"�/+X,io�p�t��H@��yҫF�9�q�Ҿ~u���	�!�yR�H�g$�C��R�w���dg��y#�?�|L�V���&!9
����yR��	i�tS���6zB���Ǖ��yB` /ZS��)%�ě1�1���4�y��9KIҥ�'��<$5ڽ�����y�� �Ʊ���Ѿs��bDE��yBe֯*0�%Y��\(�u!���y	�*[�֡�D��#N6��9b� �~b�)ڧtZ�`�E�"�Iҵ)��~�P��=9������A�NDf��3M�3�+!%����R�t�8}i���|.=��Ɩ-!�d��� ӃǍSQZ��A�@8!�QPd��P`��S�PKR#n!�D�;B,�LǪG� ���U�!��=��Ȁ�[(������q�!��-�ASbə4������;�!�D�~����u)(�ڤ��a��!�DR�d�̌ "��x��#�b��!��.�N�RH�R�����L��!�$v�i��MH�;�@ȑ�O�	m�!��3d
.��߽|��H�CC�B�!�D�8a����׬�Ш:em�,F�!�D�C#���e ˶c�p 6�[�Z�!�$+f�����3|�G�8
��*�S�OZ|�1��t>��n�D#Fy�
�'�m�T�9S�<��敕D��̳
�'�N h����{-2E���8*c
�'*�`cM��G�zd�G��2&��S
�'݀�c��)D	�	@�2ŀ���$+�r��(�x�9��E�(,(AQ""O:I�3��0�F\��₈{��F"O�˰���c�4��p�v�
 "O�����L|
��1�8X�P�"O�����2A����M;���Ж�M����ú>]�0�U'@�lN���$D���'GR�݂���R�t����'�d3�Sܧl���M�P�,�bΕ�|�XL�ȓah8{�H
k���S"L�����ȓt����p�ƥ��I�D솴e����<�* {�팈��x1�@������X��0iT+�R�:Ԯ�0( .q��	�I֨#<I���]��I6�űM��В5��_�<)�bص#@x�HS/YIx���	UyB<w���Ӟ|��)�Xo|�9�BR5F��Icҩ.I�!�� �� S�[%:͊�2�iĢ1�
�zF�d�z���C�G� Q�N�����D��UG�+D��)�(��ؽ��Y�mz� G�.D�P87��&��M��-�0m�k"c.D��HU�N+b�D�	�Ɨi ढ1m0D�,A�с;~�j6�%4w��f*OZ�i��R鄘sc�0/���t"O�)z���Q#�t�&��&�q��"OTLɆ'7B`~	砗(WiAu"O�yI炙ȩ5b�w$iAG"O��x�h��C�K��A�$*�"OR�R���-&��ka!�!�R���"O�m;j_9�܄����-?�<ĒB"O��g�$
�f���F�-x� ���"OV�c�jD�y���s"����@&"O�DC�l^�/R,!�%"۱8��Qr�"OL���~�T�aR��1,�����'#!��%J�ҹ)U,Y &�hi��	�!��	�AT��l�3	�n����v�!�D��0H(�S�G?,��ۑ��Nz!�77h��ǬR�N�~:�B(�!���$&��+��yY�a�Y�s!��^%X� ��S5x�`p����V!��*A�R���Rp$�x�C8)F!���1#
���`y���(��ךW�dB�I/Q�~���fՈ�¸ʶK�(�NB��0w��$ N��h���ϐ|����hO�>)0Sd_8e>2a
ɺw��Xe@.�O����5�M;y?��h�A�7m��ȓ=��9�?|�2���ȓ|�p)R�f�(\����M���JX�hC:�����ǁQe���x���hp�����k�M�1��Ia̓=9P@��6|�t`ۡL�)z܆�V3R�fж�*@���ӄ	�����ܛ�S�a� �z�J�Mn̔�ȓgV��	�-!��vAۊ���Ol�=�������`�B�5(v#�]�<Y&P�v���	aę=1�Vū��]�<�%$ɫ�də�K���rY{#���<�*���L]�u�ڿTtNȋuIU@�'��?��yz}3G��OފU[�>D��"SD�h'~e)�.^*4�hU��C���F{���_=s��QCu�U:"8��S�[�lN!�$���֐p
H�k��xc�Ӑ$!�$N��=
��@$p1ˤ��z��	h��H����-
��y��n7�!�v"O��rPi�xr,I�l( $�"O�X#2��<����	.0�#"OHM�fՠD� +�B �=�L��"O�6�N�&��;��Y>Ӑ�"O܅i %	{~�C5l�JWPC"OPʗ/Ɯ3'*����M�sT�Љ�"On!c�`��pHx����ZS(�b`"O�#%���d/��m4LJ�H!�"O�MҡI^?���0F���N8�&"O��{4C�h�8��=��"O@,��-��N-�DIH�X���S�"O��b �Ԋ  �T�a�ƹb���N�<I��_,��x���R24���b��K�<1�}hB�#���9/R�Җ�_P�<@��>���@��;I����kQ�<����#�����X�3� �O�<��ʛ�Z�����Ψ��Pw�d�<� m��j�:a>&	ۓ�c!ƍ�"Odth�/3�P��A+܁3
�ػS"O�̒2̅�Jr�Ջ�»2�B��"O&H�A�9%�B��
	w -��"O�HFȏ	 ��8&�Z��A`�	F���i��1� DҲ�!�����	 ]�!�dǋn�Ҁc���8A�~b4a��"O`���+@6�u�cD�ߒ�K��y����^��S@E(!*���'���yb�]�"�d�'+��r�y�Wo��yb�GP��DcQ�4���b�-�y��\e�ᙦ'ŗ~=0�I"���y�΂�z[��Ҁ�$qU �k!E���yB���.�Y��탻j�:]Y���y2č ����rW	�<�A���y�F�\��<xw�ðG!���B��y�R�إS&��Ȑ�A���yr'= :���I[;|�b��yB W0R� Kb.M�)��!�GH�y�JIDz14A��~T�ȃ�y�H�6��}
g)Y)�s�F���yb�Nb�|b@v8`���ylFL��H�V�6��`'�,�y�W��*d(s  [��AW(�y���&���"j���zqB��̞�yr"�
SG`��#��f�8TLI`�<1�oqP��`��ˁR�f�iv	�M�<�``��3}@��f��@��R��M_�<aB�ya7�s`�i"CH�AJ���2��t��;|�[�mޅ>ȓ_��<�3$�5$�p�YL��~��T�ȓ�4d8��T��Ixģӽ��m��\���J��''�r ���:@�hD��JB�$̭ k�4�(ŵzhZ �ȓD��x��b��[�
dC��ȓc���H�p/ZQ�ABY ά�ȓf�,`[�@�6WU& �6͹-|�!�ȓJ���q硆"&δu:&d��V�Đ��F a�Cc�,A�6�`�Δ�$5<�ȓ?�V���n�1�$	�	����C��A9���h�VY���S�+�̤�ȓ'��m(�Nަc�&���A�[�L�����ـ6D*hsj�27�DTK�AZb�<I����6a5�[2��]�,�v�<�U-Ørb�����Y�8 !	�^�<����M!������+S�U�%Z�<i�e3$��ts�A[)��4�HZX�<q�a��J�*p�c��%��:eόi�<Y�ˇ:p�aB�L�!Є���M�j�<��hX��n�*�E�a�ޜ*lD|�<� %�f$jj��__��{��\�<�!�.~ap�k��Vp��j�Y�<1$fU�^I�e���Y�p�v��'DM�<م�O�z��ǀ7n�����E�<P���(ǆi�&��4��1�� �C�<qԥ|����̖!fw���$Rv�<�A��2�x��h�c�����X�<�`��(���P�E1XB�)��c�X�<�i�7�<��a‸{HдeWT�<�E�1�}2��_����V�O�<a�lGt�X�ŕ	+�XT�@/�G�<IaǲT�ȸ���C:ӂ
���E�<��I�OO����%AzX��P~�<��C�ۂ�(�%��#��mIT�{�<� .� �+���he��WKS�X+'"Ox1��KIn ���!*�',B�!qS"O��*�+��g�X��G6++�-b�"O0��⊌$�=�d���iA"Ol[��?VXb���&�$66��2"O�A�mQ�]�)M�m��B �>�!�d=>Z�qN�2~��py�Z?}\!�D�#�`��Rl��B�����C+\P!�d�.qZ0��HE�[�@pj�V�?6!��J�?����&��%�Xy$�L�.*!�$W�∹3A(+��9��ܦ !�$Q
A|��p��&!���c�Ǆ!��֚Q;E.�B����!Y#!�D��K�Ɗ@���@,Y!���0d��ؐ��R�4��xH��U"�!�Ӕߢ�ƅ�Rt�r@E�.-w!�䆹W�@4��e�zM
Up*�`l!�$�~9�������b/\i�j[$yh!��ѹW��X�D. @#�i2iQ#K!�d�@*M�&�P>-��Q�NW 
1!�$��V�X�k�o�<b����ؙ'!�Dϭ����k�$�t�v�	!�d��6�Ѐ I�f��<�iV�%*!�Ċ�S�4YҡŀM�Duا(��R�!��[�8Y�ɖC��i��@0g薵&M!���VONA��8t��P�u爡qC!�$Z1,���@kmb���+5!�Dܗ[�|Uh��#O���/xO!��F�Q�rD�ud˵e� ��ƦFD!��]y")Q�-
�%|h(H�ʈ�3=!�\�Y��h�턮;g>U�Dǐ�!򤚼0x����j]#+�\!�ǙMe!�V�bz�uˀ�¬}8���Gғf5!�DV�\�@lS���"��E$��"�!�D[m��p��ίJ��IjD,R#4�!�D�J{r��LYP��}Q���!��T>)���:����X5!�d��VNQ��K�' $	"j��z�!��K5F`0!m'f�8�wBM'!��A�t`Y��;b`jq�۶�!�D�j��!�'�N�(����!�8Gh̙�l]�p�ʙ1��œ1�!��>AS�8`�:h�blxu�9	�!�$���H��]>'�С҅��!�bݎ��&��(c��E�n!��/^�Y��!��;$+h�!��L���� �	�88	����,�!�D��/H�,�-8zp��JD�o�!�䈕��0�$�B�%��X�S<u�!�ǞIQ�M�����'aD�Pn,|�!��X���f�ݟ+X�چ�џM�!��1�)����BK J�F�c�"OD}+�4$BHCq!�8�h��1"Ol�9f@ϲ��ԩ�@ r��A"O
��'�8|�H����J�h�"OȄ/��80�E�Zv��o0�!��	�(��9"�ӭ$0*�$��O�!�Q�Lxt��fG�s�|"CMY a�!��|{�s�@E�a�vI����p�!򤋞
Ș� Ö(2��t�7�^	�!�[�j�h���	o,V�� ��,:!�dD-� ��J�	 q���r�!���:+TTK�O�Y�`ɰ�M�S�!���|5LHdO�#�&$Y���!�� ����q�ظV	Z�N����t"O��*�&�	7V�T�EW�i "O�=X��� '��E�ӊ�O�Șt"Oօ�U��lf�)5�X9z�d�u"O�h�*��'v��[L�L��Ȁ�"O���c�M� `^@�sDɉm j	iV"O~\)�(M�<a�r�b�`���"OXc�w:�$�c����y�"O,d��`V?1!�	�BP�[T2	%"O�h�dY�dhʡ�� ǹ=���	�'I�%q'E�,���� @A�',h�Q�l�h�"u!�yx�"�'�d�¥ꉴE2iP��`��
�'���bC��$ h:`%���	�'��h�@t�-���V�h��'� �� �_�h!uŖ:#����'i$�P&:����Q9�<��
�'�T����.�PC�!a���
�'g�|����|Xp\�C�Y�J(֠�'A{Ã/mj�Q6�<�� �'ڗ��q��� 8%,R
�'�]`e�]";E\��B9-�"�	�'�$Ԑ!�W���h�--j�,��'x���w�I�XfȁY�+��T�r�'ٺ]�2�]�[f��a �7V �"�'��SȖ�G��t!�POA "�'�da�B��(��Qg�"D���
�'rbx�q�	`ܦ���<���
�'������#�)��)�.1��'
�4��	F1�p8sFG&�K�'��TH��Ư7���s
U<�Z��'�ν!��tt���mY .�L���'54`mX+�����6r�> ��'\��Q��,30L��%ߊl� q�'��!�D�F�Ja�H��W�/5Li��'�l��Y86$<3�D�-/^��	�'�2YK���|���f�s�&H��'#l�$%Ό,�8`FLÇ6ZE��'�>����W�Q������,yJ� ����Op��0§�
�ۣDZ:<|��
Г6�T�'�2�'P���O|�J%�u����"j������.28HC䉺E�R�͗]7�(�GeD�BC�I==Bpiu��	���Q/�	,�(C�	�9&�z�@ӊ͌ �F-��}"C�ɜ=ٺ=bq�Nt��OǴ)��B䉮a��h9R-��R����'��l��?A��iO�B`�c�b]<���"I$E�S�h&��gܓe�F�PT,�P��X���	9�ȓd�m��
�GƠ���5�Ň�8��%�g��#ae� F.�&kyR0�ȓE�>��JU$8���M�O�xT�ȓ�=�fÓ >̱2��rWb��ȓV���8E��G���Y��jJ���T�����؞�i�@\<"EL��?�ӓ^^��5��5�
-q��ȓ\� Ȑq@� x	p���>���ȓ`:���Ț '�\� BJ/M,��bu�pv�Q�3�h��4G�)��(�ȓ���RE�Y�8<3�l�4����>�l���H7�DQ+c-��PӤ��FL���"�Ё�Z���<�'����Э�0@�0h)���)`�C�ɮZ\"�[���7�b�1��[x TC�	�	!	��d�>�)Q�k�tC�)� dX���ȹV$A�q�ʶ�̲�"O�|���YT= ������ʵ"O�`��G�_��)�C�/����f"O2}��j�uN��d��={�4�C"OT�[���`
�[�Ⰼ�Q�^J�<�!�]mAP���WrNS�TE�<��oՕ;
v}(�/�e4�]����|�<�w�.{��L�%��<H���s�d�p�<Y�e�\��9�d��?lV|k���m�<�A��k�z�CF����n,#e �O���,��@>y��%F4?J�=�"��Y�h�"E1D��*穕/L���k1�[13���P5D��P[���0,�4[U�HQa�0z�,C��/n�@X�\�{̼��C�.O�B�I&���(��t]�M!�,5�B䉃|R,�pn��!�Y����ra�C��	9�����O� #�œŮڙ'^⟬�	D>e�`�z��D�Dم=m�\ۀ.1D�4³�R���E�w�ظ�ĲRD$D��I�J��(򖨪��*2D PQl!D�$�u�� eU�2\���
���y"�2v^�Ԡ$��O~5+�J��yR���%v��X�H?2��HEj�2�y�GG�6��qCNY��q�gDP���hOq�lI�!D� U|� ��e���C�"O�dpQ
@p:�X���G+P�-"3"O$"�+�\
DF�0���X�"O�UB��X�R��ɂ�D��]��<��"Ol) �l�)f����������X�"Of�c�J�1'¬�T�Z	
�~� c"OR�����бo�Ќ��Y�xD{��N�R����Bo�L���9��]�!��>Q����Մ��fy섂�KڂZ!��S���:ce�qL�A�j��!�$� V��ѐ�Ί#$:"�7��7!�$�1d��VC��<�����U�Q!� k��``N���
y��־�!�D�g�.Ӏ+�)"�`��A�P+�2�)�'E]0����@�j�,�#�%Q����'2��⥝�'��ccOW+6!X���'U�K7�0=B�$C9����'�TMec�X��9� �95�v�!�'TV ��e�0b���۳d�+.�����'�r,a�"Jb@H�83	Y�z���'|��.@�T��D�c8n��'���+s���W����U�9#&�
�'�z�IQ�Y�r���3���7�zi�'/��W!U�v�PLE꜁k�� A�'`L�HA���>d���#{F�l��'�	2e�g�5�H4��GaU��y̋&/���hH�Bj�Y�����yr��6N�F I��Ǩ?�I�G��?���'J��i�^}�� 5Z���t!\k�<A�D< O�-#Rjͫue^��7D�c�<9�����n�*�o�L���&g�G�<Y3��2[�8�	�5P}NdZ�A�<��B�q��tG(c{"xB  {�<���A���	�,�����%�x�<Q�  �-�$������r�(��q�<����bl�xp���9��4��E�n�<3�Ͽ�J�2��-C�����j�<qe����!׭5jK�bK	f�<�"��;4j���¸iJ��V��V�<�䪙x�Hu��1��ݺ�.T\�<� ��" FP�9�Ty�5l��w�b@ Q"O&��$�� �YzKF�(��)y�"O�|��Oլ��Lq������Q"O�$22�ݭn����� г/D��J"O@಄�>�<pzr��?"��t"!"O.��P�̅#
����ŋ:�R�a�"On�k1c�0hOh�rg�<(��(1"O�� ��V`��&�\��"O���dl0%ۗNu6�iY!"O��h�0o�,+��ӏ ���"O��"�L�#h"��K̠X��YV"O�5c�PE��H{j^/Y�Hc�"O�pxl[u�dhPF�Q�*Ժ�"O|,R���o�4���G�����"O�u�D��-�@-	UB;8h��A"O�`Z�aEK
��D���3�
r���O���2���"!o��5v�1���ص�N���%��i88����N\��m��P��Ș��53\
�����X��!��y�t�D�֛	�B�R��*)q�-��:j8��ƀ�<d�d
�.'zj�l��'���Q�K�2M����j3r��JP�!��h��D�93�oO�d��0�?�-O#~��XK����	t������H�<Ib��Eh�Q����B$4���j�<�צ�y©��͇�l�jۤ�EQ�<�ȃ1B���u*�1��ݪqL�X�<9� \$Ei0�y8�z���V�<�T'W�>
ʵ���B/lI9QGJ~�<�C�U
����A�M�z��$�TO���?���ň�b��cO	�T�A�'KE;�&��"O�i�D��
.������[�]��Ma�"O�$ѵ�̥d����H�A����"O�-���Ȁs�J�s2�89j�"O�!ff��.���EC
Eiy��"OΌ�U#I�_���C�֒C3teA�"OV�J�"�"%��<[Ċз	-�`f"OR8T�6Ÿ�Z ��2�P� "O�Ak��K�|A�D���R�D@!�"Oܜ���܉���Cd�$�g"O�H����(u�\�s�E�vn	��"O��ë]����b��N��Ʌ"O�%-R)%=H%���@Y���;�"O�9�qN)q�9Pˋ'0l�aA"O� �%�2�-Ѕ�];�N�U�|R�'�az"'�,ph�V�����p����yҤ�$/VP�Q��&�|+����y�-�I�d[�E({�YY'�;�yR�J�{������ku6]oJ��y�g�JN���s!ɏ]n��S�	ŵ�y���25V�1�B� \NZeb�-�y�AX�4tZ\p%��#D�ROF�䓥0>	D�7���Qև�c�x|�uJ{�<W!�{j�)v��	o`���'Xs�<��'?i�!�4+�-	P�@ K
{�<Q'�v	��(S�|w�(H�u�<�se��D��p� [������J�<i���:̜D�A@Rlơ��A�<Q C�kG��P�gV=Byv��`�	~�<�4IהX���Ygė6k�B=c��{�<iH��	&����C�6F)�y���t�<���I�X��h��m�R�ҐH!+ Z�<qA�+K��X�Nź��a((�q�<a�Yƒ�w�
�bڌ��Uw�<� ���	\y���z��g�2%��"O0"�d�n	���GMkJ��v"O0Aڂ(f�ɲ��>DёR"OF�DE�6u&hS��R�Ftb)yw"O��c�/Q� ���k,L-
�q�c"O�H���!���Q�/�����"O��X��
�>�*M1ʃ)��S�"O��8 �0/T�J��E7t�Hp7P�,��ɴ]�J�Ƈ4�l�сF!��C�ɉYU��{����pe	c��C�I�O���XbH"AX�W�.6^zC���,��� ڼu9�����̄.��B�I�6��qq`��#d�9`l�,_��B�ɂd���c���OT�����"Y)����g�(*�����ćU�%�h��8D�,ʄm�-�:���KR�2�` ��5D������2S#2l)u+R/]���hp�&D�\���{<q�&!\�?3����$D���hG<얥&�@Y��$D���  �w(��#,V��(6 !D����M��e�`�q@�, ���
?D����?k�l�!6I�-�ހ�/D����)<(Ķ ;�KH�}�l���.D�X&�ٔP����c�)
�����-D�<;a�2բ|�oF�R|xz��*D���U���	yn�H (EBh��b@,D����Q�U$���- �A=�}Jm4D�<Ah�4i�~,��X�Z-���&�O��d�i�B�L��@����R&�	�ȓA��0��N_8]X0�;�C�,��ԄȓNDzz��C58q$�;p�~U��+�Z(є�?$��(��7hm*U�ȓit䉻v���Qx�����X5���ȓ
�]��,B�+��3E��2cؐ�ȓ:RƸ�4o�l�Y��g�� �����I����I�<�6���p��(hf��We�B��I�<��L�$����g���W��l"�E]�<1U�ڔ~c�݁�n�&R��Ѣ.�\�<)�a�V�&0�Ԉ�1o)�I9��m�<�EgK2p/�����2A��!��u�<!�CWd��L��'�08����&�q�<��Z���pht�N$j�b�B	�Ex���'��Pő�:X����gO.Z�^ #�'{Z���ǉ��(������W<$��'X�y�tCD��\Rd�I�b��'���蟶9��T)�([�x���'Le�e�RD�PX�cC�Ԩ�'2�����t�U�GJ��R���'4D I�A�a*�X�%�$E�Ɲ��L�H���KP��z��W!d��݇ȓ�xq�s��ee�ݐW HqX$��:�X�2�#�~$�V���{b�Є��.� �,���S �	�t@��U����h�Ly�mS�h�`�ȓb�EJ�&�U<��=��ȓ	C�=
��I�v�*'�@�����ȓ�Tإ��u�TM�@�d& |�����c��	k����W��z���$��,a�R�n�"m�v��H����Z&�;'W�d��ʔN&M�JЕ'�a~�Iϛw����O?`ϖi�c昚�y�g�3e,à\�OjL��3d�?�yr�Y��lk�A:���q�@��y�-\'A& ��b��2�b\y��E	��d�Oj⟢|� Ɓ��d/y�@�RԤ�-�,*�"ONR@��,4�3��CY{�	�""O��cT!>�arD��Ef��"O� �� ��%���`,�o�����"O����@1NڒD�kg�`�X"O�x���+)V��L.`�\�R�"O���S��2))�	�> � x��D>ړ��D�3xX��ڄt���yA F�Y4!�>桠�
�W��p��ˎf!�d�^n�k�&�?U�j�Т� �.���'�a~��J)C��أ&�� E<�+V؁�yBc�%f�ډ���K�S?40q��ݷ�y�չ&�
<`T���PӞ1걉��yb(@�1���`)]�EL �с�A��hO*��I��~�5	��	������!�d�
8�K0�D�cLa�v���!��8d��L`r��.�^9�p&��!�D��L��֪M�v�.T�4��+]~!�M�!���RQ�Eln���eC�/�!��D��8"�i̝Wax�@�ݸ
n!��[�_�	i��K�riq�8 �Ox�=���
5���v�d�mX�@�VxA "O���2�������b'.�ȷ"O`U{��OB�E�F\��R"Od��¢�8�U�-Q���ʇ"O�-�Հ�%
��d���VF���"OYZw�Ƚ&��#�f�*T��I�"OD�����L�qY���_�D�#"O�s��Q�<��l�7P3`Ⱝ��"Od�q�O1.2-�W�-OB>��G"O�}�g �)����_%z�c�"O愻$i*aP�¡N�!rb��"O"���F��>Jb�rB>8S�la�"Ox�ke���U��p�a��w�8�"O�q�<#VV*�O���y�"ObX�G�E�2x���Ņ-�`a�a"O�V����������o�` �"O�XfNԸa�X5 ��.��Ы�"O���+~,����n�1a����"O�IQ��>K~d�Rc�L��Tz"OX �@�0 H���ޜU�r�C�"O"�xw�C�-˶���6�4%��"O�(S��AD2Re�ٽd��0�"O��A"]�h�� 9��)FBE�"O�!�nS�9	��B���8�my�"O���+�zh�#�oTA H)k&"O�S3���=��������C
2��"Oƭr2�٬'/h�p%�#e�� ��"Op4�@/�-[���A��%Ҝ�
�"O�S�R���a��D�1"OгũW� ��|:��σD��h��"O��Yd�����w��0�.��"Ot�;�Ǉ�1�
̀���?Y����B"O���FA)栰PL�Ny��&"O숑d�!w$��q`X�5[$���"O���U(۹l7�0&m�}<�Ix�"O��rf��,�OKֱ�r"O��p���Lq�3���f5�tXV"O��rc�l۲	r �C�Y2lQ8�"O*�[�o�s YKi�0"2mJ"O\�ȴ�
��@��f��>�#7"O�Z���+e&"I���
����v"O$���n�<1Q�1Q��Xjt"O�*�g��t�f	;�#�<w@@�d"O� Q��g�V�� ��A_�qY�"OF,��Aڲx����g�*+"�x�"O��9惞:��P1��@��^��"O>03f+�*m`B}��Ř��D7� D����W/����H�"?l�I�m"D�4cU��8H5�C�XÚk-D���2녫b.���@N�;W���ɴ�*D�P��E��y;D.�9rFIե(D�����ptj��]��%ʜ�#!�dԺk~ )�@�·dFN�HQAQ=}�!�I����A��92J0ء@I�-�!�d�o���W�ǿo� ʗJ��!�$D2J�*)F����R��!�K�4�f����W�=�f�r�	�!�D	�F)���	�w���8�LD/n�!򄜶�n-�W�G�G��D`r�˱�!��Ly@.���JX'Wm�(�Q�[l!��"�R�dؠQ\��;b�]�!��@j��@�L^!ONH��5�Y�[{!�(	���%4���� {�!�M�F�xQBCމu�n1��x]!�ĔJ��h�#:���#�V'Z1!�dM�kҌ��.L3_��-`�&�#!��?�P��D�c���Q�E &!�1��+Zo�n�бNR�!��>�:1P��Ύ&R��Q�l�-�!�D�(���4��'.�m�Pl��X�!��s�p�D��L)80�Ʀ�!򤛲U*.�"�.u��x���=MX�C�I1.$�أt�@	aw�5cBØ�_��C�Ii|�=j��Ԍ<�!�'"�?�C�I�E����u�x���߲V��C�I�u �yQa&�|�F�����1U�B䉫!_���.qL��Ǉ�dxrB䉊H�
t�E��<e:حkV@�>�lB䉌O�.�
��XS~ĽK���oJ�C�	5rȍx7 P��^]sc�˷Nr�C�-c2J��I�B�2�Y� �&^�tC�I�='b������N�X�Z����q�RC䉙\���&	N�$J]ʑ� &2fC�I}*B1�#�D��x��BU�JjB��
zT��%��[�P��"O�RN�2?��$�%�7mD���"O��s�jֆt�Y�'�E�j��b"O� +�
���`��@
�&hXM:�"Ob�0aL�-���ToT�R*t��"O�A�Ҋy$�`QTI�~b\�w"O2i#���B���(�G�>B�]R�"OJ��_�2�p 4FK�uX���"O�!�P�ZR�=q��R��y�g"O�9��	�t�����!z�l�؆"O�|�s�]�|V�G:N�
��"O�p`�IY�}R鐧�A���$"O��0J�:o��a�GVi���2"O� ��jS�+Č������`��As"O@�Ґ$B7b)�5�0���'���*2�'�'�B��>!a�X�<(�0�Y�1~<2E
�x�<�SF��j��Q��2���#�u�<��	&yx@��(Գ+O����V�<yf
��|�,�EN�/�@!�mSO�<��!K:v��erC���[�x��E��D�<��J�y��R�٩-�\���
@�<�J*wr=P!J�;�v)��~�<Qs�Xf�}�Ɂ;U+<񨇅�y�<� ��+Tc
������m �=���s"O\�8t��9=�ᰱ&�,<&P�k�"O�qq�ZB���AS�=�$"O�5B�,�S�~teɌ*.؄��"O|�����:S�5�v�K���2"Oh4롊@�Lj%H�r��3"Ot9H$�ˤ$δ`
Pi�/L��څ"O�8�'����D�"�K'�( �Q"O����!]7�QÇI�R�"O�)2�Ĝ�^��5���&K
�ٓ"O�бc�����F�_`����"O&��BÏ�g��u�Ȑ�A6%��"O���5��1���皱w����"O^�sCoY�Yz��YUg��HFY�"Oj��f��a�f�a��Q,�!�"OX��"ْ|�� ���*G;ؐ1�"O.9�ǖ�p�ū0��0���"Or)	5-G�tMq�%��G"O.�;5̞J�"���ܠ)i�"OԽSĭ�=<�����X (�6"OT%��d�CV�S�쌸j�= �"O&���Ϙ[1���j��y����"O�|Ҁ�h��*�X���
%"O��Ti���T����[�A t"O>���_T� G,�&��II%"O|�ja䁐j ���ʇ�D�j	y�"O��2F�ֆg�Ȥx2G�0�(�Q"O��AF���_f�ak�*4EJ�!�"O(,�*:&�D��P:
�@X$"Or�+����#M"�8vcAI�zEr"O̴8�O$P������1]��Rw"OtU2i��ZR�D���A}�zD�"O��ҋH�[��:��T�Hqc�"O�qPP��=>ߘ@A��)�N	��"O�t"F'O#w��[E��y��D�3"O���DҤSB�i&.�dv���"O,q�
�*-j񀃂CYj�q��"O���T� `b6�[�yp��ۓ"Ov�"V)��.p�5Z�Ŗa!zb"O`ui#\{&�k㪈�bRR��"O���cDJ�^��#�g�3@E���"O֔[w�=ԁ*cF��WAưK�"O�ЛhW-�e�d>6�D�'"OХYPV"\y��r霅"��B�"O��TeF@�\H���Ão?���""O����@�"9&DrV�3
���&"O�Y�Ӌ�^�P�����&в5rR"Oެ��+�,5V`C4�)�d� �"O4!�M (�j��/P<�8���"O�A	uF	�y�x�2,�"n����q"OR����@�X�	S� ��\��"Ob�zV�I_V��������7"O6�� �$eEV����J�^� "O
��C
�Fp�`�Mӓv�p|y@"O��ѐ@�Y'�Չ��Q�KEr!��"OʙӲcZ49|�T��K6_�%R�"O�țB��*R���pNI[Z|1�"O$J2m=X�4I��qR�T�p"OD��4�ɹ��E�m�6:H�� "Oȩ�6�B��|i���J�2��0"O���"N�ܔ�eB�)HՒ��V"O�9�%N�J���c��9�f}i�"O�$3ǅU�c���p��	/�.g"O�a�G����9HT�#j���&"O� F0�m�i.�h��_T�@aI�"O�tP�C�ď�A�Y�e"O��b�.J�=��+a䛡5qP""O,,R�J��-����0K1��b&"O0� ���Gr=���m��PX�"O� Cs���;pd���Y|@D�#"O.�c�%{�xaS5�� �U��"O�Ē�,�Mv���!$A��"O|D��,i+ !��w�ڨE"O5��$[�+䦑*ԏ$d?���"O���@B$+��Mx��@�A��� "O���H&?�05� �(8+F��"On��D�ǥB'@����:z�H�"OHZ�E�m�HX�H��Q�	��"O�fG9	��9�F�=.���"O�Eu�G,Az
�d�@/��0�"O�E��lQ 4�N"� �`��"O�I�G4B�<��!մ���"Ot�Д/U-$��]Ɂ!�:~$"Ov%: 	M�|�x�!���**�J!p"O�𠲨�q�����7�8 �p"O0HǮN =��b��պ
�v�"OZ%{T,՛5(��rƄ�@k�T��"O� ׏�!z��c%�A>���"O��B�a�(l[t=�ă-(2�Tau"O���� ~ִ;�Y�!�zR"OV�X0%��ab�-9�]8;/����"Oδ�T�5 �jG��HoJͣw"O.0��#u^�dn�"md|�q�"O���u�_�BUR����	|X�0"O�%�n! �u�q�%hV0Ա6"O49S`Ç�	�&��_C4X�"O疴�B��IװZY�a�"O^�S��2-�Xq0��H�=�%"O� �g�X!Ct���65�Zt"O�1g�-�4�� ��.(�"O�x�ĦC���
Jt��%"Ob-�$I�3TJX(p�I���C�"O�D#�# �*Q�G$��t�"O ���	;v@-Pn�����"O���edǣW���Ҍ�E��B�"O�!��ںH�ܳU�'"�m�"O��!"M�p�pykSǮD-�U"O
0�4�{�Bo�L�"O�Q8 ��	0���j�m_�A�b�H"O��X�W� '���$7M(�"O�i�0g�&@#e�ˢV�+"O~Y�0�W��)�U���|��=�A�|"�'g���1�%'��	�ΕMff1�	�':���qȕ&F:����:V�$�k	�'KP�7䆪Ob�4���0R��]��'��SSL��rN0'��K�.�R
�'s�ى5��(s�<��Aqx$�	�'���� �*.p�]rT.�7C�5 �'r���r���@Ϻ�#�/�?���K>�
�c��ܣ�K֎��FEY�[ ��3>��U�ݽ����̀) ���ȓ`��I��1m�j�"B�?u�J��ȓe=�-�$�?*�Mqf�>>��!��p��Y��#<U4���ȱ� ��W���b�<]Ԅi���)U,���Ed���d�Z��yi��ܧ�d �ȓ���Z�@�q?:$�DdԊm��(�ȓ\�" v��c���@�炬r2���S�? "�P�'Y������#Ϛ=��Ī�"O�	��ْ���RF�K�/C��t"O:UZfm��n08�� �v6���s"O�B0�K6�٠�^4"�3�"O�pG�W�Q���+Q���I5��"O�����;"����KׅxX$2�"OȽ�#@әH�N�P��]k�Yk "O�3h�(0hY ���<<�qzV"OB��&n�'�rdQ4aW�h��d"O8�@�-a`�Ж��5-"@|ك"O�ap�H�7���vN� �U+�"OJ�3v�?42�ӊ�\�4��"O��P����a�ԧ	vø�r'"O�}Sw�F�x*�@� T�"w"O������:��1aۀ[R�e�"O��b���8�� ��^)6���"O�(�5��Z]2e�uo[z�@"�"O���u,A+.\������Ig`u1�'���q0�-�.ē�7 ƌ���	3D�(���9?��&�ۜ �e�1�1D��C��F4?�%$�s�1S���	�y�&M�.>�@XA�K�RD�rv�1�y2Ak �u��'\�N��@�B�Ɖ�y��I'B��kH�AT�ٳ!"�y���+@��X�k�&=�h�Cϐ��x¡]7Rp7�N:d
�Ea��&�!�&N�TPVa�� �)ai*`�!�DH7T�݋��X?�48�h��{\!�$D�f��)0P!�?m�<��)9A2!�NBw�#e�׏Bp�xҳ�SF&!��t�J��%kX�4Z֕!)��!�� �{�<�g��::jh���x���1Oj�P��O2v���I�o�0��"Ol�A�&�8{bp(�(,B�)(�"O"t끅��(���bK%K� ��R"O�|#��S![��@Xfg�@�N��"O���D
4(��`�����k��3"Ox�l� �qf#ة	�Ԥ��"OF,b���⎽��"��u
"O��JE��2�@�	ʦhQt"O0�����k9А�ԏK1.���"O>���Ρ�	��OE��m�"OKF�>���3�E�d
��K �L6�yR�Ɋ^^^�K�e�]��%
��y�a��xS�nR�b�3�cK��y�؉�TCw�}�2������y��V8bNw����_ �y­��l,�g�oi *!�L#�y��O�R�����jG�Pjp��ʁ�y�D�t��H6GR6��A�W'�y2�˕~��"���'��ţѥ9�yb
ڼg���X�
�	B�۠Dߎ�y䖌?*p4���ܜ_z��`�!�y�W�9����u'�+4V�� �@�y�%�0� �0ŏ�niq��U�y�4	���)q��H��,rɕ�y2�� ]���aJX�m=�q�v�C��y�՚Kb�|q��/\A�( ����H�<9��`����Ջ]D.�ȓreva��� �h�2���)Ȝ��6����Z6j��f�w`X��ȓ����`#.���Ĝt�8���iVʕ3D�ԖX+1� E��d�ȓn��U@��K� �G�G�����S�? �);s�ىR�FU��h��	%�Qȁ"O���iJ(ZX�$+�ߧf�!R�"OF�Q��z)N�[�k^�s�VQ��"O�Y�#�̋@_��j��
>a��b"OF��@��W�,Cb
Ee�����"OșdF.��<BlS1^�N�t"OܠPs%W:xh�%!�l� ��c�"OR�` �Z
	�H�s�I��r�,�I�"ORՒ ��k#��ZT#�^pbذ�"O �`]���yyС�:j ���"O�1��@	+l�@g��b����"OYW�O�R��yG�� �D�*C"O��� W�JB�����ԕQ���3v"O�p���)X�%J� P .�X��"O
L`�K&J�
ШP/Q'��j "Ox�U��1pT�MX�/W�&�F��"O�-���ݼ4P,�D��mwT8B�"O��ǫ�E� Ô ��[P�X"OH!�vj�36�b ��(ƩkCBI��"Ot�%̘�9s��²g�+jasA"O����^,sZ��� ���d"O���P._�fgi����H��"Otʂ��f��p��S:/e�&"O�-;��[�n�|�C��l��1��"O�8�"#\�m�ހ�oE�v�t���"O`����F�p�C��C����"O�1�j��������\N��)f"O�Y�cK!,=�e���\��}I%"O�`@�_h0`+w��Y����Q"O��ض�؇Q�D�чF�s� ܪu"Ol);&�� /��5)�̞���"O�m�%fL}��Gk�- R��"O��H���i(6	 ��O�<��1w"O�±�\1o��ɸ������`Q"O
F���w ���f�4���s "O2q��#Ǝh��I�4c�Fd�Ҕ"O������nX��9EKW�xӲHJ�"OX�U�Ӹs�b)`
�Ϩ�0P"O昂�e#6e��3cT*_�م"O��3�IF�F�T���Ѝi<|d�%"O��� ���U��4��"Q"
#P"O��F�c�����f�B�X�"O�-9��Q-aFH��l�J�:$ g"O�l����HHBv�օK֌�05"OE�����h���Sv��j�\̨�"O�Z���4�fu��/��\c�"OTU P�'������ Z�6x�t"O�9��9+���ňBKL}*�"OⰂ��+�1�3:�3�'���EF����,�P�(>�<��'�u:W�ȏmc�Р)X�;^4�[�'�F�SA��S�)s�!�=5��ɚ	�'xj�A�^�h�u�;+�4��	�'&�����+�$�H&e�>L���"�'ʄ�d�Դm�Xha�LB�Iun�x�'����K�~=�Y���A+^)�	�'�R�!Pj��5�ޘ*���:.�J���'+��o�Q�[�|TKa��U��'/���!�E�!�ry�'�Dd���'"��a�L�Vic�/� ,�|�
�'�.�T�UnUr����9�	�'�̫� R�r}��uGHuC	�'����d^�F̩��I/g'�ث�'���B�+82��X�)��Y�@�8��� �|�+JT}����٠m�င"OH�X�F�9�vMk��Ro�x�`"ON0	Ł�� ^��#DB|�|��"O֡����@���C+�:�Ӥ"O���c̥E�Z�׆Y'."O�`!��h]���2�\#"���V"O�ـ&/,I�M���,X*��a"O8�f�ɖ5�r9ZE	J+ބ��"O����0��gƟ<;����B"O>��. �ri"0����h��"O�9 ,��'���"c��8؈��D"O<�C���% �D��s���,�$�`�"O��KA��c���QE"�=	P��"O�Yr�oE��s!�J�
Yiu"Oy���X)oj� �7!�mި�Q"O��y�J�E��F"�o;�98f"OjX��f��U��k�斋 ��	�"O�����
c��J�.p8�"O�@CE�Q���@5�Q'89#$"O�9�u�V�+6�Xۥe�?i�!)"O����l��T����ì7�����"O�H�$I���y;&�����s"O���ă5�֘"@���v�r"Oށ�d.]�x=�D���!7��z�"O�l�ԗ.�2ԑV+��>�X@�@"O��X�*N-;3�k kB���:b"O����a?F�����D\Q�"O0���3uO,���.�Eh�"OT�5"�4&�dL�6G�w�Y��"OI�+\�ѷ ݣ0�
�i"O��3iD��IpT�N`n� jt"O�x%��[����Tm�.Y�"�"O�y�$�J3�T��NwT�i�"O4ɠ����LL�	V�*fj8I9�"O����xӨ�YCG>��� �	1D���g�Q�as�U2C�!_���"��<D���"�G�/y"�9ϕ=�t��ą5D�iF�6yjĳC�)Z�r�j4D��B�A��J�!I"K��E�α�4D�@��`A0I���`��Fm��%�d<D� � J߮*�ȸc�����i��9D��:�nC�~m��w��71oؑ�b7D��A�4��1F�Bs�U:sG3D�P�4mٻcì$�2'U�d��jq4D�4ɡ��)}�B�f�my��xw�0D�@���? ��\��E�'*p@ Hg�4D����BB��^�a1*A�B�>�2â%D�
G�ݫs�N��_9�8�K�o1D�8�p��zY�T�^)��Đ��-D��#��ӷ3�4���!��p�s�+D�D;�ʷ7͌My�΃-?h�,/D�hxv��<}P�ܩ�L9� �kD�,D�Љ�b��I�Ƙ�PF����U�D D����oU�)�T[�DI�E��UR��(D�`�¡H_�Xz�b�2p�\�J��<D�@Q2b�'��q)AJ��~  ��j;D�$���'.��1�u"��F �1%/8D�8[�
\f��ؔ B''��ca�5D��!�ʍ')�6\��!�N�Jp��I/D�TI��a��iP�D��>�:��(D�x�ꈿJ̀J�<Sg�X'�$D���an�)#��fG8.=*�s�"#D�Ђ�\q��蕦32�&��6D���	M�j#BmЦ��}_^���(D�� ��Y�A#n������GP8�a"O�)bQ�E01���j�CN~��Q"O%ꇋQ68�^̉�a^5i�� �"O���W�he�B�P	o��ܹB"O�5Sq��9R���H%����<D� +��L��t��ѧp�P��<D��s4sV]��O]0*�����&7D�`�1��1BN\�G\)&����J*D��8eFM<-ab-+�NZ�2�d!�)D��ūW�^�eGbR�l\,�;1�&D���c�	f (Q�5"�_j��� D���b ��&���r��0|Fc�"D�l{� %A���R3��#�J��>D�$
�hO�`��2�@��s������/D� ��85�PT҄拣L�ȉ8g&)D�����H�z>�)�/�4bU�A�'D�|Sb�:2�%��2P(4H!D����G��\f�L���0���4�,D�$�`�N `n�(T)F�*��̢��<D��y�%Q�(�9�G�sa.�q�<D��9�!դl�=x2Ƈ< ��k:D�$8�GB�\�ȼB�*
a޴�4D�i��Y��6N�o��@@�%D��C0J��=� �c��cN�QN!D�$I�$͇6>��3$R�/<R��#!D��Zplө�6�$�ĭ%�hQ�w+!D��c0$�>ɔ19vLC�3j���t!D�|@W��n�RM���b�(0 �=D�$��i�l�h43K#�q��<D��4�n(�UY)R� dx��>D�p�4(	��lx���Z���ҡ�;D�d!�-�d�L�����B�P!�7D��R1� �����?da�qs׀;LOH�@�7��34�XQ��A��sF���v�;D�L�A��)�  ���@�"��m�!'�IF���ON��XV�N.\�*��W�P!��'ŢMX����zd� ;��N�z��M�
�'��]��/p|d�A6���\_�,��'	T���Y�IdA&Є[�(�c�y��)�ӑF:���CZ�F=TX��M�-q C�I�k?$`�	K�LP�8��)9��C�	�IE�9�qL�|:lY��lC�ɸR�࣢G��e���{"�Y9�pC�ɭ�pYqU)�.�m���2Zd��'(1O?�	?gr�2�H���9����Y�JC�	�m�j��T�'S��UT$Ԙ�<�Ip��໔ϋ TTB5�
�;]��� 1D�T1�o	�t��؃��g���e:ʓi�xˎ�=���9��� K������y��]*v"�M�|�Y�с�
E��i�|FlA��&�1e�֙Hg�"��	I���,�ɯm�-�Ӄ�@����󄁹b��B�	 /�Q:�c��բ$��W|���u؟�i�����=�1�����)5�'D�(V�j�Hw��,Yt\�P`(D���U�^3��}PA/U	v�ڰ$&ʓ�hO�&Z�����X�X� (#��RB�	/\\�Aj�
Z$D6�Cb�ϭS�����.�DJ�L�
 D�92� ���u�!�R�ԤI�+"]:��4:�B"�}�'����+�!�&��'a��%�x�� �)D��(���~B4ق$��zl��E�&D�abΝ �|l���J�QMh�&�/D�8� �_.���֕7�F<yv,-D�� ���2դ��!��t�"%i�"O�!C
�[�.�z4*B��
<$"O�[�aԾ'�d)׈*qX^�8��'�(�<Ad���sp�P��	?|��8�HF�<	�8z���@��$(����JM~'?�S�O[6�	�A�^�r�ƋD�1��H��)��<��Ʊ�΁�C�K:sn^ ��RB�<q�ᔚ�^�Q�+W�I�A��ʔ�<�
��,$8�Z@.���bcم�FX�$�O�3R�K�)}�5�%E§Z��@��'��'�i�v����`�`cW)F� q���'�S���C9K��Yy�E��|7�Уa�X��OF���k�-�d��fj�@�|�q�DyX� �O��9U΁�0^j����p����7"O�%��ގ+��	��NNF�4%I�O&Ͱ$/� Fn�8���70�yy��#}"�'������,D��݈��++�X���O������}�j'�� / �CP�D?C�a~U����ꏩ\+^:�H F�Z��v�>�
��P(&$��7��dB�"
���g	�p����'l$��'���
H���ӮeH&��[�PE �[4w;0�ȓTAf("V���/j8`���f���'�a~��>mP������qT��а=9�{r��_�i#��ݰ,[���D�	��y�b��+@p���0k�y�G�D���'���FyJ~UC�0`c���R�����`9&�UV�' �O��'źl��"G���@���WB1Dy��Q�ܪ��%���`Bǀ2Yݔ���g���?i���CRU���
Ul�i7�X8,�V
Oޅ���?#�V-#Ü	Щ�|2�)�Ss �LIe�j( ��z���'&n����|m��:�,J�}, hs�y"�'�,ѺצT�t��E	{��k
�'��X��1�v4��ũ:N��	�'�>��6�L'h�~PZ�C��5�ޡ��'0��@"Q|�4{Ҡ֟*8%��'������YX�P���ة�	�'A�Q�#�.<[�0��w;d`	�'�`�
љdxȅx���Eb�{�o�'<�'�� ��N�"8�
�K)"��
�'�D�(�#�#y�(�_�Hٖ�u"O���e9>���ҧ3*\IJc���'�ў��,!A�<F�
ё%���T�RX8"O<1���x�&@s�Q<Q�T=3"O�ݪ��-3[jX��F!z�޹C3"O4p�2��7 *a��F0e(���"O�h�q�S�0%KkL6y���"Ox�)�b�1V���P�I�;θk��$8|ODZ�(ג(cؙ�È.Hn���"OM�5�οc�\a:#h��+�yqP�'�	D
4��a-��%�Ш��iN�*����q���qJ�5��{��]�g�ȻM>�������|����0$� � (ɳ"O�i�'��*3�`1C�X,m�*�PA�6�SⓥS"�d�a��Q(��Q#k u�jB䉰 �>�u�SM��yc�n<�C�}"�i5>�C@��V��9J�M[tM�o)����f?i�� |��<��ů?���Q��M[�z�Z�RK�4Di�Ӹx���_�O�h[�j�p?��j�d����,�١FN�e����!D���'͈�-pʥ�QbȦ���C�=,O����Is�
W���Hءe̼8�p5�M<�O�Ϙ'�����%X���kg%��7��MQ���1�g�? ���`��:d�� pQ�R�a��٩�:O����� �慪e�>����&+�44y���$>�ĝ2$�+ٽ-�2��K�[D�~P�d�fعl|X�s���'�L=���*}��'�6�S3V� � ��]۩OVc��D�T���lU�U����8�#�eΞ�yR�T�s[>��eC�-��)���'�ў�	�䂔��y�B۠_��"G"ON}�!�Ʊ?����4��*^0���	g8��A��\��$�!ԩ�Ah�c3D��ذ'
�p1�y:��71��9�2�(�	a�'�N���'֒�܀s�Q6=��,P�'�EyZw(�'~��P3��!�S��km3G�!����`�v��I�r��w.E�l��I.�yR�/ғV�Pa���(ƈD��-WO\$�ȓ$4&��#��$r�V��)W#�6}�O�=�bE��(�Gb�C�АbJ^H�<��:`�Xh3���		���)�o�Fܓ���hO�%;F��2����L/x�O��Z�b9�X��.�E�"����6`�!�D�51I�SFD̢m��LPw����'��'��?I�Dd�"�bAJC��)&�aT�.D����d��b��AwANh �G�O�7�<�S�'��^!+d�2�C[�xp�uΕ r�!���`��0U�?�jq�U5=��o-�|�DؖtoH<�a��)#�y� hӶ�0?�,O��1@�Z���X�.A�W6!��"O���-�;+����gKD2(��+�"O�� �'l�}k��N.
�f0" "O8���LUdy��̐t�"O���&C6��5��J��b�I��"O�s��T�y�9s ��e(���"O��sASB>4�!��S1C� ��s"OT(gl��\� `¥�7�Q��"O`L)2�/aH��Eg�&���"Od!�W�s�Q��E�	w,}�t"O�e��Q7)����پ���!�Ó\uԩ�fɑ�)+�Y �ժ!9!�$���p�I�`O������˿3!��=��@R�J��߀{�,��<!�K
{6V���-�*�}SҊ��&!�$�CJ�k�	I�P�0�)���q!�ѹ+&�	ԠE&D�
�:D�`!��ϫ	�����#5.ʒ���<U!�$���֌�@�E)t�.�ʆ*k!��;y��H�R����ZL;׎4cb!�-p�qu� �<�ܥqQ(�7jI!�d
`�L�����$�28�pD(:!�DZ9:�8p�!��{��t��E!�dA�Ww��J3C�1O�Xc1�	�p�!���;8�����;]d^����D�0�!�dŪM�p� �&��uKv���
�9.�!��N	P����/eI|��)ġR:!��@v�LBf��n�\�q��<_�!�dP�`Dp��Ð_� Չũ��!�D�7ij��)��A�PD�v��?�!��'>�[�D��S�� �Vh�>W�!�d�9=�M�#H��w�T4҄M�2�!��	1Rk�5���	PE�����H�!��9��)���i;�t+u�	1D�!�d��Cdlu�B��>u�V�7�!�$Wp�dʥN#�
�Q��%J/!�H�Ʋ�����l�FY(�g��9�!��R;êm*͎� �Zh�F��i�!�� 4���&:rVѹ�LT�!jp��"O0�`�䕃l&��+˄�s�N��P蒌AF@��J9%�R�A�'�&�PnU��"�5a�.�@��'�*��4[����eQ�����'Ȁ�#�
ϫ�N-�U H�}U��[�'h�Q��ނ\��6���jy����'���"��5C������:g��9��'�1�V��&��!�^�g�T��'&�������9qV=i�ԜZC�I#��"��^|!@�̀��C�	;3S���F�A�%��1m�� q�C�xo�$�GW�:�=s2/� 0�^C�ɞSY��s-J�NΑ����7�C��0����BtI�hh�NI�*C�ɒN�0eqehAL�Lp��:*C�	}�ܐ���˨:�oʔz�C�I�s�b1됎��8�$�¡L��C䉿Mf��� ).p�؅�BڈB䉯(\P�,I�d���P��(	�B�Ɏ����Ǚ�0:��J7�X�	/�B�I���Ī&D��c��ʦ�ܮY^RB�I0���2C�=Cf��#�e�(.��C�	2�x�g�ʚJ��'F�8��C�8��Ei��ܤcq�2�K�	ntB�I�d>B)y�j�h� ��d�/�C��&8v��1eT01�Ԡ��'��Ms B�IZ�a�&� �`��NB�I�p�j�1GM6og�l��`� !�$߼pݐű$�֢5|�i���fe!��'Rc�)(��3|
����Z�W!���7<�� 5+	P9K���!�DM�i�x���W�,�|���ϋ6/��~���5��q�!dF�OS8�9C�.s�T=Xe��u�<IA��4PTL$+n�=�E�S��Z�'jV�rmԕ���~��L��p���m.N���Ya	�W�<1�������+kRl��b�#.Lȑ*\_z����Y?E���[��@�,#[@U�ҌD�i�Ʉȓn�HA���H�q�dh���.Ԕ��:��8���'I:���� ͉��O��(�-��O|0*`�C�S=�H��'��1�
��N���u�hY�Cʌ	B�M��oXI�'+�Ȩ@`V.t �lK�"�#��I�r��"�Z��с��X�H���\�Ӑ8$�u�S���M��a*��B�I[~X\:#		K�t����葵G�7�����J�&U���+�g?1��x(��s+�':�p��L�<��%�$Bm I+#k�
\"���B XZ�D:��R�6�����a+,,��;��O�|#�o2k�*�!A!\76c��'24 ��dg�ę��޼�rE.ƥK��]+e� =?���Q�ȠV��~��PxfHa@l�u���C��4��'��1�p��J Z�����r����>�8�Æ�E*'�NKA�Z�G��B��?=��ZqT2�A�5�� _U���à)\iQ�N��\4��UE,�'�~�o	�	BN��㜠G-T�Z�n���=���X���]�ȁ�7�G�{���U�	:������(~�v4�W^���c/�̺+���ã�؉q����]�eA��D5sKqO��s7ڸ'�]�qq'�ŷvG"bA)��4V<QK��8?���q�)� 9x3E�5�p?�򈇇}��xz3`��uӃm�#*�v`���<���7d���Q^,"���Q�n��hs�8�Ī�"Ϫ0���Y@��0p���SG"O��{do[=Q�����b���ŝ?F���u��<I0E`f�
)]��K�/�?T���˟�D�4u:����$ljݐJ�~;azrb�3�vx�r�?i`�u�jd0��K�̬{������A) Z�t�`��Ե5�ϨO��Rb�
�HEZ6��-ߜ�{���E.Մ�d����	�_�-q�h�5YF�z�n�S��1;S)i�9+�G�U쀉��	�$��DBR��1�
d�5ə#xX�)&��F1��"�$JM �����?a4��B�4J��}����<Y�
=��cRk�<�wf�6x��,�vн`,���n̸yb@�׉�o��� �Rk?�@�>OHh�'���S�? �)"�d��3CoK�f�d�I��'񈍑�Ř2B�Ҡ���2�a5�6�� JZ!s����'�`��3��h����	0�<��ФI�z(vu���['���\¢ʒ]�,��z�+X�0�>�@�'���vg�;V	�e���9D��R��Jnʰb0fU�%��A�IW,dJ���=ф�<�`LS�[��Ijâ�3X��8�5D��H�)�)w0� �Dʂ;=>�9��'�K��W}B�P;��9C��CO�<9e��1�d���:f����@��H�<)6�,lhP^ؔS��/`c�!��b���+sC�UY��XKA$;#FA��p9��%�B9�Ó@�'@N��ȓ@�|m;uH��|���#7��2������R�`q��j�x��	��,2Uy�#%�
ap `�!�YÊ{"���c�� uX` �ޟH!wI�;IQ��P�ᖩR�D��)D��C���:�>i3w�,�us�q�ܼ�G�&o��7��9a� [��5:��S�S9i�ȵ��_�-��A#������DK�o�T���C#�ybOK�����G�� ��{�+[��|;���~�ʓA``�|�'���6bʠS^*!B�χ
�yX�{�gC�(�"T�Ht�O�p8r ̞v0�a��a�e��NǢd��١ǀ��t��d�O�iP(ׇ0���ٕ�"���O��09��O�lj��V�mf��T�i'lz��F�4H���F�����y�'���:#��*�@��-�VSB�-p:z��� ]��R�T3#���:��<%?5��l�6Z&q`��¸	�t����=\O%����(���q�'" 1�$�6wW�ٛ����{Z�y�B��D�IC7��<�r$9�gy�_��8�T��33�Jt�'�����''2��@�Mt���D�DJþ,� 1���+~,p�1d�\;�6�� Γp����"7lOtac'���t��U��n��'f�	s�׷u���[�߅z��d���'{�^,R2&�3`v����S�T�	`$
e�T�� � X!�Đ�B>}1j�67�ZŢ�nC�"�F��&-&L�æF*Z��a�t�!V�8�O�i�O_����j�#-R$)��Ϥc���3�2��D*I�pX���EE��IبD���4+���9F_0vV�B��!X�ԲS�_�h�qFBC�^�=�3�/��4��7�����%�܇y��LI�@!$ވC�	�Ѵݠ�I�)8�$��T�+�z���y�\��ӫ���)�'m�.%���a� �r�A��6��dJ�'g���	�
����ï�&�tC-O,�{3�μp�h˓0�~�C�k��Nd	����'ꖡ��ɭL`��	%킑j��V�?�H�&�	d�ʉ��NX3����SO��sꛭ �*�r�A'(���*Q�x򂃋LU�ţE��9kZU��X$��O�ԍ$���0����,[����	�'s�|�fo�"}��=R�B�c��TgK�i�1�'H\�� ,�.�¸O�'k���(͖[7�W�.E�.�3B�,�<�sc��rr�-F���o�8O��A��ߟ(O���@d��<�����8���HB�p_69�R�ZAA��"qh�c|����	h5y�� Kd���K\�LOڤ�S�@���(
QE:�C֛��Q�����z�D�@T �b���H�D�!�4��ɧ}� h�Ֆj�>�ڢ�S�?VP0��dm��ɔ�o�RH�gA3D�t6�C�	`�/�FL�wC�(-y���>���WV�d!�k�.
dqO�n
�)ڬQ�n�;�j��c ��S����n�v!����A����O9jN��*B.��תE	���q�jҶ(D�D�M�Ffh��I�w�����6�p<��M�9$��!��.?9r�Ƞf�Dh���Nv�D����R~B��>��x��4\��dc:���H�e	�8NO�œ�ċr�O�ӆ#�mZ#3���C�T]©"C�1	LxB䉕	�r�ڂ�	���8g��#L�JP��{b��&d'��vј�a0+��l���@19���ȓ�J4�6�ޟB�����N����'�F�����yWl�b6����@9����'q�����<To*��UďE@jP	�'��Z�՚$;�p��dC�9V��y�y��)�J�%��Dߠca�haJ�	�C�	JZ�(Q����L���Uƅ|#<�ϓ��]��F�$7�T �h\Z����S�? B�Pvnڽe��˔ �k���@b	$4����=>�2D�u�U�iz!F!$LO���r�� ����'�QS��� D�����Q\n=S£B.^����T$4D��K�Á=g$&����D��DO5D�LPT��u�Yp5j�'Y\(�b�>D�D▩^ w���6��0�p�B9D���u� j�ʇ�͇o��Y"*=D�p�L�M���wI	48���S&8�O�	���~��Ɇσ�f�@1'£X ��'�EhS9e�j� �#3>�iN>�#�~¬@�@��9�D�|��J�4dA‒=�d0:W��/�$��	a��u���>S� ���9�$=*����!�"�LKpt�s�c���� �<D���5f�=��c2�"ԣ�+K��O��`C����O�@أ���lx)@"ȧ`ͤU��O�����ŒJɖY� ��yq��!�@>�4��m�!�SvNi�A�H�n��0�t_���êqA�'�e E��F��'Ѥ~�.���J��E�6��HMw�H5:e�P�&��QQ��C�,��LY��4}��i��|���K��^'��\2��Q2�V�\�R,�'�3J�����cPꙠ�OŒ\|:5���4+ĳL�T|h���8���%
���Q�P� HB�@���Od�e'#l�P	��	�'�^�c��L�s��#��K���,ľn��Q?���X�x*֌!@��xH��Bg/"������E�
ܱD:8qb�>1b�����(vv���$�';�L� �+ĸ1��,�e��.5F"a��8OF�#Ӊ
]<��BC��'<�R�P��y�ԟ��j&��||�Q��>$�����,d�i���F�7l�D��"1��
�n�R"���A�$�N�=Zq9�/�)zB��F�ŀ�@ӧ��Dx`�Z�J�I���Mh8@�∥�\r�>`4�tj�1O8�1��§p�(�k���l\):��m𕌂���ɵe���W3	~Vp"��חа<%E]�� �p�Ax�y�� �<!����`�A�$xɦ�J!�o´I��u�
;v��z�ɇJ԰BI
�VoB]���>�OFM�b�_�2�m���8IP�-x���;?�Xh�-��~B-�gr����i�m��A�9HQɧ��ʟ2��y��E66\���AF���O�!�Y�_^�ih�O��H���F6%y��V���JU�"TDy`�'��xu�Ii�S�O��	�X�;�1�t,�%5G&X0�O����/�a�.�O�>��s⒂'����OϘi�l��)1D��y����)�y$JT�V�G�.��U�R�˓
g:��`��~8��C�E[
B>��ȓF=� ņ�F�>�[e*L�Z��ȓ~xA,D�!%D��!�6�T��ȓH������N����T� �T��чȓSY���a0W���P"��%��+X8��l�S~d#B�нB+�!�ȓPvN��O�&��ђ��	?-FH��	���+4��->�d�:p��9Xh�ȓA���ȉ��cP,F�_�,���x�#ef�^��'Ɯ.r�0��*}d��;?}�գ�@�f��h��I��+��S}�J�;�H�`�(�ȓh�Di��F��=�a�
|I�ЅȓqW� ���	���UxD�B&(��ȓ:��p�W'Yc������%���A�U(��M�1�`Q!��& B剪;n�$!���2=Jؙ�,��l>D�؃����{���"��Dq-�1;�?D�X�d��Z��d{d"!z=i�H)D�$"��ǚ<�X����U�52����;D�������4xG�9�J�@�ȗs�<���#oߌ��*�ilpyPcBD�<cn�)c�����[)o�>�3�+�H�<�5La�ͫ�Q!
jl�I K�<�c��26qpb+W����Б�FG�<!�g֜N��f�ܙd�	P4	OA�<)����\�Ru!O�1�8�+P�@G�<�o�t|3'�Z}Z�I�u�F�<�%s���ʑ�(Wx$�2��z�<Qï�
�����JH&�����
r�<� �p��2��p�f�:K��M�"O,�1@��P��s��K��ҡ��"Ol��N�o��t�s�!|��b"O��R�AX)f�ؕq!
%��"O
yK�Z*L!F%27;_�2�"O�m�2́)h�hbi�	�j��A"O\�����,�@�]1Ko(�(�"Od��.�Y�֌ �eD�uAd���"O����+��Pw$�&OW�0)`"O�-��G?%y�L�`c�:A4��"O��%O�}=@�C�!0�a(�"OX�S$H�25�`��"�)(ȡ�"O����%� ��U���k��"O���6�aO�h#�[�M&��!"O�T���_-)DxD�Ԭ�!%n�*�"O�ju�W�mKE� #څ����yR��.0oyR%W,'�:��ꃤ�yb >(/�JF,/Xnij6O���y���}6� ����w��&���y�%�)� l�b��)�ċ��ɢ�y�1]��C.A�O�t�%��8�yr�ʫI����k���Q�@[�yB" jDޱ��tݲ�U� ?�y"'Д8Q�2F��n��DY�%��y��E�&4�aJG ^�)"�H�^8�yR�ٿS�&5!c�%�8��2�y"ɖ�~\��@i��x�+�)�y���5�V���۝| @���O�yBɏ+&�ԋ2O��v�,l�K�yR�ԑ޴�x���r0佚�d)�y2掼nR"����]x��2�A�7�yb)�L� l��̋9�D���C�yRgɀ=��<1	"Q���yb�/n�h��%%�l `��y�π�y�r�7'D�y,�ා�2�y���4鰁%Jެsxʝ $�y��E��,B�B�4Y���:LI�y2�Sbd(aR3M/]��i2�o��y���	Y�2�3�à �fpI��9�y���=w-Ra�i�Bm�!-�"�yJ��F[p���ԅc��U�`g��y".��)M2� �ҟc¹�0-P��y�[4����C�g����铏�y�k\�;�|�@�
�
���ؤH� �y���*��10��U�t��8˳e�y�D��:Qbad���z?
!C����ybK�$h���VM֏h���X���y��	K�@9�i�4l���#t!��yo �CFT�2�$E"�����y��(tnpM�ѷ"���R���
�y�,G��ٛ@Z%V���J���yҪ�� �\�V�Y�<99��Q��y-��D:��CN�9�0���yH�l��LN��$=Y$C�2�yr�W�;UѰ��t�H��s�@��=�N��;|�W���N�n4D3�͖��X��	��c��!9>���L�2�6��=iDHtZ@؍���B����M�1x�ȃ�	]!���9wK6�H#I�x:�
t��XyP�K�����	��"|�'2��)�$ׂ5NL� TY ̌0�'�0ژu��� ���$�0}U�� %�����@x8�TY�kU<�:���	O3���&�6LO�L�$'����Y��'�)RЬ ���D�0j0�P��'�4%e�b��<��g����y¤�
b�ꅳ���p�π �I���'+�z�Ç���:��"O"��*��S� %h&��6K�(�0��O�\\+M�X26!?�g~��˰��M��ʠs��;�fʉ�y"j�!*18�f���,}��J:L��ePrᓁ7mα��IN�p�R��}��2� �%|x���D�	<KT�c�B���~2���q�0�S��Ҏd�H=`��С�ya�0W����C��P&��A������'Nְ�m�	��?�:��:��)
E��E�޸��j/D�X��,��I���
E�C��(3_�X�="�>�#Wa!�A%���yI:D�gM
a�<���9��E��K�s~8m3�]i�<I�ر\�z�*��7`t��Zg@�k�<���_m�N}p�A�&�@�;���I�<a�D��2��u�۸X�:��^�<F��<2��)������P�Z��B��z��)1 �Ц���x!��
%�B�	�w�h0���M�#�����%�;`�~���*��+�)+�Odq+�DXTB%��C�?b��Yc���s3H��=�O|���Ⱦ`��MC�o�O��y��"Fc����Z1ex�4�b"O��Fj���jL����Y
��c�i�L]��bV�Hs��(փC��D�#�ڨJ��)�	�$*��2c�lH�I���z�`[�z�H�˲-��<A�HЉrOؙ��K� #�r�ˤA�1@��xW����	�Q>�n���Zfj�0d�("�.C2��H�=q���rt�P�t4�'��l�"�@����-��زp�'y,���$Ș�a{�3?a D��.�8O��i�,�V�X ��� %��ɠf��-2�AW'��G�Z9�4Em��X��۶tg�|hm�{60��ȓ�~}j$��
����0 pm��h�I�C>@�� �L��}P�L��`}�S���~�1R��������ҧl��H�'��(�4��-9	�R��4���Y�$,�"��="D�aU.�4��Y��0��<A�#Į*w� h�l��?��0���W�@j�T�ժ
�%r#~��oF!<�H}Bre�1Z�%p�L�h�b �3o�'P����'w2��d�!5D��H��-��U��C�MO\�qĜ�~��D�P�h�b�aa�'��}aB+�!B�E5�[0�&�8�'���q�@�b�x���+K+%m�!C�4��-0I>�d��%U7ǔ�)dMc�	��T�+
��$i��_�FD3����{k�{�(�4b:��F��(���B�C�F]���%N+&��b@mH<9rm�o ����0rj@�+w��_�'}�D���`(5�~Z�
W�pw�U)�\$�����X�<)t�ô-��X��C�\�2-�R���D��k�.�⥚>E�4-�0_��i���-7�����%ϐ�!�J��e��苄?��]����7��$��
u")�V'���<	B�F�x@�$B���R�]x��h`O$C���"���6<4�x�H!mY[��X�f���їȁUn!�dQ�t����s�ҍ|.K4 ��y�'��L2��@%8�<Z�ޖwt�A���d��=%p�A�CEV���ʦ���y2� p�)а�fA�6a���U��p�1��"F#.h;��+ܸO�' <8�va��'v��`�U�g ���'�q��<T_H$��3u�8�Rr��9hz���Ĳ :�({�����<� 
��[�.5��#V(і�j��{8����
�^� Xs֪��c�:��3f �|��y�2��	�ň�?�!�Ė
Hf��t-.y漈��\�	Y����#�>���қ���!�E�f8(�����!�;
_*�`C���=�rq�e �>��Е>��J L��>�O��b�'!���S�ٖoIb�;�
O�U���^�G[&l��Q�R�6�J�샵k���(4��'�0?*����k��1�
��D��v8�L:�o��e��:𓟔��L�R 8U{P-��{N�p�*O�����AO���R$�/ �Ǖx"�H�4Z
(F�|��d�ߗq���0lK#$�(pN-�yŔ�L&��B����v������$�DL�g�D��z|DM��KM�:֍îY�!��:F��t��,�Y����P�>�!�
*1I�5C��?.b��m�!��̄s|�UG�3z�f� ��0�!�� zM�r�
�����Ƙe2Lk'"O��S&l4;�б���	*�5��"O`��[�Q��́1CT8s���"O.8 tD�	�vH2�HlbD�"O�t��VEӺ�SF�'dN8�"O.�)�h��M��P�#kM�$]zD��"OA�cC+-9b5J�*�* ���"O|H*�E�<
p"_�]u`)Ic"O��L�r�FE���dPl�U"OP5IbCV"r¬�P�C@pP��"O��R1��5�t�u��v�j�I�"O��b�Z�����S^����R"Ot�k5,;v��rF��o�Ԕb$�'����*��x/��2g�yI����O���{�	��j�WN���ٗ2�
\E}2.�!)��a��i�9,��)�9�Cr��TX!�D2k+Z����Lp�"�T�2H�	<�l`k�7��)��3J0)��Q�Hؤ<���  �2�U��!
%!�PΔ��(S
{E��A��V�ɦ�4#f�!�2��Aj�3?�i&���>cG� ��,Q= ��{��-L\�?�#�E�:�[���l�Z���(6c	+7j��U�!HR� �E��c6��J�`��\�S�O1ƹA��]�w����@@�b����]��U�/���pk�D�i�*klv�>�r�N;Y�|���ڱ �Xy'n�<�%��1o�f��"�=,O����Y`.�e�1S6�يT4O4���f�X�Z�۬ID�'�F�jF6Z���[��K�v 䨀*�h�"5sfm0�P z�1�\ *@�� ��(�%�%/E#�G�H"�:RHk� y�"Q�6d��`�, ����^����?��*J�<t�+䨘�n�\x���<�{��|��'�3A���i�_ (�gj2N1h�s `�0�4�{��B�0�=�4�ƺ.jC����)�'	H��5�L�rb���闩KB��'d�y���D?K�F%̓ ��J�fX:�T�>����(L�����ٯC&ȕ��Ƣ<�S�Ra��*/,OBi�S�_��EK�G�}:Z��!0O�����5�n��g� �il��Hw�F�38��P^���Y����[�|���F#"ܽC�&НP�����	Ň��l2�ǟ0X�����h ���}8��m�����BI�G�i>�X�ŤM���q��C�4V�`*��!�5ZZT℩ܟ{>�DT�Ѣb
%(G�!�F�F8<�Z����S���Ij�l�����S[B��"Pa@t����-�2�
2����]���S�O	�0 E�b���"AE�yf��1�'v�ECv��J[�A���r]���N>�šs_���dB7`�������{�蚃A~!�$�(2�D�R���^�,��uA1k�!�D'7=pTKr�����A
�W�!�$�{�tZ� %aɂ@B�V�!�	�"%�wOZ/�0�o��!��6cSB�QA�_6f��Q4��6�!�dE8H{t9��T>a����햤�!��7O�6p���	qgDh�K9:�!����(��&WR�����Y:G�!��a=,�� ص6w��#�#�yM!�DL%�����C�xt��2$��'#!�ė<g�l7� �G3��XP㗘o)!����(�P�H��8���b(�0d!��O0(FA����2:���S�A��!��P�8�B@'�u̔��Ꮛ;�!��?y�Ȭ�$kĉ ���RV �e�!���<{F@�buC�� ���`!'�!�d�L2ޑ;��[�4��� ��S�hq!�51j�P7劔H(����@�
l!�d��P}�E��
�qR��C�N��!�D��2�2��4�Q�	$I��nH3/�!�ϖ}���h���#4�������N�!������bo^S,0Tr[\�!�DE �p��J.>A1w��!�!�$��K,�$qw�y�i���+i�!��Fg>�Y�ׇ.L��LS!�!�� ��dsK�9��F�%h�$�"�"O�󀝶K�L����,���C"Oj���)F�;�Ta�O��v�P1"O�1B�g![��U9Pm�{��л�"O�q�6`"*�X<J��L�h�:<�"O4���.���˧צ\�)�"O��i��Ƌa�@0��HI��.���"O �p��"w�.@�Ԫ$��"O@�1�kL�Je�A��A$�"mc0"OV�b��w\mi�#��
'"�9$D��lA<<����a)Z$Q"p�;Pb�0{��O�SU����2(U�Ah2����4L$ Y՚>�Ƀ�!i�L�|M~�iLeRr��ӏ�-M�.��� RB��_�[��YH��A$�0|b���T |����&Ul�j��|?	�C��6�:p�6}��� �5	Z�iA)��,���J��+<�S��U�@���>E�t�J��S+��Q�d҄ș%1F��j�$>� <�M����.6Mp5�ᓬL-dD����=�����#!9����b$M�-�JK�8�C�~z��)ϵ�n� �J����Q��%8�X���R�V�q��]�>+bDP�S?�F��ɜ[����R*
 IZt�	�I@��?��

�,����e@��)�GҜ-{�L�\%x�	���X�Xp4�2�}�E��p���"�f�[6�K4xB"l���Ǩx�A�>e��@�7�V?1V���L�$��@�"�lT�MNR���P�@��� ԭb�D����t@�~�	&�I�|��)FT|���umn)�1_�4���/txY�۴R�a@�J?֝ݟT�l�a��}��JV/s��!@�J~Ӕ�)!��`j� e��]I�O��Sm��T��	��լx@>�O<AJ�+Y��xn�:�PG��)h�*Tk@�@6>�"@�� l0�	� ���i��Ȏ���d��B��4,�j�N�gBҊ��	�nԛ<�?O��AH�<t��wl_�)o�Z\�|��h~�a��F�"D�E'��t�>ɍ����D�<+�(z��%O���k�����0>��fķGpe9��A�0�,�`i0.kDx�a��+� ��C��S���`E��j=:E%2�ɚA�LU��S�w��eZc��;���bP
F(�O��'� ��Hv˧V�$��o&b$V�V #����F��8;Jr�'�l:���l�����>﨟輨�.۾4�J��b��6i>B7�'��CÍ�*,�ʤa�Ɠ�t"a���ֵ
��t٣�M�h��y�Ҋ����h��}�
�Jf�qP��ˁB�xS6͇�D1xu��?N~Lb��؊lZ����)�d���ujJ(�A2)lZ}�ۍo2Ɇ�����r�˖���P�AS�6u��Lj�
�dV�Wy����
?�D��ȓ^��)c����LW�T8+��C�fD��`q�I��O$�P���	;>/&���OD�@�-�8��d�7�2%��]z����&`M��PîB�Tơ���e+��H �0�kG�!��Ćȓ]��'�7l��Ҷ��gt���>�\�':SeL�F��?^z��ȓUa����Ί�p�H�fE
��@`�ȓ�H�SSi�zP� �P::���C�^�CtH�M�����A]2.8.Y�ȓ���'�ӭz'&X�cҵQ�J9�ȓ \�}��Gεw�ACA�\�p�ȓu#jm!#�1v��DCƇFK(�ȓ	���{Q�Z�3�`4�p��o�,��ȓ]���Al %ˁ#J�%.���p���cI):�n���"R3�d�ȓ���0�ˋ�t�Υ�t%��-��b��]8q��XDpS$�]	�͆�L� '��p�������Xc"��ȓc��,�"�ޞ+�<I1$��,ex��ȓ�e�a�FH}����fV�]jņȓ"�H'�J�Jf���uL�:F����X���)��#(�!�"GW< �&̈́ȓ3��\*�k.���� xp��S�? (�#`:6���ِHƌ.�ͪ"O��vE��A��QBBH@0��i�b"O`�[��PP��eSe�*���d"ON{���a~,H�W�+jd�i�"O�av�)=��V��-�BIx�"Ov5����a��*��w�����"O��a� �`=(���	�.[3�y���r����c	H4�l����y¢�'`��
�ʝt˨1ᓉ��y��@�������aI�U�r�T>�yd��L��H��� B��8Â�̖�y�'[��D��ʒIU�8C��yr�סp^��d�A�@�$��a����y�j��7BPh1��7h�ݛ!l_��yR�҇!�8�0��_�,a�9@鏁�y"^!8�tX�G)���,(�Pn�0�y���IHbY�T�D&z�vؐu�M��yb91�\[�b��ZD�o
�y��>`
Ⱥ����"�L�Ys�ʊ�y��</�Չ�E	.n<pg���y�&r�� A'ȸ_�$�	U�H��y�3s�1��	͔,Y�<����3�y�tb��!�������/]��y2� ��l��	��n�n�94� �yr�}�B�1���f\Ą�I��yrǤdL���K�O8�))`����y��P�鰤��HB'L�h	ڒ.@��y�g��g9X�pK�:���/W�y"*Z" s@X;@�RW-E"�y�OL�p��{��Iw���y��	G�&N�z��|���_+�y2B�h�r�3��=��2&���y�'M�>�2I`�O�3;��P�Iȭ�y�޹Jf
�x�䈧%@���Vg�,�yrj���s�J}�)�����y҄��7��1�!�;�@� Dᘰ�y2�M�D���0M�70�E@���yR���Rd(J�+إ�u.�$�y��K��<� P(T�o+�Up5Ȃ��y�"�k�F9Jq�C�c?j$)ƦO��y��!�viI�⁻*�2�զ���yB���`�|xҠ+hH	E%���yb��{>��H�ۺo3�m��*�yB�o9Ry�cM�9j�H�C!���yB�@_u�U���aݮ��B��y�6x��`�LU�x\	abD�*�yRhӆf2���eӺ6g����dҥ�y�X;����BC#,�(!���\.�y�8m�������e�֬܈�y��:��A���t4����y��O"�R
� �-`�N5�A����y"M�*R�8�x ��
D�Q�1)E!�y�Cբrj��6�Rx��(��y�`%2]�����(�$�I�K�'�y�mN��������Z�qa'J,�yb�6�|s�DX�0��s�̏�y��ܮKN�	@�1�6U:�bP�y�J�^��'�8?�jXB���yҏXK6��(�hC=n�x�Æ�7�y�L%M+�;�/�Z� H �́��yr�It�.� �ũW2���*й�y��\����MKU :�������y��څEl<C&�E#}J��'̔��y�	�R��%��'S8xܔy��	��y
� $b���X��k��[9�ִ1�"O>�iP\A�5k�C-\n�a��"O�R�e��h��䡕���t\��1"O��;P�؎zMĝ�6(K�H �d� "O]�3l��&�zI��ң"O�kS���+|��s���4)��"O��rf'�'LBtɂcfR��U�&"O��(� U�C�Tu�S	��
�"O�qSV�����W��~����"O�����8�P,�6�	��9�"O������%���g���*�I5"O`�4�G���٠�bD�w���5"O�}�5�ٶ[L��y2�)�y�"O��"ca��2l9vaӼ)V)�W"O~���M&R?.����T�z�"OfH)W)N�S��d D������"OU�2%C vm̅����%�^��"OɛN�5H4��3�]�TAn�w"O +r��PJ؅�b�ݭ1�42s"O�q
�扝w;K嫐��Z�"O�`�V�Ӏ7�d�4���*�dL"O�u!��Xh��aM�G��`"Od�B�">
Za�j��b;V���"O�E���  Dz�oL+N4�u�"O*����.'�:���Ͼ3���""Op=��� �9"�m�JR�$C"O���`��b[�,�
K'h�Q6"O:h�U
��W��$�P�̴ 9\�@"O�<����¥�T��RP��S�"O�U�E�Z/T�M�Pb@�5����"O8�"�n��`bZ�q�BX�`9��"O4=�0▐V)2$c���p�8�s"O�d:�BƸw^
���]6[Vvݐc"O�\� ��S ,��E�+p���"O�[�c߄)}Ȩ��c��X0�"O\U��[��	�bB[�8�=X"OP���bOزE�G}ܝӣ"O�����������%΀�}oVB�"Oh<�Eo�$�@��*�3r_(\�5"O$��r C>����@	 
�x�P"O�4`�Jͤd�ء���6�@G"O��``��)A��B7��k5�(�"O��x�ǅ��2ex�L��w����"O^���Z�T�ܤaQ�V�uV��c�"OD��bH�}�r�P1��j=T��P"O�A�ի�1�riQgFC�uG:�"�"O�Ir�lF 1��d�
C+!��i�"O���+ X1������b"O��l����ɶ)U)%�
i�5"OR!g��0:H@�
Ȭo��D�Q"Obe��섳�����]�wκe:u"OT���#�*Yv�����N��x�"Od��gݨ�l}HA��<q��Cq"O�Dz�E!fY���fd��k��y�$"O`�җD��<�\0��ɽd���b�"OHɉ'f
3���t�̡in�� �"O|����׽9��[�ɓ.[�Xp%"O6��F#V<I�j\ң'�/@Wt���"O
�+CK�F%�PF�]�8YS"O���� ��q�"yq(7~Q+�"O����P���F/$�yV"OZ�r��J)&����&��7��D+E"O������|e�4y��pwAk�"O�#�_T�q���˯FEu�Q"O� ��k���qh)����04QXd"Ot5
W	M�(��q�[,#��H1"O�9��є&�vh�&�pe�t�"OTxf�:��	�� 9J��Q"Ox�)A͏�y�赩����"7��W"O� A��Y��
ҋ_	��R�"OV9@,B~���sT�N.��	�"O�ų���:F�1�D!��!��"O �A��̈A
������Q"O�|8��J�i�p�!��O=	�N!Z�"O�RpEPvA`���(*l�܉�"O�=���k�P��凗)>�-�"OrqRf��+: 4����08�iD"O��,M�i��+U
&��6C���y���$j��	��Ӆ*D\1'��y��ռ
EP�R�'l���5��(�y�7f�H�2큼m60��,��yb�^8VVb�b)�0d |�	�b
��y���̚%��Ƹ���O� �y�(�eL�	���Ѩ�3�Q�yB�M�L	�)RL�< h�"��y"�x\��0%�!a>e�!!G��y�̎+�n��c��щ��yRP���H��bW�I��ba�-�yb��ZZ�C0+*FKJ �E�:�yb��6hW��C�DJG1���c#��yr,�:�h�c�B-P$!���8�yb	�*2D�7 ��At �����y���";gT�X#�_�c2��� g�2�y")F:Uľ(P!(�_��R���yҩN�7x<�bo��Q{��( g��yR�N��x�A X+�d�I�,S�y�m�Pز�k��`���X��y�Ό�1&�`j�g��+	��RW�M$�yrD��zNR��!�FaA��yҮ����ӥ��򩂀O�.�y"�C�>���
�$�����,�ybo� ������R���Rb埂�yR�?�Թ2�E�8S���f
G��y�HG    ��   �  i  �    �*  �6  UB  �H  �Q  X  J^  �d  �j  q  Zw  �}  ��  _�  א  1�  s�  ��  ��  <�  �  ��  ?�  ��  ��  �  ��  �  L�  ��  ��  ��   ^   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n%�^L���ܮ*����EK�0�RP�"�%?���i��O�9O����-t<���C$m����EL�d�O�$r�r����$��$�O_�h���4j���RɀF�b0�yB�'��V�O������^�q$V]*B=h_�1A�l�f�s#��4�Ӟ�M�;U�"M����-V0���L* ��P��?љ'-�)��8'y ilZ�<��!�=�e�APht��d��<��'�$A��hO�)�O��Ѣ�АsaZ���v-���0O˓��ji�&�2Ę'������fڶ����"${<�����e}��'��=O,�)9�<���Єum�u�Q��Ar�$�'���,p��,���#��(5�'�F��7gş ��=��L؍cT���]�<�'U��9O�Til�*�~����Y;��q�:O@�l�!x�x�=_��4�F|	�"R.r�����X��-A7O���O��D�>Y~6�(?��O�B�	��|<� ���f���``�[�3}\qI>i(O���O����O��D�O��G� ���[r艎K�~��pį<�0�iG��;�[����S�ߟ�qGJX����Aȓ�c�4�jQ��DLΦ0�4g=�����O��t���<siZ�CZM�d��=8&И�iB����ZX���1BL?�I���R�a1��icr�k�b�=a�d����؟�����@�	՟�SOy"}��	g%�O�a��d5���A��9v>]Y�$�O�yoW�{��	�M�R�i�47��J>�!OE�v���� _
�)C'`�6物9U���̋#���B�<�+H�����VQ8l8!/�6g��1A!�U����Ɵ���֟��Iџ��	s��%�j]#��Z3X��P�Lު6	��y*Oz�����4m>��	��M�M>Y6iAD>*�k�Tx�.�d��'J�6���i��(} �l��<��f�A9��K�5�*�A�^�-����臬rO��D������O���O���6�:����$�A��		�~���OF˓r���PA2���ЖO��� ��P�XsF܀�oD3o޾���O���'~�6�Ҧ� L<�'�Z!'�*?���y��[�1�H�`C�?r��Z%Fݓ�M�R���S�1��D,��ol�J�G}&�Y��1>mV���O��$�O����<�&�i����ƀI04 ��
�U�~(�R�.�&m�'D7m%����$�ަիF(��M~mGte����	��M��i�u���i���O�`b���R�o/?C��4T"���ڻ��-	��|�@�'���'bb�'��'Q哚o�� `�`RV!�9����4���4|9�H:��?�����<����y�R�^d~Y
�Oڔ%�F�:�ʐ8�(7����N<ͧ�r�'%�f b�4�yB.Dh�u������gj�Γ{�����On��K>�,O��d�O��qSa�y��P�����򄬩���O���O��D�<1T�i@�B �'X�'��t1�QN�|1�Ϸu���s��$�^}2�q� �n����]B�)R9�Q�����J�Γ�?IC�
o��Sp�4���
�a��R�F��$m�"x�)֙c3�����N�d�O4��O���2����*�V	XTJ��P�L�*I�vL��?�7�iو���Y�d8�4���y-�K�)�5KJ3Wߪq�ACP/�y��q��LmZ#�M���M��'s����-��'j��<�u�ʁ0M�p�M�-��L>�+O8�$�O��d�O\���O�0	�EȚ'�S�i�I%�h����<���iw~9#A�'T��'���y�C׭���'����yFJ�.n`��?Y�4S8ɧB���br�D<	�c��sօXKE�NP C1AК��A�Q�xQQ��Fk��O|˓˜L��`��U���"fCY�}.��j���?Q��?���|�,O`ql�Y�z=�I4)�x]�w@eY�����4lK�;O|�og�M��	��do�4�Mۢ�s(=f��0��5��y�|L��4�y�B��V�������?mz�8O����he�=� ���^��Ea�M ��8Ѡ:O��d�O����OL�d�O��?��-[+l&�+g�
�\�H���-�Jy��'3&7M A����M�����^�n��$Q���!dW�;�h�~y�'��o$�M���*cI��4�yZw���G��e�H�B�@9l2Y�g!�!Y�x���'�&�|�.O^���O����O���!˦j�n-	�=I�]�Aj�O��d�<�ջi�dh���'��'��>U�|��� Q�i���I���n7��S�ꇱY��P[WCB�u�2X��+�z�~P��H�
em�&ȵ<ͧJ�\��y�ɢk��y��� �Iy�N*�t�	��h��ݟ��)�Qy��Ӭ0��&~�HI�cnG�

�I8CË�a������DF|}�ak�l!@��P�>�J�C����3�A�֦9�ش4k�iߴ�y��'�,�f�Us�,OT	��f � ������5��?Oʓ�?I���?	���?����) ���}�7��շ���m�Y��ij�&�'�2�'��y��l��&4XdрS�8�˄�X'3�mn+�MӴ�x�O���O̬*�it�Č�6�2HXW�T�.����D>>󤃄85ڴy�o�ؒO�ʓ�?	��S���r�.�'E@wc�����?9��?q.OvhnڛFv@�I� �I�	C�5�5��&�%��h��w��I�?�T^���ݴ}���"�>��������'�<�I�"���O(�V(��h��Qͽ<Y�'7���H��?)%,K+Q�$ec�6p`��e�E��?	���?y��?1��i�O&����0o#ȸ�׋M=&�2u\0�$���q���Zyr�d����,=l+A�r�P�1�m�,T=b��ɦ�1ߴ#'����b��=On��Ή�T���O��u؆���]r4�9E��;I\�qs�|rR���	��X��Ο������wg�3��3�T;`�N
$dUyr)i�J��p��O����O��?�R��	�P�Ԑ��%�/?�@�V%���T����4cՉ����O���Z�):>�P���)z0@�&O�(:��Z��E�=xbO�y�Sy��W�.����6f�_�X1�,\�&F��'F��'��O����Mˠ���?��!����Ʃݩ"�����?Ɂ�i��O:��'�¾i�26�$(�ҭI4V�5�l�#�ݣg-��Qw�x�4�	ٟ{d�JZ�dh�~yB�O��
�0�,`��K�\6l`A3E�%�y2�'�2�'L��'���iJ�Y�m Sa��B�N��V@s&����O��䦩�t��Ty�"d��O"];Q�צ�c*R�+�|�XbRu�I<�M�ǳi�����s|��<O���ҵ^��4�6I	�|`�h"*��q"����?�&��<����?y���?Af�^B��A�DW$N:vD�����?�����dXЦuh��쟼�I�`��?���	�=�u"� �I
�!�a"'?��X���ٴ`q�F�%�4��I�;U�A��c��s�n(0��88��G%=
�HCǪ�<��''���+��L:T�2@N��F�F���u��T��?���?��Ş��DĦe0�R�Jo�lV�.+���V�I�,��'��6m7��-��$��is�"��Nh!��)�5h��r�թ�MK�iV�x�e�i��D�O�|D������<1��D�e��3��O�s�꼓4��<y.O����O��d�O��D�O@˧.�TS�*!_���%l�1tHdx��i:p )��'���'W��yr�o���]��CW�S�+F���#{N|m��M�t�x�Ou���O��}�Ѽid�Ĉ=�1�nC"bTڸ`W�~,�d3�(��t%�O
ʓ�?I�WE2�����t���"W�QފI@��?����?),O��oZ$kBܗ'��!��u��u$�$y�u�6J^��O�'��i{�O�apR�˦UHe��@Ct�S=O�$Q�bT99�'�:�@˓����O��Z��%�A�>��L���1u�� '�������㟀�Iş�G�T�'�<��n#
m�ݛ���,!�I��'��6�DS��˓` ���4�P����ݰo� �d�Tk@���8O�o��Ms4�i��ƹi6��O@�`Ҍ���Ŗ2	�m�$N�)�Ht�"�)@���O@��?���?����?a���X�a���^.��	�OibT�)O��m��i�u��͟���A�s�x�1ߧN݈HTO�E0�Ǘ����̦AIݴ	������O;��#[L����+A6(-��٣�Z|F���Y:�� *j�e�'p��&���'`yP��Z�X����@�U��`S��'V�'������W�`r�4a��,Q��s@0�j�.�'2�b,�j������'��'��k����~��	mZR��0���9!�v4��厏]�b�sG)�Φ�͓�?�+�!���釅���䟸��N�R
,J���H�}�7���e'��O����O�i\��'��hy���zv$ȕ�^�.���"�O��d�OB�n��6@��'�6�4�Ď0*^V��u&�Ȳ��$��'��شZ�6�O1Vp*�iO��O�3䥁=�v�hՍP�nn�%�(J,ܣ�'��'�	�t����	<�֝���&m��T��b��p�I����'d\6m�&�E�'���'1�S�?.0ɘ��>n�f �� A�mX�o��I��M�ѷi0�O�	���y�@''�:Ǉ�\��A�5�3٢@i�- t����C��O�UhL>�0j��i^��i��_(Ҧ@������?9��?y��?�|�+O�$nZ)}T�):�/��lahZ�/��9Úcyboe�h�H�Or�nZp��@�ah��c��P�[�����4E6�&O&�v;O��Ē*s�8�Oq�)� ����%�4ֈ%�0��?��\��;OJ˓�?q���?����?)���?iMI�|�:�Vj6��2խ��Fl�E/9a���.O�ܦc>�`�4�?a1.^'Mv�C�@��i28`�"[6⛦c�<$���?M�S`�d-l�<�d�<o���B�.̽	}�����<�V
�/J����H
�����Ov���/��E2�K��Vyps!�.$���D�O��$�O��H��&HҨl���'����o�Ayw�BiE( Շ�^[�O���'S7�Ŧ�H<i���0��e�H�%JЋ6K��<���W���0pa'u��M;(OR�ӄ�?�7��O�I�3��/�Ҹ��b� #�Ƅ"�N�O����O����O��}
��w^p���P f����E�5o`��!ۛ���	W���2�M[��w��0Ư�>�9#ժP%Xp �'\�7M��:�4v�I��4��$�!������jp���/��Րg��
+��"��/�$�<���?���?��?�b�\�lp�pB��,9��Ӗ��$Iæ1��BIџ�I�L�SG��'����?x�F�*� ��0yk���>�%�i+�7��f�i>����?ɪ�A^<����5���Ť{�R���LayR�ߪ�����2��'���$F����D��Q���Ba퇗1z��	ٟ�����i>=�'�6-�#�"�$ݓm�
E1���̚����e�?AfX���	���cڴD�&�#&�˥5i�h���X�v�1�۠�M�'6t4+U�%d�8�'L܆K%�O�4ט� F��tO�VPI���r�f�	ϟ��IɟD�I�����s����AQmR s��� ��C��)���?Q�Z4�v��e3剰�M�M>�".L�l���+5�qk� "M��)��'b�6����ӭM��oZD~REܾ
������V�s
��[>�I�����!P�|�^��	⟰�	�x�U�H�fji�0cK�u�"x;!�Zڟ��Izy¨a�ҡ�b��O����O�˧4�Ҽ�2�-<.��#�X� `��'l����{Ӵ%����?��HI"F��ru`�$	a�Y룪ѭq���U�=W�e�'�������&�|R�
�J^����%*�Բf�@+M�'���'����_��۴m�5�R� ��aL6��q��?1��k���d�F}��hӬ�1��7�	��e	�&�<X�L���޴D���ش�yb�'뺽*����?	�EU�4kv��4~��X���YV��``|�@�'��'���'B�'哈U��KRcX�x���	2ǈ� A��Yش}����?����䧽?Ѵ��yg�K�q�n�C'�G�:G0=�Q��,;�6mKͦ�I<ͧ����)&A�۴�y��G;=vȘÅD�71Ѽ4Y���-�y�̛\j<P��� �'k�Iȟ�	�W�)�b*��y�� �Z"�%��՟�IןĔ'R6���zV����O �d��XA�p@�Zj�"ǀj�lوr�<����Ms��x!�a�Z���m � �!P�@� �y��'�H
۩Mi��*�<����F�	ğ4)���B� �H�aĩx��D�&ߟT�Iğx�	���E���'��PRW�Ʋ�А0� ;2�	+��'�<6�\�_b˓hh�v�4��x�h�g�������"����O�7�E˦I�ߴ�^M��4�y��'��i����?�
d�9BZ4Q�#H�|@H����΄G=�'B�	ϟP��ßP�	۟���1vQ�i�aD	+t#�`5��-��ԗ'��7�4f���O��d5���O|�����a��".�q �$ �G�\}�n�b�l����|*����EL�S��l��+��P�
� ݂,{��wO������0
�����6���O�ʓ^���a�� 
w�E �.��7޵)��?!��?���|�+O\o�U����ɾ�^�ᑍu��e�7e֫D����	�M{��>�g�i7m�ɦ�@��]y��re�`w"� G+Է�,�l�<y��:�z���h����/O������=y��A?W'^(8�c��&���Jt>O���O���O����O>�?��G �'`��	Ck����A�bJ�Οx��ß��4~���)OL�ml��� ��V&�Aī��c��P(I>Q�4ś�OXYt�ih���O �0T�˥,�3r�ؑqK<�0U�ņi�L���$��O���?����?���xt<���x'`�Dʳh�4	���?).O�mZ7Lfl���<��B��8��p5��7f�@٥�����{}��~���l�5���|"��H����s��,	�8�*҄ũ}cE��	!�l�bjR������F���N���O��4�؏}EΩ*L��9����e��O���O���O1��˓,��&�I��r-X����St�s�d��_�%���'҅pӎ��q�O�AoZ<��Y��"��Z��P���W�&�,�A�4_��V�M��'1")V(xab���1^��I�=N��Ӻ%`���3�6�IHy��'r�'7��'�RU>��+s5R�h�%M"Mb����M#��¢�?Y��?�K~Γ[&��w�N��f��]�궧 
=	�@Ӄ�d��1l�����|2�'�ZD䕗�M��'��%A��֚5�,9�j<Q��ؚ'Kl�Z��S?�H>�(O2�d�O���)A�}����G*֕d���'��O"�d�OR�ľ<r�i�t�*��'���'�N�C�"%_~�;d�כZ�*ͫ��D�g}�HzӼ!n%�ēQh�H!�ȅO��0��'�;e���͓�?��_��fa
Ԉ��������iD�D�4@Z�ЀJY�
qx'�֜n����O����O^�d*ڧ�?�Ō;l������N��I��o��?IT�i��I�Y�d��4���y�CG�d���ӧG.H�X5H����yB��Ox6��립��k�ܦy͓�?Y��R�:]��	�M�? ��B�5%�.�@A��P	�y�F�9���<i���?1��?Q���?a�ē(X=���~�:@��X���D�Ħq��$Jhy��'K��e�W��C��]��%�536PT���tyb�'֛��:��O��$�OkҰB��[FH`���V�= ̳Mþq(gU�H�V������*��)-�uГ�IX�P�;��O�=��O\�9m��8$�H�s��ܢ�1D�lx�� $0]Ft�##گ�D����;�	�y��l�	�Lj�����G0W'T�8�j�1��`��K
�nk����e
C 8�di�	���H�'Z�E�RW�٧��3�P�5�U�;1v�A���w�&�ѳ� Ԃ-�@̇-,*H���'�\�a����T�"b�!%]���\�.���c���L��1�Q<�Rxl��Z��r��^��ڱ �!خ�Y�O����O��O����OUʴ��ON9	Bk�2F�m��Eьc5�A�q}��'��'.�*+���I|�CΆ^��̨�CL1|/������iכ��'��'���'����'�� �*9���W��hg@H�m�x�IAy2�OC}���d�
9��HJ��EҲ@́[�&E��Xt��؟H��>�`A�	`�Ip���ǌ�� b���v�l)D�զ��'�T�J�!i�\��?��'sJ�i�%�v��?h���c@N�k�Ҹ#A�r�,���OlI���O��$�O��?��T���:Q���&JМ��DL�~�D6-�&F�nZڟ�	�Ӗ����<I�'��N@*���? :�=����>R
�f(N0xW�'}��'��Oq"�'��F�\33���p��	
E%�=JRE ���	П4�ɸ ��ۯO�ʓ�?I�'�
]p�R>'¤��A�En�3�4�?����?�cBX�~��������۟H��I��	��F64���JR*�dK"o��*%�Ҧ�ē�?�����{�EEX������0Cv�@0�Uo}��Ѓo�[���	��t%?�0��A6�ZE���f�Y-�(Qj���}"�'0�'x2�'*f��%Ҁ=4��j�F��c�]JB]���I���Iuy��˽:>��U�~��ӎљ
Ш���LOK����?�����?���k��K��W?��Hbf��ԃ�㎎ah�u�gR���������~y��Bzx��?Ab&�'e�`�F� 0b��p�S�,���'�	ş`�'�f"�P>]�I�ϸ��s L>,P, � D�'����4�?a���?	���t��W?�	؟\��;>�$`R�jL�C����GI_/t.�9�O���<�@-���	�Ol���?!0F�V�WnR٨1@�CTx@�сs�J���OX�`��Ϧ��'lr�Ox��k$Ǳp�<��"ͭk\-x�#U���Iß`Q5K��I˟t�	Z�cr�C���e*L!i�-\+:�)�4s��Z��i`B�'f�OÖO�)�A��)"�ֺ~�V)�����mڥ)gzh��������h�m��W>���Nj�pił�%{J����ż�M��?�3�ཐ/O��I���# b��``�� =4���#��L�O�������./jQ�J�&I<���+�M�l�H���Gy��~��B�?���Xŀ��aQ�@5w�7��On@����ܟ��'v�C�P~D�!^�C��e� 6F��m�W�D�	����?)��?1��[(Z�$��G��l҄�V)g�4�ۈ�')��h����s"�_6S<�䒧�ϡ�6�������ڟ��?Y��?A���]}򊕘h�>��PbY�>@@%{�Oŧ�ē�?�/O��ŧ4��ʧ�?y�U��p	V�״ k�x���"2��F���O���ւ*� �O� s'��K|��*q,qi�#��I㟀�'` �bc(���O���Ƽ�#Lx�8ę��N�k�=`��x"Y�� #�ӟl'?=�'d�LJ�J�&`भ�7�$ �bL�'#"�U/y�R�'y��'��Z���07�n�S��N;�(x��P�<�`7��O���G�\��b?ɐw�1,�!0�=)8�ȉ'IxӚq3�P���IΟX�I�?��N<�'J݂���_�W't�SCڭN\4����i8H�'P��'R�O��s������+d�̴��h�
_����rΟ�&z0��'�ʼ�2y`0���b� _�ݙ��Fv"
���3W�lx)D������6e5'I�uJ��T�@����vo��2��9K���ŉ���м��g�)�OO/'L�+�䝱?)�l�숎,A��Q2C��Te��[�a���hS�_3<h�皿+� ��.�7������,�5y�#�y0�	�"�0��	ޟD�	ڟ`���ɟ��I�|��dЍ?Sp$���� p��#��\�d�ް��ݟ��%�Q�\�Bp��DV�N�X�f�JQm�����PXt1c��~\��bG@8n����Ǔ<�u�	��M�G�4<�M�0��<V���DbҼby���dZ^��yB�(���n�y_��"�y�b٪@"t2fa�<6��f��y��>9+O6HC�d���M�Iߟ��O�
p�CD�:e�MkƇܥps��▊B�2��'2��_�� �[C�24`�kT�K�$��O�jY��܁t�vi��� �lo�4Î�D�]���Yb
=�6c��;iT�'!NB���)X6ɂš�	@�HGy�a���?���䧡?9b�rV8�y��KL���r����?����9O0��6k@$^АYsV-<(S$`�'�O~]�)�|T��*�?q4�#�<ON�[�Mզ	�I��<�O�X5�'���'��d�Ȇ�d>�٥,�"����H�=�l H��{�^�ԧ��'��O� ����ԭ$ܜ�3�L3E>܃&K[)���:�/�&#��J�O?�H�$R *�q�x��5�	����i"��OZb�"~�	*hu�l�g��}<��,&C�5J��H�����1.}����v�2"<�$�)*G!OV=�+*�����K�<ivG�Q�|DK�G"J�����`�<1�HXc�ԑr2큞8����Y_�<��fW���������kB*��\�<���ڂ4�!�D�iB����D�W�<qfd9qH��R�P��=�F!�L�<��:�P�Gg��S���`��G�<a�G�J� XA@�^�^A����G�<�V$�8iF8u���GCT�`#$�]h�<�GOO?��< �J
�\V +��a�<1��ۀX� @:�.۴e������`�<�6�ҟLt�k#�
e��X`�r�<)DLK0[Q�=�qB�{�RdrQ��j�<�^XS �D-fuz����>u�h�ȓa���z�Ʈ+���	��&\lΡ��u^�d�S�ͧ>6� �Ӌ��~p��0_��*�Eǲe��p��]�5����%��F�3F,^�]¹�ȓ(��cE��,)����1�B':��ȓ'�
)Y�%ٯnL��PB�~$�ȓ�U`�.��<����8�"O�q�F/�X��)P�T�����"O,��Ӄ��F��I�&Ne��9��"O��â˘,<��waA�i����"O���"ۍ	��̉A'�XJ��h�"O �,E���i`�"5y(�i���y�aJ& �� ��`�3% �Cdc��y��W��ճ�>~��E��y�"ݏj2J��0ꋦfFN%�b���yr�'Z3ZQ�gƣfK�@rE �yr��3{�(�JT
�Z�����y��ɑ{�H�{��E�Q�=��ԙ�yg�0H��Òk6D�$��3a���yR�)H�HsS�^�5����w�ؓ�yBf��v<��V#L�`�lI��O�yRN�AK8�����Q=bܺ7mT��yBgR
$p�XQ�fF�P&��ö����y�eŖ�R��s`X-=�0Yj&�R�yi�J��4�P$Ω+'��K! �yb�&���(Z���Ӂ����y����mx�t�%�PC���F]��yH�8�84�-��ҽ��c��y�
�zx+�.�-?F��#f�y"jK8�x���	�2�y�֎�y���w\p�E-ājy
�Z�L� �y@^�6x���"�4��������y��ԑp���Q��%e�@�J�y2�W����-�T�\�3�kD:�yR�A�\}B��3M-�ݙ���y�e��	�g�I�H"���Pl���y��0V��)Qh��>ּ �"��yr���$N=A5ِ0Z:��r�K!�yB"�75P�ȴ��!�@4�2`�7�ybW�W3�u��n�R��R/��'F(SR�2S8ҽD��-�Lx�z���3*�����y�n�)��"� ������k5yl����B��	�]T�"|�'���"o�?�rq��A�  Te��'Ѹ���� �)�ȟ�����Q���uP�1�{��0�>�!���B�AYvIP��p=񷌀�Ж\P.F؟D����Ĉz%.�9-�����.(D�� \�0���<����@�F2
b�S���VD�b�Q��E)i.�}��l���(!$&����d��	XC�<�3��0h�F�"dI�Ϯi��g��~s��rc��򄞾%
>�snm"e�ܙYv�͛�`�Ʈ,�ȓ,Df����ވG��)@'� ���Bl�<L;�z��"��='I '2a�DÞ[I��FG�gX��9օ�`�)+>�� �C���&l�A�N&�y"�]00��ގf��<+�ֺ�HO�\ ����h�V�SR��C���3��B6ȣ�"O����y�~��K]�q��ȁP�iS"��%'�o�S��M����Tas"X�i^�qS��h�<�c&�!WlQ���ܼFx�D��Pv��}���i��Q���V`OR]QC�
��z��R� lOh\C�hI��J'�АRi���/С	A�(�B�Ԧ[%�Y)I��S
�.�$d+j��_�f�hDO)�~T�>QEB�_պ]���P�5�~�����'�j��	:S�t�� ���M�x��	�'�L���t�vT�0�x�\%Kp��$X<BsfW�N���	bӼ`@��Y�)I����^>�$���"�;&R�{Q��[؟8y�CO�P���+e�G�"`��Ytd���1�4P���	R ��Q�k� qf0 S�F�@��!ӷ�8��է'{�Y�S͹��0���QmQ�|x�o��y5Н�����A��ю�O^؈���{��8`��Kݺ�`앭��'�.��)7�J���<i��P�vi""N
j�0�NSW?i��X3Q�9RT#�95��Rs�H?��̙�:�L��ҩ��S���K��!�� �n��>}�Pڒ�&4���&,G:)..�!��b�~�#�DE�(Br����z?A��jZE�/�$wWP���A��s�:���"P�ADj���o_�_�����'=�m cL
(M",H�(�<V8�D:A-�8#L�@q� ʒD��b�gE�3TB�1�$G�"-J� ���E8M>����=h/�R�e�u�S�_v�'�݁���e�*IRb`@7|��d��0�Z�� �X9P^$���M�%�$7�E8kR
� �Iʋ=�XQϓ"���+D��.8���G�2��'�z��q�ɷ�Z�+��H�/��|�O>��צT�'
}f���wdT�1�N�)Uʠ�C�:�JB�ɎN�<L3b� ݢ�{��"q���`��cV�	��%�[?�1b_�&��t�)����g͌f�����:#`drc�x�<Q�I�D��E��;�޹��dE�!K�lٲH����72�I��D��[�)��p�Ç�	���1QF�_v쑆�	t�ʩ��Þ���f�Y�8��_2;w���*A�;6����+)4��S�ăC� U�X�p�O� )�	�{�Rizq�4�']��
���_�f!j�l���q�Z�!P M�j��2 ��l�MlZ+{�
�+R��s�h5*��֒g̾|�e�n#6�I`"O���)Ki�=���&����^�H�T�ɸ05�{B�P�"IV�R�z���K��G�>��(��v\��$F�D?PcW��@�CF@֚a9!�Jr=�=;�]}0)�Ta^:*ב�P�R-�^K�>�t@
9D<�ȅ�T�[�9�);D���sI*P�2�ҤӦi�j�r`�e�.hA�E��������چaD��suo�*-\x-��cV;�y�kM9^L���hrI��Ί���d�x�D��-+B!��F]�V�`	1���Y��u��I9G2n���'$n���@�2�0�aX/.'Θ�'
A�2dA�=y\��#-��r���2��䅩L y��	$?EjH(3�3I��PN�rg!� n2ܱ`�N��ꐓ_���]�{�LX�=E�ܴh�&�ց׌#s|`�%N՝*?�����كN�x_|���ޱ*��(�'<�|���'����׫wO�m�1D�c�����'L2ء��o�l���)��S�'Y�!ÑdP<�$����wm��y��Ip�%;�Q█b`��!�yҮ7�D���J9L� q;��,�y�\LLEZ���K*�pL�/�y�ĈA��rԩ��N@���f)�y�˶Jtd ��M;I��10#0�yR�H&B�&�)��>�^�4�y�]<�
��a��f9`���޳�y
� �(yta�Ml���L#l�m��"O@�ѲaB7AR��BCI]�¡�"O���7Μ7����+խ�t�2V"O�y�.�A3` ۖL���݋s"O,�����	(q�ņ�Ȍ9"OH}z�A����h+�� |�8��"O��`ή1���Y�d�Z� tP�"O�\۳��e̼P��@ج��A��"O��g!��9�RAW��� ��1�"O�����"bBh	�-�
u��a��"Of����� �/a�Nm�"O@d�ꚝm�H0ӥ䋸%z\h��"OVH	T��.'w���D �JF6�Q"ORܢQU�H� �H8���"Oh@��ү~�*%&�-!R���"O��W̋�,o6�Y�,��	d"Ol(�/��Z�tIժL�H�=��"O�ݓ�䔡O+\�D�� �$��y� �����[�6>.8(�KG�yR03��$*����'��[�	ޡ�y⢜�s�`*-���n�0Č,�y���xEK���J̘Ӧ���y"'��w�T���)�$����<�yr��*K�\�H�2i)"o�:�y�ʭN�*���<R)�L]&�y���m�R���>�P��h��y����_> �Y�V
�(чل�y��CKl$I4!�~���4�y<a�y�&�&8�9����y���'���QK(`����U��y"�޵��m����/h^�tٶh[��y�-�|�6�KW늓*�p��P&���yb���Q� ��-��R���'�y䆹-B�yӐ�M .r�(d԰�yG_+6����G��~9 
$�C��y���:c��NH>he���y�f��#�Ip�m�,����y�B��VMīW�C�f�aÀ���yR�$ֈ� K��;ʞD�RB�9�y�n	�ʬr���!=*�#�(_��y"�L�\�`�A�$�fU�D���y��
7(���BQ+{�zQ��:�y�H��[]����]��Xk�=�y�ǀ� ���P'[?$��� q�Q�y�C@+	�5��K-kMZ5�͟%�y2!����)��K�K~������y�&�JV���B]���q����yZP� �D��t!"T)���"C�Ɂb9��xS	G��ݣ�v�$C��64����Λm����s�f��C�I�R�rm{pN�W&��ifi�	<"C�	� �P@�g�D+1`ŋ4�{UC䉦P��С���DYn�?V;�C�	�x��I	6�� TI�u�P�~èC�	#Z��a�M�H7��� ǟ:z��C�f�E:�+�L�!I�_QC�C�	�r �L�`�X<�,(�C��7:82���@�.�F����6zC�I=X�hF@�*h��6�V�j{2C䉍`d怣PjJ�)����G�7^C�I�t�� b©F#�i%F�O��C�I���c��.����DY+ǂC䉋]
�bD�Ǧ[�~Io�3Sw���ȓdl]��&�<&�yg��6f�H��S�? �C�mH�B��{��q"OI��`T�2��Lp�"O�a�'�� �r�ل@�T�V�S$"O�����B��
E^� �"O��ឥ_A`a���P��<��"O�Q"_�M�!����:�&��"Oҩ	g��J�05�P/��h�"O�TU�ا$H�:���l�ĵ��"O�����о3��ſw�\D�"O8Ա�hK5�
�&��L����"O>:w�J�sXr�EɧcX-�"O���eoL�:Pes��Te�C�"O~X����!l�촩f��;F��g"Ot�+�N
�HRm ����Y80Xҗ"O�!�"�O*���sr�R,Na��"OݓTK�BT����˜ �A3�"O>��QKP;<4,��ᒖ�X�"Oh���ÒH/ ��P ��v<ͺ�"O΅X�A�s/.��#NJ�2H���"O�����a<r�,W�5��c"OH��䎣|�(�;�I��0Jh�"O2�j�,_<A�z00�G	cW��p"OH��e�9]ʄ��V��[4R ;�"O�(Ś�eV4�(�Ћ#�Ft��"O�t���*0VY��蕤ɘ �b"O(����҇nl>����X�b�T��"O��(û)|.\	�,��	�j0��"O��A�腰L{�D)UkQ�`�c�"Ol��*�3
��`�	E�T`��"O��SGB�ma��S�G%�U%"O`�X���KP@�����/0x��G"O���p�J�@��FB�]v�"O����dޥ7��ᅌW�ez
�@"OR�el��d`�X�ą(uU�t"O�逕杵t�Nl�"�6qY�s�"Ov��p��r�vpd.ƄlV�] �"Of5�O���}��.�9��"O�{���~�Tl�����q�"O��Wj�/4u8�B��b�K7"O����Ȫ��y�S�g����'"OI��U�n6&� �=u����s"O�)1�ω'A��I���^�0ؓ�"O��Y�d��]{��rn�	�`i�"OVt*�ˋ*�P�mW�Q
�� �"O�s񣃒b/�Ål��Sb�q�"O�����n���Q�LlAn�V"O E�udԞ~2ȀG�w"$D`�"O�����<q�xcDmXsx(�"O�01���6���d��lb�Cw"O�(�#�"e T�`oY7EX��r�"O^����ҖBRHre�I.�0h��"OL���8����E��tk^iKu"O&��Ƈp�m҃�
����"OЁ�p<]l�ԓG��f��9�"O�J� ԟ4��[A�"~ŔXA�"OV�Ar��=;�U��1W
�͋U"O�x�����r̆!���;Ljd��"O��e�	<���AAŸP��E��"O��ۺG���q���6�B�8d"O�$r@�ѻ^��`��Fz�
#"O$�"ed�-~��bD���d~��"OΈC��\ jnh�C'ׁ;��u��"O��V��(i:-��ƀ�|%���`"O��c��O/c��r��;j��Bw"O� *�j�E)��xDS**�ٓ"O�\k��30+�Z��W��h��"Ob ����
ir��Y�6���"O�P��g�*^<�D�=P�p� R"ON�і�߱LAZ�ȕ:\s��y�"O8}EK�U�M(Gk��"O>��6㝸'.�V��HS�H�"Oꀀ�kUM�ipb�rƝC""OX4��r���i�b�(NS�� 	�'�p�� �ʦJ�$Ո���:W[Ą)�'���[�ˎ���1�B�NU�Ir�'p,����_�hse�M�K��@*�'������Q\ ���сm�����'V�i�#�w/��0�L%̴���'bd�aĝ�c�R����Ŏ �U�
�'_�4Yf�o ޥ����.%�e��'���nT�*f`( �� sJ��;�'�aᦩ�� fm���d�✈�'Vt����);�j�H�%����'M�U��a�'.���&iS��4)��'E�H�GHh�q��J���6Eh�'�@s5�ҿ%� ��&N�uZ����'���$�	BJ5Q�h�'�l��'�1c��;�i�V��Cn�ӓ��'��(7C�0:�jٸe�6\!Y
�'�.9�F�,Np���&���P�'�h$�a$CFl�l�7J]�u��(��'���	���$>�B$��,>����	�'������`���N_�NXy�	�'w쐰S�BBԀ��o�.����O�왕��`�$_'uFn���"O��qR́1=.�84dY�\��z�"O��K%5Dv<�EH���� R"O �B���?<ÄHH���v3�=�4"O����$ޮ
�	���Iq24�#�"O�T���S;?��E[ŀM/w0�l�d"O��h�� ������4J�J�"O����<F��ER���]f��"O��u)�%!vq)��F����!"OJ 4HܕC��@(4/H/I�@%��"O8h�6�׉0�(�0�N��y���� "O���΄�N�{f$��B�XX�b"Oި` �u3<pCp�F
�0�a#"O.X�U��(͈�`?
h2���>A
�CPbE��f���e�F��A�r݆ȓ07r�A�)�]���Y�*�	�"\�ȓ'�����	p�)�MJW�V|�ȓ=��uaU��t�#��9��1��;k��GE��H�\���x^Ty��b��Rf��(��u�k`~���7@�,Sd[7������?t��(��P;!a �ǚU�.yDÔ�BF�� ������)���ĉ�t��WRv@gŃ��d{BeQ�'�-�ȓb�KE@���֪q_���y�@�NΈ�!���S�`h���Í�y��ʠ<�
�p�J�A�4����y�F�:/�^\h�ئ©@K/�y��Z�{����@j�|l���yb' N�E��{Ҕ����:�PyR�	&S���R�dn�pƧ\A�<I����!0��?g���XƊt�<�P�L01E��xR��V�����Hr�<i���+��r�KQ�{Zn�"�h�m�<� Zu��� m|�5�ԃ$3��\(�"O��G�� ��]���4^��=��"OM��*K<
x��aU�S�Tq�s"O��C�.(�V�Q�+�����"O���E�z��x!`Ȉ1�t��"OH`
��us��3��tm�� 5"Oqj%Jڛt�l�)�*R�{:�䣧"O�]yw'�":!�\d��/.Yb}�"O�2�->dz�i�4b�l�"OHY7 }�Rm`i�"�����"O�0RG\�Y Z͐�CBJ�m��"O��؅V�yr �r�8;+ᚒ"O<��`]M��` ݫ%^� "O��s6AS ���r��	:�1"O1�E(ѐ�2��$d4��s�"O*��3(ڒ^�B�x��q��_��y¥���L����i|�P�͉�y2
 f�%� ��X�$s�� �yD��(�
pxą
:�X��Y��yR	��*��p
�c[�	�<���yR�)8��1T���+�0%Z�,E�y�(S.ϤdP�'O<veH����]�yb���B ��8�ɀ+qh�� ����yR&U�a�p,˷�͸Ln\/�y�.֎K��b�h1Nؠ#tmԳ�y�."�u��'T�!E�a��5�y�B �QE0��Ą1!��@�;�yBkL<"Җy��F�rT��G���y��Z']���2)����#���y���)���󀀿�D�(�n֝�y�E�J��i�������Y�y� б��(�uC�$�Duy��	��yr���D-a��єLz�ݲ�#(�y�JɎH^,\X!��<��<+����y�EN�3��/Q�-:������4�y��1����dF�3$�}1�<�y�(�]�0�j͡`Z�H35�I �y��)K��U��,Yb�b���y���b�˴��O"�ġ���1�y�	�3C����Ą�J�%�R�Ȱ�y�+�A�<�����::��)ǀ�
�y��̝i�̜�&U�H�����\��y���B��QR���o�؉X E���ybŉ'�
���� 'dĺP����yr��6¼�뇁עW�V(H�a��y"C7By���q��6Y��uK��Ņ�y�S�7�V`Y��A�LISw@I?�y���@1��ȁ�69�	P�HT2�y����Ґ{�eL�vE�?�y"K�_��Y�CK���rqp ����y��S;�~�Pte��w���2�-�
�y��YO���k��R�D� ��&O��yr��{߈  �nR2;?��)����y�Vj��Y�k�3����mĤ�yr`]�a�4��< t 2��y��E�$$�w`�&���I�yҥ	.\�����z�tT���yi�@�S!L��'uܝ��F��yREس�p:JV����I���y2B�m����'�4���$���yr��0/ �{O�j-�8#��9�y" �!n�Q�I�*hT��!��R�y��|����,�M��DjX��y��f
�۳�O�O|�وt� >�y
� ���3'���i�&Zt�$ v"O�m;E`�0g���P�=:��("�"O4�*��d�^���ăRS
�E"OD<�.��8��a�Lt0��T�<AЎD(~.Ź�3@ ��
�Q�<qdnթ�!z0H
/W!������V�<qR�;P����l�g�<A4(G6n�|c�Gӓ�j�u��l�<q%hș��-��ܦ��EQ�Qs�<a�K�Eh��Z�&��k"����W�<����Q�a��D
Q�1d��J�<��c7ms:�K$�("�,1B�JE�<1�"J9*q��j�#(&B�H�l�G�<���6D�48�vjRIܒ���#NF�<a�N��Lsd�H���:h`pQ+��<iE�b���a�lN��K�b�f�<��n��D~Z�(��ŵR�"��A�a�<��-q7&a�DW�d����g�w�<���U�j��B�6�4��F�h�<aT,�W���q�E��5����y�<y��Vn|JE@$iȹj�V����x�<a�-Q?=��k�B�?�,)�d�w�<����(؆���*X<1%N\��l�<I��FTn�XzdJ�8�l�p�@@�<I��Z�JlXI^�b�p�}�<���K/B
�yF�M�,^�u�uÝO�<A�ɛ�LXūQAlJv}�7JXJ�<Y�#j��RPpC��A��G�<ARaD�lQV�!aT�M&�t"�`HE�<�b蓘o\D�+��T��"�&�C�<��[=gˈ�儒35>�f�x�<Y���>*�q�c�':�{�ii�<�tǖ�{(�h;���A���ӭ b�<�6 
 T��@������@m�a�<�4�ɱX����2DԐzf/a�<�.���i���ܞ:d��PG�[�<�᥈>�V�Dg�0���7/�\�<Ia��=;�����\T	��0�(�|�<��֥^)�R��$�؀��Oy�<y#�^*z���d��D88PT��u�<Yuf�8 "l i����$0x��G�<9���n��A�J�8`���^�<�r���=<6�@�B�6d�	�mFW�<Y��-7����˻`�ʉ��]O�<!�� 0Q�U��M�8;f��b��L�<)&$�=�z�ۇ�*u2^4c`#LF�<i�B�q����-K��D äh�D�<i����7g�x�%,׉_����G@�<���۶/Ct��B́�ZQ�Q�7�GW�<	�L*k��m�F/�e��)P�T�<��ӎ�v�aq���Ƭq �v�<!��N�=�����79Φl�.J�<Y�)1����[�y��!QWH�<Q�LG�pM�q�(D�N�_�<��C��J�L�9cNˢ)<����r�<RMF�w������Z�Z��W��r�<�pkE����Lː�BDڥ�Z�<Y6� �<_�����=J�u ��YT�<A�,�� ��P��@Z!"�����eR{�<�!!�`�D��S!�r�<l�d��y�<�ҍ�_r�6��z�ިAF�a�<��l�u�ș�-ōM�E��O�h�<��쐾o=�4� H���S	�M�<�d�6*��H1셅�,�̈́`�<� 0L���ЗZ5��C@C8$�h��"Ou��D��T� ����4��Æ�^�<၌�J�nq`UG�>����_�<A���Ŵ�b �Đ<�*(e�W�<���	z�Yr�-�5h1��h�V�<q再/0P5�G�	X�4q�3��g�<���AϤ����Y��т�f�c�<�q-@�J9{Po��7�����k�<�4/�<CJ�A�a[�n�X���&�g�<����w�nI�CO�IL�*W,	L�<�$KB,H@�D�]4'U��Ba�<Ƀ��97jʰ`%ШTl�B,_H�<�����d��x��$��1��Yy�<)wh)0z�4����	B!ڴ	�)�o�<!r�[c�mR�K�;�ai�"�S�<�2(S%L�KӮ2��w��V�<V�ͫq �)@�N�d�����CH�<ye$Rx�Uk��
8 Z�Hd*Y�<A
oa�/��q����T�A�$q���{ȴ�I�$ˎ���KV�X�n�.M��iֵ𐄐�GJ��7��5U���ȓS;M���I�lTL;��� �:���-�T�PR!;n?����l,K<�,�ȓ\��=IR�^$sF��Wj��LVL�� ��(R戠��q"Š5�q��J\�ej2-�:d��OɁ	�ԇȓjr�(r�%�=�Z򇋇{�H�ȓD��l	�B�0>�ة��L���NL����u�Ѕ�G�, <�������q�R'4� 1	ƫU+0t�-��"�8 ��)9 �u�!��Eb�'>�@��F�S�H��Q@I^|���
�'���Jʝ~�
 a��?hFp`�'P�E�1%�7.F�[�œ9�E�'D6��ec�?\
����K�)�����'!.!j��]'M��Mۧ5
Vp�
�'�(��ѫ� 3�> a4��=6``a
�'��;���}(���ˌDy�ٸ	�'fn�	�&�y"8�JQ+�>�ʘ�	�'3��"��4d\H����ȓP%�-JBER�E���rGE@����]�R�b�"K"�\س�ļM�,܆ȓ"q���Ð(8�u�V��!1�e�ȓ{��u�����T����H氅�}�����żrt��B7>������d�Έ�j�i��]'Fn�ȓd����KN�����iZ�]sH��+��B�,b�@���8���ȓL�@��#!�b0���7h<���\y���A4�����2g@HI��#]��#ϗ.�8��A�(bx���}�����!�9;�%��F��m�H	�ȓ/�ZlRT�ѲZz���C�?���ȓSV`�q�%B�aԈ��EJN�%j��Fh��O���'�P,<��]�ȓ�ؔK��4�D�ӕ�̦|Z�Ԅ��j)�a���	��i�"���h|M���Ԓ!W~A�1��Z�@`�ȓ�(�Yb����T��ȷ_�t`�����cG*G])�C޻E�@8�ȓR(pP]y��(cQT�2ئ$��"O �Ic�I�e�Mh�!�!M�ʹ�f"Oذ�6W�����֋3{�d��\�<A�KJ�3�hi@(�]���J���B�<� n�#e�J#:�^ �i�w��5q�"O��I�`.���w����䐓"O1�m\�cޢ�1'_1d��dQ%"O�Lk�'�59:45jwK@m�"O2����r$���f�� f�h`�"O�9)rN�c�(�:p� {ʥ��"O�a�!�4��šp%�"+`���"Ob��C��Xa���s�7�b���'�(��!�5�Xa`0%T+�J���'��e���#�x�K�Qh���'��+�`�i��2ք��'�|��ubZvA�tX��A!��\��'�`["��xt��D	�ܚ��'f,�ch�7@m�V�(�bT��+��= ��G'H�mA4�	�ȓz�����-ѷ9\2���&����|��@a��>-Tj��w(���i���CX1�Z@��o��@���ȓB="M�s�'&$��`&$�%����ȓI{�@���$�]PC��ä���%��"lڽ1���Ɔ�P^Շȓ,�1!g"̺[�&h� �"O��ȓ>R��W��$r�BA���%#�4H��!�8Ê:v�@��Ս^Ϯ�ȓ2É�Z^��Wg5��a��v,�!!�u��v&�>:��ȓ@����P�ȕ:�~�2��G:p#̵��*�Z`{���W�$��+�4z�"��r���Ru`Fk[xDBh9=�Їȓ3�R4�FBǺ�E��gӴc��̇� 1������7R�5lU%F0���l��̰��@$�"��$`�����oQ�q�d����!uE������D�d����l�j��3 �3e�LՅȓ�2P�u`�	t�|9�)̭iKȘ�ȓ �<�d�^������,(>���e�s�+�1S�Xq�C�)�Ć�QX�Qr�7S��0�B��B����ȓfR �f�W-3ޘ 1�T�=��ԄȓpŊ�0���Z� ��<l��̄ȓh��<XB�5�]2�H�Y9��ȓ,r*i�ghly��] 1�,d���� X�>pH���ǿT������{�,$"!ZR��;/�r=�ȓ��0�K�^�NL3�(ǾM�p��ȓ+_�����i�t��a\?|�m�����B��P�pd:� ��v��نȓ"_�u#��Q�F��\�;�R��	v�������.���� �L]d4�-�;D�}��<D�p�H�eR]B��K';	8�q��/D�P����'ZR�����\7I0����+D�4R���xpnEX�+V�m�9��)$D�D�򢔀4t�
�\� Ai4-/D�lc��LE.��fO^�3�����,D�`�V$'pd+��9,E��Q�?D��D,P�
�ɫ6B*
t� C#c?D���獢1�mф�@,^����<D� �4C�/6��� C߽#�:���9D����LØ2��g&_FP��+D�d�0%��O"�Q�°$�N��D*D����U+&�@�+�ø+D�z�h2D��@!#E	\��9h����D��i�O@�=E���&&K�0�B)��\4�e�R�,n!���[��z#� �y�Æ!;P!�� ��Y�~�<uǚ4pY^��"OtX�V��
7ܞ�a�����"OE(҆�-��Q���ļF}JT�e"O��#�R�3�n�"6|��
�"O�H8�����Xx�MHSqfi[��d�O���Oj�;w��J���HE
^�*��)��'�f���o��'R�;Uo��z���'���vNȝM�f`�A�ϝw>l�B�'��ҍ�~@����}'���'��ybEAV�0���*�v�r��'l�lR���<E<��۠=F�8�'�l1���I���H�� ȄʓB���`u��u�fZ2)�A��ȓ� )�S_ N?2(��н]�bH�ȓ.��-��
Y�*�hѓ"U�I��`��w)��
'.ƕDڬ	�#��}�X\��e��c��ͣ~�$|pփ�)C�����!��!�Q�ld8�b�*H��'����ԔȠ�ϔr< ��"�4؉�EK�"�I��T�Q�Xi��:��o��8�ұ$%�@���v��%�@�L�~�J�z�W5�F���G�Z8�ǩ��_r�
҅	'o�9�ȓy�ع��,q��)�ACT�Н��FN^��$����Kw'�G�ńȓzLnMI���-+���E�T�9�*��ȓ+/ u+A�L�_�̱�MƎ%,B��(�����#ƫLR�1�JF
6�0y�ȓh�ɒCU�3��pѠcɜt|d�ȓ-���!��T�P:|�6��(��`�ȓ����݊a�RZ�KYT�d��ȓ5�d*D�H^d��ɲ�#F�rp��/��Mң���X,yA�X�F�h��!���Gɋ&r@��x!"\08a*Y��af������<Ft�H�c�*nN��ȓR���E�4%Cf ���>K�4���3&hy���	�c���ӀO�;gH���ȓo�X�9S�БOs���զ�7s�4�ȓ�*PbG���OCL ��O�/O�>��[8���5�b ���.t�61�ȓ?N8=�P�S4(�ڔ)���&)� ��-�09�`/R�Zd��OH�Rt�Ȅȓ3�P�Q�`��n[�$r4GҊw��l��V͖�9���%(�pm�.R@���ȓ�(���۳_fB�i�CX�ZR���i�����טPÎU��<�Ե��/֩�Vb��6e԰i2jF�%���,��+0'�'wV&��t��P �8�� >%9��ɿ/�0��M��5�ȓT8��r��';��p���cq�]���r\�`�_1I@H��I܁p��ȓCӰ��rLI;F*�s�&A?yVv=�ȓ�⭃�K%P�Fh3H��(�ȓC�|��$��!h�-��dQoR�!�?9���0|
֠R	3����G.!�H!���d�<����K� x�4Ę�r�DXaHa�<��	1o�4	1�b��*�[�<I�쎀e8�m�T"D�F^bh�L�<1A@�1)����#u���(7�P�<y�*�^������S�
�8��[W�<i����>�|��X�u������m�<��%\�J!�Th�"��� ����g�<��ģ,�, ��l�	2@ +w�]e�<�Ύ�kT�(F�ֶW����BCEd�<� ���ĕ!%@�h��J�q"O pAPf�o�J��P�!s��0��"O�ݻQ	�e����m�x�c"O2P�[6~-6��cϜ-O�� x��$�O���IB�+�
� ƕ�v� �X�aȋqў���I�+(6Qi�E	�:ؙ�l­w]B�IX�D�KEN̋} ��P�E�1"2C�	�K\1�rO��hXN���l�<47C�ɪEEr8�ǃҋq�,* �R�B�ɷ^k���$K*d���J_����$h�P��f�.1 4��$D�)�t��'&)D�(�f=R�|��%��g�(�4n(D���t�:WF,�aw.^�
$�(�E!"D���r�TyG��`�%юyK~@h�B>D��	h����Q5R��K D��2�J/��aJ�P.t�t��g�0D��!�I7s��PǪ1Kz��/.4�x��Z3(�$��9	�����ψ|y��'��83�.i��a�FĔD�FHH>I�
tC�O�z�V�ZP�òY��X�ȓjɖ��p�O�D�4-Rd̗�~ނD���"�z���vp!:A�"Fв$��AIEK��kr�ꏢG�Ω�ȓO�f����?����MJ�!-�=�ȓB���)Q�+B�Eт�	�hh��7<�h��C�>���!$��bٕ'�a~b J(�4�^�����%�K��yb�E�'����,�X��� �!Ƅ�y��FD\q�߃}z�A�'�5�y��Υ���G�6f�\]b#�'�y2�~n��;)U2�� R��5��x�V?z�� �#Z$�("F�V w!򤚧zh`a[�j�-%V�E��MS!�$O"S���e�*h��%`TJZ?!򄞂<6{���8}N��FI>X%!�E�m��L+�  �(�V����A�!�d�-!`T��V�=/ڬ�1��
�!�dD�l2�����X-�\J��n�!�Ę<Z��}����;��S@����!�H�xX��)'�_^*�k�B]>�'a|�!�2�	�B���ta���C�y��firAk�,Y4��`V�3A�����2U���ȈDp��#��2<(�%�ȓV �@e|o2e�b�+NZ����}K����:b0�;���*"݆�Bs��2�2�b���lI?��5E{2�'}Hq���"ŜQB�&ɶ&錐i
�'�r�Y��u9�	Bo�H@��	�'h@�5��7\��A2��F_��I�'�6������^)80�7C�<KHb)a�'�L�G�Cz���V�š7���P�'$b��ˋ*k�"!3����0�ȓ�(���̔�_���Pk@�6!�M���g~"�E0��]����8G2\������y�#��^dɁ�P�A��qS�;�y2���J5(i�H�#���y��č�y2ⓞ)V��3��Уl}̵{D���y���g�\��]�9�S�^�y2�L90���YS��]�b�s�I�!�y� P�f��$IfU�0�7�y��2n$f��*	�����ꘕ�y��N�4U^����*����V�y�e
)W��!*2+$�L
w��5�y2�K$Fh��R�#'�𐖠��y
� <�i�f	�����S��}�"O�ʅ�^\Y ��BjR��ܸ��"Of�1GO��V3*�0G��-t+����"O����l١�(H��Z��"O<āGA�$Қd��C�h��"O�=0�G�x��A�U�Ț��Q�"O�l9��'E��P��n�L��졤"O6�I��);�O�	ƌ��"Oz�ە@O薌I mηP���E"O&H	�
<u� =�a��$4�؁y�"OL��u��>�n
����HC�'��Q��Y�lA&C#�T�C�'����	�+�<h� �ن�p�J�'8�"V��',|���k��?�Y��'�p�iVn��3#�U��c�;}@�r�'�$���ʠDSB,3��i{	�'jN�̏-;9��0�mK((qx$q(O��OZ�}��0�����,h�V	�0�
� �vm��~R>�C�֘[�n��%�E�5��i�ȓ��WH 5���x��4 7 L�ȓb�p�kaF�W~�`A�%6�ؠ�ȓ^�zYi�P�.��$��F9W߈X�ȓ�r�t��Q}¬�U���ȓ@�D��'�S&4�TMIV�ͅy�����|����z��# �|�@IAL�
�<�3�8D�0C�;>�:���� 3LLu"��!D��R��%CW�y�aO�"g��)�&%D���F 9ig����М�,u"��?D�\���ڷF��PY�G�%n�b99+?D�dK��!`�S�MO�3�P�<��Vy��58fFE�2�ҒUݲ���(	�˓���h��d����%�ʎvevP���K3�!�&!�T�� ���Qba괧�&�!���K�>�[�ށ�l�b��R�!򄖉}vޠU�3>�p 
�e�2k�!��R����d-N�5δ��E_:Kp!�$�q'.��E��� �T<c%�H~4�O����|
�O7�H�gl����Okux1�	�'*H|� Ɛ�j(�%�>s��A"
�'8�q�������T���d����	�'qt��e�\�N��Q���Z	�'�������z�3�o P���'�
D+���Xn�a�PH�y��er�'14��G�^;\N��w�FgD��[��'����|:P���<AހI��>'#�0�t�YV�<���4f��kd˼Q��¡)�{�<����96pMb'�ܶ�J��db�a�<��c�gb��(1-b���֍a�<���
�%� �It�S�|{�$Z���E�<���I�Lø�1��V!:�)��\�<a��^+Y��W�&XZ�Ы���X����$2�
S4�'	�*IwA�A)�v����L�H9���ߍ~Tb��v�4I����족�˙',�e��/Hz�u�ȓiU*y����P�b��,��v;Q$/r�A+�.5Qsv��v�`-�2L��1xz��f��<{j	�ȓPa�� @�	<؂�
f/5Hp6��wwr��-� �N�ʑ�J Dx��	{~r/��FF��.֬z�b,�Eg���y��� *)R�["Z�m�}�u��yb�޻#�L5���ߢ<�"���Ԅ�y�h�)��X9 �K	0�@ѣ�T��y�@�L���K+��<��^��y
� T���D]D=�� �r��D"O�r���:R
�q�N�O�8EQ'�P���pO״�8��ݫZVP(U�"D���#@�=5"��P�`	t�*��Ӌ%D���3�I�yn���#�9v�u�1D��x��ޑO� |�F�\�Wn$��e�;D�Xx���'_[�y�CN�q��AIt�.D�,y��L+XB=#�M־�� pv�,D�p�ć&-������T��`�!+D�|�W�S�(��,�rL�+�\\AF*6D��`�D.\��4��H��I���a�9D�\I@e	�B��z5��n��D`F�7D�<R�n]4䜌���D �Ԍ��+D��R����d2Pܨ���#�b��7 &D�䨆�E_E���~R��ĥ$D�XQ�
Y�V�l���I����O�OC��<^�:PR4k�*�@�
\abLʓ�?��_�l�i��J�6�bF�J6s�����;-Dp �kL<6H@�鰦P3v[��ȓ`�|%�E/\���m-X��9�ȓ~��ɢ��Fa�LA ��"\�Ru��%5�łBJ�V<�F(	H�.5�Ɠ|6L��*��n$BD��z9�X�-O���΄k̥��&,�)��r���d��@��g�P��m�4�PCY��j>D��0j��m��p�Z�~�t��i<D��ئM�q�H��$��`)ҥ��.D�� Eǫb�\�.�!�E��c&D�)3Ï7�tA9��x���P�P����
|�i�E� ��`Ѝ��/�B��ȓlt��ࡗ0Wit$z���>K����?����hY ��>ju���|�x��ȓD�t� �N����(c���P��Մȓ%�x��$Vy�4¤h[�e~ƀ��ON��s��ܿ4���)ѦC���d��9\*E� b͌Z�,�	�G�*3$���;2Hy���Ѻ>�lX8�m�K��<�ȓb��h�F�!M�`��fL;I$^��ȓ�T8��M�NV�����P�x,Ԑ�ȓ���b��8��t#S�l\|(��nވ�G*��.���#!S�i��V�qr
ز�L�@�&�n��ȓw��!��C�":瘈�g�U	��ȓ&6����� Z���t��+���2A̽����%�p���<s��J0,`#  W.:� ���$ȦspD��tY��"<�&����8t4��)Z�L�����35���k*l�&u��8bPia(߂?1�ET�/���ȓ)�]Y��CQ��bǂ�@�f��ȓ-ty���¶ckZeK�(6X�l��B-�A�R�Ń} ��f�浆�b�����V�zAƠ��(��9����P�c!�( �<�p�®E����!����J��~R�*E��O5��ȓ?��bQ�ԌZ�푫l}�	��=D�d�"יTg���O<n㸑�Ԇ<D�Tz�G���1:��M#<�X� D�� �J�U�݊0e^�{�6���@3D����НK����U^4,�;D��zTĐ�?�y��[M]���p�<D����fG,F�i���x���:D����@_ �4�����<���,D�T���̃ ��R2*S�z�����'D�� \5b�gZ,��H�!��W��X&"O��jq��kײx	Ȍ<�Eb"O��aW�؈��\
'���`E!�"O���`�kE�Ih�+��f�ni�"O0��&H���B8�d��H�@T�%"O�Y*gؗA_N�[��#q�(��"O��b� �1��3��;����"Oʽkw���4R�J� �F&�"O�M�f��bӾ���	=$#f�:�"O"�A�38�С��)��0����"O =�W@!~)�acwȌ0Q��
�"O  �e�.|�LqP�G�n}ހ�"OĜ�p�[�&���K�M��ڜe"O�`Q�i���R޶	up"Ol��7�H>4��D��ܦP��qxV*O,h����n�ؓBX�[����'K�0P�� �% 2J�K�^)0�3
�'�!���:��@�$O�L���A�'�\EH����x@ C���{��a�'�=�7ˇ5�V�*7�ԅ!E��'��h�ӧ�1A�����o��ɒ8�
�'��0��K8��pHV��&Җ��'�fi��8pB��u�N���9��'Uz����+&�����c<�����'��l+���g`�(Ί�}�`�
�'�� 1K�洂�'� z�j��''�<�vn� l���e
V�>��9#�',�Q5鏕KA�c�[�3��l{�'�r�YG��N���k�ȇ0��
�'�M�$c��7]�(��7��i;
�'ؚ�P�ٌ
z���Bҿ�0y��'b.U`���@���N&u�K�'�r��a�Q�n!�E�į@$���"O�� ��Hq��d AP�F��""O�@�ZR`��8��Im�� r"O�p���E�f�z���N9vɠqx6"O��؃E�Dj"u�U�����"O���GcX��u��&؀|�����"O��0���!�Ba�䐫+|x�!�"O�����Py����7�E�x�FY�W"OV����x)�!�!{��[�"O���W���-� ��0����@I0"O�,��*ޭ*�)�Yp���"Or�Av�?�8��l�-�j��"O���/F�e����V',���.�!��	��hc��.h �� �ϑ?2�!���FC��"�Nꄝ�A��~!�D��tE�,ƥ�;u��aVMV0,i!�d!ݴ�ㄨ~�$�� ��vq!�$a�l%�foR$a���c#$�>5!�Ę�@�\�� �S�>��DIO��!�$B�pU0���g�rYR�']4B�!��-
�x���k���AL�4�!�$2X7����ÓXʰ]��do�!�DF�tT�"��\R��p䋋!�$Q's3�!�hY�RV"�#��Ppg!�C� _�yjflN��񁓠S�-Z!�$~�"H6K�8I'V�!v���A!���0t�z��-�>'�U�r�Z�9'!��DQ��e�G!2�~$8���!�ė�5;A�#�a����!t�!�d^��R��J�NҀ�U��'�!�7k�
1���N�Y�amG�r�!�	��&�9�L�m+������!�� ����APT�,b"D�ar��S"O\�
w��=+ؼ�@@Ǥ8�Y��"O
T�d*�3L��9Ơ�[o�	�'"OP]�q�Yw�l�UF�u˄b�"O&��3 �<�ly+�D�_��P%"O�)��,� C����PW�Yl*ȑF"Ob���")4G��;��zb�"Ol��r	[^u�À]|�: a�"O�ڠ� �{v���Z�{���"O�p�q���������C�"OL��Z3�RܪԢS�Hֈh�"O"����2����'�b*P�� "O�*Q�.w�DY��f�.I�=�"O�{�䁚0A�2�f4<кm "O��be\�4��kA��:�N��$"O�E�C\Khp��@��z�n�g"OI�'�\"��q�" �p�r��"O�<"����5H���-���H%"OPdud��
$�Qɀ�˵>�j4I�"O �3�HЬO1t�a��1m`NT��"O8`ꡈZ,0G
(e�$S.�(�"O�𑬁J�t!oD�"CP��A"O�qREʴc/0�nV���.!�dг<U�eB���F�b�͌�Ar!��4�L��É&�R�X2J	�4t!�dP������#�l�&�"?n!��Û:�:� Њ��z���ɶG�!�ʶ#������9�Nݪ��W�J�!�d+�J, �dG�?�����9�!�dڍ]������#5�I�|ќC�I"�����ŉg�Z�A�41ΞC�ɽ"H���i�-PFDxD,��yP�C�<T���c!�̀<�D Z��̨u8JB�I;x?�Y�K�;m���g�~} B�I%d�x��_9Y�������,B�ɯ�ua��	y��qXE䋳R��C�	U��M���LI]�1�E�՚5�C䉪wU�x�&�M�	%�� �m�(#M�B�	8�t�5(F��X-]P�B�L��K��	.Ek�y
���9d��B�F4�	F�42|��1�jB��,th���z����^�KDB�I\��T�h {��ȆB�I�lݪ�+�-�(b�.�B�C�>��C�	+-�ʩ�Ն�d��8�PkT|��C�ɚ4!����P������L�<B�#E�Q�%]�NR�q"a�1o�B�	�^�HC3������Y�W�p�
�'"���[b��h�こ�L�RU�
�'�6b�![�?��`c�o�(}`
�'�ؐ�tgY�`R��˂�:gI��'��R$�=,���Ɨ4:����'�H���Δ_����"Õ%g}1
�'.l�3BƆ�.�v���l�P�*P3	�'b%�aR�y��i@>'�1��'y���sD4)aLa��QQ0pZ
�'U��R��6c������)�'����4�_�.F�asA��-@{�y�'�����RA]�0��j�6�P�J�'<����X?m���uHU�𲈘�'s<��_�$�z�c�
(��'6j�X���	��d��|�~��'��I�C$[�j I4�;?��k	�'��mȤK]?D|8�� &������� $�F�&� ����p7���c"Ox���|C�\�#�Z p��e"O���1NO�,L��Џ!���"O6D"�ƿw"�A�t`��-�!�s"O�ڰ��IPB�ޤR�`hw���yB�<����i�}��|��K�y zIr��D�ܼy�A+�䓶�y2��bY�!������F,�y�'�<.R��ˑa�,
�R%*����y����d��P��4�����G܁�y"j,1���6��*2�2����ԅ�yR(@6�^��d΋�3:�ٻ��O2�y�H�sP($jsl�#�2���e�yr��/{ )����!v�8�a&X��y�K��N�LMP�΂��	8dJ��y���0:�u�P�E,	o@�ϙ�y���6��2��(w]`Px�R�yR�&����Իpx	��!�y����1�Jv����1���y���y�v�9P/	��\<2�*�3�y�c��x�0�D�ا'��p������y  n��p�SZ#:�$��	R��y�D�&<��qɇ`
�P�V��)�y2.5�ś�G���h�㛵�y���,&"X���ҹK�-ڤ��yb+M�e�j��emw�ޥT�� �y2��rȤq" D4m��v�R6�yƃ�?��8���7���p$�y@�sV ɷ�"6���qť��y��]�v� �!����3���;�F�2�y����m� O����ˤ���yr��i����)
#*�&�Db_6�y�
J53�̸�b�&4����ȅ�y�Mߖ2�L���Z'O��9��]>�y"fX!¡��Τ��Ȣ��yrK��IZIzw�:��l�bJ��yn�@�I`��{�l	�c��y"kC�	a����\VU�vJR��yb�%AY���3N�조ࠋ��y)$���I�<�������yb�D )Լ���������#�yb�u�ƅ�'pq��E�y®�6�tzt�+��� ���y�$A��Y��I�|t�u��bX#�y�d�2 �R�FP�pN��xv%�1�yb�V�o�h�&�e��� K�y¨J��ġ�N?aI�]pS��yR�;A45�J�.��H��E��yB#�u�xpG��[` {�n�"�y�3a�:AY�C��y&�)�	�y��ߖ5����&a�����SsϚ�Py�
�T�#���J?@Z�ώV�<A�Cӊ_Ȩ���<�l�f S�<Aw*�'��C�B
_�i�T�GZ�<��	+,���xRe�2[�j帆��n�<1�Dk�V���o�+���`&Âi�<����*������'t%�� ���N�<�P�^z 4j�l��>?"ٳ�L�L�<y$��H33�Ě
K��1G�@�<�s�ɻBa�3հ!G���%�Js�<1C` 3>&@Bb�ߑg�ج��Gt�<9dKI2)�B	���P������m�<��ǌ=ҡ���D���ف�h�<aD$���B��Q;y�L9�&Qe�<� L�3��֢R���%Η�
IDE؅"O�m8p�N�<8��l��@��Q�"O��2U"Ѥ	|�ja&�T�~��c"O�򓇙�Im|b��w� "O��V��˄�0t*_2|�*��"O9��m��ZEkħF��"O�8�6�ƷJc$���L�D�N�	�"O���E�^jr��&�L��,+!"O��sՎ�q�܄(c �[�N�0�"OZQ��iT�����l�
�zW"O�-Y��9
�&IU��'Q��8�u"O� �Ů�d�[���2ܼ*�"OR��d+ݐ-R�ݲ�o��e�r%��"O��	e�׆\�Pq�`E�-�j�:D"O����e��d�t�p��Ђd2P=�2"O�ZW�P[�j�H�)S�Z.1H#"O���2혇�XE9Ї������"O ����F.���>T�N�yt"Or 9BOS�7�H �D�gODm��"OB4!�F�ґ��B8`>ʹ�s"O�X1�Ŏ�$� �JD��|�`B"O�1�U����f	�:R�`�G"O$�[pkȕFLFHq� 9��5"O���e-�M�,�zfCH�K�8�"O�]a��D/j���DN�+�dՉp"O.���
c��#�⚣2|nثS"Oh��pG,<���7Bd؆7�&D���G�V
��Z�LX���ŉ&D�h�ǧ�P��rT��G�\5�N#D�pQ¢�J�� � ���i�$"D��)�$�2,��9A��M\Ҵj!D��uj�*��؃�ɑ�jH�V�)D��&��>64�HD�.;ht	f�,D��ą6Kn킓�ěl��H7�)D���L��Ҡ��3-X^���!D�@ e߇��Baf�
I���0( D��Q��A�<�+�j�9�q��+D���.R�}ɲ�Q�
H��|�6"$D����9��׀�8W����*"D��ba��+�M���8D�|b'�-D�ԑGc�H�h�X4�7V�q��-D���sR9v��ԁ�`Q*kV�ԈS`*D��P���	X�5�'P4
z��J0&+D���#!Wy؞H�!�_j���'D�8	Aa� E����HL� �P��&�&D���gBf=�P+�.��%������0D�@�w/�>O�a��D#tb�9���0D����P6�T��g�]*j'�d�G�-D�@���\�*��K�k,X�!�i-D�Tf���|��e�4]�py�%D��n��m놵�P̙�GN�b&A#D��@���:UM���T$�2R�� D� X�c#iB��Yf#O;�
���I>D�\�#fS�/�b��F�8򶀙�'>D��H�@ע;�H�qFE�j��ؒJ?D��@V��]A��[1���r��(8�d>D��(���N4��(����,���׮?D���&b��Ea0,�㥚 +��q`�=D�عdMۛV6�� T�>r���EN=D�@[*ǜg� �I�K�fR*m��.:D��B0�V3��h�$�MO�`�,8D�� �#�6
P8x�j��|���0�6D��h7c��5�F�H���L�F���B4D�|3S,�"|`� �D����$7D�� �l s�3�)����za|�XP"O�� �AJ.#>��cd\C��0�"OZ�&�Љ�IZ1��.s9�=�e"O4�8a'V�v�Z��ŭѠ`%
I�0"O^$�%�Q5n��騶��:F,6M�p"O�Y����.5e�5�������"O�m�f���
��j4bf"O�0��H��d��$��l��T#�"O|�z�B��W<a
�dߔNE2�"O� ��'�#?�0�I��=���{�"Of��"S&㎙ѓGA���[4"O�p���F�lL0�Z$�T�gB��SD*O�1�J�6B��h�\��TmC	�'����o>en���M���M�	�'�՚���P/D�ITc�
�����'��LA㤉 �v]Q����xI�	�'v����H`�c�E49��S	�'r�p�b�A
pyF��� �H�!	�'��@%I��q�E��	ML��'\�	����1��t���3l��'��aP�ڹu�u�4�ъ}%��:�'t�-p�ɔ�<�|�n�M�r���'J�8���iz�$���\9���'��tXF�=�А�6k��5;�<�	�'��D qH� D�pt�f$My^� 	�'D��A��-@�}a�c�.E��,��'�|�(��OHL8TK*�\�B�'���8/Aqzļ!�g�-/j��	�'�l�����-V���4>�`�y	�'�H;��:4�H*�P�:hq�'c.@P���]¨������`�,t�
�'t��*��F>?�!gnQ��j�
�'�F��&
�)ف�@]Y�@h
�'֘񐎓7jԠ�-I�]O�]��'/p��`���krmTaj�A�'�H܁ө 6pA��a�I�2���'tx��S
7Z�Y�pk!� i�'ڤbv#ݨSܨ�B�����lQ�'\xQ륉��/�$1�RDΕ|40���'`���2�O�+x�IKrdO�c7�%��'Gt�J�'mrf q��V��<�']\��#���9�a㐿�\���'�h)k��X2,��0ao�v��A��'�P��D�U���KA j��=a�'�:l�T���Y��03�Փi�Qs�'D�9�r�ݘdB�P�NZ�/��(I�'�,PA ��!^�Z�Q�L#.�l��'=�H�,S Q"n�HRA%-���
�'���¤ �;�H��dȮ(��@�
�'�-���L�h�x���A%$0L��'�D��&��'�%�O/�x{�'�D��ĕ�9s��[�iH��RU�
�'}� (��G��aJ����9
�'_PX���U_:Mr�ɔ��i	�'���N�$�q��	*G� �'ւꕏ�=jA|�b��F�#�X�'�(p�Ë�'�XcP˅�+��I�'�N��C#N�.��;n�'��9c
�'*V-�D �vY�A�Ҫ-Y�5�	�'�F\35�� ڢs� ���%��'h���4,%�(�H33�`��'~6lke��+$��pt��W��Q�
�'f%� K2aG�ir��D��
�'�1�L�E�D�) [�Er	��� $D9R���^����cd��H�K�"Ob����V�b|�P��l�^L+�"Op�q�*t�~�p��[�X�����"O ���d�(< ��@�Ə7��"O*@ b��f
�5k�e�:"�C�"Oм	�E�h�X�d��r���@"Os���"[֡j�?Pь0�U"O\�����$ie�F�W3H�F���"Oޜ���=���Xя�2u��`�"O�hQ�B��m���`�K�v�pu"O4&l��y��T9�8~c���"OF�Я�%���K�lL�]_�"O�]�&K7Y�%���&Qhj��A"O����p肶�J^��5"�"O�XZ5lW:sT�ö���	���r�"O�@ NB����C��4�=z"O���ȇ%S8��j3&�75|�(�"O�!F���#s�	��'�3��V"OKB/l����Ť��A�N|���C	�y"�K#�Z,H���=Z�t;vLS
�y"�E��vȩw��0�,��#�y��4;#���!&è�j!ZBOC��y2'M�|��D�A��pp�NP��y��N'̙��W�4����,F.�y҂גt2�K-t��o,�y�$O.��I��GW u-��ꂨ���y�+Ғ2�p��R�یv�J$XŠD��yRHqQfE�RAP��9�CNH��y2�߉T���CK��J��FS��y��P�u�� ƌS>��QT	�7�y"�+D�@�JV�H�j�@�B̈́�yr �@9�F�O�dX�y�	ͽ�y��QA�4���Y�[�\m�wO��y�d"��K&��/T��12����yb�N.l��ty���9�@�i� ��y��>Z�y�N#Y$=��Z��y�Gpa�J�A	�Q3���0�����'��dEGP�(�s�ٶ%�ȉ�'R�܋��.G�&e�EVlk��K	�'1�d[6h�zb@X�A�*f��<��'������(2us'M�9[lʄ�
�'%�<���4aꈙá��`���	�'X�H�!��1_	&XB�j�_c2�R	�'�z\�-��։ipN&Q2�uI�'i���$�n����<J��<�'@밉P�}�d��sĒ B�v ��'f�Ʌ�K%	k�!S`E5f�Qb�'��E"�A���6���](bEZ4X�'�� �)
5d&��{�LP=h+ ��
�' ���&�[�ΘkQ�20\q��'�*@�ۡ;��uh�C?�����'��(㠜��|�"�δ]a X��'�\�qj�< �"lY�ט��'�z5�A�0��*�W�x��
�'$��!��A�/��d���.�x���'F���qd�$W�,�֏N}kt��
�'�X���e\�1T����'�����'�
lva�Gv�@�@3�:�	�'�,d��*[6���!0x�n1�ʓRH���uØ1���$b9?�Ĉ��H	�u�%�:n딴ZfB۹S�Bx�ȓj6���b,N�|�£oV�T����DVN�x�bH@C���n��H��D�ȓn�Tz��D�m� !��=����S�? @ pBa��IB �ajM���52�"Oj�J��!�R���h�5̢M�"Of�P��q��S��N�@��15"O�$@I c���3���>Ԫ�"Oʙb��O,W�	�*]m���"O���a�"C]�H`wV���qa"O}"v�� 1���sa�E��@��P"O�)s�O�e�:i[�
 !q��"O�w˝$Lo��롄G�un���4"O �Zp�2�`�գ��S1V]���Q@�<��M�2eZ�z���[���U
%]��	O�)�?��b��X����j:�PAc�<!D�L�m���a��LFʌ,a�F�C�<�)^�B^x���WP�\8eC�|�<��bҭ&�n��F"����c�y�<y�+�:�ly��/�\��� &��\�<��@��g���
1?�| �e�Y�<�Eg�>��w�V�Y�`�U�<�����D\����� W�����H�<A- ko�4�G�� m$���	P�<���
v��-�P�K�K)-���f�<�E_(X{D)��8�`8�w��m�<!pN�;�ʗ�#�~�A#`m��X�>�f��>~�(��� 5�����)�D�<i���A�T䛧�H<_\	�'�Z~�'�?u�q ��;\���>](���(D��8#R	n��|��4#�:�>���"�0� Ƅ8P����^#V���ȓs0p���%'�J�#/Ou44D��:�jՈD����d�c/X,��4E{b�'�� ���v����!C?']$+
�'X<@2�j�#�n<At�0 �E��'�F�G٤�p�:��#%z�=R�'�.����G�4�TM[��đr�u�
�'Q��B2G�0lZey���&J���'�
0h��ٓf�����aT\"u�H�,��IC�xT����}q(]e�@L,�C�	9R� b��D�G�1 v�D/CC�I�}<: �aΊ�p4u:��ś0H8c����ɐ(|�4�q�Q11gh���	7�C䉬[��]�aN�6c�Zٙ$G(��C�ɻJD]`w��~8�ڴep�d"Oؙ��F�0��
�J��*iY�<����=��,(x�0�K��7�(t��^�<�Ph_�Q{6؁v �	a� ����V�<�r�\�ju��e"�_����-�x�<��o�N�Ը�b�?u��Y��	t�'�?%���)I��M��o�2H��R��7D�P����=@ 岴	��1���2�A1D�@@�K�TVH�����{B`$D�(XS��`8�������E(�=D����H����qS�L�M��ݰU�-�O,�I,Ph�P����6(%��2�bWv�v#=�'��>IBt�=C���酦�n�`�)�O��'ޞ#!E��-�L�(bPc��J
�'�(���C \�A�
K�0l�*O�"=a��5g5~!q�L>��r��@�0C!�D�-3�����cŊ��1Ԥ7<Lў�P��K�M
"�tQ���W:^�b�"OJ���A�ܨ� Z>:�a
P��z�OY�R�X	p1W�.l�(h�'�6��1�E�$�����kK�a��%�'�@�a@�2��A��gָ�^x��'�@�Z�Bž�8Y���0?����� �I��%[q��*�ʇ�H٨��"O���ːf=����G&8J��"O���1��/�"�+�ɜ�>y6,��"O��c�P�Hy"Ƞ�*��8a:�"O��zҢ��u��5�
�R��!�:O@�=E�dI��WJ*�s�l	�d�0m
@��yb�ԴP-ܝ���NmY�A)���y2kT��D{g�?b����p��5�y��ܧ8���pg�Y���P`Eگ�y�⛈�2�౪؍PR�pp( �yr͐��d;D�.CR渒P`'�yr��1p�T�Ö��2@� m˗FD"�y����Yi<a��%3}C��:�y�'�M�1R�KĐ��L�R�yb$��������x2�wLG�yrnI���J�E��aNQ�&E��y�%�\ҔQQDS�^DI�a�Q��y�7l�U���T�aF���pM���y""��(���3��5H����@4�yrfA W�F�2���X�N܁�@��y��_�	���tFK�ebl�p!!F��y�ELhml0B�nͧF��؛PR�y�B�m.IZ�+��=�D�6(U�y���*�Z���+��4+��%i�4�yR.v�� l�&3@4���F��y�H6X4�i� *��Յ�y5L�b1��0�xk��Ǚ�yRD��~$b"$DC�l|�:��\��y��/	�܍�S,U&]��������y"OǜC�\8������P����yR ���K� �>3H �� �y"���2:6����C�#9��r&^�y�BV� j�E*@�[�6kvF���'5.t*��Y�$�-`F�+\��y��'��͑S���g���'`�L���(�'�H:��(GZ�1;���<�<��'�؈�h�� � 
$�A/EU���'E~�����1��`�*����'e�9Q�Α4z޸�VLO�$ê�'~p���ς
��ӕ�$n��	�'�dkAZ�8`�M)��V.�,�Z�'�L�qa-�t�j�r(S)��<��'���Ѥi_�$��`2�<I���#�'l��{�X
7#�-p���?�l2	�'Nlآbu�h9�Ƙ<���y�'r�}�2�L�æ��,�+,Wn���'{�y@e*�G'���ƥ[0$D���'#JM��,ޘR�,�8�dYs�8C�'�>Uq�0@��F�s�((8Q�m!�'W�ŉ�ڨ�@��Lϓ5z(P	�'�А���:!hF�Y�.��,��'@\ݨ���<t�B'� $�<X�'$�<�5&	�#j� ���s�<Qh�'O����]�x�8���N� �`���'G ��aG߃t�i��V� ˒���'�<�#��A�	}�Z��ي��tq�'H>\�UDN'%�(�v�]5xj����'��بp�J�s��`���\t��p[�'���O^H>,	a�Èw��	�'��#�X+�$)��-�0�X�	�'���ˢ��798`kL�%;�Q(�'���òˋ5E��!Z#�� 2����'h�����5Z�U�+���`��'IvA�cM�9~p �`)ڜ6|L���� �!:��@�7H �4��	h��"OdXB@��N�X`�0��J��݉!"O��J�-$n�¨S�៮h��@�"O�ݘpk�P����E���"O���c@�w���P'�S:f"��"O��8�+JF#���5�/h��z�"O�E���E[t�8B� ۱*��� �"O�0�Y�y��]	dbƧz��D�"Ot���%O�JDH��c,� "O<� ��T�h'Z���f�<U����"O,<x�c�# ��5pƜ�|FPd"O���$ 0�С���'xY��"O�a�eJ0L�`(Qe�ޢB`�V"ODЂ�A�y�F�©���l°"O�q�r	�'�05Cc�F�!��I�W"O��Z����� �h��JN��y"A�'z����U�f��}�����yB�+YbY���ϕe���Y��� �y2j_@�hf��g�Q�î�;�y���}�nK T�S�V���,��yҪ�������F@�P�`�!�y�Sl?������g|������'�yb`J����J����O�\���L� �yb(ˎ@�9�#@�B�b��E���yR(��9?ꈡ'��3;������y�Yd�%� Ђ;a�l��m7�yB˘�A��7KP,7I�T�����y���+9v�����+��0B0��y�&F�tb��	Th�VU(�B�O���y"L���I��o˳L;pࡃ��y�:]�q�CX>y�H�z b��y�kޚ��I7`K�x���h��A��yB��#��p�ړ�-�ge;i���`�M��0?ɵ��w��h���N�5@ihqC�r�<a��	o�t���-=B����j�[�<a�-�	�(Y����6����DKl�<�F��Q�B pT꟠��y�m�<�REW�P�@,�G �!#�N�0G&Md�<1D M.��R�[�o� ���c�<) ��S�U����0`�|�R��Z�<�E� F����\2��U�#�Q�<���){`��G/ݯ-�Z�Hu�<1��)G�8��uj��W��Mbd'�o�<a1C&oh�0�`��nE\�Z�fCe�<�eAB2+m"�����'Z��a�z�<A�n��,AȪ�'B�i;Z�֥U]�< ���/߀��g�E_
#%mLg�<i��	�L�f�A%��m��=��ȚH�<�Vd �1ؐ%Z	L�X"��D�<y�I�J�T!!J\�:�@]�GA�<�՗��\��8R��j��K�<�ը�Nutt�"�8� �q0� ^�<�@J�$�xe+��YoܠYe�c�<��f2s�x� �� �c���1�KZ�<y�eN#n>�C�Hv�\�Q�I]�<�R/Q-D>b���WQ�6|�f'w�<�3��#>���`T+~� ݀a$^s�<!D ۙ(&P�"�\.:��aYD��g�<�K�3Eǐ��dl�Z��Ѐ�j{�<iCP*dM�e	�ɝU"�}BC�j�<�g�Y��\*E��2��"�%T�D���ƲM�fT��`�LZ�YQ�2D�����Q�{Ĉ�Ivx��7�.D�<����eْ�����|�\"�f/D�� �t{���4lxw�(�,� Q"O~2�O�@N8��O3T{�D��"O�aY&cݮς�;���)hQ(�"O
HU`�kî�� -ú,D2H�C"O��BW�@�qR �1���9@�5є"O���B/�6�
�)�yF<��"Op0�5�F3E�R�K�ОB��ɰP"Ov`
S�S���Iʗ'�?ky��"O� rc��"�6,�����f���"O�4+��B�Sy&�"F ��]�����"O�`!�aû*B 9�O;k���2�"O��ńG�*7�{R�N�n�(�B"O�\�F��8!ƍ�A�� (`���"O�$���J`��i$B9J"O eG�<w:d��O��`���"O��R�K���eX��J?��ܒ�"O:Lũ^�M�=�F����"OP�����Xul���ڛ@�x�5"O$511��\�tU�2E�O
 A�"Ob1�!7D�Ȱ"���)#"O��8��X�X<"��D��-�F�W"O�!�3�F]E!���1v��5*2"O�9"!�O)���A`��uҜ��"O8A�-M�k�1���k96�"O�j�1S�x�NG�/p��"O��I��H5���с���)��'��P�G�a�S�O�P̛�O��vo���1dK�`Z~��a"OX�b lA �����cV-2�Ĳ��O���>�ny�	�*�f	�d0%h���㇃&�l�E}�IJT�	=|>d�I(�`YcT	"�~Q�w�N�6`��ЁL "E1!�TD<`!��)"]����dR��� �Ԃ��:�X[҂VA62�4ZR1������Ǜ2AK��G\��́]I!���m�(�"��x����~+�,���ۀQ.��ߴy���? �BO�z����O�@�&94�v��&坴2���"��$�O���EV�_#�� ȏ�F�dp�dF�
dÎ��1'!a��y��FMa� ���vz��'�D�@k� �`�5f��Z�l<��P�E����w`��M�!���z9�QH^4U� !��Y:=�����'�DŐ��\`��C�ɵo����`�-	��S �7H��jk��d`�)��CE�K�u�Af�+K�(�`Y|��<�
�p��K16�@�Ѭ͉ �3�"O�|K�K.r�dm� �҉, �T���50��j�W&�2��2"�%X��4�K�p�jM���S( ��x�A 9?�=�V�M0�^���I�F�ੑ��\	5��m#�B��������>zF��p�](©��J$`��c���uY��	�lj$����:A��!�b�;f7�c���.Y~���Q��)�]��
Z����ˁ��`�QC*�o�(�v	��A�"݋f�֟4����I�D�W��.d�4"�aP�~�d|�0dN{;@�B��A�@��M��E�l�'կe������+��� �n��"E��^Dt	(qDGw�'��@铨��l���,����"����P�v�۟,�|�3���C
`ם�"��Fg�-�T��Z�h��&<s����w`�Eu�l"UEa�����yqO���ɡ�U�T:�ɐ�K�oX�Ѷ(,b�~a�����q���Зf��i�4�z������ɱe����g��*C	4��AD���T�D�QlC�&ds�^���7m�
=�uP$��mΆ��@ҖW�I�Pf΅��(��耩k,a��G Za{�Kp��(�"ѤyXǏL�2���Q�6�t�x�{����FO9\�X�Ѧ��@�A������;`�F�H2���:C��)g��Z��F|2\
C�D�TK� �uC�eO P`���	M��" �sU�<B��ʟ��\w��{�ܔ8�X�y��>q �ݘx0!�F��2�đ���<�W��#l���;��h ��6%� 4
7F�=qeL�C@':VEpf Ԓ��6�L�|��g�+
�
�J��'>F�;[Ԗ�ȅn�5w���խI�D
i�$����:4P�K���<��B��eKB�xe"��$`�`�`�nJ�TB$#��_H<�p�X*J�a;�l�8m�qʒ��b�_�$��S��p�gLU	$��.eͻ|��:Bn�!n^�˦.	�%�l���%N��G��Y�`A�� ONj�n�	^��t��k�.n�h�'�6�� C�b�e�&9���h,H����R&�ȸ��I	Y�L�C䗛R�6er&
�%�μ�ߔ=�61���g�!��U
|m�%�p���DkSD��Ola
�H�)$� Њ2�3� � �%�*X���#�! ��͓�"O���d�D�]���#���35��X��Z?J�B����I9��d9�g?ٗ� G<�z�{��('O�U�<q�]�N�Liq�F�K��	u/���?����AdX���[R�*�p��j"&h�㤝#�� 7�Z�&:a|b@�8(Ҹ!�Q�M��q��+�~���ʇ�	'.b���q�ѧM���Lek��ضC�Y�����H��(O��9�,go����ޑ٘O�j�!⟝j?��q�dI�X,�2	�'9��s�B@>=�Ҩ���n��0z��( ��KM�xӧ���aG�b�F$b���E��q�A	"D� !⊂!����)G�"D��"}2����A�鉉h�� �uh��h&����B�|�C�$����O�<,��AJ0G7�C�I�L:`0�!עd�����2c��C䉔W#����a��@�c�Q�C�ɸF�>)��̴X��\KqA�8]�C�ɞ4�������M��Xx�IP�2��B�I t�<�9#���P9���4%�9u�C�ɦpo�D�V(�&�����I1:�B�I0v9�i�V�?7��4���	�mO�B�	\u�%�%��>Mv����>L�C�	������h10L���ǂc�C�	�p��؈��	�ӃEPۤC�	T,�]�Q&$W��%���Q��C䉱Rm�Qb`�
1���2��+.�C�	�*4c�Y6�����!�>*�B�I��\��݊1��̘'��_޲B�Io+|1�a��b�̬P�c� -ԂB�	%��Ш&OBF{�D:�a�I�PC�	�jP�#V�X��$�ӏXwKtB䉅.����n�#��qP��*�B�I/i�u8!�]Tȸ@�cۮ0V�C�	 v��`s��<"+�]�sFU-w�C�ɴ���S��4�pm�Ӭ	dC�	 ��ʀ�׸G�^�b3.N�OA�C�I9ĆT��#�R����}n�C�	�n�(��Uj5�\Ej��W�g� B䉀<7�zU&W�GO���K�Q["B�	�<!>��#��84�eP�d�4B�I0�dE,�!l�t�i��7��B䉳)S&��D�G ~��0*�>)�B�I?g�:������5Bqx�g_�ٲB�I�#�rhkq/&n��JBn�'m�\C�ɑ�B�a�X8M����ca��"�(C�	i��	82c�K����F�+�C䉜��u�Q�	�b ���䇓��C�	�|OZ[!%�=�$�ۦL��}��C��6��	��.�;*�w�0>N�C�	!VY�����GG>���M7(��B䉊<>6�@��O���m�� �:2�$B�,j�j�R��F�D�hj䌷?\��D�.6j� (�OB�N4� dE�aW!�d�G��颖&ģ��[��]�!�]/DS��ȖLL��Fс`ˡHw!�D�5,7�QVL����@����!�֐y�PH`C�H�`�\�A��k�!�e+�<*�p��L*5��@�!���8`-��/F��쵙�#1!�$Y�m/�h�W�'�n� �Q��!��� CU�d0vQ�)��A7M�j�!򤑻h��5� �;+?V	��@;y�!�Ԏ.�@�ŋD�f�J��
j!�d״l8!��*���"q�Nz!�$��tB�y'@� �Y�~!�� �x�@4it$\Z���C��P��"O�uce�T;iN�9s�eյ ��'"O��82#�	K�~t���P�)�"Ot���ŭ���c���L�
�"O���aB�W�	aw5�]*2"O�u1���I�d��4 �7�ڌZ"O�l�fOG� Y�1��A�
?Ѳ��p"O�d��j�;n�)s)�(q��K�"O@�#�W�Q����^>�b=;`"O���tę'ir�es�:0�>-��"O
��ѫ�&s��8�G�[�´S"O.��̛$c(u�"E+3�`5`�"Oް�%��E��J��P.�7"Oܤ"7@.2�"9 ��/C��7"O�L�wΜ:�ٹ�d@.g0���5"O�D ��S�[g���wC�%A)l�; "O�T�&MX��Q7�J�EL��"O����$�1m�+*$&1�\QG�~�<�bK�+��P�5eU=?�1��t�<1$"U��zs���J`��PC�k�<Q�'�	3zB� "��1'B][��3D�� �O��������J=�G0D���7h�$j����(�O�<5���/D�X��`3./�	��&I�/�)�r@ D����U�me����X�frrx+a�>D�4�g�ڿptdI1Mݩ"n���+?D�t[U�&w88�P�[�R�r��/D���wB�+W=*��H̽7Ur��9D�L��ގt�ŉ�
�&�`���1D�@��K�j�@����?ht���("D��9��F�1�p��&�=�|��n.D��X��`b>dI����b=����(D���&�8IF��g	�t��ru +D�8��"��b�"���-���1�)D�@1e�h�����M�8��F�3D�l�&�U~�b-k����dճ��.D�lC�IE��xT��![bO�)SA�(D�<�!)� =|DH!�d�!O�ƅ�bb=D�D�S��&Hb�9jқ{�B$[��:D�jW͞�H�T��`�R�d���t%2D��𒁒#W16����kT��E�4D��$`��e�#ច3�$�À$D�����m��A�I�m�� �"D��[5�� =/��c��ض[/���I%D� SM�C���PQD�6'�p�r-D��K$I�j[��.1�&�(C��
4C!����d ��e��~j��
�Iܫ)C!�ٻNO�ԩUoځE�X��t)!���9­�V#�(��9�m��7!���>O (��ц]�Bz�C��׏=`!�
,���p���bǄ���I&@r!���w�P�o�q�2�1�@�#_!���6\��+�3I��@���&J!�$�f�X�P�`���S�hJ!�đ2,`J����BM�ZXB�g�!T!��
��H-Q"��bؔ�БE�*4.!�J�`��$��l�3�N�)���Y!򄁽o�&�+�H�H���@��#c�!򄒳4S�$����q�*l�UfR$ j!��fu:E�D*`���f#��E�!���Y�%L�\�D;�b��_�!��1a�F�R� Q���J�O�A�!�A�lr���4`TBw�*�gM`!�DM(�4��ūN	h�3\!�� ����G)?B5�F���+��#"O �cgV��м�p��j��\��"O��@G�@�@A�o]M��r"Oƴ��Ũ]�"Xh���<-'�yav"O�qA�W	F�0:%��	Q&ò"O�� �Ŗ1h��iku/������"Ox�� �_� p����� E���F"O"Q��i1��<��J(c�&d0�"O�E�W��8��/+�8ˆ"Op��S�E��:'�pJq
F"O��`�aA"F�����jZ Y}D��"O��0Ğ}�� b0�FO����"O%��L�6X�ʩx�ㄇ2��,	C"O��:'�?�h��њq���`�"ORq�QF������Sȃ�N�"�w"O��1�mΑP��)P�� >h���"O��s� �`�����E��"O8L���;%�b�Y�%ހ���"O�������$I��E��}�2��"O�, p'
]��R��	1�ڭ�"O��*�,C��$#m�025"Ot�vf�����,�)�$-�`"O�|���+i<��jły�"@G"Oh��#��<�%[B(�1:��}��"O���v)ȓ )lQ �gB4,xz!6"O�@�`@ΑD%�6Ǘ+�x��"OR�[���h�p)�E�90�0�{D"O��$&�o3&@  � =L��"Ov�I���W��E)�OKN��9P"Op�����:2B��"�]�;���u"OlZu�^�P�}��X/*I�"O4pA3���(Ы��d�=�U"O����D��r�n$H��A ���i"O�����Q�`��S��t��"O��c%S�p@�3�	Z�vy��"O�m�-�m��Qg��;	q@"OT�P��7��U�2��k�̐�$"O�v�ۑ]d���gԸ\4��U"O��!�أ!�T0�E��]����"OP�䙈uP��# �� ;=�U�w"O�5Q荙�^��Ղ^9Z;��Ң"O~�4 �,,�L�I��2"Oxiu��=~3|�cΞ0;� �"O��)��^
������ >"e.��"OL piУ��<` �O
"B����"O��+7+�F�<���͒�pNBE��"O����x��,��J�1)��0�"O&�Aa�)�����J̻L�h1"O�M�w��:X`��d��<6|��"O�s҄�:5 �B�.4�䱘�"O"M���#��yc��O�f( "O�$s��@>T�0Z�c4[���Bw"O��Y�`�,-8�`b�-h�^}�"O8��8=��ᢌ�_[rMB%"O�P��`��*'�%� �ǉOM&��"O���&����EۚV:Q��"O��##F�U����aM�;�rq@�"Ot(���sL���<��-��"O�}r�����`���&��%YU"ON�[��cD$#Vb��Da0h��"O���5�ʁ$�)��B��C�����"O���RI�hXN1!A�ҫ	�
3"O E��E�S������g'�,�P"O��(6���7�ʔ���R� `���"O� ���Bس1݆���Օt�,���"Or��E��5��%��Ż�"O������(A�gjI�O�P��"O>�"����cƊ2$4��"O �J�V�wU�H�.� �Ț�"OZ4���R&��f��O�#�"O(�� ��A*B��� p8t�r"ON�ё�0T�,�R�Y�d����"O"Aᢍ��U�V1 wI�n��G"Oz�����H4��!�h��Vi~!�"O�0�@WK���S��(ED7"O~���4rw�-âM��H@j�b"O�@8�	��H��͘�/��Ka"O�i��E� �e�wPD x�"Oрb��/����J&j`SA"O��'��(Y��X �G�T\���V"O.�0�Q7��h�	�15���"O��b�.�L@8�C#>&���"OfԠ�*��IJ,� fE&0b�yg"O<tk3��>4��"#	h԰ې"O�P�$���-�@jf-�}>�s"O�4�+��R����A-^;���"O�41��s���ɀ���_&8P�F"O41��wG�p�c
`����"O,��Ƥ�Ada9ǣ�) 
th�S"O���c�Ae \("!ĺ\��"O�q�ă�4�ԢU���b�,%2�"O4���h`�MK�l�:��A.�yr���i8�o�[��A����y��3rq�S�	��M�`!T�_��y�iT�{�x���i��K4.C��y�,�2w��87TX��r��ȶ�y��qx�cVp�"c
��y�gS/wі�Hi�Kc֙3vG�yB�RD<t(��ډi���⩌7�yB�:5<�<ѷΌ�{r|ݢ/ϱ�y�,�v!�p�AE�ioP���$�y�����߉\���s�+�jfh��`����J��f   �?ɸy�ȓ{�~���l���Z��剓!���ȓ~Z���F�)DԶq{�_	[��ȓ-�Ό��ҴEt5�'@W�Y�ȓk*�8a&B�3�����D�{V4��jz��giַͶ�p�An�A�ȓW?^�:֦T)w�����6B{N\�ȓ2�t�@�Ț6|؂2��j%zL�ȓC�H)��k[/��K)8�)�� W��@�G�z��J�
� mȅ��*���tb
$[���
�.e�a�ȓEH��k4� �\:uO֍H��i�ȓl�d�Rj )zp�2h2[�Q�ȓ�.���l� xN$Uy��� �V0�ȓ?�A fb�	8���b�@_F̇ȓ�J���	lB��3c^�}r	��
�H����Rt���FG5(A�����E����%VR�s�E1���ȓ��q�S�II�ʁ��i�)=����{�hs��P&V`�˃�B�PX�U�ȓ���Tk�:b���Q�A�x��ȓ P���"���F�1۶��`F����IR�|Y�����r㩁�x�bІȓ \�(���Ӡ�~"u(�%l��m�ȓ+IT\J�#Ȧ|�9�aS�<V���ȓ3����j�8&���!bm��cm�P��S�? D�&h�&���� �Y/T�w"O�0���D�@1�4`�#7*i��"O䀲jG���@bo�2��s"OL��Ba�,{:ܡ5Ė�~>�I�s"O�L񦣛�^���9�39>��W"O����3(D,$ Kӧ%z��v"O���Y�VP5�ʬY��Z`"O�]�rn�Iۀ�����$
��f"O���1�ݢ"S���,N(t+d͊�"O�ų ��)��T�����`*x�4"O�CIM��V4��#*Dv9��"O��Ibo�)X�tZ#�·a>���"ODP��LH�h� L#�ɋ�S�Z��"O tإ
�
m����Ǉ2u$;�"O脐��=LԹ�ɢ'���B�"O������,Ȧ��
�*g���K�"O��	'i&mVu�D	���5ӆ"ODXJ�+����;�fЦG�4 �"Ohp����Ӡ��e��o�\��"O�u�3�\�*أ���z]��
&"OqQ �,. u���I�P)
"O���Ԩ�6}>9�sϑM��-�"O��(��Ru~��CD�<�I�"O���R��l?��+#�/9�jܘ!"O�� b� v�,�©��eٌ�@g"OfE��'%���au��� Ƙx:�"O4����p�
&]�q@ ��"O��S4oZ*=�|U�f�-RƌK�"OHd�g�]DN�
B<7\Q�"Ob$!6c��^�@4��Z� `���"O��R4B��Q&��֤	�}�t"O$p`#hE�R����mH��6+ "Of��P�&| �O�62x�Z�"O ��^_���`��<Z�L��"O,�ڥ�W<�2���%U��3"O���s���>��#lZ�i�"O���ӤL	��+P��-V����"O�sP-ԊG	։q����O�<P(�"O0�+�N�lF�(���1v�b-)�"O qr��/?����Eй�b`�"O���20gK����R&mn�I1�/��<F�''
8��D�2H1��@BDY<��3�'X�8�@�U��ē!H%,����'��-� m7Ux�+!	� <D��'p0�*
�c�*Q��=�jI>��ν��<�}��m\>@}�rG���]�~hqr��Gyb�]�v�t)�y��)]�d���B+�:���μf��ɷ>l����.�)�,vZ�"֋ .R��AeN�X2��r�Ũb�
�*��T��)��� ��)p�m�qv#C�lRl��q�Ȕ8���6Q�<���v*���Z�"�0���IE������#<ب�"b+���`YdoX<[�<ʓ�Oc~�������mV2R��m�&�Ǹa�R$���Ͻm�d!+����0|b�I
�k�Me�N�uv��:ZR|��4%5����q��;{H-"����~�K|�uJY�P��Ͳn4}�X�֎˕Z���U,����S��M�;j6�Pt	^�1َ�I��٩t=�$i�F3�	�0|2�K�MlY�׎]{f�J�B�Q��P�X�J|j%N��l3�Da�м��D�P��	2ê��?�~��f�,1�U(���:^�2H��TV�<9��=A7��hS����H�{P�BR�<��,ܭl���3%�}�!�Wn�r�<�.ՓO|���&B[n<HU��n�<�r`��	u�0+ �Z�~�v��C��l�<��Q/b��
3鄷#z��3���e�'~ay�*�Hx<��MՋeB������y�F7&,� ��'����FL5�y
� ����$�T=k�iV�y��Mb�"O��1C��7( ���0(���"O	��"�9:��]��m�6$�	�@"ON�)�'6���(�i�'n��0�v"Öq��^z�l�	H�<@����d"ONm���ߓ{��q,J�|d�Q�"O�� �,�#`FH��̗vY�b�"O���S�ƞDj~��ɍ-s<���"O���c���	������y0�Ub"O�TI��U)1XP��9x�@1"Oȸz�Y(�2��)��5Be"O�]b.mjn0ڳmL�0K�H�"ON�
ce�@z2�C��,T/ܬ2�"O� P�'G�8�4"xJ,{"O2y��s/��Jo��&���'"O �q��N>P��MC�" ����"O�Pk��%���P��e��H7"OL�0�(]��9R����E��"O �҉ZU�����
�%
�}��"O
��AEߤ>����
-M�|"OD@��gӼp�¬��J4z��bF"O,��6 ��t|�أ���Hx9K""OB�@��}�^Q8j4��B"O�Lk2���\�s0g],+`P�{�"OV8�քS� ��P��8PL�(�"O�UYUb��U~Ri��'���Q�"O�)P�Z
7�P�M:l͞�8�"ON%q@�"/��J5�>�A)�"O����hM�C��XX����_Fl
�"O�1C�]�S	b�c��B#��K$"O<܉6�B cr@A CdB%�
m�e"O��؂Kώ�6l�K���|5"O�q����_p�(�2a_����36"O:0�5䉻i;>�ɤ"')���q�"OpK���8�D����GQ��yТ"OȐJU B��I`#��|T�"OtL�� ߏt9Z9I�O�D}A�"OL�ySG�&8���q��|�䲄"O�<X$N��]�t�igʀ�{�L���"O�$Y �ØR#`I ʙ�;~x])�"O�5���-�� !B�%>�I��"O��� >:���Q�m�|�uzF"O"�x3,c�P3ƥT��;f"O([�DU�@NA��g��\����"OP�C���<ʄ���L>@m�Ts!"O�qY"�ߕ#"V��ܼP\��`"O����+ S�TpWʝ9.바��"OhE �+ѦZW��(P|�*h�R"O��eRP�=��7�hI!�"O cC��%#�B���eڼ5�����"O,�(�=G��� ���L�(@H�"O�$�2d�h�4dw�r{̅:�"O�x��O�t]�
��* ��y��_=�89QʔS�ڐ� ��yB�K<F ��ʧ*�2OKZ��rͲ�y�m2Yih#)� I��9b`ݶ�y�J<��0�:qb��a�@��y	��k�0��a��,`���Ja���y2F~�F�p���S��AY`�վ�yr�L��� d��a1��q�ӽ�yˢ&u�����C/`�P$� $E��yR�Tbj�!��T0ڄ��,�$�yҭ�P�Y��c�%QP���s�O��y���=8��;��	�8BY0�}�<� <���׊q������JFp4�c"O�,���ŷs�ވ�����3.�5ap*O���e�9Ea�
��\`�'"�����&M���ˌE�@�C�'� ��!Q<r�� Hg��9.m+
�'�p�����7�^�&�?*ݖ`Y�'��=����-ub�	�#�z�����'m�Y��A�k���E��xO-��'8�$qJ���t�vl�4_bΩY�'�J�0�Ł��aBG�W��m`�'dp��FK��Q���H�>�E�'  4����>��Y��(:,\���'�z)1�cȧ��*UJޡ!/Li��'�E�'�§j���HD�^�J2Ʃ��'�fٹS	��,�æ�xa��{�'I�m�u��6����E�o�p+�'\X�7ɇ�ow�9*���`��AS�'�h�K��4���F�A_�d���'rh��.��x���LC%V}8��'�8� �Kګ��!P��G�M����'�REHq �/4P��gX�L��L
�'rn�`oV�ܳ@��H��
�'���b7�ٹ#U�g L�9�|��	�'6���KBt|}p��2��	�
�'�8m�sKB(���4�69N�z�'����1�E�MRp���3�(9�'��d�V��M���E;�}�	�'�N}��
�l^�Y�GL+ Q�t��'�.y��G61u���	�1u��1�'�`P!�R�l�L� �o��k����'i�h��ɍ,�~3�/ݖa�@��'�ny�E�H5*�@fk�l�����'�B�y���5b�K6�ːz���;	�'K��q�jNx����]G��q��'O>!B�l
�M����"��<��`2�'W|���/����5�ʑ4	�(�
�'h<|q&¥@�� Vk�#�f��'�J4��Ǉ*_��3���*`��'tlQ U��-��Lha�1�N�2�'ld�I `ԫ\��S�iY�_�����'� m#d�݊�b��g�5H�p���'W�|��$Ō`]n���I���'S���ǧ ��cM:q� :�'ʦ�qn�3Tea@��
0��)"�'�n=+uL�;#/��bJ�$ݺ��
�'����qe
Or�0���L���ȓS�<��`D�/t�1t��C�Z��ȓK����&\ ���Q�@e�x��X\I:+��s���AQC�=����K�>���C^~x�ۂ蜝}Kꠇ�[C*Sh�� ��X� �K��x�ȓ9O�IRp�2qV�%{�A� 40��L(Jxg��j~lx;eNb;�y��y�0�t�%�P�kE�F�|���ȓm;D���>8�r5�1�O15Be�ȓ��<��bD�o�^�SP�4~.�Y��eH����X �Qs3�-� ��M�r�-�I���� �*�z��$���a�郯9����XBT�A��5�n�EE�'*XD�@'�3������f0I��2/"Y��/Gmp���'G�<Hb�͘^^3#��1I$ʕ�����2�X��X��$��1E��I�ȓS�ư+2a�� ��oC���S�? u�A�ħ+� KO�_j�Z"O�IYB�ߢl<��Dt��tY�"O8�	3�¹h��z�.�.9��]b3"Oz �6A�H]�b�,�ɒ�"O�ظ�n��,ش��Eg��V^�"O����`�3�p�2�(�Vيc"O2H�S`�a��f�LP��e"O�	���e
�� �+�%b��d(!�$��&�Dd���~�:��T�U�R%!�.Ex���֎�'�,���2!�
.u (�#�>R��`P��I2ko!�ބW��\�AѠ��}0��֎!��D�~	,4�������r����P�!�ߓ�n����$u�3��ي?�!�w��Mp����>�* ��� (�!�D�	\w��@f'�=�X�� �!���,�t�B�'�ܽv
�h�!��E:�ج[V�g�M�T�R4�!��T!8��m�r��m��U�7�E�g�!�׉�DI�]�}��(6��Q�!�$�Ixy���t�Z�j�1F�!�%\�f�a�Q�y׊z��L5t�!�DU�0�t�QT��7<]����A$�!�D�H����Лf2̲Sל"�!�d��^�4�6EIv0�7ki*!�$1I"�A�F8F�Ī"-��8!�d��&tv��WgM/E��Ȧ�Py�ءa?�)�M��'&y*d�ڮ�yrf�
���DF�l8�֒�y�B[9viM����H�r��:�y���r�ة8B��6QE�k�E�y������Іޡ2� ��� �yR(�)o�UH���h��@���y�i�-@�(
�*	�j���3C�y�����҃��2��pi ��,�y��K6y�(!t1>�'	���y"V�8|	�S�� �@�뀍�y�<8;�q�Dqm;&��d�!�ߜR�~ٲ���%M�*�'@'�!��5G3^E�G�%�n  �hB�	�!�$֘�ȡ��d��B��mI�Y�!�dJ�!.4��+�?��(;u��SX!���Q��
0��+�����;F!�D�yw�E��̊�yl��H��!�P3slZ��«V -s�e�JJ;S�!�$�:��CS�N�ȤٳC��>�!��:wݎ�*����_HU���sx!򄄯{�����^'BR��%��Qj!�<L�
�+�n)G�(�k��p�!�d�*0GB�{��O�cj�P���6QO!�\�=�6d�C�r�"Q��aV8R�!���X�. �e���X�r�A�&�5!�$�O;^�s�m 5S���9���!�D��2HB��A�_M��; n32!��˰EK�T��ϫ.� �I�ķ	!򄊵I�D�C,�	��b!����!�DL�6���W#��*`��F�U�!�^&V��*�
��]�U` �.L�!�ҏf�fDcK�lYfx�n F!�DA#��%�V@��x��V!��X)
�jIJ'g��?0d�F+��!�䎙�]�CkW�	&h������!�J�+��h��_v��*��E�XV!�DB� ���^)2
_(��"O� �Q�N�r�% C>��`@�"O�t�Ώ{'R]�ph�FHXe��"O�t�$���u���Y���}�"O���A��	g~a�Qχ�"��@
�"O�}`��g�mIԤ�.b�e9�"O�qC#�5�]�2ꆾ�M��8D�|2�
   ��   �  ?  �  r  �)  �4  @  �J  V  �a  �l  �w  ��  0�  a�    �  U�  ��  �  *�  ��  ��  D�  ��  �  ��  �  c�  ��  ��  =�  � � ; - C% �, 4  > F �L �R Y [  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�Tn�9g*�Qq4��d@9�L��|�X|{��>?Q����'N���ĳe�����(P����m$es�KB���	
E���m�f~�7�R1�[�iR�5j�P�1a�	/^�\y�h�Z1O��D�<Q��IL ;�S��NA��@ס�$G���lړ��c�����Ӽ���:�⡛�.A�mS~��b���?A��yU�b>A���֦��QDp���I��>*��a`F�\����y��Od����4�F���lg�C� �~e��]�h:�ı<�M>��iR� q�y�;s�[�8>'�M[���=X�O0ʓ�?���y�Z�$�A��;!2���P��HQ��,?!�r�h���.�[�'r�j���?�a��(��A^-s��}`#���D�<i�S��y"�l�$���'��M�v,�@d́�y�Kdӈ�;������n��|2t�>s=���K��	xp��<���?� R	ܴ���q>�1��Ct`���OZ�%@� YV�;�9@%&���<�'�?)��?���?�s��'���I"*��#dP�����ď�}�qy��'C�p�9���A D�+�v�0�S���<a������O��{�ڢR��Y���Jbe@�@#I�9b�U�8��� h����D��Ay2��Sr�� �-�hI����'��'��O�	&�MQh�?�?ٴ/�#��!��"+�`�O=�?q���'J�۟���䟐K��^?��L��&�5����1m[9.Z�o�Y~Bǹm�P���p�'�#Pc�Rr|0��S%�!�s��<���?)���?9���?)��T���p�'�J.%�t|QQbʷ��A�����I�M�$@Pv���'h�'>�r#��W`}��$YT���|�'9�O�a`ӵi�I�O��ĩ�%�N0�7-�3O���Ecj���8���<!���?���?���۷,���Y��K:^sv�Y��?q���$��]��ӟ8����O�Q�u�� z�eD5!恙�O�˓�?�����S��#�*/�f��R�ֈny��r��D� <���B�J�*nn���O�i��?A/�DG�i���HW�:�6��1��)DH���OL�D�O4��ɰ<i��i;�5��iڂg�&X
�A�P���!�܇���ݟ��?�(O���|�&9P��B��$<Bꂣ��Dz T�ش��D�^�8l��'"���Z;�U�1��m��"��"*�0����O����O4�D�O����|��F�$$bx��c���a(Ǐ�d_�,Ęqv��'�ҟ���'��w<��EdO�T�(�sˋ��,�R��'��|�������6<O<B��#c�����8r�p�;O�=�1�?�?qW?���<�'�?�`�F�J��T�ǂ2Q�0����?���?I����ɦ��F�ʟ���ן��� D$ND��	�$Rz��))a.�K���$�O���!��]	V�@󡂛J�h��*I�x��	7�� �ӑ$��c>1�@�'������hWHĳ��Ռi��@� 	нP��x���,��ǟ<�Iz�O����e� 1Bbh�1��D���v���2 f�O
�D�O���]/,5�@���ue�$*�i��hb�I�������˒ܦ}�'�
x��� [�W��o���WC�� )��'�'�䓢���O����O��d�O.�$"IblSf�־\\��g#^r8�A˛F��6>o��'����'4��sq�E&�@��D�%I�| U�P�	���&�b>�ّ�Mq �b�I�V%l�����O��d���~yR�)M8��	���'O�ɴ�P���ջ*�5I�/��1���	ٟ4��ן �i>	�'h�7"yG��DN-s�Lѕ�ňM�X�K�������OV�`�'���'{B'	�E��AcH�6^��-��ʂ n��B�ia�	�*%�Ar����� �H��P�h��k�$/lT�(�8O��D�O����O��d�O�?=q�JfLq����"���b����������42_(y�'�?�����dV ��:"��YU��I��5�<Y����)ͬ6m.?Ifń JO�-P��$ԺA��6&x�Ԥ�OrP	H>�,O �d�O����Op�9�JԻ^�� ���-��0#�C�Or��<�ÿiZ@`a��'q��'K�S����2�_w��u2f�܉M�����O��d9��?MQ�U�v�7$�l�=	Pm��X�(�}I���|
A�O�@�J>颠�rT������-&����4����?����?q��?�|�*O��lڌ?i衡ՍG-6jQh�+~�ڳ�۟���ޟl�?�(O&�Đض�b&�B�N4�i⭚5�Lʓ}b�qܴ��D�)}�>���'$�:˓n���D&�&�~4Q�CL3$��%���d�O6��O��$�Op���|ڔD�X*L�#�^�,��,+�$VY���	��'�����'��w�B���ӣP�����>LD���3�'
��|��D��RQ�7OF��U���1�~�%!�P�X��a5O
��Ά��?Y��%��<�'�?�ǂ�'�:��Y�As��!�j+�?9���?Q���
�u�������	��P��
A�a��c��U}��ӡ�TD���$�O��D,�d��<a���T��1z������ɷcf���R�Ǧ��O~��%������z�6}��N�iq��Q��PF&����d�	�����_�Ob"��-vl�u㢨�2%��]��b;���Ӕx��d�OX���O�����!���`jH�9R%E0o��	ҟ��I؟�R��æ��'`��I�!��?�C"-�40�'��-5�HtZ nZ�H0�'��i>-�I�������P��2�%)�� �w�<�Q�D(@[L�'[R6��q'J��O��-��3p�>� D�ˆ^�t}���P�c($��'���'�ɧ�OZ�|�P�'͖Iڢ荸U��yt�'p�0y0RX��rG�	-�B�s��Hy2"�>j��J�%J�t<s��D10�'�'D�OZ�)�McFS�?�Ԅ��k�s�nJ�n:v%It,���?����'��Iߟ���䟔xQ�&'+&�l�p�j�Ȟlx���i��"{>8�p�O-q�B�.Cn�䨳"$���ِ�W?!�d�O����OD���O���;�S�������l%R#KO�c���ϟt��.�M+�	�|���?�M>�@��w��4�b�&:�x��C뙶���?���|��	��M��O���=D�J['K{=�n4z�^�Zc��O�u�N>y+O���O��D�O"@��U~Fx��#2���P��Of�$�<I��iR<@q�'��'�������D�9c��Y��F]�Hc���$�O�%��?E��o��,�!�c�z����o�H����M5�1����KSʟ�V�|2�J�.��S�M�`&���a�n�b�'�B�'_��4Q��;ݴ9X�rR���;��עޯ%%���e� ���O���'������hx�Ä6M�Q�E@"p~�	�vlPl�m~���g4H|�S�_�I�X��qUBQ;aZ*�顥K�G���	[y��'.�'{��'x��?�@EĎW޵�P���xU�0��m�Ħ�p�����p��ܟ�%?�Iǟ杜=��`�JN�e�T x�L�2k����l�Ş����ش�y"NS.-�N�"� �a���M˵�y��T&"�d�Ɉ ��'����I
6>\aX5(�f���IG��8UTJ��I�����ٟЗ'267m	�a�����Of�DS1�Ե3C߯N��y(�(1� �4�'J��'��'�l�J$MB�2� ��AI�;�����Odp��µY\��	O>�i@5�?Yo�Oz  5�O3<+� "D�D�؅��Oh�$�OR���O�}���j�tP�>w�p�P2@��"�����]ћfl	H�I���?�;,\LH8�R� }��L�?��	ϓ�?!���?��@��M��Or$�cM��b!�A�3<�]Zb�Wd�I5' H��Ob��|
���?I���?��Z���BMڄX����g�S␸
(OWc���I�E�O���Of���D��0d��\3
��l�$^�];�ʓ�?a���DȖ^�8�"&	�0�r0I3���D�2���-*� z\=��'N��%�,�'^8p�&�"Y�����* 6\S��'I��'�R���W�p�ߴ ���Q:ೡ�V(Z_�Y��
�0q� i���?���S�P�	�<�	�Fr�ZL�1�,iX��˓P���1��ᦥ�'MBQs���?�Ӕ���w� �AW�~8�B��٘)���'��'/��'>��'K����W4;�P�!0��T7����Ox���O��n�b|�'��|�e��ژȂ�1�TAӰ�N]�',����Ԋҁ):����lY ��9Rh���OݰT�d�F@5Is�+��'��	'�̗����'�B�'6NLbU��0�� H�u�h�3�'b�^� �ڴc��
��?���M�m|���s(����CE<@�	Ky��'���|ʟdt�f��H\����u8���eaF�s��h�f��_��i>!ل�'��%��d�� F�MZr �o��\��o�����	���	˟b>�'�N7Mٮg�H�12�5uZ����GçW�@16��OL�D�O&���'&b�[<)�F��� 	f�M����'vR�'4�� #�i~�	�^4Hr�� T|�f�C�d�$Љa�C�	h����;O<ʓ�?	��?a��?i����)M:B�R|�d�Q<w|��!D�,��doZ�|��8�',2���O��4�.4I��ϟ5z�p�'G=^�����O��O1�r��c�
��(��;׌ ��B���V��	�s��0�'A�D'����d�'͠�Vh1��P1(�(� �Q��'���'��Z��ٴTJ�����?��|��h�g�Z�k�[�'Ӛ*�ؐ��W�������%��Q��ͮ��lZT'�/J�r���j8?ɴ�E,&�ViQā�2��,�X�ĕ��?1�L\�TKH�K�NJ�bUh��#c�	�?����?���?��)�OD�	��@<D0tP���`#���Oho�:H��'F�4�lP��e�����Y�E� �D僇2O&���OR��	�-s"6-*?Y�)�0[���IG�-é�.GԚX����(t��dxL>�/O�i�OT���O����OT�Td��X�Ҽq��E�'��a"��<��i����T�'��'l�O2�-j���K4D�{�����D������t��S�)��yL{�Ī�D��q��Z��������/O�
�� �~��|�_�S�i6G��)z�kY&y��|�������I�(�	ϟ�Ssy�Kxӈ���O:)�B	"'縥K��X,�P q��O��:��Xyb�'r�'7 )�߈;t"�@\�[�����J�K��旟��v��@@Q>��]7C�j(��̠	HT١w��;e����X��ӟH�I��x��n�'>�>aE.;OlQ��ş�Ql����?��k��nK���t�'\2�|��)1���(�Fl��Ѧ�E�S�'������D
�F��F���
)6��+�l@=g��5c�۟oظ-)0B
���sv�|"R����ߟ$��Ɵ�Z �^m��[��K:
+�h3h]�����ly�nj�R��R��Oh���O��'1����W_�ja��l�jJV��'��	՟���q�)�A��V�q�L���I{����$�#6{�P���4MD˟�XA�|�-��3����gJH�0�x��@�8`�"�'���' ��tV����4TĤEp�@�'�J�C�mb��}�����O���'X�@��Y	��p�nI��KH���z��=o�V~���`7�T�ӵ)��I�E"��iQ�	�so���cj��#$�IXy��'d��'{B�'q"U>�Z�(����Z��V7�\�C�A��Mce���?����?�M~���?ͻE.lD�c����rb�Z�Y��?QI>�|�0���M{�'n�	x�LG�s)X��ő �(�(�'�t�8W��A?�L>1)O�	�O@}�rΛ�#���EɈ1N�*a����O��$�O���<9�iY�V�P�ɼ[���%͕�5�Ѻ��-Jo���?�.O���.��*�4XhslC�p���C%쉋eĴ�
�<qe� ˂M�I~2EA�O�M��}��h���H�/v<��G	P�EA��?i���?���h���d�}J��iW?=� ;KӎlPP�d�æ��0���`���H�?ͻ�H�NTv|lՍE�G_j�ϓ�?A���?��`
 �MC�OTuP �����R�Q:lyKW��4>lBW��+l��'�i>��	؟�	ğ��I/p������
�`B�%�δ�'�f6�PC�d�D�O��$=�	�O,�Q#�9O`J�&�
�"��E�<�������O�24�oʛo'̡�fO��_
�)x"\ʦ���V�, ��#1��ƚI�byr����0��K�[ʾ)s�R�b�'���'d�O�剺�M#�KH)�?�B��Cd���ı#it�{3bC�<y���'�����I��0$�:K �]�����)37JQ,{�doZz~���8EY���䧂���Kn�e�B@��r��`��<���?����?����?A������ф���9�ǚ� C��'db�~�v��  �<a����a�$� (Li���ɹI��!0N>����?ͧ@���ش���7a��)E'�+spL�5��y� j���?�2''�d�<�'�?����?	��.W�Zl�	�8a���A�O��?�������e��@W��	ߟȔOC��	���mRlZ!��taȴ��O�ʓ�?����S�4'.�Ё��h́_��d ��/r2 ��,ʌd��4��O�I��?9`K0��ݡ؅JЅO;<P��[b��������O����O��I�<�v�i*��=1�:l@�F�):�J�peB%O$2�'���<1��hZ�A^��X��m�Ͳ,O�����b���exP�E�ҡ�,Oѻ��ك^��<��0�j5�G:O���?���?9��?������:5
�iV`UUˈ����g� `oZ?(���'���T�'��w�2�HT�#n�*Y��a9#n�[�'5�|�����[�&6O>8��H�9$�@|#3#]�&Ԃ�4OF�CP�7�~��|BS�l�I՟��� ��j3�Ta�lF��ba�ϟp�	ş��	Jy��|�$��OX���O�8��@�*��x��D	�6.�h � ��yyr�'��O�X�54ޅ���SY��� V���`�� ��-�Q��N����ܟ�i�iR?[q�$jņ�
N�Lx5��ɟ0�	��<��ПE��'�n�r���>)��� �-"lh�c�']\7-J�f���O>�$+�i��2�����c�̜]β	r�+m����˟��ɒ&� o�o~�g�l�^��g�? rPc�6L�Ў]�z���2@F ���<�'�?��?���?��eP�5L��ʶ㔺 ��ڶć����¦U;P�T�����ٟH'?牼3vЬ���������nӐ~�Y�'�B�'Gɧ�O�0�"nؤ-h�;C"ی@��Gچe�O�	�2���?��%���< F԰6��8���L����8�?��?���?�'��� ��!�e���TH��� �&���o�*��9��ş��IZ������O\���O��R�O�cb����5k�@=�FNR#E�6m-?�,�(�������'��s"@N&�`@#V�Z���1��<i���?!���?���?��D��R���{%bB-�lm�%M��')��p����F2�$���OܓOt�O_�Sf��C)�q��D�R�$�OJ�T,���ٴ��d���Q�����z%���F;IC�U�CF��?a��>�ĸ<����?����?�u�s<zs�Ѭ"�2D��]��?�����d��}r������	ҟx�O:(��V�O���GM�sq��O�˓�?���S�dJ�pr�P�O#pȔ�#ĝ	^�$�;����JX��S�/��(]r�I=��� ��!d��f��rv�����4�I�|�)�Sly"�g�H�8�@zjh�B�˂9����5W ���Of�d:��Uy��'z�%��K�g��u(�U�aС�'���=L���������Y(nq�,DPJG�m	W� �4�v=O�˓�?Q���?���?����	��vc�h�&Df&0)�EX6Ξ8lZ�i���I�<�	_��柘�i�	�2o�*]��Z�A?�H�1$���(�	o�)�=t�Em�<	c�;��$���s�\��F��<��U*KP�dȥ����D�Ob���VtC�Ǡ�r\��������O��$�O^�5���Ej��'z"T�x#���6a,R�2����
<W��O�˓�?�����$0��0�V=[�4X
�A�X~0��'�zѰ���%��f�H��~�' `4h�H��9TkQ�#x|2!�'b��'���'2�>��+v��9C��"zNX(V�H�,�֌�	?�Mp+���?����?ɏ�w��A���>pd�Q Ѫ�G�Vm[�'�B�'�d�@˛�����Q?U�����^�̸:��̊-��9q��M���&�,���d�'l2�'�b�'bDY�s��:S��	��>1�y�bR����4HfN�i��?Y��䧒?���$NaH|[�Z�fd����nҐ��d�OZ��#��)l�����DÞE#<��O��U�܀7��G��<w�D�A�':�l$�P�'lF9��Y\���@g�җj�r�zt�'OB�'2���$W��8ݴy}�9z��rxIwm\U�Ȅ��/v<zI@���?q�R^�d�	۟ �Ʉ?j:��T�g��!�Q�W�e.�������'��������?Q�}��;�@h�	�CL�	#)�1`�D��?����?����?����O��}Q�`YM����g�(W�l'�'	�'F7�ܙ#��˓�?aJ>�vG'V�@�����R�"�ݳ���?���|�4O��M��O��BӉ��h[��KQn\�y���U� .-(ܠ���ēO ��|z���?���|h��
T� �V4"��B҈�`��?�+Of�o� L6Y�	ݟ���`��,��hg���.�z���@4��D�<����?�L>�O��-I
>WAfؑRjF7���X�t��r%`�-��i>ݢ�'v��&�H2��%$=4�q�m�:�rL '������ȟ��Iɟb>�'�,7��|����X�E@��pCL
��	��Ρ<)���'���ş��`�P�r���q�A�<T�b�
�����,�I�1B��nN~Zw�ԍa��O�b�'��5�ׁ��	��#IP�
^69��'��䟬�I蟴��ҟ��IC��!�-��˗�$�n�/E3��A��i��§�'���'�O�"��y'�T�Z-�aF��xTy`cK�?"��'nɧ�O�Tp1�iv��)��\�P	�>!|��f��8e�D��z���h�j�O~��|��C�l��-��,��B�2-���B��?����?�+O:�oZ�
����	ݟ���9�&X�g��4k=x)s �I t��A�?)/O��d�O��OIj�MM�D�~��V�˵:�dsv���:e��f<��l�C�'�~����8�E)݌W *Pa���:K���������Iџp����8F���'+�ʆK�)$*D�N�>��r�'��6��G0����O���=�i�I��Ď*t(���� #V4@P��k�(�I��,��1��Tn�_~�Ȉ���;����V�U�2\�O�~�I��|_����T�����I�%k�~r,��HB�:��Q��fPKy��qӪu�f��OT���O����4A���M$#B(\�)V�<���?QM>�|Rf��4/�����8�:P� �)*�B��0*I~BA�1SD(���0��'@剫A[`� ��͍)( �H�j�;	�4��Iϟ���ݟ��i>��'A�7��~T�D�;r�6�X��Y�v!l�I��[���D�O��X�'v���y7C�n�>�*T�*���y��2N8K�i���86UȜ�V�O�
�'?���L�<� �J���0�Q��-~��͟��	ǟ��I��D��@��y��bP����rn
�aN����?��3כ6�ȎW��Iݟ�%��������\���NB	"h(1e�I�Iџ��i>�j!�ڦm�' l�j
� �ta�F�4�;r�֊R�N��H��?1�l3�d�<�'�?����?�2�K�rR��"��zSvtK!I(�?�����ă覡�#�_����	����O̤1s��}�*�9a�W�>Mt`�O`˓�?a����S�d�N1Z��]c�d��jic�`
384�T�G�hƘp�O�)̴�?a� 8��2�d�A�jJ-�rϥy|j�$�O&�d�O���	�<�ƵiI��	p��m�(�%����"�� ���'4"��<	��Z)h�yC�JB' aQ���z������?q狅�M3�O��AH%.������K:w B4��造0�Qq׹���<���?����?1���?�/����A%�
0#�\�У�:�ء��\�EXcAߟ�	џH'?�	˟�6_��E �"p\�=+��̝�h`�	��$&�b>awD�Φ�̓-|�X�KO	�d#���{~8�̓h:�H�����&�(�'��'�jhR��M h�H���m��9��'���'�S����4@�ɡ��?	��%` ��%�0�pg#�2�
�"R����j��\%Ѝ�6mG�]!8�����	�(�'�B�إc:t]�EX��D#^��PX��'MY����[v4�!��� *��C��'e2�'��'q�>-���1R�tSΆ�m�N���F�]t"��Ɋ�M��������OT��]�\e�e���Ed2	�GX�U`��Iޟt��џ`8�����uGBX�Tg����>H��P��"�A�0'U�J���&�X�'���'tb�'���'-~��K�5�`��S;��)Z�P���41�6�����?���䧄?�j�4 ��p�!E�_J)H�+����O��d9����\L�g��?y*���
�3W�MI�o��l�'�����LJs?�H>A.O2���ʒ>7wT(`�ȍ�@������O����OP�$�O�	�<� �i�bx���'�~}p�g�.m������K�w��#��'r���<���?ͻ@$R�����sa��x��
??\��M�&�M�Op����	�r��5������	�!A�Q����!���� �B8O��O<�D�OP���O��?�`�皗o�����PR�/� \����ן(���M[�/��|���?�K>��f<$<���l�� ��%µ���?���|�
T��M�O4�9���:O@=��L%Q��a�͗��M��?QȒO���|���?��"gZ�3PK�.-��9�h*<�����?I+O20l�F��Y��ڟ���J��A�-UHtk���Ժu;��M����<q��?J>�O��pqN�h=rM� �S�P8�x�,ߊ���i�i>E#��O&�O�9;�b�Pt^��C���ɡ�-�OJ�d�O
��O1�|�u��fCޱ&�``���й ��+��k�mc2Y����n�����O�%��I��+J-:��՚:�6�[�O���	!G��7�1?!�� �X�D��/�� ё[�a���拄>3�V�ʚ']���H�	џ���ʟ@��m��
έu�J���E�fvdɊZ����	h�b���!�O����OF������O��"\P*�Z�M	z���"�w�����OڒO1�(���	l�2�I�>)�`�C��&R�0���$�+���I�?��0*�OғO��?	�|��ȘF��'�H|�u��h�PX���?���?1/O��l�r6������ ���B�R����5Uq�(��2��5�?/O���*�	�Bb��!r�����_���B&\��w��:�Z��J~�W)�OP�o�i���s���3Ɛ
0$�D:
�'&$d
s�	�츇k��p�=��'I�6-��&�z��?��wy��)���9k�q��$o��)�'��'�c�=.�ƒ�L���#eB�	ӹ=�FlH��K#	Y6�r�'39��O>���O�):'^�i��miFo�,\�@9T���[۴��)S(O��9��9Y{����L�W�M8cJ�?�p	�'�2�'ɧ�OB�{��r�P��T�] ?�\���h,X�uiGY��sQ��hr�]w�	fy��� N����GT7��ř�մ�0>�t�i�BQ���'��]qP�G2y��c��	,z��',���<��?	�XsjI�σ�}TaIDϽ;��VhϠ�M��O�l�1�T��`o6����V���=1X2X��M�9 �*H �3OX��� (%x�g
�4��d+GVq8J��?a��i��P�ɟ���(�ćB��	I&@��k��@�v(��h)x�O�$�O�;^I�6�7?��&L��
 e�xh*�-����@P�.���%�0�'d�O����Ƈ�=�~�Ӆ�߄�h�j%�� �M; hԛ��d�Oz�'X�ZC��?�:��J/:/X��'a�	͟��IP�)����c@)�cd�������>���V��M�3T���,x��D!�dH�����á�1M=�U)w�ˎz(!��Nۦm(3BS�pu��#Ӆ�y��Đ���6d6�'�����<��" �D0�Y�9mn	
⊱#���+���?a�h��M{�O�R�3o`������J$NP�*�� 7z���Fks��d�<����?!���?����?�)�¨{��̕z����%�K8%�����ʊ����rn�yyR�'i�4�4���"am�{�b��]8�yp*�O��b>)� k�ᦥ�S�? �@C�˝+��1�H߱H��l�9O��	�H���?�d�%�$�<a���?q���X*�$�@�ՓRI^�ڇH��?���?q���Ʀ)
�ˉ⟤��՟<BD�n�z@i�D��n)��T �a�����O���[ K�Th6P�2��&�6!�sM#?��X�i�Gڄ��'k����?�VeQ�7$��g��S�r��D��?����?����?I��	�O|���'�� ,�	�-BQV�Ī�O�IoZ������h��w�Ӽ�PoT�[��!�&V�)�4�yE��<����$�)��6�6?�≕�R����T�&� 0%IU~8�B�G��Ѕ#H>Y.O
���O~��O���O���Q��2@_�%��Iي(C�3�̩<y��iN\��'I��'���y� ��^k��l�n�ՠP�ærh�I����?�|���[����h@�\5>~�ГWI�sP��蒸��'�*��N
ڟ<[��|�^�q'&C�o�l����va2C�D۟t��ӟ��I��sybgӺ��u�O
�%�+%���i�?�z$����O>�D8��^y2�'��	
05�1�uo�3'MM�4HқO��z��W�I�'n>��&B�?��d����w
��c`#Ȩv��x��$Ž6�)��'7r�'gb�'%�'��t�0c�C�pD�7���!m`���O����Of�mP-@<�'\��|r��?-�>t`͜�rdAcƩx��'Lb������Y�������J�0�D���.���Xj�(�'F�'������'s�'6`�a��_@b��)�4�)f�'#BW����4O�J���?������Vl-�W��
6MˁA1��IHy��'/r�|ʟ"	�d�ͽ*�`��nV'Y�6��cc��aF��{��|��i>k��'���&�`I��٦!1��b�᜽$�8u�4B�ß��I��@�	˟b>��'o26��x �	#�n�c�K�>ƼM�@"���I�� �?�-O��D�^|��˅OX&?t�E
4��P&��Ob�p�`p�4�=��᳆i��O�t��	�w� V�ܵD���'��	ɟT��ʟ<�����	^��o˫"y�PD�³m=��4M��%[۴L:��?�����O��w ��U@���$��c�B&8�Ȳ��'e��|����s��=OVH㗤�4������&+�X�R<O�MS��)�?�� �$�<ͧ�?1F�¶gf�8q刞%�z`P��,�?9���?�����զm��a�ƟP�����s.�/� �� � �5a�E�c�S����d�O �7�D�;�04��,0Q��H
U�ѩy,�	,`�>u%��S�Jb>]S�'�J��ɡ-(�911�E�q�x��O�RP��ܟh��ß��n�O����?RXa�^����A�L�* " c� ��&��O���O��]vo���-ӹf�R���gS�Q���ޟ��	�t1�k�ߦ��'�>9٤J�?���i��p���*�X���#+��3��'��i>��	��4�����I�2\�#���~�L���J�J�� �'��7M|T˓�?)N~J���8d���\f� �0�&7��*O���OؒO1��Mq#��+:=4i�Ч!a���y!��_6��tyrE�y:���䓁�L����P�ͦ��� ��,>A����OR�$�O �4�&�W_���� `���/|b��eh#%H�|�6��B�'��O���?��?yP�тK�^��U��7��l��Ci��-�ߴ��$��.56�X�O��O	ǍݒJ��]�Ɔ��^Eb�MI��y��'v�'���'����'�����B"�X�g�J�_h��$�O��$�٦��,m>��IƟL%�hLT�c~f��A�t�S��IA�IΟ�i>!������'��o@�C`�-����m��ȩ��ˠL�d�������O���O��çu�N�x�ºG������אJ8����O�ʓEs��T�j �	џ�O���$DU���uk�c��P��	�'I�Z�D���,%��'0�^L w��M�T��%!��\��
#��a��t�ߴ��i>A��Ot�O��#�����R?B�Kh�O(�d�O��d�O1�f˓?��f�C7O<��Tg/���/U9�F����'~b�'�ɧ�4W�X�	�w��+�.1_�h9�FE8I������`�ͦ��'�ʭ��a�)O�5�1�I|���3� ��=Ya<O�ʓ�?����?i��?�������5i2��AKɋH�L�H�Ir� �o�'�`=�'�����'��w��u��N�aٌ�J%e�_��U���'��|���M�mӛ�?O�L�p�ɣ\]D���@$K���S>O�<�ׅ�~B�|�Q���ڟ��ǎZ�J��MCn��q�ꬣF
�ٟ���� ��ky��t�\�3���O^�D�O�ӑ��_ �-�V�oc�9���,�d�Ov˓�?�����M*�p�W�ETpB���QMNE�'���d,�&̚��6��dm�韜¦�'��b&�N�ׄ�A$h�s<�[S�'�2�'�r�'T�>�]*=���؅)��~�a`� 2}����I��MSB/�2�?��?AH>I�Ӽ���a�E���~�����A�<��?���)��!�ٴ���S��H@)p�@1I�┊�i�c~��v�J�����O`���O��D�O���0���p��P0�]�Č�
Xʼ˓%^���f9�ӟ�%?U�I����B҈��/�>C�"�`��'�2�'�ɧ�O �1� n}PGD�tVZI���x��e�W�x��'F��z$|?I>�.Oh%�N�~�J�ʂ��F�i0���O.�d�O<���O�)�<Iq�i�J@q�'��I`�%0�Hm�J��r0j����'�ҟ|�O��	�@�	��S���w���b��yfhL8Q�_EU�(nt~"�D��'����3��<`���hqa_�=���K�<	���?����?���?Y�����BB�!�AN`&�FX�yN2�'��nӰ,S&?�����O"�O����QX���lڌc�^a�H(�d�O��4�~��5�qӐ�Ӻ�䧖�|}��"�M9k��9����x�N���(bN�OB��?A��?Q��uʔU � J��h*r,�.4d�����?	.O�l�z�(8���$�	V���	R��ևZ�?i}������$�<Q��?�H>�O�>�;����dMZ�A�q8��bt쓬C�8�� �ib���|rԩ��d$��a��6'����^�$��jb+�̟<��ҟH�	��b>�'H�6�0�܁�$�)J|9��P�qe\ �m�<����'��۟�kD`��N�f�ץ+t�=qF�����I�>$�mt~R�S��e����ā*G�nm� ����ɚs,��$�<����?����?A���?	,�*xXX1� @�g����|�5@�˦�2@Zş4�	ޟx$?�	ğ�<n?��Q�)�n�@1I�@M�2���ϟD%�b>�BG ƦA�N�Y�3$P46lH���*� ]�'}���h?�O>�+O��d�OFHA�Իm?��xUb�,SDi�m�O��$�O����<���i��d#��'�r�'PL+C�U%9�"d�sˌ����V�d�<!��?�M>)U"X�+n(���8��,a�g�W~"�ӭ7C�����iVړ��ta�'��H��	�n͡'�M(��!��'�R�'&R�S�X�΀��^Yx5.	����A�֟���47�*!�-Od��$�i��#�O�"^:��*�SIഛ�p����ɟ��ɳG�n�t~��T8����'Z��B7��c�Fy�M#Gb�*K>q+O��d�O:���O����O4��E�v68I��#>���p�*OV�lZ4`���ԟ��	d�s� )��^�U�z9�Pg��)���Ky��'*R�|��@�[<���XL�i��[-	�k��C"����Z8,0��A���O:ʓ[�z�`M��D�n�����CG�4����?���?���|b*O}m�0[��ɩK��07ON8J;~!���,��Iڟ��?i(O�D�OF��K2=n>��D�	>�r�P��[79r�yp�l�z�nݐ�P���8�>y�u@.�M�#�ص��!��9p����4Ʀ�A�\(,�`�f:�Э!��߻ �Ea�3d��p�`��s:��蟚�@�Au�1RӋ7�x���,KY�ܰ�aH��7�~%PR��ߘ'�|-H�ޫ.
�!�P!R^�.)W'+T���
�A�9zU�tj�/kI�A���ۡ:2��[�"U B�~�R�%!@�b��`Dً=r,!t�%Z>��Ԡ��y��͈���Hۂ�¤ �4[1��z�K܁����
+F�=SU��+J��!R爇(����
tn�Y���3Eޛ��'w��'j��x&��>�+O��$��(��+	'�^�kā�0q�@"{�ޓO����Ev�˟���ǟ�
瀘�F&*��bW!/G�A�1�M��M;��#�.�j�U�0�'��|ZcT���I@- �TY�b�#V��1�O�,���O.ʓ�?I���?�(O�����Îtb�S�(h�(4�ВHn ��'������&�4���������J
�7I�,R���Cg�c�b�X�I����Iy��_Q<p�<%���!gӯ6.�0�!��6-�<y���䓹?q�H����'�v��TI�S���Ý��`�O����OH�Ġ<��"ԀV4������4ʘ))�l���[>�ܱ�iĬ�M;����?1��v�������I�EV2��t�؆Af�9��#ܪq827��O��<�"_��؟��	bj �D[f��S㛶h���sm`����	 L�N��?A�OO�}y��.h�x�F�ʢ@�VL��4��Ā�T�n��h�I��yZc��5�@���Dh�](���O��YS�4�?y�L;��B��&V������f�{Ei�`m��ŕ�0�46��OV��Od��HF}�Z��0�fܣ"M��o��D�S�T��M�c�O���'����Yh�dip��ܨ���>�tHmZ��`�I�����锼����<����~¯U,GF�'���� D�P�+�M;O>y�ˍR4�OfR�'�ˑ
]H=�f���!��A�O/Tr7��O<T�#��|}U�|��G�i��q���P?L���=7k�|���>��M����?����?Q+O�����q��A�%M�o����d�˅;��,$���Iǟ%����u��;\RPh�s��ia���M������OH���Op�a��ĺV6���h�BT;L�8� q�VoT�T��U�h�	؟t'�l�����'�^x�R�'(~�<�m˜<b������>����?)�����ܬRr`%>Q��C�<���@�D�#���b�և�MK�����4����1�Ġ�-�u�q�#�<�rE�@<�M����?i,Oֈ�K����s��9�o�>����P�?���w�)�d�<���?AO~�Ӻ{w�΀[�r�!�
��\+����
RY}��'��R�'���'=��O��i�A� *�3A2ԭX�Aѻ�^��1Dh�B�d�<Y�Pq���'׮u � �wN *��
*(0�l�� u��͟��'���U��'k� L���g	N��R��T�@U�İ�m;�Ş�?ƈ�� �<�d-�'��#�c9��'���'�ĵ��B'�4�\�����i�eZ�RXl�;���,%��vk���$+�dV��O:�$��Ș�# �W"e5'˽}+��(�{�h��%B������s��f�h� Q��Y�6Nҙ{^��j�x"�C����O����O�˓J�ls%�!��Y)�@3&6����6#��'M��'E�'L�i��C׏�A���(��N�~�ۇ�aӢ�ĳ<���?Y����K�z��9̧�`YA��6M���k�߀1�J��'|�'��'}�i>-��
,����$�.�
B��q~��O���O8���<��MD�!B�Ov�p�q��
0�ƍ�Vk�,z̥s�av���$;�d�<ͧ�?�I?����G�>�Z�H�� b�J��tӘ�$�O˓ y\a�e���'��\c�2AgFN1"Z�9C̈�(X+H<+O����OГ���؊�Ț$K��F4j��1Pбi��_.�i�ߴ'�Sҟ�������=9(L�����R2�I�\�O0�6W���I��ЂI|2M~n�Z4f����1)�00���4��6���F	����������pyʟj̠v�;8�(�܃����`]K}b˟&�O>	c�$��H0ǉɟ�X����U��M;��?1�R5���/O�Sy����0�@U���.'�H��D�Z(��tFx��3���OB���O�����F��0x��bٵ1�^u���T���	0 |T��N<�'�?I>�;�������-gg^�1d��.���&��	g�I��\�'�b(^�Z���r�ߙd�؈y�F^��怣UZ�p�	؟�?	��~��@�"l�!��U�|CB���!׍�Ms�k�K~2�'r��'I�I6p}�OU�8 `O�8(����ME+$.<q�Ov���O\�Ot��|
���p��F7?T�Q�T-XI�x��S���	ܟ���eyb�	"�l�rjQ(O	@MW���pB��ɦ���h�IVy�Ojr�~z�h��rTY��	�/d�!� �Ȧy��؟8�'��Q�)���O����h�AT���Mz4)Ɯ[
�0�x�X�L���H$?�iݥQ2���YаQYv(Q}0P@w�>���'��K���?I���?9�'�����VK�s�TP���.p��(�Ѷi�r^�|���.�Sⓛ(R���J͈)Q��"7
�06��xp�m�ٟ��I̟4�S>��d�<a��ˇp�T �ᏼb5�$����%�V����yB�'0�x���?�H�}���K�i9Q�r {+�Nz�6�'�2�'���W&�>I,Ol�Į���F�s�����P��L|+�ϫ>�-O.�擟�şX�����P�V`ee�K�F����>�M��0���sWY�ȗ'�_���i��Z'��V4�����(+4�>����<.O��$�Oz��4Q�2��2��L)�Ó&W���k��*2
!�'��ϟX�'���'?��
�I�F��2M��=�Nqp��R�'�2�'��'�r_�L1a���D@-�4Ad˫t�"����T��M�-O����<���?y��&<��\2��谦��dT��YC΄�[E~��W����ן,��_y�7��맺?��	N�\br�#9�;0�7p���'_�����	�� jd�1�sӤ��e�L�s�ޑ˵�8<��xز�i���'��.x\|X)��`�$�O�ɕ1k�"����Â�Qs�ÂI�m}��'�B�'��#�'�_�D�'D��l7�Գ'��x���_z�PlZ^yA�7!�7��O����O�)s}Zw��8x!ظ~������[#�jش�?�e�R`͓R�s��}���I+�e���"LTt±�A��q�7d��M����?i��R�Y���'uZ�6����
��ɇFLd�rv�wӺm:�6O|�O��?���c|��C�p9����-O-V�!�ݴ�?���?ip�2��	Ly��'#�d�suh��
:ϔ���Ʒ7��I|yr��)��4�:��O���\284�)�%j>T`�O�WZn�Ɵi�b�9����<����OkL\�"H��A�H�<0D�S.�p��I:|�Z�ޟ��	ߟ$��ȟ�'���!1�J7t��5)�?;��P5�������D�Op��?����?�ԩ�r�k��E,�*4۶��fj����?Q��?i���?I/O@��D�|����'L���f�
�̈`k�Ԧٖ'�T������0�	4xh��	-f��!�M� T`�:��x�ٴ�?����?�����D��!m��O�Zc�X�I�����F4Fd��4�?�+O���O���2bw��|n�!PR����#�#>LI�`!��\�Z6�O
���<�GZ(]���џ\�	�?	Q6�R�k&�")�4&�1Q����$�O���O��;OR�'�?��Or�!��d�5j��P�2E;�2}�ߴ�򤖚.3\�lZ�����4��5����&��Ι�e���ъ����U���'���^&��Ļ<��DIU�6BT1���1"z�P�p�W�M�gEK���'\B�'@��ƴ>�*OB��ׯ� T ,AA�T�/s��J4��٦9q�B"?�.O�?��I�h�h5�W�Cx�)A��5M��9��4�?1���?����;{��ISy��'��d�#m�����>�	��B�՛�|2+���yʟ��O6�d[�CU�1�gK�&��P�I���bel�㟌���/��$�<�����Ok� X�٢��$�P�(�/����i�ɝ��yb�'�"�'�2�'W�ɠh*p��!��z�D�xìԜ:�(|�A"���D�<�����d�O����O��Vb+^ȉ�/�
<	"Oه,)�D�O����O��$�O�˓nt���1�( �u���	�f��Y9��,+R�i�������'�"�'��E]��y�-�$L� ��	�<E:#��UM�7M�O����O����<����	7��O�$���AҨF}�;�(S&H�u�1�s����-�D�O��$M�a�d#}�9cEv��cHNAy�Y�ҭI��M���?A(O�5C��Aq�ğ���=c�e��ΟR6�(��&�$�jI�N<Y��?	"o�&�?�K>��O�|�p$��;
�x�A��e �H��4��d\�6��%o������O��I�r~R߮X��ܛ�ѣ(�����L+�M���?�&m���?YM>q��4D��v/ڸ��i�q �1�����M�P��Z�F�'���'����"�ɺv���{����}��(.�d���41�,5�����O���Y56�C�a���萧��;o�6��O8���O�(d�S쓑?1�'�
����H�)���!£�7�|-�޴��Z�m�S��'���'���	�f�">�|��c�1��y����#z���>9�������lӶv��aǣrѣqHl}�o���'���'"X��d�
5T�0�LX0��w�W�G�HKK<!��?N>)���?����03u�t����{k� q�Mܓ}\0�<Y���?)�����¡}N���'uJjܨF�	6�H03d6>*�T�'*R�'��'+B�'�Z5��'6n�J�QO��]��fG��8�hs��>����?����@%Gu
�$>yAtH��Z#�yr����B�E;/w�)�ڴ�?yL>Y��?�vj[,�?YO�p���*jg���g�ށ!T��!�OjӼ���ONʓݠ�8ԓ��'�����5c�=���V����r�0Z4O ���O��8O��O���<~!.�$g+2n��G�ik$7�<���>	&��E�~���RW������	-�3vM�����|�b���O�,y���O��O��>M �
ݨ\�Έi��4(.�m	�|Ӑ�y��٦���˟��	�?q;�}�
��1�z���ήa�a gJ�)\6��,��$"��>��˟�����}Fh!+c�P,a�0K��)�Mk���?��r�,����x�'���O���/�:|a3�(�,d*ֶiY�'�He2G�-�)�O����O��BR���ik����?4UzU��M�	1T0���}R�'4ɧ5V"�p�����;���O ��$�1j��D�<����?)���P��ꝪaK�^	J� *��+AT��V��O��$�OV�d�O�OT�D���i�Gўaęb5'�.Ը���Me��!ĝ������@�	XyB_�Y1R�S�(�� ���іmz��jN�Y��?���?��(^.��)��y��!����z_�x)'��!��I�t�	��4��P#�E�}���'�P��N�[>���I�,����G {���%���O˓c���&�����i����&��,��� �{Ӝ�d�O��4#l	d����'������`���BNO��\0���&ɰO&�D�O((��r�4��-Z���x���O��5�'�>�ȃ,t�p�O���O0D�%*&�ӡ���� ���r�<n��p����"<ي��MV�"lh��%/+��U�LԵ�M��
|���'�B�'���/���O�����=x$�YX�-\ ��7K�⦕�q�!�S�O���
�xҥ(�U�^�2A�őg�7��O�$�O�A[��a��?��'d,Q��h�xL���A?7$�j�}�$����'��'��DE2���i�n�f�8��?H�D6��O�U�L�	����	\�i�JCg�^/���$ @�j�걣��>	#�u��?Y��?9.O8���n%\%Pe)�",o��ۀ X���$�(�	蟔%�,�I�p���#6��=�-R�gfDIa�`%2) c�L����i�lڟ �o�eG,ρM`e�5��t��Ԧ��'�r�|�'��ɤVv6��}�ؑPl�b�0���%^E�I˟L��ڟ��'��u��"�ɟ;A`B(=o�P���%M'z�LoZڟ�Ij��xt���~�q-_a�L٢��I���$����������آ��~�4�'��O�"d	�	W�RxHb��4�b��6���O �0G�GxZw�r���	{$h�Q"Q1o�>0ݴ��D����to�
����O���w~RJ�C%|��j�p���&aդ�M���?�׆z�'xq�ƥ����6R9�@��> ��}Hg�iwXA�4�f�n�$�O������?���(�6$� | Xl ���u*^u�۴ �pDx����O��ӷa�q���u���s�qxb�צ�	ԟ8�ɀpc@,�J<a��?��'� k�
@ rX�=p�b͌HH@Ȫ�}Ҥ����'Nr�'�r��7n߆%CD����@i��XE���j���h��?!,Oj��?��۰K��	��'k��������D�$�8�v`<?����?i�����<^���Ɖ�.'�Ҍ�G�j|�����{�	ϟd�I��?�R��:<dZ��G��3����B�Y�\a�<����?���?1��C�
���O0@�k&.�2VA��iw^q��KTͦ����4��o���0�']�=��t�? �|��'�<1%kGܠ��GY�<��ßЕ'7��3d/�'�2CO�
D��aR:��0���N�6��O̓O���<	�i�s�4B�^qI�� ݘ؁ ��D�6-�O���<��[!1��O�B�O�^)�ġ�--�B�sJ�Q�ȐSG#���O�������'g�Rd#�c̟(��!��:E�lJy���'��7��J�t�'���d=?��gD�C Uh�W%x�X�y�%Nᦉ�I�|�5�3ݸOs�%���O�e߾�c���=���9�4]p����?���?A���?Y���)I,>��1XpΊ�G�z�����#_"�$�'�R����I�O�1XcA �:���WW*���DEΦU�	㟬�I�G��H�I<ͧ�?	�*d<�YD&�!d8��R�ݯ��= F�ć�)1O����O&�D� Y$�#�úY��|aƯ[�W�l�mğ�8@D�ޟp������OԒO&�"v��%�Z�i5��U��P��m��8VU���?y���?.O���R�9b,���"������(����>�����?��GS�%�Ge�.��u�%�̲[,𹕫�f̓�?����?�*O������|�㢀�~��<��_�}@yH�-\A}r�'�"�|b�'�¡�8��Ć;�dE�2�^
WH�Y�����	ԟp�	ߟ���ݟ$x3 �E�t�'u�jM��J���Z�ՂgLTYcA&v�`��7���Ob�wS��$��r�� C&��]���T
��r��$�O��wK�=A�]?��I쟘��ovd8b`�8��0�v��~�ZM�۴��'P�"}�'}�T��
7�TH��I }b�%8�4�?I��E�,1I���?���?����?���TܵO��4�Ǉ#��ˢ��զ���[yB���O�O��Q#䏒]��9 ���v3�D��
?�6���0>��勦#)8��Ā�8��$��o�K�<�e�+#*��y&�ޒ7\��H+�(8N�bc��i&�}�g߃2�J� C`�!7�	9��ٜ+d�m��)�<M�� �/6Tx*3J�,
R ��<: Z��<��y`b� �W�8�a""�;�j�I�02"��e
�(6j����=�tG��c�8ga�=3�����!�?Y��?���=&�.�O��z>�Ue��"�$����"�gL��(�#�0R ����՗T ���d�&�0��R�	T��8C��? �l�kbn�<Z�(ZB���d�tY45It�9�x���d��0K�
�xc��d�Q
�����	C�'
�O�uB7�F9,�r92��d�q�"O��1�C��n0���*c(�ȡ���U�	uy�oɠV��?�l�`�b��ġG��<�����?����5���?i�O��M�d�T.�|ٹׅˤQ��q!���Y�����8�|�H���y8�PQe��->�0�*D��,a��� $tf<��N/J!f� ��Ѡ8�x��[;�?	����D^�{�T�!���8e /A�]��yR�'Լ0u�)S$mb��L�FiJ����+��|�W�iT�[�  S��H�0!֪j��0�'��uK~�9��|�����Ia� ��V��w@^�)�lH�b�	B��0���?")��)�P�/lm0�����|����#s�~Uq��;��L0 ���$L22�9����[r�%0���O"0��]���)�QaT�b�A�@Y���B3��.���	ɟ�D���'��JA%��O�� �G�j���'�>-Xdh��s��J�ub���3�i>�����$~9hmr¬Q(���f�*\i�AlZ���	��Q�ɗfr��I៤�I՟�]"v5�em^�Hs{d��,qz�cb�i��ɷ,�j���1�3��ƿ?��-�w��89�1J�_$&�d���P9����N��q1��L>A��J9Ɣ8K��Yp���h4�?��O�)�����	.�^<�҉S�I���� B�=DrC䉐r�N(�b�#"�lH��I��jp��8�����ğL�'���8t�݅fH�h��[�\�69�k�l�~ma��'���'�R�m��I����'ZahM�4� �	jె��
�8	W��HmĐ��B�\��W%	`H��r���f�f��$���U�#aP#?�2���Iw$XJ�'2�9e�Q6
���m��4���uQ4����.Nى��^������(�DG>v�~�pfMA�y�Q2F.ƕe�1O�mL��?S�Q������N@HVES�v�((�Vj�)�����O��P�O��`>Qu�;�찑����\mZ&r� �D��"q�H��PJ�'M,���ؽC�#�-O�u��� 3fd����%Q�"8q��
P)��i�!�'x����?�,Op-��X�%�l����d~ ����D�O��d@�>�6��C�)u��dkc)�	L!���¦!�V ڊf���	�������%G�ܕ'f��QT.lӆ�d�O�ʧo2 ���D�|(�A�X7N6F(�� ���?�Sc�}0qB	v�|�����)�|�) �Z��7-ױtZ�	��D�P����U��4ZeEǞ羘x��Y��M3��'��	�*M>�ѡ��U�
#1�`;�I[�S�'	¤#a�ʲ@���ksE�+�����S�? �YY�-����,��^}�,�A�6��|�S�I���I�)�!����R�{|��Aܴ�?���?鰆� ۠�����?����?ͻK޶5����t�=!S:+�鳌y"&�!��<��͒T,<舵��k��:�e�@�Ak���I>@����Ȫ��`��w�	�<! ���>�O��A��c�@aHt� v���"O4l�ccF�WVQBq��/B���" ��PY��4�X�O�q����:.��}�̈́~"FŃ@eX�F|<(���O����O����Z�t�'��I;2z&lK��q��0b��b�IY��RBת(E*ͱ�j�?:���ã{8t�'!(ͩևM�x� ��#@�������,�?����?�����$�O����D>xlzRjC�f4!Y�H1D� ��fš!�<KqN�E��yq�2����<aqMR�����'£]�+Ǌ�b���^5Yb��r r�'ֆ��A�'-�'�,\���E�:��O.9(F�%md�B��/	�X���'׬ ����z&i�K|�!H�o@�36CsD�V�D����c�џ��Ov�D����I�䊕��şo^��b�����'xb��ӷN�p�;g�(|R�h�nW
K����D�O@�\��0�(ނY�����	@R�\m��.z��=Q��$R<
�T�R"'��b��P>m!��$�$��2�����,g!�$�_� �*��Tl�m�`J'z+!��*(+�0��C�}�^XA�)���!��$I��#6$ l:V�1�i �!� /�n��R	ӰP�!�5հ,�!���X��p�'ƈ6��ѷj�	Z�!�$ʺmդ`�2�
B�Qʅ��!�!�-�+ҋI�N��"	*�!�$Ҝ���`gBc�r��e͖�L�!�䄫Y���$��'�d�è!l!�wf(��m� xy ����ٱu:!��C�[_v�����[m�ht!�dA�ب�c�Q�aX��R�E�W!��/dQ���G�/HNQ&d�j!���v��zQc�9�8dC�d�]�!�$F1x8����!q��AAv�֋B�!�d��< �I$�3k�貄`>w�!�Č,��a(#�XLĐ�.�!򄖀D���)+Dܬyv�K�1�!�Dy�m!2M��l0���2$��!�$\Zu�ĳ#�#�d��L��H�!�d��[ ���B�l�\���V�!�D��9�D�C�H��0D<ڑ%�|�!򤆅?��A���,��`CԢ�!�N�W!�)�7B�.5���cΎB�!�d�2n�Y����4�1@���P�!�O�-�����gX�2�=Z�'˵�!�$Z��Ų�EO���R�^�!�W�{�{���PK~1�Ă"}�{2�VF<�`R��OD�(�E�g1�l�q�N7L�YZB"O*���J?�v�b6�V&<4�T{�����ng�u�����H�dAR�iˢl���j6J��$"O��0�͞B�bĉ�+G&n��#�ɜK��i�-G^�D'�g?QSF
*{�DЇ"F.�YP`KI�<A�Q�vb]*a�Н7�Z�*�@�۟x�'קn�9��'�J��OA�c�X9ٓg�O�:rߓ9qv��R"3�Z7��_��pz�g	 X�,2Eh��.�!��̸k���x��>e=�e��
9n��O,|aG�ٛu�ڝ��Ɇ&Zߴ)ʗG��B|!�c�i�!�dq��em� v�n��f�� R����HO>�7��>*U2��.��颐4D�\2�l�')
�� �D >��m���.D�L#E�I @�t�ea�(���R�,D���BAM�U�����/�x���!,D�� ��A�M,1I�!���Q�"O��R��
�Q�m�!B��t(a"O���ݨW�d��,٪R�l�E"O&=�ƠWHрH�኉(wa�Cc"OT����$�$����(w�JA��"O��+�j��J�h0)P��67�]��"Oiԥ�+$���aHN��p�w"O����)T
��-�4)�5*�;
�'k��!mƁɰH̗o���	�'�&5qp�޲K����Ҩܷg�\i�
�'���`��\>�:ҍ��Y�ژB	�'���W�x���&f��9�'3��B��S)V�,�D�V�Gpلʓq��,Z�i[�b���#�$�*����ȓK��VZ�4�"���T�[�VL��z��3w+�/�<)c��IsȽ��vp�0���/y���$c�:¼��c��\�@�܌-r� h��̛m,L��N'��*�Gċh|z��G�u�^��ȓ;B��_��*�� hPXJ�ȓY򄀒��/RUZt��m�~�<��^:��ķ]�R�QT\D��ȓG�03��ҽ(Et48v	I�NbԄ�gyH�qƤ	��,L��SL�DP��HAn�bI� [��,*P�4vr��ȓ�j�x�i�'\뺡z��@.���Q�
Q�?�P2��́Q��ȓ]���gI�R�~9R�L;v�i�ȓ{B����H��W! t��B�\̅�S�R`�=!u��XېT�d�/�2!hSA]V�<���M��(�Sҿg*���4�AP�	�{GDa�?�~��ʇv�x�`�͔�,��x9U�]G�<IqA�S���́>$-�ʞ�t�� �6ɒq�Y�E��<h|��}&��3u�&	�}3�'܌y`��p��8��1��(yh�\�F��z�x	�(�9�j��
ե�졪����0K���p���@}�<�O�~��	���Z��J	NI��@n��c�Ͳ&�ڙ[�Fڗ7�r ��I��'P��{6C�p�hQH�!{V��9�ō�c;�'^�>�DW���ͣB ��f�j\ ЄLl��I>�Ի��t�ȩ0L ����҈�ī������� I�j�ڦlϸ�~�ħImi
��'��Q��J%k�0!au���ؙ���7fdP�"v���rǃ����'WH�2G���l��7͈'t�82��>Jf��W��~B�Ec^PX9V�)u���GE^�5�e ��Q�Uޙ��˔�d��W�A6 %�y��}��'-�.x�0m!Pn�'a��d�$#ٗcp">���m�Jl�" �LP��� ><0�`����501�ɂ�0%؞	��[���yC�c�(��'��>����s~��[�=���)	>����OJ�v�	p��M.cilmb"jܬ?�vY:���O�%�d����l{���샓;g�	�D���=lOܙ
��N�~����O�x��
2ǅ�P�lբ䏚;�|ԉ�쇜@��'U��'�T��KϤ2�Xe��ݯ�43� 4�T��CW%�@zu�[�C���U>S�\%R4\�7�<d�7�X
P}���ɇ[Z���n�?sX	��AKPOX�?ᖢǚ-?L<c#D7M��<b��&N��E"_�N+�f&v�PW̚h�<9УU�x�7�ȝn���[~�g��{�\# �I�W���I�����<ؙW��@����v̙�m��`b"O�hj�вQ�����*;t��D���F��,s�韬`�K��-�q��'r����g��,95�R�Z�y��'}�)�6ǖ+^-�bD@ʺo���hq���+����.�&�$��
ۓX��Y�Eǜ'>�X�䆓�s��%��	�),Tp��ى&|牅"�Q���_�l�25X�C���C��F�Y�C�z�Q	��!zw.b���D�νK��~A�	:=�Ly��[8A����.����S�'3b�1Dd��K�m)3����@ϓC�Mi��%�$�/\��A�J�t m��!<2C!�d��<Z��.ZT�Wg�B��'\
�K�g�T�S�'rK<]���)
3���%���$��S�? ����W	�ؒ��Ur�������=[l����L�@K���V�B�[8a�h��!D�x�4Ꞅ���4b���HR�쿟4����4�t��g�@�O�%�̒C��C�I+�p@y4KF4>�T])���q��C�I�a����\9I�F���aĆ<5�C䉏6ֈ�hÊ	2il�@1�pB�Xkx�zO�.��	�L՞B�	,q�΁����0�΀B �j�p�RY���� �M�6	&������B�a㍚�R�S���p?�,��R�� �=3�a
.žc�Nu�2)/dR�s�'���)�G�;K�Xp�&R���C���K�pԉ�D���A���	Ҡ�,WqTq`�a��Ub`"Ol1�6�԰=�;enA�Nk��C$�O��h�+wTS� �0|r/��D�j�AEO4)�苰��{�<�WKV-��yPҤĳ�t�k"$@�y�t˓��M��������'�9z��i*�����$H���'"O�U��	�o��@���M�¦L	S�\�HɌP���P�v�����a�A�A	P53��� l<8!��O�L��֧�����s�f���"O*�x��L
Cla��NŨC3r���"O6Y�u��pn�%�g��nD��f"O��� D�'�}��$R*���"O�9Pv�
�a(��=g�0���"OTH2 M�Z�&�C
=�U"�"O�����^�R@(�Q�uƈUC"OD%j5�M�]��[�,�#���"O�-sv"�#A��U�d��.W�c'"O �Z��ŎP����
�U"O4y��[�~�4�����|:l"Oi���(c��i�2*�'(T��4G�V���$��#a�R�3
�''dir$/˖t4����8L�����'�B\�ulPj��tYB���H��I�'�Y@&!ֱD�>��!m�S�*|@�'c�1#J��n�� �E�M�DP�
�'Q�-j�L�$\lf�A�%DKF"�'�,�
A�M?��В�.I�F�p�'f��a��p����/�%o���
�'p� $��{NȔQ�C����u
�'Xp�c��6�L	d*��z��2	�'�6D1f�+8ޤ��sI+n�8��'gp�ZK� up��
'1 ����'�T �⣞�MM�� ��?%ƭ�Ǔ~j&AG�V�T�X7��5 ���`d��}y|�(Ҁ�J�)#Ih<ٳ�Z1:vN"`	o����f�Yw��*֞�3�͋�js�|k���+F<c?��,J H-�H�Cf
/!�u�a?D�l�F/��Dsy�W
^:j5�}y��ܴo��)
�G��x������ؕ��>q'���G�G�OXJ���-$���<��cBC�Nv�ɳ��� �Z�P�AAn�1�䇟>?!ZI@������	� 3��@"T�Q���� ��^k��D�L�$H���A>3�� ��`�2������^�.����¸�)h�O���E\?Ԡ�jj�pq���I�?��0�֍ =��`���B�0��ȃ�X�
Ԃ��c"O�|�qn�~)�k�υ3�`����'��͡�P���|�O?�s���uP���h�|���ހ�y2�J����h��ȔW��
u�O���&[N�C�+շ��<���±(��x��Ǩ [�i�aB�\���,zrH��I�CJ�c�@E�$��R�\Z�$�� V�Y�ȋ�^/��a���`ڌ0��w"(]A�@ka¯�vG �	�$AX�<���
9<Ձ%VU9h��mR�<�d���_Ԅ�E`�<��]����P�<��ʘ6<(S ��7J�P�A���H�<� �� �6�y��� cH ��"O:e7K�9tI+��OA}4�4"O�� ECWq�$��+��*���"O��o�Q�k�
s�*�b�"O�%�ī�vi�h�E��� ����"O��FS�U<������qr�$�"O�rcfнW�f��锰3dXZ"Ob�ITE�;,aI�h�!1Az%@V"Ox��C��Nh�m�愥[\l��"O��#��%e����
�O�2U!"O� �&���,�h)j�IɄ~��|4"O��;`��a|8�Y&H��xh2���"O�+�K�2r�jH�禐��d�"O|�1w���Tf��%��q�s"O�#5H�7ݾ��V��<��̰�"O$m��|`��K�D^=ju�d�"O>���S�pF����#�sW���C"O���,�'>�
�6��($��"O�
pG< ��tC�9K2��"O� g�3?�P��Ȕ�"��z�"O�}㤤�4)���u�
�P�"O,�KS#Հ �m�U@vw܍:�"O��!� �j�S�-׀vcڕx�"OJ�(�$�l�ع2�lR(Vf`�E"O֔� �?��8�lT�5H���"OFq 6��7N��s�4��k�"O�@��ք6�$�IE�0(�P�"O:�bUυ,y�����)��H/���"O��S ςފ4*��F,jMɇ"O��[ ��Y���P�)�>1hx�d"O�x����2{~Vi �(H-����"OLh�@I"��qZ�g`p�{�"O������6"�f,��ĝH�i3R"O �;��M��C�đ�@(��"O"�q2�]< ��UC������"O	k�N�n��  � 6�`��f"O��"\��2��D{�"O�����O
9x�\)q!��"O*X�LFR��OO���X�D"O���r�]�1j�Y�ڇN�4=3�"O��c�'�A���rp`�q�&I�4"O��*�+ȓh�\�	EE��|x�	�"O�8�T\/ozxHs�	�!�(�r"OziɃ*��~5H�zL5�eX�"O��x`�7m.���	�F%8"�"Ot�uDN)��`j�@,'���"O6qkY
9���@CƵ���Y�<!�ޡ�x|��K\^���y4�MJ�<I���	�a8���I�F(���l�<)C��.�D����$����h^S�<	�FáS�8y�C�͡��ìPO�<�G�֑�
�bueJ�Gj�4���c�<i����`7 ��!4J����&"Q_�<Iw�A1��R��*��,�c
S�<6떲v�t�p'O�I�m@�BW�<�Vܢ&���1JN�a2$�V��I�<�V�I�Z���@A�'F6�i��A�<�/
z��2Y�DxV�z�<y��N����qnM+Y� ,���u�<a�	D>0��pǢ��ʹ��$e�h�<�KC�)�2m����"H֢�G�Ny�<!/�<!��Ia3"&���l_�P�!�D�0f�(�Gk�>1 �̓��߭a�!�܇8�P���ߔ.d�P�_�f�!�� ��ـ�5%B\��Èvװ��"O�ca΋Q68�����|,�P"ODP��,��� {��,[a"O,Q7a�h�p���&9��"O�=�F��FK|z#��?��@r"O(5��M�yT�ˊ:z�z��d"O~���˺`�Π��
D=�Ș"�"O�0��L&ok��آ냜xw@)E"O�����X��HP�\Gݸ�"O�E�R	 P�J<RP�H�%1�m��"O��jGL�S/l����	��-��"OZ�1��9�>۶�nT��"O���N�6�x|�0�ց3��l2�"OΡAO��=N���&ǚO�z"O�]z*B�,3��ʹ{0�p	!"O��2����6��Þ>-��"O��(�fZ9��8���">���"O�a��M�>{�(eĪ��:�D5�"O���'��[�$$�QD�d�"O�d���&�:x�-�B�A1�"OV����<GB���5�P�"OJ�
�^9�L訢`�7J3���"O�r1o�9l�~��oؗ,4��Q"O�PZ�^�Q��Q�,��B���1�"O,��#;��hSs�ڞ|ܐ�"O�����L-|����m���D�]"!�V�7��,RhU�5[FL�1!�$ �5I�2���h �� 0�N/
!�D�8$���(7@F+w�\4���ޕ !��	����˜�yӬ�� �m�!�D'x��Ҡn��:����'
 	a|R�|B�\+6��a%�?%���K)�y��l};�'\��LD��y�(�2:/B��UeA���)B���4�y�F3l�&pj�`���@UӐaY>�y���B��̦%πi�Æ��y��"U(l����6.�`�G���yb���]Ԧ���(=�-[&ƀ��y2"G�&�0XZQ�H�B�x�	ָ�y�mݿ"Ob���>@�"��$n�+�y�J�,s~8M
���l�����U��y�i�^�L��Ab'R�p.K �y�+ʠjv��0ˈ��H�{����y�H͈'j��$��%(2 m�6�y���T6v�v	��`<Xw���yr�#Z�	�u
�A�< 7�P+�y�ǉ#j��q���	�V]ȖI��y�L�� 2�L�aLQ:�vqQfNE	�y��D�A�H��앣~�X��t�݆�yB��F��u��P })��i���y�MJ�DmL��N�r9X����L�yb̛.&X�2cpJ�sw&ة�ybǉ)]�L{�5_��rG���y�F57,h��a2U��ܺр���y�����J�JA��!��y�
Qk4�
"j��rC���!E Ѹ'�a{�k��C��EB��O�BhO74��(Z�'m�4K�*��`v�*7j�/z�A��4�PxrU%(>�u�!jR;���r�Ƴ�y�脺C�dh��ɭ/�Eb�M �yү��I��YFɟz�����LW��y��"�M��I�w�8�C����y2!��7�̛��8u�8hj3hѤ��x2H�z��פG#&��) ���/I�p�h��� �I�0�.X s� X=z�z$�'��Oj���1D��% ���L6攚�"O4�yAT=3�(�rCE_?MY��0�S�S����E�6M����3`�/y�B�I/K�P��ؒ\Px1����B�	�[<�[um�X���Zɉ,A��B�\�PjN�~c��spF�C �B�If��F��	i�P�Ö
JJ@$C�)?2�yW��l�4���I�
<C�I'P�~����/~���Yl,C�	� �qS��"N����M�
C��9ʹ1!��ftb�g�F�$C�Iv��}���7��d��cJS�>B�Ɉpk�L���3٠�ADhվ~rB�	�nV2�Ê+\�r$���nG�C��0��Azãԑ/�T@giA�88C�ɑ&9��)C��:2�"w �%UpC�I�L3�0�%"`�(TCa�0��B�	!nyv ��2tO��`JW
��C��P�I����-��I�� 1 ��C�	���·�E|p#��Y���C�I�O'f��T	�|�4Lyӏ%WfC䉍�����[��u�էU5,�0C�I�cQ�����09�r(�t)��ZUC�	2RK��+Uj�p�१�+c�B�	�b{��A��$Ե�GC^�y��E�F��A�ǃˀ-��I��g�y�]�r��qb��ޟ(���f.���y"#ǥp :!a*Ϯ�.=Q�P��y�FM/?� $��;A ���s�ؙ�y��7��i"�̽C[� B�y��]�3�[A��k��=CeY�y�."�LS���V�Zű�C���y�&�-N' �`e�F2"_DT���y�CV;3�k���2x2p��N#�y�.����S.�	/�iJ�f�(�y#̐�nU�ٲsCZ=��϶�y�k_d=c6��:Z:.��6G�,�y��Ȅ>`�8#1��"=��í6�y�kpIxG/��^" 	�
μ�y��_~�@Q��� �<Zq�珍 �y�	�r��8#�
"�&��p\��yB�-Uox�0��܄!�.�1 F#�yB@��nt�]22`���@��L��y��5ֶ<�6���7�|ؒ�I��yrĄ\�m��E�*�H,+���y�G��Q%X�ZV�?"�d��E��yB-�6c�N����a���X�yr��`|P��k�6���i�0�yBC�?N� �ٞE�=�Cɽ�y�ȉ;���&��ApaHF<�yR�٣0�Q� �J4~mN)��L$�yRIM�zcFy �kV�eb��t�N?�yR�R��l�Ąd��A� �A2�y���J�ݨC��$^ �����y�*R/f-2���W����H*�yB$H<t��(��Z7U�t���2�hO���I=7($E��eB�i��)�	t!�Ĉ }w�Dk�������l���	`x�hT*Oovl%�V4fkfɘ�8D��h�	�	z�"r��[V,��E6D�@�A��j�n��B��o�,L�V8D��0���Ѐ�)vfзnY@$��/:D���&P>ar��S��3t'.\C�8D�� B����/HV�م��h�ƽ�1"O̕�4���cu��hҶ�d!��"O:�i�m_K��� �O�"V�j�"O� cv�šc��k$_6���"O�����{X��]6 <@��"O����޾sR2	aeUH�t8�"O�)��H����l��y�"Oj���޲z�.9I5*L-X����"OJԪ�F!d�� ����		�)!�ĉ�OJ��������)�IѮ(�!�d #]F��!�`��'���K��K$@�!��( 2�1���p
���X�j!���;Gb\���GZ��Y�,�2"!�$�!:�����M��jx��E�aI!�� �l���J�~.�x�'˲07!�ę5J�.L ��6J^i�d�,�!�Ĝ=Fx5`�ʓ�`��+�a�!�DNi�^p[R��(��R����!�D_�<������J.9�Փ�.ϔ@�!��)^8�KrK�ձq�{!�dʎc�<(;��Bn� )� ̝�A<!�dʚn� ���"}�ƙ�%H�1�Py��5�Q��i�64Y�%c
�0�ye@tJB�pU��=w�<�R«1�y�G\T�M0��ݼy��B�C��y�I�&'vX ���y'~�YB(��yB��P����2�HHR`�o_��yR�	�.�%զq���"7i�yb� ��ycG�f~��VF@��yb-��kO��`a@�+jm��څ�yR/	�s�(��m�<%z��� ���y"K�oDq��ن$�B��\��yҦ�>/�Ivd�!��|�m���y�!�	N�2�>����ԃM2�yb�4�����+e/��#�j� �y�eS�z�xї��Yx��qs^.�y҃���`w�:TQXU×FB�yb�&
h��7�L�44
D��#ϟ�y�ˎ��L���!(����$ʂ��yҫ�,q��, 5B�<�Z(�d�'�yB��>�捰��,[el��b+���y2_|#��;��E���$���7�y���P�4�` ��`x	jq���y�o�e���P#�_�"]��mQ��yB�6�.e0�b6,fְ�P�B;�yB���GI`�h�3+���fn��yB�Paޙ���M,ne��+�'�� �%���Q*��-c��p"
�'�H���ҬD6�A�2G��d�x	�'M���Q%d� ,���oz�]H�'�T�w��IU\�1�]l����'llu@���ܪMb�14�
�'�ڕ�CAI���x�Q��n���
�'׼{�%-Co�X���ߪr��tR�'���!D�GfHes���f���
�'th|Ya�^4]��P��OD-0����
�'Z�i�!��:`����R�2��u�	�'���Y��-%$v�� ��.�
���'b�hrˊ�M��LFs�v���'���SǤ�6\�Z� J�v�<(��'oZ�1T�~S�!ڵƛ6=�r���'*��QjQe��չ��< $�!�'��E҅&�HL�<p���$D�N��'l�Y��a�":�F��� 7��m���� :Lj�k
-N���FBeڡ��"O����ӊ ��Z��ZVxer"O~�7#}�n ����;N���"O*h��R��s�F
+  ĉ�"OD�pĄ�d6 djQƶq#�as2"O���eDR�R�`��%�`���*Op)��c�Љ2BEتwB�1r�'h�� ZZ����o�\��'��$�P��5�i�1Y���z�'*�x�X=�,	���
�n<r�'ZM�@Ok5� )�#w	n, �'��x��HR�9+�q
�s�'h�eyvF�@[��{���b*8��'3�����B��I�E�ġTn����'�2!0w@a��R.F�b�����'�l	�N����U�R%ĝhF���'��d�2fF$���r�<8�4��'��I���>����AH��.f�{�'zRH+ah�><M���c�.٠l��'���xo˗ �:�3���1^��j�'*r���A�x�Y���L�x�B�Z�'�Ҩ�Ǌ�9����a�	�u�@��'s=;���pA^[q��g��yy�'�Ȕ�6E<2���0	�fk�'�a�K�#AY��(��݂`Z����'L�p��KZ��Ga�"J
�'?����"��I�d`
�@���'?,����n�Ȫ��ͣ���'D!5bP���m��^�nDc�'h9���UB�-9V'�q�i1	�'`z�:wf�#d��O3p����'.v�z�B�.w���C��ry�#�'b ��nN�(�����W0:Bz��'�t���	9h���@�"D<< ��'^��k�8=w�Ȣ� 1�Du��'V�l�6%6-�8y�'��7,`J�'�)㠣�:�`�i�� ��%K�'�p-�`Cԗ7Ժ�[t��4�z<	�';�)�E枿��zC�فs�ā	�'U�A��8XB9�.W!!�<�p�'���j0�	/3��[�F
&�@�Z	�'�I�ː��*;2`Ѓ| f���'�$����=�z`SA�N�r���*�'�Pe�%{Ġ��W�	�'-b�'����QŎ�W��X�'��<H�I
�a�@@���I��0��',�YF�>��D9��=n01�'>����=�J}���� ;*��'�q{���\�(��	J�/�����'�f��:N�\ju&���}��'�zѴo;V���1��]cvq��'>T�w�K�b�� R �dlK�'�^I��̍�����diܔbR0��
�'8$ě��ͩbd~��k�$Q�<�
�'E��pݮ	+O:�^(st�%D��0����T\r|`��'f�H��'D�4X'fO��8���>M_*8�D�0D�Dq��4A�D13,�2((9�L0D�`�7��	�^���.^9,�	��-D���� ��U�ܜ{��^x�2�&+D�좁��~1�@�*Y����(D����AܜbĖ�ñ
� v�İ�#(D���C��$���% ��L<�Qf!D���M�!7sBE�d��S�N�w!�� ���IZ�S��`�(�"O�-�s"�]ǲ=*�CDz���*�"O��p@�B!F�"1rPC\�{L$�1"OĺCa-�~���B� l���"O����/�=;��v�Aq�h �"O�̃aO� �Dq3,܇n��,aR"OL)XF��1L�ڬ�0��9}y&K�"O<[�↿9����%�ݦi�ܛ"O�h�o@�)��saF�,����"OXx!���L���F4�\x��"Oh`6��]�D�p��{|M{�"O���6�Z;DDp쑠�rFi��"O ��rf�.�����!�-1�d�w"O�M�n_2���%�4a���"O�t�K���^9���Q�{T@�"Ov�
�W�zw�H�Ǆ�A^b�Q"O\����X�AX��fG�3zL�g"O���RNY�v-"��C�_���� 1"O\������DҘ�̖m�B��"O���0��Uʑ�5����]��"O��Z�ʌ;>¬Q��3�����|��'ݪ!0���&>�(C�I�"Y��	�'7�CCͳkj��H��T���'Hb��4Ãw��*�KϽn2���
�'�8ʱ·Z[j�ȷ�ƥQQN��
�'I�5�&B pH����ܾ]:n�
�'��9���t^09qWk��%d|t 
�'�����ɇ�,���I��
�3X�u����'�2���, x]����ao�qH
�'�Ru8���3�����ρ!F�Hk	�'߈� �@G\�8����z.j0k
�'ж��B�D����Tʋ A�L�	�'�.5��� 5����6�L#:�hЫ�'� q��Su�� �hX3Y*��'#���c��=
b�8"�܏+�.�!*ON���m��T葎_&�a��f�#;!�Dܘf�r|@�'�H��E;+�!�1o+�8���ļp�Q�cJ#QI!�@�y����5/:�ib�	L�!��JRd�sɕ�T,:]�]��!�K�,�:���+]6���!G�J�!�d
��,�0�b� Hߴ�V���!�d ��[qB��g��
�UM~!�Ė1��i�p��3��CJ�>_!�Z q�LQ�I�'/s������R!���v�)��GޭT��!gI��]�!���>���	��$[d6t�5�.3w!�
�}�v]�B,��oa�쐶�I�+I�y��I�?p�a�+I�5��`�TL��v8:˓�0?a��@���䁌fh����n�<��W5S��`ô(�0�s�<)ï�;`�t�P��Ǌ��u#�C�<�w�� u;V���cF^����A�<��G�iM<�"͋<@� x1��x�<1�n7�� v&��S�)�$�_�<��H�&�� ��͝n����iS�<�!�й�%/�7�F��r%�Z�<Y�	ӭ�F<��.ҙ�z- �l�Z�<Q
�B�Z���j�$d蝘aKQ�<�t�P�*�5���@�u�P��R��I�<���!<0����]�B��e����}�<�e�B���5��^�%�ڈb��	ҟxD{�����F�DIAY��HP@\�[(�E0�"O�LP7���RPcPN�<[ʕJT"O� @�i��R��馍�;:�r���"O���ő|H4����+g�~�#�"OB9QaQ�bw�`K�`
�$�$�"OR\�$&D�U7�sM�?���Sq"O|
 ��>҄u�뗯�TM@��'ў"~���fC�] ŮP
f����$ ��yb
�d���xݦQ��qĂ��yR �ϴe���D;F���o���y���7S����bH��zj` ��yr���E�lq*Ai�/��݉��H��y�'��^���ص��%|-�0�e/�yre�&y��Z�^
K��Q� ����yri��)��"���0���4���yң�,��(�k�-->�j�
��y�ö��<���ZD������y��S�_�t=3�k�>=�$���mK9�y���&����!SR�J�GN�y�KA�pY���H���޼q���yR��=[o���ƀ,�潀�T�hOp��Dc�̵�P%@JxqOƔ9!!���v<)��Ku��u �T�-!�$F�O�i�N~�.��Ƒ!�$�:2�3�Á�B�N����*!�D�'̂0
�` �%�|�p�&���!�hT�dyV�?8���R��B�~!�D�56��A ^�Z��-q%�� !� 7ՀT�Ug[��xI31��8t�!�ʑk�.����>`�-+�c�^�!��P�@��/H� 0;S��'R�!�$����ϋb	�A!2��>��|�P"ONp�D�Yl^��0-��d%
a"O�8j�B�*�9��é!ʨ�2�O<�(f�Ub���c��c�hr "�<����)05�p��zc�I����:f��B�	�FY��'i[�)�<��" Q^tB�I�qЮm�e��9�d݋qO^�~�<B�	)Jf�(2*��+��,��
�')�hC�	�4i��QC:y�,�1RLۘRC��f�t�rK�	�
�C��3c0C�
 Ԉ��7ƒ�1,� ˀ
đI����g��8� �5�` "��
������-D�d��KV�[�͖60ti�"J7D����lJ�~ب�%Ӿ(`]��(D�<0Q��T!<̃�O�.EkV���$D��$9c�x����$� y�5D D�8"t�I8<Q�&�M�d_�lH�n!D�[C�܅"�<L
4�E3C��(R�!D��2ЮY�*U{C#Ft�*�Р�9D�����	4r���a�� "�X��8D����GP�Q���JpMφA<�1�c"7D���1��#U��C!�K�#�� 0a3D�T��ÿQ�* ��+Id��PW�/D���&Ĭt�h!j�&?+�4���n-D�DA�ǳ/f� ��E�[-��j�O�=E���ٱ��l0`���	,���5(��=��Ie�� ��a����I+�c	#	Q*ؑ�1D���c����iCE%�8Pй)��0D��2�D�#�"]��<tِ)�2�+D��&���h���\�)j��q@&$D�б�	�fB�F�ڵ!��QF?D�x���Z?D�0B�[([�Z�#��)D�"Q&ǄU�f|�c��=*\�R�!D��ȰA:8��;3i�>��l`�=D�!"B�=<h:6%�#�N����?D�� � 'B�lZ �7�*1�c"O2���fF��n���"��"O>�"�Ù+�D=P���䨐92OJ��$��	���D�Т[w���'H#D�\jt�W�{l��F�M� R ��$�!D��1BX�����8�	�p�*D�@cԂ�"A�X;�6d�M)��,D���4�TULh1
%�����e�7D�H��!N��Ł�lR�v�R�5D�@�#��p��t9�#��yj�
�2�����@icwg�0Jf��`-�Rݺ���3LON���~ЭЁ��s��	�"OZ��W�ݧd�D� a���Vʴ�$"OV��Ff��m�� A�Q&lQ��+e"O��*0h��+�j$p�,F�8ā��"O�]a���i.LB��V�
`(�"Ob��4B��J�D�k��,j����'�� ��&<E�ި�'�0~Ė�9A�)D�|�gơi/z��jͬ*n]xpi(D�\A��ɝ)�ݳ�oI�BLq(��'D�4 r�ޅt\�щ��3DF--!��*�FiAg��<�����KֹK�!�$���R 9�	
$?<�R���K�!�$Cz�Yh�0�B�9-ܙ� �	V�O��Di!N��1�ty a���A(�M�����hO�')��ԛ���=G�ʉ�7ƅD F��ȓo���BN�SfE�e!�!9�Q�ȓ��񚤍ɬU� �(� �K���ȓW��pc4��	U�h�@����uv�y����"@
��q�T�c�z9��i�K�<�c�$W�L�׃��@x��_Eh<��aӵ��`"���.�Ň��y�����+4K�<�L�g�/�y��ޯH审�d&�7یMʦ�C-�ybD�,������0VB��Ƌ���yB�A���z�f��]����B�ӕ�y��P`m�����jg�A2j��y�AڠR�г���]:�1���Ө�y2�]�pJ�`��.��?�B�h��\��hO@�����}��(�O�*E�-+v�:�!�A�L��-yUI�gȌ��X�O!�$��j�yvIK6XZ�b'�\5^!�DQ*|3���$��Q~Q�̎sV!򄀓R�l,bӢ�d3�m��Rj�!�d�=1@�!q&�D��	@ˎO!�R0;��R����v�D9`�ErP�0$�"~�P@WN,b(��%�N2�P�\�y�*T�|�zEYD��	�.��y"��d���s�m���0���&��y��B�d^����³L� ��Q�Ǳ�yR`Ӱ/\��w�]�I� ,�D��Py�!�D�襢�R$'���Nl�<��I�4:Z����̤N.�ٸ����<�����(��GȈi�B�'��(ڲ,��-���Z��L�'6)�d�i����ȓ'z�u)Q��TI���J�*(��VO�;��W)mN>0&f�$�E�ȓD�:��'�wD9x�"#zrt��u�Tm���y���t/C�A?��ʓ<���� ��xh�JHN�hC�	�yb�a��d�"Pæ�yң�[Rf�D?�L[�/	-ml�|���,+(PڕM8D���A�E�����^�O>Z���K5D��r�2L��DP�I]S�2�I�h1D�� ������z�} R͙7!	�Ps"Ot�ccl��5�H�0�U9~��H)�"OH$�%��N�\y禔#G\���"O�b��ˑ,Q��À�C�-;�E� "O�m����;,��a�Fٌ
 Z��""O�4�u��Hǔ�єC��(�n]��Y>�X�'�E��U��,Ñ"����:D���$���|��y1O��]수 6D��Xw�=c��5�"gH2g�l][��3D�dHX�'2�t 4C�q	`��2a2D�8r����{1nQi�Z��QȖ�2D�\���[�P9,ت#�=/t��/D�h��aA�s�p��'+�s|�Ѫ1D����
�+AA5�7��3]�*���g.D�(��B4[ tJ��!#wd�)��+D�쩑I�,�x���j܌Y�<�r�)D�����R�>k��e��W� C��(�$9�O�Q��IP�K�}�tJbS�@z�@$D�D!U�u.�cO�T�؀��'D�P1B��q��eC��>|�Ԫ�,9D���ƍV%β⢯� j��8�,D�XP#��6N�4��[��Q��@4�y���6:쀀��¨cP�a����y��!Kb@��� T,�ɠ����y�IA�u��i�j�G��!� �+�yB�_(�ޡ����<���
���;�y�'j�v�+ �/����e���y�K��2����T�O1y����O���y�̭ل��2��H�D�b��yb/^�YdU�Z�F�P�1Gԩ�y����)Y���s��A0�๧AL%�yr��t��t�1/ۉ=U�5 ո�y�ג^����.rft+%��y��,"�@��R��e!ϖ�y�J3:T��ׅ�Q��TF�¹�y�`H�'�y{Չ�P��P�n�(�yb��.)�]�wD����5��� 8��>��OR0[geǤy���hßT��VR��'�ɧ(�B=��J���3%l٦v)<-Y�"OXU
�m�:8�0E,�;6]0"O�,�b�� R>�@t�G�P�fMj�Or���\�Jb�1n�%L~�Cd2D��# %Z�,�&t����r��l�Eb.D�pC&(�8o�2!�7�p=���f7|O>b���Wc��l��l�(+�hy��4D� �1#�@�~�`1d�	X�*�
�C(D�H!䝗���@ ��@��{�G%D����J[(	�,@��^�d�} צ"<O�ʓ����Hl~���C���JQȲv�!��¤4�0hY�dG�h$!�kڼA�!�$��]ib%���N%cJl�0k�6J�!�Z/|;d���ׯD7�mblĜ�!�
�UB�h��_�3���p�!�dS6��TY�D�97�d��!n�!�$�'���c#�)o�,@�s*C�P�ў�F�Ԏ�F�(�C���/x����&��8t'!�G�n��閔I����ҽi"!����-S4��C*̔+��˄�Z5!� ])�ia��O�R���d>^P��'�z}�� Q=��iI*êe��11�'ff8"��ݍ)�xi���Nk���'Ⱥd I070@PE��?{+��я�d5����H6C`"<�1�-��Q8� D�T��!
�$�:5;�֗Z��2�0D�� X�ɀX4\Z�ȗ`L,'Xh�C��'Z1O���F� m�H��[8T.^�i��';�I;Bب@���,(J��$���@C�	1 �<b".MVԅ�E�^� �C�	��|H%*�$+�H+�����B�>J�F��q�
� ~��w}��C�I�z��TAL;1�ԉ��V qԮC�	p��=p5�'t�|V�G�RM�v"O�@��뛹~���J������RR�\��	<{0N��p��L=fHK�K�pB�	�%��U��@�+(.<{Wl�+ݖB�5p���VĞ/�� kHmXB䉭^f8��$��Ԍ-�EH��(B�ɬ;thc��ݭo�YC��ǚg�XB�Ij� Ua�e���j�[E����%ru�a�0/U T�k��� ��u��Iv�dpx�h3�F�N`X�gKJ}�Xh�ȓ#ʎYq���>��Y�e��g����4��d�,3.@�D`�92]�T(�'��A��hY=f����Ȝs[��s�'AF���H~�\�)@C�=r�M8�'���*��P3a��`"d�1&R	ߓ��'���P�A�-^H8H�F����pܛ�'�Ru�u�U9lfYK�o������'6�N�:uP|�C ;i�x�(ߓȘ'I���(Ҿ0Z�=;'	�8���2�'�0�vb��0���'�=B�՘�']N��4$6S�V���*G	3U�<�
�'��U��gӓl��hx���w�-�	�'����	 @�v�� �����'���S(ؠY,�DV�q�~�:�'�6m�&]��	�K܍c�2X���y��
0'D��8T`�9@;��X��N+���0>�S�O�5
N4A�ͦM8�*d�X�<����)z$�'
A"	vq�U�V�<��ևc�Ųu�ŝOں,[3�VIx���'�|�;��܉>�ֵ+��%,~x��'��)KΌ�MH\<8�"�4� d��'�qR��_8'#���a5\֌�'���qMƭw��� J�����'0�q``eYTF�qB@O�_�h���'E ``�`Z�R�戠���Y���
�'���T�(u�}a�nAN�,�b
ϓ�O��aG�U�%�,0�H89�,�"O�9�e ��P�i���2�����"Od��Lę>fJ!kd,^	f4���d"O|	"k�4�
a�C�ܮy2��K�"O�|C�O�F�Y�u��1*��;�"OHQ���կsWּ	SG
E�i3�"OF��қn����&ƕq�"O��r�/�)����0�
 ��c�"O֍YuFK�G���L@�ڤ ��"Oj0s`��i��*_(n�l0AOn�!��|�|%@׌Հ4F%�D'D����Y��f�n��l<\��@K�<��nQyUś��Ap,�2�ǍI�<	�mµ'O�a��+�-�XQ�፟D�<�䃄�<C�ˆk=���1uy�)§=����0��z� ����U���)�'?�u��,\�.��U
}�4�3�'+���b��3Z���[Q� �qT����'��%Cv�DPz�#CM�U�����'��ܱS��ڊy�!a CҢ��ʓWF� ��Вi��D�^˦�F��3� ����?��2��>����'��	�T� ��堜0p ���]�RB�ɸ!����N�9[���XD�;oPB�ɐ8o�IP�LE�0F��!F�T�.gB�=��?q���U$$�eꍍq��9iv��_~!�dr5����+P�jI��zq
-l@!�?ܘ*���/��%��&!���5��]2ŉXteB���8�!�ȰA?�ڵ��pR`��'E�l�!�$:� ,��� @NV\�w��A2!��:I�0�Ca��v�eZY�Jm��'	��#&l��2�b��.�g��P�'�BDk��ؾ6���(g(�t
�' J���o�n�f�p�^&`�4E�	�'kx,ĥ�7ͺLHG��VD�	�ܘ'�FU�GbE3ks�UZ���?&H��'qH HVdW6d���
� ����D �'�`�;G�ŏ!�U�P�.7��@	�'��=ʤ�D�_�6�����$�6eH�'B<�g
�{��j��N�c��ԇȓy?��IwĜ&x6Q*�ŁW�����2o 	i�eO%u��{Gŋ	2Lq�ȓt�S��մj>�]��"����'�ў�|"�FթU��h��Ί�
���sh�|�<Y��X�h
 ���J��|��*
N�'qa�$䕘1�fiJ�+4ɦ�	U��-�y�O�f=�x�E�.~<`ᴪ͎�y����-�<`� �+ي�ł��hO��.�#�$1 %��87[`��V���*@��ȓ����вmL����j޴B�Z0��=��x"�)�3"�b�:W(�*�����s�j��fF�v3X�J#�A�8z�8'�PF{�����*ɔd�E3:2)Rb	���yҎT�����!A)5��
ra�%�y�O `!���c��{�LQ��!ӏ�y�� N�yC��)2|T�!	����+�S�O7�9'��&f���Yg�һ<�<)�ϓ�O��A�
�&ǯ��4=���|b�'�\0ʥ�E�V��+%�PI
PN>�L>���$�	J&6ai`FX:n�6My��{jC�	(l� Y�R�ݝX�|Pq�_(E�PC�I8�|�e�\�Gd*0H���W�LC�I�;\��q¨�t
^���D�_g(C�I�V��d�&� \�P��<�C�	{Dt� �[��݂'��{�B�I�X�:�h�,Ȕ]��0�@<%��B�	�(ޤL�ֿm��`c�J�RC�	�I��`S!M*'��
�.{A�B��@�H�I�'>|Ჽb�/ߪ��C�I�
�t��<j�� �(�kcVC�I�R�~��G&N�9�|�s7 �$7�C�>}ˢ�� [Z�*��ϿP���$/?�'I4̖�c!�
<"��y@$�Z�<�FKg�NT��j�=E���*�Ȋj�<���
�d *�b���2B8
G��M�<ђ̀�yD�&����j0'\`�<Ya�'kn����"b;(����؟���V��?����N�<A��dVf��Љ��/]Q^ey
�'�>h�&��.b蔒�ƴdL��H
�'9�����>�3ł"^����'[�S�,G� �D�k4�ؠX��`��'��0W�<��A�dH��C`̵)�'U�H�f&\�B蚴�H�Q����'����7�N�@��௄�Oe���N>�K>�,O"b>� <�p)@J�}8f�K� �Fа�"O��W'vm�1o�ThUJ "OX�H��k��H��?LK�� q�'��� ��!�,u;��9��B�1D��0���jz%���d��D�,D�xZ�#H.<m�N�e�O�B�I���1���
�ڜ2T̒�E�>�?1��?��4�V�gͦ����$)��,*�f
1�y��Ӓ*9v�{v�J-�f�����yR+�)el����΂Q���yD)[���'�ў�O��H���S�1����F��Q�''�dCD��Skdy����aޤ�
�'pQ���>)��ģc��J��=P�'P��(�5��H d/)Y�ĳ�'\� �h(6� �����RՂ�X��x�,ӽE��J'��{� m������y������� 
s|��^{�<av$؊6��АLܶ?��(2\_�<Y�KF/A��W��wQ��q�[_�<��
>X����W0	�J�ҁkLt�<1�I�(b�\ ��,-mm�"b�g�<y�h� ��]�j�o@� b7ɚY�<Y&Ƃ)&$�cV�_ d�@#�-�Y�<�KW(~���G�[�B����Y�<�o�#Z-"�.�1&L���Q_�<є*�0P�5���)E�}yB��W�<�ύ''���*Ϙ��.o�<��Z_%^@P���6�	�LTF�<q�-џ����`�TTL*a��V�<A"��u�����)^�7~��a�@^S�<i�ɇ:e\>A ��A�[�`��B�x�<a&�2�n��2'�ak$�'YH�<���	I<t��B3��S�^�<�#� M�BeFJ3[���C�	L]�<��g��'��-9���-
��|��B�R�<)��'?8�[vnN53��xkT �J��a���O���)85�"����9dQ�4K	�'7jM��@�<[�z��u@��\��`C��d O�X(���F�}j�*[�.���"O�����U4F��(�H��v�#�"O�qj��ջQ ��b�g�
�D�p"O^H��
@�.'����Lu8 �6"O�,��R~��R'O��9�d*LO���lE�2v����d�,iO�9#�"O��/H	4�|�2ԅ�.e�� "Oн�&f�V�`�j�0Y���A"O����P�d8a#�+�1~9%�"OH��h��YY��%\ �"OdP�]�n���Ģա
��W"O�Lb�.��4 �)�D�܃	���D"O�cI�3C�:Y��*�dȬ���"O��"^]�4 �JLS�ȹ�b"O>��/�-S�f��4I�+N؜�+�"O�I�"�CV��m`bA�"OB-�G�D l�!��J�h�"OZ��a�Q�A�<���m�	��݀�"O��붌0s�$0�g��7j�Z��"OJ@q�R
/T&ģ��uJrT�DD{��)N�i;f���g��ԵB��-H!���.�����:P$8��	�d(!�D��jJn�2��f�4��a��V�!�$
�#@���͛w���I�ǘ4F!��
e��u�qF�#�PԂAf��:B!�$B�U������)��H����[.!�� �)�W�+pYx!��6A��a"O�A��G��?��$�f��%=@1�"O�3��K����SE̴9
	3"OJ}�!nBm:��{���F�*D��È>�Г�$Ǫ��=K�(D�誡�R�[�	�����A���%D�|2!X#N��1t�K8'ɲ� #�d"�S�'xX�*Ѧ�e9��t@��v<9h�.P�h�X��;`�*�8T��@!
�6��h 䛔Q5C�f9D�HZ �A�=̖�0���'C��2��,D�d����U�<� �L� Yx`%+D�`�U�4.�$|Y��޹���B*D�(5O�Z�̨�cX�M�eZ�E)D��� ��"�`�u�Y%
q��(�&(D���,(��<��*
e��T`&ͺ�y"��Ȝ�2�m�g�$U�����y�n�%Yre�f��Y���t�4�y"JF(�0�Z5Q�[��(���y�k��7�D��D_�M�
T;�	�y���5w-Z$x���F�\(0S*�y�C�WK�y��f�>8�%�w�����O��=�}RAM�r)�}Xg�]&Q��HA�����II���O�����'i���PG�(=F�a�b"OL�jҩ���4��WK�a;
иS"O4�3���L}V���:0�y��"Oa��o�/t��ɫ��1r�֕	"O�.؄(C��� �:J�<�`�"Of�B���E|�P��O����(�"ON�9A��,,�d�� H�/S�1q�"O��
��Z r[x@vS��Q�"O�dɳ�Ƃ6��B���l��2"O��ƈ��n��Q���bq�&"O�6��l7���TfKD!6��g,D�~"�+T���jI��ɖ.�	A|T��d/?QC$��+ﮡ�Eԍq�;��B�<)2�Ԏ@2@�3u��	+��mW�UA�<�؃�,Y�n�/[�H���{�<���?_�8X��'�}%��X�FO�<����3`Ĺ�u��H�x��UH�<q ̘�>���(޼�l<�w��Z�<!�����ժ�I��=�.����B�<a���:{������R���%C{���0=�B�ы�$U�l��P�&�q�<�f�04�9�rd�^|2yi�V�<qDH]8xF:�7e>#~ܢׁ�O�<	WO�(X�9>'�dbPL�<�!j�(��)�,@4Y"����K�<�&UaӾ���BŚ&t���.Jh<��&|s6�SG�\�9�l����Dpm!�D7}�}�w�B�X���x�	�Tў��S�]G�y+��
�|����L�b��C�I�Qs2����[#>Q���r�K�xChB�ɱmyn����� ^��ɕ�\�:y�B�I�)m�� ��P�i݆|S���4v�C�ɠ~��d!> [�LA��J-:5�C�Iw'B�3�"C ��;���(XB�ɨj�4��FI�7���p�mƽd��B��=1�D�#��`E�s�B�s��B�I�/��r��Ю4��;6���FB�ɧ:���C�a�I�*��7\@B�I�]$�T�dƏ�f�C�凜
�B�I)мa�nԶ9 TR��B�10B�I9{�}��9N��3B��B�)� �ɓ#�bɜ��fY�\�.1����O\��$�"�v�BCƯM��I��P�#�!�$
��2)a���<I�t���4=!���9 Z�*0i��-؈D1�<b�!��3B���c�.�^�Qb��K:6�!�W/Z*T�:��N{=H]���?�!���&FTB/I6|0h��s�*=!�	?��ܢ�d u�nL+�%V�$,�'�ў��<i�cC �����i��߆P�!�d�(.���Q��L�fM�Xb4$��(�!�ĔM�f��p�ɿ0�D5� �ھNW!��3J��!��zè9Pv)��"�!��Q"AE�U2E�N�P���C�b̹�!�$�6EZ�$YC��0Oa�9�AG]�!���'��J��R�y5�,��"^�Z��O����!SE�ٴ� �|�:�f�G�!�dL�<a~��։9Rv��02�T�6�!���h�	���Ɲ s���b$�5}�!���-�lU�����Gp��1� H�!�S @�x"S'��W�رka�:YR!�$Zq
�8	FFF2w�riA 
ډQ@!�# J����[�;JX��qG��!�%�z<���a�dXE��q�!������ڲ�I�U�Q[g� y{!�Ⱥ~�6����H�T�y�ФE�!��!�1�g�B�@��Sb�w�!�d 5q$��i�����b-AwźR!�1V�*��嬊6g�r-밥��:!���r���
�l�tY��nI�]�O8��� f�Q;C��@�����I[!�D��/�V�ڡψY��T G��s�!��� ��򎃣	s��5��
�!�Qb�8
k�T�1�T�%�!�̖Hk�1�e���}Z��В+��T0!�K�t0���bO�DdJ �1%��|�!�$؆S��i��_�(P���Bc�{�!�T����f��*)9���r!�*G�!�D�mT�\�4͙<!1BH��:�!�$���a�A%ɳ$����44�!��܇W��H�1o3 �4	�ֺ}#!��	!�p#4'��Fp����)�}2Y��(��@�w�e˳&�U\xB���~�<� � ʪ0Igc� r%F<�T}���0=if)��:Ҟ��$���M"����a�<ie@�n��YX�ٰb�dy�č�T�<�T✰ݬu�#��2�Zy�RLM�<YSË}�Nȩ����h���Ks#�r�<Y[�Ƭ� �	�N�I�B׷P��B����4�E�H�Z�5�SE}�B�I<B�0},M^"S��b�ɛ�j�!�M�5�)j��� r����L�8u!�$׉@~�1�T>g�!��͚�Nt!�5R��)�pH@�h�taWc� X!��AF�Z��ѽxD�;�h��!����I����|^�0rK�Rp!�$U�`R��BZ�lh�L�3�!�A�|�X`&��
|<Z��'e�J�!�$ɪ����E�6Ǽh���sQ!�$���f U�a�n�{��(!��{	�Ѳ���N�>ʒ�.!��B4l��QA�-ՊTxL�u ڹ]!�$��On�#eF(xXbѓ�@@�!��]�;��)�O�svBCC�L�!���;\�1�w�� b� ���N�!�� M���H�cSXh���sl�d#"O���P)%�V�#��CNRj`��"O)K ��?�r�8sD��p���U"Ol��0��(�С�A���K`�0Q"O�ܺ6㏦Fܢ�#�'YN� �d"O����R/
-,�� �:򔰋4"O*d�m�V#��p� �t�ܐ�"O� �"�
].*<�sFΤS%h�:r"O�EජM�*r��-��K6��{�<�&��>x�P0jS��zzpP�S{�<Q�K��z`LH)P�:��t1W��Q�<�"O��lkF�[:db�'9:��	�'��%���U�S/���cZ-�=�	�'�����E�S��� &. `���'�H3�僣X��Q"�!�A�B�#�'�`�c���{B\u	VX�,��8��'��k�J�]�����&���'ڄ�B�F�X9��'�#� �I�'��a#�
"w�h�S� �����'��h8�� �6Ն���Ħ#��Ź�'���X�Mʦ$1��� q�r�'h�-h�D^������ؿU�=P�'��]��m׽:�6���ED�^�<�'>�M��E	 (�@� Q��(�Z��'�TT�W&P���(b�m �j��R�'� ��a�>��CG8,6�AK�''\0� �9⣒6����'���!��Cx�QA*ݛW�Y�'I��c`JHH}�x�nǞ��1	�'��@�iC�<T�밃M	0�C	�'oqK���6[�hS��X7�t�H�'���Aɑ9>�-�����Y�'�$��������;��P�����'�8S�$�O���{����uBxJ�'G�m�j� ��ޯ8�`���'m>h1Cb޽K/DуQ�ߨEX����'`���Ŕ/i"�	��E��u���'[�� ���+t�A��qBxղ�'tI4
		:��5�d+тe%�p �')�P�1��<�6���d;\`�'��rC��8|^B��E/_}�Ȼ�'C蝱�+T���`�B#m�X3�'�� A4l��8=Q*@㘣]a����'`�F�=����$���X�he��'���(/4ej���"^�d<��'ER� �聬$��\Ti�YK�])�'z4�p��/�P5�s�s��ail�<!�!t���&D�>NB� �)�!�ą=/ ����[�FVL���4�!��T*��Q��\)N8lar/��>o!򄌵H����+͈1D|�3^!��W:m����.Z�C�d$3q�R�!򄏽i��S@2I��Bnœlz!�$W8{�pia�ܨe��"��_!�đ�^�m"7gEX�D8���6g�!�Hq�Y�Ǭ�T�~�K���`<��_/��q5 �w�FL�a]R�Z݆�4��� ��7X�F���Ǔa��Ɇ�J�H��IN�^�Y�c韑^J�@��J��4�/הZ� d�j_�L�ȓ@ሀY7�%D��B��Dfx��ȓ3�M��N^�	Z|���Z ,���c��)���<sz��$al`dP�ȓ@�Z���Gƫ\�^uYo��nyn��S�? �� !���\J��K���S��pAc"Ox���\���Ӡ�3D2"O2jӊ6J�z�-I�m��z�"O^}+lN?'R��W��'�����"OYC����e�<-�*2����"OD%�e�P7yɚy��AF�uvd`�0"Oh��4(F~�$l�FbDko�P�"O��y��\�a�F��ժڤv^�D �"O�eS#�#%���ag)N[qX�+�"O�Ф��
��\bozϽ3���ȓo$�fDܚs��UǈU�ȓ�v0�rKR�M�x���ˊg, ��m�6E!a�60���b�8��{�R�w6rj��@M�����ȓ:�.PP��E��x'V}�����x�|@��ݶr������ i�Zфȓ=T��UӼ^�|P�4�#M**!�ȓ9���E��G�XI˗�Yl,5��/Q>��v<%;���Y�>`��d��8 Eo�3@B�r �	�(=��ȓl�|�:�fҴ$c^,a�M��0��8�ȓf�hA��&.��ࠗ�S�a�5��j�$"�H#Cv�� �۱B�$���V�Z�pc�$0�p�n/!=и��ul���(fSt9��G�v6�ȓu� ��M�8]d���a��/�ha��.�p9(v��)w���`��Z�ZQ��6�F���L����$�]:RȒ��ȓC<��ψ$'��8�כgB��ȓthv�[ BϒS� ���l��W�H �ȓZ0�A�D��p3�-�-3�6��UZ��&MH
{( ��*R�L�؇ȓ"T�$!D@	�7v���IY/A^x���?\CVEM�38(�Bq�E�[N����,zr�BӤ��j/p���V�G�B�	6h�u�o��V ��D�f�hC�,2����ɉ+�r��G�-#(�C�ɱE�@R�����Kf����C�I�E��°	[�C�E���L�w��B�I�����!GN3��-��ㄓU�vC�I�g������({?2� F���C�IHa��
צ��2�B��0�
#EV�C�əI��T����0����;�C�ɷn��Lj�R� �:��ڒ8QjB䉃[�,L�d�9G6��'K��ZB�I�`�(Т.Y.'�=p��X;rC�ɼw��b2D��Sq�:b��B䉀Y����e�I��̉�v��B�	@"���S	|nXɃ`ϸs��B䉙�	p!I�UN�Q�����B䉄 Ր3B�|d8��w#\ʤB䉛;dz��ć�Gd2gi�_�zB�I�k�<��	مp�8l �ؓ]�4C�	�l�KWJ��D-@��1=^!�d�(��4n"1���1��\Z!�D�8w7Z��q�¹�e0���d=!�((���c�0,�B�A�U,�Py��SbD�U�gθ�%L���y2�0xJJyy���*/����&ڥ�y� ��k@ ��A8O��y�L3�yr@�]n(��?2�(��'���yR'E0��M���-ب��DMց�yR��1Lr�zfaY���q���V��y"���� 3gm�	�\��-��y
� ���d��uѺ�2aK� ^�	�E"O��UfR+@L�x���;n��"Ox$qOJxp*F��[d|�Zb"OH�1Q�فm���`Ѩ]�j��e"O�ۢJ�qArEA�EH�`���"OBd�WEV�����E��Z�P"O��B%�ŇT'�9�$�����"OB�1��ĈM�&��p�M��`��"O޽�����{<Դj'ヂe�]��'���'�<ӓ/��N��J�U�xx�	�'�>Р �j�d`Yf�ՓnK�5*�����D�da̛{ZRLY��-�H�Ɔ�%�y���F'8��$�)O9��Qբ��M��#�S��M���N�",<��"��e^��	�f�C�<I�X+;��9Y���Xǒ�	Q�D�<	�'��|�ەJ��	��ڠ��tJ��_
�yb ���<�`!傔��möˆ��y2�߫y����#IS��33Lޝ��O#J�k͊V^�P$��g9�a	��^d�<Y�o�	�ܸs�!pR�с��b�<i���;�MSE�@�-N⬲r�@a�<�n_  4���S� �P� �JB��Y�<�b�0ZRea@"�b܉�	QO�<�r�����,�t[�,�fF�G�<�Djΐ1�r������h^2a�!�Z�<���ܤAi��[r�ͼy�Za���
Z�<�g�(A���#R@��`lZ�<ABG�r��Ы<( l{`dBW�<�/܍_Jh�ؒ��	#�1�SG,D��y��.y�U�ң�*T2l�b(D�(bǫN\����bI�W<Y`�&%D�`0qJƲ+��UY���`��%A�<�����%��%�$�n�[ ���lB�+_��LJ��%�>$�b�V�]TB�	�O�P�a�1j>>�Y�'Q:�\B�&�ԼB ާ�<p`��O6��C䉣f���p���;}Hd�V��/&B�I":�8R�9^����&�9>B��/m��$C�Cܸqd��'H�R#b��G{���掙C��KAYFr:��A�I��y"�C4W+%�/S�9��.
�<B�I/-�Qu�N!E��k��.,^�C䉑�d� �aR1i´��$�3z�B�-��T2�'�2<`f�g`�3m_�B�I3~��D��H����$JOp�$C�ɄVQ�*��6�q��4�,B��%�8и 	ր;�rܡ%`��B�	or���'C/o-���b�͋�b�ȅ� ��1<6@��5c׵m��C�1]x�������X�L�%N��C�o�|	�kA��C���aEvC�IzY��
�l�{t��	C�\�~B䉕t��U�D�	�n���o�hPT�'aў�?�1����$���S<?ʞ���L%D�*��E���Ye✠m��@P�a'D�����K7:nx!	�H��I�j	k �8D�̸Vm[�G`�t�u%��'�Z�xf7LO.㟤�6l9`L ��$,D�q��2D��hnWBZ�a9�
ɶ+� ��k/ғFO��ը�:�b�{��_�z�;��Z�'�ў�'KŨ��t�
���!�U�>���'gў"}�'��yJ�8�A�[~��r�W�'��x���/Q�Ѡ��HmԥsG@����� 5��>!Հ��n����ϝB�t�S��y�'XQ��S�? ���K��4m�p0�T��z 2�"O2I��(;X���l��B�)�U��}���Ƀ+wAvq����0��I/L4b� E{J|
dV|�ʡ��&@%��]�a�_�!�E/>j��G�A���8mʩ!��#<���!����
�	�@Z9�b}H�&V�[!��_:0�`�ӯ��`AfS\�Q�T��əQ�,݋��w�5�7���B�ɪ!b9�dg�
:|� e���c����и'&�'L�A�1*ߪM�`(B��� k�z��D�Y�O�x4�W#��1(�FѰò�Ҍ�DH<�a�ȧQ�x3c@�Jol����fy�X���<	��,��I^�M���|l��E���C�ɞ,��F�F2C���bG�ŽAdʓOn�b����ԎBC@J1s�J �-�� j��x2��3C躡+�:�U��R�$���d*,O�Ȃ�
I�J�Tq�J��&� ��'(���Ir��Zg!�xx~́�iB-��=�	�a�T�G���
�<��l
B�8=�=yܴ ��c��)�|*�
�Jf:Y:�(ҭ"NJ�Qp+Jq�<�"@�	�P����Q&y#P���'^d#=��	 1
�dpX{h"!{4�Ҙq�x0��D�>��8��)\�}��K�|�X�0C�	�lm�C��-O+�`@qW�:��8{9��I_}�*?��� |�X���+hO���g�%,JP���<O�I�*G�{-C!.�XC��p��'`Q�d�fލ����Z�]Sf�K��1D�l
ƙ�LCLpzp,��^�:8���$D���f��if$��w���e�.`qTn"D��Yl�c�<�8%	�B��}��B T��	Ԏ�(gbN�S� ����>A�����&deɠ�X,�����ST!�d� � $�FM����� Y��'�R��'��8��	p0(a@�
 ~�:5��K�=ђ�8�''"�
���0Ǆ���,�1Qa�4�'�6ܳ4d�R�3�JM�r
�y���MH����T�\��+�,J�f~�$���8D�`a\�v`ӴK-1S�M���2D�PP��Ӣ���y�L��
_8-��m>�d4�O����B�z�r鎆D���D�_���)�=h�q��g��?O�����1D�P"�$w��UI�H����W�0D���c��1h�S5쟩[c��ЧN/D�$�s��HVC���27�P�0�?D��#ѭB�:����/^�Lh�+D���kB>l}H�el�A#��3D�*D�x�b�<8�,Aᣧ�o��P�%@#D����������˫n��8ր D��(�j1 0c�$u �>���<�Ǔ:��8ۥ�����I$-�k`�������nZ>�D��l�;v�dq���$v�B��cd�y���?_
��2�2ɾ"?1�����R�m��Z�p���91"O �C��IuV��7g��]�"�'�1O�Y���H���pd�T�<�Z�a"O>�8�J�2;��p	�,Z5y�mP��i�ў"~nZ�;�,iD��tr؀E�]�2B�<G[jȹ���0�B��\�KEB�ɤҊ-FL�m�) �X��C�1_c�L:#M?NP�� 3�`m�7�<�������0�̤5�&� �8��V}�R�|�}
��ԣ��Cӥ��
3NEp�F�p�<�������
�|<�!x��TC�ӂ�)��(*~��*p��41%v(ʇ��aC�)� �Tq�1����N�x�V���"O����5��0˦�ҷ!��=00"O*��Bk��/p�,� �*�O����=���I/�:�(��W�`�|I��FLX��Z Z���u�ORWouf��9�Hۃ]�t�a"O��2�H���� HM0e�B,�a���+�(O�Ov.�v�J�mW�@3�fV!���x�'���3�_	x����dEa�'��]��ƃ%�$t��E�q4<��'R�)�a��1�x�P̞
9���{R�'e(���'Y�]�bU;� <+���'m �J���T��y�& .L��'#L�T��3�VY�h�. `k�'ў"~��&Ϫ����� uH�����x�<1S�R�jD@����Rb(26e^�<�c���5`T�ߴj�iKK\�<gj��[�
��ݴ.�d�q��KY�<)�ސ7�Pz��G����A2��@�<�ᧁ�O^^D�!��Y��I�JC�<�4�	��U�ʜ#�D2Ѭ�h�<Y��L�g�\AF'U/ʨ�Ȓ��Y�<��% �v��uE��h����k�<�V �^���*��'l0��R��g�<	͙2&Ci�/R;P��LY�ŀc�<��"	����s�%���t��n�a�<�7�]��zM�EÎ�x����`�<"j�y� Ps \�%��%�AŔ]�<'K�g��	�d%8�C��V�<	f��`�I���U,u������
G�<Q��Z�F<[��z`��cl�A�<Qco�u���[�fϏS�����{�<)� +�h��އ)zd���u�<�I�a�T���!f��
k�<Q�-�04�b�H�Ś7����l�<��W&5�%Qt�r�z�`t�<�Q�Xx���p���:��GF�m�<�S-^(f�x���Ȋa��<[�N�e�<��������hDN�	
Yȍ*a�V�<qP-�ak�AЅa17
�:�ǅZ�<��P*����A�@ µ �L�< �l�q�t�^ ^l��/@S�<!�*��h��ˋ�N`8���R�<y�o�"9��<!B��o��	��w�<��J�/�@L�!O�?��PKZp�<�jJ�Q�6H`�΋=����S�<fN6'��hpE�/av�3�oS�<)��՜6N�i	�J�z%��ˇJ�}*�(`"+F	EB��Y�J=�<���9�ұ�bTuΚ�B��E�<I�,C>"XH�Ȳ��=�tI���B�<�d�S>�(��F�SF�icG�|�<QG A�0��HU�G&p�.кF��|�<I�D�6&�:0g^(9��;�,{�<	U/ۢ�Ȑ eX�wKlx���\�<�u�M2rR���BN-	�⡙W�Y�<�A4�x�U��#T�D,�!��B�<��ؓ|3W�ԛ�Z�X�.f�<qt�Z�(~�	C��@�?����a_`�<	+�[z�����l��@�T�<����{]�uʀ�ҙ[H@��#M�<��&��H8Y�şaT������c�<�H btP<���˳6e�ܺp�T\�<��. -FHw/ׯ|��P��,MZ�<���.S�T�'E�+`�JҋUo�<q#m3'�tՒ�/ʡV�Lyۖ�_s�<� |��T
Q	�xi����T�&"O���I��I�T�P��j�����"O�qS��ޠ]��| �N�4c���xr"OZ1�FЅk��a
7Yl��aÖ"Oܨ��\�V�L�ڴ�F�8�4�:��'o��x%���L�a|Z	��у/��P!UK�O����D�h�j�	�����?Ѡ��!_��}B��ğ;1d1�H�r�<q�d�b��e���՛x�ĩ[��Dܓd��5��B�$Ut�����1@��f�F�(^H=��?k!�D�!"�a�d�M,2N��鱭@>Q\0r�,�$L@�̖'�LiE�,Oj]�!���|�'��l a+�"O�t�G��?�B���>Gv�@ۤ�ʗz�9�ӪźY�D��	�3�B͈� Ԏ]T�b�
�{����$W�V��}Ȳc�(o�6-��r�r�X%dt�J!����,m�!�$�=���PE�DN�S>y�qO��9!���We���Gl'ҧ\� B�(�|�{�*�o9�ЇȓF�p��G8���˰�]�L(tKV�x�@I��^�p�<y�OL�<mͣ'9W���|�<a��F<�z���^1':�a�1F�h��7N��i7�c��'�rQ�fJ�S�H?/bP��`�]0�G(���$��X�(�e�o��x��G͒R�!�$�9J��h��Z�]�e��
�O�ģwa�(r��#~J�S:*�L,3��Ҥe6�h�Ϛ}�<)2,׌P)Fi*@hR����$#�Q�<ae%|� �)�!WZ����XM�<��Ơ7��B$	ɆP� �c��K�<���@34��Ǯ�d��xq&�A�<�/	!^d��2J�"���(��T�<�� 2�.�h��mN<�h���P�<���R�wZ��Ӄ���U f�VY�<�#%�QJ�sg"ΓQ%�@�A�C�<�$�Г�̹Qa�J�t�d x�<A!튑_ar=(d�0r����p��]�<�-Ƿ^E,�c�OƲ@��Ir�R|�<��%��0T%A�&�-zHq4J�E�<�口�h���&�<�ty���Vh�<)'K��Fn�⬛�il�Cc�<0`�v�����H�z!{v�%��IN�,_
)s"�@E	�h��ȓuc����A�|kn����
H�h��IfV1 (�ntRL[2`�-�q��x�\({TNƈ(@��{f�ݤ#\���+�����MF�I�(�e�4wν�ȓR֠��5�4m��S#�5씁�ȓ��+R�J ơ;'"N
����;�dR��F5@
D�+U'؀-����ȓ�b�W�U�]˅ ƪ�]��$)9Qbk;U%\1���'l��ȓ>��]�wj[�w�"�J�@)7��t���⑚r��%6ܙ"A�O!����I�r�d !�O��D�>]�blc��%@Xt�e"O��X1NF�1���I%��8��P��$N`)}3#E��h�~b	Z:7�0m
&�hr'"O����MZ��$XF�[��U/X�iܬE��+�~Ҍ�-��bߖ� ����y�O4	�<@A�6c侴R�-�'��x���9j�D��P��7�<�E��gM�����8���RC*�^w��Y�D[�i�L�'���'$�N]�tb] �v��􍟛z�LY��	��~���m_y�@Mc��,%�����?|�t�� NN--(�",_�p��Y��`�<���͖	���KR+P�9�~����q��֠ipX� &aV�gr���b!WtH��	�������l͏1ǲ<�f��{�p�*P�޸����I�3Ġ�4��()7b����B%9������I{┺2C��	h&@�ӊ)�E�-5�|���D?d�)��ףd��G���Axeba��:�K"#`��6γy
�0A�N�H�P	A�-l��30�����d�� (z���,Oq?%��$���Lc��\�s��<X����b^џ�[�O/'�pU���	z��]a3ez�? |{���q�N�
S
�7BPqB��2A��8I��E�2���S�w:�9�~�'m�hE$WR�Y0rI)�RtA.OX]��A�&G�,�*�!�e�t)j�b>�)wd��_D�����6�"��B�T�sC*��� �*m�`SSl2LO`=��[�	zb@*fN�0�����n� -f��� '��i��x�)O���H��I��Ӝ~��Be?L�e�VgX*�����
38J|���G�<F�	���C�]H��9�)D�j"�A'���(��U�ڝe�V�ʖ�t���(X@���ؔ��4�r�eƿW�� b���r������N%[#��Q�j�����Y&\p��KX���0����0��)K�3�4��I�	wߐq�'��Ӳ��O*ܠE���ތ�"�h�v�zPZ��kc�J�,�E�u��+=z1ꇧ@�2�@�|�e�D�K" �a�)-���^?Q2�	�H�6PA��.LO:�������!Q�і{6��q��K"�8��
}�#
Dv1�e��J�Fs2��bSp"Pı�.�'��|�∉@ء��8�D0!�eZw��E�B75nA���D!X���g��\�$hk3A��[�H,�E;��|*��!^|�Ȩ��"{)�Уix�̰�o�#}5��cG�P��cH�lb�)�F�^W,AT��$:��C�$`�rA8�fB���4X�N�*�l�O�<@��Y%(�f\*&��Rn"<���T.�<5����G^��eJd��9�y2�1��h��%�v���G�_p�C��HG�>T��=��F��O@���I3W;*Q��/Y@dm�c"O�u�5��k%�0���6F.(JӸi�R�D�����|$;�)�#��`#J�3���$[�Pk朱�'��a�LȻ3�<a�SH/���c�',�t��M���!(c���J�x���'R���jƤ	ZE�bΙ08� ��'���ꆋ�t��rrDF�4ǂ �'Y`	���=ގ�H��%V�c	�'@} '�T�~*�y7�Q�b�5��'�*fJ Q��΅8dB4�&[+�?���4|�T�K>E�$�W�J��CE�)i�p��[��!�D�I ؈�4sS��B���W��	�	����R�)�y��H.m�ʕ�v�U}�b�pHɜ�p>�5,B�&t����ۍ],�s��S���<1��G<5�����B�9V\�~�L(8��SE K�׬u ���(O�Q�f�-2��c�Ҥ}ȟ��2��%VFt� a�.m�H��'�lAB%g�S�O����TK���(��G��#V܉��ݯN��(�;~�h%{��#~���0�8��� >�4qJ���T�x�	�*�p=���[9��y��ʶl��(�d�S�~��������@��4����V�'�� ٔ*�x���c �6�Ι�� Y-���R�J8�ثf�J8$��H0,��['F�X&��.�$k1&�Dص�
f����+�	�5N�ʧ<���;�L��&d�(��cHX7��GyRع8��kDL%n�� ���	_��Y; o�Vr�Ma��X�}h�럶�B�I�>E���D-p�Qb��H�O��I�B׺"�8���B�<@
` �ň��Q4��0�J�	mr!�_��~�GG�z\�}���K��x9RR�R��$k�({jTtR�j�'�(]+E�N3d�*��ǆE�q�B�g?��ޚ�ܥjA4I�x9v���i�}r@�ˌR�@��P�H��בb�I�$O�-F��ex��]4z����@�I���r��O�ٛ���d�'�c��.3�U�d��a�i1M��:Y$l��l���<a��!8\,d��'ldCU͔$k;�`��z¾�:�V/W�FA��C�}N�ťO����G����?��AM�&��6�H��`�*�H�\��d�:�h�>qpIL�DM��F�4s���*o]��/p�D�#�_}b��~l�k��'>�u���= D^13���5툩#K��J�
/Mg�{g�I�;c���hߴo����k�����!eZ�R�D��ȓc����F�f�����P2�8@F�N�$G"�|DK��L>Q�%��R��t,X*�hf�~(<�Bfá~yL�(ą�(�\jU�9�4�WG�QEX��[*�T�rp$�.�\M;� �
��x�JA���3UmPB~���a�΅:f�!�z��ǩ� �yb��0_ @`�E��5b��4��	�9	�S�[�h��K	n���~�� $��q�p�֢CS�	KF�u�<	`Ñ�`�um�Qk���� ��2�$FS�<�1���/r
 4�~�K�p�0��6Ch�a��
.,9���!4����m��5�B��Eغ{���'��:i��/��@�.)m�����'�p����c��0��+��f��%��h��풅�=3�d�C�*�E��ҡ�Y]P��F���)Id�J���=� �T���ٗM�����e[//,����;��M�ĬZ\_��Ғ���*�\���]*M$RSBO
K� 8P��c�!�䐜~c �7e$J����@Oٚ>��$9*8m�F^�x������>2L������7w�d�!�K����q��T.'@!��/�(�B�EE3���{��>D_�����C.SD$���q�����~z�C0��-X<�Qgңf-��	�5�h��DC��x�薠� m�6I�,�%/��q�,or$��I��h�"@��0=�ox���d�-ф�P�YD�' �M��&�jt��{$�/֐�(� X+kYP�F��*���`�dЎ���j�f/T��b������z�jA2V�62Bm�(���!�)���u�� �ιA-���b>�]&L��4�֋
�.�=H���f"OL���A�H8)�Pe# m�퀠M��[��PdҢQ�Rr�Y����O65�0��3M)�����
R�������4��{��;�Q�-Y�N.�Y�COT�%��%� E��x�ȱ��o^�@�k�
��W��'�'�(�b ��)�aJ�6|�����=�vl��&)��s&��o����!m��e�"�yB&Z���#R��Y��"O葉�h�w�M��$[���0��/ޘ}��\� �[}H�}��,MY�왙�(�Fܧ�y�)D�q&��㔟
��(u#���y�M �<��|*!f��v�[O���?��L�n�9 �*7lOf�@�B�Y�01�`��C��-���'��xTkX0J�n�l��D���*�ř!Cz-z�,T�&C�� Hn.B5�S�Q�\ !�Pۂ=���7��#p	�C��>����l�T� � �er�B��=D��'��:V��!�)_�g��T#�p�"�K�HXb�)��<锭ڟ@*L���$M!O�L���Q�<B� �+T�� �a��	��`�N?Q�J]�
���č�V��`�M�#����,O"!���6_�*�QW�1֌<�a��?S�!�$X�1I��So�4x�xٲ����!�D�'��Y`�i $��
�kY�!��<�-;���5
��ѡ@O2�!��R&XH���E
	��`2AMϸs�!�8zw��*��7�|X��,ɬG9!�� :��	�%
(]���䁞!�$L�,��!�d(Ɇo�P�hU�}!�W�JLb��s��/I^��Q/�(!�Ď�UJ����'K9�t�PK�$!���i��=�'�L�Q��1p�
�!�d�>���gGG��Hkf�G�s!�ˍ#E�u.�)��+S�+�'��Ż��R=T)�)�� 'B�K�'�8�pL4{Đ��K]�o��'T�� g�&"㾕��ړ�6A)�'��}�W�4J� B�5�n��'5��9�N���%X2㐊!�T��'W<�R'a�6����c׻(�����';
ǭ�9Hh�p�ϧ!�C�'��y��?lo�!c C1�VD;
�'t8�I��}��o�9���`�'�� ��_�¸�u��F��PA�'���:gj
�5��̻��K16[\���'tZ��L�8��h�U=pq�p�'Zs��F�:x�Si�0t� Y�'cz�c�� ��B����9�� �'�ld�$I�$s��Q�6-�fD�
�'�pɊ@B��]����+v���'�Ƅ�#��>���g�DQlM1�'yh\Q�E
�.��U@�����D��'�ѣ�D>C�����B��L��	�'�X�2�D"�,���%D;�I@�'�\��Q"�-�ʰ�b灹��1��'v�E�� �>���h3ŗ��|A1�'��XS�-Ɏ?` u�rM��|�:���'溸�U*O" ������āNp
��� J��bN�+D��CeG�+f>�"OD�#"��&h�<��tb�';Q�4�e"O��J��Y���{�]4MDft��"OZ�PD��n]"���`�)bM[ "O,���2XnH��ϝA��;&"Of�	�$^;xJR!�MU�5Q���"O�}xǅ��߾��#ػ#�E��"O��)b�"H0 ��+��-ƙ�f"Ob�I77�	I�I+JoD�*�'��aS��5�a|B�σ/�v�Y[��B��6䦱Pۓ;A�e��&�5h��D��(=�e{�"@>e+>��!�Fk!�ы~��h��%Z�(�G��pNqO
�C.��$�P�s�d;ҧQ|Z�(�E��,g܅�/WKN��_� e����>0^%t�7hX�(��N�$�a�#S�hi��<)��0"�
��v@��Z��iHb��J�<1tk��"��q��O�Z��ě���C��z��4:���U�'���!ɕ88�ҽ�0b��dŪדuj6�84�@._��!J�4�AY�����H1@g$�'M��]�ȓ��1��KA�;� 㩋5d̌�=�%��j^�5lY'�H��u:EBC�{�ꙸ��
aS6\xw"O>�H �R��	��;@f.�@�Ҏ�Xa�j`yB��L����%|���@�|��9���1!�$A-��
a��PX{6%#�`�ҋ�!!t��'I�u؞`@��K>J��0��K�j�,����<lOx!���$������@�)A"�3=�!�p	�!3ttȆ�l 1s�@ӷ/�9�P�]�!��P�?����"j���<F�6Y["L�3"��6��L�!�$'OeX � ���I����Y�!�D�H�`�c�'(zr�$�˥�!�$	;1l�@Pr�&3�-�0�׉\�!�pi���@+ݾ<�:��L7N�!��,\I��[@��=x
���BL�!�DZ<9��(B$R���_s!򄁸z��� �.�ib�Q���O�}L!��O�{3T���O��8A�=��Y�!��� ~�����j)n��D] w�!�d08�'dO�u�aJr,�\!�БZĲЋ�g�$rn����sC!�,ޙ��ʔ$�����gÚ!�!�䂴ulȘQu��/
�>l���6�!�dC� �Z��W�T��]k!gH"'!�D�+%���S�[�R��@'S�0+!�N[��i�E��O�Z�q�Ï!��6\�M��ǴsK�t��h]�A!�W� +|� B	[�M8v9��G�u!�B�DFU�3B8g��h��ۆ^!�$��hA�Ā�=%�d+r��E8!�dԽ�����7BW��X�*�q!�$�1�Tz��I�Ul���R��!��K#o�.�Q���`^�!��Ǵl�!���`>����.eAdz����!���,�B)"1ի	E��D˞8�!��I&0� ���혷(1���H�4�!�d�(,�L� ��+L��w
ӥl�!�$N(5�Lt+�!3�������!�D�t5J��pN2��B��k�!��F�틆��:X>J���*2n�!򄞘-�5�EF�L�l�A�Ɍ	q��{"��U�Ȑ �9OB���� (��j��َ~�`<b!"O=H�e_cmȤc��X�>� �����:�������h�����/&E2`r�ɉQ��8�"O�&��8fƝ;�Ww4�1�Ɋ bU��3&�yy��g����*K����B�
@�pU�Q(ȸ p����P�0�)��0�.V�P��W�	C��C G��,*�Q�M�r����� ʽ	���7s�� @@�X�0�.�)��<��ة2�$�	��~R�`��Ui
y���6@�p���L�����?c�\E�vm0�Oy3��0k���I�E--F��V@�WN���o��~"�L67��
�Y�xT�4�2�O���ϵ~p��0���a���~�ּ@�z�'�ʼ"��2����.����Mӽj�P��wa��;�v��w�FF�(�æ�T�z�јs�O�$"�u�gy��J�Iн�S&��CI��!C\��[�A�gH�?��Ɠw�ꌡ�0�9<B,�{��2��[2���h�*��c��"qX8@��P;&����dش�R\h�[
"�Th��LW95��E�I�D���p�Ķ}�j���~Ba�Q
m���*��P2jX1���S .��$���'M�tA�b(�O�$�,�/rr������&2�"-�1�*t��B�����?1��R0r�R�.rt����ɿ>��ԻB�I�!�v�N��E�&�2��q�џh�!��:4�5���'z�IB�(��n$�G̒����$�rPzT'F3��9�)�:��	��d,���-�d�nP��l��1�4TGN��'�<�AN��K�O�ݺ��ݣ|����������3�Ƣw����E�~r��"2��4]x��|`��]�P�JQ۷�!/Lv��e��<�j�xq�9���#X�b>⒄�	!]�lp��]�sKP�qC@��H1[P��1q��Bቹ$�H�Xb������g�xh
g�D�$��$�<��ܫ ��8�*�j+���|�����.�
y���Zjk��6�Hi؟9��e�8��@���?|v�����zY��cT��{(<�t�tC�*X6Kq�^R�'!�5�LU�'b���QP!d��+¡|��ʠ�B�	,b��a�ՎQ$����LW <B�	"7��[�+�=rN�B�(���C�ID؍�Ħ�#�(��`�+u�\C�	�#1V��c�r\zp �M'K�C�	f�P�P��?�T�3ץ�-s�C䉜'R¨[�J�<@Y�Ujv��B�I2TBhh*Ѝ�f�Up�cª^��B��!o�:mS'��zP�@�ku"O��$�K�>�>����Ӵ?�����"O���ի�G^�Ǘ�x�Z�a�"OVy	��k>�,����,;,89��'����M�|�ɧ����M7*��H�c`��~3�M?D�\ALմS٬H񧡔N�j��ñ>�F�ʾ��d�t <OJic�"9$�ད5��|;`�q��'G���U&M&Qݔ�X��_�T�� YK�-�̋fA�T��=YEO(�OQ�k�	!��}CR��-<భS��I:W]y�+B%��mk!�,=��Su]R}pW�U�a	<@e���ir��Uv7X��{��)��^Ut�b
� N7��H��4N�>���G/p�X8��C��G��\�4��n��?�Ҽ~�Ҩ�#�H'����4	c}��@�(�D�'��$�bGծKu	E)�Q숣�	̃,tP������V��)�p�:���O�!�%ϻ<��,ࢄ�1 D�a��>S�(��C"Q8�p>�����B��� )�ԥs�F���x���/1�@����\9"o.I�'`��Z#��vB�T�O�������^�� #0Tt�2�<Q����@hF�[��0s@��W��lѫ6�U���4=c�\:5ڮ��R��_6,��U�K�"~�I3&Z�Q����Ш�S�F� �P4k�嘤jVP|��M�8�vX���s��?�t T
��(yP���FQV�P �CB?�5�I�D����*%LOV��m&�Q��Ğ2��I�^��N��F�^�hI�]cj���m{���$�yGT��wm@(Th���憜'�#�9o��ū�8�O�ͻ$��1nmj��Q�D�T���H-#�U��#B�{!LQ?I�/
��@�@��^�
c�#+ʡ�!"��"Ƃ�y����*%F��p������( L��P���!F�,[� ��TN��Xh��\�D�<К��O���Q�>�+��=���>�$A%hX{G� 5uy�QرD۷3�1O�Yȑ[7����:����O���V���0� �A��V��C�4��0h h��DN��t�"C�6��e�̕$>��heA0}��Y*Lp,��j`�''7^Q ��k�B4�w��0/�
Q'n�jݠ�c�"O��CIA�qo��@�n�I�`���� �9��&�b隥�0�3�dɽi$��P��%yx)�$�8(A�𤞵b��������I#�2$YJ����"M�t		�EC��(�D�!2Bv��c����x�'ă%8V$ё�M~R�]�5���a� 46y�Q�e�yRۨ�s����J�#	���	+u,^%�{�R*�5yLZ��~BpM��G�T�˃��9�ԋ���n�<��
�N���Bᎂ���K�)8�B���,�<x�H�f����~
J�� �)aƝ��l0��;�H�1O�42���n��q�i�+Q�&�ab��#B�
E��!�l�*��$t���D@�l�Б�1 �L`M:�hF�[8�~2d����3�m�y�5h2'$?�e���G�~���'ڃ'q�I���'�� �2@GLM��V�ً�K,	l�p`N�������?��$��KHI�(h�  �x�Х�-�yb/�5Kaj�FY�2 y�P ��~r�O�5���q	��|,p��-Z�3��\E�$��H4�BAD�D�9�@ʜ�y�C��L��ە��8��I��BQ16;X��do��X���c���	$ 5SK?91r�V�K����N�a�,�	Q�1BA�~b,��_}6y2�E�75���y$.]��$hC��EQ�d{�
�A���
���B�����\�_,�!� �2#�D�o!ʓ��BܣY#���BU� �x�����}*������!\&��bCS�B]\�B�.#D����%��)�`���L�8q���0˺zZ�1�b��^�ք�G�,y���'� ,�b>睴n0͉p�R�lv��@3�1u��B�ɧcTZ�1�hj�+#�)q�|L:�)vrs��*-f�B��Ʀ�b�g#2��yҭ��S��Qŝ"qX�g�X��=�QGE�|<�Ua�ME Pݘ ꊉX׸ ���"whr�ѡQ����m˳-}v$zӓ\4T�gsS���-�0<[��?և��e�p�2V����X��CZ�c}��Y/���9Ѓ�pG̕���v����ы9D���aD]xX��#��-����T�L�y�w`ŋL3�a�2̋)�LɲA݄��O����%A�
i�TOz���1�!�D�>y�(�����^*F�r�N��
�b)�<��(���o؞�r��R/<,L-�%� &�Y��(|O~`�b�� ���bشWd��Q�[5A6�,����=ǀ%��
c��c%ƥ<
>]x�"��|�i�?��/�Nȴ�*ҧP �Cq/'\�
�\
e�%�ȓJ(t�$O�N�(ɔ�D?Nʄ����/I7�\I>E��'��i�AH,=x1Q�F!]�hM��'?���D��-�X�*Jix�8�'y�e9�(�R��`�ݱ?��P�urAT�;��:D�ث�	�#ႌ��Yv���B�8D�x�%.���V%�`��?T)cl4D�cKύ @���m�99�U��	)D��b�蚬ѪX� �E�ʙ��!'D�`i�k	 :~\)�7��;/&HA���&D��aਃ�5���)N���`��@(D�Գ�e�;Zn��ʂ�n`�v�)D� K�O�-XvTh�k��;L��3�%D�\��L�)*�Z�zU.�,k�VۗB6D���+��+"�q�
�f,>5��0D�P�Ä�0\x8ՀG\�k7}1��1D�`6dW����{���,��<�*D�����A�$�k�-��2�xIbc)D�4�w���14�K��V�=ӞĊ��8D�@�W�S`b��'d�נ䀤6D�Tr�ȃnp�cE�dШ<[6�5D�\�鑀Px�����T%"=�ܚf`0D������!$���3S�26f޸��-D�ȉ��AX)�m�0Nn��+D��$f��>�1t�ӐL�`5`��2D��e�����%C�Ռ}��W&/D��x�Y��Lju�Ъ?��pj9D�����T }��l@(Nh�Xq�H4D� ��C�S]��[���4��ؖo8�	�;���f�ف5-A%��<R��b����Ŋ�d~\�	�?������3D�dI4��&_| &� ~�d��R�6D��QBֆ8��6��4�6��6D��9�)�9;��y/D�e�hHS�g3D������z�Z)iP��� ?f��2D���a	7y��. �<[�B��?�!���<���s��|m��b0lݎo!�Ю"�t|�5�N�B���e
 �ON%Fx�nv�z��."��iRt��/�(��w��O��$!��??)��T�2�@�ARL?�� ��x�E�	K*��㨈[�ְ�w?O&�����	1����EH�<E�TGΛDg��x#���	�SJY(t�Ad��7��	Z����S(���sw��$,d;�C=7K<a��M�wZ�zo��g�T>-8�Lޱ`lX�Ʈ�(V�P���S��'�T���2�s��s�04���'JN���o�*a�(C "O��r#�-xit���ֿ%ͺ��"O���l��-{<h8��'\"80�p"O���0Y�S1� E�_ ��"O�a�V�2V�
I��MR�1Ʃ85"O�T�q�'�*GJ��%t� `�'ϦəC�0M��� xj���'E��s�*�|}>cĉB?~`����'b�q9ɛ��Tb��|��գ�'ð��A&�\������x��`{�'H8����b���T4_��|�
�'C�eX,�wK�H�DT�Q����
�'����'B"%�2|���W14�|�	�'�~���΅C7�i�R��%}��h	�'\���_�.�
�+��Y�]Z ��'�R�Ae��5d��tǀ�� ��U�'Qnت0
�S��Z�#�0|.H��'^�!����t(��*���y2⚯y���u���*�c���yB�ݙ[C4�!�A�+^6L�B�!�y�Nʧ@�*1����)�.	�s�ؚ�y�R�C
���,(�d9v`�y��,~h�#lZ�$\iUo�y ՐB���;/�
���t*P�y���uU%t/��Xf��wJ��y�D	,E}>��w��>��`D`Ӹ�yM�VO$es�4FZ^=1O��yNθWf�����'k�E����yBh�	&:1;`�S�"�1͘��y��-|L̈�QB-L�)9�͎��yrC�;: h!��u����'L@��y�`�b?�p�§#�Rб�Y��y��(.��[W��-_"h��gN��y�#��jte8g�*ܠ����yI�`�����J$V�(|w��yb��>���GC+J�Z�ef�x�<IuD�}o���B�!��9%�BE�<��GV,l�BU�1���ȡ�h�<�䥀R����r�ؒQ����P�Z�<1�����ȅS����"HM~�<q�ǋLȅ�gIT�(Ԡ8v��}�<�@�'������2� �GKA^�<9'�`)R]�DM
�Y���E�\�<�4��V[��r�eC8��D�W�<Y��p�!�m�lu�a�&�ES�<)u@[
�j$⵪ڽUD��0�H	D�<!bb�-Sp��PL:�@�&��T�<�1��,.�MhGd5m�0�3�T�<���,E'�X�A�0:���ٚz�<�!��9L�d�ROE�yz>���P�<��M�=1���S�
�5u�PU��M�<�gAʮ#t��J5�ʴy��M�%�MQ�<Q�B�A)�bѬN�k��X�<Y�G	�h����tH^&{a�آ"��x�<AD�]%W=VT��B��N�N�*e��v�<1c�6�� j����J�b�iE �s�<9U�7����n��_F-�3F�j�<AgG"_"�h ����t�i�<�nPrP���ÿ/��6(�l�<y���/����ed\�m,h�)���n�<� ��"GÓZ\b٨��E�	�d"Oj�"���|�h���{��%��"O��6�J�7^��C��(	t�˥"O��j���6aF�A��lY�+6D�"O��
gA��q��I�Q���4"O<��bA���t���V-6',���"O�y�`�@�����!ڴ��"OZ�	b	�_c@�5b�7f�̍��"OJIs� ���x)�/z�쩨'"O I��h�t؀� �H(�0f"O��r@��f)90���tX0�"Or��T��=!c6y��H�\�r"O�\2F��	UC��9ԃ��}����"O.��e]�9��-�$b��!��"O� 2 B�.�.��G��%u��R�"O|H#G�K�e&�Yv!�,o�aC"O�!wJB�R��J�E+n`���e"O^�B�(RK#�9 �{���"O�i���O�{"�"�[���(G"OaP�iS=`����R��qs~��c"O�#��S9D���i�D]�F^�]��"O��Qw�"wq�]��eC O^�`A"O*�����=T��p��/|5ʼ�"O��2���4nX>m��jW�.���"O�It$ڑ8��y�1��.�	"OT=0��F�'^��ko8]0	�"O��S�!zv���G�Lu"Ot`����OeZ���ʁ=�A�&"O���愘/�. ��^��(��"O� �'�k%��� �' ��8"O �����w��\Su&�+iA\�"O��h��:?p � �c�F��#"O�yТS�B�pІ�J�Vv��"O�M(1&�(
G�aA�@��IB���"O����A�(=���P��1A.�dQs"O���ugSG<t�R	�%*δ(�"On�7I�B���7��?B�3"OV�J�l� ;�8���\�n��yR�Ւ&�4�)�����8�w+؁�yB�C�xy"��W�$73"�3�!8�yc��*WeAccH�ѕ#E��yR��5f5dc�I�Y8VQ��K�y�G��0a�ir����` $1C���y&] �|XP�_4/����Hſ�yR�Ơ7��=����>Y��'��/�yR�4	�e�����9t����@ݒ�yO]�5�̅1�*H�Y��}�1���yb�
�sA(5I�OɩZ�Ua�͢�yb��1Vh�p��R�V�����l3�yҢ�U�B��,�,MN �MF�y�O[1m��yw@�q���N��yr���n)IB��e���+F#N��y���8)���+�W<\L+�@��y��(n4p�	دQ�0�dÂ��y���j^&yG�ԚCg@��f��y�'P QB�҆D�g��@3�M/�y"��nJ�A����+U%���҉�y�	8tAVёw�$S�"8��IV��yҊ�9�V��ȃ:HC�u� M#�y��T��`�D'�;|"�j I��y��I9�@����>[�9z��y���2!
�k2㝌Si�@0�yR�^sZ���蓱�\$�d��*�yb�S�k�����N��2���H���y
� zd4)Η&�x��u��p�LH�"OJK���/;Dz��Dδ4w(\�"O�u� 
#sq@<�`�~��Ⱥu"O�c���*AŸ$�#�7Q���&"O0x��I�+n��ta���{K(�%"Ox(�dX�d�KMW�81��Q"O�İ��Fy�mBFF�='t���Q"O�A�s�%\�RJ僪N��0"OD(�@���N���d���a��"Ol 3B��72�f�AqE�1"p0ц"O�h��Ʌf�|;a�� &�q��"OV;��;���1/��h�T���"O��d�I�s|H$� ��5@d,�v"O��ҦϜtD�p��L�N�T�C"Ob )�̈́;C$x��� Շ1�\X1"O8�y�i+v�1���V�x�"O8qRuo�A���׳,r�(t"OH�*��E6JOv|I��I��ܸ�"OF�P1���SvXp�JQX�Q"O<� ��G�'�4-���F��"O�Y!6/��i��q'�ږ;ԒȈ"Or�iP'�6Grt]J�j��;^;�"O"!�Cj�%�V���׋G�i�"O��"�ݜ6��1��A�J2-q"Oh83�W�X�h{q�̝!:��"O�s��CH�c�'�O���"O�X"��J���Aas�T�"�̍Y$"O
�w��;7��$:B쏄�N��"Op%�Ĺ0 �g�^���C���!��NQc<���rDp���>U�!���>�����V.x���G|�!��A��Z=�T�_A�:�m�3�!�䋌a��[�O
�!3X����R� !�dܧw�L�9�m��$ụ�C#�!�$VR����%��L���Dn@!�dN8I� l��ı�|5���)!��3yr�qd&:�La�&�7!�䏋n�����T=r�,�3��T!�C��ܱ�)Ͻ_Ȓ�0�d�!0�!��
M�0��h�	L�1U�V�{�!�D�s=X�"�䛡��{c@\�b�!�΀8h���]$
��Q�`�!�dA>���4��-稠C�aJ��!��q\����J�Z��W	S�!���\�pEÿL��\�1���!�d��Q=؈�tΛ<
�R���iU7Y�!�d_�\�^�S�� 
mܖ8Yv��!�!��@��y��Q�E�BP �܅!�$O<��Y{7g���������!���qh���h� +�T�1���F�!��L�<�(XI5ƚdx��2�!��fQn��׀��))%/̺fn!�M �`PK�J�/�Hy�cN�e<!���?,��*掤6�]�%��B�!�d�1<�2L�6�(�j�AԟI�!�D[�*�\[�	����U6)�!��L
\�t���0_K�E�����!�U�����v�#9�-� +�k�!��F�>�L�`o�,J�X����V�!��@�����3v���cƐd!��٤(�F���Yz�ݓ��Պ�ȓ*~�IK�enm�U�ÕD`(��ʓ^������)bj�D�l3{�^B䉶.�D1�7��+y�^��P��S B�)� Ph��m5QF�L��Ø�AbQC "O
�H"���I�P;���$0r���"O�Ph� A�uԸ:T��+,��E"Ob�Dl�-���Q1�G3:T�+1"O�(K	�UȐ���M��cWy�<!D��~�B��Æ�� �BP����t�<��DQ�@,�F	͠����AW�<9���y��5��2m���`�S�<	���b�`�0��P��B�%HC���ȓ!G4�ʀgF{�v��ůKn[�Ą�hUhpI�H��"����� e�Q�ȓ5~���� (,� ���Ȝn��L��V���+SF٣Q�@���y��U�ȓXZ���C��Trp�,׾d�ЇȓHH&)Re*�=|�BAP��>S����QI��S��Sid��Z��'��݆ȓN!�9"�(?j�LŀW�J-ly�Y�ȓ/ي��a��oQ�h�wo)L�T��q-P��&CM2�*y�bEO#\,��ȓp��x[���		���r�&�ƹ�ȓ.��  @�?�   �  �  ,  �  *+  �6  �B  �M  �Y  �d  �n  5v  ��  /�  q�  Ϙ  5�  y�  ��  �  ��  �  :�  ��  ��  %�  }�  ��  �  L�  �  ��  2 W � � �" �* �1 9 `? �E �G  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<���C����P��1�ޜ�F�Ai�K���3bH-D�x��U�Y@�L �2�3��??�
�"�^��"D�*N��UOB?U�E�ȓ0�v���,[�� ��T�Y����ȓp�s�MӶs��yU��9�z`�ȓaZ`�;׎R<g�����;UU
)��X��qaE��?F�d�$��]�ц�rBj���H?�dg�A�5潆�%�:��(�j�  ��I��ȓs��Iȟ&�������~_����@J�<�%��"@+'I�WưH#�'�����˗0oءh�hY-O�xm�
�'�x bi~����N	�/>��	��� �5	1�#!�����:(D�D"O��B� 0X����IR+9^���"Ol����yӂ(��'<x	Z����	�j��[�M�e5根b��O<C��K�����'�a��`���(
C�	Jmry;�	('�u�!�B��B�IR�����a� J݂ �F����B�"'ޖ�V��
yH�q'$ʷC����hO�>�R��L�%����)��x%��Z�a=D� j��K\L�B"�35T��:D��qc�gN�x�&+
�E�U"��6D�ػQE�2��B
-m���颭'D���c�57.E��\�Ĳ����'D�����G�:��#%�$rR��V,%D�0%!X�Zք�EL�~4J,�@�.���<q�.uR������0G�y���X�<�bJ�?c'hA���	�$������]�<��2m�~i�FHͧ_�\Y���p(<A޴Pd��J��?�0�_^�y�ȓI�i+AI>0�L��'�ƛl�����6�X�9���&[^2��� -��T��~t&���\�(4��C��?�N5��Sj�pZ���k����FG�\��@�ȓ{��؂4�J-$,فW"L���ȓl�8E��3zAA���2h�م��zy���w�r�.������R����y�b����9���p:)��%���O��G�4�03Nx�A2f� ��xPŎ��ybJA|��|3���p�ˣ����4�S�OVxDG^R�H���ʨ$R��	�'B�T���X�T4�qk�W��
�'a,Ƃ��j�	��C	���yR��G�4�8��
R�Ip��8�y��sV*�򢫜��*����!�yAW)W�pl�4�y@��(l����	�'8�MI�,�1�6)��l��X��'^��N]b}j�����/����'a��Z��°O��Y�F��`�N�І���2����g�%;Z̀!$C�h�b��F{"�'���%ph�bE��6'�:�ˆ�	�U�ȓ!JA����T�ai�7L<��>��'Uў�M`�jC�Ԏ\%���AÈL��C��:!��M���C
b���ۥ���(:vC䉸 �Xe)�ꔹov����^;wF#?Q��iD4n��|�&�·��S�Nե4�!�.$� �.`�
ik.�:���M��H�P�!eh��`X�sdiфq��[7"OƜمg>�d�(A5&Y�7"O�1��ǜ31�U!��TF�DX�"O:u�.��LP�q���>\`$�s"O�IZ�@ͧ9Y"ݣ1&��wO�B�"O��!b9L��T�d�N�����"O�c��/Z������&��|Z�"O���ר��6�ї����m) "O�m��I HK�H�#�ߴ?���C0�O�ʓ�hO�O$���6n��+��%i�*�X���N>Y���	?�"|�`�
@�����@)j�����	��!�Á+Vl�fm��%~���I�&���j���!fQ�V
�X0@C�*���Wm�=����'�HF*���ɐϘ'�>�sqa�D�҄i�'�K�ϓ��O����
Dq˺��3�^HԼJ�"O]Sף�J` �S���!���"O(��%��Q���k�6P��E"O� � Y���;+�t���\q����$�O�YEz�O`F��	PF�=����%Ĥ�'�)�ǣR��ؘz3��"!XҝJ�'�ў�}r��>	�ē�jzr��pGWj���>	�� 1�T%�BS�k��Q�"/�\�[&�=�O�|�Ê&W�~�۴�� �Y�y��)�Ӱt!aV��W�T酢]*H�d�$��(O?��H��D�����O3H�&L��m�i�'�y"�܀Q�Α���s�n��E]6�y��^^��PrA�=;�̐��ے�y��H�H�����U9AHQ� ���y��A\5�H)�ヅ,�:(���M�yb�?>�Tm`�n�QG,䘰��/�yrEʖy�h����!I��g�@��yr��PEv(ʵ�ڞ�vaC' ��(O,��D��4�&�sOc�d�F��!-��>)J�"��D�O=���ЌK8y<P����Dt��q��D��'|��@E?.2��
��!���	�E�➨x�o��HUJ!D��B٢t��
��P�}y2��ܦ�E~b��0b����6�L9�����֜�0>��xB�H&�* �$3�6�y�Md�!�wXpp+4��6@y�P揇����u��}BشC�4-CM�$Mt���o4L���=Ն�����D�� _�ST(��w1B��qh�p]��I%��"H��U<�m:�a�%��!`��
ک%����ɷ[���B�G�dP,3��;G��B�I6� F��
 ��'�5'�B�	";�z�r@�r��Q�fl�11��'!�"=��7��g���:u��2:�hYXC�\�<���GH��,G.r��<�BX�<��N �J��i�*xטx�`k�V�<�%��Fv(��ϱp�*vŒ&"O^D@�ȱ5$q	�K�"��2"O|�k�aɟ ������}%ք�q"O`4ZI�(��T���
�EY�"O���D��՚3�$(Rތ�e"O�<ӵ����
`��dA� TR!�7"O ��U��T�V4�E��pB\0�"O衺�I��h������=,�p��"O�W�5�q�����@|�a�ŨBZ�<�uaO�o�����'ؾ�F�S�<IA@%:$��p*�
dp>����Z�<����x�:q�G��e��0c+MU�<A3�jdK�	[�r�L����O�<dG��>��M��d��I�NHH�d
p�<��	no�tЁY�X��s��'T��Y������pé����	�#D���Ƅ"q<���M�:4-����!D����a�O�:�J��@��͓h!D�h���^+슐1�l��f�	l D���С��Lv4{T�]��y��N D��K���"�!rAͬ@��ua�c<D��*q ��j�̽cP�~_�(���8T�x	"FX/ZV���ݣg�R�"OйR6� jx��P
ԨH�~$��"O���!��=.&�"#J.q����%"ON�3@Ӹ!%|��P��,y���	"O���Bƛ.~��͠4N��"��R"OԽ�#O�x|)��1�ޙC`"O�MbJ�F�r�R�oƟl��a"O�t9A�
��	��d99��e"O0̓$���n�|������K�F�RQ"O<��"��c�D��"[W��!SG"O� p���	K�׼�6K�&?��%Q"O�����N�&`ڶO՚x�j��q"O�Y�tk������N��t�.���"O� ���p�x���˟ؖ���"O.���	�2<N�D�Z/2�6Y���'�2�'���'���'r�'�b�'�<��B�x �9�bG�#*Fy���'0��'\��'�R�'B�'��'>1�gd_�a椠���	^���1��'�B�'R��'fB�'7"�'���'�B!��!_�A���@��-̆}�Q�' b�'���'�R�'���'ub�'� ����K$L��ǜ5t�y��'Q"�'T��'���'�2�'2�'6����Ёp�i!��F�t���&�'4b�'N"�'���'�'V��'6i�qȈNCR������4E=���'���'6��';��'N�'pR�'�lش���A�H%&���hSJC��?����?9���?a�Ӛlן��ٟX��]$N0&l��F�Zt�"@N$���۟,�	���Iן��	��<�	۟��	���M̎*>Y��ʞ@F���Iܟ��Iӟ��	ڟ��I˟ �Iܟ��ɟa��a���ɁG�x�#�
�A�ʤ������Iٟ������I̟���ӟ��I�X0V�����R=����t�20�I���	�H������ޟd�Iǟ��/m`\S�꜑݂}�!<�N-�	���	�4�	��	���	�4�?Q�5S��[�-�&w��(3�CG�>��9['U�$�	Oy���O*�mZ�pU�h@l
)��!t�g�%A8?A3�i�O�9O���P�&ᰰ�ށ@:�pc�X������O���6�y�����D ���OLf��U�|1��+V�>�h��y��'��	�O[^PQUo��0
 �nG��p��abӚ���D+� �Mϻh��H��D�+����0�^?VX	���?�'��)��9
`�oZ�<уO�&t&ri*r��("��<!�'���dX�hO�i�O
�hҧ��F����R?v�(]0W7O����4����ǘ')x�Q"��	iN
�XD��mg\�у�IB}"�'?O�|�~���FRf�YR��?����'0�摕>TyK�����՟|K��'��0�fdG	�>�Kc��
���a%X�h�'���9Ot�1AƷpǆ����9���49O�o���
W�F�4����s�>D��ZA@7_�.\;�8ON���ON�d֫"�>7�5?Y�O��	�)C��i�5�p�Z�{�H�yp:L>Y*O�)�OF�D�Ob���Op��k�"Wl������lp ���<)B�i�A���'M��'�OL�`��~Mȹz�aZ�k9F�X��"x�\Û�i&�)�Q�XͲPg�HJ��E��:+��!e=p�T���_툽�HۊZ���;<�'�^�
����AU$UM�X�?C�L#���?����?!��|�,Oj�n<_2�A�I�3&h�&��Mz���1*�)&I����/�M{�i�>�F�i�6٦e�S���`��eW�I�r	9AL,_��o��<�!�S.#'Pɘ�'�3T0�xN?1���w����/S>m�p���'P��@�'���'���'���'���;F�T�hp<h9��6F����OB���O Ym�]��-�'1�6-3��Ō57��b�`	=k�.\�R��X�$�\��4JF��O�6�b�i��ɋ]n�Z��U�*"l Q�֐o�X�� ��T��"�Ty��b�h˓�?a���?�����k��:�e�o�pqI���?I.O0�oZ.r����	��Iv����HX�x��,Ȋ7�
c����d�Yy��'�e)�T>���A����E	�	�8���tJ�*M*T��+Ѕp5�P�'�6�]�N��Hwy�wt�:�iC�k�<�n�a5x�J��'�R�'���O���M�DmX�d��-x�M�V�U���{)�k��?��ia�O(X�'�P6�ų]�i`���@��03�M�M��8o���M������M��O�e������M�<��\�j�"�z ���J��y��އ<n�]�P�	̟��	��H�I� �O�\,�S�J%f8d����<R�p�0pLb�b��B�OT��O��V���Ǧ��-�zp�r✋�~Iг�%F�<��4NP���!��Ԃ(��7�m�`�C,Y�&3vQ�T�w� 0n�!eH�$��4A�� ��nM��Y�,��͟�@���)y�8�C�J9|~�!�@Ο$�I�(�	Dy��aӢjg��O&�d�OP�(DA�t�1�2��i� M��!5��/��D�֦9h�4_�'�]��N9MȪx3��N�[�&���O�UAg`D�~ӠM
Ca�<iF��Z���2����;첝��E�&c�l�S��`����O�D�OB�$(ڧ�?�r�z �ࡣ���¥r`�ӕ�?���iČ����'�`�f��]p�*���"@]�H�-Vc�扡�MS�i�z7l�6�#?���\�?��	Y�N��*l�mI����@(/b�%�.O�!m�LyR�'K"�'2�'�bLݟ;�4%�c��L��E�#��	��M��IC�����O��?�h �
��� �W�#L�a&����I��0ڴ>ω��O����0��2����~|:�`�^8
���`�W����
{���Lyҧs�X��8� ��p��YjU��O`�,����?���?��|�*O��l��N%��I�VG�!���G2z'�`r!Ȁ�r�
�	�M�2d�>���i^�7m���h�"��3�,y��RK�	�sa� bwĹnA~2(O�Q7^��S���!�u���� =kҠ��v���Yↇ�t��8O8���O0�D�OX���O��?m8��K�9���dKW�8�(�)a��ǟ���ϟ�kڴ*Q���O~7�>��$�ƌyeօ���[����PL&�d�	�<��s���oc~�B��h�sd�݆r�|��&�P�gL��Q�����D(Ǟ|�P����\�	şd�AO�{ ~�£��M�l�$D�����	jy��w�,%뵅�O\�d�O��'})(� !G�H˥F]�=Tm�'����?шʟ$ �S�YSHx;D�H�'�@m�k�&���G�7A���|�'�O�:J>�7�C h��P@F��P`j𢐵�?����?i��?�'`���N���D����k�V%�Y! �Z��2���a>����Пx��4���|�Q� o 5N�<�"ڮ%��I���|s^]K�4A9�V�ӓr�6<O �DXJ�D=���.��iوn��_b�5��m�)L�̀I:O���?����?9��?�����	^#���[rdK*h.T���5A�l�n�EɌ̲�"˟���?��쟜�I��M�;����BhK�h�ڔl̥`�f���'����=��O
�T�Oo�xu�ie���{��e�R���My��:1���! &%��]���O��|��4�t���i�}����c�)J��?����?�+OĔn�gT���ܟ�	�l��,���_���$';����?�P������x&�l〣T�P����� {�P�"� ?9r�ƇS%��Gh���T&��$�?�CY�O���
%/؆��T���?I���?����?y����O�0��ҟ; 9yf�,|�Xxyc)�O�m�Y�����˟�Yݴ���y�!�L&�(����J��В�yb�'��I!<�1m�d~��_�d�9��L�\�y�fŲ lؔ��cZ���|�W����ߟ��	ڟ��I����ҍ�0e�����$8P �HyRkxӴ����OB���O蓟D��ԿA&h���m8Yf�-�a�'�7OjO1��
���.`��Hs�(a�5JӡԄY���RF-�<y�hJ�Vr�5����䃇W؄	R�]�;�(�A�ݷ����O����O��4���eě��Nb.�;
�`�)�M.R�;b/L,6���rӸ�T��O��o�5�Mc��i'xĉg�7$ �d�ݗ�th�#Î+J��f������v�������TZ� ��ň��q�4a69ON�d�O����O����OD�?�`dK9NO���S�Ҕv�H `�����Iݟt���:��S��D�ڴ��j��qD+C�j�L*��I-l<�v�|��'m��"�<x �4��䚥lD��Ѭ� ��:h�Y[��gY��?Y�O9�D�<Y���?A��?qFo�!�Q����tʥ��Y��?����ć��
�ΐ͟���ʟ��OF~��pC
 ���`��T�D�8P��O�y�'-b:OFO���Y�b}����
�����.N"
�Np��,BQ�� ��Oy�Om���#v�'[�M�Q��Z��B
P5o�Z�'��'����O��I�MC2����q�!7iR��
>��� (O�@lZR��$7�	��M���4v�i"c��c�l�Pv���\�r�i#�$H�i=���;�4�)��O�l�'���+5����I9���wX��'P�	ԟ�����Iџ��H��ER0k̬CC�W=h��cP��*/\7m�wil�D�Or��+�i�O4�mz�!
�-: ����
+kTX���
�M�P�i�bO1��]['�n�(�*4����5@�ڄX�bD�&�*�ɻQ�*!��'8F�%�(���d�'���u�="T^ԁ�bˌ(l :��'�'7�S�t�ܴ4n�D����?����ݠ ��d#ԁ� e��2�r���>�1�i�D6M�T�	%e����j+2U[�H��5D:�W0�
�R�k�X�|����O�X��H���¡�y�����C:M�ti����?���?����h�"�D�x�V�rG�e��B�M�7m����������y�my���杁DGB	"q�T`��iQnK0 	�ȟ��'��ԁ��i��I�Ӷ,��OBBA	�C�h9��+�+���BǩIF�Iky��'�r�'���'���*p����d�n���c��4��	��?��Ο��I�T$?��ɐg�l����#mz�i��AT�f찰A�O�mo���?aN<�|*&B�=y{��$�b��R�gG�   4I�g���� �P�� JOʓ�4�0���8�j��Dc�S\�H���?1���?���|"(O�!l�A���ɶ1ۈ���;m��@G��"f��M��c�>A��i��Dl��;��g`K���(Ae�b*���e���%ڀ� T���J~Z����k I)X&��I�kr1��e�0������I�����֟�'?�[�
�-�|���ΨN�� �3`�  @ � �쟼�I#�M��GԀ�?���4��f�|�d 2��Z��"%Y l�E��b��x�M`ӂ�m��?u	A�Ц��?i���%�:)�U,��d�.�hg�C*P�q�B��Oz9@N>�*O�I�Oz���O�lXsQ�IxQ�s��,-�65W��O^�Ĵ<��i�����'�2�'�哊c�q9vg�^�>���Ȗj��.�����(�	��S����g(�K����82e��e��qp�+H���<b�O����?�b>���q�v�h��	#�S%�
�:���$�O����O���<��inh�ÊRv�� ��%�t�dH<9���'5~7�%�����VЦIR`Ӡ"��T/C4>�lJ6���?!ڴ%�Z�ڴ��$y�h���f��S�? �q�L^T��ƀP�F��Di�<O�˓�?���?����?)���ɍ#>rï�A��(�-�:xMP�mږ='���'��D�'6�7=�`i��G*�(nLwv�� F�O��b>�;�Nڦ��"[���A�
~���&��Oyp�ϓlvB�@�O��N>i)O���O��ـ'�wR��d�J]s��O*���OD��<�ƺiv��rB�'�"�'�V�zdn����Rg�3z�� ��|r�'��3����i��%�Xy3G$@���P���nj�U��$z��I�N(;�-\�
^����6 �O�h���E~0w��
\��EXT�M�pW�Q��?Y��?�����?���?)"f�6x��_)J}:���NZ�v��$�I,�M����?9��S`�f�|��yW��MJ
�!�F�p����U�ۈ�y��pӾ�lڡ�M�p�4�M��'r�[,����M`�4@p-Õ Vm���O�M���%�d���$�'��'�R�'���hT��.����"�Ҫ3�@���_����4i�L�)��?I���'�?���W�z�2m�Ь�6��pi��������Mc��iE�O1���K��Ǥ'.�d��)�6;;�P0s$Nm�@MR�����ș-��DQ�IYyb�À�Z,N�6<;��ηT'Hi���?��?���|*-Ot�lZ73�6�ɠ<�ꅂ���% �8!ˁm��pl@扠�M���
�>A��?Y��iΊ](�M
��и14�I�I3� a�Y'%I����������c���i��2�q�W5%��Uí_�&�]	V1Or���O���OD���O��?�U��	x���1��K�F������Q�4FX��!.O�qlY��h<�rA�"�pc"�_�Ɔ��I<��iz6=��p�"lqӆ�q3���(�:T4V�a�\�pA�C�<�6��W�����4�����O����PF*�� 4�x�z5��|,n�$�O$�y�v-�#�R�'0"[>5٣/Rl�����'�>�i4)"?	 _� �I㟄�N<�OB�A�p�ɚS���ɔJ^k�V�q��Զ�Y�@���4��e���0�P�O��Ȇ�Õ���f�(%��J�b�O�D�O��d�O1���B��D�+\邠!˛0 !�엂=ܾձr�'B�eӔ��X�O���2�Z����F�<����6nhʓJ�P!ش���cIx�a��:��ʓe��F#W�K5�8+bӨ��(����O���O���O8�D�|
�*Ʈ%�:��� �?���'�Q�s��6M��5=��'�"����'ފ7=�( �뚡69�%Z�d�j2�3��N��:���Ş�>!��4�y����tԸ���,�p����A_
�yb��~���	|P�'��Iԟ0���u�,@l8�ir�*d�nu��ǟL���x�'Y|6m�L��d�O"���=r�؁1N'bx
�:�C�W9d⟔��Oɦ��ܴF��'��  �A w2��`d,+ps��On8Y�h�Oʰ5H��)��?�l�O���P��=G����U0>�=9s��OR���O���Ọ}2��9wd]��
�o���a�l�����.��f�Q�;.��'\�6m+�i�]P4䏾M:�C��-�.d�Q���d��ʦ�:ٴ�d��4����	!��h��+@k%�U�"ڊI���~�}0DϘ�����4����O����O�G켠aQ�E���eAV �e��狍�2�'R����'���Ƨ^$�!�]�q���c���<���M;��|J~�E/W=I���ӨT1a76����H��T!�q�c�O�)�K>�+O�u�G�XS��_ k����O����O��d�O��<	շi��RP�'�\�	fᅰx�����4����'56�#�����$ͦ�Iڴ@��ƣ�j7�\y���`2(�X��:$h�봵i��Ib\���`�OCq�r�NYGq�(0�K>�<I�á_�U���O��$�O����O���-�	7������_�$��@%'�؜�	؟��Ɂ�M�E�@")O�dn@�I��f!1$���P-`��ȝ(_�ZI<���i��6=��5Zd�~��D) ��3I�����:��0C��ғ2�0��ܸ����4����OF����<�y�����@}h���T8
�d�O�˓D�V��pYR�'�2W>���H�6��Ф��O$�S�%?!4S����ƦbK>�Oi��Ri��#-4�n���d9֦�!)����1D5��4�h=��`^��O�pI��+|^\(���"���b��O�D�O����O1��˓`��#H�(m�!�J�B����f�ٰN��ԃ��'���mӄ��J�O�mZ?wkv����	�45"�#ya�Q�M끵i��s��i��I,�X�ؐ�O*�B�(rB(�!w�r����ܬj�B!Γ���O ���O���O���|*&,F�8�||`�N�Bƨ*��C�A��DYB�'�B�I�צ��y���	CK�/��Ix��]%�����?�J>%?M�wGަ�ϓs�H��)�1��8r&�]#I�r ϓN��B�O�5�N>I+O��$�O�	z�	ݔx#��H �Ԧkv�Qz�+�O\�D�O����<A��i���s�'���'�eS�n�13fU�®��w�U���}��'��$���C�p`$�ڃ P@$�t��B}�	�;�*$��7��<'?12��'�����B]:�1�ǁvK ���H���M��ʟX��͟���T�'x�6�0��-�ʘ@3o�	�H�N$ٜI��ϛ�ϝ*��'�Z7��O���?�;�����j]D�\	8Aaʺr�V5�K������Xl�'8ioZ�<A�έ�'/����� Di�tm��r���L�R �h2g4�ĭ<�'�?���?����?i��6"�Lz$K�Q��  ���?��$����!�����ӟ$&?���9^�昲䞧fb*��t���%۬O���&�)��LA��2�����Ӣ�
���g�j�'q`��Ä�ޟ,�ѐ|�T�����L�I�� T�j��H�$����X�I���Iܟ��Ly(}Ӳx�g��O��E�q����雇hd-09OHmZX��u��ߟ��I��Md�0M�Nx���ʡH|m���ġ��sߴ����>>�,���'��O��ĕ�9���G��!J�$ �2��.�y��'��'�b�'���	�_�r�0�� u0X�f'͍j~����O�����u��o>����M�J>Y0)TY(���E�k
��������'7�7O�d�Z2sh����$���������YBl��%5�d��E��H_M�	^yB�'C��'a2�Ԙkc.�+v*��-=��bdK���'��	��M6�5�?)��?i*��H�,�=zD�􎃭.2�2��H��O�l��?	L<�Ooja�d���m@w�цQ�v��d˄fP�n��i>�r2�'o�y'�LrF��w_6U�#�,jb}Ӡ-����	�l�I�b>%�'��7��D����m���h�E��P��Q��O0��L��m�?Q�]�p�I5b�>pyf�D�b$ )bBKE7�6U�'�p��ߴ����3p&���X*:ʓ�$�2�bI!��	SY������O���O��D�OP�Ŀ|�PF�$�f�����@8�I$)Y��fU�^PR�'��O��0�O'b�{���1R挹�#=h��k�"0:^8��,�i>��	ߟD� ��ݦU͓xgx$�waVI��Ó��:�v�ϓ}
��D��O��I>�,Ox�d�O�܂��(+��9u���6lX`q��O���O~��<��i��3��'8R�'�����@�:㌩	�NF7,Q��#��ďW}��'�O���C@�mF�dB��Ƿ_HL�HA����gY�u�|���IO��t���	ݟ�0'J��b_����W|�D��E�ǟD�Iџ����XD���'0,49����zx��sP=}��$���'�v6�y�d�$�O>�lf�Ӽ�G`ϥ�LPQ��$���ӑ���<yU�i� 6����+".�Φq�'
�!�G�?����Vj�1v�k.v�:g뛛K�'+�i>=�	�8�I�l�I�}æA�P�кhf���-�^Ԙ�'��7-�/R��Y1��O8�d���3a��O���R�had�� ��SA�Ԁ���	����'r�i/�O��Oa��������@�Ɲ07����ʳ[�.TpD _%��$�=��M���@*�O��)����D����D܏M��4���?����?Y��|b.O��mڄQs��	�%��T.�1� �o�p�
d�'�7� �	=��$P�����4J�c�6�JqC''��dJv�\"?+j0ɢ�ie�	�r������OIq�j��U�`��u�┿;�����3+O�D�O��$�O����O~��>�ӻP�J|�gc6���+�#'M<����`��<�M�q���|���=K�f�|2ဃ,S��˚�!� � �EM
�O�m�󩚧jhv6)?�p@Ws��$�O +���ϫ-s �W��O��J>�/O���O���OBi�u�سL�0���,L�i3�O����<iV�i�4ٲ]����`��+�)�&�	U�}R�u���,��D�qy�'țM2�T>���O�G�D!��!��][a��	<��-�0�^� ���|ⲁ�O�Q)L>�3�\ t�N�a��*O���
��0�?���?9��?�|�-Oh<nڿE<0��8nJ��� �"R쮝���������M�B&�<��4�9@��;�<���"�
^V�a`�ij7�D�9�7-$?P���4�,��:����{65���,Nؐ�
�e���yrP�d�	ş �	ҟ`���`�O�z�1����1��� ��L(,�O �� ��L���'��ݟ��I���9VʈHs#�&Blx
Q�4#�Ν���?)�Oj�������H�Qch���If�p0�jðs�L<�B<g�p扳1�6(#��'�.�&�$�'���'���*�!:"0�pR �V"�u� �'NB�Ԙz�"W� ��4zX0-���?q���8�d
�_u�Iӄժ���bI>a��$��	=�M�v�ih�Oh�P�`ʖ)'���j��3(ļ�!8O:�$� �F���d؋��I�?�P��'=���M�$��fDU:�*�!�T�$��ȟH��۟���W�O�*���^��e�&>�Z�9�M7,��mbӼh�ԇ�<	d�i��O��<-]j�Q)�ki&�jA� &��Or�I�@��˦Y�'�
@��?A�.� ���C�2Pv�30�N�a�ԫ�n��@��E:	O��lC�0�>p ��F&Ts��K�u�n4k�&Cq�0y�(B)tXB�����D񔈝�K��$#Ĥ��tmp�	b
U��m;�l
9Tg>m�ģ>��='�T�br�S)c1��M�98GF�R��.A1rG$f�L�#3��7� JB=KL��gO�7$6�WAƈ�)b�d�oiL�qͦGi�\i��90#^�Q�gã��<��G˞ PxI�ra�{AN��Ȩ[Q��*�v5\|���B3J�@mkw���+߮Y��ʘ$P ���OH�D�<���?)�k�4���Ӛ��ac,�9e�*���i�b�'��+W�:����O���)���'[ܠX��KF�b�N��43)�Y9���?!/O����</On�cd�E���f(�*C�l�2*������R`*�b�"|���.@��[��[b��h�r��7v�4D��i8�'T��C�o��'��S����{����2�P$k�,[�\�0m@��H�Z�ΐ'>��	ǟT�ɂ�� �a����,m��25m�E٦B�i��&ЅY��	��	�OH�Oa��)�;+��5�G��g�=�è�Y}c#`����OR��O���<��7TF�Tr#�
W�Ip��ntST���'�2�|��'��/��|���!#'@�AEQ,3�Q���|�'���'c�	�U�Δ �O��RfB�e}6$E��m ����4���O�O��$�ON��%�����k��[��Mr�Ӊk��8�K�>���?�����S>n��t�O��kث̉�RH �Y��1 D4U�7��OL�O���O�4�t��Oz5yQU�4����0�௎<Z�H� ��w����O�˓*��ɱ\?��	�t�S<d��kRB"�p��ޛ��tM<���?�#��'^�)�WN�(���O\>|8d y���Z������M���?!���BgP���=���R�A�*��tA��ďxI7��O^�V�zt���}�S ݒ�PP@KM�
�XM�E,NӦAS�fܢ�M���?���BQ���'ٖ�q�O�0Ҽi���[�$[N�rwm|ӄh�t�:�����?A��w�t��5��-	ct隑+�n&�f�'�2�'�0��A��>�-Ot�䦟`�!2G�"�@��H�-�4C'�a�ޙ�����3�Ҏ�ħ�?���?��m�/1-�$i^��`��!�BA��icR��8]܊ꓦ��O��Ok�]�E�*�zQ��H&V�Y�
��f]��*N�rb���I�@��Jy2h?1�p��ƽ 2:D�����nՖ��c�>�)O��$#�D�O���&@��|[�r:h�I��^t���-�D�O����OJ�-/�|�F2�X8�H�|��Ъ��8٬�#İi�	͟�$���I͟t���Sa?qcoD�^�q��P3O�VX�"�i}��'�r�'P�I�^ݢ�q����DD�k���sP�P�)��h!�Ǳ��yn����&�p�����!���ޟ��>�E�".���i�<~��hx�,�����쟨�'!�L�~r���?I�'� ,ЧY�m���Q3����x��'�$�@�O����i�.�c#�.���n#$.v6M�<���V�'�2�'���o�>��R�Dyc�ߎ&�U*��J�1��l�����	kb�A�?Y����P����sU��$>�hE�� �M���[�.����'�'l�T�5�4�X\P0Έk���T"�L��k����	؟(�	B�i>��'�2e�)*���������Dɱd��7��O6�D�O�s�x�i>���P?���B�EY�����hvE�@˦���w�	���9O��$�Ob��B
n@�8���	`<HD��XdmZȟ�Ȕ6���|�����Ӻ;� ��@���(ʀZ�9��OJ�Iߟ�'���'c\�DBŹeǂ�)~.j�۷%Q�*�$٨t��v���H���byZw�NQ!sAQ5OR��CH��Lx�4�?�/Of���O��$�<I��]�},��19�@��1"�����@Q(�����	n�vy�O��$G�3a[��C�(��e��aD�uf�ꓝ?Y��?9+O�L���u�ӘA�ZyᰯV )��T��Î']����4�?L>1.O�i�Of�O�j�5
�~�D�I�Ōњ!�l����<9�����-�����O���Ʈuӳ��K�\Q�V^�@LsԔx��'��I!b#<�;Ys�J7�8\X���p�@h�'b
�/�B�'��'��dY���E�*5�a-��5��iJ��27��O��7���GxJ|Ԇ-E]X�sc�6_��9��O��1�e�O����O"����$�S�ԏ�g5�L:E�<���*c䀚7A��E�Gx������L��+2)ZU�� I	Md,�nܟ��I��hg��Eyʟ��'�`(��]�h����CE	h�th��>R��O���'����5~�^�A@]�˒�!k.6�7-�Ox���c�R�i>��	H�i�K�&O�+ŊĢ�,ȟ;���@f�-�$�O���?	��?�.O.�C�͂�F�Rt�s�>�"����	�0��&�@��ß�'�D��u��-'�~ɀ�eY�4Y2,��M�������O0�$�O0ʓŔ��U:�*yH�Q?Q}���j U6�P��^���IƟ��	lyr�'��矐zf�@�; �Òb�z`�1�����O~�D�OB�J��G�}�ӊ;����"��0���*]��Z �ߴ�?�K>	.O�	�OX�OŬ�ٖ��	���Z�.�3xj�4�?	����0fW6a'>��	�?�ؾ9����`�`�U��R�?��Ol˓t�&�����'��tCη[�nL&l� F�T]Y4���M�.O�x�*�E��� �D��,�'2J%��a�4j���Hȟ������4�?��p�>��"��S�����s�ܴ>�*���gR�#M�Y��yV�nZW��(�	����T��ryʟ(�qq��x٢�&E�Gh`����-Ȗ+�+	�>c�"|:�P h�SE�lpx��	�d�v5�i0��'����/Z ����O��I<j��m���*�0��%��;0�7��OR�N���S�t�'��'��]!�]� D����-�x��x"�|����\�TL��'��I�Ԕ'�ZcK�Œ�$U3����@E�/�ΰx�4'�fY!3���<���?A���?�����$��T�Y��0�Nѐ�.�Of�ȱA�X}�Z�H�Ipy��' 2�'CD����G83�L��b!N�������d�O0���O���<	w��?t��� ^�05��*1jH��!i��4�нi��I֟��'�2�'X2N�y�j"Q�ꠐ�>K^��#ŁUw���?	���?�+O @�w��v���'��4���J/=��; h�:s��1sah���<)��?q��t��4͓��$*@�R���B�O�`}�ԧ�!&!^ ��c�O��$�<�jώ f�S����?�*��ޔ6Ϫ�"v�Y�^ņ��Ç��d�O����ODt�>OX��<��On��F_,@�p�ڕ	ˮ5�40�ش���˖NYԠmZ��4�	���������"퓃c�1'(
��ţ� fb�is��'Pp`j�'��'���F���74t���@�qs�ō�R��fi�N�6��O����Ol�	�V}�^�\�P����J<K� Jgt0��i���M[�o��<���$<���`����A�Yi��G:u�DԡנN��M��?A��jЩ'T�X�'�b�O$I��m�4|2�s��-Ua��؁�i��_�`c�c��'�?��?�ĭL:"�ry[�F\�v�X�sF���[�V�'�t��W�>�-O�Ġ<���s0�Il�uk�m�	0�@e1�@}���yR�'�R�'���'��ɓ&]�!ȒM2e��d/�:,b[,w��ӪO���?/O��D�O���J,$J +Մ<n( ��R
hE�6O����O^���O0�Ĭ<�� �.��	з���Ԉ�>�~캲M9P��6S�t�	Qy"�'���'��q��'4�#��/_h
(rOH�`x�nh���D�OF���O��4U�T?��i��K2���n���@�X���ۑ�g����<���?���f�y̓�?Q�B���$�ܿ7&�,�$�ÀL�����?1����!��O���'l��HP-1�f�k1�X1C�H��sض(\��?���?Y��I�<1-��d�?��3� ��F�
�U*pTl)��oӄ�<MZ�C�i��'���O�Ӻ��,P�n����D�Bff`��!ۦ��͟h�f	i����`yB�i�ZD,�s�R#S����Q�4�ք��rҘ6��Ov�$�O��I�S}2S�0"b��9�Y�sJĢl�qs���M{B�<,O�Eȓ�<���?��A�vi��c�G�j{�#�S)�M����?a�'��x�]���'/��OdYsA�������L���XaAt�i-�P�0Ksf��'�?���?yA�ݢ��x7��a�	��_~ϛ��'O�r���>�/O\�$�<������{�@�#s ۭoR�x�d%Xp}�.�:�yR�'�R�'���'d�	Lg����L77fM�O�?Pg~�Q0Fɶ��d�<����D�O��D�O�UR#��C&HIF,��2�Z KW��,���O�d��"���OZ�	�$l:F0������VT�eyt�	K�	�iW����'V��'�����y�e�+��c�݆(�F�g�>W��7��O�I �*�O*�D�<� ܫ/����t���Y(B� yW�@$J��1A.�M�����Op�$�O�|�2O��{���F"E��� )�eF��0G��?	����$�$�n��O��'A�􌄼(� H�N�*%Qa�nʴؾ��?Q��?��i��<aO>��O�@�uF�'�%�&��l���4��F#���l�� �Iߟ@�S�����D���K{&hr�AKw��� �i|2�'J�싚'�'�q�Ľ�@?��9(�EJ@
r�i���HR+x�Z���O��$�'��	��x;���(tm�`�X7y <A��4r�������O���;�t$�
:*�ր�aO-S8V6��Or���O���u
J}[����t?���!(����T�� %��Ve�q}]���V$%?ͧ�?I���?�p荤tD��/+`�q��� ����'�"tk�C�>I*Ov�d�<A���)H�s��3!�9F�
i�GI�`}�F˫�yX����̟�	`y(�=O��뗊A#?��-�m�R���s+�>�,O���<���?9��Q�ѡ1��N�r!���
/WD�2ŀ��<����?9���?������-��<�',��p�"��,0��,�7��"�ޝo\y�'N�IܟT�Iğ�hr�}���b-Ш����	ڡL��16�� �M��?���?(O���f���'�
����'��m���E�m��1�F~�����<	��?��%Ը��|nZ r�����ٸ7u�� �I�+;�n7��O����<)s�P9��ߟl�I�?㇫Ä�uꊯnX=W0�D�'��'�b��yR�|Bԟ���@��z�����n	55�dhxw�i剱O�i�ݴ�?���?1�'��i�}I�9n�x��/	�=Z�с&x���D�Oz���5O���y���7z��[�AUA�����J�����wP&6��O���O"�	D�I���'��>k�<�4̏! ���2Ƒ��M{��[�<	L>ُ���'¬P�F�g�>q�5�H'ɚ��pÛV�'�r�'1���q8�D�O��Ĳ���gHŭ_�>U�K�,y+�I��z��O~�I���u��$�	��RA%�?<��t�E��X�)�M��&�D��דx��'-|Zc�P� ��RV���d�t���i�O�ikRC�O�˓�?A��?�.O��pǥԊW���6�Ru��O��]]��$����ğ0%����ğ�#&#�g�� S��M�~�0��Y�l�V]��pyb�'��'��ɪsZ��ОOyjDC �P��X�q3���*2��&�D��l�	�@��9@[��+"��gm@��}��e�+e~��'b�'�R_�lB�&�	�ħ
�&�`3ݪkh�CI94p����i�|��'iM0���>y)�:;�����L�_� Deg�ꦡ��럘�'�Y�=�)�O�)�z�? ��p�,)�� qFφF�,q�x��'�U�eb�|�П`���a\�ݮM�`HV�'pH��i���9o���#ٴ6�ϟ��ӂ��ɡs�ѩ���>$�v5⅀\.!k�f�'��)�:K��|��	u�z݊Ҥ��"9B�i@�C�F)[��6��OR�d�O�iNS�៴o�u�b�1G�Y7-�D9�֡�v��Ve	;���|��I�O�U3T�QG~��C�;��0�aզ������I<_8���}��'��D��>N ����C�4m�W
Z(;�F�|ҌK Qv����O
��O :b�E�b�FZ�ż�l�<�(R��ē�?1������@�2\����G�c�x�Ch�Q}nB7�y�P�<�I���ICy���#EZQP�n��y�he{Q �tl[��5��O��=���n.6Q�g̭;��K3�sS�S�?(OR���O:�d�<�A��>CV��J!Yx�bؽz>�"DOZ"b7�����F{R[���I�����0�
�0��M��p=�e��OT���O���<�F�� 2R���р
�W���X�K�'�~�F�D��M�����Op��OY���i�xdjE呝�()q�A���Pش�?�����D��W=��OC�'Z���՛E�J��PG8�r�)�(LN��?����?1#G��<�,Oȸ�rF�?�"&���x��a!�S'ThJ6m�<��%I^��&�'h��'1�D��>��R� <��h�8A0�h����lZğ�����:�	"��9O��>QC��Ԇ$�p���e��-(�|�j����æY������I�?b�O��z���{�j؃�V|��%���i�b��'��	�><��*��]����*��29Xtm�3p�HDj�i���'���H�듲�$�O���=s�a5�ָth�C0.K ��6-�O$�>/ޥ�S���'o��'���c�V��d��:-LcR�w�x���r��4�'��	󟴕'�Zc�x �E̋K��tc�z���	�On�z�0OD��OH�d�O��d�<� /���h+���&J{�B1l�k/T���^�|�'��^�x�Iʟ���������E�7|+0쪠`]�Rx2�`0?���?I���?�.O��0�N�|����a		R�v,� ��'Kæٔ'��T�������ɺ��3�pu��E>"�0��*?Ԩ4[�ON���O����<I���o�O�P��>ׄ�H��޷Hf0�b�ja�����O2���Z�Gf��>��K� c����Y���ZtGC¦��I�4�'�r,Х% �I�O�I� .
��D�}�Q�aӧ#�8]o`y�_�,�Â#���4BV���Ȃp�$���G��Yo�jy(#(�27�u�D�'���@3?�����f�͈�,��\<��K�Ŧ9�'ut��P�4��'�4 W�RK]K�g��P6�p�شA�PU�W�i�r�'�2�O<,O:�d�5�,(��P-���G�Y*7�x�	0'`#<�3����*��@7`� �F��l;DqZEl�?ntପug�^��̠�'���J6��5i_NUQ�׈Ax��[���܂��#c�lt�1�1� �PaJ�v'�I��OD��A�B��)��6��)��j��%�V���cO�Z")S$JO�K�Ȅ���K/^��0Pn�%t	N-|$�D�!cS�M����%��W��db�L!.5Z�
�\�A���E�Y��Ū3O�L��� �[]��	�����՟�*���|B3�K�&ŲY�VV/� FlO!i��p17E�+��A��/ߺR������-�2�(��Oo�X�E-�&f"��:����!�Xq��?fF�,KlP�HO<��'{��'�\�+1H%/
�< ��^5�ў�F��U�s/���7���};)�0e�<�y�G!v2^9�F h{�Vy�W�_:�y�j�
�ľ<AD�ɢg��Sퟸ�O�U� F�1�~���
r쳆���>��'�!%Q!�1�b�J��Y�G5�-T�0��&�%5%��2@̟���<IcgW�c�p(�%F=D�0CL2��']8B4@��T�йh2�����K�'����?A�������Lu��f�7$\U�!W��y��'� �s���F�H-*�n�'<ʠC�O�=ͧ
�'��]�ԇ�(a*���<`౜'�*�Y2�r���D�O�˧dH*xK���?��E�l@�f��4F4�1��Xk.в���@�<; t�8䧑o*�2b>�$(�{�ѡB�ə#"�@o���E��0���	"���	8Ix�r3��w*L\����2-���ge��2�"I�r�'H�)��/���s	"��5C۽#V���NZ�L�!��29�6�R�A��|A������X�1O��dd�����'}.���IX"��hsA��>hDx]�F�'�B�O�n�5�F�'t��'b�v��	ٟ�˱��\�8��U���;����/���S��X�%RE�q��p<���0.�C�ЀA0�IG�TR?�R�V!�F���&"U��x`��F�p"��'q`�I �L8�~���?��hO@�7�Z��+��L��ӰD	;W[N̄ȓ-D���J��O�q3��9~�p'�i>���Ey�)R1UX7�\+��x��M!�DB#Avw��D�Od��m�P�p�O��D�O�L�qE>:��$N�zl|��"�L�3eݩR�|ăG˂}�0�A�? �Iɑ����a#'�[&����Ռ*](��$P-!�'�ⵏ����`��ܷH�(�Ҩ0���O���3�)�󯗏O?P��]��@���Q̓ig�Ex��$KŔ_hT����� �l���yr�v���$�<y��ڸI5���'�"Y>�5@ጴ�R�@'Pn����1O�l��ٟ����	��p3bLL�$��Τ�?�O���34��\P(����^ VT�����#��h2�j#x>�l343�錅O�I)Tg�&X�a#Q�uQ��jQg�O��}"d�K�E8袢���@C�P�<�3���!���:�*X~�@�1�I�pO<a��29:pr��=N�Z}�1��<yƉ$Up���'pbS>��1����	ӟ�fN�>�}JӤ�}� ��M�LJ
|:��P�4?@p�����<�O�1���L~0�wDU%�.�􉔓}�J�I����J$��"��t�9��ȘN�s����pΰ�n�`���`𢄐%��1�,K1�?���?Q������]UZT�[��B$k����y��'U�}b!ԗx�i� 83x�Y�鐽��'kr/��|���Y���)@�Z�nȉŀ�0,�����?q(R�F_`� ��?)��?�ո�����O�}�F6 (	ꥯ��c1l����O<�p�'+��4#�?�ea�2+]�En�c?1�OYx�t�J ?�ʄ����:N�&4��B���1T��O�����$\%��P�HH@N�S0!\5r!�$�3}�z��V�ɷ0�`�ˆ��,cd��Dz�O��'���R�i���K�F�(M���V/Q`Š���O����OL��8|N����O瓾f����O��h�ՉLC`,#`똽W�l����'��)�*O�e�	B�GR�2�CIO���c��'~4���?���,I�<,��팃d#��k�Iz�<��L�kV�a�n�'���T"x�<Y�(�%�R�Ӣ��[+�(�#H��<�����4}b�nڟ���Y�4!�LQp�Q���Ƽ2���P+��¤�'O"�'r�a�d
�l#��O�SW�DH{㥚�1,Q�"/N"��<IS�\W��2��T
i�QR	ù�����l��� _�dഴ��ЂE#Q�0x4�OD�}�'	99���X��)��I�<�sD��a��Bfl� }�0 �%P|��K<�2 $5��c�� $#6
�<Q�%�=����'�BT>�G�Xϟ8�	Ο�S���
�P�&j��8�u�cػ6n (�IX�S���W,
��$0�-@�Y@.h
��Zo�z��C	&�S��?T�K�b
p)�+��m��,�@@ϔAҴ��������bl��D�&x��g�%]����F��yra��: T<���\�U��0��M4�O@�EzʟtaӃ�F)J0�RP�Մ`RTI˶'�OP���%G�$i4e�O`���O*�D���ӼF��)��y�&t�I��Sc?1�H�ix�� �@7F��zCoG�����e��,��b<�O�L)�`Nv=Z�c��O0v�j��O,���'6�{�m�7AT<Q`n�E�ɢ�a7�yB5?,�Z�i&
�E��.���#=E�Tj  "7�@�H=�䕀gh���I�+�D�O����OD��p��O��Dv>��5��O�����=�v� f�
���J"^��|B�����v�P�ڙk�d�6
�v��|����?���W���"f\[�Ҁ��n>j����a_t���@� Q�Sf�V�}��ȓ'��U�O Sux��O7f��ϓ ��O�����¦��Iퟘ�OpJ�R�>��L���;00Fhه���^�B�'��
I�H������|�*P�|Ɯ��B�:+���Q&a�'&jĻ�ݜl�vq�шI�:^\��?�"F*�B�D��Am�@�I	�+� p�����x��4�?�*��ᅫ�d�* ��?�ڝ�'j�Ob�"~Γ#|���ؗe5�$sk�!/��=�<y��V���Iџt���:Cʉ������t�@��$��M����?�*�P(��(�Od���O���ӡ~n4���Ih(a)��� s�q��	l�t�S����'x)�6k͸g�xq����2�����ޯZ�DB��7<�)�矘�s��2���t	�8Q�PɅΐ�>6ZI��.�M�5�iV2��O��M�0M���꧂���<��9Ol��<�On����-�p����J�@�CQ�ɷ�HOh�[�'-���D��.�ӓO�#����:*j�O��+aA��+G|�d�OR���O�;�?1��FM\��e���!{����@Ǚv��)��ɰk��zqAL?jt��4�V�剽u�uzs�.,d��{��;���r�+=)��Q�A��&��d�r�?�Ў�� ��s�fԛ �HUP��Z�}H�����OR����O����O�Y�<��Wyr�^�EWt���]F��KZ��xb�'d,�cJ�YC��ap�\�o��B"�9��|�����MY�l�#+�,�U(`y�=�u��[r�$��ҟ(�����c@I����|b7ɕ"5�N��C+_e�� �@�F��́�� [ܔ5�R$�:�ay2��72���Z�wI<+5�03l����HL�C��$cE#e/���ј\�hf�ȝHӌ��h� �*E�<��d)tA�O����O����O����O����d�B=�)c�얲��8��A�W!�D�:%����aG�8��;bW�sh��R���	WyB`V�t�7�O��D�|��5nB`���߄�6}�#��/:�\����?���fiJ\����[#���S�[��7]>Y+UX�xpQ�V��A��9��!�E���V�չh7��0U�	w��z�Q.[�fR�q_��Gy҅<�?q2�i2�'��>RkNY�52��	��僨L���	�,�	��i>F{!%2�f �9lmt=He�X=�0>�T�x�־3��@�;_�r�2H���yR��.U�7��OT��|�3���?���?��X��Cp�$7��跠LQ�ZA�oD�8ɧ�)!��O�	��^h~�E����T���[�0����]�)�矼�S�G:�p�(P�\�~?,�x�-�=�zd�I�<��͟�E�����Z�D\���t�3BPYϓ�?��i��=[��E�9L,����"ΕEx�+<�S�T��5]ℍ[7�P Ix>��H� ���D�Er��2� 1]��	�D��4;!��Z�e�@ ��ss�H��ӏO�^B䉛FU���G�^���^?t^B�	/N=�L�ji��8�R�ئd��B�I�0R������aSf� �c��цC�IY��'e�>�R�����cSLC�I	^]�a��?MJ�(;��	FC䉂=�h�w�\��{�%͋^�C�ɏny���e��1�����M��B�I[�X�{�b�"��0St�
�q�B�	�mT� �	Xl�����\��B�	'6��0�2���K��������b�C�	e��0�EU���3ክw��C�I$P��R��Ą&�Rq{ժ
[��C�	}�E��@�u]�%�@�I�'�C�	!;ИS�I9��y	�C9zt$C��v�J}!��='��s�m��L}C�9f~r�`������%Be%��yTC��|�>1�7`Q�<Ӡ��C)�;y��B��x0,���\�2�9f	�)�B�ɨ6��ڄCD&D�\�J�ͅS�B�I/��m�8�6e�P�
)A�C�I�m��8��M�~��dj�*VU��C�	<H(` ���&A��A� �T��B�	�5bf���n5�)�vC�))ttB�	�M�.�b���DRbx R($z B䉡Ya���3%ץH6���F��P��C�v��ɠ�;7 v(BT�nB��0A���9%�C}�B�*u���B��[Zx �� ԓ/�Ү�!5n�B�	�@�h|8E�͛F��2wb>m�B䉡=�\8�v�ېE� Ҵ�V�(�B�S��\8��^"�D�Dd.��B�	I$(��/�}�����@�>
LC�I�zH���f������/D;D|PC�yUV�� M�6�
D!�0yTC�I���(�VZ��,!�c��� B�	�L�ҴI�rg^̹��GژB�������L�#�B�%�.#nB�:C^.zU
X�:�+�,ܮq�TB�V,�ȃM�Li0�R�dޮC�B�I�b�6�3�� ~,>�p2�X4��C�ɓ�N�OV<i�ݳ�ԥ	7r�'R�<�c��� D�('����жFV	 �P<h�"O�H���Q�Mx~=ӣ̆8`�f�9C�'�
Ś�'�� �3+�y8��;/CV+��b�3ud�y2�?|OHǦ{��9'��j�"�N��/F�!�9>��!Y�
O�Ȑ hC/�$H:��V��z���U�$r�ɦ��H�p���	��SM� �^Q�bj�7z!��",�L�K�dK'��u��IK8h� ��;O�UrN��yB��
#��wr�Us�/��BVb���6D��Pq�A���x�� k�f\rpm�O���Io� �bd�GW�x�`($y6��$�*��Dm���=�!"���y�hdlY(��˫[h����9�,@��Ȇe(<	D+ݣ� K�F' �, ���i�'4�Yz�'
�C� \mܧ=��%{���>�f�a��M�\�ȓ4K�TX�j@$�V\y��_;$}��'�d���&�_�S�O��XS@!H����A��sg#
�'W��i�M��pX����Q!(*B�C�y��Ah�Bԅ�I�}�8sqd+u:��c	�
'&O�u���"�)�)ߞ-���C��o�v@�F�I^���`��Px"'��$�2�P!
I@0��Γ,��'�A2��޳��d&	C�
�=a&+@�2�a�8O�\��pA�n؟h��DFnպ|�ӧ$`��BE��:#v�hU��7^K0|H��	��O>E�TΜ:x���h\?J���2�� ϨǪ�������'�`�)�, ?X|��lV3�����)z2�'�M!��˛����O~��f��90 ��Nn�
>O~y�dÉ#C✀K��� ��> ��3���C�&Vz�(i(#垽(hԊG&N��2��W`7�\��aX�΄'/�H��1O0�x�Ӓ7�<x�;i��!�&֟����hD��,j�D��-���KB��K��$#��U'�����(��W@H�;c�	~ |h�wǙ*)
B�n	5�`:��/Mv���(��|�4�D�%	�#h�j���"V�� ��oӐuk��'�>E�T*L�R��S�	IW?�'&��4�ጘ�-C8���;!��Mc����l���(v���f*&�l!r�O�U<�ǋ�;'~�
�3}��E	�9<���w�ד{)���&��ʧgwR�1��h��y 6 �2L�`ٻuN˞e�
��|g���e	80�"<����_�'�E���;MN�12��#d.��I��6e�(���'� q�-^�UX�(a��f'�)�����c7� �Y�R#�bl� %s��y�(\�1�2}�oW�?�Ӈ@1)�ǍͰCp���_�[�4�b˃ E�\��#�a��6�(@��?�S�
���Z���?Q��U�����3��<���`�)~��X�w$Ю`����G(&�)��ş�. �ޡ��DBqI����>$;�� 6�O�IF����rΟ�̹5n�C��Ւ7
ٻ\c���.Լc��yDN9#���1�@;)jB���O���
~�a"E��V0)0E���MS��_��p?S�T	~�d��v�$O���G�Op�H��I-/�a�(>��5��82j6�
�?�i��	 �C	m�����G�}�ĩ�A"%�O�)�F�.V���i@��A��&��-҃�� %/��$����5�O�C��ұ�OTԽ珞�W�Z�k�Lݬ.�H���	급9��c/:��������O����p�,*(��et��+��I~?Ae�4��)��Oy����V��rA�Rd¨Nr�ZQ��*�nt+�'&m�&�� ��U��!�6�����N9/���á�P<U���YW�"HDĔ�B�\��~b��G����QX���'�4� �y�[�p��A�A�:zAA-O��������
kB���#F5,�@U ��'��`{ ��w�p`�E�#uHX�d��8z���L$��V�E[��+C�O@� e�)��O����e$��Hhy���R�+� �
����x|���X/�	�$����OPv��҄O4���(gO�_>X�:m�J?���Wx����Ŋ�A���$Ż:�^�0�cɋ?|�P1۹p�R���+������ U���	������$ʶ}}�m�u�]cb��J� W�ׅ̖=��l�q�'0| ���Fl�ܠ��� M�	�'�?i���-`~|r�¤��?�i��A-3y]�Q����21}�8&j&�O������⡈��s��ey�O�.q* �5]��;�R�����P XVt�	�l/�h��i�!Gf� w��#���kr���'�P�T�Ԛy��E�ȏ���k���O��6��x�cY�1����d2f�a��'Kb�3�.P�d��0�˟���vf!E���Jq�?ߐEo��/.���S�� ��$���~6m!��H���ɜC{��Rp�H�W0��G���9�oE׎���b�x|22�؁y{p���
R���D��,K�f��h<+%0�{� ����g֋N	��S��'p����ȏ5P2����F'~�\5��d֠��'d,�1`Y�c��A����|T���%��Ok(��`��z�fN4z[1O��:QboӶ���(��!Tࢼ8Uj_�~�T6�2����Uv*j�/C�r�Jd�T#��zQ����B�2�%�Pӧ�^���P��� |���J�^�!1#Jj�k��^)=��(���8R��Uũ��F_�Џ�$�?(�a�J�g�A��b�5G��O<����b��s��%H��I���J);�i�i҇���_}h� �"R��
2!��=x�X�	˓Z�b"`J@9M���A&L�Kr�Yt����9��M9 J����!��e8q��/��C�\�֧�G�yG<�+L��5�2�b�B�Ȝ=1t
�"m����d�C1tdZ5̎�`�;���Z��>l��ȑ�f�h�bV�cM��BZ��	�yxڭ��@#T{��R*W,�ᘃ�ͺ9�	c�60Q��XC��b\�A����%���aa���DZ�Q`F��m ��'"��@����۠)�Շl��Pw��9u`\�Ծ��P��[��(��r쌣z�.Xh�I�:s�4�Ϙ�dզ�#!��
__�7m~����
�||��,\�2$$Q�I��	��u7 \jJ p��Y,O}����jE����á�'���bU�A"�]2_ؘ;t��6s�
`v!�(�$���#'
i2���FW��K����B��\
"z���5�� q�� ��3Kx�jt�#�yʵc4�8��]2�� ͺY���ȴx��d��X�pj��Z�.&Ţg"Ä%~.Rn���vhB:��I;d�Dh@�E1(�P4c$��jֵAD�&4z��*M�f��DՊ ���Ϣ0��ȂG�ّ;�`�Ӈ2y>p,���84���`y��!��7�<"�=��M�w�����]d����c~�B�HH�=�ɜ?6���x�+���*�?)U.��v�S�E��)�W�E�+!b��V�ɵ�(���N�V���8%H�Q��MW	,<�-P�Iމ�	��y���qP$��eȢ��?�i�m(�n%~�PQ3�%V:F;t�;��5��.a��c���m�	C�IB����	ܧe:
Tc�ɬ$�Ot��̦KF���`�:���DG�*� 9�����(�FC#����'
D��$��">�452F�~y�b"�d��|�OD��˝�N堝�S�ۑ=�i�P�'1���Pʹ|���g�&I�D����cǮI"P�I��<��¯��@�'���Ƨ�6H~axF	�?����Ё�+���ʉ�~�����G^�'ܮ�@0�g2����6�^H˄J@u?�hBN͒��ha��5|O�-[%`�%��L�0��z�N� Rr ���0���\�l+��[�s��	��ēd3���j�-!\��JT�nK:�D{2*�,d:f�ضM[(�v�ѯ˲�~2�X�(�h��"M�G;B� �ڮ{��d����h����t-�
�2?��\�d���▚r�d�*Fh��ҵD�),�n�+�CV�"f!�� ,�Sx�)AѭP̒�]	cqV�# ��Iܓx��B�'�>���m��Vء� \��x!rt�S�[��G}RH�=z����$����k�!�.1E�ۭgt���.)1�@M�X�'��B��*f�~��-��.pH�;�:�ȕ&�=F���xW�1�:��<yS�#qf:�������a@��o̓q�xЃ1A O�X�%`K_�����m Y�E�*S"�:��ݘ?�����(�,H��-�����	�{}���ӷ����M_���'"�;����×�������D]�?�z@�b��cp6		PI�$��5����iFjqy�o��D}�eCM�b����N�;u65�͇r!)�)�O��f��?��E�5��(���zg(p�uM�.����6% 2�#S�%2�����RA���Փt�H�A灉N-Q�l#l+^�P<K�4\����
�O:D#�����`dR0.B�P��dBn��R��SR�,A{D��M�1Ov���-QR,�WV�.J@���x2�����T/�:=4�!�P���'~:�Ҏ7_�����A*]�Yp⯓�om�p�Q��..�� �L1x���K<-�|E�B�N�`E��( ��ц�G�j����j��K5"�/.o�I�H��a,��D]1+?X� wl'C��Y���YN�.��~,�Y�$'�X�Ŋ�W΍h��R�"�L���,H1y1�'O.�(�����P� /�=X���V�c;�ī��A~f�)F��&VKqO���k�e5bم �>�I>�3)�Y�@�&n�G���3��w��n?7���xr�!�4/b�OX��OZ�lT,Ei��=?�Q���	*���
Y�Y��h,;��ԟ&�;ga�nuʙ0�@�|���1�hҝ3�&��R��)SA���	$�=����^IH��#��Rp�A��#zk��⑌Ԭ~r�\"��O�3��������*!h93K]���#�"O쉩G�U�:��q�H�=�H����:t��
]G����l����E��ا��`g[#9������H
u"�I!��~��EE�L@�T����CTE��	��J���b�A�,����5LE4�`��0��#ʓ, �U	��69��H6��d{څEx�d_�p�XA�A�3�r�9�d.�?�'t�$1�l�+�����=*tY�ȓܠ4Qa֭��%8;J��8�Z3u�f�xe�KL� ����ȮC\�>��?u@����:�X�@��5 "!�䏌L�Da�M�1��-�G�ҏX!�Y�u���7��%�z��E±Z$���4���2��A�S�����D�7�yb@̖},�m��� Q�ꑪC�E(�yR@�1 &Ű�UF���0��H��y
� �5���)~0D�ц�A3u��S"O��X�-ޛ<��۱"�"DW$Q�&"Op�ݸw��%�/�=jGZ�X"O��� ˉZ��IHTϑ�EH #�"O��D�N	?��A��.!Y��"O��j�c�l4��-�5V�ec�"O\H�&�߮e1�c�W�;䦉cQ"OI{eh[�{L�҆�(���"O���CO	� �����/�0i�Ÿ3"O+#Y^L�P���U`��D"O�Fl�$*�<0�@�
f����p"Ot5@�iߟnhK�AZ�
��Dk�"O�`)
{܁hԪ�� ��"O��@v� �H�ptɗ���} �"Of<��Ǌ�8�F (��X���S"O>�
Q�Ҟ �@	�c� 30j4��"O$A��	{<���G��%vC�"O��Bȇ&(��C�
;Gm���"O��*��E
an�t`�`�3b(�A�"O�h��&Ջ]�dKք�C��c"O��2��=��U��-ހ})Ĝ�Q"OB���!�3_J��K��F���"Op��3��G2��q�Üa-Z�"O�	ゆ]LW&��ၐ~.n��"O,3b�ؐJ��e�t�Q�_,ru@�"O9x+:�=��/ݱG�c&"O� ��"T:;�ڤ2�/�gҁA"O�2&ET,W'� ��olI�"OJ9�g�Է.~}3BGӌ|;��ۅ"OA����))2��cFA�e~�ѩ�"OIg��/���yǄ�Vj����"O<���i�+Z`�"��W�u�"O�go�k�n�+ԠCt&>Tx"O�����E�*��Q"�YXc"ON!�5F�(}��C���w�D�T"OL�1�fMN�h�#������"O�P`�KT�\��r��ąm�p�"OX���" �|�u���Y}{-�"O*��f�ұ4��!!6�KT� ɵ"O����È'2m��yP�	'r+9�"OX�j�ȗ?`�ɣam�$4�T�!"OtuzѬ�Zwr]k��S5�� qe"O�8�â$��A#A|�p�s "O��!bͣ�V=�G�ǵ�Pԉ�"OqBK�r#ʡ�挰X�N) �"O�X�"C��J�JP0�g28���"O��S4#��k\dp*e#�,-��#�'l���ߜS�p��N��k�%�	�'���iL1�j�k��N�xO��'���FتC�tJ�#m�qJ�'r `�d@Lq
4�� J�_H��'xT�ƂZ�[�jp! �(�)h�'u��Ѣ�
D�8H�Ʀ�)�t�	�'φ��t	�-ۢ�sl͛y���(�'� ������D���#�c�j2�U��'�tU%̆ Hb�iq�]�b�by�'���7�
!&�Ic1�_�i�
�'� l��Z��BσZA��'_r���Y,(la�An^�O�L���'��3�G�U�,q��L�A�*��'�`����&/�-�g��\	�ȓtʆ����դn^�U�X]�9�ȓ.zv��Wnr���`�U^�F���gE��OR	v辑��R�9(^���S�? V́'�-�@-�5ƌ7~�0:�"O`��Ao
f�(���_�u�"O�8Ap��+Ơ���l@�tm8�"O�x8�o��[��]-|T81�"O61��ώ���Q��='7�@a5"O�5�sA�D�f�s�HY7;6��7�'l!�XMh��p�ۄ~��	6c� �a|��'�d�����x5���I�鲒��?�!�*-AF�-\=�2U�a_�p�OҢ=�����%B@�}��A�ѩ�C
vl�"O���� ��a�����n��SBT@�'P�>�I1 ׈Y*C��-�6=(!�L�oNbB�I�9Q��'��5|2ݩr��Xb �	l��� BT���5ʓ�O\�`��!D�����Q�T�|�`�M$=�x�0�9D�P���˨.�L�F)��j��fA5D�؃aB��@-�݂FR#���(D�<+#K�#������0@��M�S�%D�`@8aZY8�
G�re��N"D�T�+�=SL��&.I���!� a*D�<c7�q#q��*/`e�(D�DsC��/_�����vu~Ti��&D���S+Y�V�`�H����c�!D����Ӂ=�,� ���C�}`A%D�l���Ͱ��!:ӀΛQ�r�Em#D���H��s�<A6�ʼc��9��"D�dsFf�	=��g别Ħ=��*$D�9��4G�e���Yz6t��c"D�Q �-�xx��ʃ���5zP?D�0�E�1*�
�ϟ6���Dk=D����L!)�X��7`XZ�E;D�H��M�K��D(�@�>h���8D�0Xb�П7*�����p$�!��8D���祇;_�� � �ӺK�DXAw�4D�X����:˨D��-_�;���&�/�D1�O����:;aq��G5P�[�"O�ɣT�R8�n ����::$b��"O�uP�J�9\{tg�24�j�Z�"OX��1T��}X�&����C�"O��c0���R�P��N�Er��ز"Oh@*�`U�l=����'_**�"O6x!�Z�6��3A�O��"O! piT7i�<�J�Ao`��9B"O�Y*% �0X|��C��
L��w"OR��� >RY3b��7`E4���"O8�(v�<mu����g?j9
�9�"Oĵ���ʣaX����`�8f�vx1E"O�乕bя"��3��ַZ� ��v"O�٣`A�r/j�r@��5Au���p"Op�;ҠT����"�2F�N���"O�M�AgT$q���Jv^H���@"O��o[����C�'���("O��yF�.�t���
$y�0�06��܄�	D.���a����Q��5D���DÿA��H��#��[��b��/D�8Xӆ	��L������R�#D�ਢ�Za\3��Hn΢�n D�)V��3F�Z�qqG	(4$���9D�ȂҮ؜R&P���ѱ#�aK�&%D�P���
��RTsB��e��A�#J#D��	'o.eoB8���Ǜo��c�"D�,�G�ĨW��(P�ƍ8r@Ãh D���'�b�,�����=���L2D��Ƃ��|�� q�Bչ�L#D�� j�"֣MW�n�;c���=�S "O�,��.�"\�����,�\��"O8��c�9fe9��Ño8��"O6�Y���E����5&K5i�h�HB�4�Sⓔt��(*5�Ɉl�v����E�B䉥%��0 Fl"u�^�-d�B�I+�t�r'�h��k5�ܢtw�C��	�h�3kʪG�銒�Z�}ọ=Y�G.���1���\B134Ά-��p$��F{��DJ��0j���	WM��R���y҇��u0�t���O��H{KX�y"@�8c��XQOڍrFv�$M�)�y����$l��LF�ZxJ��s���ybfT�h"��q�{^�l�	��y���*wh9C����^x@0�EI��ybE�1D��YS@�S��4��AR��y�o�9"
(�ve^�a�&$��G,�y�h�2'���6j�ST��L��yBj�h��PE�ׯL)��8�"N��yb_��ٻ�ɝ�BAB���>�y��>`_z��֫�;g�@�c����y�'�&h�u-^0,�DPӒ[7�y������
��zt�Ñ�G��y"�	7Q�!�%�yĨ���Y'�y�E�P�T��e�<���n��0>AO>A���j�� ,=����O�<&���t7�m0�-�z�Z��r�	�<!�}��d�X�D�l�������:����?��'պ�Id.�x���X����@�X�	�'�
�i����#��!đ7���'NV(��1�J�z@�}���S�'@*(�"��l��,QEC��t�Z�h
�'܈�!U�M�[�2ܪ��o?���'H,�!'\�~X�Ӡ�#mk�I�'Y$�%iP�~�dQC(g�`Qs�'��@-H�#�5Y�䈥5�j���'��lA�	�%3l���-���U[�'��e�ʴK�MRh�F���'t�0TE ����өo%��
�''D�*F������刎-v�
�'a21i�s�>E��N����k	�'���	�>:N$seL����X�'C`mJ���z� Ї#�	�j���'3�Y���\�@�l�O���'�X�!��)�v��f�Z�IC<��'*J��W�F�L�K!��M|�̫
�'���y%B:!ʩ�M!=�8	�'�d�#Z��q$�ؐ�;�'c�9`�\�^ ��n���p��
�'�L{C�L	m`��	��քJ���
�'�̵v��eN8Id��E��5�
�''�A�)�J(J�[2���B
Q �'Q̭"��>_��<��+�|��'4N��B�*!�X�A���z<PG�$�S��?����@���`PHވ}�ó( s�<9�H�'\���AQ�υoj\L��v�<) ̓!�� ��D�5�-��DMG����<1�ŏ	*1��cQ�2d��4��@�<�g�ܸ4�bc�"0 ��AE�<A��܁`K|@�r/�4H�%	V��C�<)��A�R�X5c��ښ_8�!�V��K�<�pjϖdw�L�F�Z!Q$y*��p�<0��w�d����G(+��U*��p�<q�E /�SGH� ^��ki�<� �՚��P���d�g@�S&��5"O�!��G�'�J���L#�6x�"O���FG#Yzy{V���?�ћ"O���IO86ؼ<4���=Ίe(U"O�uIr�]v�0JC-�6B�"O����Q��xx��i�w��"Ot�W�Ά`'J��(Ԋ\Ǥ���"O�5���sX9�G
�:X��"O����gt2>	����<����"O��
�lNB���K�LZ3t!"O\�X���T< ���45��"O�Y��d�'@[�P�hZ�m����"O ]���6H����� ��+b"O�
EČ�2S�ҡJ�:���"O��҂F7Jr� �KR�|�l�"O��ن� ���Q��
�o=&ᢗ"O�����I� ��$7�%�S"O�ŀS�ʺ�����c�c2��3d"O$�)�gH�&~�1���]'��#2"O:4�Q�C	x=�� �n
$f�J"O"%��(	`H�-�J��)�"O(�h�Ā	s�*,�%C�� ,�(Q"O��9�cZ��qA\�Ԑ�
""O���a5YH�#�@�A�P� "O��S���-��x�֮�)(e3e"O t�w�� a�|�J�M	(r.���w"OlщҨP�R&��s�lܒ|�ɋ"O���W��rt���܄t�r<R�"O�
���w_>�Q�R�D����"O���A�!r��Y�@D̠/�}�"O����@C2N�<)2�����%YD"O�Ƀ�e�0s�����\����5"OB������|̭��MƎm�f� "O�h;��J:_�-C���?�Bܣ�"OZ5╘yb6��,�>pi"�T"O�I�&C���L���Jr��{�"O�}��dI��*�@���H"Oʹ����`x�5�2�144��"O�h[��_L�p�
֤)j\D8�"O�-y$���1�b����k:\���"O��$X<��f]�)9�Yr"Oz	ӷ�����k'��"AQ3"O4�:S��'%T����I�(m�q"Ojm˃� 9Rw�lᦫӽ@��eY�"O��+�'zj͸������-��"OV���-A0���TL���6!f"O��q����q��Ё�ҠY�"O�ٓlۍw�h1�%�/���C"O��˒��wW蔺r���J�Z *P"O�U��x�r��4K�B��"O��B�&��((4$߶@���C�"O�¥_1S��	9We��r�! "O�i`���5X�(T��%LiB"Oꀓ�ƅu�R0kv�+)p&s�"O��Sw�]�Yn}I� ��3Rԝ��"O�C���~bֽЂ��%r2�|q�"OD�R(Ό"<�9 �4"Ot�����@mnb�O�~M��"O����T�.O��/�"����"O.��q�[|��΁4�II@"O\��	L!6��9`�(�.œ�"Oh��ǭ�R�D4��m�>���"O>H�6d�8#�v����s���ˆ"O�p��향t��kdB-fl�
#"O� �݊�(]	8�ʨk�"%F�ۂ"O�9��^��Q0G�	�	�I{D"O��$��Bl����ؘu���"Ox<i%�����2G� S��M �"O"-�b�X�?]��X��YN�xz "O098�,c: �넇A;+l̘�"Oִ��鎍p��Ib�C�J��w"O���2�U/���Ѣ�9��h��"O|u�A �;e>�}�����i�"ON�3۫s�p(�Fo���w"OF�f%�xw���pJD� ��\` "O���ș�hr�D!v�� �D��"Ol!��j�˖Ѣ�(
�\8�"O ���@35�:I3���T�2"O�=�F�'Q� {�GE�o�^X��"O��C1�'r�ΐ����L��%r�"O�U q������B%�Q)c-,�)�"OP���O9?_\S���q�H�"O�D�@�!+�U�r)"B���f"OT�iAGr��r��9	�Y�4"O���-N��4
PM^�Z}Z�"OB��%�8JX����L����}q�"O��ȷ�@�D�p�c ��xg��"�"OޑB�j��0�F�s��R�:R*9�"O�����#K��E ��8c���*f"O>$�@�V�|\"a��/�,N�f��"Ox1�fGB<`k̑A�.��srF]�4"O���`��j�NբW�Ta��S6"OHHk�F(�� s���bx�"O��%��h� �x��B����"O|]����e^�����,)�ji��"O��%���]9��X����S��t�5"O��!�c&@Q����L���"O�e�#R�i���[S�C����"O��)"�yJԕ����s�|p#�"Ol��@J�*�tP�E�P[Z�%"O,��!�[�BLF4@�h�	B�]!t"O�4£H�(�����W�n�$"O�	��Q����a�0
�u��O�<��3�2P��}fd��-Fq�<yv�E�0�Lyģ�%�QI���m�<ACb�'���T�D%S%��7��i�<A��^�M��Xs�.ҟl4PF�d�<���X� *VĜ>u�MrԌVu�<�4y�A�'��/w������x�<�f��PBd��D����� b.�v�<����)K�֤�Mɟ$UZ|"L�x�<A�D	'�����g.����dXo�<�D�58dj���� q�����(�c�<91���&	Q���"3�%�a�<��䖲e9�D�qÆIB`��u�g�<�gM�e!����]Ta�Ax��b�<I��цG
nU���T���Uci [�<�`k��.�$��Ą^N�ʱ�Kp�<�2�Vg]0lC���of��F�Tk�<QvLն:�IrD��!yx���P`�<i����5�0"��K= 8�C��U�<A ��J�ƥӝ_2�]c��S�<I�k؈/���a��#<�I�"iMN�<Y7+��bΐ��1&�^Y�k��_H�<Fg�:�`RdB�rU���G�<�@�O�"�f�30Ύ�S�2�*�n|�<��^snRa��e��^$=#��y�<��n��a�����:0t ����P�<� ����ܑD���1���E��8u"O���%��Ut�}�f#�*�rq�"O��S���5	����"z@L"v"On@�ᑅ/l�=Zf?#f� �"O��� Ǿ!��e��#�t����g"O���S,��h�=; �I`�Ht��"O�$`&	����4�Vb�<����c"O�y��埶pu�%�C��1��8��"O�����gX+"�!C��P�"OV���ȮK[阡EP�/"%3W"O*8�Si�=h����N(��0�"OX�)$,ڪPc�٪$��'&��̉�"O��#�B�qp��byx1��"O�̎�*qnӚ`�yq!b�Z�<Q���*���0���:_���b�q�<�V<�L2e�H�.Y��#D�,ᕤӛH�F���A &܊��$D�I!���Du1c�]�T#�M!D�D�qf��7,�,R�&\N��$U�*D��:Һ��h��VQ�Mr��T(!��@�s�|�$-�5y�u[�EL�C!���
}X��tG�Hp^MA��$!�^�t�8ʑ�ϵ3Y&`j֣��U�'ў�>U��g�)e��\��`�!-D���
�2�B:�&����#�?D�lp0HE��-"w��Ng
Ya,*D�P�b��~٠ܸЏ�'2�,B�E(D���ł�@߼���܆4�΀��+D���$�@�E�j-3���*�@y�c(D����,�����ءi�(h�˲<9���?�9�za�F%8�p��e���D��ȓ�L��J�'�V��`Ǉn>,��h�`I�5cD�t���p�ZIܼ��ȓ=^�+��h��ḇ���7-�х�Rp���E.2��{ ���ȓ&
�x��5�$�D��YkJ��ȓN}HD�ɟv��%���ĚQ�Y�ȓG�
��$Ӷi��b5��Y��ȓo�L��f�
4
��x���H�z��*��C�CP���SvN�c�
���r&J�h�A¿�`I����%� -����8�<q܀MG�	v)4���	_~b�ݿTԴ�tHP������\.�yr+ݴ�>���c����!�̄��yB����r��RBnpP��1���0>9gf+��x���g
>���d�r�<�����9�g� `֑�s�r�<���jd݁�,ѷK�H8y!�f�<���V��a#3�W8@�
��!J_b��x�u�ܱ�bΖG�}�"a��~��ȓ�v �E�2j8��i��8�(Ѕ�A����?���;ąX�X��%���IB��`ҁ�[it�d׺)
��g*.D���V�4���wB��p4��&D�$I7�M�=��hPW"R'Xmn\㥬%D�����<U%���ΫN4�B�I.�O��	^X����ֺt���a#
ܹQO�B�I`f�I֩RՠHz��.N��B�ɴl�e�@,Q�h��F�B�X�B����1ٰ)� ��|8����H��B�I=nx�i�o�A�~H��i]KڀB䉣��BՆ��9#�  �.ϔ>vpB�ɒ`��x�S	�W���ij��D.扷!܆i	�`K�k^P�0��_�(���;�� ���*�lє�`��ۃV�p��"Od�Tf<������4-�Q�"O���g�^3D��0����N)$m�"O^��fZ�L��]�q���z#��`"O`}�c�\��\���dP-,��x�"O��t/��������G���O��FŐ�=sf�RVn�[-�qĥ9D�(cc��=(�M`�܍V�t�C�6D�Ps`�t���a˛g@�A�&4D���i��9�V��� �(����'D�,�P�T�E7�7�����2D���`ˊ�� �3敯{��+@&6D���DS[�d��C��n^����'D�D�t
�1nF��E#��v�I�B+'D�,"aJ:1�T���mюI~U`F�$D�� ���K.���g�ҒkG\1-1��O:�=�O��Ũ�®Z^ ����~y�"O��+���F!�B���l�B�f"O��b\r�Yz�k� %��yC�@��y�aJ6�|�	4�K��r}�E$Y�y�o���9�@	'; ۴aR1�y"ލ����S"��"6�tj��yB���/�ZI�����0�R���/K �䓩hOq�`�K���v��0Q�Eʂa
ܳ"O
dx���,�v�����=`Z��"O�X[e� Հ�C�VG��H�"O�X�х�;�bT�6㐮�4���IS�O�衡FU��������c�����'�F<Z�g:?y���p枰o��-�)O���#�O>�p�g��.�"2����9��"O�4J�ߵ
j�����i���"O� C�׎d��\���5q5�%�E"O�肢�I0"u`�)���a�.��&"Ot ��+��#̐�S'�jЊq"�"O,�JQ��7Ԍ�BƐ(�4��OV%s%)ϋm��5c�=HN- ��O��d�O����oY�M�pGӷ ,��cXz�ń�5�p�घ�}�����	N&L�@<�ȓkjQ�wOü
��ѧ&pa�g�B�<�!	[�f�ج9P ��t�H��{�<1hD/QfT�V�E��L�(b�Ly�<鰏�s��"��p���%�[yB�|���'B~�ȓ�T�}H"�1��@ǈD�	ϟ��	�;��ئ�F2��0��o�tB�	*��"�Ĝ���C�A��>ղC�	�*D��4"Q{H�)���MrVB�	�=�T��˖V��$x�/|~B�2r��:�*BhŒ��G!��3�pB�ɽ8tn8��ć�,yh�95����B�+d;��� �>�pҡ˼flB��#������
i'6Ӏd�--|B���
��MΪ궭��ID�C�!��T�2��vN�%JDF߻mr�C�IW����qӘA�A�rk�2VB�	4���0�
�#u|��)�qc��=я��?��ƥP��u�7�(E+`l��7D�<��͗t�� ��=#4���2D�låQ.	��,q�CY�0�Ę�0D��C����0�'͘(�*�k�%<D�D��ċ0u$����֢NT�x�%M:D�TJGȂ�{��*P ��cۼ����+D���A'U.<���f�5[��j�,)D�<j�ˎnyf3cCoj����&D��P���6%��dPtoR�m�� �*1D�� ��9p_!&�:��㒘Ȑ\c'�|�)�ӵ�~d��kԣ"��򱂉�@ٞC�I�e�`�Z��u<ȋ6��;�!�$ُ���S#@[�P	Is��%�!�E�+�h����ưA��hX�������<1�ɘO���g	R�w�xDY3j
�l�`�'^(xT���+�X�g�F�̑�'g��b풶=�yqg�� ����'q\���B1[p����@H�qv���
�'5��k��>����N&eB����'��=H���J���F,37��S�'��%0��f��- 4�Cg8�����O��0h�Ő���e�	�"���t7x�QA̬��#q�Q�}S�C�I������L樠[��t�
C�I1oI��ca�� �1"���,6��B��D!�����]C��z�K q��B�	�`� �z2�1Uˊy�Vݤ)��C�	�C���-�<4(�1\>!3f�$&�S�O��	������@s��=��p�"O.P�CĭU[T��� ׮�̉#`"O$���ĒH���r�O?��)�V"O��9���o׾)�.B+.
:<��"Oҽ
ƪ��_X&��("��iS"Oޘ��J7uWl9��� |�$��"Odd{�B
w~��`��H�qdd��IH�O�%���M:f^t��-�hI�(@�'sj�1��b��+'X�S\��@�'{��[uu�j9���\Z���j�'r�|�V��s�x)Vg�V:!	�'�*PƯ\-$&��RK��X	�'��j�L�
/����r��8IF���'n����ԡI�4�#bΖ�0D4��' F�I$E�v%D�@�ܯ/.X���'�Rc� ����;�f��_��y�șXsx���+��=�8�z�)��y�h<`��j K�	hBLA��+O��y�b�oA�3� ڗt����Ɯ�y⡝�]*�	Qb�݋z>�d[&�yr��K�pe�⋬p�R434G
�y2.E�/�����![�e�2���,��yR!ök��{��Vv`9ڲeǅ�y�,N�P���B�-Lq��xe�L�y��I�J�d�a�X�`x��e��y2��q�����)�
ZIx����y��Hj�P
�O~@X �G��y",�+WRP&lE�EI��?��?�'A\����2�Hl�`j�hͺ@�'4��'''���Q�.��cDveQ�':Tp��hI$�V�"`_�Vz)1
�'� k2�0���� 9����	�'7�質��zU0D�$��%�4Y;	�'+ٳdi�xR\(S�o�G�he��'�j;ӯS.j���3�<��T1�'\���IB'Q� ��$,R�x��'��5��Y�i�a�1���@��7D�dhw�W$	Fhp�g�
|� ��i5D���l]�p�	���� ��T�P�%D�88��c�^�&Ǒ��SG�&D�P�c�0VZ��V�`���R2&D�(�֌�����F)�O�z���$D��;1&�Tj||�V�#JZ)�s�#D���a�@PC�4/N)K%'<D�\I��P�"
D��4�J�#XT}��);D�� ��+4�$ny"13��O�$��"Otⅅ.bz�����@�z)85"OZD�m�H� �Z��]*Uh�`�T"OF0�sK�w�@�փǨGf�8 "ON(c���~Q.�Q���X��re"Oz�D�e5�A8qo��~�nȣ�"O�=`�斎��x�HC>(��;�"Or����4Pp�0��в��Eq�"O���#9�̺�k�~�5��"O^-��-6װ��Q�m���"O��'�_�	�D���]0eb�"OT��I3kL����ُ>ޭ���'�^�)�'L����F�,}��-AT�����J
�'L�H2�	�3��J��Y�v��	�'����D�I��yYֆ]�=uxY��'* �̰K���ߚ/�|-��')~p����h���=�(���'�09�3?�P�j����.T�+�'
��Ir�P�sVH�1'�-��'�]J�攮�$��0 	*$�*�'��P�%F-r`7�"���"O�s���D
���:VaX���"O��r�U�A��n]|����
�'w��
�F��B��+eH�6�l��'|�5g;`���R7%C&ŸY��'Ղ@�% �;)�}�V
\�^���'�(l�&@�Q�0�-C��XMI
�'�����
E�8�zM�I�f4�;
�'��e� �78�Qk�@����`	�'��`b�9b�$�(b+R�*�(ms�'��m��D+/�ʴ{V�3R7q�
�'H�	���ц v¨���^)Q��#�'�ۀ�=/m����*���"OL1ڶ�͂sxd�䗥|t2�aG"O~�����}�7)ѝbI��AC"OX�a��7;��Ƃ��"�Vab�"O�4ǩ��W�X�8ga�r$�}B"O�!��HR:ߴ��@.�&Z �<��"O��DC�J2 Y��bS���J�"O�횔$�8�D:$��@�u+"O>�C�a�V�69r�hڛO�d�!c"O�9��lK'<� ;�&�%uj)��"O0E��o��>��MAdf�_�h��S"O�<E.�%�b���Bêz�&��q"O��B��Z��H��
�_Ypp E"O�J�C��q�q�~V,]���q>5�� �8 ������.ڠ@q�L!D�P�u�Ĉs4T}�v��
7�h0���!D��8�+R5p�X�����2(��B;D�<ӥn��"��媗�kdq 4J5D��(F�Ʒ$�	"¦��1�:Q�6�.D��ኡ+.�5F�!h�&}������6��2�R�Q�ʖ)X.XE{��'h?E�CEׁY/0�`so�WDI"�2D��`�̃	Є�$�M!a�q��9D��� ��"��Ts�
�*�ᓁ�8D�D;U(�
�2�,P`�P���,5D��C�E�1F�����;WYh�k�j D����H�?
<}��iXJ�s)D�`3�/A��Вn���� `'D�8�T�ʤ!��Մ6������7D��Ar$X�,0J%��V�H�Z��#D��jE�L�t��
SF�F�(�"D��+T!�o�B�3�Չ$)�����?D�� �AK!''bt����
��S"O^�Reꐖ��"��ץJ�Nh�T"O\lR���K`|�j���Q�K�[�4D{��iޖx���l��Ӳl��S!�d�I��C�INS�4���9:�!���q��%�nB�4Z0P��V1g�!���zڀxૈ,q�)x��Jw!��N$yb�'�`��ݥ,M!�]9>�<���`�hʬ3#�9qK!�$̂|���@4��
~xaRt���!�$�8��F��
f����F�>O�!�ǕI�z%8�oZ�	�@�Hu#!�!��	 U�!L/x��� C#Y�!�]�"��t9Bݎ3y��F�.�!�$ј.
��S$l�4�Б���&�!��8)�$��e�4_��9�K�4&!�D/?�ȱ ��T{of:zE��"O"}1	.p �"h�=5p�`"O`���M z�r�Q/:MJ�"O�)B!X%��a����;? |ae"O�0�l^�X��͓B )}��XV"O2���k�����~b��[�"O�<;�5�2pa7 ��7R~��"OҜ��M�O��92���$މyT"O���(.3�S6�cs\��a"O&l�%Ș�|c��sg��8s�(��"Ob 8�L"!<�Z��s>=`"Oށ�B�C�b#��;�?>nV��"O2(#TK�6I��RGB�k<=��"O��U��0G��Hɰj�r�pYx�"O�U"S��9��.�bL���c�'�2��@3TNʻ��EZ�F�mlP��9D��;T�#pW&|��� p�����n9D��
��L��4"��.�К�1D��ceV����� +�r�SG0D�������,�Ӥ��3�`\j+D���D�=ah*ґN%INd��'D�� b
RZ!Գ3Y�.�>d��$D����� �R|t�+�nO ����5D�x��G@YH}jA��T��؃O2D�D�b�^��<9���)fWĈ�J5D�`k���,�B̀ѢP0?g�=�q(D���QT�t����0��!|��)�Eh%D��(��U�Z�۷�M0u��J�>D�X�$n�J8 jV8�x���(D������� TpFB�c�(rG(D��nª+V� �TGd�0���w�<A,{�ʜ��ct�����L�<�s��8��A���"��PmG�<Q!+NDJ�8W�-����hBi�<iw�s�.qqd�@�h��#��@�<�a�(J��1�7N�s"��RFF�H�<�c�^�� 8�t�W������D	N�<)S��0g$]����&�j c
L�<�%�2aP�����A+Б�%�F�<!5$ {��A��Ϧ.�!XĤ�B�<g�Ś7ct��f)֟bh8@��r�<aO� Z����E�f��c'�h�<�5�жf���¦���2��P��<��+��s�8y҆"HHb6��lz�	���?�~��]�e��&�L�2 �.D�4! DN��@�&n�1�B,D��Z!�Z�
,*�[.Y�:M�,D�PPB�Y�B+
e���)st��r��=D�� Ľ���
��XY1Έ4�l�pw"O��{��� �x�E`,F� A�&"O4��J�!NDIy��ъ_���X�"O:E f��0����"� T��R"OtP���1rE�5�E�a��y��"O>=��͎4Z�xү��	w�H�"O(Y��7n�z�Ba阊0Yz���"ONXK�!��PJ�G�N�2u��"OZU��N��^H�!'ZW���z7"O����k�y)�E��P�l{$"O^,;�ș)��������< "O����/S��Ha���A�P��ݲ"O�@k��e����_&�H�W"O�hS0 �wG\���G� ,��"O����Hǲ(�4��f��"��!�"O4k!�	k$��ĀW���#�"O������3e�±����3�~ *�"OF
�@ V�P)�$F��ҴRp"O����	ů�>𑣗�d>��B"OyX�@E�C!� 8�Ac7m\��y�-V6�����$Yl�O`�C�I�^`v�p�	�2+���Jůxx�C�I�C;����NV�#�Р{Ѩ�1*֡�D�8e�a�)�*f�Ź��0��'�ў�>uZ�喊Ȥ��C�^m��"�3D�XY�I�`3����J�VY���Qj3D�4�k�Lg�h�d�?}�4�+��>D���o��8 ����)�,�aC(D�pU�%J.P4�c��;���4c:D��q���Z��SA�G�8���P��*D�	���9R� 9Bƅ�[�5���<D�p�b
�\����F.Z�A�O=D�t��eX����*)L�4��$l&D��ئm�0q���%�̴�"�#D�����_�y8�'*�-s�&7D�������pd�.�fu�c��6D���g�@u����/T��q��2ړ�0|�H�g���HUiB�;\�M����X�<�p�N�H.�t�Q"�f�>���eZ�<)1��X85���VY�ꍋ�OWV�<��-'-���b��O��`�
�y�<�4h�~��E1@�V�n�иVH�x�<��K��g�P�FG�=� Aց�u�<��Bj��(!Q��P|�#��l���hO�'r�m�ѡܴ�joP��D��=�l��b��;� ��C��)�@�ȓ6�x����
*|�llٶ@'�2���~H�T�E
�D�*�` �Ī8��̇�W#`�`i��ep����"6��ȓ7�>T�%�غwE��ѰK�k��ȓE>IcІ�:�h���"^�H��Յ�Ie�'�� �%K�z3�Z�o];d:81�'m��P	#8M6�p�Z&_�d��'n�[0���8�4� R���
�'��MB��O!i(��
���H+O��D�W�d��m͢]C��ɥ.�!�� �}ZQ��0��IѦ?j!��[�'^\��v
�e��i���N!�$����e��8�t��Bd3�!�Q+����d��t����W�Z�!��6:�H�iuhC����:�U�2�!�d�K�F ��� .���]$DK!���kB�hs �����x���f!���u�� �{��i
�O!�� 6<����.ޖ���/��n���B"OuIF@%"���zS�5��"O*p�C��v`�`�A�θi'"Ou�q�O?:�&��$�H��(�Y$"O$q��ZR�촐6
��z((b�"O^ � `(۶�H�W3=EbT��"O�	
U�HX6H��0i�E��"O sr���ʲ�b$ՒO(H�9�"O"�q�����4��u�Ľ|#�JB"O��GD !���Y�hN20"ʼ�"O\a�C�O/N���NA�3'Bl"O�9�%ۮ ��9���ND)!"OƐ!bą)L�@�ju�̓;#R��"O ����E �
�aw��~4��"OT5�B'�3%��ᷥE����"O¥�­�5Ɓ1Ö(wV�=	w"OF�!e��r2�#���0VD�r�"O�h[��r�m�4��%nTj�"O�r����,�(c!���6f� �R"O�
C� z/�T�J\aDY"O��@�U�k���0JI�&�(��"O�<�� ���h��	^`�t�p�"O-9��K 8(@=a�(�G�8��"O���SF�1@O�q���<:��"O��(��@�r����$#�5!"Oz����
[|��a5c�'�F(r"O���/	�c(ֈ�SK�;#����"O8�;S�Γ;�^��T�>T����e"O���5���K@�\�˅&4����`"OV�aԺ$͖�kb��;[�����"O�}z���W�:%0C��2�^��4"OfY��۬~,fQ�X� ����"O� T�Dy��i�N�4��"O`��(G7�v���`�<���B"Odɠ�Z�F9��JTa����2"O�`:'@ڕw��%���A�K�:��"O~�"�΅�	#�z��ּ-}�0��"O챋���z(8�V-/�F�f"O����,ۻ1]��్�i��p"Or]܊P�8ҁ�S�TO���"O�bю��L?Ɖ6	E|���"OB�:������2>�I��"O�ܳ���W0�!�41+4X�"O�I�`�f��
Cޚ{x�4h�"O���ժ�)U0�ɲ"�خAP��q�"O�Ds�jB�fL�u�.�1:�$ht"OR��� �\��m��L�CCv��"O�	���^��yi��h��4	�"O(!A��e�H��v��_��p�"On���z=rh͛��z3"O,���W�h}7bA���$Ч"O�8@ ,|lB �*�^�J�"O��m��QF�z��طz}�XQT"O<�v�&`��0Cƕ�b�="O���!�<$8�eR�DZ�v4��"OL�
��"�̅��$�� ��`(""O�lfM�.U�r��Ӄ�#Et��;�"O<I��*کU������eh��b�"O���Ϗ?4MBA5^~�x�"O���*E/#���iЯϥ!o̍[�"O��3��8Ej�r4�7
x4%�!"O`XiG���u�	�X�cQ��t"Or�����$�.@8X7��A�"O�P۠/�@Lx(s5+��	GF�R�"O� :�3q�T2c�X�GL�=R�֌�S"O��l�3w��zV
]�k3�4��"O���FW�I��ke'S��z�� "OFP3�OJ���ҵ&����i�"O؉'�P�]Р�����r�"O�� Ԋ[8@`jTJ������"O����U$���A 	��\�z�"Ot1rJ�*1�����G@�1�6���"O�p %�^�N�C��j�`�o4D������u�v�sA��h���kA+#D��;�]A��v�ĮN_Bu���Oh���OT�D�<�|J�O� q&D�S�\3��:?��("OAQ�8�d���Q:D�z��c"Oą�1fJ�nPQ��(7t4]�"O�����I%k�����\$t<�T"O�qB��'	�P:��K%vr��rB"O�]�󨏮H��<��l)\Q���B"OBY��i�( q����P�Cd�sq�D2LO��#���;f��#���P��G"OrlAwȍ�[���)R%J$:���"O��p#�a��(X֍�ݰ�c�"O@��#R	�f\���-���pW"Obx�f'�2r5��Rv��F�^���"O��fl:}|�`ѳ��R"O>ń����掋$ ���e*O��2l	_l�w�M�2���
�'���G��;��	Z���$Y�q��'��R��ɦw���Y��[�#ZT��'�r\���ɉ8�<���/�;c�<�k�'��{��8/J��Ջ��\ڜ�Q�'c��H�]2q���X�dόSiX��'><C5_�erd��L�B�#�'�ҩC�#��P�*4nW�	�	�'v����/
_xĸd!ޅc�Ը�'0t�ԯZ&r��@�'ɴ'��
�'��0��!�z�#4��&IxB	�'IV�P��<���5�H��ǢRK�<���ǏSn���ջ<Hxh��	p�<��O��g�@��O�0d"��3�̏kh<���ۘ. ��a�ZX�u`&���y�R�N������XByAam��y"(T��Ί�7�Ε"���y����ca����dE*EIؐCC��y��"Pݞ�q�S;#J괺���y��h8����D�)7��0���y� W51H�Aa/'պ8:3'ۈ��'`ў�'�X�Zf�D5o��=2M9o�,��';�p��[�5��XY�J�>j��H�'��XÑ�6KE�԰�O��b�*,��'�8wa�&/�N����"{�&C��.���o�0�6����^��C��B�0H��E	lG�pfG��jfZC�I�դ�����r���!&ER�1��C�1IY��S�j�8�|t c �)!M�C�	�^�lC���y�V�H���#C�h���#���)&d���C�	)_��%�C�.WNP8��4>�B�	�`c>�� �S�Y�&�x�jƃ$�&B�I��R���/�D͘�+C�%J.C�	>e�<����A�%�fUJ5�L 9ʼC䉫N\��(�T���0�(ɴ M�C�	^�*4���XKpaӢ�G6NB�3�T2�"S�t:���˃l�>B�ɬ%
���1=�%a*�6r�pC�)� �!�π$�r��l�6����"ON��R�<X�m"�M�EN�!а"O�PxGR�^�$��TL�dh�L3Q"OL���ß:-�"����ӕw�0��"O�S���*�.��G*�7����"OF�ˡ�άHS��1D�:,�!�d��x�XA ��)�� ��)�����hh{�n��S�B�
R��>C䉠D޲Dɥ�N"f�ʕ�`�A%��B�:��1��$�Q�Ԕ���Q"��B�	94�-�Ư��l�Pc�nO�mvB�	�o82�w��>��d����0`�B�	6H}Q2C/�#t���g�
K�bC�I8���B#	QfސX��J�1�<C��!6'��fO�@O���� �u�dC��_u�,I0��\˶D��È	c� C�ɎLeP�ڶ@���w���z��B�I�T0�惁~��,1�"�
T��C�I4$a�oLF<R���K�|C䉳<��=���"��Hz�Ŏ�czB䉦0���jf�F5G;n�R��
u�C䉱g��P�O�*E8!�S�٪E�C�	�[�����J��"f�g�(B�I:���SضB�� ��LR.
B�	�m�2��_�
UQ�T��j�B�	2n�v�˲�s���BOî=G�B�,K����p`��C�x�hC�IA�NTAg�&;7(AI/�-g_6C�ɝ��g�Is�$������B�!���RE��es�$ZFd_�e�B�ɒzcĘ��k#p�A�E�[�ܣ?i��)�0@��@څ.�Q߀`�Ь�%=!�$�<C�8UZT�P�g�"<��kƣ0,!��~�4J�#�67�x<�K�>!�[�dz�3�o�) ���Y�ʝc!��� T@jc�ޖL'D�x���9�!��b+��ʗ(�2$>�؃%
ϸ1�!�� 7΁��'�|s��T%n�!��Բ�D3��P�}��'(Ćh�!�D�=��cգTb0$�!��.�!��=x<a�����r/��C& �+?�!�$ҋa*��
�ڲ~(�R� �(�!�ĕ�5�fd
���-v�9�O؅~�!򤁵����0���r`��i]�1�!�S�	�5�B�{�����"�.�!�d�X��d[� &�"�*�A�4�!�dV:����gO�5~{��C���r�!�d��=��D+6
�d=��.�<*!�$�HcČ(N�����G�4M!�҃�P���	Dӄ��v�:$Y!�$���Pȃ5̾M��yɲ杕k�!�D]����s�1]a{dh F!�Z#MҘ��	�R[>y�A�
�E!�ą2V�E�F�@6���+��02!�D4� �� č'��� �7c�!�4%+�8�Ce��G]�ha.-4�!򄐚:�֍���hS0�AA�5�!�d�11�m`d��R.a#c�K�S�!򤋇B|�@api��W4H��i_��!��َ`NU��,�Q�$D���j4!�T�Wr� *k�)	`^<3�Ǆ')�!���[Щ3�ʖf5������!�=:֡pDh�	]�zI CX��!�Y���;ģ�m���q����~�!�� n�b�b��S(	��
�tK0���"ON!Y"hň"�N��nϛ{8\a@�"Oi
��A�6r��U�Ȍs�=�Q"Ot<`Џ_�O�n�Ж)Ƹ05"OD]����)�P�q�t���"O$q�̌�@�`�"�'8
�>�`�"O���&J�.��yPdD���<��"O��I�3U��,(G�2�xAt"O��9�Hs�0����)�"O��ࡨN{[|5�"��n�}!�"ORCs的��ja��=6L��"O"�c@�j�]x!-I3#ɰh�"O�	r��(��p�,�+`�Z���"O�Y����\��,s�,|�r��"O��`S, CDQ+W!l�x��"OZ5ZgA�D��h��Í)����"O2x �M,�ڌ@'�* ~�"�"ON�"� �0c �CA�>_��=��"O�PC�\wv ĉv!�;�^�9V*Or-��ܹ?�R|�QH<v�F3�'����#!.M�PK��q���	�'wf|���M�J5\-�%N	�neL���'�`�r��fe�Ha�LҸd1d��'͊��	�=KRU!�TY\D�(�'�Ё��ㄥh?��Cu�V�gljQ�'�@��gܖ
>(���YX��a�
�'K�p�F��x����b]�Sd�L�	�'�B�J��G��T�b�Ç�:��
�'���Rj�8)|�K�恅�b��'d]�w$��b'��*bq��'��A�B�1�4���� %��(�'U�]R�B��P���!A�aJ�'�\1����;�2�6��Q��'�`�C���>>�p`�� ҏ1�t��'�:�k`W. �X�!�t�z���'	0p�D��xް�r�/�7S�m��'X�����J�Ld�R��4���3�'�tH`LH�c��4ƂZ@0��0�'���.ҽooF�����)A�h]r�'�>ٱƎ�U
��@�D;�u��';r���e�
�X�JD��{n99�'��Ȣ$�<Xn�{sƇ�u>�)��'�X豕�Ej�`��*M1m.Ē�'آ�{Cf_�G��9���R�JIA�'B>�R�c@:C�����o�3����',�(�2h[�6����B_�'X$12�'���i&,�'p����!�2#Vrt�'� ��#_ΎXi�̃��Y��'Q|�#�#/9��6B��P1��'�6��@	9��xZ`�Z�sO&��'�J��μo?����ą[ML���'�f��$�,]���E#"Ƭ;�'� �XS
1;ʽ7�>6�-��'z�qɃ@9�q(�j ?/8����'���#�ǀ{�!�d�/.o�)P
�'1�D�bZ�ƶhq"�7�*
�'j���#��Q�f�2q�A:�0My	�'��Kt�L/@Ɋ f��
��HX	�'�t�ŁMO�Z�;�k�	'J��	�')\|Ӈ ݕl�t���*�:6|	�'1`���G� 4l���}���	�'3Z�c ��;S4����O?rM�}��'k�l����m�\p	TW�b�'L��3�%2&�WI��!<����� ���&��F{��ٕ#�o)Fa�S"OЩ!��V����J?5n���"O�@��B�K��Ɂ�,ޖm0���"O��Ж#J�}4d����VlK9q'"O��p�:u����%OSRP�`�$"O:L�&��4%޴�J%�.V��B$"OE�����@`� ���r��S"O�P�ڰ&���0'o�4{�"O6E:�NXkh�Ѩ��&G���Z�"O$\`5�5u����K@��R�"OD<����5-�D����$�R"O�laO��s�N0�b�D
A��`""O��5�=>|�<[�T2w:�01"O��c��[����K:M� � �"O�p�PNx0Nlx��[N�2!�S"OD�8"9
�2x:�+D�PAp"O(��NÍ'�9ɕ�K���٫u"O�H��/ϥ�f�JV���S��mP�"O<00�l�&E؆���7/�����"O�@8��Ԓ�i� ��:D�^�9G"O�
�Ň�,��r�GܤBP(,�!���^��\�z�M�� ��u[!�D�HD���Ə]�Hp��̅$N!���3
�j�z@��MZD���ɠN!�[$�>���(Dd�y�h��e/!�Đ&ka�	±ڼTrcƉ]+$!�*����DZ�'Nxx����u�!��D�j�9��V�%�E��h��ob!�dY�qc *�ݐN�[f�74Z!� <Zx���I�=��в&7'@!�K��`y� ��\�r�6E(]�!�N�s�� �fF�Pvؕ����M{!���a�li��BU.Pn��7�ݢo!�0
}ά�EE�+;}�4�Dݑ9]!�V�.���矵*u��qsa��>!�$�;1���Õb��H`�akS��%V$!��31n��Ǒ;<��-h�.!�AKmrH�v�H9�P�N��!�D�, ��������B���¢�3�!�$H�_��p��KC�:.�[ �Y�V�!���)���`T��F~�J�� -j�!��̜0�vtS&��:Y��t�6���4�!��j����J�7F중�*?q!�, A�s#�W�2���ի9b!��%??a�2aø��a��п�!�$��aP1h�5.�$ ��ӫi�!�HUh�1��D�B���c��%A5!���� Ђ��H�
����T��7!�dR���&�Q�p+.t�s*�~�!��l�[�kQ�*v��B��k�!��]�ډQ�C��Z������$�!�	�4�ذ륢��oK�)�͊�ys!�D_�S�ع���K>U;<�4k��8;!���`b��$$���#H�3< !�$�
A�$l�iV� �ک���n-!�g�B�i��Na@a�Z�!�B�
�ht�͆{Z\pC3�ۑ!!�� �Ĭ��E�><\!�Op�!��o�.ML�.O1�R M�!��3��Dq����FG0Y�5vG!���$G�Ic`%^�%4�X�Ν�F!�$Ѿ5�L�&c�;i/�`kף�$>!�dR*-����q�,*l�K��ٟ	!�D�!`�����(�m@�Z�AÙd�!�� 0֣D�h���OVX���a"O���c�b�D�HgiZ8�n�x�"O
�BM�0D�ى�*E88�؄��"OyJ��P2|k�P뒈D/t�z�	�"O^�x�GH�|(���M�O�vd1"O���v��$��#��Ț0�V�`�"O����R4�>�1��ƛ#�V8zG"Oܨ�s+ܨ�4�� HQ}��	�"O
3 O��8I���(�f���""Oz9�w�	g3x��c(�`|\�`#"O"��8-����HhΘxr"O���.��
�3!�n[���s"O�$���0��4��
�:4:�m""O����,H(Pp�P)X�G,��"O��0� �D��)���#d+�=���i�ў"~n��W��bԇnc�����4��C�,KU��H��š#2����딺n����p?��Lqj)�g%� RP�R�gW8�x$��zU߂)����_;\��)�$D�LЅ�̧e
h�� �����i-ʓ�hO�S�.F�@"ڨz�l�K��F�B��t���E�"BD$��H�{��B��8*@]A#3>@^؀���,WB�	�
���X�*��Q X�ّ�A�p��B�IE���Ғ�"f�l�����? �#?Y��	]�.�p��g%�]R� ��)�!�dB�9���R塎� ���r�@'k��A<�<�%�
u�|�9gh˞B���P�c����'��[qD��2I�2��R͆����M���M���<���'N���JI�'a�&�u!�0���~�I�I�L#wFX ľ!(`�$v����e�����B����c�*;y��+�dz��G{��ɝ:kȪPF@X`Ey�Ϛ<���
O�E��O�Z�$lq��҅wK<ŊRT����	�cn�А�,2���Pg���hB��|S������LXaaźQ�RB�	<o4�;�Ձ9��$3�$:Hh؅ȓ9�L��ą�z���q�
PQ"����>h����M4d4�� ��-�E~�S�?nī�)K�Ș���y��B�ɸJ�F��fO6+�d0��.Z[p���'g�?����^W���5LC/J,�!*5D��ۗ��8<*�������P��q�|F{��i�W(�ȄfM4S��e�F�q�~�Y�hPX9:Jm�f��N��0[fbC��y�%P�l�`Q��JՄD� �J��y"��#L�|�4�\)<��y��
��y���?h�컃d�'CPJ�"@0���p>��gH"jJ��2I�7�|�	��O�<�Cf�2�����U�ZY[V��r��0=AKZO��ʦ�R"uրH��΂k�x���Oc���l�(m��D�$��;:�Π�0��HD{��I%H��A�źga����,\�@!�$
�i�`P��0��E^'S�'F�����0�4)ńǻU�F\�6�ь$��	���|<Q�^3�ؙ�k׶uI,�9���;��9F��o��#|zp�2�PQ2
Ŝ �i���`�<� F�>n0L@�O&��Z`�<16D8rb<i0c��b#��R�%]S�<ɔ$ӘU�tI2C��"v���RFLh�<�"+6lxP�'�W 7%^qJ�MKo�<��G [���LK��P$�C�<�F��"�*p����`}:(r�lKy�<��Ùt�-�aA�@��
2�hO?�)� ���+Yf?d��q(��Ra��X`"Op���W wg�}���]�z�6p��':4���e�Mdm�ƭ�8,78����0D��"�I�A�x���X�`��B�2�I�<Y	ǓP3��V������	�Z���z�pb����^�F�9�@|R�3^��#>��i�/����lR ;N� p	��gQ!��������fT�Sȟ�w�	x���'��d�$E��A�圿R�n%X�fM�T���<IOIZ���O���B@��%����⊍.⊅��[�� �W�O�t|)c�8]�)Ex�O0ꓺyBS"|�����Is�]�A$���'ўb>��%M�0 ��$����|�TDP�jE[h<��J"Bx��î@i�d@�K]�<-P1AU!��Ԏ5���Ӈ-�@$�ȓ1����Fiͨ Ӳ(0�̛Q~Մȓ(O$�A���?4�I����	R�ȓHDd�Q
Y" X��8vO�����ȓ#���	4a��+a�H�j�����ē���S�A&�e�#۬���b��-U�B�I�X� m����o�צ��!��'�a}��@�.1֥!�E��),�AB%葂�ybnHLT�m���X_ڸ��oW7�y��
, D]9���.L��9�c�����7}"�>%>�?t(�EO�m0X�A@�T�lq�O|��dV�6SD���<d�Ҝ�b&�'�~�\���寂��]�<@h�.�1�L���d�!I������N��	��l��'�a|"�ED`0����>����ID�hO:����Df>��ɃC�Rܸt˗.I�|h"%3D�PK�ˋ�gq�õd>l|�6,��HF{��IՄ&mRhwk��y���Ŋ;)�!�d�=��L����a眅��%��dω'�ax����J��J
��9q�LEZ�H �c9D�t�$"����#Jx��t�8D��1��P%��6CH?:��5S�D+D�\��U5]��y2��3Fҍ�fN+D�����؜&�̀�O�"+���&E/D�Y�c��f�D�Bs)Z�˦�t�,D��в����R2�W=h`tl+D�|	 �I-����`�{v2x�T�%�O���z�D*`ʞ=`E*'�C��4B��/@&�̙�m՘2Zq�d�>"?y��;�hKE��ژꢄ4D�����	�h��5��gȫ2m�U�K����C�	7��{#N^8{���P��D�z C�Ii��y��6)t�k^�RB���E
Te^m*
�K�B/e"��Ɠ�R�h��؍>�� ��K*J��E{�O^2���@�dd�}� �J��	��'����T�.�(U�G��2.�T��hO?A��åe�lxd��2z2(��N�_�<!�޹\�tI��lG��Х�T�<�d�Y,B���� /� �I�j�<1rM���Y�F��l�9��)�#�!��׈D���ݮ!z��f�^�6[!�d^'E���Ǡ�ks,��$��Y�!�<�\#���/tnN�qC  )����~oU�S�O�*�+��;1o`,qL�"��U��'e�١7����@�A0��8s�n1D��6�V
PJ��H�ꛭ8�╋D�0�D+�IN�'�j�8��8%��)�n(����
��y�X"Ib`!QҊ�hj$�ž�y��[.�����/��$r#��)�0=!�
� �I��Ar�P�G�VHG6%�"���Px�
2�F�q'�k�2<r �ߝ���~2�|R�@Zܓ�*e�b��m�v���mȬy�ȓDE`�0fݛ=r�l��D�X�|0�ȓF2�R�+�S(h�EÙyO"�ȓ��!�T<Bo T��㘠$��ȓH�������'$�I��i��1�ȓMR�P��a�>�Kn\,p}��<������O����s�w�}�5`�� *�ɰ�'�x���M'K�����KZ�A�<Y�AU�06�8S�ظV�a:r�C�~���O	�$@�èg#�`�f
�QF����'K���&ѯ2f����S�N�T�	�'�֐���	:!��3�`��Bhz|H�'��@A�Z.Ę���f�-4٨t"�'0|I+��C�/HtAH�͚Z8���'#�� K��9�Ĩ��nԘ"����'
�Z���6iyC��;&�:���'v��̣�h������M/8P��'-5����R��;�π�7�����'+M��ϋD �`�)��|��	�'�F���'ʝu�<1D��C`�Q8�'-\A ���4M�|X��'ʀrz����''���dm�7c�%��-���!�'rV���
?s�@V��}i����'~�%ʍ��a�r*��e�<}J�'q\9��Q��(�����K�9z
�'aV}�	�;��A������	�'�$�Y��ݸG��@@f��~�Ur�'ê(�wO(���V���}c�� D���*ұX�]�u�X11G%0b�9D��P�aF�x�<�"���b{6\���5D��� F(j��IAq%� D(�"d� D��R�ܶ]�h(
G�b���=D������ʉZ�M	�C.��Pq�%D��	%̖ @Rq�%	Rz�)qV�7D�$�d�k�`���ˈX��M+�A7D����kQO�%)n��0[T�7� D��)�ȗ(�<�I��T-m���`��>D���æ����,UO��t{!
 D�8y��}���*�C��dk�C8D��pfJU5� hуS5N`�SfH!D��ʀ�YVL�B�Q# �Z��`!D�d�R�
&�L0:��P�~A��<D�𐁮�7C>���s���q� �E(D���숬R=
�@䎒�1ٔ�S��;D�\��C�$�tt�goσ,�%�G=D�+��$\V������.,ۀ*:D�l�ц̒~Z�X�$�/Ee��F$b��W%,�O����I�q�ҹ(t J*k���"Ot�s
��r�0ebe��:3TD %"O��" V��9Y���:Q $���"O��#��В4��jKݏy�Xs"O*�+�dQ�,��F��`x��2�"O���UQ)�$��ˀ�Rp�؃a"O�����\%J�b�Slڥh��a�s"O�D��Fa�h)vLQ��P1F"O�()��ǌ �<�r"Ce��#�"O��c��`�b��#lh�T�%"O� hN��8�`�%��qTH�"OVy���²G�EїE�1R�L� "O.��2iD�Q\��Dd\+�|3T"O�ԣV+�)ʎ�JW���v��x�T"Ox�+��Z���`HC@�� ��"O� v�2(	��I�s���-���"F"ODXsu�މi@���ψ�j���У"O�њ� H�g���ȃ`S3EX8&"Oz!��*��)�^�YQ��~tz�"O��{@!ξhn|A J������"O�2��/c�P}�A%G�z�B7"O|�� �S����'d�-<�(+�"Oȍ���8R^QpAC�M��Ș�"O�\i%)�.e"��SD�)`�:E��"O��KƩ־@*V�rd��).�Z�A7"O�dXB�I:�V�ڇ��h���+P"OF�9@oԤH*X"�+ȖZ0�+�"Ot�Qߝ��B��j��hD"O� ɥ�ʝK�	b�Dڵ�\r�"O��I%G��G7�\�$��6>�LT e"Oꀰc���6"8�c�����"O�ɋ��:JT���\%���"OFȢQdP��!�/�,Q��Q"O4ˇd_(s	H���*���p"O�-����+?�(�2�ֺRټ���"O�q���$cJ5؀΀z��"O�����a�Z41@)�OI�`�S"O�ĳ�h��h�E&�C�j��"Ot�K��T;<q���
f��4A�H8e\��I�Fh�!�b��a d��� �S��􄇱5|�L�����C@,Y괏R
4Z��-D��B��P�@����aoՎ;+h���)�	8!@�����R<�v!����`Ɉd��1��]�ȹ���8D�HCtDݎjBh�g�ј=1�97IX�GCqO�뤬�#!�qO�aj�w���kC�ז?BD�c�b����'w*01�ʕ|�j��R+Kb�M:@'B�S�F�؏{"�H�P�Bb?���>j���E�&�:�2�	��az���pp�O�thw��P��#���?_��*��O@��l߰�0>�a��5w�ҀED�]���X�iC�G�j���h�P�x<̓7����DM/fC�ap�o�b�2@�ȓ[���5o�	;�@z�g�"q���DyBI\X�k�S
��{v��>I��B�!~�B��LLLB�gN�D��H�Y�L�6�C�K���"~n��?3tH:T$�p������54�B�I��<q��;S���O�-�DC�I73�ʱ[��X."f��3��˜L�B�@�d���ɔ>��Xk�ZP��C�ɋ^�*�3�D#,�r�k�?�C�ɨ��H	���yt��!�B\�C���9���<N���,KfC�	���1�s�
-��$�l����>��'����I�($��0��g:RDQ�'%:�aFE�7��:��� �0�{RB��T��SU�>\�`���ufܐ1C!^�	�ZB�I46ā�äɠ��۷N_9y�h3� <�I�tQ>�;����%T�?�P����L�_R�5��8�&�[V�r H�%�&�V���<b� y��ɾ@����˞2Q�,쩇�ݾA���$�5p��c�O��!�Ï�4p�����2l�v4Y�"O50�gX|�R���/F>(B�)�&�d_�"ݚL��'\8�MN8U�X�c����ȓ|���E��K�`D��e����G�+�	��H����yZHI���I�T�`��@5b�B�I*k�0B�V6Q�RAB�l�)��B�	�7�� �
�vȱq�M2!3�B䉷6��hŌ؊L��a�"�ț�F�tD�͉x�ax�b�
�4��&��t,!�F����x�"˞h�eM�4.Z���DT�g�^�p2 ?[�����Q�����	*y?�trDD�%��OD�[��%���K|� �d �OA�.vRu1��/bւغ�"O�Xh`�&K$p��-� �"�B�U�$���R�i~��>�|�G�Z�:E�e��!Sn���e�[�p2�SY��R	�$�Z�!��,\�P�r0W����[B��3�ҕ��)�h]�Xw�[Ag�E�zqk�Ok���(|�@a��A�RbR�J
a|��xSX����K�6aa7E�J`XD��lO3/��X!�钔uV��䦄�O���bM,?�����Oޮ4�t
��O�`|!A$Ծ5R��Ě�E�AY�I�t�f�2��+O�i{�wW~�idh��7������¿kG���e'?w	�zݚpy5���}�ŋj�fx
�@�'N�~hB昿4T���*��Ch]�䫆$Wi���@Ŋk�d|�`6��f�	޺9hw���A`ԡ�� 0Apa`�Z s6t��	#UL �3AW�.Z�lK��vED2�-:h��2%M7g�b5X7�d�9��+�^���ə?�����?��V)�L�԰� (�(�(���F��A�� =	�4�@%B��򨠥M�5���I��<_2H���]� HI���7Lv����OL��v���N@괕'f��k5�7+���%��03�X%(�B�۪	Ը���̅jZ�9��S<gj��b `̹���ˆ��X������!cZ@�gJ�n�����'F
	�2��?�0<QCJ&یuA�\�}�ш�B�3��1�ٶ�����ڌ"�Q1��%܂i#!,\�	~��ؼ�V�Q$fٲ�ol�ؘpka�<	E��w�d�����H��L�HB�SS`�Y��|��ď�6K�4��S�v�h��g`�J��|����<qB�/!轐sÜ��	7�A4�0>�tF	9+	�R"�-p�R]ہ���H8d�뀬�-iH�y�OԴ]�̠��?
�>��6`�u�BEG|Ó0p��2�o�h��$pիݯ�(O���"��p��
���3j��(X�K�-,:*%[�E�=JJ�E��	R�T �T6���$�K��}�/	�u�ZYs���T�Ă����zX9�ĩ�*I��n\(mmX����u�:��O� �"�B_�LMX-BP(�	(^\���'�d��$�D��0�d�-(JL$�S*��LLR���0B2���$ģ:�1�$ђ���"�y'#L}��ŀ&�I��$�@Ϛ��y��:�jP8��.R>L�1`F#}O0ѹ��A�|�J�%�p��O�ўlX�e̍K��Ђ�X�D �wE>�O���w�	�.�.��B�4X��9Cj��f�|$+D��1�0%ڝ1������q�t�Ӥ�Ҷ^\8c�ҵZ��X�K$N��bg�
�h��00��e�t��^U���,�&^��Q�>�yb���_
��S�nUcf�m
�L�'j�.��Š��A�@�i��$C��q�v�s���e�M+��܁�"K�]
�b54D�� �	O+�,��/E�0�7��
r��T�r���YFη��L�xDT�3ړ"+���3�R(:��+�m�fJ���DU|���Ɉoh�Jtt�N�X�.�~'rl@V��Gr�LQw�'����l�G�a�`��8�� �M�NcF&O��Ԡc�k&�$�u���+��l7$�
s#�y�m
@�Q#�������J�MbcH�"o���㒼;��Xa��s�b�)�dʨ4��,� @����D"O��9HQ88O�qc&,�6�́9ǯ	[?q�۳`u�!�%n9���	�{NY��.E�_�(DI�� 9��$��@w�- �ߧ �Z%�"IB�
R8E9Ҭ�43��u
�', q�v�W�$�,M�AO0�Ђ���!_0�໌��!Ջ~ 
Dxc�5s>dPPaaѶ�yR�S,A��\�seO+u��drDO�&�y���"%�ٻ�.��OB�PI�!�y2	D��eJ�B��)�9!pDT��y�<aJx]���(f��x� ��<�yrHG:L����E!��C�P�y��U�}cƘ��c��$}�й�	H*�yR���7J��i,���a��h�y*#�Ll������GƘ�yR���K������ӽ�����.[��y�*��, ����6��ͩ��8�yr(��q\j��a�X�{g�`�e@��y�=~(-��	E(��I	� ��yrfWn"����{g�Q �(��yrg��y��c�'}���B!��yrf$%ǰ���&��Y�<���ѯ�y��*��b�T�c>����y�'_�4�#Iȫ.�8Up2��+�y��2\=D	���I�u���l��y��1[�%ʄhK�!Ĕӡ�ݧ�y
� �mɠm,Un����c1d�<X�G"O�}��P.����D�6��U"ON�rL4�����G;�ᱰ�'��3&F̓� I�Q��P5 S�i$|���" D��Dĕ(+�\�gѝT�^���C??��#9�x�xM>E��"���G/��:$�Su�5�yb�7=�F���,�%m;�I��e�����'�rh��if��ϸ'#:��E%��bon��D��<�����i'6��E�H�^��h�7�Q%�%��#P6}�t�uL/�O�t��+�hT"ɰGH�l b���	3�lr���&��Ok<d��&�:�G޻`���$8D��YW�W�l�!C�Z�$g�<A�Ew8R�3}��	�d�*��L�.��)�ㅻhu!��O�\�H�mW�&��VX��OTY"R��.����qO*�vm�:���B �l�#�' "���Mb<���G��.Dㅃ�0T 0�0@F�H؟x+����ȢG�3x�@��  ��`~lR���c�����ڕ�Z�R�`���L�&���;g"OB��s	È��%R�� )��������[䢛�P>%%�"|���@�;���h�&`5���f�Q�<�E��IG�Q9�K��'{�
4��Q�=y�r�(Or(s`�0餽(��= t� C"O�8b�>WʘId�=w>Yj�"OX�BJ�<c���seX�i5"OF�:wU ���W��c�ND�<��`��:l	�Q��xL����E�<a�B:e����!U�;ƕ��KC�<)�K�)g��) ��ۣ9J�ԋ�[y�<�,T�30�m	��[�ؼ��ƪ�w�<y��:R��1(�NK�g�2H�գZo�<�"�	x��!�儭bk�E�g+�|�<9%(�>�HAz��\� o`y���z�<��E�U���Bc j��Z���L�<A@X)TU� ��`��a8��Hu�<�5$�����D?�8�vO��<�d.Q
>v��90?{��@9 Ep�<y'a�(^.�ze�Tծ�
s��l�<�B�Мk֬��(��G?��
�E�A�<)熍8�
xB�M>s��  ��B�<��.��)ha�^�(��(�GC�<I"��D v��'b&�q��P�<!�m�4N�\��r�(D�p�b���v�<����9Q�>ݢTK'<��<8��p�<�2(�,�()��+M!E��,!�JY�<�'��T��'�ŻuD2�{�ŋo�<��	�*�� ��S�C�ʜ��C�<9E
ܽo<4qK��<zQ3� �`�<	�얫C�
%a��.x7�	3�k]e�<!��T�5��4ȴ�/a��
�J�<9��_Q�� �W<�N�z�HX@�<�#�>j��b	��Y� �1av�<A�	�h���%��p��B�Br�<)�dNƸ;�����M�6��W�<� 
�D��-��mV�~�:&��e�<��ǖ�A,�X kȖc��ԙ��^�<�@!�3Q��q#����BYfZ�Lm�<�f@�+�6�s��i4@H��"Qn�<���%UB*�PD�)D⨛���h�<)ʕDzP���N+so�|�R��k�<��@�,W��K&�V>�8��D
`�<��	���D�Ⱦ\p�����`�<�d$X9v�L��9p��ѹcnT_�<!�`��"��=�P'��r,S�Y�<�$)�;W�LX�E[<-��2!��a�<� ��R��ۖh�h�N؏Y�\�"OR	(�@�,>	p}�$QS�����"O�40��W�Y������l���Y�"O�HuC�m5*�#�&�&T��`[d"O��Je��!�t��@W)<T��V"O�2!a�p��3/�<?R,ѵ"O�<� �
e�1���M�Nx�@[%"O�x�I��X�>E���D�H�5� "O��6O�.��-����r��٪�"O��ͬ=��̀Ɓ��Y�%	D"O2hJ4Z�H[rH!A�C�~,�'"O�h�����c	V���"��r����T"ODmY�-��{vaA2J;��"O`�i�H��^�����#�}k�"O���UQ`|y+���@��`�"O, �$�)3L%���[O� \zV"O&d��@�AA�1i�UB� �"O<E�%Ooϸ�(��5� �� "O�����Ξu%&�2�lŹr"O��(��c�0�jD#_z��|�$"O����!(�n�Ҧ��O�Π�t*O������
6j�B�)ג+�zI��'yh��%�$}oRd���:/�`8��'��0��#>Rl!`g��1%bx�b�'@�0�a�-c�
T���ݫ�'g�ܓ�(�%=P<�ʣ��� �dA1�'�� ��H-T���K�-_�~Ď@��'��yA�M�0i �W:m���'�4��h�-����n�F	�'#���U����U+\6��*	�'���(��m)�P����3!�.���'/lx��k@.m喅[��W�EРy	�'�|I�7�̜Ź���<�FmS�'\�(�s(�.��؃!��kx�2�'$|���'X�|��h���qK����'� � Ax��R�$U�o��-��'h|�qp!^�R�&�ScaK,�^���'AډЅC��f�Yf��"����'(����K���p�x'ݣRԢ�B�'G�����=D�Z��h�;A$���'Ⱦ���,.9�h�DcQ�H�����'P��/F*M'�$��ϠD�^@��'�r���&?�	�Eޫ6F>L��'���Q��~�ͳeCͽ5�E��'��N�9膄J�c!����'֜iA*QOI�y��,�(W�P�
�'�������\plY����( ��	 	�'��$j��Ӯ����$�
K�@Lk	�'�h6��	'�d�sB��E9� �"O��\�o�t��#U�1!�A�"ODe���@�c��m���
+��кw"O�P��-��l��H���Q�u��2"O��à��?C-LeP��ƞ�24�D"O,Y�p����T�E#:T�f�w"O�u�F/]P�UmK41T-#�"O֥RE2jv|HPk�;���"O� DǏ�V��#�Qq�"O�]�%"K��0���#t�R�"OTYٵMJt(��F�X�&!�&"O���w�% �C�c�#9��!p"O<p���EI�xHD�8��xa�"Op5A�Þ
�f���`�,u�i�1"Ot��`D�\��ŋ'�9yJh�"O���T�YU��(�*W�6��h�f"O� .���7vDlx���)�bMS�$	�N�"�!�Y@*}�5�]F���ԋB�#_�=���YB"i���f=���F��8��Q�t��\=via�ے���ςH 0zi��8G.J>
<1��	d�S�xBz��Dd�+ "�,B �N�C��C�1*�,��n�f��	
�ɯlA�˓8�Q��h�'��ӧ�O�A��FN4�B\��N��a��<��Ԥ-��HC k$�O�-C�F(9� {��ӓ|RJ�٠$\2EBhԐ�#���4!��%ŘM�NQ�3����LźOJ�i���&N k;��	��V-)޶5�`$�OhA��٦!�L��G�/-����)��e���,}(����0?\�*�Jޤ����'}��)����<A0�ÒBϴA�1-HG%�O�a�HĬ.~�X�@�&=��q�"���H�Ӛgd�,1&)M�*�$���`��"�Y�O
U2�@> 0i$>c�L�B��&^(X1��Q�w����7"ޕ*��@�B�pD�*'ʛ,z)�m��*�zY����&Zt����䯘10C|Lc6��|e�	�i(�O�AX�ː�k�����B��s��c�I�Ə�;�$��8t7�.Y.B���sB�O*��2^ �@��%�k�0�aT�޻��x*�Gp�{m%�`���yl6��q	J0V��6Ǘq�q�g�B����(��lq�'7:]�!�i�X��x���Z�r��W�e��O�����=�"=�Q��j��%L-?�d瓘@�)AE����l�3�$K5H+rc��+�D�5J(v��$@;ex�Y�cI׻N���H���X�
�&g�=�~��tHۋaL<���*�:gz�N�>sp}�t��2�x
7Hَ1QRC�ɽY�|u�`	�	r9vY�C�k�2ţ�	W&�|����(��F��~}� �'fP�yA@M���R<[<~���Ɉw���.G|*�!��,`s#��/ItXD���)��X� NB�5� ��l��(����t&��1@��gz��Ey�ɚm��8�C@ w*�� �f{��v�(���׳G7T�i7�C�2K@B�I~$��+��qMV\	5o� "�����B�^���S�O���{���<�Ȁe(D9}6\E��'�~�����s��0eƕ�C5N�	�{�
V�%� ��	u �� ЇB
;3J��l�ZC�ɹUؠ�S��@��.�J2�_�C��C�"R��i�"j[�/;\�9a(Z��B�ɼ@Yl$(c.�<B>pɡhZ�J ,B�ɧff^e#�fsPq��V2kl����odvU�80����_/n΢��ȓtC�R6��1�.rc�˭F�%��/�T`	4F��8�2ġ�j[�{��T�ȓ���[��6&V�� ��"n�ȓD��⒂J2hb�CV��;�,��ȓVw��+��Z	D�f�V�n L�ȓB�f@�6�Ƙ@"ѪS�F$�ȓ	��	r���0J5�Y��ƈ<ФU�ȓA.P�a
�h�6���A
X��@-�੄��&"tp���Ð�"gX`�ȓk��Q�e#T O�
��a#�1^��Q��Yo\�!"%ĠB�ԜI������ȓ:�8�R�9Q�-ȑY/\�N��ȓ,�� `0�aBL�H�~nv\�ȓ� ��`l� ZY���G�=J��X�ȓ�(�[t�\CL@(�$�Yè�ȓC�1�*�4"Щ؆dE;gT���+����� �ox\����;?3����$Ϡ��'��.n~ő��ڛ�C�	�g?<I�w��[�.���n�* �\B䉧W�R?�UYq h��L��(GVC�	�hg���BG'C(` GN�m�C�ɒNѶ�˵�܈O� �pL�[ tC��B�Xa���)*���C2�B�	�\�RU�v�ُGG��Ұ)�C9lB�ɣh`���2G��F�n� \Z�OK�<Qc�%�j���t�h*RF�K�<Q��5Dd֘�0� U����D�<��I��
q	��Z���L) �t�<�u�W_NMx��i��x�D~�<� ��ƅĔn��Igω�g:���"O�=[��G���
��� �:q"O����CLek�`פmD��5"On����@�3��5T��"O>����R�xځnֿe�j +�"Oԃe̕�<R:|z��ҬO9Z�"O��j��tœ�3H�����'���5`̓O `�A�K�=�~�Y�!	��}�ȓ�t5���/O���Q�I1>
��'�r���1c}ɧ�L@B��;E>\�� 9�E��"Oz(c��#��A�����1���r�DŻ��[��*���ߑk�F�k��Ԉ"iDK
�#D�bD_�o�D�z�C��E��[�B
�C��ɇE�;L���ɆP��m�G��d�8��S�Њp�أ?��	�;��ڰn/�A�i��	Z��I5,�j����J�|}!�D��Ƚ�M��.�Zat�ƇXj�I�l�E-�S�Oi� �ի�W%��HbO��*|����'��c�l#�L�ʤ�*(�|kt	.}���Q\������{�$Y*1��iP�a�7)�@�K�����?��Y(4bܩ�$8s��������b
��aǟ)K���D�*#_�pBnD�;f�:w��.g�џx�w�8F�8����m�Q�N����I�j�d�p�̝�y�E��.aڐ�o�.nKTM�1��3��D__ٜ��C,��Lㆥ��k*J�b��#:�XC�I�Ql�Y��pI$�e/�`�qO����F�0�0<���.d�:Xz��A�k�*�K&S�<�ɘB��鰃�H�vIt��I�<ٴd��2���ԕz9���(�E�<y�+�#������ ��%���F�<4lL�mg �c��K!i�6����A�<�(T3B@�CK�6W�	���P�<q�
�XQ��R.�$z��^{�<��c2RNXe�T.�#�����w�<���u&(Zd�H�u��	y$HF�<���0vP�X'-�P|���MG�<���Fw�,��GiB�|�&\���<qFω�#�5 �Żb�f��ȋ�<Y�n��-������,8��a�z�<��BZG��`��O��:�ӧ%�r�<�%����t�b�UH�XT�0hl�<�F��@-ȱ)CF�BhЌh�A�k�<�P� �t��2H*zo����h�}�<���?���H���%��
�<�di?cj� I�#uR^}�֪�z�<�$l��0`��jp�w��HY�Ev�<A��ܚ���be�¿���2` f�<ie"��|z�0[�́M��$��ěd�<�pR�����"R
}xD!��g�<��B�ݙ���_��)i���K�<iT,�i�&h�f�$9K�t� NF�<��nt�X,!�k�B�(lsG �K�<�p��bln��W��=���	�K�<����:]Hy˕P;F���ȃL�<��C9j��A�4��u�Π��&�K�<q�OF�Q��@/u� آ�A�<q�l[�+A�h@�.��YҠ��U�<�u��*K3~���E&m��!E�[]H�����_���{�e�.�2bh��
��h���&D� ��`�GVxh��ǀi���k��$S~���?%?ɉ�/^�rx蘛�c@.ð;��#}"ɇ \�O�d��$��8b� cq�%I�\�s��O�]S'8�)ڧ$���S e�T�%*<��H�I�5��O�?�����_98S�&��/���A��?�����>�`ɟ�Sg�O�`񣂦F�"gR��Ǐ5.���/V��򄗟?W��π � wF�e��h1t���`kXP_��z*OP@��@�O��a*B�SiՄA�2�U�V���"E�WPj�S����CR�	�Mҩȥ�T>v*�]u��<A�זS���<��'o�,)������
$`�E>O�͚"Y?�0Q�"~��j����i�h�閅��	�O�4-3��O&l�����<�'i����5�^%��л�!F?* "-��\��Yb]�T	Ia>7�>�' ���Tn�*B��c���?f@���I�N��I�>/�5�����$u,�5L���c�v�XYS��<Ѷ�ϱ����|����lԱfI�i��.3y1�	CW�Ch��͓?�P4�'l�y���OY����8�:�P�� 0V��������d^y
ç%�8i�@�T2���Ҕ���x��0�'h��x��4E��'��!j⪏9;~�]�u�+�`$0�'�剕!Q�b>q��@�f�J�1B��}%� ��,?1s�(�S�O��qqi.����@Ɠ�r�����dUDx��I��#/�`)�d,K�� ��8%���O�'t�q���ԟ�t��,oXÂ�a�fгw��/3V�������,Y�6���z���u�O�r�)%W(X|@H!�ϗ�nx��ɭO@��bJ�~�q�s��"}��� +h
(,��}�R��Bɉr�<Y0��,:�ֵX$�V)s|H3�CCd�<)��d="͑�i�pRH�;6�G[�<���?=�\H!�`B7()�e��QW�<Qb��QN�ӂ!�Ύ)��	�U�<9�� ođ��M!E���HN�<�� Y�!	B�Z�i\I6$A�$F�<�#$�N�ʤA���9���x2 @�<AQ�F�EC.��c�Ųw�fX2iCs�<1�
�,����%D�ؓ���c�<9��"aR�ȩ�h�+�\��V�b�<��O��w5�6��R�^T��bTZ�<��G�$@Fy�f�:Ӥhq�AT�<�-Q�q��Y�g@/@�ئ�v�<�7m���O�Ez�ʢ��q�<�t�@��8�/�  ݾ���C�<9�H�&.�V�T3���RHNW�<Y4��>�hC�З.v���g�k�<�V'Wnz銲@ݐ9�^����@k�<)q����,�p��,-\��0�o�<q䪙� �R��2i]�{�ޱ�E�C�I��qP���Y7�	Y �^Q��B�IJ�R,A�Ԁ~B����,/PC�1M�,�jc�U�OD�e@�d/l�LC�ɶ0(�� `�8,֘B��!]*:C�	;oZ����¡y>�db�m�74C�e6�Y	��tR��!#m�I0C��Ql��ִk��)�N��� C䉽sD���˝E���
�%�5�C��!*�L��Xo.�E�$;�Љ��'� m1�
�>E�Px�eȑa�xŪ�'��d�2-O�C���B���	
�>�Q�'L����˨|VN��L�	�Jd�	�'�=Kj�o�X4�C�	���e�	�'G�� #�>Ci�#fEM_8�Z�'¼�����D�A��Ǐ�0��'7h}���9�]�U�X�w�yI�'�D��-�H��e�U�><vl��'B�ᧉL�cQH�ceL�$� K	�'+X�Ul 'Y��_)t���!
�'�v4�����`��0А��	�'��嫷c�D"��d�]�
i	�'����EB`Y���"���'�lTirHns<Z3DL �hE��'��4���;ҕ����f$رY�'
��Ua���+�fZ�X�zA�'��-Q5�g������]�^1���� �	Srl�u�n{���d�!0�"Ol *��ӯoL�{qM���&�	�"O�Pb���ٹGm�01�j��V"O��f�QW�up�����l�@�"O^=��%!$X�� �M��؁�P"O�E@��7r��PI��,8�N���"O�1`�kZ�X�d�CV�&G����"On��ˏ8�2��dèy[��@�"O�M`��Q�paTC�CRXc�"Ob�P��ҌO��aEC=|ybQ"O�`��u���x"cˬnoN囗"O�<�����
Gz��-��@*
�'���0��U6J<�FRܥ��'���pABC�? �L�[�x��'½K�B�)6�8�2���"����'[P��e۽H�z�z'+�/?��9�'�X�GK�xZ���Cn��	��q:�'�L��.��"(���Ʌ$|9�'��L@�mI�Y�ʨ��@�0�T��'�kU��E�.�r��v<Y�'����A�4|�dy��C$HR�'����	*��X�^5.~ZI�'�Xx��PvN��Bq�qz�b�'�J��dJ�c�nm�gf��;�(�
�'ަ� 5�U�#V �6�Y'-��\�
�'F6q�Dݦ1�J5��a�{h�
�'b6�J'<M�@��"D3oҤ���'�x�C��LI�GW)9҉��'�F���ͫTͺA	�ɟ'"$&l��'2Pz&$��JR����N�XT��'����AU�@�j�����EԐ��'�T�ҁ��EFL��&ϊ/�"O�i � ��gl�q�A� �G����"O�ab&n�Rr��ۃ.�DR����"O�}Y�ݵk,B-_OT�	!"O�� m�-]G�	��L<Q���r"O���&H�&fV̸�-�,iVm��"OFP��lN���2�6(�L�`C"O:�c�A��C�f��1���=�#"O�Q�D��>%�V�霛X��%��"O� �d]*IĠ�@��_�: "O�D�v@Oz׼��h
�?��͸�"O�mA)��#+���2��y
�"O�qh�"�I�M�ࡕ�~�vl`�"Ov�0�Ί�L#�Ḱ���Z�d ��"O�݀Ƥ��ABp9''�"��sS"O��Y�U�y����F�9
�h���"O����=/�� �g��,M���1"OB��vMT�m�b����6^��؛2"O��S̳�J͑S/�a�Z���"OHx�ʊX'9��KEJ
� ��"O�u�@D%x�����*�5
�-ڣ"Ov�96G2�@�2D���|L�"O�y�1ǅx
]�w͉�3�4�a�"O(��"Ç� }R nł�
�C"O�X���+�X B̅/PQР"O��5��9li:u�e�\�	��S�"OTٹ�N�((OFL:F%�/����p"O�P�@;R�19���/֎!�"O*�XXz��6c��i&C2!�DH�Jwx��AC�i!$@�/!��03T$�t�H�(%�#Eޢ]!��}vfQ��!ЊS�2���D,{�!�$�'ʶ-֏� ,����'%�W=!�� .�y��� v|�,єCRD���"O�tx� T���s��C\�Z�"O�����~)�-!�#�YZri��"O�-�ӥ M�¼� �5
f�y�"Oҙ;#/Y�A�A0��T^\J�"Ol��gXY�QƝ%v=4���"Ov4x�/\�vi���М~��W"O�]��iӅO�f�h�*��e�Z"O��@�fޤGC�$3BI\�e�\�"d"O���G�<�6�⥪T�5�%�""O��Q+���,���)ʄ�
�"O�QZ5C��O��R"c�v�"O�=
4�3B��@ -1��X�"O�=#@���3.V�� �3 �e�&"O���%�Õr^@ ŏ	!l��E"Ob1bS��"�����΅Z���yr"O ���D����͓�y��T"O�}��V��
<�DK���"O0	��J�~X���g]��)s�"O���IJ�X�B	���L��,��"O�0���ͦ$ɸ���I��H2b"O�# ���+�dq� �y~��3a"O�:�K]T(�c�{�8Х"O4t¥�ϗ+�zx�lmv4�"O�!�����D�EY��A lU�A��"OV����/ T�rU��<�]�6"O���Gd׼W%��H�h
9�e�b"O��q֊�-�`����#d8�q26"OX����ԥJ�"��'D�(y�"O�봄E%��0v�̙*Zt��	�'x�ᡦ�1b��.Ҹr�l+�'ڦ�pЌ�W��j�KD�qF<�x�'�&�Zd�J�R�,�����n�D���'C�E����;������s�0�'�Ɣ�
S/�(�$G�eV|1��'sL\���FT���Gf���
�'�Y�wNX�7KLpP�I�0q����'����#�8E���6B��*�!c�'�x]��ၨS_&�1�n�X���'y08��R����նeѾ���'YFDhኆ.T��#�ݣ_�ٙ�'��q�WŞ�#2��!���6\´�B�'+�QA�Ǟ&N�5Z!i�M�J���'>X��LUN�D`*��>J_v��'�����%�a\	;!��=Q൱�'�hP��H�:�����@��(��0�'̑�ǥ�Y�ŁE!��Mpr���'Xz�S�B�.p���b�/֝��'��HBc.�.��e��S���y�'�F��r��&���;�FBH��A�'$6���G'�����ʅ�r�~���'h��[�"IȸB�c�t�:�'����'ʙ�P�Nh1¶Y��)9�'�*��c+��������%�y��T�\\�Y�C`�����;�#���y"ܚC� �r�U"f�(k79�y�Ozaejs-\�I�)�(Պ�y�`��P�R���pS���y©Z�qy����s��Mʦ+���y��= ��8�,W�l��p��Z�yR*Z�/�$�f��..�Y����y���)�<P-��*�i�&w��C��.���I4�ߘi>���m��^�C�	�Q��\��,_;]��)�g�M�K��C�)� 2A�G̦HHp'f[�(�"O�qC!J�=
.�A�,Г`W���v"O��.`�z1IR�D"���Y�"Or�h�cWH�ꎛt�1�"O�a���B'@K�ISDhW��zi�t"O�c�`��9�SfZ=o� R�"O"`Q�T9���Qt��=�k""O�`#DeP����R���u�(K�"O��Y	��W @up1�=,p9�"O^ɂ�I\�Y>ҹP���W�}��"O|���cZ����Qp�U 0C8��"Ol�	5f�%fO�xR���hY`��"O�\�.R�;,��ؒE-�ypv"Oā聧^�b�9�2�R�8��"O"���.�y޺ #��vjj��"O��.1S �@*���.C}s2"OR�%�
	n�zV�gT�i�"OBD�a&�/���Z6dEy\���"O�Q�`��{��AӰÌ"nq�e��"O��p�Mի>z��B��PbH!�q"O\h�Ю|��5�F�� �q"O����XPD��M�K2tK@"O��P   �P   �
  '  �  ?!  .)  &2  i8  �>  E  CK  �Q  �W  ^  ad  �j  �p  (w  m}  ބ   `� u�	����Zv)C�'ll\�0"Ez+�D��8��M�P��<iW+	ٟH�hǺ��o� -���
6��x���;d�N�M��P�H�V��	Aa��]>b������Ӑ2J�mJ�A�Qd�jC�I����F `�}y! <vhX[�Z4Q�x��_wX�R��OvR�ľs��+�� g[���֦ԶA,��aL
��䁷�$��3-N�8�lZ�~1H��ǟL�	���ɒ��I�5G��]�6A�-�]=���I�H�ݴ-?Hؒ)O:�D�[�����O��dӗ�>H`u��5&�(j���5x����O����OF��?сbք�Mkt�'���H�����Ձ!�BI�� �I�HF|2�i�D5�b��*Eܩ���y���0aç>i��Ĥ��CBKB$e��S�3\��a<%S����~�l�D�O���ON���O����O�˧�y���^�<�� X�5�앰���?i�i^46mO�ٚش�?᣿i�PFw�@-#f��O��'�_�);�Yb��I�|FU#G�M�'�j蛎��n�÷�s�j�17� /�M`�,X�|[�q9�H؉s\�0�BFz�
<o� �M��'��blT����Q�C�(���Ū�2<��93"��h�����*t
�hQ��g.��r�#N3H�J''��e��6͚�A�۴~�p4p5d�R�4�$�K��j���'Z�P�!rC���y�to��BZV�	/N[����, ��d��)}�%�g/�a*H�z3]�	��`_*?�B�	�4l��(b���ء/a �P��
芸{^w�!%i
�������dD+��i�^x����y֧�h�L���'�Oxň��߱-@�s��080�s�o�O�����ǟ� ah�0�McʟzAŦ��F~Q���T�1> �2�'}�	������|�	ߙi��Ժ�O���͖�b��fn�tW��kf�)@����D�.K�=���/a&��4��O"�yv�ϧ���BR�T=
��H!�'x:����?	�T�@�<4j ��[�E,L��g�OH���O��b>�ϓi�5�To�$>X��#�K�f�����Mk6%�&��y��ȑK)��*> U���ė*C����B;��+gJY4H$b�*�C�'�F@�ȓ-��"�)��?�zPj`g�m����(ܬ�Ru�Ũ֤�@�ݔ:5
l��v� ���c	Mϐ�auO�A�����b� ,���^���:S��B:�ȓ'$���ș� B&Pr[7�p�I6qb"<E�d�&���,G#Q�Yɒ�^�!�D�3JJ��h�c�$-x��^��!�d�kV`�٩w&�P���$.7!���6�ʭ��%N.%~p�@�Ջ!�0HZY9�.C��ZD��(q���6u!�Ȁ&F�'d�Lp�c���#3��c�<9���?q.O��'��$�z��б�0!kX�x`�� ,��w� �K��}�y�xI� IU�`h�C�ޡ>�T��%��7���
w@\� �8��0k�n�ўD��cH<Q�j ��*c�Y��A�X���æ�+��ľ<��O�@u��oyr�*Q-��|�0щ��'�!�dҦp�dL�敉x�B@j���T�BFg���	ͦ��4��I�74���lZܟ(ϓH�xC��:��t�B�N���cy�'Tb>�f�RV�+1����C��)�G�ԁB����}�iE
G�"~ax���'T�0m�C��fV�I��P�ra����N��8{�%9@��KG`�à����UFyB�X%�?Ig�iՒ6-�O8��g
�0����]�bM&i��E�<������(�@b�ė�e0�L"!v�AD�	p�'?~6�-g��qF�i&��$��� �8�n�c��}3�s�D@���
`��% �����^t`�`b[
�yR� 4or���X9X�^q#ӎ�0�yRB����R���d��ɫ1h���y�%��?�� `��F�&<���.�y�͉�q�����8�bP:��yR� �o�M��G<���JQ)pݛ��| ��%��$�'w��'��7)��5�`�M\0��C��SΒ�.�k�ĵ���O�ej`��2o��'�O*t!�#� h=|x�N�6S��*�F
6\򙉥E��w�64SU��?V1�v�Z&g�f}�G6]��q ���va�3���?A�T��˅��O�b>���O��Dι,vr5��gρWn�JcH�Ӏ��d@�q������Utl����	�!z�'�h7���U'��S�?��'t^��`f��FE���mޗ>'���j4
g�7M�O����Ox˓��'VHH�	��N�g�F�r�B3 ��<�8rEEE*mk�=+�E�Y�����Y ��%�P�ƷVR�{���4e�t( �S*(Ъ�"&�	=E���{e���HO҄�'�ȏZ�[b�B�K!�E�6-��'Z��p� ��?���?����?�ΟP��c�5jq�.�t�x`P�"Or��M�=�hY9�K]c�`���|�`Ӹ���<F�!�f�'�S�y'��* 4�37M�D���'�؝��'��:��i��'>1O� ,�@�1L�N<C��Y���ZW�'�R�s��d��p�Š�.�97��zhax��-�?!W�|�%J ���z.�*NL8���y�DB:'��7��8�޵���Xj�R��OD����:W�8�
��ո��დ|�-Q94���?1-�Ȭ�ć�O@�x�ˇ�1�X��Ȅ'8}�$d�O���B!�X�@G�t&���O(ʧ��ɋ1~(�URÇ
"����d���mW�!*2��X-%鉣~j2�xG%:��~zL�AG�:����49�O0\t�'[��k�H�1§RN@[7A�.�$��[Z�}'� ��A����'��yQd�;.D}�"nS0&����զyjٴ��Œh�eM�zf䄂�˅�N�F�iP��'�e�<(�� ��'��'K"=�xx���&��X�%���1�Q���	�U?��I�~XS�[��Dѩj�b�A�U=^yL���&U�u����(:�;��֊W��6�*?iR�����S�'UH-�2�Ŭ �E	e��Ij\�CS�p���+�OT�@��pbA32!S�D��`s_�tp�O���6���ğ�O��4J���c�ԕ��P.�t��#�0#;:6��O����ORʓ��~>)Y�"�6&��a#`eH �T�ؚid(�b�i+8��Af*LO�H7ꕻz��l��KLJ���I��d�R��u�,*�8=��Ï�i���e��(O�%���Gs���nƃL����it҉z�X�lZğ`�'����"hoN�T�?�(�P)��TD{J?!PE*�y+J5&^C�2��4�WGC��n�Jy�O�7��������3�+��]�Zp�`ZƠ]�4����uyR�'�2:��
�"��~�	(	1�r��}���&		$��	(���4�ax�ݽ'&��Y�h:Zq��g�I'S1���.�����gW�7��q�eB�w8�]Ey�cߕ�?�ķi-�7��O�5�u�˗g���a��:]"�(禰<�����(��� D���~�l�Ӕ`M�L\�E(T�I`�'~�7��!
�n[��ֽ!������&W��n�Ny�ҴKM4q�t�'��OI67�m��١�����\p)ݬ`����ӊ0?��_c����Q��b'$'���Ǭ�x8v�@����:�	5�S�OP�ib��?
���Z�)��KY~�M,�?!d�|���	�������`�J��Ä]�)!�چ=���)΍2Ȱt�`2�џD��	
�Qԉi@c�o��8�cԠKq�6#�D�!6���?�'/:dqEN5Q������$�=�y���0=�Fl�>?o� �� �M��F��C�2"���	�U�R��6.24_�sR�ÄVv�-$��SR!�O�c>c����B�<��� @�_>�$�v<D�ܢ�-P>cDɄ�<O��p7ʽ<���)�'��勔��#�v�)�$'�L�W�V��?q��?I����d�|B�O�	�q�0��Y�,TQ�ti�a� �r�z���I?.��4Ju$�/+GT��EͶ=u<�K�'�c3��A"�s,�zҮ�A�`�%��4z�c�N
(o�E2���?���xr�'��|R:�|trУǧv�);�CJ�!$�2"O½�a+�-~p5�$�� �(���|B�q��m�Vy҈��@@��'����=@V�ƪQ���!%.aRP�\�	ğ ̧An^����>	��
��tj�	>l�BeG��/�݈Óq
��B��1�ȡY���?1�fᑂ�6,1��X%��Å��0<a�a�ğX����M���z�8�D���[�j�ґ��x c+O~�D%�)�'L6�p�2�N�PS,�55���'�ўb>I��4 ��0(T��2����A\�P�Bq�i��	  Ū�b�4�?1,O�ʧ�?9D
���e���2��1�Ũ��?1�Ap�P	\e���ٟ�:3.�!�tE��jǭ^��	�RE����i��7��":(�	aWf�u�O���j@��W^,d�@��M��P��O�\�v�'tp7	�-��o�O�^� @@�!a^�SA䇫S�l�M>1���?���ԟ:�f� 'W��;� GB�H����I��M���i�'�^bc�t�J yw�SQ���`��'�>�� �4�Q���`j�RdB��ek�2~�25�Fi2D�4�p#Ţ��J�E*
$J/D����	U�w�.`B���O	� 궈2D��j�Gߧr=�hk)�A�j%�d`&D�TzU�ĘF��r1;#
1d'D�lbe� }��Ƃ\�p�x�'�<�w��t8���1&��w�Pu���2j%
�%D�� $A���U�%�C�A�5sN�jb"Oh%��_�&��H�� �ZB�s�"O�����W8�����
)\@N,�Q"O����C�7 ]�%���հ���'*NK�'9r�[&o�����Ĳ.���'K���#�Qϊ��P�ͪ+�N
�'�N�1�����2�K�'�<lN���'�FDjT�Êb� H��c\�H\E��'���Dʕ��l�'b��Q���	�'̢��^�:�����~�$#��dG�}LQ?��E(͌j,��06G�1�y��:D�`@ ��Bd,�]�Sצ�� 5D�<� *Ѝ=G$䲢��(�Dq �>D�8��C�"ѣ!�hA��3�"D����i��X�mRP#�b�"D����R�a�(D+Ԥ�������O�x���)�'J�8(y��k5�� r���0�����'�J���!O�3��@,�6(���'pj��숇2Hh婳��v�h��'0.�f^:?:`���n�zSv1��'�%;ǅ�a�b��a�y��]��'�YADj�`�)a��p�t��)O�}���'���ȴ�\| ��0�N��9S��J�'�v�3a�ղJ�p���>-�hqp�'�p)�&��2]��Cg�*�̃�'?��@ƋV�2��V�D9�ĵ��'=rQ;vo�\��V�J�7,b���HӜP�LAzY��A�(�Ƶ�lM#*<��jF �AV���K'
nh�ȓ"��9��bx@=Aa耟/����e�j����Ȅ+��x ��RB؅ȓ^�x!�4F��T8��pV��:ͅ��������9�e��s��YE{�j�Ǩ�<�S�
+"�rܒ�4��:�"O`�Z�ߕx�A�Ώ�^S̠�0"O�\Q�k��)zq#d�L�r��f"O^`�qF%jF$Jg͖�c����"OJA�Fk(n$<"����)�"O"噃	g�!p�U�B�v�'�n�����
;����@v�htQ�;I7$��ȓ)�= ���J<la����ą�8kB�Bĉ
\�V8�uO�;|՘@�ȓNؤ�#�M�wK䘺��6
�y�ȓJ��dZ5A��R�#�Sx�|$�8D�$�H���жD�%���i�ƣ<���m8��3�M1n6�B���x
qU�<D��P��C-��t�̡qD�\�p�&D�@&��^y�ajabJ;D�zr�7D�Z�3E���p�ڥw�>�(�)D�PSC��gg,��j�kb�Y��#�O�T�w�OL�K�F�HFl6��
��]��"O��ANEuWll��Ǘ�&�����"O���`����X�F�!RH�B"O�)�p �(?��S����ҩ��"O�a:q䏖;T=�	�5P<耰"OZⱋ� ,��Q�/mE�q��I8ix��~:۫:���VK��]�̝��Q_�<I��t��ʰ��F�Jܑ��\�<�CDɏ,]�d��,�a���B�<�Cc�:3���s&�.
���ONG�<�$
�"-@�n�]�^!� h�<QDg�4v���u� �g�$�F�K����0?�S�O�Uh�/�:�>٣FJ� ]�d�s"O�9b�_:?m~y�W�F�A��u��"O� j����=�� �������a �"O>�â��c	"��[8g�Fѐ7"OʑhwH  =AJ�MW�E�\�"O��� �1����6���W�j�`�Q���q�$�OrH�Bk�0��;�ұkn^�K "O�$*���.aĈ��.c("Ov��%FM�*)1�X�YS~��`"ON-�q�VKZnU��Y�&C��js"O�U ѹ;���xD��eF|�e�'����'T�0�RhB�(a'	�4 >����'�qr �P�4Qj9��.JR���'w�����@6�:H�6K*4��ʓb�P0��9d���"�I� 9�ȓo� 5: Ȁ��v���<(X1�ȓ�t�+1ǝC�8�sD��n�D{�M������h{���gl񈓬S�cU�1`�"O>������K�T�MϣI�&]�"O�ų�̣L�bD���+$-"���"OJ%`#-��u֠3e˔:Mv�җ"O����왏C	<E��M,[%^t��"O,("�C���0A�W�4�:Y ��'��aË���MHxx&�-���I���r�$@��p�z����^������(�<e�x�ȓ(9�b��y��Q�4���&����ȓr�T0KWꊖ[�]{Q	�qUȥ��I ��g��(�$�(�	X�dB����y����t��(>���������'�\����S��ޡ[ ��Bs!���]��s�\Y7+N~�"TΗ�0��ȓ�v�I�+A��*D�R��?_��8�ȓpy�1e��R��WM�:[@
q�ȓ69��;Ce5���'%��m��P��I
9
�	�M$2�����#�R\�Ê��B�ɧO+��V�ڣ��!3BBa��C��;\{l-۶
�#� }r�R�B�	n���C��k���ʲ욐9)B��	*KP��F�Z<Ja�a�hm�C��#h�4�0�d�b
�hk墖�a4��=��T�O5|�VΛ�Qڹ����[�2D"�' ����
�j ]�	M�|u��'��,;�NR%{�@��@I�{�n��'�ƠR����e>.�1�LUH��H��'����W07H��j4oӾ�65Z�'�Cw�m,,�FE�lAF$���H�Fx��	]�(��}xe(n"�5���Z�@�FC�ii	Ћ�<9�B�,g��"O
�2�cO�ָ*�$Hs��!S&"Oȡ(G�5\X�2$� H���P"Onk�M�7��9 ��.SߺZ$"O`|�DKM��-�� �0>t��cT�  @#)�O
��f+E&�:$�����3G4A+s"O�Q颯D�I(��%�?>V�"O4e@�ҧV$�� ,�(? �P��"O*�9M�4d�i4�w{��!9f"O� �a_�ؽBe��RQ�E�P�'��	�'�e�S��<���##(�3+�i��'5F� ���<K�=+B�5]���B�'��[��*&��)s���N��3�'JRh�s��}�F`��$�x0�t3�'HҜQ�"IT��b��:w%̹c�',�,aF��~�ԀQ�cF�z��찋�$�4I�Q?��e�?���i�쇁l{��Qp�,D�P���W�?����d%X��	%D��JQj�U�MY& �.w2�` *"D�� r@ �� Iwp�5$ͶT]�T�#"O*�
�@R#�	e��>oBh]S�"O������k�X���J���B�'&d�K���S�Uu��Cf̀�3R�<� 	#tx���'���Ƙzc�M*��P���ȓF_���@��fV�񡏜�z2 1�ȓ_��1��#_7��5�Qy��(�ȓ0����$�Q-0Qd!)�#	�5��&'��p%B5T�9@�Ҍhtf��'*��2�`�C�g�T�5����|w@�ȓk��]Ѝ�.n@���[�M��ǀei�iQ�v.����E\N���~���nXGhp�i�C�i�A��b��������"����Q�&�e���4Y�z�I|�T��P(N�L��gG×3�C�ɿt�Ђ�T,?{b�Q4B�];�C��	W��@bB��J��a+Go�0}|B��b�iB���q���&�5�C����8�������k%E�C�ɒ	�-C'�x�! �L��Rkx�=FK�}�O���J�H�*����ۅ
���c	�'���8���c�:�� .���F��'\�hC����~H)�`IWH@X�'j�HQ1M��5����F!�=O�L�1�'�vXDlo�a�f$��HS�Q��'H>iS�W6o�� ��ڕ LdK��j!��Dx��Ie�) �+��0D]b&)���*B�K���t�ˇSo�th�����ȓO��yȚ2P�fx�!�d/`��ȓ3�f���HD��p8A)B�p6|Y�ȓyy��K�I@,i��]�1K�9
�=�Ɠqp̌X�-�\�D��B��r�lx�����ɜ��$D�쒯O������ͳw�hxq;#J9=�*��B��O
�H���O����Ox��4�͕#9��:e�F"�zT���Z��uX��Lā ��i��$�"�I ��O"��ed�(��a�[�4.�h����C2�;�&���^�l��yGN�'O�����?y�����18�J� ��	��E�&����D$�ON@RL����"0 ��c͘,�ǝ|"�i>ɘ-O0�[�h�C�>]�֯�"!����X�<Ч�>�M���?�.�z���O��d�5^'���k������UA�#/d ���[�d����MS���A��-iF��'��O	�5�&�Px�8��k�'��؛'"N�Hv!��߆d���h�E�D��;AU��
k ���a8�y"e��X�IY~J~��OZ���#!�@��ϑ8�zm1"ON%����hY�=�GAS J�
�R7�D�O8aEz�OL0��g�_�u���r��V�LE�5�'���'.�b�G�9\b�'r�'�Nם���&(#~|��Pp��S߶0ړiȐX���tT$��g\�\D�g�'����0*��Ab栲�D��Ut(IHS̷>���ۯL��@�B���O%� ��� �/�d,z@h_1H���^2:���O�=I�'y��Bĥַ4�{4�H>R��'��݂��#)���S$��M�Q��7P����ԟД'�\��I��
v��	q��8@�	�(ˇ4K��I�'o���'�2nz�!�����ͧp:(�ũ��i������
�D�aŢ�
l@�Q�5)C�(�a{�腬^���pe�[/�.��ץť-L8�
рN�9@���a�>lO�IG�'&���NY>�Q"o߷Y�̨S��'�ўdG|���?XTH�c��ķFL%@0�N��yҧ�r�L��K�r(x!:7.�/��IѦ��	j��׆ܥ�vT`�큮�Tmb��<y��Ka"OtՋ0m�gH ��a��d�}g"O����^�9�i(��>jx06"O�e9�镑q�Z��I�_����"O¡����_�y� 
�;O�D�R"O��ꠄ�?�65 ���YMԌ2 �DV%.���Ok���`��_��І�D�ƞ�:�'�#v�A<8W��K�����'m�@����?+��UN�A^\){��� ��*�aO�i���ŊQe�(�"O<���_��t�q�<4,$�"O�A2.�!��-Z	T�؝�"���O��}��C���a"��mߢ�Qܸ6����ȓK�v{�
�
�\�(�n�3a��m�ȓ;���#�^'UH�)�E�U�*�����رT��ےv�%�<����$D�\qT�;l\4p���$�w�&D��5'�j�l��S+�29|ҵ��O4ZQ�'���� i� �=��&�:��'ɸL"@KͥI��!���X���'�2Urŭ[9�480"G��M���!�'v��Xq@��U��,A��7�@�'&�sD��"������2l�qk���H=1P�l�F��#P6@9XCM>�&58��pG���'���'Q�c��g|>ЃD��"q
	��?�O�Z���iu:��e׻<�`����y�@%���l�np{G�D+���kgM9K]xP��%ە���ʧ���-m,���d��x�"�'���'j��M Z*2���O�;]��uK���U\"�'��O?����\�w��܂�+�)}�}�!�Q���hOHl��M�2mB8m��\sPj��|�!��:���O(tb��O|���|�����D��J�`� 2�Ƹx���¬�f;n��D$�/[�X򢊇1k$�#W��.F�V��?���u�	F̧��<�n]}��|;�D�@��ɢ�i�ٛ/��֝7�b�'��D�'��ăG�Щ�v`��`�Iӳ�F�E�8]I��eӠ�$J=h����v��H�?7��4|��5��ܘa蒌7��Bs�[fZ��pn�O$��C�;R��ߺ����?y�'�?a�'�A��B	:�Ѻ��V�YH�d��Q��?)�CMd����y�fB������bV?9z��������&dlTKc��O�P(�'�bƆ��~���?q���*��7u�#���;H�xp�t-��|(d4â�'�ι{���?A�B�?)�'�jp��M�;�N��Ql���rS�9ɾI���׈�&:O:H"��'	�`����O��D��C�.HV,Ҽ-�^��6��yI��`T�r�����Of��κ���y2�۠���4K��#m�ˠ��mU ���Ղ;#ӛ�?O��Dr�ul�k.�����:�V���E�/� 5�l�
E��<��i�<���5O�UY��'5��O\">OLEq26�8U&�!�Lp�ƚ�.�0E�Fj~ӨЊP��O�ʓ�?)�S�g}bE�#7d`�b��[O*���-�yr����t�2Ƌ 6U��x��A�M����?9���?���?���?����?a�#T16Ɍ)��B��Z´�҆��R����'�2Z���IS���$"(D5~����G�!8�UQRe����'Q�''Q���IB��E��ºbf�A
`a4D���+�f���roӕ[h�����3D�� �⍸`/��:��D�B-~<��<D��	�@R\ZqSD�n�d,�'�/D���A�'`�إ'P�X ��M"D� a#�\��YK�bM
`r�D� D�l� �](��I�#B�N��� D����I�iI"�豅��l|a�'m>D��G�;3pD�:%H�/��	4 =D��A\U8L!s��۟dZ������6�y��J�&�˓L�![��@���¯�yb�C�\�b��A�3^���EB���'��M�����`)�%&��[�Z�:ïݑQ�18�Ԃiڐ�U#�9A-������Z)z�{SeӇ�r��S��E�@`J�%�9���c�3�8<�d��1���Q�!��?>�K#�R,�����o�/Zh���;.�^�����6�DH�
((V�E�jߞ(|db�40O��#Q$1>3%��43v�5#�'$"B�I�rW����H�,O:�*c�VL�Zѣ��L�*`�ǕxZ�&)[&o��S�'k�H)��iY�|��0dm�F���&��QaH�O.�o�p�Oڛv�m�!J6Mp��;0��'������S����a��k�<���JZ����x}��
*���\44u�)�΂Q�!�!�I�c]���O8���D�1=0 ���$�x�����[!�D��̠eH�|�Vt#`�� �!��]l|@kc���x���*�<�!�ˡl�yq��8L�����
˷ _!�Dֹ2w�|��Y�2}n�IG��<u]!�dZ�[Ɛd���p����ݽO!��W>]r�AfE�+k��	bg,)N!�� ֹ1�  �=�.9���8ZP��q"Ox�:f�9j�R����A�T6Xل"O�8�L�b0�U��.90�Y�A"O��q�Ş<"�Z�-ȇ{+�dS�"O���peQ�q��Qf��(qj��"O�Hk�
C�@b�qH��D'hQ�,*�"O�8����5h1�Ad<Ї"O�q%���$�àO�4N阶"Oʔ��Nm� �� ("��2"O�	r��+&)�)�V����"OB�ʃ�[$`0x@�2kZw����"O�� �-�4"� ���2)�<�#"O�mB�#(1���D�2:� hH"O�S��q�.(�C�7R�`�"O,pTf�p���b Ua�D<j'"O,1Y��'W(�h3O��z�d��0"O�E��C]� 6�Sfϖ�4v��"O��{� ��|9����X�|,ä"OPA�3�� (�`��yxv�YU"O �a�L��eX�0�Sonٱ#"O���+�����%��%e�d�"Ov�S��A;~�X�YG��"O���*P�>�|�A��9�7"O�z�"�k�x ـa��S Z|q"O��$�
Z��<"���fﮬS"O¨Kр��'�Y�RN��[ "O���Q�L0/ ���G�r�fi�"O�4���
~�4�[4[��S$"O����Ӡw���ӭ�7N2�U�"Obm���]�^J�b�L<qD��x�"O�8�`�Z =M9�f�6 1^9�"OLu�s䛆u�Ղ��E �|1�"O��1G�|Ċ�+��*B}r��t"O�Hj2$ܼG�L�녔�b#�"O>U�3�O�>�B"��-$�I�0"O´2g�-u,�8jg�Q�A�HP��"O`�b���4�&��7M�r�
�G"O(!�biN1>j+\�L�*Y�s` �yr���z���#SkɊ@�*�S�hǽ�y�E̯x���J�D	|ax&�-�yR�G�ke|��׈U�P�N��1iң�yDכ1.�3M�D��l�4(��y"O�5~2Zqn8:�����N@�L!�Bk|�}#���QM�m�wg�^�!��n;���3�_�H�j�I߄T�!�2�AB!��'>��a5"ޥZ�!��ϸ �Bت�@R�W�~����e�!�$H�U�8����=�v��"UA!�$J�Ƒ�ԏ�2a�.�ՀP6M!��)�к��ݗ*u�*`!��U�8�dqs� �k�఑�DV��!�� �z�3���7��ਅ%G�M�!��i���[4
T�.�Xlc@Cߵ|�!���&U%�Sl� 6�U:�h��`�!򄁳m �K�:l3�����!��ʃbKn9�A��I=ޜisC �!��U)Լ�ąƒkET�c����!����,0�T�#W?d�� ��%�!�H-d�v�J�O�5*t�"��I)~�!�D��2�QSӄ�|�%���
.�!��
/�vD���V�t
:�Rd�#�!�D�|ư��E*�B'�	#$��"`�!�_��R|B�jM>�ݚ��B�(�!�d�AE�͈VBg�*�ˍ5!�� �A�g,_B�Zd����8�Naz!"O8d�4��
h��yzC�Y'7�क़p"Oޱ	v�N�wc��[f�N���$K5"O��2�#�
G�}�T)�*7�X�Qg"O� �Ţ����H�;s4٨�"Ol�0'��AQ.��"�	,~X��"O2E˓I��3��D�p��$b"Ob	AP/��X��*��o�HЈ�"O�9�p@ �k�(bp���P,�"OB�hCK��tn����N^�N��z5"OX2��P?��e��CǓQ�Za!�"OP)�s �(n��X�b˟S��dhf"O����Nӑ>��y��܄�ީ�"O(`x�	X
��d��b�o��3"OJ�s�'˞V��;F[}nQC"O��X�B�G,�)��&�]RH�P"OUT�/B0�#�J�
#bu��"O�Ep��G�&�	�D'P.%V��B"O�`uӗUQn�#�P$+ �@�"Ox�a� L�<@�*^��5��"OBL��!����Ƈ�%5�v@qV"O�ԩ$F�*-�U����>���q"O�� ��4W��{R��X�"DQ�"ODa+��	p� D��+X�g�0�J�"O<�j���!4�<ڇ
3�Z�3�"O"r���,ed��%�J��e�a"O����-DꞜ�@� �Q`�"OU�
@ojA��bǴC
dІ"O�0��~�|@��C+�]�e"O ����$���C�*+NU�A"O�A�b�%|����� �6���"O,�9T�
4hPT��ʀ1��M��"Ol��fo�>9�4j��׽5m����"O4�j��#*޴�:��F�*v.a#6"O`��B��W옡G�\&t��	�"O��,P�mGĨ��"�8��  "O����#Nn����w���F!P"O0���dا+:�WO�c�b�J@"O�,C�]� ��݉$N Tr��c"O��!�ʗIY��͚]���(a"O�,k�)��)�4����|�\B�"O�Ȁ�dM-J�e�Iܫ~	�X�"O�횥�I<9ź`�Y���aV"O^I�a��Pߊ�S1��#�0�"O"���3' Rtk�Y
���"O������
�x��B�DKr�`�"OX�@D_�J�dxUHS��"`�"O��4�M>�JYCrȕ�Z�Kʍ�yBI�l	���:j�V��C�\�yB�U�:r�Uh��N]0�㗶�y�I�S[6E��Nېy�R�
�yR"�_�4(@`�F̐�㌏�y��ko`��(L,=��U�#/ȱ�y�n[�'O�l�ŭ�3��H�����y2���Y��Ea���,%H����*�yr�B
�$\)���#J��f�(�y�ެMj|
��]D=@��(d�B�	f���V�6��t��ͣM�C�I�.�Ե�g��hЌ�i� ;�C䉨O�<�p"̚?J�:ec���3�lB��6e�b�qtM*�"ɳ&��Z�^B�I!@��)���f�\��7`�0/��C�	+n�n�� Ɯ|����+R"!�ܓ(�N�X�%�4��!B�08f!�� \��A* a?�m�I��N�:c"O<�1��_�`N���) ���5HS"OM�愐�g�h���ْr��u��"O��P��O��2�Nʜ9��"O
�
�*ЬH@ȸ#d�A��8�6"O�8 �/KH��!g��8W`��˧"O�����Y0����ĳ���ɨ$�!��3�l���(g���ЎH'T�!�$�<�l����"%�e���!�$]m�V����Y����d��!x�!�8\���s��Y����
]�P�!�Jc���4,�"�����d�!� ��5%̀	Z���J�y�!�D �~�M�V��(��Q��A�8G!�D�W��`�
�+�OO5%!����)f!"P*i1��!��=���{ad�� ٲ��
,!��4<��+�iT�H.���!�.6�FH�2n����q E�5�!�D�@,z��t��S�4�kG��!�d�*
���
v�K����q+��!�d��vr4�)��(Y
�H
/�!��"�s�}U�	�/� ?�!�ĝf���0U6[��-�2s!��ڮ��ܩuK0�.�#N�7Gd!�DL!~7�]��NQG��9�*ڨT!��(J����V*�)f$����!�To2TZ2`�.&H���� y!򄍽@��<I�feN��1m��!�dEkz��ҽWf9���D/9!��G�v�p,{6�[�g+ֽ��j]6gD!�ǓK`��i��s<���R�>*!���? (��ҎQ�@����4�!�E�j���R�NԲ>�hAZ��ƋR�!�ğ
	x�Pg�N�����l��7�!��\�|Q����_)=�&@v����!��j�F���] y�Q���2�!�D
R�D{Ăוq�F��$��>f,!�D�tC�P��7&�0�E�\*!�� ��Œb�F��D��cY;(!򄋂4I(Y��CD	���6��%�!��W�\@�<y%*[Mp�(����JH!�Z�K_u��m��ub��Ch�#����	�R����'Ӗu��}A3����y�(T�e���Ԯ_�_;��cBl�y§L{B�@� ��R(�YP�H��y�����`h��{,�m(rNF��yB�W$X����B>"�rL;����y� U�n��:�P/[��p���y�9���ҐD�P`�!�g�̀�y�!�2`���3<��K&[�y��[ I���`/<�VTq��R�yr�ʒyeJ��&*�/y,yPdI7�y"���K��dC��H� :Y�u���y���8q�r`xǤ�6�Jl̑��y�E�_� ���gG��o�yb��^=��0Ҧ�4F��T#D!�y��i�jYY��/>)P8�S�ybH̿Lg�%��2��[B�ұ�y�,�bȠ��`DJ��͹�ό��yboU:
�Bpx�JL~�F5��BS��y2�]�%�@�2��uF�E��U��yR�]�e�3X��9�U�L�e,8i��W&�����,�ye�y������"lB@z�I��ɥ�y
� 4B�g�%H���oR�R�ʵ"O�E f����r�L�9�<�1"O��C爓�.�\a��X���!: "O�D�u'�HO��CC�W/g��9�4"O
� c��D�,�RK�/�¤C�"O4Ej�bH]�L�fHV/��3"O,�Ѓ�M	+<���ါ�.hY�"O�X�܊el%X��˗ ?d��"O.�x�M��>Un�Z!�%/.(�'"O^�3�%Z�;3���p"�R"O\䱵i��Dc��bi���S"O|�(j�*;2]{�c�l� 8re"O>�Y���~ڰ��t�
�c"O�I���وL���{i&@z�Q 5"O�Y�k˱%S���ǲSu�J4D�؂���.t��t#ªJ�����0D�����;;b��k7e�%z��,	4�;D�D�Ν8�Lq�h5Y��( o<D�(�"�[�(�����Bа P��$D�����	��C��L�R�5�?D�tN a֖�j� Ȓ7B"�Q�<D�0��C/'hI�+�:cEFt
�l=D�0h"���k$��j��('&&ʑ@!D�tkB蘰^Y^���Ij6 ���:D��3���v�Ҽr�H�*!�P��$8D�`Z6��������<<8�i*D��a�+��T�Q�Tr�<����5D���@�K��$���L%2�i�o1D�\Z4���Pґ��U��4i&�<D��Ƀ�14�B�HC�.��@m:D��hF�/&������=���9D���qL*znڸ���*a��� ",D�L�W�E�
�Ȍh�I��xu���L)D���U�8���ʤڟP� 27�7D���4��v�6��� X6vu�V�6D���f$�@K�h�̂-;j� �5D��ZdEY1������h���G�%D� 83�%r� �Ɓ�gb|i��(?D��V0x ��c2M�v�L��'D��� D8b�T�1#	�2 0�� �'D�����3e6L)���h (�m#D���@C� �y�+M�dZ*��g D�4rt�ۥy"�P
td�2g�.����,D�D)	��/S��ʆB\y.�; %)D���4g�%� h�C��[��I�.(D��Db�,dB��!2�S�3�] 5�7D�h{�-ΟZ�TX䐡�^��5�2D���k��#"^,0(2Q�<����%D����E�'�օ���T�	��!'"B�ɩ;�ذS懆�
�j�l��K�,C��*}�Q23�Z�8�ᄊX�xa�C䉎z�v���Y� �}��n�?-�nB䉏N�nfgZ)	 �\�'"šW:B�ɮ+JF���ň/_fn r��FBB��:(>4�yR@ڳ	2hFC�I�B䉡��=�4*�4M:0u&��A�(C�	�.��T���
9�$�3TDM�bL C��0׾�:d�0�GώNQ��E�1D��`�$N���ZeE5�2DM��yr�� F뎡phɢUb1���=�yRO̩l]��2�,��H���$�S0�y"�ǆ?�f	#GdP~)V��-F�y����%���1��é?+N�$C]�y"��f�x���HB�o��Ÿ ���y
� 2��U5O�`�1�C7*~� "Od�#�ȝ���H�H��b9�U���B��g��)c��QA/יP(��v�������@\Z��1�D(��
�v5PtN�1�>�i�\*nG~Ņ�4*�-��#jx�(I�m�7�4���n5uٟ~ԁ���%`�40�ȓ[�ŻH*W��� �?I� ��iզm#�dؙs�j��o��/��i�ȓRIj�i1��;fN�9J�ǔ4~��I�ȓ.Ȑ����)j	�˔��%b0�ȓ �
�Kҏ\�,̐���eC�R�L��ȓ#VPۇ�G�(18�[Р��Z!He�ȓA��]I���$1��yD��9ⱇ�?L}���ʠu�(e���=T�nц��nxq�$�6\����C��_1BI��a�Ν;ƈ�2
�$hPCE�`�2M�ȓ%���K��\c(�#�����q�ȓ5�b=�	x&��5&��d��i��H���6ꄕL�&-)фhI��b4��˜:5��	5��so�A�ȓg�(Dp�*���,�`e�ȓV0 �؀-	W��TDȊT���e��`@����h�� �~Y���ȓ:S$�!���,���(�Ոr�!��K��a���{��� �BA�'}t��E�,Hh�˄=+(���?~�\�ȓ(�=��A^��,���@54��ȓ>`���F��,�n��ƛ�D�x!��m�b�Hǎ{�d5	R=㾝��xaJ`P�ɓ�eN���5.�79�2M�ȓ�|X���?9(ăE�HD�����J�lA!��t���9�*ӄw���ȓ\�}�(�"]{�ag�D�`h(�ȓ)L�<��:!�������>8��w�p ��0Ղ1�̰{NV,�ȓ^#6�xdl��Qg`I�!ǋ=�����)����3�lt��ˑ@V�Vr1��uz���4m�90�4tK�*��%�ȓZD��!h�z�v�@����4�P��ȓ]5z��t��#A1���GC�*>z=��6!x��/��8;7���3+�<�ȓoq�<�T�֓r��������P�ȓR�ND׌��f|t��3�A:2�M��	�\�egF3�Vq�@���~�����8R�,�Q�(<�d`�%@����m����3O��"ٓ�a�J�b��S��sr��0R�V�P�<?25��HM�� ���jnD��@VN	��$6x�2�`�*X�x����$�bi��^�TZ��#c	�xG�	k8u��|�v}���sgJm��;X����,�f���@��j�3f�8�<��QK(}�ufD\����䉄�dmI��r�����-S7}��� J�}3�(��\�|���2E6�@�ߦU��фȓ	���2��P��L��h�.r*��m�N��'*ĵ]6���l^(j�t���c*j���R�F�� 3�/��I���ȓ{�Ik҈���x�A��?����/��� '�I�)������4x���\4�qJA�8�4I���ˆ!*�Ȅȓ[�҉A�GB�b$���m�n4�ȓJ]r��-<�H��")	=jP�5��S�? ,H�k��CU���.��*Ҟq��"O��
�LͼT"��Sq���𕢶"O������5�<���cךX32ѡ1"O�Y�`�DoF��P�U�f�h���"O Y[Q䒋<�|����T�
(�y"O<p�Y��d��� �T"O���ȨfNd���
5#ǔIj�"O�̓�����j�>s�i����#m�!�T�Y"l�"a��h�+�$I�!��@�:�:�i�]Kb��׈�u=!�S�dgp�Bf�=E� ��%]�w4!�߰4 ��1J��1tM(���g�!��سOdq�`FA�K�P�9��S� !�_53>ʉ���,(%D|��|!��\� �x���_+2� ���M�!��>3��q�@��Ln��*�G�!�� ��$;sA��`O[�×�!�$˵~Qj��W�*@vA3s�W'�!�� B��(��g��#�����^��!���)��-�f�P�#�nQ ��(f�!�� $8��f�z���b��&&!�5�r���ґ+�V�!��/�!��_�f��Ũq�P�0���O��U!�D�	(��(����2��
�G�Ui!�䏆h{P��&I�t+2(�G`AM!�$ޚ��{�����ӳ&cX!�N�v8��ƬN�M�,Hj`#B�!�Ѵ?���2��)mϮ�pϟ�_�!�䜬%���C�[0�{�cޖC�Ɍua������x?`��ǦB�\�hB䉈}����ӏ\�⌐�L�p�C�I���Ģ�j�vm�`���B�S��B�	
S�`�Xiэ!���p1bM[��B��/�а Q� ~��@ˍQ�$B�	-r>l��pD@8j�J���ԁZ�8B�I�d�>]�׭5(BMZB)/B��3_Ҋ���ԍ=��B#bSv�C�	�=� }�o�:A�ys�_�L(�C�	:@mZŊ�l����:������C�	6W|�P��l(�I��*H�7��B�ɦn���@�?x>�]��� \��B�I4�}�X}��
 �Ӿk��B䉌5����9j&>��5	q�zB�ɩ;�6l0g!�{t��B�L�0�JB�ɗpz��'�6&�j�Ʉ+�zC�ɾA�Q�1��nA�q@��/`C�8f�U��¿%� 4M�70�C�85�<� L!8�� �t¥o��S6H杚5�!F���� �!��d�숖�[(��|��S'�!���"s� ! #4�4,�����O;!�DT��A�a�>y��=(�$.W!�<�\X���'*�^A��j�$!��Evx���჈�X�+TD��K!򄈭ft(�Ő�m:d1���^!���	��Xٖc5��y�w��5z!��BVaV�u�	U�<��2�Z�s`!�DҮ����%��y����b��"c!�Dז$_"aX�h\":p�Z�&r!�d��"LsJ��+u���4��X�<I�$-�xB��/���۱Hi�<q�KB�n�&m����)'��K�F[�<�e�S tln|a����;��s�<�[� �[�Ϭ������>0�B�)� �����B��l|��+-C �%�"O0p2�̛~��1�,s�0�"O:�0 kA��#d�+�4$��#�6pQ`ɹ���L(<O �@.�k�"0@C�,��y��"O�+���6M����N�$�*QxF"OLX�����d4�n�%4�<}��"O���2->A|�T,�0^^���R"O�	H�F'/<v@�G+�f��e	 "O�����8P*�՚aJ�=i1�<��"OƤ8�.6Sɦ�q6�JR b��e"O�X�u�ɰj���1�A�{�ѥ"O���$�;_��5y�)�<��C�"Oj�rsM�<�4��IS�U�%"O�#�VN�}��犬JQVM3�"O��Ã��&�nUcA�[�r���"O����O�?0�!���m|Ux@"OЌ SdURk\��!�� ?x��v"OJ��7ܑ�i		%��9d"O��3��ʪB�d�Ȳ���^�K&"O�p�!iI���<�a��&5���c"O���AL?\���G�U�B�p�"O�a�� �S���r����PS�"O�a�#�|{���G���	 "O@��!	�u�tps�B¶�b,�V"O�9�\(+oZ=��@%6��0@�"O���TDŽG�,`*��-�"C�"OV�a�Ê^���U�+~⡸�"OES�D@�9p��*M�xh(H
3"O*QGDX� �F�:`g��3n)��"O0�j'�ַ{^�X�C�x$��"O��R�K٬|���F��y|�]J�"O���!<.������(]��S�"O��2�J1Z|]c�i�*Ӓ%�a"O ���"9\�R��S�*B��"O�H�%��y����&q1�"O>�⠊�pG`���j	(�"O8���ӫK&����L9|�\��"O�����F6�LQ�D[%_��Pu"O���@,��CŌf����"O����Q9M�܊��e��ɨ7"O��7C��;p���b�Q�F쀥��"O���(:_D�+5g'+�u٣"O��9�U�-��qQ B�l�x��"O�P2�Q�� M����DA�̊U"O�E�Uè�����-�,�p�"Ot��UB��|hh �6�u�RX��"OB=�e,\-9lfLIЭ�9�v��$"O�KR�-V�t�pl^=�F��0"O|�@DI]�-IǪS�!E���"OZ|/Y��(�A*�!�X��FU3�y�ʊ)H6�`��dY\K�$�y"�@�@��ԧڋU�҅�GL��y2��<�l=#s�^�?n�x����y�腌0m�ط�"8(8aXwꗞ�y�l/�J��bl\	`atX�V��y�.0_z�kGl�Z��vƐ7�yB�!z_�:�Ώ�Mn��s�L3�y��\"]����k�8բ����"�y��n�NT*`��'-�ت&iK��yR��# u�d��"�NP`� ���y��2!���׼� ���́O?��ȓ4���!c/s�V5)���2:�V9�ȓ��z�D��y�p0 U2&����s
������.1PUZ�#��2� }��S�? �9!BݝFx��g%g��|�"O�h2�O�*G28��@7c��(a�"OPu&O��`�0�2��t9����'x�@`c�ŌU,�A
�j��4ʝr�'JA��	xUF��IH4$W��@	�'�d�;1e��W=�����S��0#�'~(H�����lԺU�L�w6 ��'14Ab�o	�$��@uDSt\p	�'1<��p���}��@N�e�f�(	�'�X���%K�m�L�IQ[LyS�'��y@&؎W�\i���]Le�
�'ݚ�H�A�Gc
ى4�;Y6��'Y�T�W��M�4	D�BXL�	c
�'���0w��'� �@5Wx��a�'�(8#T��5r�؝�#�R�"��'��an؈\V$��%��Wf����'�ڹ�E�B)�Z��F+T`Ņȓ*���2�@�p�h��P'tV5�� � ��OuS�P��b��~��ȓR���0G(���Z�m� �l���Q|����su��b�i�y�dY�ȓ[L�A#`'օ{~耴�ů*����ȓJ��H��j��0� ��bmL�Zi�Їȓ\!I���	?}6�pA�� �zi��e
��h4$]�H��u����6�p`��J��l��� ��X��+%�¼�ȓ#.\|y%b�9�\���԰s�H���u�����n���}�DDD6��؅�#y@y�P��6
#�M��i����4+B�ÔÅR-�Uk����SܴY�ȓC�� ��ݟ.4���KZ�P�ȓs��:�O�֌���>g)T݅ȓ���*��m�|�
�F�7B:P���p5�� �䔪r��]�w-��5��݄ȓ}$l�0V�)p�����̱Q*��ȓ5߀HJDꈊi|�TA���!�ЅȓJ�\�D���@t`��ЈP7�-�ȓ�d�V��g�F�&gow�Նȓz���H�/��[afP{�n��9WX0�ȓpB���@Z�����R����zBV$a�#��5c�*e�i���� �tb��7F�ir%��@$�ȓ+P�lid���cRq�#�����܇ȓ]�>�C�d�n�Qòm��Ӫ���B`�zD��0K�=#"�B�aA�e�ȓn*(�3`��P�Q���P�_h�@��?���3���H�CR$>��_���ǩ�3��� ��'��܆ȓ3��i3Wo��g�N�8��[�t<��ȓ#EF�@�,|���@ �6X����6��1i�H��1u܁0�lGTjp��a~�� ��EC`�9�UQ���ȓB�D1�h�,fE���(e5���ȓR������a�켹��˶h� M�ȓ
���̊8)B.x���E+HJ8��ȓA���x�^U���W=n1���ȓq�Z� adS�9�e�۝\0�ąȓC�qx�Kڗ'Ll�	�K\�J׌!��yU(P��LK�.Z���@�
�'\ў"|��Y���IboK�����B�<)�&��A|q�c��Z�hI��A�<1��rd�^�H�<��"�Yt�<����,@��X�FB�P��%(�s�<���"6��1gn�zQC�m�<� ��qGM�w�HA�O�^���3"O����F�B��r�΍�z�rP�"O �±dߣ5jN$z%�#+�pX��"O��d��"�(��p�P!*�V�["O���.��$i��@OS*��"O֑�G�W�Ų�fA�֤�*u"O��KB���|��E�'3�4�I�"O�1���|��Ey�D��� 1�"Op0�*߭���;� 
��@�B"O��fшX�,�`��6E")*�"OFi�P��٠�:���(�R"OR!��{4hJ����1�d��"OJd��%��H�=Z a� �*e�"O��kUw��(�/k�T=�"O��UD�%X���`ρ1��5s"O��[ta�+����[c�R(��"O�sV��.x�:����-~���"O6���&J�N<!F�JJ��YB"O��@�#;?��a֣�C+� q"Ov�#��q&Լ���Ӆ���"Ot�c\jL�zEaĶ;��8���A��y2�[�:+�Z�F�AV��P!��y"HJ5ehR��#ں%��|U+@s�<ag�**���O͍�F���E
X�<��o�S=�t�0�[�I"��e�x�<q�EٜN} �EQC2nTpE�Ut�<�,��[���y��N$�.��4GL�<ɳ�G�7?���Ǣ�:����Ph�F�<�d����@>h�biᕫ�g�<�#I�?U����G�'�� 9�Ma�<�Ӭ�1f��}X0IA��� �#��H�<I�)U�D�Pزdb��J|�-�Ռ�H�<fDŕ={����,�'�)���}�<�0�#Q�JT�e�;%���8���{�<it��l���T�ضG�,mxQ��z�<1t��^���Q�����e��u�<���,?=����L�&x�l�vALK�<��N�H<�1��@�r�Q��k�<���3u�<��G�[v��Ȋd	�g�<y�m-^~���@1�f}�v��n�<1�eՅ'�i� X�e�B}�eaMb�<�e mfa�fa�%b�`i�7�f�<A���w��a2�g�:
�HT�1 �c�<Q�O�GsZ�Q��93(r���Bu�<�S�_���90/Z8�K�LY�<���ּ<{� ��U�+�0���QI�<�����:bbP��I	�d�_�<�RIԣ�����gR�Y�0�G'WZ�<)�셹 .��a@�,P�1x#��J�<��nԘ8o���Ќ�2-΀�i0�E�<y0�LV_X�z��o����ď%T���%��:�Esv�E{�\�)��(D���v��
D�
��'��.�2���&D��FeK�X�*�Y��E��"�!(D�P1���'�@ᚖ	��2L̴yc'D�����C�଺Q�ߜY����o/D�$�C�8e�%�^%�f`�d�+D�LR�oW�k��	Ѕ�ێr��Y�Rn=D��Y�l��(��w�Z�#��x�!8D��X�ɷ*dj ،�V�S1�5D�ę�l?IL����� ꔬ3D��l�K9Hi��ǯCª$�YaC�I�VDdx1�䑶:f�2�� ��C�ɼH�|�V&Y0 X���F�C�)� ��Q�Q�@4K a��v ��{""Obp��폭P/t�:A�2��g"O�-��%הmz"yieG�д8�"O��-��'� u���:F@k�"O���DQ�T̛�g)=^Ni�"O��v���p��f
	cu�,�"O�)�E:��}[U� �\��3"O����A�}<�y�Gj�gI�es"O�uaT����J�i��6x w"O��T"��[XT�A�H�&NV5z"O�H� ��lz� �⭆�25��3�"O���ã@NH5Q�OW�;2����"O6|��G�^ݜQ&�_s ~��F"O�P�`��#e2%;4�SjJG"O.@�4*_�so�u�&,��"O��"7$�a<���G��t��XIG"O�aC�NT�5�䲴�Ņ�:�"�"Oĩ�G	H�<�ɥ��6g	d�"Ox�;fFN4B���C��1����c"O
��P�^�p��g��9��"Od��F�����^%,x���b"O$�ۅ[�[�]R�i��f�܋�"O`�ڄ�ݭH�Q7�7�x)ç"O���{ b���
�>����E"O�]x�I��Qz��!`.��ʴ�f"O������9��Q��M��.|^�z�"O U�d�� y��+3��8^a
x�s"O�`�TBțtB�8
#�Ag,�)I�"Oti���r�	!��T<H�<Z'"O�a�g�Y)Ԯ�ӊ�(x�J y0"O�T"�%�5isV��婏�)�4�s"O�	S�+D ��a��狽V��Bq"O<��r^$Xm	�f�6~��`"O�A0��%\N5*����K����"O2A3�K�� 0�#�
sT��E"O��!���xQ�S#�?0Q�@�q"O@3�~cl����HT��в"O�%1#� �H�v�:~�d���"O�i3EW
}Q��R�J�%9�"O>0��W~!H�B�g�L�0S"O����Jh����T��7�h�pB"O��� .F/_G��Q�`H�m�e��"OZ�b�SPS�� q��U��e�4"O���rkA/ :!≇9;w�9��"OBU���{q*0�WGG6uh�H�"Oȉ+R�[��D��'g�OOlX+�"O�쐹zp��(��T�<됍P�"O6P�sGD�a���y�nk�@�"O�]4̔�?�}�Q�''��� "O�1q��@�,�rH���ȵpfh���"O����yz�f�ǡc_rp��"O�y��勮y&�$����6GtD�"O��X� ��?��#���.r�<�kG"O�]��b����0����"bB�qW"O���q��4���c(O�T���p"O�0jAKա���qFiA
e�hhI�"OR���	2FG$4���f��Х"Olp��Z>w�b��c
�A��A��"O������&���'�lP�a"Ou3֌Ȼ,�:#G�+<����"ORt�0#��r=���V�X�ror5R�"O���ՁV�ݞ�GNߔ?�$A��"O�PZ��6:�����&)�d"OHm:rʇ~���D�+�D�w"O� @h�W)'5>�=h��ИaFRmI�"O��H�@�P'�4((�m��%!"O`�Y�"P�QB�ѰA��\uLpb�"OV	C��u*�A�`X�i����"O4��d���A��9VN�d2�"OVe:��W"4��͢��1T�,CU"O���3Ȕ���:M�9>MP(�*O*m��DϪ|�	Q�i�!�Le!�'c�Mç�T ^58���A�D���'DL1�`k۽)�,��%���g��{�'�~��	!7��(j��2g�Aq	�'����ɳ0���B��)3���'(��8�a�6WFH$�PE��q`ư��'�[��L q��lR���m����'-"05O*��:�#A5r�>���'sr,k�e2gN����L�3�l���'(�}�f
00Vt���-I|�
�'D�����ۥO)�Ax����_~i
�'s@|���Ζn9|	y���X��h�'����fs~:�:�\�s܆T{�'�A�B�(ԾX2#�&h�,���'f(�yC�ї=T�x�HO]��1��'����a�"qZ�	!�ժV�ڤ�'��|Z1���$�1�U�U�bX�
�'0@L���=D�|�#QxUN�`
�'7���S���c�	�zk2H�	�'�JU�U�vǜ!c3d_�r��M�	�',����c �X6�ݳn���;�'����%��7T��OͯB ���'Np�D��\!C��C���'��k��I�p�H���y/ȅ�'Ɍ)X0���Ѧ9!#G�@�n}��'vB�Cor ��i�/�>�`:�'�4��*Ab���C3�� ����
�'{�����T"$et��)B�~z~yP	�'���:��^�v���j�I�7j�=��'�Zp��oǏX`�@��U4<TyI�'B�-�`Õr4z<! �R*�T���'*ʴhV�˳S�&�I`灧W٬<Z�'An�:F��,�2�����S��E��'v6%rA�q��-{Ǎ�	HP 4��'��uk��X�~8l������]�
�'��E��*
.-(a:V�C�,���'���Cڿj��	&�K�mu��Z�'q~D`	�~HA� *��| ���'T�E҅'Ϋs7����E�'n� 8��'���� �
�m�IRX���Y�'w���aA�x9��P�Դ;��x��'�֕i$��+jh	 ��H]��a�'n���T��{������2:0�	�'L�}"S�5���!R��)%�!)	�'����%H
;S�	��"�Re�'�(�A��֔S����!oC�eHs�'�HĚ��C�D�Mڀ����(�'�ڽI&�%6����$V _2;
�'Q��q�)ܜEJl|H��0X�:)p	�'9�d ��?>��ua�)=B����'��X��:8r��!L�;�@H�'p��j"U�8~nPy��*�����'8�H3�B�!I�v)����V� 4�	�'Վ�1��!e>���SȌ�B2Ԩ	�'z� �b�M�`�0���d��x0ޠ�	�'���[S���w���aa@k�l�'P�us��L���{F,�1vz !��� fM��c݈����FE*qS��2"O��3bɟ��Q)C��X:8�"O��aPᗢ^�&���3l�hU�5"O�H��%�?�����C��4˾�)P"O����t�fH��)́s&y�"O������L#\��(�w%mG�VX���ʐ5&�T+r���x�� �3D�����؈*b�7�\�U[��]J�<9קėZ�͡e��7���r��{�<��j�z�EH����a�jCJB\�<�]�\26T���7af$Ò��r�<�"�Sߢ�ҲDر^; 	S�� C�<Ц�Z;�-�$�ͱ5T�����@�<�JF��*��kƨ1�a���\w�<y���?U�ĩ�V�EԄ���{�<�ˑm(��t@\�P�2���AQw�<pBP\>.��#jђl�*����h�<�1�R�1v���ېnt���e�<��*�;���;,��YcBēe�!��4">6�����w�@;�g�Q�!�\�-�J��Wb�i��;� ��4X!�@<?��p�v��"�8���1U!��˸>Ǭ4�ևN(f���qp�A4,!�D�y)20)�ƩK6��AJC�R�!�]$q�2u��@P���z�kY�!�{֌��$I�+�̀�
ނ0T!�DڅW����F�������#!�d�2r�������7�
�A�؀#�!�dK�A�"i#�N·5�
H��e�@�!�d�5$���f�~��ӀM=�Py�� �D]\�{v�-��D��E��y����H�q��cR�
и�	�Ԕ�y���/�.`a�f����tI�3�yl��*&��F�,t?�L*���y2M�5��1�:h<�8�����yr ٶ;��6��6M�D0k�bO>�y�jڄ!b���$Uƨ�!HȞ�y2��';�<��C�`Xhґ���y�L���b��ǡ��,��]9�'�y2Bvg�Pq�(^�^*%{�!�1�y���Y@��h%�ꤻ����y��ۀLu�lxժ�� A2��y��ϼG
��&���1f�+�y�MR(��c��u^�i`Ņ���y�蚁P�j���%N?�-��;�y�`S;5�Q7H
mR���*Ť�yRnJ>7��p�X�i�����@6�yb$�/�<�����|�B0�C]*�ybd��Q��!�E��
���JB�=�y��V'\�bU�u�,3xzag߂�yR��1�m�'��*�����"�5�y��I�t��sጋ3�]�Í��y+�R}�Tc$
SԞ 9î�y��ּl)��'O&�hs�
��y�NF�s�T(�&ʝk���G�V��yre '��Xb��m�|e��J��y2̊����_~�x�A��yR�W"K��0W��0^���0�O��y��$#<Ty��R�
�$IC���yB�� ����h#L[�@x�+��yR�ȕVц�i�C�w�qz0��
�yҏ�$kX>`�׮�p�:x��yR)R?M���cL�bL~�ꙁ�y�Ɛ�>e��D��)5LAx�E�y
� �=�A�
Q<��;�ᅜz�!P"O��c�����ꜟ���Ґ"O�X�1��O��p��B�	�����"O��Q�E�>Ei�N�3�hU�Q"O�Bu`�|I�J�*�^�ptJD"OH���� � �:���h"O"pKW(I�j՞T!�ӹq1�(C�"Oڐ2ōȺ?h�Ÿ��_�4'�x�P"O��A�hψ+�+�	��Pv�hE"O���� �}���CGB�G�T+C"O��z�˟5�H�8#����J��O��������M���M3�_>�q��T����������
%:�(���I�F�Xq�e� \xԛC%́	qD6�U6U�h賂�N�+��)h�Y��m�9�>��'�"2�xBCn�&�����آ�H�g��7;�����֋Dsԭ�~��$�J����!;鄨B�.��m��U$�d�Ѧ%�,O��ޟ�����bơ�+�/0���?�~B�'�a}2��	3����&��) �<]ⱮG�(O�Im�/�M�J>���u��Ʉ{�}ct�Ǽat��`.�|�d�O��T��:�P���O�$�O�ͬ;�?��>�01���M^HcB�HVZ��`''N�҄��DU���[��:�&9�fJ4���jE?=�H��u��?���q�c�)�F�{�Ț�v��`�0��~�'$���'!V��UOY;�ȅ��V�%��(�O`�y��'_$6�C�'��$w-�lK�#�0�B�s�vL�O>�
��X2p��%n[���@�BǪ-m�Ŧ-��4�?Y��i���O���\>�����0���b�I�pD�}�Vȕzު���̟��	ߟ�ɠn����	ݟt���S�n���ՕZh؁�ƲB��Њ�q�T!Qf��(톸Z��U*7Ñ��:UL�����
 $FH[u�ӈn�1�*˶$Dh=����m��y%a��HO��z�'���c��0����&N�~F�v➾ ;��'������'�p�I~���A*Nx���hh��r֊���yR(�K�>���Fį]�h��Ν�]���$C����4�?�@�irV$ag!t����O���w���r$���J���������F-k@���O��D��\�T���%����Z� �ÝO��@�41t�p���� ��p!���ê|cZ�!��W�#�UYã�wf�ZC��qrZ����0��5�bh!ݾ�Fz��Ը�?)��i*�7��O��'�t({��Ȝvja�M88vv��`�'��OT�}��Т�
5(�6=puCW���g�����٦��޴�M�2D3wk��"�'ͨK�������~?�Ȓ;a>]��?(�N�9s��O�dd����#��)��t�F���jĖ]� ����Ƹ;!�BQ��E�ל9sI��ݟ��'��]c��lXP�E�|"���SR�t�ߴ)n�ૢ
�tDX�@r�O��-�S�@8 ���k��kV��ρzB��P�պe�FM�?��ilF6��O."~n�Dd(�Bh�4ų�G]" M�	ݟ��	{؞$��,�$x���C��Q�q�d�&:ʓ`����y��O����O�HX����3D�̨�D��C>~)�D,�O
���E�xT����Or���O ��Ǻ���M�eŐH_�@��M��o;rp ��d5��(w�Ε~�p�%��H���O^0�Dx���8�(8"���P�ȠdQ�XX�6L�Y#LU��+n}�y��p�ĭ�)=�c��
�N]-��T(!���{"��1Q�>q��Bʟ|ٴR\����'k��h�B�ET�1!��pT�'fay�fȗU�*,�A�L��bB��jx!mڕ�ML>�'��H>�۴-�<� @�?�   �  ?  �  �  �)  .5  �@  }K  �V  mb  �m  �x  q�  ��  #�  ��  Ơ  �  g�  ��  �  A�  ��  �  g�  ��  c�  ��  *�  ��  ��    � �    :& �- 5 �> G �M �S Z \  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�Tnڇmp�Qq4��d@9�L��|�X|{��>?��i��O�9O>�D�f
ȩ�%ѹk���0���Xt�$�OV���x�����D���N�O��(���VQ���Q��)�y��'��O�O\����W�T�2H'"����p;��fӲ�1��+�ӧ�M�;�@|r�R�!���56� ��?��'c�)�*R9��m��<�`�GBؒ5�䂙� �&MxbM��<A�'/��D��hO�	�O��'+B�e�ݐ�h�	j����<O ������d\�Ř'�F� �#'�fƊ��x526�d]o}��'�27O~�t�e�qEϘ��t���U�	PD�'	r�J;q�H��t�
���H��'� D��D6�vIz�l��i���ؤ[�P�'���9O�U�����{ӂ� �,ͦ?ň���2Of�mZ x��}T�&�4�2�+�B�f� ���Q b1Od��O��$Yg&86M:?a�O�����!�����R�P���W���8J>	)O�)�O���O6���O���0!�#���[W�U����R���<	�iŐ)1%�'v��']�`]��)�j�	Q��:�<�m�U}��'��O1���£B��Ig�v9���Id�����<94��#���P>�����V 9nY2Hӱ(�d)�@K�����O����O6�4��˓i���Q���$%���%�X�!@(GN�"C}Ӗ⟤X�O����O@�$U3L¹H��ˁ!�p�B��W1c|�Xؖ�|ӊ�^���1Ō�F�>���q<00�&.F�N��1��1$��I����ʟ��Iܟ ��^�'&���Q��+ �Q�]�F8�4$�On���O1nڂJ��-�V�|������9���z�V٘&*V=,|�'�"�����K'Q��֐��qGf@ q���i�!���"�Jp�Q��O��O*��?����?���Pt��jY�gF��aaӴeB����?�(O��l�_E���Iǟ���s��`�:@e�Y:�k�Є��T���D]D}�'��|ʟ�M�����h%�Z9��H��ۤYZ4��4+��S�i>5r��'�4P'�`ش%�3F%���-�&@V��v���������b>�'/V7�7U%�|R�I!�PXhEJ%�F�(G��Ob��Ŧ!�?aQ���I�C�f�j�-���쐜Jτ%�'(����i�I�j����`�O��'~�c�A��x�a	�˚.<�H�'������ʟ����L��~������ႃW�t$)��ΘDK07mA]v���O��/���O��mzޡ���!CX8��D`�0l����U�ڟ��n�)�S5���o��<9���,6�aVCڷ��C���<�b�c4��d������4���$�A�,���I�^��\��M�9�V���O
�$�O�8��V�O>i2"�'�Rɓ6d���Q�X�4��#�c;A��OD��'��'��'��iX"��1�@a���D��d��O��bg�A,8�m� � ,�?� ��O��seB�Y�ȑE�*��1i�'�O��d�O����O�}�0��(p"&?I<l�qJQ*c?�5b��:R��Fm1"�'{�7-/�i�5c%��`�nscO]juEs�.q���蟜���z?\oZb~b�Z�F�ޡ�'q^5C�F	�G���+D�@�)A`!�J>	,O���O@�$�O���O�uÃ��?-)#r�:zfȘS�<٧�i�Nh�s�'��'���yr�ׂ��踵-Nfm��Rk�K\~듍?i����S�'1t�4d �o9(�����2Y<�ʶiR"G��,O`! ��Y&�?I��;���<Q��9qd q�-[97�^�b3HI�?!��?���?�'��dI���w�Mʟ�K�ԎwO��E�ی;.�;�(M���pߴ��'0�듹?A���?�Cۼv�2yS������X�J��4��Dѿ,~��ڎ�)��� ��P�o�\�A���M0&pԒ�9OD���O���O����O��?u�F-��)l���������K�$�	؟�Pٴ6&`|�,O��m�J�	�RW@H�&ޔ;��k��&0ɚb�D�	^y�.^"kC�v���+0v܌����?n��BI�x<s��'��&�(�'���'O�'�"���U�<�L���-�VP#e�'"�Y�\��4�bq
��?���)�6r|M��-��{�4XE���B��������O���6��?)0+�nTPD��Q�K�ܭ3���2�\cu� m����|��j�O\�aN>�c٨��dJ��G�"YCt	��?)���?���?�|b)O�)lZ�t���b���)�F�1��ۅ:��d��my��x�*��1�O��ğ�V'؜0C��0��� �H:+s�ʓ���4����	(t�;�� ʓ3�� �'��kN�|Rf&bv�͓��d�O����O,�D�O0��|�����x2�	�W��&* 2Sۛ�,�!��'����$�'�6=�*��c�_� q�Gԅq�\L���ON�)���Ϋ�z6�h��K��Ȁ|xdi+�k����Hv���D�4"{ky�Iuy�O�BƇ8���y�#ܮD��<i%aJ,{��'"��'剢�Mӧ"�?I���?фm v�J��oR)[�]Sj_���'{H��?����Cb�D�B&O�2?!"��<B���'d~$C�gB�p����9�i���~b�'�`i�f\�y��)c�9nZ���7�'pb�'	r�'��>��������ՄL�2��4j$��<���I��M�q.��?������4��q��cS�q
D�#�$\�N�>O6�D�O��T�{��7�8?AW-��H�iˏ8�.]�t≈72�c�[�=�x��K>)+O���O<��O����O���L�+�k5 É&�8Z��<�g�i��}�pW���	s�'oO��#��1�z,�ҩ�wP6x*�T����䟴'�b>�p�ߡX���؆��#6���C��lE�e��Yy��<lNL�	�Z.�'i�	�)l}�u�V	GDFHU$��S�B��I����I͟��i>��'27m 	|���ĕ
2ti%��>��K�/�*>X��צ]�?��U� �I����	*|pJy�Gm��"��MABJ:<�[s�RҦ��'!�  t*�?y�}b���~�#"��$���ŉH�j�͓�?���?q��?����υ�C���NN{b����nܽ{12�'���n�d�(e��<�7�iU�'e(�Q��5
��HR��Z�UIw�|R�'��O�����i��iݕP�J�+CV�5J������ˍ�@��ɡ$��'����0��ퟔ��A����  	�b��(Q�o���IڟȔ'��7��if����Ot��|J�_;p090�(�q�YslM|~�ϱ>���?�H>�O+�xz��րL\<��7�\�D���[���W��W��:[�i>�*��'�H$��vdC�J���`0`�C� ��Co ֟���ßD����b>Y�'\�7�ܗ�u�(�z��IA��$p�L�#R
B��?��:���d�N}B�'A�5��#?nh�eA�<�<q8X�d��*�Ц�'���Q���?Q˳\���@L���T��< pd�*i�\�'���'��'�B�'��S(�8�〓Xit5 �F��I��X��4i��P���?����'�?)%��yg��#?��2���6d�f�6B�f���I��X�p6my�`ؠ�ѭS�a@�#ӡU;�u���d��:%��%<�ce�DyR�'R$��'���14�Y�9�	*#l{I�I�P�	ɟP�'��7��2@���O���Xqu�`(�GՄ"���޸�㟴�O��D�O&�O��q!�ɑ1�pH��`@�Ds����0��h����F$m�S�i��$C�����d�1*��4,_?T<���Qmџ0�������D���',�u��$C&��|��?tDȉ �'~R6� YB����On$o_�ӼK�B���`��C���T� ��s�[�<	���?i�0`���4����;(*����'<�i2e���^,�-e`69�n�'/��'c�i>���ϟ��I�D�I a�K�d�}xN]р�������'S�7m�^��O��,�)�O6�2p�۩������.%H
�Pl}r�'|�O1��`�&�{�0�s��Y���� 雜A�`�G�<Y�hp������򤕰
Z�B��u{Zm⤩Ң}|���O����O@�4�"˓D����H�	��i^�_@���1)-7�(ػ�yb�i�0�4a�O��$�O2���^iI�@�w&�y���M��v��7;� ��g��aJ~*��;
I� �E��$����0V�qΓ�?q���?)��?�����O�@؂�.�B�����+Ϸi``j��'�r�'��6-זz��I�O 9ob�?v߂dp1ƪ
JX��B}X �'�X�I��S�k�t,nZ}~ݣ e�A�N�\BȌ��)���AD�_�0�5�|W��S�� ��џ𙔁O�xD��W�H?��U+��Lʟ��Iky"�bӲ@��'�OV�$�O�˧C��Py�C<S-����	�k�T��'�Xꓫ?9����S��N^YO��k�s��Y�&M��W�䅐u�\�Aq�X��O�I��?��1�$3��ՠ�c��0yTH!�ͮ{�<�D�OX���O���I�<q��i��M	��wP�aS��^4;��@�2�'��6� ��3���O��dY���Q�f �5�rd �&�O��D�%B6�%?	V/��g}R�>� ܈�U-A'al4A����:��5Oʓ�?y��?���?y����X3}~Ԁ��'KNK<�lDh^��o��%��l��ß��	p�'@��w�qqfÍ�������^'�%���'�b�|��4cU��8O��:4��ݒ��=oK����e?�yR�΂'�*��	L[�'��i>	�	���x$��9(��J�l����џL������'pd7�:=����OJ�$�)��9@�
S�5���5���0x�O��O��Oz�HE�rj�Dh���Lk��j𒟀�p����u�Z]�S����ϟ����B-�J�@�IȒp��������D�IƟ`F�T�'�]�P��0I�d���T�#�� ��'^7��	z���d�O�o�T�Ӽ3o�#@�4\)D�%B������<���?y��IWH�4�����H.�lP���!P�G�F�efIJ(��'o ���<�'�?9���?���?ٱjϏ7uh��%|�ȈVcJ���$ۦ��c��l��؟L%?}�Ia�UI�❦[Lbp����MU�I�O4���OВO1�l�h�D���R��;&����f��2z6�LFy2��64���䓏�ā�F)�]�1]&(	k��R�G�:���O����Oj�4���U�VI�0}"/M7|UQ����U�pi{7�r�R$q��xA�O��d�O��$W�P��DQ���g��9��-�5[�D��	o��,�0ճ�E4ʧ޿��
֧
I��R��_�X���7dS�<����?I��?!���?���D��)J)��AGĳP(�!���a���'Y�d�<�B"��<y�i9�' �H�D�-�\��3�#��h%�|2�'��O<�B��i��i�!ҔƏ�lEd9���A�bȬ܂�%�-G|�d�	�[�'}�Iğ���ß���2��x%��lvE��EU ���ƟH�'Cx6mC7B2���O��į|z��[*��ǯ)�%Rt�WE~���>Q���?AH>�O��=6ɞ m��� ւʪG��L���߇aT��h���4�����8X�OX̠���R)9�!�e�:�@'��O���OT���O1�ʓ�f�[��n�(`��Tn�I��@7X�J��G�'�~ӂ⟔��O,�DF�qF�m ��K~��r��+�$���sݴ����k������Uъ��|$+��U ���sHGE`!ϓ��d�O ���O����O��Ĵ|
2�O�/�vh�`Ȗ�dp�����;��vm��'�"����'�6=�x���V~�`G�
*O�!���O��D(��IA�eZ�7-v�d#�+E
lc��.�0t�"��7�h����DO!���%�D�<ͧ�?!wGV�V��D 7̓>m�L���
Ѝ�?���?�����-Pe���	��`�ņ�71Ԑ��ɜ�o���a�FF��4m��ן��?��i�������z�.<�f%\~��ͨ5�vH�U�
/D�O�r\�I.D6��)Z�*
h5�fJ�Q9fEI��'��'!��';�>���0��UJ�A� �`PT�M��$�I��M���ד�?��l-�&�4���G
�k� vÎ���j�5O$���O����u8�6�0?��ꃁg���
B�� �Gg� =�^HB�bL�2jD�$�D�����'V�'$��'�d )����\���˥-ڛ1"ƀ�]��K�4[+@�1���?����'�?i�H�o|���� �RT���\	K���ԟ�?�|g��\��'��%
�a�H����$A�����O�9�ZXc��CF�OVʓZ8�p����B���3�Ľ,�"���?����?)��|b-O�5nZ gH����8������(�27��]kD�Nܟd�ܴ��'B$듥?����?хǀ A�<��6�����R�ߐ�^�hݴ���K�^C\��O��O�g��"$��1��!h7�I*���y��'��'���'�b�)˪nw��pm�|���
g�I5���O���I�Y��f>��	��M+J>Q�G6p�(U�6
�&$�ڑ�E���?���|bF`�,�M�O�鑄��5f6(�4'T�B�Q��j����Y;��Ns@�O���|����?��K�����kV6|�m�5-	)j<t3���?y.O�hm��;��!������W���ķ>���jK�"4��it��*����V}r�'�b�|ʟ:�J��x���5R/v!�b���>�,l�O�U+�i>i�b�'�VD&�,&��+Y�I�u�A"`��h�V���	ß���ܟb>��'��7�)��#� E�^�H7��!$2�U��N�O0���ΦY�?!�S� �	z��8�G[	$�8���]a�a�'����i���/M�]��O\JH�'���Pr�
[��e]N~�ٞ'!�	ԟ�I����	�|��C����=O�0���nH�*�������h6mڀh���D�O$��3���O
nz�Q�e�����d�F=�~�K�Kݟ��	q�)��?
�o��<	T�E�(�^����
[�u���<�2�]�w����b�	{y��'�R`���i T�Z����D2�'B�'��	)�MC��F�?Y���?!�	V��a@A*�z4X����'�V��?a��S���p� �q�^����$ 4�B�ѕ�� ����R���"�"��!9��%����a׀�i`�j�<�D�O�$�O���?ڧ�?9���5�|���nj%���2�?�R�i����'��Ӹ���
��ɷ�<u��իG��������I���A��\�A�'��x�JEG� ����#�dK�ȅ$Ҁz�05H��9��<�'�?����?	��?飆�"�yy��R)Iּ#�h��������)a����	ҟ�&?�ɔN��	!�e�3�2����P&S�� �O����O:�O1�t�"���86ĺ|P$�͇w�$&'�09N �3Ó�H"IN>awW�Iy"O�	,|��L�Nf~1���W+)�"�'���'��O剛�M�!���?	cB:=�԰�$w:7M׮�y"�g�*���O����O��U�& � 	]pd�{���>`6�����d���4��5��(�AJ~Z��D�������u&<9DW�q2�̓�?����?!���?�����Od>���H�,���0emÐg�H��'��'�V6m�790�I�O"aoZx�	,/�Uyq��y8u#��Y�Q4b�t�IRyr@�2ms�F���2��-l���K��k�r�#$DqO����'j,�%���'x��'|��'�*�a��=�z)S�k_��-"��'s�Y�l��4?٠и��?�����IX4of�b'�3ZbT���A=5(�Ʌ����O��$&��?MjЉ�,3<�����n|`U@�@B��h}��U�Z���������4�Ҝ|R[>P��pM�ud�pѷ"���r�'���'���R��CߴjW�0 )�	
	�퀕�V0^�h���F��?��P؛��dWv}�'���g�� !Iʉ,[�tZ��'^�O](:��攟|yaƴ@Kq�ҝtJ,?� ���
 >�4��3O���?���?���?������10lL�R�;�����X4��o�Oh��ܟ(��[��ܟpY����2��f-�穟~�%�2���?i����Şb*�4�yro܈*����O�v�@�d����y2��9���I@��';������//��*���+Ҙ��E͚�4F��	��t��ȟt�'ê6-�O�B�$�O���ـ"����w�)Q&K���'I�㟰�OD��O6�OJ� ���=
{����\N`��[g���Q�'�;�o�w̧r:�	ɟК�ǐ�U���@��i�B���J��� �	ٟ����F�t�'�d�S��w�*,f�A�xb�	�4�'�6m˥G�*�d�O��n�F�Ӽ��@OvБ!�.Q���+@j�<��?Q�[�����4��dճ`�����nh�L*!ꈵ ���P�S>��'�*��<ͧ�?9��?���?�Q�Խw�(I`Jӊx�� 3Ơ��ć妅i�C�ٟ�����$?��I1r�]�ԩ̑F�2�`�D�=(T�x+�ON��O��O1���	�S}*�z@8r���R�K_̹aU���5��&p�b�E��gy�c�h����EK�	��a�F?t"�'gr�'Q�O��	0�MK�	W�?���;v��ab�m�ڢĄ��?Q��i?�Ob��'���'�R��XZ9���-2z(@"��:����V�i��	�v���D�O�q�h�N^I�lTbF7o���������OZ��O����OT��%��3W�Ҽ�gIF0fZd�x�fKF�0�	��4����M���|J�m͛v�|��̫7�J3dT�h�NݸR	�,z-�'R��D�#�����0��*6�����z���8��I9���2�'��%������'0��'�����"$�<;%�ܞ��2b�'�Q��[�4>t�{��?�����	��Z�@��E�2��@�;1�I�����O��d.��?����P0�<�!Gn��i{��è/�
�1F�z4����$�������|���.�]�O��m���òʟ9/r�'�"�'���D\����4n�V��U�L���� �P2�#��?��iz�Op!�'�&JOb�{rHP�i(0p�Ą��'��Y��i6�i�}z2	��?)pFP�(���*� 8D��mli���a���'3��'Y��'Sb�'��Ӭ1$`S!��;���`%V����4(ᢀ����?i�����?���y'��@vvȠgAF(S� �F�(�b�'ɧ�O�2L)��i���X�4Y�ুײ�؝[fi��T��db)[��`��Of��|��0����`�j#�Y��C��l1��z��?���?�/O��lڅ.�.������	�KL�L �c�5G��<�%fɠ#�$�?�dT�L���%���fh�)��M����&��@���$?��M
�CW�Š�4�O������?I @�d��\�'ʕ|�xX���=�?I���?���?I��I�Omq�g�y�	�@$��.���O0Ll`R�(���`��4���y'�ۀ6c��nR�K�fEK� �?�y2�'��'��Y#u�i��I�Y��ȧ�O	�H�����#)�te�#VD��s ��D�cy�O���'���',"�kH���$E{�%(�f4��I��M�T���?���?�L~���w-|X��)�(6�T�5��j�����R����͟@'�b>�B��]�9�tkB�P{�\4Y�
��]0�6?y&*�\^�$G-����fq41�&ĴH7�9�b���O���O�4�����jO� D�q���3#�� k�B��R��|� ⟄*�O��$�O���v������v+����AE�8���3�e�J�y����C��<u�N~j��U�>PA�'T�	HA8QJ��gj�L̓�?���?I��?y���O�����H��\�t��-KcTP��'���'��7m��|���O��m`�	�O>��9�OXoJu��fL�n�h�&���I���Ӽ3|�l�]~�듛� .��1+�"-G�ā'hC�\Q"D��J���?�r�+�d�<ͧ�?i���?�j�/�&Cri��v� ��"���?a����D����`fE�ӟ��I��T�OG�ɓ@�C�J�v�BAD)ÞU@�O���'cr�'@ɧ�	�( ��l ����!�dik�Np�!I[�P����@��(���0�|��@1%�!8�ϕie��h�_��'���'p��S���4U�����IT������Ůnpd�@[����Ʀq�?�Q��	��E擱N�2�
�@�)�*L�S �O:�d΍>��6M+?��c��2��,���m�ޅ�%f\56���jR�%�����O$�d�O���O��$�|�dݒ>�T�c�LuuxIڤ��Bp�փ�~i��'�2����'�v��wt"W	O#�(����E�Td9��'���|���A\v���7O�	؂`S�W=
�SO��nwZq�&7O4z�CB��~B�|Q���	�9���	G�p@{��@|�HI��Οp�	����Ay��w��Y9�<���:��Gg��;j�xC�_pm^����>�����'�lT �.�=/(���0��&����ORh��!7gU�0��6�鉷�?1���O��Y�#��'
��P��@%]0$��+�O����Ov���OУ}��V��"S*�9�V��|n"�
��3�F�����'� 6,�iޅS�C��٦��Wn:q�Ԙ;�mg���I��Ɍ5���n�f~Zw���+��O3��F��~V씛��	��|IG�R�By��'��'*��'jBi�=���u�|C�1���e��	 �M�WF�7�?����?�M~�t��B����֢�#�%�7_�$�	ϟt$�b>��(_7��Q#ǗQ~�	
��27�0Mn����dP�U�����'��'���'M"�X��ސ7�z����ݓP e��ɟ������i>A�'��7��6��"QqL8r�c�|!�mI=~�N�����?YP����⟔�ɖ.hz�h ':�̨%㘘�9B5hݦ��'`�-����?��Ɠ���w(iJ� U�i{j���$[z�h�'B�'4B�'G�'4�I���#]��y��ض=�$A�F�O��d�O��o� iQ��S�����4��'N�Uib'K'yUtp�$�֡B�\-9J>����?ͧ#�:��4��ĉ�iU�y���5)�m�s��9B��q����?	��;�D�<ͧ�?����?!Gƌ+a�2���	��	�9{�
�?�����S�AѰ�䟔�	Ɵ��O����@
1�����+2�(�Oz9�'[��'ɧ�	�.��
V��x0��I��R0��BKo�7� ?�'fY*�IA�	�L�qy��ʉW-�MJ�돌 ��1��؟�I�0�)�ly��b�(���H�a7* RAɊvݜX�K�	;�����O��lZQ�"+����X!����@J��si�1 �ȓៈ��+	�T@lZL~.A�!R8���X����@�|D�"�%�(DqP�Ŋ+3��<����?����?!��?!+��i�r�/t��(�gF޼$u2Q�"��ꦱ�I[ZyR�'��O�"�r��ˬr����0c�c��s�  x�D�O�O1�.�� kj����	"z�q�W#��c�h��{_��I�xu2��q�O��O���?����fABU�E#
z��˦�ߊ�~����?9���?9(O�l�@��%�������HK�D����(���0�CM�t�?�Y�D��a��xJ��˲��8��z��D�^��'5p�9��݆ow,�����Tȝǟ���'~.�tcY6 �RU�w�uC
�'���`%���l��MHv��2Ydʌxq�'|
7��2�D���O ImZ]�ӼA.�D��o��0���<)���?��%�����4����*ꥣ�On�	.��0ͱSɩp�h�v�|U��D҅Ҩ/?�� �ƣ{���� F�,���Z��	 ���ٟx��̟��J7hYM``���&Z]~�8�BP/y��I֟��	x�)�ӝHH��ڴ
�	8�|�; m�-����U�M����'Jf�Y��⟬r�|�S���F�@�%��x �čNF��:'G.�O
�n� ���ɸ$Z0��F�N�[X��C���*����ɹ�M���>9���?�������PbI	#�X�v`����V��M��Oށ5����'=���ﺰ:g��"}��e�TN��B	��2>O����"Q���RW^#B��أ1`_12�d�O��d��MS&ZǸiB�'��k�`��M�����C�	,)KҐ|��'i�OBN��V�i!���*����KI�!2�Bř_�D����[��$.���<���k<9����Z3`L+���O��n%(���Iʟ���Y��&�j�=�4�Nx&݀�����[J}��')��|ʟ�$�R�^�* �ⱇ�8y:-ifbH�	U&izQ!{�����4h�J?iK>��k\� ��h����ׄ�CPD<y��i\v),�0���=�l;Į�T��`Y!�'�Ok��㟨۪O����O` �ĉї5�Ή�BǛ�w�X�D�O&�zU�w��Ӻs�	S��Bǲ<� �+:hε�FGQ.J�LC�K�<�+O*�D�O���O����Or�';�Ef��!a$���K�<x̩��i��l1d�'{2�'��`lz�E�����	n-#�`$LV��O쟘�?�|j��&�M��� �t�$L�'$aBI��mzJ��2�;O�|���?��D%�d�<Y��?)o�1$�5C�8����\��?I��?�����C���I֥�ן�	���r�	�]5Z�0�S�	���R���l�Z��	����?�D�+ J�A�f��k"i�Y~�&:iL5�A�O��O`H!��O�ҧ�3ev,��D�	̢�A%�<rTb�'d��'}���ߟ������%Ѣd�S(M�f�z1��ߟ��۴D����+O�hnZX�Ӽk�:	=6<#W�_���
b�Q�<����䖈]%`6"?��]�%��	:S�̵ۃ�ˍ8E���l�)Q xO>	-O���O��D�On���O�p1��H�\�ڶ�,<���q�<� �i�� ��'\��')�O_2�F�⌹S�8J�!)�GՃB��ꓒ?����$C7^>����%�o6�Hy��Ϛ[<�8f9F�I�?]n�h#�'�q%�ؔ'��1ЩǣXwf��ʻKp+W�'�"�'WR��$[��)۴RB�C��G��x21 �\{��v����q������@}R�'���"�t
���)(��%�u(K+ӭt����U�'�LA�����?�i��$�w�˂Q`��z�N�0^*(Z�'I�'���')��'���"7m��#c��S��|:X�����O����O�m&��S���3ش��.��l`b-E�U� �a��BW�Hq�J>a��?ͧ;��Z�4����'n)'�T�J��H�=[�ap�NԒ�?���.�d�<ͧ�?)��?�gh�5�2@K�Ꮯ^���C��?�������˦R��Hϟ`�I�H�O^�3�K\� �p|8a]��P�O���'�B�'�ɧ����TH@���U��)��o]lڜI
Be�2f �u�ѕ��#e�R��c�	2�,\�0�S�4(��f-e��m������ן�)�S[y��j�r�J��9>l�.*�	!E�2� ��'���xӪ⟘8�OR�[�Kv�h�v���v�"t�bɌ�q0�d�O���ln���8]�` ����O�����ݰW=<��T��<>_H���'��	џ8�����I��T��X�D(2[
�\�T���Q<H��Æ ��7M�I�����Ox�D0�ӊ�M�;U��l��B�ѣrM�W�XX1��?iL>�|��n���Ms�'�b���	�l�d��#3�Ш�'<� ��l��2�|�\���3RJ/���a$�Qˎ"������������oy��mӜ� ��Or���O�z��V?�P�XP��/��Д/?��;����O���'�J��\:�HVK��;$�ɔb��I���t�p�Ɗ)��b>]�0�'��D��/m��A��)Ih�jpâ	!��Iӟ�	�`��`�O�R+�$_.�9� [;�케#eE04�"�d�0iI���O���Ц��?ͻb�,��v̐�\��Q�R������?����?��.��M��O�Tƥ����Fφ"����ŋҁl�x=����2^��Ot��|j��?��?��4�6��¥�3.��4���#8�|b)O�$n�y��IʟD�IU�S˟�JG�ƺEN�d�u��7:��l!Am/��$�O>�$+��S>p���o�U�����O� DH�"�k�,�'Ki!�aBW?N>�(OdmA�D� i� J!�X=bhF�A���'��'��O;�	��M#�j���?a��[^����`ơ1V�D`�Q��?Y�i��O`��'#��'HLw��UɗH	
<rap�T�]��qչi���R�jPџ�����
�l�pl����K� ���!�i4�$�O����O�d�OF�$ ���M�n ��W?>A�#)�=�d\�I����	9�M�n�����ߦ�'���S��)25��4Z{�4A'`�	Dz�Ot�d�O�	�T,J7m0?�%�Ρx���!��25d�DCԃI��g/���%���'v�'�r�'����f�d�E�f'�.xp�t���'R��۴x�U����?����	�3d3�� �hi��T�� ���O���'E��'Nɧ�i�0���r1�S�v�*}3�K��3n��	aj��R��7�Mwy�OI�������I�I⪼i"�����q���?���?��S�'��D����c�Gل!�q���T�hdᬌ�L�t�	�<Aݴ�䓅?�Z�x�ɆK�$)1��] '�0ط�%i��l�	ҟ�3u
�٦��'I̤i �H�.O�(#��N�{"�S��&p��(�=O���?!��?���?����)^ �cR,�/<(sF�]�(ҌlZ9:����ş���}���<�����\q��V"� 8~��v�֭�?����Ş}G���ݴ�y"'�%/���}�f\�S��O��ñL2���'��'A��@�I3j���Ӡ���8�w�*y7r �����ɟ��'�T6��2BFʓ�?ѳe�d�؍p�F��H�@�3�������?Q�\�����`&�Y֡É46��SW)֍s#��	��7?���Y��j�
���d�D��?�@jO2t�1�f�I2����?	��?I��?ي�9�M!�JE
Ok��A�*��h�A��O<dlZ�$n�,��۟4�ڴ���|λ@ŌH��IV�7�q	T�ߩ8�m̓�?y���?�Bņ�MS�O�ԩ:����4?M� �0B\�?
݃��W)=
ȹI>�)Ol���O����Ox���O���N�@j���/�l����<ab�i�*����'��'}�OrEY��p� %wƔ@EG\R��?1���ŞK���� �x��('g���f@�	��$3�`a�B��'JL���P?	K>�+O�䚇��"o$�2��M\����e�O����O���O�<��i8��R�'2tYd��&C�����!5I<��rB0Oh6?���Ot��'~��'�@�[����PΓ>6
��ɣ���"�t=�F�i���>
.�d��՟Z����C�"���"�&]�<�2fC�b��O��$�O~�d�O��$$�S���9𥊘�cZ�� �	�)t�^�'{R~�<���2�
�D��Y$� �2��*8�bh��l	�@sz�a �B�	ßh�i>���I����u���m�&�#�S
uP��bV
ȶp��1���'�0�%�(�'a��'��'3tMRǮ�Y\�Q��-Լm*���B�'��P�tX�4~!ʭ��?����	�4R�yv%D-w�.��N�TB����D�O��d5��?�:����
_�Q��.O�Budz�c�#��8HC�X٦j+O��~B�|��A�JA��L�6� �"$�G<F��'\r�'���d\����4��hV C�&HŲa�ˠ�Z$bO	�?q�����D�A}�'P�ma�C�G���T�ɺBYF�C�'8�ȒB�֗����9F,�)�<!v�H>3�te���Q�[�=�T)�<+Ol�D�O8�D�O����O��'م��&��˳�U�m�.\5k[�B�6�ׄ}|��'������'�d7=�n3a_�#$��Cd��L=)�'��Op��?��T%cW�7Ms�dq-R
G�phj�lEWjX���k��p�"v���#�ı<���?�)�ZSl��SF]�K7,M��d��?����?������ئ}�ǉD�����şC΀/2���h�8�|#�A�nE��Ο��IX��8���!/�\�g�p�E����!�u�1o���'9����Ɵ�����H<�)s�D?	�L��i������ʟ��	֟�G���'fdL3�jv `EЊ�Ʈe���'��7̊sP���O��l�g�Ӽ�u��!vZU?,Hp��L��<���?��!���޴��d<��<3�O^�x����`A��A�_�� jt�|�Q�X�������՟�Iן���C�=��}�g�SsE8p�Lwy��x��)B���O����O0�������J<��e�/9��(�4b|��'k�'�ɧ�O��	Gd��5��h�N%o7�̈"	U2VЛ�Oj��J��?�7�7�Ī<��H��v�p��l�3^��i
q�߼�?����?���?�'�������'Iܟ+,5>V4�2�M�]���Pȑ��۴��'����?���?1�/�j�bF(ϵ-D~(2�`G�0A���4���P�5y$���'�O���e�E	1,؃5�� Z6�8�A���jb����8R����$��h����@%v8C���.FИ�����2҄1��:4M��dG��F���Y�^�',�ݣ�e��VE`��5I�#���9���4(zb<�<9��]4*B@y��#C�P�Bϰ)D)I⅗�K5vm���O��{��>j�ە��-{f8d@ʺ=8��`���gi��[����Ӂ�HG���ʆ:b�	� ۓ,1 � 5GA�ּ2��&"�miR��\oL ���M�����D8:-��q�O�@~�������y������	8~Z`��O�˓�?��'�65K�DՊD�J�x�nX�.*�i��4��`���B����'"R�'��D�1���-ڲ�&�G�������v���Də!�T��'{���$$�֘�W�T\�6J��UԠ�׊A>r z�u�<�������O��D�O��l���X� �|�a�I��� �V��!��Iy�'`�'�'��qzu$�U�(��a�:+�6�B4G$�'���'
BX�D+!+Ѧ��$A�U�QlM�]�F���NV�M�)OP��;���OR���H���ɹ|S�� �A� hb��W�Q �Z��?Q��?�.Op	�l���'R�����%�Aw��(Z�5�De�r��:���Op�$�O���$6}����1l�D�U��K�L������M{���?)OmZ��X�t�'f�џ���V�W�����	��\	�s�x��'(���B��O��ӊ�8T�U.�~��}K�),n�Z7��<����(����'�B�' �s��08����ڮ�0�۲� @7M�O<�ă!w
�H�}�e�:!�hr���$r�ʭRd�@�!�v���M����?9��R�Y���'��<R��"c�-�$�*cxӲpҕB,�Ij���?Q�E=LX\���(ۅ{��}B�p��v�'b�'�T٨��>�(O��d����p�N�D����&�-D����p��O&YJ��a�ȟ��	ΟX�����H]`eL�8�Xe�䇐��M���C��Y1S�L�'��|Zc��52��W�R�����B�nM#�O&�rn$���Ot���O�ʓBȴ(��Bci�P�ۊ;di��ί\�mhI<����?�H>�.O�־[�2�ؠ��Koz�І��x}���'6�	������ܔ'�,����o>Ɏ�p�hS��b"2iЕL�>����?	I>�(O���Oz�!�6h�J*[&�mK�H�S}B�'���'��I�V�Be�H|
�M׀���Q�G:���A��?���'��'�i>a��X�i]>~N���'<= 4�sa	���'U�W�`�u
����'�?����H�?I]���1���K �U~�oy��'�R����u7@I��� !�̕NX���#����$�O$2�E�Oh�d�O���꟦�Ӻ{s�^�6ɩ�n�$0C쌡ԮX��fy����O�O�b$�M��]y��J�.�^�:ݴL�����?���?	����?b� ��R=����IZ!�dq�X�|�O;�S�'�?����#��� gΎs�v1���ӽR}�f�'�r�'{
@���/�4�v�ĩ��YA@�M�v��3���䱱Є`�^��:�$A��O��d��t��(S�1vPؒ@Z0y��ź�'a� �$�%Z�2	�J�G�h�B��f��4�2��>����x�Ç��D�O�D�O�ʓ%Z�u��
	`�t���ހ��|��g'5h�'R�'i�'�i�թ�/̛oAd)�L33�HY"��bӬ�D�<Q��?a�����m��Q̧"��{�C"O���T��BU֬�'�r�'w�'��i>�ɺw��`�`n�g2�pe�2�$mi�O$�D�O��D�<��l �O�<tyEJ��L_F<�3�
M�g�p����+��<ͧ�?L?y2F�K�	�v�
`�F���y���D�OLʓua�K����'��\c9�P�g!�'N�LR���L�b�M<�,O��D�Od����0�@*=jtJ��E6,{vd�@�i��	8"`�Y��4,D��ޟ��������0l� q��ޢdyR�a�I~'��]�(�	��\;I|RN~n�Ao���*��xH����
�$6��'Q����O����O^��<�On�i�"�t ��G,��v�$Q�@ʿ>���@B���8$sai�;(
d0� Q��� #������	ʟD���j�����.}"�D�Q�0Ɇ�M�2�ˑݾ#<	����'�"�'Fi0�c�|d$
��ѳ{��	1�}�x�d�b�J4&���Ɵ�$��]��D�6E�\&��'�T< �O�$!���O�ʓ�?�u+�v�|Q�&
]��U �� �Y.�h/O@�$�O�⟠��^?y���<��P�.�F=r� ���M�e+?	���?)����dU��ϧ?x��s���L�����HC���'�R�'�'��i>��	�w/�XI�MF m�C,Q�=�<���O~���O>���<��*�c�OT�� a�_xDQ��G,�l�b��d/�$�<ͧ�?	M?)��h��sE��^iBI�Y>�V�'�RT�t!dD��ħ�?����\iR�����򲙪`��E��]yB�'�����u�Z.b��@���B-��	ej���$�O�<G�O��d�O���៖�Ӻ�S#�x�&qЇC�Io�T��,\�����dy�J͐�O�O<�p�}�d�Jak�2=�h�Qܴ.t�<���i�2�'jR�OG�����6Qk���X$��<��O�~�n��N2��۟��'�����<"��ࣃN�tW����c�  9(�nݟ������h�;����<���~rÛ.1ӎ-��%�-s�B���D(��D�<7��O~�O�"�'���i��۔�D 0XD��_����lZ���s�&5����<������Ok�Χc90���E'�~�XbH�&O���sf��Ry��'������R����رB�i�x�Ħ�*
|�-᡽>i/O:���<a���?��b�d<,J#��S�B[ ���%f�
��Οp�I��t�	���'c��F�y>����[�`^�hJCgT%8��b�u��˓�?I/O����O(�$I9]q�d7oX�sǪ��2��F�B$1�)�>y���?������ ��l�O�rG�9�� �%J2�N]xW� ?��6m�O���?���?�� �K�禁��NC�Z���'��_tܙʔ rӰ���O��D>tP1�Q?m�Iݟ@��?jB:���	qI�ebC�E�v��(��OL��O��֤?��$�O4˓��D�̄k�@|�qC_�\�Ba�Sa�&�M�(OxX�ʘަ���Ɵx�	�?�ȫO��C3�^|9Ĩ�<����G@L#3Ǜv�'�r���yR�~���O��l��$]WH�Vh�(e�:(�ڴ0*"�;ֺi|��'��O?\���܄e�`9��H"M�V-��g�Zmlm��@��Ij��T�'�?a��Q�l�t�If含���1��a��F�'���'�8��c�>I.O���Բ�+t/�$�o��\YQ'�>i)O�ԐF������ҟ�J�$��!�^��D@��s�@�M��Os.�C5X���'��[���i������Oju��ƈ 2��
���> l��<A���?I��?�����Ѵo�B�!G!/>P���ñɀ�*+�o}rQ����Ryb�'�'���"�1�n0���ц0�x]+WW��yb�'K��'�'��Ɋ	��5۝O����HZ-��Z�)�&L���4���O˓�?)��?ɰeS�<1u:@0��hPL5Q� �AVh��	���'42�'�"Q��R����I�Okl0	���R��X�z�h��Һis�T�0��ԟ��I-Hz~��B�ܴ�\;r�צswy
֫�e]f�lȟ��ay�@�p���?!����p-�-��p�',�h� ���Mʑ)�	��@�I՟P"fGr��O�П���e`T�SC(�z @!F���k��i�剣W�
9y޴�?���?��'[��i����Υ5�*��5ɽC%���gM|�"�D�O�@P���L�'�q��,���i�.h�"!F�'Y`iє�i:����p�����O6�D����'O�� x;b
�/���!���B�=ڴ@�H�'��Ip���?QwDB0� p�Dt
d!B�QE]�6�'e��'�:\�!ǫ>q+O��$��h�#GZ��T�*�<p�n���b|��O��6O��$�Iş֭̑�)|����G��?%o(XBFډ�M3�ZW�p3�T���'�RQ���i�� 0�9��Q n�	�#I�HU�9�ǲi�bA�)�y��'���':��'��ɏO��M"��ʥgHα� ��K�|��Ѭؚ����<�����OF���O&aj��'�ݠQ���7�&�Z�چc���O�D�O��D�O�˓� �1��!Q�oݵMt�A�@�B>�Tq`��i"�	ޟ4�'#��'yB��y��kO��;A,-Ɖ���U�6�R6��O����O���<�7�ϖr��OI� ��!�<yR�d���v�V���-p���d(�D�O���ȃl��7}�	m�6x�e��
1ޖ�1�K��M��?Q)O����Yv�ܟ ��m*"��5S����d�p(H%8K<y��?���Ք�?�N>A�O�DзjNt�@+3av�<R�4���|@�o�(��	�O����p~"��0t���"@-2�۳F���M��?�t�?�H>I����Ǡ�DQE�	8x$ma��
�M�UG	E��6�'Z��'��$G5�ɡ�����	#s�44��أI����ش8��@�����O}��8uS0�7�ι��+�6�@7��O�D�O����h��?��'�aȐDƋ �e*��7�LX�4��?�v�S���'.R�'2L���+n�z�ӶNő)CT)+� eӞ��ҷV�&��>�����3C��l��h�E��"��q��XI}R�ԕ��'(r�'��^�t�B�v)Xy⳯��|�DY�#�.c��zO<���?M>����?���Ր\����/�'4�I�!N�,�L1�<����?�������`beϧ8zy ����j$��z%���'q��'��'p��'�
��'�<-��!��G^��$�ԲX��3�˩>���?�����͎g�T�&>a�a#�%��hѦ	>��-��[��MK�����?A�N��������ID�^<���͚U;�B�,L#h�6��O
�D�<��OH�",�O���O�^��E�Y�"�D�����R�:G�'��O���9��7���?�@���
Ӳ������Ր�	y��ʓZ��(�i���'�?i��^��Ƀe�(M���Y�&�6�`��λGjZ7M�O�d��(\�d-��2�&g^��Q��Π�$����X��7����m�ៀ�	����Ӈ��'Y��T9e�B� &�'&�΄av���-�`>O�O��?���
P���2蕵5z�ᩓICy��p �4�?���?�$��r�'yB�'��dW�W��)ѦO.^Y$� Ŏ�����|��J��v���O@�ĕ�tE��pc���l�ɐl�eجXmӟ�q3��3��'�|Zctx$UM���D�:���	i̼��O�Rg3ON��?!�����ORѨ�A�W�-ʀNU����N��q ��?9���?�H>1��~���?LZD���͕_���tS��Mp�Tw~��'B�''�	J�25R�OѶ-�@�ݴ��P���ZHz�O����O>�d2���Y�8�'l.С�!�*��	�I�r��'���'_��'�+�(b��'��2 X��K�TC��a�� �6-�OB�O��<��*�w��)ԴU١L�vTc���	� 7�O����<��h�ىO���OĴ�!I�/ඌap �:K'�r�1���OL�D ���'w4��!l�]F�`�s��i�t�n�ty�� {�~7�k�$�'C�d�7?Y�N�� :
��F��&4,-*6m�O�dŸ'�x�}r��=XҴ�`U�X>9�4y�/�ŦU[�k�M����?���bw�x�'\����ۨ���(8�z����b�z�E�)§�?�c�A�1p!�RщC�|�0���7���'Zb�'�8��q�5�����u�Vm��N�H4��[�n9J�}�>Q� Lz��?q��?Q��Q���xBB��}�@� 
�)���'�v�[��/�D�O��d=��ƶ��"�>|��k��̔!��{$U���AK4�	şp�IޟX�'�z���ɷ+����&�� �B�<N��O�$�O`�O��O}�������8S���*Ҽ�c��1O>�$�O@���O����C�:�����F�3P�0z��]�4@_�Fy�m�ɟt��矨'�p��gy�+��M{���8v���cхĥ�T�!��L}B�'sr�'V�ɪz�0�L|B'�φF�^�ɦ�̟s{��3	,2қ��'�b�$��05����p�'έ�Bq�`B�;��t�i��'��'������'R�'/��O�������%`y"��s��ZCŋ!���O.˓`	��DxZw(���V�79e��i�_�W�]��4��ĖD�~�lZ>����O����M~g<
� �����x��%S��M����?�a��e�'�q��p�E燛G٢�yUaOr�rd��i��xC{� ���O&���e�>�GGM8'����+�D(���kQ�yi�f����O��?��IŦ�*BE��x�6Q��vOLaH��ij�'aR ��1�O����OB��(Xԍ��-�V,rE��v��c���$�3�	������dQ^���a��T
�$��b�/��$WR;��nyr�'+�'��� %����Dr�T,����;�D�y��I۟��I��P�'����\.
x��P$ȘD�,�c��1��O6���O��$/�Ɉw��@�0P��1���M0!q�Y9��<�	��(��Ο�I󟄺v�՟�P'�(ڀ!&k�44g�%ࡃ�M{��?����䓱?�-O�Pd�� tL*�l��V=2dD�*<��a^���I�@�'�R��L���̟0r�AZ�C���"��>g(!! ���Mc�����?i-O´�x��ҳ"o4T�1ҵ8Cbe!��,�Mc��?�.OtA�Q�Sן��ӷ"�ڬb���K\���r�V�(���K<���?Q6��D�'��郠D��9���Y9z@l,����2��X���C���M�#P?��I�?�!?1�n��R�
�h�]Z��T��i������pm;��O�z�����(v�T�$�T�
�K�4D :���?9��y����d�|JW�X"Cx����I�&1(1(WD��j��	 (�D#<�|R��\x`V�+��T�0LC�
B\�Xsa�����؟x���L,��N<�'�?��{�FRT̗5'��%��^�4o2��C��� }�1O ���OX�dQ�B��91.��/���1ց���p|m��<����Ry��~����,y��SÁp\|��
�uhFpyC�x���#����OD�$�O��*�=Z�a^/��`�D�O(�rɞ�	�O~� �$�O|�D� vx�B⧈���1b�dr6%@��O����O��4M�͙�8���� ��<'0)KTl��`Y"��CW���	��D'���I��|ѱ��>!u	�Ae�� ����1�n|j%�X}�'��'���'�J�J��'6��'z�����	J��wȴ�7�-8K���'��'q�]�D�Q
)�D��?����3��z�Xi�Ǔ>td�f�',R_�� 6`ߥ��I�O���ꟾ@� �M`�xܪ�D�
��5��Ȗ�?���>AK;Oxdu��A'��@b`�æ���쟐��KRş���ߟ���?��5v/��7�����cN�>p�a ��M��M{������p���x�u���I:��"l��:��')B��g�:ga|��,� a�tK@8J��դȤ�y��<Z��œ`�02Æ�ʤ  ��Μ5�];nY�s�ݠZ&h��al�6N��eӀb�>.��]
%�ڞ<C$���˕���e�V$�W�vIѠ L�R�"ֈ>q��)sB��CnLؠR,R�
0X�N\�<;���GF�H��{B`�Ud���4�ԗ2�Iv��)�6���ܟ ��ܟ�{^wz"�'h�)�}��z�ُf+����I-��r���GNV} �$\5mZ@�C��v�'�B�˂G�((��Dr ���q4�U�/{�a�	�7n�Ё#G>A��U�q�/���ѣ��>$�g&>DP�M8SĚԟP��t�'��O8���ȕY1t��ƯN,��|"O��"*!hk �0,�-Vl^x���Ҧ��	fy�%ψT���?qPn�w��I� C J
8Y�I�2�?���$��*���?��O��- �-P�uiJ�ρ(,��Q�)��Q4jV ����c�m8�@B7c�nI^d+��?߬�� ń��d-k�,Ȥ=�C�"�4��x��ٳ�?�������4;v��"R�#�֔�%'�<y�1O���䎌4���&`�&g���4 C���D{�O��7�ـ +��P�#Є��²����$�<��טB���O��]>��7O���(���ͻZ�����[2T��p�䍔Ɵ<��F V�:V��x����s�@8�?�O哬1��yO��Q���̕S��'m�lꗧ����������yc�Y�O_���Ԧ�E�0U���V	z�.$0L�|�6�O��-�'�?���D�?_�yy�ʹ�q� t�<!�� t'2L��OB
Y"� b�/�hO��v�'��a%fC�\*����K�;jZl��Oj���d�O��d�3	�&<��j�O���O�4��!!e*a�uadEH� �ɲ ���Oءëw1��'"������j���3c�	'!�
T0�Ā�w���'��H�f�A�g�	�;S�Y[r��6j�!5gG5��i�	y~B
��?�'�hOv�R���Ar�a@�Α.RHzu�U*O�iƥ�p���"N�R��q�O�-Fz�O*RY�P+2��NĎ5*U*���@-��E�9n?"U�4�㟌�	��l�jt���?I����	J?a��pdo�B ����]�i�� 1�nUW�����V�j��F�T�उ '�p�H�d81Ȑ��/ϗ~�a{����t�9��-�8@:�l�h�V]����?9�d�*�.\0u��gW(}:� �s��'�;���(�Jh@q��c6M��7��+�M�J>yw�ƵV���埘��M��9St� hXx�)#����I�x����h�'0�țCa�KĎ�#Ae-�M �	"��x�1jةF�l0�B
�e8��S�fʳW�ė�b>��"Ǧg�T�:񩛩W�����Y	r���'�X����?Y+O^���Iǡ*�DI�U�;%3d$�����OL��K�rE�
ϝ`�\�0v"�-~!�dV�����i?~��"����������'
HP��y��d�O�'M͒5`�}6X�B&μ`#8h����j�(���?�Ff��J:Zq��ƙODX����|�' �
I��#�i�j}�9d�E�$����@N@�<�DL���7F�|%�!�;��IY'L}�LZ��Y�i^��	W![�j��1׼x�	u�S��k ~�P+C�q`�P��Ә}_�L��S�? �E�����`g@ϩK�9�2��|�鉏'�RL�����my����/F�.�p޴�?����?9 �2�f�����?����?ͻ]:��ѤE��2���^8эy����<�4D�o���5���Du(vM�R�\�℆�	��<�O\�<X*� ��$vZ��<!@����>�O �S`NƃM�T9���)3�؀V"O,�Z%��=���i	]��9П�*��4���O ��B\�,�x�2I�b�:�	60-��U��O��OP�t���'��iғ'��\��B��
nL[MåXa���/"�O����,�6(F��s��f^��
u(�5{�h����6(��0�HS�F�9f�
S6�\�f�'"r�''�S����f��<-��C��Xέ'nA$:������:�Z�+̠$����w�t���<��P�̕'�T$�$q�l�d�Oj�"^�z���HJ'_Lr��4/�O���ۆc�����O���2Lbd�9��~�I2�l�5O��0��@�N�IV���Dܢ�c"[!$<��8��ȳoc��yq���;`�@�g[�H��ԨҀ!���@����8�۴�?yd8>�-Z�4)�V��������O��"|�B퇿j��u[W�H�B����i����	��M#s!��i� s�� j4,ٶ�F���	t�'Z)siI�q܆8��] �b�k�'a�ܢ�d��I}6qA�q5�I D���H�*�@�[Q&ܖx7�(�D$D���d@HpL:Eyt ��x�����7D��x1��[�
�3���O�x���!D��R *p��#�&�t,��a;D�`�Ѧ0=������#M��	�!�8D�(��V�f����d�׆VD�y�tN6D�����M�$��L�S�ֺ���yGF6D��ik�+�9+�J-��1�
5D���R�A1`���9��5Z�pIC��8D�`Rm�$(\� ̅� �l-�" 6D��"��G
W�R���,u:��u�2D�`w&/(�8rMĢs���&,D��[2$�'=�<���GĎ0���نI<D�L�B�!0N���RF��r�����9D�@��@��<�hū�HM���}��6D�h�b�U�<����X:�4D��KՃ5,Q�ڔJ��O����v�.D��:����da�M�B�<A�,9D��!�K�0u+���%��TJ���CN3D��5`��{6¥S�� O�"�1D�P�6��m�p�"&�[�p@�b�0D�4C��J�E����F�`�F.D�J� ɖF�<˱B؃h�Nࡤ�8D�{g��4Y°Z�+T�Q`�i7D�$ٰhT*T$*R(��p���*��3D��i�⎴_��4�Q�M"#����2D�Lۓl��)��������d	1D��X�H�Im�����H"�PPQ�/|O��ɤ�	]���	9R�9J�M�9�\��"	�}�B�3=�|P��N��[�B0��I7�\��a&�)cr����S�Wx��_��DK�*Rx~$C�I��>�JfH Kf�DY%�F�;@`� �L�xG��'2����1!�`r�D�KlV�y2c
&.��PlB�b�Ѐڔ� 7�?���C:
�6�i�
,lO�)`�^�4����KVB�Ȭ�'�ta��8$i�(mz�T�;������$�(i
l��ȓ-�V�i�_�,��Q9�kP&?���?�D���:S���S(�':q����8�s��A�T�ȓ;��pR!��/��(��M�5!6�'4(#=E�DN՘X�CKߘL��Ǎ��y���]��t��.̖MyZ���/���y��'D>�!d�%F��,9U�]��[�ڤ!��f��t�"AN'�\���S�? ���F"�;QT��"�ϑw-�X E"OHЂ��&Ht����%E��w"OȌs�F9|�8y� Ӡ p��"O�!�phǃc%lpA ���w ,��"On�5�҈X�؅d�uW����"Oƥ�U��Ҡ�$"C�.T6��"O��"������Cv��=҂"Oꤋ4@ڻ^L�B E+��'"OJu11��2��0��4���"O�(��L�;�pЊ2F�"V�N!	p"O|`#���`��A�eW�
Ԫ�"O���D` ~���Y��ґJ�Z�Z�"O� ��#V#d�R䊕��U�	�"OPt�4BR0_��)���F�$�e�6"O�0���̨�k�5xL��A"O�i
���m�H��3�^�K]ґ�G"O4�*c�˜�,lX��ДKP�9a"O|)�D�̣,J�,Y��>�B��c"O��y�L�1p+^�&ȓ�q��hs"Od�r��C5���suI�AtB�Z�'/Lx���V+J׸ ���1�`��'l��g��^�2e(D��/:��Xk�'�|L1�J�g�V�����eV��k�'Ӑ��c�+o֊(��:s��8K�'�DI�R�
$�P�F��e[(XQ�'t}P¥Ŝm��&�ɤ`\ ��'ў\�#�=-1$m�"ŀ�A�Y�'��hH�!\���.ޖB�`��'����o�f�J��VLӓ@�
�J�Tź�{bH��^��p�V�ǢgB�i��i,�y��t���C$�ޙ)���*dn���ē7[̳����\<d4��(P(69��Xsh؊�yBB\{꬈�rZ�B��0Ed�"�D����J� ��%]?7���L>�7�@m�����%6��`NE<�3�Y�Ex�YSB��Hm�I�7�8D�pK�E��Ћ�*�$CX�@�@�%�tx�y*�d����mȒ=��n�t|�d��'׾I �X�#����)� >r^��u�p�DH���uxl�psHӹ'�HA�K��mr��O��}��!����2������(I�7Z�b�$CI�8�$;�H ��!����"Bc��a��b|>�3Vb,t���[�H4�s>lO�e�`d�$l���(�h�ກ�0.G�l�Fl���B˦����j#�O&�����n+�ElڃP��1Y��<�djB��=&�<���O��D�Ѕ��+�� 5B�0
��@��6}�)�4A�84۰�%��m�K%FB>m�I>y���S�EȖg�<��	V�F+�)�@�	�1ʶ	��ԧg޼�IVd�!�H��hӓd̤Jf���)R����V� ��Q0G\�l%�$D��A�Uۓ.o��i�!2>��ϓ}i"p�F�F� ��� !�tTؕ"
'y��(]�'(+j�X���L,�p��q[�xCœ�;nr����s"�P��$E���h�'Κ5Zp:a-ʐhuXMS�ʭV�b�Z��~���U�	�nX�	��q��Ĩf�A ����ܱ��ЙOP�aa����8^$}��×*�����&Fͼ)��Iʧ��<YŨ�^k�8(pa�:=�$:��V�'�x�k�صa+��c��p��0�\<r�;5���6�}h$�^�qo!���))`1Xׇ����ܒ�M���	O����##�\�`�4)fk�#|b��K�^Ե��L�	� }+��v�<Q��L�b�(�FI7�<$��=E�J�(��J�m�b�S2Ȝ��}&� B#�Z��xH+�c��xI�u�$%#$���"f��P��y�1B*W�h��c��p�9���|�$�q3�6lO�R$h�>=^.l�F@�Z��D��'�6q!$�T6�"�c�'�.y���[� �$0'�ߡT�,L�'���F' Q��@�P�_"�X��}���(s֪2��	�ݖ��f0s�h9��C3m|d!+Pmm�����F�[
��aC�F1d�
����2<O�!��G3��Q8�|Ѣc]�`*� �i�;A�
��x1��J
#Z;����U�+;$T$���b�T�/3qOq���%��U�b��g"@r�P�"O� �K����P낆��2\�b`�@x�*Xp��L�d����i3j\ї�I#zȮ1�y2F�����z�ӁI�������~"�':P -��Z�����@!m����	�'��!2b�ݘ> 0��R��I	�'v)��NLVځb�"`^���'�DВpH�d$R��"�4SU���'�ra���O�<�f9���2P���1�'�vE�#��&XI���%S@�S mVV}r�K�+�>7�>��3�	�L�1CE��J�l�dC�����$1 "��Ff'O8B���CمL�$p!��*{dVQ�#�{��XI��<;/e�Bn#f#�(P�;�P�x��sbQ&*�&"��~"@EŜ��%GZ}�X�b�X�<9�h��>�|L�f*ї3���үX?dcK5W���!��ĕz���	D�x�����\~TP���'H!�$ EK��cG!P�t0D�8G�,OD`�R�?.�L<%>c�T�K4�aTLJ.\e����&D�h���
)s��[�E��Fn��ٲ�&,���R��'��y��GO���56����ۓ�0��F��4��� hK�E��^���7�!D������#iwN<su B�f_���!D�뢡Ǆgڔ�����S���g(+D���sKYd� ��c,)T���-D�6��4��D�?�*C��`�<Y��}`�I��B�LS�I�fDv�<Iԭ���㡇�/�f�⇁\w�<���<@L)�كz=.�3"&H[�<��G�2N8hK�j�X���iEc�<�`��.�u�f��yEJTCtFc�<�v��\�E�M�.�	q��?��"O���
T* ��b@[(iRh͠�"Op�AS�P-7�:�w��*H|�&"Ox��$dP�/��]���UO**�f"O����Z������G�g�Y�"O�d�����5��]aD��k�`��"O��R���X���(��ԏ	�̵�"O���Aƚ�V5jQIr�F�~����P�r���Zu���EƟ���Le^��a_=��|�kR<��d��Av2M�u�����3���"+��ȓO���� ��8J�`��teS���X�ȓ脱q� �&)]2]����5�V���3l���dEM�#S�
"ǋ�O輇ȓ/�4x�C�лs贼1�ȅ�Y����	�G�ށ�rƑ!�v�0��*	$��f�
�F�Td2�c��l�n��G#4�Բ��?"�⧇�ys�K�m;}��N��k�ڴ^���A��F&J�������o�PQ"�ЎH'�l��"O��0�,�)�J� T�VN���!,Kw�r!ز��F-,A e$���q�0O���f1^v��7׈!6����
Oj�@SFX2j�")��!N 5@�H
�H�lm��6,� J�$�ď�H���dʠ:�8�8p<=^�u�U�ˏ�ay��<|r�T�«�3�mYԇ\�x�J��2�Q�.ǂ��ơͻ?��u��'ptIC��SM0ŹѪ�w6R�"���Y�@Q�e�U��O�ᆌ��bn���w�	E���'D�:V�H�Y/�lB�c8��Ai��g��t�u��$ 2�ӧ������^&U`�&!��PۮX�-D�����`{b�3���2�Ȣ�<���-Hbz�ࢋ?,O�P��K	����A����' N��Յ�1f`��BK�C��� F�O(�9J�c'$��y&F�k��|��B�"�N��'�;D�,��D��_	fx;@�K%,�|�k.D��BA%U	hx�#C�?�l�k�A)D���e��P%�R��%
��b�9D����&(dh��à&��4ѕ6D�� 6d2�l�+}(�` NG|��"O�|�gL�	A�ZQjr$����r"O���!�2�M��F'	��"O
�)0b���&��v���E�\��D"Oti#�K�(h�8!��J��P#"Oƴ#����,����Q�xߘhsg"Oj� �W��y(�+�QAt�$D�`�"j
ɖ�d��7h��#�%!D�lI���
4;���[Z��a$D� D�Ù}��\ڃE�$��3�"D�P��H5[�\a�`7'"� �G?D��$��z�p�ń�,��Y9�"<D�(��Ó&ӂU��,²&��Qu.9D��8��D��ѷ �:�t��2
=D��dl��� �7oQ4F�B�'�/D�p3PLK3W<�A�aHt�2`3��-D��J�'�=�>09S�!X�Ѱ�.D�H!#4_�2	�%#����#�>D�Is�
a���2��O-X���c*D�|�ge�	���Qk�f�~��u$)D�L���K�>�b�\:Zٜ�@�%D�ģ�j L�Z�b0�I
R�.D��#�� -`Hl�3L�_d��J�1D���`��#K2�{1dH�m2����-D�(��OT%���'Z�]�H�E�+D�<z��_�0��Lb��ؙV��[�/D����g�G8>Q�&E��i�E-8D�H#d֦��<� �f�$�6�!�$2s�~�j�c��R�x+VJ�>{A!�DT�N	d��&p|�aR��1��'mbY��_�'Äd�����'rΙ�$�D�(l�,>{���8�'���:#�
%"5NE����(y=�@�
�'|��Q��Ɍx���(U�n��	��'�d����68�T4�VG�q��!�'�8��U��F��!��^�:x�q��'�H�K6��$T��tm�4Z
���'�I��@[���P���-�ޕ��'� C$�6a||�����>d��U��'��m[5�)�QCEB.�n�J�'�r<7"^1N�Q�7�2�0��'�P���	Ĉ����ݕT�,��'��`E� WPt���O^r��
�'�y�Êê:gd�3q�_7�0��'���	TfM��e{��F)����'j��C��:���8 Z��b"�'Uu�bhR�=�j�3��E�=�D�8�'d��Rb�7k�1cg�c��9��'t�2�<E_��7�Ҏ-U��A�'�=i� RnQW�V�1d" *�'z&�G��h�����"@5�	�'#�|@��C?k����6&�ɱ�'��K�װ.�U�r�H�<�8(+�'��I��3i`&����!0�y�'.5 "IԜ/M2�F���c(e��'1�u:G%D)U�@`�@Q?N&Ac�'��P����K��BM�S���'��TY��=�d��'��O��\��'�����L<<�p���8D�`�2�'�
m�)S@K��Ý(9>���'�1�a@���� v�I꤂�'�5�$��)�$4���˘q���3�'&ڌSa�-uEd9YWHW
ʊT��'&P���I^ WGbY�C�O� KJuR��� ��y5��Ue�\hB�Z�JJ�`�"O�Pj�@�����W�m�x��%"Od�つ�o�6�{��5��T
""O"��"�C�&K�pʢ�2�l;�"O�-�E`Cn,M�S�M�k�=:�"Ol�zQ ��!-�E	�A�3E+�h�W"O|d��CZ�/E�9s1��5()��"O*}�*P�2�2E�M�W�xM��"O~��A�1R�^tȀ
�m�PeX�"O�U	��Շ��XQ�K�&����s"On�p �� j[���A�-�(�"Ol���Js�I#��y��堔"O&�a��>��[ ��7d7D�d��m���V�Q�R�q��1�u�4D�@x�׃	K��Ӑ`�Ur�i��+2D��S(��q� s��=k�cr=D��!��V&���'��"J�d��:D�@jîB��#�)Ғ\��=Rp3D�<R��I)g2P�4�-J bP3D��ě=�+n^��U���:��C�	3���8���VRH�ɦE��1�C�	�W� X��5t<!� kؚD�B�I�[`-�m�<R��`���9ZnB�I4S���X���+N`9qu)�f*�B�I$i�n�Y"o��H.��i�_�*B�ɳo��a�?B�L��T�s��C�.sٸ����Z
i^�.�`��C�ɗ#V8��GDC�.������U�ȓm�v�Y�g�;bR�0	�<����,;��:�b� #]����*5x$戆�q�	X�&<Q��MPr-Y�I+,}���M�?�>�p* �^�BT	��*C�	�N<\=2t��4Z��ޗ$�B�	�K���z$4�P& ���B�	8�Bd�FIF2O*a�$��g2�B䉁/OB(�#�d��s�V�Hk�B�	�v�$L$M�P7̈æ�X�o�ZB�I�
����pj�A����� �/XB䉊nМ}����)զZ�R�J=�C�I=VXF,"U�ԒTlx@T���+��C��-� ����%;�@t1V����C䉷gm���F�7.�`bG���B�I�� K�$�3R�>���l,/K2C��9By��Q�\�Ԭ��i�.x�JB�I2c���@�N*&Ȱ����]l$B�	�$M
e� ��W����t/ŬPNbC�.x�tZ$j��b����A��IÌC�	�(F^Px�ڀ�1�];(�B�I8N���)f+>1�zT��06SnC�	�c\"0�Ā�wp$���AW@C�	8 �6}"5b�M�>�S�4�6C�	�o���Q�S�Q' �/3��B�	�2���s��
h��*S �-"]�B�I�%���Ӎ�	D��Q5���JؔB�I1:�r�#MXL���(@hB��'s��ĉ��<�툑g�1	������H�v������
R�P"�J�"�B�I�!"ܸ4�)P8�r���!~6-�d���X�$@E��b(-8�3D� 3�lڢ~���R.6-�X#�$2D� ���Ug�!;Vn�d��`�0D��kM�bz`1"�>
�Z���."D���A�_�ҡq�ΰW�<́B44��is ZYb��I�����B�)� �M��⋧�����'?Q����'��ObyB�*X�i�6�	��:1>xXR0"O�8���E3#��p��o�f����<�S��8'%~�06��?I�"y�p_.U�B�搴@�ٜ_��-c$(ЀW$�B�I=b���]���&-~��B�I9�L�3f�af�cT.�66c�B�I�n�E1`��/(��c� bdB䉶=#���1���RF����� q@B�ɜ_�
PG���MH�`	���VN@B�ɏ
2�1�"��Z5p��&�ʿj7B�	&�X9��d�,W����M�;��C�I<B]��h�^���]�<�C�g�"(��%WTL�'1W��C�I�z0q�E�C����M�NA�C䉕+�6�17�]~~Zq�����B䉟.���c��<"(2�b)�?زB�ɲ.;e(�F�+OE���B�	?\4�!���Ӫ��$�Í`=�B�ɡB̢��e6mr��É�>��C�I�2F��vdX�]˦���>�2C�I+ ��H�� �'?(H1�CӍe�pC�	 o��cq�ǚX,�`��҅*>
B�I�U>��&#H<Lìu���Ҩ;}8C�I�-t�C�ƶِ��䩌	��B�I�%`k'g���AM��w��B�	�R��ia'��*�L)��k[�o�`B�I	K �����t�|-�#رLB�ɂ]��Z�fB�T�,8SV�0+��C��AI�i��^�W%JHˆDH=> �C�I�NQ2Bgq���uaG���C�	�.|x���H��J�� XčѮR�rC�I ��))�	��aw� 1$�0p��B�	+��Mhn��eh���'q̈B�QvD���O�3..\� �+m�`B��(�BMH�.߄J�t���e�#�C��F�����e"fAf�C�	(
�P<Q ���c.��0CJw�B䉢n���G�&w�$i�,�EydC䉚q��:#Ŏ,B����A⒆|.C��B�B�*��=>�\��p��>LB�	�w�I"e�!�<���[_ZC�	�{԰Ѣ#�^�A�X5�FE�2C�	�v�\�s�ף<
��i�B&%GC�	��4I�Y'(v����U�N8�B�I����d��"*}��1�Ȃ]z�C䉕"+4���(�/Ҟ�OZ�-��C��3��� ��m����b���B�I���pY�=b;ʭZ� ©&��C�I=}D.M($h� jJ�3�ݭ��C�IMJd�V@�fP����Z�h�C�I�WR&���(d�H���;]�LC�I�K2`@��۰$6b�q�,B�J�C��J�Y�˂d`t�a�� %E�B��4��$�&� [1E �
�4�C�I&oZ|��V�µ ��8�H��v\�C�I�%�,=ɱ)��>���z�G]�2H��=I�'<hp�D��m;jY1��9�Nd�ȓ@��E)gI*9;�|� P� )��'�}��ToW��� ��|t5[�$J>�yD�Nl} ��	<��!#�0�yb�yZ\�*7��?moHxB����y�+Ǿx�Xi���M4n��M�����yR��^�6�A��NXF&!7���y
� D���Ez5�a�cD�_�1�"O� ,��X��Pǁ�	�4�"O�Q*q�W� lXP����T�Rؑ�"O�uYƀ�40�ի��/G	ԩSg"O�� �	Y�g�"�q ���X�z�T"O@�֩��>J�A Q
̎G��̓"O`\t�\-m����H{� d"O������k�6�"Ƌ�?�>�Xu"O�����ft�!��d\&
��h�"O,Mеh�J�vB��U@��y� "Ohx3�BF5#J����,I����"O���2L���t�ϳy�K�"O�a��"޵b� �u�G=�J���"O%9"��pD=�Qi���y�"Or`ԧG 3.U�%K�9�^d��"O,�Pp��YLD�����VG��	1"OV�%$Ί)�T����$c09+R"O�%�W)K�T�j��QYo[�7"O��ې`� h*��@�4*�4%2�"O�e�H�樁�`��K�RM�5"O8 �#� j�(ph�GR�Х"O2`
B�!��Ag�mܲu9b"O�11dc��I\����V��r�h�"O� b�H��w��#� ��E0"OD|	 GW�x�����FҼ^���"OD���W�C�&� $�j�Rw"O �̺&�Zh*N4�ŋU"OPa�A\Ku8����e$
� �"O:a*㎚_3����j�Til<D��	���{�ک�@��7�����%D�H�aI�,P"��2�
�Pf�L��o&D�xC�g�(FA��x�ַ�{��?D�e'��7X��S�Y���ᥤ#D��(3#͎�,%����/iT��/D�T���ʗ_o�,D���$�<�� �.D����jJ8O'0��PB� � Arb,D��"u�'$)��ۆ�O�=���(&*D��{�\<$<�:A�'smq�r�$D��d>c��@F��"��D�&D�|�rEC:�H³�Z&aĚ�`��'D�P@B�1Q}ڰR6+����
F�+D����AN�OS�|Q�U;�咡�<D��@T�H�h��Y����MB�m9D�lC%'�����'R�D�	��7D�h�D��Olb��d�	FXQ "D�tB���4��\�ӥҒv`�-��-D�t �G\�#ͮ��`)��_��!��'-D�D0���Ry�a*�n�'�}��C,D��-m��PP�nP���}kVmϙw}!�ď�*����ONm>���]!�dԋaQ�dY�
�-z�rp�əGZ!��B�H�+ a\? }p�� a�G!�$[���aC�P9Wd"�BU�S-X)!�$�=%T�X�u�Ҏ$Lb�S��]��!��C�5rrgC�o���Ñ@O~�!�$�Ԯ|�Fᗈw��� 7 ��p�!���
�J=(��P<Mu�H���E�6�!��ҪD�� [�-^�iB���C�*|�!��Y�	�@@4L��	�(;#!�dK�M� e�֮Hh�Ax׭�K�!��RW�V�Pt�PG��Y��M�&�!�䆧5̅+a�'4�Vq���#G�!���р}k�H���+��˾@�!�)U�(Xb�ٗQ5V\��)U�!�� ��ؗ�e�r��T���;�|@��"O,uXU��!���l��1�.Q1"O�X��#�>%!�9��	J��Q��"O�R�ϋ)"�<l������s"O���b옸�4�ڀ⅄o�dl�"O�A�����Ah޴ࡠ��@�Vm(E"O�q�� �$�`���Jfl8䃥"O�1�����vyءH�'���"O���&!��ܢ�HK� �laP"Oh]:��\��4 2���q:B� c"O���a _9��}�E���	���"O���U.Ʌ�A���F~D��"OH�N8W�l��ϝ/5Y֡c�"O���(Q7W.
&Oϲ?8�8�"O�,C����H})�GDޤm�d"O����΍1����� �^��"OJ�q�@M�R������J!8M�1"O���K#��l���A?Gf�
3"O�p��\5ͤ�Zgm�44�ч"O��A�� �x*��6̙6Wp��"OF����r�}�%�L�ni�qq�"O�@�,�2Lj��b%�02O����"OM+��U�c�\q�dC��1洐�"Om�Ӡ���HA	��'P�~�h�"O����"�@+~��:0���k�"O��@PaĚH��I�#���:�ۀ"OfXA��<Z�� ������%"O�]�aY'j�^���4���h�"O�PZE�ɵ�t�`g!/�`i�w"O�I3F��'�,	rOP���9�"O~�s��@�<��Z�F3K�W"O�u�s�\ h�N�/Ɋ�xx�"O�Q���Y3h�vI���v���"O�i"$�Ɨ.���3%O>gm�L�U"O�y ���Q;� q��V�u��"O:M�^ ˚�xA��/x��m�"O�šu��7<�������Zi����"O�z����pXt/ďdM��!"OdA��E�+	d�Ӯ_�7/,��"O�}�6	�VN���ڵMfh5"O����0Wt�A��NH5���"O��p���{�$���+�x��"O��%�F�p�@5��%�+X� Uɐ"O8d"ԇ�w=|�*�֔q�`Hk�"O�1qhHs��;�շ+���qf"O��p��#ĘtҖʅg��I�"OR��:"�hᥬA�?��5r'"O�)�`��d��\��*�Ey��qr"OX�F�T�.���J�O�c%:V"O��aCN� f�����ϻk"��"O���-C �u#��]�qc>р�',|�v�~N`0:v��,<j<��'<�Y��!)*�C+^�L�'�0=��i2[�\��GC�%t*�B䉨y�T);@�/��S��?� C�	����Q�G�~T���j_�C�;�x�AJ��������4E��B� .�j<��F�d��P� . �z�jC�I���)�ւ֡[��m����W�FC�n-:A8�!ѱ0J�1�ш�g�hC�I3(��9(�B+rC�Y��w�B�	?5Z��HC'�0�ͺ'C���B�ɫ�Hi#�M�Z�V�8�Aӵ_�B�I \���F��v*9c���C�)� ���L\�%�e�͚%��13"O��(LU�q>��G�ϝBrg"O����D'_6�l����8�%�5"O,�KEL$��쉣Dݕv!�t�c"O��{BX4F���˄��>4&��"OZ� ��0 ��s-e3�PS5"O�����[4t��DbF�J#�!F"O��Z2��hC�)�f�5�|��G"O��V)�94l�fk �D?�%�"O"	��&Z$lh�dR�N��U"OL�A�2T@�Ȕ�D��@��V"O�� �ß�� �B@�6��� "O�#3JW�"��vk��'���"O\e����b�\xҢ�&`u��d"O�HGO̧=܌)�\$lXR��"OV%�ReS:s^����ºW;~���"OTM����x$�ѕ�Q�N>:hb"O.,����$v-ԁ©m-�%�1"Ob.EC~1`1(C�RbB=�y�N�0j)��EK�0>�`�ˍ��yr(�?vf\s"3�x����Y,���0>ɴ���O��}���H/A���e�<��*�ZpC&�X%F�ɫ�c�d�<����?�hڥ��|/��ۂ�Jb�<9C
6�����,��D (��Wy�<�c���:�AZ7:�['�|�<q�;����UJȓF	J1j�!�{�<�eM�!S`�R����\_�Q�A�o���0=�q`��9nD�;��Ȏ'�x����S�<�&쉋A	���֮B0T��E��S�<���R�>��YEA���0�R�<�!e�R��Sq��)P�v�����D�<qu&�@��yY�.ݫ4�MSf�[�<�J׉t�8�@�(@��9��Ao�<)u־�<��$P=A5���piDy��'��ؕd�6��+�*��]�Zl��'y�Lz�E�	l���3�%Ԣ!�����'��)(�FF}k����kE�	�',e ��ś	�9ya$ \�����'�����C�`di���Yi�y�
�'�{�f�!;!P�w�D,}wh1J
�'R�	P��D�&�c��$Q>�	�'��urF�H�w���u��i[ ���'4����-.��1���g>j�h�'T"�13��K��a���YN�tI�']���A/�A��0d��9�,�
�'|>5a��Pϰ�D$ǚ2�d��'�ڹ�5�K��e"ծ�t�x���	J�'ȐHG]�gPPa�,�Tϲh�+O"��D�W2r5�$$М,~�K��
!�d�<f6B�9d�ׄtT��)ߏ!�جH�N�7JJ�'d|��fR�J�!�$� m�����׎_F�}��>�!��O: 6��ñKG�8�H�"3-���!��ӡk�ْ��2���6K�+}�!��;����G�Ǒ
��ȓBGX&="!�Y	M;�<��E�-L���+H0-�!�H+j�f<!��f�\uIQj��!�$L�2f�(�꘠h���dHהL�!���R���J�6�����3N!��?+v<�hK�:��rT�6g/!��,O4�1S�#�v8����s�B�)�'�ژc� ���3Tk~s�`�
�'�\��� |$TiߙsC�

��� xD�ƪ�@�b��c�̸�B�!s"O~�+v��af�	6�D�����"O�xAᥜ�_	콫D�e���"OQ㡩�)`ْ!����b�� "O����iU�~�4���ʜ�%���v�'�ў"~�T�%8�"D0r��5�f��5��3�y��<l��B0F!/є�5$��yRL�y�| ��P�|| j��ٓ�y�g�{�ٳ7�щw�|� ����y�:Y �R�㙾j7Yc���yB�����EB�9c;�!" Q��y��"t�N��qeʧbT����/�y�m(�~y��oM6_�*�螑�y���CJa�� ��W���M-�y��Z)I�^)[w囫V�ܸ�Ɏ�y�S�n�r<��dC�&�RE����y��K�e´<���<��	����y"��
�x
�.��ء*M��yBNCϖ����)r6a�d��0�hO��D\��/	4n�Y5��q�!���'J���c�)�����rx!�.;"J�+�lųv
nܐ��ơ^l!�dU7
��rJɖ+�P�Ys`KBb!�$C��<�������p(!��'_!�$�D� ��5 ^�l�5i! �qR!�$ݧQ�F AQU<��nB�ep!�$V+ ��\���sN��P�,I�/�!���>(��YT+@�sbHU���v�!�*������QB	Y���
C�!�D��H1¹�q�9	tYC��.>�!���:(�@M�2`z�"����Ah!���<�L����Y�$6Ui�#��J��Dգ,��0P�Ak�����Š�~��hOQ>EV�٤-�ҽc�M�
(��C�&D�$��M�0~l�b�*ҝV<>�Մ0D�� Fe)W&̼:e���n0��dB0D�|@TG,b��¯M�&\���0D�(H��#bx�H�n4(Ҏl�/D�@z�OG7 ]�9�v�K���t�c�,D� �"�@���L@�Ɗ4{�I�L&�O��?#����c]�O� �m��B�	6o���H�hU1T&t���[;I�C�Ɋ7�HL�w�
F \�H���l��C��D/�$� I�V�T9&@�	C{�C��*I�|�q��,�R�k�1HS�C�	b��Y��C+x� uh��O] �C䉶��5C��F�R�><z�&m�|C�3��Aф�X2A�IJ��.�C�	+Ơ"�M?JB�y���_�f�6B�ɴ`���ٕgL� d��%/B�1)B�	�M��J���2��'J�M��C�	�b�l`A�Ӷ0�� ���o%�B�Iq��R 朇E��ps��1��B�I%DG:���M�]Zl� R'�t�D$�S�O�W���3�K˥{(���%/�j���ʅ�#�:�r��ЉTh#D���e
� q��P`�cO�(|B, F(5D�ȚeOU�g��5�"�NQ�p�5D��Hr�ϱ���#�9�� ti1D�X���M1E�@�V�������b<D��@!蚟4�5�#E�.Yے�Cdd/D��&@	-zܘpe�)	}r8jp�-D�$!�&��*�����Z�R,�$�,D�4Xt��7? �����OtER%�.D�� ⥐��B�"p��eh��R��
�"O�9Y�ˍ��Aa7Ύ?�N�)�"O����	
u��C-ߣ�ޝ��O�$�
 d|U�R�
�s���j0 ,D��1�,Z��le�jG*u4��t�(D���6h
�j8���oE 091W�(D�����V8Y����TF�>z��"��'D�����#6dRq�N@�N-z�:�&"D����/�,�JxKb@��8�@$���!D����D�B���7W~ƀh"�?�������RT%�`�j�/8I�t��$+LO�Q��LM�sq��x G]2YEXً "O6)P"�ǯ������zc"OZ����	[F�$�0&W�:��(�"O�ܪP�ٜk�r�E���s�}�"O.��wE�q��4i��ȥ|��R�"O�p���*j��P`(�����'L�\k��*+�\�s)R7J�vIؑ0D�Pˢ
R����s#+ �p���/D�@peǏ%#.8eRE���D	@����,D��:׮W��`+�/��"���C*D��p���n9J@KW=K6AXQ�)D�Ba+�\�r��T%�)}>�Zw�3D��A5�
voެ�b�G=^�Ȱ`@1��ƈ�����I�R��q��^m�@��'��' ў�O��`���^�lvi�%��"�@J�'�H����5d>l	�ną�*��'���;�Ük����5�?	�����'�2�i�	ۅ7������O2�$uJ�'��ʖ@IkC�d��b�U��5��'�X�9P�1$�I����O�,k�'�I+R�U�#�|}��Om���r2"O�5�ԳI���pC!E!p��˦"O�H���K�4���V�G�T&�"O���bR19��pN��t^Q�T"Op�C�G�J, �e.DHW���"OF�R��5C�����]�tZP�ؗ"OM�aE�(LTHb�Ԟj":�AA"O.��SCPaŨ����`�ne� ��y��q/J�i��"4��M3;D���T ]'jd���Ň+`��b'<D�$
�(��`ܶ����^��*�D�:D��CW�J34ՠ�Ì�	_.*h��%D����	�ch(�p��?����%�!D�d	g�ľL��4��r"X�R&f D��6�-#�@=bs�˥J*���"A�O���S�O�hy�J\]���ЀC�&��d��"O>1��O�*xRlɄ�F�r�\)�W"Ov|��뙲K�65��暟A6B���"O$Hړ��a���b�?�Ma�"O��r��_&T�A�c[�H�Hp"O>��`��n�~p�DAA��,z4"O�!�@�M0�9
#�':�b�e�'!��:(��Z�6u;��
�!��epT�`u�S�[���c��l�!�$�!���۔$�m�Ff� �%�!��A m<�����"y�c��)�!��E'��J��=yjU�5ś�j�!�A�=��Y
���@����QCLN�!�$F�nJ�Xb"��^p~l Sd�`p!���O�Y��K]�Cb&����Q�S"Ou9��)j�`�鴅�z&&<��"O��&���U��!�0��@��"OHL�UH�( �N�zwB
�2r���"O� ��IpA��D�"ႤN��C�"O����H&!�}��J�R�����"O��)�_��Q2��U�NG��4"O���B�� FJ
53�J��
�'��c
I'v]�,[���^Q,���'!�Px�A0S8L��Q�OG��j���8���Rc��7�8!Sh�*0����"O H��
Y0T�)	����?/(�s"O�	���I���0�̒�4���"O$�H�"*5�:��7i�l��"OppA���������^h��!��"OtXuR�+��[6%��}���1"O�#`��B�\�UÀ�A��e"�"O��cPL�-�&����9�-[�"Oȑ#�Y3@�M����m�b%;f"O��:6̈�"䈈%��#φL#�"O�ّTJj\;�2-혔�E�|B�'/�9�	V�TIa�놴?��]`�'���*wgS?	�p1'�n��P�'#��C6⋈o�-�"P�+N$B	�'^`��#��.�� �����F	�'��Pg(�R5b���n�u3���	�' ��!�h�b�a 2��̈�'w��Y�@�	�y�A��zb`/D�����ڇC�RL�5M�a��勗�7D����#�<zRlQAɕ(��=%'6D��q�O�p�Ra��ϟ^!h���.D�,xǇ�a����1�K^u�!!��-T�$JX�am��P�Ș2/=[4"O�4S塁�[Ψ��ŴI�j��w"OrXB�m4Q�� ���U�xqp'"O�}���E5nA.	���	>�6,H�"O(����^�3?�e�!Ę�"�A��"O�x��/,ʔ�5�$X��""OH��aD�^޸�9��x�@]2#"Or�"�D6#5�U 7��\���ZW"O�pxt�ھ6}�t���R.B`!y�'#�Ɍ	$(��m�d�R�u
I����4��S�`������O3{�L���л7~�C�I8\�J��I�T�k�ؒf"O�e�P*N!R��X�v�V�\� M�#O�	��O�3଒n�A�6y�b=D�����V`|9���>t�4��O<D� {��H44Vf�p�d:q�� R(|O�c�( R�֊x�f]�"`���n$D�D0��?���F���p4vE��� D�T����Y�d0RS�,fHS<D��b0a�I42H��+�<F�.��s-<O�ʓ���4��Isf^,	r�qB4}H!�$0�
#��k4�H��jN�+�!�	9y)��c���*-,��k��[V!�|��$J�D/q�P�
�L!��P4'�@|�v�[�Q���:�cA�@!�d�3R�����x�=Em�(�!���1K�,�CMهsGFA�o�-ў�D���ӠI_�	V��( �anO'mi!�<���iH�<�)@2�j*!�D��������^q.�"�j� �!�ʣ~2j)3K�#jD(� �օT�!�@	Yr�Y�2��)4����)�(�!�[��#��r���6�Փ�!�$&���X4�0�$K�WR�)�t��j�OC�Q
۰Sl 	�*T �lI�'m ��ڬ4h%�v�ՃJ������� j|p2*۴d�DXJ���stxy!�'�1O�� M�yKء�w�J��v�A��'��	(p ����)/Ş(���R�X>��$qə&�>M�������֬��'�>�)�G�m�ĥ�h��FE��'M�����b�l��!ȅV8��
�'���X'��B�̌Kg$�5&�A��'�@;d��2;�.�ɧ�݁%�b��'�����(�.UR��q�A�.O���ȝQ�|1A�6ZH�e�5���8�!��$E8�9��D	{�E��/N�z�!��82MT�z��� ��E��>�!��=#(-`�"O�F PZD���!�$�;*��0�K3o�0dq@ ��ew!��K�j���9��������_�L��yB�?%.�8I1 _7D�T���F����.�ɅژU#(O�g|�X�Pf�BJ/D���O�00�6=�G� !���"(4�hb�HJ�?վp�a퐜	!r�fJ�<��p�<��a�մ	��gG�<�q��+����� ͎_F���C�<�Fɠ1�x{�׋9�J�1��v����<@�VW��QF�Y�e���[5g�s�<���~���fс\(Ҕ����g�<� �J�+�n���?{����Ga����<y�±k�pȧ��$z',<���f�<)� �#��HyB�"i�9���I�<�/��$W*�a�IX�AN.M��G�<���5I������� �Q��z�<i7b9S�>��6��r�=���<ّHV�P8�pPF�x�9�@��{�<	!��f�T����mC�	x�����Γ1����B̍�iqJI�è��#�0�'����	�Q�J@���F�*�A3&�1�C�	 �\��Ëǚ8���"�B�6�C�I)�y�t/M���<3D�^�m���d:?����j,�#ɮgg�i[Pe]r�<���UQ���U��r���M�n�<q �� ~*\��I^)�� ��0����N��?��C�j�̆�$�đx��E&�	S�)T!�ȓ�Hma6�7�X���Df��ȓ���s��P�P���#�*�>h���	u�'����ƏX�)��|�v�V�>@��'�4
� ��G�6n\�f6�M��'	z\�rꌊsDj�����^���'׼�2�/��@�&�r��
��Q�''<�A��M�0��RF`�'\�%kG+�hŔ�"wǐ�ug��z
�'2@��B��Vz~��+`6�� �'��!`#�T����D;G�FtC�'9Y�����Xa��-,�u�
�'(����I�dI\�K�G4	~<]��'�|�3G�G�R3�-@��ŸU� �Z�"O�� e΍ B|�H���'k�,��"O!��	�I�<�BeX�;��l �"O�9hV�	����%اD�ܽb�"O"U��  ?!��E��/�N�)5X��D{��Ɂ�[� �+��ݾ[B �'$�OݔB�	* �Tc �*Y�Z={�N��h�B䉽Q&&���O�%9�a2���-!8�D��5���C��(LMy�@H(C��C䉹Y4DA�d�E�f���my�C��%#ߤ�B�.���&AlK<�?ь�� "p��*�/Z�6�a��@�p�U�'��IV-
�%ФE���P6��D6C䉎�
 �Oߋ'{� y��jC�	Q �ȡU�Ƽr�n	�T��X��=��?���	O# ��¥e��T 4��lU>c!򄉄sT�Y�S��0��G��?!�G�'���3A��}�-� *�%N!��@�pyА�b�� 5��9V�Q�lL!�D���!���J�
ݰs�WH!�UD e��L nn$(I`���(C!��ڭ\�x9'�0+R��B"ā<!�d�L�����3�m���A�
3!�$وgm��S�j�C/�5(��+u'!��ʮ5�<hk�H�N<�u�V�*ls!��A�	&��Ń�B.�p��.Mr�{��d��O&ب�B� 8����0���j{!�D�7E�z��ׯ��?�l���� G!�$�6x�椐��B�T/�����¨{C!�$�\���Q��{ ��p��8E3!�Ă�M�$!8�&G�U7����b"!�$�T�B�#�V�_�p��`2!��e����A�t����Q�L!��#at�Yp��.M΍��n�3��	K��(�"�).D�f��@QD�&�I1"O�A�%�6<�����-t0�1(S�	G>}�&L0��N�j0�0Ģ)D��S�g���2r��$ 2��C=D�d �`!L���c�
�z��A�<��?9��I�4:!��*��6z8)�ls�!��M�l���!��h�C�X�!���a��MJg�U2@x�t��+��K�!�DJ�{ X���x_�3wj U��'mў�>A�OG	��K5�Ȁv�Y��;D������ ް�bE�Eo�!:D�a�ҹ#�6|�Č�7on�4D���B>E�,ə&�0]�3��<q��哣�e"dL�$|��RV`(���d0~���dd�*�f����G ���&�����h|�k�I�#/O����/'c*�Ot�O�=��]N<�����Ia2��k���yBCP�C�%3��Z�KxPq���û�yr�S>z�l<A��:It����ּ�y�b�?SN	�S!N Am�4.̶�y��u���Z�`N�+�^4cʟ��ybl�LSXL���C�FĹ��U�y��ߓd2B��&�NO����Ҳ�y�BR<M��������I��\���M6�yRE�)aQ����˴D�
����=��<���K;h˦�c�K֘C��Q��p
rur�AP&{�z�(��Q��,�ȓ_�$}1c$�u��l��I������|�ꈤx��msW̅62p6Є�Iw~C\�?XT\a�e�8�L`cu���y��Q�p�B�o-:RBD�$�M��y2�GQ��`áͲ,gM3� ���y"�VZ���M7;r����yrmA}���ƞ	ـ�$C�7�?�����'p"�'F�'�	0�B_6�����8Q}�5��"O����.b(�, A<c�pdۡ"Ox`ʑ�T9x���ƒqb���"O|�!œ/gz��r�J�0\Tmi "O�(�Fe�NP&���TY���E"On`u�b�����pQ(Q��"O��*%'�,)�0���N�J_2e�|��|�Q���|� �܃#�>%���3ՋK@q�"O�L2��ڑn���ᤃ�y�b�p"O���P.}쭩僀�8�2���'�09�mۢQ��]���$"!��#D���J�%~2lٖ+���]��!!D�`ۖ���zq^ �E<6z��,>D�L ����\�����WILѐ6�;��?���O�@u� �0@�\�c�
��J���'�d$����(�i� �/F��8
�'�)���9B\� �Qr���r�)���S���*�+\?(�����$�y�fҢKRN�C�&WE��
 �ߝ�yjZ<�T})ԥ��<�d h'�/�yb)תyF��u��⥪C@Y��ybb@6;�8�A��0$�y@�$��?Y
�'ݴ��͌�{��p���|�VM��'v�ɹ�bޤv�l�&"m���p�'h��x�n�*D�t��.7q�T��'[��Q5nI�$���V�F�c�e�'_t�A��G�~t���3n���'XR�y�����X���Up�\8�'�>XSg�է]޸`���\%֕�	�'-ʴ��$�;m^��0!�2t�4D�	�'EʐK�g�AC~x��C�s͈���'�Z�%�,Y�t��2�@!>>V�z�'v�4�c
L*M���bC *	&�ݱ
�'�t+�&�D� ��W� `�	�'���Rb�1NH4��휒�@�(	�'Jh�� ��9wJ��f�W�,��8�	�'�p%�fo�3SB��5 �>�
�'P� �4$�%�,1�Ѧ'҈К	�'�4��(UA�����b%B�	B�'�>H��J�����O��$�^}��' ��{w�Vp���f)б1�hDk	�'l�Y9q��d�)(�IA�T�(�I�'a��+�?	n~]���Sy�xK>A���IO�4@De�寓�Q���c�*��,X!��Z�X,��Ŧ 5R��ͲuJװGў0��	[�v�&���>��؂4N�VB�	6<���e�$1�@��P�giLB�It9���SJ�!���+�� e�*B�I�:'(()v�޸ ��uyȆ+�8C�82�6U���/�eK�,C(�����	�RX) ���:~r��W,����B�	>r�b���H�,���=�B�4Zx�O�~&��	|�|��"O�Y1&��6�5�t	ظFt����"O�LJb�7rư��肀NN�E8"O�M���'M(3gٽ?AfX��"O�阆��f�Фۆ �5h��$"O�X��"��2��D�� w1�d[�"O�U�׊�$�,�1��ǐTG�r�"O|d:���w�<�"�g��:�%{"O��{��'��ia�C\1��@�"OހJ$?<�4���}d���S"O�YH�z_���g]"��3"O�0�V.���&,k�`#Ҵ�u"Or\[ ��w9�DZ7T|�(��X��E{��ɍ1~���%B]��Haf��S�!�p�  (�7�$*v�9Ee!�� 8?Kt�Z��Q<I'vP�4휩8W!��_��u��m�7�N,
Lʫ4D!�DD]0��[��- '%��i)!򄈦�:$1Я@6j���h n�2p!�� L'IJ�7�nI:#Fۅ���r�"O��s�ȏ1U(��v��2�$)��"OԈ;�[�:u8����80�x�"O��ua�2Q��5��Љ ��s"O0DC`%@5�&Xcf&O�vzh�ڶ"O������4Q�8R�Y�.q�"OT����߬OǄ<x�b̄gY"�Zf�|�)�,_	��˶�1\�2�j���k���-�<�V�e8%��×xOH*D���C-_>4s��F��<m.%���&D�L���.�� 1�T.n1�Vd*D��S�CrTL)yS��7z��\��-D�|j�a��� ��g�(�L�`�+D���@�=����O��IS�H3$e(D�����H9t�hc&N>Rd�#�h8D�Xу�Ǳ>�*���0>o4�ٱ`7D������o�,a`&PG,pAK(D�PH!���M�2KNH��L(D�D��cH?.bU"쌭Z5����'D�$ytə�lS�	�,��\�9��*O$|R�hM%
���X���r**Ѩ�"OPy`&'ɁvW�`P��D�J�0#�P���	n���O��h�@�#Ub�R��nǢ�����?����	!pn�0CaJ� ����̗s�C�	��,B���4 W/�B�	#Qz��c3v4-fC.z�B�I�BW��p0�O�m	2��S�0c�C��
r� ���>��"QLN!T��C�	�!����F�Ai���%�zC�I�
�����f�@�4T�H��q�:C�9<�p٪���j�0�3�[�o�"C�	&�
� tY4p�)�/'�B�ɗj�(ԉ��b�5��
]M\�B䉥J�>�Un��e�����Ǚ*��B��\\9#U�PYLAC��P0��%?AAj�.>\��DD�_"����E�<I�C�y���*M�&���1p�@�<��>Հ0�@�аc��QD+�}�<!$�7-%�e��J�OG�P6��z�<q��Z ���SM!Q�,`!G�l�<��ީ,&<����bA��p�i�<m!�;o�Xɉӣؕ-W��X$��g�<q�Z>����];A��a��e��0=D� K2a
�4 P���(O_�<�򀚓$��03F��.�jp0��	U�<�ǏƐk�h �3n�}"`��7"�f�<a3��(�1�F���<xtX��x�<��BS�����C 㞡��B]�<I���= ��Uۑ��;.����EYh<�6Û�z{���e�D�vml���CE��yI�S֊*QcR8z�+�m �hO�����/,��J�Ԡ@�ㄆ�c5!�dY-$��A#c�0}�%�!J`!��$0����n���@�Ș>|�!��S�
�@أ��L��.�q�PG!���(���C��%F�6�򒈉�%9!�ĐE�.(!�С�ְYf)с�!�A08���P���D�s��v�!�䝾U��*�J�!���P�תi[!�4,����CF&u�u�#jʉFO!���Z����ˁ�}���O�)1!��º����>��E(��9~A!�$�[Ӭ3c�&+�T$��,F4>!�U}����Q��
�-͘v!�� ���EdA0���Ճҵ�������Ox��$�4D^�)V#v��� 6f�c�!�$�V5:�#���k|~�3�dY�9�!���b���Q��/+?�C�1!�䁂 �XYg:X4xա�2�!�䋜NfPDQC�i��4Z'�ܱl|!��/Mΐ,��	�'0� a(��".�!���5]!ZtB�i��C�����7��'�ўt�<�$�4z_dH:'ϐ"7�ma��w�<�6lB�w+��A�iנG<x�2���v�<1!a̅P>�9;�ԛN���R�~�<9�J ��I�RCG�t�@M�d��@�<��X� �p�&АwP��cma�<	��]���0	��Y�,�BdSY�<af���0X��A5JDIW^�ac]��0=)�&""Zl�vc\<Ф@���[�<��+â�����/^�h�@�[S�<ѷ��6w�-�o�i�Du�H	S�<��N�(�`0��<[�,Q��QO�<i�	��	��!d�4z�X�C I�<�Q̌5y����N�D�޵+�A�z�<q�	E+T��3���*v<�{$jw�<q�ZW%�Ib
��XQ�u{�<	ϣ,vjL�&e��,��]�<����=D���xd
�Rq��w�<���,I
�u� @�̄�ԃ�y�<� �_ت,�$ID0Rfl���^�<�Caܤ)��dj�hE�'��,�7��X�<��	�o�дY#-���|1#�
X��0=�p-��Z���E("{��C�k�W�<Q���G�(��&�q��s�W�<��ۈN��L8��û
����e�DR�<��&�:<w�yS@�8��4��G�W�<��\�h�8yE���B���]R�<9q�G�H��E�t��(��P��O�<�bȭ~P�M�Bi�H�|�K�VH�<�Ŏ�)"�D����#2BG�<iMTl(0�f�%iI�J�/�E�<1���>-���#@��6o,��Im�<9d��j^By`��G�K�U�@+�k�<#���(��=��I�\��=���jx�ܕ'����lO�YĲ<�)_�K#^�"O2@q4��!K��Gܛz��4��$8LO�3㒇K(j��G�����"O��H��HI՜ɑ� �tؐb"O�x���ȧ]��]k�^���t(S"O4!X��#r�x��A2~���"O��;`�5A5�@a[?�̡�"O��2�L�"K�����X	�d���"O|�h�G :��bk�)�搀%"O�(��J�)2Tɠ� �k�>Q23"O�y���U�}��0a"���6��,��"O�-"�Rv@K����S��ȵ"O�I����*����y`����"O<D`���0 �l��Q�B:ev�ж"O�i���P.]`*\�Ѣ�cNP�2�"O0��Dmϊ:A Z�j�VE(q��"O�P;䆣%�4y�!�L�'��H0#"OptiW0+�T��C o�XBU"OZ�p'J�L�b��!�H$`�"���"OV��\+�0�	e�z����"OZxi�Ü&<ԅ�6���vt��"OD�:��\.��y��	[�oǸ��"OV��c �2d�6�9�邜_�nI8%"O� ��a�$�2 8e���;�B�s0"Of��S���xܪ��U*��̪���"O|5DgJ���	(cG�
�y��"OٰF�P(l�<���X�5��"O�H�vD܁@�QWJ�d�3"O֠��[��0ɻ��6�zȫp"O��2q��$�� ���(,����"O���`N�i�X�W����6�K�"O�@wG+|������ܳM�R)�"O0d�a̞S~|%xR�+v����*O�����=tT�0�#~����'�0��AY�v��l�.X!a�Xi��'��S�:���4��,_�(�c�'.��ٓ�L�
�z!����?o��"�'M��AA�YB����&�=*�*�'vK��4��/������h�<y"��.ja|�%j�0%c�1��e�<!O��t��t�-m| �C��v�<����y�p�լ`Q䘘D`�K�<9����[ش�bY�=8��E�<�m��RQh�(`��17�	�I|�<�6��5�s�m���8�H�x�<i���N��,�SEp�@����It�<ђ��>C�%k��/=�D�P/�t�<i��!@fm��B.��03*�d�<�Sc�2#��(Q�K�#���']�<��N5���q��C�F���zQPb�<�UN�1)���ǇŽ�h;2�L`�<9�O��b2, ��Ǐ4Nb��B�<���>�V�(b�Ҏ(�؜R��~�<ibiрaNP�L��T<���|�<�!	�L!#uoT
��	4�P�<I���b�*��!��2�SV��U�<�2ꉑ*����H��_�)�ס�O�<yCO��f}2���M�I���As�p�<�����s�8p��?h���	��IH�<�e� n�H����� ]����M�x�<�1��lB4��]�Py�Qq���K�<�!�J�!�vU2�цUJj4	�AK�<IU�qג�B�j;����q�<P"ՂCјi�l40�D��W�<�W��)%@P�Ȱc� �e��S�<�"HVj��8B��4ztqh���I�<!��ʷ\�2�T���D��` [G�<A�Ϙ��6��Tk?q���ȓ}��@�eO[�n�Ʊ��Q%r2�؆ȓyޔ�ˣ�A�(�R��"%��E�ȓ r-bwAH?��Ũ[8q���=a��$)�[|(��l°||���ȓW��A�%�7�|����QMzl�ȓy�<5����n���;��ץ���ȓ~���Q��,
Pbq���BEf��ȓ^�z�dk�e���tHJ�l'��",*S �aqЙ�E�ź|Ȱ8�ȓE������A�VT��z4Eн̨�ȓn�R��e��,�ljS�0l���ȓdu�d(QՍ67>T��ҝpsVe�ȓ\�LCV
�(\$�j���e�R���P����c�=	��W9b)Ȧ"Od1ۑF��+���Q�&��O�D�u"O!i�G�֞��d�0*߲L�"O.�c���0S�|�iqO�4�0#1"O�`�£
�ļ:D���6˪�1"O<%z�.�Or&!cfP6�4u"4"O� ���B�M�6��G��2�~��"O�,J�LF�� ��.G�2�,ٶ"Oj���˅i���p/U��^X�G"OJa`.��p#�5��Õ�Um�i{�"O��Ӓ�).N��#/A8b	��'�"�e�u���B���T��'0�4�&�1}�|t���"j���'s�T	4�0�SD��Zqd
��ǟ�y�FD�I*,�J�(��&vJ=�7g4�y�.�@HzEj�!?�I��yr�8�����?�H�iZ��y��G%0h��"2j!-�F���*��j��\:H��G�^|�P�ȓPY������.����FD���ȓ �\�$�Ԧ�X�҄��%eV��ȓ� 4�fK�0̪��i=2���T��� ��hH�uʔ�
�4���Tڞ%�C��i�ZYJ�N5U�H��.PL�� >~�<퉅�ߕ<�m�ȓS�zQ���ԵX&�����K*p�ȓ"�V|3h`���Q6bA:�,��ȓ{���E�:k]h��υ�trj���Z��X�
��
/v��Bn\�Ix��b͌���R�O�H��'U3t]�C䉴r)��sJV�f�、1"4C�	6,k1���\;AL���	M�8�
C� :����S=$�00#��:c�C�ɉ+7<�paZ!O�0$L���B�	1@���i7�78G���BQ8P��B�I�a� �k��c��,t�Ћ|��B�IU<a��=@Hd���L�hָB�1<��� ���c'{��C��B�ɆO2� f��H��I�&���(�C��=
B��3A�P5p�����-T:C�ɻ\vᑲ��,zqti��_ 9 C�ɋ{�L��dL	�5H`��vB
�+�C�I)��US��ݩ�0�hqeԝ%��C䉴��%�֨�t��ْF�:Bo�C�I�K�r��b�261\" ��2�C�I�n�d��"��D���;0�I%O��B�	�~��qaE��j�БB�K#}�jB�I{lM��(�:�9�Scׅfg*C�	�F��f��!��JQ"<\r.B�ɜ:_<��R^:�m�Bg[!O6B�ɏZg��Q$˫K����W)m��C�	�^��8[Ul�6dڰS��S�a�C�	�@�ʲ�)"� �w�K?C�ɬx@� S"BQ���	a�N�e&�C�ɉxY�={`�P|C�\X�	�%$*B�	�qw�:�"�%�� �K!.�C�IR�:Y�`/��T�DIb��U9[DC�I%@^��9�!"~��CgN�I�B��.ю�J�DV+��D��eMF=zB�	�M���i�%S5	n���.JY�C�I�tA1��G�|q�H�!�E�IW�B�	�H6D0W�X-U�,zf��8+іB�I�C��͐��'F��mz�f�9dJxB�I)x��樝0�͡@�_ XB䉧6�T��d��EWp��Sgްk�B�X6`فG�;F��+���L��B�(qjJ�R$(�/TX k�ڋ:�hB� �R!�5n�E=R4S��T���C�9$�@���jD�A:ԑ!͕!O�C��(���cϘ	R�Hµ���;D�� 6���gP?F��(J��vʑ�"O�D�Da�)��ݻ��O�NpT�"a"O�q���J���mF:JO��t"O�Dq���td4h� Gl<��"O(��/�~0�[7X�W:���"O�0��%���0��(8H�=��"O`��1�J�70"h�,�Se��w"O��2�#0b�JDj�
Oa�P�'"OŠ�*��#Z읓1C�%�[�'0��'H��æݺb�؀���
�D���'�~�ժ�&@��Y�A]�J�D�s��D��HD�Ĩ��[��Q�_+��#���y"e��lƠ�3n�5Xs��#i]��M{�m%�S��M��+@�+f��hsO��2��G+�w�<qCGS�/�.X�$/�}��L9�k������p>����0�^Tk7͜�B4�1��,r�<�Ǭ��F�R�Z�d:zz�`�Äv�<)�":S	V� #��v}�-@���g�'_�?��Q�+�:A���w�P"�,D�Т�BE�p�XPYkZ%"`�\�b))D���uŌF�|��Aܑz*-�tG&D��A���Xd�Bc/�1�BzE#D���&ܡq�����FӚ~ M���#D�X��J��H� +��[�&�@]qce>D�1���)g�]�2��9<��DJg�=D�<��M�4�F�22�W�9ʺ�GI<D�4�dMW7WiΈbF�+���0� D���6du(�X�6��~n���uc<D�$R��,4��#�M�T�Ԣk%D�#dR(ːTC�'ԥ.縱zN"D��"�NM5�Y��e8��1��>D���RPC��ؒ�͎=��B3(�<����S	J�$-�"E�~����T����C�ɜkaF k����`T!b�0C�	{�X9[u������v���W���Јy�JX!u�ƒcD����W4#�!�;_20���J�o*����n��!�$�x�JɃ��/;��iU#�3-�!���Gs�����D0�tY��+�1O��=�|Jq��D�6��.._�x8��k�<�P��9�vA�uV�Ԑ�!��Q�<iFÂ-W���ōTU�b�w"Kb�<A��˟xʭ3���X,b ����a�<�5$)L7޸���Ǐ}=ƥ�D�T^�<�����A��T�C�'H�]���\�<�`�!W�>͠��F�#8"���UV�<q�[��(�ką�1����ClAL�<`DI""�|ʳ�ȯ-��T��Dl쓇p=��&��/)�h�M�+.�J����q�<��`F?��iW�)
�r	o�<f�=p�\<÷��%@ d���U�<ѷ��o�e귉ѠL#�!��CV�<�2A�q.��e�S5S�X�B�(OX��&�S�'>'�9`vI֐u�>�Pd�.WM�ȓ�|$�˛(0�8�&Lۦ��ȓb��{ԯʋK��3`T�Z�$���kf�0膠"�����$����C��:,pA�!F�;����f�m3X���J�طM]�_Dfu�@G?l���Ez���K�Ol;'̚i@Q�G�w�����d6�S�t� v-MZD��(Bڐ��n�<��$4�S�O�,��Y*P�)K����>5ˈ�d1O�e+���+t|65L�%t�&l�"V�d��'�$	�* Y�,t��$�I,�M���+��~
� ����d��K'�9b jݫy恸P"O���R%QY�L�0��S(ᶡv��j����А*��9$m�5%��(�D�1O��=%>�X��s��)ëL�%v��&���y"oK�V�l<s2c�~U��`V�K�O�"<�L<��Ks���r��;��z@��~�<�u��?��#���I�.e��Lr�' ay"�H�~}�������D��l�y2D�"<��aŊo�(����Θ'��$�a�?�LA6Õ+]z�-��e-��"?�u��	I@�q#K�&^�L	�R��FY��O<H#u�N�_���r�M�t[:x�CT�<�'�1O@0�}Ba�c��,����8M� K@�=�y�+>s��5�Q�k�ʨq�JN��L�
�=%?�(�M��F�)5�M���4�� %��)wB�4[�H�	!�N.4���JQf�>#�ڢ<�˓Po����A�"���k�C<�q��	���D:}B68NȤ1W#�<Y1���G&��hO����Ɏz�l��2q���"���(�qO�7M��ا�-�
�Y� 2O�*l��f H��m:6"O�\�
�8DP8A�o=����$
�2�HO.�D}�	6������~I�yYDDشʈO��c�b?�7K�K5�j�r;��C/D����)l�����p����Er��'�>�O�>9 �� .�jE@F�rbl)�d �hO����7��y����E��A���F�5�ay����z�r�#��3��=���D�!�(B䉧_����	�"o��IW��sA�B��=Uf��)A�	�y�)�f)��uZB��;,H�Ժ�D�dc��ǎ��"%C�	�����
�o�$��D�-��'�ў�?Eٰ*2ZΘ�孅 jC��K''D�$!�E�;���IU:i��M�1�&��!���#��?���A�D���{"�M�5�8سO�,KO!�D�{T� �'2ip�t��!�N�!|�R�O�,��jb�_�t��{�i'�H����'�W����#hX^Մȓy����ǘ�t<PT��'�t�ȓA1����[���M�!{�)$�����91b,*fD+�>P�UN�	f��=Y�Z���cSH$��$�g��ȓK-��Ð�N�,q,�0�Os�t��n����T�G�brR�:걆ȓJ ��F�M����"u�<2�p<��{��I$$G�p)��	�����J�&5xP��Z����C�a��,���f)�փƵ^�Ƞ������
t��b8.�x�aF�|��xzSK�H��%B�	h�'ǅtԦU (ӳKih,�=�'\�x+ϳT���@�'�@(9r�ۊ��?�4�M��i@�*w"	�&�T@�U��BR�<�l�_ߔH���Ȼ%�("w��Q�'DQ?�z�$WC��%Z�&XN2RI�O B�I�- T�h�O�J��!��+�� 1����5�	�=��D*�e uߌڐLT+l��C��(N!Xyڧ�+=PPu�!e)i:b7,�S��M[�ƚ�� �A�$���SUa�e�<�t�Ł=a������n
8Ȓb[�<��-B�:�p�Ώ!fxe��+K�<I�J�2r�YE�43��Tb�k�ɦ��i��(�,<K
�ǧV�K����?!�Olʓ��OԒ�����D^�H�f�N��4��'+Iիq]����^�kf�M<!4*<�S�'A;b�:q�'4b�p��'Y��%��S�? 
4�ak�0U@�3�CJ�NÃ"O�0ٖ�ɪ��x�D凴3}��R"OB9CgOH}�b�!3i�uC��O*ʓ�=!B�V�m3rI�Չ͓Q�bu�S@X�@��Y�ʧ�O8�F2�,[ ��PM���"O��D�72Ԥ!"��(Y޴!���N�(O�O0�
V�?	0��Âv���J
�':�QZƋEd484#E#r���	�'�|���Q0��Ó�2o3p�
�'��h�� K�O<J�SVe��� 혉{�'j�>M%��QcB�5ry�� �F�<Q4�/"�؅i�:V���ېfEF�<1pOԊ�1DA��d+�1��J�<���S�1Q��)�gV�#wz�*����<B�	�\�lA�WC�{�L9�үD8�2B䉸J
4�&����*P.8�B��:lHzf�1PM�����:V��C�I!A`fY�d�ѽTp�Es キ1�C�I�+G��j�F�7�6p94(��J2nB��B�;��c{���CA=A�FB�	G��Z� �#4h̀
F�,`�8B䉥'b���4)O�SA��Z���C�ɏ"]1���	9ɒ� w��*��C�	<�L22J��1l\��/ٗ|q�C�	M�����E�/	+FذO�?]�B�I7qR�2�L� �h����H	�B�ɢe� @�A��u%�=13僰�B��0U-�E`��f��U:��1ie�B�I�:�ЁC�L�6�ahD�qXC�IE���a`Ϡ-��y�Р�O�C��:!�F�2`F�76�;�/�8y��B�	�9Fp����m$�5�&�ͨ6b&C�I2s]��g�G,Z��Rs$L�z
C��-PޭW�@�2���a�E(:pJB�	'ojl�E(B�\���Ʈ�xC䉞��))�"ɟ$>�1t��&W}B䉛=��ء  �.wtH��t� )�C��1W�,y{��*C�=�vC��s�C�I3<Cd�;@c��E}&���%�K� C䉙#D�[�K�&N�)�Mְ �
C�I�N"�|�U�έ}�13G+ 7�B�	Bi�����I�J�E�$M��,��7fp��b��L�P@q�O�7����?7L��m�;<�i��C�
�DH��h�<e���K'0 u�q@\�L��a��	�"��4Q�i�dИQÌ�6@Pԅ�9/L�@�D�u�^-+r-�7W���<Q���X���"V�!�q̓T "�b�X/8���A�8�݄�6�%R`�ԩ{Vl����-h�l1�ȓq(d}i�nՅ4͎�rs�Э;؉��\�$�b�h��ٙ"n��0���ȓb��1A�dtG��pk$�ȓr�p�( D��M粕��h����P��R��CP�>�zEIG�K(�vi��ˀ� ��\'��j�R�b��ȓ��1v�[�Bm��p,�u��؄ȓE�Rl�1F �7>~%b�勄T'�q�ȓ%����XOF�2���]�8؆�f(�p7�� ^����Iu�
��ȓw�-��,@����H��?
݅�&Fŉ�T3<Y+�n�snJ���:�H�n��,���%�P�"&����wF�"צ&M6�)5�):�.,��(c��s��ʷ�$���vi����S�? ���N%O�>��%R/�h3�"O�=!���(թW��>,p�W"Of(��
�/˰\a�#V	K���%"OzM�3+M�{=��r�!C�~���:"O���T��7?[t��Iyܤ��'�,ua�c �D�a|"��o��p��G�<�Y�O��=��'�Ie�ium�O�����G7B)����'id��"O؝h�*���нD&�.dʡ�u�$ɗ0����:�R�Z����7�̃��(=�����4[F!�ą�pQ�IBp��Y�ҭ���"(L�X��& a�(�'���D�,O��k������i�K�R�$�5"O<��D�T
)���BBI�5P���H �SH�Z����,!��U��I��4�P$�3����0�V�r2�����6;9 ��%/�>6-
�^���
��<}ȩZP�E��!��r�)�ƣpi�}��^5qO��B��d�t�S!�'0��b@�ڂB<��baFY� \D���8�g�$fd����/Pt¼0!�H�FuV@�`R��)��<�waZ�Dv��
��fU �Q a�N�<q�M8a�ʼ��aĘN�TkCbG,Ԑ#VH�iJ����'q�e#�g�#I��<c�	�lg���g:u�M�� t���:5�t��"�E�C_V#���pm!�䙮:dH���R�KV~D(���/n@�Ot��MH3\w�"~����=Q��ΟZ�(��D�N�<��O�5f`E�v�GK��$SE��E�<q�G�j������<c1
W�<�v�� F�Qh 	��y�5��c�<9���=�jU/Ň<�ډi���w�<� &J-	�(����<{�`���p�<��͹{���c@�L:I����C�^o�<����ՂU	��1FTؑ�G�<i)Y�^k�(+���w���L�T�<Y���;vX�+�F&h1G�U�<Q&IM�i�p�r���i� ɗ�K�<5
� 	������u{ֵX0� F�<�3���%�����$"��a��k�<��[����d�	���!B$[�<A��A�I+ze���!��E�^Q�<y���7e�,z`nޫF��x%!�H�<�ńD��ْ2�
,�P`/OE�<y.��-�nA!�n##�T�#r)�A�<iC�9AR�1㴋�l��0p'�~�<���D�|�b���D�Xခ($ Hv�<�����8��) E�]�^ɺ��RN8,O\�[�;Ƙ'�2��",ԋj�R���x��i�' ��k��zf4�؂eG
b꾔{,O����*���J��|ҁ΁>�� s�^ɠA��Ŗf�<yq�`tt ��L����]�<ٵG�wo^���%N2j�|��ǖ^�<9�JN�i�@q��$ޢy̚���X�<q����À�	�\��Ƭ�C�� ��׶f�X5#Sb̰�n9[1����%)!�@�=�ε�ٽ|�JcaF��OZ�kR�$&�2��)J�c����n�4��􀒎��!��_%D,�j,����H�M�"��Eb�A+7���c�'�	N~BTdǢl��'9�����]�jR<�1��O�b����
������r-v!��O�,��eW�H��p2��W�.�.�q�LҁoZp����H�q*z1�O���Ou@\��'�Q>����L�=np����'?�c��N���v���qHP�v	ۃO�P��u/�*�4��6�ż��!���^����x�|�'w�U����W"��S�Z(��4��4����<$B�!��H1�I��nХV#q�k,Umh��A�ʩ#2�%1!DM'=�R-��&1:��zBc�R؞X�)�r�$��hȻ\z����A���h����#���ەG�����u�r�*��wAе�>E�b$N�5�-9�Ŏo�N@1�rX��̓dT��Q�T �l	��Ҡ+�n��)vBIA2�W�,:d�ᱡ� ������'�r-��'o�p�P?��U��,&�<�Â��P�]7i=��y��M�!Q�.�6��$��,Pj� t�S�-��zH���f���It���C����'�_�o���#h��-�~�'֭yrE�(>ui���7=�`:�4�y� �+���C�ƘJ�(�S�KR{(��\c<~�re��.qf􌐔��|����£(T�|�B���OCR��ӓ�ʕ!��T�r��i�eK�/@��p���t(!�jM;x�غ��#}U,�O��u�e�K�B��h�q�KD�$���D�A�F^5$hm��I�IC�P����ɐ�1�$��f��M�#�c��`aQ��%C�`9��^7?3�I`�m��'�����b>�)���<9�0	6�G�bT�>�k��XK`dنӜa0�gՒ|x]��E_�4�,q�WJ�9<:sX nQ�1jÌ��y�xК(O�M�h-���$����8l]���N��w\���O�<��׻��m�R��`l0��Zn�t�È�lM�T�J�(��r	֏�~R�63W�Y�Ш�V��$X��4r/�}RE��ĝ��K +.akw��%0Z�����rH�b>��Q���pM�4H���a���0r	CVA��Ї잜-��Bተtv<`�dJR�K�v�A��&KF�a��N�*u��i��"0p����7A>x�$�W���t-U��-3�'N!	�	!�0��<9��N�
�(Q�� �X!�aD�8l�E�E��2T:0*��
�"B����;	J��#���4�����7�p�$����;5�z�� �88q�(������S�lqE�ɬ�����1!�D��,���u�]�:�<���됁^U�����8]t���'�����8�3OL��J�N#.�@]���+D�4�g�ܩ'<����(�Ju�UH|�.�+��ǡ6ܒ���GI��qԭѼ�:�*`��{`.P��	�s���c�O�̢�aۘd.Bb���<I�F"O��S�G���� !hE�1+�1� "OH�Q�ːN�]ه��2^��
$"O8l��(P4F=�sF���²�yb�ٛpf���� 8)����Q�˧�y��?`��R+�$�:��A�yR��=U�]����	�d�0���?�sE]�Z��ՙH>E��Ǒ�x���0:���a\�HR!�ԍA~E��Q�3+BE2�f�4%C��5E�(�qA���6
�y�ț�)	�|0���XV���,ԇ�p>Qu��2Sh0����oᰩ�')J/wϲٰ3��zd�6N*x��~�f��Y,�X��V f��k4���(O8��C&�\&�x�Qf�d��c̟�!��fJ)=�f��5��~tq���'k���.FH�S�Oj������q�\H��@�:'
Ҹ���X��Yz�O��j.�K��:<�#~��$�0�0d�	97���p�M^'D���L�����+�p=�A#��kKȘ#���Z:�M���պ<�I��$L8G�Q�e�5/�H��g~r�Y4,�F��c�5o�T}�@`� 8�~�B2D�� ��I<]����L7P��#Ă=n�0ƠM�0[|I�S�ݣ?Xೆ)?�g�Bu(�8�'-}*��E����M��v��D�S��=��m�B�NI�̥��l��ʧ#(���қp�̒�N B�t9��
G4�Yw�Al���O,x��>�X��!�ͭk]����F`�۱m�����w�P7)"~��� �D�$c�h�\T�V-Y���I�D�p&��!0�az�@�&M4�0�R�2pء�Ft�dCL3+*�	sg�B�r\����L�ui����ǀ�0��
H^2����
�P͸u"�ORŨUL�//�TIa�*Z���Ԡd�RH�81
���$��)�M?��	��� �MȎZZ�b$\Q��
�8uC��]@�ZpD��w���d�XJ�zPd��T@֠����d�U'�L����`�!�M�B�V!`�>I"��c���>��J\�`��eo��H�^�1O�������x +sF���錢>��T�!���PQ�4�%�.+~�I �F��2�m���U!P�y�����$	�"&���2�-}҃�eIT�+��[��}�b��vӄ�AI�+�2�:���	缽[P"OR��!j`�kD�z��B7WN#�� M�<1�.	-�q��'�|���Ѿa1�m����|���8�'��hQ!F�5Y������6�ȓ���*n� 
㥘h����ϻyI@�b���4%G�	�I.O�51%�ФgۘI�O\�����2�P��v��z�|@	�"O�ȱ!���(��a�+�7e$F�BC�>��֗l�F����OB4%����O����A�N�����^7z�'qJ� ���HI�d��){�rH�T��ȟܙ��7K��Сǎ���Ou�Kvd�� DmO\��K��t����,E�2���<�G)،hm9q� �+z���r��Ѱ����0<�%�WpJh�V��4/�J���A�M��lp�Z�a:��:���+ ��pa�O�>�F�)#@��Q���2*������)� J8S!h+v��`��� X�X�P�	��R����k]*	��,�`B0[!��X
�bW�̨l9ڴ�S��(^P!�R�yJ0��X�`^6��t������ n̺8���&!�"�h'�=# Ў���f��NГ/L�:Uc�5�!����������̱��!����N������} �0��~ c=�ɼA�t$�P�w���q��/CUL����P�e��l΂;�V�B�D�햌�Q�O�B���ӈ�)RD|q8q����0=��ʺeİdqG�?���d�^�'gn���
�`ȮT	��ć=����Fi����H�=o�cf�2����U�<�6�*�ESv$� �P І�kA4�y��5`Kzh�Hāo/$���D-�M�|�;*�\3�NҘ����!�Ĵ`�X�ȓ"J��qFB��0.��S�(�p�Dq	�D�c+�-r�;A�F�Q�K��?�a�X 3)���<Q_SP�2����a�5+J|䣕�'�PH���<^��{w����DC&(�|�	��6"N�	 �ŁjN0p��,c�`y3��' ܀�D�H"��z�I�4z������O6rX(�qɛh�N@;�j�k)�l��\!)��H�ba8�h�tB���"O��LT@��:�Ƌ�-�h�3�9�Z�P��Q�Rn���B�ȶ=� ��Nܧ�yw����`��U�
%U'T�I��yAۙS���1$c��AI���$���?)�NE>Nq#�/lOmчɀ�{"��S�^>`�b ��'c��C&h��
�em���Y�G�lm�DK%�]
�.C�Ɍwh)3,���l2G�>�0�3���'�(�B6�SN�\�ɊF����T)��B��PzF��c���B������+��Ǆ>�,M$�"~�K:��PC֧"�~��҆Ƕ$y>9�� 6���y�T�H�@�2Qd��/�d���$�O��X��}����r��h�ʃ�y��%\O4�!\'��@�kӧ�y��2iez�	��%N��ݻ��_��y"�Մ�8@*R+�2)���#� ��y2�( 8�	��Y�Wfxd2c�ظ�y2�
w�:,�u�	?/�4�B���y��o�Z��T�5���J��y�ܐ���Q韒p�8Lt���y��K�lڬI�ϫr��T�C��y�']�e���Sq	_$b+ !�"/�(�y\4蘨�`�2RF-s7D0�y�n]�g�>1[ӈD)W�J��1gW�y�IE2�Q ���Ht^0!��7D�$SR�Υ{Uh�z�·#g:dA�U�2D�����#9~ ӧ�"t�(W�/D��T΅('��-&��3�Ru!�-D��Q/߷_�=�w�C[A��3c(D��⢠A�&� p�"���,K&D���o��'d��Ŀݬ\�í&D�L`�+DC:A% C5wE��� A&D�4�!g$=LHS�B�!	��K��$D�t��ʔ	^��� I�,񮬀@�$D�P�1� �٘tc夘�)k���#D�t��$ʭW�̪G�
�	�m�D!D���v&���|$��A_&-NR'<D����I�(��6�$gWPŐ�� D�,a�N_X�"Y�RM�o�V�2D�,`�
˹*�"�a�(M��k1D�䊳� Ǫ���3�	�f�2D�$RFhB�+�����F�.���k.D��Bә|\D��#�H�q	/D��z��̮J7Jr���9��(T#.D���Z�FpQ�C�[z�9 �)D�p�K���5&ï7fX� 8D�������J���6Ht��g8D�`ZwNF"$s�L��An
��v�:D�pҀ�B�NEPb�ܒW��٫G(%D�H�'⒚p��Y�ڕS+��`�%D�� >l�a?;��tL���(ሆ"O��0�V/FR-���R/�F�`c"O^Q)�.�$�r� ���UL��"OxYZD��.O}�ʰ$� )И��"Ox�z!�T�M"XA���� �P!0"OR��6Lx7�L�w�S	S�PEb"O4	 ��#LL(�a/^�m����"Ofy��V2�޴hq���&�h�K�"O�Q�9Tў5�R���4z`�'���S5�ٳ+4a|����,�2L��o��2$�Y��=���ڡY�N$�C�O0���l�r:���fF��t"O����Ն�!Ћ�4PzB��
h&!��W�L�4"}��㓜m�����ءst�#�/�y�<����A��Ļ����m��ڕ����@K��Ͻ	:��
qQ>�q^L����5z��C�Ϋ!��T��*�X�׎P�_B�ġ	Ol�Q��L4��90e�Ba{�� .^�Й�D�5�0�:V���p=%�,J����!���M��+F5]v��[�Y�)�Ċj�<���^�+q�a���)k������d��N��'�S�K��I���))^|jFb/�$�v���!�d>D:�s���+�� ip�A�aF���9C8���'g��E�,O"��v��	@(vy���Gt�ѣ"OP�9Slإ��ջ�����P=���2��A��Ϙ�8]�L��	�%��%a�-�71Ǹ�h e�-����Ę��X������?)�C�s��p��ޥl^^q�f�`�<�b���� �c����p}���^�<���N����5[�,D+f���b�j�"`\�3W"ONAJס�
,ɐM`Պ�j8D��"O��@�� ��5�N n�]�r"O���,٧Q2�{��*\�Uɰ"OZ=j�ݲdN�(�ٝjb��b"O����M��X�p
�w�d�Z�"O�(È',QĈ0���$�$){�"O�I#� �n�@���d��"O�V�
@e�K����v��!��oI`�<�%A�mOn��b���  �AFb�<�!�� %�T��� 9&ϰ�ӗ�O\�<!�o�@��sE۶%��A"(F�<��P7?0Ds��Z0I>N��2�	H�<a"��[E���W��,�$�aG�F�<1c�BR���
�$ۯ36��c1͋C�<�P�B�wn�����^xѡ���<)c�^��	��@L�0���� Zo�<I̜L4l����܅��hS�<�U�Ҿ-8ntT�C<Q�� ��'P�<�������w8:�*�Vb�Z�<�`)A��\�����o��)����W�<)��G1 �ݨ�	�T��A���d�<�`J�MѸ�Ap/�]���w&�<A�i@�|�F�+��L ���V%t�<9&��6H���yq��Y}�QJ���_�<�7T���/��[�3W��a�<�WJ݅~�Nm���\�^P�M�@�V�<I1N٩��%X��U���Z�[L�<�g�̠E�@3��-r�l�r�M�<�$����I�rF�%&���RA�q�<т�j�	�%W;n���(�!��<[Z�cg�"|�$h��	>p�{����wID��7O�����ơA�  roݏ/Nb�	5"Oh��,1h��b���)|�p13��$�4^�����3�h�����4o��*�!Dzw���"Od�C��?ᨄ��/� d37���2c�U�C�
xy���q���D�LYX���%�`�l�K��6\��¢���#�)�|�X�`�ˆM����R��G�@�0�1�إذ=� T8��ܳ*��tK�L�~6M�Ti%�dL{<Y�t�~���Y��H�$	�F�~�C�J��7u���7g��u��i!�.�O��kת�JP�(�fY� \*ԓG⌆K��A�dE�~Bូb$h����'.e�dR��O��(���~�EO^��Y��'0����Om�'p=Kp'��.x�̓?�j�{�@��+H
����!s���9����B�N�ų&H\C?1b'�=|V���	!L�A�F
[�'�i��"n�j�mT�g��c)���v����6E���O�^���D0��P��вY��t2P���T,3��i�9�ӓ��`@V��vv~X�b��z<H ��'G0�(ǧ��/W���g�BE��N�hQ�d[�Oφ���@J����xQ�d�Y>�ɺTk��?Y�� ���(T�@%4$����l	9N'�h���Ap��Y*LƎ���B����p� $���w>��'��x ��o蒼чA�W�|E��K����ƟƟЂ�*8�jPҋ�0w}��0eǆ 'treJ���%�� #w'
Qt�I�_����\oH�p�\�m�Q�j'�ġ�'$��6Ń��pD�I�<�Y`�";`V1���[ nĢ<���0��T%�D��O��q��*v�"	ӓ;���ZI�,���E<ᰛ'���1�J�~�x,� D�Ņz�r,�P�ӏ9��V���u��ZFO��� a �N(<!a���d��R"(+��	5D�A� �[&ˠ�\�`Č)"h:�Ox-�=��O~�d��BI)t�V��1��!D��[�����$SvvA��B�D?����E�#P�E:�'�QQC!�)B�Y����~��M��d��1� 1��DEӍw����fT!��ũ�] �yR��m�8Q�Bw�
�(Ǟ.�yb+V�SJ�b�!Ϥh̜�䌑0�y���8x$d�Y�^+���� ���y"�D�"@�Ʌ��Zj�,a�@^��y"^^������_�4����yMO8��(��O�p�S�+���y"�M�w��������" i�J��yB%�6}�ɐ�Hǯs�ؕ���W6�y��L@��	#È�ai��2�)�!�yb@\A��r��E-\�|�����yb�:��`�_�нE�)�?��i�w,�i�M>E��ء"ܬ"UL��DÄ���!�DR�VT$x��L�B��@�2�����I-e^�*D���y��St������O12ṷ�C�p>��G^3�5�4��-N5����d�P��˟}kp��t��.I��~�`��~$0*ρ=�$l�b�/�(O�R �{.GO��?�,d�ʟ\�&h:{���B%I�&�0��r�'�©�Ln�S�O�N���h�l��"m�l�Q�\,XY�@��5J]�1�.��g�L#~��2@cI�%iĞ,��[;g��� ]��0�p=a�M��9
J���0HG�Ӭi���3p���8@�Qs��s8,Ѫ6�M�'9(ŚFO�>�pm�e�D{c�����
CP��B5�Rp8�H�SJ�7L�tic�`ƶ赋��W.�pQf��*�hD�� �9;���
P��ضC �pr�ӧ��8�̀���F�䐔`��R�Q�0
��d!��@\�"E $�ȌJb˧y �p�V�ܖol���+D0
ڲ=�'b�m��]���J���O�L���t�f���U�#��3�$<
0=x7�֛"RX�k��@��"~��@>��$o̤E!����g���I�{d2r.�	f�az)���8��F �����������>Mtj�!�a˟B�ب�����-x ݁�#�&7*�ׇ�'��Q���i'���C�"�O���c�>y|�Ku,�)�
�I�L	�$��l�� �V�|����Z?�擎�RF#E���{̇'Kc���tY�](t��ÇƸXc��$ٹ_-~��㧦�\
�%_&��w��4N�\X ��|��}� Ky�]�>񔁀?�,�>�$�V6<��9:��=P�Ɓ^�1O�5
p�F�����> ����/с���X#/*4#��	A�A� T,B�I�)BD�MLZ��+�G؀9�mJv$ x���)c(}�L�;�"i�#�FP��kv��2�x��eڗ�*��4BPc���Ж"O���`j�� I���eC�;O�F�:��
.��v�r�x�>�3�dՅn�|0p�IJr�``C�0"���P�x]!�E��_a��!��.M�}R��dP:��D��teA̙7j���@� !"Ć�	3a΀yCk����n��}87�6}�h<)�d}B�ɤN�n�JcBS#"!�3x�'
,6���d�8��\kH`���i@�Q���{�[�n�T+�\�v�!�#0�c���HHX�*B�]�0:��03h�`
�5�*0��I-}
� �5@Q	ܷ^/&9s�*�%���wO(q�IY,ZKY��W6?Б#(��1��ͪ��x�r}����;���𤊕A�T�CH�(�D䓡��`M�~��ؒ.\A�dR�l(T�3�
�t�<�;��F	zF.�ȖŊ1��8Yw�'���P�����7yhx���d�=��{�E��a��&ׯ3�����T�z�8�7F˴���fX3�y�,[�51���n	���G Z��~�I�5Y�D�g�<��rv�փ.۞�E�tmD�-�D�C6���c��ap���yb�8�}x� <e�h��ȍ�.�R��a \�2	�{VG�g��$>���D�R=p@^J��{��8c&�~"nX0< :3��=}lT�bS)��v��<���ȇ5����)0��88�+Os����Í:����$��Lų&�?ʓk���@aC�<����f�c�T���+^�< �W�U�9�X8z�(�5(݀g8D�c�d�R2�$*5,�T/<A��0wI�|	u�̠T��a*U"S�r�=��Q7�b>睄:+�+t�ثl*�i���ѱ(ƎC�ɸ`J��;��Yc���2Q�B�plH�;&�^91�)9v��,�<<[GF�����#��`��c�L���blU���إd&Nh*�C&|O�Mz��70hT��܃N��}���_%|-���@8 �D�]�?(�I��"�X�r��(>��x��ԇq�P��*Um�OP�RM Vv8 ɡ
�(猥xs�+��gq��E�I�>�j�P������C��!+4T��EĜ3@�l� ��2V�	���T�:ZJ�)#I�0�-kU�\!*6P����D>�x�ǆ[�s���b��K�ߟ�yR��@���}��p���?I��ls�����-lOl�b�+�'Hq��M��'�H���'�|�:���~�d�n�&\8�$�1#;]?|���L̑�RC�?C|�D�@�D7�:���I s�"�4��|��Йf�ӟG���KacR�@̇�UC�	\�JdjR��4{>$y��aV��e'$��H'�"~�YP�B��AIf�Ck�(:6���J�F�S��,O�싔J_#A���~*`qb0E?�O^�R�oս!1��D��!�|X��"O��+J�.X�VeJc��ل 3T*O���u.L�;JK�Y�씨�'e*I���X�H�x1�� ^�E��'s���͸4�QOP�I"���'�$b�����x0#L�BZY�'<,��K��GvX�W-\/^ؙ��'Pj��P 0n�X:tS�k8\��'CJ����Bt��+àڿW����'=|�p�$�Y���d�4Iۈ-�
�'�����eҶa�SD$FN��
�'�ڬ"mݘ@1�XP "�1(�L�	�'�ިҕ��	̆� o��4���	�'4�AiFD��b����*-���'�ج���|,0��F&	/O�B�'gDd*�D&D����4�h<@
�'>̙��g��{7"-�&	���P
�'��sUɊ�J�\!y���� Q�'�P4�f����UP�#٪	���
�':�-���2	>����&^8q�nDI�'���@Q58���C�E�@�;�'Un)�ZI"|��l�60��	�'�4�i�LE*�Խ� 8���'��q÷	�"H�u�+>O�=��'Q�`F-�D�J9���@7��-��y"��0����E�f�,a9�MU�Ș'�v(��てy�8��\<�$��'��4PÅ��ҁC3�%-� ]+
�'��(gG\9Z���S��<%I���
�'-���KC�BMC�J	�(�
�'v&x��إ	K���3aWz��
�'��mX�x�8��QNҰq
�'<t��aZJ\������y]l�	�'���	U�I"-|u�@�!hX���-+{���H�������������D�R�x� c�<�X�OJ  ����22HS	�g�? :<�`+8X�BN�5aj��2O 4y��E�*�&�Y��<E�d�6\e�5R�׺<�0 	� �*e�E��%.r��^���IW0,:��F�U9w ,2�<r[v�⇃oU^�x��g�T>]+d�X�X�tPۅ
ߛ~j����5B��'k����4�s��sӼ�y�/٥oe���ی$�c"O.<Z�Fڼ;~���tς�A�Rq[�"Ov�S�gS'"�rl1 @6,Q9v"O�`��Q2����E'�%	�6"O�\���}b0�XQ�x��2�"O���֮N�x�Z��GT/a��"O�"2���~�p32�� H�ф"O̕K���\���I�N���6"Op�j`O \�JET�nEld�"OF������ 5J���@(AE"O�����ˮ4�4�d
�J[��v"O����ސ�Ă�%f(��Ib"OT��ES�c��J��M/o	v,k�"O�!�2�;�2%�A�'�M#�"OD���^�~�E#� p� q*�"OӱH�B{�u�i֯Qr�L�"Op�1a�^��A��
Q�eX�A�u"O��P@֍)k8��F�R�qH�ɱ�"O�l�V��O�V���ב�<)`�"O�9K��E-p�L��)��Թ�e"O@�s���EZ`��q�[�q�n�"O�kA��t�"�p�	?B�(q*�"OH�c�,JmR��0�A�(�轳�"O�-�&�jf�i��H���"O8��"dڅ)0��*���
~��JP"OD�9d��3$l�V�\�?}"= "O�ԛ�C���03-��^���"O�%��"�x��黓╪�8)[�"O8��D��j-
��r���`ִ�u"O��0���O,�y��Ɋ͢衣"O��i6��1G�u��,ܓT��U �"O���䇮=~�P����$��p��"O����)lU"��vkY=�lm
�"O@1���ߵ#�P(3�I
@���z�"O`ғ̞G���I��B$�g�!�G�)V�)ZD�>�N9��V W�!�������S!����笓�Y�!��
�<TUJ'L�T2J�@��V?Y�!�dZ�oNN��񆏕�!���R*]!��F|= =����7�:�C�&%�!��!)�� ��+;���#�w[!�S!Y�\�G�TyD�d�<T!�D��"�x�4M�R_8���肕Xa!��@�h�{�`V;+i�H�!&��&Q!�D�"_P���B�![��Y�A%N=!�$��46&� �l.U� ��%֜<!�d�\8�W��Sn��PCF
�!�ĀP��dr1�ۥw�^|�eaUF�!�(+y�ٷ���I�v!A!�`�!�X a@�f�ˁ��A�D�A�hk!��F��8jW�0D��ذ��Z[!�䕖*���[�.
"S��(��[#\!��#N�6|�A2zj����	�!���qSj\Rp#м$��])$��*�!��U�s� �bq��3�t0ע۱S�!�d�
"L��DF/ڬ��d��as!�dR�+"� J�g�,���i֪Z�RM!�Ğ5@x~�b�Y�^=p�� +l!򄌘~�D!�F�'<��|2��X\!�$əV�ԉ�w��4�D�p̌,B�!��  ���[d*� �ŧ�Q���["O���H@0� ����?{�F�"O�ir3b$�Dus�f\�\ע,:0"O���F�"KU��!!�Ԯ�ιa�*O��!p�+A�Ё I0:$�ՠ�'�"T�gmv�����2NZ
�'�$���O�*�y���%[��y�'=���̌',��ɻ����p�#�'��93�
�M[r����ِI�"8��'�x%p���~�UC��(=1D���'I:)C���a�{�lW�Gx�I��'Kn	�(�1v =�rmвD���	�'��-��Ho?���dҕ'h܉��'\$�K��
o8�����4i2���'g����מ%Fθ2F�EFw��'�JDI�"�D�y��0.<ɂ�'��1j�L��|�Biީq��q�'M��y� �P섟?�l� �'��qaT�`�M[�/���t��'���c�(пh�� ���u��H�'�P} �(�#0[Fg#�5t�6���'N�D`� e��KG�H9s�����'��db�#GK��Q��]�"�BA�'װ��oR/l�v��ж?�PX
�'|
���H�2r��9#ՎR		 z�
�'�<t���Ţo�x�ħ�>{����'�(H��U�$A��O���'�n�c���P�����	s���c�'�h�!�Gۙjq�A� B"i+=��'1�a��z��1���K�f�@��'6����ՀT�P��\�)X�'�\-�w�B�9M��ڇ�)��iq�'�,�򗉋3"!�dSgJL%s,�P�'d�*Sȑ�Zd慰jM����9�'��
�텢P����e"+l���'qh0��j�8�N4��D�M�]�'pV�T)[a�P�`��[3�L���'�6�F�]2|ػ��vU⬳�'���s`�C!~l��(�jon�c�'o����H�}�eGK1^�I�'�@tr�L�k̖�!UB fH$��'L��J��
��<k�*��L�dq��';:D	���(*�8�âݏV��	�'�Z����5(��\R`�b�@�	�'����3&'?����3��[4|`+�'WHm�c��������S�ZH
�'<c6���x�:'`J��2	�'/lZU�K324�@v��@i�x�'-�� �C�	Z5��g��?bl�C�'�6�3_"�@hQ,ƺ{Ƞ�"OL$�֤�2 �m�	B�>Ls�"O���3��
"�ƽ(Ʃ 6l�� E"O�0�R!�		i"9*C.��2�X���"O�\*#D%0qq��f]�0!L��"O��gK�\���&ء�r���"OT8�e���P�`q��ˉr}H�(�"O�%C�&��dqx̋&  (Ml����"O��(ţ�;;7�DzTE3\T�q�"O���X�AՆк%�h��֮ĢoW!�D�4��U��o@*D�(tsvm��W�!�d����!7b��-ꤤ[`��	P�!�䕁6��@CjN?:�(H;���c�!򤜅QSH<�1���,i��ݎ�!�D݃R���֮����K�� D!�� �(ιy0ڹ.�6/�x�Җ"O�UY��^������3A��X1"O��b��Y`��݉3nSQ�,��c"O�|:�T.C��|��l�5^��EZq"O� S��/��h&�"���a�"O����ꓸ,*̠%�ώ)k�I�"Ob�����B%Ēm�� ӂ���h�!�DL�.z�-�V�M6ܦDS�dC'�!�đy���H`�V(QȘ�� A&�!���k׺�@bӽ]�&UB�`���!�DǛf��3��@�DB���SI;�!�D�,�� �գb92�9�(\_�!�$؅�@i���+H������!���)��(��a��>3��SC	��!�Ą�>�u�N�Yt�ש]�!�Y%z��A�/>xX�"党�\�!��v-����	i��"��w�!�$�TD�g��#D�:d�u���!�Ĝ�-�Ν��ِ�xK�Αz!�$�4�m�&�݈0�(�D�W�.!���	�^ ��M[6Q�)z G��7v!��X�&��r����j�J��2%
"f!�$�w�d�vNh��2�#ԍXd!�յ� ��NѻH�( �e��XP!���$B�˗ N2~���F��QH!�Ȍ45n�+פ
S�贘t�
�D!���*����
b��T���Q�fK!���L��Aq4�N4>0Q�@�s@!򄋰r�n����`��A� f3!��KO�<XS�K�3/�л�K�!���E�)����r�b����{�!�ܾ,�b�dMN;O�l�끦 n!����Ե��[n��8�Ӌo`!�Ğ�$�\�wc |�3��)$\!�uј��b��c��(��V_N!�Շ\���Ҡ�Y�����0)6!�Lq:^$#��_  ju{���h�!�D\�<�r�b#�ŰV����Vf!�$V4	>^�KF%��EoDtR�͋C�!��-p�Uӡ�_0STD�����>{�!���8*w̌�Ǫ��fN��cӬ�F	!�D%^�%9�me֬�RL�!�B�l[P�^?(�(�/��C�!��Ưg�T�&�nG,Ls�(O'j�!��X�b� ���ܞ#;�)s�g�� �!��y�TX#R��7:2t
��@�pT!�
�a�ʈ��b�O6daʓ��(=!�dK�H��H�-�����8"�!�H���Y�Z&�<� 1MM$�!�䅵4�-�l��)5L�I6KJ�G�!���W�րDaзE�8�R�	4eT!�DH3��R��^�4���ȃz!�[q44�1%��,綨rӇ�Mb!�d\)+��p�K	�o������;2!��9|�>��������A��=!�ƈ"���S��B�d���;d!��c�Pa��G�O�����˦0!�DÃ<6�1�tɘ�E���4,B/X!�D�am&LhaH��'�J�m�|W!�'O�J�F�ѲXx��V�ޡ]3!��:[>��`�/@�H�`}y�
�?�!�Y�0��d@��H 	��̀�I
�!�G�EnT��bY�[��42�H���!�d��a��i�:���mOu�!�� �E��C�B,���#�����"O�D+��&%Wl$��e�0W���c"Oֈ	��! �y�B�ĸsZ@频"Odq
��?�X�8��чOR p�"O����OL7|�=���M�b�c�"O&Yc$SQ��!��y�@��"O�ph��5aW� �N� h-��"O�0��^����J6��tp�ٙP"O��: @ɧ~��¢!�)U	��'Xh���=q?V�`�M"!:�4C�'x��Pt�I�&Nr�G$�OWL���'��8���#Lй��Gq �	��'�:'�9�ih����W�D�"�'�|X���59� �'�I5l�'(��Jw)Hd
A:V�],�:y0�'��h;�� A�0E2V�F7r�B,��'���8�ӺC��@�/H�h��T�ʓe�.tڕg\�3t��8�+[� ��ͅȓ
��A�G��;DVTaЧɩt�䌅ȓB��<�JѪpp�W���?��8�ȓD%�!  @�?�   �  w  �    &  �.  �5  �;  &B  hH  �N  �T  .[  oa  �g  �m  9t  |z  ��  ��  A�  ��  ș  
�  M�  ��  S�  ;�  @�  ,�  p�  ��  C�  ��  $�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��~~�:ٶ񩗫��Ɍ=[C�ՙ�y�Kɮ�f,ȳa;%Q ������y��^Q��a�:��Z�	��y�号i؄�կ3H�ܲpd��y�K�[I,���K�&T����B��y�~�N��r�@���Lq���yB(��1 �@��ޚ��M�����y2a�B��%2e��*P�#6�ܩ�y�C�?դ�C�f	�{V.��&�0�y��@W�8`�۱r����fô�y�#(k�P��8=�4�R'�	�yrhL�:AZ�+V ��&������J��yB��KA$��A��[Wb����з��9�a|�Tc�I�ҭֽf8m��c��y�7<�0�8�/��Y��'E��y ��J�R���?E����\��yB�ҳ!�ccK��#K* ��C���y�U,>X\г�gòe�����`Ƃ�HO���Ӄy�\�&��u��!꧎�h!�DE,CtY��.���Px����S�
O���,R	z]�a���&&�H�דnqOR͋�J�?1Zrxdgu~��b"O@p"�c�*v-P��]�q��)R�"O� \#@�D!#�h��(J7/�@���"Ol����T:;�&��Qf�}�m T�$7LO�����*Lsj}��J�?Y�%��"O24�nH;	�v88Q���S��81�"O��D�\ v�2R2j��|���q��'���E��,.@B� T�9W�����'D��	cGW&<��g�7mV�Ё�%D�@#U�^!>D���
��x�`��`%D��Q����H�<���\4�z�	�i(@�ay��R��b�r$�0"��$b�-�+�yB�([kj�pǂ�^�L�2l���?��'o��9�D
:�e�ϕ�U,��'���K�O|�^��4 �/X�@�'+�����_'S���!��9�8�'��d����C3v|+FO	)d���
�'n��'�ޫfn2|:rj�)�z%+	�'X��P���c:l%�R	j�a����ą�1���@Kļ� ���<$!��I�^�Je�ԐQh�)�nۗL#ў����5v������ن��E�zB�	�*�L5���*���0���B�	)q'
�sá�V:(��`�>C�2zŲ�J�jŦ��!���RC��G8��@v���"Z�q�E̩8�.B��1NQ*����(a�J��C��C�<B�	���Y�կ��h�<�"�ɷ�=�	�'A�~�G%�9�:�o�~B<��ȓJ�	awL)Z�$���
��&�ȓN�l��Fg�i޺(���Y&Ỳ���1F5K4I���rc�:p`��	ꦥDx��I�r�a�1�O}X��ǻb�8C��80�H!�H�!�
�c��1�dO�����9t���q�$�c$�)��ÞCw�zR�>��'�f�s`�\�.Zf �1m�.i�EB�'s��D�_��j�� 6��s�i�	G{Zw���;fE/oY�8¤�)}���'��uH��W=M��uH4_>/���'R�r7.=yf�Ƀ@Ű*'*��ߓ��'�b�x&
��#�m�RD�
)8���'�y!�B/"t�$��9���aǓ�HO�idk6g	@�B%��>w]�eA��i.��Das�3�-�%/˼Y�i;i~�Oy����)�N���ʇ3�ja��ՙLy!�Z�L(rO.��!q�c�P!��\4G���q�?r���aÅ?<��~���u�ۨ`�S�Ő>g8�kd"O�Y+���ěg�ԷSb�a��'���,ѵ/�	px����g��9�B�4C0D�ȣrŎ��j� F@���3�*�O&�=E�d�ԍx�l�RćO�Z^59��<�!�D��ք8+�J�'Uk�1���-�!�-Q�0�!�V?hh����ϖ�E�!��O�	!� ��O�1V�#���1 "O`���^��I��j��[b4��"O�P�1b9(�4�&�B7)-Ɲв"OvI8�˕31*��5�Ұ,R�Zt"OT� �J0S�IqM� >�x
"O8���k�hA�Ƣ�+.@�����1lO>i:6쟮��aѣ��$+#�3�"O���%!V�HB��J!�]mAB��&"O<D�oĬ$l!BD� t3@L[�"O�ͣ�+��k�܄��ɃǦ5P�"Oxq°,O�hĺ5ٵ��QJ�P㳐|��)�Ӿ ��8�U	P&O�i�����C�)� �"u�Qw���awЄC+^��"O����݋ ����BA�2!�U�2"O���5�1�6Ɂ@BO�j@!"OD�X��V{T Y9��_I�:�h"O����+QQ��[q��Z;���c"O&}J� ��Dj1і)':$ +��1�ŞE_�	딢�A>�Y��C�����T|k� ���V�x���T�z͆�Ew��C���+�<8g�id5��(� �+aK4G��e@�%��3�A�ȓQ�NhI��@�S��<�����7K�l��`�� B���$� pI
�I���_>���/�>h��)��9�Y�Ԏ�>Z{|�ȓ#V2����dD���Qb���ȓ1^&h�'�]aج�C-�I��Q��b,���C҉YU���p&�>!�@���&��@qA���E*E��:s�h�I�'��m�Pa�*Ɛx34FǔV��e	�'��8"��H� ��T�0�E�[Q�|A�'6v�k��W�la���j���'@�@� KJzta�d�;L�z�`�'��uh���)RqX�KI�<��u���D(<O��p�h�_L��a��Xw���"OιV�N*P�,��.I�p]Ш�W"O��$i�#;,���JL���a"O��Q�)7>��p) P��"O����I~��*��(~�h4"O��A�I� !�|�'�#�Y"�"O( 1�
�U�d���m�%+�2���"O�H�Ǝ�y���ǩ�6A�"OT����5~%0�j҉\v�@X�"OF�(���<u�X5:,�hQ"Oجk���[G�a�T���^ ���"OZ�� ���_�x������"O�)�abR4o�n��"�)��)�6"O�0���}������Y)5�!�u"O�q*�猥bD�]@�[0
E<x�%"Op����u�5��熍E&��9�"O�"4 ��L�p�p�� b��a�"O�@�� ��	5��
 �4Y"O�� �Ȓ�4r���!�K�O����"O,9#�_GR�4�"d��P��2�"OƉ
7 �3{�j��`ʧ|�^`��"O�8�jۈ]�ȍ�p��s�;�"O�IR�ֶy��x����-G�,yv"O�`	��.�(x9�)iغ���"OʍIT��a/D��GH=~Ϟ�9"Od��V�J�S��3���D�B�"O�x���C;(:(� ���pg"Ob&1�����?5k���sh�8�!�$ߔd�p�3��u��b� '!��Tؖ����D<��ݧ!�����zpL�M��c��!�D_06�Z���k�Y~t0�^/I�!�D˗I�9b�N��J������#}!��#Ъxi��v+�%JS��wT!�d�	��	�E�c�ey�'�k�!�׻NV���H�^�X{'GU�=!�S���D���>H(�F�5e)!�d �^�
Q@�f��]��DA�d�(!�/����$L�A>�@�$@;]�!�$�3.>�C�XqD�wd�r�!�)!j��`���9 �3�B߿'!�D�EK0�`�D
&�����Ms�!�� �u�$�E��0�� ~r��!�"O��J#:�~��f$<W0["O:���,K�ΉA�% M�i�"O���E	W�iˬTR�dBD4@a��"Oh�����EfTk��R2L�`t�'��џ���ݟL�	ݟ,�Iʟ�; UR�s/�l
����9���I����I���Iʟ��	꟤�Iٟ����{�h�I�M�v�:��Ϛ%-L�������៼��͟�����	؟���8	Ǵ@0V���jq�vm�K��I��ß�����I՟(�I͟(��`�I�X߈��挑1$�ht*�d�������ß�����|�I��(�	쟬�	ԟ��I�h���"��@��=xԪ��0�ި�I��	ş�I۟��	ßd�	ҟ���)�����C��
����t��h��֟ �	ןt�Iןx���D���@�IS�xS��t~f�ۂ���j��Ɵ�������IПx�I���	��0�I~�rq��̐D�	��`�������|�I��4������	�������<�I�(w.y����D�ٖ�������I�����ן��	ߟ�	̟H�Iޟ��Ƀk�Tq���A�,��ƞ�RLm�������ǟ��	ן��IٟH�	۟D�I;�,5s��L�xa�7���������\����<�I۟\�	ן8�	����	�"�����I
�(�s��"׸�������Iܟ<��ޟl�������4�?��R����^��-9e�P�J�~@2U�D��Uy���O�HmھO_]k��0�r�TG<V��XB�1?a�i��O�9O��$�f����_ H `Z�˫i��d�O�Ԑ��`�����#��O�L%P��Yv�����
) ��j�y�'!��r�O�f��T+�#Z�q8g��)iY��dl��4"r�$9����Mϻ+
�|���=7aj�*�nO9+�:e����?ٛ'��)�?P�mZ�<�@��Z:��Ӷ��+FL<0EL�<ɝ'������hO�)�O�T@��� V6`��eiۉ�4pr>O����(P��ƹ˘'�����Ė�h�R�୑v���x}��'��:O��'�#�m��]�1YŅ�?2��'��-�$Vgd$@����� @��'�&�8�IŁ��]�B�\�Dt��Z��'���9OXu��ؿoh�간�+�B�cd>O��n�0F��QΛ��4�0���n	8DFL�`E� Wx
`6=O���O0�DO1�6/?��O���)� ���ӇJ��rWdl�����]Z<Ԇȓl�T��҈E�����0��M����D��BFU��	U	^:�%i��Mfa24�tdX�Z�ȕ@s�R���� פF�Ts�UI�[.�Bũ�J	'���2��>Q��J��ְ6�j��!K0� Yr�̇�ND}��.U�ܱ���(}��
�Ӻ"�:uQ�H�;NR�G�а�|�bF	�*�����DN��r���1b���ٓ��Skͻ���� �PX�!��/I>��WkJ�b5��=1f�ub�'��;�m�uI�3-N];5��,��`�Dg��Z��p��aѾE�B�ʏ,)A q��Cŕ9�BA���~�3Q��V|9�3c��Aw̄:�j F��-���p��b�d���.��T)�H��q�T�AD���"��Fώ]u��Y6D�HR�'HR�'�V�'�?QC��{L\m�A�+a�������������t$<jUo�k� ��'�Q�,�p�G�F9� 4'ȑ�,Ȋ�"H)?��t���2D ���5(GP�ӳ*=H���{*�aqn` c��y��⃕5��ǆ��~�L�n�?˓�?�)O��p���?�X������B�<��H�X�Ȑ���.>p��8v���pq��pD�쟐�'�T���q�Aa�DCT���h�� 7i���(�hOԟ��	ݟ0�I�r~�h�IʟP̧J� �)aUk��j��$�j,���4�%���1pz���|,����ƫP�|����|���s*�,�RmC$C������,� �`�k;ʓ��}��ܟ� v�ڂk�����`D H��ջU�8D��d��8?����
\x�"ae*O��=Ѵc�3`(� �vCVG��*C���<�q�i��'9�5���zӸ���O�ʧ�0�:��:�ڈp��/!��]y��*�?���?��k֎5 f�P�%K�I�O�b�	��D�<��qP,�M{`�x���N��bY1H��p�ʛ���$B��h��A9�L����Y�EQ��x�a�O¢}�#�S5/Of�b�AY��đ!���<)�\q��!UJӾB�	ȓ���'�ў擞��&�� � EgI@�+^�R�Dh�<Iߓd�4$�� �7AH��4,��Z"��ȓ|MZ,�m_3Q�q�q�E/JʈT��r�(p�)ф;��|���.�ε�ȓ N t�Ɛ<}����Q��J)X�c�gO�Y�ʰ�7]x�y��G�  ���A��lIC+	+9!Z��ȓN�H��d�?, !���*ɼՅȓ-�(���k��Cf�%r�`ۨV�^���S�? �$�7)�!��a��L�d��"O�lX�$RuP�i���*��1{5"O��B&T�i��q*R��8!}��;�"O��PR"+X]UHV�L�i�����"O��b#V�`�����e��M�����"O��H��QrLx!�eU�
3`Ѻ�"O�ss��
��MR���� �Ã"Ox�і��.;U-KF@]1��Q�"O�� �ĕ#(�z�lW�C����"O��`���<iР�!,��-� %i`"O�8�T���;��Ă��ƠM�^��R"O>5Yq�ܸ;q����
NV̬ �2"O$As��Y�%k������t��C"O\5(% '��y*#+Y�x�&"OB�S
7Z44K�陹L�ȹ�"O����4T���(0�B�!NH�2"O�a�-#Ɗp����8CC��S"O��AP��=.�8���V�T<8�7"O�B$�L;$����+�e�X)�"O��� ,r��Ԫ�D��'�<��"OX��OR)2�1A���6a�4�{""OB٣��Pr ��2 ��<�����' Q�t����-�|�5��`1�tH0�3D��*�MN�5Ժ�3��ڇB2�8z�ǳ<��ǘ#+��OQ>I"wk�f�Z�7�M�mĮ�p5�4D�H�p������P�/[-y�I�N4�dO�X��1��'��I��2K2��J�@��%��8��,� �#ņ�tN,�JA�ē�^�p ��
&���J��R�T$L=��ɔn���Q�)�ot��Fa�?�P">��%�:~J>��慞]Q(���Z?M��^����9�<���!D�Lt�Ѳ{���j���$6�T���+`�,��cٌV*�L`A�=Mp�Ӏ5��ܓ�`��v)���Q��5y�<B�I8u0d�Ly|X��/t�F�WS�<@��O��@���@�d4FxR
Q<0I*����S�s�ҸJ�m˭��>I�eۍ%�'nډ?:f\{0��0�P��7��3Kb����k֕G��`	�� 1�1�]E"i�6l�&y7N�EzrJ�.�Ț��b�|2i���M�' =�C%G @"Ʃ	#l�!�&���p�I	�`Q��9f��6TM��m#p"(�$Z�qG,ڂ�Y�q��6�s�!X�l�&G�D8���F1��l+D�H�b+���sT��>�:��6h�h6���e�E���נ��(��g�'F�y���D��p�ǂ�I&���	�S�v�2��K$y,�X�ڱ4F,�J�T�=Q��j�%~�Ig�'��@B4b��D���J%���m�l�S���O2F-�� �)��%�M�d剤MQ�MӢX�P���5FD��y���<2Z�U�� D<z��y5M�;�y��M�x�Be§oI�ST���!�' mX����=K��ぉ�huF��ȓ7H��&�+_��d)�əw�x��\� "��G�l�68���^���ቅ\���;ՃMWbh#!�).��Ą�@,�0�-�E/�M��A� -RT�6�N�f��R�
�${U��	�Rx�q��>cL��A�6NW #>aV�N�T�Q�o�� 	�*���� Θ}�	xᮞ
X�F��T"Or��0σ�;�QP��I�4������'s<���%x��JWR�"~�w�o�D��]�
��$3�A �y2�H�(��ʔ	I�2�Z��ɷ����&LI����vξ��ʍ^�tD�𩔭u���u���^Qa}��c=�A�ݴt��|b%$0n��!.��$��ȓ;��q�@e�&��ԥQ_u�Gz"�ȽJ���F����# =�Dz���z�6ڥ�J��y�'^ZG����h�4w� �`V�S��M�D�3������6�
�h�MjV�7q�
M���ٟ�yRNø<���� ֩1�Ic�L����G0N���	�p�.���˛l�i�M�5(�����
X�Pe�L�$�;ֆT�. �d��!F���]��@��0#b<!�,_ B��%Gz�'��n�d"��� �aT�J�<�� !�\�m�*X�"O����'�9a����J����k�i��e:�(\�8�ɧ����@�D ܥK��2�
�A��G�yr�
�p!c���ki��A�LL����H����)LO ��S暍�dŞO���
�'�l�iJ���@�7E�b��֏��1m���χ�;���'�9i���W�di��FD>e�Pu��O����ŝh~�A.$&^"|"��"D�#�`+��͖q�<�"�(n���P��L����
�n}2��2\�d(�E���T?c�tSQi�O���KV�BY.u� d:�tQUaڒZ�<m�D �'ii4�cO_�iN-��O�i���^��d�cʅ�1I �z�R	V�x��-O�K!�ky�O���L��t�Z�S�(�q����	��� S��Z�<�4�^	ZFuȃ�M %I�+W��S~�� ʒ�;�hP��S�h�$eh�F

W�0b����?BzB�I���1vă>+�)9�!(l�d�c��XK�@�	�? ��'�@`�O���cj�hh%jE�+�܌j	�'2��-�/�����H\�@�=i��W�M��]���Lγ�MkD+Jj��}�E�W�HL0G�	?�n����+�0<1Aj���i��M��ݹ gD `~�)��+���K��ȽK�F ��}8�E)I9:@h��K^�6琴��+.?�"������ �����>9��]5��I��z!t5rU��l�8�D$�=�!�Ĝ<I<����ǆ5HV	ʁ�<\�ɑ���h�lY�(O�q3�S�dh��\8p1���^���gD���Hb�%�v�U�'#j��q�_�1G�%3e��?_��Q�$�ݶ Q�6���<���J��,����.�	#��0�u�Ͳ��TA��O�3h�#��4�KJ0����8���"�L0��4��yc�o��
.�K`��`���a奌vzM���X�\[v*��O��dI4�.z�@4��>�b/[�	|p�dЀI�,9�G�GyB��<�'0�p�1�X����A���^|����A2EM)r���aBz��dC�T��'t��˚��� ~�&u��cЋ�7W�*l��×VL��h�j�s؟�z¨	/̸*dB�v�2@����K k�i�DG&�ybP�2-�ɔbm��:��Ζ����OҪ=����G#�]��ez 8OV�[���H�ddЇ,�v0��G9�X���H�����>2~a|���kD�R�!<n	�Eۖj�#�����O��p͓�v�9O��I P����F�(��Lڲg!�dqF�hȴ���A�v�
F�X�[�v�c���<�dǉ �Ի���x�wQ ���&U�%���NR:Ȳ��y؟ 3�	�٪A�
"�-R���2�bH����y"*-�	�k�x#<yf��=�@*vd��1���{�'����B�c��y*2����i�O���9���N�$�����Z���),���!a��-�d
S�ȋ��+Bx���e�Q�&LN�=\�� �s�����R��0��	Qt���Z!��
*�	*��G�y���-�gͮ�P�ȏ�<�Ӣ�oQ��xҔ��}b/c�~�C�&�� ������?�b�iF��Bq��dЦ����I8���@�Z
T'�XCe�jX����(��"B`�C�Z�_Rf�r�,9lO�@i�Cڌ����	�t��HǛx<�#�-��jC�)�X�x�@�=
ڣF��O��*ǪE	KҔ"~z��A"JՈ��D�N��CW`Wl�<�+fU�7Y���T�p�<B@bR-�X�	r��~�+[.*$�U0򧅗7eTy�����y2E��m1��	��H����J�gX��M�%V|a��2�'3>���D�=����ǝ�[�k
�1๱r�5��&�"�q���/�������) ;!�D�s�|��b�+C:��t��"1�O���D,�ef�"~�Ņ��2\xqG�
c ��v/�p�<�mM�J�fxb��ŀ5�0�B�N�զ�QA�,�ا���#��2z�(c��X�N)��a�T&�yB Ѿ��1j�@�-���
b�����A�h�m��I	(?�i��	Q-d���F�L14��D��i�a���gᏵs�d�I�DK�E�V���(v�B���;�R�p�RZ�*4GzR�	-t{�"~B�.74�64��eJq�7dZ�<� ���GK��5��xx%�n$���ixh��
�n�S��M�Ĉ/�z�+�b�I����"i�{�<�
��v�f���p���j#�P}2��x�p���-��r���sE�p(�S�&�a��	���(��)r��1 �6O�iq
O�Ƀ�"OD�1%������)�#U������ɥ�r���2$��8���[�f��t��m�B�ɦ,�,I��$Q;E�D����84�&7M�I1%�>E��4=�ٹ�GZ6Y�����a���	e
�b�זN�bЛ��I�˒��'6u��.�O�l���ۼ:(�LwFÁ\��j�'9����&r�Lڣ;n�"��iv �h��&D�`W�Y�$�J!0��]�M�l���1ғ}M��(��Ӣ1����0�?{w��Y�C��M�C�	�3k�tE�a�x�{Щ�/i�7��]U.��>E�ܴV��91@l����:f���6�,l�ȓ43�щ.�N�<��&�ai�'ڸ��
�Z-��[��_k��A�� ����ȓ*�u�R%�-HQ��3����f�z]PQ�Z#f�ThD�������h�����6
7�}Z�C�+�.��ȓ�ܽ��bV�j�DPJҫ�BɇȓrO4i�q�N�A�����C�p?��ȓj.�A�$� ){v��ѶO�O��=�ȓ�9f�H��T�	u���,"��ȓ�6���$es�ЙC��'"�0�ȓ��t�qB(/�Py�
�<n�LQ��"�4P�T�ռVZȘx��&�L��j>��6	Ia���3�ޕy��مȓ\᪨��I\dxܛ1�DV�r���A�J<˒�XjE�rg� �|@��"��U���@Ej�ش�HȈ��ȓWEm��iZ�f���BbA.-��ȓ䈰�*��JNjiR��t5Ft�ȓ��A@,��)��	��W�6Մȓ����v#�>G�`�Yq�϶c�)�ȓb���4�V2A���!"0�:\��p Hg�ݸRp M)�`��;��q�ȓ1N��hWh�f�� U�����FV���4*Fy���Q�&�T��r�A�v(�?H��f+W9����&��2$4#q#G�54�|��*	0jb��<RzMbE��p4�$������f�0?���LPp�H���_D����
*S�qX�Ia��Յ�;0q�G�)<��-W����ȓN�t�h�f�?9>���e�	�]L��0���2��-B�i#�G.�P	��H𺱸��ZOZd8ۆ#�:�@���[ҁ��̕�OM��R��Y�^#�U�ȓ@a�fJ TM��oY�\�00��n�$)ӥDi�l� T şo�&e��2�����I�B�Ly�EEHE��L�ȓ^�)���,u %MZ� ���ȓ�� ������)b��5Rp��lȚB�RX�4M�Q�ݪ_ȄȓT�Lᅁ
fh����C��5N`������ZF��T2)â�S���0�ȓd:���E�-��Ay�������ȓ4�Bu�ǉ9 ��\#B$��-j����S��pI��\2B��q�$\ 8DN��ȓPT���5v�:�kWJS?�ޜ��7sD�x'dC?p
mC/�N��8�ȓ,�2m���}�S!tJp��S�? N�(��lpꁋ�]qlI3&"O���Gњ+�`b�WW��j�"O"=h6K�S�\���T2C�2�0"O.��ܘ>�l�Y3�1k�2tP"O�͂��� y㸘0Rn����Ёt"O�1%�2"�­;�J g\��"Oh��힌'�R�C�`K-:Q�8��"OX	v�ӥ-�����6>�܀w"OF%�II�H�dQtM�X��d�"O��qC��5��I��+�?:����"O4��ĥ7$�-�EKаI|@��"O�ah�/�7C����t�H9Fw���"O�Zu$Һ{�Ƽr�	$��-Pf"O��P�&�?f<������3�j�#"Ov���7d�
��ʹ�21�F"O`H��g!G�H�+t�J.k�:<;�"O�dc�I��i�daR/N-,-|t	�"O����0Ql���.�v����"Ofl3%n+Et<�J�,�@4�q"O��D��tf��ن��V��`��"O�q�jQ��"d+��)\P�PG"O��h% �"�J����%m[���d"Oα ����� U(��-E�P�"O�����	c�h�� 
�!���"OR=q�,��6�2�IU
���"Op�rWn��ƌ��Ǔ�(`�"O�@���֬ݱg_�@�"OJA�k̤��4���_�t�ؼ#&"O^�`� �1�1 ��%�P�Q�"O X�Śf��@"Q���t9��"O�qˢ��
\`H��T�_�Q�"O���W�-���hWf�?��|
�"O��1���X�4��dX	o�~�K�"O��C�d�U�Td��"��G��\��"O4k6�G*a��3l��.�h���"O�щ�,\�hᴹ�)ϨF�8"Ov�R�j1,�Jy�6�Ʌ&hl]JE"O�mq�G�x��Hv��S5N�b"O�1d"v:����#�u"O��C�� �Z̈�ktaٳQ2��@t"O� �agT8s�͉�n��'�aQr"Oh�@�T= ��h���*0��}C@"Oڡ��L�
��92�g�?x\K�"O���ڱz+�)�� ��J�"Od[Ʉ ��{E��C�D嫅"O�K�]�0��J��F�~􀊲"O�ȷCH>'h��Z��\ t(+�"O.(���0b�e��=2m���"O�Uȥ�͏3 *��셂U��HX�"OJ��� �%��k75��� �"O�H�V��$�P�l���@�p"O`��!Z���� �*�,���d"O$A1aQ55��7��Gf(�2 "O����D�y���"�OɃ3L1�S"O�kV��3lpZ,R5[�s1,�Hd"O���CǞ7m��H��, �p�G"O>]ZF
0�zhp�i�07D�"O�Qу��Lms�NXK:�a�"O8ЃT���3	ڹYv.B
9H��'���F?26�mx�/�<�j]J�n z�!�D�DJ��PKܿzȮi� ͂��!�7Y�z�)��#3���a�,\�[n!���$qD��G�V�6~���@Ԣ?�!�d�2)�ʹIB	�8
C*�3B���!��  �H@-�#f�4���(n��"O�1��I)4�y�ٛk �M(W"O�<��Y�HJk$%ƍB戙#"O
0'�@�bY]����3"uA�"O��T�*G|	hG�}#�}��"O���(^�TC��d��)���`f"O$%f��&�����0�R��2"O�����a�	�L�$~9b�"O�a�6��i{�� ��_�9*�9�"O��IQ�G'Or�
�Hfe�7"O,� e�K�d�I 8�9��"OzI{��ѐQ�JAI,A�"O�1kV&�b�:�C��X7X~��w"OF!�W*��+
v���E�z%R�"O�P93
(e���!���n꺑1�"O�ux'ΟQ]��0�\X�^L:E"OV�ꒆR�hA��3�+L*4�V%�"O��U�>M�m�f��<5�f�C"OR��j��}Xs���č�"O��8W�R�&�p,�1�s��9�"O����AH�E��y@!\�_
���"O�$(�EP��~��I�g<!Z�"OY�Rœ,SL��	�#ʞ�nZ�"O�U�À��5pt2F~w�]c"O��P���,4.�D��?�~�!F"O��� �F�  ���㋹l���a�"ON��T(�
X/v�K�l<�~��"O�񄍉$`�����jI�oR���"Oj�8e$;�ThBT1��0"O6�a��_���c�F�:�X"O��+f��]s����E����jt"O�ЋC!�~��B��ڑ�L�`R"O`��"�o^dՈ�&Աq�ƵB3"O�.ѨT���Q�-�=أ"On�sDƓM 	�5o�����C�"O~�����;CV���߳[�,8q�"O���EkH�f�����"	�����"O�L���)���)����Ԩb�"O�(�U�Uv-_��R�A�/�F�'>�?];���/����5��	4r�(�t� D��%���9��N<!x���=D��T��fffmQ���'_�ӱK8D�ĳ f^�=���"�nA�5X(��8D� ��F.yD��p!JM�N�4�� 6D����g��K�<�0���!]eJ]���6D���B�J'\�,%x���:V�"ꃫ6D�Ѓ��R8RX",�A䟁:�
5D�d�q��=hGl��.\*%-ܮ��C��%cE���戋hL������:��C�ɚ,�x��4� �i�ެ��gU�Nu�B�,m�#�	�(
�<�¬��1�B�Ƀ:j\ȹ�a�L�p�ҦR�!��C�	�Z%�����L������C8��C�ɜ+�4��r ^�s�M!���B�I�Ah���ca.˦L�tn�65�B�	�d�ԘP!A�0i�����c��B�	@�
	����xn��HYA��B�	?<m|,H�2lyBu�eʋ g�B�	�a���R��NQ�׈�*5*B��(6�Z ���E�K?�)A�=-��#>����#h��{�
j�����$�	[�!�U�d�q"��.P�����/�!�$�R�`�1U�ʧg��5�@�X[!��s� �[��H����0�vH!�� ��˰��l �(�zDت�"O�)�p.~���G�iF�]:&"O8K"l�V�DIQ�c�"OHp��)��@��� D�?6Mؔ�"Od��a"߁'mC�#@J�	
�"O"���EE&!5n����F�]I�uy!"O�	��"ΰWIV`��Eqކ��S"O<��6�{��@�Ef"jݞE(�"O�Y��	�\�^|z�E��<�P u"O�Y�M�4'K¢%�JQ��H��y �"6x�5��'F4������yrc�@��i(��@@RK�Ҵ�yLP�,q��S��߀8��`�$��y������*U�X����y���r�dx�kHS������ׯ�y�b�:��D�#�کD��-BgCY'�y�+J0����!L�Q���17�C#�yr`g,t	���rdd����y�k��^��YF�:d��H#F��y�F}�](�
�Ym�a��d��y��-t.�dR�k�$O�,���7�yb�ӆ.T���"M���k��ԛ�y"�XM�����I���1M\;�y"��?#u �؅�F�@��d��y�.�=:�x�i�¹j���I����y.�>c
.�1�H��R��]k��A��y�&*�ʴ��QZ���R�^�y�L['?K�pi��4JW������y��j�.e�u��A�n�XI$�y�dԔ���v�P�9p��r���y��^��3%�-DBP"P�L�y�%�4y�����v�~�j��C��y	^=r*�1��e�>���n !�yöF�И8�՗.c P#�(Z*�y�l��XB�E*;��ŒbhF$�y�+�F_��Dë.�L,�aM���y��O��}� & �`!��0�y�-�(:�M�������b��y��/��-�t.�
��x�h5�y�m�U`|XSrI�|Y�=;��?�y�搠*1����F��g���Œ��yB�S�l����*^7֜��^��yb���4�I� �L�(�d��y��\F�pǠ�|�L�7���y�I�5��L�dg!��ꦠ˖�y���D	0D��CZ�R�kL��yB��%dJ�P�֠ʂ.g������y�1v�0�G�H�(0�Lj��K��y2�_S�N	��+%�̀�e���yR$[*c84	���J0�YQ&��ȓd.���&�9$3���Á}�T��ȓF�&l
Q���!pl�a�:t����vӐ}��(��5y�m�7&q@�ȓ�D���iX�D� H�En5C� ��'�h�x�d�	�<P8�$��eHB`�� ���R� �X�{��H�aK�q��O�b9���W�ME"bu�܇�^�޵���H&a-v��06J�I�'zNu;�B�L���aȒA�`���'�.��IۓVZ�9����!1��}��'�̸���3y���� d�)
uI�'�p�	ƍ$]d�[����
G��h
�'���Dg�=c�g����
�'�N)j�@ؙf�v��T�}ɉ��� d���.B��	ͤH� �"O��-+�P�ə:M��Hb"O���'-;����P�T<a� jV"O��P�D"#B��3�XX�
Uv"Oz�*o؂:k��0���\dD�'"O������)�t�a&	Ej��Q26"O�*��ުY�� ǅؒ.�l�"O��@b��w#��04���5��Av"O�tȤ(͍V�����[�Y���"O�ٻ�U�Z�X0��<`����"O,���`ީn(�TKN�*����"O���	ǕX���zlW�d~��"O��C���	5�X�a�(ur�E��"O�Hh��������^&@��"O,�{�:P���S��P(���	4"O�q�ʂ� 1��C7G���J�4"O��i/��{&�}��6i�� ��"Ob�� ����.�"d~ZU �"O�}1ƃ�@~��§��0P\@�"O8$�ÅG�	h87��^,��"O왘�Aن!c�p#U$��#!"Op8�%�:@������Sq�x��"O��)�A�5{�
T���ǖ7�8`"Ovu.��1VI�`���蔅���y>!�\��
�R���tl �y�'RNE;�̖Kܪ	��M��y�h��`/@��	"M���G��y2ʅ1kb.���?F<�[Ee��y�F�[^i�'�^�h�:�:���2�y��
8�JPpR' �nq�,Ec٩�y�#ʐ]�����Gb>Lx��Q��y���(+�dۤ�C;+dƕc/H<�y�߅=���b��۞p�V����y���K�Ҩ�`ǁ*J<���R�<!�'C�VRY0�R�Zx�DCҨ�Z�<9�MJp<� �柍e�:�s�Z�<�!��,e�pH�q�W�^��1�JQ�<9@�+J���C�	A �J�gFK�<уb�
6��1�+LaQ����*�O�<�5B�@6���M=+atL"C�GL�<y0㒶p�i�W�Ƣ=��F�[I�<1�+�'��]�ǝ5�Xx�f }�<��-�1#��9��%�9���T��}�<�D�o�)�EB׍#7b�F~�<q $�622����(С������A�<y�� Ltp��&l��(�=3��LV�<��*�
O�t$U-p�>- `�y�<9qh��1�#�R-@g��c�L�<A�O]���ى���?��0��F�<�vOE�2lF�cb�f������G�<YBd�<i.iedʉS��8&o�<Y�F>pM��!D �è�g�<	d�@�/�hQK�o�"jbֹ�g'�[�<	!U)Z頖��'�����p�<1�^1�.,��Z;O<�� B&�f�<��傿C�(kD�
�OSF�h�d�<���@��q2ԅ��6"��c�<���ǿ�����M�*'T��Pw
_�<1��4Ar���ՁH[��x��X�<�$o��#���AI��*���`$R�<��+*�Z�y�L��&�r\3d�[L�<gg����]SeΚ�g������IJ�<y ���w�|�ɲ�))R�b����<QT_ִ}�w��:o,��a�~�<� ~���$���=[���l��	�2"O@1Kpň��潈��"uL]Bs"OB��@���h��Do�x����"ONzti�pn�UC��{�,5y�"O���sE]�m�Z�3���&�v}�"Or �1�W��z��M�,��b�"OF��C�	�M\l��@�>WvB� "O���-`d<��e�bI�A"O�a��ЈH�
��Ǆ�Wt���"O��2���+K�n�9�,މB�sd*O�iɐ��z9�M�լ]�����'U�6M��9萬ţAdzM#�'�0�;W�Ԡ@���䫛�|g$)��'�ޠB媕/F���ª��}�d]Q�'
��� <���� ����'�Taf,>:�fA{T�KI�̬�'���H�@��`C.ٖ*�J�z�'��=� "ŒNn�r�"��#kll��'W��'�N�",S�aܞ�&=��'�*ӂ��/u���	�!f�	�	�'LP( v�Ŝ�dm !��#&����'Z�ı�,V?
����懬�����'|^�K��28��X1�X<f����'8��Y ���=Oʙ���
W'ހ��'���j���k��;�o�|Xؕ#�'/nًS�ԡ8m���5i߈_����'���@�f�,�q��+X{JH"
�'����荍�.��D��L���;
�'�bu����<jAB bDc�pzِ	�'ࢱ�x��HDiE R�Ty	�'�Y�@@�����SoT0�];	�',^��m�"9�is�W�_���	�'���c�_��p��C4[��X�
�''���MѬ6ﾩ	�f�!�Xp
�'�L�3%Ѿ���Ѫ���0�	�'�U+!DT06�k��F%��`�	�'.j�1j���J9��ǀ�p�n-��'���3Q�@�0
���f�mnJTj�'&�I�k�2�݃u�а_��A��'�Ād�Ϫ3ZQ�D��RB�܈�'0�TRd-W#�쁗mܠJf�L
�'ti�G��.��h"���;\�p��'�RP���m�y�ܑ DH���'|�Ғ!�-F���cq��a��B�'Ո9yKP��fȺ9�i��'EZ0�I�~(e눂y-����'�\��ˀ> �!x�B��\�d�	�'����@�<[����ޭUz���')��ZF)0��5I�@L�@_����'!���$3���ej� Do̡�'9�Y(P,KE0PU���-��	�' \=`�+Ȫ9�ҽ��Q�#����'Լ�9vw��ҳ�0�-V:D��)�IC
q����7MP"P���d�(D��b��Gtơ:Ch��(�J��$!&D�(j�瀼pKR�IP�S�.�x���i6D��POӕw���mP�9)�݂�"6D��Y��h�t���˫X8\Rň(D�(��� 8��d��!ʛ!�( �d;D�<8¦=�H���@ӓ"v�r�M7D�0y���8U�����T�E�
тr #D� J�a��lbpJ�$e���q�&D�����G�m���n[C��8�&D��c�ET�FZ�yJ�$ߚt\��8a�"D�� ��S6��j��u铍�X�$i'"O�(�I��|,8��[�F��ᨤ"O��:F̚=<���r�*ɘ{�"�P@"O���e�/)��p�! �Б�"O�1UL_)8T���&0�nUb�"O>���+̄/3z�2��U�-qh	�"O4�n�5k�I��s���cH��y�-�D�����V�6Ub)�E۪�y��]:�`!a@�ڸ3�N��'�?�y�i���7��zH���Μ�yB@�p�P����ʦv��qc�@E��y".\�j�s6b®nḇc�����y�Պ`�*�ժ8�.i��C˨�yRK[:r����'4��T"1���yBFM�r��93���E���y",�?6��jY�w2&!�5���y"l����UX��-8(ֵ��
	"�yb�;rh4�3b�9,�܃3�4�yb��'mId���,�"�DLK��I��y$Q�K�<��GL"������#�y�*[�O��(�UO5!`�-8$��y�+"�l���(!m�aI��̊�y�Eē5�<{��ů|�pɢ A1�yr�֐%��9�Y�Ԉ��f�� �y�ڵR�����:��Ʌ���yra��&���k�4yȀ
`^�y��Ȧt�r����o;D��p��	�y�nG䎩3����:�^��E%�y���x�iV�g��6B[��yB(_?s���ن�bZ\:�i�$�y��E�%R�n�����R��yҨH�%4
dQ��ҏz��m��yc0e�xՠsG��j��QhԤS�y2�U��]���P�@�8U�̰�y��V�WDhc�ɐ��i[�	�>�y�;0^��#ҷ!�@x����y"ʎ#�M�GI����eK��H��y�e̡=����C�<��iy[h��	�'��]`�Ơ(k,�� g�!�\�0�'��H�HK
`w��.�5&���	�'<�RAO�!��ID��l(�2�'U^Ԣ ��0$Ϧ����ϧh�05�'���H��+׶�a��ݯZ�>@�
�'`*TT�[8<<�"���e�����'�.`���V�^>"r�"a�f)�	�'E�Y��Z
�TH{���g��	�'=��$ !9��3񍗦_���K�'�� y�_�N9�$�0���2��Q�'�-;�C�5g.( ��`C?����'��W-ȟw���QÝ;pZ�c�'�Vi�FX�Z��Я�8�J��'��q������9�R�'Y�\�
�'e|��
u��+AI�y~`(�'�&�z���'V�60�e�w�ҩ��'X\�����5%U�t�'x����'�
�Ғ��*lƄ�T��4mQ�X��' } �CT�):n���(�	��'���5��
�aR&�����'l�`{W'G;r�|��e��or(�B�'��I���EA��qq&� k�tii�'V�M���@�R�� �Σd�����'�b)�Fď0y�Ĉ@��F.$ջ
�'ޒ�XF �:6�"����Ҵ;�N�X�'#l�)���7u��R�FW�-Ǭ����� )H3��Q=�ܐ�e=z��8�"O�ݪcG�fe^͓�dה0��ES"O�A�Ƥ�7s<�HD�l��q�"O���T	̙A�慑���*��� "O��9F(�b�.��a�ȗ
ֶ�8"O�H7��	o*�FD�H��y1Q"O��c�� L��p�J�s���"Oؔ��D��|<���WL=D� �"O��#'*>c=�-?$ay"O~�P�Ǌ07�퉁�P$�!{"O�1�0�WX�����e�8,��"O����C�lM
ԊÖP�X��"O\l�r�.-�Y�A���:A��"O�� ���%Ig,��u�Lq�"OZ�+֌Y�nW>Җ��8R�x�"ONY)�@��U,�!5	2с1"O&\A1�+z�
,:!�ަ.���P�"O��-�/�Z��I�-	�֥ʷ"OX����(!;�IH�I�I��@�"O�X�	U7]�NbA�S>�@I�"OBeJ4�E��!I�!�8�&��"O��q�VT��;�M��&�>p"O�$CW���K~E� G$�Z�k�"O ��Ix�R�o_(<�4B�"O�l)�n�im����Q��ţ�"O*�v@׿�.I9�
W�S�D���"O��i��Ԇqr�9 H#<�r�"OBT�c��(p}&R��#-:�5�S"O>9�0F�6,4��Y8X$���"Ov��dC�{"�Ԣ$�1B�9��"O
�6�� skhC�W)2�I�"O|=�"�(|��S��B�;qܿ�y�l[�^���j��"<3���>�y⊒9���*s�E�I��g���y�hQ+A�����G��@�N�I�+���yB�09����s�þ7B6��R�K�y� f��ȑ�LQ+�u�!H��y���2^��aj�{H����!�y�X
Q��2�L��tv<��X��y��C�v�YF�£9�B�C��� �y�)Y|�����C!Ao�PaGb���y��؆U�0<),Ҕ<��i�&�Ҙ�yB�un�����:x���e˞�y�� 4��S��G�-1�DX��y@TD�"ؚd
ݽ@'���k̑�y��^�R5rMŲL� 6����y���('��`P�6T�� ��y���;p�,�b�0���#�y�M�7ZEd��& �)X=�W˖��y�iخ_f`��a��	�Ԭ�g)� �yR���|��u�Ӥݦ�TEaW��.�y�L��v-sW��|�����Ψ�ybo\xwr��U�I8��I�`��y��:*ނ��g�ͩQ��A8&
���yb/0���P���*� ��y�B7)$��hC���t�
`��B��yRHD.7���'芬_��dH�(�y"l�}�lK�B���dj��y�ۏo��q����ƌ�^�yR/�d�$�*�48��O�C�@C��,p�T0���A�l�LSʀ�7�PC�ɟ�����-��Ay���`F_�5�C�Is h8��]����r��<5��C�	�qQ�
,, ���jEB8�!�� ��yN���)����2*0"O�h� �M��0يƪ���m�0"O,�ї.$C����Dr�0�J#"O�Xb�-�AxPU�gBŁ>6�;t"O
U�FQ<���0�x��t��"Ob��r�� U���S-�*L:݂p"O4U1���
>.ECA�Xv���"O��!�I��3#��	b�ĢG"O���*�f��!w��JY�"O֩#�MV�,��m0���y�� "O��j�����,MY��#�G@:�!�d �X���
%B�@�R'�*�!�䗥FQ��1�n�=5��<�,Ҏj�!�DX�?�"H���������ډB�!�D�PGzu��A�V��d�a�)5�!��+$b,���"�5=�����oK<!�Ą� U���+�5 �ʐ��o��\!�$Y4p����G�$!�rJ�9O!�$I�n#�Ȓf�p�L�A�`�3*:!�dܭx�ƱsR���qyz%I��.5!�L�{�51�Ϛ� �����-��d�!�DǆD���Ѭ�<�2a���EYr!�䟀!Ƕ���l��&�����LO�Ap!�R���zׂ��r��+�*Qm!���H4�9�i2a�V0���R�@h!�˻%6�l�'G�H]0Ђ��pg!���G�,��o_/��9�$�K�<\!���cA.�i�KԀa)�ĭfA!�V�L}���s��/Ӟ���^�"!�U��;q��|���U�X!!�d��5�� Р��� �vDM?!�$mE
	�o۽���E�V�!���Q[,y� )O��AqA
/!��!�(d�Z�`i����lN�1�!��H�,�JU���
g 99��w�!�DE���@W��-a(6�hB '!�^%`{$�GB��1A!�_�!�S4��9ІF���u�%��y�!�D�Y�$$K�*t�z�
Fb�5!��K
@���K�.�H���I!�Fi��lad��4�~ "�]�.B!�$&R���Qbܪn���g�#�!�d�,�&Y���W�6�D����0�!�dS�G��̻���2<����Y&w!�dB9�v�j���8��BsK߆XC!�$�'C�|E��-ֽ&�d��5�Q�d!�d�5��0!�[g� H�%iڲn!�䏭r�< 1ԍ�+��rAj�0B!�d�W6u���0i�p�sr�As+!�$	�~�a(��B����h�5F'!��d�A#�ǀ�k�ԝ�"E�J4!�$� Ҡ�;G\S���+0��0!��5�n�ZU(b͎ЉR�A�p!�O�>1=�R
[�$�f�� B?9�!��!K{�Ay �ߖ.s���� �%R,!򄜠,X��#��>oHp�E�T�f%!�d���.�%��*�Nt����/;!�DA��ГW1���ZC�%W !�䇅��a���7?ZmґHT�Y !��\�8��ᗤ->�8��̜ Q�!���)��Bp�S�t/��{�!!�D0�-��ѥ%F
���%
�f!�DI�Rn��!�"k]�	�Q��!�$�"M@��&���!�%`MD��!�� ,]�eeԤ'a�����ȣ�"O�-���A��Z0��n� X��yi�"O�5�fU�y�vݢwL�6�q "O��i�%πQ��!&�>&}(c�"OpҠ���{Np��O(=��"O�u��� ����b�9_�%�C"O 1��A11E*�{�H�9 �vaT"O@QS!`�%k��\��(G�@�l��""O|�)��".w$����	gа��r"O~�8�a��J&Ú���B"O����@|g�aJ�ǾL
��Q�"O�mzeǅ�E�\U[��1���9e"O���i��c�x�en�4W]�"Odx(���j�����Ҹd�4�;�"O��{���+U�H@qEV���x"O��X��h2�DXW�څ��"O���%�&b� (��@�D�ʽ�"O��ՊJ�Sg����49�̰E"O^�!"M��%Ǯ@�2��Y"O:%�cĦ�\@��bM7e��(g"O�Ś�iЏ����2�N9{� ,�""O�ѣ��s7R�	A��$.|t��e"O�iYC��n�$�㧡�(By`p��"O�thd��&NI�ڨI��U
U"O)ѧcG�P�� 1HW�{��0��"O~�p��	/4�nM�d��Dr(�b"Ob<P4��"\�L��A40U-�"O��mW	n8�ЏO�ymj��0"OJ�-y����
T' �TҢ�ʤ�y����r��6i���m�"��y�N� ����ߦ>��$�Q��y���P�qZG�ʲ( �Q�e&�1�y�fE&P�$c'{RȪ���-�y��ƭg��� 0�D/jn����^��y"�� c��]��Mlv�a�%�&�y��s���A�f](d�R0AäS<�y��O	VV~�mV8��Y���R�����J���U���H�n��x��]{���� 
��$�C�fB��ȓH�֭@s�#h�{��%p`�����x�k�ڗw?��HR ��V��ȓkb�ٻwkݧv��.\��9�Re(-��[��(CN?o�U��2������@,$� �������1�ȓX�`�H��ĝud"hࠀY�99Ȩ��s�d*��J1N?h�sg�;w�H�ȓg�|�����q�ۢ�G�&�xM��V
>��d�8=F4bS�����ȓ����$�H�5@ ��7�.���W4��4ά��E-��f��ȓGx��[:w���D��;��ȓa���R�)&,��@���!�����$�Aq)��`Ұ`�䕊4GHa��0~�1K�	!q~��0�I�4�ȓ=|�DI'ꕗ*�-	���t8
��ȓ'�f���΄�^�^4閁�%R̶Ņ�>���	��0��HjA�#e~u�ȓxc��{�nH�`��H@}o6T�ȓ>ռ��TR��~Ese��OƬ��ȓ8������D�A�L�5�t��ȓ\:�1f�1�pp`R;p�@<��[�>4�P/3i����H^�Z���kX(� %��L����2q.N������h�C�4�sw��S����S�? �¨גe���u��jBx	�"OV�ڤa���"Q��x"Y#"O���Aɽ,* �k��	����p"O*}�G�3�>l{���
�4��"OR [�$��>A�-���F�C鶬"Op��c�6�ک���:��U��"O$��ClN�\��b�	Y��0w"O���
�({�����!D+l��-��"O�a�7�Z}�`�SP��=c�=Ѷ"O��Y4�ԥ;�^�3≘W�y��"OX<��A\��ݰ�(�G�D���"O��cD%�<^Q󆔹ox:y��"O��e�	u��6������Q!"O�����W�rL��D���)T��[�"O�]��N�=�ʉr	(8�-�"O*���@�dr���,Jx� {�"O�u�Va6�<�!O2_bR�i""O$A�5AJ�n�
���o�I��9P"O��f�_j�1zc�K�*����"O�q���Ȼq9HŰT�D�p�)�"O���%Ԋ�3�T�����E"O�剡�<A^	p�j�a{p5�"O������*��m냏��Q{N��S"O`}y��?�H�A�N�0k�pb�"O����ゥ
�. 3t�R�Fa�3�"ObHR@��n�$��@յV$��"Oa�T�Q�[P�A��H�_�I�"O~(���ڈ)AJ
#FE�]:w"O�U9DgI�	U�(�愴fRƝ��"O�0%�%X��� �0`"�,��"OZ�ٰA��UB�֮ڜk`�Q"O	B��ʶOV�i�f[�E��"O����P�m�h˶B(6{Xhɰ"O�Pk�`�O+�M�U��hz�i�"O�г�'�3z8&Da��5t�\��"O�@��.&�!5�٬7]�5�s"O|!CƋ�L�j���B?zJ��"OXI	��ܤ�])E�͏(��9"O��1 ԟ]�"�p"'��#�`|1S"O|h`�m�!`;� �,D�Y�L!�"O���1-�P�@3F�/n�����"ORY��U2Jn2R�߰q���QQ"Oa!��Ϫ*NF-8�e�L�R�t"OtT��B�o��:0��&��I�"OP����%H�\�ԄJ
�,��"Oؠm�>���c ?׬��p"O��P�#Պw�zi"�BM!o��h�"O2	�#��'>չuH8?�zux�"O����� P�]�D&�8N����"OJ��4MN�.&�-���N�!4h�"Oб���
l� ��	:2vl�w"O���S��x���B�Kdl�9A"O.XcՈ;�&���I%.$�A"O�d�E
7�8�a�=k}�q�"O|��&�0U�Q��-n��f"O}�t�LʪhKC���Z�(�[�"O�H�s$�=,E,KN`�pMX�"OnIH��:��)́�y_֐A!"O(�#3�j1�1�g��*$�p	�v"O�QA�C�:x��5��~ٔ,�R"O*�
AM.{wX\��j߉@Ζ�ѥ"O�ɠ�Fٰ��u RI�&dn �"O(=[��[?�H�Ř(HD���"O8����3A������% -��ʕ"O� �-rp��:�8���%t$�Y"O�h�P�Ĝ�@l �iZ?84��"Ol� �f�ô��e��s�Sv"O>eZ�g�;
� �S	N( qt��"OvѻW��e�\�T��/]n}r�"O�]�̎�	�l=��FK�Cv�P"O��Q2b���!�e��Q�92c"OhY',�xq���VT�-8��"Oڀˁd��Q�����"O�y2c�V�WQ�xPƂ�r�8@Jd"O�Ar$�N�X9��U��"O�|H�g� ֹS�A �N} u3D"O���cj�#���T!��l�x�"O4���D����ϖ�BGB&"O@��TkR�D�&=I��ġ"O`��A"ON���c$|iGDK�{(恛�"O�Mb��߸b������<�6���"O0�G�}Z>8��f�!&{���0"O6D�p+�8j�� C�'n�p"O T�U��j���`ƁxH�J�"O �$L�
R��� �ſ*^�1"O��k ���P���P�K!,��@"O��`F@����!$D�B�^6Tb!�$�|L�C&&	�sXڅ��BfZ!򄖐Ş@G��m@�c�#��8�!��օf
�hX�ګQ��y�'u�!�$�7I(�8p $|���/ۛo�!��pM+�&�	T�I!���*y!�	���j�#n:Zp"���;@i!�6�`uZ䮊�W�0���F?}e!�D�?d�dLasc�'tAd��g��fl!�ād ,��	A\I�!�Ԅ]u^!�D% ���ӿa��Eq$�Ķw_!�䆆�����ϕ8|���;bE��k�*�93�4A�h���̸ j(�ȓ+F�a-��L�l�B��E� ��ȓK��J�0:n<�dȌ ^���ȓv:L�xv�
u����2�\�'�܅ȓ ��Ѥ�ײ!.~<a�H�ƀ�ȓh��0Ȥ Ph`� ���|H]�ȓ7���P&���0�u�G�B6�ȓ;q�%Ѿd�=@B�����I��V.T.��c���w6��ȓ)�
��p��=f����蒋5H⹇�E���5���]`��Q�b8����a�9��K`��ꊨFu��ȓ|Z���ME	t�H�dæJY4Q�ȓ����%E�:�<}�F�"�h���H	` ���j�M	�O��9 T��ȓG�L��C]4d��!�b� eop͆ȓƙ���ʨoNI�TO%K�8$�ȓt���:���klְy���h���ȓRP��C��C�"H|�	�EN�`Ԡ��fb�%�vK�F�y�_��Q�M�<����>��ٰ'nތ���p�J�<qӌܽ%�S���7��Ы'b�E�<Y���2E�a���[�Nঙc1��g�<)`$�k����ML�JU�A� c�<9�❕/�>ݒgb�'�8��Q*�_�<	V-�'X��q펢�J9q#�d�<I��A2f�5�ĕy��x@��d�<�Ä�i8�H�gҎ*���S�G�c�<	w�\;���*��yk�Cz�<��o�*�$8e��.lq�t+�r�<� �J��:v ,	���*m�j��"Oq׉�v���bܾM�$�0�"O�ZT+�6m��� ϼ+0��v"O�|� \'Qt
�1��s.���"Oizd��V�b%8s	Ԧz�"�D"OZ�kV�a}�
���oNV��a"O.�!�m��I# f��D0I�"OR��І�6d�8(2bEY����"O"Y�W�P�E��Ha�E&=nTZ�"O�8h��\�%��)p�ߖ!}�pu"O��a�M+Kt�PrT�E2Hdh\ST"O����.��x��-!bV��T"O�X(Í7д1���8�r���"OU�N�e�i�&�ΕS��ht"Oh��!�UQJ�5�U���Y�.@r�"Oz��v'V>V\��q7c�#i�~�"OxItB�
L�@�,:-N�+�"O��Sp R.LƂ��� Dn�P�"ODTÓ§5Z�c�E�!j���"OD���R�\�I�mI�f���e"O�0SשS}�Q*��W�WPN��"OԌh`��kVx��F",*C|��"O�(�'B5l�|�q�
D @7�|� "O�U�w=j�$h�P��#9�T%��"O���F`!,�� �]�C�P�*�"O���u�F�& ;ƍH�xܝK�"O�����C�<Չ�,-~[�\H�"O�Ybt�����lQ��/Htz�"O��2�j�a��"�	N,��"O��!D	�Py��V�(�D�"O �P$�ĚY*�ă�L�ފ�1"Or)�	�V���� E���	�"OduJ�-��-h���&@�`?�R�"O� ���"wHA!"E�7zPvXCE"O�xrBk?A=���d�sLt��"O���C	�>$�"��#E��ހSa"Oع#���>��<����%�6�j�"O���/��G��4jT� �Rm�#"O�:�Kۻ0|v���NZ�
��Ea�"O�e��3*(a��T�x܈(�"O�L�QDJ$V*u��(ҳX�iE"O�CAL�F�L�H�G��X�����"O �{f�B�&3'L<oiv��"O�$���*(W\`Sd
�aN�$"O�}Z0F�'>�Lp���>?f�U�"OTY
ҿi$�'$T3O c�"OD�z�ƞ� tT`�I͟R3���"OV�r�ɓG<�ٖj֊;:L�"O�� 	LY�L����r'8�K�"O%�V���E[_�fpPA�"OP�(���l� � ��].k|�l*�"O��jէ1@���
��W�Q��-IF"OB	@���1�Q�&'	#��� "O��Z��E�N�&���*���Ʌ"Od���7-t�C��RyJ�p�"OV`h �|���be��9g[��d"OL=Z�
°OYp8"v���kZ=��'2���H_�'7�Q�d��C��!
�'\*Q`�
��q�sD��R��a�'�����nߔ���;�O��7 D��
�'�Dt�$W(X�Q����!�'�.ؠ�[o  g�C�g>�%p�'�V�;��,X!	�f���H���H�'���ڰNP�O'��u�];=�±���� �yX��5;Ú�h�$��p0ňf"O�P��&��Q����s$=s	T�"OR�I�d�C�$򄅑q �A�f"O�i�f/X ���bČ��B��"O�@�%�� �`���3d���"O ��T��16��5�M�f���"O,�jb��d
�`�,J3�8,�F"O"Ux�%��%P��T�D~��"Om�.�i[�|3�	�6�B"O���$șb&���fȈ�vz-�"O9(�iV,U�.��%���ãz�!�̜`*zMSQ`ڦ=��,)d嘓dH!��:���[d$��W9V5Je1H!��R�-ب��SIT��rlD�K!�ě�e�H���)%��P�A'[!�dQ�*y�� [r3p�X%� Cd!��8lU��1ŏ?��]�U�/KW!���zt��7F	 �J�*ݛU>��D�'��4	��]�ȴ��y�S�$�٣�ɕ2Z1
��c���y�c(���-=;l�eg
�y�ύ:�>\H�6����ed��yb䏘1b�]������BS��yR�L�AWX$[���5�� ��޵�yRmG'_�0{A�
�qt�_5�y�+U�eLX�P���dD(��(�y�I�E�E�#L6ږ���B�y�&�8|��C�Y;)�zĸ�n�y���P���"�$Â "�-yQ�:�y���G� ����a8B=RaE��ybH�'B$ٓ#FnD��u��y2쎋�Z��UA�:���{����y"���,��8�.4 A����Py2�0%���s��#p0���^�<���H`����%�A}�L��ES�<Q���;9?��էA�I4�6��S�<���f-� ��*��=#�iJN�<!ЫU���q"��ƴ+�*�@�<�u��S��}�$!���̹b��@�<!�Li�L+�d>k��xgN�{�<�˜%)B�:��Þ"J�����y�<a��9F	��1�;`t]R�Lk�<�OZwN2���*�/i��9Tφj�<A�!8��
�8�FVk�<�4	�<����AM/N����i�<���_!_$��FD�r4&堥kEA�<)6,Z�*��� �7 �6 
eDW�<9�o@�&��JǊ�0A��a�%��h�<1W�_0�lX`�/�TaR$�\�<y���	h�f0�O��p:���$An!��TC'h�z��+0�$x�*��9O!�Dъ.��#���"�����d%F!��0�(E�C�N�t֙���W;)!��Ey���#��VU�7��.d!�Ԇ>��H	'�r̐�' 1O!�d�B��ץ�f%9�HF�4!�$�,J�B���?��YeAS 0 !��?�dh��"�VR��M�w�!�ą,���Vj�	:t �T	�d !�d�U��X�Ñ06fA�Hb�!�$�{��5�CFG�옚u��41s!�Ǘ7� Q��O?^���1g�1�!�Ĝ�덀�cяQC�I7�V1:�FC䉗��!��`hA�0G�.C�)� ��E�N6AZ18y�V�ir"O��Ö%��(�Lk�1�H�C"OZ]�&�B*]S�8S�j�<uQ(�"Of���]��P��g*<<j�aQ"O�|�KS��P�)B{r�x�"O��!�ᙽ�~����`�ݚ"O꼘D�^�C&xYrg脽R2�XP"OD,���+�<�A�#����"O
���(�
 `%"¿}���Py�`D�e�؈SA����a�7TR�<��hP��
4 ��e�Z0{HH�<i&N���l�M�`���.��<1W���N�΍w�A:kX�Z��~�<1��ɯu�
��ԑ_��QA�	w�<	�GB�
�H��ι{I�`��k�<����5���`!���s��|{�~�<Y䀞"4�Q����l�ySf�}�<Y���.F��K�M��Ka��hI�{�<AC�âC�U��� ��� ČIo�<���}d`���&"$T�7J�f�<b [���1-A�	�ʴ�b�<��/E4?4LtB#��ef�6.��y��2g������pq� �y�&M9$�y�H�	t�͠�嗨�y⎁�; ���h����ٱ�k@��y2ǛnD*<��Z2`�Z�3C6�y�
��|ʶ�`�(a{�n֮�y��� 0t;U �_Zl��'Y��y��80�2���-F��ƑaB̆	�y�M��&yR��%�1�8�����y�
:�Ҷ�W�2�eYU�T�y�,�5�p�S�*���(A�yRΗ1&�Q�#��!u�Ʉ�ՙ�yr�[�b� ��Rjŷ:-s�)\��y�HR�r���H�@�C�c���y���:V�q��4	�N̸ e��y��.�&�!"
�(	�X�cL;�y�DL�-�~�p@�ުX}��(�	���y�A�Pu�0ƌK����6Jہ�y/�*-2Dء4mF�G���y�'G�y��R�D�W��ccb(�y�*5� daH�-PBI�dX��yRY�jҌy���/;+l��
��y�¹0�1���9� ��4��yBkݨM�J�"S���8u^� Ta�(�y�̡fn���� /
�[R�\��y�O�1�Т&l(�t�� D,�y��"k�f�#���;�z��͌�y��ُ"N�Kg�XCj<�y�bf�)�1��O�� 
���8�y�&N�OfʰZ�k͌AH�H'����yBgU%?W�a��ģ3R����%�y��}66��CK���c6&��y"�-h�t�"�U�;M��5 �(�y�뇅<নq�C��"�^L�U*̸�yB� :G�4Dq��V�qDH􂈨�yb"�*��5�v��8N������y#E�#����En��CX0�p&f��ybnʭ@#N�a�.���˅ T?�y���M���a�;i"���B+�yb� Wz�ڃj��H0���L��yB`�2%�\�14�V|�lX��Oȥ�yb+�"Z$��ӭ��v�:�kw��y�(�R����'h�2`�r(��P��y
� �m��f����pIq*�6(�A%"O�8�V�b�V�J	����X��"O�0�,Հ$~ԉBu����U"O�\ò�l ĨKgCzZR�"O+��O"#����TF��cX��"O�ݡ�cH��Y
��v8�E{�"Oa�B+Z�
��D� �Lu��"O\�U��7_y*(�ו�4�j�"Of}i4
W\h�+ǞA�z�s�"O��@$GޥTl*tD!:h����"O�A�s��
y�)k�oF�K�}5"O����V-p@�a�o�"D�"Ox)��!
�X�Ӊx�h�rp"O��!Ұ~|����Gƃ*c|I8�"O$1R�k��	x,�����@Z��م"O~u��o��2�� ����1�\��"O�}�T�Z�9�ᢅ$O�_��as"O0�(�!ɐ_��)�i� ��y0@"OnXK1'ٸ(d3��O>�l��"O�h��ȥ&9��XG���g�e�"O�TiR�C��A�Ά�f�0�V"O(�����#y:,�Q-�G��� "OD4 �"�t�[�=V�^��e"Od�RVA0G��[��G��p�"OZܙra�ʊ� $M�=~,�"OdQ�����d�����<v��8�"O�A�K��%Z9��DX�K9ж"Oz�J�oE KHr�@�}��=[�"Oni�G��4�`� ��z�����"O�@� ��Ԝ`���Ѳq�
��V"O�		�J,�ј���&@q`��'"O��#㙲U+�mP��o��}0C"O�����I0z�0�����3F�g"Ozuj�,�hV��ÁZ�I"�	B�"O��8��װ>L���aظ)z�	�"O��I�J�g2�9cT���I�"O5�7�[�i,�]�ԯ�`F�hp`"O��ӣ� k���B�AN5@�\c""OH��ƨ�lV)
�(4:~HA"O�9����\��0���U4$���"O��]*��@���A� �q'"OD$�`�>!�ԑSa"ޏ~̌���"O~�`�/�I�깩�/?)���"O�(Z�b�W<i�B\*� �"O�	; ��e�:��%��9�n�K6"O` �f�>'>J�Цĉv���"O`8zT�ޟC9H��e	�k�H=�C"O����r���G�9B�|y�"O<�ie��Fo��2�cYg�@���"O�!"A�~u�1"�TdZ%X�"O����͚:rg�q&�%9���"O*�� �P!��r6�ۅG,�4�"O�E�a�_�R���Ia^�Pm��w"O�eP`�Ȣ���j7n�8 ���"O�t��]�5-���$L�5�ӤI,D��XBDΣ��̪��	DV�!EC?D����!��UX#l��rל� ��=D�Ԛw�I�4���`��H�)�M�'�>D�|c���&���fȋ|B��� "8D��Їk�j@�|��NF�y�l�Ath7D��9V��5M5f���Ŋv�2ap��4D�4�2.��<�*i�uʂ$I�&��2D�D�XbZQb��?N1��v�2D���!C^��NTW)�:3��8�3D�� ��A�"#��S�j�����"O���)M�.{����/�����"O� ��eOqKD������U��c6"O�<�RA�LT��v��B�ՙ�"O�x�P��8@�Z���b�<B�ʌ��"O\��'R�F}�Tr�&ϖ8~h�"OR1jW���1h��X�E�=0pLQS�"O�
���1,�rM�2$O$tC|%�"O��rA/,Q�P��u�Տ]XD��"ON,P�������ɪ!L�lQq"OP���fc�����8a,�)"O�Q��h���
�aQEȤ&���"O>P��̟&v�(�{�-� BB�`t"O��e�K`�@�qV��P�.�"O�Q�n��DR�Ex��ͨB"O��1Q� �ph�!2� 9t�x�"O|���&?d�b.Iyb���"O�ix��ίl#��gWgx�r�"O�����4��ܫ�E� d�p��"O y���3_�q�D
P�0�"O
Ab �îGm�(3��9 �b�"O\x(4�%0��/��V�iB#"O��Y�Ȧy,� E�"�lI��"O���gŋ8bF�sD���H�2@�@"O"-�@1\�r��ӊK�9�����"O�y�7⌴q}��
s��#LR�lA"O�1`�h�AH�$ �
?r,90�'��	
�ݬ��De�8N��k	�';���C��+�a�ԥش.%>�	�'��$8���
7���!�aN� ��]��'e\9s�J5�L��h�.�9a�'gfAaeK��8Jh@¡�$�'�FEr�Cφcz`���IC}^2�c�'�0��"D����7E@�"��I�
�'A$��!���<�G�r��	�
�'tЕ-��G�$�;�"@�.�Y��'�R�9��bpp��vMR��Ԩ�'�UkW��m��AsC���f��
�'V�����ŗ>`N�@n��|�Jp�	�'e��C^5<�*�r֕BCnY��'��lZ&�Z�+��T���W�8�yC�'J���qڇ0.��zf�N9/���'k^-I2��J�D�%��,Y�`ER�'�Ωq���|>����l)HP���'ԄM��͙T�5�� �l���'J����"W����B�9����'�R�����0�*P	�V���9�'6�Ȃ a'"�r(Ї����\��'O�5�a"�5��tؑ�Ejh��'���8�֜\JDaOKdk؝��'�1� �[�}|�䉐]K���'�Y��Aǔ^q��1��D�")��p
�'�Pr�d�<"�\xj��r��	�'��+pn��3:���g�x���'y\R���6c¼!��bJ=n��Z�'v̀kI@�%G��!����t��J�'0hT��D�i��5���d� �c�'���'�%F�lQ��Ƹ]�Ri�'������'JV��w&�.]�� �':@5z�����ǆ�O�mA�'$x��R�?Sk^eQR���B� Hx�'��Z��ۡy�j b�dD$:��L`�'��8��a��4�r ��Nj�j���'�(���B3dݢ1�˄oA<;��� �l��/_�c��d��"��<���C�"O��R�Í�8X�aYO���`C"O�x�1��h��81f�؜�x��$"O���'�Z3@X�!��/؃{��x4"O�4Z6�?e�ˢ��;:ZX��"O��VlϡD�|,	E�T��I��"O)��*K<��(�E^�+�"O�ɢc�Ğ8�q��"΄)� ]��"O$�
������,3�8�+�"O���E'I��㣁��h-��"O����J�A�B4�� �tV=� "Ob�!��Q&w���� O�Yk�d�"Ot��6��-Zմ}��N�v�p0"Ox�ŋ��
�rŞ�xx53�"O����j ?T�Ac��%t�̚u"O
��7��b���+���B��}�g"O���K0Kv���7Ύ��ĕi"O,���	7:���c.hҾ�b�"O�A�/�n�h��"8�|D��"O���`#��F����珊O�@�"O�k�O!����!.P�"O  ��$�4g�iP�g�kH�H�"Ot��1,[�2�)2�/
���"O���"�c,HY��$�3' ��zq"O�;d�7�(3D���D��e"O0���"	�@r|��B�)�xAy1"O��5 ש6�
�Bk�}<r"O���`ĄT1l�s�ƽͬ��$"OR ���D�U�$J׫Y�]l<� "ON�ɵ��)| ���d�^�dUc�"OXp+I�%[	��a�"��Y"��2"O�Q ���'0V�`Htb�!2 ��Ұ"O��:Ӆ�2&��+�B���"�'��.��)2�����P1��'���{p/�>�[0�S"8I��P�'�~�R�	�]i�5He�S�]p�m��'#�ͫ"#�j<�LH�.F�x=��'����� �#=RTs'7K;��(�'��pBd�_"h>Q��+�5l�f� 	�'R��e�Q�����𢅖:^�=A�'DJ!:�k��G<<I����~e\\��'�.��[.����Q�Xv�v0p�'XF�`��ѨS�n��jjȤP�'������= C��2E
��_ E�'�^�����[����חLN�*�'YxiJ ��r�x�x�$P<� ��'�(-�:^�pP׌ɺ�ЙS�'��2�۱oG��C�oA�iEV���'��BW�ݪH�jA3��T�b��h�'Z��Bϖ�"lP��e��V}zC�'$E���">U�Eqb�CJlFa�'�散悟; "�AC�A�?p ��'��	{�JͳU�Ȩ���5�jd��'(z�Al �X.�`gl��f!	�'�2T�� ��5S��uI~c��c�'B5�6(YRw�Q�M�pj���'G��2Z�
ʦ��Γj��f"OU
��6d�����ݖ#�d��f"O$�&�ƛ%(�ǈK�@�z��D"Oz�+�K d��UY�'�7k�
��#"OlS�[�V*V���O��d�"O��A�4.��yi��|M�� "O��*vK
b�*Ikg�/@)�YI2"O*pZ`mϱb��Rֈ��?�͸v"O� 
��`��2�Z��T�&�:U(�"O�e���x<b��姖j�bx�3"O��r���
\��L�ᬆ�
ִ�C1"O �*5`%�qH�-��oϔ��"Ox��T�S�yj8-��j\���D9U"Of}BC�	?!�HQʏ"p��E��"O8�Bel�!Xd@�8J=��� "O"I
qf^@���PT�S:�h�ˢ"O�4 ��[x��`ԫW��Y;�"O�@!�Ǘ�=�8h0�e̘��L"O�|B�Z�2��x!n�$a����G"O�ͨ���a<h��m�8d��P�t"Ozy�vH��`�b�0⬌s���p%"ONm�1��cT�0�n&plTQg"O�=�CI]�F�p0��.�4gV��"O"4+�I�Y�B1�p/_�8RL9�"O���CI3o���Fś�(?�l�"Od� �ǌ;�	��#לD9��"O|4{��@-7�v��!,���	�'��Zb��)
w�ti �қ%��I�'0��Ag���R�>�����+F��i��'MR�� ŀ�\� �u���;�h�'m� �5c[n�RH�5�I�dRR�#�'�@����S۔T@�f�)\$`�'~,�W͗�ji�㴇�;ZF ��'��h���̸@���T��"w��`�'Y���m.���c��*E��#�'�T��%�i(\Z�-&?��$��'>�]s�Jɇ+�0hb-��j=��'� �9�I�>��5#al�  Ũ(	�'VB�:AI�1-���CPN�!l���'�Π���ڽg�hQ����4�K�f�<!wE˕b�"}H���:,��;���a�<���[�XҼYQ�L/n��U�Gg�Z�<9�nr,�RqdM3 >��KO^�<I�oQ�U`e-�+2]�uR ʌc�<��˖��p�2dhƌ˗͔_�<�f��}M�Ū��m@�b��Q�<����M.��R�%I` �P�<�sʬ9�p�B��Nw�TكΊB�<i�%�Q�Q{'HS�tc�
�C�<�<5x�� �σ*�Bq��(�~�<���K�O[�9ä�X<5� �0��v�<4CN�X"����>c��Ha楏p�<��o�(M#$�h�
��W�Bi��Wk�<!4�Ww�\�s�	N�o��l�׈�i�<�����dh��v�U;=����b�<�!��Q�@���.C
E1k�^�<�%��%VM���W՜H��8A4�QY�<i7�̭9Vh�k�wV��w @�<�0'�5$1�uaM�jM�Q�ƬJr�<!bE�r�U�3�V�Mj�<��C޹M�,�AFa�b��h�`%�[�<�S'��r�>��B�	&�P9�
Y�<�uj�WE4�Ѐ/M�5��YAO�<�K�>Rn93�@U�|nhɈa�u�<YIM#].��F,P�_vX���]�<�d&Q	T�v�tjO�"FNx ��S�<��LΊWhj��a(���<@a��d�<�D�J2 &�b�Ђ��K7#�u�<�j�6
�v�)�M���� Հr�<����
�Vة�'uٰ�P���k�<9s�܉� �Q�ߤe!)�k�<%[#BC��Ņ �F3 x��Y]�<� �e��K��&���J ��YX؈�"OJ�b$GH�`D���ܘP�\"O4+�-̒d�B�9v&��jm��"OVy3���hPd� u���	�2�"O����̲Y�.���N�#[��!��"O�HvNʡ �h8A��9o��b"O<%2�b!8����aL-_�!b"O��;t�Gc�]�o�%0I���A"O�z-�1\2���QlF�@&ʭR""Ol��el��m���p�%~�q"O�aY�I��N�N�h@I � b���"O�sr)7��X�fԌ�-�Q"O�9�IN9ݼ�Gf
)�|��"O�P*�cǇe ��ᆏ?x4�A"ONp@*� o/ Q�4/f =`���X��TJ��W� x�K��H�*�RІ�{r�$��aE&&�f͛�R?\DQ�ȓS�h 2Dmȭp(f��'�4i����ȓv,lC"�Q����H�-TTP���O�XpPҩU�Ǹ͡�Y'��̓"�D遇l�]��IM�H�FLD|"m� D
6��>�" ҤG��y�&�o�6��#T�(��M��C�y��C7aU���S�B"�LI����:�y��U,��1#�M$@��H1�&�y�ǚ	K hA���H�,��'�"�y�!7;�"��!�T�{�����y�m��/�n�����4L8���1�yr�V1B���p���
E�P��yB,��C?6	����ǌY��Z��y2�ߺJ�da��	Ж̺g#���ybJ��dT���o�$��t�6
��y��IE��6� [$f]�&Ĝ��yRG�:f
�j���>M3���,H�y��P�q`F,��@xd}�!��'�yr�ן#������ P����N2�y2�Ǹ|��Bw)����I�0΋�ybBۀ�Q6n[~!��gX
�y��6&Q�ٲG^�k�����a̒�yr�8[6��X7�NZ8���n���y��]G�$��ЪʛO쁤�^�y�@�E��4��Wt�� u���y"Ң[4�����S3�@1�H�y�P3M�5+�\�f�h��ԩC���<!��ܺg�j��O�P!4)
E���p�@�Vd��"O�d���KUw� �T�O�s(�@�x��X�p��@���=�0E(G�˴J6�i��E�Y.��"O�Y�k��'@���Ĉx���p&���R��X壁�6�3�$�uΘ0�(�/SF����  �!�dÀsؐ��F�e��k�B�� ���k�(*m��*	X�|��J�8A��W+}2���9��"ڄ�ېX��1��CW`��hQ��� �.{|���&!Qi�<�4�89i��8g!ϭ\�X�9�
�dy"��?�f:��)h�<�����ȇi��i8��1<�9\O��e�ȓQ�xY	s�ޣ�Nq1HI�
�B�y��V�3c�9b��T����`�U]����U&�cfL�Mnj8��F
������M�5
%Q�bI�,��҄n��O�|�!ϙ��X���ީK��u��@,�O̰IEؓO��r�ƨ/\���c�ɛ?�ƨyc�XL�؂A*+[����On0�zG�X�7"�ȓ�nů$ �L�	�'f��G��4K༐�e�Q��v�z�ƹ}�Q�t.�(Z� )���)dn�G��w*�!�&JP�|a�$*�[]����'�b�VO�5m�F�H'�n^٣&I��h�dI��Op���QFT���f�t�'ߐ	��B�Mn4�F�Ͱof8��ߓj�����һjԆ(Q6�)K��4q�1nn���mZb:�ʴ�1�r��I�y|�]�d�	�K����Z1uV�P������iW�@��EcF�V�a�$�3� Z�ѵ΅<3�(�ڷ������"O�@�`��HQ�1�+�8Z:A��ހw  ]��ٓ���S҆\�P��+c��;��\�.�����AA8�h��!D���T�]?S�W��Dz
]q���8|k,�s�oG~��3TG�0� ��g���t�~lEy���U�Z�/V5i��kӥ[�p=�em��,��X�f ߝQ<J1�6�J̖�;���L�f=��lӠh�rt�T�I���|B�G9E�����5S��U!*��'�ْ i��D2��0D��#7��� ܭ	�T��.iz��P��PKL1��C�|ԈB䉬T\Ђ5/{�u�7�M',Cr���eĮ_�l��a'�}��D���V�����w�5iѦ��A����M´/�@�c
�'�IA�&�T��1`m]�.��<��)��Dj�U(%l���y����Yq�E�'\*�Y��m��E�0���j�8��x2(S![��$@��F��h�CW�%��x���dM� !�6x� A�'��]�V,ӦE!jբ�TQ���{b�G++��;Ԏ7g�&12!K�c�p��_?�) +L�50�Q:0��&d�C�	�h$�rE�)Cl����/U�J�vi��`C�S=|�r�	�^����G�O����;Gd��;U	X�������&�t�ȓ.�BX��I��~�JCG^�qR�Ȣ�;F�Ȳ��+7s�e9G��ɺQ�	�E�J�!a�@3@��uc�K���D�;_2jȉԎ�G�L��g�ɐ��u�a�M�j�B���Ğa��'� }���E�y,�@��'�$EB��$@!IL �d�g�>��"��#�KPM1zT"�N3D����U�S�� ±g�-*���"N�l�X(����z����R�Fm8(C���M��9(���y�O�4�+�*b�8�N�'D7�B�o��`��B+#�h��i� P��B�I)!�^������cNz}��'(|C�	9{���2d%�RxN�"�e�-�C�I<h�hp�D]�H V)��/��J��B�	�wI��{ӡ��2(m�F�˦)���$�&"��Bր[�6!�� @x�!���X�.Ś7��0!�!k�!�!�!��
\�^�勁{{�E�NνD�!�>�&|�E��!P�}1⋌jq!򤇀1W�T�V��B�m�2bT�\N!�X� m���q!^< �$�Z�.-*!�$߻4���
P������]�C�!��@�f���#�,D�>��Gk�DG!�Ęr��$����%#��d�M�x'!�$ ���ۧɐMX3A�H!�dΉwc��B"�	\�DU�t��d�!򤔡y��Ѫ���H�r=�Ղ�D�!�D^hִ����0�n�{ �K@�!�Ć��(|c1�9X٬I���P.Y�!���0���!�NH˂�9���!�DH�_/Z��@�1,�R�a��ѐj�!�D�+E��e���-����%�:�!�B�|���Se�B�����d �r�!�O�?fR���h��:x�M�Vߠ�!�Dח?�)kTmP#h�F��"O*Y�0b��L��o�*~����"O�A��!S*d�6�qM��]^UA�"O¨�ĕ�?o�iqg�+�
LK"O*}�� �N�rd㤧-d���"O���Ȁ-&�
f[�X�p`P�"Oμ�tB�9�@ғe�Z�Z�Q�"O��i1D�&8"���2	���b�"OF�y&Ʃ�����Hıf�`��"Ov	8@��G(=	RlX4~t���"O�<�@h�'o�$x�%ʬV��"O4���Q�PC��F����"O<Ř�ŏ1k�L�!ޘZ5�h! "OPE���ڳy3������"�= �"O �Z ҡe�ՙ�OG�N���S"O� ����NҔ��u	B,	/rT�p"O��s�K. ~	�V']c�8z#"Ov��`���8���6������B�"Ot$bh��>KH�˳��Vv,-ړ"Or���Y�QT����s�J���"O:=A�<9���`��IQ�3w"O���a�ɋx5�쒇��@#ƩP�"OL�d+��gaRx�eM̎k.����"OȬ�p � 3���Jb�޳#���0"O qz��ׇj�<C�#�`4"Oƈ� ��!����e/ڙ-_�Mx�"O܍�2�/]e;Rg� GDd��"O^ �5�
����"/%<Hn� 2"O�y0�  
�<r���eNBui�"O�Ń��W1~ \�h�ň0t& �13"Oz�3�A�C?�� ��E�pJJe1�"Oxԫ�װH��@��Ү�&(��"OP4W
��.Kĕ�hH1mR��y�!�?)�����ᆥv��!�y2��|wj�J��Y���)�.F,��'����BZY�O]��s#���uV�P��%`��'<���'3~��H`����*P�x:K�0��<���x�D���$�4 �\ph<Y�-���1�eY>6C�R�F ]>L�
`]�%L�!�a{��܍)�&�)�A9-e��c� �Ұ<Qs�C2p_�P��'��1��u�݁P�˸7 Z�5�L�E�!���|jfM@a��)v��&@�*Y�'R2�ȗ� %V)�b���-)Q>}�A7=�)*l��#k���7D���g��	�|]qNQ�+��ɱq���~ڡ�Pj״�ű�͜��T�>�O6���@�@�.=�T��E� UzR
O�Q��!I�^�2�K�`�J!�A�iNmѤ�ĳ,���:&/Ԣ�0=�U'�D��<��Z.�T��Un� ��GQ�k�`ɨ�,Fh~傣IG-Bt8 ���Rq�؟I��Q��`<B�i ��F�s�fΐTZ�u�'�:�B��$������*6�����Ʉ�Z%^Uw�݈b��{w��nf!��e}u��.�-p܀�ڦ��u.��+�Y�\�"���oOD`	���|B� ��F�P!,}�ep1/O��xRb��:V95��9 &|TR)���I�
Wf����h�<�E�bx��j�뙑8LV�C 0�̬�`)O��A��J����CX���,�"M�5�˴B�i�¦'2�C�	'F�B%���C� ;P	�r)-��PB~�"��ӆ/V<�d�R�g�t ������T�K��R8B�|�8P�ؑ�y���>�:���
�@�l�o�=O�,|���#n�,���m�(������|�LT�6� &#��9��Y���Px�b+kR���T�nd�p�'��F�_�JOH9��f��eT*y��!k��L8�I@W�h��c�[����Đ� V�C�M�`qJ#���69�!P��XH��Ɉ}��P
�'	<�x�W8eI�R�4/����I<����jX��˕��˔���G4N�mZ�*²IDlL���>!�Ě=p͘d^� Zq�@/�͛Qǐ�KE�-���7�X4)���x�o\�<t	C��Gm`�8t�ٮ��x���0r�p@�Iš~t��1��_��GV�\�g�YN؞���Ӱh�pE�ԯ�
p�A"\O8����;c*�|��'�U�A��Q��*�&X<����'dЩЌ�?c	��af�F�S��H�b�^��ʤG�tf��q�d����R���k5 O��y�*N	dK.�`�D0�����G�-�y��2~	��
/fa.��	��yr�4UD����/+����IӮ�y�Ϳxs!q� !E,���ybh�P���y�Ԩ��6�yR�O3J&ryJ���!M7��k!�H/�yr���M�x���o�4�d*�Ó%�y2��)W��;��I("�aw,��y
� ��tJV�pA"�cvÚ1|욈0"O����]I�D���(�d���P"O
m���
�^A���^��E"O zϏV�j�8'*��$��	�'"O��#%ݨ�ֽI�*A�-|�X"O
�@B, �����º&x�=�"OĔ��J.S�D�kw�X1PQT���"Oȑ��b�gs模 D^�t5�Eӵ"O������h$�����5"O��'"�=�bXے�ݮFr�: "O�%S���� BF�rs�K-y��S"O�=q�Ǧ0c�I*������"O��q���7�d	HF�4�hI`"O,�Q�I]�s�(U�5V�+�TY`"O"q�$��MSV́ � ��H�+�"O����E�&:68R&�22���J
�'�>rSBG�{b
��#��9E<y�	�'3"-��Z70$H���l��6�J�	�'<5B��ʢ��YPɁ�I:�1	�'��	���4@И��wJT6s��!�'��p9�K��8~��j4���
-�'R]׮�X3&tc ����t��'������7�̌�N2y����'z�݀�	#FY8��͜�l�*���'x4��C�?�x��H�Xq$#�'��=��ٴhN ر�ʀd�����'���҅��'G�������P���X�'l|��#�T���tφM����
�'d2��e�$�:e�dlT"Al��
�'�N�x��T����D0T�&m*�'�! D;^y�����ؠqtlH
�'U�D��A�j�rE���(�ƈr�'
�0�4+�oZ�����%>��k�'ɸ�tJ�5��� �	��~���'�P��S/`xZ���
�8{'��J�'��@�'�5�da��(s@-0	�'g��"g��r�X��R3&ft9	�'�x!bA�*(�0%��_���'񮽒��9��=9�	S)b�@���'��<��I�7�RD�q�M�u�|�K�'��h	�Y�q,�H���i[����'��hpb�E7����T�ԁ�@��'@8G$ŗ�z�+�����	�'��5�n�Z����vj,\ͮ8�'�֡���A&.\YFDO�!*�k�'��%����O���Tm�"q^���'t���$�Na��)G�X:'���ϓN`��9g�z�$Do�i3c΅Nt�������z�!�D�r��� ض9ojuk����މ'q��ʖ�� ���	��
���B��bJx�Pb�E�^W!�ā(�z���e�xLK��/�F���'?����*SY��>�OdIڇ'^�~��88�Hݣ2y2��AO`E���C *��8B�Đ`��hsC�(�0�9�"N� pL��ICM0�P��	�Zy��N�X�?��E6/~�#��X9l>���w�$����]#U��0��K�Ԥ��ȓ>�q)4�p�)��T�T3���'����%�VJD�H�;娟ʉJ!nά8���foX�42���"O�9t�-wZb��+(��k�`_�E�L�b��� �$�B�;�3�z��e��n�"ycWB�qEhЇ�	����ǁ�=4�hY�E�,��JV�����-U�I�Q�˻��|��;}�x0�l[���g�2�(O-�hS:~�dxb�\��9�
�r�V�X 4v�#��2~H� � %JE�<�uM>.o���GU�C�4��A��[��ۂ��zZ!`��ҳ֕�50���thпm_�P�KރA?>��F�N�<� �iD.��q�diU�@W���&B��:�MR���H�EMn-�TN���(O��a1�	J1��P3F�����'�!���ȉ	��9���>s�u�tJ��bU���£�0��K����N��i9���A�#a�w|@���ՒA$���?IrHD�)�I���+�6���	\)&�@ ��z�h90�.ݑX��у� eVD�ȓ8�r�k��B�7�������s�t<��<c�2���~f^tQ'(Ƃ;�v�?�`�wx�
�C�0:�p{� �<sI����'Hf�!u��Z�h���F�s��W$�S�\�� I5(uv�C�,�vHd�I�]�'���E�^�<ى�&߿Gd��דOu���W�Л���*ċ�9�"T�ER�!�ty�fM�;"Ն��#�YM.�9B�'F>aY���1�Lo�� �H���{J֑M-��Z"�
!+��IІ�~�~�B�?U�0��30�k��
�s[��z��3D��#�Hs6��P0�ںtW�=����&�=I�cY����#�E� y,
���)_	�y���y���$H̶k�H:��
8�y�#I�:��XY^DѸ�o[�d a��T�P��Ҭ�=����fӄK��i�/%�*�d A��&d\0��
�r$��뉙�]�/�ڑϪOZ���A��i�����_8�∲4E�+2$@��t�H��BN�:>��б��g�L��=Q�H@2@�ȉ���_wR��) gG�4S��\��fo�,>6tݲ3ᓹ�)�F"O�A�wM�/X^�AAP�0	�-ڱ{��y�b+�A~H t�̃.�����i���y��/uZ$��c�6q8`㠈 �y�d�E.����۲'�\bs�P�/M�mY �;}�1C� K$4���ZwX#>��f�k� 0DΒ:�v��e�ET��$���W�^�R\����b�A��
�:��V&9|V>9f�U���Đ�b���;Y#,�T1��4
��4�v�� Y��a�G�-§W|�hB���m���;�阴V����HD3�ȣQd�H��EWZQ2	Ҁ��4rL�4
U�)���O�\p3lE�] }٢�۽P�^�b�"OT��e��F�����1O�r�	�"O���#B��9Ō��r����r"OF	*t�7d�d����!'��xY�"O�Ѣ���U�*Q8T�Ó7]�3$"O��R`N5�.����l�p�h6"O��-�:  6���*Ւ6Ț\�0"O)�eE�%{~l���E'h����"OTI��)U�< xX4�b�r��"OH�x0m\���K�U��BR"O��U�D5_��8��*�h3t��g"O�\;���Rڸ)rž��Rw"OT��39�@�х��$�"O�Y�
�_H𔡳#
�Y�X]�U"O�3�Ɉ,4���P�1Kwf��"O��.�^ ����~ ���3f�!R!�IcuV<"@ᘁZܼ�v)>7!��HN��P��˒&J~��G��L!�S�P���Y*�5[Eϋ�ed!��&�*a��O�/��9A�/V!�]���t��v��K��WiP!���	�8����8W��a*e��9L!�d��S�jl@GHC!e~& ��E�"�!�$�s�<�{�j�Ok���0�825!��ӐpM:��䀶VP��qDK
!�>��z����%`Y���P�'�����G�s�	s�	:H��'����jſ%�"�Y�+[91>�8��'�|��G�J_*�B�*�-��H�'�0��e͆,b@�b3�M�q�z[�'�n�8�:y��h�H�v��Yk�'�v0bu�Ȉ9 � �2���]���'�L��"�!Hʰ��P�\�_���)	�'�dL�u� f]2<�w䗨H�����'l|8���I�(��I�g@9]�2Ԩ
�'�(QKT'�#ix������P�
�'ˈmړ#ɏD��p���p.��	��� �m�v�B�X%����e�t�V"O,�VOK�@��Ex�n�!�H�"On�6�A�R��#�lɘI����6"O�i@m��XJ:�w)۬i��qc�"O�9�$=�u#�R�|�H�w"Ol|����5���ǉ�Mh�}��"O����\������X!?%Z��s"O���V�9r#�c�e߿a�h�3�"O.(*d�Ͼ 1F4�nł:���I`"O|!Y NW~��
�L��T�8���"OU�Ɨ"c��	@D����J�"O��A�%40E�4E� �z�@c"O��S�ڧO��!1G�T���g"O�h�k��x��À
I00�*�9�"Oؙ�`XQ�>M�v)��-��d�2"O�h&d��8��𚖏P)���"O*����\�e�x�F�wpR�"O��BĀ����:D�͢ �,ē�"Oz�0���U�����P�4EI�"O�(��dO*fȸ�T�х5�\ d"OX��H4P���E�r���T"O�4k�C)9�����c�!r��*�"O$h���S)}�ج�g�H6���c"Or�E��:�x�ϗ(���j�"O�({p��'i�$+��4=	<��"Of�'	�C��pZdGv�"i�W"O�uW,��f�(��IΊH3�K�"O~�c@-Q�o����%�;(kg"ON<���R�4�ƫ�u�l�C"O�Z�?���B�����ѧ"O�\T��;Y�3�-ʺ@k�"Ojyc�閟Mp:�{�#P/s��dX4"OPUs�(Q|�1IG�C�V�"4�P"O�I�e��vJ�,�e����P:�"O�A�#ėO��y��`�>`N��"OT��`�B�5T$A�ҙibm�C"Oj��e�gJ�  �S
��B�"O^�GE�[��{�f���6�6"O�\���� SU�`#A�X |�ȃ"O��@�Ԍ{����ЁS�|&
Њ"O�٨N�=Tx#Ï
$o�8�"O
 (B	�k����ӈ�h�,��"O�j0G�<����ܳH
\��b"O�����H�h#ɇyT|���"O�#N�hqD�H�bQ�[[�j�"O���vJZ�OE��x��T�J�ny20"OJi�
�6��qg.I
JIbq��"O��҉�aUV��G�z�xu"O�10�)�+ w��C&�V��4��"O�H�������ⓗ^�.�8�"O��(dMƏl��Tj�m���r�"O�8��A(�H�IW�;$.��"Ot�h4�	[�)30g�T+""OH��"Q,1D��Ck�"-��"Ovxq A���Q�wj�I���"O�%zL]�'A����莩��"O^iڡo�b�:���	$w�F5V"OL]i�٦+JX��F�J�J� &"O|�����,l�z5M�M�Y��"O�t�I�%S���BxԦ���y�5D%�)�Ç�B<��R��yB�w�%�G�^F�rI�7�]�y("�z�[�%����.Ў�y�%��QTj&�zܸfd���y
� Hp�W��PLՙ1��0B�0���"O�\ 3g�-2>T�����&`��ܫ�"O8��򊖃iL.��6��}b��&"O����(~h���YS��q�"O����)�J�!�LX�h3"O4����jh��&D@"OFD���0#�Q�i�<�P"O���!KV�z�$�b`쇩�Z�d"O��)��4
�>lX7��Hz�,C0"O:���j��
j|zG#��z~~|�0"OVl�!͓�c�4���#\en(���'uxb�MI�S�]��J�~�l�c	�'fb}s`I<\HL�#�F�b[����'=���4��4n`H0�I�P�Fћ
�';��Q�䓯H�� �ɐn�t�
�'���!$d�Oz\�Xp#L
��͂	�'�Dj���R�7垛��]X�'$�2�F�,m�@��ֈ�R2�I�'ЦlC%P�'d���%��<K�Q8�'Ю�ڗ�_�L2J%�GĊ1tɣ�'%��q�_=h@"��� 0O<]i�'��mבD�`���#/� ݫ	�'Q��3�׫�ꨫ���>�KXs�<	q�@3|L>@a��N�tdĨ�AI�m�<M�Pe.ݙ�$��7���H$�!T���Qa� W���0s�Z��\�zH4D�ڔ�K>U�,�Z�6	�@�O�y�AP��#��� .ܤ�:�j��yr߳v4�"�����ܡs�ч��dZ�S�I�U-F����|!v��p �7���#Q��бƂ��S�ɠ<i���cs��%eY�V�>�w� ܦ�jdLN�?��(���1?E��l�"4�DgAY#Fyȑ��=[�T,JS�
$q��'�a�����r,���ī�ujdf�܈[��� גx�9�a��(n��e3c���n*�R�\�O��[� P(�\9n�a��,��Aa���C�b���s&`ȵ��$��7��T�ԟqOX�9@ԩ'&(*��^�M]j�d�i� �2���ӝ�HT��4|x(�eiǑ-��aQ�x"�Ο,�SI�Ot<�b-^kD�*1����8J��pEB�O(�y0�O�h4`qlܵ
�ܠ�N	Q�*���'�!X��uK��BFɌL>�x��L�c�`�@�#��hExrJ�yȐoZ)v`��bB-�?��O�z���D�"@L��J����2P��@T�1 ����ሄ�.ϛF&
��0|Z�B9hiT#1K�'l����Zu�(���fU�����CpDcXwQ?�H6ȋ�m�r�L z�~%9���O��޴|ր-
T�/���<%d�z����2���У֌ L�[�4P.X�C�U���O	��0Ј�:e-�9�T�Ql���`���ڬ[��ԟ�c���F�+bi���
M{�h[;jl��}�����Q�_���d�۔D� �&�qzUGx"n/�΍���$h߈x�G[�?^�$���ϗ'���SX?��=m�Z�y@O��	�]���\�ɚ	�5�?�~R� ��HU�ݳ��K�P�Q}����O�>�����!ɾER��Ъ%�-2C�O�|����j�i�%K[_��� ������\S��%��;j��Y#��d6݆ȓq�,��8<����%�[�:A���ȓΌ,`��.p�$�R�!n0�ȓ�� k4!�r8�B����ʅ�ȓw�Ac��|J)b���N�م�X�-˄���HO4����	�,H���r�isD�إ�&��բP�ȓ<��	)���B~�T�W��8�l��ٶu���vq�{a�:1�C�ɜ+�`IKv�CC�Zu���mTC�.+東�M��T��3�eÛRL�B�I�}*P��3N*w���gFvZB�	$��#�ʒW���2	C�X�C�)� s6N�:n�nȣW����P��"O�T��)_�Q-(ř���b໕"O���eN� �Ɛ��G�+� ��"O4Ƀ�b f��K��b7@�R"O�8 ��']����N95�0�F"O��rD%F�Y7Vl����h�"O����ޒx�X
�(2"O���+� D@��ԨR(���3�"O.QZ���
BI$�eG�4��T�w"OP�QC��;Y"��1GȦ�R�0&"Oh��	�����+0e��3��ɺ�"OJ|��.�o�T�a�� ���:c"O��Z�`]�\:�����(5"O\E�,$����U�Ů(��H�"O����cF�rt� �Q���!�%Y�"O4�ST^�\{�0BR��^~j�Cu"ON*2"�?EV�%�K�s@A%"O�8��)B�S#�A	��OEj�a�"O�@��d�vFİe�'$�l �"ObHQ�D`�����B7�0�"O�X���/��Б6��v�)@"Ob9r�a�$bJ��:��3#�YY "Ol��FeV�X�7!�3: �W"O�x���Ko�p���(��1r!"O2��g ��|r�<	�)�D߰�9�"O�� r�2 �󶧋�pk�(s"O�uk5n>�pPY�fI(MУ"O�x�w��Q���&D��Z:�u��"O6q�C��d�����ZDz$p�"OH��炨L���k%��74C�,k'"O�M9　�:����6C���v"O�A&@�pϢ쑲�Ӂ�ހK�"OD�I2)����g�!�����"O�=b�cT�o@L��b`¦����"O�( �>3�&\`�O���3"O���`�&)Gt�������"O�%����Z��#��p�x��"OFY@�֎���p�"�E�R�S2"O�hR!�		kj�P�o]-4�(��"O �c��X�9~����O�g,l�r"O�Ĺ���7?p���S�@��q�7"Ob�yS�ȇ)�R��儸z��"O��"1����L�dؗW����"O���W�_*=���#�B� 5jr"Oą��ƈ�$�c[�{|N�At"O<a���b��@�oԙd�p(�"O��4�O�|Q@�$ը��W"O�:�E_:k��E{`�(9`�h��"Ol�� (_� �T�1�$F����"ORXr6�_57�|se�)�P�"O�,B�A�R�Y���&v
p`"Ox=yq��2���I4��6e�t��"O�-����rʚQ��J5+��2�"O�Պ@B�F��ƠϣV�@|`�"O�*RL�'�$�CIɻ[yt�B�"O��y��ѤL�!���)wr�|�c"OȘ�5�SlS�*�I�a�01��"O@��� ˍ.��<�T��6^��ģ�"O�X��к�ʀ$�:JOļj�"O�4Dә┼S�Ś7"
���"OH��4���B�rA�Vě�&,��p�"O���v��|��Ø�>�s�"O�SoS�*�e�f�>)A0�i�"Oh�y�,J�L��$8��iY�<��"O� )��ɪS��Y2R$�S��Q�"O�H@��Y�w�n���Hƽ{��i�"OV�"!C���u�[V"��@Q"OF��dO^#v��(�D�λKH�&"O���F�d��#�Á���#"O,���H�y���{��\���D"OL�;�d�J!�X��n�:ܙ%"O�CiE {t2��O�S�R�+1"OL4�e�K��y��M2,����"O"8�wdR	#eF%8�� o�Ș#�"O�B���v@8,PA#0�i6"O�HjU�H�V����d�1B�z��u"ON��A�8��������_�z� "OP���E�+2/�m��#7�,�"O��CrBٸJ��[Т�"v�&hA3"O(��%�N̸�5��H�+�"O�hIC,w��A�$�L5B�4�`"O���Aײ/c~�pG J�3�P`"OjP�Q���H�9z�H��"V �a"OJ����)7m�ij�!��;�H��"O�D���-^c���V`�X��L{�"O����Z&H8SƇ�p��%:"O������U^��3�M�3ӆ	��"O�����S�Pр1��мW�� �"O ���G�#:|��$�5�`c�"OI��fM33�(i�� �7&� �(�"OhQ!� �+[дA%�-=gV!�"O�	[�-��>3�؉p�
-g\a �"O�druc��U�rH��*Tfm+c"O��t��%]d̃�)Q�\?H5�t"O���#L� �9B�Li>+�u�<�$@��*�}�VL̛<�t�n�m�<Y�o��$�8���D|��c�C�<)��@�X5���B^8r�����|�<!�+�5��б���26�2��]�<I�\�T�|y gY�v��q�r�<aqjȡK^�q�/q
��P�N�p�<���҇7���	c�y@�B�W�<��(�t�����\���`�wI�<��&^"��G�N ���u��\�<Q�B��!4	C�݋7����\�<���@8D�L6"��]ΐ�#���`�<��㎷]�0p��ôC |S&�W�<"�1���SD@جtjc��l�<	bK &B�(j��.\���i�f�<�0��1`�,�+S���`��_�<1�H�'
Z]�1lQ%����S��b�<a1" �E��y�1B
n��@y���`�<I�� ~i(�����DS&�BS�<�������:�#�7[̚��BG
P�<兂�J��Ƞ�M���0Qԁ�g�<A_�^z�L�t%��,��q�լO`�<� �V�~�0LS���"�R5�`�[�<v��[g`�C�^u�����OP(�ȓ��bíF�)Z�AI�Nr�ȓu8\#BA[�c�R��4聾O@�@��!����.*������`"�ц�7@��Cӏܯ\�\�@��{�>��ȓB��x:�cȟUcttp�@X�\��ȓ1�(j�NL44�,���J�s�b���l��P��,G�P���B~G4х�a�"�Sa��0Z��7b�XN��ȓu(�K�$^0F��e�r����Y��s�$ ��φ�NԂ�q��. 2��S�? .\�eK���( ��^$�"Op�Aҏѻ".���3��Ă���"O��I�"/YM�Tp,Ël�t�1s"O���E�-;jT	#���M�
A��"O�m� �]δ��!�,~�  "Od���Jӯs$p���7~ڨ�)"OU��˝7^'֝�rX7/نHSp"O���X_MQ���8c�J�:�"O��!��S,~�QVE�v�<��"Oҥ3����2��%�F%>�0���"O���t�&\&� #��!7T�SU"O>��@�7G�:M;7��\g|���"O�(� �=!�t$�
K����"O�� !�ύK��I�璀/8�"O�,�s�P��a��L����"O�H�e�F4 -���LӇs��T#P"OYi����+�<HHG�եVK�8��"O�(�E��1 y�u��i��fD݁�"O4) !b�*-d��!�
(@�mi�"O�b0
�-2xF��P�'�� �s"Oe����L�R�E�s���5"O����=E
��c��+>��
�"O�uR@O%>=��hP3=�0)�c"OR%��U:�By���Ts.��"O����C�
/�p`33E�0J�""O����j0и$_<����"Ol���8qh(�d�����V"OD��u��i30=8�
"a����"O����^�e �2�O�d��Q@F"Onja͉��j-�򊃇OHE"Oxqxp	�.8�<s�'�]f�Ա"O�������<��f��%Q�ݡ�"O4)��Hޖ����W��	U^ ��"Oα�5�ylX԰�eړfe �hV"O�й�û�ִ³�R8(��8z�"O�����OBA�#d��Hy����"O���2N(Y:�DK]mHH��"O
hI0��/�~�  �(7��xx�"O��K!���Iq��q�	��"O���U��K�Л���7皉�"O���u"#^n��!9z�蹧"O<���㒭o�v�!���JfbE8#"O�������T�eI�2UH�;c"O�@�O�WtYIfd� |�^,�0"O�m�"� T�ٓc<Yr6]�F"O��b�T;�J� I��`�W"Oԁ�#
�/<W28��.Ǒz�� �"OB���l�C�x�ѬB�K�j��"OH�"��b�cKB	l�訡�"O�E��A�J�ؕ����6�� "O�u��
> ���P�Q8v��)à"O�]Q�,��O���y�Y�"x��"OXR!�	�>t �%
ɩ�"OD`í�#f=�=I�A�#P���"O��I$�
7@��4���t�ZX��"OH�+w���$���ذ ͔b�"O���Dc4Y�
}��D�l�� 0"O`UI�    �P   6  �  $  �!  �)  d2  �8  �>  BE  �K  1S  �Y  �_  !f  el  �r  �x  /  !�   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dlӊ�Ӕ;O��JB�'� �aE�4_���B��O򽙶���A��#p��cap5q6�ݲxB�02�`�q��@�?5����?�S��g�ra*U&�$[a���똘+r�U���5^%��5JA�p �0aA��&�u��סx��T�'HP5"���#d��;M�g��1� a*j~Qb�k�Oj��a�,p��ZU	H�Q3��ߟ��ɟ����i�膸&���ŉg�JeH�H�쟠�I"c�a�4���O�4�T����OH����F���-1h�S>J�;r
�O����O,��<������ش$��'V(��)�3)?�Yd.��/�6�����_�'�k�!ɶ��-�"��JQ֮DT&��O�����)���?e�A�A�V����ښ<4I���O��d�O��d�O��d�O8�$�|�w���i�0 4R乥䎪Cy�ܠ��>��.d�.�mک���K���"O��M�5���?)FźA��h��LŎ e.�`,��eg��(3�B=�'���_�n����%W�J�(j�T��Bq�ۉ Kr���%�Mõ�iYT6m�D��3WC����/�4�ؐ��`=A��`�L44�Ho�,tlHD��	�i���~��R���n�,���4Y���d��3�&ϊ�[!�N�]���# .ʹ02`�p�Lݗ#Pm�%�M��i��-p&b�T�j��D qI��eOc�ġ[=δ�	��`�}�0$�H<��aj{Ӳ�m2�M�FJ$v�ą��C�L�.� �d��qʍ�v��:�n����>0�Z��i4(|JT ��?���XV�̛B�X�7�'e�ONh2��L�S���DZ�(R�S��O��h����@	K��Ms͟BUB��ތ{�ժì1z�
L���'��I��I�|"��ɅY�l�j�O��$�~�>���^�s��gm=lW���dV�f��B��!Q;����C�OT�ă\AtL��N�7���!#�'��:���?� _��c��ѻ@Ux�n�}�=�V��O�$�O��b>]�ƨ@(s�C>&�>�Yv�t��0�O�Dl�g�fHb�23�	��M�<ú�J�4���1%���m����_��k�n��i�8H�N�iς>HMu@��	���'��L�Q�4#J��2�#X�8�Og�*�Zas���`ƒe��@R����m8?Y�-L� r�%a�$�*V8�J�;ѱ�&�3$�8����iD{��9�����7��O&=o�$�H��S�{��T���'c�Ix�`� BW,�O��=�}b �5'��J@�Ժo8�8�g�u�'��.o��8lz�	�$�~����ԦRGD%	�J�-�B �� a�0�?I�g�'C�<�H�f7�y�`qu��'=L�)��]$U��ǆj��a��'!�dkE�3p.hYb���c,8��'	x����W�z�<ѱEk�Z����'͂x�Ď#{np��f�NpfĊ
�'�r)�3F۴.�\V@\t��%"u7$��	�����Iy\>-Χ�z��(ǲU���M�&� ��+�/�r�:
���8��숹�m��ۍ�� 7�D�x�TL�R'�>__�U)�l��F����D�#�:�P3	F(Z�x�uA��vVJl�c�'#h6-�P�'K�IP~�o��3��f�
��B!Y'�?a�'V~s�AI�1W����#��Z���K�v6OR6͉��O�L<�eӘ�ds��IÃ�-f��$H�֊�P���O���joџ�ͧrH�����nt�Ȁ��Ɵta2nU=l��E�'���0�����"�T�h�G)�&B-� ��H�&J�aԬ�� ��9Z���R���OϪj�� #�ӹ"^Q��#��On��M��L�q�ۯlhN�w`�-:pm�.O���9�)ʧ3!��@�&����l�afG{"�I�M+"��4��4�` �V�"Ÿ�I�X���|�d��bO�b����>�Q4��P'V�+��T���]�"�5D���χ�k�X���.�����/���y�N�_���cZ�=9Q��K��y��
%�sPc��~�E���y"��+%A(l�e��0}y����*�y�F԰,r����÷rp���^�Ne���|R
]��D�'�R�'��I�1x���s��H$�ig��m^�)�@�0�4�	^��1y�#�J�t�	/-x�2��X�)[�L!�K']��prA'˥a�D山兼^���#�4(?f�ӬOJ��2a�����i�3r~����'���,�����E����	4��n�=��݊�`��}}p��B-}x�ܳ�b�B(Dn�uY@o]�
G2�t蕧Mnګ�MkN>�'��/O��z�,ĸorMk��^�]n���E` �-�@�o�����ϟH�'��O��0eD��?��cLR�E�6�
�F��Y�P�-���+�'�D��Ǎi��Y��J�\��b��^�]vVԡ5͙ e~��뜯t�$���)�O�dc#O\�&���+qĚl7��"D��daڴ��D�O6��O���OZ�A��H�_�tԢ�#䒩#"T���*�X���a�J����Č�|��m&��ݴ�?I(OޕҀP覅���L�`ilN�tҳ%D�r&�{������I/}�Bh�	��ΧO!hd�', �.R�
�ɑ:9���� �McGȐ�/��������mQ�'���@mA���<�vI߈u��"�'�%�4��Ӏ�1b���o��0<���ߟ�K>�e65c�T9���?����Y�<a��!-�~|�)Qp�Dܺ�Ǆ\��hO�����#��Y���ҟ1��X1�+��[m�'����p�����O��'2��
�|>�dbFd� (�\�'m�h.��k���?���`������O��g�䊧m�n��.P�=�4�X�^�#��I5N!�R�:�)�'8����rT�T磃�FT
t�'�d��Q�����<Ys�n�(�{�./�<ٰe�`-�S�O6��hF* j�H��/#K���	#��D��9i�O�x�`��N�P�3 �-���ܴ�?���?A���A8������?a��?ٝw>l�*d�Q�\�:`�7 �-���*Op��_�tz��D�X��T�D�$@��r!c� $1O.A"!_�7Cax��\�#�bٳAC���	��Q�7>�f��`�'��O��+ړ#R��4☢Ty$�h�	��|k,O�jS�'��Ӳ�	_�١�׫V�"t�+O~��'P��O��OtʧHn@�s� n��1j3+������46�&�'l��'���w��0��Ȳ���I�|��Y!?F��[#�˷D|�X�vúU���'(r����X+�E���@��N�.��A�nJx'���:t��e�^*��XEy�=tu�Q[�� )�-	�Y4����iG�F�v����<�����'� 1���5{S2������|{dhks��/�S��E�j�T��Y{�HA��1Th�'��Atmg��˓J��z���dm�t�7�VaTn��e$�*,눁�#H�OL��?)�����BՎ"�$h���!P x�k�[.LR����e���o��]�	�4�*�X*_;U7��
��Ω2H��W��l���W�I��iK3KɇE�V\1�#�b�>��ɛ�M�t�i���1��T#�M�z�L��#����	��\�?E����1���PT��d���R�C/�hO�=�S�i`L`ʆ!��Y�H���ޠoD�E�`gd�*�C���Bn�?�H~�R�iw�d\R�eS1D�f��B�h�I58��"<E��k��!���9e�AR�21j���$Ԙ��"|b�*��LQ$H�z�8�BE�I~�Ȑ��?!ӕ|���ޚ;��4:��<oh��э~8!��X @ڄ���ͺ8bx%;�%�/6џ���	�vHN<r������p�%�>&}�6m(��
�
W��?�'�sO�+�X��S!]��d��y��^:�0=)gJ>��<��ΟE�"HsU�]̓f��؆鉮i"�GA
p�$�����7�ę�,�����*24��Ђ��fN�Sg�U�!��ʲ8�@��P�nѻVB:^��I-�HO>��U�[C�b�3��5"�DpҤ͓�6#���	ȟ\�	����'-�S�|za��%k� �!ʶY�zl�'H�"��Е"�O�a�NUAJ<���"H� ���74�]��⌮n'��	�eU��1$��r���q� U)"�qX�ǟ����ē�?1���䓮���֟�Y+s�X3Q�(�`W�@4�yR��/	���`)�1vOd�H�#���u��kg�r�p"�Ls��?�'=!8�%1#$}JFgA?f
pQ����O��dq>e�4����xR%��*s�Dn�@;DR�fG�D� f�>K�n�ې���䰀ٴz:r|�`/�8���[3�̫��'�����?I�i����2���f��/���V#��w��ϟ��?E�숦�(�86�S�b�l�P��ؒ��d8�S�'O����ls�)�(��	���\ #~�7�<��F�P���'�	i�4�'���4b��N|��h��;�Aj�'B2j��&�\Y�3�>���OC���P�\.3�Ӥ"�n;P�����\��O�s��qdo�kp�(�����	�q�F&�S ��x���'���$5�\��X妅��4�?���	�"%bD3�n܉}0�6��`��'��'�ў���r��ۧ�\�[�(R�B
�z�Z�?�ÿiW�7�-�d�5(:���Ȟz�ļ��շA���D�t��3�Lzr9(��Z�bsh�\,J8ؔ�ȓ���q֋�G�l� X�,ܙ�ȓA��;b�� iv]i���&M��ņ�r1����Z>p�8=q!��\n���Y�b(� �&�f�YqA��F<��_��P�i@Px�R��+pp$�'�Ż�>��հF�vϣS%r(w%C3(!�� ��R��#~B8�{���%#K^�0"Oȥ��$��T�,�٢�T�X[6�c"Ov`À��Y|�y�0���WG"O�eZBL������ fc ��%�'��y�'�ޕZg( �"��ز"	�0W�%��'������	E9��2	ǩ2���'�`		�����Q�C*0����'Cj��s����\���S-����'�Ru��\0�mkE �����3�'m6 y��HT߆��⊖2<b�����$r�Q?Y8q�A�6� )ƻ>#�y3"�*D�4�i;x���FQ�.	X���)D������S�<{�M�6�D��(D����N�=��5�2N�!���"�&D�𱑂��U���b�6:\���b�#D��C�^| 0Ys�k*az��VF�O:��)�{��@�E�>^�����ߺ]
F��')�s�<3C�Q#	��]�lX��'��$r&�(�\\:c��>׆���'B���쎢B���5:�^Tq	�'3�c��E�Z��0�
.�4(	�'�Ҁ����-rx�R	 �Dल(OH�3�'|�5-�7j�ق�>����' �Ab�N�'/�28��đ96L����'�>m�CF%jy����Ȇ E�%��'Q
���eq�ri_H��G
M��y�mS�~��Q��J�v�p#�����>�1 g?1�1|�@[Ad^��ȅ�f��X�<1�(H�,�����j�;R��|ٰS�<y�G��_����IF�,�\Ia�Ov�<�E	 ���L�qd��i��Aa��n�<���(���a�M��<�@Dj�<�ւö\z��s&T�N`x7j�N�'�DH��	�I���;s�Ɖt�"4����!��F%3@$�ro�1�ȹ��U�<�!�D��$NYq�'M�s´�I!�Ϯ�!�՜3�� ���_�-P���K?�!�D��a���y��D)UA�L@K��zA!�d��jh�J�o_;8��_�=�	�%Q�"<E�t����as 't6F��N
S!!�^>'jI!�_�[-48[�i�(Zo!�č��JU����6'd�C�*S!�$�2C�l���U?=�p��hĚJ=!��L�P��88�-`�'��*%!�
N��)2�U
۞4��e�3�	�(�����{T@A��=v~#qD�)W�!�92nV10��,qG e
���<�!���~^N�x0c�*���g��/<�!�ĀJT����8	�.��4 �=_�!��% 9I2n�*a����#��}2�@��~�$�G`�M2��]"PX�|3�����yꙥ�J�J�^/C�e�&���y�Ě	}lh��1:�@�g�A��Py�J�}8xb�뚗/����X�<م�֔|l�T[t��R��T[P�_�<�P�ͽ핓HS�y^��3�U�vuў(B�K2�p��0�%Dr�:|Y�$�,I�ȓ:A�}�@㝲*P��y���U�ڴ�ȓQhn �`��2ƨ���AX4��ȓ6l�Y���-|ItM
a��> ��ȓ
�Z��DJ"
�0q����%���f*�<qW.�'<lr �S(�2� ��	��"<E��$� �&5���ՖIvv ��X,X�!�d�(fИ��I�#r zd+�)w�!�� ��:-��*�&]���؀H�U�p"O:dA��������b�Q"O��4k�'|�t���萜�"O>�!"�)��E�b��!w����X�1��5�O~� tȁ2j̉�JZ�k��Ģ"O� XQ"B,�,h�uIH�3�b�"O�!z�*�|CH"���Y�eR5"O��"�Ǔ0�P��X�I��9��"O3�c�M+�HA�)h32�'=d���'ɠ�;ǨH�պ5P��_�i�v���'T�U��22��`���?5,���'$l��a�:d��s�e�4��48�'�9���νM�,�ۂF�%x*6��'���R"�1DA����e���'��q#��by��CA"�_]Υy��҂ #Q?-k@R�zT	�_s8�� J'D��!Do��He��r��2��q��%D��3h�3ku% p`XL���S3A6D��ssH
'�4�q��ԩ+���3�4D��Z&+�ԈUA�D�|hc�3D���Fxz���"N+N�hd�Ѧ�O�=�w�)�' f�,U-$�"Kދ�b=��'��$�Kٞ+�<�#r,J�]����'����1��U���0�O���`�'$|�BrG��'�$0#f�*Oo��s�'�8��
�86��;D��NKFx��'2�Q&!̸sn����	�LF9-O0D�U�'M�5A%�æcպ ��M�#P�&���'�����m6`�BNG����'��Рh
�ap��!8%ֱ��'TzЀ��� -�����*Ȣ�3�'�$t�uD�����阚���cv����KA�e��CA�}�ę��ц\z����G�ܪyt@���C�-S9�ȓ �fE�N�d��u�����$��*���H�j�e��A��J�4�ȓ~���H0䞩"�"Ur'S�
�b�ȓ2,
4S�k�y� �"�
�]$��E{bH�4���"��s�O)z����LF�d� ��"O�mq��ҭn_*�H0��H��3�"O``��"�$cp¶k��(�D<�u"OFad���^b�p�v*�Ty�` �"O4���*"�����Hf{�!��"OƬ24#��cx��`�:kĺ���'̬$��ӌ(��QQ��m�
�'*�AX͆�D�9�[wv�k��X� �ȓ��e�WhyD�(� �:]馹�ȓ4�h����(:&���h��np��ML)آ�C�|����M��m��yt�t�Ө��$[���*OX��'l��	�FE���A+�N��g��	b<Ն�B�����F(��/��{l@Іȓ{?:ԡW�D�{���������1��}���VFT
 C$X��*޷}�0ͅ�@��Mh�Ŵ)�&��èQ�U����	*
��I�F�0��?� |�!��HC�I]���0�N*tP<���(wQrC�	(/�؇LίL���X�w=HC�Olx�p��$���)%���HC�ɑ�	 G��jn��S#
1�(C�	o�^rf��3���F����=�s/�U�On(���e�e��ʧa�/N�Q��'Z���'K�RH(�ff_�]�S�'6ȩ��� D
Q��Y3Y���;��� ��{&�/\]Z�뱭��\�9"O�`��
H�t�e/Db�2��"O�5�S�V�%M~l���`�:H���'Z�h����S�F�h �"B������@͐2da��>��"ș[���S��f;h���R��Y�/�)�
�a%Zs�@ ��\�lI�`�C�z��Z-fX���A����쐺B�<��Q� (yT�p�ȓ;��P��߰Cp�b$I9~��|�'<��:�l	n�y�aԈ	!8x2 ,�go�h�ȓ.2�b��[(��(�5�tL*U�ȓT�� c[��2�Ʉ�J�A$1�ȓNx �e�/a24��.XyB��ȓ	�YӤ��D"�}��I
jB@5��ɵ����$D"��`�ʵ
*�%�Ǌ�;��B�ɏ.zF(�V�HK<�a��m�1<7�C�2�Q��+A�j���*% �)W�C�I>Mn^�1��`R^Y��P9#�~C�ɖ �eI���=V�X�)�
�I�C��Z<0��C��V�P�̛�;"�=q�o�p�O����g�����j5f��.��
�'�.`yV���B�c�+������'Z����N��cc�K��|��'8U��U�[��E��J��:l��'[NI0�	T��lʶo^�$�Ő
�'����0.^��"¸ �d�5�F�Fx���R�^
�ࣰ ѿ�B��ӫko�B�	�
��g!��	��\#�җ�FC䉭K��c�B�]/Ƽ��Ak�B��:a�|A��޵Cr��J�d��N�PB�I�o� ea#�ε��I�PjԔxO`B�$B�D ��Un��mK�G�`����{��qy�d�=��to	�u��'����v~d�SG�<.��}H��[����ӵ1d��'n�ԤLW�����4�8�Ieb�5�4m�;Y��ҷn��w+��BQ21��=F|"�ϧj�
�*�h�*X��
t�\$s���]�	[� �dc��,7`}	�#�*8�">�aKޟ���I�'��� 悅,r��!%��v32�'a~��֯X��m3�	1L�)���-�䓌hO�IPy�D���@����".�tIڰ��DȻP��l�4-x �	k���c����'�na���2u����o�&6z��D�'�J���*{���R�`�[�����[>��|bCʚ="}��:�m��@��q�OD�<� ��5D���:�a�@h��6�'�x@%�M�z}lTB���4͓W1�d�O��S�X~"�A��ق$��>��`J�-�yR�F:DM:@d	pa9 E���'6RO/��|�s��
��0����%/���Ph+2������?q�L&x�Z�'�?���?�@��4�����W�D#an\𐵀ָ{�IëO���pd
��
]㒙?#<��Q(JMTXAf`U�R��%וm
�	�4R����=�l�g�' �D!C h�l��a��>��y�O��"�'+��I�<ɑ�)P4t`����T,�k�j<��yn�\ؑhN0�-���͔A<ʉ�	:�HO�	�O��?��q��fY�}5<d�qGBo���A�G
>klt��,�)�?���?���
�D�O0��h�(�oM(v��W)G�(�HLh`�[GR���F������'��
�o@��yA!�[�|��E)�U�ʼ�e�-xz��'�`8��3�'̤��w�V����o�-���H��'FўE|	�J�����L\#k�u�wL��0<���8�Xd 2D�'���h1D<2��	��Ms����'0
	�N?����ψ2Z�b$�B!�8D� ���0=�'�A�S��y��7D��q���1<ĜzAD�do��B�f5D�@�C�я ]p���#یs�E`b�&D��r�cАU\���؝=����>D��cQb�n����&X��� �;�I ��#<���Ũ ��NC��{� Hd�I��"O>��-ЛJo4hQg���)�c"O���Ԇ2o~�$���A?s��B�"O� 
$��_X:`�L�HR���d"O:2�Q�e� � ��Z2S�8`�R"O��ѡ_��\���1rX��3&Ʈ�O8�}�'B|`F�0�x�2�(�4�&����pP�L��>4�xf@�#O�̅ȓO*��Aꇕp��<�sL������1�搑�D�Mz bO��,�ȓ[��E�A���N�E�#a����� \+�CՖ6Dd2 � u"�	
-ê�������I�/�@�ٷ)ׄT�!�dLw����$W�Y�N��t��_�!�dʈ�5´oF��M���|�!����H���L�s��ZE۫]�!�$�. pQ�!䁹{\��"Ԧ��sџ�K��F�M�J>	�X�x��FA�;'��|���,��$�O����O�� FX+N�`��'H��R�n>ɢ����/�L�X�G3Q��qi ,�x{����2%�,�U��%>"� �V��,2���p�RR�\D���5b/�8i�&3ʓi2u��ӟl����$�'!�,1�*\��,U�1�D�H����ٟ`�?E���^�TP��>89�����u��O��=���i��7̀z�	���T�j	����F��r�˓�?�"B��?������O��tV��'eH�f���v��w�D�Y
Ó�hO>p�ā[�1��+V,B�oը�Y���2�'�1��q�EX��*,D��� �B-�JV˦��Ʌe�H��abZ5�	韘��ߟ�ΓԢ0(ԥ� L�5����?B�TI¯��Mc�ז����yb������{ę?��%O�!��땟,�8{��Ǆ[<Qr�'��"�2o��a�a����|���p̓t�,�����N������D>��G���,�� /$��I�<�Ə�Xnz�A ��B�!�s�����DX�|�#��'̍q���?��*Gz?�S쟐���?��ɰ�d�c����B�Hj`%�'H�:0���e����I񟸂D����K�����+�uW��"ZM��BĤM�E0sc��4�y��Ĉ�?��n����O�r�'����V E�9�@�z ��U8I*F)"#=O�LQ�'��at�A�I�<�4mn��E�4�ᔛ+��i��!��2�������M{�'w((�$�i�6�Q$���?e��J�j��+A��^}A�c�4�<Ճٴ�h��'nl��?a�'�?�'g�}��O����t�A�!�l�E�&sB�y1�i�$0��'��	ޟd�)�>�CDذ�f$	��_�#��A�n[C�<��FR��+7n�!a�Hr�������	��t�	ٟ��	ğ�	矬�	ޟd �fгB�,+r��#���[$�W7�Ms��?�,O���=��p����KI?�� ���m쓮��(O���B<�Z�&
zw���"OtӲ����L3�	#&hz3""O؈� �w�
�ꡅ�)��I��"OV���(W�M
S��I����"O�H��	��Hc��=OO"h�p"Op���޸:(ѹ'��U����"O�d����&,�<r3�_;Z���K "O"-�w�1�*$j��F4d�D�0"O&����,k>�drv�I(@�Ne�5"Or���iΐR �`2�R��JĻf�	�HO�Sٜ����
>�$����C�I&|�Q�v��v`EHB��u?2c�`�c�N�Z�y�ۊZdH�	5@�1��� 4(�m�t���ML�`����J�S|�M"���>�������J�TZa�9h���KA�T�6���E�o>�cV��$'����\).�T5cV�P,�`0*A)�����6l/��h�'��>Qq���P����*�yZ��Q�),PP
M3:P�ȓV/���"ᝥfh�������V{p��]a$ikU��%3-����o�V�݆ȓD�d��O�, f���]�m9<ņȓl�8V�+CD�	F����x����ǵm��.ʂ/ƈ��Ym����F��Z�!W(T�>���t#��a��y�ĉ�1j\�_����ȓ��X�&I�A^�z�I� Y$��?���c��=d���M�G�$����k5C֨d�
�������ȓ}PTp�F-��4�1	�t�h��{��l{�P�lvX��5K�Y�<��S�? D�B�/F%�eKe20e�@I7"Ox�qw��,����ڿ[_�3"Of�
�`�I���!Mh�"Oty��Nr+J�G�Q�{���"O�q��e�.!�@0����W��e��"O:<jG�Ϳ+�B�sd��
�h�T"O�Qp�[���ԂG�%��"O�\R�
9/�*��T�ϗtꬔ��"Ot	�'���A�`@LE��t"O؅8��՚V�/O4U8Z�"O��ig�U�+J�]�f�:h� DJ"O��梏	#��)�兿I��x+E"O��y����脒�d/G����"OD��������Ą�=]�؅��"O�ೀ��toD���z�H��q"O�3�`S�vVd��(��Ak�"O8M*�o@���pۄB[B��f"O@�+��O>{yL�ۅ Ǵ�ܚ�"ORx�BF_��x�A�Y�>�y0�"Oʵ�Ed�5vDb&N\�(I��"ON�����|+Vj�wņ��F"O��ұ J�D���i���K4"O����C%wِ�d\�(��l� "O�c5$G5EQJ�����(ӊuR�"O���)Y�CB  ��G��l��1"O������.!��iE�K�@�����"O�U0�&�&
�^�9�ǟ����2"OơS��I��Nd��K�-M��0u"O�� �	p�b���	� <o�#@"OFT:'��!Z�����[�{bRd��"O`!QV��O�h�T+ӐkN�Q4"O���'�5#2���ק�	Hݔp��"OT9���=J���a���1�*��P"O�|��o�
f"U)fd����c"O��p-�'��Y$F^>"8I�f"O\Ÿ3��_;@��H2��)R"O Փ�a����q��&	���1"O�둪P��բgfj�yb"O�Q����vO:r!&P`-�""OL���V8e�p@��@�f<Ɣ��"O���&V*pv��q���g/���S"O��D�_�M�ҭ[EQ�Y"Q9�"O`�� ��	ON��j�i
?��]S"O2`�BKM��W)M8hg�q!P"O��0A��Z1�mVBC-����"O�Zt�A�dq0T{"�v�N�3�"O$���>Z����ͳ�(�jS"O�˒FE���e�@�:�Ѐ"O��e�GR`t�Z��2w*�%��"O��*C�Y�E�j��%@�>�,�2p"Oz��d�/
q����Ņ~�n�9c"O2��c�J�Xz�;BG@�4�,u�"O�`��f�Pq�p�O1'�l8�"O���`'Y1Ί3�ܣ|`�3�"OĐ+��Hf���i6��:�T�"O:���بt�`���!
�NI) "O��S��VP4q@F�c��8C"O�\¤)��PQCOD
b�����"O4 � J�D�(���\�9�2U"Ol�+��!m,8�I��E(�UK�"O��X�,�A���#.H�0�"O(][�O��l����U&X
z�2%"O��J�f��-� �PsI�5��!w"Ol�CC �q4踉�H\��ò"O� �#槁�OO��B�4JU`p�"O:*���ӚxJ�mD��q"O�DЗ�	���ɛB]�"O�y�ҫW�@HA�c/�8@� s"O�e�䡇0s��=Y�K��p'�`K�"O��p㆛V�r1��$�l	p$"O�0�Bu�H���"������"O�d��ZIF��a�����"ORȊ�־�uR HIF�R	��"O�d�4��~%�9R���j�~I�W"O������g:$H���X�3����C"O��*��p��@�ƍن0h��2t"O�����Z�{Vs������q"O
�����k48�tP�4�P�SU"O���6�J�[{�򅕬q��`"O�A��Z�)�������Xȉ`"Oh� �`ƜM�(9�&c/z�D�*3"O>��(»�>�c���o&�!�`"OPq��2�
5 �h�(�W4�u��6�N�s��+Y��HR.�)R��a��|7�� �)W O�y�R�ˌ0�.���U�1x��v>����Ā�x���g�5�s-�4]h�BH�	V(5��s�6$Q����a��o��w����'Q�x���9i�I4��sb����'3j$@�S��]���PrI��'����:+J�{X���ʰ��`�<I%�8Rr-��� ���z���\�<�g�J����ԍ6�l��2FY�<���MS��z�`�'9�ՒPPL�<�3i�z����M�bO:���B�<�׃L�F}�l���Ut@M9�#�~�<� EG�d�RtQ`� �x��he��e�<���ѓja�tk��ٍp2��Ŝb�<�2��
��P p��x�A�	I�<�!�5�X��B�ĕA ����	B�<���ؒ<:��`�FO�Hw��KN��<�T`���Fi�c�p�� �&q�<���t�68�%�֯O��-ZQ��r�<�%$O�^�����[2t�*�ZG��p�<	P� �]�D�B��K0n�m��c�<�GD�:Ex����[�F��ud�<�v,�7w�R&̊\X:�ac�<WG��S�%��EH��8���c�<�C��]�z����,�ʐ7�v�<�Ơ��S�ā�4��)|"�1��Os�<��9N�<d�ujQ�-�����o�<�PO�"0d�-��ʐn�D����O�<�q�9g/��R�N� �t����O�<�q��.����3�P�b�����S�<a�
b�N	@�C��/�x$�G�N�<���>��sI�D�T��y����=`b�ܟ?R��6�޹�y�أ�h!c��@(7/��C.��y�ɇ(%T���`�4�����8�y�y�"�Ӷ�K.a*� �$ₗ�yR��Q����jP ]��9����yB,��@�xU����+�*g���y��(�ԥjQ"�S���v&���y"�������2DAډ����/�y�EH�	�¼����-N"�����y��hsX��R���1���y��SF��
�N�(*�RV��;�yR������6b
�@,9cg�y
� ���W
�z�)sf�ƣ]:�+�"Oȳ��ޡ,A�5@��ѱYj^�q�"O�x�OC�%m�z���%0_�P`"O 9P,Tm�\@2�Ö2���H�"O T���Ї&>�);���0\򘑀"OJ�;�'F]�l�c�S�<K�Qp"O|,���U�H@�19cf��/�0Pt"O�h���y��\��	�"OV�{Ef[)`� ��3ǒ?U�� ��"OT�Yd�0&�Y�����<�|!�"O^Tr,�4�Y��ILP��%�T"Op�����L<�k���	p"O����F%/!Ԅ�T��,p���S"O�=�!G�Tv\8"IP*\��Z"O4��抍<X|�[�W5u"�	�a"O�@ivj�3��@(F)�T@(��"OX$*T�ߝdK��U��Ƹ��"OplG��/�a�M�
�`Y
�"O֨@��nn��k�7,��la"O�K1�"}|n�H3�CP�*���"O��R�HY.sq����N�U��{A"O��2�g D̙�&�u�i�"O��yC$��B-�k���1!���)�!�D�+aQ����K�:���ە@�7u!�䚉ӰX��R��y�FN	8k!�d��.�����F H�����!lk!���u�F\�U��'l���U��zb!�d\�eM)��B�?�u�0`ݐG/!�d�8��2aN��Z��!C��!!�
+.7�liT,�;n@(�w�W�!�d��"����.��K�u���!�� �i,:���-���\��!�#BH����@�Hoj�EO>2�!��'�$�J���s�������!�d�B.v��犂�L�0� �Gl|!�dU�j��,Q�>��m��[)a��P��\b =(�j\���h���g�ZĄȓx�V4GC��j�;D��P�� j ���"
�,��pC�F1 �ȓ~5t1�%�CBЪ�U9|�~ԇ�,u��Cp8|�� ��9|�x�ȓO�����D& ZuA�3ir��ȓ��l�r.O�p�ƍ[�T~�U�ȓ�,q�	�
�$�����V��ۦ�O�}0 bff��W���ȓYy�q@��6�ȡܸY���'����g���"H���ջ��AX�'�@4EG -�CB�I|�8 �'�l`��� H�jm�Y9,$�2@"(D���`DC����� r���R#&D�hfф"��ai�lZv�P��'D��X �S���H��͌'R��q�&D�����Q�N8�劯e�Ԩ�1�6D���P.�Wr�3w$N"��؁� D�d�p���q�%a�ЮJ�Hʤ�<D����!��`4�Tە&�/A �o?D�r���8��a��	�41
5٧2�I�8��� 혳?��X����O��{@
X�(>�a��W�p6�\"O�툵�-5S�%���&}:��"O�h$g<2��@��vڄ[`"Od� �G]�,�F.ˏ.��E#7"O��A5�˳����,@�m��K�"OR�dG�A�"1��!D�:(�ٵ"OXA�
�4h���'K�F��&"O� �����ͪo_zL���ݵg*58�"O�<P�2>v��Ѧ��a�V�P"Ol��C�R�p)�u*��]}<T!b�"O�ѩC�� 4��ʴ�K�^|��v"O�@�'�� 1xc�	��j���'<����"�'Q2����� ���h�'ZH���5A�ZiR��ȱ`��I�
�'I����W5���h���6Јd��'͌a�.\,fP0�*P��'�(Љ����t]���4�EK	�'X��B!�J��Yr���d]��'�H-�D,�g�"]0�7F%�L��'Q���`�]�D̚�ڦj��9@�'�Ds *Q<\j��E-V����'���
U�]$S�`���#V�e�'+����Q;cy\�P��&L�X�
�'[����X5�� (�E}8��[
�'Ԧ0��Į=E0��J�!�I��'��0���&G��Ç/�R�ޱ�	�'MNL��ה�h�b�ퟢY)�ys�'��ai^"xƈC"# K@�`�	�'����L��/sV]C�A��U2��(	�'��MG͝�$�P)`qaZ�  `��'�p[�G��ʾ)A�Ќ^�<�a�'�4C$�͙x��E�PnK�X^���
�'#Zi+�c��-���h�m��kZX*�'7H�b�N� 0)Qj\��,)�'ޅ��#�#>���w�J�&���R�'$��1Wo���J�)'�HhbEs
�'h9q�s�a�c��4Y�'��}��8n�Z�`��\,8�J%��'���eAʥ%ޠ����EV^<��'���ק�!E��QtIBQ��	�'U�uKǧ�6��0�ԧg�
D�'Bl�1m� ��L�䩇���=J
�'�f������!KT@L"���S�'�U�����6�
q!F�A�8�{�'�xP)w�����Q�! ~CxA��'m�x����5���jvg��qd���'��)R�P��p4�+��hy���'�1� ��
6�@\)��b�D��	�'8 � ��1O��C��
r����'���������ǉ	����'ќ1��A %	s+f]@��d�4�?D���q�ʃ��Z�P�}RE���!D���Mʏ~��i���Ƀ pB	�A /D�p�7 P�rx#Et�>�`�-D���B�򾁃�H�b�!�G/D���'�H6Z�T����P���Y�A/D���NL1:C�!�t �!|QB$d"D��R�P�n%Zí�8\�<0S2D����A�"R��n��F",S=D�����D�:]����]~��{�9D��BG-"ax����o#-oz1��A4D��3c�Ĝ��1��v�F{�&1D�1����.�ιCBǐ:5��"S#$D���%c	�	Œ����������G"D��µ�[oH��mK?#��$Q6�.D��I�jB CS���D�H�Bf����-D����2^,x���F#^�T�Y��7D������9��~�(E���y�	�<7��0�ċ��g�z�y4��y2���D�$� ��b^���!�y"țK��Y�μc�5���<�y
� d����T��#���-o�EJ�"O���oEe�h�1�*V�/�t���"Of�R���Q,��
=��Q"OJy�Ù�h��T��i��Q�@�&"O�iہ�W�whVxb�)�5,�٨�"Om����Q�b(��.wp�Ce"O�T�0���L}�}�$;*u�tB�"OF�����_'��z 6$BLl��"Oȍ�$[/E��\�U�V�\�Z��"O*5��M���[T��:.���w"O��#��3U���2��Jm�fA0�"O���A��$�td*�̮'���"�"O��ئ��	��m�C�L@��/D���U#��Mf��2a�)-�8D˄*(D����d �pt�@wA���2�4D�\��B�p�:���f
>"?��S�2D���T�Uc�7+G`��F�d�<	�/,�T�AK��P91Q�V�<Q7�-6=b�fd֭d�m��y�<$e$�|\q�	5�:�Px�<a%�N6F���*� ��Ej �GI�r�<y��2o�t�K�$x$3��Yp�<IgLO��hEstH���$�5��L�<)JP�7�ҏ�4A��(��VR�<	��B�9*0��uo[�,��8T,C�<�����d2�%Y�R(��(�"�]�<qe#���a�����\@r+�Y�<A0���5>! F�ݴ$XAXSd�`�<YҊٜV��l����	`ׂi��AP}�<)�B_�
�>����^��uH3��x�<atMЋb�h	�+n}�}:��Iv�<)g`�6a��9����1��p⑤�p��R�Ơ��		\?n%a'd��(�ވ��/Q�z�"��$_"H��uCL: ����㭋�"R�xS�j�4_�C�I:��)��^�-c��
q�WE�r#=1�##�ܕ�p����O�0r��:rv�%k�U؎m	�'�� `s	��_�6���`�I���q�4D�. R�C�Y�-Z/O?7m;"��x��� �Ou����P,!�D�mI�`5�C�E߰�P�RdCD�$��8�Y��0JU.4C2L4�o���Z�*0�	���:X=��E����� �� �hd���R�txX�s��6:��0��F�9�,4���0,)�q���!�F��3�۴,2�p���P�!�R��2���6�Ps���_n�ݲ �PȬՑ&��=�y"g��4ǐ\W�D�O�Xk�˖-��Iw٥0EN5��a��6>lю��O�$;��-aV���P�5J�3�"O�"��_�-�)��ɐ;�X��g!O 2I�t�6�"���E�8��<�Cz��Q�@K$p�)���*��퉄B�4��F�s��� &�Ńk�(��E�:n!pa��!0X=�r�@���%ߋ3p8d[e�0S/�$Ǧ,��+y�ư+W�϶<����e�BL����!+�䍱*����l�����"O���O�Kd����a֝k��a��<p�ܲ@N���f�K��N<&O�>1��/b ��H�
"28в,O�^�����d8H�Q.�/wrzI��kɍ"�@�+�Xe��p#��$8��*$�������0G �����"%&

G��{Rj��p! �{ ��pǸ�j�" �`�b�j6��|��i�1��������+�^DXgI�#�N�� ˞���f���(���޲
Ǽ������N_<"��P��K�FP��ʶM_�y�E�?o"e��	�:F�~��gb+�$�`�00�+�?E��'���ݑ2@@�C�y��'d�q��Y3��ˇ�	��0sD�>��4S���c���}���HM:I"���
όy1�P#�p?)��]�N� ���!G_|S�*��x���1q��D�09�X�W60HrХ�WQ���$��5�pd���G7��q� �(F,�����y
� ���&�/�hp�`�>�}���O|�R�H��G�1O�>A���En]|����2Z6�1�)D��jp�"*��a��Y�s�@\��)��W�hgr���ɉv�|��"��8X(P�__F!�D�M��`Ս��X�6��v�\��!�Ą�)�͛<��(æ�_�E�!�9,`�5셈h��E�L�g!��߷>G:P���8K��Rso��!�	#0c�| �fW�)�[H��T-<�!�<�M3�-L
{e�@�p���x�!�_��[po;1V���î�898!�D&Qrb��KE�D�M��LH�!!���H�.U+�-�u�F���U!��*<�:ʀ ¾A��5�橂h
!����%��N�y�0Ic�� sV!��Ӻ7V���j�����eUe!�D�2O�T@���;��]�N"V]!�d�	��1�pE0h���R'-Vr�!򤅶PBЭ��-ʥ�F4Cd�Nz�!��T� 5>A�g�W+'z����l�!�E�?.��Q���!�0#I��!�$��O�� �����<q�B�M��p�!򄄰+k,�Xv(ۘ~A��Zg�@�H�!�]�p�D���J%N)��!V�!�d��g��A�w��W��(�.I"q�!�=ᖭ��C	�?d��@NH1 �!��ܹRk�d����Gyxp�B�۞y:!�ғl:.1�!`��A��3��@fS!�$��q��m"T��jD�cGG�)A!�D�I�Yh�NE�^Q�"��Uc�!�J+)7�H(bȄ��Re�BLή}�!�d�1����򊛴w�*�*���<e*!�d�t��pqDG����ܓy%!�d�xr)�Q!�"��1�b!�D��w�BLA�6]zv�����!��ǀ+��xGi��~]`�̅8.&!��/EO�X�D	Ճl��0�f@�.�!��-���"���jH �"��V�!�d�$� ����
eH��T�E��!�R$p���k��F�&�~�T��/*!��R>}��JQG�W 4�vL�=~@!�l�l%G�"���qC@&�!���(t�4�$��d����3��!�$&#H(:�]Y��p���{!��X������KvI���Zm!���STܙ��̶g�9�H	R�!��Z�}�=Q �̌fw����ݏj�!��� l���	�`K����V�^�!<!�$�	,�D,��T+e�P�����"`3!�D�&��))�M���ź�ɨI�!�D�	(�աdjV�3�R$�RB�d�!�l��s��9n��3�����D��'��j�땓 �2��WL�����c�<���!cW��	C��8��S��g�<񥩛'�t�2�fѿ4�h���	�e�<qת��s&�Dr��=^�N�pp�Dh�<��ᔗ1+��!'l�=E���Ѐ�x�<�"^�瞴�!���{����Ɵu�<��2?C�xQ3��M�A�V��M�<I�&N�.��tB�с	���r�-ER�<�V�В^���K2��-�e�+@lܓ6����$ޤR����U�Y�T�%�0Rv@��h2�����pm�8�D1D��$�\��$zT*E�i�� p��+D�\cs&��;���t/��	5z�!G�*D�� +���&R���zT�K9A. "O�-�FcÏ$����c�ۓ[Lڅ&"O6I��ʔ�"�fmx#>x.d��	�'����O�1``�q͋[��	�'�>��O�M�x�S���\�� 	�'�r����V�9�Xs���(j�>Ys�'f��b��N�;����fȌ�M	`,�'0�˱hP�{�}(���0�-��'[�Ƞ�m-���GK��B%r�'�>)�6,i�ّ��	*q�h��'���`�i�<>�z0LW-;���'��<�!�P�8����W �	%�&i�'�ZI�a��@GzaZWA��N���C�'�̕i��TU�
���L؁Jߦ�`
�'3�!HU+l�l�C�$�ܐ[
�'``I� �$F�
%ȀG�<�+
�'1t��`�	�������r��a	�'4���wb�e< jdμ�'*�+�y�W�,���A��޹�mL��y҄�h��p�g��{�Ѕ`�G��y��@�	.�Bp���iqv��Ti��yr��;/a~�P��S�a��4�yc_�2�ɱa�}��$��y��%zHA�J;7"�
DC�7�yҥE \��E�3B��'7nX�h\��y����Ha�E
�V��p���y��'��
�j[�ȶ��$˖�y�)C	�(���L+% ��)&�:�y�*�(.��9"Og�
���y�f���<x�1	�^����.�y�'B�G�zX+��!J�P�����y��<7`*4C�+ۭ?"h8y�/�y"	�7 ��m��@N ��2P���y��@d�� 	�Ni��"�3�y��8`��C�b`�����yb-�8��}��EY(u8����y���������*_�kJ8<˕�,�y�a�;H�XR�Ό�sѰ �T�[��y҈�(���jr
��8�y�N��n[`�9M�^FdC��� �y�l�"T���ɢ�ցg�<�j�#�y�FK�e�b��� ���Aw�E��y�eO�J.��"oA�T���P�D��y"�0����Jl���!��%�ybb��y��@�DJ�\0T��y���(١��Ӏe�h8����=�y�!�������k��,�t�A�:�y���.�V)⑅��716��фJ��y��C�����65jLY#Q�ӭ�y�����5�'f��*��Xs�@���y2h�1N`���+'2�\8�Ӡ�yR��Y�="e�T� @���y��Ӱ<��FٻzY��17����y#����y��O�rcZ��w-\�yBg�%U�����Zn(�;��M)�y"�	2�u�F�� 7L�fV2�y�k��j��s��1�VOF��yr(P$T�jM��GD5j�F���C��y�M�G��Gc9Ȩ g ��y2۩s���Oɱ_.��׫S��y��N� �H�3m@/dh�H�r� �y��)F�>��2j	�]Ɉ��Qj���y�ȗMw�}KB�##�Phqǎ�yR�� qh�SK��b�����y
� ,�ˢ/¼�\�5�ʣs;����"O�2��N�B��xh�c�N�@�"O�ǏQ�U��2�V�v!#6"O����.QF�y+#�&o;�$ �"O��(��ŋ��Hz�"���"O���� �f!eއ^@!�"O؝;�(�k�"e�ĕ����b�"O�=�UC�0*f�ӧL�!L��2"*O8H�Oܖ!��z��II
����'�B�8u@�l��d��J���'�T�N�<,�ѣ�##�n� �'2��A�Q:u�{f(�t�x�x�'px�OG��8V�@+]6���'�j-f`F:)e���F�6̩a�'!=�r\R�Z8XFh#G ȓc&+�����+U��"/��ȓ��h�1�L����DH�����fg^L�d��T���PA�Qi_x��A�.�1gܰ�$	 CƐ� D��Dʎ�Y"FJ���xEF�X��D��7 ��[�FĻF�`�'r"��1�h����P.Q0�W�Ҍ_�jH��zVb8#f��h�c",Գ$R8���G�����O�pT[a�K/	����vՋ���gq:�R��1J������d�u,^�Bl��ڠ�-���ȓm���+;���*7���
��t*h|�;EDe� �W"FJP��'&d���	�.|�Ř��SJ�ȓ�J���@�"crM(�H[?ǤĄ�$P��K1o�}��RD��H��>�b9�T�\/u��k��8W'���ȓ?��@Sc�Å���H��2�ͅ�F�9��j��q��E
Ɣ:�R����pl�Q"�T�>�{Rj[:`:)�ȓ�h�����+R�ܫp���e���ȓC���ڦXv<l�aX)cP���� ��,`��Y:* �-KB+ŝ��Ԅȓ+Z)�BҏO��m	"\!M�(������� �9@�.��pD�G[|���=��l+3KǪR
&���#G�H|����Yѓ��@
z�wܲSN�]��Z�D���6(�T���U&y�F9���|\��=v9��#*P�~�����7�
d{W��������f�+�ZI��og*��Ǐǝ����ڨ>�*ĄȓE��s��V�hܻ�����ȓ&�Bx(��X?�p�Ӏކ!ݖ��ȓF	��3��ɢ�($�Y�ȓu3�@{���)L~ t�&h����.!��J��Rv��qh�9��(��ŴTI�ž:6��&H�	L쮼��kv�DlE>jl�m#�oI�/���$,ړF�HY@����1�X�>@-�ȓ38z�Jp� n�)�r�E�W���ȓh�d-+QC�Lb���N���f��3HEQ�m��M��=r���C�	�8�PZ��V Qa.L�Tl]�m�B�i%%K-�%��D؀#�p=<e 
�'��Xђ�B�}^��1h�s��t�	���$JzL�0I4;* ��0MJ`�<9נ0;�̃��3{\���Y�<�W��,x´��(b7b=kFW�<�Ą�41\t۲�!?k��R�<� �iР�W�l�:�&蔤t�Z�J"O� c���3aZաp)�$V�di�"OB8ۆEI�b����h�/6Т@�t"O��K��ɰ=PRd��'�S�b)�"O�t�BF�k
�����:Ѳ�"OZ5��� C�0X�;�R0�e"O�4�#K�>�47 C�"6�I�"OH��U�U� ��܋c�[�C��@"O�}pϔ^�H����_���ZC"OtxR�	+�y�Ӣԕ���r"O$���f��إ�����6,m�a"O8P�3-4{���z5��"O�h��ѕ;b��M�<�ti c"O��3�愖d+F�!",�,n��"O~��F̃�{室i7d�zs$�9�"OrQ�b'_=<��(B-	4&��� �"O�U;fŊ=>ٚ�q��0�����"O�YsJ�ZԜ
�JF�(�1c"O�12���Hj�'���TJ�"O���P��� ���Q��8�C"O摫�-͍"0HX��e��$�B�"O$U�ä)m5���g�_7H���"O��i�M�<�*1��ĉ�2��9�"O��"��6l�P�"֭n"��#�"O�-���OI{����a�=^a�C"OFM����5t��%�"�O�.Ё�"O,Xw��0�6c��TH��"Ozubw�H�5G��bf� �x���"O,�Q�J��<q����6쩁"O<���H��+	�Tk$Q��{A"O@D��H�3|����Նh�4�"Od8���O���dFQ��a�"O���͝�]�؝y�ť0ƈ�h�"O�-�a�v��j��ٔ:�x��&"Or���O��q��[�V�J�"O�q�&�+��|�3���pY"O��K��ʴx�t�2���!�&�[�"O��aiȀZ�l�f~쒀��"OJ�+W��`/�<�F%�0ξt)u"O �2nH5^�4����!�� �"O�h�DE1T�h���p�bAP$"O�)p�H r|^4s�ՂU�	�5"O����`�Kx|�RH^ &.��#"O��Շ݈Fu<\	Gg��3�4�"OX���)�_�~��ƃz��"O��ks
��`�>D�c�W���� "O�0�@H�p�L����,T���"O��b��J"�x��	FJE��"O���.�:p	��'�2*b�PW"O�,1�'ҡf����UA��4��b"OQ����!)���� �Ҍ�#5"O�d�!גGG��*&�_�\�2�"O2� ��<V ��2&K�7�%�"O��wCS��[Q�T6;�L���"Ot	P&�?B�̹�3%�u�& �p"O̔D�Y�pB�-����i�H�5"O�0��һy��@ B�/"$���&"O�J��ۘ"1<#�!ÏZ��S"O|�Za�W��b%�R"S�A�%"O�� q�^�fj<���H<K��qQ�"O\���F��0X(���ݧ}�Ҝ
"O���)J�'���2o��ɮ��$"O�xAt⏸j~��3C�Q����A7"O�`��+E��uq� r]ΐp"O� 
p��M���(�G���wD�ѐV"O��u,T+>��GW_2�X`�"Ox�P�胷.6�E3����:}�V"O\�	a)�<q��������D"O�����@�fm��W�d�P�"O�U��#յz���R�Z۴4)g"OH�#���	����c��0�'5�1��@0�4�4b�
�i�
�'�hU@�j�Vf��G�?��e�	�'6ꗖ#$6�YWMǳ/���Sb�o�<�!��3����P��R~	�O�l�<ѣ��*���OF8z����_�<���F�5��,��F�b��Y�<��aɏa�f)kfڂ����B�W�<yT��=p�34g	'"��ء^�<�T���1J�4�.ߋf��'�b�<���܀d�J�G�G�mCd�IL^�<!Q��4J��}x���0h��ٺd��<A���$P@�s�Z0E̾��g��{�<���]�n�8q��@J+c�ܼR�F�<adH��f�*�@�`��C���T�^w�<)���],c���4?̔�AYv�<9ei�.0��glųl/��Z��p�<y��ۻ_H�#r�+L<>Y�d#�l�<�QIO��H�ja,��q�
��%��p�<��(_�1k�Y��׏JPH��.�j�<�#l[3M�<��!�@�N2Vl{4�~�<	�gT�!eb�c�-%���@�e�<�AJ�#��b�*(H>:Ĩ�x�<���;9�)��/&m��ِ	I�<�6��Tj���OJ	�~�����J�<Y���1���2��Ĩ��J�<�Ӎ�FIf9�@���sڒD���^�<�P�8b�<Ұkڗ%YLxF�C]�<!�j
)hE�)J���Si��3Q.�r�<I�bK-D��R/A};�m��&�W�<�r��i}�g�
G,{��X�<q�dQ�'jF�Y&��O2����&�_�<aFj� <�����]�$@���Y�<�$�GU���G
��b6��c�S�<a@%��7n�Dq�MF�?�܈��L�<�7��eP� �6!"�b�`Bp�<�
�5P�\k�}�R�� ��m�<�Ed�I	�!��Ö �B��lGk�<�r�N65�Z��sB��K>���DWg�<���:c]8(s�g�
S�6�+�D�d�<An��c�:9JTI�E���#B!T�4:����|P��,K�֬�(D����	��{0)���WQj���%D��ᅋ;yRb��d얧TQ��Ѡ�$D�,�4S�\ҥ
�b�B�n!D��ku�R!��i�N<!�
8�É#D� ���ۅp�Z���6F��=�Bm D���WO(`$����ѵn��Ib��<D� YBIՔ,����qD��g���a�5D�x9Co��~�N ��M�):Ĥ�e�4D�0���]��`2�"�(���2�3D���G��'�<�����X�l0$K0D� �y�X.ƒ[w �a�,D�0����H����K��=n�I2K&D�T�Pmހ{t=JF�@v��� "/%D�\�0�Y�:K��P�l��XS�1�(.D��@i=R�\4�� _�	��y�/D�h�u �Qt�b�ʐV�H��D :D�� $�p4iQ�iL�����Fg&��"O��K�+�\w��z��@��bqpT"O&P�n'Y^D�q�MU3$�X�е"O�I箂"J�����)qvU�'"O�a�B�6�$��#Oި]�d�"O�c�@E�[�h�3L1B}y�"O^�:ǃC18��"G��B?c�!���fKz��I�>qb�H%6q!�DN4n{��4͊�]Iv���j\!�$�#�ʤ�T��Y\f�[��1>!�D��l4�#��Z��C-�8%!�B�O���ץT�r�rH���&!�۶�����1&�AS��^`!�ɯYH=�r��z��j�)�!�d�.*(h�Q��,cD��d���!�����W.A$@AĽℊ�Tm!�$��<^� d�	��UI4J!�d �V%�TdD�1�jp��(�&<!�d��_�\{�b߲Z�޽y���H!��n}�����;u���	���.8!�d[�+��a��� ;�"�x�aŎr#!�dȰ�HtP'��&Xq�Li���pw!��H�<i�I� ��*hlz�ᘛ6c!�2��d��L:�*�O�a!�$��r ����CS�a�th�4	��U!�D�	_8i R�ʡ��e`c��kR!��
�u���F J#��Tѧ"�=f�!��ƅ*e. ld��9��� 0�!��U���Yu`P(Q�nX�K�"�!�D��N"�´�;h���Zu˛)._!�D��W Ԛ1�ӸI
�pid�ƛ=C!�D�;j���1�U�L�X�I�"*!�dA1A�.�
�FK3lѨ	 ���L!��!`x���&6^>��IY�!�E!�za����#G�@�@�J(f�!��ŏ���ʀ�(SZܡ�f͒A!�D��t)j�W��5����J?B7!�DY�w�P��/,�t�U�$�!�G����2+�$o�ȝ����F�!��$�T��!Һb�ƀ����6�!�$�h�D	� �+�|���0}!�D�[��jt� gi`��CiZ�<~!�DTcK|=�Ī��g ���2ӻ|s!��2d�VA)bH�0VLFsV��!��;�� ��$�-Ta�\�b�$)�!�d�f���j�c�cR�9���I�q�!�d�	���ˁj[5CI��y!�v�!򄋳S6.���3|J�q �`Sy�!�䍀0Ad�`�A��xE6	H�o��I�!���6q��� ��]'N6����_�0�!��z��%�e��3|R�m�Q�!��A;ʔA`GE�r��s��v�!�D3$LPQ�W��k�PTy�	�k�!��Ee���i�Z�}��<����!�dɣd��k��\D8E��M�4!�F��6a� gӗob��@�&�<>!�$I�La�XѴ�	<N$ B�Tl#!�$J�;j�����B ���\!�Q+-���ôՙb&�	@!�`!��N@����1�פ%������6�!�Z:;ؔ�Tg:NB�]� �H�z�!��h:}9��)R�&�s!˚8I�!�D�to>�q�+�C
��fcz!�H��f�	e����	�"��{�!�� ^�C�"��"�^��V�_:Bx�@ʕ"O�(�N�F�.��!�N���P�"ODq4��Y�h�J'PC��t�r"OȊ`���6�Y5l�=?e��2�"Ob)�d�%~�H�@ O��4�ˠ"Oި@��?*����o�p�����"O�������-`�B�p�*0C�"O�	[ k���t�vfD�n���u"OzYsD�A�B��u+�^���"Oԣ�#���2`r� �H+�uC�"O�%R�N e��h�〔)�=��"O����V>6��X"�!܃s6|��d"O܉�`�5	,�l+ �B��h� "Oq�h�"p6mKd���<�X�"O����>۲�CE��i����"O|Y�n$�����O�mӞ!"Ol1#mL6���g����B ��"OnRga�{�<��1H��z9�"O&�AF�3Ih���+}��3�"O�Xb
-V�X 1�UH�l`�C"O����-Dz���Ӊ9��S�"OB!H�@�5x<E%C:�ЭC�"O�hC�-H%,]��'���E�"OL� ��ϰ,It��Ǚ/z(��"O����* ?[�lɁ2	C��$	��"O�a�F ����m�a��B�"ON�bԠ˲� ���2�$Y��"O�Uj���P�Ԕ0V�'R�Hd�"O�-���C�]����M���e"O�!H�o@.�RU�gOW�J�~��"O`�\;#�-��L�} ��i"O�p5��T�	Y6ꀾ�j�e"O�W \V�Q���;���v�D�<���5�(�u'��Sh�S���~�<YbZ�����<�0T;���w�<�W�#O E��텚B=T�z`�l�<�Ҏ�� ��+rȃW~��DAN�<�g�P2��5����V�H�O�<q��@Z�U0Tb[�kU�hH��T�<q  HZ��ƫ"b�k���P�<��G�2	FA�ɦWr~t;b'K�<��f��a����B���zX���D�<�SG�:2��H������ҁ��B�<I�(_�c}�eQ�\�VrzA����|�<���W�u�f���E�S�B�iv��t�<ɠ�8b�x;�bw���b�IX�<ɇ�ۘ<�$ԃ׈�2CCH��F�]�<�燑x��J�I�#f�8DWoB]�<A ��:����ݙO}P���MZ�<����pfJ-i�H@#������W�<� #Z�O��5�Djڕ_>="��Q�<IgȀ'�����l
���#CV�<9�W.`jLL���ÎF�R�X֮�Q�<���ɢ)b4��BE��Y448�O�N�<����/V6���D�!���K��s�<aF��~��!֣1����!�U�<!W(H{�t�����%aR�a��BO�<��I+���i�K� 
<Y&iL�<�S�G'8�9SF�R��qY�
�r�<����+�B9��o�`�R�6.r�<ql�<H�8b�fQ�gY F��o�<��D� k��3��68�q�@�<adm�F�ܤ�t���yD0���iy�<���R�j�` b.�Pj��y�<� (y�u���@4:d��b�L㠕�""O��SV ك[��P;�'���$�"O~iC�"I�oÎU�f'>A�Jű�"O&Ș��`��d敏Xk��0�"OP��4
�+C��J�ǟ� c(�������h�,P���'���\?9��MEj y����e��,;V%��x�t�0���?Q�k����KCs�7�� G�@��K��|rb.Q�"n=�"��%؜�3��E�'�P������ G��V7�j`b�s�J(�g���f����/�
d.�a$	3ғH�U�ɋ�M����ľi#��H�̋�>����1�U�����3Bߏ����]B��?IJ_� 0(���Ɗf�L1�NTZ8��C۴%��V�il�k��҂c��Ӑ�S��(��'�v�Q�|�����O�˧��ea��?��4Q�uHW���-��L'/�pe �C�8��B(�mn�C���(knx��������X!4�pS�:	��Թ��0*v7��
X<
�@�[	w�A�! ��tZ����� �s��	���%��Hpo�����H�vӒԣs�'F�7-cyJ~bɟ���ǿksو��۶u/v�Z�ꈷ���tyB�|ʟ�	�R�͸�E��X�։�#� !�V#=	ݴd��'�7�|"]w��yGo��X�Ę%��jE����*�O��dL=�@eiQd�O2�d�O��Ժ;��Ms��W�p� ��2fnyH1�U���aIA�X=��00G�0 f�uXa����&�1�D�hs-Q:��F�0�E)"BY���jv�ڧVWI�C�S\�t
[3$��c��� �?��q*v�1c���9��>Q���ҟ4�	���?����$Ɓ_N�����C���q�C�"A���O���ɝ,���)T��4w`��E��-̘�Qڴ����'p7M�O�	��˧F&���8����Ѥ�5;��,���6Nm������?���?�F��?���?�F*��]D�E9`MU�pv��.m��耠�<2�����Z0&����C9f���`$(��S�bm�rK��G�@J�K�4a�^ŋV�R�Z�P���ʿW�T��u�[��HO摪�'@B�+t�\0{Pd<�3`��;`�YEE�B'�7-�Oʓ�?���U?	P���y�B�]rT��!D�8��2
虈�!#ߨ�h����ʀ�D8�Mk.O^�ڑdQĺ���?q��l�� �;^]af�G(ب,H�F�;#`��֟ ��}I��0 
�6���e	) �@�1�4��ظ�cپpK*��pD~ꁳ��?$�����%�>1���9���S$�.&sV�У��5i�QB��Y>8�pZ��䐂9��bӚ�n����O��2!ˡ0و%F�CK���Ԭ�O���?���OD�cD�;��"�����|;g�'��7����o0Dv�)�/\�1q��a`�\i��!f�pD�[� �d�O��' x��	���?AߴJPxˤ���7`�a2��O:A]���ĝ�{��8�`=(p��×�p)������럀��>o ��������eM���6�G�-ߒ�P���?h` &�W�e�_�k�`b?�o���
$�ȥb��@bLh��6M��[�,l�5���'���iUZ �)жx-:U���>c�y��{�)�IT�O���	U�nZ��a�'˨s�Q�p�ߴ%����	aݕ�m|�H��e��y��!�\	���=��/   ����O������d~f�0	�'�>H�e�!��X0��&��TA�'4�\�ī�	"N@y�"�
����'��L��)Wvr��ɓ�p�� ��'F�ۄc0T�h�!`��g;��y	�'%B��6� � �ج<Rh��'|&Y��H݌C] �Ȳ��3c>�'��p*W�XOQ@�8��Q�0đ��'�����i�@���c�8�B��'l���b-�:AV8�Po�8�����'�t�tϱ[Ed�(�X� ��t��'��Hr'���y�Xچ�0p#��J��� 8��`a�Ѥ���ʝz�-Z�"O�h�ŝ*�rhe(ɕ5>�Ic"Ob}; ���O�f]p��[�:�8���"O�)����R`�r���F��q�&"O�X�L,∔�pk]&��P�"Ox��kŦ>���� �(&�fQ"O` ���Gp�.�+@��%�Ȭ*�"O�+%)�2J@��VA�N���"O�2qI��B�5(Rw9�,0�"O�"���<Q^�kw�2$���"O��"v��=?�AF�"V��"OnI���]�{TP4K����"�9��"O�K`�=(䖡kW�ْZh�t"OP�t��#-Hp)�|�qyC"O�,"We�:J��QV'��j�҂"O.���`�`Nh�/њ#�<�d"O��+r�O;�6���+B ��"O���4�݂{+2��s�ڐVg
|�"O>H�82<�t#�;�l�"O������9k�e�w��^Mm9�"O \h�C��Gl����ӿUp5�s"O��ԧ�� :.i����.'�"Q��"O|L 5�H:�E�ƍڧ�bh;6"O�m�p%��8^츙�+T�{^�C�"O�-��I�\.��τ .jY*P"O�0Pg�7r����n{�#R"O���7�� �:���c,�7"O�\P�G�i����p�ŮYa
y�`"O
�( ��
XN�*�Hܤ#�" a�"O���v��\L���,?����d"O4��5 �u���f���1�z���"OvU�Q		|m��E��+g"O����)H����DM ���!"O�� VJG�oڬ0!A�[�jpD��"O�`�p�@�]�Y-ye��cC��y��a�ڈ�4�҄hOz��&�yr�8e����-]����{����y�L$7K��B�^�l0Q��� ��y�E5v���PS#����s��yB"�qI���GU�{�1j�D
��yrX�g��$[1��+��x'�y�.��V6mY���Bi˝bid-��'��Y�T�:�y��l�����;�'��=H#FX�e�b�s�O<
�~<��'��[�L�yL��Rƾ7���'�x�H�߲j�b8�F�g���#�'(��wdYVz]ఌ �Q
B���'�fm��c�(_��Y��C�,I��'?�\�G�ԛd��  W愼x��;�'0��Q�]�iX����(k�e@
�'Zn��P"��!_$Ջ��K(h�a��'@ʅ)C���N�3��IXR����'<����C�,L$D�+N�J&�i�
�'����,�(�@�����E˔���'~����΁9o��I��D��X	�'u��BB��~_")	�BP	K`b���'$^ RuB�(\���i��C�F��	�'����g�+"ߊ��q�T��m�	�'��(b֢ˉ/=�82)�+F�f�'�j� @ͼ:)���w�H�'Q|-���[[jdH���E��|��'ӄ���&�����B��|�����'|����G�:���/X�u��'���x��π�U�F�`H������ �Qs��v2��b!ʎ�͌m�e"ON����lЦU
!�W<O(�P9"OD��Ǒ� 6Ԩ���'P,Q�'Br$�AZ�	+��<�!�'�\Ш�JɵMؖH�#���E|H���'~�`��t 4\j�M}kz�(�'��X�q'�.��x�ąP0KgP̉�'6́4�VUxL�gc��J4�Q�
�'��Ə�C�����AH9L]��
�'�<�e�T%D�jXZS�D3A�|y��'�FE��� E���qR�)��
	�'�0�r�� -��&�A,ʼ�	�'��+�kF�Eh��S��<"�'�Q��
�Bfv���Cu���K>���0=I���ߘ�d�	,�^�J�h
p��$�$*�b��d�ߠ=f�ys�ŉg�4 �,�JH<����D�:���V1'|�rg��L�'��/��N9*p�Q�	M7l�襓�CQ4�x�-nP!�dO�p���sg�$%��Se��;q����<��-���?7*l�S��M{����,ł��!��7Z�EZ��V�<q�j����9FɷN���c]3g*�'
�#Ԑ}�@��(q��4�g�'e:��
��'W(���F�H�ʥ���jDS&�r�N�KR"I�t_z�0�!��m�riL�d���J��'��F�H�Q (�y�[�$pʌ���xa��j�
� E�ޣ]
�OH(MQ�G�e��}:@ I�L-Q�'��Y0���D|�3F��\+�X�E#j�+�Hԧ����)ؕ�h���()�Q��0x��	�鉶�!�dȓu������J% ��4x�\n��=[�.<	o�U T�Y�w/ȴ�"�Oh��:�눨��Mh���&�9�tD0lO�P��h�g�	8q��1)K��@��:^�^����>'�,��L)t^����I�Y�)��"��`��t:6+^c �b�̈S�(j�
e[���,
�L`��h��+�0���g߉8�Q #�$+-�B��<2������
�f����ùH��!G��,���h�fϽqp8�9�t�OȖ�	������Q�K=�"u� C�C�I�fPd���F^`�X#a�\-�Diڴl�v�`��,_�$�ᖣ�v�ɒ5��Y��Ў1�$�c��E�|��d��$��õ ��e�*xI��݀TH��`�e<p���
L�$��J�,H���bG	�	Jb�Ac�ț
�ܠ��"�ɣ[PP:�"�24���
���w��O�.�d�2j�	r+�=0�
�'����@�E"iX%F6�+�OH,E@�
qb�����Ha��~RƲ��]�ㄗT�bT��Lح�yBD�u_
��Ӌ�&e�9(�0���J8�c�T�8�����'�Ę�3$�����- $H�q�R��9� ��%�܌���S�[U�Sh:�xZ6��8QaB/*�����;&h1;�&PȈO��C�h��v���p#�	�¼\��N�owɫ�\�?�!�N�WOt�Qs��;r�4wG�a�L;u�$/Y1w�)�'��9�)Z�- �4��-˒B�k�'(�q�0�n�`q���!�����O�(��*���v���9��1��ڎH�����)j���D�u�rq1��\$�TD ���p�@�Z�<ѵ*����:"���B�� �h�ȓ�Dd�Ti�n�t��B�Yz�<Ō jTJ`�cbY�}�����m�<1�A�#�����D�j��lħg�<�R��1c��ci
S5x�Ť�N�<A�M�
�4x1gʖ�
!�|X7.�f�<1���9:� ��˖V1"�z�J�{�<A(�<��(��chͺ��y�<��!%��K���!]պ�r��n�<1��5h��IB�M%I[��1 �	i�<)��D�F�h�ᦄ;f��p����c�<!G���(�yySd��%@YI!��}�<� b-EN�[uGF*
�(�҅�Jr�<� �L�
xE���AL\��"O�L��AS);��I��^�'& !8f"OdUELS�0�ġE�ܻ4
� U"O�	�g�`�!��iU2��XK�"O�� /�:�(FR�;w��g"O
�r%by-&�GB*.]�y��"O���'h��m]��jW�X�CBj���"O��f�5�r�`q$H�^���K�"O*q ��6����%�i�gjO�<ѐ \I�m3&�J*�<RפN�<	�d�x�"$��ĝ_����Ī�L�<�di�5A�p��g��G�PA��V~�<�#���4��%	�p3}��l�w�<!�YZ�"�	b!@?7�� �$�u�<G��TF~�x0,�LW�ň�{�<A�ܭ>�H�9@��jF���,O�<�F+� [���z��I2�T�H�#t�<1��N�*�:�@0E]*���A�p�<	AP@����J
�!A�Sg�<	�A	�1�R�q���/�H�E �d�<i ��\��0�� $��B�	u�<�%bɬ��<	S��|d�ѡ\O�<�7�4\]��cF�%�99g��A�<	��� 0Y��.�ypP`k�.�\�<A�ܫx���u�EJ�������q�<��#Z�!����2i�9>"��j��J�<A�'
#�`]PU�2H����,�`�<Q"o��9v!�f��:�,���^|�<�Ī��v��GaH.x�8yH�%Zv�<�aJ�);~�Ę���L���D�}�<ypn�(ق#���yt��fFZe�<Qu"P 4KQ��J�2���堖Z�<Iϋ�V��}QQ��.Um&��!�X�<����襑�Ń*% �t)�W�<�&"ܸ/�})'L��e��Z�*�x�<I�̊!"��H�ښd�~��Ҋ�z�<���(r�D���LzƖ�1�Oz�<�4��0�Pp�*e�p���]�<!֌��j>��nϠp&ؤ G�X�<ᒊΒv��4{��=5�����ȋn�<iI֧T5f��gL7o9N��W��t�<���B# M�	Ƭԫ\��Q��'
h�<0���t��iv��o�@�1�k�`ܓ`�n�7b�y,��5�G�{Ͱ}&��Î��l����T�8�7D��;��V�.�N}⃡ȜsV �#)D�a�L� b��zB��"�z+'D�|q�$�!"N�� �?�����?D��X�AC�b�&�r���%���0�?D�ȩ5�ĴdI��y���h�z�J�(;D��Y��w��I�A^�76�]h�<��O�k �2T��*|۲z�<��b�"Ҏ��'!��zk �Zr)w�<Y��R�  M��g�_�d�0�g�<'��XnFP�� M2i����Y�<��G���H2�F��P��U�J{�<! �ȋT�����G����ٕ�z�<��J4"+��!�iD#>},��5ĕx�<y5̗�a�|)��i�)iQ�`QR�q�<��/�,��f�d�h�$MWG�<a��J;a*d`dZ69t�Q�iC�<��/�G3��N[/`R���g]h�<�d�_52>��gc�|�  Z�<�����vf��"Q
ڑ{gp@I�N�a�<�2��3�x�-��Ȱ�G�V�<� � :0�S�r_�E��x���"O���	M=	l��`'���s	���d"OnB���.f  Em��,�
,�"O(XSMC7%5 �`!��$� (�A"O���E���^0�hwD;/����"O~�(�[<!&��$L[.)s��a"O�#F�B�AQ�<҇d�fϊ�w"O<�q�$@�C��-����[4��$"O�]�&��7�@L���;.��"O4�G�°k*)�K�q�ձ4"O��:Ǯ �2lq-�A%���f"OB-zq��<�$��)L2f`��"O�M�VH��e�3��4�G�.g!�DF�^W�E�DD�3!1�P�7�@�J�!�Dե	��3����x#'�9D�!�I	)D�D#�'P�O��˴*E�!�ܲ\f��3j��.j�T1u�B�.E!�$�&EBI���Wq���.R2�!�[�c	�\�蛦N�J#�4)�!�Y�e�J𫲨
!i4��爌\�!�d�T����A�|�kp��N�!�D˳"<hXgE�����Ғ58!�$حg�T�phG�>H����!��Q>���Hgg�{��h��ۉx !���`� ۨ+��\��kG��!�D�r�h��!�j��i��48^!�D:��!T�Ú�`�3 N!�d�W7���w�j�Yk�!�(�!�$�Y��� ��{J*I�V�5#u!��zI�LâoH��]�4��%"�!���z�� ��-�%��"�!�$ZJ*�*�Uu��]R�#P��!�$^���Q5+�f����7B!�$ً<�b);��]L[r0�''�,-!�dߝ?�p:��6ܤ-#Fa%!�d�s�¡g������3�f��j!�d�����]�9��$���!�D]\���3q���)x.�'d܀#_!�dP41���jE<(Eta0�u{!򄋱�E�� 97��p��6Lk!�P5@4j$x!�:F>���U�}}!�DMb���@�;G6�ݹC�ңU�!���SP(lA4�^";�,�5/�!��K��M�4�k��a�H���!��>V��cӫ:YB M��Iæn�!�$+�Չ��W9)Ԫ9���Kw�!�$R�:��DjE��p`4u)�g�o!�䚹,b�A�
+Ly(� �g�\!��D'���Ke�V3f�D�qdˉO!�Č�r�����j�[y3�����!���NP��El�&NV�2� ��r9!�$�(*ʬ�2�־B��J��V-l,!�d�
P�BU��c�\KJ�S���>ft!�$�9f؋��?f,����� �`r!�AA��1X%�]�^2}w�R�s`!�Ԣz2����F�d!�E,ٳ R!�$��%���A'�Z�\���Z0�ʁ�!���(�2��-p�쫲��+iz!�L:%K�uI�F�z	�M"0(T��!�D�T�&�+�BG�w�j�+��#[�!�] X�6�HEǙp�A�A�O�!�$�&(0u�F�.=������&=�!�;N~6@��aV�X,��oQ�o�!�d�u���	��&_I���� ڡ"�!�� �x(P͐%beyC�N,F��U"O���1a��S�@a˦!4x-S"O�T��\��8"��q1��"O�Xȥˆ�hШ|B ��1x�$)�"Om@�E���!`L��0��Q"O@��NC�dP���)�X`�A"Oh�B��a�F���G����B;D��
�eC* ��B�Fr�H�`�p�<�c�
?K�D� s@U�B�Nextl�j�<�R�Q;D���B.Z���E�j�<��H�pFQ��F��\<��DI@�<�s×�TJy`�"Ƙ6ǆYa�i�x�<i��!p^-�0�K{-��Z�-�H�<���	2����Q�W���A�<a�]� V�ĉ��ҎI�d�)��~�<�Î�?�����E�m���a�|�<i@�s~ ��Nԉ`��mb��`�<W.�B8d�q�:f9	
�v�<�Ĉ�f�R�	��V�(�S(k�<a̔*���8���9H	�,�Lm�<�WO�@߀���B�X6�D��G�T�<1�)@�n����G��I+�<���
E�<�F�8L�B�@�G2w`�⋟}�<A���:�z�ׁD��4��,
z�<I�b�ر��&Օ*t�ɀ%��t�<1�U�sɆ�HB��h�}�U�q�<)��(&��$�Րs�xH��l�<�1*8E�����Q
ؐXsOQd�<���*%��ҝY�n�3��[�<���$�B9�Lʨ]ȱAW�<��bD�@(��[W���b�g�<�R�'F�Z�#�`�bQk��h�<�f�ͮ{y ��r���aAN��6�He(<��4:����& �Z�pI��D�-<��ȓO�m+c��;��@v/� G��d��=Y��C!N�Wp�\0#�B( �ȓ&��4ۃ+��6�D50� 2�zh�ȓ@�F�f��L��a��R�L��W��uˣo�B���RlE 6���ȓ~�ܘ�%
��#����̣��$�ʓyz(�G#��A׺8���-["�B�	?	3b}p���MNڸ��		�H��B�I�-�F�)���.\7 �x�+H�kS�C�I)#!���\�@ �i�Z�V�C�ɠX��˷��P��%�0O�8�C��*k5�!�(L�I-�y�2�Ռ/pC�	
i�t�ԎǊ|���� ��=>�B�	���m�ײ��`��(�I��	�'�p�S�ӹ,�j%��&C�<�+�'��l���m�����:lk$<�'���Hb�%>HM �$�{����'R��{�eF��^�B���E�Z�S�'�|��rM���6�`C�?m�\h�'�z�h���*I�$��'']��td��'r�c��V)�%crDCr:f�H
�'ێ�B,�"��"b Sl���	�'�8s �s�,BJI�jo�{	�'���Do��,E�l��C�<ѥ��"y`�I&7� ���}�<��b�!��U��cH�L���L�a�<Q�n��qPc��Un����[F�<��䟽0�҄9`�ŗKI����X�<��d��z\�gΑ��4�0h�]�<�w�W$��PlZ�'t܈I�g�W�<� ڰ���&:����<@��k�"O�'�aD�I;�%�	��Y�"O�K��Y�N.h�����2X�"O���1�_' ���$�ל���"O�)��kT41q�ÐwB4�p"O�4��OP WX}�bi+b�2�"O�8�W#?"���/@<A$݀�"OV�q��Put�� 3o���f"O`�S�G�U"LБ�-x�u$"OЭ�B�Ħ ﶑�VG�r��h�"O���fkef�čQ���r"O8(���)��aQ�M
&_��I�G"O`-�p'�8Br�Uj�
�lW8=��"Ou����[�1�tO�-
�h0"O�{@KA��ҍ@ 00"O� �Ì��s�쑕���z�b�"O�eiTM�	�>L�l�#'��$"O�� ��Z���C��'�"�"O>L9�eâ1y���gۙ�\��"O�ݑj��M��J7&X(A�v���"O��0؄Eդ!�b�$��ѥ"OX��r�� c�x���'ǽ�&�� "O�X�����H�d�AQ��<Lm�]��"O�СP��%X��!�R"$W�a�"O��*�чc��p8A%hL\�7"O	0� A�bmR���Ĕ/k.�|�'"O^��@ _�E�������9�4Y�"O� @�]f���iFb]����"O��*7/��D,��7��7��)�"OAZ�E1;eTH!#i�`�^]��"O	� h�I/�H��HM�@�L�yq"ObУ���xV�i����:�r0)q"Obl�U)�X|D�$�D%���Pc"O�u#��%9�Mɓ�O�/]$h��"O��r�����@�g�?�\�T"O�g�I�;���[eMU�D��LKa"O8�Ƀ扚�<�2��4:m�X"O�)�g {j��Pr&�\���ذ"O��I���օx&�7?�(�8p"Ol�: �	%�&����)ce��P"O���U�ة2��{aBxd"Ob�!��0�4B�-�qc���"O �R� R�g�
�����~OҜ�s"O<��� +��I��[�$h�!��"OL\��A[�e��L;���&1º	��"O�-��
�	x���#�	�,�"O�(
p��(i�8�!X&=� x2�"O��@B�*&\��ʵ�r��2�"Of=�3D۹/T�p��m��mA�"OvI�^�i�@+,X�\���"O���p�Ih��P���;9��L��"OJ�8��1}:ՙ�`����m�"O��!����l�q!����@}�e"O�RHI9�@�&��ꩀ"O��GX�S0𴃑�O�eN��!&"O�a3o�vy6���ЈR<�8�"O��	t�V26l��a3,������"O�U2���R����SM�-uz�:r"O�[͎"H��h�sF"k��a"O�6i�~������a����"O}iQ�a:p��GA�Aef@�"O>��r��^pp��%Y�	K�U[&"Oy�~<��E  ¥:B"O�Չ���6���r��q���g"O� ����_'� eP�HT, �ݐ�"OA`J�H�( ��בy�z��s"O�ᨓoUuq��@	L����f"O��PR�[�X�`�H"i�,���"O�m�sG�z�Ű�@�"�0�˅"O �`GL�$8��CZ=6����"O¥�7��L���	�(R�r�؅"O�Q�6#��g;�$I ���T5���"O�� �K$9`@P;{=d�"f"O�|! E:
.($�手&}���"O.]H�퍍.�"�CQ�.���U"Oqs۵q^��@ [�~�qp"OV<�fM9"W��׮ے��Q��"Oh����&��C$�2/&��%"O*X"6KÃQ>�ِ$�(r���"O.}:@C_�={P�$Şm��@�"Ot���!�#��@qcCA/\݄�3�"O����];.ٹ�,
�6�
�۲"O�p���B�.B�5�ܼr���"O�yr$��	���΀k�j!*�"O�ԂvFK0�����l��<q@"O#gI��-��̐P� �rղ�"O�t��l�+Qʚ<q�͐�~��K0"O�1���	a���hV/��:m@���"O�i:D��$�V�(�oY`�j�Rs"O�¦L�~6PC�'4�|<��"O��:6�ڊцX4��&13��P�"O���A�I� ����|��c�"ODE��	�/A��[ 牟+�����"O,�9(�Fm:���J��8S�"O����}�`�^0~&1YS"Op�p�\�����t$W�͓�"O�,KA ҭO���b$�Ѓu�G"O�`2���t)��˹1
r��b"O�̘���N�8�{ �_�<����3"O�P�@�H�,(0
�/2�v���"O����L�1���bp��#m` ib"O�D+ ��2sF\��!�٤@S:�hd"O��k���R��9Z�GЉu��q�"O,�hWQ7c*٩a�K��!�"O��36N9!�����׽]��[�"OR@	օA4�PsƇ�
yڸ)j"O�I2�ˎ!j �87揎\�Ή��"O��#ϕ
�@k�D��&��Y`"O<�x��U�lء�#�m����"O,�#3��O `���/}����"O���kT1p031!W 0n�U��"O�x�Ae��B��W�Y3]�d�$"O��sE��7ozU��咮O邴:�"OE�4kN'rݾ	(δg�lx�"Oՠ���7�R��S��S�4}��"O��r� ')X؈v'%�Pl�&"O�A8dl��Cwh]�0�ȶU�^a"ON�k���[��͈�yVɑg"O��!�ώ*�00�ڮW<���"O���@
�i�X�{�*ҧX~Ic"O��[��l�au�U�	]攁#"O���e���U~m2�IC�wE��b"O�˖�F�
f��"2�̢V"O���wc��-y��Dl��E "O����g�d`�%]�,��PJ%"ON9R�`��C�.�q�<N���R"Ot3ӌ�N�8B���!f���"Oҝ8 I6+�Ę$�H	Y�bg"O� D�v)�.LhA���L�TR~��"O�:�KT�U�|���(1:Ѕ�F"OЄ��Ο	�ҽ�uH՞�"O����*Fj%h-�ӤW_�D��"Oʗ*V�%��␰&��+� C��y�X0J)��(�-�(͘����y�j��6��Rl�4%�t�ՍY=�y�\�tU5.w����P	�yb����6�*C�ٻS��)���"�yb$��R���L�(H@�r�^,�y���}��pTl5������[;�y�$�/���1";2HL��bi���y"�Ԟ`���Ɠ6+r�IJ5�y���DX�쐖��5EHH<J�$��y��=���sJ%h��Rm���y¯�0Vk6�@��p<�)	2���y�	�*#h4#d�ݳfnP�2F���yB�M�!���7�Pt��c��	��y�''^$�8ql��n� �ꗨ\�yb��^>1E*�l$�[����yBK_#\P�!�_�Np�N#�yҤݳ%,����B�ЀY��dY��yb� �C��p�0*ڐJ��Q0g���y�͓�L=
=��L�^q	���;�y��		������F�wJ����!�y�^�'u��� ��!E�ԍ��C�4�y�
�(b<��Q��7�4U�[��y��K�J�,�����4cֵON��y�)��}*tcF1����G�y����4rܽ�����\{t�9�y��_$�BГb݄f��q	$薘�y#
�ꀌ�Q��Z��[���;��<��7�N����-}���;�(�>kY!�$G_����kP�'��݉4B_6C��C6���?/��0��c��,�7ツ|��B䉊qj�l+aH��qQ���F�O�,��b����ha:v
�m�
 v%ܱD��]�ēZ�$�3��	�1�e��3=��Yp@"O�� ���"'���X�� +��'�j�<!pkI)m���p�^�HKZ8R��U�<q!�ݰuO8���.q��� �{�<Q�b�����8 	�.�����Vv�<�� m�L�3��/���r�/h�<���41���� ���(R*xJ�" P�<Y��ٔM{�	�`"S�<�(z�
s�<�w�[4Sq�t@�� (u�	Vd�p�<IsDS�&4<��MM#	p��˳ �k�<�!B��R�ťX��bo�B�<)�;-����a�n,XI��(�{�<a�ͯz#���c�6�J�`� ]u�<1wC7[��}�� \$JS�dꖎ�U�<�U� �Pj�y���F��R�<��	�2 W�X��A�8�Pt+���D�<���K�s���2AF��Eߌ|c#@��<)�>4dիG�S�$AȽ:��}�<QT-װwV�����Q�1LH
�%z�<���O�fz�U���<c�!B1�@�<��m .NU�1)w���;�J��2,WC�<9FoV�r���'I�r��`#wd�{�<1UmؗF�����N
�x�`[p`x�<I���"E�QX����n���jr�<���ߟ|ƪ��L�6|�9H�Rp�<���@$bRp�D/�Z諧o�n�<yƍ�d6�Mq�!Ɩe�Lu3fdY`�<� ��2�.�7n���`�ˍWm6�[F"O���4�L�S�Kc��d���V"O*�U��&(�q#�
H�h��"Od g�'��ak��h�ļ�&"O`;�.��\/��C���]�pI�"O4�P��$j7��QAϡ	��t�u"OTY8ň��+��*t�E37wx�0F"Ob���
�N�����χ6nԱ �"O���f@~�1�J�sT�Y$"O�	q�f�:�|3���%�H)�"O�\�V�ۓg�|��$�@�? ���Q"O6�G�
2hۇ�I�Q�E�w"O����Ȍ''t�q���8݊���"Ot���OI,F\L���nE=��UJ�"O��:D�R�bZ�%@d :Q���{"O l��E�r 6%�!n["Y�`T�!"OFy��*L
j�bi�@^�$
X̺B"OxtRP�A+�,i�����.����"O�E�bу�z�d`Z�"��q�q"O���Z�d�H�.�$��q B*O �+��7-`��U�R]�D@�'�
]{�dI�"&~vE
[���:�'��A�$ �>�QA�D�Q8N�S�'�T��Lӟjt���;Ҍ}��'n��c�O�>�8���W�4�>
�'�V��c�
&��,�aS�2�%i�'�B�ۢeR{��sQjʖ"����'2F��P6\+g�6
$j��e"D� *�B #�x��!�N�P.L(�B.D�k�)".�8Q��9�&X��� D��y��4��(�&�y��أ.�g�<��N���R��fKРs$b�<���T5 XDz��tE#kXd�<� L
\y��aD�WR���!l�u�<����=`�i�ȁ�k����$͋y�<��$_�+����ɇB0d���#�j�<�S�F8T�d���I���h�T��N�<YG!��u��@	�-����G�<�Q*+l�b� q�8�a���@�<��l#r�L��VR�,ʒ�
�<�!k�j�D���[�4rm�}�<��I����i���v��X�W@b�<!���eTL�J��Ā6�`L�ł�_�<��>��{-�8e����R'X^�<acH�W8��B�U2:�5�BG(T�@���c�
�p��דO4�DSP�0D��cC@52�B�al�(٠P�3D�����|���B��h�EM%D��;q$'16Ȓ0hEib�l(�!D��Qj��#bސ{1����1E�$D�V�;V����gJx�`Q�c!�<�O ��["VHq��4��O� ����\:~�@���E�4T�m*�{2�'��5�%���:!�WL�'E�$ ���|�'�V::�T�S�D2M�,�� �f�'�Q2ViՆQBQ�U���"�� sӟ\���j�.#�T�7lW&q=$F�ɰB�����צ-��4�?q��������m��KP�\<�0���d�'��)��hqĭG�c��_��`� ��o�a}2�i
�7�pӮ�c���>��rnP�7�R����O��92�\�j���$�<�'t]�Ɲx��И�Q��� K+�Ձ��f����fh���؇BJ�qiŋ���O���;j��O;E��ea(\��J�o�*M�&i�N�XDL"�Z�B��$������C�{���iqmț)xR#�ii ]C���?D�i�R�?5$?7팖86:�"�m��!�M�{���O����~�ր�"8*m���z[Q�0�4p6�f�|�O��"G�Rx���\=28���^08�'���v�<��DQ2N���bJ*ES���"`]�b2���'�C6x�{w�w�{uD�?���)� .8uAC�Jǈ��rg��T��8C₪AT� eʆ ����	F��p�'�D�ɖ�Z0C@~��� �I��Щ�)�O�;$�O��$����Y���I��Dl�!R�,غ�i2����Λj�NJ�'���!��>]�Q�ÎU�9fz������1��4���������}��!�A���I9��L��"�@QiSf¥t��d�OBY`��>0T�ɲ����cpm���2!�� 3�T�R��E�[�m���b���΃W��0�Յ��hib�Ivd˪z�:�1��� ��䣕�VGj(MNC�'f� ���J�6�
�F�2.z`���A�g���%�[�XT�f�'!�	�4�'4�� ��F	g�ڠQf�
�J��1�"O1�J׼9�����d�Iq��Od1n���M�.OV�K7l���IU�7pQX��D��$m�ɲ��U�;�������d�~e�1�<
F��jS�؄{�x(9�Ȝz@H�)�}S�L� �>�(V鉡C��YG/�Z9IW��Xv���O����!K�H}���[^,؉�D��O���r��mZ���Oh�Y0AS�T��PעF����f�O|�b>��IZ}��ͨP�LHi�U�(��h��@F7�p>�2�i�7�m�T	7�T�8��:��X�K��M˒FG�z����'@b�'��D�%L�"�'ԛ��v�*�c�5*�H����~��e�'b~!��W��yB�'���[�,Oy�'�%oj�mp&�I1`�>�ң�iY$��냡�<�8NW�G	��1�&K�0X��k1��:�J�-�,��q,W3%�~�*e�iH�ݑ��?��i���sӾyppAQ��#�-`G�t��$�O��(�	f�5��9s�G&Z�$\�@�)0�yFybOz��o�ɟش�?1�'�u����ݎty2I�-^�(*W1EY�Of��$�?j 8  �   f   Ĵ���	��Z�Zv���/ʜ�cd�<������qe�H�4͒6R64<�b����%�0��-�VEC�A3�0�qC�MӐ�iU��q�ؔ'��	㦱�1��9�bY�Qc.��5�L�}�F���K�L�
Tg0�o��'d��q��˕L"�F&K&�ʘC� 9 ��d�6�����U�B'�����	R}vp��3���=V|U����b�T�Q̖�x��dW(��M�#�d��TĢ�OV��'�N��4"�6Ʉ�v$Z9�:]9��َ=����"�+;�`���]?��	;\̞l�7C�?eNѹK�mMV�y�T��g���?!Q�(�赁GJ�O���	�@���Dj��}�Tʓ= �Įj�i���65��)�B�$M*m�F?�I	j��)S�I�r�H��j�H���9P�T�O��������dQ����˰H~��[7,6'��#<��-�	K_y�fm�@�� #��Z#J6ԡ�OҀ��X�/x�pp�_4�zh#&�#�����$W��Op�2�Op���X3T�����d������_��ȣ�ɕ��O���d�;M�n��w*ۍ5�:�!Α�O:8*���[��?i�g<1����Y������[̓m�d#<��-"�$�,F6�E	[>G���	��hi��U(�OJ��J<Y��O^PJ����}���QN	�H� H��'7V�'���Z�I]?��O����t"RX�$yӶ��?0a��s�{"��g�'$$�O��5����4oK�2�N��]� � ��d���9�.�,������8��a���5D�� H   ��ł%}r���&"O~jai�3�HI��٤uU�i�1"O>!Ȓ ]#0s�h���2Sp �g"O�|@�� \lH1�t$�e��F"O�P��(׮cYZ���,��_��"O>�Ke���@�٥�	2eH8��T"O���A�xz��q��D�G���"O��3��Q/6��!sƭ��=���v"O���ťl`�t����A��Y�@"O�p�Hϋ%"���vH��"O�$o�ٶ��¤K�}� ��"O إ!G��Eq�C� ��h�"O��*p틎+�ԱH׃	�F�,�b"O�ER�n�R�S�?Zӄa�"O�s���>殡#Ǉ���Mjr"Oԥ�$��)jƃU==x�"O�Ő�E5j�R͓�䗜/�ȸd"O�hA�bv��UP   #
  �  @  �  b&  �.  �4  ;  wA  �G  �M  VT  �Z  �`  "g  cm  �s  �y  ـ   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dlӆ�>O��JB�'� �a�0�R���%S�A��$j�醊~�Lhj�E��]��$K�W����aݩrGH	�?M2��?�Rc��Q��M��j�0KƮq�d�5@�ԉ��7@�D�՞U�R��7�	��uGiГa����'�������o��+⭒�Z-8�5�̦C�"Qi���O��Q"m�&�2��S�Mզ庠+Dȟ�����������P��	+/��jC�X
����
���'��O���Ҧ�����OL��Mn�4���(5�pȡ��)DL��%���O�1��@|���'�D���Ђ��M.I���S��7<_n��	-ғȈO�6M�&���r�G�v�X�7I�_��m�'6���H�5�w�0* ��\<�UN�tb�[���ϟP��ٟ�I��0�����	\��3���"�Y2_.@qb���H����'M�7���Yشx����'��$'H6휓:8��d�'�$H��`D�a�(�>�`B䉁Q�>}r�T�dP���`�����c���Ϛ�0��#*���o�,�M�r�i����Ofܭ�'ID瞅�B@L5�l�F��5  ��:��y�X9�&��*�HB +.g���b��O�⟠jr��?=��T`N��$�`@
ڟ���D��xX�j�v��$�g�@��p"7�*���?�����O����wO��L����A�1��!�,O�=E����2&�pX��M�m(���SE�7A�r���������M�ʟ��+X�Oɼ����¦�L}�0�'��şx���|��E])E$�9�O��$��}u@ x'���%� �r͗�m���d�#iU����XR�\�b���OdH�6Nߡ?":����5��]R��'�
����?9�_�4�� ̬W�2��0L�z�y ��O��D�O��b>1̓ �e3䧁5���8�^�`��ć���M�� �5$|t�
2��):\��C���t����=/(�⟠�Ӓ44�!��"�6Tȹ��@��d�d}�ȓo��<TaV�(��e�[=^o4%�ȓ�C3�dc,�R`�պ+E�u��0Z���u�ʅ=@�@���}��@�ȓY�^�&A�.�@ b䡄n���ȓS����VT#�L0�C��E�	1>�"<E�tj�o��4a$�:�1�	R�8�!�$�ʲ���w$��+'�)-���ȓ*qh�3��͎��UZU��$KђI�ȓ`V�MA���@2�e�s*D(�������	XbN��>��PS&��썅Ɠg&�CS�¯Y�(QA���u�� ��R6��$�O���<�-��瓯|��Y�D�N�^�B�╣�A1�1���ɬp�.4��	=G���KC��J�eBA*�r|�Х��.]�x��C�='�֙b�G��m�hxG{�mE5?<���z�V1ܴxun\��d�Ӧ푉�$�<��O����*9���eV�<ծ�17�'�!��JF�$uy0�O�"TF��фF�!8�Gs���ͦ��ٴ��	ǃcJ��l��̓%��uS�K7~�н�0i�'JȜ��	sy"�'��1�f��
Q"U؜�����Pl��9kdڠ��ISz�1��1ax��Ț'F8��E��F��sd,"�TyQ@h*(���;���#�lٍ3�ʽEy�ܛ�?饷ij7��O��c�uB�Tۣ��V��仆��<	����(��uY���[�@<;T,�LTE�	@�'��7͌)N�y�QG˩L�|�$��3��n�Y�'-U�2�]z��JG��;h=ɘW/Y�R����6�y� ��;�����t�^��C�:�yB*A�E�Go�s.�=�ҨF'�yRl�q���hfˍdw��R��yR�A:�M�r-�\W����#�yR��6^�5!���5U6���3�(y����|��T���'��'A�	/%B�L`t��W���ڀ+g�f�[ ����(%� �ѥ�Jt��ɍ2�"q"��X�J�@�mմϨ]�p�^� ���	ؗ�F5�J6��M���کO��!�x$�dH7$�I�"!16�'��yd$Q��R��p�I՟0��G�@1�a����
X���bVQx�`���J- �2�{%&��$M��@����Jߦ�ڴ���|B�'��D	
)q���DHk�p0q��(�*q0����u�IΟ@�	ay��D�9���g
�U�Z��t�ј->������I��qF*Hz0az�ė<<��\+�K�-�l�ؓ��,)A�	Ȗj�!�L{����ɺF�_��"=9���Yvt�f�+�0���#al�	��M�-O*�$�O����O�D&
CCPS�L�f+By  G�g�<�Қ8�. ���T4_�*��-�M��M���G��L m�B���s�d��FO1��4rm��F`��Gx
� �iE�@��U0A\6č5�'A|0���T�<����� �ݓ���-?:ax2O��?Ad�|�+�-ݜ\ig�Z-w�W���y�d�>I��[�p�v}��M���?q�'A�s�:\�������3I>aD������O~��je�+C��!��^_�R�
�O��� �)�'M#�4Sˋ�<@�I3#��.!���'>^�����\�y�BT˛֢��x��'&<,��O3ɧ�بՄ�CJ�aB�L4[�(9V"O*}X�4<G��!�3k�0���/�h��DR/݋h}�8�sAқ+Ű�a6 k���O��kt� �3}mZ/s��
��4
(*U*ԭ�+�'o���|�(�.3^)0�![	P�l<�<	0�VP������X@֘��
;@Jf����[��:BJl��5�3�,_�����@�>�A"�EŪ�0C�*��РcJ;A���ʃT���Vґ�"|B�-T�\��ŗl1h�Ye#�%+��ոi)a|�
;b���҃ͬ#�Q[� =���R	�'�$󐠞4x�a��陇���q��P"�x� �4N�]�L�yK}2�Lі;�T�b��UO�"FZ�M\
�P���bt�3mD��ybJV�&�֭qaaǧK;��"T���4ıO�f��u�'�PIrj��J9��x�L.N�D�K���D�O:��O��SA>�$�O�4���oi�Dc��"��T�[�\Aax���#����;y��A{��'@��N�=(�B���L�I{v�(�r��y����M�X��aIK�o6b�E�^+�
�a�O�<����=��T�t��ܓ�̒iu���f��"�?����D0��|�d�'X��B��j���L�a��R���ē�E�9lZȟd�'��OYL�H���7`O:p�&V9)U�p��h�Ǭ!�S�O��qK��g���];�+j ?��N�i���:X�"BL N�AB���'�Ĉ���������O&�%�"|*%ܢq=�8����p��R@�Bs�<	��M<@G�d��
�,OJ�z���d�'��}� �H0p̤۰�C��f�B'��"�M3K>լ������I4H:�iS��0#�iYs�.s��c�t ��=LO����u�(�m�"0��ʈ.|az���#P��\���c@0Ⴏ[�:��'H0�����Ϙ'(�Ei%��a~,5���;*�4�
�'��d(���,�(}⍄r? �)O�!Ez���N>(��q'�8z�Q�d���� C�O����O��<�+����
S�a��h���E�g �T���� �y��~"N�%]t����Jl���:f��M�PaBY��}�db�E��P�#܁�^���ˌ�\!��۲ b��$�OX�$�(����$� ͧ(Ϣ�І+��{�|x��(��?D�dAm�T��a�IߗȢLZ�;��覥�ܴ���5A�p��O��	�Z�x�����F�,��Q턇2K����<���?q�Oᠤ��?}��'��z�iXu��%ٔZb4\A�3�'��4�Gh�.;�ت�,W�fn�7�&X��k�F�`�
T`G�ܻ�ax�h_��?��j���'��`�KFV�0!��bZ*n(��V����O�S�O�,��O�T�Z h�g"���*OX�=�|bղi.�a�1�H,h��2�t�oZ|y��om66�O ˓����O�(�d�� 5���LU^����O���N��Z�`A�ZR}2�'u��U1�,2��E��$�j�4���/ ?��.E�2�0�c�eR�JP1��T\���⎄j�vq���>�6������$�Mӱi[r�ӆX|�9�Z�3;JIS�o� &+L�OR�d�O@�=��Si�=[�U�����0u\ mD�c�|�nq�I�?Qd%زK�D���:��U�%�U��=R�N	�?�g�'�F�"L1��X�/'�f��'��X2�D/]T�
�S�^���'w&�3��@�p���B�Eo�A�'Rr1�扅"Z����%O֪O�J��'��{5���m��	u*%r����'����e�:��\a�l=B�Dؒ-O�y��'Լ���A�+wb���?�ā��� ��S�Hׁl$�+�"��d�v"OT�CAR�\�@�[�S)k�8�&"O��Z�(��Do��cЦ�  �@q"O�����o��Mq�D8i����s�'f^=h�'̂D@4�#f����B $a6�k�'�"��O�]N�i�G��u�M��'��rfB�^h�HBh��?�p��'����7o\�-:�$�f0��r�'Ty���T+R+�hd���!}8���'Blj���hc�1D�Œ'�@���Z�$Q?�AV�P6n�l G��N�\��O"D�Ԣ!�1�E� R��h1SJ-D���c�*#��0��D�\J朢5�-D�� +�u@�p�N·j^�<�u�6D�D��/ԠGo���H@��a#�4D�� 7�Z���P�B�`1Z�2fG�OP�Z�)�k�<�h��S8_R�*�N�Mn����'��}iȈn�te��,��Q���' N�Y���:o�h��J+K�����'o�����si��P7��D���
�'kB%(��߼A�A���Jz�J
�' L�b1���kD h�.�F^��A+OP��W�'	����/>-�={�FV�:�B���'�X���G��f��pU��-����'W�T�Nʐu%�x9�H@ #6t	�'�T��#h�8`t�4(U�W�J�ш�'�I�ӈJ�H�4Mʄk�n��@����%6��,����Ju*�h����NlpH��K�|=��Z�B��=D���T��KrlY/�P�ʴ�h)���F�v(���߈E�l�:
u�>u��vy✻ƎY�8W���E��3����ȓo/�����ƣD��m����B0F�E{4ݨ�������Zc��)���	�t`�U"OFy�#��*�b5:f̅=i��G"O2%��hZ�7Qx� F��<�L{"O�uZ���GPX-y����Q⒑3c"O��1%!��0�R�Šѹ&��T��"O�<j���;=\����.��U.����'u�A(���5���C��V$=R�s���(���ȓv��\B��U'm�Ƞ$��R��ȓV�����H;�м�� ޞ6�$�ȓ4����D�H$4�p��
��4��o��$
���F��WM�f�指ȓ+<��%BH�۠�kR%D�
��'�x�o�^9����G��BL	S#T��Z~��q�jH�D� ���S>=�x�������X��9�Ro���ȓ1$�����+e�`��A����� E�<�WL�e�i���;�T���De����=�j�I�.ʬF��:1)ՕZ�B�	)_�ܹ�)�5���׀��=B��!�XZrL��@���#pb�nB���nɱ�Jܒa��aE�ҜjFB䉛��;� Sl�|b�*s�NB�ɲY��Y���D�!s�1js�=�G�IW�Oh�اgŀ%'�\:U�>��)�'�0mi��4ntb�`eT�bm"̀�'���)u"�"*�pA&K*iD�A�'*��@TgS<��� "��n��0�'��}�c�R^rl1W��kn����'Q�=�����a"�U[� �d�}����Dx���!�P8��m5�v����W��B䉻%����f�rv�@��㔺��B�)� �ʲ$��-7�|���2�6ݪ�"O��*ҪU`�L�VcB�IRJ�	s"O��3�O�%
O|�`��I?<�DP�"OXX�D�
MP���G��,W9���sY��b !�O�����i�@$(�DX�1Kи��"Od�*eL�K��@��#�.oܼص"O��*� ]�"�*�x��A><��Aa�"OZ,�%�Ϙ�n�2#�ǸXVB�!�"O�E�B��J,T�RK�]�`qhs�'c����'ˌ�t�@ n�h��L�}�h��'�4�@�7&� �+
KFN%��'�\T"X�;���'������'2��vIM&a!ށ�u�X��l)�'K�.9(�4x�a�(P\=��Hh�<�D7x4JUR&i̥T�����b�'u�����)�
D**E{'B�n�R�������!��A�������Dq,���bH�@�!��֟nyB,{��J;�8�8ϑ#j{!�D��q:d 1�B�v�����^��!�DO�c��[�Ϫ���g�<�!�d\�6�ԠBS X�R�V�RT	!R�r�ҕ�O?a�3��2��hp�kùl��9׉�Y�<�B߈�`
���;{�0�V�q�<	��=/N���'B8!�؉Z�-Mm�<)� �W���2�NY�#�h�<i�ӻ@�n$��	�ܢ�
�~�<AUi˓ Z�}zR�N0g`=�G�|y���p>��� ="��@#a݅6�%�d#|�<q��/���QR�@�����!�L�<�c�I�<n�;Q���2�D��`c�`�<9S,�+n�f���՘i��y��Y�<Iшڒ7�ޑ!��֔ i������Vx�dbgc�����A"s� ��)���iQ! 7D����hY:7�
�T�Y�G_�%��h'D�|R��K�b�q $�7I8^�Q®1D� �W�	(�0"�˖,?�^m�s�3D�S *����X+�j�1G�E�@,D�h"�ً�\L�K�3�D\p�,�L�d�E�T�E�0.������bSb��y���j)f�b�Z��Хz�-[-�y�L��m�>���;_h�3�O�y��#!p9R1��7o����yAJ�ĭyR���5Hx� �_��y2B�&*�5�i�-��ࡌ��?�U-�\�����x�  1l*�'�NH,8Yǧ+D���)P=]���#�
ȓw�;D�L���3�b�r���/M��0�'D�x�t�
:M�EQ��-���6�7D��K��	G�a
�c�rX��V	4D������?Kw6�2JJ�s�l��c%�<!��W8�����ǓA��X�Ӭ�5R4$��2D�TB� �~Μs�N��S�,0g/D�XK )L�I�+�ޥ;vN�	 ��#�y"��b�1��H�4�5E����'���-�5G�6�Ar"�&3h���Y̖`��q; ya�	�K���'k�7*5.h��D�<S#�V�+:��qbj�$W,����(��CP�6�Ja�g�U��x��ȓ+��ж��lD�.��T���^�Z����wl~Db珓��d�ȓ�D)��:"'ܠ�Bfw�=F{ߎ���BT��M��0�p�a����?�  ��"OD����25�U���u�J��"O*�ŏ�90ZF��$дq�"O� �`����V$pQwB)un�)�"O����_�3Ѵa�1���M�L�"O�@I�@�oҤ��u����VQ�V�'�� ���nR(iQ���4�xǈζrunфȓIc��1��TB�Ѐ+�lٮ*nX�ȓ:��*��Oc�u#QK#?�y:�hd��TmMc�Q�h�p�ȓ5c��W�E�d���zT
�&��ȓWX��Ѱ͈$ZN��r(�;	4��'m����1�d�Q�c�¤��=���(�9�dMQ�0��kĮ�8�ȓ+�Zmӡ�Y�&$�Yڱ���Tq�L�ȓB���CB
LI����'Y$����E��i�����nd���$蕸`�~0��IC��ɺ1`���h&ec$�;�O8$C�I�zd�����,��|�P���aQ&C�	(`��[�Tl�m��!O@C�	�-`h�;ƩKK��h��n�bC�I�^p�$��-�
�j�h	/
�XC䉔v��BB+pN�UxC�ţy�$�=i�J^b�O�~DxTHR;<N�B@&�1� ��'�x�R��6e jL��ɏ
n�Y��'!|����[�_���O �-��1��'P���4�1jAR�C��Ѯ"ef(��'�0Ad���=�mH+c�q��'�<������7����H�i��'��H����S� ��C��mp�c��2Ķ���X߬�����<��aDP�>*���g��IRg�7~,��s�KM&#����N Խ�� �҂ə��Q:$R]��Ғ�#��<^�������6b�]��@�A��<6��h��Ʋ*h,!!���	2����q}��%��m�d�c҆ϋ>�!BG,=�|B�I/�tL��k��|��̚��C)bB�;7� C�L60Yƕ�WH�^�C����y�C(!w��	�
$j�&C�	�?�`mj��D=t�-JѢ�u�RC�ɉu��X���5�Ƀ=Z*㟄K�4�S�)��E7^8�K�3]����j�55�!�DY����׋�<S���ҭv!򤏭w2���h�v4���
�'c!�>xٸ5['HЙ4��8�@Ћ�!�S(i@���O��7�H�k�!�#�<�H�KO��Ua�성�^�I���"�g?�a ��B䈘��G�� �-���V�<Q��@q��`qdH�tt�kw\]�<1R`W)U�������+ U�#��W�<�P�\�EM����Uz)�em)D�<@A�I�"<�p�EH	/ъ���*+D�ȋ��
+�6�	�'D�!y~��Q��O�]KE�'��IIM�\��P��cЈ(jX�
�'�\�aH#�t�A 若/r��c�'.ĝ	�;l��q㋨%�h J�'84���"�N0P�Ol|�'p�Iم�%2�V	"���<�� 1ߓO��O�� 'dK�����ǃ�"(nؚD"OH��7�m�]1&�\�|�z�Y�"O�؁��>d�09��C��bl��'q�(�����p�~��'�A�e�8�Q�'�j0"h��r ��)�P$�'�r`a��K@���8gMʬ����,�#�O�'f= 0`q$��<5�ja��ņ�`+���a�ٓpG(���8+����^Nɸ� �7RH(<�� ��1��S�? � �b��@�)7h\�V��"O �xcCX?W�N���TgB^ �"O��sAǤ`6��`Z7E$d�2j��O��}��XB�(Jwdֲ(=BA�%\�2�8�ȓ\�:��o�z���ˡ
��f���ȓz?
���E*<1�S�IԨ�l5��=q����g!s�d���f�xRbP�ȓoņ���T'��r�J�, ����M��� �@Z���!�.A�h������~�����Ff߈����-.��P�k^�\�!�d
+d��8��n�:f)���
VVL!�����p�$�ɵW.�JQ�b!�d�2&>(e�6E
�g�.����ho!�䀚��d��L�{����n�ł"O:)Qrɍ�,�(�v�ŅPъ��f"O��[bZ.G��ق�[&a���X�"O���V��H��g�<�LՉ�"Oz)�T��Y���� ��W����"O,��/Y��(�%�N���c`"O`s�m�1b��j�
��|�����P�(���ؖ'��j̧�M�w(�2w&<�E�V'`:xp���$�0p�N�K{f�W�Y���Q�?��@�	B̧/5�����Q��L�d�B*O}*��C�i�j�	��P���'���'���hR��%�24J��P��
��,���c�.�d��z��y�P���?7��R ��5f �L�­����I�����H\2@����� �Tʅ�<aXwVr�'I���'���6�D��6�,4̼l��ɦKu�mi��'^�ȋ'UB7O@���ޟ�^w�P�'g0.�{V��T#܍C���	 ����>d�����O�8��O���'���O�b���A��3Ī�QJ�|j�d�
�H�䞳CSr�'��g�'���Q����u7�m�Ѻ�Nl���PD]&w� SeGeӠ�	�k��D�O����?1������4;:��a�
�@b�][���XLfy����<a�Fʟ��'�u�'�����is�,�Q�(m�T���W��M���!1|7�m������O��ď"nv�S��G�ޝ�C�R�2M�u���C3^�`�ߴ2w4�!�'�xx���?!�'�?�'%��ɜOu���!��nX����Rz�(��i� ��'�������)�>I���8-=2��1i���X�o>B�I-A���N��Q��B� ^�26m�O��$�O��d�O��D�O���OZ�D� �αp��
�-�r���V|��m����IMy��'��O���;}�
��B�N����$o�,^��b��'��Gy2C:]�2AC��Nm�#R���y�iE!�89䆆�sgP�S!��yR&��L�hc]�8�t-p@���y� ��y� �� *[��w�G)�y2*��V�#7�ۅ��jF���yR"�oR�Ha��u�%���y��A�P�ber�rL��H���y�h�<�������J@Z�[8�yBa�,��9�Q��aV�1�i���v}��Ò�o�h���E̝Nхȓh�z��o�F�V��%NN�=O�$�ȓ��d��khIá��fA�d�?9�L.#$�#�4%
Ȑ���A�	۬��B7�h�"��8Ir�ٰCH��3�.X*P�s�F�/�$�bN���cf��"}<q3DG �l�Z�
�4l}�Y�ņ21���xR�R|((����SxQ���-!���dd�u#٘����XQ1�|��� x"�
��|T	�v��y��+B9l��mt�l<����y�OS�'T�\ٳ!��gFp5ap�Y��yb#N��čS�a���*��5�yr'��[�����^�'��`���R��yR'�0tc�DK�
��%.dy���yb	�}����J�|x#�ފ�y��Q�K^tܹ�H�DU9��K.�yR�� 
0�\s�����uH�cͩ�y҂]k��0��O�>0�WX��y�EZ1{���c���M)���B+Q�y��$'̬��Q�R���Q�E��3�y�۪_�8��v�ȕ=���v�6�y
� �J@E��RS���4���|��Y��"O�ؙ��I�e��i����znX�Hu"O�|ja��/B�����Zk���"ON!�Se�Uj���-R (Z�"O�2��S�\�ӠBT�:�B1U"O�43��O2?�azq�R\@|U�P"O��7ODZ���8KV�P��I �"O2��T�.�ȟ�Zj�!"O�I26�?L���Y�&�xM68)�"O�tp`R70.>P��E���٩�"O����*
�5$��Q$�s���&"O�(IakZ+�2-a�����HG"O�5c
A3�	q�B�-Q� I��"O��(�*J&D�Ef��h��(�"O4���C�L$!1t⎚¸]�"O�ͫ3��4c���s˅,>��3<!�D���RϚ*h���1d
�CU!�dD�hOx�J�(͜U�&	)ͫ\�!�D��J����b�Ѻ$��!)�hͩ>!�dI�Im@� ��CflNt�@HԤ�!��Q�Dm&X�fL�X��æ��'�!�d5@�HQ7ꏒW>�(��%j�!�$BQ�4@���k�|��$AW23g!��& H�����ޮgն	��N�-H!�� ~��-Ps%�}�:�Q�-
11!����x�TKK�����Ǣ9�!��,\3r����I�4�!aƫ!�$�5=.��Q��P,?�~E���G�!���"i���W�&f�=�IEk�!�D��k^�&�Q�@I�e��,R�!�$
tO��QbȎ�j� Q�TH��}Y!��Q��f�#�I�>D�6\	���^s!��>�d�R�ֱP>4%�����k!��q���5m3ve��DK�m!�$�'Z�}(梐u�����/g!��l� ��'n��K���� �
5+!�$�7:�\"f��!��lX�Ȍ�mo!��,290��A�]�>��fJ��n�!�d�΢�����$��8��HE�H�!�)|�9V4��tYg��#.�!�$յ:W��
�(W2Ր��9sl!��ݐ���aǗj9�T[��� 6!�D�3<D�#F�W4B	��CS�	?�!��wj��Z�޾�������!�$UP�|��Πp9 D0%�ĿO>!�D�>M�@�u�Qb��.!��Z�S@� ���u�!����T�!�d̰|���3ժTJ�`i�%]��Py2퍒Lp}�]S�-�PaP.�yQ�U�pd���"J�X�G�ۑ�y�n�8�&x�S	��:�N���d�6�yB�-��)�ր� 7f��E�Ó�yr4�I��E͡2��#P�Ý�y�3�r Zׁ[�8z,X�.P�y��⽀�E�=5�\��F��yb��5��e+��Ћ]�ȓ�� �yBȋ9o1r�K�kT�(8���aZ��y�e�9TĘ�0�E''F�D�&�C��y�π���`�E��4�x#�͙�y�Z�zx�2c��$��2-��y� �:e]��Rb�x���r"��y�K�a�����A�o�zX�@�6�yɉ9X��B*
<{�AP����yl�(�u����&9�$�ѣ���y
� �X�e�2+�u�%�_�U[��	b"OF��R�mS6�XrjF<�D�;A"O:%��q���y�
��v�� "O���t@��J��K
����Ʉ"O�y8�$Ƌ+R��Jt(�]��}��"O �`�����xC ��/W2���"O"���]
���Cń�=m�H"O�-� ��h:%���;wr�ó"O�h���ѹD�لb�_��E�"O(1j�'O�z�v�rt"_//�bԒ0"O�Qi2�x��@IS�b~Z)�
�'��9Q!GT*+�Mۀ��0�y��'(v8�B�ȼ6��9 ���#-�d[�'*�p����Sl� e.ʑ�H�#�'��ct�ݵt�9�'�Bw��)
�'��=(Ba�Pft�yvj�g:�=��'^����) �z=J�#I^U�'�D}!�]8��I�4��-�te��'�,]*�c��������0��|�'�ƍ�`ưYF�x�TFG�����'�^��G(gk��#!B����'��Պu�&�Q��-3,�C	�' ��l��3<�EJ��&|�L�Z	�'��g��RA��c���B����'�NܙF�53,�Z�ͅ*d�����'���0�ג@�(�����^�4\��'�Cc>T�l�Y��4�D�{�'
@�!� S%:eaၬ4� ��'B͋dF�
K�4�x�Hă<�ʸ�
�'�z�2Ύ7Q�$�3ć=6(�"
�'Cz��KU8��Sd��
Z6t�	�'|�L����h��L	�|�2��E�<Ypl
?�v 0ƐSl����~�<�Q�%E,�:�&�U�2�t�b�<)D*Z�RR��@&#P�M���@�.�X�<y֬�25/�I����+UѼ1�+Q�<��P�b������*��=�roXG�<�-̙F�^��#�&.����RF�<Y��~fT���R�8��e��D�<���Ђ�����D�>T3��D�<�s�޵+o"�j҃_	6�R|R��D�<	��T�#�bD�燈q�� kU�@�<��ŝ�Z*��N=H�`�W/�<�p��u��� b�Ճ~>y�Fw�<!u̞"!���-��sw"��F+�{�<A&I��{ڜ��(�<e�N��(W`�<iGcҷ<�$�`�D�)�-P�G�X�<���5I0��z�AKk�fyB��J�<�U� Xh��ƟK䈈��)X]�<�bjpL�#�FJ�z%%LW�<�ǅ�h�@aPb�v���S��T�<��W�\���cU�!r�`�	B.�R�<y�5-"�яßC�ĵ�s��W�<C��h� ��o�_�LQW��X�<1s�˒/�Hid%A�0����s��P�<9bfJ}�t��xlv��g�L�<QƭO�*�4�q&��iP>HpVJ�<i�I�:6qa�*[J}�t@�br�<F	��Y�F4s�(I#�L�x��s�<1p	Ė)(���t߻m^JM�e�q�<A�C<9zbY�#NY��8�'�Bm�<It�f�T8�g�<n�5�u�o�<I֭ g$���@�d��Q(���B�<�t�Y2C�~����Tz�A@ge�|�<� �5y�+��4��U��s.$�"OH5��� IC>��A,��^�	r"OXU��k_�8��h�'��{r"OxlKrh�1ur)�-�#x~�g"OLxل��z\�0��O|�RQ�1"OlU�	Y�:�^�1�}Ӱm�%"O�I��
20lِ�N�]��4�3"O�`@��O��Q��6 �q �"O�I�t�G�}�9'�>�!F"O|A�����z��e��&�$f��+�"O�j �1y5���F�>lS�{"OP1
\_1�j���7f��"O�5#��ɩ^�I�`���R�J�"O��K��(� ib��`�D��"OR�2蔫4"!�D΍x��H�"OD [���:xT%���N��S"O��(`�~1ذ����6,B�9A�"O�$���<��`�޲8B\��"OV]��0�����&�,\zԐ�"O�}����p��E`vD\W�	��"On�0F�ݢi8X��bO�G��d�0"O��Q�"��2���G�������"OB�Y�+�??N&�J"C �B "O�1c�
��W��S����(#"O�ѓM^�]�hP@�ѭ	��*P"OxȘr�X9}R�$��O��	��"O.���F��o]~U����V���"O��t��"5�� �5#��Fb�X�V"OB%�a��(Z�B=�왱?^F�S"O���sĀ�8�Tpr��ɤdC�h�t"O,�:&�ڳd��U�e2�D"O�D0����b�u)��X�~��M��"O�;`�I[�*yc��
~��"Oʨ�F�J�E�(!�� D��a"Od pǪ�4���ņJ�x�V���"O��#`U	w���Af7vp��"ON�Z�>j�0�9d�P?X��"O���������������"O
��eY���MAV��4"O�YHf��`Q�-���A�EѨqy"O����N��GѲPx�͟���H"O|	huj9S��Q���o��L�P"O��c�T�'w����i��S�xQV"O6�2%���(̻d��8Y��P�"OD=�&KH  �2W�P�8�jH	�"O��L?*�X×f
Oۂ!Y�"O���w�H1D+<􉤅I=��YS�"OT�cC	�6v�fQ	��þR�� �"O�U��lU�&���#B�
m���"O*�Ҷ��&Q8d�S��̭�DQ��"Ol��C�ī8�TY��DY�7�z]	�"OL��Wf���d����-Ԯԙ�"O�y����04�H)ySCv��(q�"O�}��g���� HB�>Β!("O�1SíC�6h0�Г1��"�"O�ya��<t�e���� Lҥ5"O�)����/]ƴ�ccZ}G�D���$�����TKY6n��3�a�8��'���"Ad:e���"gS�n>��'+n<��݉,��UC�d��)Y�'/�];�Z9��X�W�V�nB �x�'�ּ�@Q?ln�|iPO��g<�)�'5^w/͔��`�E�cg��;�'��`�E��vzV ��j��P�x
�'���d��6?�%�����[r@U���� P��LÊ*��[AP�҂"Ox�c)�O�"Հ@����t"OjU	�@-P8�`*sg�8���9�"O�a&)
�1`
���Z�p$�"O�$V�@5�~ #��H5T��h�"OtP"M�b<A����i�|�i0"O��)�'�N�*8�äM8/&�0r�"O��Kv)�;b<)fD��S*���r"O��g`�(����*�;G+D�c�"O��bg��z��
d*�,Y ���"OT�{ h˥��q�j�"�dЃ"O:!��-�Pې���ʹ#�NT��"O�c�a�-&�A{�N�6*��rp"Oj��g�>g�tRƮJ9���i"O1�.ק&�<$��v�؍@5"O�d{�)�3��=�&��\UpLrr"Om��]���}*`���obB�	F"O�<��-&b�����9�"1P"Ov(vgJېౕ��+V���V"O~,��WfS���ρ�{�d��w"O���tȟ���)�ωt�2�8�"O�jK���胷o��D���V"OTey��Y
�t9�HQK� �D"OB�������,���ʀ3X���*O��[�-�H��܉�ܾ[����'� ��ܥS�[��C�J Y�'����!�z_����F&��
�'O�� q/� 3�u'��wxn��
�'^�,���QyZ|9��y�X���'P�0*�S�jNb�ڤ
��C�Ph(�'����#�;[~�U�!/[�Ag܀��'��!�3!��W�H�"�AFq���'<���t�F��|��ʕ:D>���']�!O��F�z�E\:hڎ���'N�Uk�Ο�Fd[�J>f*�1����O4?�iab��nv�	g&�b�<��9u��h���h���®D�<1�]ʸۀ�з3�͢�_A�<�!/JY��J���^(�\�<'�.q��a�f�)��Y(�+d�<!%��	�H�P�@@މᓫ�c�<	#� =Hٛ�L��[��E���t�<� ��}�r\�vѦ�!�u��i�<�2l�s�r�"@��9���2d��@�<�W�\4g���)Am��Eu���h�t�<��̋h.��tǊ+^�896I�r�<Y�IԈA��\�sjƒ�"lpI�e�<���X�<�pZ��Ն�DI Bl`�<��̗oD��b� .�`���<��Fər�`�b��B�h�*��E�<y��جq"n�c��fk
��QF�X�<!S��.�!GD�.�\�x�\�<�gI�)G%̻�Þ.D�<����UW�<Q�N�)X��-9�,�:��SE%@W�<	�ծ
�|�!�eĿu�XU���\Q�<���|���C��ih����EU�<i���[��A�M�=���1�e�o�<����.]��(���Ё	U$k�<�ģO=N&z�` ��z]���b�Fc�<Q���$B�ʀ�hñ<bly�n�h�<��ԍk:p���ی,�nQ���X�<�򯖣n���c�N� 8�qa��Q�<����2wph1f��'��2Ǆ�h�<�`Q
P�|:f�$��ӂ�`�<� P�r��_�V�P�d���"O���G�����:p��">D��� �&����e	�By�p��G=D���`hȵZ�bցV "�����9D�t)�֙B�0��!�("��6�*D�P�,��V;��s�׾b�	�@�(D���m �\�1�҇}w��6D�@��C�,�Z�j��%6�(q�q�5D���0IL������O)K�zT�)D����_0<�TLH��;>|2쓅�(D�8EB�#�b�TA����4D��)T��*'U]AG�Q8��ѡ&3D�����&B�TZ"
u��qj6�?D���$G#���� ��!@���?D� ��	�ɂ HЧ�}��I��<D�<	�R�*�Kq�T�dN�`�D/D���5�D-Z��q���Q�6P@`#�9D���Q���(찰z�͒�UX�́�"2D� �� ���S%�ђ2?leP��0D��P3� :^X�{@�P��F�Y4f?D�y�e�N���g� |��C�)D�`ɒkH�}@�-��jɑ}&�"7D��yP�"D�$�BV�ö2=�Fl5D��c"i�;`2��F���4�����'D�0ӱHЖT�f�q0��=�@�:D����'�D�n�!����8���x��-D����ۨyl]Z��7-_�@ش�-D����г/�<�ZVB�����(��6D��B������1z��6u�beH�i?D�d��D�9Q~P�+c-|��q)[�!��R~���h�$.=�E�ֈ8�!�$ӯ������	"��SGo�!�P �u�䢚���Q�1�{}!�K�(�VA�7O�A��̋�@i!��u��y�M��-�nMY��K�M!�H�t� tX�H;
�<r@�+0�!�dM>ReJ�b2�0.��:v�!�D�M�~Q
�U*��A����s�!�d�;1����oM�x4b�&�;�!�d[()��=S��re�S��;�!�%n7r��Ü/w(@y�I�"4!��@�x�lx��N�Q�l��"�؎#$!�$�,r젲"I�D�2a��@�!��V��tbS"�j��4��(O�)�!�	�m�)�����~�sD-  �!�ɾ.�T��R�I�\�(��,��(6!���`�c�̰;0�<�3���C�	;�R�)t)@�Y^���E�-�B�ɋe~��J�ϊ F�����,�B�,̋�C�	�^�B��4*c�B�"t�.uyp��'�>t�Z+4DC䉕m�X�HNJ0�nE:d28�C�	e~���2F0�)Խ�B��2j:��+` _)L�Dief�~�B�	�-��m�El]��qU��HCRC�	�SLD�й0A�f�0TΎ�A�1D�X�@cЩØ�0�#uHL�tB"D����lT�R��\���SifqIT�<D� 2�-��<b\HD��&I��a���&D����>n��aW;?�d��!� D��P�M�
�({�e�����h7�0D��Ӥ��E�����S�]2*̪&0D�P� V3/ �e��S�"$�9�`�8D�� LכE� -�`o��B�<k��$D�� v�E�h�E�W�NM�Ѓ�"O&���DF����ΰIe8��T"O|�0�/�f����<�B��2"OZe�S��۬��&��/:2"Oh����N	(��3��(��:�"O���GJ�$��պa
ǝu:�*V"Oڤ��#I(s��k6i�3C�-;�"O�p��C9�j 3�ńv{"�"O�����"M�0�c���\`d �"OH�a�K�5<~�Y0.X�3����"OX���f�\MB���&
K>|��"OT��`L�A0���W�����"OLI8�څ:�戹�d��B?,��"O:��cD
, ����
V/{B0��"O 0�2��/S���p��M&1u>���"O�I!��9��Ͳ��$.�$���"O��#ׯ@����Ri�x�&�"Od��`�4.ZT�s��0J:RDq�"O�L�U�ҽ3R���%fť'>|x�"O �⠀�_12%g����H#P"O�0C@*
X-�YCe��tS�9��"O��CBg�s�Ґ�0e�_����c"Of3�|��
�$�$Ԭ�c�"O���Gдfi����DB�\<���"O� R��4Oyv\y3j�wx�q�W"OLlxd/I(Z<"���J TY���%"O�R���D\FM��ID<YF���"O�M���ß0� �(�ț�b��`�"O�͘��A:b����o��g"d��"OŐq/�r�N`'D��rH1(�"O ��v#�5&l0�B���W"OT�s���gyxh�n�-2��
�"O��І'� ��#-�?�@�e"O���rkV$(��K�U�`�"OX���Ν3_k�كsm�{&48�1"O�=���Цhj���*�����"O����N߰%��`�eMά��`I�"O�i�+��tZ<�[�#H<D��3#"O���r�B�]Ƕ�"%6T�ё""O@xK��ϡu��`�bLKT.���"O�e��*�%zzj�8��\�X����"O�[�E@�um��C	�
C�Yx�"Omd�	%$�x�A-(B��;�"O�Q��+̊[�u���֛��ɥ"Oj�vN�(o,6���L� ��x�Q"O$�ä��D2��j�㈛ �tzE"O.x�����K�]J�"�k�V8�"O��:rO��z`�$a�ƒ��2"O�p�U�sXJ�:Dg�j�Fx�d"O�;PE.b�2S�ܢE�ؚv"O���.�Hp��J��5B�"O^I�:O)���C�{�{s"O$��,�:eMd��A�S8d��"Ob}��&R?�����4g6�3�"Oܵ"��(1(��9��G`'\,�b"Ob�!��L��c�Hx�Q"O�Q�3��!u~Xx(�� �ج�c"OX��C��.e��mi铯F_Vt�0"O�e��O
�	�H�u8�H�"OV�H%@�f����Ϟ>;4bi �"Ov}��(�.Y5�h	BoJ4�P�$
-Z�( ���f��ɫ#CC Z�'���QSo�z:ư�R�P�U�l1�'�܁��S�Rs��x�,F8Q$��'ń]��n:wl���q�BV����� ��'N�)�� '���0L2�I4"O���"���g�6库�38����"OP̐��Ax��� 7#����"O���@$��0 ���_2v�lk@"O�<z��=h��x�a�N0|��'�X�[���8�pX���n��'�l-2@��HW�)b)�PT&�b�'F%a���O*,��w�.Lx6���'88����<,�WkVG�6x�'�I�p�*Q��S��˛D��[�'� ��%J����i	S��A�Qh�'f��7�J�%`�<("d�4b���
�':�+��1atj��q��Z�V��	�'��,Q�m��t�m+k�&&ư��'�D����
W
��c���<���'�"���N%%����臻_]��'޶� �	�!Dt8C�]Tʠ��'�ȭ��Ce�<k� �����'��XB��-v��9G�Ο�@=;�'��!��Bĭ!/���v���x7p�x
�'t����΁�K0Y1��7{5hT��'@�,KV�W���(!bB�;b�:`��'I$�8QC�7>��dj$K��
�'�~ɓ�˟']���3tNԺ ��3
�'x���P+��4<�YV��y� A	�'z<�؇����r֧HZ�����',"�eǇ.aw�I�vL�Llxj�'�va�C���^�t��	\6V9�K�'T��FbĠ�6���@Î5Y	�'_.����9Zޘ;T�_�bx����'P M*E%Q�zf�}h3d��C���'M6���b����KH��A�Zu�'�ZͺW��+���ɑ�7�^�h�'���ڰ"��A�IcPe��&��'q6��7��A���(@_N�0r�'����Я�Ql`S�H'�
(��'m|�q��׊~�ޥ�v	�Y&P��'Դ������_g�l+��A���'��3TD֪h�LH�`�[#c�Q�
�'��'h��@�lT�p��1��Q�
�'��Y�aɍ*v��g/�0�F�
�'`�w�[a:� g��W�T)��';�,��V�\�v�ӧT�fD�<i���l9�4���P
�,x�%#K@�<�Tć���	��W� ���#q�C{�<b.��V��m�o��+vg�B�<��nT;2���6�G�V�K2�W�<�qjI�MJX� k���B�ccBS�<��J\�D5\�j��n�Hp���R�<1f�l	0���he<��v�<y�`�
)[����3K��I�{�<�r,����AZC���x(�t.u�<�"C�-5�D��$�f�1�AmI�<y@�C�U���(�oQ|Q8%� �Q�<�D�H�/��|�j��Fl��� �P�<A�`ت>��`�O�<~|�cF�Nt�<�� ���X�đ�|�[�*l�<Y�)MC��#dض|L.�@v�j�<�%A� ���,�H��Hp�bP�<��%o�2�3Ǐ�S���"/�O�<�W`T,B�BE	ۊL�R$C��
C�<��e@�rN�@�Q@݅%]�+W��B�<17�N7R	Z��^�-���:P
_~�<y����UJ:���E��0�f9aT�s�<� &���0s�����	�)�n���"O���� <]pt�A���1U�Hȣ"O�9�6
�R�-SJ�.���Q�"O�bP�ߊI�����_�5"Ox;��l�Zԩ�$�@�"O�2�I�a8؜�b�4SI�@�6"OP�yרN�w$���PJ=:?�$!b"O�d �K���H����/y��9��"O }�$@1�j����8q*�yR"O�9Y�E����I�ɚ&� ��"OR�y��ňl����I�xT��"OPM��aܘ]	�t��ھv��$ �"O�a�+�/wW���g�0u�]�C"O���LB�.�εX���{hfypr"O0H�ϭ����$D%i[f(I2"O
%��˛�~ڸ��pZ�x�"O~��*� �D�J��N�LX��p�"O����|��@ϧC!2�	�"Ol@`#OQ�{�D:7D�v��l��"O~� uE:��]+�mV�S�����"O�H�fě#�&�a#͆ [~^a:�"O�pb6��?v$]J6�,uW(x�E"OБr�'�>
W�t��&D�ZV�%��"O@$pg*U�<\<xf�S�\ݪ�
�"Om�($'��!�fI^�T��V"OjAa��(��`��`��!ЬE!�O�p����:J]�E#RA�v�!�D^a)�Y(!�1aX�-�I��!��/&`)���y0lX��DһW�!�䍕|�m�ӡ|.��"�05�!�B<���MûLoș˖�^�o&!�@�2�RM�6�e=�0G�S�!��?�H�*�D�"�#���!�A+w5~%�u�I6i4i�[��!�[�ޜڑ�WJ[Ry�h�"R!�̬H!��J�̙�"at1i�I\�X&!�G�S@��u���U���qG���c�!���$��1��R�K�h�H`���"!�d��|M�惨[ܘ�ӇE��!�� d{�U� ���>�֜2���Py�j�s�:��DsF����yB�=F.���cV� L�B���ynN�B =�s�B�i�6�3��B��yJ�\��$C�-�2��QH�yR� B���(5�Ob�H��́�yb���<�˒������F\��y�O@�{C�(�K��h��_��yb�_�{��S�P�}���vo��yr�Մm���!����w�DI�.Z�yh����e��"�z��=2�\��yB/͞�]��R�j��ls��X��y���	G�qQF!)UR*���\��y2�7r%�(��MD\��EDH��0<!���Ըh�PPȥ�σ_I��L�y
!��O�H��UcS�;Mvus�
L$w�!��_"!+�����J*l �j%
͕FS!�d�߬��f .3����� �j�!�d� �Ƞ�fň	�ڹˠS�?�!���ox�\�p�T��h�C�{!�C@� ؂��ɏ-z�Ę���O!��]Gp��!Uf�+5��>?!�)j����)~S�ܱdA�4!��~1\�R4.@�S��-#� �'}!�D ��]����yx� �$ty!�� ؁:�:�n������ �
�C$"O윸u���U�ȧ*����"O~Q�ۛF��:"Ϝ�x�N��"O�L⑍�+���B�L<�Jt+B"O¬zF�p�@��f㞟~C�mX�"O���wO�3A6(�#cƂm7x�3"O*d#U�Ĝ�5���:$.̓�"O2�s�J$A����!W�U@@Q�"OT@�P̝'H��#R+��^�D̉"O6�sC��@D�@��O9~��qv"O��CP��g+N�Wm���`�P"O�a�Bo��/���+��Ҹ�&"O C犋)T\:lH�J§_r�)�"O29�G�Ƕr�L�*�J�6d�i��"OlY8��� ((�bv�Յ-}~-K�"O
Xc���!���GbB�8u`�s"O��C�6��
���n\�Kg"O���ǫ��L���R�@�I]�,p�"O�@�f�,�����0?X`yt"O�يe@^;�ؼ�非!;�3�"On-��Ύr�H	Q�.BF}��ۇ"O�\�i�&DJB0࠭�9P���
�"O�I�"�Qm�l����1f��p��"O.HP�.�/����#�JǰA��"O�T���6���0�9p����"O�]�F���S��Y9�F�*`����&"O��BoT+-�r���F�
�^`�"OVe���,=���`��:M�!�P"O�T@Tb�+-�qP"eS�E=v �"O�lq��1��8�U��,3�A�r"O��`%���MVf�����!.%�@��"O�=P��"Q�p�RaQ�8k֭ "O�#1���G~�����<[c��AS"Oz�{�$N=�NL�#k��TL�8�"Oj�ʇ���U��yf��`��2�"O �r#J0(R�,�P*[�}Ҥ"O���rML�9_��c+M�CF��bP"Oj��CA���$ 0��'D�t�"OH�"A��R�艢�n�w1�ڂ"O�ѣ�#M�X#\�qD�®
���"O��c������>NEc"O>��%�|M���]�D����!"O�=��`��L��\9� ��"OJKtc�"�n�P��0g�
U��"O��EY	h�`Z�M�a̖��s"O��� 퇸l�`qc�*Wcظk�"O��P�Ձ�,!3�P�:(d= U"O�H���(D��\�fX�y`��`"OL4���+g�ɓkP�3+ L�R"O�ea��20FEE�I�pz<��"O�Xu+J�.g�ə�E&Krƭz�"O:���O����
�ReV�q6"O���"�T�)�Z	iSc\2o]��$"O�D�r
� [���S���l9�3"O�9@4�8iZ�|i2�9NS �%"O@e@�D2YT�Qo�=}D��"O��c���8��7�.��,��"OI�JE�/E�l�E$�"OF�hF�Q�6Z�����p�r@:T"O~��
,�����"T��E�"O�(@/�:)`$KE�9>�3�"Ol�)��&B5+�ݜr���"O\x��T�~wZ��D��:.��UA�"Op�b�KM�3E�E���K� ) 5"O� �8�ҹ,��y��BC�3�r1��"O�x�dJ1Pڔt�&BA*�N%X0"O蔨R��,:Kj����)�~$@"On}ȶ��e����2Ǩ�*h�"O:�iFC�w2��2�Ƶ��-�w"O���v	Y�t���KB1\����"Ona���� ����YNh��"O�9gG�HJ5�3GӶF�$@H�"O@9��%Q����g̓<o����""O�A�DD9S@dё���6��u+f"O��!ߟ}U�Iqg˦vin�"O��8$�tC���F�,g�qC"O��3Q�[�p#BUɖ䟪+G�Qj�"On�HD&-jB��c)>_^��"O\��P���l��1Q
O>%Ƭ��"O�D�l 6
:2��K�Z��V"O`�0�Fw-�a��<Դxc�"O��XVi,Ф�ڶ`ѳd�d�!g"O��[��ˀG��e�7U�g�����"OΘ���ɳ�
���
�Z���I"O�uHB'nYu��Ф=���V"O.�s�j�41 ���)�P"ON\�V��%'���ݨ�B4H�H%D��� +���ݲ��%�x H�a?D�i�V���TVm���v���9D�@���Bov���B+�3�0mya,D�\���
K )���HF�|��(D�@�V�M�g�Le�Ug\�i��D{��0D�D����TOXI��W=�@�+D�\Z��0	��8b�3�آ�*D����n�MD�ɵH�p�����%D��s!!��TV a�B�)Ĝ32
$D�X���-c h��2K��o�Lݛ�@$D��"{��sr�((��pA(#D�l#�ů3���8�'Z�H>ƨ��� D�pQW�Z�e���d��08e�#D����e�9S/,D�tU6iF�=�2! D���� 1,��=C�CT�%�$D�����"̲�2F��"U���j D�h���@�R	�(#6Oۄc&f"A�1D� [�C��Fa���"O�5�JQ��m0D����,͘��ԾkB�Ų7� D��"&��>7>t{㉑�(��% dd*D�� so�-)=�l+�+Ϸ�n��*D��whD1L*���GI�$� ��%D�� �Ǒ�63x������Q+�>D���$�`�!�F��E��:D�h�%(<4py`%�-D��UȆ�#D�h۱dX$$~VdY7h.FuV�!v=D���/َ`�ع��a�~!|�2#�'D��AEL	6���g�?a���*�$D���֨.��\�'�ݜ&Kvm��F"D��rա�1)�b�xׯ!�����!D�8�W4��TϘ-Aͺ鈗�#D��3e�[
�� Y�%V&u���G.D��9.ׂ �a	B̉13�ޙkT�(D�(��!Q޺��䦛>9� �#�(D��R� �cR�a��N�x�2t'2Ox%;�F=Zb�y���; � 	�'�,����/pJ�� Ǣ�[��Xj�'@x�htA�mƪd�.��L,��C�'���:��"s����ˇ�{��p
�'���c��T%k]�h""��ct�1r
�'��}+ת �0��z"!ڶSL�]���� ���l���r���׾���#�"OR�M��<��! U��c�^ [�"O|�� ڭtt�U���P�I�"OI��"�+�fe�IOk���T"O\����/�:�[�K�0���;�"O��b�Z�r/�aQR���v�:�"O�����o`iJ��{���"O�%�/��o�fySA�`�H�C�"O�;łЗ�D�K���m�4=q�"Ov��qΏ�A�v�9�χ��l��w"O2Q�v/CX�deY��/�tE+�"O�)ɠ�[�C��M�����K�N��"Om��]��qI�JW�q��M�W"O�}8�m��?0 ,z���&a�S�'��Ðj��m�\À�1)Tڱ��'��䡒Ν�UΠB�N:%Ӫ���'��ЅR@����h��*�'�l˵Bι0��i��A����'��Xc��̏9j�Z�JU�
�Ё�'�d�dDX@x��w��q�F.D���)�9@�S�I0���b�(D������W�@�Ӷ���0bX����$D�`��@:�r���/E��ذ��%D��h��Ѷ?5>�(D'��3��X��� D��ъ�;m�tr#� x����2D�����M�"�J��^�r�����:D�t�Ed�mI`���P)M����!�4D��㤆�D.()��M*��03b�.D�T�.��/Gr�Y`� B��4R2")D����B��b�ʣ4v-�Bk&D�\��H*f4N�9!ɆZ�T�u�"D���-��e*L谢l0c���@h#D� �g�ئ@��*�A���3�&D�Ը1�$@Ĺ��Q����$D�칶dʴ`Ԏ�p�C�5!w�K�b"D���f��`����N�Lĺ����+D� �d�_?,l�d(	&n0�&�%D���U	��x��(H6D]�B�2���#D��H�!��n0DA5(�$j2���,D��iS#SƠ	��O�������>D���P�څ��	�b�ƷG��8�%.1D���ǭ̋@L�̀pj �0D�t�qn��f ����U����.D����عA�����S6Ps`�/D��	7j�����c�@�P>M��*D�Ȱ��gg�(�ġЏ7J�`e�4D�d�@�X:j���в��<2N��r�3D�|�A�����	�*�1V�b�h�C2D�,�f�F6'
H�t@C�Gk"D�H��G�:�^-*VG�,#���!D�\�0��~Wf�ȥŨs�m`�� D����Ạ,)����^�PMr����#D��� �# ��PQhܭm�00E�>D���'F��Y�N��N�%Uu�@A��?D�u$�v���xÆ1������>D�H���un��S(�) \D(�'D��� ɴVU�eá���3iZ��)'D��i1�N�<	��*���QT����#D�(���F���3��ҡ���h!D�H� ��\��X��Υm$���:D���r��o`�`�̩>�&X{u*O�dS�
-1)91�ȟPV� 2"OR���'�7 ��1f�=��܀�"O��3#�1�4�h�O�{��{�"O� �1w�\�"K���-V�~�T��"On�����	MG,X�C�/W4�ҁ"O@|���SEXd�E�!rN�q��"O>\:U P�Y��H2����S��2�"OFX:��3�F�7.�lh��"O��S�/ޑa\Č��#��'�����"O��ċ
8[��yAbZ.|�h3�"O��XT���8ՋU
����H�"ONЧD�'r�f�U�r�K�"Ou���
�T1p�D�����"Ob���.��T�ht�U�6��\�"OlL�U.K}�ԙ;�JI�)��=��"O<l@�A� 7;f�(�T�N���"OfQy��:?�0)as��+"��a��"O:�@/�o�@̚-F�X����"OlkT�V�~Y9��4>s�<"G"O��:�G �W�BԠ5�˱`^4��"Oi���=QmX��_3Pް�"OfܺSJHd~��h@�7M�U�0"O�)ZQI&\ή���>xޖA��"O��'���W\�RoӼ�J�s�"OR�AF G� �����lŘE��ܚ�"O0�<"X�v��9[��9��"O!8E�2-r�4 �H!���	�"OL�$ZM� ��/F����X�"ODMZ4���"(���N�e��	��"O:U)�"B�b�� n׋����"OM"��-si����v�"O*4����a.�(��� �T"O��Zv��'oǸ� ��4+�F�2�"O�S� �%�L:Eg�"Cx�eɔ"O|[�T!q<dI@CM;aqi�c"O.�U��3��t8G�K+M z@XA"Ox}� ˏ7k��]�2ʬ���""O> R�fp�����G�b��T"O>p�F��)�L��E�
=�pg"OT��ba�r�l��ƺn+vH0�"Om��D>B ���dԪ^RѣD"O�<�,ވ.c��9�Y�i����"O؅q��¸y��� BN�D���"O:����"�\4p�I�i��t�*O*L9d#V�Z��pd�E�K�J�'��i$�� r�@S�ϋ:��(	�'o�@����<z�
�}֎�(�'/.@�a#�<{ia�N�$'.r	�'<.�
�	9��4ң��)~�bm�ȓ<���S�ѓB���cqEW%k&ԅȓn�^���JB�0o&P�L6o�����
M�dY@ďwZ�k���;?�͇�n�ᲁ�R2��f�8xY��U0�j�.��R�,$kP��2B@Z��ȓ��0�#Zn8�����ؖ?NҴ��L�8�k&���$���Y:�Z���t���B]���+D�N�R<��"���3�	9N ��
c�R�rԄȓ[Τ�W��XN���'�:����_LPz���!D�� jWh
&|̆����0h��%m*%�1�]���ȓ%�������11�  R ANli��ń�V�:��{�T�8��<��r�l�����k�y�P'�*���oO�0ڥ)|j��*G�_=(؅�bФ�r�E3t�`d`�eBD�����d%�sh\��aP��K�?m���S�? Z�ȑ釛8J8xD���^��4K�"O
 QU9/�D��b��2[��%��"O�m��,�DhB��  �Z8:c"OR�9�a5.T�s����8�{�"O�ȩ%d�6U�pܱ
�������	ߟ��GJZ�j����'��T_?���A�)Vȉ��P t*)��M
,���?����4$��G�?7�V�{94���|b��M���@Ji|���l�'����!?gr	R��w>e�G�X-fTL+�D�w�����L/b��u(�&/ғ6{���I�M�7��4�i�pǙ�iS2@�Ca�?m=*m�p!;!w��֝P��?�ײ��#R�k�P�+-��ݙ�2�OJmn�$�MKٴR/@p��lbA�脠X�4�rs
Z?q5�˄M/�6�'��V>Us�'��T��Ӧ��u��0b��K�AC1?U�C��IR�J��HK�}����_'f%^D`�I�?!�O��T���|	B�_2"�(u�"~�0��i�M���g�@�CWn�H���^$U!�k��t�dH'肕&\�]禓'���N��?��iS��S�c�ܴW�T(���	.*��4a��[uW���Of���S�,O\��m�5K�.��C����IŦ=��4�?ٲ�i_�غ3��Yd������?,�`���1s��'�P4	0f8J�2�'���'#���xmZ;^b�a1��8#:����̙4A�]� �"~��ㅳM4H�bU��ja7`�̚m���*1�E�K�I�
�r���0^�� ��dg�����e��CG�Fb�t`rd6%����T�:����/�>9L^�����:���?1����D1�mi�/�b�HCq���3��$�O���$C+i�u��Ǥ2*uA��F�2,(ڴB4���'�6-�O���T�'O�\��%�#TV�C��"T�̸�↕PdJ�A��?Y��?	צ��?)��?CM>	��4K������r�Wb�^d�ղ���)z�1b�*�3t�uZ���Xx 
��� f�Y{`�7	�v�r���`��p@�)0Q�����	�v�(�ă0c\���գ�
�A 7a޸f>8Y�¥�����qy��'��O$�'jU���Р�}� ��5BM\����u��!�7�Y?5���H��Q�V����1݂��S�i��	6�豩^wr�'���i�:ɢb��!G�z�#&���ed(�D��,�?���?�&DK	pЊ��A�H1v�z
��1Y~���M:b0�߂M�z� �&ߥl1<"=ɳ�N�!��C��Ϯ}\�Pa	\6/p(гR�E�J��ACC1�1��ΗS�������O4n�>�MC����Ʌf��y0�#�\�uh�I٤ �\t�Iʟ%�"~�	<2%�ӆ�=q*�
t�R�4nz��dʦ�h۴�M��	�s��*."	��m?A.(�qY���?�.����E�O*���Z<��aB�5t�D3�N�<|��� ��'Ap��Zs�A�1��i�� 8����uן�˧��\c�>a5䂤M�Ĵ���^�!x�ܴ�Z��E���nJpQ�#Δ6��}`!lﱟk��(G��dG�/�h�o��V����?!��i��S�SM�ܴK�ܠ��cB8����Ն�T\�=�����D�M�Y]�D�7�[~��Y����(Odm���M���Զ�,�ԃT:]��x�*MnYhBg��T؞�S�   �   d   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4͒6R64<�b����!$My�+�D��`����M�'�i[B�p�\�'x���͓_�������<.p����_�/Բ|ǭR�K��у%�	�.�' %�F�ҞK�������,���#�� ��B)\5���I�X*��+�>��Uh� YO^˓y�� ��5ܤ1��l;Fr�Jj�s��lڲJ��`�}�V�{�.�>�?�fE����GX��҇C?qix��㆔�,�~��'����	(�X�a��b�t�'y��c��3��4�׫eÞb�I�,<B� ��Vt~r���>���C�
�?���'0�����
,?R� *Ot�9ӂV�"��\Sc�X�W}*�r E���'�|EEx"H�&��°�K4CR|���� ��#<�G+�u���a�B���< p8�O�""B��O�ሏ��_��'ق,�J&N� �P*_h*R9�4zU�"<�EO5���*S���a;
2�aԴr:���u�q�"<�'n"?�G�2K��=�e�+n���q��my�WR�' `�?�D�"C�	26%G�"Y&+J�#<�"�6�wS���U	,B W(�#@��3Ζ+�1OR��DO*��,}�����A=��i����m�	�8#<y'!!���F?adn�3<� A�DX�'�0������8L�@��9�'���?��6�"c ��c��T�W�^�r�;�	dP�(�r�>Y!�	,��Ek���C�B�ԉG[}�!�D�'_6�Dx� U�"�!v���S2XS�Q��y�� d  �Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   ~   Ĵ���	��Z�tIJ(ʜ�cd�<��k٥���qe�H�4͒6R64<y�b�l`�V. 'Oo�tۖ�h�B�h�#Ԙ26-�Ԧݘ�4B,�D�<�O\6-c�bb��&��RA��M:d�R�A�F�B�҇��)�qO��H<��"��"�v�2�4x j���><v�Z�+��[i���'���(���'�ȡ``J��]\0��'�����A�9��;W-�1r0�ӒI��_��
�4y��5s�'�4�v.\�<���|"�MZ������z�b�Y.8$4]�P�άyq��-w�x�i	�L���:^�DH���;��q�af�!9�V
%aְ���#ď%&��ImE�1	��l,҃�O�ye���[׶�q�S����,�(zb�K�(W�G1��Q�BXp�/��R�qOҹ*���[�@�|���A?X�^�"���+�,Dx��Bf�'�P��'�D�e�ȉ*yZ5��%;�
q�N�Hi��!)�qO`��
�
o��y f��6�q�2�i-^=Fxr�T�'��I���ط5��a���hk��_�'��c�����$ ��?!��p��	Ŭ.F�q_�,�`˓k�D#<!s�)�	���4�A�V"P<�kV 8"F-Iq�	�%��t�B�'[�-�u��(i�4i��l�J��yR�Rb�'j�%�,��kP$��Ġs�Z4[n����@��s��i+q�'����7O�"	��I0�d��wf�>DJ0��MyR"^�[��%� �|r�@?�-A�O׾�a�#Z�`E,%K�Z[�O�|���%�(Or\�N�(�.�K�Tܓ��!O+.��d�>��!�4�#<��
�T��qC�Ap8��c_|�<qR�� 2  ��D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"    %    %  n  �!  �'  �)   Ĵ���	����Zv)C�'ll\�0R�P��I� TF�؁���TR�	�8�RB�ɖ�>���چ?��aC�]'^H�I�!nB�Ύ)h�;0�E����~�&n��,�h�Q��X-J`�I�mE1nN�h�u��+U*��>�,�"a
,�^A:t�_�X�J�
cLP++�p�m�YC�uk�(��*�\ңbM	�:M��W!6L	o1?�rԁBT9u��'a�%r�=K��O��d�O���@��p��¡�~tb��E�-*��	i�i9�����|�
0�6�+�NErH ���*���$J!"]l��3�'���qs���P�՝E9�/OV�{��'�7�7ړ�~�I�9%����:�e��N��D��oڇZ
��� K�f@��b��=�n0���ď@�v)�>1��l~�O�^>suK�5_���r�7K�.�J#��;	���k�'�^�Ƞ8q��<#c�$V� Ԡ
�'� 1�D�E�Z���ԌT]L
�'��3�n"G<x�G"TP�'l���ɀ<,)[�;{�N��	�' ̈���i�v��P��z	��Y�'����*gl�=��'�l�(�'���EO7Fz��'�B�f��,��'MRu�Ԅ�! ��t�⫄{r��	�'҂�:#���6����`-�Z�
�'u����6i�l̉uꈘ!h�I
�'��1H�Nկj�(�X��/ �Թ��'N)w�σI<<�9ՠĠ<��#�'4�\�v/T�b�V�A,͈<����'�XЄ�S8�(�A'���a��@��'�L��t
��s�5�ViG/���{�'},���6iJ�[F��;'x:���'�H���q[�M�r���^����' �8��Ұcu�ёUc�$TF�}�'���6O��[ʄku-��UP�4��'���	  "O� q�4G�R{:d{�'�E#g,C�\R��LL�|r�A*�'.�Q��C�kC����N(m���k
�'v�bF�p6
V-�^ޝZ	�'�j\�e-�,���1G�;����'���W%�x�T �b�:+�5��'-^ܲ�C9����F#7����'l< �0f
lA�cU�W(
�@�'6*�H&H�Wp�����"@�����'��l�@��/lH�p3#�z\t�[�'��)��@'$W2�Y�B�n�,���'o2�I�D�?�.0����h���	�'C,�ò�7g���1��3�h�y�'�$)q�����H�Fߤ2�.)R�'�ܺBԒ�� �X(,�N���'���V/ƽVSm.Ala��'`� �e�J�bB�? �H<��I>D�D
TJ�l2���a�P�=�,�D�7D�8& �A���Pk HU��@ 1D�<�գ�6*�4$���ܣr��	��<D���vf�� v���#Z�9x�P�O%D�Bb�J�d�P	�,j4)�D(%D�`��
�,��䯄�7�&]x� D���˜�"�,	uEB21�6m#D�D��d�j~�QA&�A<$� �I��!D�($I,'��	�!�� ��
�J!D��*��NSB�)��̨]���9f�.D�� r!�
 W���%��Rݼ-Дj,D�$�0�[�fHdOT>Z-�%�+D��R��?d&�|2��НTv���F�*D��'�M���`�qI��:A;!�*D���冈b|0劄k )�I2D�(D� ��h?�(�Ђ�,z�,�K�G)D���Nmh�9D��6V�M�R�j!�� 
��aD$[�V�Y�kU9v(I�T"O����]y< ��a�q��"OHhHD�
�*6&�AŔP�L��"OJ5r'NA��	D��R�DC!"O0 ـ�Z�.Pt�R��X�L[J8�"O`TZ!����ؤ�-H-tV82�"O>�Z�ǈ�$�H"��s����"O�(A6�C�nd��E.��14"O�8b��ΝN򆡲�+B��Ti�"Oz0qs�}�*��MQ_]h�"O�C��7l�Ȍ���=i1<8Sc"O(:��1�r(ऀ�j'2�"OV��7�Zl,��P'v��P6"O�a��OϒL���U��e�8Ya"Od�AE[\b�p!q��:{��1�"O̱ҕœ��	JaF��	��1QQ"O8���QiH����O]#Y��y�"ODPӁ%Z;xiD�'8��R "O>И��P'-�¸Pg��CUҽb�"ON��d�Y�Ms(yk��^�p��I(�"O­p��|K��Av DPa��"O$! V	\����va�-CV���"O�����O�6�Eˇ��@��"O�qC�T�`W `�0� K�z��6"O�̸�e\�Z{F�za�X����"O����#�2��\hĄ�-r|���!"O&�Q,J�3�H`�!P�4{��r�"O<�q�D�8Z�ltkA�%	;�1a"O$ q`�ӿ%��"&�L��C�"O�I8 ��;)X��E�+$k�j�"Ov0�`�.`��2P�SN��j�"O2$�P!!� � +נn��|��"O���_&d(Y�b)1{����r"O�J�NU(l[p��r��S/�p�"O��A�-��t� ��~(9B"OB ��іs�R�VU=� ]�5"O6Ҩ�n�|pJ�JޗL�&�f"O ����4���0ǢL/�*��@"OH�� �tW�p��H�Pm ��"O}I��ՏJp\�P�j0c�T�)R"O:���-�=[���)u�X)�f�+#"O���fa�8U3�YQ��P>U�f4��"O��P7E;"�J��/���"O��X�MP"d|f��Iǅ}�(��a"O���e�	4��D�V%N8A?0��"O�A�P W;D}Z�d����At"O�uP�k�*=4�7"Xر�"O�9f�Rv����@�=�e˕"OXr��+�f����6�
|*��DB�%\��Su��s��dJ|�c��O�}�!�D���ݘ#�/]�)���)Ct!�4��m�	�Q>˓5����)[�ci�i�s���.�|���T�hNG�&���hּz�v���O��Aat�k�b��0>��*�+Ԗ�8'(�o��]3�̇yx��:# �./a�\1�ė�<��� ���N��z9S�,�j�<9"F�^r�0W�c��u����m���GF4��f	߿�ĉ��C>�'g�^���<C�.��blLq~!�ȓ-���$��d�*��@��6�����A��xKB�'T�h���y�g�/g��8E
��B͆pS��x'C��'}���c�U�DTD��EǠE�"� �y�^TYELU��tX��'x�ti�-�`�F8���(��4Y�/i��1ʙ6�hD�p��|ں5ꑆ��K�Ω��+Lj0��5�c�<Y�˝�L����dN�*jqv�b%��~y2
�]+���1���ozV�p�+C	b�>Q���eضi�`�%v,�zN;D�� �t�N�ML�[�"�G�,���_�jad�����E)��s@��2L��O�1O�32��b���%��m�� U�'��16�/Dژ ���oA�l�Vj�#9��@���^i�L�ܖ)%az��N�R�p��֑`�*T0��Q6��O0�He�Ͳ���O�J�X0��j�p��s0
T/ ����mU3On�庆"OP�[/.�Pc�X2Y��@W��Gm�"IXe3"=z�AÃ�`�OU֌����*�Yѥٓz�yk
�'�%ǉ]d,��,�(�  �H0XP�A�R <O`���!��Ϙ'Odp�&����J�����'�drT$� ?��్ŉ$��G���f�"��cQ*^[X�ʴI�k��<rbEC�`��P�cJW�p!ęǓ�~����aB�1%��$�[�[����`z�1�C>D�P`F�zN�3��@!$zDRǇ'�I�j�����[t�>!�G�ào�6�1 �N0�$(D���S�#f$��쎎�<��JF:~Uj0`Bj<�$�l���~�4�5f�Mb��t��=p�!�DD�8<h����	eɠ]�U/��'m��0;�$)�O0t�&�@4��}�w�Q��ΐ���'p�1(��9��D���d��*�L�,	C���*�!�$۔M��$�^�m挜���4w��OV����+���p�Ć� ��a�g���x��)�"OpM�+�( ����!�D�, ��˴"O����Ԡi|y���ϮD̊mY�"O�P���'q����@<� �K�'�H���	��c��%�� ��%J�x�<�f�ӹm{�L�!�P;g_:��m�t�<�C�4.�j�2��O>��L�
T|�<1�C�3T�H�gʹ8����a�z�<�奀�72]�0�6��z�<Y�'��n��iL���8I��Mv�<y�䒉Gr �궦TU"�\�<�,M�l�2A����OI�9$�Fb�<�bh��h�C�0@��I�EVT�<1�+O�k4�-s�F��:F�M��Lo�<ႊ�-:�eeF9�PH���d�<�,^3(����e �E-x<�CAJ[�<���?x� 1Ǡ\�dn~}ӂ��Y�<�e'S�0L$ep��[,O��]�S��a�<��mƶz�x�#�¥-;
,#ě�<�d��0���3��)�(�v�Cx�<y��S3Q��4.� m�|m�Q�N`�<������	���m��Y�G�{�<�&�ϑK��u+�l�N���A�<�G���bq��Bc�i{���h�<��M�+�da�b��
3:yʗ�By�<��S���X��-G
_: J2�x�<Ʉπb�h���i����&w�<�'�>Ym����;f���U!
w�<��(ͼ\�0� �+�4|��r�h}�<�	�(g���"�і&���&�Nw�<��
'�TAkB̄>`���G�z�<Y�.Q�)������o<A�w�Kv�<��+�u�hj�a˯%j���Ee�L�<���	ZF�BKB0���c�<I����Xqt�xd��a�ٹ!g�<�����P	S��O86�̱A��$T�*���,�P܋_��l�qk5D�p�7��9,�Mj��[8�&��q�4D�d3+�	v��#f$#�����4D��GQ6�:`zuZ�j����7�'D��`p Z�P��8�K�u�Ha�$D� ��"��X�U{�kȢ(��l�w�#D��G��\ʌ��%cI5.F�d��B$D��E�k�4���V7Q��0�)$D�� �a
So��%3���%�YK�ppC"O��˾E_����*FB�"O����J
i��0�I�|��h��"O��	���s�X�Z!l�]Pn1�T"O�E���?:�F�1t�Vx	�B"O>����)~��i���6v�˅"O��Ώ9;}J�)˾r����v"Ovؘ�Ԍ#M:Q�G�v����"Or�����1@i��W,~gpA	Q"OҌ�,\�Oz�S.�%xH.���"O��k#��?{��קO�L	"O���B��@�FF�
D�Y�G"O���Fcu#+/��2��Y#��TN�<��������͕Y�T��fG؟�2'D	d���%S�m�0�C "���	�'v:�qb.��OSl����?28(	�'7�x3BJ��5�@m+ �]'fbqA�'��{�+*.k�%(�mL��Bx"
�'m8�3$@A��̀*L,D��'��𖇐�]w^$��쎢u2��'(U A�X
1�9)� 0w�TL��'_�P�Sc1g����0g]rP�	�'1(�cХLG����F�.bސ�`�'��L����G�u�4&j*�<��'r.��cH�b���A�-�#d�Tb
�'s4��'���^�C@J��#�',��3e�
^�}�5��^�I�
�'��ӗ�c�0���H�M��AQ
�'Eŉ�h��v���#$΃ zł�i	�'�Z�rg�#�u���I�m�:J	�'uT�s&N��αs !�qF�M��'�cGe�AY�)q�Sc��@b	�'wB��D�C7�"�R��F,ƃ�yb�I0��x��c� X�=��6�y�&ƞa�����HK����Pyң1^T1�u�� ��L��L�}�<��b��_R�h
6�Ħ�x��h�v�<)ƫŗ7�a��V�V<P\I��EJ�<��V	{?*��ŏge@��P�H�<)�B�=Pu0����7}LV�Xw�MB�<�ǫ"@n0�C�@�Q�� ��U�<�s$N�M�T�$��	ZXqR'��y�<��l�<bN�	[4�o�@��G�t�<1�њx��l"����I�R�P��Up�<��>7�X�TҶ"��� a�o�<y�f���a�Q*Y��"'�k�<Y@Z-��)�"Ȯ:���Λg�<yp�!B��ʦ	� B<Ri�U�d�<i�k�h��f�A�#'�]@i�^�<�u����Y�%�#	D��q�<I0�C"A!��5���\���Oj�<�)W�.т 3�Ŏ,l$���Ph�J�<iW���8*����Z�y[��aQ|�<1�R� �Z�S���4 �� �M�<Ib�1���yh5e�FldGCn�<�E����|0��
C�`���If�<Qtݜ"(D�A0L��3/�0Ұ!b�<���L��<���f	a�������U�<�S�K�!�p�o��5���n^W�<��o^��e��*X#rb�	ubTT�<	�G#_���H��� BW��S�<тoY�t�HY�1-�Cwt82�Z[�<)և^�	���q�W�8k�xH�O[�<�1�/^MT�D "���JS�FN�<� *< nQ���\��i�"O(���1\�����C��`(I"OtD�%��;�A�&WZ��Q�#"O�{��3xڦ��%�٨N&��I�"O���S&Y�܁ZbI�,�h*E"O��*J]N�^�iA!�5U �l(�"O���w�3�4�/�W���s"O$�s��va4]Ѳ�ĆT��a�"Ot܉Wh�=v!��s���$Ir `�"O�@���H�B�q��4 
� !�"O��u�L q���uI��AE"O0�!v'Ӌ�j�!�h��$Ȑ"O���Q�!�ʩ ��0�ب�"O�1�o�;K�����N�Ը�"O��C��AM8{bH^�	�"O�);�ЖEҌ ��D�]N֡	a"O�쩥� �|���ke�ƺq���"O�!��
�2���3�g��(@�G"O|� �^�`��F\ ���8�"O|eq��Y/B����̱�b�h"O��I���5O�! ��ƜEʌq�"O�ziJ#e��}P��ͣM�n=�`"O�0���ïi:��S�2��ك�"OB��@L9��-���#6���X�"O��iF���QH�ٷ엦|x�P��"O��#cC��r$n���[0	"O�9X���=`4��cJ0�a"O�u�F��p	\�#$.0:��H&"O �ɡn- ��$��ℌ0D��"O��ą�g-p�I�K���,��"O��k�&�_���V�
�1���p"Ox×IR�W�<��@��&�]J�"Opl�#��X��%jW �k���;�"O�a4a�_���V��.�tH�e"O�P��9�b�G-����_6�yr`�P�c�ō�0dT�ug�!�y"GV�]Y�YsMۼ(1&��dd�	�y��˜S֜$��C�r�UQ�B�y��XwS\�xR*[�^?�Ёw�[8�y
�a�vi"Ǆ�]Ѣx@�aK��yr,8^�n ��玢j�e��8�y"ă�'F''Z,\�ỶO�H�<1�"��wn4�AYs � ��f�<1��Al��8p*?��j4m�d�<�`��n��@+QC�<h�:`�a�<��	_�K�����Ύ/-�@I�a�<9�!Zy1 ��C���v�y�<9��:$S$Т&ZVMP��r�<90�:1�RDra��m+R(�VM�x�<���A9p6\��6���K� ]v�<!�F�;rL��Sao�
�8)��JG�<	Ce��]!�2�k� e����DbE�<aqᖿ%���3
�;/L&i01&~�<qq�[�>���YdHA�H�y2� R�<�%���67
��e+�0AVn��!�LK�<��%K0�taU��\ĩ�6�R}�<ɦL�$������X�JӶ]�b	�p�<� �N֞�h�/j���J'+�l�<@cQ�e���5$)��L:c��g�<9�LT��M�"�R�I�T�c�	f�<��ʈ�f|PW*��YW>��_�<�bVo��I�WF�y�(�+���Q�<�t.%<�4���=�d�W��y�<IL�߰u���b���y�<� ���$��"D��o����"O�K���_�@�P�C>b��a�U"O�Ѓ�n�5
BT�3a�W��q1!"O���0g�6����/͡B&���"OX-���G7y����M�4,��"O"�����5n�6�0v� ��"O.�"N�Y����&�\�1��"O:�K��C&J�Y���d
l�a"OQ�qnX�41��Q:<��"O�����'V�����̗[����D"O\̛"�G jl&���4]s�q16"OԨ��O��rb�����_�G"O�%h$*B�:�������V�F���'���B�wd@��F��O�u��FQ_!�	V�@�Q;,2l��u�H&V!�º=5�0��%T�xs0dЩG!򄎜$�l9)��ñd��D�&�;r!�D��jU6�(��ݺ{CVHj��η]�!��M33�5`Bl	=?D�6ʝ'6
!�3b�lc1��]"�{��G�( !�D@a��m"v(X�7��E�䁄�h�!�D�8)T
�V���K�jt�!��]ўPR��o�"��Fź�Py�H[A4���	=i+�x�bf���yb#����I@O��M�z�ӢE���y2��b�}��`��G��X�ٱ�y�	��U�%�Df��M617�'�y���?tz�	V�:+�M�F&X��y"��W�C&� ֢}#��y�Q��*���֥.����"���y�O�>-���^+0�L�¢�8�y�EJ�3�
�H7m	H�P�@݃�y���1F6���mW�|1��T��y��,|úLR���	S��K2 ��y�*�m�,cP��O��ȁ���ybf��]�(��B@�?ѬyRCQ��y��>T�ν�&1�`ͳ�N��y��Q���[�%A2)b��IƦ@�yr-G�cn���$C���F��y�J0-�L�vL�-2P�b���y��>4��2T��;����=�yb�͂;�n	Y�c
�5�θP�&� �yb43H(I�NF5�VxѶNQ$�yb���ĜшDc�Jw�|������y��"�T%�O�VD�"ѥH�yr�Ń_=�DI��8�%��*2����z�z�cFG͆;����lH���F��b�Q��f]��;�ze��" ��Soׅ	��z�G�:˜��ȓ	�YJ��h�	�dh�B�����	���"E�,8�� �la��� ����z�P[�o��U3�L��=̆��5�Z7c�TR@�6�̬�ȓSR\���V�/b��K�0�`̇�.&V��K��+�24�T��*6R\�ȓ �L-�'���F@E@�&�쉅ȓfg*9�2fZ�ic�ȡi�q0 1�ȓD�%p���E8���7j�.�-�ȓX*��$�~��+��� 7�x ��_.�2��!YN^���V�+���ȓ���5ɟ"2���@o����X��`�TqsD�F;a�<��OŸm!.m��dZ��1D��+������5,�.����=eȂ(� ܉��ԗFb=��S�? ����/�+����%�����"O��r�F��T�ֽ�q$X9���r"O��4�ї	(�#�I}����"O�2W�L!:Z�5���4G�N�q1"O,�a$Γ�=��)�� ��\�LY�"Of%��`|������
:���	"Ox+�HM**@���K59�\բ�"O �`A���a	8Dã�Q̄4CR"Ot�+��,yf��-����"O�@�����]{W`��4��"O�a�ċO��(C� F�LF&|��"O��C(� �R�˔ED,"&ͨ�"O��XMb;��Ǣٗ��'"O����S��w�͛&���K�"O)(�h��q�v�*�*�ނ�T�S !�d����ÍL1��ӭF!�K�("�Z`�W�tS�Q�g���>Z!�ѐyo�A;��
>.����.`�!�d�� �  �   w   Ĵ���	��Z�tIJ(ʜ�cd�<��k٥���qe�H�4͒6R64<9�bʄZa�V�OnaB��G�M��h}{4�B(+�6�UΦi۴U���<Y�Ov7mj��De�z��d��/�\a0A߸.w�Yc�.Cr��=
��8p4��c�d];0#���ӐI�0 �������#u�\�w��Tzb��8��-�]��(�ȑϕq[Ey� ��2�|�V��2�%ذ��y�V�{r��7�M�҇�y�*ǗpTm�V�OL瓭aݸ͂r�F.�d��\� ��ESe���8 h���O�q�NƉZ�xX˟�ڶ;��a��;+�,/Lb)�N��Y�r�0G	ɐ�?�&OX�%�x)�E-�O��	j��Ti_�]�rʓs���r�!�uU)�����0�#@�c䲠C�%4�	r��8��LS1{}x����'@H�dZ��OnM�����-�����8I�p��k��Zgz��r
����O����U6��':칱&��F�X#b5<�L	ڴH֚#<I)%b	ܤ0d�ߏ'��|*d�ǀr�D ����N�n��#<	��.?9ƉH�';8D��E�s�\́�E�Uy�f�h�'��0�?��j
Y�&���ة � ��S%�A��"<96(*�o����ȁ޾�3���e�^y�0��d1O�x ����ēml.%�h�X$J=O���"��0z��I4Fp�'���6)p�(cgAsk��r��_�D ��UMyb�	H?!њxB꩟�#��q[r�S��7(��,:�J�8
���=���#�\U��'��y�C�K�z ����9�݁�O��[��D�8�OdM�	�D����a������d"O�V�  �qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  z  �    �*  h6  B  �M  fY  �d  o  8w  T�  ��  �  R�  ��  �  )�  j�  ��  �  e�  ��  �  r�  ��  ?�  ��  ��  v�    � t P  �* �5 �C `N �V �\ c �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����O��=���Y�+�F���eIq���JK\�<1!( )�%p@�ř'#�ܙ�TW�'w|��I�E�J�����{�)"�/�F��B�IX��-Iӯ�7�ة5�Jba�u�	�'XJXw�
P��-��I[� �l��
��� ��{�*\">d 0� o9f�:�"O8����e����!(�"R �R"O
=�kZ�t�:f�C(kA@B2"O���1aT�l��yj'&�8l��u��"O�"3�	K�,@A�˽\u���%�'�剁IQ,h�A� 
��T@* �L���'!`5MV�+�z�i�ݕ.G�P"��HO���Q��cD������z-�"O�܂���u�0"
]�8�Z���	��0<��	XX���0��r;�}k�c�F�<	E/�����b��B���t��E�<��NʭZ� �被�������j�<�R�)����ɀr����F�e�<IcY�n��,��%�T$IUF�M�<QCK�@�������Ip��EB�<�e'��%�!A�*Q�)�THX�@�<Y�!]2yΈ��� �I/�P����p�<٤H�<��y��фk���Bn�<�1�D|L��a��=�m0�yB�E�`+X����I��A��y���':�kQ��h����y�+�F,|��Z�0�i���Z��yRE�!���h2ԋ+
����y"��;(?�h��c�!T��	i���yB�N4�M(���M��9�����M��'7��b)Ÿ4w\��!��=L`����'@9{�`4Lb�,`�թQ���'���(6�Ӿ�x�J!��:����'*=�� �g�H0�- <PMz�'y�0�q��.)(�� ,׃
��"�'n�؋��O�7G��\�*T����'>ys����?ڔp��o֜��C�)��<Y퉟:��|�go�)r)l����b�<!cn�/@���bd��u�*E`B��x�<!2悑D�\)��D�2�svMIu���p�{�cY>/QB��e��0"U𥣗�y򥟏=Ҧ` ��Ns�X���=��'+ўb>i��C��0���2���?� 	 �M7D����ǔ` <2A��c�� �V����xB�Zv�L$��,Ωw��TI2KK��y���c�:|�!K�>̨)�d0-M�=�'9P�	Ǆؑ0��H�Pm�;R��

ד��'��a)�A	>#�����9!�>D�
�'�����I�O��� 䌑�q ��'p��˲d̩��,�@f�Յ�;�yRK��|��� ��wI���V���y2���q�h���F�.#Z|XƬȻ�y���L�\�c.M�%�������yRdհg_�Tٗ"�>�IEfނ�y2��^r�9�%�/�0�0e`Å�ybOڪQ�n��T��"��Q�տ�y�gS�+�T�sdo�3_04Aլ��y� �?/l��nK� Jǝ2�ў"~Γ�j��q��	���[�
�)|R��ȓEA�y�h5T����Mȇd������?9g/�r_8��֎ط1�@PgDx�<�U�ъl��fS4+�8 d�r�<!�B>p� K�V� �z`��$F{���Ŕ<M\�0�	��j�d%��7�6C�	����b�)u-&�:��]5C��/}����LϪm'��9�Fߟ6 D����<Q��-se��#�_>v���z�<�N�	s��L8'U��hS��t�'#�?�hd/� d,��7\�xiSp�7D�� >}6�ͫP�D��#�շc�`��e=O��Dz��IG	�������������D�Q�!�$�]�X�k$">n�R(@'.�&F�Ї牑I�I�@̙ �`쏨V�C䉪&D$![a�!��E�	��B�	�N�@�0s�E�$$K�	��(�pB��Z�Vi*R���N���F��C�I�q[�0�*��Y�0�I=��B�ɷ)�b}�r*K��
�ę3�ZB��8Z���B���Y�&�Q2,6�_8��?a�@ăD�X�@'�!&^�vc�}؞� �Z��j�41��p���-VH=��<���ȓTZBmqB��*J�����i�&�m�/1�	[�Ok�̸��&Ze�πri�	�'~l���G�E]y`D�B'T�
�'R�}Q��8k1�X#��)3���	�'3ġaǦR��jY�ťܱ|���	�'2\q�Y�&S�$T�BvRt1	ϓ�O���#f;�6���F	{eܩ9�"O��x��Ž��,Jc�ךw}�!㗟|"�i�2��>}ȱ�U?Eɴ���Δ��@�1�Cz�<�gC� 8�`�_'/��I��u��u�p�$�>��O�X��̙ƌ�(1�q��2F�zC�^�C��R�z���!@ǐdJ˓�y��S�\T�d�����C�G�q�:C䉸:��br�ʄ0�l��G��dC�əZ�*!h����`�H7cǚd��B�	�>x֤b����R6� Aj��(��B�	!g��F�P�(��q�M�(��B�<6e��b�D<h�p,�y�B�	e�̉����<>�Xt���J�CƲB�I�Y�X�;��ݡc� �;e<]�B�ɈZ<��4�T�����$�B�	�Qiڹ�R�D6U8���_�K�ZC�ɐ_�Ȭ�JK�QT��wR -�"C�ɷ8e��X��F��Ԫ��"6C�Ie9he��Ԍ��ȉ���3lg2C�I�6��$��CT�P���:�%�7^`�B�ɶId�h� z��L�< ��B�I
T-� 
���d(fp(@��F��C�����
�/"�bV!.��C�	�	i����S���t��&��nz�C�	)��4��J� `��f��6B��.�����A*b���ʒ�n4�C�lR9
$�I�T�شk��B�	�+� � �BO25h�!�5N��Fk�B�I�jhy����8 �!�*Ћ�C�9S4�@��4&��p@�*W��B�ɑ�H�CA�u���+�d9�6B�ɹ!hآ�R�tȐ`��=s_>C�	�~���'*�=;*�P�`*T�-QJB䉠6]D�jt�9:,�T�k�?t�(B�	8Y=��Q�N}�,��lN_#�C��"�*Hs@�C�l#����L�4/�C�� X�@Y�cƇH��<�Gi-�C�I�<�Mp4!��F/�dA�f?\e!��� s.�IeD$-,��GŚ�@/!�ă�C�5@3l�})r�⣍:i'!��%	�4Xg@\*&$X�c\��!�DΛcT	�m��.���!@\�!��]e���ZP���J}rS���0z!��P��[���;w��P�Cτ:f`!��6�$)B��.�:�P��<w!�d7%6���bސ����v�Mb!�� BQ2Vk��48u#��5[����"O����(ð��4���Gߴ @"O�X��/ݷ���ÖHڤ6����"OAQ͆�a)��PDʜ�_Q.eS"O�Ժ�坎z	��;��k ���'r�'���'�b�'��'a2�' ,x��u \aZ��S�+GT8h��'q��'C2�'B�'b"�'���'�T��!�	�ȼRm	%xmF����'��'�r�'���'�2�'g�'�&�Z���=7Й��)�
	���/�?���?���?����?	��?a���?��E�)���Eo͕v.�����?	��?���?��?����?Y���?aAO�+P`�|8�LN�n��p�KR:�?I��?	���?a��?!���?���?y�$�3X��[��[dd�Q)`D�/�?A��?)���?���?Q���?���?�� ȣn�$s�[�S�t0��Y3�?���?	��?Y��?���?a��?��׏������[Z�*��D�L$�?����?���?9���?���?����?���C.8b��"t���b�S��?���?����?��?q��?���?Y�f�L�� ���)O�z��TL�3�?9���?)��?i��?���?���?I�e�N����ݰ\��	��%L)�?���?���?����?����?���?ač��d�4�j��@�^��,r!�E��?���?1���?����?������'�B�Q;`@ah� ��0�%�m��B�˓�?�.O1��	(�MӒ��5m-��*�.I�$-gAOuL�X�'��7M<�i>��@����/�v��,� V4ȡ1�����I״�o�b~R:���SD�)��[���f�G�E�TC���]�1O��ĸ<ɏ�)�$Eڐ!��J�
)��͈î:�%n�N?^c���Jt��yg ׂg�H�Ok��ږ��cF"�'���>�|�D�@%�M��'��ف4i&�bT[�&@G-��'�����Pa�i>�	/��l��冲s���ȕ*_�O�0�vy��|B�a�����_�>��#�㐈Tt��M�t~���Y�O���O^�Iz}bO}x�� �Ds�q�U�Q����O�A��*�#4l1��E���4l��d�i<�#W���h����fZ;���D�O?�I�(�&Q��!̫e�8�ףހ8���Ɏ�M��MXg~��o�t��%�Lx�Uɀ=%$�iRb�%u(Z����I؟̘�!�����'m�)]�?-31�<6K�D	W�2@%aH;a�ў�Ry2����X�*�������4������Ȧ](S�2�I~��f���$�H�sn��;& ���
�R����០���'�?i�^i.=+��F�( �AЗ.C�,!8�rnߧ-�j�'�U	��Is�B#T������	0%�9т�P�H�"�9%v.�d�<I)O,�O�lZ�f�͓U�iˤ"4��ʳ�C�2y�X͓J�V�4��$�OJ���O���Y;�
�#	 �(�3GB�J 6�f�ts�ğ!6�O����8(��H��s⍍EB�Y�#f?��)��<q���d�<E�4j�6g�����'�6g6Q���\��'H 7�~��	�MKJ>�0 \�<��1���.��j3�� �yB_���	̟���3��m��<i���?��Ѱ.�J\�`AV�Wnn��2�o�����hO�ɵ<��hD8Z��	̽k!b�
"j�����5q�&
���'E哜T�l�N�5e&ֽ#sM��2��m�������	�<9O|z�A��x�t��X\}ٱ�$G�.����#!Ƭ���s~2�'B@����g:�'M�<��ؼ-r�r�%�X5&4�5�'���']��Oe���M��$�2� !=��\ʁ��2$�=�(O��nN�9��I��M#ɝ*����)�� �Q����mZɟd��#�a��?a0O\�G��1�1(b~Ϙ!Qhlp�V�%%��Ώ�yBU�����$��ڟx�Iϟ@�O6�����]�Jl�a�(U*,� `���ʦk�O��D�O>����DΦ��3���ӂ�A�<|;`�Ө;`
��4h_��0O�Ş5���ٴ�y"0a��Y{�H!n���Zc虅�y�/��E� P���ݠ5��'��i>����F �$%�%x�bI)�V�DS�I�	�����ğH�'.7�F�|� ��O��$Ux�(4#���1��yH�i�$#P���O()o��M�'�ɝ��J�
�"t��)9e�G�3�
�����B'b�P�$@:«"?1��8�٩\w����v��	X�K��~�*rf��Y
���O����O���|*1@�N���'��EL�Zy��e��&)�hX �'�"6-�T�(�
z���4�������ej@r2��FX���?OXHl��M��'P�-�ߴ�yR�'f�<A� Ly(�I����Jq�9ᤍD��De�a�pN�'��i>��	����	��4�	��lpbQ�s����߼X]�'��7M[�q���D�O��<�9OVj�x�D�(v��!�v��>j�NU�'�R7-MЦ���ħ����$#hX��(a�J����߮�
$;s�9qQ���'dEj��'A��n�p��Vy2C]T~0�$O�@���D�@
��'r��'��O1�I��MkA��?9��������8��2��33�����&�'Q�'���?��4�?!FA
4r�^<�E�6�2X�IS4��۴�y2�TK�29H���Z�:���_wo�]�q�? D�S��@+b��r�M��g0j�;b3O��O��$�O8�D�O��?����K�̄iA��-PRP�92L̟\�Iڟt��4q�m�)O�lf�	�������U�u`�!N������mٴ�?9�gE	�MC�'$FY��ě-�=j���t�"���ϙx$x�G!ۧ4.|aJg�xR/�<�'�?1��?�ģM,R~��c@Y7U��!i�4�?����A⦱S ��8��蟀�O7���c
���t�u���m�n؀�O\��'3~6�����̓��'�*�ʋ)���z�N�tq��K�j���82��q�t��'���'�h���Tz�K>���G�\8U=&eX�j
{=����ܟ���ǟ��)�SWy qӨ��n��DWD�J�]3#��Rt�C�|���t���\s}s�,yID�ӭ�Ha���&=`��4$�զ���1�|lZ�<���J�}�3��H�(��'-�)X!i$q�h��J�)WI��'��	럠�I؟����L��F��Q�&��mٖĆ>a����6)�,7MX0:ږ�D�O���;�9Oȩoz�M���5�p�@d�5�V�ː ɬ�M���i��>ͧ���XL����4�y�
�*��5�` 
�R�= Y�<��e�2`�!�U�+�N�M>�)O�I�O�E3�Kb�89S׈��a�����O��d�O`�d�<Q"�i��c$�'4��'��d���œsvJ����g=�Uɴ�$Fy��'#��2O��
]�	�M.v{^#`N�ϥ%w�x�	�=����q`��V$R���d�­�u���O�պ��˼$=
�Ci�訃'�O&���O����O*�}��
ܜ*�%N�s�-e$ѫ{D����fD�v)�)e��	��M[��w@�)&�>N���UH�;MnԘ��'�X7�������Gq@nZ�<���FJ�x���V��Sq%�C�6��C&75�m�#D��䓷�4�����Oz���O��ēz`���B�!:c����52Д�z����7(��	ϟ@�3��$K�dɥ��j&�]"` �7��I&�M�'�i���3ҧQcF� �G��tG2��`�4�a*A�E7z���'8hH�t��ʟ���|bP� �R%�1Frh�(E�b"F=;�+Xğ���ş������]y��{Ӕy�l�OX�Ǆ��!�|`$ӕg�f�ْ�OB7'�	���O�6m�O������Q:$���E�.Վh���\��7M5?y�M'?h,�	0���56�۫w_��U��&
`ޡ�D�֊�y��'j��'��'��	κ��e����<#�HZ`��/2"��D�Ov��E⦗�#�	|�po�J�I=4� I3�
M�#�CV��$�ϓ����٦���|"4�8�M��O����E+�\���x��"@*M������x�O��|���?���i���pd�K�h����
�F�����?�.OF�o�/0�Zd�I��`��b�d�'\�A#	B34k���2�����O}2�r��o��<��d#A `�9�L�
~�"��d>r!d
\:/?�]+�O�)P8�?�WH!�dB9`Y*is �ya��s�4r�����O����O���ɶ<��i��5��ゾcG���ra� yD�8E��i=�	٦��?ٰT��ߴ^�"�J3�]<ob��5�
D,����i)�'�y��8O����(����'?���C�B�c6�R�.�\a�f ^�"��zy��'�"�'���'�i>Ї��4�(����^����D�T��M{�ɋ��?y���?)H~j�'���wG|yK�ʎ���A��� Ö4*t�w��m�<)�O1�b,� g�*�Ʌ@�D�C�M�B�(� G@4��I>��|!��''4D'�x�����'L\��
X6\��FR�
��iR��'�r�'
"_�$�޴cV�|K��?���r���kA�E#�9v�݂P��!9��J�>鰻iKB6x�@�'4�Z��2C�aB���"A�����O�4Ò�M�:������	9�?���O�$CD��pT���p�� ��#��O8���Of���Of�}���#��Z�5:�xH���w��4Y��F�܆j�����?�;i���~^�AP��V!VXHΓ?���Kk�Z�Ā��Z6M2?)���GV��� '�b��]C��G�X805^l{J>/O�I�O���Od���O�	�aTuT�t��@�i���`ζ<�b�i2�pZ�V���	]�'=uT�q£Ĥ:�jt��e��+�����U����4}\�5O�"}�F���D��U�>���D⚯b���ñ-�}~�ą_��=���{��'��	�>i��8R�N2D|x���/S���Q�	ɟt�����i>ŕ'��6��h�6�$ �(o�i� ���p��6$���f�⟄�(O��{�[o��L$���+ ��)*��A&
Hhź�1(��H�Z%����>1Yc�>�{�g����dׁ���!�'~��'Q��'���'��H3D8���ذdC{��s�g�OD���Or8m��lm�d�'�V�|���( 	�u�[��f���I�'����c�4�?��l��M��'�r�7(9���4�:pD�D�0x� ß�Q�|�P��ş���֟P����X�*L���	<fw4�V�͟\�	]y2By��x��O����O�')��Yp.G�s�0����y����'�*��?ܴ�yb����Oަ5��� 0=�!�ei�B�T#E��ԉR1�؁�O��i��?A$�2�dƀ>NT�u�C�\g�c��;I���d�O��d�O���<週i�$GH��7�̰�A���<�*����*p��������^�	:��D�֦}P@Mڱa5���C�X��(��(�M���{C`���4�y��'Ɇ�{�(��?�c�O� ީB�G�66��:A`ċQ|���66O<��?���?Q���?����i�+Ό#5*�5z��`؛*R*lڍ~�D��	�0���?���~��y�չsۼ���c�;")��Q-0�X7m�֦�̓��4���)�O��h��i�T� �N98��3���d�C��8O�rퟌ�?���)�Ŀ<ͧ�?��L.#� ��ş�V2��@�R��?i���?���d��XkLПL�I矴����~�^��� ȴ[����A$j��z����MK�i��d�>!"�Kb8$b�)�i7�!�aÊH~B�S���5C2�F٘O��)��YE�%*#���r�R`NL!#(�QB�'���'���ן0X ��@��ȋ��?*x�p�`E�����4)�*���OH6M/�i���f�-��ղ��a�j,��`�Бش:����'��Ң��=��d�04��q��jD��:���,a����Gi+�37�:�$�<ͧ�?����?����?� ��7�~�;��
!��(�FNO��$�П0˰��<����O�`�L;s�.m�2)!����>�A�iS7��q�i>���?�
W�L�b���(Do�
_zPE)H+�k��$gb�IU��<
Q�'���$�8�'��s&oڋ$nIЀc�/n�"`� �'���'m2���DZ��ݴ]�Y ���Hu�P�P���Z���3��)��M[�R�<����Mk��R��*tʝ*�f��U����D��M��OF���.A������`����K:M��H�8���,A��$�O��d�O��D�O��;�S<C7z��A@�0E�\"E`�*��ɗ'7"�w�v�*�>�d��Ӧ�&��8D��Ti(ŀ�ʎ%��l�F���<Y�Ov%mڦ�M�'`��,B�4����!2�(ɺ�+�Op��(ãК&PH�Ycf��n/8��'��i>A�	����I C���Z�-��-=�e02�Z%~������h�'��7-ߦg��˓�?�,�B��A�`���QoٶAt�=�Ӕ��OB0l�MS�'ñ��5p@�q�ij @��_Z���e�[f��P������i>�I�'$�'��{�k�ab��i4��'~��������Iȟ��I�b>i�'��6�=kƆȡ�⏋Bx�@C�F�~��Ku,(?��4��'U�����Q�ExJe �<-Av�b��8M7��Ϧu����A��?Y�ժd��	���D�m����G��^Y,xBp��N��d�<���?y���?����?�-�T��p�§�F�!�C�`B�dQ"�@ݦ!��韸�	ޟ�$?��	�M�;+�$k��4�,Ԑ�)�#0�Ʋi�:6--�4�����O��F�u�|�	([�N$)��9)������{ْ�ɐ"Z�Q�"�'Y�t&�@���D�'t>q��C�h5�Qb�;=���ҁ�'l��'��]��ڴ<��	����?!�� �p8��˙o(9�!��b�l-A���>�@�i6f���' ܙ �J��lա�� 9H�yÞ'�b�V�:c|�H�n�=��������oHB�$F�3�$�!��_]ȈWD�:W��$�O ���O��D!�缛��]�6d��[��'`X��"ʸ�?	�is$��$��m�P�ӼS ��"	{�E�'�:)6�T��<��i�.7�O�����u�6���papE�))��tc�j��"��/hq���U�_��'�`���$�';��'f��'Ӭԁ�'Oa��H5���K�l �^�Ęߴy��Y:��?�����<���h���%U�~xΙ��e��\��	��M�Էi��:�)��N��N�qKr	�򁕓u�d��;%X���e샠?����w����'W�&� �'�p�ڒd(eܤ(�g`��N	��J��'*r�'^"��DQ��A�41��!���KJ��SS�� ]M���+��&N q��M��b��>�W�i-�6-�O��[R��x�� 1D�t$��'�\�	��i_��O�A@�$W��r���ӣ�5��Ө>��	Vi;c�$�I
/�y��'�2�'���'�R�Ɍ��|�Eg̢i�h)�aJ�`!�ʓ�?��ihP�ɟސn�f�I�B)I��:�L<���WN�r}����O07=�j��dh�l�H��)Z���΂{!:]n�2�fB�]k��$�1����4�����O��$W�TkT�Q GD�i�Ɖ��;d���D�O�ʓp����95�2�'�r\>�8ï�2	rh;qW�
�1��*1?��P����4Dn���|ʟ��@B�K��y��C�@ΩP�A���~H#���s��i>%���'�T-&�8��Vx�n����8^�ppH&���	����՟b>ɖ'��6M� xW&l!u��h�v�����?�$��e�Ol�֦��?�QW�ȱߴUꂹ�fCA!-F.y��EK	
{5Z��i���ΰH�V��h���P�"����~:ƀ,B�:I"���8U�hH8�AN�<),OV���O����O��$�O@˧=���ƄZBB [�(���L���i�hm"rS� �	_�S�<I���#c�^) �ޭy�R�
A�$jC(%�$|��Ij}���bI2-l�3O�H���$|��UB�@�;��m�7>O�I���?��N>�Ļ<�'�?��K��>�A�D� .�~d��L��?q��?y��� ¦ik3' ß ���g �6np��v
]�Y��J�d�^�[���>�M�d�ir�>�,���Ȣ�!Q�uP%z�.Ec~�!CB�hq�5@����O�jm�I��C�1-�|؃EV:JG$T*5��4Sab�'��'���s�-�����r	�%j+`t CH���"��Z����':�f�4�\�a�iA* j$x�=p���9W��d�ꦝ0۴p�mӏZ���0O���3�X��'	�� �BQ͎l��hZ�e��r���+&�D�<����?����?����?��E<g�.�S��s��B$,����9�pc�������%?�I	q�����+�7PVA���2;B�h.O��DkӞ��s�O��Ȑ��N�zI1�҆H�ظi�%ղ{_�<h�O��q�&*�?a��=��<i!+(?9���1-B@6L��?����?y���?�'��$�ͦM�Q��˟�0�oJ<�(� �B�6-8�c壟\m�J��4x�ן�m�ȟ�1��͑x��a��S'WV�A��UU�
�n�^~���W]J=��k�'=�k,JKPB�� l
��}{�O�
���O���O@���O��� �S�he�`�AL'u#�A�ӂS����	ןD�ɮ�M�"�Ԛ���x�|�OL�
�$�#s� �pq��h���t�0�'�6�Ȧ���N�~�l��<��W�-y�\Tܹ�ȏo��e���
��'��$�t�����'q��'�x���E1f5���2�$��-"�'2V����40D��i���?y�����\�(by�FB�_�Xbe@ J��	������4�y�iFU� �B�"����ĝ��vdAFŗa$b(:Q���ӧ1�B�Q�ZAȬ�r��!
(JԹGK�����P������)�SIy�u�ذ�������1C�ln� N������O8�m�W�E�	%�M��ٶ
��)��$(��3ŧS!"��'1�Ұ�i`��O<��AD����x���J3n�##�ȿ&?�y.i�0�'���'�'�"�'
��1I��A"7�E�]ghY�N�mJ�K�4@x�����?���g?�����2#Աux�!��@c�<�4�
/7·i�d�<%?�84��'iT�ɼ(a"�G�K<�ڝ�f�=R��Iz��|���'J&�%�x�����'^$!e�*gRHQwD�0x����'�2�'�U���ߴy�:�k���?1�;qB 
�.P6��E`�
�N����>	��i46Mv���'[���酮0��8#ӯ�y�ƨj�O6�qP �G�
�I��ID�?Q�K�Oh=�3�R<J¥��H7���rw��O���O"���O£}��o���� �O�?V�����VX����v(���:O7'�iށ���ݐ!��1W��d�(q�Jh���4����'��S��B'��dT2�4s�'_�x9���WU�]+��ӰKŚa�7��<ͧ�?����?���?i��ū[f����QuO.=�C-&��D���	���Qܟl����$?e��<0��$�Ѳu�0	7h�_b8Y��O�oz�޴�yR�S23K�T�AŢ$rz��h>��(f�T�o9t�*���@,�O4�RL>�(O��Q�;t����7jZ4�Zщ�O �D�OF�d�O�<i@�i�F!�4�'
����E_�c�.���2W�'՛���~}`nӬ�oß�����	A�����,A��Kݕy3@�o��<!��]��i���'?���r�z�Ε)�Q@�)�F6�B�J}����֟l����4�	۟|�
��V��
��#�x�Z�� ���O�oڮh����<��4��'��L��a@�d� !1d���&�F�A�'��	�Mkg����@��-1�����uJ���թ$��#Q�jؚs��\���#a�'�<&�������'y��'�X�j�$�B��ؠQ�H�U*\�(��'�\���4sU�"��?����	�"	,:���L
O)�@a�HZ)9��I��D�馡@�4�yB�)^��qJ��.��Y�v'��U�G_�t��q���6*��w�	�Zb�*�2HN�t[�&BD����|�	��)�Scy�cg�� w��+[^E[�'՜g������V�j��MˏRj�>�ŷiT!p�h�0	jd���(Dj���@Cq��䟇1�7#?�E��$1j�)0����Rgf\Y��Y�Z�Ԋc,U�ybV�`���h��̟X�	ӟ��OT<p1�*�Є��&�:0��+�b��q:���O����O����t����AWXp��OtP�r���0H5o��MÛ'��)��3�:m��<����9��Y"��َv�.�2�O�<�3I�%3X�����䓳�4�����m���`M	�3B�`;d���<j���O���O<ʓ}��6�	�!3��'9RJ�p��q&�Ӭd���fζg�R�|҆�>)��i�>7q�x�'A���ub	� q�x��-b �3�'w2%�8W�ꡊ�
�6��d럪�{�|���$�7B���7x����rbF_�B���O����O��:�'�?���پ2�� ���$�z!8�F9�?a�iZ �2��'���xӖ��ݴZ2H���DG@sTQZ燑� ���ɘ�Mk0�i����7wn�F��lZ�Q8!���į�>�Q_ux��R��'f����|B]��ϟt��柸�	����k�`�޼����S$��ᰍ�ey�y�xxY��O"�d�O����|Γm]Bz"ߋs-Z��ϝ�?"�&W�p�4�0O��:���O�rЎ�@��T�'&c��q�T�����l8Ƃ��BQh�Iiy���*m���|��ٲw�H�M2�'	��'��Of� �M��ˆ��?Q�	�<�V5��;� bC��W?Y�4��'u��5����n��\�U�V�@p(�0h�ޔ�G�],rj�4#G�r�.�	П��Eb�0����0?��p+k�X3��=hU(�h��''�,f\���O���O��$�O��=���s'�H@��2^uR`ƀ��H�`��˟�I��MdZ��dr�P�OF|���-�`���H�*�ͱ5�d�0�'������Bp�������g1� �py�O�-��f/"�{B�O�?�C@,���<ͧ�?9���?)KE≮Dc� v�M��͒)�?����?9�8�d����?Y���?1���4A�2�h�W`�>c->�C������$iy��'���On���JQ\Tx�$��)7���'�OϨ� %��D3��O���R
�?�2�&�C$V�J7�D��|0B��X5�����O��d�O��<���i� �����t�n(��Zi�&�0]�*��I��)�?�g]�P�4RX��Ʀ�$.��U*yP�a#��i�R!��G����pcSeR����~jÀB8CO�5�F�2���� �b�4j�%[`h�QC@�<"�Ȱa�I�hgʕ���8��`c�	J���a�X��py��nG����K��+�VE�Ў�e�ND�`kJ��h��S�� �h'M@���d1h�1<���o�`�g��<�BgO�5���`�6eQ��L�!b��A�b��t5N�Se��LH��L�!��a!e�'?�@*�/�"�� $0 >�xв�	�<��!���B;n�У�`�3��j-�>�r�s�'
:4��X�HS�q�	�FƜq��@�a]�)HD�NЦI��؟��	�?yJ<�'XuN�� 
�*�����Q�|�F���`��'��G�s�T��Q�E��AҰj��,�����V� �޴�?��?q%�_�I������'���͗s�zl��i!SV,ŉW*3O��IWy�����'���'�b���X�0��
!z�rjeE�.�7��O^�pWo�N�i>��I��\�'�X�02��`�VR�lÉP��@�x�b�D˶<�1O0��O���<"b��Q���%��,�t�ӱ�84]r�XR�x��')��'���ϟ��ɾ:qFX�#M��@��@�ֈƷ,&�eC"�&�I��,�	�'�L0aci>�9�G�Į�(����")�`�&�>1���?QI>9.Ob�afX���2�� ;
L	d�B�@�Rq٣c�>���?q����d���<P$>�b�ˉ��dR�KV� ���Єk[��M����?�,O�D�Of����	�7+�4r�I�dϐ�+��Z#9�lZȟ��Iry�������k�ּ[�(����T��!�G�%k�'��ɧ1�,#|��O�fbѫ#�4Q[F�3@�^(�۴���-�,n����i�O|��`~���3o.&��f��.b�ԡ
��A��Ms��?�A&
���4�@����'͎��:H>�����W�'�F���4U��s2�i��'e��O� O�I�j����"J�$�`��#�4ja��mZ�Q�����D;�9O��<;~6h����<O"�b�v��%Lh�N���O ��P0M�T%��S��2;���"�K�iµJ�=�6Q�']�I�T�c���I�L�	�4�>��4
Y1"{*�8�`N�C�����4�?��#�dd���D�'��P���+�	��*��T�"iڂ���M��Z����<���?��� ���X�	�7f/�� ������S�j�N�	����Id�'���'��!s��
]��1pP�C�1Rx�&>��'!��'��Y��Bg"��T�>�$8�����0k��ݲ��?i��䓦�Վ	�ɷ4{:����-o(v���t&���?���?9)OXE��N��of �NM�&�1aI���ٴ�?y������O���RvP��^��H�M�&AC���7H)D�9b�iG��'I�	�EDjL|����1C�`�8&'M�c��<�wʇe$�%���'�ȵ���)�?�J�ؠbf�Q"���S��I�Q j�`ʓlȘ"A�iQ��'�?I�'f��I�8df����ɑo��h����1�d6��<����L~ʟғ���m�	:�v�4�03�q��̝��M�`�����']B�'M�4M3�4��avFI�W����O�	_�U�����C��5?y/O������O�P�n�x�8D�!���<dT��N���}�Işp����-���D�'k��O�PYC)I�`YuӥƓ�2jp � D�j�6�,hכ�D�'0��ORM�M�L�gü>!��	`�i��M݀\��	�I���=Aƍ��Z�xG͛�/�z ���}bmT9o!
�O���Onʓ�?!����AH�8�A(ɺT��$`JJ��ݑ,O@�d�O��D0�	���a��~j��a���1.g�5�Eї*���P�5?���?i)O�����Q������$m��d��|ʒ�c��_ ;�6��O��d�O4⟨��=$�4@(� `�T��Fm��>���;�d�C?�As�R�H�Iӟ`�'��c��z���T�6퉰1F<a��+���typV���M���'��a̎��A)J<�i�Uq��(X�%���	���Ijy"�'F�t��Z>!�I՟�Ӯ	�b𪇂Ίqe�Aa��(2�"%�	�<������b��' p�1���c\8�3��X� ��'5�#�5�"�'��'P�$^�֝�~\>��F)QS��҄�|M�{�O*˓kl)GxJ|�����U�b�rAP�%Eb�P����!7͝ß��	�����?}���d�'#�s�	@"����JV�B�F�Y"w�"�x��]
I�1O>��	4 ��4�S�-��Hr%j׏3J��`ݴ�?����?���	��4�&���O\���s=��!�$I�&�2]�lu��y��Cd��f���O���5��0;ƬݠQ�θ`��� vTx�R�
��,O����O��D1�uR�����h�:�a����szJ�#�JM�!F�\~��'r�Q����f%VH� �D�F�t(;CC��3�E�py2�'e2�'��O�d
=V�!�����!J"�E.����Z�6����8�	yy��'�mi�ܟ� �ܢ�!��fKb�G��Йٵ�i���'�"���O���FH�6�Y��e^1_ںe���\�����O��d�<��qN�#.����N�(��[)�JL|��E� t&�n����?��*�<�F�h�I!�������5x^�sfF��27��O4˓�?q�D���)�O������9�-�jcBy��٢[#�A ��m��?Ydk�-?+Tp�<�Ouԙ����~J��"��)Lh�O*������O����O��	�<��L��Ҁ@�m��:GLk|���'���0o�ƥ�y���J���R�*ч�<�^�	Q듓�M���*�?I���?1��J,O���O>�X�l�<3kr�2�EZ�L��9�3B��r'�Jc�"|j���~)j�b�:q�
Di�bW>E�N��лi���'���U�i>1���\�g8� @��HD(2���(r܀Ȋq�D�>y�~5%>1�	՟��E����&Q��iU�_�B)��l�����sy��'���'�qO���uI�:R���@�ԭ`�W���&OU�%Z���?������O0�d�B��j����Zs'�.H<˓�?���?q��'�4�牖�7���R���W���	ʵNa����O,���ON��?��ž���ɂ
 ��ᇁ^���S+�;�M���?����'B�M^*ٹݴ`+�P`��2[��@���&@+ND�'9��'��ٟܰ��]���'`(��!�b����G��-�m�!�h���:��ߟ�bm�&WHOVM�1�R��Y�́�LRH�h1�iU�`��#T&��O��'b��b�zf,�h���T���G(�8�c���IJ�eJL:�~
 ���C�`��į�1$�F�b4�Ds}�'�v<��'uB�'���O��i݉z��b�����!�|u�d�>���#K�A�DTw�S�n�*d!�I
,�Q�T!E��mچR�0�����D�Iܟl�Ky�Oy�#K �N!�"�؋D�A�R�S�|6m��N"��f��S��:ՎX1WRx��h�R���v�׭�M����?���!��2-O��O��Ķ�0�f��f����=:����CҌ��'��q���-���O�$���D��'�:�A��"o2���lӺ���<8�ʓ�?����?��{�$ �M*x��eL�Y(�Q0�f�����S�"5������I�|�IEy�I6��ġe�ݴn��y����z$iC�-�d�O���*�D�O����W�H�YդƸq[`�R Fo*
��N�O��D�O��D�O��D�O6�D�S+�	nڭ9���y�DL*��ؒ��06�\�N<�����?�2B �=/|�JB��I�9#1�Q7Hƴu�i���'1R�'�剞_��1��P���.�6�i��0L2`�E��o�ޟ��'�R�'{�A�	�yr�'��$O>��yS��!d��I$�������'p�\�������)�O��� �PB��:��9��LJ n�T��jZg}��'S��'S:P��'��	5k��@���E��M[
��U�`�ۊLz�\n�cyMF�;(P6��O�d�Or�	�J}Zw[�$9Ue�~	��H��4�?���r�Z���?Q*O��>��@b��(q��WƐ��HE�u�i�*УE�ܦ�������I�?遫O����)�G��e������!��0;�i�b�`�'�"T�����p4�@"�$��ch�����7��ղiE��'r��[\6��Or�D�O��d�O��B�)�*9P�G�
kh�k��^�X*�F�'��	�29��)z��?��)ߚ�o�/x���QM�ĳi�r�/�6M�O��$�O����V�T�OH�'	?u��9�Q�Ǚ":(��[�P;�$j� �'���'.T���J�s��X�pa��]�Z�q�cʏ
��*�O���?a-O��$�O���Z)7�C��;T��M�w��5v`�5X�1O���O�����O����<������I;E��Tb�f��6z��$R�R�&X�0��by2�'���'\��!�'��ј���l��8�5*�-%���?8�I�_����IΟ��'l��+�D�~��D�T�Ϥ[z���	�-5t��E�iBZ���	� �I.b���̟����m��ar�*8z5>`<��n�����	Ey"�T;0�'�?I���)N  ?���R,[o�0M9���8���֟|����`���h�p%����
���*L!~�`V��V�f�nayR�%2��7M�O��OZ��x}Zw�t�%%Տf���a�Z�g�x%��4�?��l !� ��S0Oz��}�����0sT�BkN7��Q*�C����*rCN��M����?���g[���'�D���˰y�m�Ձ��B"s��D�ہ1O2�O��?u�� ,�֍Z�lX�WV���lȍpA���4�?����?�q��b��I\y��'��$@0�:�js�ȬoD����M�."��f�'l�	�r� �)2��?���0��$`��	i�����,͈�ã�i����Qش���d�O�˓�?�1=s!�o�=0��`��0�Ҵ�'K\$;�'���'���'@�Z�$zu�[�$�"qC�X�R�������S�O�ʓ�?�.O����O�����<���TJ)6Ͳ�"�ѵ;�}�s2O��d�Oh�D�O$�D�<)k����
q��2���:��"!CB(5��^�P��My��'gR�'��C���WȘ6d�N��w�(J�h4�i��'�"�'��i��с@^?���B�����I6n��E�����n��dZܴ�?Y.O���O�������O4�$��~�3wlT��`X�&�S��<x���O��$�<a�
�T���Οt�	�?E1� Z�h'��.���qE	V�&�-��T�������I,_����?%Ac`��uc�X�&��T�>�c��s��gġJñi���'b"�O�>�Ӻ�r���U��J�m��\�G!�������h{�(`�43���=�ӁCM����LW�k͚�k�J@���7�ϭx*�n埘���P�S;��ĵ<���)�n��V�U�����Ձ�O��?��I�{���۪n��Y�*�lq��ܴ�?���?��D#���jy2�'��E1A&�h��ȣJ�h��fA���V�'�剧L�)���?	��1A��!OE�6�c�'G�8���Ÿi0�G�/`4�Oj���OJ�Ok,����ː�T�e\� i�	���"�L���EyB�'���$�Ag �8�f�J�Vys�,R3p�*��i0��O��1�$�O���90j�:$�C
^"�ز�*$#�Bh+��6���O*���O<ʓx^&�K�=���qV�����.5��)�N�H}��'�_������ �	�"��r4��фdN�6��YB@�Γ\�
��'v��'nBX���܆�ħ/hH0��@#`�h	��R�3��a׶iq�|��'pbB�yr�>1f`C���K��H�̌�`ud�ئ�I��'�XM:0O<���O��iA8WM<�9$�O�T"�&D�0�:}%���	ȟ�X! ���%�p�'j��CmH0 T��f�=F=F�n�Py�0��7�Gl�t�'O�$�>?)�N�*xdT9ʴ�E9tv~�{gdTЦm��꟠�̇ϟ�&���}�g�8_r�Z� �2�r%H�C���W�K��MS��?1��*�x2�'�`���h�7_Flx�*
h����r�α �7O\�O�?����q@e[�oϲ�B��ڨ�F��۴�?I���?��N���O����|0�b\�\�%I�!P1(� dz�Z�O !�E�t�SƟ��I֟�w�G(R{�Ih��B4�ڵ3%γ�M�EJd]h��d�O8�Ok�W�C�h�ô�ث0gܠ���ܓHH�ɐ%�p�IDy�'wB�'�ɟr�ق�݆Y����<a�@�1g���ē�?�������O����OF�J�ə!9;8%�穁�4��2�&�l��<����?L~j�	˛(C�I�� �~�P'��?eF>�����-%�������Py�'���'��й��'BR���F�9�2�+���`Ѧ�qK�>����?�����/5d�%>	�QM_��.]�5KG�'�`���+�M#�����?)�^.�� �����~���͕!��x!ĕr2���iH��'��I�!b@�N|���B��Ϻhx�hAƁ�L�n��P�H�W�'���'<��K4�'�ɧ�)�7/��[�H	�|mlY�/�=SO��V����҇�M��T?=���?���ONh@Jɡv�v�`�K�H�u���i)��'�Jp��'�'�q��ِ�K~�U��n��� !����/W��7m�O��D�Oj��Iq��˟P���H4B�@ Q�S�B��˕�^��MS�l���'����R.V�;�%}�tRT�FHG
�m�ៀ��ß���H���?a��~rK #����܉t`$���#���MSL>A(��K��O��'�҈��L��8yTGA��M�c.).�7��O:���B�r�i>qGy��3���q����Tnl��sT����Y',�t�D�<a���?A����DZ-��e
�˙#_DJe�v��E�< ��f�IןE{r�O�A��I��J��k'�P-sBց)��i��'�r�'cB�'j員k��	NȌ�񶅏5��b� �f��M�޴����O�O����O�)�!�]����
@ �T��,�y����%��&��D�O��$�O4˓zv>����4��$x�M��Pf��� 2��)�7��O>�d4�ɠ~6�c?m�g�Ƅ[Y�4;1��'�hȚ7�p�<��O��d�O�@hA��O����O���L�`���Q����G@&���B`��П��������&�~�iaҕ(���Q���0�j�mZR~b&�^��v��~����"2��@���§�irA|q`��i�����O�i%�)���b:���+K�D~�B��ǯn�`���	z�6��O���O4�IPV����7G�4Q�\B�mD�C!����̘�M�q��_���F��Se��Qd-Y
J� �S.�l�� ����@H���<�ē�?����~���x레zf�	��T�h)ބ��'�j�+�y��'��'��y �G�.>�:C�":\���.q���ā uf�&����۟0'��� �R԰B&!p2�`�n�`��H�ܜ�<9��?�������n�٨5,�<D����J%�A�v�;���O���<���O���E����a�9r	,�K2F]�=J���D�O���Ob�(4�O���c�Mx��� �5�D��O����O �O����OT �U���r�F�Z����,ϕRC��SD�>����?!+O����6YQ��ӟ���j	��޸q%k�_�n���9�M������M��	��xL�~;����`�SM`�`�쑿�M����?	(OF�����ϟL��~춬�gl�9D���Z��U��� pL<�-O�����B���N�Aq ,ҐlX>+jpEc/H��ݕ'�x![�Az���O��O��8M\訧��3y��Cq�,uܐo�Kyrh��O���abУЕ'�bJ2B��2\��rP�iR�l�R�|����O�D��'�<����� .p���]3�%�f �gl^��ijBx����۟����Y*��z��% �1#$J��Mc��?��^�x,qלxR�'���O�)�i�p�\�#  �
�����$TK1O��D�O8��צ ���bl_{��H�f���"��n�ן,�������?Y����r��oQ����D	=>Զ��j�^}r���'r�'�]�Q��.=�qBd��n��y�)B4R��K<����?�J>�L� �a��X5�`@�=iIŬ+��ɟ����8�'y�iCE�k>��,�Z�
`ـ�'}�B��N�>A��?iO>I.OH0��R���W
߽5�p�2Q���5`�ɓg�>��?����S�'��&>���m�<z��r@�ހT\������M����䓾p<��)59>4�$��!2�n@J�`��]�Iӟ��'5���g&��O��)�A��d��:��Q�����'����IƺA�a�������1j7�<����64�&��~����Ԑ�̙��R�
��1�Î�s� ����`��B�	;:R��TO�x-�V���_�7��"M��Do�ʟ��I�����+���?���@<�z6�ך~���J2#_�_�a�'�x��!.��)�$���	l�8�p�l�$�Oz���N�&���	ߟd��)���ucR�d�Z�I!�V6H�Bh��؟T��۟0�1	���t�f˷>��3�gB�M���Thi��?�CT?��w�I��X\��F�D�`� �۽:)���O"��][g.�@"N�W�l�OBL�a��Tq�y�ᅩ	?l��'�~0jk67�28�'@���[��dI�g�uC�(�1{	��J!`ٵ<�Vd�6�ֱ\3l�jU��l}6m0p�T>� �kt@��@���h��p+[dUA��ݧpkܘ����X��q��[��-���Yc��q k_��Ja1"��,���WJ��d�ҽB�/�->��`��
�C���n�)Â� р��,����Dr3�̈�̈����ipoڞ
8="'�'���'�Qcf^8bLL���%?�|���WE���׋*C"�� ҿ%���T�A�'d�Y"�%b%�Ӧ��d�	P�B��-��Po��l��1R��; c��P'm�E�'�p]����?���d��>	�B��׉f���q&/���y��'��"�,�l�S��B�gD�;� �'� t#"l�0Ft���c�7����'�Xȑ3D�>�����\�D�P���O��$�0p���HƢ�,uwc��"NRIz�H�n���qn�G^� ��|����O�����b�nE�����m��T�D&A� �5"�>h �Y�𧈟�	 zl��1 �+������ ����'3"����F�O���Q!&u٪l��aѠ5�l�XR"O��Y�$�2Z��Y��Vp�i��I��HO�>y��c��q��%����8���I�����@ ���	۟���͟0�]w���'n��r����D�ѻ�B�MM����Oxu뇨��{��t���U'�������h=��E��'�R")׺H��4�I>o��� 1��8�������$UgP�%8a�X7E�v\PV�M�%���	C���'[ўt�'~ 
d��Z��#�߹���`�?D��b�⊽Gi
$�����(��]*����HO�DyB��~�X7M�6}b,�qK��k�F�C�O��D�OZ�d�Op�Hm�OT��y>�cW,Z����Pӻ:��be�� ��d"�LB�6��9� / xx�$[�k���$�ˁ��O2E0t���|\T�ck��X��M���]x�H�ck�O��$ƟzK<�&�#F|��4%�,{ �=��D�m� E0�	�c�\����@� �!��< ����+Ȍc��S�#��'��d�d}_���5Nɬ����Ot˧u1�p��<�>	�ucO�w�&}Y�#��?	���?��^bT���r��-4�􁡵�b��S�C���s#��5�Bp��T�+簢<!@H��u�dB a�/8���$�~���CPc8�Phɛ$z���UH�'�V���Fb���0���9@�O�#p����q`S'w��	Ɵ������qxPc�#tm␰�f�	AC���d[J�I|*��P�
R8 ߪ�P��`����1M�|��ڴ�?����)�1U���O��d!0�D%"���?reQe�D��1���;+
}c�9?�O�1�2�γfh݂�%R'�,�k� ױo�z�u&Z�;(b}뢙�"~�	�>�H�P��4N�*��(Xv���'���H۴}䛖�'�?�D�.*"�Q 6���NnB�����;���O���W1;؍�qM+)VljT�T�rn�l��V8cnr�$-x����HK�^��8Qr�Z=I��d�O�qqSY�����O(��O�<�O���X a��EJQ�,YNv@3&���d��#�z�+"I4��!���n�ذ��+,h�l�sd4.n���C�)��]�G+�
 #��r�?�=�tX&KS��y�Nگ>���Z��J��?�$�	��?!�iUV6ݟ�̟��'�2x���*B�����$��YX
�'��`xR$)����LL�	-|Lj�D3ғVe�IlyR����=� l`� ����iRƊ�8�@y��O����O����{�b���O��S�aF��Oz�r5ކ}T:��G*Ck���;5�'n�k)O�́�b�3AV)	)9f{��"T�'����?���@��kFǘ5N�	#�a����?1�������8ax�x�v��	GΘy)C�=(!�$Sw�"hp��E��07gNd���]y}2[�|ʰ/9��D�O�ʧ@A�4��,�18�;bHC?+d����U��?i���?���[=O����/Y8 Ro�#��0uD�Yv�ڕ,�>-�qM�zQ�����!�8e�ԏ,����B�?	ҡBO�7N� ;t(�DN�M1� ʓ0� h�I�M#��	�����K !ն*�^���KZ�$�OZ��$H� �� ����*��Ȃѫ�G�a|"�)�D݁N�x��M�z���L�'	��'��Q�'��\>	���Tݟ���,��nD2�0�A �1
(�W�ՆY���!2�5k��"�D�	�?�O81�2��, 4�e��i-
��+��LCq{���	�F|�1ǉ.E!����O�99����E�C +Ɏ4�aYr���$���,O�O ��U�� �%��/�z���Jns#�/D���b��^�)��ο{`~�s�g(�I��X���$������%t,TX ch��2F�4��.#Vm^,��˟��s�K�r �I�����ɟ�������A�\h�&@�~F�l:�!IL,�d
f�<��Iui4 S<�8�sK��E]L�	r�&Lq
�7VΘ�LX�6aҪK�!�
�z�S������?��S�'x�V��p�f��I�9�A�T;�Ҝ��g D��[�F�5x�(c��%'���3�B�HO��n~��}��f�ͫO�N����lw�!�A�S��'�r�'��U2��'��<�6���'�)H�r�:xPqk�wH�1cV��5�p>15
Thy��
J3����G18_t��+�#�p>)�����3�xU�`�Ȅ̰���[��C�0{�$ep ֔=���Y����4�pC�I./�F�PKA�,��h"ą�(\#��I���'φ57�f���D�O�˧tQ*��ddN�zY)� ��(x(�HM�
�?����?	�c�V�,�b
�8ոٱ2Ƃ��(th��a a߿swT��D�*0�<�R��1t�pP#Ö�D��׫����T$8h���)�F-0Z̄Ey�AL��?Y����ڨ0s��izh%��@�a&!�à6����ѵDwt����A6p�a|R:�dI�t��D��6\�\ ��۰T�1O���K�%��BT(��^T"s���>Q�!�䃃y������J�\��`�	��!�D�D���ؐ��$M�zP�Ԉ� o!���9����Ee�Tֈ��(��B!���:��pP�F��*���S!G!����0<�IU�ړ8�$[��6]!��0V��B���6�dE B��!�D�6 㺀qSʙ0/�ơ��G�!�Ą�4K��ӂMGu
�K$A_�2�!�dI�~h�J�ǝ� �r\1q�ݯL�!�D�W4:��`!�)(ơ���!��P2}fq�"�vhq��!�d��~Qб8�L�$�5�'M�T�!�H�N]�D��2�5��'5!�G��pqS�m5 ׎HB�	x!�dƊ7�����
Ia@�Y��li!�9r{ YB���(Q8��%D�Q�!���g���K/U�����K!�DԟwM�H�&�ՄIM�eBd���&�!�d�V���1@�Rx�bcX�{�!��^b �`��B�lXc��)Is!��QwDm`��&����"k� qb!�D's��ai�k؇P�F�yf�`!��{� b/E%{E�H;#h¥8q!�$�H�hYj��)�~q���me!�(p���f�ػ��`PAfB^U!�*D�pz!�>1L|�s�J<X^!���7���!F���r՘'/�[U!��OJ���kƄt�8�"��	Q<!�� ���DA�A���h���Ls"O�6�G�6bf�OF/5fx�'"O���C*#|ެ����U)@�I�"O�e�tWt*)�����lHsQ"O �ɴ
ӎjByX�n�!?�9�"O��b��3m�@�wn�"k�<#E�'�̵	ϙ-
���'R�Q�R	s����� \�l)h��
�'X���넏DĄږM�Y�d��O���%�^3|��0��Fś��X�N�H7�إIYv�ȓ�>ԓ�*�"]�i&E<uX0y��S������rZ�Q�'Ҵ�Q��c�
��\���d�>w�FII��X<a����N]�4 ��(a�̏}ˎ���o3�����
�?ٱ� �A ^|�0���4�
%)�4<�F�;J�n�J4�:O(H���P~_�PPq��<Ʌ�ޝ`�$*�_;zk�A7攜<Hh�
�HY�r�~���
!��<i��V&]q=��
�03���GW~��
O�v�Y`͟0n�Ɏ6h��ڷf�%_�85�r'�<&g�=�v`�&p[%$zӾ̄ƓeB���Q�׉dhjTP��"l���DL�qm�5�k��I����s��OD��
E!?y��@ܘ���
0�(����-v!���S�бC$.��f�\�Rv�����h�+d�BYk��]�\�DϺ&8���&��&l\�g~�Q��&)���د{2�H��N �0<i2A�fG~ܑEL�6r �B� ӧx�,��vK�AS��8P�_�C��Ê�PX2)Q�cu~4;
�[��!(�Wb-
��,B�"��'���X�LDzccD�R�R�%i�����L�v�P@�^�: 8��X#CD <�LݽfH��f��A��jA k��h�@ �PI0c���j/���)D�1
��	#Iz@��f�i�D ���nN�Y�rd� ����֧Ջm�!�d^�`���$1p��=�S<qDN���eԾQr�O�3p�<�A�ܼ^����,0=�< �#�d��I�mK�j�)}&� ��
�X�ax�eK�S�M�7�}��İ0�и`��E��*ܤ���׷p�"�U"�;L���'�T9O�|��'֒�e��%��x�G��3� Ȁ�Ov��2�>� ��J�4|�7l�<+���,h�H�
c}���G���j�;���*��䂅Y�>8��b��6@�e�D�Y�>Y��ⓓz��+wU�U���sӾ�d�@�a�U��Լ6T�C���dLY	�Y�F��Im�0��
�s��+ ��z~��S�q�┡UJ�S?�O�5�׎G]�a����A��=�B��,g� 7��x�Pt��D��{I�}����c`ax���d��	F��~$�]�=6^�+ ��X��tzF!V$u�x���딚F�j!��Y�'�bDPc�'�^�)$�7�i>9[�3��[�aZ�_c̔{4N+?��Ӕv7ֹk�`�6'k�U�fk��?� m����Ė$b���C�3B� 8p'@��zFl�Ȣ8,��>E�����E���C��J2�,�slT0YY@@�4^�����O��-�wdD+�y�eR+&�|��1�Cq�����8��d�?���ɷ	-�M��D�r�V�P���"�&���c'�+=�m�kJ�d�t���
�"/���ݤZ���oZ�Wv�(äL�&V�Q�vK�	����UX�0@��9�$��=v���i�i�COP�*��?R%Y����V�I3�ՎB��!8��'�+ea=�i>U��L�^��=��I�{m�4a��9�j���b1�u���f�8���M(.[��(���2C��V�հg���/p�є-N�>�j4 T@W)y ��;Y���w�V#�t䓖�o�p�)§"��D�� \�{�\�A��-+��	��CL�ÑM�?=.~�+%F
����'�\�jSB�4N��y�Hχ7�AsW��3����c��1��>�g��Y�}z�뛮=��� �!K�1
�T8�-<�yBi��f>�hR5ɍ�(����q� �HO h�0�F_�4�|�[9�����)ђI�1F�Dn�<!�͗US$8����?��T�����b�$W�%�"~n�Y��`��_��*RMU��B�I	A�LM�-Q''��T��JR���(	:8K�����p=1pk��^V^�{E]/<������xX���-S1�n6M��	�Lq�
�	����C���!��%<�P$~���8C#
(]đ�� ��I�>}��,D�x!�v�J�8�c�6D��!��3!:,xX"(N�	��TA���O�1��2�O���5	
xyb�
`9�X�6�c�̫ dJ+-�!�̈0Gh�	��noJ��$J!`y�I �~B[�h���O~qyW����I�C���;��4m�p�dΘ�0?1cD��?�'�	_�`a0�Y|( �#�	��r��'�8��G	�<A���O[h�#��v�X�b�af~	��i�h�+7�	�y
� (Y�@'��H{b���"/-d��ض���L�"����'�桳�g1F�X0q0��{�Xb�'�Va��x��4��Ƅ�R��q�韾*������;�8H�v��]��c�܍l�r��	�'E�ّ�d�lV8��˄gr�9�4{Ґ-a��i��r%͈�=e^5��G�a�y��gO���N`��g�s�(�iP�]$L9C�'���#t�'(@q���S4#y�lp쉟r]���od,eqo�EO��kS�.��)��|�6:�x���L���AeA!�^��Ҫ���OR�;�A!}R&[�V^�6��@c�탶d�8^�m�5J[;���J���<lC!�c��^���A�'�m*@A�*0BB��Z�d�ѝ'�ā �>٧��%��J�N��ū;sda�6�DA�Fe�T����}�&�W�VH<9@hN���1���#>�n�j�]����j���M�p���_��X���=J�r���J���5Y�\b�;E������`E��0?!S����?�'�D�B��X�#��	C��{:^h�� �!�Ψs�� GP@�O`-	�F�1��<�b@(g�Z�%,*��X�&f��D|�ON,He�"���i�0�Q� �#�x��blIe=>M"A� |p"�F*Ά�V�Ҷ��<i�J�l�bW�,�qqao�A��$˖�e�>0�M
ț���; H�b��,�v���%�b)�Э�Uh|�蜨L�B�
�'2��J���b��Fa\k"Ԕk�4鴰b��ic�pZ�
1�J�&+�4�"���Ne��Ƥ ���l_�t!���+�8,���'����$}˞�i4�X3�,d����G�1A0�؞Bۜ!%�S���a:D@ K��SV*,e���;�D�3TG���A�ԫ	��S��S�JL��s�☓9���x��'J�qR�y�@<!Sm�~V�25�8�����̍6�F��a�-W����Q�X�[�ay��U?l�&x��bA0B�n�I�mВ�?�bc���!����,���EߟX�Db@2F�~�	mѐn�HՃ6!N����!��=�D��E���B�9P�)�aE��|}����?a�7%��DÂk^L�t/]9w� `ÛGq$�f�I�����^HC�"�0#Q�ِ6��f�|d���'M&��&��+)X��T� >\@��/Ոv4te�T�	��-�CŻ
sB�*�KV�J}z��P�O�@��'Ũ��X\�B��
�Y�
}�1,ՎW�d,Ez"k"l.F��GЌ �b׋�ybbU�ܥ��U9k0�7	A0q�\�e�J��1�ۄ	�bX��P�*�*ᚑ�J6?�xM�O�pKĩ�Y)��c��'PT�R��'�:���K27�98�M��"Q.� ���`�ɞ&��h�	"��xO �S�LF�,^�z&�!�M��� =
����Z�TG4b 	�:&
,�'h��|
�D�#��1)�x`hfl�0(���P��"b��?����Q@^�/Z�����O9��9'��Fa*����^W<�Y���,iD�����_X��1E��S�	�@��Y9"j��6��� �@�#<!`�Jl�vL�2K�<"��h}�b
�>lԋW�"�ޥ�2�9+�!���G�|�pAj�\((���	˓��M�pM� �SF���Q]��XD'�NW$	R�O�%��(�m_n}�I��{��	c�N��*sb��m��kQ�4��$���ֹ;1_� <����HLC�h��l����=���e�b�`�E�;kI@��u`�">\�A�'��y�*�G3У��29P��&���`(�i��㊣>8``�K8/4����=�O�x�%'�Xg�Y��-�A`����  y��mrF_�%���X���L��!�3��G���[.O"=�@�3���nX�44�� �8**:0;�k��M&��U.�g�':�D��	�4�DU"��kM��'��7�|�d�BpI�+T��U�1+����|�+O@�R�ƮV
 �r	:]� |Rf�Ĕ7�>�I��R�&E� K�L}L�s��R� W�i1aC�I2����?O>���I��mХ��:���	W��%7De����/NP9C�G\�-�\�CU�Nbآ4 4lO���EH=/.`� S�fl�j&(��IQ��mڧ�~b�V�"
��,5��X:ua;Gb-��5v��[}J�i��P�6��IǶ�8��Dm�kJ�8����C<BK�A��F�u�ʨ#ԁ��@���a0��$�~�S����(O��iM�rjT" "� 1x,��߅���;`吒G�$���s�'��x�D̝O�$�1���e$��sӀ�m��%����Ê�F������O(X�~�YVQ��B�4;�pM��fX�9$v��0��*qU���W�gW��ҠL�]fX�S�;�xzrm�MJ�m�a�u���9��|�&K�0-d�!%J]�?ƈh!QJI�	I�U�r�L$����匉�����^-O���d�H�=zbd�7� ]�w�]�*)�Ȃ0���<1��~��E�j�L�:�d�S?0|��䬟��LՈ�bz(��"�L�;*`a1�'�j�S5�a�2T!���'�^��@�Z����o��d�� 9��J��d	`��	!~�KR��c0N��S�D���Pbg�� �!{6��i�$@�l����ח�OT���k�]���6
Y0f &���<��HM	EHP�+�ϹfW���g,�(}�ԕR������)�	�8N"��GI\+�@�i���[�X��\��BЯ(&�͋ �ψ����%��K���fjΜH0��*��'��,3�O�RQ��ʐ:\�<��J���`��O��Q�揍?C��
0S��M��V����G� ���#g�>w��)r��v�b?Ak��W�`��3��R�����*D��%@M�/��q١���HI��X��U�����?�$杴d���T��M>�w�@�� }��E�����#�\��$�+>�
�b��D��Q4��ai����`V�C�f��
�����<� TX)R�	�N=B!v�B#6>���I�g�:�
�l�K�I�T�^<U֊�7��N߈�B��V{d����f!�M�YD�A-6C�u���U!4�!�$Y�6��vnƅ+(t(`l4`w!�d̑�j�I�k�;%����&|!�$��Wa�A�VO�|Pa �Vq!�䊭a�U��(�-2h �V�P�bY!�$��� ���NT2���i[Fo!�D]'F��Q�YG��1؄8W!�$Iڬh�D��;T�xd��� %2�!�T�e��:�NL�@�L�A�R109!�$M�H�tMr�iÿF0�ѣ�տY8!�DćPOf�R,R�b|���.��$X!�@�it����4�^�Qg.k�!�d��de��Z�l�{��i:��:�!�HW�}b�-�T�����o�_�!�AJ�q����6i5+G��?W!��� �ni��/�,6���nK!��#+� 8�D�;l*tL�+ԣY.!�X�z%�I��/�@�|SD�T*�!�V�v��]�&m�"���|�!��8���@�${�(;�KQ�T�!�D_�7�4 #�a.Ĺ��.&�!��N�,�j0��ͩU�N�y`A͍^�!��ȱQj�"��"?,��k�x�!���B@�U/h�QB�GW"!�$B�}�TLB�eS�Y�BA�]�E�!�D��B:h�2���zH��mD	!�d@"Z|�9�2��|���,��!�P6~MV��(��/r�(sbl�s�!�J�vQ��ҀŁ�<YdMZ�@J"8!��H���)��'�� O� ��!�䇡O�	�`P�h/�)NQ$u�!���&N�8!�f�W�*'���4b�{�!�ͿIʜ<�� g	 ���U�" +�''<���A[���P���<��'�<,zd��[TT�;��Z�{�4u0�'�H�20�βZ��$sw�$!��Q��'h���cG ]��A`��b ̰��'��i�d��r�Y��Ȇ�,�x���'���"W��W�%qgǗ� |	��'��@�!�?��K�H�D`�4!
�'�X�����>�L�h7j^$R���	�'!*Il.jXV���,�mu��		�'��x#tIM�1+?8>�;�'�d��/�l���;�K@�1,p��'cx�!BE����Y��TX���'�~��f�*-�H�$��4Q8�I��'�~�Wᑈ~�ؽ�F�6L�K�'"ZŢ ��wFik�
�>�$�����!K��	f�+�@0Q7���<Y�O̭:W�u�L�EW� ��g�<��A�I���H���7rx��3iz�<i��N�$\|ŀ��R�Y��!���x�<���7x��ido�t�l��'�n�<�'���!���#�F���gMi�<�7*��@Ȃ�"]=�l�E�l�<AD�\�D�j�����6;��c�F�e�<I5�Ft���W�U|����K�<����B���
#��3�]'�o�<�P�"U-�s���)(8�����j�<ѱ'Q�tn&�aA�>sf�P"G�e�<	r�Xx�L|X�(��_��E�b��_�<١���v�5X�U�k�^�<� J\هDw ��#b��)���X�"O(��K=si�D�t,�^�T���"O�����J!c��g���ZE"Oح�g�/=@ �A�U�D|����"O�ب�R%f�2�gJ��r� �"OY�$�͝n�0�Ce��b��T)r"O@|Aa�/(J��H�-��0�(���"OV���Z�M_|��R+�g�>���"O.����ȕX���k�	J��<E{�"O��A�G���M��(��=��ړ"O��(�냄:�ЈHP��ʼ-�G"O�H�/���J�x�Oڈɲ�z�"O�� �AG�����2D�a��"O4��ᜧ@���f�;���"ON�0d�]|a��lB
	���"O���RNO2�2u�F���业"O��y4gȾB�Rd��}�A8�"Oʐs�M�a�6�"�Ci��� "O��Wɛ�M���CCX�`���"Ol�W-�"Y18(�@A+-��R�"ONMc���4"�,jc��cĨ���"O�*a���$����C��[↩;$"O|����a�@\94I?W~��S"O�\��F��2i��:#�fc"ea�"O�U�6AH*11e13�޵FX�,�C"O��e�"uߢ(���2r>^X�$"OH��GA�_�`��aW��n(� "OrM��.kk ڕ�Fb�|�j�"Ol<� g��i�H��@�U�Xta"O�eؗKX,��񐁁�N"�&�X����¯��ª�ha��QbB�Z�N�y�/��fB��{�G[�Y1�تe�@�y���vŚ� �.&Z�u"B ��>Y���y�ٌ_.����$m(�R� ��y2f��Q����!`
>$S�텨���hO����{%�5�@0W U�}~м��"O&(H�ㅑg�p���ȸ_j֬2�iR�"=E��4��uɅ�)T���	(ڐ�ȓ[V����1�t����Y�H�ȓJ�,L�t�]>�:Y	s�\&E_�y�ȓ[uz�rj$j�ɡ%`Z�(��A�ȓnӼ}R�˅�Ff�Ճ�{��|��f��ĺs�R�"`0S��-n� (���T�"��1H> ��V'm����	J<1���5QJ PR�J��,=��/�I�<d�K���	��TmZ�)Q�_�<�F�kאհ0mOd|ht�ǬE�<1p��#Iܡ c��V�"�� F�J�<9�K�M2�� ͘3
p��O�<y���$�c!��@؂�0GN�<ac�X6F��i�hQ�W���h��Q�<�QBԉc'�A�N�>�x����EN�<a�b�2�T�   D M�*�K�<�4GӒ@�"��<�2����JD�<i��`E�TrS(6Y�9�&Ɠ�dD{����2�H�P��E%X	�}Fl�<i,bB�E�^����4w�L3W�4T@B䉚3�&|SK��a.�)l�$gf��d;�2}=
9��dV�/��zŵ9wrC䉣��qv��9?|\��T#ˁUg�B�I�DV�sp	Q�g��{�C\h�B�	(`tN���偽Z9>�Ae�,GfB�	�	C�9*��	�?l��.S�@uBB�	(�z=2�-��y�ޤ�#�15�B�)� X�VL�$`hb�m�x�ɇ"O�q����fH�x�߾
�>)!�"O y�'�ؠv���b�۪J��L��"OT1��t&�P� ��O�HD�"O�!(w��*�M��ΪOj�L�"O,�#�L���ҨًlNv�0�"O�5K� ��-8���^� %"O��R��1Q�ps!/F�8`�8��"O�@S`�
� ����G��-I�m��"OX�xvD�Xf 0���V�0�ح	T"ON�K�fU�U$ht�*H�5�	"��'��$I54��7ɼ#�`aRc'ʯ_t!��P�N.�ء���x�^�0l��yX!򤖻�0��3\^6�`21�!x�!�d]��\ ��͛�_�|�ðI
v�!��
j(�K���aCG���P!����֡(�JD#�Vl��g�y�!��Z1��*���N�p9��%�� [!򤜬6:�Xr��Ž(�~�B���
q=!��WL���%&ڧ:��a"��V��Py��CP�`����Õhq��`��Y=�yrJR:*F��pAL�V�jprS���y��%$�A��k
�<�\ѓ�� �yB�\�9"E��%؛��P���y��ъ=h�����"���7�0�yB	�{�DX��+	u�RG��yҫ�	
��S��w���aq���y���t�"�@F��A-jY1F
�y q ��ECE�b��� ��M���	V���O^�|Cv�>3�:����ߺkL.�i�'z��֣��'�Υ���7_�0�
�'��!���&	�ԡ�@�Y>����'���d��l��j�L�<M�����'������F�y���<G����'���yW���/��"B��̸ ��'AY���-t(����V��$R�'3�ej���_�:��ČD�U:�K�'B I١�O�cJ���ҡ�W�`�"���8����NZ�>�6\``D̤��h1"O~]����w�˅��w��PQ�"O0�"�IÒ���:%��/��``"O$�*3��m�P����ȓj��u"O�Tp�Q�&l����,U�;���v"O�8�­�/c�X���AO�w��9�2"Of ��B��C�n��ӆ6�h��7"O$���f�ԤHunT+g�L�["OUTl�j���� M�q�v!�"Ohש�!F�� 6 ڑx�"O���sG��Y�`��D.v��#�"O���最$�|�ȦG�t����"OXf��0{o��1T��:�k�"O�a�g��%�6�pF�(Q8��"O^y�"C�&kC�\b4�ć��"W"Op����<!�"�u��M�@"OB�zuÑ3�8��゗	����"OL���@H-C�Zd�V^"�K#"O�)"Bf�>�(-��BP�*�a2�"O X����82��!��kg"O�X��@o/`yJ��5|g��A"Or�k�M��8�0�J$�q*�"Oh"��P�_Gd�AAK<]��1:3��8��	�es�U���7Ga@��*N?1�NB䉯ApU�v��e�z�ڣoN�7"0B�I�-���B�	)QlԺb��$nC�)� �\u /��}D��??��q;�"Otɤ��)S-
p��ѵ��Di�"OʔH㤛�U���!1�2���*OD=
c'YP��j�ʷ_q
�'z�a ۙv�I�c��[	��@	�'�y�ӪV��3�ν&�P�X�'��[��I<y8�j�hA=���'<t|��FN��$Er��)"��� �'��c��'�~����IC��T�<Y)�J�������4_�Tu����b�<)��Y%!FRp��ʔ�6���ɏf�<)�Є ~ ���(�ԁY�<ɕ� (X^v|R�'��[�8�!� ~�<!��.�XكO�v�6���x�<�0�
6��	���J�4�CAQp�<���� *�@ �1OK9i/�貧�v�<a#G�56�x�ȍ25�v�
�B�n�<FK�8.��)ub�3�����
LP�<�e������V/%'����j�b�<)���h�fWJS/�x�D
�]�<�T�U9A�
���M�N���+���b�<JK�#�ԙx�΄����8��UV�<�ʋ6����T�((�x��2@h�<!���mMp�J!�C�3� �$�l�<!b�ک7W�t���%"`T�5 �a�<A3�%g ٠1�
���R��a�<� ��,ۼ�1�K�!-��i���[�<YcS�=T�a	�-��Y��	p�<�4�E�;Y�Q� ���R���Aէ�u�<�`GZ�T�L4�R�4=�
�ea�s�<���	��ֽ�'���U\A�Yn�<��h�,��i��2m���l�<Q.�$<�y:AmD>��-ZP��e�<�I>N�NxC0+�(M�	z��y�<	�c٭�T4�qf�Y��L�ԣ@\�<���!x�� �GjXFEre@XY�<�DK�6��UB�ԓq���HY�<q���J|��%�H�4��Ĺ5��S�<y�%!M�y��Nӄ:�0d�C�Y�<qq�Ԕ(������?�xIQ�MW�<1SoP7-FV��aM?}����AG{�<Y��9$*R���=-����b@{�<��H���9 T���*�k�<	� j�M �O�o�=����_�<�e�R�D傸XЃ
ABb�K�"�T�<��F��C(Q���
=na�$K1.�R�<���=Xr�H�4}6`}�q�H�<�P�U��(ATL�0u�0#�Y�<Q2-U�cJ����-�.~)s4��Q�<��$'h��s%�<Ğ�Z5�^f�<q1fF�~E����Ś�J����GH]h�<T��!1�D�b��K�N���4��n�<	G ��>$gN��.�j׉�m�<1c��$e@�9Q'�	� ��s�<A'-�/�Z�#�_ƸZ҈�r�<����&U�1��E�>i�PHQI�<9��~v9c'�[78P�<��fLp�<�̚,�r��/ݵr��Y壃p�<av�Q�
����CK�W�R<J5��m�<Y �[�o����A)2�d�1ħ�f�<ᠤP��0��IȤ~�����e�a�<Y��\�J�"�� �*L٨�����[�<i`χ�O���sW�$\����1�CZ�<I"źi�ZԐ�gG�r�H�J�<� D����"�.�)R!	#B�`1P�"O̸����3���`���-eɚ�7"O0�
5"��00�⃩[�8�;E"O�5C�Ő�"�A�g:qW!3F"O(�2�c	>���`ԼL��h&"O"�
+�=!U�E�@"S� 2�D2"O�R`�V07
��ȅk (o"�x�"O>�в(��G�}0"離- R`0"O~l)"��e���8�WOZ䊑"ODU��e؟���"��NKJ�C"O^9ȰoD2W�f0;�BX�A]�9�7"O�f�Z�;ش���Х&Gܕh�"Ohd!)�=6�	��nqV�y��"O4(B�!�<^M���@S�"U�4K�"Ox���B�u���2�, �xP �r�"O�ks<��5H�F�P�5Y�"Op;VD�<:�8�`׀'A���"O����R�e	�<S�6J�}i�"Of�b�K�0h�ޙ�U�͙zG@L;""O:����J <���G6nG�2�"O8r�e�)	�8��CV:=Lqr7"O�,�SK�4Q�!�LR'W$�i��"O�4�ߟ?��@3@�[~\�"O�8x����Qi��I�	dظ��"O�e��_?&�B��!�J�V0�f"O���%2�2=( �� �
�d"O*1Y�S�}�h��aJ��(I�"O�X��NHT"X�F�$h���"O6��D��{О�)e�i.>Ԫ"Ol�S���]օʷC��u�H�4"O���#�H
j[�i�rȆ�Z�C"OH�s坵+c��EgM�	B�8�"O���,�@�>��Q�@9m<LH�3"OR�s��u��Jd�?��"E"OnDcs䝱{1�upG�+3h�K "Ol�jpn޲��@#�K�[>AZ2"O	��W�;�D)���R��QY""O�u�!fK�X{�(��@
�Q����q"Orؘ��X(3 �C����"O(�3���?T-��RIZ!w*Z�"O((oL;��0R�HH����QS"O ��D�@</H�Cg��`��}�"O��CEҜWj�)r��Y��d[%"O�ܨ1

#^\5����Wed{D"OZL��	Tn@�yWJF1J~q�U"OJ}�@ o�,;�)9q+<Dq�"O2�kYm�VA�.E�ܫG��d�!��D7 � i�#/���͉�-B!򄏡�l<�e^�n�� ̖	=!�%^*���%!�o�}Ѓ�ǀ�!���`<�p�ƪ��}�p��	�?7i!�D[9j�Lq��
3 ��1-�!�D���#t�3l�>Y)"��.<z!�źX����,�z�t؀ǟ�i !�J�g���Ü6ܢ����\��!�D���a\�1:ȁ�U��.�!�D�DZ�N/4#�<���҂/�!���+�>	�B&"g���rڮd�!�Ĝ%U���qr��>�I���δ^!�Ē�`��9���H�"�� �79!��BN��$�Ō�
s�괹��!��F)k�yA��-'
�8�'	�y�!�D� D(�UJ-;�r�Jd(�4-�!�՜I�0���P"씱8�˄|�!�� ��iA�ٙNCVp�FP5_|l�8�"O
��W��H����4#@�`�3"O�� ��� .ɾ�0��+]'Ya�"O��;ס���D\�n�m{V�a�"OR��U���
�:m�-C
	��"O�� �C7-���G��{�6���"O�h@$�Zy��1�l�&�fq� "Ox�r�+YjB� �H�d��|""O Q+"V2f$a��@-a����"O&�5��sL��,]!p� �R"Ox�XDIV^U�E%�n �"O���(O�#����}���J"O���QB�7��lz��
%����D"O šq��(����AX6Iy����"O��'�J��a�� ^v�<�3�"O0jr��
������#�R���"ODPF��>O���o�&5zDܺ"O� `�K�&<ȡ�s�G��:�HW"O�A�b�=q�\D�Ň8��0��"OZ,ɑNޏu=�<�瑳"o�`�"Od�[T��8Q���r�e[B�)""O`t�����0�K�kSPL��"O���숧F��pz$k !S�N�С"O��:A�[�i"�A��@\m1��0*On�r�ME킽 p��4�$�	�'�P	�nDU�<��6L�a��	�'.& ��Q A�ɋ
4V@`�'&}�fK��՜a�6\�����'�z��㑶~[�(Zs�0�K�'����⭉/R��[�`вd�X<��'��ª��R�岴��&WT���':0����?��ꖯ.P℈�'f�q�7"lX;V��7�l��'IFPq& F���<8a�+�, *�'kЈ5Y)��P��r�����'$��(�/I�a"���ƫ,_�`	�'�`��b��]�����
!A�T��'��QD�.Gg�)���� MV���'�X�T���I���# �xɒA��o�<�>)G䰻�J�R��"� �j�<9&���,�l��d�MF��Q�oE{�<QPpf�9 ��Bi�a�<ф��� @�����>�j@�v˞s�<�J
w  \x��b����v%q�<�b��  �3CJ��BDol�<y�f���4�S�HRT����m�j�<	�瞲!Ҫ�*LR�T���f�i�<����-z��ɒ$�G!X�.u�4cPd�<��_��L�KR��(�8���^�<)��%	� ����p��`r�M�]�<I"��#�y4@�>s
�m�� o�<Q��J��4IҺ/4Й(c-Vt�<	��71�ؐ$��h��i�S�\q�<��Q �$�Rp[�Fv1 �c�i�<��k�j�h��c� E:Reg�<A%�Y�pi"(��fQ�PP E�K�<�0*2T���d�v�D��@
�b�<����FFK�U�;!l�
���^�<QU�K?S}F��%T��Q)&D�<���&z���V	�1�����h�<��e ^�ܜ���ѡfY���7"O̓��+�5�rS�N��z�"O4�����	n�x�D�B (B�t8�"ON��㎶��ɹ0!R�656�H�"O� �sf$#���Au�ҁ'p��D"O�){�G�.��{��;!�!�0"O��aP��T���0aE�<r"��"O*=����Kj�Z�C�P����"Ob�@�%PN�`�`��NW���"O:<;�� &[�pT��A*H2��e"O��p�.ΰ~Jp��G�[+бiP"O���mK�?F|�k��ԇ{�HA"O.8#� ��bQ��B�K	cX<�"O�yY1��;_�H4�#J�+|��p�"O��X�.O�AK�m!��0E����'G&@{.��X�`���4�l���'g"�I¤Sj��|ˢ�і+���ʓ<Yp�S��2�f�1r蝚T�Ru��652@�a��byވq�ܘoΜ��ȓ�p��7^m�ޡ�A��(�*�"O�8�G��*:��0��:B` "OD`J�,����2�`Q#N4r"OH`:�O���,�h�iބc��"O���cPjptHΡh��m�p"O	�Ӫ�eOL9�b��- ��X��"ONm(0EP�jj���e�0���;p"O�=��� Q @I��M�6K%"O�2G��(h��A�7/}DT)�"O�-�A'@P �S�Ϛdy��9�"O:)���G��q2�2�@�`�'4��" o@�@|D��e
m�
�'l�P'�	"!�F���V��	�'<���"*E'[�hp��ゾTxVA��'K汢ק	�9vx���� N�H��	�'Ӵ<�G�	w�ЈS�I�t�B�'"4��iٿ}�HIq!o�Q��%��'�:A;QeW<Zi\�I ؝N����'и3"+�(�I!�*�)����'(�Bfʄ�*6�@ke����'�f�!a�ö&lA�fއ~vT\k�'�6�*&ڔwI,���ĺ���'S��;��нb�js.J�7�!��'T �0��P> zjX�ۭ|
���'$�б��	~�@�:��ǭr;�8��'y�����J�b9�G\�`���'Z�����B?L�☚�*��N�,m��'�H�*AA.o��A��j�M��1�'2���f��4,�:3�;J(�+�',�YAp`�;%g��Rr��B�� `�'��\��K�Z5<����6r�Q�'���̈́�l�x��V�X���K�';��Hr�_"S6��pӂծ^C�z�'����E��>#�0�q�.��q�'�Q�CCݰ(b^�
R��-*�H2�'����@(	���C6��S�5��'�MCn[�Y?(���kǘ��
�'2�ö&?@��$i�(Zi�ъ
�'�n؛Sb�����G�73�F�	�'�tc�]�ot)�7�]��-��'1��ӓ���i��胆�қ_C~xY�'�nѪ�"��h����E�C;0�
�'���
!S�����V/=7����'�D��7�~�ҕ�'�#2�4�p�'Lt�s�&��Cd`���'Wh�q�'�l�;��#5Ǌ�1!��T����'���C��4_�,��DµJ'f5��'	<A.�$mG_�x�DX�'j�i�d�_K�����ާ��	���� ��r``�$K�ؘS��I���@$"O0���@�� �ds�c�7��p�"O4
���=R��'A?u����"O��R���<R(Հذ+���h%"Ol|�-;.���O�2�����"OLX�Q	�S��C<p"��t"O,9�,C5I��@a�+�ZL��"O��
1fM7R�dS#,_�P���"O^l���K0A�PjD+T�?Ҥe��^�xE{��I^%�:-�#�\?C�^����ƻ7!�$��N�0����C��U( ��"m�!�dF�a�,Z��D<1)^��-�!�$
�.n���T�h��sjʽ'!��"2K��b�Իwt�U�E*ɫ*!�DX������4`V~x�%����'�����Ɛ8�\ S��H6�|RH>y���)�	�t��]Z��G ?9���D�;L�LB�I,{"�D����Gаq�0�R-j%�B�I�Z�Blk���%@�@]X ���i��B䉧|���qƀ�a|�QWC΋_[�B䉴"W����#�L9AS��ǐB���ީ!�.R�,A,��/��w*R�`F{J?�Q�N-��(s��]�#�^Yx���<���?q���?����l�����V PJ�B�H%;�!�'A�Αs�F�S=����^�5t!��l� ���5{�`x��(Ğ�!��'y
, �D��=��E@
n!��ӑx�~i�fK�2M�09��EM35!�^h�T��Gy�	s��!�d+�:Y#S��?s���
�@��!��9�>�2C�A�sPԫ��J"�!�$�!��؂�C7 =��SՌY�B�!�Ğ�F�`:��  �m�gč<�!��E�=0��Z��ԍ��wkQ��!򤗕f���h��znX�۲J�	O!�Q?J�,ذ��(_aH��R)G41!�$��b%�}i�D�z�i�-�?:R!�$�5
ūj�&�=S��5_���ȓ����o�b�f3`��\0���l���ʻcP4��rI{��$��n5|�vj�00�8����9H����(�(ā2ČX@\�0��x݅ȓJp�Q�F�&�tL1P�V/�t�� ���j!�@<f<�KnFuEb�S�B�bz�P<����B�"GnC�ɉkF$���A��B���Å�VC�	6B�� Svk#]�ٻ$��C�f@,�Rb��"m��Mj�%]6wVC�>1T���$�:E�бi M�%" :B�	�l��q�1Qw�=˄ǎ4:c�B�I+e�z{#ɓ�Q���2�f��'���?��hOzZ��t���W.\2*�X���)D�@�	�|ވщ��UB�ɧg)D�J�'�=���A�A	"���-'D�| �ܛF(��|�[��L
�LB�I�xI�0ДoZ}�z�xÄ�T�!��U�H�jN�=K�l�I%�$N!�$�@��(�G��%�=�g��
 4��)�U��us�"�2�4�Ї�Β鎰�'��4����-f �`CG�@�m��'n�҅X�R� �J�M�����'�5;�g�6�4����܆PN�'��y�'ID�(�;�M�#^��
�'���`�!F�]:rJ�<=���
��� ��Sd�X(2R��%NO� c�բ��$�O��}��"##2��;,W��P�u���ȓe|�ꊱ4  �7�N�f����ȓp5��3�,��>��&�5$p��ȓ�h����w~q�`O�.P�����0T�DJ�G5>���@H�7����_~�p�6�K?��88EM�(q[z��ȓ?���Rc�+Ym����!D�v���Iu�''f��c��'9d��F�/	�f��'������	o
 ���M�yD8Y{�'�@q'�H)ڊ8Z�Ț�p��!��'.��i�Jގ	���jѿa��M��'��q2D��Sy�Ѐ$茒1�d	��'���)��/*�x�R-I�V2vi��'��il M� �("��<Q��	�'Y�݊Ġ�:(pbJ �]&̻�'�p��D�Ua2XK�	��g$B��	�'�0ԋ���.-�|����S�rh	�'0�3`��#Q���j�H:���'[D]h�jY
���'<_�4x�'�x��O?�$�"�%N��'�n�ʂ�L�4n�k�������$�'~F��#i�}gl��',#y��ȓU�~CQd��b�A+Yt��ȓZ�2 QwbQ�q��#����ȕ�ȓy�(Lz�`�<T�fe���=E����L��K��J�]��s���8'��!�ȓxm���6�07(��� `X��ȓe��\�����P���	&Qq�X�ȓ5X���):��X$͝i�:���9�@d)D�����X�g�>ö!��P��D�)4�V�y��= ���u
l�iKC�ʁI��ـ:�zi�ȓ!�N�j"�A�>��f B:h�>���i�B�9�a�zYT���Ǎ�W����ȓQ�B����0Zn��sa_�_b��ȓ1��Q�!A�Y��bI��{Ⱥ��ȓ^�-��M�s�DyQ!��x��y���.�9��#�xQ��� �a�ȓ[ά���ȿ+CLM����;ô���()hJ5`ΌL�(�����Ar�̅�Z
@�XP�#E#0�y��EVD�ȓ6%򠢁Ł9Z(�pbN9����:3���m���F�������t�$��J�;t� �"�G��N���_� D�6�9n��*7.�48�ȓW��XK��l���8��_�t?X�ȓcA���Q^
�@�Q�*�zمȓu��1:�	�b�"d[�٥a��U�ȓr�$C7+���VpZ!�S�?B���u�nu风К��,
5hA��e��fS��Є�ݝ?/��r��M)D��ȓY<�0K�RU���؟��Іȓ[�|� ��H�*��T�K�N���@���0A &��Ю8`ڜ��E���Ԃ�g�J�JT��)y����q�Z��AF"+����٣|��D�ȓ7�WcQ�W��0#N*\7\��ȓ|�����1w���'�l��i�ȓS�$`��v1��k��P�i�x���cs*u��&��i�b�{�(�%`�L�ȓgO��%j�1a�mӄ ߚ]����ȓg��)~}���`W<!�ԙ��i�VyX�E6�DLռ�f���S�? �z�FވP��ĉvC�Q�v\ʱ"O`Hue�+����S�b�t)2"Of�Q�Hˉqq�G�{fz@!"O��i����P���3B�_C�`�"OVm3�Fd�>�p�A��+=0�"O�ɺ�@L����C�ʜ�]/V}�C"O����M�_L. :��+Or��"OxE:��_�+G>ڕ��9M�M "OXXcu��Y�x0#	`��D�"O��#g�M��ݒ7K�29���k�"O.��vn�!OG��1
��f�0�1"O��$B�4�*=����'b��"O��oK�r��u����΂��4xJ!�䃍Rx�
6����| Ӆ"hC!���'2���`�)$׀T�P���	3!�D d�TH�Wg�N��鍪$!�D�.4�h���@]�x����2I��!�� .�K��Q��EhO�>��9�'�X�񂀬�ҡadJ�7�:���'%"���G8Bv����3z�4��'�N��4�P<jϠQi�`�w�J���'Z��S͞�TW�i�0&�j6�	�'88 f)��b�x�)#j���B�'�,80�"��c�X=ۇgC+b�$��'����A�4G���[�!��o��p�'t��KcG�(�"(�F��<�̙�'`za���54#hl��M�/x�	��'ۨ9�!��-!x���䃤+�����'��DZ� �-��0��]����C�'��l0�"�w4��װ�!��'Ϛ�+�
8/�!�hU~�ze��'N�Kvi��X�v�i�+�,z�(S�'.�!A�F��ū�D��RL��'�).��}�n-�Cȹ
�����'v`� A�Z~� c#�
^\���xR�V�?���ד,��=Zज़��y���`)i��+�A�����y*:�pX��!)0֙��N��y,��6T�1`mϔVlB��pd��y��csJh��/?5:ѩ �]��yb\�J�f��d�	:�������y���$H��������s��C�I�e�qɒl;F�H�!�U"oc�B�I�X�Ҭ˳�1=T� ����vh�B��(܈��F6*�̙���QG�B�I�M�A�0'  �Y�'�ilB�I�K��T�ϵZ�-�2B�I�l�!)�4��EH˔e�
B�ɵY���P��
�U2��Y�`�6q�C��%c��ա���K�e&cEI@�C�I	��ж���>�bģ�ÂZ�C�	�V���J���D�cn<r܎C�ɣBIܭ2�(^�.�L��7aPC�	�op�5�����dl����dǷp4lC�?HȦ#��W�+L�����I�4ZC�ɏ4}49��R�����\�c�bB�Iu�<� �e�H8�&��&8B�ɾ @���(h�4xpg�!
UB�	:#�ԋeڰy��`�͈�q�C�<P���Q�~���J#I��B�Ix��`sjѲ6	|��&*H$3XlB�	1%9���vF��e�!�i�SU`���Ob�Or�}�0�-b�	�,s���&��Y��Ԇ�m�@=#���!��P�"�6�`��S�? �� ���:����N~jh P"OH�{J۩j~l!�ʳo���8V"O@���'_3V�n��"O 8����2"OX uBh`��N6�*���"O��)�C5t��@{�ᅮ4���Q'V�h�'�ў�O�$���H�YlH�K�x^(�[�'��a�Ga�6��C�	Ԥl5��K�'��r���wb}���^^@�Y�'�V1��/2�Z��m�Sshp�	�'O����eN��0��R@���{	�'���RJ&IG
�s�'L|�	�'V�D�K�m��̣S�H*���	�'��Q��\�h����&�C�Vps/O�=�����x�\;
�^�x�cPK�98TJ�y�G>D�D�!��|"|����;���J�!D�D1�G�_���r&F��`���@2?D�<a���!6�M�7��*�j��)D�lr��p�<pG�$hl2,�r�$D�LC��P�x&Q���CGc �+.D�0[�̡�N� �&��kb/'�����虛-�%��0妄� �~��"O��`�b�[Y��Z� cg~�R"O^�#Yq"$���Tk�z��{�<�nݒ#�=AW�,F�@6�[P�<�  J�o��AJ�+��`��x�<I��B�n�����5̒@l�p�<�t���̙�Bj�
��p�R*g�<!a��q���t��	d|����c�<��458�aE��^�.#6G@b�<) N@
#�0x+�,�|�d$�w�<)BD������bJ�t,�x�M~�<��PjМQ󂀁�.<�zT�ph<��dF��`K�O4H����Ƨ̙��On"~[� �N�2M�eS�B�d2�1��y�@���o��EZ��S&=��ȓ0t���	QW���`�%x�|m�ȓW�7n�EF�!Fl�$l6@���*��'i�8 aaP�d����yy ��:1Nm�V�C�/0���ȓ�|5X1�K�HȢ �6�ت"=>���Q�|-`4���B�u*��˭.��ȓp����/��%¬��CX3��ȓXLlp��ӡX	ʡy!֭K�lU��=0>͚����zfi���i�n4�ȓz�A���9˰$�R ��0[�%�ȓ2pF#��@W'j���(�+CLH��N���1g��(i��1�b�}�f��ȓW#�i�F�Z�{��S��/F�0���ė'��d��Dx̬za'F�?�����D�&�!��7R�6yړ$��:�0}r�,�}�!�dB.<�̑����T�ȁ�7	-�!��G�ڀ�v� )�[�M��!�	< ��m����(�>�s��	�!��/'��ڱ��2g�@�� �Ȟ>!�D��nU�qC�1dwb���G�|e�y��	6Iq�A�[:8����E�ͼB�	�,l������;�:6J@�a��B�	��$*��m�H\�� "�B�	�^��� ��E<��1oF�B�I�D�:��dP[�H�!�#7-hC�I�r,�����A�!LD���J�nɘ�Gr�q;��An�YzΉ�a���R�C�<5®��EM0w%�@����C䉜
��sD.��g�x����7��B�)� x�Z���"��]��!Ex�U"�"O&y@/��!�p`���݉2�N@"O�Yx�OA�$!����%pj.P�`"O,�PB�AAڇ��Ҩ�"O81#"B�GX��!$��%P��#�"O��Ԇ�(&����ҖX����"O`U ��X�"9�a�J�<T���"O�z��;v{0���ƼQ<�L*�"O T&▍C��2�mX��A`a"O�M2��R)�f�b���`e"O�T�c$��4�j�r�k���RV"ODڧ$ۼ4A����ʚ� �:���"O�����:fu�(��	o��m�"OVxbE҂tE�适ʗ\���BE"Ol�sU�� (����+[�(����"O�푣��/���CL)�Q	�"O�ͨdlx��r��ZR�I"O��D�Q���ȶf[|��-J�"O: � Qń�Ƅ�E��aӶ"OXEr"�3i$�i�Af�6s��pk�"O��BnK[�^�u�I9�l��"O��Qr��9��m�fDL�y�&,i"Oz����ר>T�Ӧ$z��I�"O��Ѩ��x�Y7#��T0F�S�"O8���'�{���S��Î^+�	��"O�h�`�LL�1� �)�@<IP"O�Q���,9����ےWZ�(D"Ot�F�.?J�4sq��u��D"O��ǣ��y�0�9�B��iRF �&"O���!�%M�0����!)M@�Yb"O,��6m���5�ۼdAv���"OR�� �\�D��B��F�]1\Q�"O��FIZ:�d��/@�)�� �"OBGj����tNӭw�~$W"O����I�Ti���M
&�h�y6"OĈrD�
�Vi�G-�l|�5 D"OF8{u/��0�5)v�N�GSp��"O�%���LX��k6�]�"O���	!;˶�*�%�A-���t"O6x���I����`2��A�u"OX��RnΗd�����S"ODD	�n��,G��!�`݌S�Z}P�"O����^d��Cb
�N�R��v"O��K���#T�zeaQ�T��D�d"O4���H�1C�Y��iX"d���f"OBP��OK�:)�Aà�����,�J�<�u��2I��0	��hy��b`�Hy��)�'|�� jt� ��0��ȝ^���{�&ݛ# S�V"@-�ǂU�(J���q�D���MI3����bpC^��ȓ-(��!PB^J2��y$`ԕ+ڈ��{�Ycn�Y9ʬ��NP�7�]��,�P=���)}`���~� Іȓ)µ�wa_J%x���I�H��ȓP���α1�
1B���3�t��BY񑔡
x%�R��_"��E��wB6���W�h�r��V�%�~ ��@l�J�Kι ��r���'D�p��fe<�1��Q�k��%���ĜF� ܇ȓ@;�x��D=ypν��eƀ,̰�ȓP�,4cF�r�|�1׆�uiP���sy2�'��	ly2��˕�L�Mb& ?o 虲�f�4\�!��0'��Db(�XK�H��� !�$Ϊfͱ�̅�|�䈀�P`�!�� r  F�Жt	���w�X�2"O��R�Ȍ4@Uh�3k��й4"O�᩠,B�G.��pa	�]��Y��'�ў"~R��/P8�L�/u<D��b�,���0>�լ��1��rЭ�:"�� �Ly�<���ЄAO��Z���&���d��I�<�s��l?z4�eȞ�dV�iA��B�<٣B�D�D��BN�&4\iG�A�<��k�넕"�,T�BäX��.N@�<�P��~d���~��ܸ��Zw�<� j�Q3T�bc+_� I��P��Ο��ʟ`$�"~2�^�c0\  B*��9��戰�y�N*N68S�i #��g���yBM�*�r�Z��Z(�*��$��7�y���sR$	(0nBAL�RĊ���y���3l��L�f�\�,�,L
�M��yB�D�kY�9��Q�$^\�r�Ʊ�yB��f�����l&l��ř9�hO���I�X��Q	���-/�-���X,d!��(��|{��{�8�W�,�!�@]=2�XB/8D_�USBK��.�!����(�8��.�`Xl`�!K��`�!��	��BE>|���`�O
H�!� D�@��@M��4s��v�'�2�)���S�D�I�R�*��i��*����O���$�'
�D�ӗM�00�єҁ>�!��>vO�����Vz�AjV��8!�D�\��#�ݾcl��Ȅ�҈N�!�$�3F:����܂i����	�Rt!�$�?I��ٱ�ڏ_Y��ʶJ��=r!�$�Q�����5YYA����#�!�dͪ=Zx��!A8?(l��a@?a!��E� �qF��N!b�q�K�,K!�d� 9���9��>r�P�[�l�!K2!�ա/�f����:U�5�TKG!�d]ff�H���~ƾ�SViю5!�Ě�W	��AFi�S�-�
b���ȓC+��p�n��+*lC���*�~��ȓIBT���Ǿix�M�d͠cVP1F{R�'�&(��$%��
�cY�M�����' X\�F/�ER�U��(Tn��'�l��Bჵ5ܒH����YN]�
�'�}h���;����UL� (J�ā	�'�8س�.4R�e1`��-�� ��'L��c��&;[�p�D�\������'���j�@Q�]�XPt��@�ZH>(O ��I�,s��'�� P���Z�*!�$X�=��c �n��S��0h!�d�_ Rq��g��v6U�E�ƤpX!�Ğ\��0���A=T�����\}P!�d�����6�ꘪ�f�n�!���-)����ΊTڸLBe��U�!�D�h�FHR�JZ�9�8�i�BG�L �'3r��7�Ʌhf��F�	�T!�K9'B�	�jk���E��F�r {��'��C䉁3`m��Q=���t�N�y�xB�IҤ+1��+#dڱ�勽sAC�^9 ���nΨ;������T C�ɺ_o⹊�؅X'bB��"��B�ɟO��4��b���t�0���}�BY��@y�'�ў�O�0��Jh1��ksƈ�R�R�'7�A*GE�I�����47Ʊ
�'e�\"�¯O���h��34pI�'i�z���L�L�сǬ#������ �C�e�)�� !�oP�v@�tp�"O� �'O3l���^2n�Р""O�AH���7�PQ'HJYh�6�|Q�@��ӧj��0��#,$m�S�K* o�B䉰c���H.P���sԪ�}��B�	� cB����D�#���ȀbO�z��C��&�^H`v��	lV��o�	�C�ɩ@�"��ՠ� �z��F��#+D�B�	:L�v�	S�w)��(P;R�B��2 �{UO��	�^Y�`M�V�B�	#|1�,;�E�>>,���/aшB��3\ܩ`l�`�(pa�%+�C��eQ�]�s�Y X� U���P�\\C�	��$K�C�U� ł�f��^�C�I�"�ͣ 
�Z��iy��F:ve�C�	�x���wa�UX�Z 	�2��C�I�5dvU�I�(Qi��6�O�T$���D����� |��j������;�""D��	�b��W�H�ďͪ=��4S�>D�Jg�:Ot9�����-����@�)D�� `�݃:�L@􏙆^�b�pC�%D����$�����
]3��ԠF!�B&��\��$*��)gbX�!�Ac.
����k�*%� o͔?pў���K
ņ	mE:�D�*'��B䉱V�a8�E�9Nֈ!��*��B�I<�RpuI�����H;��B䉼/^�e�Ԅ��`�l0�u	�'dj�s�@�5Kȕ`�DG' (�
�'�)"'�j
�1Z�K��U�3
�'�ŚgiF+�*��G�|���'�(��C�8���!/M�V�Zz�'(��x�dʴFߺ�+�M�2a�'Hd���k��|���B��܋N��h�'�`����?R�V83�t��'d
T��$@�2�JQ��H�'Y�)
eN޽	(���?��XK�'	��+�O�e�����˳u̘d�'���sFI�0?����uL�r�'�:����O��&dShNt	�'*lT��-]>A���"��>Ø)�'����3N�W��x�#/� Z}��'���35e�Cc~`24��%C ���'/<�����+w0���g��x�� �'DLq⑪�IaH��rcD�q��<��'�Pb�"�.���+�ۚ|c�x1�'��i�Bf��c����F�yJ%[�'�NU�B*L&��T�V�r^� ��'�"X"��~�42�����
�'�];P��5<�0z`ƥf/L݃�'���1V�M�x5:P�8X�P���'�c�gE(���G���d�q	�'h�q�bB�b��7�a�k�'���뷃șcݒd���O4JN,x
�'�fSa��T�9Ч�>NL:�	
�'�&4x��B�t�XtϏ�G����'ڦQcD΂#�M��Hŋ7V���"Oؠ:�V ����h��1�p��2"O�F,F�!*�颷�ڜ��7"O�5���W�����O4VP&e�5"O �p��ִx�@����{瘨h6"O��1G��~ʦu��-���"O�PA@����
Ԏ߾N��H��"Oș�d
�] ���$��n���S"O� P�c�4'Ȏ� b�
�B=K�"O�"�k�)�쨠b�Y�!6�Q"O�`�c��<E�qQ���
b>y
�"O�q����*a,�����Y�?�u"�"O\��4OҾ�\h1O��_'I�5"O��
ư}[~�u�T�j&^��3"O4��C$�u!b$ݞ	����"OD%Z��.�6L8�r��Ѱ7"O��P/J)^�ڴBI-��e�"O���2���2��ź�@ڿp���"OA���!>=����׌Y�&��b"O&@��Ǒ h�̌�$��n����c"O����0���C�S;8�j���"O��̹B�<{wBٯ_f��0"O���"a�g@�~^��"O(�@`[�E��(2�	+kh�E��"O
�J���_�F��4��"_P��Q�"O4Q���\8&(T9N���R"O���P�Y�&,�����'G~��"OjP�FΧ���Ƈ<l|�6"O���*�z�Z����0��0�"O���ŮwjԸxe�F^gҴ��"O��sR�/b�r%�ʣ'`��s�"O�-����4�����
�+QlH�"O �'*+�Tv�G+�6���"O*DK�C&}p�X7�H�*��"O�؊�CG}�2hR*�$*e`"O�D���
��U�刏�f�=AB"O �bvb�R�JӍȳG�h��"Oi�Q�(�6��$gӚs�T�*g"O���PT%]�\�qc�j��5�"O\�q��fF� 	.@hU%T��y��e���W��l)(���NW�yb�)4Fa�'�<W�mSW�Y��y�����U]4;�<dw(_��y�["XȦ�bUK��7ߺ�ba�C��y,�n����E.ؒG�Y�𥑄�y�3�D�S"ͣD!�us��X��y���0x|ZQZ�+��Bp���Q�׷�yb��(|D��"�]/V-�JG��y�+��j>`������$��<s��I��y�6'0T��ϗ�#9R�aЊ2�y��yT����n�/�����^�yr)D������)��(ͨ�(��ߎ�y�,V 4p���%�)3�
V�ybE =O��|�S��P�%k��R��y"f%F(�b�0�iʇ%�:�y�h\(���t�08�N�*�!��y���`t��!����3I�E�Ō���yBl�/p� R�
��x~��"�j��y"@�Z�h		R��4Z���R#���y�DD���Hk�U @����c�^��y����[����#��
<��\k�'�9�y��O�Ԅ��e�F���0�jA�yb��ri�=DER������y2h��>��;��W�<^l�P)���yb�?AY�QRNߘ-(�5B��X�y��Y'1��p�7V8n���N��y�]�`�:Q��|ڎIc�OP8�y�J�N��I�d�.tP�����	�yb��y�v�R�oY�sx����Y<�yß :�|��$f�o��M �S�y�kа ��ɹ�>R5*���yr��:�}rMK��|��b7�y
� R�����~���#���MG�y)C"O���[�&|�C=!��I�"OB�{D��Q�`��e֡x���"O��"�L�ef��4�8�:y�"O��*Z[���q�^�0޴�G"O��`��M#��)ŭɟ����u"O�(B@�O+t��@���<<����0"O���OYN�:t�w X��%cZ��y�iQ3��)�bKL7h�&��ΐ�y�cL~%c��8KЎ��'�ý�yR��Z]��i!4Q)	��Y�',4  g���� J�Hz�:Y��'���q�#ӆ8��[��2L��	�'�B�����7"a�d��m�0Q�
�'��	�0OX!'��-�R�$O�X�	�'ќ9bs �t�A@b�0A,$��'~��q�J�L��ZfO�<�����'������*�qau�̞4o�5��'��ұ��3+�N��D�3-r�Aj�'U(E�FT��~]�р�%x8J�'gp+0��� iE�t��`
�'P�uS��-uZV�y��G�p�j��	�'�Rq���8X6(����rO>�K	�'L��"2nP?ݰQ �gvv�2�'(H���B q����L�&o�~M��'U$h#�
�S������a!�	�'g�1+G�
'���BAO�ia#�'ŀT�f
'+ :ABUIJ���E �'�T0sU�4v�|�!eBү#d�1�'�pi� ��j30lID�Źq7"���'��-��c�,Q��{�$P���Q�'l�'$2Ѥ˦,�&� ���'.Z�С̅J��9�V��8�
�'|�,KsT�5��3.�D�gϛS�<�ą�8f��d�Ô^2�`��R�<����]OR�h���Vi%h���d�<Y�Ր_v�pp�Cх7T��)	`�<�!. :�t����<HxZ��4Ϟ[�<)���8���(�*
�T ��p [[�<��ƌ����=�|x�TŋT�<��Q��Kg�W���z��]k�<���O���q�ܖ5�z=���N�<I"�UY��ag!�"��4Z�	�s�<q�e,U�D�bDf� WYfuh�S�<�B-P(@C5b�H Lg����M�<�+S��>�;���"<�p@($C^�<u+� bv�q�t�)GQr���c�<�V�^>;�,�������p��� \�<a��[�c4��Hbڭ:�\��*r�<�m�[����(I�]�P��Do�B�<�G#N)Q�����mm�JF�<Q��˭	%b���O�>|.���$�<q˂�k��)&lQ>WJ��Z#��}�<�E)Z�C�����h�f�����U�<y��lg��F �,8�	�J�P�<���3vL����Ȓ& ��2�LGI�<� �')�b�ʄ�]b,q
�j�B�<� &]�u��̂SF���1�T��A�<��.?G@�5���DqY�I!@z�<e
�d\Dn��@�a�2�yr(ښ3�<91��.=n0����y���x�3�]�7��,��IS'�y��ܭ>	�	C��YfA�fX�y��������@��V�T�3�݈�y
� $u�E�=A��<@�#YTmHP"O��5N��>|u!���V�tP��"O,�a��]�_~@E���E.�Y1�"Obl���ʡw��ZqnM7���A"OVk�K3P�tM��#~<zS"O$��69S�9��?2G"O���*i��"�t�s`"���x�<��˅k|ne�G��~��}�x�<QҊ�:��\ٱ�ދ>�v\���H�<)���.�f��� ��H�D�G�<����*u��Ը5,�1�� ��Ai�<Q%��
)謴�R j���
b��h�<)V��5	�|г�53�VX*���o�<AɺNK�@$Iǧ|�Iz��l�<��-%��)��)�#C�8-*gE�p�<��+�F 4R� �^����3G\p�<A���7'�QSCF�8���W�<���Ҋzt�����]�
�P͊A�RG�<qW�J,Q|��$��p��գ�<�d�ӕG"�ש� a�E�"cV�<�C�ݯ��Jf��m=����GZ�<�&ǟY�}��D��*�4 �P��<�ݞG������l� ɱ�DD�<)
ɷ? ��u �x��p 	k�<�F�AB�p�/��#tf��B��j�<��H�3F&��vX�ln����@�<t�V
�����Vr���B�<i�H�BS�$�fn�>bC Y1@�Z�<��Z�F�-y(��u�YY��M�<Ac�9�0�%��+R%&�8f(LJ؞�=�a}���J�E^�B*dH���E�<A�փSI"qٕ��.+�r���NJ�<If�'հ�iiԳ7�F�I�n�P�<��A�nf��e�ƭ��}��N̓�~R�~���Ĝ1hf����F���k���K�<1J�,*���`l��h!��ǬGJ�<���[�t���K��	�l�yp�SC�<�����c�΁���X���H�<)�AL
TP�N�fĄ�E�'�ў|�' I tTq��B��U*M��'�:p3d�D�g�(�j �ԍt���	�'�"�:��)��(��v����'g04�s���Ȱ5ywA�g���p�')��`���� ��� ga2_Ɯ"
�'GtⅯ@�Z��J�[�7-JUI �&D���挙pXIJb��A܈t#��#D�0��l��=�R�,�/c�| �D�"D�0с͋��x���o/^h������'O��Y���$J�4��xi0��'J�B|� qӒC�I~4dYBW����!̃�}��D�B��<��O4�@Q3lgd���K_�jx\Z��'��'*P��kv�Y����&=�<��y��'B��	,�'^��QT�\y�[W�޶Ʊ��	2!��O������ `��O(Ԧ8��'�ў"~��O�s�ję��t_Z�Z��'5Z0��M۟'��)�i�/K"� �tL��l�r�m	���c8��o��F�����Ԑ��F\9Uh�}�'�ĉ�a� ��~��~⨚�g��P .�e�ȁR��-��>��O�����D�f`H��ŀV��ը�U����ɿRd\ �S�D�F1z�J� %O�~����?�"��9]Y�� ��i�d�T�<�f@Ihdś��T�_�ty��Oh�<ѕdȱD8�u��C�PX(U��H�<q�^+�0�� K�1�ِ&Mߺ1`��m�L��t�S�? "��b��o
�9��
-���ku"O,詡��_�`�3����U����C�'��OpE� �*qu
v֨;�~L0�O���ъ}�̊5B�* f�h�^�!�$�"骍�&&�8N��U��O�!�(qy8�@-"��䐗f�	E�!�d�5Kd�Q���X�ct��^�!�dܖ?�Հh�iڒ�!���={ar�ON�`j���T\�C�=��{R�	�<���	J?a>d���� w�:9P�)ךz�!��?���u�H�x��Hպ-�!�#x�z�L�6kA,��g�^�!�䓊;%�S4�Ɠ.h��g�/w7�'y�|�e��%�l�K&EK�?J�����y����2 �Ā�����Ԃ�<�yb���I��:.
�ܻ�
	���M+����Y�>�H�ǃI��dM!��"R
�i#�P��r����&!�d�i0]9�BX�w:8�!��U��	�'����I^?+O��a�D"L� �� �E��)�l54���7��@8@�{0a_`jF͛�A6D��hA,�rn�{���G�%�&�7D��Q�Ex��
�%�v��P��6D�|[SD�),X[BHDb�t7")D�4
A�3R�"�����H"�Q�s�,D�����/,��s　�q�`�2�&D� � �1��a�iD�N�j�Cw�"D�@���"QzR4S��5kAXeBRm"D������p4���+@CF�xSsI"D�t�C��y�⠚%�ߞ�@!�S�*�d-�OPa�`^1;��K�.�*���T"O�HY҅�#]1�\w���t^�m��"O~�0A�]+?��9	��S�R4��X�G{��閅=���B"`�5vLM�c�֩bs�<�ߓd��xgCWm���w��.? ���IJ�+�91O� ���ᕿ� ��k54�%��2��BwL�w�i�'V��?i����@	�(Kq�z�H�H�ġʲ"O,8�7i��q/2�F׫n�c3"OF(���,o� k4��V��y�"O����߯;
t:���O]�����$4\O� (t�T(D���B��BURUhg"O�P! (R�Z��b��HT
�"O�x��F�l	�	h��y�"O�r��L&'�|u)�A� Q���`"O�Z5��v.B�W@�LGt�A"O~E9��N�!�����(� -�t��	h���	D+*k�p�酁Yk���N�"e!��m�Q ��)��Y�'(V�G�!�K��m&�� B���3%�$<�a}��>�B*�6`04��"�����A�<����'5���B�cneF�^����?1�fWg�h	��b^NT����,Xz�<Y�l�x�&*���.m���r1��Z�'	���O���1�E�l1���Ύ�]O(��'��.�0��I�Jn��A�6�y�C�΂X����(O@��DL��yRo^
/~��1�S�n�I�ui��n���$L�$bn�[UIЗZ�P��%���!��.za$Jr�،���W	�!�V�8��8�A1��� � �#�����?�H?	`�dN��x� P>n�񘶤0D�p�#�	!��`�cBZ%}8>e� �,D��"0�B�y0��p�3r]M1d�.D�� ��)Ѩ�v�љ��S~8�C#��0�S�S�y�h�vܲj�X@��@7ekbC�g[h�ZU�]�.�
Q^�E��xx�'űO?�n�H��a�'>����n�.i��O�':�O��	�1�KQ�^��`#*�� 6"OH5BPk�!����#�5Zٚh���|��`~B9OL�� -ǯ^�TI�1!>t�kB�'"�'6<���)�_;h0�����@��d%��HejS���RSn�Kv.N:�B�ȓo��T�N�>:,^H���[Æ%�'��'��)�Y�:&�'aP����33����1�O�d/��>hJ�H���&�Y�@ٺ�E�'�,���p=ɀ��*E��m���Bh��cFf؞��=с���S���BU��}��T@8T�d�D&\���ز�+�l��U�r�,�È�$q>��nڸlPV���Ο��Ԡ�iU6\C���FX�6�8g��U�#k ��������Y����G:+���s�Pr�'鑞�ce��B������%m�*���9?qF%!�O�ɐ�X0���Ha�՟| "s �>���)�S͒0�A�
鲉�ta���ʙE"O�1U���m��`���vd��X�ϓ"qO�#<�Lޟ+9��y��%WR�P�*�Y<Q�֟�f�����V� %�hX�~r�E�ȓ��9LZR��d:1)�>L,D���o���B'D�,2>tݣ���;0�ְ�ȓ0�@-�qOZ�,��5��a[ 8Ol���{1��a��G� ��a���R ���ȓ&��Ljf'��9�U`kZj��`�ȓ<?��MT(�l����&&�2��ȓa�fHq�e�X����7Ț��ȓ;���3N�56�=CV�1�XĆȓ�P���	n��S�(_�fE��l������;�]81��*E
nH���<��`I\��pb5��9����ȓ2�f��%�|���+Tfƥ�ȓ��b2 �M.�:�#�	pپ0��+}��E�д\cu2�,�t���ȓl���@�\-�`� G��!8�4��ȓ�,{��?<����M��Ņȓ]8����J�X\x�d��K՚؇�Bh<y�0d߷n��5�P��9,6���R��E{CQ-v��!G�,�xT�ȓ��k�, �*8�D��s�Շ�:�}�0Iy�̄*�EJ)L�fi�ȓf����ǂ�\` ,���ʝ,�\І�&:rY�S#�7"�ԩ��^�~'PɆȓt��|i0ڶ,ji�a��?"�\��_hN�!Ƨ�
oij���^�+�̴���<8"'[�9�ڸ�(�5J�!��%Լ���B�&�8��y�HC�I����aޢ4q$�xb�O6*��C��WR̄
7�:(���F���Z��C�I�b˼�)'�˓.mF��t��"��C�I/6���e��X���HʷTp�C�n�!�ѷ]\
X`Q,�k�jC�ɅC*��q�E\)�1C�V�@C�ɪ7%8Ey��8#K�.�s3D=D������eJZ�#��3�6%���0D��"U�H�y	x��N���Kcl-D�0�O�$e�v�q&*�6�ؔ�E�+D�� +�1�8�a���S��cc)D��㓦UL�N���e>5����V�g�H���]Ux�+���/n
f��cF4�d�Y	w!,np-�a	l��m��S�? 8k��'8x�A�eʫ":~�ɴ"OL$�r����Ph�Uf�c�A0�"O�I�@L �F��d��K|�D�G"O�ik��?~ո�S�Ǝ�O~8��"O���f���:��sD�0�x��v"Of��W�~����<_�v(�g"O�uB�Ƅ�2�UY�fɎ��%��"O�8�F����Q�.��s�"O�!��C�+N �H΃�ԭ!�"O��a��A�:��2��F�8��V"OZPs��ԃQ*���bݭ&TD�p"O�x`�%��r�X%�[�94H���"O��(�ߜ��XX�o'D�4���"O��#�=Ԯm���Y�b�ԁ26"O�PqV�K�Ah���a��]��ce"O��$����A��.h��(c"OLIS�I�qĤ�QH�qh$yP"O�Q
�-�|i���r�V�O`�#�"On�K�Ƃ���lO '}�M�1"Oƽ����1/��I�.˂����'��Y���{��=w��y"tm1L�I��c��C�ɖ+Al�i��߯HJ�L뇏W�V��'��Ё�o�/�6��Ӥm��ͣ��ǇK���%7�pB䉢m�-��]��+�P{��=�F���<��кS ��'+�"��Y��3���3fn�+!8����V�2���!3�mx��1�ŭb垨�W��=	�	4�'F��\1e�G�~AP�����Ab�ɱ��	YO�zE�4��'��g��H�#/�W�|�T8�2���Cb��X^��їEN* j�]�O%܀�ƈ���X��w�� [s��E�͘o�"��!��6�{���0�+�wr�\�宆�8�uy*��j��]8��M�Y�z�C��|�&Kut�@��9�ט�X�v؀��O+e��=r�w�B�I�KxP�2%,��"ޒ����9[ �=�Ǖ�S�Z@bm�@���E�Z#H~X�2<O��A`��^,�睑;H�A�weC�m�"ʖm�*��D�S�:HS��I� ̢Dz6n]<<��*��ǲ^�f���c�%d��ͻ�ˈ �?�E�95�p��>8�� :�{��I�����+,��pz5���O��� CD4I�L1m\PU��\�nt��B�&H���3fS�&YLP�� �<t!�x�`K�;i �02��	4ȇ�	�h��1 f��w�|Ĺ�IڙBY~	��i,�7��}���yWi��=�t�1O��B0���YB�LH�.���4 3D��`ToҲ%�Q2MBŸXR5GЈB�*1["K�"�4�@�$Vp�0ԏr�f=J��/�Y��O��IR�L�)iF�l �#UM�di�ff��� ��v�'���겍�9&�-p��L	m�hP1S�W�~�~�:��c(������2�r�ҷW(0���a6��h�zD	#ϗ�}�t�
�O��	pG�Ҽ��b-4K���B�5~TdY�����!�Y�5�[�k8�P�we�:	�K��&v����ϖ�L�)��OU37��@:��_~�j�ɔ.�n�P1�'0�Ջņ;bK�/o� cs�
5i�`��"��/�\��6��12�J� &�h/L��b���m�$3Ӭ�1`�L�F�U�*��mB�^"ⵥZ��ֹ�/]���}"���!_Z��|�H�0��@�3�I!-�� #�H�8*���g%�
� ���M30�ν�B������$�B�̳1�ڝ����z^\�����!/�֘{���O�H$c��WZ\`����c\��
�2��OrTq1!�E�XťQ�׾őwJ	Q���ȗ���?T ����Z�|���X�{������
а�ɷ��	Q��Ĉg���`q���!C�^����*��.ؽZ%�"=!���Y*J�gN��b�'L��Y-�%��Jp�h���}��H��19Kd8�T�V�0����h�`�  �ㄆ�Oh�CN
x��`�JC0;Hb4�d`s�4��É���n��V	['�5!�Γ=?��XV�x��4
$�-qW.��:��cЈh����𢚒p�u����Ib�*T'�~�����[�
lH��ԁ�.Cvh@�A�ٻ(�m�&T�(Oh};�˅:�H=��S�\,���ip�����漴�`ʚ"\b����W
.���nJ���Nɔ��=��iF:�<%0�c�+�D��LJY�|�ɓ�R�@:`qD}�l@(˴@���ƞ8rr8Dk�D�&t���C&(�h����D�ơid��z\:l��v���`b�3�jm�"��Ǧ��UoWJ=1,�2Dpd�g@jX�D"8K�B;�"��c�6ĈT���M�QɓcE\<+!�� P�`�RXj#��V�+bghU��5,8�m�"	jd��R�F�S�D��X�n+����Z)fn%8m@�=���d	#
^�T{WC4T�  !Q�;;M��`�4v7��:On Aw��C�ؑ�n�k��!@�"ь�� *�↦H�8���f��n.��Q��e'xD�MC)Og਱F����,Jf�ǤL�2��DF��~B��}M���$�ֈka2`�2V��o� �aMOT�ѓ"�
4��Q�邬��d����;+��H�o��BOJȹ�$��x���@�%��g�~d{d���L^y��,�fX�R�o��FG�i�%�U�{6�j��ԸJ����KOV�41��	t�N��d�]=Z��p9u�h�� 
1�Q*w�.����,� qB���
�)�@���hc�K�Z�
q"�R;C��1��J7�ʓH�3 �Ѭ,:�4���"��Ď1�5����.$&!��X�j�����eS0���bS���-�'l��BDdP6��b�R����Ǎ�?&X�eB�-!I#�e�2AR19 +�B,4#D�4Yh��d����"�O뮄�[�2a�d , t�p���B�\X� ��3��@��d��Go����$ؼ2�(H�K����ef��ZD��s3쁀�p(ۑ+ۄEh������I���Z�9 �b�P�S-bAI��r����# �,��ju�֕9 U�f�۹38����R/x})���i����4��m���`莟*���1N��MY(�f������ ͙�%�?��ċ>B:`�;D�r�a��Y�	0-
x��x�&$�1�s1���ޔ����5iJ�=3A�N8\�=X�m���X���ܲ�@.��&��2��U�,*u%N+��+R� ����W�}�����'
��G�Ǻ����,*�^l� E�H���3�HI{�т�ŷYx���o>!����a�/-�@@�P�֛K���k��	ڼ�ˌ2�(��e�ؾ�#�ȟ,c ��
_�|HQ��OH��&X��I�6m��,��,5���ʕ�� Nx�\�V��{�.���⏬Z9�tGʦlLi�7M�;"����!��L}�L�v�Еy� �s�*�IƲ,�V`�	�#���'k�Ob0��*�P!���!b���zP�1�M�@�D�4B ��/փR 6�h��O!z�5[N
�<�DКR'�;a���H2g��6�l��pGM�e���P"�I�V���S�넑qutCA�V�0�B r�JL�A�\<y��V3ql9�L� W���k�KD�ptt	k!V�2�HR���>�U�C�F�|1���V�aF��@�\�;�f�1˓U�"���u6l�J5��mR�0cN΂R��x'c��VԸ��2��8ݴ�h� ��Z7�y�F� �2��w�hX��d�� ��!�U+ש�`��]�ĺ#3� ��v
@<@QphIpg֪*����-A�k�
�#d��uz��r�^�������BW~tq g��/����Aٟ|I�ە����Xb�I�-:�9Ӥma��ۗ���䖍[j�iۓ[A#����B%]�Y�Q�վ��g��t$0I�OZ�`��/s�D��`g"� 0B�`0#}#V�2�N�eF^�ml�`0/E�V��A+1̉)5
t��q���R� 5nv
 c�W䘅h@@K
"TRvFI:A�2`iu����G�D�P%I��&x�\ʶ��Ph�D���M�7	�n�!I�U>)��IߧR��A{�d��x�2'�U����GυS��	"�D3�OXa;4F�j\�P��,ç.j@�0`O-���A5�^�o�,H�f��l�*ۙQ����&�"�W�uz@"ϛW��X�$љ`Q>t�%��iUo�<��e� o���#fT�:�� )���	WH9�f�O0]�2eAR�Q	P��+4���� ������M#1@�{�����l2x@h@�)bM�,X�Ǒr雦-F��S�lțD�B�\
!�p��`��W���Q�DO#0�ԝ`�F,����._�%lv����[��MH	ߓY�E��n�(��`��QTL�T@�%0T(M�B ZbfH��M6Pb�e��(	��HЦ��SZT��`�5X>e��@ۏ�5�D[�В��6��+z\�a��_��O���k	7-�=	�9�?���>C��@��� '�*`*�'П=��vlé[\��C%Etɡ�n�c�:�.,����9���aw�U1��䊌|��iȢ�s�:���+�`���W���(�< ,g�B��1Tl�#��O�y�T�_�H�R��r��!X�j�s*�$5l$���ݏ
)xݪU�V�:��]b�F��U@��,P~Ն�I�aND�� �b �S3�ĀL���ɗh4-k�$ bL|Cb�k>9C��Y�&bAf%;�b߈T,ܴh��!}9�<�q��|��h��-,Op<Qr��.��cA�DBS�ĩ�,�%|/�t�'�4M��)T�
(�
P��K�/tHY�4a�DZ���r�'~)�d�ڴk�,��J;�D]r�¨u*� �끼1A���?��;x|b��4jO�U�Xb�O@�髓+�5�.5�ѥS�I�.��Ҩ�='��S�)R"U*����C8-� �c�4�(9��œ<H�(���X?�	*4��@bΏa�f�`��S�C<Э
0#,��x&o�O8�*�]�4��P0"��`�b�hЄӪB=��݂/w����#�;�b��&ϵ#J%�ɉJ8��cP�W�'a�|���B�'�������O��Ar���-G����K����d@�":�����ШA��y��H*H���E���`Y�US}�� 2ÿU/BT�IADcayRL�|�L���� *�����N�W-�I0�-<�fى��/��PQ�b1��DV*̀����P!�y �	�%=R,���ٽSȵ�"���+�qOX|��̕�Q�>��0B�/��� N��J�^M9%�r��b�k�����C�c���J䡔� �pM��̭:H.�Fn��"~Γ3�8���_�?W8��V�5�h�.�8I��5��eS�l��M�7�4��ԙ��`��y�����jD�QY��P�FcU��~rC�9���0��6�uF�B#H�]y�fX��9��\s�8P@r��m��(1a2J��A	��!M�AA���
�MKf)}ݝ�$!т#�-c�����^�~�����:<��Ҋ�D�6xg���cy1j���_Y���$��`�9 ��7���$H�*{B���@H���rQy��@���.0��� (��T?1��>N�C#DN1XB���G1�d�`�����b�B3�#�I7co��q�뉛y)�4J�C�T���B^���%ɥ(�m���I< ,�S��ے]��S�O�ҵ�qI�YP"H8rc�g��Ę�g������e�B�"4,1�zzʝ�����٦=7��ͻ(�H����w�RId �O��O�
��@���<1%�,mԨ�k �E��E��FW�cRB�i��!�Y��$�z�K�3,�jI��m�/$�M�=���:`�t;�ㄸp4�3�b
[X���&��t�r0�NĖ5���p�*b	Z�KdD�t8������Rr�j6��9AL��z��_Z���h�U2Dؐ�އ<�p`��B>�d=~�ɘEĿw�*��
���@GY�)WN�;�gѨ|����ЄT�1�G�R��ȓ7�¹�HV�gle�ĉb���(#�]�i�t=�A��0R�Z�`6���1�ҥ�6�|*A�3u?�N�7jc��ːa9��X�R3B!�Z�zlB �w*F?ȎIɠꇂ,5��GfE3y�f��3Lؕ�z$�"c��xiL ��jǛ;���������Uh�(��0��!e�&<O�YH�ȋ�4��l��+��@7`��Z�];���8t.<�Q�
w�P�ժP7'�f�[��'@ԁ`�,�ki�8��CC�q�ഒJ>��#C2s�b��G��5���O�6 K���+DЅ`ĥ@%P�x�*2�+!*�q������y
� t����N� 1�j�E��"�>��T��I���0�)&^�)�ҫOxd�����}�D$�S��杭6�*��a+�-48cL��TΒO6<s5���O�x� �P/fN���@|��z2�N6#r��q�(]	&6-�=PL���6�Π]?"�KA�8���η w ��`�&	CR�B���/!�x�yB/.2e���dU(&���R��$����'��a��M�Ca��q��A�A�h���\*��Df��5/�4�'��y�Ow�q)O�)�L�fEB���>Y ����Q��I�x�\�a�*���H���-J�X����%[�Y�RJ�˟�	ׅ�?�|M�&�ƛ_/��(���p]����mW�l�b�ѵ�
�~���74T:}:���(l�\�PV��_�&A�ҥ�����D�`������50\*]�B(�u�"�,�l)Üw�*I�U��;	۞�*P.	9m�Kd@��䗀vA8�)3DXc��{r�҅^�nt*R�P5xU'Q)�r��#
G$ 1qQ�Gе0r���o�;�zXB�c�0pA#c�-�l����'!\�xz�$\�Ϭ��woM ��`sS%M&5L�Fy�\!Ǹ�؇�L#��tC�̤0ڐ�ї�?�(u��l�>
��bmH�y�����S�k��A��+-ӊ�ѷ >�,e�,�;���D��@�w��0^gZQ�o�g����'�Ƞ��o�	� 	�Ԛk��pK�)/��M�P�S�V��F%M>w2`B�G�"����&F�;S��[G�V"j A��A�kd\�E�~��~B��:/R0l���&u��

�N���Ń'y�X�a�5k�x��+T�)^$L�W�	 a#0����y� 5[���!E���8�۷�ȧ
4Y��	��Qlh8�A�:{ǚ\b�g�'6A��)K4�2v)� '�BDq�@��� @�Ꭱa��<p2�q�+�)
 1�,r���%�\tY�l ���4xCE�{�X1��mT##�|��f��9_Ѐ�w�s�'��A�F��h.EC�gY�+aT�C��<e��CfAF�9x�����j��֠Y?a|X���-���q]<g ��sv�F$>r�����?���D{���1�gD&r�N�il+}rF�N��"�蘗p�h����57l����+5��Ea��'u��Џ��� ��ʮ�xg���s����g�������%w�?U�# �w�
��t���W�����a��y5(� qnN�8�nR���+0��#������!����;ZV�����rU�H!���F=$�i��;{ɬdA�e���;DCٺK���ݩH���j6`�$I	�Ѱ$�� &K҄�d(J�d�\����I�X҄M�I���r M��uW�a� 	�*"/J�!���	 żT�X9S���5$�-<ڕD~�
�y�ȝn�Q@�)���J�cJ�!{�� }��-�sd0� ��ٲe���k_�>CQIc!dC�vG]�}��!�cT>�QaG�K|n��eb�a;d9�*��ŎW	R����P�e�F\�Q��r̩a@�� @j�a��eQ?i�m���n8�&j]��Y��+!�&tlX�ૐ	��� v�8}R��!���	�z�&����c�p�c�oGUٓ&O-Ĉ5m��(�Q�b�#ը�!��1��OL�);�&%`$��'W`\��'�JpRUE:"GX"�!@�_�(�����A*��"eSd�O�([�k��Dx�h��!g�����I�^�ڠy欟:e������$D:#Ni��i�uB�7@ڃ�y2��%#~Xq�Y	{�~�[�\+��Qb �����O�"~�	�7�x��{��dA�Z��|C�I�z*�h"�M�
��H%C�5&2˓I,`c5lO\u��IH�h%jSǁ�AM>{u"O�@	�B �BF1c��##�87"O�@�%��/��Ӏ�(CR"O��CC��G�d�@���V=���"OD��*�,@A��UO	�+^DA��"O|� �!W��`	�ΞpC�B�"O& �s��'C���3pÍ� ��I�"O���p΍8kI��y�%M�J��I�"O�i��Uy�!�vi;�0�B�"O���Ǩ� ��iR�)�[U�Yr�"O��� %��Ra
#fʒC�hi��"O��¢nUH��Z�%	_�R ڦ"O4<��KI�]�N���ܛta����"O�hP�c��<��c]�_�%#�"O�e"e�6.�U��9/<��q"O&�
�h��2@8\'>�B%"OZ(K��ħY@���d S�.'�a)�"O:P��"�,f#и����(���"O, ��Ȇ<G��`��/T����D"OT�A��r`kql��O�2 �"OLD���%I�H1��aƧZ�����"O�����O@�m Ǡ��AS$�+V"O��`6���� ����&@8��a"O.�3p���$g���CY�ycP-�"O`䩀�H�Kj���኶z��'"O��U�ܒKf���K[���CV"O܀�`T0�|x)�W�
�"O� x{�"̈�H�c��Y�"�13"O�H�-!��!�m4�f!�!"O�|ի��`���XĖHٚe��"OX��p'E�;�@�Q2@�.?��l�!"O�-�Ixi��:0ԃ
�nD�"O��+Qm�&w�p��_���� "O�ђ�f�7�F�
%�{�pJ�"O<�($�F�-n!��cL|TJ��"O�q�tE½0�p�z �/G�5"�"Ov�C ���
$�]r���F,Hap�"O��km�FWBD� ,�34��#"O&1`�kH?��]��J(9��)7"O$�F Y�O�n-◀��u�,�8�"ON�ʂ'D(	���U�F�t�1��"O�Iz��?���i�Bi�N�@�"O��䮕��M0�R�e��,�7�7D�DC� �4���3��)<�1���4D�(�u�O�I|ѐÄvz�	D%1D���G���d��NT�HT!W�,D��yAՎl�A'��}0�@�'D���/���@�
,Ej Z�H"D�L�������WŃ�Q>a�Ӏ D�RE@\�q�(��LL���	#=D�L�lF�j�&t�K�<D�U���8<O$p	$�4�����Y��e�`LX�R1L9LH��S�B�V�G%2I���3?�4��O2l��߫f}a�'k���b'˭J]M򃠕�uN2��
ڵDQ�_ed��μ`=
�;��  �yB��&n��+�Cо
�>�G��y��ъ]ʨ��F�H&�h�Fh<��>�f(˼s���` 3d��1��-Մq���Y�D�j cFL�:�P˓9®1 ���1|H�"<��k=2�xɪ5M67R��R,�s�'��u�e-^�d�j�ڦ��*_|I9���k���
|����լ'�z�MN;gx�}��G~RZ��d�Ǡ���I�/P�9i�lC�j�p�0葮mC����e��>��O����ĉ,W�-I�,C���͖:

x�����Z�҄[��v�<"F�b�Z�q�F�Rt���+4%;p���>�|�p�Ǎ,�JMCR�F/c�\�I�V|�Բ�����&=_�h�Ŏzt|5�'dE�Գ�<%�<dÐKʂ7�^C��(.�V����ЩZ��%@�	1�z��"�'8��U� 1�D4 ��|�{�F�++D��UW��~4��A��O8dʔm̠RN��C+C-.�(FC&O�� j�`��V���Sn��R�HMscA��}Q���޿:��mkU.��p=1$&��F��t3@��4 �=�E
Ba�D+�i	�Ze�����[P�|f	5G��x0�5�5D2v���H�n���:D:�Y�ȓ/������:L� ӈ ���"�p��lI�Jᶐ���ӈ���ܦ)i���P:PJ�`�����E�uw`�CK�;Moԅb��B]`8Jg'&,Oڤ#�H��8���(4�#i�!�D��"q��KF�F3	pt���Iv�-rA��;g`(Ӡ'��&c��4'آw��c&����T����5�B}1
�qa^����S��*I��=9N�.�r4(c�v���ԯ�&��&�@�N���ʁ�z���YAӸm.~}XĪ�^���ʘYy�!ѫ�p����%���^�"@�H�FbI> �mQf&؂i���`��
�l,��;q��ge�1��ߌ'J�h��B�<
�Mi6��k��\��b�*F���ፆ\j�)慉�+,r�m2��2ˏ���g��Fѡt`ӌ+���@�>l��ԝH ���Z=���3v�`���K4՘�A�?	,p�۱cƋ�Jͩe�D!�X�袂ٿ��{��ی^\4QrN�/(џ�2l��l4te@�D�Y�LL�anۯY4�� e	�@���%i%����cȍU�ĠX�遈X�BP��X4��p��
D���U�ǆEَ}��&N.3���a��#k��I��#n�4PY#g\�h��$��03,��A؂6W
�X�'P[��aaG��"�HE��6|&�PU��y,�"a� 5R �p��ҌQ_��I1�-#�PsJR�ف%�̆+�::��eͩC��ܪ!���r�oZ�Ү�q�(О^9�L���up��!͊�QF�����S�C�8�B�ꉍ7V��H���	h4�dӮ���(Ӆ�
BA����&]�'\fH�h�g�q(e�[ "�:��4 *}+1��!�HtTĒ&yb��*�bQ��X��
�4�uǉޘ,����٬c>f��@��ms����֑���ZFc�w��>�'��x�|5�q��F'���.����a�.�%q�n��<�0���W.(��rL�A%����0
��qղiS�z�HD�>LH8�0��T<�<+Ç�+9�0ř��D�&:�� ���hTQf�o����t���<X�eC$
��0T��9x�,Qc�_6>q�*��@��$��'��$1*|�գR%��4(+��<s� �c�Z<*y�@C��3!ˇJ �@��P:Б���7�\�T����y̓<P��&�� ��V��*� \x��F�-[�	���Ԗ!�����%�t�2�>�Xy)��^(z�<�b��(P�%�S��IpO�=]�����`��v(�CSX���_%�$�d����I`H�+p%H̓t`߄I"T� '����R8��azூ���<1e-D�g���*�	��d�����I
V�R�9�H�,S��k�*);��q坟�2�u�'�%��� �]9V�Q_D�p'��p���+#���aT��Dۃs��n:xb2�Ӣ,�"��\c0�5@�4�Ç&9*Ǡ�WG�	*���
7Uj��袩�xrH��R�iy��˧I���y�b˯{��[E0��`�$��F��Eb��gf�sr U�[p��(@hE�Y/��!�f\1$N����P��U"�dc�!� ՜]��x�(�_"� ���4N�2) gGƿ�J�H��Y"9İT��i ut�a��ȟ�]�/�2A�����N
A��c��(�B\�UՊ����$o��{A����	Cu�
)�L@�F�:ӓ#;t�D}s"�%�|��g�><*�K�4^��CQ
F�)t��ІC�8F���S3�]���4(l��@�_+P��h��Z�=ohl����
����¥"�&�*�k�?�6�"(��[%bPlӭt��̡S�/%�&Dڵ �<�B/O�$�P�W�G�֝�?`q2q˷*��d�s�@�a��l������L�M9�XV���;j}*!�˵/��P���A�d��X�qC���^$*�Z�g�|}����\��-���Ġf'�Yh�O^qC�#]C�DT���OU�4�5P8�8�MDLM|��5���C�\U#��B�L ɔDV/Z]�bT(ԶU2�0��D�KFv��w�bE��폩`l��;�具G$�� ��)����Fظ"Z\ҧ������"Y'^�� ���X�����������X�AQkT�=�T�A�+�)�P���R��#�����2�Y�M3��� ���EXG��M!���s�˰�jm�bF�&d��Uha��{6�����(g�pZ6�ۆ��)�M��x̙'�]+(�ؔ�UJL$$�D�Hz�ȑ���^��,ir�,ғpu"Q��*�%��h�E9L��Ig��=��,9��+_��$�X$qv*E���ȑ&��t��P8N��]"''S���2��]�,��̓��9`Gq��((G�5�2�'w�X��n�,$�w'X#o�%@$ggjT����"~u�	�&�i����lM���DO3@�*c�8�r��@���-��^�%@��'�|�C� ��4�3���C`|ق�$Z�]u.�`D���9���D&�,JO����G@�u�CiL�@epź��ZY:�(�@ڇ�?�G'Y8}�n]����(�pvG�|�'v ���9y�~}�F�ß�8�0�G�>��kdf���4�Q�f�0��Al��韰aA���;�f�Z�'D�:�bT72�d��#�)�~	j�4^�P�҆bG�)�jlbeB٭E"����+h-r4�r/�$����/b�9���5��ʰ*T$���k4�P#)�:ą�I��z��$��[D@�P�h��&ڀ�p��4@p�5��e�^�)Bm�|��`�%�BAǈu?a���]0����bN����S@X�n�8UZp�V�}s�ٙ��������lզ�|d�ׇ^@~e!0	�-�LY�щF�~x��E}-��Ph�ǃ�yA ���k��y��_!q>���'6�U�"jx����3�_Ert�r���6)�T�	�,(�.X��
�� 1.u� �[t�>$���iWZ	7 �e��T��*�8�!@��Z��L���e�Z��gG � �h+�CV��ƀ���Ԋ|{ `0��4%7|E�`o�2X���*[2\9�+��G[���u��^��{���]�fxȕ��}ڴ���ƈ���Xs��%q�b<�'��,f�P���5fVnlZ����}߾���FH���|#%�'t�z����PQ���:M�ӌ����\B�ɘJˊ�ҎU&>x��' ���,Y�&�By��سv�ֹ@���D|��	g�Y.%�	7�܈r�$k�G[rr�]�rB��r�g��1G{��� i�
�<8��2Ԩ�$��+a��g����(A���1�,uP�'�\9RԎW��#�J��D�[�\��|K�F+�>�X+�O����]~�� #���RT �Óp^�����;!���Pg�+���d��	x�͇=�\-x��,[N\HfN�Z�`��q���BEŇdclU	��Om�0�R��``v�UX�HyPe 7�8)�`�/Ҧ��te�7���8V,OO���1��+HR�Ma#܌a���!�d�?޴���%��3����i%�����UX�T`�{ �Cq��)ΰ@�ł��0�Jf	 G�&T�ҟ̸P��1Lo>!�>))Q0A�5.�\���� ���r��E���'l89"�P�(*] a��~�e���q"�.��i��GU
(YX,JF�޲+X�2���NxR����Ţe��	�Qb�.��a��g�
)[Z �;���3�L=D�ht�Љm�t���0�ȑ���%Fz���M���O�-W�;��:@+V*f���$��qt��˱�Z,�x�2��?M��t�[�
��W�a�ԋ�o��u}&��`��ʝ����9S�P�nӬ�
��dU-q��)�T��\�����L<d 9ĕ�S�Ö��>z,��ّ�F�!CX����m���g"3|)b�5���ɒt�vN����8xu����
=8�(��7צg��S��?S��Ջ�̓�������B(mc�c
��b��3�0H~�S4s4�pR�����?E��'P!4��"EJ3d�\
.�&YB^>��SO� ��2�Ŗz�:#�b 8��O�"Ub�wST��P_(������B�1�'���r1�%a���hUJi�'��#���'g(�q�HM����;u��Er�B&S�����	�M���h[�d/�i:�47�>�'B�[D�ӎH�yö��=�p&�t�>倌�D�ET�st�����c҄�u��*CdI2U����Hg�O%�ܑjTa�&P�8(���*ڃ�ɡu�YȵY��(c����(� `U hҰ	� �.�&����ӯ7	>u��e͗X�TL
H,�R��s١F�}����Dǟ�8���1S�d�	�xBr�aa�#	��S�O!hd �J�0*(�C��3��ZT��V���K�"18wD���/FpL@�����i�!�1�;/�����)~X@1�d�t�v��O���B@���<Q������d��pWP`�$˽D��uY1�	)H<rUY�M���m���´�����'�RP9�	T�j1��f�,f�!���j�"�匫^3��J�TX!B���8�_�m�C�a�^�1Ė	���P�Q�>�"��D�m�(�±�F�MQ ��4�F^�'��TXs)��4��#m^$_:p�p7iˆ0�<��A«<���y1��5I��P��*/]H�s D�`���  �ݚ��S�4� ᧮_�CV6C���,hy:�s�*@�{��=0$��2�өE􉣟w{�uk��ք*'��r�ɪr�V���'�^<�ul�6G� ������$����!�Z�|es�����Y�+]-(�-�l�4B����� 8��t.R�>��m��,	
n��It�'��}�,j���y4샨N�lux�غ0!�+���Y��kֆ���k��ѹ����ד6�fLa�Yk��E�r��|$����M�q��`X��7�A���uU��`�H��4�dL1��F�aÆ(�dkت@V� 瀝t�<A�C��KN����"�ܥ�v���&=N,���;H*(z�)+h���JL�ӻU����w�h��VEP�R����sě;XQ�X O>�c�;�E�I�=����c�%1�u�ƦS<?��mY��ߛ=6b�IrcǦ}�ק:,/��C�'ƭ?Mh��`���di�nߚ?2�%C6 ����uV�Q���2e�Q� � �8;YЁ	 ���d��={v.�/O�  ��
%`<��0��E�����T�K�0��D*�cʌkX��N.�����R�i>Ia��D�F>�a����|��3?9����)��/Y�*��h�� �4�!��^�l�i��x�敩�Q�=��96`�$�~���l�{���#kߑ`�@r �O?���^�6X��Q�(k)�p¦(św"�Q(s �����&�O'k�J�Y�_�2T��q���	ڠd�[ 	�!��a۷I�J�ǧV�o��ضU�Ԃ�?:�|lX+�qO�	�p.�Qk\�d�M�"����G��my�F��H�,T��I�`l��� �TfF����C�O�,��!F���Q��0;F�jB�W%<� R�DY�o"02���)�(OJ�J2��':�2dD�0i2bS�J'Q6r����G/:��Ȼ�C?*�XB�#�(j��S�ȾO<���Ү$P6v�����/8������˿��d���=cD=Rd��D�Z���c����;7���2s!��?��h��g*B��#(��2nX���5_|���M0 �	1,�J�li���ؐ2���cS�d�jV�z��	���O�Z�eK�xa�h� �H0b5���P�O�@P��g&�<k��M	��<"D�ʝ|f�d� ���`3����:�<M�f8xs�4#f��13�H�o�_jp��G�N1flPa㣛�P�����S�\o���_D�^�@��,dEb=(��Y���y`Tn�2]*�
��� 7Ê���ބ@�P�`��R�"S�d�^��� Ș\=�q	`ɚ�%�����)3���#�W�'�����FLx`&!�B��Њ]�M�^1r�m�
$�y�q �.��A���T!R��ұ0�! �,��m�t"T��8�!��ӻ[��5�^�v2���cmS_���'�`���'-��YG�;%6��un�_~�M�Bks����Q��7H����YZH\�����(�(S��ӄa�%ĄY�*�q�#��E?i@���?G�TbFg�	T�Q��:a���SdH$esF���%��'*ީ+����;@�Dzf7��I�"]��[��_p�^���f^�khѤE�<G��	)7�.a�����AHS�կ���O�$"F�ч�4u��6D�N�P*��b�iX��S&M��pc�D1�,2v��0}�\w��Sᬃ� ���*�HSg𨅀��Ղ�T��0
S�~�$�XF�H�'��(�J�Ħ��W��gh�ab��\�K�2� �������_'��ٛ���0E�������^g�E`���M�6�`dX�~�响#�ⅈ'͆�ܠ8`t��M9v�?�7b^�} |� Q�{0��U�+xڐh��F.u�P�/D�
Wȹ��I7L�t�����&�H4�P��;�H���iHTHx��W3qb�B��Ë>J�'g�̈��ǟ�Z M	�	��>Mr�*�z�)��J��������Y���.3�`@�0�_8|������DӟH�R�AV+U� K��cS�L�	�d�V����Tz�MG�;�1����	v�ݨ�'Ѳ�pS	�'^���#��OB:��B+��q��^7
�`k玪M��p�~�R���2R�S7z�t�
��Tx�<bA�]�ֽB��.Y�^|��ʴ! ��e�Uʼ�O?��ń&��p���ܠ�Z�+�!�dJH�&��r�\(�nU!
�4l��5r[�ĲE�':QJ��5�a��
Ue�L�	�' 8;�i�7m��q�Ռ�-D���:�'�bm1�%^�Z��;�C��U��P�'���ZGg�0�dBX4F���'��`��8d.X�Kƾ_*�;�'a:�zvJ�@ʎy[E�E�Q�Pi�	�'�$-��nȷ�q����Nբ��	�'c���'�ޛS4�]�F���8��[	�'�j�0��	e*�eAvmV
DĜM��' �A�5n�9J�D�ҀY)U��5��'%Y;R*@5p��V�K���'5*q�Ɓ��x���.N��{�'ru����>93�+��,+ T0�'Q���dW�~V��S��$��,H�'�<D��E��1��YӢ�\�w3��[�'��X��k�L�1ė�cn�� �'w�)�.<a�Ը�VꉿQ��;�'e���@�X�%֤HUŔ:Rܨ��	�'�u�M�4<��`��ױJ�P�	�'���?rƜJR&�)Eܜ�	�'Y$�[1��$;��a�Q�X�?�xH�'� �'%�$|�q��Հ&����'���{C�:7L*�*E?�^�
��� �=sd�7]!C�C��L�e"O��K�˙�d!���UJ�
'L*��""O�1R��ث�vY��AL#0��"O.-�E�޹x.����̚='�i��"OJL��A*_9f�!�sL��W"O<	c�D"�d�kݬR�.ub"O�չt䐼X�Q��:0�iٵ9O��@a����{�[Z������8W<6�p�͏�6Ÿ�D��]"�{�CC�w��l�<%>i�a!� ]�6@�'C��% w�Z����� �J4̙;4)��M���=��(G�ƹ�0|Z�ܙ¤%: H��t��SK��M3#c�4Dm��s{h���_y�O������X���3�J�|���	���L[r���Ό�3�V���Ȏ�0|b�ӿ�bDɳ۱M�82#��F�2�c�<ڲ��ȣ!2�ͅᓤ |RXs`�¥r�MZD�����L�ŵG(X"'Θ$E�ʜ�k-����Ռ�9f��m�7=�����\�J�K�A��x�C�Y>*�a����	{�i��S��(Y7LRT�2���߆H�:���O��ᓙF�|�+��&An�@���a���=Y�0�?牠^�@5�׭d��Pg�ٶ`�jO�ñ�H�<�b���D�F�d��-P�lUBeI҉()5�Ec�(WX�
�4J�.M2�'5du���(�'����=��(����l�,Ĺ�D^,�?Ѳ�����f�[I��R
�',�jpR!�R>�d��hM�pF�����O(�[!lV�Z���	M�'���>S�ͻ��֦^\@�Z0�<,�R6 9y�T�ҬO^�ˢ*%�'�N�]Jt�͉ra�u�Д��>gx!�Tg�>y��� 0���0��OX29�B�F3O�����V|�O��s�$�0O�����h�OY07�@<�����u��	�<E�@�K�<>�P���p���)�'W��c�f�� �7lO�Tl*��geɻa14U`��M��҆�I>�M�_�E��X5Barh�d%B!p�0���?)�JW ��)�5 ���8�̀	THBEI&�.� \P�Ο�H�d#��"�O#�DcddU�+��[$mQ#[D��#B���n��s�MS��Vy ��j����f*�9p����J�i'�-��'�����^ ,N��fB�r�ϥOu*jE��JJoB�d 7�Q
	mV��'`�1���8F(&�Q��9OY����	����Z�3|��	�"O�i��O	�d̜���0T�<�"O&��7�N{9J1��m�gm.�"Oz��F+���j��*d�0Ӈ"O�@3�	uQ���;0ǂ�8P"Of�
��@OZ�T��J�´"O`���@�M��BR�+�Y��"OĈ�%h�xpi���Ă�d�"O�-�`D-��|Qf@J�^�x"O2*2��#A�̼z�	�u(i��"O�(��KƉ>RxEP�ko�a�Q"O H��N8�Ȅ�u)WsQp�Q&"O(�K��D�.���H�t�4��"O}I�o�?i/�Y˒���j�A�"OF����
Z:x��q�M�p���6"On<�u�JJ�`��R�H��$�� "O���@��Li���O]$(.t�&"O@D��l�-d��ٸ�`��?/�+�"O6�`��c2��r2��7(t��%"O��w.̉]����n��U�J�"O��9���5s����4-��f8�I
s"O,D�Մ��Qj�q�,WI�*���"OMj� *3?�㦡�M�̠{�"O�i�g�{@�%kg D�HP�"O��pAcؖ*Ұ�xRO8�&2G"O�P���
?�:��1X&f!��"O����#ަ81VA3E��0�&�
�"O���� ��8
���0�M���2%"O�c�P;>�6,����~��Y)�"O��Sff�=_�FK���@�V�2""OZP�di��
:x�8��-^N|��"O�9sfLU�l982DÃ4H���"O:�k��֕<jĔb��ǄJ߸��u"O恁���$K>�=[功�~���c"O� T�Ұ�K2C(�Q�	�e���(`"O��"�lC3	�A ��Jg.4��"Ox��&��N���@���^t5Q"O&��T�-�h|��AĝK"Vٴ"O���b�U��pӳ�ʳ	�I�"O8A2�Z<-1� ��`�5�U"O4��!�X8>��Y%ݛ%1��8�"O�M���	�� x�U;m�a"Oƅ�BџX~+
� 4	~��3"O�!��B	m��B��z�t�s"O��y�lŗ'6ت3oʄJ`F�0!"O&�����6Q�`�^XWT��"O.�+@a� 4�]�SM�:H0-�U"O��"%��6`�e���(K���"O���*�O����r��{��L��"O>�B뚹�q�q�K
j�졩c"O�RB��3����֫Fs���"O&� �Y�b����t'ىP��ə�"O����D���<��f^u{�(RE"O��	sP�/��ePr�����D"O&���*��j��l��$i��IھAc!�$��\��Eb ������m!��J:
X�<��	����b��ȯQ!�8S@��J6(ɐ@h@ �'�Ac6!�D֙lb�1�"͘�	�ry:���("!�Ď"r����f�r��i!�䊘�\9�W!:�R|��!�$l�!��Q�nYn�:�)�z���z� E�!���Jr�1�k�W�f|b��۝v�!������!�銀j���:Vn'�!�È�ʬ��X69*"N�
!��+�"�*7���<����O�2b!�dͣ_d81���V�0i:�oT�/!�D�A�@iyeKȨ1���)þ>!�d�n �NЛ 'b��d��{�!�$�='��Zg�]<�pt: 	�2�!���|�&�#�D�Zn�c�O"V�!�B�0e4��(�^Z��#���' �!�˰K��]�?X�Xf`Ǭy	!�NQ��,�)�nqR�«+�!�E�3C�H	�͌��h�ĥX�f&!򄄟c�aѠH�=.��ADT!򤋓}�
�b�E�����d��!-!�
8d۔=���#��c��S>`!��Q.���C�S�	ᜉ�$f�!�J��;��S�����`"�z"!�Q�aԄ)RC�@#�`U�W,O��!�d�<v�4]a�@�[<��p��� w�!�8$|(��
�d9б�@~!�� ¾`k� �6Z�
=#ȹ�!���!A��oL��+�/K����'�4ŋ�Ė8����f.ȭ�i�'������Y��
	F9� ��'���Y�(֕�(@��� �>!�9	�'g:���B�9�bQ�Dk5
��lx�'0`�I�-W9S�Xq���D\5��'�:�c�Q'!���� �ؔL��%p	�'Q��2��#A�(�F�ːW���r�'� "�)�T��4�T��M���	�'�v��!C��6-��b�"R�K���
�'hx|�T�jġ� �·U��A	�'�lzV���viF%����r�	�'W,�����!d[G�
pf�y�'`BP��\�W��f!�ؙJ��� ؃�"^�����K�*zjܰ"O6�{���vL�ö��
R0!�"Oԭ�) ]<Pi�f�hj���"O�C��A&i&�҅�S��ɓ�"O$�h�-�Te�ҥϢa�M��"ON�`D��=�&��t1,���"OP�g��6~.�}�b��5NJ���"O|h��l�^D 5�G�����S�"O�y�����m� �I����"O|�a5����6�s]H�"On��֤y���vf�,m���%"O
5I��]2E |B�ޔ+Vnl�W"O�,p����S� ��a۞_>��@�"O�U�N����Q�A+d0�e�3"O�斑q7jxtA�~wH{�"O�u9u��3���A�@I��c"O�1H&��c& ����97�2��"Oڸ!��X���!��+u�!��"Oʵ�t�ەN�=B��P:>�R"O A����42�u2��Q-$10��"O��@�	�vY�P ��R6|�a@�"O^���T-M~����,ͮ8�v�C"O�5�`dGN8t �޷TC����"OBlB��� �\H�a�ɡ+MvԳ"O ����8+�H��bgǁ疴I�"O���˴f��Բ��	�.��"O���gX%7�"|����>��ՉW"Or1���M�ԜxF O"&{���%"O��C���Yd������$�$�g"Oy1 %w���Q�-�"WR�Ra"OBa��;h��ip'׏pLx`�"O0U��&˩;Fܲ#�B�>/��D"OB��L�z�8pe-P�}z���"O$hҗ�	���uaDQ�z��!�d"O4�Q�-��Q�X}h��ԉ*^ܨ��"O@���ҫn���eޒ%�|�Y%"O��;��N�r�Nɨ ��t��ɲ""O�PB����M*���%�"%�G�,D����^�5���C��?�(����)D�pJ3�ՒX�xH�Ȑ4��}ï)D��"���=d(P]���Y/V��U�&D�X!牨O*$�j��D�*ef�!��"���%l�$Ŷ}S�Ա!�Ĝ�sx ��5�xE�7� 6�!��7$������>{(�PX�!��Ћj���Ì�9,q�h��L��!��,���� ��	�2�z��J�K�!�dE?8�r-�Ť�6e��a#P!̀8�!��/	��`��P �m�3aD
"�!�Q8Ȟ��^>�j�O?Ne!���N����c���p𰤘
(�!�d�>t�`jg�739�y�lF�|�!�$�S��@��!N
G�y3P��0e�!�X><8�YL�9)2�C�)N6D�!�D\6�Z�
��N�c������$f�!��z( IQ,�b�5�/�Xo!���� 	� Ǉ�b�8�Q�d�!�Dͳ���+����DN*c�!�Éy�~��oX%:��Q�N# �!�Dŕ^~T��blV�;����� ւ0!򤐒A����FZ�i�R���`�7 !�>v��d�/�~L{���-O�!�D�6��Z�GPU��+�م^�!�$ۗ(в����H�ShD���>!�� � `�
VT��Ա��RZ�έҷ"O1!�4�dL)��I���DB"OF0h���9Ѻ��q���,�r9˖"O��HWA��~�ܸc 92�(�"O
�:��*<,AS*�7����w"O �j"`W[�Kթ�AP5y�"O`�ڳ���R��]
��� X�֔�'"O���e�o��)�RƞS{PA"O�,xQ	K|���AO�:gvtp�"O�y*���9�|5��"dm���1"OV�I��� k�X���P�R^�A`"O�T"�cе4��#��� /N���$"O��iٗ"����"�ɓG.�M�w"O��f��^Jx���@�&����"O.�����>0�92������"O@90v�֑[p��,|�\A�"O�8dD[�T�p7Q�)#P�3W�2D�Pq�@�I�V�B�l
�-jz �o2D�8ʤ��c�T��aL?F�@Dc�'$D���k�N��� %j�  ���/D���bف$�
�K	"D�hZ�.D�`E	K�c@v�����V�bp�*D�p�r���W�hu8���nQ��/)D�0ku�W��e��iQ�?�VM�S�:D��d��"�9����B�@E� �5D���%�5r�� �.4)�q���2D�8�2�+)l�l�����Pݰ�d3D������$sC������'s���0D�Цg�Yp�!�R�;�dP`�G4D� j��m�H��AK���|���3D���F�0�Z*��9�b�L3D��I��N�G(Q�蜾���E�1D�l�G�l@б�aY�I�qǇ+D��� ��WD^�wGٕ){�T!�i+D�T��
¿9� U0�F� ���)D��rs$˩b�2��R���E/(D��Z�   ��   �  ?  �  k  �)  �4  @  �J  V  �a  �l  �w  ��  #�  Y�  ��   �  O�  ��  �  %�  {�  ��  ;�  ��  �  ��  ��  ^�  ��  ��  ?�  � � > � �% =- k4 U> cF �L -S pY p[  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�$n�18�srʙ�2�<I: *�E�+n���D�O�H�'Zb'O�I$�	�5Kւ=U�`�aC>6�'�$�b��i��I�|���O(�j߸��t�ޫc��A��D����<I�����3�'^x��k��=�X5`\ u���aD�i�ҽz�y��I�O��L��y�bnV�(�BY��/��y����OL�	E}���b��^A��1OT0:��"*�x�ѡ�Ɂu�6�k�5Ox牘�?Q�N#��|Z��j�NlI��y�,�F�.c6BH����;�Ϧ-�a@1�	�q���й8)4�k4*��,~�U�?�*O���O���V}R�������wI��'~����
-��d�O��Q	ߕZ�1����Z�h��Ǧ殜pn� 6�@�%I�:�|����O?�I$4�wkO�k���׆G�O�d���
!?�������.��EC
|�	�
^dа%I��y2�'Q��'�����i����|RB�O;Q�'g��w�`	����~�2x�6�Te�I]y�O:B�'i��'�r�h�6*�E�k�4��Dc��I�M[ա����$�O��?a��B\AT�����	z�H�ʳ�VyR�'��O1�|�je�."�^q��4�=K^���
��<��~?>��:����U*b	8Q�w��	_�Tb�Fw^����O(��O��4�������̚/��N�C���X�ʁ�{�F�£f@��y��'��O��?Q��?	�B���Ą�$�sB��G��"�
�4���$Dܡ��'��O��ߡ[�lpr��<g�RxY3)��y2�'	�'���'���iW+pn����!��fȓ�0|˓�?���i���ȟ��$:�d�d4@�;�[�L���;V[�/�O
��O�	O�{�07�0?Q #�&�> ��"� p�R@�0��Rl��4$�d�'"��5�4�?�E�)�N%��Ȱ��`ם�?!���d�ɦճ㢇џX���O]L��3��:A54,���,����O���?�����S��J��(yQb�f0Is����D��A�=c�X�O�I���?Y�j#�dȺ@�x�	 �ƞm�|t2�a��1��d�OT���O��i�<�s�i����%�?4���-�N��ra���YV�Ɵ0�?�.O,�d��t�eZ1ZTV�tm26#�˓&&
�a�4���J�`Q����Bצ˓	��u�4G�	f4Q��Ki�6����d�O��D�Ot�D�O��d�|BD� p����&K�}+�
��\(��@3V���'-"���'��wq,�E��:Ok�%��V����'�2�|����
�_3Ob���! \��)!/�i��9��3O� b�؂�?���;��<ͧ�?�A&M�&ŀ!�θ\iJad���?���?�����Ĝ��*2O���$����XR5%A�tG�@����9~f�ǈe���$�O`��=�dƫv}���R*$�<D���[�I�0`H���O��k%xb>�÷�'/x��I�;�ص(�뜽���z&��L
���؟8����\��\�O<��U3x�r �@��6V�;���sr�bӒ�i�&�O����O����!�m�tD��)k�|����$qr��Οl�I�0+ ʃ殮�'�0�8u�C]z�.ڲx�$8�	�T" ��g#������O:��O�d�O�dV?s�*)�pEX�<7*�	ÆBuR<�ye�V�T�6��'������',z��)]4�����&���^�P�I�L$�b>I�g�Ǉ9�X�٢��$Vļ#�F�5F P�ú�˓vd����OL-�K>.O Q�I�<	T%Z4�P�~�ŀ�!�O��$�O*��O�<)U�i�eڀ�'K:�ɣ�_�ex����U;}�v!��'q��$�<����?��LI��F��&�*����K�P�wk�8�M��O,�2���(�4�� ���O��C����Q �"�;�0O����Of���O����O��?�xӡI�9�|�$���^�����ϟ��	՟x��4p\��'�?����->�)5BH!'qƥ 0����P)�<!������&P�6�)?��"EK��t;p&�	6����o��Qפ���O�O��(I>�,OH���O���OȽ��*�PT��A�͹y�ِ���OD�$�<���i�0i[�'dB�'���W���%�N��(�1�����O��d=��?��0�G�n�8|�Si��-`t�9����z�k%mA?���|
���O*1zH>�C�EI�c�M�aHN��� Է�?!��?��?�|�.O��nڝ���2b�*y��� P���bj��\�I��?i*O.�D�F���� $0����B	y��G�\���4����6�Ը!����ʓ7�@�����PB0a	������d�O��D�O���O��$�|�񭜸�8�x������dΚ����S��B�'�"��T�'W�w�Ll��]�'rp�+��V�zzDL��'���|����A�d*��5O�}�$!ڐy�� 5��f�t�@2O�9����?1�+�d�<�'�?�v��)�� ��JO�$���zD�?����?����d��%���DٟL�I��z���P�b��F��7rNi�K�m����ON��;�dY)Xpk�d+c�,)�u+ϐuh��&V���ʦ=L~�ui��(�I����K]�E��u�`�>h"��I���I����IM�O)�ձ$�ش���]�p=Iu�݇q`�h��@ٷk�O����O����5��8�N��p�`�2N7T�����x�	̟�3$�̦M�'1�\�4-�?���ܨP٘�2gC�}�Ri��b
��'��i>��	П���ǟ�I46oP�u"�sJ
&KM1�ʉ�'[�7��Kk��d�O��D-��#�� `��>/��YU��*���':��'ɧ�Ov�A�RFD:`������Q�����蟀e6D�;^�tZ�M�~��Tj�Igy2��8мqpDҋO&��p� �u"�'�'U�O�I�M�d��:�?�����(g�a16cN�]�4*��R��?�����']��Ɵ��Iܟ$�Si��Ay��WQ�f��TB�� r�xl�@~B	Y�.��D��\ܧ��!��C@�� ���5ks@`���<1���?����?����?9��dI��cP\KD
�_0���èɜ
�"�'�" {� D�B1�&���O �OT0��D X#����Udx`S�%���Ox�4�,��$z�X�ӺÅa�.I�ڈ9$)�Ja6]R�eJ |XF���F���ONʓ�?1��?��(��mH�$^7+��)�t(ȪF�����?�+Oz�n�'�4@��ܟL�Ia�$�	Ġy��� ��\
u#/��d�<���?YH>�O�����H�8A�bR�`FI��!�9py\�QwJ
�g�i>�a��'N�$��#�H(8�Fɓ�a��>!<C`�ݟ��I�����b>��'u�6m)�"۰G>!�|���.�RH�ல<�����'����@��HP���xq��@^��"gdy�\4y����� EH�b���Oyr�߂�Ă$G�,sQ
McreE�yBZ�@�	ПX���L��џؕO'≰ �4p����� u�6tr�{��5����O��$�OD���D�O�n
(�`�����=��M�2+&�6�)��8��	n�<a�A��t�,-�n�;��\�g��<A'�"'��d�5����$�O���)qN�"�%�c�:,�զ{���D�O���OV�E��&���B��'r��)/Ð��Z9i�b�xK۝N��O�ʓ�?���� �L�Z#�ǧU�@�h�Ă�'�4h�V�B�(��-)����ϟ)�'��X8���)KwY�%�Ӏ#�z$���'���'��'��>��ɖ>A�P�BD�8
x�gM��L��\�I��M����d�OH��] "��DB5E̩L��	q�C$d@�I���I۟0z�
�֦��'oB��P(Y�?j2��༒Y�@)0@)�^��$I>)(O�	�O����O*�d�Op����	+h�< f�C`����<q��iC.ة@�'�R�'��O����&B6�����<g��D��.	Dx�I����?�|����hsX��3��?x	H�G/�����Q4'���$�'"R��V�OZ�-�f{����&��� -�$���Lҟ��	ޟ���՟�Wy��n�\�P��OܱY6�1R)�⧢1	
^m;���O��-�	dyR�'o��'@��1g�5F�*6��hP��S*܇/����Hc�Db�čc�S��IsG��ఽ�an�-F	�0�l�������ٟ��Iӟh���D��U�r����C�%;r�Z��V��?I��?�s�iÜ���W�`��^�	.U.\! /�!��)1�E�v�&�(�I���Ӻ~�&lo�j~�KU������&!��M���]0�*���Ο@r�|�^����,�I���S�ȇdJ��G�؅�ZM�蟔�IZy2Bb��tj���O��d�O*ʧ U��"���1\����
X$28H`�'x�	���	k�)�0BR�^LKת��oj�
�N�
#LE@Z�[��������K�|B�$ iC���9�J)h�r�'�B�'����Z��b�4^Ƽ�p2��;ua �����^��<��⚎���Ov�T�'P2�O����3�=]`���fW�iC�' �8���i[�	�.����r�� ��a�E��-x(@�l+h,�M�<O���?q���?���?����iS'_��A�Κ�3þ�	kU��V�n�;��Q�'�2�i�O���(|N��I�O0�0��@L+W�|�$�O�O1�f��A`���I"J�.,�I� [����F�e3F�I�*��H�u�'e�%�X����'n0! � �:��Ip�ozZX��'"�'��S�����6ޘ��ϟ\�	.w�X�u��,������;"�H��?q)O,�D�O�O�p�A�S,w���r��/���:c��l#@�J;����&RH�<r&ڟ��槗��29�h��'�Q���ݟ��Iן��	ҟ�E���'��P����Դ��]��v�'z67-��x�^˓�?ɋ�w�a0�N�[����5EL3]:8�'B�'W�+ne����T�I�Ą�/��+ ��L4��vH��e���&�Ԕ��4�'���'�b�'-2����I��P\P��
�C�)��P��#شT�^J��?9���䧄?c�����2��IrO���&�@�����O��:���7AЈ="�`�>�M�"@�'~PV�`��t�Ԍ�'<��r?QI>�)O:�KՆ�B��7�F�M5NP�4��O�d�ON���O�)�<��i|~u���'5��Eኩ%�~��`lF�j'��
F�'����<1���?��+�Y����1W���$�3���j�'	�M�O�0�+ˆ�(����Y!ZI�قF�@�v�$��a�/6����O"�D�O����O���'���l�Z��_�L���i6��q1f��I� �ɒ�MC��|"���?J>�"iæ�VT&혟 �����EB���?���|
b��#�M��O�.Ȧ^�(SI\58iX�!�,	>N�vEAE�O�U�I>I-Op���O���O��*�U06�I�EG"�
W�O@���<	�i��	%�'�B�'���M~�e�F5n�*��N�!#����O��D ��?5{r��k�ԉ�G�Sf�&���,ڳ'W%F�y����|�$��O��cI>�C��2�
$9SA�.\ؘ%�B�_��?q��?��?�|z/O�`nڻf��e�P�H�	l���9%�L�$h_Gy��'��O˓�?AQ؛R�^��N���k��#���Q��6�4?!5(<u�~������J�V��t#Î��y#�ꛩ"�$�<Q���?Y���?���?�/������.� �Q�ԃ}|�8����u8C%����՟@'?�I��h�jw��H�F�Vn�_�����l%�b>���ڦ��H�D	�e���Pdr��M�͓]F�)�h��@$�������'�T)�F��2�Z�C�v��A�'���'��T��޴-E��P,O>�D%o&�SS�O
#$�Pʲ�
�a"�T�'���L"�:��	^,���i�	тXw�I�X:��h�]�� �$?�x��'� ��ɫp��D���
jJ�E{p��D=���I���I䟴��{�O���T5R�%9��Q(.	��P�͚%��&}Ӵ�A�E�O��$�O���]4$�ar��F��@t��}���	���IşLb5��'��0f�aZ4+�$x��=o˅�"�I��)����4�B���O����O����%���!�Z�k�����/ȷ��˓r՛�@�E�'�B��4�'�x�@��IO�pWl��Ȍ�]�<�IQ�ŞV(b�`�*�/^h}QFlG;lP�w���3�� �(O�@�_�?	��+�d�<�tj�/�t�X�'��@qҘ��i��?����?���?ͧ���Tצy �@�(A���bh�ҕ��	g��37�ҟ���n����O��4��Tc�1��i�@-b�%aD�� ^�7�2?����
8"�SQ���E۷�K�YnB�M�+��(�hx�P�	����	��4��ҟ����פS�H2�lX0N�9A���?��?9��iH�W���	k�d�����'�!�̳�m�6�\�%�������Ӥm��m�A~�&�9b:n�+5r�� t?}L8�����8Q3�|�R���؟���Ο����G>` ʤ`�nB�= EH�ş��Ily�qӾi���On���Oʧ6�A	Sǈ<zф��S�Z�hh�'4�	��T�IZ�)*&�MW�����ԸY����
b"���T I�Z���� 埜"$�| @�[:�5�C��2��eb�K-|��'.�'���tZ��h�4J썊C�JOJ�٨�܃:�
Q�E����?���?��Y�h��6g֊GkK�%9ǎb0(ɖ'�0 f�i���j�x|���O�(��'�l�q�Œ_�BL��(W�vND]�'��I�����������C��C�%|�@�a��P
�Y�f�O�	�6��9�(��O���&�i�O�4� m��Kӣ(����i�x�y���O���*���B��7k��3/p�� ��>��!�a	S��y�m�b*���������O~�ƢPlad�Ѯ^v%W�!M���$�O��$�O�ʓ<w�&�ޓ/���'zr��W7b�ـc��X��q�^<]��O˓�?��T��(�D J�L�5��Ξ���� �c��P�&�c�0���X��a���DY
=���'�Я�ة��2�6���O����O��d?�'�?�G�J�)��X�s�#}�d�y�'ڜ�?	S�ix�y�_����X�Ӽ;�%Ϡ;�Z�a���eS�u�PB�<���?�o����4��Dؔc]0���π ���qI_�66�� � Z9@k��;�ı<ͧ�?����?���?�u�ͽXrj�����0n��g����d�Ħ�J" ��(�I��%?��5=h�G,ش_>���ß�I�ܖ'R�'�ɧ�OŖ;$��K�t�k%�۾cT��ɷ[�>�X��O�	�oA6�?�O<��<1v)��%��va�'g�,��!�ǘ�?���?����?�'��$�J�A��\jU�yG�e8�iޡ3N�0�n��?a����'����t�	埬3Վ&%R�c

:B�t��/	�C�2�m�S~���$�H��Ӌ��O�7B�= ;�2�L[�w����2*ؖ�y��'�2�'���'}2�������8�K�H��� ��>#<r���O���Ʀ)��g>Q���8'�ؕJ	u���+�e��N_R�R��$����'v8��i��ɀ]�4i�J�+ M~-�န�)&9�FeP�g���P�IRy2�'2�'|r��6:{*���l��Hׄ|�f�S k:��'��	�Ms@�_�?���?�(���3�T�A��ԧG�в�ᜟ �'y��'�ɧ�	��{�JTjAGʀ �|�Al�$xje�EOGHX�'�<�'s2�$���&Kĕ��iܗV�t�r�B�3��;���?���?��S�'���٦�针߱r��1;I֎e\D�Y����[���I���	Z���D�O��ZG V����7d��.��-A�F�O��ğ�7m<?��EЪj1��>9��⁘e�j|��$�%9c���d�p���'���'��'���'f�<L���C�M@��K,>�s�4g�>�Q��?�����'�?��Ӽ�r� ^���Y[c8]A����?����Ş=�t�ٴ�y�ń�Fm�!���*����$�y�A
rwz��I8�'u�IΟ4�I�?P���_�8k�E���|$�����IП �'��6m�&1����O���4:u�xMڝW��0Z6M�n�"⟠�'("�'M�'j�ACH�"� ����b�|[�O�APs!R*n66�%��&T��d�O:Eqw�����ks�D�{��ڔ��O���O,�d�O^�}��� -Ӄ��^g��� �_NX��#�V%B�Q�I��(�?ͻT
�KLЛuD��Xe#7gA�@Γ�?Y���?�����M�OD�(�-��zsL#]���܅�v�˰�f�F�O|��|���?���?Q��M�9���B�I^��Ef�E/Xj*O2�m	�: ��ӟ|��J�s��)[�J���+ �!�L�р��py��'tb�|��4�@TWT@�@�͞>�pEd]�z�\���B�����Ⱥl�$��hJ�O.����� H
3���*W��~��T���?���?9��|�*O<�oڕV�����w�0�:dBT3.��$Ț
,ȉ��ݟ�?�-Or�d�OT�d=D�:��� ^17NDG ؓ>�xM��.|���`O� #Q����>��ݣ>|�ڶIE<v�@��J��*zb��쟰�����	䟸��{��M�h�w�S�C
��i���#CT�
���?Y��z$�&c��S��џ�'�4�5f�$T\���g�V�{��	U�Rr�IԟL�i>��Cf�I�'�r͘vC�2e��=H�!�H��x�.W�0'<�I�D�'#�i>��������_p�l $/[0R*�1g��B^\�	ןԗ'R7mD*\����O�$�|B� ��+m=�G	T�ْVb�C~V�H�	T%��'R��Ѫ֭X*��;UCuU����T0H����AŨ����|����O2M>���E�v�P"��ȥZ��X�L8�?���?9���?�|�/O��m�M	�Ȳ��ϔ)o"=�B�36S� 	�B�my"�'��O���?�2C�?"�3�!2v�A��T�?�N�\�ش����%���A�)O�P��dB_�T{��P�v��0�?O,��?��?��?�����i� nl� �iL���T�J�D���nژ_�2,��ן`�IP�ןP�i�혵��2,�e�ŗR�j��s��ޟ,��r�)��Y�(�m��<�b��$s���PJ�C>��f�H�<9W��S ���B*����4�����_(�4͐3!6� ��b�.u �d�OR���O�˓�֮ĒGB�'�BcA��쳥,Ы&��-X�C	0�O�˓�?Q���M����	�>,�P��䣞�ג��'Y�`Ռ/��6��X��~��'����5��2ޜu	�� ���i�'��'1��'��>�������j��ۊU13SL����I��M֍V���D�O&��|PX�!�Ҝ8P2<���Fe����L���H"���릡�'�����d��?iy��΢!���1AQ}�t�裀�5}��'��i>���ן���џD�I�
�|�y6� ��m���A���'/�6m�(���O��#�9O$̒6@ X��Ҥ�)T����K�<����?�J>�|t��# �y�ף��.�)I3��`_�@![n~�f·#мL���\��'��� 	�`1�����Am��*w��J��8�	ğl�I����i>�'��7m�MO����B�dI���=5��x�t�6H\�$�O���'���ygϙ�~�堅���mD\��P�C��0�B��i��ɕ_~�c�O3h�$?���"E�0�ҹQ�|��&o��n��I��	� �I�����~�'4�VؙF�֡ ��50�EZ>N,��R���?i�8r�F`��^h�I���%��z�o�<d~H���21b������o�	�$�i>��r�ڛ����z�j4� �H���l�$�
�)�2�:E�R)˔�?��m"��<ͧ�?	��?�0X\�4��#�M�>�e��?Q���ܦ�Y������L�O嘑�`Y�z:�P�j�r�����O�˓�?)���S����[3~L���R�w;)����,�E���b	.�C�O�Z��?i�H'�� 1-=Fe�N՜Fl̨*@�	R�����O���O���i�<���i(fQ��!��x��3�n��%������'���'��O���?ч*�5|��\R�N��":L+7f
�?��pr�P�4����r\���Xk-OL��p _���yk��q�F�Ŀ<���?9��?���?I.����,�ը3�M9wG�
��������ß<$?�����ݤ�D���3}��<��nx	lM��ڟ8'�b>a�0��Eϓ-n* A�AB�7� �B��Y�O��Γt�t�s���X'��'��'	V(X�'L<ZD�t��!PT2���'C2�'LP��iڴ`2UB���?���y�lb���Up�q4�"Ƽ����_�0��R��X�1Z���-|����'�$U����'�L9s�m@�E#4��2��t- ⟀���'J�
e�54&����0)�,�J��'l�'���'$�>y̓]m�,J!��;h�t9zUȋ(a�u�	��M{�`�.���Ov��]=@�3R"_�$f�= $.�"0��џD�Ißxa�����u�+�'1���T�S<f�pR����D�~�<1&���'�B�'�'���'  ���E�:�y e	�tU�P�cR����4e׆�����?����䧐?�g �w�0�#��,z����D�O���9���(D�03�(fȼ�!�bj�R��}��%�'nhRsi�S?J>�,O]�D`S:.��d����6S�4�T��O��$�O����O�<�ǽi�.ܢa�'�h�bd䈼�ʱpDA� 2�؂ �'�"�d�<���?ͻ\�Uڥ���M�3 �H*`�Ī�Mk�OJ yB�U:���D*��wޡ�$�P�;��C@F�q�B��<1��?y��?����?!��TA
1E��)C�ʌ0{z1��c֒s�'��$rӦsf>�@��O��OZ�C�}(���ԇ��
�~���Hܚ�䓺?���|����"�M��OX9)U�.}N���ƊB�j��Fں������uj��O���|2��?����.p�P�?��u3� \耄Z���?a*Ooڽ$ ���ӟ4��n�$�Z29DT���:mM�X�⧈,���<���?aJ>�O���Iga�="��A0̅*3��!����t.(���io�i>��$�O��OrYТ(��g� LO������On�$�O����O1��ʓD:��@	�g,$0��7)�$S2�;d��`�PV���It�����O�0 �(%oεp�G�q��@C�M�O��䁈#!b7m>?�B��y,��)=�'�y��Z��"5�>��I��yB[��I����柈���P�O��Y����B��r��5G�(I(��t�r4x�A�O@�d�O���F���O��ݿ*0E8�cϭCG��֧]	)��d�O�O1���Q�o��牝l��Xy��uX`恘� ���ɕW�ڝ��O��O���?�8]q��_�U����	0Z�V0)��?����?,O��n�b����៸��2�L����:%�0z����-�?�.O&�d-�ɽNMı��B�=�
�+1��f�{�0Α�#tQ�M~R!n�O~Q���<_F��R�5gk��;hF$`��̅�%Br8��π	@�*��oR��91��qԛi��|�b�'��4�}06CZu�H�C���8Mp�I�4O$���O��dR>6�*?aC"Fh��?�ܪ�aո'��E�v��=9� �&�T�'�џ��V�߈&������5/�:Z��!?9$�i/�� X���Io�'^F�!�dVB�ɳ�Ԃh��t�+O����O��O1�� �gG�I�`dc��S;h�Α+Ѯ�7�P�˴
�<)G�O�r�B�dҪ����ď�b��R���z�����a|҈bӬ�b M�Ozt	��-	h��k٧8��!q�;OP��7�	zy��'���'�tL����Q7�ā5\( ���*ՈYw̛V���+��>���@�_���ъ�nߝ#X>M"����7�L`�C�o�؅�	�D|2�����8f�n���MU#"̤��ϟ��ɧ�M���Y�4�'��'d�����܂{�d�e
�?�:)�b�|b�'��O���i��Ij�+�!��c�];�.l�s&�����'��'��i�)h�R͖�FXj,J�g�TM�Gx�)lӄ b���O���OV˧Ww ����X(QPF	U0jf�'q�	ȟ���z�):sK���Vݚ���&M�.�!�3�$8s���M�']�擟��d3��D$����G�>�4�BӣD�]!�B������!)��u�1(�y�x8��! ��'���D�<!���*�Ӗ��b�(դ܈������?�dh�M#�O��`���݈��D��M��R��!�ǔXizE0Oʓ�?����?Y���?����iL?x\I"AFn�*�*E��l&ؔ'���I�O���9u�f�I��i�IY1D�*R���d"�)擽!��nZ�<� Zq���U?H4��p����Ua6O\A�dB��?��i1��<Q��?ip(08z��R�,۶~x��W)Ք�?���?�����d�զq3I�����	ş��o޸:�80;����tT�W��|����d�O�⟄j���5��%�$ �	W��͓��6?A@�A��9S#�ٴ��E���D�4�?��]O,��Ǆ�2P�	;S�-�?i��?���?!����O��SJ�; t�壓0P��j�Oo�[�~d�	ß���B�Ӽ���4/��3��
D�0�q#`[�<A������v��6m!?I�˕2 ��)�	B�L��z�-�Bͳd �,�cI+�$�<����?9��?���?�I��eѪ���̄d�XRDM���U��5�GƐ��	�h&?�	 �H�V��9*�Ѐ	�+�T�zЗ'&��ɁdY�-:�@{��� �9+n��p���"Q���D����6c�ONe
H>�.O2͐1#�z�(�b(�*R؉r@�O:�$�O��$�O�ɡ<'�ii�)��'�*1RW,�2�#؂�X�1�'��Ĺ<����D�6�fP9u�,�ZaBg���5�S� �^7(?y�'��6�I�	�䧉���,4���<>^�I���<���?���?���?���T�� *�QxS�ӣ �L�q��E�4���'�Jq��(Ȇ��<)���qD��K��2�M��mɧ|9H>����?�'6�����4��$@)Q,�sw&� $��X�64�yH�g��?� "�D�<�'�?����?1U�I�9j��f�
]a0C�o]�?1����[��9�'�ɟ���ퟨ�O�
D�A� �\���f$d���p�O�ʓ�?����S��J ���Ự��x����C�8���a!� %~i��O�i ��?� %/�$�J�
ar���H�b造���	�����O����O���<	��i����	S-� �)dLA�_ϬL)s�:��,�?Q.O�DY��0F�W�'��ke��xYt���O���q�b���/%,�AE@�N�O�~���ք��a�[�Xi^ [�'�	����I�<�	���IU�$您i�p�ڐ�R&6B����
Rv6�3T��?q����y�(_;jìl����0o�{�Ʌ�2�''ɧ�Oa�Y���iw�I5�RA�a��W6`%q��[�r�'� !0�&��Z�|�V���ǟ0�TOG��:�Zs-�h�:�(���|��柀�I@y��c�tq�a�O���O�Ÿ�Z&N�:�Ǭ* �ළ?�	Py�'Gb�|r �)���FQ�t�M�����$��(�qe�ߍ"E1�u8��'E����/ $��d"����$�G��_=l���O��D�O��$;�'�?	A�]�(َu��f�'jX�C�e،�?!S�i�4��ݟ��I����?�;M`mXb���2*�r�f�-�l�̓�?)��?�M	�M��O����
/�ҵ�]
�!�)ՉHiР1!��qړO���|����?����?��z��q3+�;����%NJ/�*O<|nښb@D��П��IK�П��بb�tɪC$ĜD�t]�A�Ky"�'3R�|��t�٠e�1A2�{b\� ��
A�&��U�i/�ʓ07��'I���$��'>�Z�(Դ;�,	u蟒8�ũU�'�r�'�����dY����4	g$����x��p;v�9Sj����?)�b]���	�8�I�B��9 �g��Ƕ�3�߈[�T��m��Q�'"nRՏ�o�M~z�;K
�0U��I�t37��:�*IΓ�?����?����?�����Oe�IZ$��v.,�3�!!0e1�'�"�''z6-� ��i�O���%��D� ,@�#N;�Zd��,!RhH�O��$�O�
�fn�7�6?9�)-�d��� ��V!3tF�5�]AR ��H%�8�'SB�'/��'v�	�D��R����>�z��!�'��Z�\��4l�i��?�����_gP�R�F֒rWzq�.�7N�D�Oʓ�?����S����}z�d�փ3]b����Z=�����E�G���-�<�''#,�	F�I2!ښmrֈ�d���kZEk���������؟�)�Iy��m�����Ojg� Qr/D�P�P�W-C�}�����O8��-���OZʓ�?����a֔ڕ�ς$*�m3�M��?Q��%��q�4��dE��^a��O��	;��z��Ɨ�E	Z�<�١:Or˓�?Q��?����?���򉆦���C�����0(ÔG�n�;k���I��T�	N�ß��iށpd�ͅ/:�	Q�*@�xۗ�
؟\�	p�)�ӈ�0�m��<!F(ۢ/g�R��92��s �<�rfH(���IL�	Uy�'����
)��1�wo�U�,	���)}��'���']�	<�MS���?���?�a�:r�(�n�<�(��ƨ҂�䓍?q+O����O2�O�!ІjM a�I��#�.0�|hJ���<����-H��]�4�d��)I���C��T�lW�-a��!eB��:6�@����П��	�@G��w����פ�!}"�|� O
��Y�'{b6M�}���Oz��/���O�����&�C"&�,tB�����O����O��a&�{�r�Ӻ�BT��J�-E�^��V&F�M��%�P����O�˓�?i���?���?��/�X��t@Rf�t��A��Z�fI�(O�oZ�A1����ƟH�	p�ğ��Td��h&��G�Q+<X���u"Wuy�'��|����A��� ������0̔H)&��f�~H�Щx�5�'�04J�b�D?!J>Y)O���G^Oz���IǾ=\�i1b�O��d�O2��O��<Iq�i��9��'�P�x�k�.�������� f�' �|��'����h�i��ON�b���*��q�tp���I�{� �mZj~���>'�l�������3����caD�{�.]�#$����@�<1���?	��?��?I��D"
6d��p�ņ� y�@޸ 2�'2"�u��8�2�R���O�Oĩ�%�Gz�
9� �n�LYҗ <��O��4��qe���Ӻ'���D���c��s�ܜ��˃�)NAr�c��OB��?)���?Q��n�J��Tв$#��:g�A�v�0(P��?�(O�An�2FbT�'�r^>�IdnQ�LH�5Α1�9{#.!?	)O\�D�O��O�Ӊd=-���MsLic�?6֙H���
"���nڛ��4�r��'R�'-���	��e�: ���pX@���'�b�'��OH�I�M�F/�����bI�>;��X�dݛZhT(���?�����':�I���)�dG�+"����"0#T�QlL̟��	�L��l�Z~�(��������
(ζ)"b�&+�´�c�λor�<��?!���?���?q)��( b��n�T��D������"�ʦ�(�+����I֟�%?��I��1JL�!�]�e�*�'�+����ԟ|&�b>����Ǧ�Γ&kD�:���&u��@��Bӟqy���Yxm����&���'�"�'f�����t��A���҇A\f}{��'g��'�"P�\Aݴl~f����?��,�
HٶgI�d�맊cdL��bP�l��ݟ�'�H�S�7[� -iPi��ZGt`d(?QҠڪ~�I�4��O�����?	�� 0w"P	�E�	�x00�7��?����?���?���	�O"�;���9�=� �F T�*��6��OR1l#*rB����D��k�Ӽ�@� w|.��!��\�$�2(A�<q���?��:�U+ݴ��D��	�j�O� ��*�<2�g��}� H��|�W�x�I���͟��I��4�ԃЄY���q�+�ӲE��dy�Dp��ex�m�O,���O�����ɾl��R�Q�305��!�/B�˓�?����S�'Q�aA��ǡ~\����n�py@�%���n��'�ԡ��G͟� ǟ|�W�� ��8� �F�¹17^ɟ ���D��̟�SDyt�V���O�4z�h������fފ1�4O���/��ey�'E�'��[��C�2�6I*b9�q[�H,Y�������hE�|��4�)��\������?e
@z6�C�H����$K?3��S'�q�T�+�H�r�$����1c]z����F�\����`&@)TF�²*��d�����\�q���."�Z(�&�"�0�T#��c30t
3�
��'2|s铮w��kȐKB�y�b����G�X�L�Tyе��=>���㖤c�����˗W'A9S`��V��[ōx�*�JbcM4 I"�%��-���a�/��.��cѧĳB�R�0�l�Zl��`J:arLˤ������T*� �٘�*�:\�PQ�L�0Iԛ��'7��'j���>�)O��$��P�B��=B1f�Y�(�$�CТw�N�O��z��Do�S�����ğ�itɃ%�t�k���*J$j�����M���O�N�sY���'�|Zcbz#�JP:��d��J�!�O�����O�ʓ�?���?�+OBЫ����8�R-���	8\8Rc(H�	(�'I�	��$���I�
a�Y�d�wl�e�� ^�T*�b���	͟��	vy��̀x�T��N�$���7qG��rT�AM7m�<1����?9��cJ��@�'�n����
Ap����&���N0�O6��O����<Y&ɏm��Sҟ���P�v���t�G?Sր�r�,�MC����?I��)�}����I�i�>��pgA�n^*�"�T��6��O���<q��4��֟���S��IM� 6J����!(�,9pa/�`�	�\���M"Z��?��O�Ԍ���X�B�얰Vծ�H�4��
`��n�ǟ��IʟԔ�yZcD0H��'"f*a��S�BzƵ ޴�?���f�83��	�j���c2��"��%�!�e�F א}��7M�ON�D�O��I�|}"R��C�̎$g�-��^(Wec0�Յ�M���(��'��N�D�3x_�}2h�Y�qZ��4���o���I� �b�ҏ��D�<I��~B+ :n����ӧܴEb`�ف�MsH>y���%�O�R�'@��N9^�H�1@�Z�U�Fh
�Ƈ
ux7��OH��J	H}�Q���IZ�i�au��"���CB�G7v�V�؀d�>9wI���䓂?q���?�,O~�J!_[ ��1��̂'ʄ�X��W"h%� ��՟H$���uW��O��.bF��5�&�M+���D�O�d�O��l1���3�D��� u��!&+]�M�|e�2\���	�`&�����T�'؈:୉+,X�R�����E,�>1���?	�����G�(T�Y&>}k�(��b�� �=5V�q�O���M���䓥�4����(��"Z(��KuF�1��؉��A��M���?�*O��r��T�ݟL�s��Wș�p� aP�'-O�:����&�d�<����?�N~�Ӻk2V@��j��&Xm*=�FgR}��'�>�bC�'[��'���O��i�y"�*m|DL��C	9�mg�Z���<q'��ħS�X}K�E�*R'$���+�#^�om�����ȟL�	៰�nyʟZ}� ީ�5��iì�)���`Y0��7[����"3�Ş�?97 ��dtP��"�XS�MF�4����'}R�'���H6�4���D���Xgi]6&L��t�}���:׋r�z��$�$e��O��d��lB��ۗ+�浊pJ^=r�aQ�>�`��D�<����[�b̌!b(�m]Dd�dMŎd��ODu3㖟��	�\��uy��\:�Lu��B�=Mt���i�'�L����4��O��D'�$�<��,gp=2�`���8�iBހq���o�`�'���'��U�(D�� ��TJ�>,S�0��d[$4�ށR�b�����O��d4��<�'�?���D�xm�x*3�0�9bĤ��!��ٟ�����']��둈/�i^i���
��\���h��&�lZ��$�����'��v8���@�ңE5\��j�PN�oן\��Kyb�����b����kO���r6Ɏ2~��!Q �5�'���ǟ��x�s���8pr/Ӆ�0��v��68��6-�<��a��T�����~���
B���j���4)�� �Ō/l�b�m�2��?���h�O\��M�&&V�P�@IєO�x��Sߦ�q��؟0��ɟ<�I�?����	V�-x$�s�lC�&��2LT6l��)�'��z���}nf@����| �(Q�F�1U� d��4�?����?y�J\ ��?9�Op�A���tj�Ѥ�3��t ��b�';��6���O��$�#\,�u�P�n�D���NA/yop�o�˟�S������|�����Ӻ+�k�!�,q��}7�4#�Nv�ȟ@%����]y�'��03�A1JF�0�J�0���A��L�3�����	[��?i�'�h�c�&'_��Af�V*\}z�4]���'U��'l�Y��y�����D�e��He�M&S?d![U�A�����O��d9���<ͧ�?9�l�y�
k$�ƤC��AS�)��XP���(�	ϟ��'��ɐ��6�)�n���Lʄs��x�L�	)(MmZПD%�T�����'��'`$���+F�ߺ	JG�.���l�����	wy�ֱzL�*�D�kL��(��M���"���@	< ?�'D��П��IE�s��ݤl0+VA�;���* 0vܐ��?Y�� �?��?�����,O��[ l�jR�nS8NvJ%�a/ױ?ԛ��'��I�Fp"<%>�Q`� 
�Rk��Q�B� ,�x��H�CA��!��������?IJ�O�� ����	,d)!DFн' �%g�i-���'��T������=�d$�a�5/��L2e��2�VH*'�ib�'��ē5I�����O�I5b]1�vk�zdBA0�Փ0�R���H?(z�i>u�I����	Cl`ٙ� C�\��Gojt�ٴ�?�C/��w��Iey��'��	�֘$6.� (Z"���#��(J��BXb�͓����O��D0��OJ� )�&�ɩw}& �Ca��C�N�H
OB}�Q���Zy��'�r�'��$)�Kۖ�| ǧG�Dk`�p����y��'}�'�"�'��Ɇ74� )�O�fa�E"�a�h���UR��޴���O���?i���?����<�R+54,�t���H%`'���.��I˟��	��̔'g�0����~���4,n���aGdx�T;�J�������i��]�������	��c>7��7�^�S@ɝ�n�L(b�ۘ����'6�]���H�!����O�����4��g�������{��:�%�[}R�'��'����'b�]���'��Ě���,��Q�Й/�zXmZVy��S�JZ�6��O����O��I�Y}ZwĜ�`T�D���q��c���dGi�z���Ot�ѕ4O�(��yr��L�3	���'��8X�>�z��ЛAI��9^/�6M�OH�D�Oz��T}�Z�pI� B��Mi�6��$J ��M��� �<9H>Y����'t�����9���0�����i�`����O����N���'��џ��QZޕش��
z�t���ǡt3 �'��.x���|����?q�w%6ă��֥7������
Y
(U���iqrd���ҨO���?�,O�������k�Bi�m�@�T�(�PM3D^���x�H�	�0�	韸��Ty҃�n���WC�2k}�pq�BR�U�U�`i�>�+Oh���<���?���a��dh�OT����Z���+Fw�pp�P�<q���?���?�����X�G"̑ϧ&s�
�
-$���4H��oUy"�'�I՟\����D:���X�
3�X����_	�� .��Mk���?I���?I-O�5�o���5�S7k2�Sób���(C��M������OJ���O���1Or���&�pbܥ�D�K��V%�׊oӠ���O�ʓs�fAӰ^?y������8tޔY	3��l@*��Pz
ݓ�O��$�O��ͧX��$�|�����>!��
$��1.�R6�M�/OE���ঽ��������?��O�Y���lЖe.4F��i0ݹ2X���'������ħ<Y��T�,|�$�ȦJ��OY
l��=�M��$yڛ�'�b�'��� �>�.O�tJ�SV�Rb�� Ht�1@UȦ�iS�"?�)Or�?A��@� ��f�d��Ks(VB�P@۴�?Y���?I�EZ�k�	Py��'��$(_�ȢE�=��]@d���}1�F�|����yʟR�$�O��$�Y�.�{�"�w�X9En�ƀl�ş�C1�V���d�<A���Dȼ� �!A1#�p?f���Y�m^�[6�ipB����y2�'��'xB�'��	� ����	�)k҄�WC �8v�� � L%��$�<�����OJ���O�|(�7KGZ�`rbJF��02h�'d�d�O����O��D�OT˓#Dv��0��+A�Z�O��!K�
;8�(ubd�i-�	����',��'�����y�@	w�N���8O�
L9���Q��6��O����O�D�<��fާ�O�N+�A�]�G���{��т!a�x�� �$�Oz�d����7}R��$�m;�+S-'�P���_��M����?�-O�u�s��R�۟ ��$��4���%b� SмQ��S����?q�R�x`��������+8^���&G���B��5(U��Ms-O���	Z��|���j��'�d�Eđ�x���(M�` Fq�4�?9��
�����䓠�O��<x��)�����  m� ߢ �4�?i���?�����O�<�W�ٌYh��5�� Mɜ8���ͦM���l� $�4����F3hx�#�թw�8���G��*P�Ѹi)��'��fȄJ�c�0��v?�&�C)���}2�|:"�Gަi$�h+ �b���?Y���?�P��Hh�=2�n�;������?3D��'�F�y'�4���L'���o� C�")��{�A�xoP�I�� �<���?1��򤛳\�R��գK&$�.Փ=�mH�)_�	���	p�I���I'4h������q��˴��8�Z���-��������'��lc�>� !ٛ7�zx0�R8��1�bͰ>y��?AM>q���?ٔ�O�<��,ʲ)}.ػP��
M�(=;eO���ğ(����t�'O�P!�;�IJ�M"�e���4��;�D�u�X5m�⟸&�����䫗�ޟp�O�u���0��{Ӫ�^��5A�i���'n前/��iI|���2�BG!z�����ֲK���Ժ>T�'4R�'�i�'�'|�I�0�P��5��[$���Pq�V�ԩ�i�M�W?��I�?�
�O���DY<#MD�q�K�J�)¶iCr�'���w�'D�'"q�$)�.ʅgjtL"0�B�#>)��i#�`�!mӨ���O|�d�ҩ�>т��$&����A,ï 3̈3h�����,ʧ�y�|����O�R`=m�b0	�^e�"�B%����	̟��I�:��M<���?��'�&%2��4f�P��.�]�t`޴��M���&��4�'���'�̀��.��c�^�r�̴:�Z�q�t���$J\A>��>�����{��)��z��I�W�U�G��^}����y^�x�	��x�OT�	\�P-�� ��u�� ���E��|���'B_��Ik�ҟ��imt$B��K:(�)�Ѣ?ތnZ1;���?	��?�*O����͕�|�mT1m��1�OL�`\�)��aY^}�'��'��O�!x�R?��RiJ"k�T,q��˔L/����>���?����?���E�x9�,�����:�ܘ���ߙ���§�ݸS\�l�ß�'����Cy"ˁ�ē�T x��%/� �xqOO�ym�An�ßT�Idy�#R�c����$��t `!�\<9m<�˴Ê�_Uv%ۖÞT��՟���
`R�#<��O��)r�!ތD�n�`Üs��	Bݴ��X��`�o$��I�O�	�y~"A�1<� ��ƻ0N`���?�M3���?ɤ�BE�'�q��]���(%�|XP�۬20��u�i֞�E�q� ���OB����4&����'	l��L�5mlP@�,����qݴJ| Ex��	�O��"�e���i�լ�P�ơ�Ai���	��0�Ɋ*�Y�}��'x�D�?5�p9b�柒:p����i�j�OF��A��O���O�P*�䟣?��9G�D�P@F����� 4�J�kN<����?1O>�1-nX-+p�إUD0�Z�bͽ`N@a�'�2lj�y��'���'j�	e��k6)ՠSFyK��WzQ.��&M��ē�?I�����?A�	��b'>9؊�1+D�HKrD(�G�J��?���?����?	v�Y���ԤL 	ʹ(��MN�8�F���ҿ�M+��?��䓤?	-O  ���ix.�:���) ��B��BuګOV���O���<!�
@$%Z�O���9¬� I�����7rN -�g�r�X�D�O⟤�J%�/j�a��P2�h���$F@�7��O��d�O�$ʇ%:�'��$��7��+mb���O�AF��1R��t�	ߟX�'{�������1Ea
�[�ҥ�c��	4�vԂ�i��	�S1Lh#�4 ���P�������#^�L2waQ3~�(�g�L�v�'�2g2�O��>a�/QB����uᒻM)�Qoa�  �P�Ҧ��	ʟ��	�?�[�}�+Ѭz:� ��L�v3:��	�y��7M�&�������0S�<��cC�f�|0$��-(���[W�i��'��	�u�O�$�O�	('E���ǉR�1��dk@-��od�c��*�5�	����ɟ1�CN�hl��r��'m��#6���M{��B�h��?1�\?��Ig�	�hf��@�p���
b����iM<9�+�u~��'xB�'��30qB�
4s
8eH8I-�U�C@����?����?��B��a��e�cN�uL�I�ků5I����y��'U��'�B�'�!Y�ԟ�Y���D,E@=F
�.Y��Z%�iv��'�"�|��'��	�<�7� ��'
�g���VI&2�$Q1�\�4�	����'��%�/X�R�'��OԊT[���r�	^�ʤ�G)	/L$^7M�OΒOJ�d�<1�ɂB�I	a�ڤ�`�V�:a`����;`�7�O���<��.��n�O\"�O���pC��.�m)��G�^p�./։'��'+k"���� ʧ.��3r͐$>h%Ȫ�M�,O���!�覱۬������R��'�ހ���\�T�K���OaD�[ݴ�?)��MR�FxR�i� o����6�6�3��!%�6c�RH��'#���?i��Ο��'bެ� J_[��%��ذ�>cOOx���O��I߂_�AE�=A�9��R#{��7�O��D�O��t��t�i>��Iӟ$4K<d6a�!"����2#����'�D��y��'�2�'���Q�ȜD�X�9���PbR��vJ�>�L�9�?������O��OH)d�Ӥ?�jH��`�?s�؅*Ak]P�	� ���?���?i/OhH���Z :�ʩ�������ȠA�>M\�>������?���g�  �f#<f�:��i���$C�t��?)���?�/O�HJ2/M�|z�*�8_�n� 'C��`0�SoH}R�'��|B�'������䈠H�B�')U3g�Y��Q�=����0�	��`�	䟼�㥙A���O��B�ɍX��	5�Ҁw���[t�i��|��'��Vh�O�s�8.�Jb#��x�qu�i'r�'H剖)m�ꯟ��d�O$�ɉ�/��鳯
ox��S ȵr�v�o�A��>�S��$��b/��}��M���\o�ܟ�	�yA����ğ��IП���L�i��@�Z�O�����@%]Ä�B�wӸ�ĩ<����o���'F�P����S�����a,Lb�0�Ir"�5�f,�G�|��!>;��98�� ~Q&q�B�1D��AK�q�B����h�8񸖉��t嘴���G�+�(Y�
�q����N�e��#��t�H����`��P���w�4�	�/r�����e 4%��7�@+�X�B��� ln0����c�dd
�!n��!�g ��`�ūZ�V�c��@�+��\�F*�wF@`�����	�������ug�'0>��`��ϝ�e�j��6㚂t�� aw��R��YWl
KRr�IGOEL�!D~m§y��(Z[x5P�S�ja�L��N��z��"p	�E���E��-J����T�!�aT�Sd��<YW��C1x-b���ʂ�� �Ic�'��O�U�C쒷u	J5��5�t�)�"O�$�@�]�'4�h$�K�;d���c��ܦ���^y�:]���'�?�Th��V����H/bKt�Y����?���1�`�����?�O��=S �[�]-4��ݫf�֨`�W�q�~��Ť�UWx �o8�؃bLڈik��0a�L8"��e�U�̡30A��@
40ݑ�/G�!��xr���?Q������+�Ve{�|�@ysn�"�1O���D�XǮ (�Ŏ.�ԋ�VD^�F{�O�7��%b��$(���}�l�P�T8��$�<��^�/ț�OQR_>���՟�'��
f(H�b
�1W���p��������x�
�n�$Q��"6�?�O=�S��R4��Y(BV������f�8�'�r�* ��f�2Q�G�1�B�Ǩ�RH�O�Ip�eA>9�� G�	a �!K�tyA�Ob��$ڧ�?)�J��_��%����-�p�F~�<)�.��^<IP#�ŏP�ZL;�g��hO�I�p�'�����*�P�zq�Pd���TIhӢ���O\�����ʧJ ���O����O�nJdT��B	$W,h����S7sN�	��bI���$��d!r��|���+�p���	�>Nx����'��<Z��J@}�ƈ�!����}&�S����`D���t�yk��C����'� 9���|r���М6����O#dY�]�B@"b�!��q�2����ʧ_;Ș��#�0@��	*�HO��O0˓�ta�~T~�0D���t)���Ё|{�L����?���?	�����$�O,�S�tk�P�!�&z�0��!l�1`��!UzB%M=�O�,�� ��E' 92'g�G��ʇ���n���`��Z����ɝ}����>w���S�"h��B���O���������G��v�
1U�)Ta|b�|B!�{�+�`�6$d+CN���'��7&���Owұ�OD�C 0�%��3� �sd
Àe�'v2�'�R0�����:#��U;V̏� k�6��?�����j��pNB�Qw�Q�`�x".C7j"�q�A�3qKH��7�i�j%acT�B����=Ib�8�R
}�	㟴�'=��M�Cclz�̈́�=:Y��y��'.�y(�=�^�j�m��N�Ҕ��x��}Ӝ}��,�7Sٞ`b4�Ǩ�J�����O
�C�U:5�i���'t�S'P�~�I�i'N s� Z�w�̺Q�%&#J}�	�4C��ǵ�c�P'�|�S�TY>��b�L>+P���'�)�Ib�#>}��C=HS�䊇oʧo{4�
/:�4��d"�h��
�/N�WL��HU>�	� ���I]���� �)�Sת=�æ�1\�� R�M1zB�)� �20l.d�&m���_�fHr�;��|"p鉗k�:$���H>3�)����)2�p�ڴ�?Y���?Q�L�3�q���?Q��?ͻ�^<)$�5's��B��)=����y�2��<��gP�Q	V5���*�n�@CC�T�qش0��	�*��Yh�HI5#� H�F�e�.��<q�F�ʟ�>�O�Q���7l��.��\���Q�>�!��}�J�ڔS����z�-����HO�8�d\�_�(��GK=8R�F��FΖ�0��۫����O��d�O
,�O��9�����&4yu�E1��r\
Z`����B,H��Pq6b�K���+w�"}=h  �#�O:TqbJBj�h��ܛd8Ή G��bb��' ��'�	ꟴ�?�vK;?��Ědg��>A�j�<iv E-�h	�`Ä�&� �'-�j̓f���nyٔh��6M�O�$P�*d�����,(ˣB��z�D�O>=��J�ON���Of�Ҁm�(~�Ƽ&� d�?� �+ɛER�Hw�/O�y�`��EĖ/��`@�B0o6�d��*�)��)��[{�\���+H���d�O:�m�� ���5f&`@8աŠ#��f�Ryr�'��O>]��M�"L�э�23�4X
�C"�O*�E֦1�w��YrD����E����膢��M���'�c�����S���e�gOE6pn���/&�����5�p�"A��iX���H���d���q.����Ղ,T���ȓUiT�� �P1Y4ɻ�G��s����ȓ|X0%���Bȕ�"h93�͇�78��eAU�A� �R�B]L�ȓ~RaA�.�p"�BFL��`Ї�5���(H`���a Z'%L�ȓ�h�s�h���D�a�KG��Vu��~�b��Q�߁J:� @�K�5nu�ȓ'�j���� �J^��M�)f���ȓd,<�{b�$l�����~Ϯ���F�!#,�j�T�
���3�蔆�Y�b���fðT1�A��
;	�Ԅ�|W��sbH�E�`(�`��g�H���L^-+���JD1نn��F���x�Y�q��?gT~��`��DHvI�ȓB �d�P+Lc~����[
>e^��6�(�q���+}d:R�O�=��%��_���k�VY#���c�)�d=��S���T�6n`cdF_�
I�ȓ@2\�2��ӋC��1NH����ȓ{�����G�g�|�1L�K�(݆�d�8�Z�L%]�5��	�sF�9��a��q�w�-gM���!�͜&���ȓy�XTv�W��q�"�H��5��(R� D���_�)����>7���ȓcYYIC@�;�X!'�^B��q�ȓ!����3�śqW��X��A�/���Y��9�4�B�RtA�ņ-f2L���IPQ|�"��9�?S՜!X��j�-ڕu|EJ��A�<)���.m�8k�k�I�$�I���C��:A�;�
D�Y��#}:JW+;v��ԅ�h,Ҝ)�
C�<0kГ(� C�E[�9ɷ·�Y 0 T��h��$�st�ũ���Q;����.�D�!�d�0_�(ppS��7m<��sk��N�B�3*Y���X؞��@ND o��r@H��QZ]a�� |O8x���B����4R��ƪ���Z}��.�'h��
����p�U�ڎ���Yz���?��/\�5dѻ��#�'*�$Ce��w&�����
I�)�ȓ,F,ó�i��1��QD�%�'�#=E��G�U
�a���̙C�.y� Nň�y"K�'X�`2�&9�% �n�'�y�kő!S:�h�iC�V@�;$���y���T����b �o�xb �]��y
� BT� M�()1[�ʩJ
D�!"OQq*��B����c��mXS3"Oʉ�Q.�(%�L
���
6�	"O�0�B��6s�P�3�B8�H��w"O4Y9�@�$[r���Ӝ�+F"O�y��U�Y��!����M�a"O�cu��	e>J0��
1'���'"O<�I8U�꽨%Ԭ �p|�D"Ot�R#�L"�^��S 5��q�G"O�+s�i�]������� "O���#-B� ��L
�-?y����"O�9VEЧ'�pY�g��\j"O̔�F@O#\���FJ�^���"O`A1����5Ԯ����}pX!c�"O�q;�ǰ<�}J^T����"O>�ȕ��.n�&\I�/�P
�x&"O�M3T��7u���%H�8��"OZ �Ae՝O�DU��� �{ˬ���"O��q5Lк6���C�ő��*���"O�p�FJEH1|���C��mx��"O*�(���U�~)�f�¯�>�a'"O�)p���&n�8���_�ȕQt"O�9zp�"ÖPSs	<��@�"O�@Q�HMi;,	(�Bލk�P��"OhM��ˌ�M-���a�8M�ER�"O��2�@&�X*#@�Je�ɳ�"O�u"!.��Jm�hn�6�z�X�"O�<s3n+��-�QL�<����"O��w��2D���f7����S�'���a��$�;{\�$a��VY�P���!�DI BmB���1V��fR�o��'k�X����ٝ3R.��ǧ˖\�(��]�@!���GG
��w�/ܾp��#zn�sp���>���P��� d��r���|B�˻�0P�b��S�����xB�ۉk�TP�+�r�Ѹ�P�2'�ƾ�=S�'�.G�y��	3bx̛�@�1Qp1O�S�{�:('$��X�׆X�(ۄ���X	Eٶa�ÎG�R�d�"��4�d)�@�6A������-:�X��-!�D�z�Iv��?�0$����9����FJ~"j��W���0�Ŝ�p���2(ҡ ��c?Y�5�ֹ%ܸ�J�s��ݒaG���cƜ=T�x��퉾$f�A�I�Y�¸r�j���z��j4��q#�;'hvy{�?�)�c`fY;g����M[�mC<��T��K454��%L���c�m1��(Ί�X�cSč�'
���Y�.Kb�{���v���8u�������2$�z�a��!�)a�ٶR��m�T�æÈO"� &(��B�,9�P�̀	W:T�p B�\$�Ĭ��Y��/ģ2������U�H���j!�g�IR��?�fF tV�EZ�B+� �3&��<AcmE�	�E�4�����bV�����$)�S
qm&���k�~��x�� >GH��Z���K�`�Q؞��gթ&�\�у���/��q#�@- �V�h��<=�����r!��O��SM>A �>����4l=&��c	U؟ ��j.<	�M%z�`b�� D|�)C��[��P�c��a��B��'�����ԥ�n�ۀ���x�t�����W��#b�F����U�W#��I��R�,�:���������� D�p0W���t�ւ{#��It�>?锥fvF5�� Nf�ԁЉ�v�O}��WԗyY0y#�-+���'s���CO>7�]�剆-h�R�17�^(^���qF�Ohـ�!<����i&8#���8:[< ���&�z�ē@NrQДϊ*1މ!�EC&]G��@�$%y����8r�4e��E��| DG�bA~�)�D�� V�����`?�A&�Y0k��$��U8��[GFҳ8�^�u���h6!�K-V'����M3W%����/��O��	�N�'n5Q?���M�LE�A�B�h[�lڽ��d���zf^4can���;��Ԩwh%�����{$�x"��66��vm�$�����E��y�Θ}9��E!�p��HZ���%�`��H;�)��������&*�H3TG�t�fB�)� ���To�x��B�*�u2 jܓJ�*9@��L��&J�9^��5�2��'D�T{��.sp R���
j�4-;@k������2)��xa��l�5�A�ϟ|�C�I�P`�@�AO�e�|�� �K op�B�I�dk&l&�
8� ą%i��B�ɫ>���e������	V̈́B䉋���j2N�!Z�d��(�,A	C�	ML��0O�x�t��hϘ%M�@��P��c��R��MRD*���aI+q��E�����������p?�Ǣ\�!��� eI��S����e[�
��^T^��4�'���7�0#^�	rf@ث�\���Dޚxk!s⅟"c�����ɱ���~�BaRP똚Ȗ��u"O.e��X�J��)����.R�P�p��O�u�4O��:Ff��⇱�0|��,R;UBY*p��w�&�20ʞ|�<1$b?S����a�1!���"G*�˓?@p�AF�Ĝn����'��3�A�@'�L��F�9N�S�'�,���O�s~�����V?�pY����[�d���I5@�����犚f�p�+��Ι[�V��$,p����')�Y��05�bL��@T҉��'���,7V�0h`�׭I�,�Q�'�f�Gb��=�N���E�1�@��'@f�)��+� ]���.z`i�'��TQ�f؜s��(��ι���R�'���s����iq#���:�,k�'At:Ë�v=`��I�nq�P��'�ڨ�G�T:J}`��3i�eT@�y�'���� �ڣ���:4��5A��z�'>����Xp�Г�G�)I���	�'Q||y �@�h�8�[�L�2i�
�'�lɦ(\�}��;i��d+	�'�r=����:�:0��8lx8�	�'R8� W�A��U;4-�5t��E��'�V銅˜�c��i��dތ���'J��`�Ⓦ !�8Z3�2�vl��'����%;���q�勨+Nh�
�'�0���)�sܢ����M���	�'��K��9����P�ʡm�>���'$�h3
�+�<B0m��p����'*D�9E���4@�U��˺�� "O�\Jp�7��ٛ�k���^�J0"O��2SB�	5C�(qs
:$��0� "O�C�$k]P�*Ɖ�$d���"O�쑦���=���I��C)%]�!��'j��#6&ܤ
��Ta䆅�:s�I�&�4�J�2��ŠD�����>��x��؋<�`h�g���,��@6��I�;Ny�	�hҌ9;�I��T�~"B�@*{5���!�;2�h����s�<Q�'�R��a�Ǆ؜4>n����,!p��a�N4|D��	��G�_I>��}�I<����B�~`�ҧ��>a֔��Ni(<�b�ʢ}�����d��N������I#�p�w�Ϯ9G������K�tp
˓6�ؔ�"j�<x�l��g�R��}��Ɍ}���D��"����Tf�V�t-RB&a&e(�HJ�~$Ƞ�L6$��QQd��,tj�n�: N�� �.�>}D4�@k#�
c?�`�a�>,G��T��>s�i�h-D��r1��&'w�Tp���N��a��O�O�L2�'Ic�Z�L�"~b�@/fN�<��[I	̙w�B��yr��d���E?���GDL����B
���o��<Q��%6�x��.���x+1�\���X�g��l����u*~-:�	��+�)ѹ��x���D�����ޝrL��ن,�:�yBƒ! R.�Z D�L�C,ޫ�y2Ŏ�1��k��T�` ��3E�P��yri��5��3��4$��H�����y��Dp�Z=�r� "���IP;�y
� �@i%-@�X�,D���&O�0d�"O���u������ H^�Md²"O�<QgK�86	|�J�F�#D(q�"O:xAФ[O {�Œ/��3"O��rd�ԟ=��K.�<�"Ov�+�d��9��u��jT7"��=0"Oޤ�	X�N7��b�'W�3�.<��"O`�b�o����(Z'g�r��h��"O̐3$��)c#�T�0�Oٸ�!&"O� A#/���ʣC��"1�S"Oz���R�]�l����D� ���'I0*0���N�2E�(�ƴ��'o�(2��^|���g���qWJ�;�'�>8����l(��#��eI�=:�'��u�`/�0x?ޔ�,ˈ2�Q��'Ж`R i�s��T��o��-d�8�'�$	��ׯT��	覀ڸ*z<�x�'��D��Mدt&鱧�P����'	�MCU������6�_y��]��'�t32�UI<Q���Q	j�� �'s��F&�#\�:��[� ��	�'�-آ��I�lEk�O�R�FL��')��i􂋩d�ʘ�K�6I(��S	�'9���EKV�`{���A��H�ps�'�D�ȷfM�R�H�L���A�N�<�ӍУs�|p���MY�dR�q�<�q��8舩�5��A��Xo�<�k��E'��*�O3w��ĉp�i�<��D�ҴBG&D6f�(�ڶ��<Q���2!��i�àʍp��bpk�}�<!��1V-��⇌B�*�*�Dz�<���2&�8PƊ�}��8�djM\�<)FOُ:��E	�+�P;�@���Zb�<�����RUOS��)`PjĸY"�B䉮Fgb)W�˶�l�6�"O�B��.���B*<8�:Q��J��z��B��/dÒ��VCLlZUᦫ��[i:B䉢
�qe���<#yh�A��+�B�
0yV�V.
��:Ъ_9Kj4C�	2g�<��N�R������&P�dB�I�$m�!k0.�4̩7��l@B�	�9 �((����l���Ǉ�-x��B��mV&����A�!��[se
7K��B�.c�X�ٟU�����UՈB�I>�,Xa��	F�����,"�B�1xL)$	Ƃ�������hB�I�5��E�l��t�S�ۮ�8B�ɩ�N�eW=��`���؛snB�	;x(Lc�E6,�C��zw>B�0l�$k&/Ћ���J�@֯;�@C�=)�����^XM�����ҵ%�B䉧 �"�W�Y�GkF܊B�I^��
�F�|��EZ ��N~B�	8k-���̆��֮_2f�DB�RGX5��� U��ѳ"-��2QB�a@�l��@�6��r���8s�C䉣�B�����=Õ��n7�C䉭YJ���(ʊB�8u��P�3�B�I�t���K�,s�8EK%��N�B�	�q�X���9�N$A�YӲB�"F��(�EA)K5��GG�#J^B��$0&8a��Z�T��@��C��M�2B�	�5�"����u��H�@���Y��C��27�YÂ�߬Q^$�Z�7IK�C�)� P�h��=u����UǊ� �-�"O8`��%H).4 �悚KZA�r"O�]�#+��C�����*V�W��lb�"O|��U�5{
���J�d=	"O֠�狂H�:\�$ǝ,]u�"O����\:49!5 [w�0��"O.��	9{s�����f(a`"O��T��}��j E��dS��R"ORЈ@J+腣���43Ih<*"O8}�'o�5]���#��wb@鸇"O�eK�(�;r�ڔ����hC�P�"OdM8�ʳFa�X�f.܁�"O�p���1y��|0��tZ5:�"Ov!��L��Y2w�B	����"O�0U*L�s{��#��ӘN)�XQ�"OJHB"@E)9��Y�e�W~�%*"ON���S�4P0�9 -x�"O��� ]?>&A%�A��19bj7D�((T�׆Kx@�a �
29�z�c
8D�\��-L>���Q�d Q��6D���W�K
)�x@�vaЭ��Lf�"D�03�F�7DFU���ͨ;��0� 5D��*%DH'O�p�K5��<r�0y�-D���t&K�I�Z���o��L�`�+D���vl�S�H�2ĉW�t�� ��F(D�HsҤ�/G�`�+���$��� �.9D����<7��XT�Tp�����6D�����9H��ٸ��?T�f�c��2D��+VMJ;/=di���Z7Z��B�1D���d�[t�L�ң*�.�Y��3D�L���Cv�H�0��0EN���!�1�O~�Ob�v$�R����(�/QX�Hi�"O�|�wc[y� �Ibm`*
�Q'"O�[��Fpb��F�ÜuhU�S"ON�G�UN,����I��1"O��#3̒\v��a��Z�yj<Q&"O�-�T_�s9����L��aq$�'�l�̒/�bI a��<!�LX�'�1&��R�v�( ���{�h��'�|E��Ǝ����@�(�D��'& )5jO��F���� .ZƩ)�'�؜J�$	*p� i��qߠ`�
�'e�`!�@.����Gkި2p,%+
�'ef��6�^� ?v��U燂���	�'#\�s�iX5!�#�E��U�	�'���C����I��?����'��� '�K�u@~y4�E�}V@9H�'46Ĩ�F,Km������=xj�,��'(
�(`�؟<�\���0�ԥS�'0ҽ���Hzd+�J�wAx�'u*�h�쎇.�СY�m�:s����'I�t�����J�0�+G=�J�s�'�����!�ZQC�.��:�@A�'���GN�!��$�w�4�����'�$M�.�'F������T�4=�8 �'΀\�'�[R0lCV��0�V�Î{B�'�JX��ꗫS/��CdLĉ?��ɠ�'f��3��M�#8z���R4=�Qzߴ�Px���4G���f�@�-=�q��!C�y"g�)��\��b��*�}8�D��yRč��@y�m�'$�ѫwk���y�ӺW��x[���r!��a)%�y���-t]���C��{�����*%��xB�L<3�"ei���T����Ƀn=:����� 2�iu̠�~�9��A�?.���'��O(]�X���h�B���#"O�YID+�:tA��ɲ�ٳa��qs$��6�S�ӓ[�p�- �F*(�1CȈ/�B�\ ع���1tFډ°	"~�B䉀=��tg�L�V��������*ٔB�ɀdh����
f�q��#A=�8C�I8#0� A"�,U����5_=6�B�	��z��N�y����B¡R�B�IJ���!L������A��B�	\�,�WI�������H3t�C�I}L\ˣ�t$&ͣ��� ��C䉿N�T���
��Ea&U�$"�<FL�C�I�ڈ� v�w�8iq��f��C�	 <ƌ�0�W
��a��7g�B�I�4���`F�ԤTl� �v�B��]k<
��?g~� ���9K�B�	�mp�����	JvxP{%�ʮx@�B�I�;gKp&P�m�v@n�H�B�I7��"Tgρ'�Z8 �M'!d>C��u����ҭ'FT�Q�DJ�a'dC䉫6�P���Vt��y�4�F_2�B�	.?��e�`�R���$�P�B�Ƀ*
:|��ġ@F�N�����"O��(�G+I��T�ÀI��u�U"O��ۡB!P'V���IO�&����&"O�e���A�$�2��F�1e����"Of,�K�VĪ��K��FH����"O����	J�ty&h� ���Q�"O8�
EL�,D	$T��F�.~�n8KC"O���Ch��X�h����\����"On��dلf&�qAN6S�Ѐ8T"O��P�O͜^p��b_�c��'"Ov=Z%EĎI?�$y�U�\L�5;�"Oꐀs`- �84�D��8|H ��"O����+�N���K�, x�� "Ot ��U5��5�"���d�8�"O� a���`, �{/��2�-��"O�)�l>2C<�i�	qd��"Ov�8���NL�0;�a�Sh�(��"O�i�)�c?���V�@6nO^D�"Ov� ���k}����ş�?K��h2"O��Z��̀1�	��W��ax�"O�h�g!^�����%Ջ,��e�`"OZe9�]1?h8x�`��%P�)��"ON�pU��59�y��I�3���"Or����N�k�<�GƈZ��4"O�EqE� /���Yc���p��"O�)Pe%�$}*ܤ`P��5JĨ���"O~ ��)w� 5�'��,����"O�!-Q�r��k�@(|�ֽ�"Oڈi��t��k�U�Tn*Q�"O �Ƒ�v���$�ui,�1�"O4�(SFū4_:5x�eL�BRd�"Ot���J�ga�d���&ot��"OT����>Rd�itၺW�`��"O�H�'C���riуO�2&v*�%�Ii>�v�1v��B5�]?
��0�n7D���dʇnL>�@0"��h��QS�@;?�
�^��0ŕ�CFNA�dV�8a���ȓK��`r3�9���+	5\�,�ȓt���v�V'X���bS���9!`y��?`!����	vO��p���/.08��{�T�2�	FZ1Ǉy r���S�? p1�,�]�ȝ�d�<:�z5"O(�� @ݹHl���Q�B�OHH�"OB!1ƃQFs�1�#��,Y�P4�D"O�P�o�s���{@��.�HM�"Oxi࢈�l�Z�A��Zpx��"O��Iv�P�x���q"�]h�(7"OT��O�m�ƬJ��3%�Tc"O�#T�(.Na�g��r�:�c�"O�MkA�b��w���T�u0`"Oh��d\��w�O�+F�a"O���5��y����3L+�ȸ�"O� �,C�(�(��~nv\��"O��Z�@"��L25�:��6"O8���ǏQ�`d��4bFIy�"O���Kɱ:w��b�����d���"Oj�Aő��>�zF@��=���"O���?��-�$��O�"��"O�(K��J�p�v����A/�α�%"Od�A�P�MQ��u'J nu��zu"O���U�^�jtӂcވDo2�)�"O���+ģ1���A�)V2U#"OȀ�Ѡ��~d��h�MT�oF�a"O2sl�0�8���aծ![��"O���'����Ph��O�App�r�"O���%�Ĭ�Ѐ��%]8�)�$"O��K (\�nh"3�$ϖ:0�q��"O�)��-b�^�6É<>�p��"O�<a���:h�(H\=rM�8
�"O|L�dI�U�vLU�ؐw$��Ӓ"O��S3�JpdhL��D�,~<�t"O�-�:Jtx���r	����y"�1�E���B�+uԽ�����yR��4���bP�J^H1�E���ybG�E6��3S!�eR@4�7�V!�y�]>}�� ۑ�ن[ئd��ɑ�y��=M$�����̼^D$�E���y�l3MT��p�IǅJ����1�N��y��O@���ֈ�2@*&�jN	��yrCǱcB.0`�LV,l�YѠ�
�y��$wS< 	u�	O#�IU��y"����K5�Ύ-���eʗVG!�$C�T��EB��ZaH����)=!�ې"�<�*��9]R�@��;K!�P=J�A�a#+yG	#�共>�!��ʞ[M<l�h��0������!���2H���"į%<���_�>�!�dF!vzE�����j��#��T�!��4<��=�`A_k�
)yG/P�{y!�d�77c0!�M�Z]��7���;�!�Z�@.nHxe �
s� -x4!@9A�!�䎲|*��H��J�`�H�ڈ5�!��*ِ����=.2�ITn�j�!��a�N,�Fb� �Z�;�N	&%!���'�������s�){2�4�!�$����j��#% ��$O�4�!���͚��cΟ	���nE�!�Dه9��H�A��u�p��-
�Z�!��D:��C�f�}����6ʑ�w�!��4^�e�Q&��B�(�)��ԡ�!��Wzj�2��V�2�o�%w!��R�E���b0H)�,,��͑;\!��H�IVh)�,��`�4��r*�m�!�$��$^�b��P�Nui���y�!���2i�B3��ݮx`,@�
���!�� �闥�9p��D�慒)2�N�"Oa�
�9;� [�I*2��L("O(Q�u$�0���c׾<o\Q؀"O(\�U�Q�p�pA Ҭ��GO��Q�"Ot̀���+��`ô-�>Q�hZ�"O�8���C���	%�V�W(Np�"OCAE�H�c���t�!""O�<a�a>
�
�Cs��d{�$��"OTi)�ٗ0,�R`&_�Cf����"O�j��
1|�ղp$�	t���"O���D*eX1C#�Oat]Y�"O�@��$F-w�|�A%���o�:�ʧ"Ob�K��q����?2�FP�g"O���"Gο4gX����$S�Z`Zs"O�X�坳:9�dc[68vIjd"O�������$�bͪn�@a�"O�|·�N�"ʙ�P*71?��"O49����h��Z6+0�ݘ "OFDQ#B�9�z0����J���"O4�K��)$���`�Qs
��"O���ԭ���I���ab(�!""O�8�©F�NpZ���=\`��D"O���u���*Q�T{`��DUF��"O��)Q���ht��)"*�"M/�xS�"O �p�!Wj�v()2)��L�-z"O.l�cD�Q&����GP=,�a�"O�D��N�V[� *% 3��22"OP*2�(�61q��C�F�)�"O<A�d@�\8|�)��ǗF��u"O��B�#G�!��t���*���1"OL���
�?��|�C��r�r��"O.�@����H�V�" ��� "O$0�f���}���i%eC�(j����"O�Q�$Q2Ril#7*�ڕ�F"Ojɓ�ƅ�@�d�X�ɉ(1�R"O��y�`"`<^���I
L05#A"Ol�r�j
(I����DO	�Uc#�"O>��W�^��B9s)�0Y$�<��'�x$����9�(Hs��P1���'{� ��_9E"�eX-�:q-��'����.WQl��E��v�5��'�r���"Q��s��i�b��'^|��7$R�Z.�	Y�ːK���'F�Ԓ�����I�ˀJ."��'�h!�&'@�gr����5G�����'�z8�$`_�U���"�c�<C�N�K�'b����8\�maa�#7����'�Z�e�,Q����n�.A�ȓnM��jǅ
P=PP�n��a:�)��#�@9���ƆP��˅�+ؖ\�ȓyߪE�gW��!�R�J���ȓ.4:P�5nHc� ǦF�bt�ȓ5�n803�U�!o^���]������P�@��N24�3�^'{�橆ȓE���b
A�\ˇ\"��Y��"�R����>L����"�����SZh=q���H��W|6���S���ܻu�&�"�K�0[���ȓQ�� �dn�2E�:�7dO�6Y�!�ȓpE��j��/R���7�U[������)���PQ\��`�Xe�$�ȓ4��=�Ti����xz6��� ����ȓE�D�і��S�T��fN��|@��r�� b�M���aF P�U��S�? ^I�EG#f���B��8���(�"OFr��:�hhГ�HWvN��B"O�e�͎X�buQ� NjT<Y4"O4���D*OK�HPh�S�x3"O�2w�U�'�&Y#�ֳN�+"O�����'H"r�٣�I:m�Չ�"O�9j $�P��:�Z1m.M��"O�9��ԧ/�l���|_F�9�"O��#D/�14�D�"�ꀴ��8 u"O>����᮸��cL*[�<*f"OX=AiΊ	�P��a�D��4"O0Mʃ��1h����Hbu�1��"O���Ǌ�E��3��HffF���"On(@�� &E�`���W�c~$�R�"O�8�N7���F�R��x�w"O��)��
�Bfyʡ��S���"Oz��k��I��� Q�Z��U��"O(�Y�fU3l����@�Ėպ�"O"!b^|�&k":�0ځ���x!��N2E*�(b�O�$nҴrP,�L�!���^f�g�$P9�\�V)L�&=�'ca|��K�|��1
aC��'���P�ly�ȓ36��s)��h'A�Iś;ڥ��=�>�A�fV"n��)��iA�@Ȁ)���8�:'��Cc��!���-�Z���xҌhJ��A��U`�A��ͅ�=� � ƥhAN�d�
�Q�������� �O�!�rz���
wn�?��y���P6���'L�����K�*��ȓ&��b5��40 ����l�Jf8��ȓGOt�k�EΨT�X�%._$(rLŅ�P�J�H��  ��q�RI�!��0��D�ĐE�����6J����\�ȓ	F��!��:t�����4�`!��u�$�1����jiXe�L7N��'a~BmːSPې̈́ӌ-��i��y� ��)Ba�ZU.�����?�y��N5\�5�� J�X�c���yR��>S?Vk����E�(����Y8�y2%�|ՒQ��fK���y2�պ>$ij3�8xsD���(
��y��}@=`4`�Y��Yq W��y��?�}��I���P`ĝ�y)ςl��$K �*���`��y��̟?��е�C�y�j�P���y�I�An�4�M*'�L@ǈ��y�@B�Rb�)<�*��m.��. ��PA =B}0#%�2E��Ij�'��-���2܂)1�#��Y�� /Ov��D��S���7g]2\C���f� X"!��0S��IDœ�9�ڥ4J�|!�DG�Ki0��R,��"�Y4!���T����  �.�`��7!�D�[b4����;	 x��H�!�dN.&�@�� �t�pfe�]�!�đ�Q�EB!��`�aā'�!�$R�[wؐP��.ː�;GDߋm�!��A�DD�� ֳa��p�B�k�!�	[]d��k߼F���PQ��;4�!��ޘbVB�s�#&�P�JA�u|!�$\�e�!��n�o{4�8�lQ�g_!�d�7���ui�6Q�"QzU�Q��"�)�d2���XC�X�l8zh+��=D��J�@�B�.�7"��,�ĩ%�0D�� r� ���#u����s�P `2a��"OF$�al�8�8
6�K�A!��"O�˅)V2*!�̰�
�`�މkP"O����� Mx|1�J˺f�3�"O,\�b�L8vK|�f�x��5�'Rў"~2g��]2�}ZDd�V<(�a�yEB�	�rج ��gȽ�ڼ�%P5Z$B�ɨɶ+��ΧKЈ�ţ�}�B�ɼ\��⅄�;frƜ�p�֘O��C�	"h�N� 4L�5Pm1��0��C䉻d��=x�Ho/"5B��SbB�I1S`�<�6M�q� 9E㐈$�B�	� V*Q	7��Yvt���'l~�B�I%O �g�dB��P�Y�77 B�ɩ?�t<"�H�&h�b$����.��C��L� 3��=%`d1��Ծz�B�	"jI��`r�/[���Q���!]��C�	  �pHJ���=-h��� !��f��C䉴^���S���] ��ⲥ��=	Ó
���A�#��	mI#Q���Ͷ��V�"p���xqn�\
L����l9wC37��*J쬡��<���S�Q>trE{�`Y�!"��1��t�׳�]Ђ��M�om!��-l��Y��ߎ�t�K�Z!��UR��T��J�	X�&��S���QU!�D�1<t��r�HUu�����/�3N!�!dyY�a�Oݸ�1��9^E!�D�Z^�z��;k��y�C��T�!�dī&=�4�p�ɴ�
�VDǇUW!�Zy7f�ST�7��UZ� +�"O
%�&�S�Tt�H�
 �tݡ񄍌Kk���`
!My��0��F����hOQ>ixsQ�e��x�4�*L ����d+D��9� �!;4T�C&jЎ�ҽ��-D�p�&�Dw����Ǝ#�ڌi&�+D���Ո��F�5(0��>s�tPh��*D���$�:���Y�ʋ	mx�$)D�L�u�Τ*�$��bϊ� � 8��9D���׭ }�t
0�	&W7&��t�7�O��	�.��0slR
.��@ ��� �tC�ɘ�ݚ2��)�|"'�/]uBC��>Yd.��Ť��[\�l�BE��!��D��tEЬ*A6ɰ��_\>!��Y�>ΒA���hDl(s���d�!�D�����[ ]3rb���IM)!�ĕ�B`|��JܿW��L�6!�d�+sw>���#��«���!�DB��J��3�+�F���IW*UE!�D�*z*,*��� &�h嫅+O�G)!�$�>�Z�S�ˏ1o�,��
��!�ܠw������^R�H��5C�@�!򤅦6�B���u��q��E�!�$�VBR]�fK�2e�耂d��Z���)�'!%��yDB�"� ��(���/O���$��#�P0aF�ù��0C��gy!�D�q>}#b�3c��m�=?g!���9�t�ʢ&�&/XJ ��چ}�!�?t|���#�IH�a�ń+�!�ľ����Gƕ8�6���4;!�d�?:Ph����k���'.9L�!��L�8<b��"'��o��i�Ο�n�!�Dͤ^��]S�M�-��p)�|!�D[�m�urSB[	0�, -xf!�� `��䠁�x�E�a�8BP���f"OhCQbjV�A1F���GiT"O@[Q�5�X-��n�&�xDJ�O~��D��,\�%���]�)�*�"+>D���S��S<��ҍ�'T$`It�:D���A��b'�$�3�^�iu�����,D�d�B�� F�J"��>E�5�$�,D��k#�3B}\����;*F:X�V�)D��Tb��L�ڱB�l���A�"Գ�yB�cLȀR�F9Ō���lف��O�#~2�f��v��B��,��ƀr���0=	�	
_��G#� U�0�S)�r�<!��̧`@�Pj��T�IX��Q�	q�<�a�)w���c��E�x��z�Yo�<�b�V�4���#�`�n̺��q�<qv��#�h���[X�	a�c�<�sj;?��9���#L]�$���[x�$Ex�#�$�����W~d�Q�F�y����f6��񃀖?q
d�ʒ�yBk�9�١����J~L�����y"`W7<u�0�6� <�j�ӀG��y�7.N���R��2Bb��@S���y�蕣JZQD��Gֶ���G�y�S� �����GէR��X�� ք��O�"~�`*T@u�q�ܣTz&�Z�����%��G{J?̓1aVE�qb�70�^m�:D���1�B7��@(��7 Za�Uh8D� �R�[�POx3)��!6i���6D���N�#P��@BAJ�d�r�4D�*S˧KZ��PCA��`T���$D�h�0�E��� � <�`��2� 4��U5i���2Nil�c��U�<�Q�ر#m�92���h�z���M�<�pj�,�vm��Ǟ�R��(VI�<��-[0 )DC�|(�Y�C^�<�Pj
�<����D0nBE`�<Qҩ(ZT�*�LO�}x��7jR�<�(ڳ�j�S�O"O�t��,XG�<QFLY�wZz ��+�mn�)�KFy�'�ax��vD�W�]�9�¦X��y�(��pQ�s�C F�b1���y+D�w���:!-�@������y2��!;pT$����%����-ʸ�y����̸�$!�A���7�yb�L
"���s���א��-W��y�΂�CL���m�	2n�PF�ϭ�?�,O"�O?��Q4hx
qS��8=�F�OS�<���
�T�����>/����WH�<	'�,(0��� F�3�6���NH�<I���2�r\aRn88x�I��
G�<1$DJ&I��kd
���l��c�w�<I �W�%�I;`$�&P*�	�e�z�<A�jQ�3�и�#iK���HJt������"�V��C�	�?#�es�B �\d}�ȓzD$C�*����Rbg��tM��R��͸�F�9RTyC��d��̇ȓ�0U��N�@14��Un�i���ↈ�VSS����K y�ȓ>��r3�]�Q�l��"ư��m�ȓT�>8sp�
�G#.��4��)؇ȓ�͛�B?IB��@�	 C@x����x2(߀q0�4 `j�)�T��"jĵ�y�V�.�JI��ӳyG��2�V�yR�V�G�M�$-v��XJ���!�y
� >	;҄�����P��}Yu"O�D���t�XJ!�ȗ'n��d"O�Ha�d04S�ٳ�K�W�n��'iP) ��#+jPX��l��aG>���'F�Hw�\���;.�[v$�A	�'[Й��eY8a��=��g��T�̽҈�d&��ai�ȕ|�
�;�ݿ\/�� �"O`���V0�6���Q"n�\��"O0ț�L��U�Z �-�0����"O���1�9,s��q*J��P�t"Or�qu%D�W����aCK2�޴q�"O4��+F��D��b۞X�&D+g"O��A��G�ZC~"� ;�Z��b"O�0ʆ��LU9a�.���*"O���Qm�%��HVd�y�D
�"O*�c iF+ �9§m��RtRe��"OZ����[�gU 1�t)BI�R�[��|��'�L�c���X���)��W��%p�'��xV��8RY���6O&�Q�'b,�p��n���EB�]����'����G�5T�PӁ*��.��'~B���Sݜ���,�+X���"�'��KFԱ���s�S�KÔ��
�'��PfeԃGXН���K�J\x��	�'\����!���74?a8���'�z�*�o��ީ3���o�q�'��
nB!'�}:�EE4Q�����'I�$�mݛe8nY�ad��L�}2�'_�pS��%�,ȠɁ�V1|���'�0�Q�g��HC��t���zr�$6D��Q��.>p]�q�����E�'D���7����)
��܉Q�|�8pE'D�ȉ �"�Ztxe��}�D�v&D�x�T�C&U8"�8��ÂT�R�7�"D�ذ��TA�� ͲR�9���?D���>wB|[Ҩ��z, T �/�y¦ߐ"����GFH��L]��>�O�a4�C��@H��)-�fhzdU���'�ɧ(�+�U�V�ࠩ�K�;t��He"O����
0�歹Oά)i(���"Ob)�Ǖ�/���z�I�iL ��O\Z7�OO�Ɲ���	^�bA�5D�c6/ҡ;�4`�0�?^�6txj2D�(�@��c��a;�狙0�hwa#|O�b���"��'�0�Ӵi0[p�����=D����R�V���o�%5<�)9�o/D���� K�*�U�B�K���#)D�4C���^qp����B�ַ8�\���<��O0)��j�{�@�J_8B��K�"O����DO"*�i��*��LqKd"Ol�8O?	���y�j�j�"p��"OH1�H�>*qt�k&�R�!�B�;�"O�SpJX-z�l���ʈ����5"O�̃fZ�z���H�G�����"O橢�������*c���k��I[�O.���'O�.���k�*��4u��j�"O2���j]B��b�ױ7l�\�3"O�D1��Ab� �����\�02�"O�E�l�`v�N2`�22��#r�!�d�'�r���F�x�D��0.V&�!�ے��tٰ��J�f�%&�!�D�T��-9Ћ�?S�������f�џ�F����2h;���Ci��%.6�A��V��y"	k0F(�e��#]Б�4�C��y
� H���/O5'd}��c��-�����'n1O�P���4<��`���{Ex!�V�'P�I�pW�aC\*"m��;6k�Uv�C�5tL�C�!�#|s��#��|�C�;n���;bjs߮Yk��h��C��>/���&���F�Y7���Ms�C䉡ou2,��HO�7H;�BP�z!�C��=�� W.�V���F�f\,�ȓe목b"V�=n2�)��K�^��'ja~�.S4�!��̩0��a�dP��yRhʌW~TKv��T�a���yȊ�53>����N�t�34�;�y ��^ɰ�%M4��yæ
��y�
Ր3K���A�
�p�P�"ڬ�yB�����hC'e�rѲ���<���dO�V�*� �*�4g��i!r�A�{2��f�Z]��3���m�o�!��O�L���,����0l�59���^!RZY�R���(��!�I�j/6B�,#3ZP��.˰7�E+��J#X�B�ɉ*I�ڗ W�p}QA��r�:B�I0U����	�u6~�A�G"t����%�qz<��uc�w���b*ĘM��C�	�z�5#�n�:2Q��{�E�dzxC䉟69��DS�2r8�B1��
Et���;�	�yԄ�:E�'k�nE:����HC�ɨa(p��7��
������nbB�ɇy�v��"�Z�Z�d5Z��Fd�B�ɴur1K�瞹 �����B�I�2�1��gձ+:�#���6Oz�B�	�s����M�`��dKBZ�B�ɂPܾ�p��I&%���`�E���Du��1vC�3�
i�gǈB
a� %�D �O�颁B���f�TAے�~� "OJ	��#�JvZ�F�_
��(�P"O�yH"O]��P`��L�a�,I7�'��	�h���� ɻX��Z���<6�B䉿<I,D���N0����V�L9D�^B䉱i#�a� �U0��q�o�Q�JB䉩f$���	��3���XG�V�	�B��HLH��qN�+�d���%bB�I2���w�j�J(�6��01|�C�I�C��)`����4���pU怱1"���$!�Sx*�ʘ-H��f��:	�����Y���pW�&�$��U��:0j~l���B��PN�&*�:w#_�o�vM�ȓ;aFd���!�Y��HS�%4܆����إ
�;�����'^ڄ�ȓ�Ld[W�U��j}KA-D&9��t�^��e�WD�����<'<Ņ�|F\�f��.С�b@���ņ�}B��+��X=!�쥩���x� ��ȓE'̈H�fA�@��`��v�Q�Ɠ
GR-p%��Z���qrC�20]K�'�i(�%���S���%�r���R�JUCS*S*��gT������/܊� ��c���񑀜# d&���8�řD�~�b�9t�G*Fh ��'3ў"|�R햪yj��&&�=#�@�I'�7�y�'ʝm�p4s�J�e��+�H2�yr��:(��X�wHR�����֋B���'�az��h.��p&N-���	Ё�&�y�d��wnhT�$X��3#V��y�愎o��}�"떡 �H�h"�M���O.#~� \E��T+�FQ$�D�DS��'����0j�� ��^
^{�Z�D�(��C�	5W��]p���52P��2�����C�	�8	> Ů�4]2l�UO�""�D�=��?Ɏ�J�<Ҩz��K"E̉(V���
!��35Lk'�H�w-i#�^�%�!�$ b^@P��I�~_���gB̙9�!���Q�
�cez�i��ܥQ!�ǔ\�(�bO�_�r8��'P�9!�d=cv(;uD�W��Q9㨑�A2!���	ܐ y����g������g�!���ZvJ�����khj��H93�!�gb☪g��"|�d�Q �!���5��@@@�2/`����O�`�!�$��mZj1�3~��@@�\?�{��d�
	�ڝ�T��wa�9`�n�Q)!�$�'�mi���3#�8H����H!���ƁZ!ȑ� �/P���]�i�o�6�01��+�z�V��ȓkl�蛀�O��:�2凃p� 1�ȓv��y���sn�:��͢6D���R,�ekF��ON�1Xb9D���f��-v�� ���
���`��<���S+Ml�3F-�$$tu�4	b�C�I�FKV$�b&�72�T+ )�c���=ç����H J��h�e"JS��=��#o�}��E�"x^���vȅ�i9|نȓ4�g��C2���^Y�ޭF{��'!?I:�߸F(.u"1���c5D� � c�6�~%�7@D,V��S
/D��hW������1�&�u�PF�1D��6Lݲ��p�b�6
��@D�/��$�S�'�bP���D9���Cwش�ȓj喐�e�d����[�A��	�РC�Z�H;09a"�SN�ȓt���S䂋13��8�O�n��X�'ў�|��"IC/�q�����zx�,Gxb
�'h�z�	�_=�XP*�����0>����!�ڄ���.^�HaX�e�p�Ib�	`�'��E�D�f/�<h ��P�h�3"OR8���X���yІ3\֒�U"OP�8��"#!TiFkE:nǪ�("O�� �D�0j��I��k�*aa�"O�|��ܘ3M.��(O�0�� �F"O� �휤!k�2����0i��"O.�Q�ٸtE���tn�Z����"O��CQ"ֈǮ4�-ݥx��=P"O�0&��/&b��@�ŁCJ^i�"O��+E�,84�7��`9E�"O�:�ˉPĔ�0tA�PX���"O�� lB6m�B|1�o�;P7�҄"Oj�Y��	J@ʃE[D�|�4�'C�I%[@���Fѣw @"p�G�rxC�I���E�T�Աc���Ƒ�//bC䉪����E����Yz�hˏl]ZC�ɫ-$e�	�h�ҥ�T?j|C䉖-9�&��&r����"�����O@㟤�I�&��"hV1�!!V��-0")5�A�<!��˹c^�U���^����!Ue�<iU��?p��N���@�B^�<i����I�Nr��_N!��P�<���.$ b&� >���	�O�<1v̘�<�;7E
�0~��rD	Id�<�� B�/�H	j��NhL��)�M�^�R�Zyb�� �4Hakǲ$���-f�Ͱ�"O��[C��C��e��E	!}+����"O��q�폥�Ι3��>����b�'��h⅄�[�}���%^���D0D�lH�lݔz�^�H�`�R!�cK/D��Q�b��qRI���W
	�U�0D�8(�
 -M����a�A"@I�.���?���O]&�x�) X-�#*\��V$`�'S�A(�,�h���)��I}�1�'��15O��8UI3nP<5T���2�)�$iS�xg�B��05�)hɍ�yBܻH�*��P炲 p�m(��ҿ�y!�:o�qz�̐.!�6 �B듚�y2�A�jT��IЭ#z�s�C�y2L@5e�BƄ�o~�i�a���?�	�'Sdq¤��vf�1�0c�2��0�'��1��F������k�l9�'b�E����WY��C���
��'�V8�\7n��y�7Ё��'�f�k!���0{�a�"Q�w'xQ��'qpD���ܧ��A�e�X�r딬Z�'�0�Õ�øX���#��C`!���'�Z�Z���K5, @6ǔ>W6Z��'����Ɨ5�DI��I5d�v��'{p���FL�Rg�|���Gd��My�'uF��J�,ĖA���ǈ2���'/^嚠�D=X �kV�� _��B
�'6�0kG.����W���J�����yүЦ-O��D@ĽI��0Ѥo��y����h�h�N<B�F�3DԼ�yb+F
Yl�����6?�ћrjG�yRڱ'|E�E�_%\.�ڶ�E��yr�ͽ<B.a��̞�V�:tK�E��y�ǈ>M`�3��U�f��Ǫ�y��&zE����c.f�Qnʧ�y�&��y���.b�*����N����hOq� ��7ǃO���Bf_��|��"OhX�U� �Lܻa㍠��q����L��� n� [��:���
ҴI��'D�`*r��#;�D��9��I���%D�H�C畖t��(R�5-L�0قf7D� )�jN� �x�8SD�j=����3D��KR� ��������j��Oh����
rX�4i��V�k�倁�ҷH{!�ͱۮ� ��T%~a�]��"Wd`!�$Ӄ���vaU$tC��D�Bf!򤁧0�J#I/j��iZ��	S!�ĕ�_������MQ�0�Vf�#&!�݀PA �Ո٦O��-[�8(�C�I�a�80�V��/vy�9�)��ZzB�ɋ(����RJ�#a���R-Md�C䉥k�x��'���!:���D6C�p-@q���Hy����6`^�1��B�I�'�P�Jc�2��d�D ^*BzB��=%�ْ��K�!����U@�~GB�I4v�~����"S�ƹ#��Z�]��C�I���,��$0"���ì�o�C�7���H��t����wʇ*R���hOQ>���#Ķ`�����Z2l�\���>T�L۳�Ӊ)��B�l�G��7"O=⃯X *f��� ��N���!"O��p4GF�A��]1w�I3�	��"O���*��HZZ��,�"y���"O���!ћ5����X�@����"O� ����.��a�ȭ�a*ɦ?9ܵb�"O2�Z�E�ߔYR�H��~��"OT��&eǉF������ ᘩ��"O�4���|��]��.hf�0Rt"OF Ѩ��L�8�.X*j���"Of�!��@�����9y��s�"O|�-!1�U�D��^�XM�|��)�S@8tm9�Ǆ<Q]�"��Cl���6�,�@|����	2̨�*�);D��	T�\�Y�P�[����2Y��k� ;D��#��e�Z�s$.� h=X2�8D�8`uJ&7�>q��B¥C��Ԡ1�4D����Z�Y HĄ�=��|��A.D�<�t,�/,�Ӄܤ6�pQ��.9D���mP�}��c��L`�Ͱ�a1D�P�[f�.���W�uG��3Ui/D���a͔
^r%X���38��3s�2D���Ԥ\�K��X� #п:���Ӈ#D��cD�l�,�sd��3` h��v-D���I�\�V!D�`*HQ
7D�����˺Q3�K�c;G�h���@ D��X%�
S}$�u#L�E8U	CĠ<����hOq��| �NT�C�P��@�E�t%���'����=�r�����-�\���
O'�`�ȓVAx��f)�)�T������u���D=9�-Jl���&G��ȓU����nN�}�Z���J��x?v��g6��FX:>�y��΍7zL��s����v��{�)!�h)/��ȓzc(ĸ5�m�� �%�բ��ȓk�ܽZŔ-*�
$�p,�_$���^�j�#��GbQ	��X�g�P�ȓt��5�BO�($T%�2<�<�ȓDEl�E�H#(��;dF-�ȓ!���@��	A]�Q.�4b���k~2�O�E���2��Z�Lmp�^-�y��Ph܅ˁ��7Y�r0��#�y�ǻ
�.TQc�[$MX�YPWđ+�yB�������D@8I�&B�yrcH�,<ɖ@�;>\�0���U��yr��>J����>�ڰ"��?�y���:2Ӕ�UD=�Ы����y"H��~�z�8��R��C� �?��'�azrb��9�f�	�ET����-�y�j�d68�H�-
	`U� su Љ�y�h^U|,U�U[��D!Uɝ<�y��55�:$Q"FnE���y�LU�S�h�i7"�-hwR�[UL�ym�;D��1�N�]x�'商��xB�� 7�4�Q&��n���r��P�!�D�;p-�	;�i�*e:�٪��L��ўX��'+�hHEn�.�8ـ`	�{.B�2H��co	` �q!F�H.	
�C�ɎJ��X�Ȅ���Bk��
��C�	'f7�1EcN�e�VLKǍE�B�	%Y��S�G�BN0x3��qxC��F�!�\,1U��H�@��%bC���*�q��'"��hh���"fC�I�"��c& F�q����J�l��B�	�xXAm�n��qBV�n��C�	�?�pǃ�-�,�A畗i�C䉆-�Z�)��[.�<(�Tf�B���~;gWO, �e���8C�I�w����e��1�.a ����/�xC�)� �����oM�	�(�3y�L:��$�Ov����4��M0�$X;Tܐ� �m!�V�7#��1�h�_@|����a�!�������n$r�R�-�9r�!��/|��4�3d��#4 ���Ky�	�'�P��Q�ɎfX��dG+t���'.n5j"N
�'���'ދ9�����'9X��H�wad=b"̖�{��=	M>i���'�	�R+�$C��Z.j�7�܏"^C䉟= ��RC-Kp5<H�S!�0,��B�I�1�:MYv �#z����Y#��B�I	<,��hd�2^�E"�Wi�B�	�
[�٘4�P!*��5�TB��DאB�ɨJ�.�;��,���Ē3;Q�B�	/��X��l�(K�$��(Hq4�4��0�%ȇ@X��j�x���T%C�ɏ��H�e�6�4(#�dY�+��B�ɼ��D�@b�tbpL�7�C䉺WU���EB�{�j�)0zC䉲,>� ���C�:�Y�U0xNbC䉊0<�9�ʀ5k!���R"!��B��*u��F�-X��Jr�\�B�	8f�f��*�#M����.�jB�I !ƀ��OI�%���R����;��B�(��A����G���[�!��5� C�II`��c�+0�`�`�Z�C�	��� 2���:��� V�WtB�V��q`�/��7����
�Gf.C�ɚF�X��(�����K�M�㟔���5\�^H�Ə�~d����p��B�ISH���98��8g��}�B�	���i��ܪU���1.PF�ZC�I8���s���&֞i�)͛P�lB�	�xH\�0�.��Vˀ�	hM��
B�I%W���V���	j��#�B�ɱv�d<�0N]-G�]re*�)q>B�9@ �A���&7ܴ��	�
E& B�	�Y��wM[8]o�`B�O�>'@C�ɮs�=;e΍�{���@'c�� C䉳h��!b
Vy���y�MBK�:C�I+8U��(�`��?q���̞3����Ĺ<ir�Ͳ8�@��)S� �WHΩ�ybFO������ O�x���K!��'�az�@ɳ?���"@�-|0�X*1���yB
(�f����V�-�0�Õ�yr���E0r���G]E�\��n���y�l�2a��Li`�I�A�����ϐ�y¬ܿ[��1�c�B�хI��yb��,T��M�BN�)�4�k���9�yB��-=�Z�k� 	 ��E��g�8�y��&_ $9A#�h;�R��y�n�
`ٰ��B� ��0!�Ǻ�y��vZ��#��!.���b��"�y��F�"�I�'>�Yxΐ��yboLE$�T2�+�� �
	A�F�	�y.ԝ p�z�.���(���y�A���dE����/*�s�b��yҀ�8'��x	�+��Qإ�@��y�T�qh��A��ۍ>J��'��yR��+z`�$�ϒz{��A����y��L�e	�Hw	O�yR�8����y��,^�j�Q�LS>}ͨ�sC)���y��F+"TJ�
������P!򤊜�a�@-C=p�����o׬V!�� F��Ў� ���"�j��$ѵ"O�D�F�»y��R���`��"O�볇���� ËK��
e"O�EBf΃KqҰ23��5̠��s"OXq��g�� Y(́`��0�2"O��hs�	�����E�K���C�"O�]X�iP�(\8a"ʗ�q��8IA"OPMrҏO�;�=�C)�&���"O0�I4�
�@P��5����"Ob�X�	[�� K�ނT�lp
%"O�t:��y{�<KЈ�P�b�"�"Oz��.Z�UH^�@@H�#*��Y�c"O��c�e�#V�)�%�>t���2v"ORA{A�b�b�*�.@*^ű��Z�<�c�OS@Ma�C«�Ȩ`�Y�<ْ��hټ4�P�'�hӁl�~�<a�m��c"��j@,�09�f~�<�ffN	�V<�CoB(�<(��c e�<�iA��j6��	:�\��Ru�<���s�~��f��i����5�\�<!���#����E�H-���B��}�<�F�ݨyNx����Z��,{#Jv�<�'���UTD�g�@�o�: K��j�<ɷ	� ��5kw��v&Z 	�� \�<�B�'W��Ysh�h��m;"A�m�<�����83wK̬L�r�B��t�<Y�e�q�B��ԃ���ʐ"�G�<q7�V�h�6BQ�v�F�"#��n�<����,v-n���d�p��"Q�Na�<A�Qiv�1����Г�Y_�<�4CL@����ԨW�N:B���D�<�uk̾e�u�Q(�#(֌`�iW}�<1p#�X����T�'�%�,P�<1��bx5��K@�7�L)��%�B�<�Biɭ<|�y�O*�:����N{�<��m5��DI���F�Z#�M�<�Ά���˦"U�Z� ���-�_�<�F�n��s��xJh��#X�<qt`�2(C$X�F(��:3R����~�<)�Y����-ݖx�Z����|�<��D.D�i�(�.?��rev�<a��:�8� 񮅭��i7nr�<���P#$�\1�ʙ���)�m�<�!�.e��굈ءv��ҳ�Ep�<���08޼��N�\�p�spI�F�<���ړo���%O�4_��UM@�<aW��h�l8ģS:<�P���T�<ѦF�3c����ӡdq�0�Z{�<��$7��R�cZQ` �w�w�<QEa
�jf�s`b���Z��E��I�<i�@�l]�
g�O���8[���G�<I��=e�B��Ȓ�B�p����F�<�g �����s��L#(-*���@�<�H��& ��kײ*�z���G�H�<��4qv�ɠ����oC|�<Q��1_P��S#�.4;^K�Bu�<Q���2uGE����$�W&�t�<�r/D"2�A��Ǥ�¥2a�U�<q׋@� �h�%����kתIw�<q�E��:Th!��'l!elѼPy��aM�)'��$N�p���7�4���j��-����A��]S�f�2�^,�ȓl�D���e�e�(�u'�#�̆ȓlNTRF&�H BLR7.W��S�? ��KfO�,ʎ���腯-#*8��"O���]�n�dHQCg+n��dZ�"OzT��;K��T����`��d "O*%��k�n1�A�F�
p j��v"O��)A�5�A���E�h�=��"O�q�D��P�Н4#.xu0U "O~I�PjV�M̞�C˾p�]Æ"Ot�(U�M�~Ͼs���(fq����"O\��+F�}� �Iq��BbH�3�"OҹB�lI71�8ꐁWSzD1U"O���߃3�0���EW�H��ac�"O��+tcǝ�lݘ���u�ޅ*�"O��G<��`"g�̜XtxX�"O���U���0ej�Һxiʴ�a"O���5bX�UP�$�w\$k�"O<mJ�C͕M,����X ��"O%�΅*~Y�=���ԧ V�`"O�싱�\0o�&��?/S	�E"O������Zh�2bB1f@���R"O��#C�Q��#T�V(C"�9a�"O}c"�A6	��ɪD�_��p�2"O@i �����h�T�֠~�3�"Of"7�g��G@}�k"O���!%��b�@X���ߑ" ���"O��i^���c�m��d:qNV$!��>S�m�b�$4th�{c`93!��6�,B�+NqBQ� ��F*!�$E�:�e �D�+$[#d��J !���>D���e��+�&Q��K��l�!򤍇cnĲRN�@6�%�G	��b�!�D�*����EX�* ���I6=m!�d��V��Z�� ��EE��$[!��fw��p7x8��9��W�2!�䌤�v���-K�j��q�$�)x!��FH��EJI�\dq�غK!�	|n0Y�A��&� Q���"-^!�$ڵH�9�&-$�ЄY)RE!��='�%�t"�p�#�_+!9!򄊩8F��FɌ��
�PKZ�2!�ؕ(���7�MP�ܐ���ӲB�!�Գ'>8�4+�)�t�3늜5!��	�L�p�]��`�c�� �!�$ɷp!� G_<�̙*V���R�!�[�r/�C�@�|ͲT��G95�!�܇"��z挔�~�N��f� ��!��F�ɒp��<��F�`�!�Đ�}�i�� Ob�����¹C�!�Dð)W~�%�"��AN��;!��c2�yCl�=�d��KB!�Ď�i���a7l���e��&^�!���5Mf&�s ���\{&�(���'�!��/86qUH�Q`Lp���ͮSv!��~Z�)�2��	e��*F�Ѿ\�!�䘼1�&��*�2����[�8�!�đ�C|pq ��Htt႓͈+E<!��\aT����+/R�/��|����ᆩ;st�� �X45��`�ȓC�8�#���!B#i�c��,Li�y�ȓ��k楐@Z�]0���&{�����@~���g��*��@�K�y�\��L��y��/�G浻vA��i\�e�ȓB|ĳq)��e����E�!֬���V<��c��9Vj\"7�BZ�p��' *����Y"�1"!+M J����S�?  �g۲x_N�kthC=Zc�t��"O,hb��*6�=�t�R60���Q�"O��ᦕ�'��-�nR��zU;�"O�}:W��x=�Q��� �����"O��ţY�%_r`z_'c�`ѡ�"O�5���)H.�W'��-cb"O�dA�%�	-��h�c�p��Y�f"O��1���XF)a��� �Y�w"O���D�  H)�Qm[!>�����'BF�'�6���I-gd�XW&��[,���'\T�g�ޠ@�>�:�a��H����D���G��g�iߘ�h%F��o���� �yr�+NP	�5dQ�`\8Q����M�ĉ$�S��M��m2Bܶ	����}b�܋/Or�<a�E"e�D=B�6d��Q�<��'&�|�Ē�g���[�f��
G������y�O�$��I��@4wJ�f�.�y��T�61I�-Wt�hU0Wȋ��O�#r�AU�B���T퉱8eՐ%O�C�<�E�h���!W�	1���*f�{�<���?Rd�,SQ���$���ǫWy�<��(��_�r��gͅ&X���.�`�<�@��+|�,��o�;_̰42��g�<�(��p*4�@�I��V�l}s�]a�<��� ��|�J��7i@�2�@f�<��]�3���0)�x�:���W�<��n@<M@�I,TB��b^Q�<!���I4�yp�kU+֐��f:T��P�������{�$��c\N`B�
)D���	��X��6:�L�!�&D��Q�F_�uVjDj�*5T*nd�*O"���͆@O�SWhGR�6�b4U��D{�򩙣 �B$�u��j�ukS�_*!�D2J��hW�,A����l˲0�!�$ڟV���A���|O���S����!��9oP�(�g�Q�5 �H��z�!���*U�$j��X�9p�sd��)~�!��8�m�ч q�V��ɭY�!�D�$�8@`��A�qɆ<!5� c�1O��=�|�ᄓ�C6Z�K%/�# ��P��j�<��@�ඥ�T��!6ehAS�P�<I'n�Ųq�(�<�b��&i�K�<a�DB�$�\�bʰK���Je��G�<a�����,%%��0Z��B�<�t��nl��Q+�����Z娏H�<qq�W�
$�<�E�O�q3�����]�<�5䝜-iH1�M��IcZ2Q�\�<���'7M4��q煦�
`Zs��^쓸p=Q'\�$�0p�f])x6Ƶ:�f�S�<a��\#bZ�-��Ť��╧�N�<�6��UQ��h%
\�^��庂iNA�<�dk�A:`� �"@� ��Nz�<�b�ՓgkB9� Ǟi ���@���/�S��(��\���M2K�j�Q�$�ȓ#I�`���{��r�o!�X�ȓ ��`OĨ!_��k�S�`�Rm�ȓ4H���,7�p���,ו}2"���	I�6��΋�,i,�y�=m�ꑆ�9��  +K?W���,���fDFzb�Ts�O��운H['3�<@��.Y2����d(�S�Dn�\��aV^�1y �����D)�S�Oɂ5�ˀ�e.=��Ǥ*L.����/Orxye�M3�(L���>:.e�\�\E�'�]�ԅX��%j�1D-�����+��~
� ��y�(\�9���0ep�h�"OR=J��	�T�|�"�
ӛ5�Ri���Iv���i:"Fj�LP?}��K�iZ�1O��=%>]1M��W␍�6`�=�
4r��_:�y	cdt�7ƌ�B
B�8 E��OP"<	K<YQC�b�h�Z�O�5���Z�<�'�֍RY@Y��k���"�$S�'ay�n�*�~�A��l����1�y�g�p2n��v��/�hH
$̛��'��$ ��q�	0Y������ތV[ ���h�?arX#?���S/� �I���
iӺ��p΄. y ���O��(R
�5m�r�CA��/���\���'p1O ���}���s��x��m�^�������y� [�yqgԒQ"H �'L���v"��=%?a�U�Ƽ;�e2W��1с� � `��U�]�jpq�!�xLad��K)�<Q�I6�x�Ș�������M��	����&}�d$q4Tk#A��:��x�HC�hO2��d�;L#�� ��4��E8V��#�qO�6m��ا�+��I�Q3rH�83�]&~���S�"O��A� W���s��/qа�1E���HO��D}���5�h���J���c5�ǫ��O��lc?q#W"g����֎V�V0��:#�<D�tI�	�j�b���B�=OK��Bdkx�4�'D�O�>y�3I�"Ĵ���)��p 0+G?�hOL���ڒK|lQ¨�	Y�Q۷��8u�ay2��3A�ȍ�CL�'����ۼ/C�I=.򼂱F�_"��)�\/�B�	�J�ZS�PR�n)� ,��z?�B�	�#~��)�;m����`N��B�	U��p�1�µ7��)	E���v�'ў�?]:@$�C��]�'�G�h�aX�n%D�l��$�'! �k�fкs�Rk≥���a�'rG�"z�LYa�(��A`~�ؔ`�(?w
C�I+s`C�o��Wڼ
5���	�B�	�$����4'�`�h��L8���c���'�T���J��D ���"[}��x��'Lɫ�픴j',#�(J�b�!��']40Pgʘ�X�цe�k��L<�A�����+�@ s��p�2TE{��'.�iӹ_l飒�lҐE��'sX�� �\$��	�X�a��݀�'��]cpƘ����Y��%Yg����'hz1�7k�-?�2����?Rh�	�'*(|ⷊʆr��ȫR-M=H��x�'�t��"ѝ$�P�A���>��'�V����>f��(2P��
ϸ([�'��PHb@ |�0�@�-u����'<����Z"V^�����U슰q�{�;O���Q���sG��J���b�;sa2�i'�V� 5>F ��J^!ԕ�gK-�y�H�Sd�ś��
Wu@�j�����O�~jQ��(T��P0Kݑ)���	��쟬��� �q����֚i����K�RL��x�pd�0�ܳ �b���&܅�K���"`锗"�\�F��O�b�mZB������AB	z����U��&J�M�mL8�y����{B�ñOy���a�4�yҩ
�d�EڗJ2�x!�P��y�	M�Q,�ڷ(��R�r�C����Mk�'�F�*R�P.@��� j�l�a��Y�D�'�q���K�-�-z�ys�o��d&��u"O�%#ӫ[ ��t�� 3���A�x��Hk���O�XI��I'����t;��+��� .�`ťOl� �C�,.����"O���vb�6S��`��)�*$��[�"O��K�LF�\�Re��hҴf(���Ox˓۰=�΋;i�*mS���\"	��}X���R����Op@I5��Z$�1�皔M�mh�"O�(	ňȩ;2l,$jLдdV1�Ox-����d$]�E��ű�HћybZիܾ�y"#Ϡ^���S�*�o"���ŕ��y�!�@\܁p�C�^�$m(Rk� �y��[�*�ӡkK�Z�Њd���'`a{�$t��p&I�]&8h����y] Aa����E5Om� ��̟�y�-��p�I'C^�R����R8�y�)�'��a���P��.Q��-�t� �ȓ~eиʢd�D�r�p���$��<����=3��L[84X�K�u�Ʌ�Bm�����S)�
u��K��`���>@���AW�T�Ѓ��;+������V�f��Ӈ�4RΘ��V�d%:���B�d�ö×*�ʕ�ȓqr��A�_�f{���^�4���ȓdH��ʣύ/x����M<<i`a��$��m��yax(��Ӯ|�I�ȓ �x����po�dRP�Ģf��]�ȓ
�X\�D�_�� ��,��sn���ȓ5�Q��*V 4I�|���z�
��ȓz� �zphǜ%�����^�\��L��r@���O��{L��t�.,���ȓh��0��(/�r})bC/`Y>؇���9Y���j��I�%ʰ5�:Q�ȓIN��p@�G�hG��tj��8���P����t��z3@�A����
}���j�8v�U=1G�q�*�e6����AԜ�PP��7e�M����&-,��ȓ��� lݟTP��hQ葦h���ȓ/b:�8�e�2i_*�Bl�!@��� !�݈jM�=��1@#M�vOHx��F,F��R �I1������2B��ȓ'��C��#M$$jǋC�Z����#h��"��6,p�lA4)S3gt������G期��,Y�ڀ/����x��8*ƽ�ҋ/Z�@'Q��y��[i�8m��E���1F�J#�y2��t��s���85 ����y�kR�u,�0��Ĭ$����ٰ�yb��1^=������]Ƞ뇍�y­��%A��c!�T M[�\��* #�'T�`����d�4�#⤚�}T9��yǕjYƘp1���u���#�y�E}��5�! �Q�Ȥx"	��yr��2\�T�۶dR�u�D��
�y���#��:2E��Hg$�y��
?``eBŖs341*��@��y2ETJ����T��n����y�f?%	ޥȄ�_�u��`��&���y���|p��D�H�b; ٢�)���y.� ���6i�� �P`1H]�y⢀:�F�:��՛���+E�y�d���Z�ѣ�Fx+Ƒ"�f���yb���*]���킟DӬ�RC���y2���yda������E��?�y"AU ;MR0+�%�^n���@����yB̟��B�ե^#��"�.�yn�"%� R�AD�U���@�_2�yb�[��X\PAGA�Q��X@�G��y
� >�p��8�����/�J�5:�"O (cP��'La�E��R�lʌ�"OΌ�b�Y A��!,γB� B�"O0 #�Q���p��H�-�sC"O�t�L�"�L�t�^&{��(�'���� L�H�a|��`@j\�&P�9����6㕀ΰ=��ӗ�l�2�	�O�<K&�à)z��%ɝw����@"O�y`bJ�17Z��uʑ�O�6����dC'L�l}K�/��Q8�#}a�ڀ$�(p�P�B >��$�Q-�P�<qQ!܊S`i���fǲy�B�$օؑ7I��
C�Q>�Y˂���-�>b=lD��FMAjɅȓR Q��%��X�xĪ���9D�j�)%�ДV�X�φ-H�a{�ϛ&0<���nV^<1ga�?�p=Ia@�e�U�?�Mr̿jL���\�4��}���
u�<9%&jV�D��$'���J�"Gyܓbsz	Q#�*7�nD���i_/10
��RbN��Д0u�TO!�d�'j�� �$����!hY!&�P�a�(6��'�D�D�,O�a`��X�D_H���G)s��c�"O�Q��I�g��ȧ�4BA�-�cj_5)U�(A��J�o�I��	�B�
�V�Au���%��l=b���T����-ǌ�?q��R)8���� ����g	N�<Ⴆ�5=��8YeJ��r^�up�e�J����@�E�;눟�LHu=�@)�7`Ȃ����"O��0�IF�iN�9�G�N�|Ј�"O��u�Iડ��e�b� ��"O@�Ҧ�*G-V�y0dІO���Q�"O�!tm�+C ���ٵWu�c�"O��f���h�"LK� v�l!b"O,�pţ�Q�X% K��j`��q"O�Y!E��4�4)��T��s"O��y7�U��Ș&H�#�@I��"O�l F//lk>m�&ǜ.w����p"O�)�4 �7Hp%0iJ�-�ʬЂ*OD�pG�G~P�#�f�W��-J�'�ּ@R�Q�?~��RCE^(E��x�'��L10ƕ	/�+b��PU��
�'`��1d+N;KL��A�=��B
�'5~��r.<HpP<���ͭ4qH)	�'���QdnO�Kg<ɠ��ݜsfT�R	�'v��p���j_n���J��a��H	�'�-�1�Q.l��Q��!\\jŐ�'A�)�D�y���®P�!SU��' wdJp�V��G؊�����)T��S�'(执I `Jdn��H>j�"���cvC�	Xlz�{�*��Fx ��¥5�H�D�n����
��ҧ(�F|cTe� ]H8��%	r=ӕ"O��Ҧ r���S�^7򪤱Ħ��m���2>���������3�	�L���҆+��M��TI˘u(���DL�bPq��U
3�Ё��鋃 TlP��~cR�c�ݨ����d��<�"�	-N4T̅���)~��(`ק�<'�ٱ�@ʸ�v�O]>aJ��%,h��RC�##e4���'�6#L�5�"A����."� �1�bL����,���B���s�4�~3ąt���S���(3�4�qʂ�y���묍14�MRБ��dd�[����򲬍%!�`1�*p��'����������@:r�@���o<v� �S��;�a}��	�u
�9 �_3/Z�|���b�\�3��//����%)�P}9��'!�z���0(T�X�O�O{Δ���͂�qa ��"����W�?b��
��`M�x�EO|��\>4�C��+#*(��;����?Ա�)OJ��Y�pS��͋i�v��MC�
<�Q*g�>�Yam�,=w�]x���U=D����#���p��-�Ԙ���%P��6g�
Ux1�bo��@"��'�\X��$Řh#v��1EЭy|����D�;OT��v�.Y�aF���Il�x��1�Эzx����9���XCOؕr�nt�q��$c�1�I�F=�^�f$��bJ�#����Ǹ1�� C�Ӫ/��*Q�Ƚ |�#�H�6�&����̠��$\\O��''pƜPN]v��H���(غ�Fz�E��:e^�P� 8f� ����m\f7͌H�? ��"�˷^1X0% �2���Gj�$#�L����"S �_�Q�H�~�'��Z����rRdrP$J�t��Y�4B�,�%n�I�ty�O?5N��9�AX�:�����\coH����υlDt��� ֈ]���Ļ��t���֜y�~P�Z�,��7˖:' ��@R�`.&���m�)z�d�{��.Z<}q&"{��K�0l餅�K�|q���K�hh{0癘z���d�1��}�$A1�2��D	f�r�j��a��=���ͨb|&8ʀ�,E���3v�nƄ*�'��
~�z�Z�t�p�0���DW�y�F� gf��o.@T�mS���O��*r�T���䒕m�(��e�C��-'�dP8�����)����K�H�8�AG;��JR��	���L��91�,D
/*A�ER.k��ϓS�D���⁐7\(�)�L��%-4Z��҂�Q�'2�8���8H�@A!ơ&�0,��=l�Y:tꊰ�2���Ĵ\Y��0BҢBut� 3�;>�LDÅ%�>%4r�'�2$ڨ�c�~RD�N.aH�y�g\Ⱥ�2���(���wą.>Zx�X����?��M$	�,#�P.�U���Ə�p�m�0p��хzb�pѩW�I�(�������5jȉ�/ˈu#���U�J��p<�1>,"��"���k$��J���FI�{N�Y��,أ)%���'�\8{�"��X�m�q��T��ڍ�đ�](f�*��D��A��P"�"��K���4�	�y��17��µkM�bŨ$���y���!wڰ���#(J�$C�yb$�9r� k�+��Q��%�y��R!Q����u�1 j�R�iZ�y��E�U���i���0�4�� 	��y��£P�F�,�-�� �E���yү�l�&�*w���dIB��y��Q;P��`�	�B��Q"��y�Ax6e�P�P1I�w����yBei�p���+�6�!D.\�y��F.B��e� ˮ���X�?i�bԋ^�	xI>E��虆����0�ٕH�6	��>{q!���H��%�ҤR���'���`��I/0�,�r`l�>(��y2��)��lH'&�,j:2���e���p>� /�&�К������'ɝ�t}�Tj^�2��ka
�{��~�EW(�z �V�8Y���(O��-�ֽJ@���T�0Q�̟�`K�þ'� �:u)C�)� �� �'�<�k�K�k�S�O�l��dc�B	K�(mn��aŖOA�PV����p�����Tn#~�ɑ���@�K�����.opb�"��L�5F�-�p=�ƅ_ �X�RӇ��k�F6�[�ڨ�+`�Q�Z`�l��M]
[f�ݻ���d݊Y`���a-�? ~�0E��.�N���AN�,�x�	�8��T�"A��Y�HZ1!�q��U�Ru���ФID�Jg��U~���N+*b�N�y�T>5	2jA6� lao�#���L4�=�HY�*�4�,p@���&�ѕO����4e�ސ)1L5F�X��$�ݎMY�q�A�ɐ��)��XBC��3J��z�aŝp�<]�剕�4�dY,@@!��κB�6�ʔ�2���r1�\C7r������Y:������#�'c $h(��'+Ё
�l[3v����T�>�DiR��2ʶ1c!�ػ#OF}�#i$���O�4���&S�؅xWj�8
5�M�p�U�5ɀExR/jq���'PjI������K�b�'F��X�F+�Z� ��+�eJ�o���� N�1Ĕ���S���ɜe�s�"K
KxUp����B�{�G'd��y�����H�k�O`XpB�MNg��F	G�K�
m��.�v֠�t�b�z,�L��Q�)L��q���	7~ˌ鑕��2O���E�'���FA}B��h�QZ��u�$�+x�^��g^�9�,��K����>�`ةD)4\O�H�uI	�D��i�V�G��L��>�$M��i��g$��")��� 3�iM���e��rMb�P1Jb<�[�'� ����AȀ�B�hH�pA3��>"6����|�C��%iA�J.��c�KD�����̊��U==�����(v<�:�D[�N6@��! �Op�{񂄺8+�;��׏��`���'��0��4[9��'�� 	��z`%!�#ӪJ�q��'O�@KgÜ�j2�3���E�h�8L�,R7�K�	��Ũa�'�h�Cv�b�%v�p`�hX�!�)��-�Zхȓ$���QE(F���"$�<��i�J�O`<����.@򵡑�X�'��	1W�J����P�����δt�B�		T�� ��=V��a#��Z>�Sň��M!�aS	1���S|���U��
��Ȑ�B�yM��X �+�O�ɢ/փ1P� 2�O���
Jp����U
!3rH���Q(����� ���6ŉ�-n�i����Ĝ+����mT��H��Ty|�Z!�8@*���6��J:��R3���k~�qr��]!�6(L���K'n.��ċN,��d��DT"M��	ߦ\vhѸ��ƚ��tx���Mݴ����&5i�)Q遇�!��+Xj��aD���8��)Cv�H�����-L�|-[gt�4a���S��1O�!��\ a���We<���'6��Y�ف��Q[d��y� A�0b!8�2$��h�4G1zA�G��$���+�=��Ȕ�d��D�Q0�<E@+ ��bHU�j�Ц�W	(�*���S,��`nS�8��!;�CO 4`�B�	� öe�����u�/���r̛�S0��ѫ�Z���QL�&Ϯ%*5�#�s��j�	��@��% �In5� D���@�
c&�H+�-[H�$�#@ P�l<�H�BO7BںUД�>����a �T��;�ɚ��0Cv�Z�BO&�s��<C����$B<$W��c��]|����cŤY��M�N��C�h�9�ZD���O:�Z����;LO@x�f,�a�+�l�1MϪę���;����-=#� (♤b��A�ca	nь1��c�Fs<`k���2=��s*7D�<ȰlZ�?)�h:wQ-e����"�����3Bȧr��Bvn�/,�4ؐ,�,��O[�. �?����N�����3���=�!� �%8x�7��J����ۀ�r"Cx_40AQ�l؞��w@�@.��	��F�m��� �,|Ol���@-����ߴQ;��K�&Z1��@rTVh��"��f��f��	s4�^�"��?a ��C,��>�'5E(�!c՘[)v��eY�rYf���XV(౬E�E�lᐡC	.o�쵈E���R�QL>E��'%�a�A9&w�2dS %��H@�'x���FK��i7(�u9��@�'7P� {��c卞�inXq��V�N��ѱ��6D�P�7��l��C�ѥf%���s.!D�D2%B�h�P� �*:%Q �>D�܃@^�0�A9
�� � D�tHtX�=O<�vJ�:h��Ds��;D�t8�I��E�¤����wBt �U�9D��`����f�v�%��Yxۣ�4D�\#���[1�|@Iəy�2�KR5D��)AM��/Ѡ�@�=UL�Hը9D��j�$��Iq: �b]& ��FA7D�(�`
�����wk^�	�ܺR�7D�<�&H�uàe�tA�6�6D��/0D���ׄ��]���f�
�r���)E1D��K5Cև���J��W�-@b\�U$(D�4C�o_�m` 	�!�W�O����H(D�dB0��:h��Ď�gJ��1ԉ<D�X�bʑ]\9��=x^x%�r�=D�x*��A(9gu1�(�%yTF�2tK;D�����D'��M��g^nP�ңD,D������>N�]Q�ú*6���%.D���E!J�A�|�VGA�>4Bu�ri1D���W�3�<4��-��Q{T��&f1D�����5284�1�v�hdk�%D�H!�/�lXk�/�\����<D�Hp��9��e`K!"Q&�#$�<D�� ��˔Tj0Yx��6�$�� 9D�\�@��k��!gU�$��5D���1!H�e�HX�/^���)5D?D��C�jܡ!	.e�����)VtXŮ)D��ۂ�̠��l臆�&M@,H%�;D��@�HѸ4l��3�
 ,24Pq%,D��&�؂L�&�Sv(�+��!i�++D����Ǩg�~��g�
95��e2D��rQ+!�R4��m�>z�<�F(7D���b�s��)�柦���Ǝ)D��Jӭ���Ͱ�I�?i�K�95!�D��nMLRF��<���@�p4!�T�K�*�G�37���6�H�o!�� h��R�ظ�(K�1��p8�"OB�z��1NT�J�(ԍq���"O,IA�8&�
��(
�DR"O�5Ir	4s�4�+�D�8����c"O�]S2�4�<05�H&A0��+�"O�Q���
4��T��Mɢ&�YqF"O�݈��O�!�d�b�[,����"OLi��`E�h�h���+Y�]|���"O��0��ܼf��}3�)N�_��s�'���{�Y7r�a|B��!+���#l?�X��`��=i�mG�I2�@��O��\�I(PɳǗ�/����"On<�"f�>IP��@�Ћ6�d�  K�Y#I�3A�"}�A��$��g�שG;`���.T���wL�k������L�vZ{v	�:|ͰI�fH����$�(�剴LMbM��ɛ�$1�Q�V"J:N��B�ɟ2������&i?zM"ƭH*GS4�9cK_
;B�\�VC�%�='.�;�p�!�Vmq"e�篈E�����ZO��{�����׀�I�>��`剭S=,H&�!D�����(�\i�*G��<����3�ɉ�t����7m!��D���y���,�1
%Kd%�yra��Lc-aw��60����4@�;2P����u���1�|�'��+��܌&!\q��M�sxP���'�@�r��K.4��)�j�h���.ԩ5ʰ�z��>�D��D�}y�m�d�O�1c(�C���X�a{"&z-�ͰA��ΟSpB��m}Z�jW(�IPx��)4D�Ԑt$W�V�fE� �)4n$2D,2�ɄA��M��n�O�8(s'NƝB�`t��B�$|���c�'�&�J�Ϋ�
�P�?$�܈�'���ĭT#j�� �ɽ'��m3�'�4�8�#T|�l�s"�</VLT�'F|�7RK1�� ����5b����'}�D2c�ۀEUT���^�U,��'�@��2��A@-��j ����'�B����
@�м�`ܱ \T��'�p�ҧ�C]{�k��}Kx�#�'ɠe��H�L�Px� 8�2���'=ʝ�c(��!ލ��C�
#�A��'�DR�D�L����o�Jº�3�'����I�,R�L�v��F`���'Xh5z��ӭ7�l�K�$ՋKAh�	�'��E�`��
�5BУ�.�>��'n�@�$R�֔3�H��{���8�''nб�n�$.Z9�R�C���	�'VZ|���=�r��c�ˬDed�`�'65h�D��]�r����� l��'�$, ��$�Y�j�3�ZtX
�'�$��N�4ꔐZ�mP��,��	�'_R�AV�Ոy:@a�`S�{-Np		�'���;AM�yQV��%\=f�L�	�'� ِ��1�e1V&.(
 �s
�'�⽠��'�`�
TĂ�-�v� �'�Z�:��ܿ<a	tC�7�����'5�Q��&�'|�Ȉ����6�,Q�'b@4����.).��� ��Z���I�'R4=b��g�jU���8[^�e��'��TI���	2X�	��E�S�zT��'|J47�A���z@n��C�����'�N�#s�q��t��d�#�N��ߓ|O�1�Ю��y��տX�>T��(ѭN�V� 	��y"@�#��}b�C��L\<����(��'q"-)d�ցo8�dF��よM��c�L�G(��c��̩�y�N� b���#BW�G�ĵ@cd�.|�Zf��/< v����|�'
H�"_� ��(�FΗ�.V�i�N��A��/<\qO�vx!�&��<��t��� W��=q�lPm�њs�ɥK�4��)� l����	j��*B�!����&�&�#�����~ڗ땆'K���C�Ԍ`��0�摸1�ҙ����7.�����/&�O`��q�4!��H,���)rI4#G��3�~r�ְf�X�3b�:_���p�O�!�e��~J�*_�� ��oW�%L�p27�I�'x�#䓼Y��8͓K&Z��  �O�~�ab@,ʐt�bj^cOؐ�m�#L�R��O�CB@�g�gy�� T3���) �B�*��e�_���%*��0� �?�$�U�#�p]" �0�.H��1��'7Ib��SǇK�`��)>v�Y���O�vy\���߇�a�@�F�j6�ܻ�	X���u����x\��Ê���嫇�~�p-�{:*����=>�A�ϋ1�:��ƅ\8��p�6�Oh�yeO
30����$@�9�s2��NU�c����?�@�Q8!n�T�20����t �>y�(�&(���ܛZ%Rػ����B�*DF�:�џ�h�?jB+��'�R�c7FW
>`ʱ��)�F���G�a�6!�S恠�n���Dmy��Ι���$^INQ���x�y�j����I<@P�&]�8���VX��`Dḑn�X躃�==�-B��F<�A��4���ѱ���u
���$ˍYk:��ծ(��d'�ρ"����0*�L�ڢM�q5���	�s5� �KYk�-���$K<l�K��v�a90
OXZ�Npur���7X"l)P7EA������~Ң[-����`��?UP��D~>eF��x,pl R�Oq��+D+=�Oj��@,D^��(��bP4	� ��@���z0n-���-�8:g��"��:2F^�<K��Z�G0��Dl�h�(�Ӹ}�ԅ�0��D3��CfT�5UC�ɓ���(Z'1˂�+�AR#/�B�I,IV�$PW�R!G\���Giŕn��B�I�����V���nZD�Ҁo�@2�B�	�zߤD�2�	��HhAw⁚�lB�I+;�Db��^?RbR����"�|B�	�?\t�a'� h�<�႕~!|B�I1
����)��m�@�k�~B��	���� ��X�!���IRB��BpR�j厯tT�M�RA�7�B䉺}�fH��N68��0RcA�,U�.B�I�~H�ͳ��B�5Ơ,2֧7,'*�d\<
�.�KC,*��b�x��v��qpfЬB%5��C����#=G�,)1���� ��'��)j7�ɐgaXA���F8PV̂+P�R0���ٝ*������eq� S�aрL��|���ΜXfr`� M�7Q
��Q�nN7N?�ȅ��%#cJucp��-j ��p��6j�~�<��(�'&i^]3�h�/o*��P� �!;\�8��5jX�"ۖ��Ýş��5�ӫX�qO?�����3a��0�LŽ���3LK�4\iӦ�
u�@�P���.)����'�l��F��9o�FYjt��pJìO�q�gj�i�|���I�\���8b�HJn�)۳J�Y^�d���!���$ƞ�8���E՟�ɱ9���5E	�]�BQ�d�ˢx��ܘb�2��5C��'�Z����VX"E��h�-[�Ꜫ��X�jE�A�F�T[����O�����X�3�u�%˞���|��Ϝ�>��s1I��W�=j)T�'��Y�u��;��K��N�]�)z*��$ �=��d����4^��&_�B�-�㩍lM�S��?!0
; ��R��p,�։>�4�����)*��0�A�j�ˍA��?��m
yۜm[6 �~�4S�bX{?ɶ�[����;�)8LO�- ��ўQ��<'$�S���IPH� 1?�UꉢsF� �JL�����!��+5|�� L��tR� @�`q 6n��0����8�K˧G'�bbJ�&I��H�ы��
��r4��%�e��'�D �@���L15h3}b
/E!��P)��Z^`����>{Aa�hx�p�cH�:�J���N�.ED��'�J�y�J9)���X��\���9z���'�������H�矜@T�X�R� �*H,��X���9�	,��P��_�Ȋ�*�3RKr1p�?͋$G�FSQs!AՓDpA��>��ڊ���(
דz�t�R�� >` �s���9ٖ�O�TG� Ly�9#��T)ζd��o�
c`��U�F�����w�R��B�	N�t�JvBƏex�I�_ V�ؙل
7}��Ծ����}&� �a��3)U�Qhמt�p�Ba(���$����A*�l5�)2�%bK(pr���8�a~r��;ô��SaS�8N�bt�B��p<���O�H��0U�1?�J��mL}�%�ķC���Q��E�<��d�Dy6hZG��)3߸"��D��J;Q`�mR�^�?��hOL�b?E�� �=8��
��SZ��Ր�l=D�`;�-�oO���T�SG`j�۠��"���N�Hp4ea�=?�b?��O� �QP���',���#���n�&tÔO2U�����2c`����ՊG�U��#�O�T�� ��4"R����3SD�|r@�.}�a1�ĭb�~R+�8�X9I���AeZt(���JeRC
�pz�)D�Ň[<�1p�'��zO�-&�B�Q�L",���,���.��)���{��a-�a�qB��쭡ҡ�
N|�������г��"�Ĵ�v���"@j���|18�&�7@�)2KFZ_@��g�!�'?<I�!u���Bhe�;����y"��%��h0%Ɣ&��`� ύzV`���	�[jHA��(���O?Ͱ��$�>�0j��_0E\�p��y�~b垇e��x $��>@D#��_��t�	F.���p�31xP��N�w��|(r�F0Y讵(�k�hrr�Ҷ� ʓmy
t8""�2_綉H���kxj��FgA!"h�SgY�MN <��!bR"(��C�I#S:�XR��ċ#��񌗗/*0"�Τ�F�����vm��@ U6�pj��$�s�}�0�	�
;`+ּ.<�m���?D��ԭ]�d}���
J)>�t�	��Z�I�̥0G��(�������נ���f{����*��>v� ��m4 �P��SiՃPZ��DE�>�B؀eU�u�H����a�"�'�C�'[�w�L����1���<s6�Q�?LO�P[�BƗAb$$HpeԘh%��Z�n����&�-��\`Р�,�%�f��kj\�(C�
�Mٌ��t�	>�d����'D�����7p�I��-��fGR&�)I2��G�5{�vPzV�0a`����ᒚ��O��ΝO:Г�
L)52��ˡiM�4!�$,D�� N|9�݀�HV(��Ԝ
��P��c^M؞�p��X�th�Ë�U�Ҥ�ť!|O!hUl̈YT�`ڴi����֏Q�Lbؙ3�k�9fĐ�� �䀚��&^F���Ϸ^�B,�?��+�	G,�)�;�'S����D�_�M��E.,���ȓgV���o��a�1"�!A�pv�E R(���N>E��'����)B�B0M�|u�'^�}91�:T�:%����,@z
���'�ԩ�i�d�(�(N�;jb�ɡB�{>�p#5D��y�]D���nкV����.1D��c�!�.�B7B�,Y��	��,D�t��C�J'0R'�΂O^t�8� +D�pp�d�:�FL=9'�s��*D��g�Q�>�iɗ�̍65���`&D��XR��m�LQ� 4F�tɡ-$D�h:��C��.d��b�P�Ȣ��%D�p����fȲ=��%�A�88�@H.D�c0n;Ps>pi�e��wj���R ,D�܋p�ї7� ]D��${F�-D����/Ƨƨ=���3o�<�ӡ,D�����z�F���n�X��H�&� D�����cǬ}(!��8N(q$!D��*b�/�rI��d��(��� D���%�ͨ(�����A+��㧤0D�,P�/�Qy� �7[I_�$���=D��z��W.'��d����!b)��4D�d��*�����`�f�8��d2�1D�����y\��f_��P���+D��)WL�9�\�@���,���(D�4��]�6�`@��MU8@��� �)D�T�0�M\��$:GF!�N+D��s�"�\��Y��������)D��x�bB�
�Ҕ)�吳����&:�I0���Q�[	 !8��`όeSc��a�� l�T��f�I�,�\Q�(=D�,QC挈IC4d�8m:	��=D�p34��:"�,59qɉ } Mq�,:D���"�JYc�I0bZ���8D��R�$X�?��œ�+φ�y� *D��S�n�g��]�W@E"fN�k�b5D��sUg���*ac�6�.,�D9D� ��["g|p�va�'65��!)��&�O0��;�$��%��@�J;3L�}��q���w�<��'��)t����}��3� �	Cs ]�D3�SA�=C���2�9O�!B$C���|�;dh�<E�d/�
*x��a�E0VPC`�B�G������ٟF�uXS����E�<���a'�mf�D�M6q^�Ã.�w��l1��g�T>�	�kƒJ�䅠� A��Ҡ@
 ��'��ڰ`*�s��s�H��c ��j��9�&�V�!�|Y@4"O��k1g<(^�b�M��-��t��"Oj)��ˁf�d���>^"��w"O�QS�&C�ڄa&���7����"OTٳQAS#>�`�MҾ|H��"OF5�TC�L;XJ0,�Y�B���"OLj���12i��(A1��`�"OP�: �}�4�0�ـ��3"O�tH��-5�EZ�&�)k����"ONeH��ý�Bẖb�RN
@�G"O��xՆD�G�p�i��Id���"Olt�$B����!+a���t"OB�4I�jYbU2&���V"Ov��3�;5R�A
�KȮe�LW"OX�R@��^֌��e
$q���"O�Z��#��Xȵ���c���"O"l�@�_��Nu��"�/��\��"OP��"���C2�c��q�A"O�=a\W ��N�<?d��`"Oz�R͈֮3e�Q�3ΐ
2ZPPd"O*XZG�W�'��1��F(FUd�JW"OR�ە!֙}�FUQ0���$Kր*�"O��B�m��A�ȸbdZ3nq
�"O��I��8��ZGJ	�c  {�"O6|�&ǅ�K� �=\��E"Ot�g�
h�`�r�C)S����"O����	�g��{�K�@�8��"O�Mֶ$� �n\�Di~6���b6!�D�NC�(Q�o�T}�m��(�5!��ϛ&Ҕ�!	��^�C�Ǐ��!�� �׺�k�UyTx��؄w�!�d�>=�eB���<r�Y�vL�7!�D�y�<����RZ�lq7I\M�!�$�765���·F�R���(A��!�TY�aR6|��Q��nɷ�!�dE6v'hԂ��E�ZT��F�o�!�$
�,��кd��kXɲ]�!��/FqR4��](o����RM
�!��R	<�2#�Z�(tn�a#��6`�!�dI6CA�zQ�T�XY���t-��'�!�䏘�h=c��H�u(�	��fOH�!򤎸����a��,m\DK&���!��>��ᙣh�1-�Ңō�w�!��X�(�2u�!nH�$�YE[�!��3H�haz�#��n����w�ã6�!��.Fր���%'7x4Bc���]�!�ކ+�(M:'
�}ÈԫH�Q~!�L*�����VX���Cο{r!�'y3�-*׫ƵM�(�1��d!��PiW�Ms4��6;6�qr'̾\!��4�ݡb�
�].Td��
6U!�$��s�-�5Aȕ]|R���c�kE!�Dȩq��T�P@�)}and ��"/U!�L�^�>qh���q��4�6�[�!���(E�2�S"lG+2�h���ķJ�!��G#d|$�:��${ �!����,�!�P2G��,��i_*Q��ш�A?!�ݪs��cچkV��3�̏�a!�z�XqfR�	�X��끊m�!�$I�2���E�@+N�5P�*J";�!�� b��@��m�$��f��q�"O䈀b�Y,1OTt��!)�t	�p"O0��d!���E�|4�+�"O�,K�1.2�L�`e�xcB�5"O ��@�O->��������RD0�� "O�����[%N��2$D�'�x��"O|Iru�P�'M49y��И:�N!J�"O� (�"^,�1%"î[�j�ô"O�ь�9%��x�� �h?@D��"O0܈�'�ʾq�3��3X��R"O�}�ģ�2t�d 3CęX�:0�2"OJ8:e�P�	2ף�%в���"O����
�:D���Y��q�&"O��h��<6�\�1��i��E�d"O��k7k/�i��N�,y�쭚U"O,P��␲U��Y�U�Q�)�ԁ�"O�=����v $�s�[&@�h�r"O�@�O�8XD<�Fi�7t����U"O�y�fdJ`�  �(ܘ�~�ѧ"O<��2	ޙD]s��Ϸ�bY�"OF̛��(Nb�R%.I�TEKs"O>i���8��A%	�\l:��"OL	�voU4m|2����k]"�"u"O\��v�G�b��)���:TL��"Ob��U�\�,~�jb"Z"k(|�)�"O~,rR�A�YHTu`�`J3~C���"O"	�a^99_��x�Aɭ���9#"Or��	�� C؅X��Ŧ��`v"O���GӁ
u��0���
,�p�RQ"O�y���.(���J'dї ���"OZ$�VXW�R�9d$A��hpB"O�K�.|� -����R] b"O�iE�ă0ۢt���� dR���"OL��ԬQ$(���cRb�=N�<``"O^�Z5G�fX�[��	"���"O��q�
7��];d ڴSX@ a"O^�A1����4��Մ�9� )r"O�,�!�&xA��a�m�����"O ���X+G�X̃s��&'%�Y��"O"�3��l ��QG�43�e�C"O6Y(��=�B`�!�C�\H�Ц"O����H�[��]�l�=�h�J�"O="
�2_����[ǘ���"O��8����c<��d�<w�ޤS�"O���"cۻl����ەn����"O�Lq+� ?8� x�� ����$"O������j����̼@$"O�5��`�*6:QB^�t�1��"O��pu�E;x��0�S��:����"O,iDA04^� �#��(� �"O&�#��W�_��0�Q�ߘ
��X�"O�4��g8N%���!�($�!4"OR��m�5����� K�8�0Y#�"O<�	FM�2&2�S��Z�2n�"O��Cj����W|Ö��1NN��y������yQ��m�Da� 익�yb��"�1����!S�<�yR��!���∘�`����A��yr��(cW匫,�D�S�*�.�yRN֜<�h4��g�:&2���u�C��y䂦6��T;F�ӠI�L[����y�m��Sq@y�l�+sz�g�̀�yR�Z�7��Փq�5x~���֎	�yR A�r��"��ڍG��$� 8�y
� �л��G�~b��������l�g"O&�!e�I����/1��F4D���O�&L\�͑2hg��0S�2D���S�,?Xh:�)ٜ3��*�@0D����@5~<P i3)\HZ�8Ì,D�4Qu��N!����# -c��.D�����պV���l����@�)D��+��4iA0�Z��&C̬�`�+D��`�$,�\�a ��{�  e)D�hh�XBT�DE_�hA��rto1D�da!_�"б�2& :j�e�֢3D�|�3�Ӻ%��.�;j3���b1D�|���M�2���IP�#�-� �0D�����]��p(a�\6?e>� T�,D����Ʌ�j��׀#-g�|�w�5D�D��I�1�n�B��!��4D��rG%ǪRP8j�mޱ]bNpÐ 1D��Y�3��!3���"z�k�!9D����51�I��&Z�T0D�<D��:W�R�j���������#6D���$�B<�oF~+�Y��o3D��s D�l��,ѱ3嬕j�
-D��H@�
�n��3#��Q+�m>D�8�U#��5ξ�x�B��k�#7D�����E.�dK"dĩc��:�4D�|�3��Kk�5@�Ă!&Zʤ�3D�0����0b�#˅�	ܒ�K6�/D�d��!F5�Ue��!dq{�;D�8Q�IML�i� �e32B=D�T[�@�<ls��������5D������"/TSqh��^<���Ub6D�XPT˜�dZܺ�9u:P����5D�<���0N8�@��#�<�h%8D�4����u.���T��x�C5D���' S���8C���4��q��*8D�� �/S�T�r��W5��(�!+D���~<��I�ː�r&�`�4D����gVc
xc&Y�����-?D� �wiV�d<��FE��v����D=D� ���Z 7v���f�"�!x <D�Ⱥf�rj4��԰$�Y�5D�������^�"Ep�+���p5D�0����Kʄ�X�%&3�Б��b4D�c�	�{��m���Ok���Al-D�L�k�>:��LZ���3Ȭ��-'D�h�dդ%TLsE�نw � *�"$D�X�ы9���+l�)5�z�.!D�$��)��~̾P�b"/�}��F)D�̚a�R�(*`�`�V���e:�$D�\ ��*�C�!�]��X@�#D�����	)�x�rc��z���>D��pb%f�f�b!iщ4�Z��� D��zd-9hTp�1"0!9$+3D�d�̈7s\��D:��!O/D�Sr��
i��H�5@�5M���T�?D��9R���jt���M�Q��)xW(3D�HA�@�:dpę
���M�ص��K0D��f%�$2֠�kQEK�n����,<D����/���B
<1G����B8D�l� �Z2���w��8@)s��6D��&)�,@bLaX���,�PF!D�P�D��� pf���'[&C�I����q�dS�j�A��ϛ�9!C�ɧ=E��D��'�(s��XvDB�)� ,$yë�\�1cb�ъQ�&�9s"O�!օ�6"�8+���L\�+�"O�{d�� w�>-*��1?1�ԛ�"O���%��<�f��ǅ$xy�E"O��+4O5=l�IÖ� N��C"O����9/��y����I�`Б"O�E��!eS��
�$�!�Ѹ*O(���{�*�8QkY)c�0���'�t]�h�y��40Q���[��)#�'°8#�ٖ#�������q�'���I���$��"b�Ž��P�'�Z��&� �x���QCL�5�f)b�'���FP=\�dy@�86�|m��'"����=z��ҷMQ0y��
�'�T�,YM[(uS���.搹�'-�10��
p2�!6�L#+�И�'%� �7��nݞt-�.�� �'
�L�Ib3���P� ��	z�'B0Q��$=\��'�X�=��"�'��<��WEDL�q���sPL��'���J  ���   �  ?  �  �  �)  #5  {@  oK  �V  \b  �m  �x  b�  �  �  w�  ��  �  Y�  ��  �  7�  ��  ��  [�  ��  Y�  ��  �  y�  ��     � � � b R& �- )5 ? %G �M �S 2Z 3\  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6-\�c
�<4�d5h��'�B�'���'	�'/�'�B�'���k'�M�=��Y�A�D�S��܃��'���'�b�'���'�"�'�b�'�t�"���#H( �TQ)G��ڟ���ğl�Iԟ��I˟d���x�	؟�QH��&
ga%@B�Z��[�$���<�I�	ӟD���������5i /;N`��M`�
$��J��	���	�������ß���4��$04��)�¢�6���N��|��埬��������p��ٟ�����D{ ��n��0��/�'j��: *]�l�I̟����8��ן��I꟔����T9���Y�`��DI ªK���韴��ퟨ����	ڟ���ٟ$�I럌aF��sk��C�cV��p��ɟ��I����I����I��(�����I˟�������H���-�^�rA��Ɵ���ɟ����p�Iٟ��I蟀�Iğ�yD� XCbE#!�0�� �����Iϟ��	͟�	�������������Ɍ|��Q�C�%����A��)n ���	؟�Iʟ��	�����㟐�	������Pӧᑘ �􁣃�ȴ1������|���X�	����	��|�۴�?���4_J�2���7[��R�Z"Y�VH��U�h�	Qy���O�$n��k8�srʙ�2�<I: *�E�+n���$���=�?��<���=	�(%i�=1�lӏ�$E{F���?����Mc�Ox���M?5�؈1څ�K�*I���կ&���'"�>	q7�S6Ig4|����?UuTip���M�`��F̓��O��6=�|�aAP�B�Ra�"D�?�`�	#d�O���w��ק�O�v�+��i����*���5q=�i�2�);�D~��/�=ͧ�?1���kؙAADX�/�XP�n��<A)O��O0m:H�hb��6�׹^��3&eE�_�Z���Q��#��韰�	�<	�O��b3	�-�>|[&A��0*2�����L��,= � 8�!6擬=!�!V��l���Jׂ��r�^�}�-8�'�Fy�[�(�)��<I!Oz,-s&F�5�t+1j��<ye�il%��OT�l�k��|J��Q�/�7��~������<���?A�U�4���|>���'Gx��*(.P�D�#[P�r��!�d�<ͧ�?9���?A���?a2f9<2*="#Ԭ]aʐ
�1��d�ǦR�(Sǟ���ܟ���͐>.��u�扏���â��:���ǟ��?�|��/M%��ҥÆ6���{B ��y���T�����	���e"�1Cv�O��g"�V�I0B�E[1��R8"0����?	���?�Ӧ�S`y��iӘ(Ѡ�O��11��%o�>�v�¬<L��ˤ?O�]n�f��1���ݟT��ӟ�҃a� �ba�u
;�H�3'#I�P[b|l�S~�Ϝ�$��p�i�'ݿ��H*c���V�W?	��=�R���<9��?����?��?����\�%Ԯ��h�0o�JT���]>d=�I�,K�4/�%�O�68��3}D`d����18Ѕ�TF!&�N�O�D�O�	�7U(f6�8?!�L5^��7N�f�2͸g,�� �
�YAc��&���'��'d��'X��+��ʛS\ 90�N���H��'+�R��ٴV0H���?y����iK(2��[6cC3A⠀PH��S��	&��D�O��$=��?	lNP�Π�fA�/�����J  � i�a[	e���������	R�|�+܁=&�mX�	B^4�pCM�=���'���'���4T�(j�4_��9��h�s,�E�'ғ.�j\R� ؃�?)�;ӛ����t}��'LTMvb�?��3��U�r>rP3�X�,����i�'&�I��_�?Q+gW�P��N�b\âF �>��Au���'=b�'}�'�R�'W�ӂq�^$8�f�Xe��P��'p���x޴Pհ(h���?�����<���y�#�3{���,X�}�VYҔCr���'�ɧ�OE2�B��i���>y2�H0���R٦��g°%��D�	��$
�}$�O���|��p.� ������4��ʈ4/^S���?i��?�(O��oZ�)[���Iş��	�(!�Y�����`���K� ��N\��?I�P����'�p�� �1aݶ�"C$��r���+?�EN�?s��&L�h�';r����?��bG�7��`j ���@�z��_��?���?����?��	�O���#E.E��-���/;�tD����O"Tn��(���IΟD��4���yG�2Z��1Vnޑ��CnV��y��'�B�'�PY�a�iK�I1����ԟ��sbg!.�^X�g��!`ZRD���&��<����?��?1��?��@��_JD1�)҅<H�Յ�����%�q
�ɟ\���&?�ɗxL�8��(� OE;^�qs�O>�D�OޓO1�ĕ�A��`G�=�PϞTn`����<U�pZ��<��EȎi�Z�$.���򤚇Ƕ=�� N2<�Dc��ώ�d�O,�d�O��4��˓� Rg��/�fTʍ@$�ø)t��Za�Q��y|���|)�Oh���O��d4eyH�	T;���hW#�*M�,� C�e���|�h��-9�'��� ����O,VPp�J��Za��9O���O��d�O����O �?`�7m�Mâ㋉=����q��Пl�	��H�ڴ��;*O�dm�E�	K?��
��[=oR!��L	�b���IkyR%ߢ}@�f��T�� ��<8��[f�	6\�~���i� Q7�����'ØD&���'�R�'���'��Y�%$X�A���󂨂A�'B�S�k�42 �t
���?����iH�#�Z ��dO�A�p���0-�	>����O��i%ɧ�I1Ѯ��e��rM�
�(V�%�6A�m҂`I�H{'����'�RN\�I�2<�	0�Ҥ\`"\��M;2%���Iџ�Iݟl�)�SPyR%i��T3S/=��p����U^��8d�X�3���{�F���|}r�'�v�▩��:N�l���C"?
�@V��:E��¦��'�:a�CD��?q rW������|��ؠ�F��(�A����'���'��'s��'>�ӵ�2�x��!��鄡�
�ڝٴ8�r%8���?9����'�?AU��yWg޷a���ah¯U�0áK[�u���'�ɧ�O8�a  �i���u�S�Ko�N]BR�F���^7'%� ��!5�O���|b��>e\��%�UI7N��2�Ƈ �b���?i��?�(OX�mZ{���Iǟ��ɯI���j���p�pP	��ͯl�\��?�]������X%�,�2╜]& {ӆ��a���J�&+?	��J_l@!�4S��O�����?Y��L"4�����c�`8Au � �?����?����?�����O� #�h��@&,��2TrD��0@E�O�Ym�Dm$����޴���yw#ȝlcЄ�6��� ��������y2�'s��'��Q�ұi&�ɯo_v�q�O}���3�ѐ} Xxa1b2u0�caVx�	sy�Of��'���'��	�2uv��i�U���WM�Y��	��M+Cf����O6�?��"��	|J`:3��6ܮ�	q,P?���O4��/��>_N����6Lb��ߒA��A" ��4���~K�Q#'i�O�I>	/O@%���?ې�ȁ�Y�=��F��O����O����O�ɤ<A�i&���2�'�Ic��j���w�GN:\(��'��7>�	�����Of�d�O���P*�-
f�ҁYs6�!R���7�>?�`���k� �)*�����A��f�z��/�J�'�o�L���P�	̟`�	ӟl��������c�E�|!��+��?i��?�E�iehI
[�@�ٴ��=���fm�}�` �eF�C6��K>	���?ͧx�Б�޴������!��2�"����� GjU�!��0p��dS�������O&���Or�DI�&HL�����pZ0�1������$�O�˓j����$��' ^>ej#��=��tʴh�^��m֢4?�Y�l�I֟0$��)���F�(�� ��нZ�y���]��\���A2��4�X}s�ɂ�O0��rJ�8�̠V혇�=Ѷi�O����Oj���O1���T˛&�Ňp@t��G��O.L����;}b6y G�'}2�bӜ�@��OD�d��+������;�<����"?Xʓ4���ݴ��d
k>
���B�� �6I�'J��$�q��cX^A���D�O��$�O����OZ�ļ|2Q�a	���@m�_<%��(�8;l���W�v��'9����'�7=�N	����e�>�x�	A-(EJ"��O��b>`����̓]nr(RY�n!���R�e.  (��y��xe�H��BR�Py��'�b�úa[��[� ��R1���b*R0f!b�'��'�剝�M��)�?���?yG�	a=X�P�B%wr�Hb.��'�N��?���!�y�vB�ft*m��%P "U�'��<۔���^�@lR����IǟDR��'dfPi�Z�z�^!���Q��y���'��'���'/�>����R��7{P�tFT6\ʬ�	,�Mc�IM��?��r+�f�4�JA[���:��i8Ӣ�^��>O��D�O�D��L�.7�(?Y�������)�.Z�J�4eD�=����G��:��(�M>�/O���O����O���OD@k�g�'f���o�>>*�A��<q��iw��I�'�'v�O
��T�\ ˶�r�~�z��"
޲듵?!���D�W$���! WS��aj��@.:p\�`J�ɩ=����'��$���'����	4��y�ѤI���4�?����?����?ͧ���Mئ-1p#��@��(�}z�d�d��N���nv����4��'b���?���?��.H�����QZP����z:�"�4���O�*�L ��@����6�.<<��p��&� ��?J��O��O����OB�2�S�e3j!�j�� rh����FH�j<�	џ���M˶��ϧ�?i�iX�'nB���l�!0�
������xx��|��'@�Ot��RS�i@�	�P�����b܋"�z(��䐈~�v��R@C�<+��b�	^y�O��'OR��?*.�P㬁�O�Bb"`�>TP��'�剌�M�v�Y
�?����?I(����Lĝ0h�`��)C��qyÞ��)�O��d�OT�O��K�|@PPFC�ua��j�b��@��D�H�h�Y�F#?ͧ�`�$�����܍*�+ME�N��@�bҵi��?i��?��S�'��D���:���s7��s(��W>�x�^�B�%�'B\7- �I�����O�a���-Ms*e
�S�l�Ź6h�O���թ- V7�<?�s��M���>� ���d̸CJ4��"f�+t��q�8O���?)���?���?�����'~�zd���.4C����q��nZy�>��՟L��]�'n��w_@�+���3L\L��'�[�@���'���|��d�9P���9O�i���2:��x���h���X�;O�(#�)��?�֩-���<�'�?�5���pe���τ"0��9��.5�?���?�����YҦ��WbQߟ��I��(�`Ż�楚'c̼t*���v�L��x���˟��I|�ɬGg:=��)K���@��b<Ƣ�+)B�3�	�,x���O~�N�O����/� ZT���>@�9��zd�$�O.���O���&ڧ�?�E�U�A��3`᎐:X���f���?�u�i��hr�'�"�`�f��ݴ^��Z����H@�sJ��J��I��	��|�6DP��1�'���Sa�R�?��7�ؒ �#��\�Y�xp)b� Pb�'��i>1�	ʟX������%�tAs6N��\Gd����e$�і'n*7mY7^
�$�O���+�I�O��� P�c=���A��lg�Д
^^}��'=2�|��Daȶ=�XQ17�G�;�
�krm����Կi��k+\�H`���H$�,�'V�$AdJ^�����!��
�©�S�'�2�'!"���4[�D��4-Ch��*B`u⴪�'��јp C�,92q��
������j}2�'��'[&�Cŀѽ	��|� �DҺ��,M0�ƞ�L�2(I�Q>}�],64�)�f��j�2D�Щ������l�I��4�I�x��M��	�qzD�PH��P�1F�Q�԰j��?���ߛvT�V)���M;H>�w���a �}�&��ugέ���?���|�E��M��O���IU���O>p��s�U�V�U3tE�O��KM>9,OP�$�O����O^�y�fPB7��1�ߺRJF b1��Ot��<�@�i�0�[��'��'!�S5�VB�b�T�*����F�2��`��I����I`�)�D� I�� �4�
�]�X`E&FH$� ���S3�<��$[�\y��|�"x���O>(Ȩ�#WH��'���'��tT�x(�4A#0��/Q�k��`��߼���g)�?��2ٛF��v}"�'%6���EE��t��0n�pt��RX��UF��y�'\Tܙ�	�?
�S�$c#�׽'}��ʔ-Á)�J\�Bd�ԗ'��'���'���'{�y�)�h[50 �@Â�[Jh��4-_�i����?I�����<	c��y��
dq��=�4�y N��, b�'�ɧ�O�^�X"�i��P)bup�1�k�W��K��V$�$T�nIh�'��'��i>��I(�dp`C�� I��cp��(?�B���̟�����|�'�6���_]����O��d��kxV�����m<�b�,�A��ț�OV��5�I�o����(���2���4+2�xQ��ه+�8'h\��J~����OV����5}n�ˑ��}�
����G������?I��?���h����9&Y^��a��8�� ��S�s)<�Ēᦁ��Uڟt����M���w�1	��,	)�E�7��6"\4B�'\��'�2�	�TZ�束�;T�Ȕ����"��Q�CX_�I��CZ����O���|����?����?i�O��u9��S.-V��DԈ*O,	l�?8&2��I՟0�	h�՟@����%H���-��Y�(�q�ф����OT�b>��!i��-
hʰF�5�vA����H�B�ty�3w|P�I}��'q�I76�S;$� D�#�;40d��Iß������i>U�'�|6mU�3��$�F�(�4����.Z�i�����Q�?�X�8�Iԟ��q�`��i�)���Pʜ5!���Ri��Q�'ׄ�jsfn�H~���Z� 9��`��=~��"��4"6���?)���?����?����Oz\=[e�h����pz�H���'`��'��7MR�_Q�)�O&dmZr�	(
Z��`P�T*]��p�FLU��&�p�	����f��oZc~"��b������*�J��B�p�H���Pȟԡ2�|�_��Sߟ��I����)E�n�2)�ш:4��V&����Ioy��}�,4X�B�Ov���O��'-��ݒC���'î�A�IƯ$�q�'̄듔?����S���8T���$.ZJ^6�"߲r�QCի˕W���Y�O�)��?I��+�$ޢ���2���Xj��`�5x�����O���O2���<	v�i��sr�âZ\��z��	�G��4��ǻ'C��'a�6m3��8����O�<����^�A��͠w(��Qƺ<ɢk���M��O��0A����R�b�<��F	���.P�\Au,�
TV�͓��$�O���OD��O���|j)K�|�R�
���b�Ry�6"˙���D�%VDr�'���D�'RD6=�pAkEnV�X 3�Þ�O���@�O���%��iV�"�$6mi�8�倌�v(����ˁ+��� �r���a�-�$<��<��?)�K�?h�cCۖy�U˷�	9�?����?�����DϦE�MK�����܂e$͕l3��qS�G,'���N�o��[]���L�?aI�)Tt,<{B�O�Z��@"Rg~ℊ3��PӅ%1��O���I$1����1K� Qp �L6|zE�Z�(+B�'!��'���ߟ��'�u�Hd"�5d�����bF��41޴f~=�.O��oS�Ӽ#���g���S�H�6����F��<y��?Q���R�p޴��d�%~m��I�π (h��%h��4�Y<S2��t�2���<ͧ�?i��?���?1�mQ%u��i���C^��+E�:�������j��x����&?}��B�<�x�D�]�@��ڛ^��+�OT��O֒O1�<�ZЂC8
}���P˟i��u15����� ����bo�BA�_�	zyB��T��7
�pS�����-���'���'H�O/�	��MCs�V�?1r��S��e� ���TS�!l��<I!�i�OT�'	B�'D�-��_�f���I'aä1��:� R��i�	�F�\8���O���$?e���pz|ۃ%�V�!V)�?�(�����I՟|�	ޟd��f�':��`$ސJ���@h�hl���?���$���nL���'|7�)�ā�p����R+���Q���<i1OL��<��>�M��O(�����"��򩂧O�X���Z
Q?���(���Oʓ�?����?��XQT2�o�>�`F�Єw�.Uj���?*O�9oZ�,(]��П�	{����%��]� ��.V�Z�!���$_}��'���|ʟ<�1T�ԙu���b�/6��S��n�\�B�B�5�&��|���O�H�N>Y͌�h�l�1A�ù.1LM��	���?1��?���?�|�(O��oڗt���w+[�;t�A���U�LY"i�ݟp�	6�Mۉ���>��c�<H�¹/ndIc���z���8���?�C��MK�O@<�q���O�\p4,��I��y�5F��i@~�(�'��؟$����8����ID�D�D6Z�ȓ*�U%d�`sE_�6MZ)xZ���O���1���O��mz�	���E�pb�TQƂ؜e��ȕȟ���U�)擯0̀%lZ�<��/"r�0 ��Ƙm>]�3N��<! G)`���5����$�O^�ݑ_b��c��ƿ[[�3��h����O����OF˓WśV�K:-�b�'Kb���ѫև�,N� �! =�O���'Q��'�'z��r�I�Ԫ�"a.����O.�T�L��6m<�	���O�z�̀-<-4���-�!�j@����Oh��O���Oh�}*��O?8dy�f�x���;�'ķ@*̙�D����x��	�M���w/2�a�N?K��]��cM }�R�
�'JB�'5�%��5}�6���XSC8T��4�E1O�r�94�3P�\����z\�'�����d�'���'I��'G��RwK�J�A� �4�f��2P��H�4SC
����?�����<�S%S�V^��5��~�X#s�X�}T�I��t�	[�)���Ö�B�:R�h�)ůeؤ�q@�%lc��_��Is��OҨ�L>Y+O��Fn�iJ�R��%_�d���O���Ov���O�ɷ<Y��i/�� �'Bx,I�̈́z���
�ð/i�T97�'�6m2�� ���O��d�Oy`�f�<1Yn4��D�CI|@�egC�M7�4?����A��	-�S�ߥ�o�K!�b���:D��h �m���	���I͟���ߟh�ʃE£l�)�f�>]��¨��?Q���?D�i��A��Ob(m��O�8�ņG�7�`���#�s����D�)�$�O��4�t�b�|ӆ�$Ṉ���I� (VA����E�����ԙx��$��䓅�4�����O���O�$	He��Q>?�ljǌ�c2��d�Ot�v,�V�����'B]>m���	fn�R��ݬg\!�g�%?A�\� ��Ɵ$��'mx�
W
P
dNb [��K}�X ���/{����dǏ��4�����?ԒO0)��
.���2V�Є6��O���O����O1���h��j�4���J��u|~$��8?��A��'�"�g�|����O������a0P�Il�M+��v����Ot�cփt�>�Ӻ�2��-�z��<	o�iX���	\Q�L����<�.OF���O��d�O����Obʧ7����DS� �F]q7�v�Ȥ��i>~�B%�'��'l�O��&x���\�&ٗ.�6MV5�fS� �0�d�O�O1� m��dx�
�Ɋ!xh�Z%(AQ� ���c���	�U�@e�' ��$�H�����'1�P�#]�)u�!��ģi݊�b��'(��'tr_�`(�4os,���?�����R�o�	/�FY�H8U�>�É�"�>Q��?�H>	��G#�Dx;6�8����dǇH~bl�80%���i�1�^�;�'@rA\4 vXPS�j�5�ܥb ���db�'���'�r�ş�����n���yFɃ:2�eZe��ʟ��4k=L}h)OJ�ll�Ӽ�Ujلdb sA�.�N�ؗmF�<I��?���6�:�4���J�I0�a���`��3ǠJ�{���mT+,s���7h(�D�<ͧ�?���?��?iC���{ ��ኲ?a���٢��dMϦ]j#.K矄����L%?��	�"X��b%ES�Mu ���;%g�� �O*�d�OГO1�� �W�ڠT�+t�� } �E ՙ|�Ş�H�'�@.3����A�Ioy���(����P$3*N��[�]���'|r�'��O��ɕ�M�EM�.�?��a�:�h�Z�
:[�:�2%�U��?q�i��OZ��'vb�'��I&R�&	��M+W��	z�! �8�6�&�i>�Ɇ F�l{��OJ�&?9�ݾ ��l���kL� ���ц!R��Ɵ$�I���������\��5y� *6Oկu�DhsK ��r|K��?9��<��F���'h�7�/���Z)@�*�	A�Z�0j�N�G�`�O���O�	�&Sժ6%?�ũ\J�? �%Ń�h��͉�k|� �2�?�&.���<�'�?����?QC�GI�=��b�,�6E�j\�?�����d�����矬�	˟<�O�dأ�lF�Mb��:mV�P��O�d�'�b�'�ɧ�I�:fO����M
JG\}�ƌ
�Eh�R䂈)<���d�ğP���|��Rs���8N94�g��.����	ӟ���ӟ�)�]y��w��xD�՞D��VoO�g@��+AL	FEP˓z����ND}"�'��ʠ���q|�����9a��'h���u������ex�����	-]0���4Ԃv����$����	My��'.R�'��'RU>͑�!�b�q�X�;�I� ���M�t�K�?9��?�K~"��(��wU�L�h��"l���E�8oz� �U�'��|�����7\�f4OМ�Њ��P��u��KԑZ֢�C0Oz���~��|�^�d��ԟ�� l$5��2���������ϟ���ɟ�	}y��d�>��l�<���,]lAs%�B�N��B$��?:9��ʧ>A����'���ߩ<����˛KA|���OV9�.�(�@�*�0����?��O~JR�ôu�s,ȼz���2�L�OX���O���O�}���n��0DD� {�\�C�(3�ĩ���Xh���U+s���'^6�6�i��x�E�c/�a��ռvP�j@�{���	���	� ed}mZ{~Zw,P�z0�OV$�hլ��I�J@h�N�zIP��/�]�hyr�'�B�'��'W�.�7p͞��TP 0�~�z��M�c��I�?�sȝ�<�I�$%?-��7�J���؎o�<!�)�^�,@z�O����O��O1��$Ӑ���z�L�
F��E��$\�l
~6m�{y��7Y�`u������D��K�fٰу�6�����+Y?�?���?���?ͧ��$T�A������l9�$[	.�V\�cσ������֟���4��'(���?Y��?)0E8��)ғ��o�H��bj5h��}s۴��$��T�"Dy�'d�d�� �.�.�<���(��`��gȉ	����O���O����O`�D,�"?�0#���WT�5�5�N��-����ɝ�MwL��|��e��֗|�oU�N
B�r�	4���B�̤*��'�B��� ��0������[ա��D@�M��ȅ[��,�|�H��џrq�|�V��럴��ϟ(hD�]R��f	��5 m1�Οp�	sy��a�L��U��O����O��'���)W��0��)a���i�L�'���?!����S���O�G���#��ϋJn�I������ytk,'������S.���-�D��T�{ �'0\ ��.�j/����O��D�O���)�<ǺiQ6h�M�7=���ǿ<���s��΍1=��'�|6�0�����$�Of�R�
#j�8a c�����[�g�O���ޒBh6�.?��>E�i#���ߛ�J0�p+M#r�u��`X��y�]���	ȟT������	ן�Ow����ˀNX�#1�ϛ=0�s���|����O(�$�O���.��R��ݴ���K�e��&�`��&�<,��������&�b>QApO�������m,2Q$���A���Jߦ`x2����%�0�'y��'��
7�Z?j�U�D�э&�>!�r�'���'�2[���ߴ2r(H���?��a{ąqR���0��F'ϕQ���"���>q����'��u� �P�'O�D���
9��O�<9%&��r5�ZrJ:���?qrj�OZ�9&��&X�t�G�ۊ%(c"ODɚ���'P�
����{�����O��nZ�3����	����ݴ���ywձIi�Ղ��=��@Zw��2�y��'�"�'L�I�Ծil��0"�����ܟj�#�u� �ǦKB��Qǌ/�$�<�������񇒞u��
P-�Y��	)�M�aJ ��?Y���?����J�
LɗM�PF�a6I�hL�꓌?1����ŞdFy8��ߴ;�#��
x
)�FEH+��X*O���̙��?��B �D�<�e���m�d��&��Hzq`�b��Aߴp,��[\� ��C�ZE�8�W"g}�!��7L�6��]S}r�'�r�'.|�Q�@�Y��9b&��4�y��I�=c�Ɣ�tBD��^d�dfVp���}�@B�F���i J��n���I�7G�\�L}ZVT��c?=� �I����ɸ�M#�N _�tk�ʓO昂��?=X�Q3f� ���s,.���O.�4�,@y0�s���9�`|�оf?@Q@	�"���*h���P�uy"��_��P	vJ$�$��jٝS�����4B�k��?�����gp�\0�I�,��8�'J�?Oe��3��D�O���-��?y)" E���p�?`I���Ǘ"BR�CVO�֦��+O�]��~ғ|"��f����ڄ$��i;�dն�x"k~��� l\PDQ����y��]��H���$�Oro�u���	ȟ���j�@��(���U�����I�#�4=mJ~Zw��x
��O�u�'|�E�$lD�_�0xC��W_��ٙ'��I����I۟��I�,��S�4���	�����^�e$,<�%BQ�(s�6�6q
���OR�$(�S��M�;b�8h�J�at�d�!/V�!�¡0������OR�r0�i��� �s�E�7.�bFc��%�:�w;O^��ϫ�?q��:��<����?Y L��D��`ʰǓp<�`A���?���?Y���DR�r�i�����ğD��ˋa���&Ą��v�b���t�-����?a�a�e�0�X_a|l��iE�7���u�2����Fo� O~�7j�O�h��LCN\x� >e�`1B!�݊_����?���?a��h�6�d�#=f�`"��&C��T�%��0���PǦyzq�Wy�k��杘1�L�2e�.{�Ÿ@�P�,���	ӟ`�'�)c�i��	��ے�O�L�U��iQh�S�ωF*�L��"�\�	Iy2�'��'b�'P��O.MΪ-[F@�#
��+ёJI�	�M��n��?i���?yH~r��^l<(��C�zBv �f-(d�4��V���	Q�S�'b9���Ĉ��t��V(6-Lj��ġu�"<�*Oڴ�1�̎�?�� "��<�c�ʋ��y�ʋ��Z�����?i��?a��?�'�����y�l�ܟ���瑯uo�僱�C�ܬ��ޟ�Pߴ��'����?Y/OJL`7bM���E�9p�m�Yxn6m*?��X���O�X'?������SL�*��iBA#Y���ϟl�I���Iן���h�'c������U�F��������"���?	�g�����$�'n7m&��E�)s3�۷��*Ύ�u���O����O�IV��V7�#?��C[�=����o:
�Y�H���<-r3��O�N>y+O󹊛��':rfE�}�f	���A�2�R���b�*MW��'>�	��M�p�>�?����?Y)��Ep�.Z�?�(���˜H�J����0[�O
���O��O�ӿ,A��C�O�x�BD��m۔&z2��AP�2.�l���;?�'dV���7��l�.\���S�l�!ŊK�:A��r��?���?!�Ş��$����Jp��'��� �%،\�H���k 1���	ɟ���4��'?r��?!f�;4�.��ڒ)�湘d9�?a��X�L� ٴ����co�Ř������D}�u�b�M�P�֡�9)9r�	fyR�'�"�'��'�]>ف��נm��\��I�/�Ise���?I��Ey��'s񟢼nzޙr�	�%q�J�x��B�*�� 2)����	J�)��7)B@m��<y`镎p�x�&��,L�ȱ��G�<w��o��䊜����4��������b�P�B� �F
�l����Ox�D�O��@���e�-e���'�*H>E8@0[��(lr=[҇�i��O���'X��'d�'��sS��w�`�!�'A�d�L���ON��B@ܾ@�&��A�	���?�A��O��gM�+;~@U�2&�s��e�t�Ol�d�O*���O~�}���E���D�����@��H��R��|��'�6�5�iލ��̔?�@�*���-�V���a��������	"Yf�dlZV~2F���y��1S&NݪwA
' �Hk�H;���3q�|�X��ß����x��ϟ,�*N:6�pXդ�d9p����cy��p�$0���O���O4���d
�z�@��S�O�^�������T��U�'>�'ɧ�OiN��'�Dތ��Ł�a�<�Ia��N�f�<I�AF
z�d��_�|y"��8�:�7�/R������K�2�'���'��O��	��M�R����?	���-G���R)>Qy���&M�<9d�i[�O�'���'����`����ֻoB��mʗ
��d�i\�ɶ)*�	"ڟғ����ASَ��Hç2&:G`U~����O ���Ob�$�O���+�S�3�@�K& B�j�Vp�S#�e�q����4��9�M#� �|��ԛƞ|�fݖƌxq) �~�VrD�]:l�'�B��d&8�&���Y�a ��.Rk��){��*��5@�q �O.�O���?���?�E/�x�'
�$���S'M�&yp��?�*OT�o��wC>���ԟL�If�� �hŲ@�F#��Iv����`@ �y��'@�ꓧ?����S���qҜM�U��:H��Y�ФyZ0�G��vK���<�'s���IR�ɹ�D���Q?$��Z�,�?���Işx�I����)�Sfyr�aӞ0��I�!�x(*�D�"7���s�#�����O��ow�ϟ��On���U�"Є�i.�=� ػJ�H���O8I�fv�����4�S�?!�'4��9񬝒}5&�c!V*q�`�*�'��IğL�	ܟ��Iܟ���|��ꕟg��Й2C9"9��6��1$�7�%Rl�d�O~�D5�I�O�Qnz޹ٲ�^�Wb)I���`���hp��˟�	R�)��| �n��<��O`�4�6B��?������<	�@e",��_�sy��'�2N�I�nb2e��osF�8s��"��'�'��I��M3� ����d�OH�����Z�l�#��F�:L�8!��4���O\<�'�b�'?�'�h�Y�A�4���C���i��U-��dSS�B��2��_���b����ZŐ�D�]6�s��G!W,�P��ہ"����O6���O���=��S��ѥx�d�!�I� �����?v�iQ0Z6R�'��6-8�4��.�0c�^����w/Ny#Sd��S����O����O�8#n|���Ӻ�Q��b�i*/ 
�����d�����N��Oh˓�?y���?����?ɞO�d��ҩ
�x�-;�
N��&MY*O��lگ6O8��Iҟ@��|�ПxH����ZI�P�D~� wc���D�O��$%���6-�� LiPbK�%�xs -/-�J�@�dӒH�'xxi�tCs?�H>�)O<�PoؼD�ie���de��*��OL���O��D�O�	�<�f�i������'� Ǩů�L�XEC�6(nm���'�X6-1���O ��'T��y牄!G�@�	4I��;��i��)SQ8�Hc�i~�	�L!D)*!؟���4��´�ņ�q`�6�Y�!���O����O����O��D$�S�9����= ��耏��0��'��!f���9�h�dPЦm$� �`h؝54^�+��,h�)+�@�	��i>�J��Rݦ��u�m��T9����8s��;�E�<|�����'�^�&�ؔ'���'K��'�h��t�G^���	�V�`���'��P���ڴt*hJ/OD�d�|:cn�(fYt9�T���BԢ��`�Em~"��>����?qN>�O�n]K�J�dQ�|��c  9�B|���֥t���zv�iG���|��d���$�p8�C�/pP��`T�6�L�#ԟ���ܟ��	�b>��',V7m� oC����\�}�L"��5x��	'��O��$��5�?QuX�L���.��%����ڤu�WF	�l���ҟ����֦��'J"�(�d�wb)O�H�7$�	�F5Y,�\?�,I�=ON��?!��?i���?����¯[C"����	#�FM0P��LLnZ�}�,�	�H��G��t����Kc��.D�v6e��}�y!���^)��'ɧ�O�ZpF�iB�dX&
d=3!�/YU����D~�d�33b����'A�'d�	П0�	OꜬISm߂n㮜���K�l���	ɟL�	ʟ��'�6mnVZ���O���#'s��Qc�`V��N��ff㟄��O�d�O��O��A6�� ;�$e�/x��!♟TL
:�znZ��'u��IݟD�s&K�Ho��R���?4�PAJ�o��� �	������� G��'�8�;'����5�V�\%K�0��b�'�@6m�Yܠ���O2tn�h�ӼC�Q�V~ECTmh�ԈHP���<i��?���`]�4��d+":��O�N0���+�������jBt�Q�|�Z���I���I������$���0[X�����h�P9�FGuyB/{Ӭ�����O����O�����DJ7�����A��pB�A;;��'���'	ɧ�O]� ���H�_�%��(۔#=z�)��Y�}T�,��O~�rQ�3�?	d�+�ħ<)�'M)
GH1s��׍� u�H�?���?���?ͧ�����ڱ��h)@�<����bo�B�t(�w'�֟�ٴ��'�D��?Q���?��`�4����V�dA&�ʐ9��*�4��D��C )���ĸO��#�l�s�fY�2�"1� Db�=p��h�w'_��r�b�X)�vn�g����,-0N\`�`�7d�NU�#7T(X��$f�ȪK��&��A�#�������CΧ���(��X-+18��<)�-)X�l+w���*]'J�3-�V= Eḏx� �x*מk��3S��Hp�������Z�Y�H�99����aǧTS\�A��X��@��V�5ᾕ��DF~������S�e��m\2{�&�_� �t��%S�!��	@` P41Y�H�	Q�%��`��,�Խ��4�?���?� ׺s��I^y2�'���^�4�`+�����®�d��|.�S���N���O���~Ɋ���I2Q�ue��{�"�n��AfnƓ����<9����C�̂�.�j90����kȨ
��t}�7LS���I����ILyb�O;^�ޔ��lA7�e3!��>�taꕁ�>!/O0�D'�d�O2��"4 � Ǟ���f�)-��#C��O��D�O�˓r�^l�<������?�Z!r���k�vI�Ľi���ß�'����ßTHw��e?���)������&��ϝo}��'�'��IK�ݚ������%��4����	,hT�Uc(_���n����%������dCH�蟘�O�)��Ȍg�=����u�t�i]"�'1�I�/��Ub��j���OB��02}di�.�:�������Ov���O �%/�	~"�f��B��hy�d#�ʜY�� Ц��'� ��Պl�n���O��d�|���ET�-=�U��%łB ��ãIͦ��I񟘪�)JS���O7��8�*�4��)'�؎Il���4"߰�ⶶiy��'%B�O�����!B�h�c�̾"�j	�ŒJ<�l��D���?Q��4�'I�i���W?+�t��r̙0�r��j~����O���L�cz���'��	��,�d���B`�	X��8���K�r� Io�M�	bl0e�N|���?���0�r��B#�2DR�m���6�u���M�	�4@�OPʓ�?�K>��l$�xb%��X%4VB%�&2���6@[>d$�@����<��Ey"��,)ș�L��b�:�K�iL��2�<��OR�<�$�<�;c"L`�B��ä�3f��)Y��n�'}�'2T�<y� �$����@�+�Ъ���c��m`d�J����O��#��<ͧ�?!qœ�EEr�
Q��3n�XUhU��k%�	ȟ���X�'ܐqF�9�IQ�,�2i�q���|Cl,���aK�lZ���%������'��b�B�	!/�BY1U��&��tl�(�	hyRŐ�zI�����k�G?n� �V�;N�mI㎚�
�'v�	Ο���W�s���'�1�W�G�;���� �5V ��?�w���?1���?����)O�ߘu���PN^%7�%�ѭ�'Vț��'�	2r�"<%>�J%�K=FW�BT�9ұ�"�wӔlxՈ�O����O��D��S�4�+� ~���[� �sk���X�$���/�S�'�?!ԨD��A�4,ӆ7ʛ�+��6��O4���O���C�]�i>��IR?��[��)�F��`4I��ۦ��Ir��.������Ib?	�/T(Zy�����HD+�{:���'�X<��[��ө�㟀
�$�*֐��ˌ i�>�)�����ē>-��'�b�'HV��r��>l��)�q
���H�i��H�N<��?�H>	,O���/w��y	5�Ω�ԣ���}��&�'��՟��	��,�'dF��1�v>I���Z� �bq㝵[l �!@
�>1���?yK>9(O�I�Oj\I�<Y.�҉G�K����T�{}R�'o��'o��)78Q�N|�%/B�O��
4 �+(Lآ��Aϛ��'��'1�i>��In�IK5��!pE"#^ ��#�^�g��v�'��[����� ��'�?i��#sed;��c��)vh}�c�g�	_y��'����u��@�4�v�:��,�̭��O˲r��<�
ֹ����~:��j����2�j$W��##B�{����c�n�R˓�?���6w�O1��M��Ŀ>��\����u���u	Qݦ��uB���H��ڟ(�I�?����Ŀ �]�����&"`<
���;��p�'�:���ᓾ+Z04��J!b"�sdnY�!��qߴ�?����?�W@T���?��OfPJ�L�'_�P(S���&�1�A��Z�'�v����O6�M3W��������)�Q�ϸW�<Mm��� ;@�ۅ���|���Ӻ��n�.Sw�i��-B⨼�w �Y�Iϟ�%��IZy�'���9�\;�|��
üj��d����#��� ��v���?��'��	�&��X5���4��Hڴ&���'J��'k�S������1�����18��Ĕ��\eh�m�&��$�O\�D#��<�'�?	7��$��|�1lơ)��m�����^���ϟx��ɟ�'��1��;�i�,F���iC&sҔ�5���K��@n�џ`$�����D�'I�e!�͒�lZ
X�!JFL�C��l��$�	}y2N$`���d�klK�2t9W��_�L�Y�N�$z��'��������r�s��]:Pj"i����A$8|���@�z�L��?a����?��?y���)O�ĜX�H<[�C�G.�\���\C��'*��8�#<%>e���Z0K��=6��; m�,��oeӼ��w	����Iٟ����?�;�O�ʓ+ծ�[��&$��i`W;s��kC�i�� �'Lr^������Tj�����W�� /	򚙄��٦�����	�y��!�O^˓�?��'��
�	��;T<�'�;�����OF�F����d�'mb�'����>Y�1p�Ҍ>:hDb#�}���$��\^T�'*�	���'+ZcFF������*����l;�O��
V:OZ��?�����<��E���N�?�bE��O
�c�(q�O�T9�IMyB�'��	͟�I��̱��F��{�嘗 y��B�u	����|������Iџ��' �Y�}>a�@�=r°�^2� l�Tjz���?,O�D�O��D�f���]�@ᐃT4D�8@S榖$4�� �'���'��V�0�`����	�O�@%�Fb8L���%�<�,E�5��Cy��'(��'�����ܴ-Bd���ޙ@�,��bm� �n�ş,��eyj��4��?������Z1>���skĻy2����ۓ+��Iܟ��I柴C�i���	|yB՟������,c6!�.�EX���i��I�l��P�ڴ�?����?��'VX�i�IX#bV�S�<�$�4��!3r�t�F���O8Q�3Oh���y�)�
EjY����)`�ԁ�J���eU�KX6M�O����O��	�K}]��R���X��5NMy.Ds!(��Ms ��<�I>���t�'�:�����DH԰��Ҙv�LL���x����O��H3�b�'H�Iɟ��<�>�h��[�6�|Ah�a\'��'�������|:��?��O8Z��P�'T��y��W�N�N|r׺ibj̱9�X�����OH˓�?�1[Ƞ������)��IN�n,��'/�-��'qB�'���'�W�`P�X]�x�����| 2fM	�,��ʭO@ʓ�?�,OB�$�O��ڡҴ�Xv
�@�jX�e���hq�<O*���O����O����<1�B�6.�)
N܌[T%�>���u�J�/�FY�t�IjyR�'���'9h���'��P�g�h��lA7���2�	b�����O����O0˓wv^H�P?A�i�]�!Ǆ�*5�	s����b�&�D�<����?���/`�͓��i0Xd��C�A��J�(M3X���:ش�?�����$�1?-b\�O���'����¤ ˜Y�B�S~x81����yn�듲?���?�g�_�<i+�����?q��F��*T�x#��q�*q�� }��ʓaBd��b�i<�'U��O�*�Ӻ3 cB�!|}��E�G:4����I���1I"?�(Ob�>Ub�j��4�@AI�e���Tc�:01��EƦ��	ğP�I�?QӨO0�J{T�)1�]�.�@,sC[��D<ғ�if|�9�OT���O@�`��/�NI��O-]� 0��쒷y�6M�O��D�O�X�$ �R}�_����d?�U��&q2�!�%a��X��@�W��Φ�%�T
աg��'�?����?1����mGHT�Q	]�0d��kC:-���'�Du�l�>�+Ot��<���� �P�"��o"4�J�A���� �i�ݢ�y��'��'G�'剷Z�I�El���t��0H�YM�LçN�
����<������O��d�O�=PtC�-g@��b��>�@Hs�h> ;���O,�$�O��ON�T��-Z�?��M����( ��Ժ��Z M��]I��i7�՟$�'6�'Wk҇�yBC�,g�B�j4Iߐx�K	�[zPe2�i�b�'�2�'A�ɨo1��	L|�"L /&�dY�iڤ�.&�/%֛��'z�'K��'�Ms�'A�tfV��Bͳ"��D��,#vllm���	Py2�Ϧ3C��j�d�v�q��[t���C�S-���t��P��ҟ�I5�N��	O��s*�HVi��g�	�r¸�0�J�̦͖'x�\F�gӬ��O���O�~�?���*�x�ri9���elxl֟ �	�l˘U�IL�	n�'le�`	G�ɇ�¬����%�H�l�>�JT��4�?����?��6�O�`��&ٺ��IkG�F�e0n�����YI��z��$� ���D���C
-��"%N�"�ց�Ѽi���'�RaP�˜c����v?�PC�L��pऍʿd.�k�ǋڦ�$�܂��k��?1���?Y�`țP���#$�˾P����[(�XW�i�B�}Y�c���	R�i����Զ����S��}���[��>IDP_̓�?Y��?9-O8	�T�;Ty�lz3,��&i�l�wJ�'�X����&�\����g�JP�)2"�~�����,�U:�x�y��'v��'"�	?
�TIۚON�ȕ�P	uN�@�R�B肉�O�D�OؒO�d�O����?O\��E�	=F��!�Y�k�|���h}��'���'��	$6�0J|�pBĚhe�x�&OR�g<⽨fmH�W���'��'��'�����'��M��`�D��0]8{GH4�lAnޟ0��@y��E�}��������`�!IըTp�9$�0}>P<+��y�I����	�[���O�IN���:V��3,�#�l�֎B̦і'�� ��{�F��O���O��"��Z�	J6��us�M�3V1��lZџD�IZ�����t�	wܧ�l����,`�����J�6%�:�l�s�%�ݴ�?���?A����O�l����|�*�2�Fv�(�ZFj��� �@��$��"�aK�H8��wh$!�6K�#;x1P%�i���'�bHR�O����O��	��}�A)�S�F�z�$c�7�=�$���'>a�I柀�I:fv�;�� �NDqw��P�Fوٴ�?�ǉT�O��7���D���� |0�F��/i��T���3
z�|�'�"�'��ݟ�b��4�@�Ǫ��M����G5 �  �'���'��|��'���Ho���2&N�'N��E1fۛB����O���O�˓O#�=� I3��Ieς(�1ʉ-P!Hx!q]�8�	ן��II�G�0��O�����@jA�8 �l� 2H��O����O$�d�O��$N�[h�D�O,�$��oI��G
B�m:Bђ�߉S0�,oZ� $� �	hy�eI+��j��i��ċ�e�^	�&ED�T�Z�l���0��ky���
m��F����i��H��m@P�� Q�J��W(EH�	����	�Y�n#<Q�O���:��ѾX�<�W
̯�~�ٴ���-`��lڕ��I�O���PI~�(Q�1�&i3�%�'e�6����ɋ�M����?A�SJ�'�q���+6�B�r�0�%�	:n"���׹i�Х��w�H���O�������&���	�	��I"+�!�(�Qf�%5c
11�4�jdFx����O�$���V�X�~5Z��a��0���Sۦ��������[Нq�}r�'t�d��J�l�q��Z���䔇Z�O������O����O(a��C�e��殏�<<p)��h�Ȧm�	~.�jH<����?�L>�10�x�-&� ��ğ�9ڠ9h�L�>Q�(Qj��?��?�.O8p���{1R�ȣj�UƎ�J&��&��%$���ݟ�'���ݟDے�#n�Z	�!�
Ӥ�9��{�b����ş�����<�	 
|	�I#nY�Y����0m�f�ҠN�-t�p�4�?1��?9M>9����d/S��L�Vx|QA�/����g������O����O��i-d,�Ғ��o�R1�&G<�$K�h����7M�OB��<��\Wdb?� CG�	^Nd��\�{��ංx�X�d�O ���OD���O����O�����Є):^^�8J�61D���b�i���ĕ'c�,
���`��b ���<)e̐L��T�i^�I�y����4X��S͟����� �kUlt{��FB��Q���j��f�'�����O�>ݣ`���m\���eᑣw��(u�~��J�M����I�����?i@�}r��%9�Ej�+�!7�I[�*��u��7-��jX���r�1��)"@/}��z�	�X ��c��ij��'Lo)rԲO���O����K�3��0�J��#b�c�T��&�	��<�Iȟ0���!)����"iE�tȐ��&��D���	gy��'��'����-	���'�)+�,)��I6�%,���џp��� �'�n���8�����/ Yā**�n��O��$�O&��0�	d�ؒ �?L�v��� �\E��
 ��4��۟�������%�����آ�ԩ/`��C�	�l�Zŋg�ȹ�M���?	�����?-O0�+��� �mk'E�C�f��B
�-�|<��Y��Iߟ4�'�b*Ғs\�ԟ��"Bd�(�-I5 �b�KW
V�M�����?�*OT���x�*�+-�z�)5���|��x�q�%�Mk��?�(Oe���HV�Ɵ,��/-���܎0��X#g��3X� ��I<���?q7�_�'���U6I:�PH7� ��v����&�6Y�0@ADŔ�M˂Q?��	�?���O�Q � F�m!WJ�T6�@ǲi?�'�h���<�Ӓl�t��
Z�-ꑬ�^8,6���3*��O��Dg���<A.�X��FFU�id����S��u[Ջ�G}�*�9�O1����R=���R_��Q/֌"�$l�������!��!���|
���?�u ����J�7kߢqФ��%7r �}���Ϙ']��'S�*W���"�� 'H�����bq�7�s��s��<�#]?=�II�	�?���Y��R&���y6F�JP��IN<Q�Sy~R�'"�'
�I8��A��UT>��u�ݤX\�B珃���'�Ҕ|"�'��K�oDl�Yf��%c!v���"i��yk�y��'���'�ɲ>w�9 �O���iC���	� ؂īK%K�����Ox���O
�Oz���OԓT[��[����/_�B�
u Y
�n�>���?Y���?Y���� ����?Q�$�H�'�\�#�����"Vn%	�i�r�|�'��I�`0O*d��J�;|D��!!C?.G&Yj@�i�'<�I�
/��r��V��Ob�IO�[2H���7���t3=>�oZi�N�>�CM��F���fGB�/h�o�����	�V �h��������<�RyZccz�� �Z�k��9
���S����4�?-O�`�7�)�)ϫ�i�j�
tw&��6��d�R��K��H��'{�=���G3�	�`�1+�1;�'Ɋ�N�v� Q��iG�+�`Ф���{��$��0 �.t���W�0�Y6K�b�p�cj@�7�T��%���o�f���C�"����>�`|�&�+u(lI�����y���q�6I�FA�6,��P�"�0����!a��Q1���X�}�2*��	�d"�J����'�"�'�"�{�e�����'@7����mT�3�楓�FM�l��Y"�CF/��	0�">Ԁ�E�ҿER��8�v��2�<9s��3M(�떇��)����M�#
��3Ф��Xh�A�ö�HO�! ��S�V�(�c6MR O��RƯN��'�ў��?�QH��[����ˈ%kv�qf/{�<����>}�-1�O�I�L����\u̓6_�f�'��I�Y'������Dك �@��XҚآs�G0t��	&�'��:6B�'���\(2���K~5@�	MK[5ɡ�HT��`t�QfM��0����%�&#w�ɑ��O�wM���EF*p8��JB���!s��3O���P�'7�_�(ѱl�Du+r����>�IY�����_�����+*�p=I�J?��hO�	�ئ�K����S��
�>����[���'0ư9d�s���Od˧k��y#�~�P܈t�!>ּx*��A�M�F�`���?ac(�:Fƴ��m�:"��ȟ�'��I�:X�R<)��J.�\���HB���tS��eU�c��X����?�dEY�lR��'6rF�j�ȪA�I��������O���$�'���۟�@�'�A�`i+�$U9$��A-D��	�$�0���Qc�ȉ1O
U�����6ғ0&U��8��y��<*f� �i��'F������0�'8��'��w$��8�֟Dcnh9�,ް*�2- �D�eߴy�'�X�Hg������k���$ŲIR@<�U� &d��ӠY�$��kI� �3�Ğ>(���5JH9I:(�$��d9?i,�����'n�F��%H0hI�F_�F9��'�ֹ��F�N�<jCㅞ��p�O�Gz�O5[����a=yhb�b�I�ak�I�l�0d&hY��)�� ��̟L����u��'�"5�%�ƌH1�\T�V�So$����K2[���jS���q�a|2�X g]:���O7N�@����Ig��RՅO�)�d��"!lO��钀N�z_ܹ@��ƶ3����J�1S��'yF��i�I$@<A'�ԭl��Hk���	:����U�dCU32Μ�<���ie�'_M�Ve�~:��N����b	T��B�D�VШ
���?���,�?�������h1�HR�	  gc`{��i�n@Kў%��OD��ZǓB��UL9P��h-_?�MCR�5OT�$�a�5> ��n`8�L��(�O0��<A��B�j����$��s��]+���c̓�?�ϓOx�pJ�Δ~ު���
Ѵ_
.���0����S)0]vɂs-G�!� |��LˉEP���'�2�M����?a/��%��H�O@�´⏊BY��C�;O�D
�F�O>��M!H]����gE�y��Dm��'����{BZ�D�[Z��,��o��B�>񳭜�%�*��0n4N�V	5iD������1B�e�.iv=� ��G,�i�-�X�� /�����jB|(�1E�'L��{6�6?u!�� Ұ�1
%�҄�O}N�AJ�&&��|z��I&p�J��6�U�=���bk��rdzl
۴�?���?q����\`�r���?���?�;�&��G`ޱ@���+5��'�6!9�yBK�<��<��M�v$*@/ȼQ�����Qܓr5�i��I�V�^P;�D����}�M�oZ��<9�M�ܟ�>�O|�3��G �+�I/X���"O��fm��]p�[FK�Y,.��a��Ɉ�4��Oh]�j�Bl���AS�������h���O��$�O�$�e�d�'��)b}��V�!@bDhSOf���@,�Ob ����	sH4�5�J�4$
�R��ʬY����	sUPpc�X�^8 ����A�X�cf�'�B�'��_�\�Iv�¢pS�I�.��É'�f ��1#����ٳضi�$��\�ڭ�<��T�T�'�L�ʕ�y�v���On�
��out#�@�|�o�O
��E�;7���O����;Y���b��M≹kr\P5cX�l�"ʠ��'\���d�S�lY�!�#����d�(~ze�����Tö�� w��A;��vL�Iǟt��4�?�����|�P� Q59p����3���O��"|*կؑW<�D�Si�\�5�Ҫ�y��X���M3��n��ŋL-.�%��f�8Wi�6�w�'f��JF��d��1�(Ҳ ����'��hӃRU4v4�S�ͦ%!8D��'ז�q$E�?!<����B�H�B� �'T"}�5�͞
�`h���>��+�'����Y��L�KZ�e�¡��'��Ÿd��8#TbKU\2��;
�'g�$	� DR]�,��9T���C	�'Ƕ!+!�I�A4",���D��t��'n�� �J�A%�<�1*f<c�'f����"��x��$j��J�'Mv�QwJ�&m���2 ��I���		�'\��ï�.Z�z�'��E�)�y����8E�pI�2�N�
�Ċ��y2"��w�ҕ�u)��\r0 
eiB��y����uc֕h#'*Y4Jl�T�G�y�W�(��[ �@�B��%Ѥ��;�yreςc�ȥ1s���2��pg�"�y�U`^��D�'#��SƧί�y���Y$l�1jήH�l�h� �y�F���v)���؉<�dIc�*�yb�°fN���J�;�Q rn���y"���U�����?�T�B��Q�y�DT���C�D�vq��05����y"�ʛ-nF�ȰgY�j���T�W��yB��@�3�#� _��[���8�y�dűDy���ȗ1Xq�q�CE��y���7݊ ��+�"p�ձ��з�y��O Z���j �K�_�.D��]�yjP=c`Q��E�.�-0� ��y�&�.�\H������a�e)�-��=Y��$^���R�'D��*��ɭ��,�W@�U|�Dp	�'��]cEg��0��؅#C�R��i�Ҫ[�'%��F��|�O�ҵ��^�Ms�q�f"K?A���'���j�ފZb`"�#�*/��:s+˯����F!}������as�-.��8r�$'m!�D�@|�Pp�A�j�]�3D�3Y�B�'�
����g؞8+oO�gY�X�Sc�=���eM;|O���c
�^ޤk�4"�|��d,NU����-�~S�؄ȓ6����<7�މ�aeDU�z��?�"�]-e%zP+�'?ђ�K��6]uP����K�?Q������� F��-Y# �59�u�'��#=E�$��.S����ą	����ș��Pyb�uzW��4���:` a�<� �Q#��Ԩ� ҷEN d�q��w�<���k��a�ʅ� �l5�t�<� �!y��߹�ʥ��_�
�(��U"O�q5/��0�J,1�χ(�j��f"O��Q$� *[��iI��g�ʴ"O�����]*{)c �?V�f�b�"O�	RF�ҡ���HG�_j��G"O���ס�|c���BZƘ	��"O�P�Dٿ��AQ��-��x�v"O����֧6	�Ջ���L�"O�Uc����m���������"O,!1�̉VhE ����E~�P�&"O⹂ׂ�I�V��AjԲJij��"O0�r�ߧZXl��vk��zs�\�"Ol�{���\MZx�,�/t b��"OB(��a�$^o���uX:2}�"O�KwgÕ��y�g�
Z���a"O>e{a��)s�R�r�
(P��js"O���(�;0��<�qjE3
��2"O�h#`�7���W�Q����"O��y��ł^��q� ,�K =BB"Od8t�	5�̍r$�[?��-I�"OP=	�Oݺvqb5;T��+.���Z�"O�؁F���>���Y�fkJ�f"O~x��ԫ\Z@��)�ZL��!�"O�z3-Ֆv���f��!9N<��'��+�Ar��#Jʾ)8�9q��v�<��m�K�@�t-�8���dŐX�<��:o�Z��!�Ȇ=z�I�tf�P�<��M_ �rSɗ9�P�2�JP�<�Ga		e����H�,Y�I#�bX�!���~ܓb����� ^�&�� �iB[g��ȓg�����0mQ���ԗ�Ą%�P��e�k�S�	�p���&*i�!pg��S�)��q�ƌq!�*c����Q�x$(C`�8W�h�0�c��_�n��N�R�g�Ƀ���Cq�ɔ ��!E�>rbB�ɣVh`��

R%�r��|�@�ˠ�ND��s�(E"hwz1ʣT���Ą�x�S�䉋�Na�yh�nնQ2TE��0<	��Z�����0���N�̩��M[F#H�"��[�a�n����a��у $�ٛ0�|2��Oz�k$�^�$ZuǖT�
����DX�5��mJ����P'E�`��H!(!�әJ���"��7���Y��X&9#���]Ϙ�y�%�X؞�Sç-q� ey�T+�BĝQ�
�Q�B�G�@Ű@#� �\��@���#�"�L�۴)�$`BQ
p�0����pV�A�����&u`� W�.!�-�	Hc&����ƱP0s���#fb��0n�O�l=�013Q�&��O<���K� y�b�ڕ�ؚ8�XY������U���"cE�5{R1���Y��K�:`�Pb��P�n�l���$�N�Y��"B��`F,�5��|���r��\�G%��y��a��(k��)#BՅ��؛�*I�}��l�Ĩ����Z�ta#ub�⅊� �9�OX���-Pta{��V�^�`��b'�)@�(����)}������>m�����ڨiپ��I?e;�/��[,?<�)`U+fOLA�Vf�1/7a��Ƈ8��Z�*a�|��BH�
���:"F�Um"@B��(nt�T�Nx�p�4=B��x#3y�֥0�m'�(S�	�q�	�$L�X�ʈ�]��E��ȷHl~E	րE�
�P�v��=�y§=�d��jA;��*�L�-��dŢB�v�CQ������ÊΡl�>9H	^�Vhi�A�o�!h�"3D�P���U�R�f�H寐TR�1�*�?^)�fV��?AA(U9(b�>�O(�St�L�7?\y�g!��Y��4�TO���?
��P�mV�q�@��@��4��@e�`�R�'���閭�3C�|iS��I�_��E2	ӓ>��P���5z"���(���ϊ+}?�Qbc�\/+DXL�ȓJ�Uc��;U|�)#�G*$���>��y�*�E�ԍ
vdy��ώ�T
����РB��p�G7�OԉR���|�R��6O � N����'�B�ضOC≨u�1"e��R|䕨���	w�C�	�jF���� `Z�����Ə���O���f�Ǎ����O�V�K!(�?{�ə����M���� �]R���h��U��l ��`	���gܓc��dK��L��(κ4�dx���(**tD(5D�C��'��1�	�=c�8��ɭ����4_?@UyR%�*&��"�a(k(bC�	 p��I�oR�;xx��ȸ��C䉃KF~�%��%/W��81AG(EY�B�I�(YFܚc��k��d,tV�A1�,D�Xz���(H� ��Ժ)�>PZ��=D������8#e� ��Vt(`mȭK�ɂx�����4ޖ���'���Jr�\<!���'a�iF`�
�����*�\���5�վI}���6���W�ف%�^��~��������m�(
�����O�軷I��؆1���K�i�`�"22��X�dV�>�(E�T"O$֧
�/����TZ�EX&�Op\��>�`��.�0�0|����49�	;1��;!�R8��P�ȓZ��Hh��'ks
m�� E�Cc8�*�<i4m_E��Ԕ��}���� 	s7G��Ёhā�y��0(�6��BV 	�^EA��ޭs��,��kI��D��Q�,�0lc�e@	o�YБ';lO�,ha�t�1�����jM'b�0��7'Ŕ����Q�r�y'�"��0S����t��GH��F�\)-l(���2��܇ȓh�Ӳ �<,%b�h����/�!�ȓ����U��9�NĘV�I�=��Ԅȓz�x�I�bS�g���
	��ȓ;0�MVCE�;���e�A&G�<��'��YbQ�����uPI�~���ȓO�TT�5V���eڢ*�����x�A��6��A � 
"B`i�ȓQ(V���	Z? <�����Ćȓ@.��0`��mVT,��ߞH�D�ȓ:�U�%�
NjHL֦(%ȴ�ȓ.~���S��Fx�#f�!* f��ȓ"�L�0׎ҡPF�]s$�n^x��ȓP*a��I(���٣[�C��M��Y��p��a�  �G�ѼM��ȓ^��LB`GI:>\���H�;sH����6i�-���(<���CøD�l�ȓe�(ĉǤE4[d�ꅛ�����P$��V#�2\\�4���"L����k����F�4@�Zu'�~b����1�8�B���3p>z}���f~�P��f<<8D�E�2$�52�������ȓ>��}Ӑ+ڄr�Zp�'�8���I�l�1+Am�
>"��è�0w� �x  ߆��Xҳ̈́�.T�B$#4�P�Ǌޫgm� �#�Hy�X(5�4}BG	6
��,��j+�H�;u��`t���5	4i�JߎYc���6#�0"O��Z�Z2YD��0nK�]Qz���Ș�!���aE�	�$���Ƹk�q�O�a&f�#�PI�tK�	;`�j�
O�!SKC;rޤ�u��PF� q�
B�$���L(]ώ-A��
c8��u�(�	�H��m{᧞:
�X��n�
��v�N?u�9�P�t��"��_�
`9Í�%D,� $�2I��,�C���k�8(���^|*�E{bG	8 �.�X�3�N��l��/HH"R��(� ��ȓA��а���+���Q�#wC:��		3(i���a6�S�Op�k���cL�C�T�"O��X�J^�w�4���,��\�X��%V� ���ޱ0�b�#��'�i�CҖE��E˂ㄊ@��)
�r��-I�I!v9x`"������歚�i1�)#O����E�ƴ	`B��yU�%Bq"Oj�A�N#=cX�c���&y��k!򄆢(�	褮�>R�Y�Ո!hd!�$��JLt-����0��g܍Y9!��0�y���V)reu�Ԙ`!!�� �x�A�)9���z�b��;N>�2U"O���i��N"Hd�灋Km��@�"OX<;E �>UiVݲ�@Me@�� "O�Ac#-?	�ȃ�m��8F���"O<�bqF�*�.Q��*��>���i`"O֔  l�#(�E�P)��}��*�"O84���AY"`Ͱ������4"OҴx�m�0�� �H!�r��3"O8�'��-kӦ>��� F"O�E��ç~�xUk@`F�=����"OzX�s��.G�fe�1��A� X�"O����I�a�+ʉ�J�RI�&DX�<���}�T��	͚H_lt�"COn�<1��*Kǀ�Ȅ�U8N9�	Mk�<!����X`�CDg��1�h�r�<q6�:l��o]�q����r�<	3F-[�P0Q��S�� �a @Jt�<q�h��* Bc�X7&�lp��$WJ�<�W�F��a��>���+�ÝJ�<��L�w[��j�aE�d!��bdk�<	����Z]	�O!|&us�Gk�<��Z��x�p��5�@��n�@�<�4�T�!.�H��T�m6Z�q.�|�<���ѭ4� q�NȡO7��S�x�<��H�Oh2�	H�`���C�p�<a�c�q2�AE�I� �@H�<)dh�bV�f�zi�k�����ȓ[��6�H�AX��']1'b�m��~�����G�V���㕨-/𺉆ȓ0&4h��J�!n}������1��ȓ1�,)
ED�HK�X1󀎦i��a��g'(1��R*���� F�|E��H�֜���F�!Dn� ��<��ȓ$:I��O�s�b9h�Ϙ
>��1�ȓ#���QB
�i_R	�M�x0���k�$�	�_�{�3�DL�	pd�ȓ[���)Cg
 Tk.Y��A���ȓDW�8R�'�A��cu���A�إ�ȓ2�B�@�&�Ҝ���B�M�v�ȓ=��,) �[.0m�d�=n�x�ȓ���U�C�K.�}��֠��نȓr�:@���+?����g�,�����(�I�4W���v�_J���ȓ)�� ��̅�l���EV�a���ȓH8����#�4��D�ĩ (H�ȓmD�[h�?�r���F��(&D��ȓ�:�Cd�];~���!V%<0��l���@��֨[Pȼ����ΰ�ȓ=�`2�G�G�.!r�g?���ȓ����wą�_\ڀq����!y�4��_�H�#iضp��Q5��/!�y��rQvԸ�L؂[`�'��*����pj���mޚ^�����dߦOo�1�� <�<2����5!���`�C�	��(K��.8,"�"�L�S�B��"2��˕�M�r���G	�p��C䉴w��@�&
7#���q!Z�B.�C�	<K�0��ɐL���SP��#�C�	?J���2�Jˢ�$x�m�H&B�h~x��Q������	9ZC�ɉs��(��a�,��/@�u�(C�;���P2Z�QC��'@�]��C�	�:2�0"�I����S�(7)�C�Ɉ/�$t��nT�c�vuІD�}V~C�)� ���C�k��xڄ%�7(ά��"Oz,Q�E��`�y�DY:R}@�	"Ox�򳣘�5�բ�D��#KPt��"Oh�`bW�N��QUS+�<�a"O�q(��էOԢ@"a�T!5��`G"O��{�<"�nH 2CZ (:0�u"O�d!W�֦aq�1C{�	��"O~b���l:$Bץt��P�P"O`����>�4�z� [.�%h�"O�x�w��D.��1aHQu��!7"O���C/Z�b����}m�I�"O�i�ֈ�J�2ieO��S2�+ "O�����B\d Ѷ�ƃA�ొ�"O�qЩ��d���B�Rk��IC�"Oʄ��E�dBq��tٲ�Q'"OP��K�Q�0��JF!n[r�a�"Ovq�!Щ#P�Z ��
p4�"O&�[���!6
��f�	-*\��"OĠ2@
]v�y&O�g"��b"O�1v	ޚ+o���B�G�I�E"O�	ʤ/]4��T��/нL����"O��4��+[O���b�j!XC"O J��0_j��A�I�vlP`*E"O>\9��/k�a���^_���"O�x���� *��gǆ
a*`�x$"OB�3��^�fӀdI��Ptn�`�"O0	k��,_Oz���?S-�l� "O�c�D�k=
E�'��;rG�1�"O^K0�G&u�����)	B:�#"O2��P�L�o�`ͥ3>* "O�M�J�sx`وe�^�=6ȭ��'��'L\�� ��4yz\�o��Lq�'�� 2v��d�2�/ $H�R�x�'~ē��FmRd�֢/KFp���'J���s��7�0daSm�,nB�0�'���a�'6�z8���+㞙�	�'�r�'Q�;B��AkQ6NTI)	�'��Q��Ӂ*��K�T�qܸ}��'X qP6
V�D�s�Y�f-�u��'.�(rh�?�) �(S&Z��-�ʓ_pt����Y��P�Ȇ�m��`�#Ռh�T���e��ȓ"L>0����K�>	��.��8��"#�����;|b*�H���xشل�m��$���H�HrP�9 c�[\i�ȓL��h�mBa�j�P��uf����7�"T�&����m�si�I�Bu��dvR�b�]-H�����HK�~KfB��?�%�d���ae�����C�g�B�I@�J̻#L�����dͣx�nC�ɃHC6 ����+��� �h�f2C�	�gl\XI�j��fkz!J�)#"�B��>Q� 1@#�v�  �dǒZ�B�IZz��4�؉�/�*1B�J�EJ��wQ�}@���;+2C�I� n$` 'GZ!ɘU���� ^Db����ɀ�8���P,U96U�E1.��B䉣������Z�.��T��.\0�7m?������;���T�M�u�t��Ѩ1D�H����:�r��g.A�VPZ��L1D��٧��p�������~�x���0D��÷��^L���.��b�	�!/D�(a�01P�6�݈)����-4��kѧ�LS�IՋ]lw �Z��+}�B�)� �\x�%��o��K�I���!(��'*�O��g�	#�`����ө�>4U"O��"�a,5���sEE9>������3�S�v�g_�L���1	J�>�"B�7d��	cO�(��l���ƓDB�I�T�L��K�W@hD[A�Ĕ!V�C�	�pS��A)\��8���-�B䉿Y@���]�F��!��͠%#�C�	���;Eʍ�*�$�"�N��V��C�	��#J��?���P3	ˣx��C�	9% ��W��(�y�lI�a��C䉬L��x�C!�w�6�3'D\^F�B�Ipf8p�c��Rn$�YE�U�?�B�I_x�a�P�.4Q���#��B��tC�����s����ӌ$�B�I�e�A!@o�}��`Ca֖qhC�	� ��$�',�*dY�̋2�I%~fC�	�L�b\{B¡F��p��Z�E��C�d `��b4��M�PC�ɐ)$�x���z�-��KM6C�=x��E �,Sw�D#�e�TC��
;�h�2g�Ȑ#�`�@�Se<JC�� 7j4��'�4����Ҫ��w؂C�	�&`�If� j�Q�D�R�*߀C�	*����J+�d�´f�%Q;|C�B��| �)I�k.�*$,�;IC�
!M���u��,HZ �־O�C�ɥ�D�d��� ��Ӹp`PB�I<n�,���-�T�̃�-�TFB�	��i�3��r�,�6��XtB�	;2�`Ђ�5l�,�h��M�@k�C�	�\t��y�F��<� �*��1G��C�	�%⢉����SC�I�*ǾKp�C�	X��T�&�;�B�2�D�c��C�ɤf���K�!��0�
2nu���7D����n
j����^</�z��Ԏ6D��HT�
H��+�aQ	L��`)D����gR8Bjp	�t@T< i#��*D� `5�5F<}�����t���g�:D��+�Q�Ek捊cA�'E9
a3�.#D�
S��<�p���"�� D�$�5���V|�,BGn��ny"���=D�(��΁�I�'g͉N@ �<D�,��i\;
�J��#�F�*Z)��;D�p�RJ��G����c�!k�N�ф�:D�L�s��)	1�Q'N�!t�A�� :D�,yӆS�fP!gސђ��;D�$� Pvۂ���ݶ|�Rf>D����Jׯ����eF��*-��@7D� 8á0	t�l�D��^���y�f5D�HSǔ-�%pp�/�b�� D�h;ΓH��*��*_XL) a=D��1&x�,b/��7d�}�a�<D���Xoon��Ƣ �H�:H;��4D��3N=,9�XʦD�pr(��b?D�����|@d��S6���>D��T(��RV�X�&��v�0m;B.1��0|�B�& �h5�$A .��I4�][�<iU�\�.@.]qe���>�����`~�'�lj2%Ĭ&�ҥ��B�t�v�P�'ذl���^�L�6����B/hd��'g,u����Qhp�Q ��0��1;�'6���(+S<�YA,�+6��'d\���4���@*�����S��� �!	x��K�	�#:�p�w"O���q"Y�s�@�p��o4\���"O��qm^(m
�$z�S�=�(�A"Op�1JX�?��;LJF�3�"Oj���d	!�.�)cHʾO8L��"O X�P"߼�:$H L4�&"O4�[/=A��p��MN�X&��� "O\(�lE6OtaK�ӚL)����"O@ؙ�%�<�%ɰ>+´��"O�@�c�:�˕���rG��	�"O����
t��Z�ɿ&,��f"Oh�PӆWW�x�K�a3}(0�:D"O��H��Z���rkV\:��v"O�y`r ��)e���b�8J��@��"O�2䀁'$ߘm0�`R]�l|2#"On`��CT�A b����ɒ���Q"Op�F�N�5yhs(IzmJD�"O]j�&H�z#؉�'���KO�%��"O��q̗33��`P`LX0|3��"O�=�®*pJ��$Q<K�8""OV@�qc]�mBq PcX�5ƶ$A�"O��瘲S�2����8��eb"O���ھi�p����R�=���+�"OD1�-5�.�R�獗7}r� "O2� �ՙ !���W	F0mt���"OxxBD��K�\�p�HY:Eb8�1�"OPQ9�m^'L*��9����e�6���"O~�R5f�,_�<ث��� �z ��"O���'�[�P�Y*q�C�[�h�ȑ"OJ�q����Bٲ򧚺Hx�]��"O��7�:"0@aa�&dh`��"Or�C`	 �Q�My3�BT����"O�Eqc��z��ҥ���?I�=�0"Oxlғ,�d��z���T�\x�"O:�����;f�=��@�$�a"O��3�!��Ju��`��o*\�"Ohr@Mݎhv��C���&�B�"O�|��o�pp9���EB�	KR"OJ�@6�$���,��!�v�z$"O����޾�2�o~La��"Oj�3��4m^x%#�)$t�Qz3"O���"�> \�3v�-���a�"Oz�4j�X�l ���C�u(�"O��c񃅇��c��Ʉ:��m�R"Oll �EW�%��Q� �,� aq�"O�es�C�x���CC�=-�B�Ó"O�5��M�M.bl��N' Z�"O��T)]~������\��"O�,�����!kE��; �&�Yr"O����@�MB��X�UZ�"Oܘ���L++��	�'�r�a;
�'�� e�Ԝۤp�o
-iZ�!�'�d�IaI߼P�qV��?2�1�',�Y
�N�	̦H�U������'�d��։]3��a)E��*X� ��'�[����.l<���3\2*p��'�����U���a�#V�ZP��'�f0�2借{����ʒfİ��'s��za`Ҏ^9�<sUb�9\����
�'�T8y��rd�2K� XD���'-d a���9M�P@V'ڟ[C�M��'ۮ	��n�`$����hH�=���3�'Vj̒���%Lcth����a�̹P�'�rhk�L�7�uB-NUC�@z��� ��YA䇼w=j4� �N1��1�"OTB�$%\h��9�e_�I��6"O�3��O��`TJ�I;6=��"O6���H��wU^5K% �Vp�X�"O��'��LI�� �L��>�2"Or�9�OY�TZ|�S��)3>���4"O�I+1嘥4ct!Jt��7VμQE"O�����'��-x֊8P
��"O����DG*/�Fxrt*I���h8""O�0���*j��t)��vzY�`"OL�7B��7����ۉaP�T "O��A��k�
�a-�A>��"O�y2ǫ��i<��
�ƐC�@��0"OH�j��\) ��erAHP?h���PF"O���.�#G��cGu��I�$"ON���%���)����,�i�"OF��6�E����!We�TBq"O��s�%��E��J����X�"Oh�)���!@��]��M�>.n�9B"O�|{ǠQ�@ٚ�S!��,z�cu"Ob�+r�'6��^��y��"O(���S�B����D�g�&<�Q"Ob1H��V,j�� +`��$$�(p��"O�ź���.�D�)t�F�.n�a�V"OΌc� �~J
��V�5��P� "O� �d�љ]�A�R"�9�t�ғ"OB�A�ϙiК�BA]��0�yV"OZ@��b_/��p� 	E�$$�u"OԊ!㚽"5.-qF�:۠��"O�J)"����\�"�e��"O�T��-�$5��Pēw��\�T"O���^�F�t( ��&�����"O^������+�b��`�f`6��E"Ov�2$nXMS~�b��L-U����c"O���)�hA�" �
�d�v"OTt8�(߂AO΍1���4r�x�
w"O� X∐�.w�c"�ӥk��u"O4�+T�@�"�l�2l���8�"O�T��,(z��Pi#˘0^w�8%"O����� k���0j!zh��3"OJ�2�XnX>�iD�o���Q"O�Q� ��]K�%˲H@�� �0"O&� �́������@�L�D) u"OB�{���)��yBq�?��	�"O2�Bf�A��:���/�
C"OZ���tb�������\�֡��"O�1�,����YA�W4f�Ȅ`�"On�q��		�*0X�Kd��+"O��a�k��|@�ӅۤP;#"O�\q���nZ���iB�vk��Ң"O�e�������7iЙ`��yg"O��)ư9�8���ϟ$���d"O:A��	�<	&Y�AF�|< ��"O.��QB�s2l�#�V�zh- �"O��1�S�w�*`�V��]B���"O8�k@埵j
�(Q��\]>1k"O"�5-e�@eѰ��P����"O������CP�SjEU̜2&"O&T�ҩM)�*X�pɛM�m{�"O~��@W� �r���K�!W"O\���c��Y�A�'mZ�Z8��(�"OZ���!ϭ���#.۩id(X�"O����
,]J#�
/yؕs"O�ĻF��%*xl1���|�"���"O� ���	LK�iV�R�A��q�2"O،Zq/�/w�����%H�|�5"OrD��ǅ(WP���������!"O� �jA���"+�yx��"O�h
4�76�Z=����fz$�"Oз'�		?$�Ё�ܚ&터kv"O����N�d�BN��'����"O��Y"N�=Qa��12���"OF��7��+w� J'� ��k�"Oz��&J�t�8Q��Ś��L�1c"OB\8G����1b��te�Թ$"O��j�5v���D$��VN���"O�]b3%}��A6�T'a��\��"O-{���7���8�.�v����D"O�5Xgǈ9:p�L��E�8�0�;�"O(��!h��x��(�e�7����`"Ov i��ڝt5��xw$ث%U$��"OX��J�[��M�`�u`��5"O�P0�'I�]аd��-s��@&"Ox@ju�lA��0p-5>�����"O�b��;;4I�PgK<X�4��|��'�(���� �P� 1�q֌��'���%���� ஍&9�&�i�'$h�(A`��a� !P6>>Z�q�'��hr���
%j\�/(4� ��'��9Ŋ�?  ~�3��� �|K
�'��� �D 4Pd!p�R>s�)�'*)��/�2C_,�E���H��4S���'��I��=6��e��*V�nQ�'1�xc��;�P,�qF��P+j�c�'�>����[?�H�!l �\�'���'��>����
��	�'�"̩5%];e�ARr+R\�U�'�6�9��Ƕˬ��W�;�l��'�� 1"��g��u���=0�VL+O&����7YÐf�84��w�OS!�YnB���`S|�1�2#O�D�!�$ҕZ7���e�׵{^l!�w�L�!�$� r�Еd
�y��y�J��!�]'*4���w�\��
i�ڎ�!�J,:��(�i�K�dLӆ,O!�[.*�B��F�/���H�~T!�䏀o����W(U�i'` R!-!Kp!��Vp#:4�;LVR3]�,�ȓD���#Iόaj�x�uƇ�o�����2i���J^'b�\ك��	 _�؅ȓR
��jP)��"�֦
l����A�r���'��XK4 )���J�ч��`�'�D�q��[�][�$C��H� \܅y.O��� R�NXze_�Oa���P�$!�Ęy�,��L�)���z�+!�d�2ad�����L5�0�S�H+_�!��#��AY��Ɍ'��8��_�!�d�<M����bnӧ{�Ne�f�B�$�!��9=�h� ��m�0�(q����!���Z#�[ëP��aFN8]�!�$αG���R�lL�dǖ��r",T~!���.�ƕ1�C�z��-k����!�^QBa�t�~�2F�J�p�!���:��)bfS�[s�q�w��B�!�$�0�J��7��b���듯�6f!�D�yy�k�f/��5��F>�"�)�<g�8'fRbt��ᆆP����s�'�.�ja��_��ึ�M���{��� 
��0$�)�!�&� �l#�U��"O�F"�9�e�J<;�Mz`"O�]�G^?m����T�Rg,M��"O�9�"Z^N�Qr�E1cde�$"O����ɣ<��KQHͩ2Dy��'�ў"~�G�@�K��ȓ�oݸM۲�$ڬ�yZ
H6�߄(��6ᑞ[lY��	$��h�AQޤ�yp�ȓ�hQ�#qު��DO��"* ąȓ9��)z)�6j$�J�$�g��ȓ02$�fgW�4/�+V�x�p�ȓI�`8-t����EN9)�Uad�C�<I�hN-
�h�(�D�~L��rQ���<0H�+��A���)�����s�<���ZT#��S�+�rQ����k�<at��$���B�"ˢ�q	�h�<��e8-j�j�)/р�{#Jb�<!�Ä(f� ��N�&@d�t,�]�<�BRe�4��fc�W+���G�T�'tax��߆'��-q��W������BԶ�y���I\�ȷ��:?*��RХƶ�y��]5�Cj��8o$pAըB��y"�%d�v�Cň�!\��A+l"�y��K�0�H�(eAG�g@i� Q�yrm��!�����g� 1�>� fF��yr�G�Y ��h�N�&�������y�ɑ����S%�`��.�y2���!��E���К��i��
��y�� ����%� [z�i��<�y2��0(���ɘ?B�e*�m��y��>�����E��V�ć��y�7R!p�ANå
C���[���x�Q,LH%(q��/����a디��	f��(���� \��x��\|�z���"O6�r+Q�1��X��#T����"O������mo�t3�����X"OX<[b�cƶ���h��uO�a��"O�]i C�8��I�iЂsA|ipD"O�4)_26$��Ze�<�`t"OV\H��Dz�)`�-F�-�e�'v�$�t��RG�Ӿe��o��f&!�$�T�.��� ˱P_��[�_�U!�1^� Y���]�tH�i[�&�!�� >c`]�5��zS�`�"cғ�!򤑳Q�n�8��`N���A��+�!�d�eXꁨVN� �@�0��<np!��;t "�.ߪ5�~Hq7J�U]!��L�]��8� �ɘA�:�f��]�!�$�X@�8�S�R�4���#�'�ЕJ�f��j	��r'V*܆ʓv`��w�ڀ/����KǓ�X��@
�y�PF����w ����]9��^�|�����W���f�,�x�ڕ�R��ZQġ��o���� 5:����#dB@p�A�*%�4Q�̣<�	�zV�`��"9l�DZ��)(EdI��2߈��@n�7omQb��$59�ч�p^��Rg���C����@$R}���WNz�"s�Z�0CjyC1ښ �$���$�0`�M{��!õJH��9�ȓ}M*A�$��"���.V �~]�ȓ �bH�b��8A��y6M {�%��n�N,y"lQ�m8�
TF�;M�2\��h?�d�bE.R$�j&�J ����S�? ��$��d8���`��8?�,q*�"O�4��߰ 9��k%
YE�:i��"O��:E��+��AQ	�7#&��uO<�jc�(ȼ9�4��<�zE�QC7D�T��C��vq�PKud�	=��ǭ8D�H�@$�)��Q
�G��k�  .7D��{��)(b@݀��]5e���5J!D�0	f@����ۍv���:d&!D��Z�I�dL�B��&|	r��!D�hSE�1~۴0��mЫ M�	x%B?�∟�p*�K�	���`e�q�� ��;LO�2�#M�4F�	1*��X�X�S"Ox]�gκ2�B��
�x��(I�"O@�S�Ξ�l��U1���8���"O�"Wn�b��Px5IܹK$]2�'���8��J;�((���D�$m��'�f�+�O^�R�F��C�B:H��xKϓ�Od��v�&�^�CFq��r"O�Ȉ��ʜ�d1�4Ƅ�A��w"OĴ�1`�eg�2pF��Kj��"O��(�i��Q��j�E97 �e"Opq�v�Y�v����F��J[�LH�"O��X�ȏ$�@��Y�^zЭ��"Ox5 ����tC��Y��:�������F�OD��u��>CJ��F�_�������hO�G0�cC�C0���B0�[��ȓVٸ 2DÊ/q���ꘂ�@i��"9B	��"
1K��]�P�� R���ȓC����+d�`��DѺ?RT�ȓ�Dt�eD�#G��A׭�?X�h����ԑ�aa��9L4I��N��Q��$��6v�K�o�]6�PR�'˼f���h�'S������z��Ӭ['\���'s��9��	�E�Qx3M�y����'����$L~��h�@����	�'���ueӽ8~u��͜�gX���'�0�Bs�0)1��1b+�� Ո�H�'E@�E_�.��Q�%P��l
�'g�#��Fl�(q��R�S�����&Or�#��/F���d��2�L`�f"OsdƏ�r�}��N�2�d)Yt"O��Q���tYzS�G	+|ʘ�"O�4k�e��m��{��7=c�i!e"O�S'ҵ���`u��vD�a� .D��9�F�j��@S��4܌�A�/D�0*�lD9b���ص�=࡭�Ovʓ��S�O#�٢5<���i�JC,xȬ���"O��2T�L0,���I }�Z0ڰ"O�"BE�8lvV�=;��x��"O�0:��f�P��l�
*J��"O^h[��3d�
�͟f�\�%"O��y%f�R�qʂ�# 6�v"Od9S��[6�"��Q�V�j挝T�'g!�΀~<��Sǅ(_��8�E��<O*!��[�"�µ&����Z�̏R!�D_�>4=��bF �l� �e߯\�!�N�|����r��J�@���9I�!�)��)׬M�]�a�qd��!����3��*�~q�1���4�!��j��Z	�d|��+i/r(c�"O�4Kņ�|��h�k�+^u�����'f!���1������1+�H�I��@&6�!��`�~�)��h�*!�7��!p�!�d�_�n�h�N�+!ƾ+�:!��S�? @����J�b-�ʖ�cQ.A��"Or�;"����p�#6.8����"O���C��9�p�'B��/��b"O��DÎ3?+r��C��8���Y�"Ó .I�}}��C��l��)�R"O��ۀH#OZ\0�ڡY�r���IP>10�LP7�f}��W�k�8���g+D�ٵ/�%�"���!�;.M��k$D�̓OڟO�xT�4���F�,��p�$D�Ԑ#�,�>L'P!�����>D��8���0��xJp���k甄I�)D���%�_#C�؁�ec� S�T-��h%D�b`Jܐ ���@��.p�A��)6D��pEi�'�HI�MB�R<�)�/D�����W:3԰QbZ5��`�g�0D���R�R� ��	��#56����H.D�[�k�X�&��s�ĜY���b �7��!�O�;c��	�T��-Y D؂0'"O��K��E){�A�lҤ'���"O�8y��
-Vl�U��9�b�@"OMCpO�<[t.Q@��ν:��E�"O�M1E.R�{��l����x�
H"O���t�٘)��913	����d�a"OZ(sB�07�F@���Ϟ����"O��f��->*�ȣ-�-�z���"O�QZ"��3�t�E���P��E"O�e�F�)8b%*q�G;G��q�"O
���"R/0+V�X��3^��"O�a��F�G֠s����1"O4 ������"�ӗ7�D�"O"���(HKgnZ"� at�U�"O���@,[��L7A0��g"OL���'�+Hq|,i���2b� �Q�"Of	�/�79�.	s�*��4���H�"O�X��ق,��@8gGػ)��I�"O�����=s;���po˵q��C"O���d�U�z���h� X|�U�'M�ɧ,�i��oN-���S�(�����D2��37%��P�9�� g�Z:�C�I �p�!ˎ]A8��[F�C�	5,a�D�O���< @�LV��C�I2�@�¨Xʖ����]��:�����4��K��i�\�`p!��3����ȓbr8"2�	+u!9P' y��8��O�K�$9a�)�9�@cK�=@_����xph3?�rQ{���9����ȓ-���QP��-�d������ȓ8��Y � *|�}2%#�6'<B,���ty���X�V�\^�"�@��ҿEX��� D�tY&D��g�BKBv$��##)D�ԣ@�ǥp�
	���	�|��'D��a'�6����Jրy��t	��#D��#gO�*X����d�P9r6 ��>D�XPd�0@��4�q��:q �uK�%;D���4JE0o$���-LB��i#�:��蟖(£�< ���I��ؠ)Ej=D�`� f�Eg�bHH>	�{V)D�\yC���NH��G�_�䩲�'D��w�͋y,��.J-������0D���+��B����1j��R�^i�.-D�����O�J�`T�gPM@ҥ%D�� a�ޢVp3#�;,���'�刟0�;d�{<�З�P,oqXa�3"O�b��@1X��  ��	���q"O� Xٳp�I�,`~���fW�z��q�'?1Ob�+d"�#6h AF^ �ر�'�I�x�fܓ��!vj���A�dB�I6Hq~�+!?18Q���̊f��B�I� 4��CʼHuv�B�+�G#B�ɏ'SR��RL�D�`��帞� �'W2�r��(= <r��B?j�X��'��%Y��ۋI>��3G͕@���
�'�Y��&<Ap Щ؝?���*O�����2Z~�*���^f��T��)S!�-w�Б�n�;#	��q�琔�!�$���ő�h�����Z�e�
m�!�$R�'���q��C�:�t%�"m�!��[L��	��
K)i��E��4�!�$�<���&�,=�x�3�G�k��y�ችZ�0����G���E�\�u���$/扂D:���AK�o<���a♜ ��C�I�]?\�A�`>H`�͙�(q�C�;c61ht�U�C̲�8rm�'	���ȓI�]۔�Y��X�-�!g.�<�ȓ)�r ��.0(�Ƙ#�ƀ��'k�5��KJ�
�����c�1�M��I_̓5h��n� E&��Ч_7����"[�1�s��V<hS�D�>�v�ȓH�VeЄ03nԕ����{
l��	I�nج�Ub��)������,����ȓp4���b<����*������ȓwg؜��fB mX�A���p��ȓo<DAj��Y`�(�B��;d虄ȓO��\p^2OD�8����S�͇�\����k֑cͺU�Si܅�ƹ�ȓY���QiΤ;h� 8D���[n݆�I�<����x��@I�h��Q��'Kj�I~�Q�I�*��hj¡�??��0�H2D����K� ?�p,"��Y�#]���N1D��R���lI�VoJ���0�9�O��E#�ݣv(ة0<(�3�
;z�l��ȓg7n8�f���q�H��8v� m�ȓ
��4	�a�2&����l[���ȓy�|1�J�~N=(V�ըE��Յ���uPG¯YXa��q�`0�ȓCL�E���*��10Ҡ�bm�Є�U?�a�g�>JL�q�T�D�����P�'��zV��Q= 0�i -O�$��'��U��b1^T����4L�^t��'�\�Еd�
�X]c�lҮKت�3�'����`�Μ#�4��h��?50��	�'�nxa���%L�=S@�;1p�iz�'�Z����_�è�����#%�,��'���2ƀ�)1����������'�� HP#�<f�0��)�;#�tYc�'����ݲ@D�:��"!X9�'u8�{�^!P]���A_�'��`
�'�)Kt�Z:�0���$�,9�q"O���\(�e���Y ^��@�6"On��GG]`ڌ�� �9�r���"O��A*)
��A��aq�tQ$"O�C�&_(��K��3SFh�R�@E{��I��%j, ��ǘ�KW� cD-�5|JB�ɨ6��p'a�EW��僉.TB�68 %sr��0jy�`%X�F<����I�kAa�$ *v�6� '��#/r�C䉭X��y�t)�DF�3��B�	';��1*3%˽D�$�i�(%ؚ�?a��� �,�rLݭ��e��h]�f6����'J�	* �L�b��:Ѩ�(��J�k�DB�ɘ)��U�����5�n�8V*SfB䉱"�`ɻ� �	�\�%�)���=y���?i��ɗ;�)ӥ臃�4&ͮ!�!�d� ?ډkt� X��ō(�!�D >�DUK�#�ZAiq�
�l�!��.=����P�]��a�u�Vi!�W�x�2b��C��b���FP�Y_!�Ĝ�)/����Fݗb�~@���\2sn!�$��2��ҋU��d�b�%�E�!��&~�Ľ:���9B�B�d��!���f3�X���.аPѡ���!�d�3/��a�C�
�8��PՇ�4�!�/U�t)ɲ��@�fq�ug֧U��{��B� ba8#̔�\�&�g���!��%�Ω+.L�p��]#;�!�[3�xx��,F��a�	�u�!�$�Ke4�j��T��1����/x!���t?�37)�'q3�|qu%I>�!�d�"W�r���ƩE~ՙ�c���!�$ݼA�zl �K�r�4�"D�7S�!�$եm�ܘ`� ߢx�z��CɠF��H��(�"m�[$�@*$R���L $"O( ia��i{���DHF8`�r�d��o>���iڎ}jv���
F����U�1D��!����w�9�G��g�X�[CM3D����Ⱦ2��QYt�A�fZ�C�D%��?Q��)�>�>�K ,Z�s�Z�:/��!��,�D1�ծ��1��x2�Ǉ (!򄝧y6P�#Q��*H�����l!��\��%�˖i-���rl�*om�'ў�>��1�Y�T�)�G�e|��%�)D�� @�Z��\���
wR1�U�)D��� j�׌Q	q�.?��䉲�;D����w��S��D�V*R��<����Ӽ>:UXq�-`�XX *�k���.n�����»b�B�)b,?�&����{b~��eI5)heB���&�O�Or�=�5���=3�Y1��� $������8�yb��-9dZY��GY�R	���4A��y��]���`VR!Na��c�g�5�y��.-�d QdD\�D�<1�,��y2��8k�4�I֫�1$`�J��yrC�(9p(!VG�+��d*��ى�y�FIr	�]AΒ�*<P��V�T�yb�9��Ap�Ȁ2�ԩ����y�j�1n�4��ǤL�E��(�G��y�EɜidTB6e��2�0�Hw���y2��+E
��1%�
2�ʌ��b���yҀ�hu�am�'Z�"$XV�C	�yb�
n9��dƏ-R	h�������>��Ol!$�>C�9s񈘶B�z���"O�����Crn\�P�T`�d��"O���W��%�p��b�*�{@"O���0�U!Qx��,͡(�����"O�Xp��E .hla��,e~}3@�'K����O���4����r��3�Ϗ9M�Dj%�f�C�	�/�z��j��∬�Bm҂�>C�1E�#%���u�vtH#�u�B�	6uo�T�� rV���C�.U�B�	�Kq 0��\>�����ؔ&��B�	�nE�cv	�&P�����]ÒB�ɹv�ڱl�Ez���T�\�P�O��O,�ۘπ ��ҁ֎?�����/��)8e"O�����L/���*Š]R�)�"OJ���g�=d���cPKF��7�'v�D�&܈g�L@Jv�քpc@�4D��%�� 3�ʨF�W"} :<�, D��bR��&��ˇ� A�Zl��j#D�p���3#�����T/1
�ĉ�`4���?����O���KbH�]<�c��õ�`��'i��0lQ����EOuJ���'x,y��   
��� o��4* �"�)����|6�l�քњo)"БA���yRV46;T9�c�s}��M��yB
m��{VoG�r��%ː� �yM�M<~�x�d�.u�z�+#i��yC�l �@�*i���X�9�?�	�'Έ�����~FМ�p�(�����'�tHQ�X�	�^X��o�%"�xI��'Zp�;�Kч#��A�⏳��ȫ
�'�I�� Pe^�/�DE@����yγ`��!�1DR*nnĴ@���y���/S�y)e�ȯk���Z�
��y��7��p����j/�`:�I�I�<I�) �O �
�ǌw�����M�p�<q� 	=�u;�a��5b�L�w�Vk�<AE��"F/�i'�ϒ^��Dʆ��O�<a���oN�|�쀩p�q��J�<��`̰4E����hĨ'Ҁ��'	F�<� �H�Y㠵�B釚<��|)��UV�<�0�j��������5�Pi����}�<��EM:�phb�K�*��9�6�}�<)� ��Z>�1(���6L$����M�<A�c���|͙B�@�`y�����RS�<!fS=-񰁠GcA�? 
(�!Ji�<��$�>kY�y��7���dIh�<)�%V&E��=HW@N�#�r�ZV��b�<�q�׼t9�\#]�g]�y�6c��Y���O�����BK�\у�Y�S�: `	�'����%L�}��@�"�
":����.Oh���u��4zs�Wb�}��"O0��G��6n@�٣ql�,�`l�t"Ot��V��?� E�a�۰}u��Q"Ot�q�o\�7=�ŋ��
�&�E�"O��a�5J����k�+aPu��0=q�(Rc�jHvj��J����̙V�<��A�3���	��M�D�vq{M�R�<�Ae�O�4�;�6l�B܋ �j�<�C�I�?�(ak�3".,��ƃh�<�-�7[fvU��MW3tL[gǓf�<1 � d���{sވ}��Q�Ia�<)�ǆ]f$IP�薇$�f5I��\d�<)P��=d�,����RL�dm��Wb�<ID�$K��$�����$���SX�<Q0-�
?Z2�#e���iÞ�p3D(D�ĹkB�4J:��T@��
���`�	,D��p�����I)3	|�1��(D�`˨=��${@��"(Zu��4D��*V���r�����-Q�@̀�M8D��3!����Z����#��Ro�<q���S	}�$�$��?��u����
��C�?=:6���)�"oa^�㪉9�C�	��~��g���0����#>XC�	�"��p�X.\�F���"C�Ƀ0�՚����p	�Ȍ �8C�ɉ#�L����L�h<�&ʔ`�hB�)� (�!Ї�7A^|�q��=
��-K0"Ox!�UL߬w8�c_�6�Z���"O�<��.��ެ+��LB�n��"OF�@�_1Mh�<�5�܃"O�`#��'j�1C��1{h�P�"O.�AU0M� i�e�^*x� �"O�4!HL�nn�M	#o�O��AB7�|��)�n��]+C#�i����*D�� �d>����%lĜD�ܝW�@d1��"D����&���"'��"T��!D�l�Q��?8)$�:�C%0A�I>D��#�ԽAb%#�$�")���0D���E�ˤug�)ӓE�3[}��6:D�Pi�H0@����hG�#���r&2D���bC9�b�"p�ĦL0���0D����2�U� � 8�<Y��F-D��i���;T�:�!m J�T:�c/D���.�&��Hs��@�V�ֽ��L/D��i��]�A�<-�V�L���r�G0D����J8j���#\�Iy�QH�l,D��%g� k��	�@&0(�v4)Vc?D��z�(L+K�С�f��J�8L33��<��hOq��hK%�H�)��pDN�*v~���'Tb�D"�~.2��bgծ7������^�ȼ�ȓ[�a���L�[P�ˈt[f��ȓ
_�<���'"F�5/2����	�8o/�)JPP��u\8U�ȓkrp�rDʅ��p�!⍨g�q��Oʂf"ހj��S`Q�����K���p2K�)T��f�[M���ȓ �ޝ��A�*�5�r��TANM��[��I�[&���*��^�R"<��_��:��Jc���j4�\6"'F<�ȓ)f)�c� 0����&]�n=�ȓs�ځ!Lݚ ��e�fʚD|����	O~(G_��ͳ�MU?SƱ-ߩ�y�/V����3tɁ:�"�"��yrjل�65��΁5G��-���y�ǙALV��a��(t����y�U0<W����(H�t �	��y¨	�(s���FOA#;�B�Ε�y2ʛ64�a��ͭf1 �! �y�n� �N�Cd0
DnP��b���'azr�0!�!1Fj� � �ń��y��܋4,�"Έ�a�|�P3�y·���¢;C���I��a[vD��'6����T�db豱��,Sm����'Hx٪�#�~�V�B�Qj�(��'?0��h��$��$!߀Pof�!�'ڊ��F�յ �ʁ�ǻm�h`"F"O|E��fM�,�ơpf�~�a�S�	F>�kr��6�z4�$�K2�`#D���s���4@�s�V�QT�xY�F,D��I`D�-�jt{Ы��E���)D�Ȓ�5�2X���3PUPp�0�&D�\��-�m�2]�TH���&Љ�F&D����O�vtΰ*�"�S}
0	1�7D�İv�$a�X�8�B�-M@�wA;D�|�!�R~4<*�/�%F��jt`7D�L�JؘUв ʇ����t;#f!D�x�צ�
 Y���f��4(��L!�>D���F�>j��]ҷ�P$}�-Hã&D��؄`H/X��$:B�ϡa*~	�a D�|S���"$��IC�BYc��=D�� ,����L6s)�x�g��!<��pIB���O����ݚoA ��P9lfn�C&oO�v�!�&X�"�3%���MJ�fm��n�!��I�<����a�/R5vYʴn�_!��7{nA9'�����ּxd���U���-Tx�*'Ï5{�l�zD7D���4(U2$$4�������� D��r�X�L��Q󠀋Y��X�' �� ړ��'��͚�ǖ0|(%��R2��I�'	��ZAk�?&� (±�޲'��(��'�pvJ��j���OH�q4�
�'�d��_R��(%.W����
�'4�  �V�@��e�N�)-<��	�'B��Q��5+7��¦��r�.�A	�'K\ �C�^�Vmi���>_j��x���'+&5���v�:�2",��)��'w�Љ'��Gl�m1u����桺�'r<�seOʱ�T�b�-
�,�h�'ňŘ�HH�u5De9�閎2%xe;�'�N�z���R��)�	&*0�\�	�'�X�{Ck�`$yYr�X)�0�z	�'�:�jcĘwY��x�"��t�����'�\�Kǎ+(���9m���j�'�$���Ҏ|\t,��*�T�D9�'2�@B`W�e�p��A���D��j�'������X ^��(4O���'j�DKv'�5u�V�E�HGOfd2�'�%pR��>���e���K�,��'9h�B+ܦ
U���#��]Ȥ���'�"���B�|=PSͭ4I@A��'�X\)b�+H�E��&]=+�|��'���sWKH-S�V�r:<�{
�'�ۢ%��x�24��X6c䵛	�'�P3"����r�cV�b?�
�'*.������#�ŷX~�Xi
�'Ξ�E[�sP՛ĠF"� |�	�'�`�AТܺL�����(G7���'G�h���ϧ�f�H�=Ǩ��'���eF1	�E�"��@<���'�Xaɡ��d�(�r��C�h`D��'5�1*��h�����[��j���d��$P5�@� ���aⓁ;_�B�vp�EH������	;b���鉒��)�4Cɼ��ѩ�<j�B�	�P�
} ��(y���EÆR-�B��()J4z��C-/���g��B�ɭrSF�z��;f�������rB�I�>�<<aˑ�8�Z���ۊUpNB����E��H� �2n[ d�B�I�+7�L!���-	|X�!��6=B�I5`S�(Z LʓeGP�ۗ,�)W�C� �񃖉�E%0��O�/(+C�ɶD���鐕��Q��OOR�B�	~�.e�� $�Q{��5�BC�	d���h�5��y*0'���C䉸�BM���Įi^��a��,C�	�#J�P�V-\작�gD�0��B�I8; ��5ɐM/J�ʦB8pÖB�IhM�R�@��pT[�#U�B����d����H�\�A�;nkrB�I*%ΔQ8�ĲY��r1.��Y�lB�Ikz���CY�tӚ�(�h�l��C䉚4�����bܬ�A]D4B�ɳqo쁩$��W�8��&�� �bB�)� z8`�%�>�ɠ���-����"O,Lb�홊-��l���[�y�1"O:��ÅY�0"1�.p���1"O>���٦6�^���� �{ӎ qP"O�H�s�G�^K��3n�lYQA"O�=(�`�"D�Pl c��,��"Oh���>L���7lO��ڌ9�"O����Z�$ɬ%�$�@�e�l��&"ON�zw ���\� �ַCo�x��"O*D���8gx^YiCn�"g;���q"Ou�����	-�( �ǿ7, `�"OJ��fb[�wlJ� ���y"�Z�"O黴��5�zdw`\�(�xq�"O�R��H�R��Lh�M�>J���v"O�P2cT��~���)�Pcґ��"O�}��HK
�ȉ���	22�M�"Oz1�a �,jؒ�TO��kD=q�"O�ɵ R�&�Z�K��T�\a���""O@�8�J��Vg���l�f�B<+"O��r���#Ӕh���"�哐"O:�
�\)V�R�Q">O��3�"O�#'I�}RD��Â�=jf�"OLtJu��z~  ��q�hcR"O4]{�HN05� x%���F�4��"O�C�@�I��Ȃa��@d`Jc"O��kU/*TƴH�ػאv"O��C�"�#J���ԻI�6t��"O����/���� r�ٲ����"O�q�&A{U���3��/4'2�[�"O�����K�%Z1�gO�z,�ĈG"O4����Al����E�-�����"Onds�oQ/n���Ía�05�e"O��p"A*��H����D�hA�g"O�xQL��c.�JcɅ�N��m��"O"勇L�.,ʪq�c�;V�����"O�8[��2Y�e�fSz"OD�2�K��boH0з��J��#�\�<نϑ�^�ꔙ&,�\�)zW��T�<$oG��<���K(4�腠@g�F�<	��B�K�yPG!�`�����X�<�JN�<�8� MB����H�S�<�CD�-3�!K�@ .S4\4� `ZD�<	5�E�M�PX��g�,0�xY�����<��ʟ73;xp �g��PO\ P� �b�<av�X�x�A5�<!�բSu�<�"[o�xȑ��9,ń���&�t�<ق�ޟE\�q	'c�8"��o�<�d��L�hDP偂�_'�x�7KYs�<�`cW��Fai���3d]r�@�u�<ّ��#q��y�@�0R �T��Qu�<) .������9�'p�<���� f�XhN�5�81cW�^C�<��(
��X9�$ٻE`@"P�	B�<���@�sD$�p�.71��e�[G�<�0��5/_⽁��ӟx\��A�<I��-xr�Ke�\w���`Ӈ@{�<
EG�����A�T �a�B>D�@i�H�&�9l�/�ՙ�@(D�$J�O�hS�����6d���6l1D��	�U�,��mH5 #.��d��+D��ԍU'
j ����¤_f��m.D�Tp�)32�~�H�\@R�5G.D�"�%�Z�M
V��[t���Ff0D��aŎ�+8"q���(/<*+D�� �ّ!ګ�>M��j�>t�H��"Oġ��#?ErA3iui>%��"O ���ͤL����l	dh&"O��ѠR�K1���R&��0	lؓ"O�	��iN6l[�aZ�n�M���R"Oh(+�b9)6
�Y2d�k�6t�"O3Ǒ	�x�y�?e?��HR"Oȴ�����ba���3��(��"O��(1f@��YE�ǈn�b})C"Oڡ�U�Q%O3!��+O09�j���"O�&�<�q0`!���a��"O@�(�zٸ�jA��|�T���"O�=�e$=+��HKQO�8Y�ba��"OrA�Te�g"y�d�km�7"O �:Ç˒敲��
�%��٥"O&`��YC�\��U%Ú4��lxQ"O
��uoŞc�P�R�2^	��D�<��MF:B���MmJ���B�<	�ۚK AA2��6��Day�<97o�9�p$b�/��lB3��`�<�vQ��.�c���=����v �b�<9!�A	FLpiߚx���1�"�w�<��Гx��rB˅w��10��p�<�d��fJ0ls2Ǎ�%�Z�	�kNj�<�1L�-J�xʆ�T0?@t�
&��k�<�UCY��o�bQ�S�\N�<q�ǂN��O�.}�P��NI�<��B��@�D(ګ(��T�b��}�<f�W�5OB�k#AE.q8rp�h�d�<I�o�k�f�ga@)����EX�<�vi�.���F"F<�c�	[�<���;����v`]�:# �W�{�<!6JL5�T�R&@+s8cP Lm�<�r�۷��oC���B�k�<�b�>B��v&��^� �25(@S�<��-�r�p�Bi�F��u����T�<i`�yYN�k��O�ԈIt�{�<A`F�8KpD���]0u�kPb�<����J$�8����5��)q��a�<���8��1XpL�:��9Ї��t�<�V��������,�*5��kW��k�<q ��A�Hc�߃Ίu�a�c�<�vă�"{	��)��T2Z=��Nc�<��D��`_�� &I>^�j�z�.Y]�<a��U�k���L�[�䘂COc�<�J�i�nqpC���Ez�,�R��\�<�A�[�6&�Y}�Tb�@ Z�<a�U&}:�i����cX�p�`��`�<Q�E-)�Ē�)��N=����&�u�<�5�1����q-��y�B4��L�<�N�7��Dc��*	�:�X��L�<Iť���P�`C%8dP��B�I�<qSB��������P�2��J��M�<&�"	HP�[�,̨T�l����c�<ɲĜ��n`ʗg�h�b�RM�u�<!2��l���q`���Z4AÖr�<AbCS�]��}j��ec�� ��FJ�<���ь��i3@�7'Tfh���j�<ъA�惡�D)�ޞH�"I�i�<ɷ&�<]�
��� �p,��7NPz�<) ��,a�ZT@!(��EF����Uu�<9�"�UmT�w�b�>t�SHo�<��CЌ(+�XB(���4��1,Gk�<y1��N�:dR1�W2w3pY�7,�e�<� $l�We�b�uIRaS"�0\�"O���5�Q��-b��wL��f"OF�"���/�a�E*�4��"O�LY���2 <h�	�M�o)�(�a"O��B1�ހF�58C/*(�q�"OjHA��E�ĩ�s��*��!��"O.�7�K�m"aj��$����1"O��ů]2(yt �[�[���9B"O�`rO��|�������'p����'�~A�''���	�=X|)
�nGp�c�'ج���e��<�=�f×7A��������XE��g=]�~|�f�K_�tArE۲�y��*A�$;"��h�%#rW��M�$h$�S��MkȂ�\����1�8ѸǦHa�<ɧ)đO���M�4QO}�O�<A�'��|2n�'-L8�RAЗo�d����%�y���� ͂v�L�e��P�w�yU�j$�C"�9cŀ���lȕ��O�#"�j؏�@lC��Q�n}�#�H�<�aF�V����0懖-��(X�N�F�<)An^>5q!f]�!6����Y�<��̒.��bo&�1A�d�X�<y�M9s�L����i|-!���T�<Y-�
). �Y�PRB�A�N�<q�Å�~����d�;	�E�F�G�<�ɟ����tb��v��m��&D�<�Ѭ�%.vmce�<W��!
�|�<! mõP�,��$AՊiAz��3�y�<�DF�<i����B��}��!V�[I�<q�!m���b܅����j�\�<��j����Yc��}KZ$�Ć�A�<ae�ِ"�.��%�< �����hy��)ʧ02�d�'S�4,���nD��^Έ���&������E̅�_�p\J����'l���P�+���^�:�(��f�qrh��T|,�ȓ�����͍ZP̄!R��8d����;n%��
.pEYCbҍ��Ʉ�/Mh�r$�@Bu��}�~E�<���	*u&���I��.��m��P�|!�DO�Ɉ����=Q�PX��`Z��Py2��7>��]���;B0����N��y�A�]�*H3!�4�,�JVώ
�yJ8����ȝ�1��J��Q��y�Ɖ{M��9���uHr� �#Y��y�%�?h
`�#�fzX���I\�<�Th��,��C��,
���WLo�<ѤN�h���餂��}����h��p=ɢ�V�+�<d�&lH�f�媤��d�<цe�u���!�KѵKZ���Ui�<ARg�	o� ��O�N�8Ȓ����<�W[�'�><�P �+f@N�:R�Za�<����;+pIbaE�(O<�E�J�a��$�S��I�����R���z�#�?�Ȝ��)�� 4��&G���vJ����ȓu���R��!X^���,W�7x$5��N��E*��j"Fl��
3L���g��@�6����I�@�N@,qņȓ3-�+����
0�T&�~�Fz�`U�O>a�t%��G���UC-�@���,�S���.0��aG�W��i�&)���2�S�Os�q��cU�/�(�xp.�J�9���'O�̣�
��� -:�%��5�����]���'\ �a�(�$�������N����d>��~
� �d)#��ov2AJ  ��+g�#�"O��c7-U�
�0 Qʖ�Y},��Y���	Ң5K��i�T� ���a�1O�=%>E����f!fk7��6�t�u͌��yrA��0(��ڒ��9�\XQ�Dʶ�On"<qK<	S�,%�N]; !�IJS$e�<� ��?i`=�'А+�f��&a�'-ay���ڸ�rK�=Avhڔ`�o��B�ɵD5�Q��"2%�n���W1Z�2b����͸'p�'��e�T.&A��$�ΐ\�𙣍�d�s�O���%),��UxfISd�H!2*MYH<��'ǞE�(�d�Qaǰ���-�cy�Q�h�<���"��?@�8��͖<��Az�`ò(��B�ɃkΙ�PB[6f�e�a�%]s�O�eӊ���Ă?0vXC�b�I�L��LG��x"�� 0�J�"�K��@獉�OЁ���6,ON���Ɋ/Ȱ�HgK��*�*E�W�'�r����
i`��y3 �bv��1�Z����=�ÓeF�*I�t
��h��/>�D�=Yڴ^>b����|b�>����/��JZ�R��Vi�<��
Y���c�k^NLP��"t��#=I���R��hЇ�f��ـkQ�	��">��Ox���tƮ��	­�".���7����y"�(ur\�+�ߒ-a��RenN��y�P�0�I>E�TB�nG�h�6.�6$T�cl�nb�=�
ÓL�)��j�ee$듥S *��T��t�'�DU�%jȒ[H�	
g�+�P�<I��� �nY�k�-qjJ-�@�M�<���;z�A�w �'$��X:�d�<I�F�q���`�m��[��a T Fk�<��@�[s�z���u�l�A,g�D&�S��C&��P#�]�Z��j̠i�0����R	##�?��$[��߆�%�\9g\�8E|��''4щ�I��
3M�Ch<���u�;$��&�V F��!T$�c�<l
��1D��b�#��z�������#|O87�2}"K3Bq�!J�z�j�JӼ�y��K�yu��)��
�HA�-K�'��y��ߗb]*y��S�@<2򓦟����p>)�CS�?+�x"�$M{\}QE�u�'�axB�ݣ���[�ȊD6�ءʒ��yRj�%n2�YūBQ�Uc!/�y�KQ�{B�\{��^(D8���@c���y2�?L�bd�H���l!� ���y«f�3!Ӆk�X!!C;J�<��v{ ��w%�U�ft"�J,<� �ȓG.@P�G f0����S �!�ȓ\�0��"M�4�(�2'S���ȓmO``�n]�a���A�l�΅�=��'��xB�� �F�(3�A�<�8$A�?�޴�M�ų=_�TC�b]n{�y� r�<�E%E�/Gt�a�@�K�>�bu�Jj�'^Q?��W�V�Ȣl�t�ػ\�R�w��OxB�Is�Ț�C��:d@)�vFߙ=����;�	 '�n!R���	(��B�ޫFӜC�	�`!���V灆m��h@J��A��6,�S��M��"ߤL��a���֛ei�x�R�<!&� �z��!��)��&n�G�<)�.�H3��1�j��Vp�p���l�<	1��X{n%x�oN�,B�	X�c�榉��\���〢_�h����YA!�5�+�Iq}S�@�}�GE��'��I���0O��L���RQ�<i�����T����r��KF��XuQ�b?�0 g_.E�8e�ą�Hrh �n!D�� ����`տ�@0HV�:s8�!�"O�,�d��F6�4�����;�Є"O~�2&%ɧ0,�"�I�ܑ��O����=��-�Q|�X�̜�G�\�Kt#�JX�Da�Z�����O�9�Z�Mxv*\�@��U0ŤD�C'!��~۬�э��pu�2�eNN
�O�p�����ۯ8�A`鋯@c0���(�y"ƚYƌ�)�I�;�n�	5IZ��y�E1U����� ($<ƄY�致�y��A�{SH<8SI��K0���Ѕ��'�a{BH[�7EZ�R� S5��bs`���y �
�,��lT>|6�j�.2�y�S<�I�m� ��QB5���y�)��H@�r�ک
��e�v	�&uˮ!�ȓv1*1�����zz���� t��ȓW�@���2nD@�#X�x��B[ܻr ;Cb4��ˍ</ά��ȓ��AѢ��.�vdy�.Ӱr�Ɇ�))r��.�
�$Ѣa�5D����ȓ)�pQ�⋾��@�#�-i���ȓ��H�+R$L\�9��)�a�)�ȓ6��6 �){=��A�$N���ȓ�p���:Lj-i���,N<�X�ȓ$>T�����˾����89��q� `�u-
� �z(	"`��U�l���g�r�r�j��lO����J�9j����s�>% �f��R�Ő�)�x7fa��tr��Am	>8
�H3aS�0

�ȓz�$u�3�^y��-H��t�xY��`f��"%�dpD��G,cڌ|�ȓ)�"T���B�q���`��v�����h{�\h� R3pM��
$�(���ȓ	B�0G��2Z�*���Лk.�ȓm�y�́=|'�8K KM˚a��.�����V8-��}� )�8g�(8�ȓnĶ�	��Z�)8�!תߘZ����-e�M�fO�(n��)��Sq&�B�
6�:����X�4��d�gA�s��B�&-�����į:a@�r�c� H$�B�	�?��i�6��>�<��B77��B�ɳ>4�X'��S0�갊�>��B��c���QB���D�������� �L��z�
вg�-}+�I�ȓ����%ʃ9i7���SM�'`�<��]�U��]�ߤ��®��SB��ȓ2M����=t�������5��9��6��`ƞ%LŊ�YACʋ��}�<!����A�aX�i�e��L�X̓m:��qu��rg(��!��!0�h��n���h�S(db���ˋ>{B���ȓ���1��C��UXW��"��E��!�H��ED c~��H�N�;&m�x��xz�d狶e� ('eГ/�ȓc�R�(�e
��}�4��q�j�ȓ9iBd1�+���B���ېsq~a�ȓ�$�J�Q��r�g�]�RهȓR����ٛɰ�E&	�~-,ه�( �s����TY�ӇȗL^���P: D2�)B��<1�1�R7ee�C�	���SPiק�9��E�#+�B��H����S�%[$�	rF!y�C�I'AkP�{��3&B4"�i͑@גC�	� �#��:|(�$O;�DC䉦_ϰ�De�Or��J�NJ��BB�ɯ=/ꕨG��ؐ��e+L*T�6B�)� ,T�b��K�����Q?	\@��"O � �ˮi���z$G+W
���"O�D�HĽG!�H���0;�Ȉ��"O��b���D���AQd��}-�̛ "O �z�⃴�(�����ZE�a�'.:@��͒=>a|�8{�����;?�v0����=y�G��D��B��O�p�Ĉ(1\f�#�'M�A�E!`"O�|h^�R�X���!	x�A�����ĘâB�#}Zv�E-A���R��L���#�%T�<�Ai��Y"��Ħ��Mz����-ߓ���ʅ�J!Hn�	�~IQ>˓�hÑ�O�T�΁I�H�5X�dq�ȓ (i����<8�x��P�Y��$�0�@�0���C#N�c�a{B,L<�����ȟ/@R`��,D�p=!����xkq�H��Mc2F�[B�0xq)�5���RD��M�<��[d�t%�W;$�§�Qܓ	M�dIN�v����޼Q���2�A��j8DHZ�70-!�d)Q	����gſ.��㥫�+�F�B5�ˉo}^��'�<�F�,O|���=fr�kb�Y.u�}�!"OJ��SKF*pp)*s���{�Lխ�-<�h��r�W�1��]�퉂/�j�k�?O��}Y���P���ҵ-n8�� ���?I�,B�u�L�h1�1ql�V��\�<1Ќ��=�"��7����`[P��#|dB���������AFX
�V���3 2�)��"O�u��2/��92a��E(J�@�"OT9��ĂnfHy���܄p}#�"O��"F܉� t�DH�{�(�w"O���'g����Cd�S%=�N���"O<�AD�2U�x�b�S�!x4ـp"O�5
"�����K�C�	iX�"�"O�ڧE� kP��¦�>YSR��"O�Da�-豠҉���>��""O����㞓Y�6�ɆȜ�us`��"O�����W�Z�|���ݶW~�ط"OfĹ����wV�@����[�"D��"O,,�VII?'b��WkF%ri� p'"Of��p�X)w�\4!�	i�X$�E"O����L�:`/c��&���1�"D�� b%A�C����p���(���G$D�<H��Z!��t��
.&�x ,%D��r� �k�t�8�C�?=�A7�?D��c���82�5�K�'p�l���/D�PA�a1K`�$�@A�(X]thi�H*D���=YF����2��q�k7O�`u'S�ؘ'bi�ⳤ�9��ѭ34���"��o�<� �5s�4Yx� ��ּ���hyr��	�$�B�N�O���+n�:U�s�p�вiأ��C�bs�p:��@�����C<�$0&�� �%N�� ��ǐ~�?��Q�ggr���I�]�N �b�Nz��p�FG�-D����� �#��0�V�	< 2N�P��:X]� �KLcx��i���}nH< ,��Ag>�:�H[�#�3,E����@���w����M���!b��:�!�$L�+<<�S`R�1ZMZ��!(?��3? *(��Ԧ*R��cb�O�������Q�F �B��6"OBUK����*�^mH�� �q�,eA���4&�|��b��V	 �Qw�Ӕ3�s�  ]5OQF��r:����<:h: ��AձHX>��ɪb��d0�n>2FdP�D�!��@� �dX�$��IL� 8r�Kԟ� �GHxh�Ԕ>%>U�`cM�2?(`!�6.�"mQ�B0���|�1�(�H�(u��$r�O�q��h5H��X�����p�2�ц+�XIk�Ļ<!��+�gyrgʞh�@qȆ�>ܤ�%�M�#[����GڗG����Td�h�k�B�~��Y5X`4��ꎱPK,ܩ�Y�P�DH�e��x؞�{"l	r��� eGKcS@���Eع#�l�8GPq�\h�ŕ�]Q���ME�J�`SD�����&�f��-��6�N�*u�t�4��m4�O�eRc�۪t��1�$$/�(� ��%Y�����"_Mjl�2m��5@�%YL����')�"���-�|H꬟,8���Ѫa���&'Ҭ���ɶ>@CcM���p���O�m�l�۴ie� J(�A���W0Ա�%�ǂM��$ �d4�*�C�:X �dA�&!���~�'��iP���5���P�I���iܴ�r����,�i��8�0����Ǳ/�!zp��\cXNTzV�L��Db�,3�P�j��D�d��L�0�@'P���"ӓ,��H��F�{�z�R���/p�1���
Hb$�wN֫2����AY��;]���KL˅^hV���bU�v.`磜��� �k۰��}+��Z����H UR@"��.�:��W**Hے4Uń!p��Y�2�������mH VYX*�]��K��U���4䖯sE
�n�
Lr5�e»ڈO���5n��L���	B�d?�DP'+ɮX��h�w��1_��:էϊN+2���Ϸz�NYHS���Q�ɖ>��U���Ht�
R��8@���?�)�!�&���O�8i�a���BhI�S��2H�|���9Aܬ�*F�����s��JM?�F�װQ �@���<LONͳ!	�*�%���
���B`�T��������*Uj���/%�'D_��:��]	@��;I��i�%�ˠe����)�*<�>�p	����e��Hĕv֎� �g]o��� �)�-�BPyG��OԽ�]�C�����h�U�L<�O�b�#c$�7Zj�LSƯ�Dx,@��j��#m�>1��ua怊��W'&Kba���֢G}�$��(�PxB�Ӝ\,v㭍3�dtB����Op��7��O�2��åF�p,���T��.R�,��'O
�q��'d~�jd�� 	.@2�'K��D-e��1�P�1 �(J
�'�Dd�a�_3�<�B �=p%���'K��B��=���`�@�^�H+�'w�$���.A�a��S��=:�'�����L�9�D��B�C���	�'�h�ek^,�p�"ȵE02�a�'�q� �R�,n݀���$��j�'��\�'n�-�`��aG� d��2�'��b��4���0��"sh��
�'[<� r��I�tU���w|�S��"�H������S�ODF-���z貇)�+ΘzA"O؍{s�VN�Pر.F,���R�t�w4P�p�'�h� �$�%�HrqU	�ze#�TS.���m@�:�VaB7 �0r�L00�B�)bL�9k"|��'����w.W6LX��g�YN����.����nV4O\��@����	�$]6A�b�K'���F�؁w�%��-Ď��=E���J�Im���c'�������)�����fH8z�����0Ĺ��*��4Qr-	w$����Y�St�u��F�>)A�>�ʔ�דe/^�Z�Q�F LhH�`δpE��v"��4��9� ��P;פ�y�'�D�D�f*Z�˟/x��y��H51c �bS��w8���0�L!������Z�X@�G-��T.�q��*�>'�-{@��}Ѷ����-X(8��N��'	�t!���3�^� �):Y@�Dy����`	�ɍ0�F,��/](��iG�n� ��b�:Z$���$��N�v��fM�6 b��U�>E���9ê#T��(n~�y/���@�a׆	��Զ<ƶ�po���E���{B��Q�� X�D(�3A٭l��I��3
��
�j��D5v��S�m��$�1i�4�`#��%�.4�ˀ#����^?�	,�v@���8l�Йf�K?y	N��s'�W� ��j�mx���*
�h���;Q�úy��%��+OL���Ȋ=�2��7�ݲ�~�/�	FW�H&��Z��'���1;, N�1!! ����c +L�����I��K@kU?	Q�c1��!��&B��1��*I�Q��	FcZc�q
�	9}̆�7��9�}��0*T8�91�X7�$[�G#`:�c� K��#a;�I�K�t��&X�> �Snx�7��Ј2�Ɏ8�� ,��P���p=��!��9�@LA�gS�9�:s��z��'cy$�����O����Ǧ��/عF��̻eb,
EѰ�8D�h0�C�Z�#��_ ;ƨUh"��@;��'t�M���h�g��w"~ٓUmA�w)�a�E���XeJC�	��bHs��p��kԭ�>%B�J�j�77{n"��'ڼq 5'C��Ր�
��^v�١Ǔ  :��(W~�Q�Pq�3!���h
��Q+w`✅ȓ9��(9ĭ�f��Q��Km̧OΘ���$���%��=aB�,�1�pR���p	�7����C�I=ap`���n�u�.IAD�k4~��'��r�N�E��јC7�Sy�D�BBE��IU�X���'���040��.P$��uG��,cC�/�?Ib�߶sS�iQ .Of�i�gX):�XGΔ�#���*�'�\����4u�抛8|��+�E� ��3 ѧm�������SZa{
� ���E��'3P��0�U%�5�c�I?\3>MR�AT�qعq�<����ECʲI��(C�&։P��tb%V{!�d��C�R�Q��%akj�aږ^P����05;��$
Ѽ��-�`�� Ј�	��\��p����	��Y�:R!���Y�ĔI?7�<��7�+7P�Y�E͛!z��{��8x���2c�~�3�	�$K�yf�'�<8��շ[����V:/ڊ&iԪRdJ�W�,,��14Ms�^�FvI���0=��.5�����L�oaƠ��hI�'�����	�/0����0΍mfҐ�q��,� �D$ۤe��)E�-��pV*�R�<�`o�1H(�k�i��E^���	��M"�;F錿CR�0������(�$�~����%�<��Pp@�=H���c�O�<�c�%=n�H{�ڗ}�A �&J<>�h}���7@ �m�w��ub���S%<k�TCd ZV��8�2�kՑq'� �H��rK�х{�$�{d��6�:5�^��XLp�OSYsFgK6P��zPL����d��u��|(��S�a�F� �D�<^s���el?��2��ݛ� �&��Q�	y��0�k��tub�#�	x�h���c@�q����3$�y�<�s�ҽ^I`P�����|�,��϶>�8�UDǄZK�`�g��\��l�S�R�_Hq���]�B�F� �蔍I�T!S'�K޼C�	"T!��a��U�.��VMB��f��\�uuFqqR��=�-�-g��<�N_?
Ot`�n�|�����$�S�ի!�i�����O<;UX��fS�jT��'��d�TE��5XȈP�],ytL��2��;Z������X�O��Ȳ���4IB9��jq�b-��'�n �BOʬd�~�R%Y=h�U�1��-��Z��|��9O.�Z2`�p�vIR�X�x�b�j "O�QS��
.62t����j��OTx�����0>S���0��&�G{��ib�l�{�<�W(�k- �b&�
1B�I���h�<�m��&��a�3���hՎ�a�<���Q/��&�U8tp�`�M_�<1R:�Q���9Og��`SlUw�<�Q�ϑZP̌��@C�v���&$�e�<�Í�V�xp�+M.G'��ې�a�<q��Խ?w���Si�N�|�4��z�<��-'�a��K�������X�<�0���Z:��h�!��pa��P�B�<aE��/`�8��^K�ŀ�(�}�<�c��o�Mْ��h�ҵ��n��<9�e�Zw}
dHCU�TM�G�w�<�V�ޡ ��Yt�]�؉֡�m�<Y@D-L�����k<*���Nd�<ib(ư���gO]�" ��D��K�<�ȺzU� ��&њ=��� �F�<i��	l�1 �.�\liG�<S&�"v<�#0)\�r�SP��D�<�f	ڊ)����#I�)�N�K��C�<9$$Ǥ9�J�)�,�9�͐t��~�<1M�&+�<"d@F�Y�aʖ�t�<i��E�kY��
� �6��l�G�l�<ٔ�S.R���rd��U���9���R�<9Ǎ6N�!#f�5G�D�y��K�<���ڟ֤�"�,H��<��N�B�<!�!ѪgRB�@F�mH!4er�<AW'W�n�N]kDT�Oaz����No�<�S�A�x�e2k�>/F0�!��Q�<����1�F=��ԇ����s�LJ�<��� �v�"��gJ�$Y��X�!ˀO�<Wo1?��|�e�!t�&!�T�H�<�V��M%��h"GLE(LA���E�<!���1ך=b�΋#�B�M K�<	�[�����sd[z�4�	Ly�<�&Ň�0c�
OC�db�<D�Y��܅�E�$�^�Wr�Bs'/D���Q�J*�Tk�,�.?0r�s?D�� :���oO:p��@����q3�"O0�k�K�6�H�����ro���"OH��T�
�_x�ʆ���"_�U�"O���Õ>���3c�F�^�����"Ol�"�M��RK��9�Zhsb"O
�a�)�#�d��,CЄ՛v"O�ɻ�F�8%�+�v�Pї"O�)�"�7|�I��	�b�<�Hq"O�!�0"�=O�h0����!5zt���'"����̆3)�a|҄Ğ9]�3Ҧ́�D�1��
�Ӱ=1�Aѩ4c�L�Q��O��(�Й|[`��� � R��Ia"O���G@�7q��aّ��Wc�ЙV�dL+3D�P�3� ȼ#}���ƬL�I��
�f.���F�<Qb"�tZ����XS��a��!,�)H�T3L�	-9Q>�&����/��!*��� ��㘝��M\>pIv"D���(�B79��EÖa+Z$� HH3	#a{B��O/|���-8j�������p=�Tn�m$�EX"AC8�M������a 0}��J�	�_�<9�퓐gq����3q2��v��mܓ9@y[�a�h��(���	\�0|8I �B�y�F,蔩�1�!���	'�L��韀xZN4�(ߒu�4���M�|���'IV�E�,O6��&��6����_.���"Oxi�J*:��\�&o�w�z�W�w�X��#�m�b��ɰ!����ɤYF����nh�����b�(�	��M9�?!��ѧT!-��T2uM���- H�<Aō^G��aЉV�}�AŊ@�"�\y�ʛ=����/E�ⵐ$,g�I�B[��yR�˃l�F�#@�e�"�Q�P��y���+������+[�^��4����y�Bx�n�! O��L��aWA���yba:L �P2퉮N���Y��y�ײ*�b��@�G��(�5��7�y�+�;\��,�&�J�0Xx��#:�y��B
f�I�f�?����EF���y⊈8]ؘ���	1U� :�A��ybj�cˆ;q�A�!��E���[=�y�[wȽ�\"�8��G��(�y���8PJ]���BV�[KN��yB�(d��)����!�"e��a���ybHO��%8zj��@A`ID��'�1cTc�3� s� �i�U:�'�t�P��R>`8Y5��(m^f��'�@�0Ȇ{�¼��B	�K�T�s�'����0f�!y:�Y�Ԏ G^���'04uHs�<��\�D�I*sur�'D�s��ׂ��axD�Z�#�z	��'�XXrF,7P�,���~�1���4��r�n %�I,3�����-D�ܪgbD��ek��@�+D��AwhӰ��)KG�x��i��'D� ��$+g����W+�>��*��8D� ˱�M-T����Y@y)�C#D��[`ԥh�xy���cJB�P� ?D���GĎA��Ңϓt� �<D��0���>4��1�˝N�
ij��=D�(��L�`-�VV�07������y�GT;/��V��/��5�0�7�y�N@�Kf��'�jҬ9��l�*��=���Z��z�'�ҭ!��|���+vK�\L�y��'����a��4(�E�D"NYZ�}��ST�&a�3g�}�O��@��CA�S'�; ��-s.:���'J�y�DG�$4L��bh|XRZ&/Gz�aRa�<�A�)�gy"��u�j�X�qqIW6�� 3H����l�mqO�$�q�AZ�%B�x�%�3l��AN��m�dX�#^Z4��)� �z��E�`�v�+�EA�� �-?�d��� Ý~j�K�Y=�1Q�f[?B���`�� =��ţ�L�q�iÖ�?�O��H�
 F+����$Q�P>b��J�&e��=Y��~cߖS�&��ȡ��Tr��O���i�~"ө�%u�I����N��Y#Ь]A�'��9��I۞&L2Y�v�`�4I�9P1H���~Mr����9������Pq���O��Q�̔\�gy��u*L�	 D8��˴�U���$�#
�(�ϓ�?	�d�	Th\*" 1�7P�tq��đ6��c���ZCqe��~jZ4	��Q�3���ëQ�,q�k�8n\Xp�T?^i2��I���#`f� �^ų�~� Mb��K�T��y��!	�KFd��Jι"d�{
+�O�l�D����b��ܸ�$��z���!�?) .9M�2���J��9JVE�>q�I��ZP��ڦ�Nx��g#0JʼY�b,&�џ��a��|��0	��'����v	�#/.�`6�Ĳ�zp�#��${��Rb^{�+�gy"�	
I;��$D/3-��ZRۮp��!����|��	!m��9:���q��k�
o��$�Ƌ�b̧�����
 |�x0#�Ād�����gG\ٓ&�#'����w�2lb����ԭa�+J���I&|��1o�6�����i]�4�����
;w،�+�01(4��%�:F^JT�c
Oʝyq�C������(R�bP����}E:�q�'�@��gcJ�z���X@qO���<���3톋HJ%�!��6~H���$�6B|N5z���NE�� �b�/0���!��U?.B�I�Jg4y �DMDF݊�e	hl�?�t���6c?Mw-�p�V�k�bT;y.>�P#)D��z�,+<��r�F� ��4:�a'D�t:fh�|��>&~�� ��f[B�I�g2��HS��$KQ��r$�C�	3 e�-�%��ly�$5�A�Vm�C��y���ѳ�	*H`��_$NZ�C�ɢr�� £�;M�Bes�ޮ*�C�ɻ���!�$t��ɂdqBC�[�nY�$bDF���H;fXC䉗sA�$1  A�e��E�g��#�ZC�	/U,3�"� f��ys� ؤ�|B�	!��x�+�4'��#�&�9C&��	71�VEQ�-���q }AQÛ$"�,���M{jф�3�Ȱ�4�(S< 2r.�
s�F��'qBq����q�R����!L����T#V�)�w���s�
��^	x��� 蓠vM��%&��g��� 	3@r�A��J�X`�m��	(&�|KP� $z[�X���3( ޣ<�B"*#�T�M %x^�L8��0da�>���q�5W���d��t�S�(�qO?qj1G^�g5���$�g!�yd�ݴq�*��+lMf�Qv�_CP�Ec���'�R����+@���`
+vZ��O.P�Pb�<Q"��d�B[���#�R�*���1L���%^[9��R�O�
\r0��ܟ��
Y~,����CZ�8�7E�|4��ׯ����'�|���E/)��Q	V��H�*h��f߈�]��.c���dK����_�
d+C	�����|��`׬G,��A��{T�P�@�W�'fa�f V�B&��)�,޽}^�D�(��T��IVMt�А��M�W䑓%�n�pu���͌+��S��?��QU@֌igL�dM)�ad�^��`u�wʰsvd�L(E����'nL�r�/r�������o�d<�'4r���%L7!�vu��	2lpl�;R���5WV�W�9f��fGƽ#4�r#�E {CЀ+��~���i�)¾աqbL-a;��{�kO:9QH%�_���>�߅%%��6e�0[���Bc�
��K�*R�H2åۼ,U���^�^\��$*��m�O.��b��$3���N�ab�qf�<>���
ϓa`�Y6m��~�T4d���pn	�O<�sU��\��r&�G��D��{�d����%)����$�(�WH^DK`��dO:9�<A@�ReM8�C�ސ(��Y  �Z�k���ƎRgv��5&Z#���'w@���0��z��ΣYR(H�ԈW�PT:
@"��)�T�ȴ`�F����C"�M��B�&A�գb�H�x;�QA
�Z�<9���7�f�DO�4����a���&ߢU�O���C�$����s2�(���(�E3&� T�֡��
�Fqm�X�>���e�N(�<P����h��#�O�)�-�5t���m�h�-x�xB��:��U[��Z~Ɖ(Z���C
aZD�8B��*�y��0y½�r��	PQ�9N�7����02�ܣn�fϸ6VJ��~�%هb氺ֈȤC����l�l�<i��*��(ɴ�I���c�t�,�$�N��P�a�/J8L%�~RN�� D�+�uHA���K_�8��O�A��|�*�YP�`�Xx�,��f<9��g*�9fOE� ��dN�#f(ݫCoЂ!�@u��J�|��~��ߩ=뚰1soۮs�����	��Fz�ňu��27��:WkM���{��'l��"�e�"$�X-��A�@����Ċ�W�""n����yѡ(]h��"���4rb\Y�P�G�vT�8 hC!�y"@X/ni5�X�2s��E�� �~R�C�D�D����,Kb
�)�gɭ�0�F� �p��|R1lF�Gi6�Ԭ��y�O҇~���0�A�83@E�! ��&�(]���6�ӁU���ZJ?�3�G"4��y��P�S��+�,�~���
�Ȁkg.	y*�mY�S>?��AA�S�p����ܕS�&�Ӏ��]����4n�;(`}�  A�&v�@q�% ʓGZ��d�N9'xA��%|�|t��*J��$3��*Z�6�x�G۠��'�%D�XY%�U��<�ӎ6eoL�[RIǕT���x%�N9�PP3V&�>&�lh9���V��b>��%PP$qa@�U�`��QJ����C�4�`����}�V�C�:`3dIp�4G�����:A�<�S�����h#�OO(~�Zc���3Jũ����p�9kM(P9p#8|O^��Vă�?���C�E�^D�4襀�W��TO�4N)�%D�\$I��Q�I�v��e�
��a��Eڹ����S��O`XҪ8+���cD� ��cS��$��ò�
m��j ˆ0xzs��
*V
C�I�
�
��`j���Տ�5�$���.љ��P�IA�[�j�Y�HҊ����9�)r'߹^dz�Y�mV�w��"OR���&@�i�5���u�ڼ�Q�'k(�Q�Z��0����>G �)h1�ٳK5�1"�U�H��d2#�ؙI�?�M��+(k&����� pz<�f�}�<���O�P"����B]аysD�M��6m�ЁA2�F"}����500��P@�.X�����@�<qw���}������5�����iłw����lO���S��y2)^/���QH	%U��x
r��y"AI�i;X(�%���1�e�)�~��/pԄ�Ɂo�u��7pNDha��F�h�VC�In�dx��@N� t����8-\C�&o"�mZ�HŞo�z!gI���C�I�)�&�	�aW�LbݹQ@ލ5��C�I8 �0<�0���MSH�3#�_N��B�ɕP`��㔅\0�(1zf�е;y.B䉼]�����'сF�
ɳf��(��B䉃L@l:t���Xy����e�;F�B�ɻ1<4�l�)�ژ��D��X��B�ɌvW�l�7ȂXa;�ڕ[��B�I�F�>h�c��|�
���J�?>B�I�o�S�D�/��\��N�6�TC�ɧP�l����m)�T�d/�,�B�6;��	�ܷS�И$��+TЪB�ɬ_�ȹA��,�Ь1%�͏6�nB�I���
S0����B\' �$B�I;f��y�g� y*q���d� B�I=fR:�@`�gk¡�PW�G�:B�0@ƈ�`B��)��a�.(3,C�I i+LФ�Ėp��Y�4NT9H C�I�sn��.��r��'	��l��C� �du����n'�xa�[��C�	2���)rc��dN�4��nJ	��C�	�.06�T�B�pH��s"�)a�C�%Vd�򤀖�!f�`�.d�c��FH%)k�eZ��G�HvU��7�	d�(QU	_�I�Xm-ġG�VB�4�ʩs3�P#dVTɊ��A24�*B�	�9j�бg�ÜY��F��X�@B�Ɂo����B�4��G�%4��B��-�hX%�����4/�;h��B�I�'&���f�R/�l㷯�)��B�	DS�,7o�)~P�p���@;�C�I�?p8�a%� �ʈ�(�7*�@����Rຫ�A?q:u��J�1~�!)��ɽ<�~`Ju�G~Bd{xn�Ȅ��]>� 8���N� ��s��8Ԍ�$9O�X@�816��#a�<E���K:�}"�e
�\=
��Ņ7��`�#!��2^����Z���	�&yR$��	�3hbaIu�8X^�l�7e�m���q���g�T>��b�
�@�(@Kp�i@�O.��'q�mH�o<�s��s��	e`Nm��X�� [5U��yp�"O0�k��IN�E�3/*���'"On`�C�۴h����ós>��Zc"On�r�-���h�����Q"8E�S"OB�`�۰D[�P ��(vz�5��"O�8i��+�ƨ�V���)h��"Otu��GY�B�����a�n�*Ӥ"O��[�l��[�(\҃�̫���z4"O"!چ|`Vx�U��v���F"O\]x���Y��E�³g�fh�p"O�a(!��Y�FM��J :���E"O�tzq/߽6� �YW	�7y*R��"OJY��H�]��x�'U�C�րې"O��x�n���c'�/-��3"OP���&:�p��e�n��n,D� ��
h�����} ����j#D��
��W�UDc#��)+���+�/!D� ��f$06�Y�C �=?2�ⷠ=D�\S��ҟuk�,��@_?zj�2tn8D�(���P�-��ޓ+;.�(��7D�l����vC�-"r'H�S�(5{��3D�p�2&Ϋ���y�mY�S_Z�J��/D������0]���>l�X�#��0D�D�g�!l�(Mzq,�V�:��ŉ4D�Lz H�7ض؃��� ҁ�G�0D�\cEcM�}�V�P0"�h�j@�L/D���f C�C�tЛ ��nc|	��M"D����#b�T����؋5\H�	��:D��궤�:cv� Z��U�#�qZ5$8D�`�S-�<%�d|��U�D�9�C!D�XXeᇗX<�q%�F+K��1�<D�P���˾T�`ܩE"��cv)�&�9D�Hy iY>=)����+Ҝg��H �b8D�|B�n[�t\E��eD�%@) �K;D�{���7fWr����$E�.A�G.D�dJ$d�)������� c�а���8D�x�&�P�����i.	��	��:D��kd�=H�
�JAX&<X�je`9D����	(L�F�+㕼-�&*D����/�42�!c�:�p�Z3c+D���4ϗ�s�����Ӫb��b�>D������-I����� ��l�����(D�HY�[Z��1��
�I����1D��C���H:�0�X$sz�Iv�0D�t� f���ץ	�$"��:G�.D����j�>po��j��#�8񈐋,D� @�����s�
�N|
�²�'D��`�N�"7�UT�ݽ:}kTm&D�I����5j� ܍g�(��"D�� B��f��iu����M��>D�4�$�xk�r�M�m�Y�C�0D�L��K���I:v
�_v��ږh/D����J%V��1�ߤ�.�Б�+D���D�NSt4`a��~��Q�(D�4�B�(Q��ٜ�Ȉ�!�)D�0�r�L#qv�Î$`����))D��a�"X/sEF�zr߹n�rH���'D�Ȱp��	R��b� 1rP���$D�pr���w�Z��UE�,~FfLK�G$D����"9TΤ��EȚ�A�Z��@�#D�� 3�!�13�2}C�	x��9r"O2��&�@�]�����J=P�z��4"OX�A"��^��pq��Z<K���"O}�G�Q3Ell��](=��:�"O:���K'$�"	3f�&���e"OЅ�uI�0�F�jgb	 0n����"O�ɠkͯI=~ �v��r��"O�][r��*slt@�tK�x4���"ORT�w�P�Y�\ sc�@-+�Eq!"O�(��kG��:7���H
��1"OpQz5�/S���U�Uj����"Op�
B�Ϛp&-i���K��ç"O �Q$��!Y�Qu�ՋTѤAҗ"O.Xf�ȠNv�Q���$�0@��"O`���.8�2<�5I�\u��2"O9Yr�Ή=` <��;uL���"O|�1��!@����&C�3�]Z�"ONi�EȌMV �1�������k�"O����è) ���M=x��у�"O����J�>Cϼ�8�A����"O���,L$PL �����6�� ��"O���bL4,EZT� �E7C�~@�"O@XGH��4l�4��Wf�����"O6��U��Rh4�H�B�9�A�'"O�ṳFr�m�L���(��f"O*��7�+C�lD���9��;�"OV�3u"�+.HTM�,N�)�1��"O�=����l!�Ī[9�D+�*O������#R�,y��Z�xP(�	�'� 4�E��8x�%��|�5�	�'��Y���"Z����G�I5 ���J
�'f�UJ$�W�	RW�?%}&U�	�'��5�Y' V�h;�,���"`9�'Vԑ9��2m��!�ӄ
�y	��'�8�	"U3����Mp�K�'�K	�z}�g^�$���𓡎n�<A'�Um��8)�̤PI�h�)�m�<Y��a���`�� ��P�]g�<�fHLq�zUc@�T�C��6�`�<a���'�,A`��P�V�30�@c�<a���/�T�	�I�{,���� `�<����^���%-Cg�Ze�0�X�<�$�'6���1�C���K�^�<���@�Hc�m Ɯ�Rc��W�<IbcP�60`�醬Q��ļ�rj	z�<AP�%]�1 7ؖQ%n	`��P�<���Mg����f�gN���է�p�<Q�ά3���3e��R�08���p�<��
G�<�\�b �İD��B�<�E�ՂnJ��rw�E�Y,C&���<�6�%B�N�	���q��D1�`}�<qS��i|�q�ؿ8Ǫ1ѕo�}�<�&�+&�ґ���4�:@x�<����#9DV�i��L3- i��t�<IӋs-<��q(�q"	�eo�<y�� 1���h���|(��m�v�<��1Tr,�_��l�C�~�<�����+��q�憁a3H�G'Np�<9#�Ԩ�P��ʦIܞ����^l�<1��ºnJ�2akA=*�`��dk�<y�䂘�
�h&�38f�d�r&�m�<�	��t����aV�VV��9Ul�m�<�Ŏ�5H�那��i�����h�<�AR(z_\��1h[�So����C}�<� ��քu�0��ǈ�\�8Yr"O��3&뛺7d��f	�_��Z�"O*Q�.M�\r$�xb+��,�̅�e"O������Trt�_�V���p"O�kd��,���ȭ+o���$"O8�[�F�&FpM��1rf*�J "Oʙzh�=�f��`�؍Urʙ�'"O����]��҄C�)h(�3"O����IF&]JʽyBd�&8:a؆"O�p�a�={܄Ԛ�-z6l�`"O�ܩ�`˔D>�k��٦z5��� "O�]�X�%CLe^��"O* $A�7OA�L��1ib����"ONe�ׇZ� #,��a�D>,��B"Opi�-Aq�~ ��O#D�⥑a"O�h��IC�{�\�HƩ�8G|�x`�"O�QAg�W�|�;�&R�xԔ���"O�y��L�s��&���̡h "OF��n�����v��+1��}�f"O�Pg ��*�S�K�w����"O���ॆ�q�Č�cX:�άsd"O��@a�.�*�r�HBxy��r"O�P� �vV)	Jt�*"O�<��Ĉ9�h�f(�=0d�5�a"O��sueLDFx�DL/5>ބ�"O�ĩ3��4M�i���67��t�""Ods�E�(����T�U�Ȅ"O�9�1�.��vc/@853"O.-P���(c�)�C��b�"O~1`�/�IƜ5�m:-�&�"O,�I� Ojn*$������"O�Ř7M܃T�mh�d�#�l��t"O�m �FI��$��	�t����A"O��v+�n�(y��蔴K�"OX�jB$�&L�Qk�a#j��Lб"O��*wCA
��#���p�&%B�"O.�u ��K�D}P��"O�4��546���cJ^�Ĺ�"O�q�n�A�t�ba ��F�
��v"OLT��L�FŦ�[r�=5<H�"O�sm�"z$X�b��u0�-{�"O�	���	�<�P1��e����"Ojh���6��y�cf�5B�.M�"O�yԄD8�l�$�̢(kb	)b"O�	E.I�7��c���b��Z�"O4a�H٠fЩ��Q��"O8(p�Ġ]�TT���Y5N�i�*OЬ��HąB�hi��b�8+���I�'�XP�jݑ(q>a�u�Z�#�f���'E2�/[�mA �B��%S�'���%�Rp���!V��
�'xX��A�J�R�1@%����
�' �a�!#Q��C�Ã!I�Pt 	�'���j��B �5�4��/;��@�'[2����-.���;���,�q:�'������@�wf�hඋ^yh��@	�'9�Xp��Րx�>%8�/ݘlE����'����OI3j_��+�*�	O��Li�'w*mH0��*'s֐�gA�JX�=��'V|ڣ��<9G���F�����'�"�j3�۳6����'@	L�d-@�'���x��?R^,4JJ�J=����'�T�H��,�v�Qs@�G����'Ά�0���Pf�QCN�
md�1b���  U��L	�\\��F^&Zq�"O^�2"ПmezA����
Dh��`"O�@���H]��؁�'-280�"Or��S�L֎9 M��?�b�)�"Oh��靤��L��&JD�6"O�:�i�C�D�C���
8����"O�X�a��W�̼�uJ�@쎬r7"O�}h�E�/V�ԁ�#��h$ r"O��ْ���;�ة�Z�
����yBI
3
�lu[�Z]��� e���y�o�+tDb�C�$XrY�Dҽ�y��ђ+f����R9p��aD
�yR �R���A"�q�F��y�J�dw�A�N�'���L�y"n��x��%�2o[2h����O�'�y� ��Io8) �d��wz�d���J'�y�o�
(Av�R4ŝ? ޑ"ցΩ�y�%�fhSDdV�"ߒi!&���yR��_�̄�l�;l����I=�y�ퟒb-i0�n�T����y���L @  �	<�䓮?���|Z�[9�M��O�NE�	�&eh�-b���fC�=��P��O6hL>9(O���O���Ox��1���=�n	�ч�|��e����Ov�$�<AU�i������'���'��	��4���G\�DXDo�����J���ß��?�O��h�g�Y�T�a2 ;Ą:#������HU���i>Ợ�'`V&��0D//񃧇��s�F�k�%�����I���	��b>I�'nT7��p
b!��.�x����c�@��!�O������?��^�����5��cÂ;_�b�v$]Ey�������Ҧ9�u�Ƃ>^���$]@y"��Yc���q ��eܕ�JD�y"V����|�	ԟh��͟��O��l���_�h1�m£Lf0��mlӂZ�K�O����O2�����Ȧ�A��{wf7$��i�-�<{���I�P'�b>�� ߦ5�=Y�խ��Ig�ds�bC)]�đ�^�vh�dƬ��&�p����'�:̒�oNg�����G��9z��'�b�'�[�,��4;��I#��?�����1L�?���"�k[�0PI>y��.2���x�Is�I/Q�P�")��
WZY`����\���6���ͽ*�x�O~��i�Ol��RO\��c	�b7�}�!
)�$����?����?y��h�D��ِ~�
Q�d�܈�<)��Q�S��������0�	��MK��wό�����H)�P�	I�\=a�'KRW� ҩDڦ��'�I�D���?��� ��r�g�8/���Z�f<�!�%��<a��?���?����?!QO���Rd�6�B�9Ƹ��B�>���禽�i�ޟ��͟x'?�	�!�r}1��@.���i6u��e˫O���(�)�<)M�a[���Q"fd�%%"�:���e��'�� ��lʟ`ל|�\� CD��{�T$�B�_#"��2�E�����矬�I��SEyrm���0�x>iA�1� ���K�SD�u���O�l�B�&:�	�Д'yz< &D��F���R�)
K�&m�T�� `(����,�ԂӜ
�4��d������3#��������-K��*rNr��Iן����I����U�_4M4��&��AZ �� (� �?Q��?)f�i��i�Oc�(jӞ�O��K ,`&���=xI��G8���O4�4���ĤaӞ�Ӻ��V��B��
5d����a�uF��cM[x�މ��o�Ym8p9dY�5`�l��T�.���YB�u��/�I�b��3��%ymJ�[��
**�����D�sA.7���F�a��ɩ�B�]%1OXx��c�-�~Ї4kpy���(=��JA�Ƃx$�qˆ!�~_r )B��D|(���z,:�A6� �<��y/�<�4�c��<L����ŃQ�j!j��&hn�bg�Lvl��)���0"&�*`B��aE���E��ݸ")'U|�:�荛i�^��a�S����b�h�,P@%L
0I��a��iAR�'�"�O�Ũ`�
0xM �N��x���Q3+&�$�OT��Q"Yb����s�X5��8��rf
F3'D�m�ayB�S��6��O���O���DX}Zcm� �c��#�
X�CC��������Id��Ix�S�'c|��Ϟ�G��1
j8�m��j�����4�?!��?���|��Ixy��C� ��4���Ӫ3�v�0.���Żi>��0��8��ǟ���+��8�����T�aG:�MS��?	�*�@��U�<�'�2�O�5"�NW�B��m��"��dQ"�J�i��'3⁲�'��O^���OʩC�dPo>���H?�Z���
�	��;��8��O����7�5����@q���4D��M{P��1w�lM)�W��xBM���0�'B�'�X�����X&3G�9�v��vx�@��ˌE)�O�ʓ�?�K>I��?�����W��(���zQ!����6�jM>���?����D
(��ϧqjK�`�,d�����fUuiҝo�byB�'��'�R�'�,����O\�I��R�z(��M#'p�P�\�T����ByR�ƚ�맇?A�@A�NL�t��5}���N�rś6�'��'�"�'�6�Z��dŁ�4x�q��'iN�P�R)d؛�'o2]����������O��գ�`�)*��ؚ�D8� Y+F�	r�Iɟ�Ɏ-�(�?y�O@zu��:����im�����MS+O�eؑ��E��۟����?]�Okl*jtܽ!�J��:�>�9w,�5g��V�'�b�Ձ��O��>����ǚ8��Q�wØ"5Vn��o��@�g������՟����?M"O<�'M?\� 'c��S�h)�(^)�>����i���'�2�|ʟ�D�O���1� k��M�4G
1S�)��&Qܦ}������ɚRdڄ�K<ͧ�?�'�ภ�̏;L]j�
\*]����ٴ�?�I>��S?�I�x���4��#.�h%���!���$&��M��FB�P��x�O���|�%f�4Kt�Нs��U���ӇY4�O���,��|Γ�?���B�l�"Ƒ7&�n0aQHI�@T!(O����O�㟔�Ip?�0��+�:��$��B] ��T�����m#���L�'��f�	d��)Р�Jqr��^>�@xV�Jڛ��'�����O�ʓ5%��mZ�(b�ˀf^8#Z��#��0w$pO,�$�<�P���*�|�dCTNJ���/(�R٫5�#`���my���?)/O�$Px2C�k��
D�<r2�q�끺�Ms����OD��0l�|R��?Q��%�X�ϼ|�G�Rb�KP�5� O*�ĵ<�a�L��u�cļTg���gG�.�
Af厖���O"�F(�O��$�Of�$���Ӻ��F�Q���±�
.�"�Z�/]�����Ry�.�O�O~�i	$D��@v~��;�4U�������?����?�'��?�i�E�$fT`ɡ"UJ/�t�K���䔱jV�b>A�	$¾���!�/<B9��I�`F0@�4�?����?)�"&v+���D�'�2�҆�,����T~`�$�D1iҐ7M�O���<�\?��O:�O���7I�/J��Ĺ�![_u�`�P�i���8V�	����+�I�I�~Y��G��	����7,S� ���O<y��Y~r�'���'��O��,	�!�#JN����[o���&�(���?A���?)+Of�$�?U���T�q^d�h��|�CfDeӀ���<���?���򄕃C�\�̧ ���2�L�C�,����נGZ`@lZsyr�'��	��������a�(+�
A�l�ޥ!gi��*c�ǖ���O&�$�O�ʓd�`� ]?I�	�l��4FjL�Ajܠi�Ώw����4�?1.O|�D�O���W�Kz��O �	j���q"��c󀽲QD�5:b7�O��D�<)P	5 ��S���I�?�v�Q����̀�
OR�
����O���Oj��C�?5�'o��7]���/@�y��=U^��S�tz�H�M����?����
�W��#��)�%N�&��i�P#ѥU
�6�O��D��2H�Ifyr���'uD��@�J�N�
��f�23\�6����Z7��O����Of�i�k}R]�H#
� �9�P�F;�N@�rk��M���p7�i�vi��'T�I�P����� *��	!=�z]a�o;r@}A��i<"�'�bKC8/�V�����O�I�$F&�!�NיU�xzD�Z���ܴ�?q/O��0�4O�S矀�I��$I^�j�@Ð��~t��0$C�MC�pp$P�_�䕧oZNy���5FKS(�K�:7G����H>Gr(��'��1��'��	�(�	ߟ��'�|�V�P4g�%�1�r���ʀʀjM���$�O���?���?y��X3F�1*V��m!��ƣi:���?����?��?i.Oॠ�h�|"g�8Rd6 �h��`��d������'��Q����Ɵ����?�l�<n	�ƀ�N�`�2V�k�J�lZ���	����	IyBJ@7xXD�'�?�%`� y���Ae� �0�\R5!&h�6�'����D�����Oi����M�q)ÐT��S�4�����ͦ9��ğ�'�����~r���?1��C6��C�S�s4�уD�������R���I�<�I���"<��O������>A����$գ���Ѧ��'eR�c��~���$�O�������קu7��е	6IY. ]RҥX3�M{��?� ��<q&^?��L�'
]�����%���2�]8��<o� 6Ri��4�?)���?��'qx�I{y#��< `�!�׶xBhl�� &|^7�T�(w�$(�d$�Sџ؁�(S%n%0�s�㎫;���;�k�,�M��?y��/��P2S���'Z��O�=�VL�"��x�HƯs��=�i�RT����x���?����?�V�; ���bHB$�E�����ش�?��n
$ez�IKy��'��	˟�Ohą�%c�&�H:c!�:'���6�����$�O<���O&�d�^t+şR�L����IeeVu�#�M=���dyR�'i���,�	ş\;Q��/^y��F3��z��/����ǟ��	�<��h��'%Np�e�f>��3oI��x��*P:k��@դy����?�-O����O��d�1l���*�(AQc�O>P��j���&�oZ埄�	̟���Dy2Ƕ'��꧌?��<��� �M��ic�����Q~�o���'���'�b��,��	����)�P��M�6��Q�v�!2�yӤ��O$�}��p��P?i�	����Ӣ��Uq�֚ ���숀Q�Tyr�O��$�O���*%��ĭ|Γ��t��[�5����=+�XqӀ̂�M�*O&IP�^ۦ���ן0���?1p�O�nC=<�����_ds���/ӛ��'�2#�,�y�c�~Γ�OH�P�G �<����&��
 T�{ݴ&��b��i���'���Ot���'B�'��Q�ҧ�9t��`��"@X �Bf�uӶŊm�O˓���t�ߟܨF��̠�p`#�7\}��PQ V��M����?���7����T���'��O�MZ6,�|Jp�zfk��[\ ��X��'��x�O���O���O���/�$~�r]���W<��C�������I�_!T���O8��?�+O:��ƞq��*
:b��i����Zq��[�,�wFd�$��ğ�I�����y��Ӆ&�"Q�6�U�ڇ>�vQCA�>	.O��<��?q�m���2��^�b�,��D���IjƘ{1��<��?Q���?!���d� �A̧9~�M���=��[���1#G�}o�syb�'������ş(Ѵ�g� �4kKo�t��L�o��PQ%�'����O���O>�EʁI�]?Q�	oZ�`�ph�
Il��!N�F�6`"޴�?�)O��$�Op���=ZY�$�O6���^�[���70#^]�d-�����n�ß���ky�l����'�?����Qo����P
b;V)QElT�v��	������t�W�j���y�ޟZ!!w��b&ʸh�f���T���i��	�z�=�ݴ�?i��?�����i�-`eΡ1�t�b�0B�Z�I�Cj�.��O>�9OpH��y"���P������:-���(W2�6��W<�7��O���O���x}"X�h�E�k���q"�d������M�gA��<I����d4��џ����W�"-X҉ �,^H���k!�M����?)��_9���3T�,�'���O��y�B�nՐ�bU�V%6����i��]� �p�c���?���?q�Z�w#bQ�JN?_0Pě�!��C���'����gd�>y,O��iU���"�heAPE˃w�h��w V�#���HĨl�����O�d�Oʓ�$$a�޶J�n̋��$��l
:(�InyB�'g�	�t�Iş|��_�u��_.TMVi���Z��������蟔��ٟh�':r�� �v>�[�/A9�0��A)�%|Lx��g��˓�?1(O��d�O���)7���^�����>@�ZHX��	/Ѻ�l�ݟ��I؟��	wy��שY�"�k�Ι���)�H �*�&� נٿ2�&�'��'*2�'l<��G�'��,b�����@�E����,A?��\l���d�IXyB/ʟ1'��������[C���!��i�~�L���_}�����	�~՜��x��ʕ�Ȇ%���Bɋ�Q��m�Ӧ�'�0� �fӨ<�O���OJn�W$p�gŏY$̹Hpʦ��ğ$ �,a��&���}�$"��N�@DA6��
�Д8q�AȦ���k�$�M����?A��R�x��'��T񴪕�!ܴ�0��n�6�P�o|��{���O��OT�?��	�V�L�B�kC�Ec��6��'H6��޴�?���?�����l׉'�2�'���E��~Y��^��.8SC�HǛ��|���6����$�O���C*,?�0x���5N:*�"$ɹ�-n�П��kG���?!����� �YB�oD�t-N���M�k�`��U����v�P�'���'�R]���5L��dM���AK�5r;|��Ǔ2/�xQN<����?yJ>���?iu�]�FŸi���α���j�p ��͓��D�O��d�O�ʓg��@02�l�!4��8sD.\���=`����$P����ПD'����П���%�>��/B���� %�*#gB���{}��'��'���.BK�dKM|��P�5�ib�!P����+���%q����'��'���'���'d�P$����0�1���1*^n�՟H�IFy�m�(�v�.�$�����O��0鈩�ա�֑ɰ�\�	�I�K��-�Ip�I~2����XAb!�J��V)Z��U�'��Y2l�"E�Op��O���4���{�%�z�h�P��PEto�ߟ��I/[��O�IMܧT��H�qN	* ��H;�jT'@Cp�nf�eZ�4�?��?���0��'9�G�6����˿<�6$�Տ�Z(�7�O�*G��4��&��˟,��i�(brvE��h�RS`�i��V��Mk��?��]en�j��x��'���Ob-�t�@!E4�L�2�@0 "A@��i��'c����)���Ob��O"]@!	ǹY�>�(Ď�/��t�Ԧ�Ŧ���B�ڱۋ}b�'�ɧ5��!$�4T�"$�&�a�� ���-*���<	��?������	<@��L��嘃a�2G�v4����T���h��}����l�ɚG06e��l�M6͇kĎd(�τ����?���?�.Oްy����|2Rk�=�ˡ��f�B��,���O`�O���O��)� �O� �@�]�Uop`�R��h�U��}B�'��V���ɳ~on�O\���C[�����u���°A��eĚ7M�OV�O��d�<���y�I1|�N�#�.S!4��:r�J`Y��i���'�剫}�� M|:���w���c+h�y��˖5?pEq,�d��'j��'��) V�����RB�(/U)ݴ��� �'�\Mm���i�O��
T~���j,���B��N�RO���Mk��p?Y���3X�0���"��.�0�)��ʦ� �Oӳ�M����?������x�'�!9wm�4.W�� ���
�a��g����	u���?Y����
6iz���q���O�� ����'���'��{S��'�?�O� ��A&ƺd�L��f���h��-�	�I�,��J|2�d£O�R�!D2O�ŪB�� d,�5���$.�h�� "O���C���6�J�N�R��F�'İŸ� �0a�9�g� k��� �f]3h�B��%ϒZ�vӇJZS��c��B|���d�U5w��Q@udX9|���J� Ąv����L�G�J�A��Y8�@���х1�6Yu/�^U�us���cF7J� ��5�*��d�Ѝ�F��$:L�an�.�Ԓ7hG�A�r���ES��q�'�RjنP��'x"�y��|Γ?a.H��q�,!,�h)�p<9�H��'�H0�G�W�wcP!��%-z���@�td��c�V$��񄃅S���'ɖ�C��jw��=
�fE#�\&PVj����t�	R����O1b]���Er��ݫ�A��D����'�D7-�(#^
c�J�AJp���86�Pm�Fy�	R#���?	(�p3d#�Ov丢�O�xm�\I�8w+#ˢ�?���3̑���Õ&I�s�e�<8�*�Dʧ=�2ZS��3�z���*4o�lѥO�I��o�=x�bY���\�v#}��%����D�쉎V�,���WM�D�r�'G�>���$st�19k�9�R�{dL!qC䉐:�΍j�ʜ�J�zUx�&����E{�O\$"=��"@#Yx���V-D�-��L�ą[1_��6�'��'�����!ҽF�r�';���y'�%1��e�vΐ�8�.�����u<�RKR=]����'$ap�[6�|���%pm��f��.�J�KR���NTD��$�kh���=.�\z��T�Sf�������°}#&4���Y�������ą�(�O�ўx���*]lh����n�x��j2D���%�
�2��EW���֮k�D�	��HO��OZ�z�rX�G��Q��h���� K��U�@l���?A���?�G��F��OP��c!>T��E\�a�iZ�2����#���>x*(a�����=Q'��V[�9y�
��/P�;Q�� mJ�V�X�d�����'�l[��+s�l�٢D
�Izg!�"�?����hO�� c��ޯ<Ȣ)�'�
�SH�Y�0D��b�cV1CB��� �]��$P��.�	��MC���Q�_�m�ß��I�,�U�fX�%�"� f�K�H��h�I�4�"�ɟ����|
�`���$�� 'ϩ�,��L�L�n0�W�,Ox�33��DE�h��-4_�Lɑ�#=o}�x����?a���򤀡V�1��G�'��ac$�@y�D�Ol�=�)§1�dQ�4(M�a
B}0"��93�j���N�6������2h5@��f�غ"S����ߡ�M��?�-�|t����OT�h��7v���@f���������O���H�8������d�|B*��U�ꉬpV=0���
�j4�ԝ>��j�E5�i�O>�� �D8�̎�\_��I�!�#��Pub:}�U��?A��?�����O��]ó��e�dѠJ��j�ļڎyR�'��y�̝�S�:�ٵ��<Qx��խ��0<�#�Ɉ]Gn���K�4`��v,I�ި�ݴ�?���?ِ��M"|����?Q���?�;G���rF˗�h��ٻ�>��@§��P�|�8�{- ��Щƿ��	:�ɾ=<��c2l��u��it�,gk�X�Pe�#��=�!ךwdܣ�f$��3<S �j5O�и���"NN0�ⵍ",7&�@�d�O�nZ柈R��F���>��?I��U�
S����ʶB�X��!���=�I>�d�\E�Q���hT�`j�F�<���c؛^\��|��
i��P������/g���hX�t�bV	>D��"� � `�@+Tj$u�NȨ�I)D��j���o�<(hV�N���ѩV�'D��H,'�  ���Ez�5C%D����._�'�[�I�fCx�#��>D�<�T�X���qG�ŪF}p��'>D�����#X|�4$�hL��D$(D������@k�`��/>o���w� D��q��(jүd��d�V?D�hX�S��rED���rUn=D��K�Ė�i�,�A�#A��Yx��<D��J�Y-�!�;-� �(.D�T�e	p݆<Y&�#��(jw�/D�\p�j�F܎U�a�ùg���3��9D���&�ۓ/�$1"��Ý���ZP3D�4�V�Q��lZrI�5W� l�41D��x2ϔ$>��$p�f��p�� *��:D�0:d�ؼ m�X8c"��D<D�L����0(����	�� ���<D��R���q��qM��<J���8D�ܳ���Kc�\� ��q��dm8D���Am� b��4y���=`C��d�04RŤ�=&�h��s�"C�ɪ(M������4d�͖�U�C�ɛj;��AE� 6��WA�>J)�C䉇S|��Y�$�/��y@ Z�dC�I(GՖ�
)��L��xv���B��8u��+�kR1���ħܯKV6B�I����!�&�|(C��+B�I�d�>��!��/,4�Ц��#<�C��1,\՚k��c�āZ�M�C�Ɍ^K�E��K�8=�U��$��y��C�ɯI&a�+�%��ђ4�fB��04H�cȪ_��1�6�C�	�C���L�〽!% *i㞰R��p<)6$C�R����,��`�h�](<Y!ϏM+�<yg �}!jX��E��t��ܘ4b/��k�B�)��d��JC�y�P�$�0O��k�)��'4��;"@Q']n�u� ��}�&]�
�'��Up�'�_�h�)�,$qmF��J��2� X<L�qO��%٥�Ђ#䖘�!��׶Px�"O���Ζ�Cw��ف!�,tj��[T�D81A���>�!j0�Z20�&�ܖksj<��� �8ፈ�.K�<�	�=1@�Yڶ�^�֘B��0\��%�О
��x�ȝ3q� ���<�I3R�� 	�̓�~��A�[�O��B�		^����>l<!3�!&/�B䉂 � �J
��r�ܠ�S( ��B��>Նܹ��g��6� �yҋ�������]���&�u�<��eȣA�H�V��z�؀��e�<a���Y��@i�E�=��E2��^�<B0���B#1�y6&Z�<y���N��1m_<F�Ay&�QW�<��[*y�
���8b�0=)$�R�<� �	 iH&D�R �_�,B,���"OF\ T��%-�!���#L1�#"O>�k)�	�I� ��l�z�"O�I��T�4�eJ֎ۙ���D�'IN�)8�	� ,����B� ix�!�R��cC�I�3�����GY�g�yfϗ")��:⋉�?��f��c�l�)�矠C�lL�X��� .��G��HƎ+D�hK&M� Kk�q)��cfL*�Gk�����Ba��,��M��H���q�X�U�ȑK1(0��&D�B����A%t���4u�H-!�iÒV�(�CcB�e�2عd��F�&B��$s�naD@
 D�))��A7y�"<�"G� 	fV6�- ]����J<u=&)��&� ��&ބ�y2G�	H�D ��!؀ע]�y�ę� EЦ�r�4���s�(�/%0cT80��ő:Szl�� <D���CY86|b!��4xp1��}��a�/F1"i�f�*.���i%�!�-E�7�4�ٵ��
�ꔇ��&c�d��W�ik�0ڰCV��X`A���<���2@j�	3t����v�^�;�+H�R��- R�Q�k1�UExr%��jmJ��I�:�������g~� �n�~1�L���,�y��[�+Ӳ����Tp	�`��ܼ�6%�~�ӺK�e[���5�͏V�܊V�a�y��f�y2��>*&P����A,O�(I�FՂ�yb
�k����?��큣��'��D��e�,�Y$��w�
"�Y��PR��2���K���L��{�V>�[uJ�=�Ƞ{���pG�Ի��f�N貃J94o�XB��ٱ:7�ܲ�R>��>�%�ƖU�۵e��J�#�ّxrH��m�%u�'��OK�>�M�u,��>�!k4��6�� e����]�2 h0��>vl�!aၧ�����N;�dB\c� ���$u�d:�J ,������IP�FƁ�?�փ�m� S͗,�9��$*��=�x������bǸ,�<ٕ扎"G�-I h�d�ģ��/��'.��2�Ɣ7�t������fKN8W��Mgg_zT|��ț�q�䄕O���R��ZFؐ�O�I���/&Qtۦ�J�'9d���i�H�`MW�-:��{�K
��L>yΟ�rD`}6��!�ճ	�ع�Gp}B�WqnL���_b 8 \?zl���d�
�8	y��?O/$�*D혜���������'���Q:$��k�$�U��.����vm��TD�����:5�����/.W�xJA�;�|¥ȫQ�j�!d^%6�&��s =E�0��%D_��?awcҿy���Q�'��0��;�~�:�����'6�FlҕC�-\h`��NB!�y��H�B#�`������ʕf�9OV�S�\�
��3X�T�(tlb����ʐh� �"�<��A͌ћ$]��:�Q��kOl#���苓�j�����`��2*N�9{�V�/ZЩ�v>�O��'R=�;�)O1���s�	/~hD�'9
�aG��W�hy�E/�^Ȝꐫ ?6�qO�%H"�
�urmc�i)Y)ΐ`JK�db�A�T�|��	2��hJ�@5EiJ)���9v�� Vʒ�Dj�QP���l�`�ac��!%qO�	Խ��;$�X`���ͪf9~�v�8 &�ym+LSԵ[�$׏��v�&�j��
C�I6=)�$ˢqܐ�#
y��c���'(9�Չ�lób�q��D�43�19��)h� t�w�[�
�y��	(; u�s�K�J��Hq4kv�ah��C1�t��b�+��@e��<��'k\�B��򄊎@Z�'{�\�D��3���⴯�x3���L>ᰧ�78���� ��%T*=�t!Lܓ13f���ND�S��(#%�(�j�7k��XjD�{���2+��#<�$E�(���[��L�~;Ph�`mN��R剖�Șu+���5�)�de^���1�cB�u���(�Λ
y�)�DiPC�&�Y#�Ϩ"i���I=P�&i(fŘ /����� S�]Zu�<��C��tqg��"֌�>牁&Q*B��Q;,�*A9�FI�����AlE*@;�N?	|�j���7R��B� }�$����A?���z'�	T�p�#�O��JQ?��$w�1�O�<���aF�_3� ӡ*t�a�r�|�
4��`�v���f��1�ݸ'y�������?��ذ&�BMNL�O�����'���$Z>�Gx���������)G-v���%[�`���?]_��p�j�H�S�)K(�5޴a�:8�a%��^�0�#+Y�v�b���X�R���Ui��8b��ʼdc|)	���Qf�@n�M���Df.�)b���W���g�A�/�^�ʅ�.�~�p�x����)Ƿ(�d��I7��Iۆ6��L���� @�q(FD�� �lj�{"MG����o�%E%�W�S��I�Hq���`,F^��1�U�'"��d�?MFb���ujp �I�2�����'��豈�"oZZ}�Sn�~	t-�ÇP�^�)�ŗ{ev8�Hǒ����O����	��!:��9�	�ʺE��b �0�0����#��!+���S�.Q&�!%Ï(��$�4	EwD�m�;���`��\�OP��t�Pt�S�\c?ppA�9?���	�gS���{�y�o6
���=�|2���8̤�gN'�hu�T�	?gpht���d.�3zq�� "I0��<LݰI�aQ�p(�,�$cY�%��R�)�ӂB�"��OB�a�"�M���Z�I�B+ě�~�gڷ7�(DE7���I2cSZ�9PAڈc��	 ��8Rw�$12�վC���:��OƐ����O�s��Z�J��'ٽCό8��-q5�P���T�=�Q��9�Ę�^\"QS�O6\��e*C|}�7#�#m/�ܚ�f������ fܖ���gVZ�4�Ѐ�[�
�l���� ��*#�� E���('8���fiPV M	��Z^�@
�&h�	�?tz5zŋ"i��I�R�P��W���)GD�{�,M)Y�3&@U;:Ѫ�p�H�wHҕ�'*�Ћ��$ό��xc*h�� �8L�AG�<UL-�3����sdB���fb)Fx��

|����A�~7��W�)J��ď^l��sܮp�쑰�g�'y��j����O�&l9�ɀ7y*��B��DН1}4}c�n��.�7/��8��cݭyƒ�YU H�AU�I�57�I�nE�`�T�nZú����yo�(�B��8��M*`,9}�b��<)d$
=(bܒ󮛒k�ȃ' �D̓>l���Fc���"����ş��'��2���jf�� �6��t�H��s�����Y�<xe�`䀨
>��KBЩ>L���'�G�O����+8O��
_d�}K�-�PLV�QȀ�1�,�nښ/ɾ����
�
�1Na>#>	�'ћ�U��(p����`8�|�Ra/�1O�!V�\�x�8dC �S�$d�n	�p<���r�L������U�qꚫ��Q��ҝR��)y�j�X���+�b��G-f��u⊋Z�D���Ի"o�	x⫗�1%
 �<y棇�q�
��A�>@�)�Ί`̓z[\�`��Q��ɡ �=j�Ԙ�?�C%�:Su��(�ɀ-&#���GPB���1��#���:����D�%��''bH��7 �n�az2�81q��C|o����
�FCވ���37�>%��n���X�}�z��,�N������Zm�d�=Y�`�����ɑNlx�� ͏%-q�,���F�����'���[rܧGt��/P��j�'ȄJ��+!�����Pۓ9� %�����mD�yٜ$p�Lt�����63�\#<�b���s�8K��<nh ]�1��A~b�D,\7Z-����gS� )q�A��'�.9
eʎ�8n�X���N��N�0��a�X	��b�.:I=SA�x�&���Ț6n2�A�l�U��������BӅ^^�0x����x�gYt��T�1��'^أǓ�>�y�J��
�|!
0n� 6�"w�����9�*�����(5��+S.�L[���p��<�^�Pۓ:���/���1E�H�gE�̐��1I� �#5?�%/�g���<����+�:T�]e��hp���R	Y������=�k L��q�-n��Y(%#�1U5�͓[�����1��2��ܨ�r���*1!X��A�h��ɍ7�Q>�	�)��`F)8��i�Ԍ~Ű�I 6�d���ɿ�@��S�iK��S�'�����.<��lQ$ƅl�I��_p�;Bo�`�.�b��'�p䃧��;d�S�\4�0�aW8:�����Q�}���CDk����4���� ��)_�Pu;Pn'&�!��9�p>���C�߁+$�b>����R�V
��܀Ҙ@#��_�_/(b��3�	�s @L8Ğ�KD��K7�^��#>aw�Ig�ّs���4i�p�C�?�kw���,�PiҀ@�8-�� D�xp��l��`�XE5ٕ���Xj`+�$+��(Ơَt��F��������
�x�JE�v�X,�y����s5Z�
W��;^�$7��y��
`�t(7�J���Cm\��y��f~�Y�'(C(C�<�Q���2�y�"�#"���˅'6�� ���yR��4���"���hq�T�y�B�?�� ��B�b�1p�!?�y��΃wڔ�T+Pz}!�n��yRd��|N��TM��&��32����y�	�1x���%%�XQ� n��y2GM�?dƽ8� 4J	�W��yrKE%tG��2 g� YƨqT�1�yb,�&���� ��F%;�y�O�7w%��r �Z�~U��+�_�y�]�q�����DD:@qSe�ٟ�y���<��P+1BN�;���'J=�yb�_�V�B��*O8����ą��y�"X5'}��C�m�0�޹����y� Aky2��q�L�+�J��(��y���b�ɐ Ā7r6�l�`.��yr.K�(�rį!g�:E���y
� 8��A4��p��ͨa�JQ�"O��0!�.R�x3c�����d"O2$����1@��Ua7!@�'�h %"O`��և	�gx*��m�����"O�QYW�]��D��u�.�`��v"O�(���&?*�+�e�G��9�"O��y��p,������)d�`���"O0��[�I0�,���,ζT"O��xn��@�4�:�އE��R�"O�9񶃒837\���΅�D̖�!�"O0�k�2K2��4.�>����"O.|��$�턔�K��"	��"O��	q�Z7.�T�{`��	T
4�W"O�ؚ0k";.4iA�\=B�\�ɢ"O�ܫr�@<<$��r#ـ8� �x�"O�!Z%%��|����S��E��\��"O���$��7�IFk�5D̎���"OT���F+<'�u"��ڮd��M��"OR×�Ԝ�U����G����AJY�<�2�P.ɸD{!�4&D�@I^o�<�4�^�,�B�+��L�?�����B�<�dΈpI�`��.K�/.&=�ψ@�<9�`��="�sq��y� -�G�q�<��K�7݂��DK[O"��F��o�<S��>q��X
4@V�蕈2b�h�<��h�c�
9�C�]PB�T��e�<���\�@��$�w%�u�䓷�F�<񐮋�A5DQ⏂�L�ZX{�@�<�5�D�f�%z5BJ�I��|�aj�B�<�N�4w���(+M厹�n�c�<і��	i��H��c��{� H�A*�j�<�G�D>�
ؑ� �<N^)��	j�<)F�\V��B�I¡]甅�r��k�<� l�
1�&Jm�vyJҁh�<��A�|s�)�"��2���d�<�w�B�������X�����\�<I3.�0T�|�I�,�C`@Q ΏU�<yAJ�EY�`MA'h�
U����O�<�aN�6b��HXp��#�♩w�N�<�u�T+_etY34	T.5� �3G�K�<�F�*bFLі@�!Ƥ�Ȣ��H�<q�e/?֖�[F�ܢ<��40��B�<q�i�:8d���*T)���B��~�<� ��"oX �N�"��T�ǡ]E�<qb��[���y� �"����/_K�<Q���#��вNȈ��qH	E�<�V*E#"y��Ë��I�<��AO�U�<I�.ܷ/-|���%Q��ږDO�<�t�ՅjX���ܷU�>�{�E�f�<W�So��I������ @C�X�<� �,1r QR�Kd��h��U�<i�k^�mTr�S	I(֜ s,�|�<�q�+5)�b���mX$T���s�<�d�X�mLu1���&0�-���{�<Y`F۵j0�j�/H�d�0��D�x�<�h��L��q��86�ب�"j�<Aĥɟ+0A;�� o*��!�d�<�q�S�R��U�# ��2Zh�bE�z�<)�*�RYp�LP.[yY��K�<Qs! ��"4�E#^17.e!DH�<���	1B�l��Ů��H������L�<P�����ӣ��		>���l�<aA/@�<�$ c2n˓} ��/�@�<W��6��5�#��GH�����<� �b��B1cJ��Ҳ� �4��b�"O"M� �H�IXތ����5v��(J�"O�1�
= |�а#�)i�P�"OIЅ��0l���$M�Y�r��"Ox	�	6O��@eŇ?�:�Q�"O�}3d��~b8���Ē&��1��"O��1��ĥ)�������g��p�"O�����߃3�t!LW�1	��"O�|A!bL�y�.�ö)�\��(�"O���a�Nwی̫�G�d����""OPY0�ӭf%Zd��*�`�2�"OJ#to�`t�\1pBN�4���[g"O���H&"�pu�v��X�J�h�"O6d��f+�Ԩ��A?m�4Ȓ"O��2t�ӝP�ZU;E����$(� "O�D��O��&�:��I�(����"O,�q(#@�n� ���3��9s"O�9�ߺD?d<�������]�3"O�TK'J����+@�;
�h9�`"O�m:�N_�w�9#�%�%U�i�w�~����Һ)5���E�2L`Xb��Z�n�!�D����	s�:BX����BR�c�!�dI�3h��H��sYp��X�x�!�DݦV���U"Y�^����vE͊e�!�$��Yu<�!��#��Q�MO#�!��u��eb�U�V���Hb�_e!��n1�0��&Y�� �,��:�!�W�.��@%͵|�Es4Y3H�!��Q��B$�l�¡�d��!�M2(�����)O8!@��W�:^�!���y%"x9�n"S[��qU���^�!�_���tE��kN
l���گV�!�ċ� {Q�([1�lepT��	�!�䋯��'���Y7�DZs�Hd!��QYQx�Xw��(Ҋ�qc/��!�@0|�����9V���C%�N��!�d�./za[0�}��!��lˏ$�!��Y�t�De�(ٗ��pᶫ�?=
!�N$4Ǿ�X)��}�bJ��C'���,����k2�� #D�%�ȓy� ){���L������'T"�"���s���"��?���"F�d�t��*3D�T*&�Иt>��O�MK`�Xu�2D�|�(Uv d�b�@�g���U	1D�H�5F�)�́R���*.3���*ړ�0|:�(L�K�,Tt�����#�pB�	�r�,8�	��
@��"ܵv��ʌ���O��0W ��z^:I��ǒb*���q"O�����! �̬e�@�,Z��@"O�h;�L�6M@(�хI/H��UW"O.�aD�E�����ҸQ� ��"O�(Ձ����dBJ��XH�"O8 ��㊆�Jq��H��0��"ONm�J�x8h�qc�{�@�� "Or���LV�L��5!��K�%���i@"OX�HcIZ"R)nAQN�
ǶLR�"Ob�r�o�*��\PC��6
����"O2)��E�G�|�ӫ��II�@�&"O��ED�v�*��L,���w"O �� ��:��j��z����"O�Xk�&���,��T�W.tp��"OrjB&P85�d�:ak�h@fL�"O�I�u�7�8(Bq�\2VI�q"O
Pbd�.<:^4���7.��%�"O� ��ᤉ38MR�$����*�X"O��(���Z"T��!�E9(��}�"O��R��_1��6��[�N�@"O�x��솩j��R�-����"O|͙�,b�)�%ŏ�\s~�K�"Oj��b�Ǻk䜼)���z{�tb"O�� �A�"#�́�ȇ,���I$"OV�;B��g���h��G!Ј��"O��c�	Veʁ�a��|�x���"O�aCoԵMt�˂�ͤd��mA�"O:����`Ů��vFH0U�����"O�´�^Zp���z�(;�"Ot�h�'�:{�9
���z�w"O�����	"��htę����A�"O&x�Qb�t���q��9}��H""O8t�`�! �9�@�N�.�r��"O��� �S-v�� �&�?	�v�Ò"O����n0Cmh�AS�V�w>^���"O|�F�?7�D�����gF]�"O`����/��	3��[�d��"O0P�C����� ��\�j��d��"O�Y�ĝ�Ӿ��vnĉ/�1�"OlD9��9���ђ��  r���"O�Qp/5mDkЧ��.����"O��y��٪XJ-�F¬s���7"O"�PE�(lP�3k�[Aʬ��"Oz����s� �Q���p0�X"O��JA Z��L�!r�ɟ!���"O��6�>x/|t��( Y|5��"Ox�I��X�Li��P�P�H�|k�"O|�gDG1`�@�!�I����@�"O&)�`'q1�	����%�L�v"O����d�5��.�r���F�>�����S�@�@Č'LF,M[ ���7	!�d+�`@��	�dKfհrN�'!�䒦3�P�2f�,�vt��j\�S�!�D�^qh�a�;O�$�'gK��IM�����EGmt�i��O;D��"6_-v=��b�^4�339D�p95n��Rt���t��h0ܢsM6D�8��[N<��#uf�W-�ͪ2k1D�X�eOBpX"(x�P1( ���0D�\S
B�0E�`�E.�&7��eI��0T���5�� ~CʘS6HЀ�(9��"O���S��	<��12��h�E	#�'Α�Jbȅ& 0��Ra�!1����0D��Su�̴q�ܐVE�:_���aAj3D�\8S�ݨr�h�H�%ڵ>�^� �H1D�`eÝ0&H�����;05Y$C1D��B��Q�e6��q�)/�Ż��"D�(��Z�TI�H=x���� ,D����M ��n�[�0!���!�a/D�(��L�*��e�:`HѠ2O9D�,yp�>h��peCO�D�Q�T�5D���c��m�±G� }'��44D��dC�MeL�#剭f���#g 2D�l�� ���������PF.D��K��R�y�ހj�kʨ$Er� a./D���sW�9QZ�$K }�F@!��)D��XT��3V�TmhRFJ4 ς�c�<D� �7�ʘN��ip�\=S5̨��>D�(A��	�<�xS���1����>D��r�혬Or��nK#h�@�	7D��*�$K5���a�ȼL�2�0�4D�� Չ���I6\}���[
�����"Oi����K��0�S�E�C�X�1�"Oԅ��=f� ј��_"q����"Op�ESh!��rRMC�U���H�"O(�MB�@<��:�k9)�  �"O~��b V�Uߦ�B�ȜB�$�$"OT!)��� �0� �(X�s\43�"O���GF�+, �F��2��2�"Ora+qb�9m8��ׅ�4����w"O������p�GoԞC�6�0�"O�cA�
>�n�2���e
R"O�! Ҥ��Lgh���Ѳ#J
922"O4�)��>?��Y�b�x0�Dsr"OT�'�H�W"������{p��F"O������%8Y����u>48F"O�L�bK^)(r�����PPr���"O*�B�˘|n0#��DJ`�bB"Ol�!���+�Q�"ՅH����"O�-�&�m�4�Q"O�8>dv"O�*#�dܚـ��'�H8�"O�93S��@JxCA��ƥca"O���͐�9�x�p���,1�L�1"Od������t��ఓ��b{��y�"O\�#���6lxCD���wg.1Z�"O*Y�ժW`��L炠LT�l�1"O�Q��O@�T~\8�c�Ƅ��#�"OƝ"�?[��rD��n��"OL�ju`��*�ǣu�b1Z�"O���C
�+t�l�"C���B`"O��+s�Z�h-��q��?J��4i�"O�p�1�[� � (ـ"O$��n��M�b��OO�Xd`La$"O��P&A�
[����.>^ܰ��"O�"�Z%l0��C�ϣNN��zV"O�(@s�ƾXl$4�6Β�f�e"O<��eI"6��3͆�L(,8��"O�;G��O�Z(�Q�\F�	Pg"Ojm����]�~ /t�qE��e�!�dZ4 �(��Gȗ6M�fe�p��b�!��A�y/��g$ȽS��xgM+�!�P9 P$��v���"$�91��p�!��W�_9�|��×�?7䛵��0�!�d�=���P�|/&K4K]�"�!���9b�\�W`�,&s�J@/S�!�oԊ�q��O�4�u��T!�䊻	������/��M�T`\ WO!��Ҋ,����k� a���Z6R�R�!�DO�d�ꙣpc�%�~Q�*�F�!�D�<����)�(q�:�'��!�!�d������&H}�a����$�!�$�%w.D
s��$%Tf`ȥɉ"�!�DĴ&z�M�xIz�3��@�zR!��%@�vd c808��QF"��y[!�Q�D$�B��,n�n1���E7mO!�$�u8@���&Q�.��p���kF!򄑏MEN�Ҵ�!=�b���`W�!9!��̸+w��Z�o��_���U&y�!�d��"�ˢ��J�9�DI#s�!򤌎GA�Li�φ1B�Ed,[!�$ԝ�,zǊJ�*#�\�CL	.[�!�L��С "�a-*�@��X{�!���u��9��PI�*ek!�dɌa��|Ԫ�	jM�A��>�!��[���b$�!�� �CL�*!�� ʤ��M��$L�)PX�m� 8	�"O��p%�6Mڶ|� .�0<�.��"O�I�A��(氐W'k����"O4�� ��>| l����R�^�@T"O|���.u� ���5;�M�a"O�8i��޵[!~��d��y�v�ҥ"O�t!]�bӪl�TI��>ڎ`�e"Or���LL�H�P��j���T"O0���L\,^�9�@�տ:��p�r"O����m�5:���$��e�v� �"O�����9��xS$"�"Z���
"O�Њ4��'���@`&��b����"O �[Jԓ|�xD��D�w�plI"ODD��)����0�D�j��ط"O$���]�%`���~YP`�b"Of� '�X�d	P�!D&hc��ɰN0D��;#ϺI�=�Sa�<���6�9D���Ŋ#�4ݸq �u�����9D�t`���?_4\�ꀷ
�ε4�7D�d��j��?&�8���R�}]f�#�o3D��a��ȡN(����l�`�i��2D�r� ^
I����a/Z�}�<iTk1D�|z�!O�vT�ъAA˯ml
��C��
`�4,� $(oxP�#�@���B�	�r(�4�s�ȣ3�x]3��HM�B��	kt�����N�`z�/�MyBB�I}�5�䉙�u=�c�(S�B䉶p��SPmU��9"s�Vd�C��A� a;ᅏeXdy��?G.B䉔{ \u*����Z�{�'�#� B�I�>��"��͍FG�!�k̸^5�C���kTE�ogځ�@e��H��C�I ��P�_�]A�T;�˗O[VC䉏F��Q(�

Q�|��	�'��B�	3mHnmk�na
-��fՎ@�C�I��Li�dɋ�]<�R�Э�B䉉R�Y6ɀ	�(Q ��RM�.C�ɢ\��pM��:�
5��00z�B�%H�$|�/�1-�(��e ���C�	��X�s�j�/�t'� �D@�B��*t�(���ճ����Ph_�:0B�	t>E�� R��H�%�.&�C�	�77���V&`Nz��L��tF\C�I���i3ց�v�`�cf�J"�B䉋b���NX�y�2蔱!�DC�	�#���(�"� A��\"cᔩ<z�B�ɺr�P��e�Ǟ�"��j,�B�+d{ 5��'s��h衉�\�NB�I/\r��hE�x�U�S�]\*B䉺h��	�� �H��t�O�ge�C�ɔg:AQ��4?z�*��\��C�k �Mb���B%z��5��C�	&t欥�V���R��`� h]�jpC�I
L����G��	�A8��r�B�I�:`LA��(;���Į��C䉗qa`���%�Oj��@�  I6�C�ɱm?~�k2D֑7f��T��%&��C�I�+�bP�v�RLA4ap3%��X��B�	�%)�i��h�]����ةhf�B�	%*Ѐ%P��A����*f��B�	6,�J%��%��q��ÇK
/A��C�	�vu`�B�*Uh2���b���!g&C�	+%�,}��-Y "���I�/�]�B�ɡj>�1p�A8F��H��\3ӄC�)� ����j����`!dY3m����*O왺�MQ-��+QZ3E@�|��'��v$ƭ��x�q��!��m��'ߺi&�(��y1ɒ�{����'D�8�$��c���0(�q4L���'(�D@��ͿC�x�'�+l%��	�'
�+�I.-��]v�ůw���'`�%�b��2��5�H�GV͑�'v$L�t���X�k��h*p��'��l q-��%�^����	Sl����'�tC��H�Q.��a&���N��i(O$���̓x>��(�9)^�i`NԲ0�!�d����#'EʲLF�Z1螑�!��#+��i�)%��IB逐�!��NP5N�	B�'M�uq�S�@�!�W,R�H�� :[�B��d�51k!�L�kS�Ƅ�� 3;#XAR1�+D���
T�8�X�G:d@�����5ړ�0|��DA�(.��H��(S�\y{��\f�<yRJ-S��}ׁ��G�<��t�JJ�<!����nG���G��hϊ	G�N�<��kʞ�v��T�K�n�ـf.M�<���2Uu���7��B��8QN�F�<�b���L�|5 �A��?�0|�q�C�<!D��3�^JA�Fi�D�z� �j�T��9��RJ��Y��H�k^uՄ%D����Dy~N=Q$�E*R�&1�f/9D����kѠI��		�m�����Sb�p�<��'SR�@SO�K�5��Tm�<1�cP�1y"�i��ݨN���I�DHf�<��e���5��4(�IfI\M�<95Ǘ�nޠQ2A_b�X��a�<!͢\� q��D�1���WGQ�����8>/DRf��i?�Q96BI�}dD�ȓ5`�b$,/��(�gΦ̈����2�ɵ}b�m�t�]�ږ�ȓ/N4�1  &d I�b��*�^)�ȓWr���.^V��qn�o&���>��D�D���m@��rFQ"J�E{b�'��(!��5�`��h�vW�+	���y�#�$ke��2fϴ�h2� �yr�kڽ�g䈰Z^N�p��Y��y��?���PÃ�;DB���UC3�y�A�-
Y��@��G�7�z������y(Ɨ����(>!%����$ 7�yR�++�l�eIJ;��Tꖥ�y"ko��L�bǝ�~{���ǘ%��?��Y�����"Cv1l�R'L�6���y��xRA��g0*�
�蔫j��=�3'T�y�Ͼ+��Y���=e�đ3L��y85f x��8M4Qg�?�yr%����5��Z�J�\���a���y�ܥ.�h��\�?�Ȥ�3
����2�S�Oa
���wL6��ʏ?W�ey�'!��#G��8����bo�����^'�!�䜯s#Ni�&!�33m\L�� H�Q!��2�^]a@+G�vg8U��ϛ��!�d@>G�Dy�pNZ�(���� �!�_9^��	��!-6��	Г�K	u*!�ѻ~�����S:�TT��b�<d���)�'p�Jq	��2*���#�
څ��'Y���*�f�� @�/I���(x�'��Yh�JU�P�F����D<$ƚ,��'B��x��	�77z��d��'\=��� :rqi]%[������\�*�1"O����Wf��R��*{�6��0"OBЈ���mi�ep! +t�3�"O�%̔j�*�3�E�����y��'(�$V�$l38oe$vGm2�M����t�T�<�޸"#f=]~y���"D�$�Mǯ=�(�e�3W��aV�-D������$� R��F�lgz����=D���E�1_bX�aF��t��88t�:D��@FY�s�$ՠ�m�O�a -D�,*�.I) �2��⁚,Ĺ3C�&��'��|��O^�� h��1(`�4�:�ZQ�"O���aH�	����؂Ԭ���"ON0q���P��y�-���Y��"O�X�մUm�샱+Z
5�"O6\�⢄�UuJU����$=*�"OT�k7O�j�����R�e ��3�'���ܓ0@@��
yę�!]$��O��$;�g?16�"*j�L*�[�i'��xA�q�<ဤ�-^
�K�Jн}����k�<i��(oC��)qG�=\O|�R��c�<Vi͜4��P�=Aѐ�J�nCi�<�A�ܲH��@U���h�
ezu�i�<��O�F}�@"��z�*Q}�<�E��g���d�M
�#�x��0=�S�В����a>x`�8���Yy��'O`q%���\h���(���
�'��P��' Rh��.Cd*�
�'B�[g10 �<#���6�RE��'=�AHK�K�J�
P�^!11BX�'�Z�{�@	�e5�t�G�U�0Qԑ�����C(s��	
�Ś/��j���0]��'��{�L�E6�a�RK�a��يp�ܱ)�!�D́!(Zɒ��v��4y�CR
17!��{���I�$�x�������:y	!�Rf���U������GJ��!�Mm2b(8�C��Y��	/;�!��֭L�x�� CՎ;3��s(�;k��}����aţԏ��a�Ǣ;��9�l�<!	�-�,��&��_�]�@S��5�ȓ[rf�����W�>�EC�#0\ꬅȓ@e�3���Zm6);��_/�Ʉ�G�*`Ӆ�ۉ<>�p��Q}�a�ȓ\$2$;q&Ǹo���� ��*̆�.��MK�_'�雳uL��:J<��@��*_a�`fA�d��$�����R�E^�f�&����͆o~���ȓ\ϖ S#h>�Z�� Aʙ5��d��\'�d�����F�����<#^d��,��8I�O�}�(����a��$�ȓl{Lh�l	�$�Z$�s-��q����*Mn�xV� |HH2W��
t��$�ȓa��դD1/������	M+8i��,2,I ��
eF��ȇ�k���ȓ?z��k�OG��V`E`B�nc��������a�ˢj��x��ʓ�2��-�ȓUV�!L�bd	�#� T��<���p�� ��@���CA.�Q��0�ȓP����fYA��i#��C�=z��#@*�ك�($���"V��7O���ȓ5�`�t��*)f�� h��7>�E�ȓt��u2��ޠ��l�Ʉ�9�ظ��-^��3�@�_,�3�P�tN����r��P�����Y�Q-<b ����S�? .<����\��Fg�O�DH�W"O`+��Px������	�@�'�ў"~z�Ӈ!j����T/J�́�ơT���x�b��6�ĵ3Q"$P���RP �!�䁗9ᖁY�BX,%{Vл�J��t�!��G5L	B�х(�Ph�d
�p�!�+I��#R�֊�(�srdA�w!�d	,�h9�R<B��L�Κ^Z!�ĝ#��˥T�2~��J�"�8��'cў�>e��خ3=Z�:�aO�%�	)�-4�O���u<4]��*�) xԀ���u� ��0?�!�
�9�|0�bI�`�	���F�<��Q�b�U����+G(�H�$]y�<���\�k�Y3я�$s��T�W�Ms�<y���oЪ���H�f�Pq0n�<���s��JA�m9jh��"O�	��
k?��A���?VN��	����L +�R��F
Z�9]vi%��N�!�D[�X��	�,��sB4#�J;�!��,V2$���;�i�o!�@J.�d���1`� �  	�W^!��ބJ�(�����=_t�U��({>��P��(� �K�㗡,{@�9S�H�>���V��0�IŖ	�6I�BXV3�!�����q�\�ȓ�X+#ʓ�b֢Y���lɜ��'�a~�dL- Ȃ:���&�jpZ��H��y��_�Y��C�"��^l��B��y�IN��,�2�,ܜ�q�[��y���1|Yk�/]1u�2-�  X;�yR(Q(Pb��B�� Y��C����d(�S�O^��Q ������!#�hȀ
�'�Y�Ŏ����IGa�#X�}��'�R ��H�@��逖S���
�'�6)1�##<|~pL��G=��
�'c��H�йbq�<zSC�56���b�'��p%�]���x�U�+���	�r�|�ᓯaaF��e�Y:_����m\�a���0�Trg��0ڥ�[�O*��R�3D��'�ִ��+D�ĆA~��&i-D�|1�⒇U��H��ĒQ���"�(D�|�0��F��m�B+A�C�P���'D�>��ᗯ�6��M�%��(n�C�I�w�F1Z2F�֘(�(0gU�C�3�N`�#_̀�1v�H"58�$!�S�O'�k��>0h)�%�������"O����(P�(���j�%�q&��'"O���W"~Ђ��Dͷ(���W"O�I�w$���x�@���Ӹ>L�B䉷q�XT�e�P8_��YSf��Mq�B䉠�^����� d��Y�@پ"��B��3C*p���	|�W'0��q�ȓB��H�%$l�" ��A�M��=
��+��}NRi�ec��E�(�ȓ ���ŭpNf�*�%� ���ȓ-(�����}�tjW���mB��V/NE�D'��<� 5����mfj݄ȓ��1�j�7�̼��f_�>�tфȓJ�����L\�԰��MTy��-�<8���&�z�2C(��N^r��ȓ}��03a�ƣi��g�ߏu����IR5+F��c�d9R���dI�ȓ	�p�D�*
,�b� 0�(I��hN,	v��'(⠻kU�0�ȓF�4�6���Na�c�� �X��S�? �ف�m�%9X��� M���(��1"O��,L��8LIfK0�X�3�"O,�¥N�)T��� �M�v�BA�d"O$lS�e�����|Nލ"4"O��[�e�(ڑ��V�B�M*E"O��A����d�>�x%I>=:v�S"Oa��C��i���'m̽,@u�B"O`p��KN�BP�����D�W"O�zbL� �3�cT�=��"O��[&��D����R�ܮ*y���5"O|Q�jJ"��̩�@���a�"On�! �Z�	�V]��a�g���"OT4��	Ļ���f!ύJ�"��'"O��4(�2����v�V2m��Q"O
�F�6�|�1�0'��uC&"O���ĢG�B�ؕ0�bAd�q"O|m`P	�?m�����	�$Ez�QT"OB���-"�xvg��B����"O���BX� ��=a�E�7l�H �"O��k!���vOx�b�������4"Of��"��TL:P�N,?����"Oi�t�"d�s��.85�@h"O0��(�&0�hƺ,$ �f"O�YYS�L�fWv$����6��"O xCc��ix��p&�"��h�"O����Gږo"�K��F�"��S"O��d4M4�cg��m����`"Of�+��M�i�3/έ%�0L[@"O���ѡ��wR|T�@B�����"O^���N	Bx�aO����"O�D�C�ش!Ӟܨ0�B�\p67�!D��"�'8E���q΅�z��\s�c?D�0Rg�=x}��h��а1��"0��C�I�<$|H*��A2�0�A����C�ɺm]����')�ղV@0}&�B䉫K^�<b�L��X�#Mq�B�I?DA)p��(?��4��sg�B�I-]�"%qrOZ�H!�U��$L?C��B䉽{�p�T]?Yc��@�Șf{�B�p�N���[�G3N�y1�E6)�B�	oE�РgoS=�ꄸçY~��B䉭i� m�FM7X�%�%L]2��C�I5�y#tՋ�)�V� C��B�	
<v��E-A�t�Q�� !j[�B�ɗ%� y��V�DeI�.����"O�-�T���\T��)�&G�tL@�"Ox�z�v p�P���);�֔H�"O�=k�-M��|!��*-P��]�e"O
�ЄEM���Q!�GR�4m��"OD ��V�,��Y�O�� �TY"OQ 򤕾[ d�Bo��R(�P"O���aj��-��24��Q�.H�T"O�e�$aI�*
1�F��"B�ŋ1"O䅺7��s�`K��T�[B��#"O��3�F�=	��ԉ�'ے�"O�<��S��v�z��*M�� ��"O��ar�B0'q�h�����(���"O
i8E�I$S��	��g�"N��)�"O8�s�E<K���3�H�(:L��"O>�S��Հ8j�Q�01�M�u"ODh�TXȅ�vc�%*�9a"O�h%1D5(娃�1)hx��"Oh �3�/z�p-��y8ڔ`�"O�Y�B�d[�lq�e_�$��
�"O� :�ȧI�<m*]�5�76{v��"O�-��d�81Q띃l�lYBR"O���`B9Z6�-C����cq�I�"O�djuE
�<%&�9�(�Kh�V"OL�ғ���urRx(�b�\���
�"O��ce	ʰ�p�@C��`&"Ox!2�Z�$1 ݑrG�$%��{R"O�[���&wmV��vɴ��UG"O�tzac��{A��.9b���4"O�`P��3�|$;b�� h:��f"O�=�7)�d�������c �U	�"O�!�1,ʬ�J9K�i͟/�~�`"O)��o׎���(w�b�B�"O<I!rCHd�Ix�#¡l�ʨ+�"O�	ff̉;���:�m�N�+�"O����A�)��j�09��!e"O���v�W;S+�=��A�l�:4��"O�y!/8P�������\ S�"O29�焤n��t���e�(��e"Oh���M�R2%[E�^�m�:�G"O�<Z�kW��<�AG�mR8��"O�i�ޡ`��u1!�,[>Y��"OV�SRÀ�:��TPad�#=��p�"O}ۢn#>��PQD�<�콹r"O&eIf�_9rXd��"N�[vJ��"Of�!e� !NԊs��&J|*��!"O�]��Ya�e��;�t=� "Or�xb'Z�
��h
��O�`=��"OV�zŬ
�V��)���9�J4�Q"O8M���	3C�����,Ӗcl����"Opœ���;q�lɦ�S�<z��"OX�*@)P�dS��Z�L[c���Q"O.a�U�S$D�j����V5J�"O�l:�(F�� `"��I^��t"OXxr�'7MFNYb@C6B>I�p"O�<yDI�J(�)SϏ-��"O�)��	%'l��&N�4]�2H�"O�q��ݿv�x��jF�}�P�""O>1���<]�>T��)�mkԡ�"O�H`$'��0�<̓�(D	�f��"O��v�Aֺ-8�"��{�U�s"O�	ȅΝ	*�ȴbU�na���"O���A�5xPi�`�G-[=��3e"O"y�a))��8��1o'p"O��*����V�%)\�*&"O��Q
I;FF�
��Fy30-� "Ozr7&��q�X ��&J�O)�%�@"O�m�􋀺�uz��4<����"OB4�b΃�qh������$I���%"O��&��/Z��4�4Fi=�5;�"O6h��7zf�\)�/
+\+�\�"O�ڦo�V֮�x��(�ij�"Oxl����_Rt�g��s,��6"O> �@�Ǳ"���ǐ��D��G"O� P�f�|�"�F�S�:���3�"O�A����Dy
�ɴF�j�NY(�"O�ٶE��EԠkq�:o�J�q�"O���󻤈y�! d�-M(�y���#9R�4�2"��N�Zd`��қ�y/��QI�P-L��X4���y�d�!_���:b�הI:�d�_�y��\=>LK0���Bo>0��)��yr�*q�5y�2e�@���,�y2�ݲuB�0���12�H,�݆�y
� ���ӭN�����T�˝(8�c�"Oz���*B��,T�� ��|���R�"O�X@Qȗ�u�!��!�!�ĸ��"O��0/�������9u��i1"Ol9��E[�2��y����G�l�"OL��T�!Ȩ�����b�<��b"Oб!aG�u0��,�G�lyyg"O�C2�Ӯ7Da�aƍ�p���qT"OV��Uf^�`��D��!S5�@s "O�$P���:(�����K�.�C�"OX� U� K���P��ޖ~C&X@"Orx�Cg\0C��������1"O�����#��Y�eD|�  �6"O҉3��>�Z�'T�F�"O�I�uf�N=� �S%c� ���"O4ԋ%������Dm�F�d	A"O�0Q�#D�S��O2ޘ�"O�zf��zΖt���̙a�eR�"Oڵ8�K��Y��+��|�P&"O�X�6e�"V���P$�`���"O0�3�"A�D���ߥXr��!"O��x�?c�ҍ��lSLT|��V"OڭRa-�&28�� @J�:�"O��@�	Nd�h9�jN"d5sS"O����	Գ!Iu2����|b�"ON�H�WW�i�)�S����"O���᪟�X�����)�
ў "O0=����bB� �犰9��6"OZ-:U牻7[�I:�� �z���7"ONX�D�Q�Z�V��+V9ʘ�W"Ovi��_�?.
m �%S�=&rI	"Ox�rp�2/��S�n�!
�x� "O�0"�N��di���/�#�	�c"O�"��;P��M�c�G)7�6iP�"O���د}�xq	F�ˋ9�F��"O����I�:��2�0��=R#"O�`�#- 
f=��M!����"Ol@���7y���O�$��{�"Opٵ�Z�jW*�i���tR!t"O0Ш�n�4�D���P�X&"OB\ �$H�O���X%̹SM�Lж"O��8�N�1~�mIE��,TVPU!"O�A�R/��'*"h�\Ｙ��"Oz���E�I�V {����n���G"O�4!�!�5�����S�N<�0"O�����ZT�V�h�+	,���&"O� 
��,f��d�'	��l��d!'"O�X1�(Ω�b����ȔQ�
�`�"O��W#�2�pU����| p�"O@i�s�̭��(��,�{���K�"O
�tLӧ\x�
���l~p��b"O��б�N[���1��|ڮxA#"O���[���� ��b}S"O�7
Mm�
�8�Ėv�
��"O�@ �nۀD����䂾}��	r""OjM�� �(k�m��b�!�ȸSw"OH�q���3\n�����i��t;`"O0��u�	�Vj�K�J�1g�NiB�"Ov镫��B����#
�˴H��"O@)�F.C�S�a��(��(�9J�"O�P`�-ôg��=Iw� �p��"O���v(��o���!�gE
n��Y`�"O(��a��.��� �?�D5r4"OBIP�,͗:����k�1ɖ,X�"O� 0}�`�\�4�����i�b,�d"O8-�/� o�r8Vh�
}�lr�"O�l�:�nx�� � oh|��"O$���F7Xa��j�o٭-�2m��"O����POآ,�1Owj� �f"OhQ��nN��L�N��8c���G"O((c��	�@o�D5.&�|5r"O�}(� �:�Ф����/����"OFT�aΘ�~4��� �4��"O�8Jᩖ1'ƺ�b!d�8$�r@�$"O*\{��	�,�0�$�s�T�4"OA!d������ �N�$Nā�"O2l2���1T�(�z�Hˠ59؝��"Od�����R(��Ң�Ԅ4��"�"O܈bC�<d,��;@�W��D`�"O>4�Cյ5qt��2�#Ḍ`T"O�|x�C�����SaN4��@X"O|쩡*X�m#�DSrG�F˞9�$"OB�)���Y"���G�N� �H�"O��* B��TR�p%T�t89
�'��=ѶR�a[�i0E��:Q��'
����i*k4��5iSa[�'JY��.�-zRe���ۧ
��M�
�'���COF
萨Ğ|�\Ղ
�'ML�3�����닑zs���	�'�8L��h^�{D�(����c����'��i��&	�	�4��,�����'~��A��B���H�ǋ:%O0�P�'i�5ʔ�&w�Pʵ/J�1��(�'�`�ٕ	�!Հ5�q�Q�]����'G6���/0�HB���j@���'�$0
fK��+��1�ώil|��'�by�C�L�{�A�0
[�p�-s�'Y�%���^,l�{M=�$U��' �Z⌉ZG���q��h3.�	�'���[dc�/,!ny�!�P���A�'bT��i��D�Ht�ڧC��c�'��h;BF�q����Ӥ�;���b�'lQ���-cܰ�G".8��9	�'U2T�wJU�~�$l��`�4}�x��'t��IC�ܴ��AjZteV�1�'��\+�@	��*��_"f���'[��Cp@T�,R�,��#�"Fv`�
�'����M�++�MPդ��-c��:	�'a���4�˞�*-Ig�:7���(�'x���vղPr)����5V�x(�'��y�Ț'e���u�?%c��
�'�,��_�%��Y�t�ӹ2��	�'�V������kT����ʓs:����ک}N`x�k��E`ه� <^���jR8wv�2! [	<7�D�ȓU.pa�EeI7$�ڽdT�L�bP��L���Eć9�ބ� ���m�����9_`D[V��sw\M���pu���xT�c�H	�N(Kv�� z���
�����(2f�����u�чȓ���A��*e< �
��	
(��k��	ɢ�ˮb�րrpJ݋uF���<��"iX=1b��0�24a�������)rP���i�?dr��ȓ~��,Pe�?ٶM�ť44� ��bkP<� !@=�87.C�Po�ą�
��h��*�5��X#�Ϋ'>�ȓ���Ə�?"�F@�ZY�tĄ�S�? -���
�/7��3 V>����"OF Z���?6�ZQR@��챰`"O�}[�\�,��� ��/�\�t"O�(�Ad�f6h�vnV=��=��"OR����l^6	��HA�>��3"O���G:s�I��L�r�:�aT"O���W�4��Xb�؁J�
�p�"OdL�`��QU�Xi�
GS�6A�t"O~�h�O6��-%�Zr���k�"Ou�aL"<�`+Y����t�<a�䆠W@�8�\�%�ꨪf�Y~�<��偮Q��� ��"F�ݒ0�Tt�<����,D�`�¢ÛZj��
�!e�<1gNN�D2J1��.��$;Q*��u�<av _� �n�Pr�Z�_��=J�M�|�<��B\�&��ѓ2�(K�b�� �u�<1��Y����'P&q��!H�n�<�����^(�Eͪ�=)'��g�<��Ӻn���P���� ���hY�<� ��#J�|@���'Zs8,�r
T{�<Y��C�6�*�GeD'.=hC�}�<I�FY6)������.�@�(��SO�<�w@�>�%��c�]�5`���I�<!A	M�b��V	3���i�E�<��@�U)���KѠ�&h�rf@�<����8�:0��*��I��]*�(L~�<���<$­)*w�dP��.JV�<��oI�d*��r���|B�KL�<�"ń"I��B"	E�[Bڌ�vf�`�<�w�0B+����~Ŕ"���G�<i��۰o���
@D�b6�x��GB�<A�IV,Ă�9E��O7��{��\A�<���?<�i��/�s���҇�A�<�$��.@'�-�P��R�,P���RR�<a�f��<�|�%�W�#� !��W�<Q��ǝ�H��D�7e*�WbBP�<1�G˒j��A��*�|�"|Z���c�<�7�!]�r�N�R�8�а��J�<	�"p�v�(�L�m<kD�SE�<aFFv�~!�6��I�V����
C�<��	G e��ip�CZ�T���CT�B�<�q��\G>hs�#Z/˚�@TB�<�1��MҨdif�ݪ<��hv�D�<��4oށ���Q&n{�@X��z�<� c�f�� � �H#0j�:D�w�<ᠲ�,X��̀9�L���G�0�>B�O�q0!��:X�0f���[��C��>�pn��9�$��V�2B�\��ȓw���QÛ�K:J�1É0;�~��ȓl(p�j�,�\Lm�ċ�-]^��ȓa�����@�H��m�`��\J<|�ȓ#�n�J%H�?��Y(�〣.�~-�ȓ4E��� 8N�jHH�a��P�ȓ*���{B�,�"�B �̅@���?X����ʦN��<�$�M�@��}�ȓ8^
�҇*\�W��H��} �x��=b�%��{ւx8t%�aUv��ȓF�Xd��G$=*|�C�
�at*��ȓ2b���֦ɱ8q���d�doL��=z\=J"
�@~rB�Ńub�ȓ��bE�Q+v\����=-�L���Z����!����� �3}�Ȇ�q�Tk@hǛg�H19�!ٷ+��l��A��y"�U08����#��0O�6��S�? ]��E�k�6A�aȦc"dl�d"OBL�ȭK�����M �3�"OґZ���-����������"O 4�u+$&��dESv�� "O����|j���������u"O�S���&�(@�$v���0U"O|��C���^]"U ��D<-�@e�v"Obt����"�6bv��G�ʥ`"O�0��MÝJ��rI��l����"Od��B��lb��nD,�z��"O����LD)%�h�b�ڂ8�&��"O��e��L	�Q汲�!bCi�<�3F�)e��!���-"؎\�0$d�<���&]w\��4��l�e���b�<q��_:��h4�T�o�j)"��W�<�u�V>+����'�;gX�y௓R�<ѳNA�Z��U���Ĝ	6Th�G�<�a��1{j��GK�-?l���BCA�<����eҙ�I�\jl �z�<���َj�4��C,\ Zk��#��s�<ivA�W���10酸"�|D�U�<�T��8�2�閇¶]���m�S�<y�h;F�xPe	zEh= рZ�<a�Y�uZ�]��S��
w�V�<Q0"�,T��1c��
uM��F�Q�<��	C4��hq���H�,��F)XP�<!F�K�:$4�l�>%(̐*&��F�<�Q >~H�f��=P��0�6\D�<q��§v����6�l�Yfa��<�V�J�p��-���O6u����|�<�v���Y�d%�H��l��D�<)'�T:��iʮK�
��E���<��J[7UԲyq�k^+r��EVF�<9��O�g� :Ц�U�|��D�E�<�kL�S�ΐ�s�Qq�z�puj�D�<�v ��1!d=����/�����Ng�<���[����35 =��'A}�<I��{�(��ԫI�E5`���Hz�<��K�5(B�+�nրg�ʄiY@�<�"�X&ƹ�H=Jz�s��z�<QT	S�3��-�膺H눤q��^�<i�� $꼙p�6n�^�8u��Y�<�«Ќ_�
�%�[�b�����'�S�<��R�f�t��e-_��\���Q�<9���!�������'T�峁GJT�<i�H��PD��ʔ�]�\'X	K�L@Z�<%�̗bF5 ���>Ax f�U�<i��?�T��Qs<R�s@��F�<��l9^%���I�	��+0L�Z�<�� Ŭ@e4��c���v�Ƅ���[�<��Y�v8B�a0�Y:d$Fh#��ZW�<y���[`��868[��z�<i�,��f��K'n1^'�	a��r�<���?�hK'�E) 7R��a͒q�<�S�եN��-�%G���D��m�<����@]�Y��HP"	��L���]c�<��ᄢd�>4��i��^L���d�<aqd޹ފQG�ٖ
��8c�a�<���<5�j�b��a;4�b �\�<��̎wD�!���l	0�"�T�<�q�B�*��1�
79�V�� �Q�<����O�L��@JPL��ip'Es�<q�j��`^51�ғk�ܥ�Qm�<��+I��Л���'4���Oo�<� >���EO�%��"��M� xӴ"OT�a�2'XRܻ�U�K�p@�"O�-��N�6���#Юވ9���"O.�*��3�JT Q��T���q5"OH!@āهR�`�S��ҫ=��1��"Ov�b�Z�z.���
�)d�$��d"O��8a-צ��a��:o�Z�K�"OB0K�ID�LؠT��A�*V���C�"O9��ܞB��+�oʸa��Q;B"O� �fŅ#�b�2 X�.���sE"O�9�	65�\T�ծ�9�(���"O��]%$�Du�S��?j�!�"O�E��%�yQ\�Ó���]��"O��Y��[�,���*ROY�b�LɈ"O� �D�ŉR�JP��8Al���&"On����]Zj���	d���C"OJ%���� �LI6��hU�"O��#��ܧ{���\�dl��q"O�P�aN�B;FD����*"THr�"O�mk���|�Ɛ��L�Q�jX��"O�i #(�c�.��ލ?����q"O���5*�]?�ءf��4�(a"O�A�#i$h2Bd��	�^ʄ@ "Ov����{�X��Ƅ�=RT�``�"O.`�G�L��x��7Ê�FCd`J#"Ot��� �*,����=0ZE"O1@5a�[��*�B�<N5���"O�P�B�\-�ԡ)c�K+.@h�"O΍rW�V��܉���9
.�qf"O�0c� 'W_<�� ��nx ��"O�\���ب��A���ȋmn&IP"O "*E�0"�*cG:��0�d"OV�p��H�Rq��ˀ��� ��"O�|24�4�fXxvf� N����"O�1͏�X�v�r7���jXqb"O�⇣�/x����AѤ/�Ti�"OX\�g�!����!�Bf@�7"O`�x�eO�&���P�L�qd�}8�"O��Ad(Α8paawl�#af��D"OhY[��<R���a�vI0�""O<\�����d�q�� =�`�"O�Un!B=q�N�	`4:eb�"O2B��>�@����$||!�"O���Si�J~H�iǌř[��z�"O�]3%��$Gu �1ׄG�O�WLw�<�Wh\E�~]i5�͒P�~#�Up�<A��_0jJĳ�M��ZsX�
b��h�<�*Ψ,>4�b�l5�j�
���i�<9���:�J�3$�V�%A(����O�<��'/jZ�Y�F	LH>���E�<����W��E���'����_l�<)*ܲ-?�}�ь l��AH��RS�<A�4��%(B�йf�lQS�nR�<�Ռ
�-&�y����}iz #�	�c�<ae��zܨp������@���B�	�L�6��q�,`��2C�
 ��C��b�4qsT!ɤQ�ĝ���H� �B��8o��)i��;b7LP ���Jp�B�I�+-(T��U�TXJ���.:C��|�`p��_%�lQp�^�-�C�Ibq�ʅ���2�&8��HY�1��B�. FY�#�D��0��0��B�ɑ`,��ᴀ�C��M��3OĘB�ɞ=��\���?K��c��E�n�lB�)� Θ�SE�bj`��cQ�&�ta�"O���k�4����� >�Qf"O
=�Cmʠ}J����λm[<��"O
x{��2�@�i��P7W�x��"OFԳU�Q!_��`�8/&|��"O$qɗ%��(Yc �!� ��"O����՞H�4@�+I�.�m��"Oj92���r�x%�f�+�`	�"O0ly�+F8e(f( 6d��	Fi�"O�!��%�1�íqc`2"O�����ÔD��=Us��x�"O�}H�E�N,��"EA�B��A"O��!��y�8|۠ꇄt]par"O��)�`Q/*[�a���h=6<�r"O`	�f'R0x�\��	�,Q3��a�"O�X�fF�e)(}�R(�
'�m
$"OD��դ�)��JR��`��ZD"Od��AM�JxF��E���p$��"ODL��cê7����a�X�����"O���#�_
=+��A�an�;1"O�Ȫ5kP �Q���$4��Ip"O,$�
��e� \����D�6�j "O�+�+u���4F�l᠜��"O���M59D�)��X7�=["O"@�V��9�	�1�T�`�D�ؐ"Ob�I����B(�E�0�L��'"ODhH��B�x]��`�?���7"O�1:���-w\Z2��
S��%+�"O�8{�E%(���.On�D��"O2i	��P=��(�J�;}8��"O<����6aB4Bi�,t���"O���Ќ;�.���!�H_��2"O:�k�˴�4l�p �cJf�"OTx(�!�����^0iv�(�"OJu�$iM����KH>#B��I�c)D����C�F��)��D}��U�:D����CtmxP�Q��m���N7D�\��&үM�Qҷ��;����)6D���uˀ��!����L���U@3D�XX�E)�X�r����G����>D�,��ʀ	%*1Q���
l!�!1D�гÏS������-LZR�A��.D����Dt���A�B�\q��-D�H3�[�i�j�J�_�G�H��,D�x�U�O;Nk��Ȣ��Pt	!B>D��B�J�o�X���)~Fj�;D�\cg��)ꐌxb��)�2�{�A-D�ܳ6�@�W�X᳣���<[ju�ծ*D�|8#@�4��R�D9/��xQB;D�d8�G�3e����������m=D��c���5> �A���~���Qn<D���!�;�vi�������9��,D�d��E]��؅��1A����7D����2 ��� ��Y�"�֠:D�(A�Җ._\,���Ѝ�T@EO:D������nN9�T.M"�4I��$D�@+ph@����A�O�]1�4�q�"D�H���O�����76�6�I�";D��(5�B�(��e��h�n���8D�\�$�^32J�c�mY3H=�M���5D�`j��M ����S�2��u҆�/T�H
e-]�|c�u��N���<��"O��#��״hƪL�+�,Jʸ̈C"O^���;�Ztj�(
B��(�"O� �`P���i�4I%!��^����"OI�R��)|K�Ǝ�2C�Ȁ9�"O�P�6b\�tT�=���K�'��E��"O���N϶�C ����8���D:LOL�'�)UG&L��@�jĄ��"O88�U�D%h&n�(�jL-
��@r�$4��0*�Q��ɇ���Eo��gF�>I���.��'"٪����k�$�"I�Ce����'��x�����؅�A��7A���K<ѪO���DG�4(��S�V	+!�Y7&ւ	x!��7Uf� ���7�l��b�?#q����F�(d��E��b��������e�tM���qܓ���Y�Aִ|x@ ݪ%<�	�'�h�����("`�	b�0��r�)�$m@��|S��F>~@5�2&��yrF]�u����%\�y�VT �hW �hO\��$͂P�TBFB�:��5�2F�3|!��G�*X��#� >�J��w$��
 !�$��ԥR��8,H�*A�2�!�D��7�N8#�L^-c��Ӈ�T?!�$CB����q�M�2F��g	6	:!�$�$`y�s�S 3r��GG�<�!��ӻi���"�m�y�&[���D1�S�O~@�P5댄Z��8�ck�cx��'��,pr�	�(��ux�'j��܀�'�
�S���5W�2p@���Ԙ@�'��a��(Y�:���Ay)���"O�}0$l�(Z&���m�7[�X�t�|��)�*#���a��ӌp2�U��%& �B��w���$�Z��A��(d��6mU�Ity�	?�B���C@�w-<�f �!����_�"��Y/ƪFM5`נގ[�tԅ�QY��;'١?���`\#��>yU�)�I��b����ߣ0�:��B�K;!�������M�~N %YW��n�ў�'��а�����.�!��&kh�0�:D��%�μ���+"�Z�<�V �S�7D��+�g/zQ3$ŋ2e�;q&5D� `�C�B�2X*�e� vA���/5?��d�|�b�{��$񆅗
@�\��t%�x�`VI%��ht�[��P���|���acB�o������������As𤟓wb,�X����}e��ȓ|����� �&f���g�11���ȓi�z�ae��9���@��;;X�e�ȓ>�Vܲ��6TD�cwOT4e�D �'Ya~�jW%0�`����&l߈����0��>	�OJ���;!��eIcJڍn����"O���We�09���@��ӷ3����&"Oj(�h�>�D�U8m�J�e"O�%Y���#V�$9֨ <��ر@5O��=�~��'Ð���mǇ40`=i�%{-���	�'��
gJ�2m���'��= � �y�V��G{�OO4u�s�̮/f��p�DB�<^D�

���> ) �@'8]S�i
��'T���$��5^�ޑkq��.p�x�3��vL�O�O�#~R�4�$x��Y�a|����]|y��'�8�@��-Ƞ, B��U�Ɏ�D�r�'Tt�'3�\���n�r����$�-K��-�ȓV�R�����Wm�qE��|�taie*�j�	c������[�u�����	Υu��[��%lO��pP�mڣBB�pj�� �Zs�ՙ�"D��z�ʏ�N�H��6� �~���9��!D����3E��!��*Uġ�"�3D�� �y����5ҊAsU��
7����'=ўD�"܂�6(�w��zͤ݊��*D�����I�����aD1?x���<ʓ�hO�ӓ<��EmH<6��lc���$�����%?�N� M��`�%Z�	#n���nH���'wqO?7M��;�d����'�����9lў����'�L��X::����`Ah�M��}�%��}�!A��[3����NÛ�HOT��sI0ƫ����;a�S�h�c�'0�xb�B���ԌQE���'6b%�ǧ����{��Z�xC�z	�'Ĕe�2Ɛ&1Z�su���p�2̨�'��]i$�j~��!U��>V��p���9�S��oͿl#����C���@�]��y�Ŋ:h�aG%��+F��`-J�M���s��9Ӫ��y��0��� ?�`,:6"On�hB��#7s���iG;�P��U�O��Dz����� P��sG�� �͡�ޤ�!򄝎8 Xע�X\H ��_k�Q��SH>��Wj�Zɔ@	���􁆃$L!�D�����cf��V�XР��K�T1!��$�~4�'B>_�,�{u�Qt,!�߶$pb4�`@�#�8��H�"�!�$C"�)�5�^8'��Y`�5|!򄕂��4�%}N^5kS�L�L��C�	�y��3���7z�=�Х�J�C�I�
� q0�
f̎M�W�օkhRC�ɢR�N�s�U�W��p*�ȑ-L>C䉜��١s��\T�)Ad�3Y�C�r`�a��׀db�[��Ƌ2�RC�I75`�p��o�^8"*X�f���>Y�b
%tE�����.B���K0N �<	���Ӄ6E�u���8d:u�3C6J�҅E{��9O*L	SFE�4�t�g�~U4�R��4��I�P�(�=� �'�H�lj6-'���!��x_mLn��9��9D�| U�X�	��Y0(I�I�٠`f1Oj�=)F@7��!�d��M�����^}b�'!�� �'	G�ΌQ"%!Kj 	�O��=E��dH��zā.�"�L��$϶�y�m��B" D��ՑkTX�����0>��Q+0�,|au�[�Cg�ģ����p>�H<�wbM,��!Q�O���v��<1���O��I�B�<!(�(N:m9���B�5D���� 
�H���e(0J�\E���5D�8��4��)����S>�P'-?$�܀��W�Sw��G��
K������y��_)���Ra���J*�1x�hF1�yr���3͌��**l��i�'j4D�k复�Q��x���%lXp	a��1�@+ؠ��3����f��� 2ͅ2j���j'k Z�!�&{9$@��O��m� e�a!ڤlS��<�
ߓ?�e�%�.����!�)������|Q��*��4ȠBA)
����ȓ*f� ��IIQ~�c���<����=a��'�*�Y��)i�!��ѭB�^Q{�'���'�jH�lx ��^`j-)Q$�L�<���b��A;ێ�8`d�<Aӏ�� ��d��ί�^t %i�Y�<��G43���P�XO2fUHQ�[k�<A��~4B���� ;8�fx��O@�<y��֨g0Q�VN�34�.�� a�<Yr,ٯ2! �h�`��,4�M�b�Y�<rL�Z�F-f)��!i�y����<� ��3��vHxJ�K�'Kt�q"O��3@"�5:K�(hce��f��"O
�A��K=Ap����)�p@��"Of��d�;�P\��v�h�"O�m�'�8S����D�|�b0�"O�l���E�@���C5~�v��"O�ui����q����H�=^��E�"O���fkXA���Ӱ�,g��&"O�����B/Q���@@L�L<|��"O��(�e��7g$и�/ʿ۠�I�"OhD��-�P������J b��{�"O<���#�Z$G���m����"O\,)���R��#��ςC����'"OR��gIF:@����F�&' ��"O���"l�;y�T��F��#Z�b�"O0�!p�]�]X�g�8�D�"O����3P�@��S
2���Q"O*I�U�є�B=�'� &|A "ON��`��O&A ��?�����"O�P��	��,i  [;l�"O*����8����CQ�}��qa"Oܕ[��d��8C�&dv��:�"O��a@)��2UnH��Bе;v�e�v"Oj�y���1����7)C�� �"O�����&h��!v�J6F���1"O8���ē���-x���&3A��� "O�y��d��E���GI�z�v��p"O�D�T��:�.0��h�,^~2T[s"O�y�Ɖ�b�֤�e�-^�k�"O�[����dj!	�.S�� "Ob遗���i��``�H�v��x!�"O{s/ٙ��Ɂhɯi�X���"O2y���
}�603�h��	�`�e"O��
��̮Q?�8s'Æ4�`(�"OH�6�Y�X�6�1�*�
囲"OȘ
W*+����V<r�v�Zv"O<`:��Z�Z��Y��$�2ɾ��"O т�B݊$�@I�FԸ#�V�9"O*�5�.r��x������"O4�(��;P/D��%�T�R�F���'O$� �^(0��.P�s �H�'�l=1��[�F���ꍣb/��C�'��M�d/>Cr�I�Q��6R�i��'��M�򇋺6#X��1	U�S�h`0�'Fֹq�I<\H	p��M�|
�'���@7���Q�(�ehI�D��͈	�'�8�k�p��A��a�)4v����'^8�)K��
U��' x1�'غ��f��O������Z�haj�'�*hqkY����'�a�t�[�'��XCD��	d0��1K�3A]�Ņȓ!X����I$NL<��N�0���R�TE�!��[4��Vm\?[f:Y�ȓ�$Brl�D`|�1��֭ ��ȓ_op��`�Z�?���sM�B~X�ȓ3���+'��@���!I!G�v݅�Pdz]�EąI�6HpK
e>���6�� j���9X:x ���]�8�ɇ�Q�Azwe\8V�P���r�<l�ȓ7����FcAb�{ �Q�	�jq��%$��"�?V��K�o��#Ct�ȓy�������w2���ү5�����m+�钋 X��p����l�t�<��&�]���0��Iwpj���. s�<� N��3�  �M�g�.ȫ�"Ox���DĔ{��(��=�@X�Oz����0H���q����,�H]�!&��+xL��'�PZ���8�Đ���Q/m��Z��D�>H3�|3c�/�)i�x��'�Y�a8�HB�(��VC�IJ�:�6��>r�v)(��[� #8�y����ƫ��N�PӧH���B& �3cG���4����6"O��吰T�օ2˅�W�� (b!}B�
A�Pu0�$���M.-��25-�!2�"�:eHZ�`a2B�YV"��r�!7`��#��: X�p�Q"�-�F��I�C���b�́�&pȒ#�>w��#?�'̔�i���6��X�4C�Q
kӂRp��C��ўp�!�D��:�{!��1lh18�`�Q��I�+��\�5�I�"}
�ʕ�i�P����2���KVn�<��eD�r^NtiCJԎ*��,��/̤��	�S	�Gޙ��g�~� �U�7�U�w(µk*l��	�L�(4j�Z	-��a�wn��+���Oؤ����'����5S1z=ʉ�����F)��WN����/�SW����/.W��P�aB�#M"C�&]"�A��-莜
�n��(���nY�)5�=�)�'&�v�C��ԕz���uG(-�5�ȓx�J��QKG�p��t�pDA+q4�\��#��`�2�>A�q��!)����/�uA�KHJ��y�E��Re��"�"�����n����eNNF��`���������	A#P�h����}�B����D�,y�IЋ
q��U�r�r��޷;F>���B 	����ȓA���uE��X�H����Zq�.��ȓR����s��v�.����S����R��ѓ�Ⴃ<#h�傀 �B�FɆ7H,Bቆ-�4d֎~�dx�ȍ�5�v�?�[>�1J��4�
�]�N8�Cf��V�h�bR+�y"$��0Θ$V5K����C+����"��E����y�ff΍D�Ԯ�"E>T3!lR�H���C˦�y�-��f��s�I�Qx z�띶&ܛ��\�Vu�9QJCE%f�㖔�4���s� $���J�|N�:t�Pu<U��	'�q(pǊ�m*����S����	?{���F�ҪN�>��kK�R�����H<Z��'�<uZ`�Y�h��E~bB3*і��	S
��U;���l!T	�L��=as�]�wp����0A����i���ȋE	��sBͣ{���]� b�͟8f
�;T ��n�6Az��������$��2������Z��-C�O3�y2���
�eҮ[���2Ơ�h�a	�� _6��E��-c�l��OW��X�\����>�1,ǩ^�-��c��"�̰�Gi�_؟��c��P��h�׊�F� Yz��?F��b�ȗ}���P�ѧ����r�
ͬ��O+�V
,��p��f���Qz�+[�'�ָ���
-��d��&���M:3k�x4~��� V0��toC�g���Ңӕ5ۼB%3�O�X֩�"^jb�`%����E��g�<�W �d9p!��KX� )��[`p�Pu ����w;dU+`�ٌe��i��`@>Jl���'������	AJLpB4�w&zl��-�(Oy6�@4��%C�\Y'�ǖ��$A�&!45
`7��6�)K��k���h�,���է%���yZ��Q��R�i���G�ig����NH�4�i
���=�$A�6fY�_�ȃ�C��6F�a��I��u�旺#�*�8g��Q�	%I����gO�+��H�D��	E��'V0��IF�9�,��IV�W��i�K�f��!�2M�h� �I�?$Tqt���>k���f��5z�P��cF��æ�=l�ay2���+�@ F皮k�D���s�q�ҋ��cq�7M*��MBWN��[|�X���7^ܼ�RH�?y������IR|v���SJ�+o�����5�D��$�h8蠳�Jκ�$�DjC�\A���'|��@`D�M�O�aU�]�|*��
�#}��� N�2��T�Q#E�XU ���8�j��'R�@� M2�=&�
7?�`�g$~�n��&��*߬xo�Qଠ��]�]�-a5b��"�ᰅ	L����M<�G�P�3��-`PH�6x�,�!э�qy� � t����E4_���	ĪLp�&ϗ$8"��R6M#W�A�s��,��˅�̍2���P*�8����]�Z��S<,O6��e��p�H�1�_���`Z�%R�hVL\(�t�B����KŮx�MK
�T�*@C����j#)�?)��ѩ
�8���Ӏa��9pJ��p?A�dO!BwJ]	wMүp�jq�ԍ�M�I�g��r� ��Kپ\�Լi_�ڪ�ly�̟���b� V�htB
50���fګ$�Z 9��I	+v��tck��tb)��es4`M}SX�:���Y�D"1OԈ�GE��Snb�.�� �	̾(/V�b�|�/H�r���	�t�&��1i�����¤j����JF�,��?�lZ0��:שפO��@��-K;p���kp�_<�x�,��	2�!LO�m��� ˒��e�@�c�D��%�;����a�N��ț�T(���O,� ��K@���C�i�t���'Hi�֌ÎmZ�E�7	�$H��
�dG�i�<���D9�dᆚ6��5e4f�8��b����`��p k�g7.mꩇ�c�P�8�!U�Y���B%�.4<rD��v��%�"Q�RW�	��'"$���g|b@ Pބ0H��j@�V�l��T\�9p'��Թ	Ü ����ȓ}W�0��iFx���!
f�����y��8J�@�>Ulyk�kڃ4�����r�`lK�L�Xf��D�&�!�'��D�@$�s2Y�.K*:H\���'��2u�ә ����l��:�����'�"�0��	-qV"Yp�Ό�7t쌃�'��%��Y4l4"%����,Yz�']�8s�^� .�������!	�'�%Z�%��	m$	S�ɀ+�����'1	��ŕEE���Oݒ�m�'M��Z�'~ݠ���bL�	�'�đ�7�ݾ7]�A�oʗH�R 	�'���c�QP�T'[F��ƁG�<)���)-xSxً���h�<�2�){+���#�8r��;bBNgܓTP�!�3���WɅ.߶��T�9$��la5"OF��� � T�D��w���4��9"���B�O�1��3?Q��* ���ge]�+8:%R��_h<Y�aX�!��Ҁ�104��`��	,7��"�
ˡ����$��F���S�:��aˡc�F�y�`Ә>��I���OY}2���2ٌu{d�˘W�r�j̎�y�n�ArN�UFBYN���s ����XK��볠-�#��e�#v�^��EF�2y؈���F�<y��0�F�+@X�21p�H�d=`�����>���I$����	=t]�"j�W,��%b��У<� O�<v�}�%��*�|D*��1yy��0�LmG怂�N�&q�>���P:nh��c4n�,�pp�	���֦�Y>�O哏{֨����@�Id�IEz��'���g��|�'�_LBC�I�_qJ��RdZr�z̰��"�r����/C�9W-�Y�4���'��	���O���s�MѪ ��!�5͂�Dº�ߓY� ���Z���6�͌"�|������]����2fY����'��Y2d\>�z��p5�_�d�|�acs���?�3.Q9$���*(ҧ/`8Q%�R�ɂ�����X�b��WX��ɝ>x��χDr8]��GH(qblȡA�@(��hXL��D��'����sb� ��5z��7&��p��'���[�	_$.sJ����2	�����m��'U)�N���T5DU)��UmU�q{O_��{r���c�0��u,����˅��1�x"�d�7J�99�J6D�P�ua��;[Vy��_�%�ޙ�L5��;2t����+�0v�>=[T��S]RĻg��1M����i9D��C�S�(�V	����(��{��8%M:q�R-�p�)��<��FS� j��J���:��E�]o�<����Q0
��N�-��ar*m?�q(ذwt���DO�j;r�IQc�w\�C�Y�]�!��/N������W'����@�f}!�d	.%
-C��B�4�I��@
$Y!�$��^ظiʄe�;ځ�N��J0!��9=^�x%H�6F��Ip[77!��Q�[L�0Rd��~�zu&,^�$!��݃��!��n�%�hI��)��!�$�/��-K���7�:�R�\6]�!�� �Zdє<H�q�Ԇ\�F���"Op����W�F6|���-� �Ű�"O�!���*a���+�Ip���"OD�c)
�7�*�hADR�u!""O��9� C;yTH�a�J4(��G"O� ��NK#g�L��&M�80�b�p�"Ox����ZoǜXxT&�|��XyQ"Oĵ�w���0U�	�K�|`h"OP��v�Ò5""���D�)K|*�0�"O�0!ЂT'}�01CI)89���3"O�{�M}a��B7l?��YR"��y�!�$���@�+�c�Rt�&�S�!��U�aW��/�ddr�	&��5	!�$Ѕ{Y��a��;Npj�q��,#�!�$�5| �����>{�$;'�*K�!��{���"[�0b���C���!�Dω!Z��STOI�aP��
�Â��!�D�&& ђ�̶3�x�x'!�7�!�$�%R�`t8q�$����G+`z!�d6D� ��2*C� ��ԃ�'E�Y!�ɑ����h�U��Ir�JB!�$��;��yh3*��fypQ�J
�52!�dӧG��e;���Jh�˖I�!��B�!�H�3 �͊rB��P���r�!� �
4B�K� �2DM:dA%���!��V�$����rS�-Or���j��?�!�&s�����.�->��Z5��(T!�$F1:tuk�H�;< ;6f�;7M!�ѱt�N�u�K�q�Q��O��,!�$G�e�21����#N� -�"x!�D[63�L��S*KW�pp쒑n!�-�\dQ�eƦP�
*
o�!�D��# >��GO�8nLX:1��Z�!�D�1�R	Bo�q��"��L�!�l3x0i�o��<�(g��9`�`C�	�sр��匯&�m��,B�nlC�I&;�xPG��5��pˡ�.	>B䉮p;D1��P<l�<⯜:��C�ɂ^�aQ�m
�dB��Ã�� �C�;]V�1A2X.��Q�Y�C�ɋ5�h�Q�	�A�\9�A_"+rC��/r�n�[#���M��xY�d��iG�C��1YD�|�0�9�I��e�C�I�-�z�(Ӡ1)�a���BlB�	?���6.��D���M̡q�C�ɬP�^��$��("Z�0�U`�-c܀C��9p�#�O�:��=%��C䉽GMNI8v�;�`���li�C�*+�A�1/�&9bX��GJ
j�bC�I
z��,s OY� �j����F(&>~C�ɾ-�� )�O7T�(���<1�B��:?m 9�U�|'��$�TG�B�G�0y@��a�ѱ�ո�hB�	�p���(�N���q���ռ0}RB�	��P0U�V44���!@g����C䉯'ax}@�A'2l�
@!�%7ߨC��b��B�Nڽ
l�� (��!U�B�Ig7�Ɉ��+zR4y��ݑ9ߊB�I!9m D�k$;=��0�ۀ`^C�I�NF���\�e�h���[�T�C�ɺ۞,�q�Ǒ�� ����]�C�ɇ�!�o�>/I��,d�EP�,D�8��@�+*�B�iV$K��w�*D���eS,�lQ���Bբ�Y��4D�� D� �� �f�.9��Τ%H:=;e"O�MS�'�#�4�sR�R�125"�"ODR��8El�@���u30��"O�(SL��HWN�벢%.��S�"O��$��JCB�sÆ�'&� �"OƄ�G�?xz�9�B��D�
�'b�����9W: �f�μ�a:�eS�}T���� ��όA(����IGJ
YD��1[�в�	V�0¦�p��?qP�y��\=4
!�D�>V�p��L6K���Oއ+�I�e�E�@��~��S�O� �x���a��`#a�[����'5�H ���ĕ-Q��h�p�>1�c�)^�n�ᢑ��}��D9O�t����[�����?��C�t��)�D�4-��Pr/�&p��2v��H!����Ǝ B( Ŧ�}����ZΑ�92��1����5��$A]\A&i��B�_���{s拄�yB�NI�%1�l�Il���
��d�d�vx��KT��)�'I�d|�X�Bn��쏐S�
��}�$��O8ZY�tJ�S�mBH������%��y�L|�>���Mk�v=��N5<ih��c�^؟t��7��ѕ�Цt�����>���")\h�RN�3p!��QP��=1� �g����O�F����b>�U�:�<���xi��!��)D��`���=g{����$!0�,�3b'?	��H@b�"|"q��y^�8�&�؅�r%�4��|�<y����?PtQ���͢|�'`�~�<���ϝ7x>i�L�@B$����z�<� �H*-���V�G�\���t�<��BD1v�<`�ñ4R�p���\�<�G�ѭ|*
��R�4U��	�c�\�<�L�Qc�}
��,m� BJ[�<�Eφ�i}�ae� ��a)rEHT�<��L�,r#�i�r/�b8,հsNU�<idh�κ�Hg'�Ut��$�TL<aD(��^O����%�:Q*܎f�@zM�B�	�g���1�+E�'�Nt���9yc�?�FT/ܖ<3��D��my>�rd�o������L�<I�c��1�n��F��Y0~`��NCO}b�7I��Բ�C�D��\���g�%Ixm���fC��7P�����+]QP��.S�\E�O&� �<X�f�&>c�d�A�
-/�,�O��EĪL//�aB$��X���T�|����7*{Z9���8':4�*�O�{O�0hRI���
�!H(tx��Iz4�9S
S$6W�Oa�\����$W�a�%�Or
��'�ʈ�@ĉ�c�v�E��-2<A��O�3�Q,*��y�I�"}&�Ж`RXU��/)����$�T�<����f�)��Ɛ�4�r��!�)��	!aoz��1C����g�zy, ��U�Rf�Ւ�W
N��ԇ�ɝ{��D8��ѝk�j9C�l�RF �q���@ɩ��'t҈���������H& �Q���䐥nvր����}�𬣌�4��>YK�`A��zJ,M觌�&�y2E�+;����̖9Y6(�чJP�eR0���m�_�h��EÂY?E��'&�+�D�9(*����w��(�']X�"��2^E�Y3�͢v�25`Х+��<���4qn���|�L��k��ӧ�R�� ^!��ǻB�D�� �D}���{�C r*�XP�b^��M#q���_������'gZ�B�-��<��ꑪhzL\["&E���4���QM)�D�9���0vC�-/.����
!I�[8ZTw��A�8X��GW���S�*�(]����i���!�i\��/??J`�V�O��`S B�t��	��B��C#N��.ő�DݤS� mո<8����i3���$�ہ.��*_ky���'�L�S�t�`��	s��b�n�+A24���) �O�m"�Mұ <y)�&B.�L0ab%�� ���'��c�� b�$�$�Ǝ0�:Cĥ�6\ ���'�`џt���7�@y�f�E��!�����:S�0L�:���R�a�)c�'G*���B�L5>m�`�	P?ͧ{BM.R�'lRD�l�[ښ�YvnQRn�Œ)Oj}Sf�غCCP�����$�M?�Z�n�0%6�� ��H����3���!B�hK#hQQ?I�'#Y:�%)�;,ODc��2I�2 [��,5U���2"�
8�4c�f飥"ǢLz�8F$��`�uP�';}��O� q�F�P)��;�1�j]�L0�O�,+d�/WW����
�:� �3V����%��Dm��!�~RF֩��i���'|��d���d�q*�F۱^������� ^�GiP�o�~ݖOݤ�����5�ԁ�
��;���H�'y<sïc�:��S_��S>t$��&�����JU��##
T t��hz�H�<y�.�Sމ3�����(�\(�"��8��pZv�~�d������x�N��01�_�3az�kL=��p��Hc\�3Ac�g��'bX�Ý�Ϙ'@n<bT�Qٚ��炒!>���
�'69��$��(��@ݺ#0Zi�'��_N�e���I)�)�Fͅ�td.��'���ȓ�y������S�="'M��C���'?'�6q�¡9G��P�ȓ�L��6��9J�Lre�T9�I���p""g�����z� ���4��:�&�5�ћV�`�W�]�!�(�ȓ-��x�F�Q���S��[�P=��H��#�g4��C�/�I),�ȓe�Zy�wÔ�=ô�;�d�~�:���r��}�'+��oZ�X'F�f:�5�ȓ~)�3���g~�1��/L�	��8���0�Dӟ&���JdC/�t\�ȓn���s�
 �B|�ī�qF&���l��	qDÝ<�vb���GB]�ȓ-gX �%иN�^<Z��2)���h.���J=��0Ď�x @���@���O`� H�΍'W H��Tp�8�	{�p���C�RGR��,�f�S�
�&u$D3�GGoJ�ȓhF���m�4�>ȳ@frn���ȓK���a�Ď!50��\[�T�=i��̮,U����[2zw8�Um����!oU!�s�r�PWjD�:����G��8gS��
'��^8eV>�)��l"u�:Ɏ�ʵ�� ����M!���|���Ӓ*[�8 AQ�Q,�Ia��'�O� sɋIǖ�mIT3��zv�'Ş�襽U#	j}r閩,&2��0�A9M"�pJ��yR��L���rw�A1jR`��P��� o\H�pk�04"*A�@z"H� [���ŖA�<� �P6��"���H�t��UE�,Jm)ő>awK
����&]ܝ��A��h�����Ɖ0h٪�<���
&_ޣ}b���2��;��؀U,̱��J`Aө�: و��$
<>�k�CT{�r-����6F���cAû:F�O�Ss�e�HO�4��������b޴a:�,ȳj��Q͌B��!]�D��D;w����FJq t�dԜ"_N�K���m�*�(g�G���	މO���Z����G��{�ޡx�f4
	ߓ6]�=�'-G���6mS v�f�9��Jf���P�!t�d�O�( �3?�p�\!�Rh&��*�"��r�Ao�5[`�ea;?G`#}���8�(I�s�0��o��Q�t������0?�8"d ��N@�C��és|D�k�Ǔ���h����$1����*DM`1�ȋ�!�d�z��h ��ô	Uc���Im&��v@~؞��uf61��t�7���j��s�E4|O�Z!�>"QHѱ�47!�-@��ɱ!���K��?�H���K.<�+�ļI�İ!�ׂSÀ��?QPʘ��R` w�?ҧW��)9э�Ss���ff^�cll��6 5�C&F7�\�/1"�V�hC��8ajyK>E��'�`�	�㉏`��Iҧ�ӌg�"���'p��"�LJ#p��H�&��/���'S.�Sz��%�HP>^q*F�^�nA.̫�	<D�@X'�*:�<�p�`&
D��c<D�[B��.��p
]'HǞ�U�(D������L��Ʀ�B�
&D�� "����L�DU\dӒ���"O�TqΏX[�A9��I"g��A��"O��HP� c ��E��~{zh��Y���aT�ܢ"Ez]��˰8�2y�ȓ>����ԗE��3�L�nX�ȓU�"�ˣ�F�q^HC5,�m@�q�ȓx��Ma�iI�wd�@@ &֫hcF��;�2�p�-G�dU��ʁ������ȓD9���ŃN�А�$͜1shP��|պ$�un*^nz�:���z�Ҁ��+򜼉qA UD���@MI,���ȓl��h�D�A�x���;U|����e�Ȇ�Lm&���0'�;9�6���v׆,ꗫX�(-�SF*Dw�A��8����Z����@�P	
:�Q��<N6e�pmB�L����s$x��u��KZ�ZuHB������C�e�I�<��jB�1�x� �+����gF�_�<	d�սN�:`sb��8=��M@O�Z�<�Tf�"$�@q���3R4���#�m�<Y2ŕ�?�A���}��3dQ�<�doD�,�"l�P/Д���&��R�<���n�>Dh0���wji���d�<A�0����U��'��l�FOf�<I��y(-��f�T�<��gÙ`�<�f�>~Ԫ�Qa!Rk�.P��o�D�<����,�;A+�'cNy@��@�<Q7�8m�i���ޞSB��7��v�<�v�4)"��`F�m��@�T�<�	@?&z,\���V��Q�G�U�<��뀋1'ax�R�i ��Hz�<Ya�ձQ�� .�h�FpP �Zv�<�rEJ�8��iH�'�2AW�}@��Lz�<i�M��<���X �P� d{�<Q��]%F\�p�gO�/YJ�Y�&r�<��Y�8ܒI�v��|�����o�<���Ć7r�M�&�6���6�~�<a�CA�\ш�g�_0�J��2�G�<��ϳ?]�pJ�������B�<�W��L�=;À�+y�Y[�.z�<�Cb��ʬ!��Bً%R�[�w�<�D�Z~$�!->sn����J�<��C�5R�l�T+��^�؝�����<�gN��Y|\G+�9/L0�R�PC�<1�H8�"Q��5"΀���a�<QH@}��I@�H4R (D�V�<9��U(#��#u�Kd����Nv�<�a,�Ă
"�ҹ�4'EW�<I��ݱu�
�b�,�M���nNw�<��]l� �@�R�38�J�<P�B]F����,|U�e{���k��p��J ��	;�Q'��!�l�FW�C0�(�I#+��%�?%?]�6��7}#L�j��!
�d8��&}ѻB�O1��	�RnV:�H�K/k��i1��d��@ �$���O�� �{J|:QE��\�]"��R/� 2s�	C���2t�)�IRa>t�9#�}�T�P��^�&S�'�p�Dy���L�#p�V�01��	P�	2�J����	�(O�>�k�<d2LY���^��x�7�k�bɘ��N8�_|Rى3���C�k��I�K{T4�bI�
�0|Pb·l(�j I��
���@��	v�
���H���ą�-�ldzrB\�/=�����E*�yB�F&'&������S5Wh�a��U�:���닦iDH��ّ�\a�C�z?)R��k⓺A���4�>A�\4&Ujy3H�G^T�q���P�AkB��1����˪5����Y���BG���ӊN("���U�a�T(��O�&�"~� �P8�H�7&iЦ'\�.C��ʑ�K#��"}0��4��B�OՊ���$L|�f,�I�޺�
ç#������XnU�L�`��]� �'�H���?�qO����"��6���+�ဗ\bȐ��S����f���S�>�g?��ܙ�E ��KN��b�*A�@6�|r�H�@ b��>��gʛp� �	���#�tt��#D����H���H4A ���7�!D��h!cɢ(y���D�d2x��?D�$�쒗��%�B�O��P��C<D�
gƛY~�{�C�r^( sS9D���l�#=�R�U!F2i��2�6D��S-II�رX	��i�y�s�9D�t��������O�"(>��BT(8D�`i�$�k��ո1�-p�,rr�6D�|����&\��� 
[�'=�PD�4D����8p���e�3'U��� %D�|��D�jK�LÃ,�561�<�a$D�����JJ�m���B?H)��&k#D���d(&N, ���4p	�P�&�"D�x��P�]NT�{�&ʝY�|$�7,!D�Ԉĩ�!f�<�'�%uy$�C^�y�{��8�֕(m�%���&�y2Ɩ�Y0�mC�#=x�tC��+�y�hW�_A�Y�/ �N�R��G��y�b'Ƅ��Y;�XPU&R �yrO�,����g��^\��D)Ӓ�y����&���@�� P�d��yR.�K�(��W��9
�������yB�ь+�8P��˔�uܜ����y��ןL�zM� �F�f� B��P>�y��NWL\x��\jNɹA��.�y���5���H RN�۵)��y��?<����ꕣ>�6��4����y��+sL�W#6�J��tΚ#�y/z)pr��lЊT�R�Z�W�j���8e��c�qTD�ed�4�lL��^�M����&�e��\:"��ȓ	Er���٤94f�8�C K�h��\�^MҢ��kf�HC
�-"����M9>�RQ��/�����-k�R ��Ftj��� =i����F)oވ��a��`�C����=�t'�.T1&�ȓ:�ڨ�4�_+r\��S��.T+���~��Is�E6tQ��iGc�$6X�\��?@�ı�MD�7�\�9��"] >5��4�t�p�c�+R�µg� t�`��FI��
��þw�j<���#x�hi��AJ��"�Ɉ\����2@TI|����M��9����Ri^�y��C�RՅȓAav12bQ(V(,��.�6{�lT�ȓ*�Z�I���f;E�.G�V�E��Ne� ����q���$���EѠ���9�)��Vnl蘤BA���ȓH:D�j/r	�E�Z (�J�ȓ/� iv+L�wG�9�I_:W�لȓr�4����A��2b�6*<��ȓy/*��Be�P^y��a�)���ȓ�����1���3���A��y�ȓ
�(҃١;�:�c�G/R���ȓ �$�%��$��Ÿ�D�O񊄇�a��P0L�-5>b���G��Z�d���}k��@T�U�,Ő��2_�Tl���e hi��ف�����Y G�D!��'�n� 
%B��u���9Bg�ͅ�S�? 2�����2>R��FX�<v����"O�]�$��
J^h� �!H�}Z�"O&8{7�Q�Z�5c��ӶM+Vu�"O^Y"g�[Ac6�yV��&!$4��"O�h �ŵ~�h�%�I/@���"O���*�B���)�癬T2Bq�$"O��02�F�"�H-p�� �"O�!��	�6�"�ig�C�k�k�"OŘĂK�:��j���g���E"O�(�I�\�h-���C.G>a�"O�Q*�� �P��q�]�1��a�"O\�2��6`[��VH�����"O@���*H�A��@37gףF���"OL�˂�ڄ��i:���eg�=��"O��+@OXK� `P�^�7b$ͩ1"ON��a���Vڸ�bu,A�w�}�"O>��&�+����\�, S"OT`1צT93��(BI�nb���"O�]JF�͚A���#@b�M�V"O&�pCR�4��qIw����HD��"O��'FASV����U�,Z���&"OdX� ��5:̪�G'N�t8z���"O��p�5q|<���fѷ˦AK�"OL�d捚 X�h���'L����"O�	Sm��IE�sM�m!�3�"Ǫ2uÓ<�ѫ;,�֨�d"OА�@�u|��Ib`=��"O��cÉ�<f����fp�;�"OB�ò�W�>�)@��;bS�"O��aAJ��9�W�r�6t��"O�ٛgV�8�n�h��a�l��"O�S��%��$�t��#��0��"Ox�1�G;I�p!���ߪԺ�"O�����$�=���L=T��&"O���� �� �d�I�O���T"Op)CE]lw�8��q��f�>�y���%g����Vk�,���0F�Ԁ�y�#ڿG�i:0k�!qa�Q'�c�<yu���#�&kD�3o:������X�<9�(��7�*i��L�d
Δ���X�<��M")Z�T�DHH�Ms��uAW�<��M�J�2!`E�:�Z��w�R�<�"$�5����,�0�"hB0CXw�<�A"|dN0r��-J<\J�AVj�<�Q*g�t]r$��N}j�h���9�y�Fd��Y��O?���`t�P��y�F�`{�\�@�*2����+��y���3*��,#�*[��l2U٘�y�!&�� ���M;��Q3����y�K�?�e��ݚ%Й*$K �yr��[}h��FM�# �a�GF"�y�+�?h�pa��O�)IfQ��Ͳ�y,��y��&A���� 6�	��y�P�ri8�p���F�
��eh��y��'����Ĉ�,�*}�u���y�ğ)J����1+߇���lJ��y�i�/P�����`ȪX�yB���y2����iŘN��9��b܈�y��b.4Ţr��-J�iEI �y"��/F�)�UC�G�h��E�3�y��?0��*�iR-9wb��d.�<�yb�]�vp��3)E5"���5�'�y"�ܴ ��'��� ����yRf��8�y�D��-¬���J��y
� �I�1�Wd,�ԡ!eƎJ��l0�"O{���`�u|
�2�ϝ2Z�ܡ�ȓPb�њa	đ MX]�$��:%b>�ȓ��p��E���KӎP8]%��ȓ{�r%#�,i�H��H[�9׺��ȓ/����� �c1H���E7.���ȓD&f  H�5H><X�#Oɰ/V`�ȓ(�$��e9s�! $h��5"�ȓ|FF��+�36'�0����'Py�8��o��H��4MT<ii�,*Tt��s=f`�Vŕ>��� �>�ń�=�,e3e]�8�F��b�� nl�P��?��1��AH7�����]k�̄�/�v�@$��eL"HK$ꟊ5��e��nB�rb������fϭp�0�ȓV��;RI��~	ĥAcT�o6���0�}�O��J�fE���B������"��6U�ByyG��MGPu�� �V`;��Ÿg]����c��΀P�ȓ��xPD�۫hh �*�?�A�ȓv��4P�&\~�p���g����ȓ�V�h����0j�rU,�;,�e��ah8�k�l�#vdzԇ;� �ȓe���*q��_A��a��?t5��ȓO����Â7d�fQ���8+�؅ȓV����
�i$�����F�^<ⵅȓ/d��B�?�x%���H-�H���o���N��]|�#��Ϭ-����T�� �3���V����D΂��݅ȓ/�P���"Y>������m��E��I�i���X%y24�E���W�N��ȓĢA86,GJ)��F��}T��2�\�U�}�|a����2�Ȅȓ&> �	 ��!
����1��M��p:����13tLB"�G.bP��e�~a���f��udb?b+@��ȓZ���	`�T�A��'��3#� ܄ȓH"�3q �Px������Y
���ȓ9�MI�KѤnRqB�!�r�p%�ȓ]�r���o�#@1"W(N�%�r���:��BF+R�wZ�IP�ߛ+pԅ�#8æ��
Ϥ�8En��V��Ʌȓ,�mM�t
	�jH	5h`�ȓ`'FQH����0�4P�&=�l\�ȓ.�PJ!���c� 8S��:��=��s��1 4���#�BF��D��rzj�
R�G$���J��T���
y��-	�&��T+���c3 ͅ�G- ��  �,��5�B��g,�-�ʓGpH����>`v��ٱ�[�@��B��4pƌ��hIm-���j%�B�	h�y"�nL�mk
�,�(l�B�	� ! ��[�%5�`�d�D�'cxB䉨��	����3Mk���#�0�&B�I$"qVe�te�5j����ã�cM*B�	�(6䑫m^=;.��n���B�Ih�t�X$)n��8�'U�B�I>���w#Z�<�!��/vFBC�ɤnJ���c�x�8�'�&z�C��| @���u[�(kqK�^�DB�=Gc��ۧ�* ���X�NdB�ZcRڞ1.|M!��C�_��C�	06��MB0$t���j��>	
�C�	'w��X��ϓA�P5[��\�g��C�)� &�`�dN�?(e&,Da�A�"O s�ʞJd��Rk`%�DE"O�Ի�I������^��8ȃ"O\+��C�_�����'!�����"O̅�D���qa\I�,�&D���@"O��;�I��U�P���$�.<��x�V"O�ܢ�K�a>�}	 �+�f�"O<,c��U�(V�Y`�Sk�ڵ�T"On�#$��%�����/�*ͩ"O4͹'.��i��l�a�ք72e��"O�u�   ��   �  �    
  *  V5  �@  �L  eW  ~^  i  �r  ;y  �  ۅ  �  b�  ɘ  3�  ��  �  0�  r�  ��  ��  ;�  }�  ��  �  7�  y�  [�  I�  �   � z! �' �- /  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%_�Q���m���R Q�t�A�,�Or@���A0��, '"ѽv�d��"O쌩��9al��;P���u����"O��d�AR	�N��>����3"OTP
0U@F`�q-�#D��`��'�I%y��]����Q�}���7i���$�>Q��ۑeK,āc��/:TR	еO�'���,�r@k�� c�x�x�iY+bB䉇KxHA�ׄӏO�jM�6��TK��	��'"�>�Ɍ[���zA&��D�Hq�2BQ<S?P̐�'��L)��?z�(�4[0�`��ٴ8!!�4��'�
*m�������q)�{��d��\���䚀r�V�+�;<��{��)Z��K���ѲBKG�,�4��� @�<��B_y�NtCD៙n���S��զqE{���i����j� ��i�1B\�#
ϓ�O�zP@C!p��2�"��yv>(��3O�E{��I;Z7��@'�4r}c�N�W<!��6
�\������椚�2.�P<">�J>yPmS�e�f��N�(3�v q4��H��p=�!`�=Ԝ�J9$���� ]��hO�'
Cn�HRJ��Y<��'A����mM(<�p��=�q��ǹh�����Z�<	���y�>�1�L�8`�B W�<�ЄJ�H�m2w#��x-�%��P�<�ތ��̀�ʘ.f� TO�N�<�#�	n��(�%�֢$Xd���$�"�hO?牝��A4'��Hh;@�*`u�C�	"���(P�"xyv�[J�Db��n~���O�Н(���O�^,
c�Z{��AI���dE'�2x�%
H�ض�ʵ����'?���'��x���7:R��g�'Kn`��d��?q�'ȰY쎄 ��G��n`��'ή����D�p�!Q�P�v4� �'�H�b3�Țe ApQ�\��{5"O�M3`+�`� � �^�4��g��Ȅ�ɖ;��2�.�2ye<Lڔ̒�7sF��d!}��<-.YS�%Ԁ	��l��L��y"��!!X0�Tc[O�2e0�N@��y"G�:?���D��I���RD��y�hHP�m��ȈF��Y�#E��y2���}qx�b��R�����'��?�����1Vj<CƦ��?��0�2,7D�dhAAڒ ��@I����Nx�	D�3D��9��4WS�ț���	2���A1D�� �YCu���~ۘ�!��t���zA�'�!�d�j$�8��1���c��sp!�$���`���ݙ^�&P�&IҮ,T!�%d��]��a
R�J����[�QF!�dZG ����]!���&@�>!�V?�N�؅	���H�-��O��8�S�Oavu��䎘���N2b���8�'-����<2��:�'��M�~("�O���I��<����O�7k�ڔ��0���>A�`ٽ����]�c��p�uj�ޟH���vx���F��:|ʢk�rΔA��F~���]8�E�C��c�P�*�'��
^C���i���9�A��T �~��)ڧ&�q����1��P�W,�4F����ȓ2�\LA`�W��<ё$O�<��)���hO�>�xe`��5���s�H�s��p�6D�\�r�H�<��u��؁B��g4?ɫO����!V���sЖ�hA��:��~�T�l2��Az�y��'ա77 ��%F0�IA�����&��@�y�&�U$j{�dA�d/D�P����� <Y��(TZ���A�?�IS�az�h],8T"(A D�?e�Y�B)�M����s��x{�f^&�~�*���?Z�ZY��"O�X�T�L�.AV�ZG�Α����1OH���df���5K@��B��Z�k!�$/Ei�M;�䂅}��0XUfܢ_!!����AsE�e����߅!�ѵ
]f�ȕl����3/�!�e�V�
�M
+����B�"�!��ǟHH4Pɱ@D�d���QQ@�y!�Ȗy�~��VA�tI�'mӳ>f!���1L�0a��3J��(���k�!�E 1<�v�τW0(��ѳV�!��$pӀ�b#��K�pl�-���!��%~�H3�M�&�N� Q��I�!�D�"Ap�<i��+p��aaqO@#\�!��³m��x�pk�.vV�)���x�!�d��00b���J=nY����U0�!��6C���l� �� ���$�!�d��"-�ixk�<���ʅ��+	�!�d���̺��
X�����CJ�"}!�d��G�U��}����-�!���o{�e�$]�d���1�wb!�� ��2�2R�`D�m;�]-@_!�Ę�D~�1�t$Ϋ �>�{�Ãw[!����Mp��>#�
<i2%°l�!�����`��7�$0� ��2t�!�ć���2*�B�l}"� �,�!��=F��n��Ҷ׊F�!�$ӽSq6�x�%%au|�o\/X�!���
s�� X�nQ�� ��-�#!�D��;.��q�#�4����"W!!��͏��+S�P�|��кBQ%R7!�d�����A�m�{�ݻ`��&!��rC��C"J�j^6ps��6`6!��@���5 )�����K�y�!�Dޙr*���&�m}h�����!
�!�-u��ar�[5:>���d�D$]	!򤘩~��l��`�!����7��!�!��~�8á,I�x(q�G#�!�D�y�hcB�ޅc��	b3 �4�!�$=�4�x��$�B�N-i�!�D�E�!���E����2�R�7�!�dB� ]Ri��GC�4 UB��K�h�!�� ��aY�X����H5� �10"O���A,M�x�x�O��2�v���"O��W�	-m���^i�N�2"O �bQȃcY˃��gf�x�"O����T*�^�5�`T� �'��'or�'}�'��'	��'@&�y�@8� U�
O��N���'8"�'���'o��'�R�'��'jMe�L�0��o��K[�� ��'���'���'f��'r��'W�'���N�.@~��p�6�#V�'��'���'��'��'d��'��t�$��hk� K���-~Pሳ�'U�'���'"�'_�'R�'g.�B�_�^��A��49�ae�'��'�R�'�b�'��'*�'���Ӽ�ⱡw�k��S�'_b�'�b�'u��'�R�'FB�'jV�1!N�vw��I6��+��lSd�'���'c�'S��'S��'���'�V ��Dޮ�B��0�̈O�e��'���'x"�'�"�'R�'��'������.-np
�G+Q���2�' �'c��'�R�';��'���'.d�P��C�k�Y�0�*$�"3�'3��'xb�'�b�'$R�'���'=����"
�{r�@)�ǎ%I~A���'2��'b��'Or�'d��'C"�'<�e�B�K�%���M 2 � 1Q�'���'�R�'"��'M"�m�����OR��DR&��q��#0Pt�u'Mxy��'��)�3?iU�iK0�RE�!)0b@��EL�`r��7� ���d�צ��?��<���\qp��QaW�^�l�@!�[�)������?�vd��M{�OB����N?E�oA5ձ�̀2x���J0��򟬗'T�>=i0L�+q[6 P�� +J6�)�(���M���F���Ob�7=���%)�S9�H�e-��젘�4%�O��Dk��ק�Oa��v�i���f�(�:"��@ ��z��l��+��r���=ͧ�?y�:F[�I���o���D P�<i,O��O�ul�`�b��N�:��m�4D��pЉ�P�3������I�<��O��JP-j}R�{e��G�&�Bќ���I$ڈmH�b&�S�$�Z1��l�t�Q�D��79����_��IUy������d�=(��$�!��2��@�GĴ9���㦥{b`>?��i'�O�o�}���I�u�<�A2�T�*�$�O�d�OX�ↀu�����d�ꟾ �A5u�eCL�_|~����������4�V�d�O���O���Iu
[槓�V�}�t&�'#�\�h��6H43��'����'�Hl0g �m�V��# �t�Ԍ �-�>������O
ְz�bT���P	 �}�,��bަ0]Fъ�]��� ���x�+e�	Hyҫ[�9nN���h+{GJ�I��Y��0>Q0�iK�<B��'��xx�!�!8���nY�f� �1�'	7�0�I����O���OT��n��TA@�Bpj� x�� ȑoɉ��6�7?Y O>_���Z��ߥ���l]2�&<q����w�D�I�L�I��(��˟���P�ו)�>DC�I7t� =�eE�/�?����?�'�v��OP�6�4�$6e1�uX���\���7��(pJ1O����<�r��6�M��O�`�#9���3�J[x,��U��X�Rh���!�&�OV��?I��?���be����O�.
��4�`݌
�,����?(O��oڈV������D��D��k[�D9cr�*d�����y��'����?����S��.�|���B��$%2��oVH����g�_2�ha��W�擑>"��L�	�yrL	C��o��kP����!�I����	���)��ry�v�N�q���aNX�F펍v6.�Z5�N�gX��2�V���M}r�'��Q��QA�>dPC�H�	S� *%�঍�'>�t��?A� U���7�(� 	�Ŗ��X�;�d���'�"�''��'���'��S�lc���pl��C�,@S��d���4q_T�����?��䧂?�F��yGj� Cӌq �_�Y�aj�٢d�2�'Uɧ�O�S�i7��@�k���8���H���#&���t�Z�)�'�'(�i>���4�H�bk.6JPq�0�F�n��ȟ��	˟(�'o(6���^���O��D�{&�=��P�m���Y`kH�F���lA�O2���O��O��:���?r�� r "���������C�����&擝�"��џ�*PI� Gb�4!�%W��M�%��t�	؟���ߟ�F���'��$CA�0q��E�ŋ`R����'5r7-�q�.��OmZN�Ӽ#D)�[��0��J��E��,H���<���?��8��4��Dб%)c��A<�1��9?�|u�iJ0]|���G.��<�'�?����?����?ARG�&>�R4�6o��.�fu�FW���DS�52 ��ן���ݟD'?�	�R^tA.�*��Y��(,^o�@¬O���2�)�SJ&� �GĀ2b脽�!oC�Gg�8a&@	{A�	�'`EYs�������|BT�H[����5�F+^>����W���$���\�I˟�ty�Ik��ܱF�Ob���ƉJe0�q�hBt�V2O@hlZF�'���h�I�̠��1����N �.T:�
^)J"��m�A~r�D>x'����Nܧ���  L(�c����UF�>j��L�=O����O~���OJ�D�O��?e�� Z�^�I�+��M`�A��I��۴y�h�,O: m�x�ɥnN���e�Bh̴Å�[�yxU&���I��S�e:��lf~b������#wP�|HFU�7c@�b���YRjHy?	H>9-O ���O��$�O,9:%�S?�(��kQ$N^��G��OD���<��i��cZ���H�D�z���
��hr�n�<��WE}��'4��|ʟ2P��n�$/��� �>5�0�J�l���5)^
(���C*O�)]$�?�W/ �D$(���ɦ��\벴:E�	�h�D�O �d�O����<9f�i@4`���-;��4se�G�<��͓�p,r�'S 6�!�4����'��C*D�U�&A����BԡA�b�'זm�t�i��ɑ �rŲ�ٟ���Ћ�)��BIɅ@[W��͓���O����Oh��O���|�"e;=����C�@�\dAC���&�K%wB�'c��d�'p6=�\���A�X�c�H@v�q��OD�b>f���͓SĊxPEh��[>��AE)܊o��ΓU��I�ţ�Oȭ�L>�-O.��O�h	�a��in�����'@��!��F�O���OT���<I�ip~\Q��'�b�'�Ё[�e1o, ���8 ���B��p}��'�B�|b�ʗRͨ��߁[#�LE�����tPu��|1�fp��|�����j�;F�ʿ�D3�9^C�ɮq�t�j4%X�|M֤�a�����[޴^}ƨa/OFyo�~�Ӽ�%ǚgLmpag��l�|�����<q��?���w�}��4��D�1(����O��[��к��@�Z���|b[�8�I����I���I���+�BR,O�<%��������P��vyB�f�f�{U`�O����O����Ɖ{���c�%O��0�.��?�Ph�'�'kɧ�OĘL��q�l��F/txH�@�\�8�)�S��!�I�s�\�	IyrH��S���Va�6d����q��,`��'��'��O�� �MS�[0�?q�-X+'^41ō,_�b�0d�Α�?�2�i��O�x�'�b�'�"�\5o� a$ń! �\���V����i��I/Z:pt(g����2$H_�RaT��@�
/�H�R�w�P��	�pe<�� -*ז<"��R�F�8��'��Lp�*%Pԙ?�J�4��'�P٩�-�;�$h.zʲ,�bOS����,�i>I��L�ݦ��'N���cY�c����%@]$����B>=-�e�������O��$�O`��|���ψ�WO.�P�X[���$�O�ʓD'��Ʌ/�2�'2\>���ؼ|��]À��)���#�6?yVR���	ݟ�'��'@����Njd�����lS�=�) gF�	#��=��i>=9R�'q��&�����
%t�,�z�͖�On���@��֟ �����Iܟb>��'%(7� -iv���'��J���h��GB��t�<9ǰi9�O���'�b,Ԃ��]�Π@^��Y#�� "��'����i����y�T�c�On�'R�	��f����E+�nG+9�Xh����O����O��$�OB��|.U�����,��l��aks��l�d�YܴN� a���?���'�?�P��y��ƸwVtږ!Z�)�fl�6ib�'�ɧ�O�z�;��i���D�QX���LS�QP��G)c�$	b��	� ��O�ʓ�?��KT>D�F@1G��RO��y\�X{��?����?Y/O�l��NЙ�����	�ʍ�q�[�ez�2"�v]�?a�P���I���&��B��SyNhh��
�"vT.!�%�+?�@'2 %�BݴИOIw?��mY�5`d.��k��<��E�_�8�*��?A���?��h��������^� dFS&�X�$W������D�I��M�M>���s��Evvy#��<)�\��Ƅ��<Q��?���?R��ش��$J$7c�5��O��,ITJHx�r�Q��4�N%�0�|�[��������I柄�I���#g�O�:6ĹK��}�īB+�ry2�qӨ�ye`�O��$�Oړ��ɪqp��V�p,�$:3����X�'�"�'ɧ�O�hT�ӥQ+@���s(�^(��YզT���OTHᱤE+�?i��0��<��ۀʨ���ȀX�nĠ�D�#��D�O.�D�O�I�<��iR�Py4�'�	���1/&���H�/&Y�Me�'��7�%�������Or���OH|�fOV+��<F�W=QA�A�����"7- ?I�ҋ^���+�����х�}��t(׉[�~�����q�|��ϟ��	����Iϟ8��䓧s�X4�cҗ^-�m�u�B��?!���?ɷ�i��T�O�b�`���O:�T��}�ite��i(����d�O˓j6�,xܴ�����[�ҹBC�E�Fn*!i��R�&f��E#��?A�;�d�<�"�ݐ@Z���͒]gJP�flϪ�O�l�0 y�'j�\>�PBl٨�����cY�s!tmp��!?'Z���Iן�&��'q���S��@!p����jTI��q Wn����U �	2��4�>���#��OZ)
B�����2k��~�z8�0C�A<ǼiS�):�ʟW�bQ%@�2<DD�0�
)C5剅�Mk��@�>�B�^]r.Ҕh��T<�#���?�(\��M��O�����4��^�� ��i�j�_���ioV�iF�� >OR��?����?����?����I�?ib��$�ʒ ��L{R�B�Ij��nZ�;܆L�'r����'�7=��� ��j���������#�+]B�'Bɧ�O����R�i��d�s�>A��N�$[g40dZ�}<�D�@��yI4�O�ʓ��d�5sdqQGm�&R����hR�Q4ax�Oc�f|0e�<��?	��Zb���� Y�"�b��鹋�>Y���?IJ>a5l	�iFUؑ��S(1���k~�#YNhC��iPȓ��0�'��aݔx��9�܀HQ�U�`ł�H8��'
b�'v��SƟ$i�*�XĈ YW��54F�� �Bџ���4@o6Q����?��i'�O�N����!��@��F9��{UoT�t��$�O����O�p�hq�B�+��ջš�?���,�2����-X T+��LY�	myB�'�b�'���'[�-��n}��6��q�woW��i�oZ/>���I���X�s��"T.nV� B�ߧŰ� �������O~��$��F��QB�g%|*��n�k���r�%Q��I�5��US�'�i$�X�'f�����Y��1x��U_֦���'��'3����D[��Aߴ:X&q#�o�\��vn�/pY����.2��%�fڛ����y}��'���'�Z г�_���]Y"�ګ��\��� 5C�V��Rs��(�4�����aQ��W�0�� �N�{J�;O~��O����O����O�?]��M�z����k�&U�
�10�����	ȟ@cߴ@μ|ͧ�?!a�i��'�5%�A�^ �rT�ŕ|�FÁ�|R�']�O��Ah��ip�i�]�T(�D��C)�)F����IJFL���>9��'E�	�����㟰�	�N�$UZ�Ax�؜yA��O�X�	�0�'ϲ7�P�L�|�d�O��d�|^ұ�Hԙ@�j�q�����?���՟��	z�)�d�)�8��#"�L�jf̗"K�P�
�Û4-"&5��D����dj��|��!O&E�5ȀV� �HI�J���'���'���dU�tڴr����@B&���,�l|�!
��׹�?���&�Ăs}�'/�0��JW�<��dom�6�:��'R�[؛V��T�2�յ�q���1�'��s������!$cT�s@7O�ʓ�?���?��?a����%<Z�����Q)�pj2լ-�b@oڮv��8�'������'�7=��h�CfLu!V 8�)�
5�� a��O��d$����|7i���&��
�PX�F��D�� �r�g����Eh�$8�$�<�'�?�g"�8�� D�6)��@�A����?q��?i����d ��	b4C[ڟT����L�W�Х'�"Ј'K�aR����f�e��3���ݟP�?@�@���Ӈ��@Wd�`��`~�8:9JD���C>H�O7NP�	>�G" R�y'*�)8Њ ��-N2R�'�R�'���SƟ\�3�Y�:�uF/����(�r��$u�<��e�O��QѦ1�?ͻ>Ê�����wܜiQc�[�Dϓ�?y)Ol�iӬ�5�ԅ��nៀ�0�c�$Qf*���E�>�.��F�±�䓿���O�d�O���O��D�8<в=#v��F�B#��m��ʓ&���I�)���'�����'@�45a�n��!g���B ��%�>���?�M>�|5��/�T=3ք���$	��m0hII#T�򤂷��-1�U1��O��DĄ��E:�츰*C*v �h��?���?!��|�*O��o��P,�Ʉ�pم�އfLzd��KI�	�M��e�>)��?��}��Z����HX��D�e���gÈ4�M#�O��z7�^��Ҏ���w>B$p�,
U���r��g��ű�'���'���'$�'O����`AHzh��V�f �ti�O��$�Ox�lZ&A�,�Sџ��ش��o��`7G4�̋b�e��@�N>���?ͧ?~)�ڴ�����L��jm���ź"��+��F�A�*��׶������O����O`�dE�aa�,˴·9z����le����?)O��lZ�N����Iɟ���K��h���0���N_pTc$��2��DHp}"�'�O�S:�D�9�'[�Q��4�%�>�V!�3OT2W�d���Qay�O�X=��6G��' ����.�/$�ܼ���/(CM��'�R�'P"���OA�I�MS�@�bQTsӅ�U�]� @��>���?A��i�O`T�'�lڇFB0L�W�P/MA���P�N�AA�'���t�i��i�%�̐�?Ղ�Z��)�%�6Ѵ�6�c�����~M�vy��',b�'���'�2P>�R'������kY�E����M�'��0�?���?L~���dݛ�w\�V�]�[�( �Cm
�jڈE��'u��|���UZ��6:O���_�l��	q��>;b�PHw4O����ܐ�~"�|r^��ٟ�ە��Q��t�Ȧ,����!����I����	xy��|�:L�c$�O��d�OD����ӜV;2H`D�U(��8���4���O���'>��'��'�v!KWR&UH��J��߄3l���O�|ї���#8�kR�:���?9R��O�*��]n�u�#܀5aBf��Op���O����O^�}j��> �ҥH�1����;��(�����_t�B�'H7�#�i޵���\��E򰈈�bux�S�i���ITyB��	������+6�1����&� n�����r墰�Ӝyh��?��<����?����?i��?iPŚj�h�0^'�0 ����ۦ!ZǠ����I̟�&?��	�BZ8��M�z����W�qíO"��8�)�S�I۲ i��/�=I�K�B�D���-]�F�l͕'�
91fG��t���|rV�8�Ie��q���R-YБ������L��؟�SXy��n�|�gM�ORU�2�K��0���GB�����i�O��oZF��+������'�,���BD. 2HmCc�E�a�b {U�U�曟d�a��$J����^������������a��3��F�r�(��ҟ��IƟ��	͟��23h�72Hx[�]�t~�xـDb��'�2
gӾ��8���D��&��g��(H&��S*|��M�%�k�	��L�i>�BF��Ц��u'�iƊE�b@�>	���^�I(~�r��W��Ƒ��I�fZU�gDʲb�V����U���gU.dr���'�R�^�ΐj`�L/S	��REk-$��`�vj�<�$$�V'D�v�<�[�&w�l��nE�vC(��<Q��J�(D6E2l�<S�}��@�u+���"�S�'����e۳i�,���#H?$^ 5��Ӵq��;�O��a�$+B"F�[  �qg�W8w֐Ss��H��F�NIz��!0�"�����%I�oh�D0��Z/f���	� `�$9�&1�S͇|�s���,5�0�1��"���b`үANY+�*�Ӧ��	ӟH���?E`rj�'{ j�(@����r�/�����?���'H���ӟ䘚dg�4��s�@ #��&Y��#�K]��M���?i��ʇP��X���$�&�D3N���I�:��6-�O���P	#����;�)�ӹ.N�@��u,*���p�6�T�o3�|m�՟���ǟ���#����<��%�?e��Xe�7=��@#��Ƨ^�6�Z:��O��?���2I�ȉ�+��b��G�E9	/�\ٴ�?Q��?�uL�/#��Ky��'|�$C�%8bx�&n:X�\��f蛦�|#08�� ���O��D	h�,�Ҏ�#�T��
Q�\^�o�埐�rE�+���<)������`��.�@�$��	,�`�)��Bf}"���e�"]��	���ty�B
�CS�q23 ���4X�v-Y }3�I�>�-O��7���O����^KR�s �T?�B��%@��x\Z#b5��O��$�OJ�l`���F9�n<30�ԛ9^TkD%�'m�Xt�d�i�	ß�'���Iß��&Xg?)q��',�\��u���ͻ&�m}��'*��'�剽j��4*��J��ҧ=��I�Ԫ�bv�AI��[�@�nZӟ�%���	ӟ��%e�@�7�� "Xp����ʇ�n�p�n�ԟH��|yY���'�?����"(��L�UM��m���
7}�'"�'ܱX����?� �Ǥ8��H�@�� |,�*�ho�b�v@���W�i�R�'�B�O6,��Ck��!�:��gi�,H 6	K�٦��	� �`�g���O� �$�ؔ0f�A4`�;�b0:�4�#$�i]R�'���Ol�O�I�$�!�#��2r�O��`$lZ����	ퟬ%���<��s����U�ܭ  �	�ц�!	������i��'>"��S��O�I�O2�ɗA�9�4H� j��I��\�6-�O�O�%��yr�'��'���/R5q,��s�	$xs�%�Q�i�����kw~<%����$��
h*X�zE���V`ڔ�ē�?	J>�,��D�OVŚ�	�o��0q��w>c�@6r�b��?A����'	��O�	00���F0�sQ���ꬻ�i��-)�y2�'���˟��&B�}�D��L�,�8&%�/B%NxZ�*�ަ��	ş`�?������^�0���"�.*Ȝ�b�_M���
5���?�.Ot��D���'�?�EeJ�rT�H8��[^� �'O� m
�F�d�OJ˓!_�$��)F�٤)T�%�a��.H�P�@�t�p���<	��Z++���d�O��Ƹ���GI�}�,i7�]`�X���x��'��ə@�l"<��gj*i��|�q)b��-G
��'�R���k��'�r�'��TQ��]jwN,vF��l)��SC��#O�7��O�ʓ}Y�FxJ|2qg�l��sU���=��	���-8�˟�	�����?����I�-��4�eKl�%�Q�N��'�훌����O�4ڰ�=+��MJ�J��v[$�����-�������0�@N<ͧ�?q�E����t��]��Š&�R]��i���'剜��I�|B��~#]�m��1�`�:2M0E�$?��7-�O���"b�<�F^?-�?���TI.���ďU��&.Zxȉ'U�}��OP�D�O�ĺ<I��)m.��HRG0a��p�s,�=�p��ђxB�'w�'H�Iݟ���j�p0��Ö(��;!��� ��n�Д'��'�RS�<�e�֭���ㅎdE~9�rJSv�&�ڴ��M�)Ox�D�<����?��tɐ�ϓ�<J#-�,Q��OW(r���c�V���	����Isy�h^�J?���?A#'�Bi��&�F��@�<u����'���ǟ���˟X2�nn�p�Iz?� �-+h�����9fM����Ѧ������'lBT��f�~���?a��KP�L�6$M�4p9ڐ�[����S����Ɵ���0C0��'��$�?uidi��$���hƂ-�޵�e�q�.˓3<Xh�¾i��'�r�O���ӺC��-Ek>\{*�/|�����q��ǟ\xp�2?�*Ot�>�2��f�ĵ��g*C��{�arӮ��ƌC����I��p���?��O��C}� 0�ӅI��H|��7umlL	�iu����'��؟����E����`�
4� ���P�+~��`�i��'�r.��������O�ION��'B�Ow�0�r��qD�7M�O@�aǐ��S���'���'NN$�T��4m�C��ʷw�r�ەp�(���sibP�'��	�'�Zc�hL;f*ׇ;d�Ecg�N�[�����O��1�>O���?A��?�+O  �T�2E��SH	6NgZA`u�٪3���'B���0�'C��'��G��Z�`�sb��*2�Pc��cc�5a�'��'�"�'��^�АT�آ���S3T��3�Eڃ7���S վ�M+.O����<!���?y�;*� �'ߔ@�ᆒs���2i� ��5��4�?���?y���D�	*ET�O�R �	��krŢ8�v��
?8
7�O���?����?����<A-��vΛ����Tb��@h(Dí�M���?�)O�i �͟K�4�'��OZ葓�ўzs��p42���@�>����?��e=BPDxrݟ��c�%�m ژ��I@�S͒	{5�im剅J%hap�4�?)���?1�'p��i�i�"�8�L%��k���^5y&�sӆ���O^�"�5O�p��y��I�gF�����C�[�,�RI���f"	9RI�7��O��D�O,�)Vz}�U��3rH�-:�	@�B*yF�5��Î�M�����<QM>���$�'���p�"�OI
�ۃ�]&��y� k�>�$�O���Ȳ|��i�'I�	ɟ��}2V/�i�P[B�8a�Tm�� �'r�Z�����OV���O0#Ҏ�	6����߳S���'�ܦ���5� `�O���?�(O����FMQ��M�,��0���2�.���[��(i���'�r�')V��q�M@(��¥C9B��9Y���-Q�T��O�˓�?1,O����O��0i�,�p!��Y;T�9��7#�|�k�>O@��O����OJ��<� -0+���){.�t�1��m�4�a����A��_����gy��'?��'��dk�'�\0� ��ǒ-����"Nuƽ��`hӢ���O���Oʓ3���*�^?�i�a����gv����.V`�`�Y�gpӒ���<����?A�%e���Oy�6�1����)����ULV��V�'�2U�,�t!���i�Oj�d�X����8��}HƢQ�3���gf�`}��'��'qNUj�'��s����&�U*��k��:��+w�Ąl�DyR���^7��O4��O���k}Zw�������D���5 �|�l=��4�?i�Bz�|�d1�s���}*#�ʙ��ģWF��*������BC�?�M���?A���"�'�?����?qs��Q�>Аb)&*^� ���1��V�T�S�U���������$�]j)�h�7xJH��#)ʽ?�nunZ�� �I�D��G���d�<���~Bě�fF��S)=��)&C<����<���U~�O���'�r��$&aΑ�".I��epqaB�@6�O�Q���c}RP����[yB�5&/[�l@�J�e�:Pd��T������c���OT�d�O,�$�|ΓX�X���3<��T��~����s���fy2�'������П �e�|�Ь���pMU�C�b�I����I��l��ן��'^�[�p>��m�;�&�9cB4w�m8֠oӤ˓�?�(O���O��D�(S��ڴ�0��R�Ѣ~QY�E�	$��'���'�2Y��h7���	�O2�����GY�����}�@P��-�����Vy�'���'��t��'(��'������,b	�%�6�F=F�j8� �p�R�D�O�˓�� �P?����d�&����
R.M�@`"׻� �ˮOp�$�O��	�NI�|Γ���o\?i�X;�/��!ʀ%9ӂ�&�M�)O~0il٦��i�7��O�i�Y}Zw���e��5s?a�b���5l�9��4�?��S�V̓f��s�l�}�5mP1|���B�=�Y���H�e�/��M���?1���RX�ܗ'��C��N2�C��Ɍ#�@q ef�8�!�=O��<Y����'�l1���Ė�D�1ǥ�%�*�A#�oӒ���O��d��*i���'�������3�(��Ъ>��x
��k@rUlZß�'����i�O"���O(!5�O� E�1+�-�*Լ��W������ɒa�eH�On��?Q(Ol���Z<����,j�.tXS�K"}���QgW�D@�$e���'@��'>�_����0�|rUN��6C&��Ǎ!0g	ҩO�ʓ�?�,O����O��$́ H<��am_�f�T����޽Y���E6O��d�O��d�O����<1��R02��R��̙�$M5��(uؙbЛ�R����my��'���'���'*�|��E2X��ɹq�X�V<�-���s�����O6�D�OXʓy�0��A��\c����>Y�q��C�Q�ݴ�?IO>���?�s"��?�K��EM]�HL�wl�G��x�'w�����O�˓� ������'�DL��!�ޝ�ǀyH0�IG�A:WO����O�1@�3O��O���G$`���S�d�.)!WL�R��6ͨ<	�D�
���	�~����j�����V����BXIa)�����!)kӈ�$�Oh��R3O.�O.�>	�W*Z3`aB"�b)6�C$�hӠ�:����q�	ʟ��	�?�M<��P���4dF9JUv��k�o����$�i56��U�'��'��4�Ԑ�D����� ;�n��\RHd$g�0���Of��Ė9�r�$���	џ��C��p	�U�)���lܻ5b�l�Q�	$8�bI|*��?��� \�uS�ͻ#J�������
*0�%�i�r�F�8@�OV���O��Ok� ������8��%Qć��*ι�R��y��c�X�'>B�'�rU�,����Y�A1�a-И��*=��Y�M<���?9N>��?)��Ӌ>:�Y�$n	+]R�+�K��\hhX����OX�d�O"˓Ǡ���6��|��	ۍ
Ė4"�P�h��-��U�@��ȟ '�D��ȟ��D�>a�G�� {|*$�R�*^)ck�X}��'�B�'B�3k����O|��ɂ}���YF&�>G�r���ĉ-囦�'��'Z��'����'#�,O �iaC��Z���[�	��EoZ����	qy�S'x����d� ����4y����{��\z ��o�	͟��	�-�*��I@�	["`&[ez~m�e*E�\�� ��a�'︔��#t��|�O���O�D��.,�UH���r��(O�j�m�ş,��2#X2�Il�Pܧel�sb��Ny>A��`�	m��8o�^����4�?���?y��j3�'i��B3ĽI���"q�X���
��6�<c���D.�D&�S�8��+쌬A'�=�ʩ�I
��M��?��i%�MÔxb�'��O�11p��"� �d� f�L���i �'���%(�	�Oz��Oܱ�*�2X����A�n�Z�+U��Ц���0�2ٓ�}��'�ɧ5��ܗ:���D,\'tT�u�%�$����_�8�$�<���?!����<%���'��Ho��[b�A6>0N=@C�Em���O�����4(�jEfg�"�S5sS�C��Wk��������Ĕ'��H$am>iҶ��t��"���.F�����*�d�O��O��D�O^9�֊�O��!�L�gB�]�[AEt4���{}�'��R����>W��i��Ο��:�tȣ��e2�E �(��h�۴�?!K>������}�'���DS�*�d�&u��I
۴�?�������/Z��%>m���?���*�(��Y1�n��upu����;�ē�?�
�<z֙�SjM�!|�X�T�K!ڔn�zy���2R��6��`���'�� +?�4��tyD��w��h�)J^ۦ���H��\���'�Ґ��M�k x���NmӔ`!ᄉڦ1�I������?�JK<I��I>�͹��U =����֯]�H;�ɁǺig���6���,��F�4k�D�0���r�~ aC�ˏ�M�����D�q\�S�����F0�f�d(ޡ>p ��F�ܿ@��)�<9��%?Z�O����ΣvX�ɦ{�x-XV�#�Έ��e
�J�xB䉷+�
���� 4
qJS�H�pr���C�C����"��ն�Z0�(%Ǡ8k�,�4b���rZ�8x���yl�E�W�<@���'��=�y��\s	qb��+*�9����g/�lB��WO�X�BE2d3�����+nu6����(7x<�#w� }��摟?�4m����HSP2�GB�wld��%��H:� ��N�E�J�����?	��0�?9���?���?�L>i$#��\��@�n|B���\8�Xks
ފnp�=���-=��d\LVX$� �ߩ�FYce/�0I�x��0�?I��B�����NaԦ�8-�y֥��T�f�	П���T���O!�T)�Ƅ=@������sOj���'��6�ɾH�dY��l�(xG��J���p�J�o�ay�ȽO=���?9.�8� ��O��a��j)b1ڢ"O��B!Pdh�O�$7^ 8���U�l% W�Ɵ�'��)V
v��}��,Ψ5#8*dkف{�y��	���09fPCș$�H��iK#��4��@��BR�m�v�>�Fυ�$�I|�O�bJ�v��� )U�$���yr��6�d�����ăĐ&�ў�S	�HOv�����	���4LķZm� �@�Φ��������dl �j͟���|�i޵R��;�Ѓ��)P�F!p+܀���rE���?�7�
�5ق��|&�᥉ܥ;�0	���Q���a!N�m�Xɳ ���?�vjK�P�>�k���F��Ę�B8���c$�Iw�p�g�U���$,?٠�ȟ�T�'�44����.�<`���-��)��'ܚ�p"!E{������U=���'8B$%��|B����� �<Ɉc�IF��2�([�	҈=$��F�����O"���O>ɮ;�?1�����ŝ�>=LMe��)`�(�hѪ;�b!� ٌf����=lO�:̒�F�r���O�z4n9p�MDd��iE�3=�$��퉿#��i&AC3M����6$����OP�D8���'Krȡs+ɥY&��m�	<��3�'�L��C��3�.�XUo�i�B��y��sӦ�d�<� ���F�'� �4\�`�A��H<sV�HRV��'���r��'hb3�"��'��'���$��sz4)x�U;���;�=�.}�?!@�P�:��(��'�V5��R8���s��O��$�<��/��W� ��7�ջ <i�f��<q���?i���ٗC�`����^9<��5dH�!�D�WM;���CRkA
k�D�c��"\��v	ȵ�M���?	,��s���O�������@B���U1"cN�E#�O��$FD1��""IC�|2)���{寋,k/��X��ϗG�Z=7�>Q3�ƃ�L	�O>�� Bm�'�Ǘ�Z|i1K�-\Ժh ��>��bş��I���IJ��8���'�G`N�%1�J�Uuء�<I����<	��]�g�(�J`���Fr�*���H��X��d��4lBR�ϸ1�d�E`I	�TYoZƟ��	៴1�
؆#�:\�	��H�Iߟ�ݬ�PY�5+���������Xg���I!��}��.�l�t��ɡ>�S����̼w(�WZB��0�ݫ&�����L3s�|HB���#xY�%ӛ'��hh�(U!F���	&��3 �����'DB7��O(�z �Oq��	��ٔ�:#����F�~�ԕ��nU��\$��z��˔P_���׼Mt\a!��c������M{�i[�'x<�%�O��I V�	C͟x5� �k�/M�B�I>B����ꜿ6r+r價-�C�ɂT��q4���7:X� l�J��B�	���,���J0HC%�̟e��B�=K|�`��%�-�$�
 ��k�zB�I�lv��
�!�;%B�qa��C�	"+D2ղp̎�d��1�^����0D�Ģ�ԔDR� pAΎ�.����/D����cɭt��,ZS�R�u��ؖ�.D�8@��zlL	JQ�W�aPg�-D����tޖp�#� :�䓕�!D�$ȲbļA�pY��B6^\��[�:D� J5k�
��=8O�J����9D�t���ܓ^�=ط���4�Ȍ9'd5D���k�`��)�f8�����&D��#�b�c��|AF�L,���7D��)ްi� #�ےQVjp���5D�,���ۅ.�h�ٶN 89�a�s�=D��CW>k�@�X�Z?��*��=D�4��d5�D�g�էxĝ���:D��X��%#0P���$���b�7D�L�@J?=�4��@�t�pP�l8D��X�#�	U�a+vIʼT��T: �5D�4�تA��q��.Q�T��n0D��mՌn���2.	4�D��/D��cq�[GV�%3
*r �	��)D�4�TO
�[�r��i� TXsA*D�K7�J�<$�2��Z�vK�@ꃁ&D�0���PqXDB�kYN�6�Y'M#D�p�l	�O3`	u��2|>,x�L6D�@�eG&f��Dq'MǍw,���g1D��r�gV�x�V9�eǔ8^P���
+D���D��:���褋�%}��'$D�drT�ϷB�Q��ɋQA�()!D�p"�eM�s�n�v�I/1�`�=J�1�-� ̲�V3^VŨT
�>��Yv�"��ӎiV�� �ג2k�m���E-6D,C��/���F� 5 bD�V��C�6�����Q�yRi�g�l�4̎BbȨa��<�y���*@�4��q������I�Zae������1-喕+A��Zd^B�	߷\�!�d8�L��W��	�<��w��@]qO��{D�W��0<��']̸��e�zYP�cS�Tg(<I���7g� L�V��Tu�T��ij:]3�#���_5���g�\j�u( l/|OVb���o�<J���X2HA0�X1��(D���2&�w���j-v�ek�)"D�<�e��9i�tآjP�C8D�?D����n����@�+�"\� DْK=D���C�f��!C��L� g	��9D��*� 5���8�D	��Y��c*D��آ� L-��*�==��" f(D���2,�8|�S7	��d�1X�-&D�����I?K%������"q  D���f�\���G�(�T��g=D�� �<���T=�Z-��G.9����"O|ة��\!��P�
6Ԙ��"O���q���2qA#�Jۍ+��}�"O���R��p	Ǜ=��L��'yh���"�	�q�2�AAG�'	o^|S#撥P��C��=����ڝM�Xh�����s�^��?�4��$���)�矘Q nR�j��be#�c�D��H0D���m��:n5�g�L0'0�TIc�l�H�'�F;��f�.a���	c�f��k�O�ޡѰGĸ)�l����}��Ls�4g�v��٫� D*£i����bӘ,ԈC�ɦ/K]@hn�]ӕO �*#<�WmR�ߖ7�U�S��� �,�ऑ���-C�D5����y���->4�S3�ɵ6w8�P�����Gk�ߦ�V����s�P��%Sd�Хp��&]�HiJ�!D�����S-PP����UhR�s1 k�� �-a�6
L�p&@�ታ_l��s�LPhx׍�}#���Dӛ.���ݴ[d�A� 6��͸�M�E.:��f����B����dPza혋�r�R�CD�0"<I�`&/�����3/���|��HE�<t`;�,^�{7r�ɒ(@�<	����6]b@Y���$�Թχ��Ij�-6�iݱ�P�JN�� �ޥc����(D+ظ"�Z�<���	��m���&f��:U%C�<�b̈́�N⟌ِ��K�=�D|xTf���fHX ��@ԧ�V�se��	��RK�Ov��(��-�3<6�t��.O.�>9i1�i��A���V�N���Gm�g�&,Y(�:b��3 v��S�[�d$��yPBթq�PqbC((�D%��K�$��7���k��G�Y[�ab@άٸ�Ц�A�>T�$�!g&a���(��;�|J�E���y��XL	��Ԏ$�������?��(д{H�J�����4H9
%��O�S,1�>48#�<j>^}`�ÉxQ��<a�ө8���S�s�̡��%��'`�Q	�dZ�`�8Up���� �4������'~�S�*9`��I %�����"��5�U�b �ݸ�E Ux�ij"��^4)�έ;�� P��h>�O��'ZCt�z�Nŵ��T;s,V�Q��|%�T9w$F��}�1LW�jT])��8�"BM:�H_!آU�(��$��)�%,��3	��O��}��+Ϡ�(cJ«lrcG�Q�e!����r&$���(6��ʧ*K9@�w�ZyaP쏳H�|����$z����FE�9�������=apj	�_�B�B	��0ӧ��Ԙ'{�2ׯ��'��A�Aa$*����	V���9��і�V)��)��y���FV(��'in��b�3c Ijd��w���W�Ԡ01���V��r�Y�;�E5��'��S�P�^aȧ�����աOe�x�O���ѩ_7%}x4A��<Jj�����9-|�g�@a+�dC�0h1���ʗ>V�'��>���!.���J��P� ̂aO�^����꒮</4	��XvqO�*e<"ͻqY�AP�60�`j����5l��c��|R�����=9rFˠjf����b��@0 WƊ'@1SΚ!B��b�Y��<�6�����\�vuq#C�Rx���� 0%vts'Kɲ-�l@�#N��.G̭ȖF�, �X�N�5~b4�v�̪,���I0R��<���7���P<פHұX���ٳHJ+�t�O�۷@ZMtT�wE�]{��8�d	�	�(�"��I	Ni����	�w2������$�3od˧�Or��P�E�D� 1�ES�R����%%G	O5ZEI��2�4t+�{ʟ���!�w5<x`�㖙R�cC�
����ʓ'V�n�+A���z��{�^�pt�����F���!�1OF���a��	C����y��=Buo�?Zܠ��A���<Aqg��ܡ� �Q��Mm�(@*�d��$���*,�Ƀ�� V�A8��OQc�6�剤���O��U���PS!ԉ(�ʘ�4�FMsT�|��tFLqP�LN�3J���'Ȳ���A��~���d��@�$[z����'~L)�\>1Fx2X=p:܌��`�,ݣ"�\������ݸ�ȰUH�]�S��L��5�4mj`҂�n�]��%ɭu(\Ң��!f��0�B��E���P���2}1Pb���#��%�"�B̓c.�$�*;�)�T��f�m���Q��j�/�#}vֵc��v�����6���ˁ{k���`,���mO�U�9�l�;g,��{�������O�.�bd��؉���8U�Ы!b%yF �&aF����Z���d2(�fuⅉ�E�����ɸ'�V�S�E*�P!qԣU�KW
�I�d���@�R2�Z��p������O����+���	kc+DXh���B_�`�HQʔ��t�FH�=E���M�U��}�W)��������Xm���Z�χ:�	x���/
.��Ҳ�U�5x�|�Q%��wZ���'ΆI�rdR�(�>yd���d�PQ�9���`� �)�ʜ�6,�&$���9�ʀGYd��?A��iC�M�So��s��O~�C���π *9JTmV!o;z�+u̓�K u	0���Uf$�@�h>�W����Ojb�*]a��%{���k&���~�ɏ8\�����D��ቡ_7�4�2`�=$�c��[���q_3o�6�Q��O�ܘ0�ϸ'0�LY����b(jch�6*4�`�PDԼ|:��'��VF�mD}BK�I�D̩ůSk?ɢ �+C'�\��%W��8��枥l���0pJ?���f������:pV��`�y7��#��䢢�Z.#0{���'�0y��<R�x<D�����0�ND�o�r�3d���y���7��d�p"_�Q�����<m�j#**�ӟ.�Q9GK�b҆=��ͷ7������34d"�O��{0���~���'�HI�"a�+e0�]���&@�A(���d?�'ᒭ{�� �VZq������YF,����ȨV3�q� ��*�ȩ�a�Zy��h1�
7N@h�`e�ϸ't԰�CB�<�m3�����/fH}j�E�6cU8�*
�~�H|h�M�U�6��R"Ix�T"`@7%v��A(�OyR��!1�ܕڑ��(��,��L�Ո��E��M#Xw��QH��3����hB�=�}
��ʠ��'��|��ڀh1�-2�b�� 	&�؏y­�E�,� .ܱ>��ɊBř�?Y��J!�B��c��(�ԝ�ĥ�E[,�&�Q�9O͓&Ю�,�c��
s��U�A"�y��E�R��2���y��E�Qw�E�1�۽C�t�%>��7���&}�q������;��X��2<�P
S-��S��#Ok��pUb��@*eغX���$�R�P��	M�<�fU�!3
�H��'�&5�hZ�5��*�+�L� �nռC�1�&gC���4��D_CH�Z7��`��)٠>��`�g�)�&��D�M�y�+�7[�H��<y�#�`H��f�8J�$mr��	p̓�\$�(,4J\{�Rmj��9��a�S����i�TKŦ$�� ��A6Z���S�>��þa4Ŋa��c!�њ�K��l�8�B�A�8���:�M���C��J � I�9��,@������q��B��&����I�5����O�/1�ԭH�ϑu���Z�{���<@��5y@�Ѡ�E
U>���CH��Az��R�$,O|�Տ�"w�]���|X��Z��R�BT�@��r�~��'9B!AP&�/~װ8���]38ΰCS�U(H:!�\�x0��I֛\�p�c��\#d*"Q�pJ6?��H�wF��С�#_�� z.�^� O�$ۗ+��o���s�S�>�H�OR�:E��+K����AJ%���B�)E��x�� C�+��U ��	dax� �݊T�@c�L<⑩�o^�W1��ԥX5H�����+�zy洇�I�$�,={g%�92�&逦�¯s�tJ&�"�7��!�b"扛v�p=���0� (��(e��kc�'��  ������ �nV8-� �",%�X�{���y~bMH6|�8���y�g?y���0hf�DB�x%��z�%�7x7�Q)�'Q@�'HI ���/���je�%�'a���@&n��:�N�)&��Xa�L
e��#�sm���p��|Γ0�2-cG��. �������&a20�64�� �;\I�ib(�pb2,է�O��}k@�Ԝu�2h*�(<���'%�ѐIC�lD���$O�%�sɝ?^��X �E@�Sl�4��*I2|���1ɟ% ��;�Z#L.�3�i>�K��T�2}H#O�oNڽj��D�d��|򢅖ҿ��jZ+��+VnA�5�⸛'mȰ.������"e��>�g�
�dZ�ؐ+8�	��Uo��)E|B)δK v��pA�(�EQ��3g�8ٖg�]��FE�G�<�cH��@B5�M�qnĳ1%C?� �9튍�t+��iI�3����/>�>,x���7*?�eK�ȇ�o�!��Dv��\���FpZ�([GB^m~!���&�"�s�h"e���G�	!!�dѻ5�X)+0��v�F�[��9Y!�Ͽ9��LHA��-B�)CÄ[�B!�$͸~�@���GH�O$" :�Ð�d@!���`u�Z��J�coԀ"ւ�V!�D݂FӘ��1ɛ�,j�:���=p�!򄅲O��2����6WF����P;Wh!򤝀4TP��ǋ:Rtt��o�� �!�ؚ>���3�*
�g�!Rq��6�!��\�1���:!I ���!��)�!�$��<�W,?l@S�J�,r*�u��"O�Y�h�����B�7~�t�q"O�q���� i[Jh��Z	sϐ�HS"O�I�E�4��聃
R;0�VB�"O���ï�36��cI�"vE���"O�a���N�n��X�eЛ,0@���"O��G�ϤUk���/�f��"O��3��q�x��U�)ҷ7!�d01�Ҕ�aZ�6R��+�+Y!�� B��ri-_qԴk7�C�{����C"O҄����r�0��  &����s"O�����6C�n��'�� [��KU"O�  f�I�==L`��Β>/�T��"O*����D�w����d`�2Eu�p��"OD$��&X_�(R �	$?VT�)�"O�eh���!
�4�3(٬Za6���"O%��,�(��I�$�� �C "O|y�4)�]P�3����#Q"O�yb�A+��`�b[ep�uBv"O�3�@R�Fl�����f|��B"O.���G��_f��ף\y�(�aR"OF	P��T[$�S����� "O��*5��B[�k!�80�|m�"O�=�4f !^��Xq`�)xd��	"O�I�u�29�f���m�N�K�"O��'CՄd{�볍S5F��J�"O��*I�O�t�Md��h	"O�-���Rn&����Հq��"OBg	�T�9��ʅtl xD"Od���H��F��0"H dq��:�"O� {���w<�@�)Z)�7"Ox�+v�F9Py��
FςW�f4��"O~��T���w�� #Λ�l� ���"O��h�˄�$	�m{!�07��{a"O��+��܂{��V+� L���W"O��`��6)�X�A�٧))�<�0"O0gG��M(L��
	�
�i�"O���G�XbK*u�0O�1���U"O���E��f���C.�=��uXf"O�x��E���a��,N0�@��u"O<=��,ܛ[�&5�P邺3���c"O|�A���X�D��R"�7�V�4"O>Aja$ȴf�ؐ�k}�@ ��"O@v��B��:a�8q�*'X!�0&~p��
;�����Z(+g!�F�H�М�#���.�8�J̼b�!�$K�K��pO2f�@9�c
f�!�C?f�,5��B`���7C�
�!�B�s$�2&�=۰�����9�!��� rC�(^n1�v�A�1n!��`���
Ӧ�7@N|D����.u_!�$׊Wﶜ�V�Z,A,! �mص
/!��^?<�Rm�	K�;r��-�!�+V<
�����k/8"rL�.!�d�	B�~��A��?)x���˞�!�DB�v����Z.���Ȟ!�3r�Dɑ���1$�����荎[�!��Q�.<����O��Nਵ落|�!���,�ZQ��G�~�fq�ve�AZ!���'�k-�:t��⤣�G>!�]�VO8tУ��(DL�b���G�!�DR�3(�U$-J7�]��`*[�!�ý�h\��/��Rr��,�!�J4#6� �wBX ,Ha-
�q|!�d��>0�#�CU�4,�f�pn!����'zf�A2.]']avPyB�2^!�$JO��v�L�>G1�E`�"�!�$C�7���� ڃ+�&��(a�!�S�(���dm�5R �ъ�
�Q�!�$��@�bFlǌ4�L�)�:i�!�$�-w�rx��߿^վ�s�Hź]m!�d�;d�Q(�Q�tQ�p(�(L�!��=�B�$!Ψl��y����a�!�� ��iV)
H,�8V(��T"O��@r&�	ٜQ1�g�'Fܸa��"O�t˱䘚P��r�_�P�ѳ�"Ov������+ų�$�Z���p�<祖�#4�d!�:>��1�p��i�<Y�CI	/*�\1S��m�$}!�|�<���҃'�1?��zH_B�<�ĩħd�RPA�á��`���{�<I�h�5C20U�g��+d��92�Yv�<YWl��MQH[��T1"��e���o�<iwCV(|F>pӷNV�2��h��mt�<q�@�QZ�s�Ѳ<�n�jp��W�<!EGMjUY�M��F�
�Xn�<�P+X�2~����0NpY��%	p�<�k�op"�1��)т�����c�<��=�	��HL�K/����c�`�<�Չ�@�BE;�h�S�ܡ�`��Z�<��h�7NF��X4j̗Tջ�kT�<�����s�&0�g��k�H�C���L�<���V� �n)��$�2yA�D��eF�'Hў�'+�*I���B�Mf�ib"�M,ҽ��P�:	��,��Ib����fʾb4r}�ȓ,�,Y"�*V�2n2d�0MľM�ܵ�ȓ�LU��	�`; �qc&��1���R���h�ABR6���Sq����m��߭.�NY*���0w�X}��4��𭊌hnV}6-Y�*KjE�ȓ\<�!��#�X�yAT+bg�$�ȓ^��!cJ�$$�Ҭ���*gH��J:�TH�3/� ����+a�N��ȓ	���cX���!J+�م�E� ��󦍨�h ���~�ąȓ/�T<��/�h�L���ȥ<9p(�ȓ:f�<�F߄L.�8�kܦ7�%��w���yՈX�l��|ص"��;X��ȓ0p<��[�����Bƥ^�\}��J-�Y�����&J8���I� ~ e��"%�Wd>+����J�P@����+�[T�÷
R�xqoݯm��ȓ!B�x[FHđW 0q&B�)�pP�ȓYY
qRV$u
0�A�7� =#���s�)�� >>Z���ҬO�,�;�5D��p��3w(�%��3#�<�UK2D���Ӆ�H��M�!��S�tب�f<D���*]�K���c7�Ҍ_,��G=��0|JVH�]IB�Z�B��JB�A�u�<##�o�4����T>P��0Nў"~�	�.� �;2�� �1ǵ!�B�ɷn�n�
�#��OQ�\(�d2 �B�ɛ!�����đ)'� ;�C��C�	�7Xj뗄LU�ܝ#�b��s��C�R<�Q��'v�d�q�jʥmF�C�#ZE�۰�q\�J��ǺB�C�,vɢ�s2�V:�J5�
��
C�	�=���5=���B�eƎ��B�eH�9��b.U���X"ٜr��C�I 7�X��
�~����PƮC�	�8X�A���r~��&���q��C�ɨD�7둖y��eɲŬ	��C�I�T��18�$�ZP����0B�	k�ٚ��k̄����C���B�I�$p��H�!W���uA��-��B�	��=�ì�1M��H0'���B����h:#b�7<�`	�ëO#z��B�)� hE'��!���#��W*Z��\��"O��	K�L����C��&6��"OF���/�4J��*֫N8qr�"Ot���l�*>�@�I��p��� "O��C`Œj3E)���V�B"O:-��O$m�s���(��"O<��R�Y�C봭Pw	 U�=ѐ"O�0d��7`vB5�'�M�d�R "O04Ă̮t�i��KL9Q Є��"O���b�>-�*}�qI$L�PYr"O�!���"-xp-��Cw�l|q6"O,q��&�&7V5���ފȈ�ӥ"Of�ӄ�[?�)��B�E�F`k�"O������Qۦt�C��Esz$s7"OH)L*-\�#4n��pF��zC"O�����6?���F�I�Q�Z"O�G�S�EbJ����^2H���"O*0`iM�o���j4럐[=���@"O�������$����h%�,@"O��6�ÕS�Q��J�G�Iؗ"O&����D���"у��_!Z�z�"OLX�L^�.���w�� 1����s"O*U8#J�l�T �.鶉�U"O&<!Q�ڷi��0�k �@�a�"O�\i��G�ޭS3*G?^��;4"OZ�P��5"l��.&��
�"O�(J���
w�$�$���i��ӥ"O��`⑖e��\����7ۨ8�F"Op<�Bހ9�(��0mW7%�&��'��z�њTz�T��aK����'vt��dI	�v����D�ƃ�4��' h�Ǩ��x�m��{A�y��'��,JT�j��ͰS���S��mY�>a����C�bm�DPAH'R@rDj��7 |!�d�%F�𑂆�ډA�D3'�5�!��;���¢ǘ�m|1c��I��!�d�w�3��mh�gS'}t�	d��h�U&S�;t|�p1���>��Շ)D���"��##Y�e�b����:я3D�Z���~K&i�#�YE����l2D�T����K�Ph�A$��x8�q�0D�H "��0t�X%���e�b<0�c0D�h�P
��_��P�@����[��,D���2�ʵ%��Ѓ3 �4D�� TK*D�lz*��Gr�asM��a�"(O�#=9�A�5�P, �`�Jň��`�<�E}8uSl��H����_�<	�E�Qn��'������X�<1����&M�Pa��E��!c`�V�<�g:�Ԭy1i# �vq��f�<��J�0m3�}�g,�W�x��`C[l�<A���C.����L9�j�\�<��흴>�.��@�C�{�@x�e��Q�<ѕ'W�>���
4�Ά�$� �[L�<���(f����1�Ƞ)5�Ѵ21!�D��m���î-�ȕp��N�=!�DA�{�t `s�;9(�))��^?�!�d[3�ܵ� �۝Q#��P�حr8!�l*8Ȑ�2Aꀑʱ�Y�7!�DL0��9S�$��R��1CVŃ%!�$�;f|<)��_�sx$X�s��")!򤁫B�, 9�!�rsV̳t���!�$E�|��xZ��Y�l��"O��Q`�ݡ*��lk�ثlRf��b"O� �����YM���#@=уS"O�i�q��:Yt�31�]�b��3F"O��Յ Na�s�߂���	"Oj(K�cK��j)��R�n�bY3"O
U�g��1k}�᫴^Ft�x�2"O E���35�&<�sB�FG*�v"O�x�VKL�U���Z��O4|WR�*s"O,�����U�ؘ��AU�<�z�"O����.8V!��|�n<�"O�UQ�Eܷ"d���޼(Ւ<h�"Ot�c����~�6� P�>�J�"O�K�f�sD29ql��nZH�c"OH��`g�h�V2�i)9� �4"O� b@�?]^vdd���t�U"O�-rH�x�1�ܒ	��D��"O�Qx��#_��9K]�~�^Dy�"O�T0'�ƜLP�
ЪZ*��e��"OٚTFO ���"p�@��"O^@Ф�	0p�r@���D&�]�"On�"/�:U��x �`*�Yk�"O�����6~"|�S�ʖln���'"O����֟w�DI�ժA��FMs�"O�I��P ؀��#N���x��"Op̫b�Cwr����	�Ji"O���ЩIk-lp�'�I�r��@"O�p{@�Y'Ne��¡�_5ld��B"O��ssIM,P�H�dO�6Mft|�""O`�b�N�
*2.)���v��P�b"O4!�RG����kҬ"�jDK'"O��Ӄ͞y�Bȳ<YyL+�"Obi ����iA�ʤ�y�F"O���?e#�<�@Ǫk��|8�"Ox�yF�Կ
��g�Q��W"Ot��d�S'�ҵ1�@<UY�x�"Ot\;���	BϲT�UM�/!H�(��"OP���'�%7���P��x= ]�B"O
X�`Ęa�U�V�ר_���"OX��Θ6cu���능cfHrg"O���0`Y	�XU���H�=�`Uٵ"OKӻ]r=�BꙆ>g^�HN���y� ��0���;/��԰�F��y䆃(� zQ�2R�@��]��y���0"�L��j��C"(�B�K�>�y�(�"�YC���<@X���P�˘�y�ϋ�PAX��$f1��-�T���y��zY���G�
�"UtAJ$�
�y��O,ҙ� ��[���"h��yd�R���Y�e
Wg�9������y��`ˈ��t#�W�t�q�Ҧ�y��ðz�&d�2j�M���('�yb�A�BPؘ��J�~}�7@�*�y��'|4��D�.,qf1G�Q�y!˱q3N�V隰����n�0�y2ʑ6$̀HEĭ	sJ�c���yr��=14�թ0��5��T�ā؜�y��!l�P0� ��-b
�iD����y
�4V��Ӈ�؁.m��Y5gӆ�yR%�d
L����:��b����y���5D��e�FBH|9X�r!ײ�y���:K�� ��q'�yse�X2�y"g�f����`�Q��5��&��yBG��qm.̈ƪJ
zN�ٓfV:�y���Fx��Y%ř t�\yÉ���y�'ͪEYJ�!g$�d�Єk&Ш�y
� �՚u�ۯ_��d�׫�"�x�"Otm{&dM�*@��x���+��X��"O\EsѥC08_x��RG�:{�7"O�|b�
'dP2钂G�J�d1e"O�d�4�-a̩h N�q�P�v"O8Lx��m�RD �,���X�@"O�u�SkI\ ��,�1����"ON�� ���"�%�{��L�e"O�p3TJڢc�n�2aeD3:�<��"O�E3Ȋ'Rvj2�ڵ�~z7"O6�j�BƭeR�u��I�.��d��"O@D��E�t��E���X5?Ղ�r@"OP���5?�>����T�X���BR"O�1˂ ��x�VL��HQ�H� Q"O��2)��B��c�';�B��"O��ab�Xe<1Q[�Xp	�k9!�D�y��< 0�G8d�@ �bֆkA!��	���*Δ*>ČE�5���Z!�T1*O��X�����xh;q�op!�d��EiL�2��E�=��}���Ҩ�!��|��P`KU
��5Cw�I�!�"S��ѷ+�=\��p��X�!�D�{������v`��t�+G!��B0�t1�*�!	1��Z���T,!�O�!3<B�i�6$�,\���'!�$P|ڜ� F�.��Չ��I/�!�d��R��pC��7�&��&�n�!��ʪѬ8! \2Glm�Ah���!�L5%��t0���dd<C�G��7!�9G�<P8�y+m����̗�(#!�䒒l�V۶�bʎl1�H�;;!�D��:�
a����N�T�8�+J)l8!�d�$���t̎F�����F"p)!��\�8�� �X
�|J�ʙ%6�!��Z�ȒZ�"����j!�!�$ۅ*8� ��B��P�VI���!��7H�Q��W�'n���S�8�!��5,q� Ӯ�	;YbŹ^�k!�O-�F� J�,p����eJ�n[!�$H3i9��X�A8|��p) CJ5*N!��n"�M
�l?yb����aM--^!����!I���sC�D3QK�D!�D$�&���Vg6`�jD�-7!�D�)���ѯ^0?��+��Ճ\�!�O�!���铌� ]%jP��-�=�!��U�GHބ���.$$H���A,0�!�$ٛ3Jx���W&�=Tc�I�!�+DD�1gk��	C�Z!���8�0��)T�~����ĎK^!�МP��ab�$HK�$A���dI!��_���9sF];1���(��D�r)!򄘪 >.�GU�d��yHd�Q 8)!�D�X�BMA�E�2=a��Ɇ��N!��U����Rn�� �")�o��!�(	�� �A�D�Hn�J����V�!��� #
�<"��>6��a[�0�!� R��C��"`��!��:��"P��s��a�1̍�R!�d�jx�Q�����n\�VK�5o4!�䗺�"e�U�9��vJ�y1!��R��F��@�
ejUpz!��+��  -V�[���z@	�di!�"�x��Z�t��8*
C&	O!�$�'7�
����2)�Y%)J0!�� D�Bp� �T�����*wr��b"OH-0F�؈d�ġ�"��7Bs�p �"OZp�� ä:&Z5K���qu"Ov1�M�/.t�xi��'��e�"O�qa��؆i��<"D�MЖ�8�"OtYH %��J�hDHv�N�XD"O��1�&V�PF>��lU1���"Oriɇ,�$d�X*암5+B��"O��AE��6o�E����-|�(�P"O�*%eY%`ՔAJU��9����"O�袦'\Ϭ���\7��a�V����I��j�@0���T6�#� C�MB�B�I%ut�:E��$c�@١&"��
J�B�I�P9hE�ԯV$�3C^�"E�B�I^���c�_$t8m��@'	�vB��>��4h��sa��F�
�I'D��� ߩ[�A��Ɔ�)���I#D��Y��4<�a�d�Y�)���qg� ړ�0|B�J�����+�~��+ �_e�<��o[�2������gIB!{�(�^�<��ĥVi>1����;kи��Oo!�$�g�0T���OF�R�B
�B�!�DK���2���*��r��Vd)!�d�Q��<�P�T-_�^(YQ�S�!!�D���i�2��Wɬ���΁7|�'�a|�N�%i�Q1�cZ:ah<�-���y��
S)F�`���^�v��! T�y��
w���t�^��ei!k�8�y��ې|�H�a�+�Q�:E�O�y�a��Kn(QhU�I�NT^! [>�yJ8@���c�K6NzH5k����ybH��`*���H�6f]���%�y��K(u�Z�;&��A<�EX��R8��?��A��o�=F����ֆ��z&�2	�'����h��|�.�i��"y����'������,-���b�b�%^ ���'MhՋ���ktP���Ì�G��Z�'Tlk���y��P�SB0z���P�'�#��

2�H���ځ)� �	���1O�y�뜟A�&L��f��4*�����'e���ix�I�\Y���8v!�$�2�z��䆜�w��$�S�΄D�!�D��m�4�y��X.p�Z\!4�ˁEA!�Q4'Y�Ԡf�<[�XD#t�Q:5!�ݮ���Kq.S�?�bѠEQ"O�)Ѡ�,¾8Z��.���9�"O�4����&4J4���	q��'C¥U$#��@�J��s	�H�&��Op�q����9��oG;rQ,K�"O�9��IԖ���A����37"O�U��2O�zD'�&,֬8e"O����H� x�Ĕ���$~��e*b"O��v�ְT�UA�4�<�F[��D{��iG�cg�h�Щݘp"���G܏�.�� �� 1�L-U�,T�G�

3�e*$�4D�zQNG"�:��֨
�>��q�3D���#AB�:_~��$�C1^a�w�0D�t���9j�3慜 u�J�˶�.D�02c&��Gi<PN\�V(����-D�H`a����%@]on��Ök�O��=E�4���+�P|�Fc���Ҍ�3$ !���	r,��e����D(N� ~!��P�0�-��-KSo�S%-L6!��"g�p�H�I�8�� JZ�a
�`��S�? 4�;��"b���C�NÜ`�"OĈ����$2��;�m��Ş�c"OΔ0�Eȼ2�(���.��tՐq�"Ohh��I�a�
E��Љ]��%�D�'d�Ξr������	�H(T�C��P�aV�If���q�ɻ�4Ä4���e@&D� Q�[/0�|ٺ��R=\T]C**D��z	�9	&ayD'�H�`$D���	�:�b�=6�p�"7D��a�02�\=��b��@�z�?D�� �L�pW�t�
�<�6X:�&=�&��|R�O<��Q,w��$i�)�C�"OD���]�8>�S�Y&<�Kf"O���3V0�5G�{�ީ
�"O<A��P�V�܁���5��8"O�m#Bg۠]��uR��ɔ%>�"O�ċ�#Q1x��\X�n�p��J��'���K<b��0;so�DҞ�[���0��O���1�g?1T#Ys�T�d�8��A���i�<1�$V)d�'k��ڜ�fM@q�<�2�a��@�))������i�<�)�.��B%	&;��� �L�<!qi֮z�PU{�LB#lkp�|�<A�整*Ғq��չR<|��F�c�<9@dہ.��l���\�R��\��p=QWl	l�8 �Ud��_� �;Gf�<�	��|u��������TkL�2Y���ȓe�hђ��U[���6B$=��'�0d)���h�H�&'�C�:L��\��l�r�Z{>����{�9��m'l �@��*K���ѫ�G�XM���f~�U9z|Ey1+Hn�Ԡ#hM����=13�.dl��Ѷ��.T%�FH>�yR��E�t���U�I(�h��%�yrޅ4L��4c	)X@=j�(	��yb�F>:J�O�=�XM@Ua�(�y@�!����e��/$%e%��y�-+� L0gZ'S�� �*֠��>A�O�A��њ7	�}� D�P�����[����ɗEDB�q�g�]�� 3Fǐ�i�B�	+J )A�KΈ# ��#�Y��`B�	2
��mi"%����8C���NB��'��7K<�$��b�-'�C䉼A\�mo�\s�����F��C�bV�"UL V��`��&R�B�	j�,�EI�'��;P���r��B�	}��$�ĿI&�1Р
�!^�pC䉾^��9w�QpL�G�.QTC�ɑW�`a1b���V�~hW��5,C�	;h�So*z�`������FaNB��,	{�$�#��?B�H�OX�:9BB��!�~lhpG���6d�5ZcHC�	p��[c铹��I��%�j/@C�� t� �2��>A�a�b �6p�C�	�b�0U2Ea��Aw���7+�3רC�I�R`X���*��l!��xx�C�	�!�w͚�[�����7�C�ɍ�� +C;n��X���� ]C�ɰz+F�
��V�j�Tt���40�B�I�z��m3Ê�"~�4a#���ml�B�I�B���ȢBi�(I��Vet�B䉢=3�p�ш]++�9��h��fB�I�nŊ鐵�x�9�"��v�PB�	U���ƛh��}��O�FB�)� �U�1��&a�P�k�k
t���9@"O@cd/NW��H�)�+M�*����'�ў"~��M��b�I��Ae�٥�G/��x�.l����!{w���0D��!�d$0<���7 i�׃�?�!��?�P;v�ǹ;L��ԃ-K�!�$�03�$`w�S*슐�`#�=�!�BMP�P��ú��`r 㜻3[!�DE�S�<�r���	;��(�bR~:�'�ў�>-@�+ջ7d@T���Ĭ:,8`��&�O��$��Z���$K�F�	Ï��%�:��0?1�#ЯJ�00y�G��"4z�Y�<i���N�u�M:P��%%�j�<A��I��
�' �F�Hd��~�<!�G�/%���2d�L�huxF��q�<�Pn�)QV\�Ae r԰�Sb�p�<��La�kG���&��`sV��dx���'
�=�	[u����m[�^���
�'�!���~����5@�Xɺ
�'{�Y"dĎ&J�~�²�F�%)�0��')2�1W��8�t��q���\B���'�1�o�I��I[���	z��E(O��=E�-جE���
Ƞ;^�S�C(��'��ONb>� �[e���u�T�d��ua-D�HS�H �VT���3<�9u˪<�
�O�.���@�f�jŘ��H$6�r���b|�*Uo��1~\ܱ��uH�ȓa�H�®�?>�Q'H��+$���M`�� �OW�vf&$h���9����ȓ#��� T/*z�hSv�+t�^d�'�ў�|�CKƒ�Z�:2���9~�ͻ`(�X�<qW�'9f�Ċ&���h�-�F��y�<	�n	v�4D1��2��L�K�y�<�E�ɰf���Ձ�L��,k3��k�<1�֏� �����[���`�q�<�#�W�+������4�1��H���䓀���kl_�zec�eޫdN*l0��'�!�Ą�|��@3�"YMj89Ԯ��!�D6i��l �*M�f�`��~�!�Ĉ�^� 0�f�4c��\�E�;:(!�P?��P2��IU�A5!�$غ2����W>-�L�I�F��{!���,#z��P�#$T��k�LC�`r!��ޙV��J0�Y3_��c�%:���)�'@n�Y��(�~��6k���Ax�'������t:��4e�z��d��'�<c��Q<B#���d$Ol��P�'J������%���.ڪ^�L���'���Ƞ�G�3�za�s�'W����'_���U͂
��lJ�.�2P����'�PYya�=*2@���ȎS����D"O��9V#Mf#v�:�	��:�&́�"O2E��(��1�.V�Ja&�@�"Ol-�5��(OVxb���C (�"O
��'F��y�nG�F(�c"O��è����sΞ7z�V͈D"O>���ېnb<hF'��-���#�"O���D[xZ�"u��?�d]�"OVp˲i�t�9y%B�R��0�$"O<؃��#�neb�#��+9n�sw"O�}��i�-�P�x���'3���"O�h*TC@9�UA�Q?}T��	�'Gfd0f�ܑ�I�UB:.�i�'fD���Mԋ�)8�@ݔ*HdZ��� T�H&�o���2� dsr"O�u��+͵.����^�^ p�W"O�9zaH&mz��ȁ"[ʔ�5"O����)�� [�	*S~�j4"O�����7��`IS�ʍ8; <��"O����lAM�f}�&+)�dr5"O@-Y#ā,���	ȩ���"O���I�8E-�	�Ch\�R�	x�"O���,?q��R�g�':��i�P"O&�23c�?n1"���d0N<<�"O$l�1+Ҙ[v�M���sB����"O�c�A/�b9 ��6=Ҍ��7"O@�[U,���-�G,j�6-��"O���v���(���j���;�X�4"O:�y�!�� �rD��搊9�<��"O��@M �.ܢg%��x�h�:a"O����J\2\��kC�;(��d�"Oz@{I;|�=��>w�<[�"O�\�da�,@*�˔�ɍC�CR"O�44��.1.�2l��DI]qw"Oڼ�cִ �!�5O1_�d|�T"On����Nab����������w"O��HGٱ]P9��ʍ>��	�w"OXxbađ�l�*ܘ���a�}[�"O��[� k��Y�D���a�dA"O�;��	�\�j�'�?�~���"OF�ѓ)W."5��L`�\��"O��V��E��	j���^�� C�"O�V.0�0�4�V�B㋕l�
ņ��
�{���F}�a�[�Y���ȓql(��#)�8�BՃ�~}�ąȓ5��8�C�	�P=��%��;P`��p������2�~���.R�wSRU�ȓ`7Zm�Vkۍx�l�kV]J�ԆȓX��hqPn�%�VQ��D .w���ȓl�R��gA��'xݚ��Y |����ȓ<.*}{���,�v��	޳
g���ȓF,�B ѳF�L�t�Kc�j���t�6���H&>m�4���Ń=��0�������2�j���`�>[�0�ȓ 4�PC �}~@ț7��~�l-��/�f��DAΝC|P��s �(y;�	��b��1I �M���+�޻;��ȓe m����0P�,�ӤU9�z�ȓ~h�%ء�3; �c��-�XD��Z�$Z ܆N� ���$d�d��Ą�����$b�\�r.Ԗ����ȓ4d�r���%
X�Pp��K��1�ȓ!��AZb�L�c4�E�d/�
L5���ȓ��l)`��y�<�:pcW��(͇�1�\ј�Aژ]�Ɂ��TZA�%�ȓj�;E�(�d�	�D\.wڕ��Zh��hqm��TQ8���ee�e%�B�<�%!�"1|(�gkZ�Rdd�X�"�e�<iV@��6YF�A��A�6<r�)��Wb�<�u.ӗd��!(Gm�!X�3��	b�<1�ϙ~<��I�9,�*�ti�[�<a5Kq�4ᱪ�N���AU�<�5fA�4�ԔZϙ����J�Q�<��ᎏ����c��x�`�r��X�<���P�fdj`g�(&�ye�l�<�$d�c�:q��"C={������i�<�d�ҹ`��9K��#�N�d�<�� ��I�<�`	F�+v*�C�E_�<� &��`n��8v����:�"OZ���A�]�¸���9K���F"O��[P+*�0"�\^��!�"O�]I&%BMMt)�cNG���"O����NHł����)�ʈ(�"O��sG��D�b���eu���"O8!&��;��D�d!�2Z\TA3"O�\wJ�YPPy3�W�-I.��t"O�$�"�	L�$��<C2�!�"O��#2�?'Bi�e� �=���	�"O4x��Θ7g�L�-M�}ܥ	�"Op�aR��-g��8�6�F-u�"O���"���0�7��=`z�f"O<�+ԯ!��P��߈`D��"Od�	u��<}c��R�sG �Yp"O�����>tr�Qj�����k�"O���.�:! ԋ���nph� B"O�ypb��⡩�⍯��@I`"O�4��p���Ñ�|�fe��"O8mYu܇);�Mx 4�Ld�"O�Ԁ��͔|H ʎx�^��"O|Hz�F���ɳ񋒱w�Ȉ�"O |K����@��h&�X�i|�E�"On� ҡ�/aPd��I#
��Y��"O�A�p�G� �� �Ŀ+�T��"O�p b�d�ޠ� �T�6m��%"O�t�AHX�e��|�.O�l����"O�|�ˀ�#��C��ORhDQ�"O��#�ܩR<9�̜��T5x�"O��'	�w2Б9�mF�o�@Y�"O��q���=��4��
��
&"O4�B��׋I��r�@�ײ� �"O���g���tI���q͔�kA"O�l���/g�5(�$C�O"�sS"O��y��@���ٺ��O�~* h�"O��0ܶ�"��P���t��͚"Of;��" ,BE�̔6Jw$ɴ"O���p?�$�ϺGc2m�w"O,���_><���JFP?+%"O"Kt"\�=�����Bd&X��S"O2h��Նr	Tr@�̨LF�`r�"O L��!.M�0��4���?!���"O.Ԣ�[�l�di�î)
XS�"O�a�@ #yE��V[�j�]�C"O��ԠR"3����쒵(�vA��"O�ف���>Q<֠St�h�P<8�"O���ah[�Q8�-[C�6K���"O"��fm�%S!Z�@
��2��� "O(�%B�_lT��L�NHR�"O�m���)М���/�W8�r�"O��j��D�V�Ԩ����9$�22"O���25�Z-�T��hXݪ�"ON���G90Kr\�B�:i_,|C�"OX@� �3b���3�-BWfhB�"Oj	��Ő�Z�L��숞o�pH�"O�qӃ$ԑ9u2	pD��7�ndp�"OL�p�� ���9��~��0)�"O"iu�ߡ*��`�eO}�� s�"O��Q���/!���q�2h��]Y�"O@���T1<j¥��CG����[s"O�0ì޹mxܽh#l�;r>Բ�"OԽ2�]'_pVhi
�8Xҥq�"O> бH�>���#��wB�i�"O֙� ���
��XR��Z.`.X��1"O� ��+�톪#;F��O�/�B�s"OJu��G�;u?�Ī�M*4�ް��"O,��v���1�v1˲̅�&Ĩ�'"O��!Ƨ�;�� �0xd�a�:D�,�g��^�J�a��$4CN�Ru=D� ᣉ�|��۶	U�?vz�˧;D�X�!O	dT�0<�}��9D��`gO	3w<���DLu��9D��(A��2!Q�-�U��wg�X�`4D��D�ۛ ��j����l��l�p�&D��iE�/5���:"�]��h��eG'D���Qm�XgVp��#H�����'D���`��t-�i�'�x�$5�c�'D�Pvn��j}�����1D� �@��$D���G im�����/"���Vj=D���ƀ��=$���U�_��4I�<D����7�����Ϣ4�Թs�j<D�<�i��i*�	N�����w�;D�ę$D'� ��"#�<�n�B�;D�����A�-� @!g��#�F��W&;D��"�$I:kR�3���$F��s2�8D��KF��+bZ��mGY
pg�7D�h �]�{����D����c l�<I�Q�:8�!@oՁ['⨡�	�i�<ar#߱|���H���R[��ۦB�_�<qr�M{W��E��<j+0Lc�ƞC�<11�MXN��v�]�J�8�H~�<4H��6���[j�c���h4H{�<�f�ʄO�����;��谦�~�<�r�V7}�~��扌��Y BM�P�< �"6t-iD+��/�~	`���L�<YPʟ��T��-�$P	 ����S�<�gL��;����ٝ#бs��OK�<ApnH4"�B5�����")WK�<�E��>}`6�Qjܘ@ Zm���D�<9�G�p�i{���m�"$BG%D�<q�/H<p�,LdD����������8��2�(q���ecX�ȓc�L9���=M�`HcEg��^���=�h{Ҍ��7�1�ӆ2H�q�ȓ%<j�c�$,~��n /���ȓ~�Ƭ�a����:��Cz���}�t�ru�(]� �J2�ќi �"�4�{��	������^r��ȓn�:���C^p�)�IUlN@i�ȓ`�y�G��.D��H�ٍc�̰�ȓ1D��(�f��D�p�	
:y��S���R��֕QV1(�[�~���2Q���U�XFȄ)׹��B��?D�t0gj�9��e��;8lޜp>D����f��WC 
T�:��Љ�
?D����R�5���e�N��D� >D�ġ節<z��cށFN
��<D����o�Jc&H)mx�E�C9D��@��RU8�J��=TL��I�"D���Fa�0Ҧ���%ސ��5k?D��ʰ�Ɗ9Fl, b��l=���;D�pJ�� 1B)"�+P���3��2�/D���aͨCvE���N&o��t8	-D�@i�_!}���cdL�r���J�B D� :�#J$��|)� 	6p�j�2/>D��U���_JH�� d�2x��=D�h�&�9U������E�w��4.:D�di�E\:l�q	��C�4�=0�)7D�� Ȉ�!"�������,&��L��"O��#aF׽l P�w!�B��K4"O.�YĎ��9E��q!�?��;`"O�� �~"H�r/15��X�3"O a�)�l~[w�ώ9�6�pu"O	�5ʞIn��i�L�1��)��"O�����T�Y�Θ������"O|���F	 HK�Q�M��x��)2�"O�dےI�(��܋�gƶ�d� "O�iԀ�6S�b=@��	0-�Th�"O���鉢R�\J�D>|�a	�"OD��&l�+:�)BE�0r䑱�"O�� F8x����ȧ
��h�"O�8�w��4�D9z��G#/=�p�"O�ZU��?/���R��@�m2��JV"O�98�Y� �\U��&BL!���"Or<1��ڃd'f)b��ܺg��I2"OpL@�H&?�HL���;��eڣ"OXI��)Q�F�L�0��.m�F��5"Or�I3�ڎNLfu`�+Ԗ3�`�@"O�T�,;�0��%س&<P��"O,5�V�Ϩ���+œid�H�"O�(z��N6kn�D�G��
���'"OD�R�ھ�蔒tB����sB"Op��ƦK|�D3�'��2"Oh��S#�0����I�'a~AZ�"O���V���LWL)@`JG>��� "O�I0�A˂O�2ղ�kC,�Ad"OPy�i� � i"��AxBؠ�"O�a������쪃�`Xr� "O�Q�"�ĆYvQ�"�˘rI��Q"O�\�e>n��v`�![v��"O�%yd���}�(y:3���mS���"O:����Qx�(�"��A8�0t"O�}�e�Y&%� h���g�h��"O�Th����H:��Ȥ��/�أ�"O҉���(5�r���[�\|n�
�"O�0«R
q���3���PvP��"O}ہH��L�.��V<�.-�"O���CO�H�d*������� "O��Z���=d�.49�E�A��"O�|��G��	�A��U�M#"Q�p"O>�3B�C=5,��@rCМd�D-p"O�ܱ�o׆I�DPF#I�P4p"Oj�s�X�KU�b#F��d��%"O�EC僑�+(Y)��3���"O�Y���+ׄ>���� ,�V`!�ֳ
X�ȲƏ[+d���
�E�(wn!�&��Ű'I' fBG.ĚR[!�N|#����,��Q�������<�!��m�FXQ�5)����er|!�$;}V*���l��Q/�/c!�$D���)� Á;3Ѩ�ct-�J!�$�w�P��	rb�yQD��d*!�$Y>=�$��pJ��iY -	�bF"]�!�d#S���E��,Xs@1b�'N�.�!�>[N��Ы�]�(�Ɵ.A�!��҇j��(:�ʣ:$j(���Bb�!�$_+�VY*�̆�BC�@�1�]��!��ڥ��`��Ast�ȗ_αz�'rQ�Dɶ;�HP�
��T��'C,�ϗ&�J�S��B�'�EH�"�2Lp�A�Q�<a@�'�4\��o��y�R�j�	�Q��)��� ���u`�]�"��ф<�0Li"O d󇈑+m3, Pg#N�ph�#�"O�y�v
�1��á��3`F ��"Op�����b��T�ƌ7�ҙ	�"O��s�KV�������OTA"Ot 3�I�<��U���ظ_mR�yp"O��c� �8��=�V#�3��h�"O<<�TK�h�����@g@���"Oz���I�i;��qՖj1�P��"OiR"��3.eh��,�K$f�Sb"Olu�S����������h�"O~3���$�� 4ᒀol�Di&"Oj�;Ҩ�$X*�D���&_���"OPl��'Ρyo�d1���	c��b"O4)C%�oH�����`�"O�p�S�n��l�Q�Ý |H]�Q"O( �u���B���A�I�{l��k7"O�@�O "'�0qUb�c���"O��ㆵ8�8
�M�)NzQ3�"OR䂁�]�v�$Ӡm�	f�BY�w"O>l��h�3g��4L�	[��H�W"OdU�2�
'���p3�?T�`4� "Ob�6�7��H9P@�0��1&"O����ŉ�piB	Cျ�$�W"O����NʓD��	�W�g�P���"O�u� ^ B�J��0����5�"O�IWΏ�����u�Qby���"O*����G�ؼS�@��R�ܙq"O�ih���� !Ι��EX2>])A"OL��K8	�zԘ���|��A�"O&ɱ���=O� �7��7�H4��'���rW"�4dy^��`a֒X�����'� L�0���H����X�6���'HfXk@G$8�`p�ζWᶰ*�'j��(�	j�a�X_{�=�'��C�MG�%��| �,7W�R$��'�*a���
wB��ʈ [K�� �'�
Tr�G�R��� ЫLw\�*�'f�q�CS�~�
����OV�pl��'
.�@��J�4�x1��5T�:Ř�'`:}!�(C)0c�A�:#��-	�'�N�����UOąy��%�� �	�'�$���BO���Q���q�Lё�'�n���;1<"�y�(B�b�ua�':�Dp5	-8n)(��b��h�
�'�� �c�h�̋��.X�&!��'8�H��W�*=��;ԣW$��@��'��]���P>�h�`ۢߤ���'^���n�T�8d���R$�by��'PP�ჩ��V|��i���|��'����͊?::��VbO0	��'�6�C�L�~��d:���(X_��Y�'M��@LC�K.�[��Q��U�
�'ΦU�P�I�z�� �b��BE��S�'��c���:�����$F�栳�'i���ef[�kʔS��1>S>�S�'�FL�r�Q#��@A�6�`L!�'p�0q$�GiZ�}��) �%z@ls�'d�උ�"����k-��)
�'��ȣ�)��Wh���7�����'�d��Hs�@�q#���`E���'P>���<p� 3Sl�)����'�4H)!];~t��`�W4(Z� �'[��H3$N�,��JvG��&������ \�J���1�Hcs��F2
H{P"O$�s��ڳ*6�ՁU�=8|��"O�ĉ��z�<�ö%́2_zl�"O���C�( ˰���.��9� ��"OJ���I
� ��v.	� ���c�"O`��g#M�?�؀{�̪�0x!c"Op�w)�w7����jS�Kf\��W"O���I�:E@��	�OČ b"O�I�'|���0�V�R�Nk�"OFa8F� 'xXX}ȢAV��px�"O$Y����9
8x���{��93f"O
�)�ERr�y#V ��*�Y�"O�����r�x�kDj,�L"O� ۶=�()��ޣu�
-K�"O�<2%�ڵ3/���G�<MZ���"OT��a��n]��ǑF�J�"O�p��EϮT`v�9gV8]���#"OH� � */�f͡S@M	�Z�`"O����&��%�� �u��B�2��V"O�,YTMK\���Ţ�"h�p�b"OHL:��X\��PdA.��0�T"O¹¤ 
*�|a���#6}�"5"O^�Аi.q��q�?+̦T��"O�E��DѵHsv��N��D@��"O�Ғ&
%1T�8� �=J���Y�"O$$�3�IEq�ՑÎµc��M�"Oz� ��Ie0��� n��~>���"O
�����	��%��"|4���XX�<Aa�	�.�A�!	Ok���K!`�y�<!l�`����$�A�Lr� �`�t�<�d�C����)-J�0 P�hPU�<���K� �9��?
����ck�Q�<	��.tͰu�B�R�3�"q�q�P�<�P^ϐ�s���:X��G�L�<	p/�4n�� �k��YYd�r�O�<I$�½&cpt?�*���K�<Y��H9�*�5�N�=�Jł���a�<I�C�ZH�`0�J�҃G�g�<�Vd�0{�R(�W�ų3��X�%#�\�<!�Dʹ7ze��L�	�%����T�<��¹,ȁ�UI�U1���3�P�<0��c_��[3l�	
ƅ�&��E�<!AnR�h��9%&����� 
L�<A�h�	5��Z�ā#,Z渱jBo�<��E�Y��@�%�88��qG�i�<᧌ۀI$B�3��5K����PTc�<�$�&v4�	��%L�?Z�9� k�<A�L�#P۱�үE{��d�<	3g�=�P�'�0"R H�N=T���OV�&C8Q�a�հ����+D�t�B��D�����ҲJ��;f�(D�HK��X�;�-;�E�?r�Ȣ�%D�X+��{���/��^44t�'K9D��Eʛ�Q@R95$̚uF�d;�8D��9@bؗ6�
��a\)y.���f�2D�HЗ��S�8���ƈ:�x��,/D�Xjn�Z�����F�&c��kf�,D�R@��F��I�'�Uo���� ,D�p�qb��3��=�h�'3	p,8��>D��0()�r0���]�e0�vn'D��W.��`��p�0P#���f%:D��$D������2;�� �5D� A�X�0����R����I���4D������N�w���_^l��=D�� (	�$a��P�i]�TH��"Oxk�l:Y�t$��[�r8C�"O�����	J������E1�"OV4y`b�@�h��F
�p�r�"O����kD�PC���-h���a"O��b��� d}6�U�[��,rT"O�	1s
�)9����d��%��k0"OX�1f�/G��YW�٨nl��p�"O�y�O���b�Y�0=����"O0]�&�ѐu,��rg��I6V��"O,�H�E/�*5p���;GN)PV"O2��`���q>8yXg��,p,��C�"O���H�"�jqj�O�H�(�$"O���e�<[^�t�M�i��I""O�iS��)�Q�Ǚ|p��"O4�k�
'!bx���.^2���"O��Z��^7�����W&XF���"Ol�&/������҆	�j���"On<��Ig��D�B$����6$�x�<�5�H�c�ٱ�eB5�((ICʖo�<Y��тq�.$�p�W4Yu�	���s�<a�(W<bR6��&�聠5�Al�<q�  �z�v����tx@b��k�<����:mRd�*D�Z�X� ���~�<1ti@�f(��{}�� L�w�<�C�� M��EY�m־R�l1{`��v�<��)�5R<p���נK��t˲ _g�<��L
{~������H��R'a�<ɇ��.e+$��Bl��a�b��B�U�<�* @����⯗#�r��$ �G�<p�ʄc>�u�2H�6C�����A�<�&�F(���Zq�ؑoh���m�t�<����>�1��k�|1�lyr��s�<�4�@
���#�C� \|�k�W�<�2'N�g����m��q8�Zr�Fk�<���ҡ�4䙁A}���	�e�<qq���s}ʈ�4D�l�0� �GM�<Q3'�Tp<0�]�M���yG��E�<9�ƕ�6Ҟ�k�2�F4�T��V�<���T]��q1�gQ�y���2�AG�<	���o��z c_"�)a3���<a�ł�&�\asc��V�AH&j]a�<��gA,О9ʒ�I!G����e_�<�s冩Iȴ���W�K��㓣q�<�W�Ŝ��@X�����zU�G�<y�N�^�|�`��^<K�X&�h�<��됣u?ƥ��L�4n�B�Ko�<qӋ��\Af��N)���" �i�<��(A�)2��e�[�n�r�![b�<a�'�@�=���P%?����f�v�<���.tS���w��!&�Ft�V�v�<yT��	1-�����\{�|Ӱ �r�<q#���H�� pA��]X���Cl�<Q�����m�&f�8]����Эf�<ɱ�\�yvl9i1-��ݸFE�{�<9@>796�b�eG.T����C�P�<�0��mm�؋R`Q�PJ$2s�KV�<���݉+�t}��D�'�:@Z�h�N�<��Q�*[BE�%�3	j@����e�<�����!�G;�v98��G�<�!�ӆJ�T-6��66+�Eà`�Z�<P���`�,�P��I�j��Ms�-R�<�t��
��2�&űc-�9�sOH�<Ae��l�4�g�-~��a�(EB�<� ��6
�D�@�C5j�\AbQ"O�[��_�m��A���!��]��"O(ŀ��I�v�f��QBN<�J̚"O��x0�C�fDN��gˇZ��P�G"OHMK&GG�N���S(>	�+R"O�J2!ڈ+���YǏ��i4SQ"O�
R��9%|`��P�S�����f"ONLc��df]I�fޙ>���"O�
�YQ��1f�n&dL26"Ol�%�S�DMI�e^�ڼ��"O�hR�'�Z�I 䡜�r(�ԩ1"O���$�;6�@!CA�74\�A6"O���CƜ4A� S�� {Y����"O�ɫC^3N��h���&?���"O�R$��t��i@ �(,H����"Oz���h�C��T `�ϥ�L���"ON���H�`�'�H�i�ء�"O����	W�Q2P����.[P��B"Oܰ׮��m�);/ �=b�"O,0`��I/qtxYb(�_'�H�0"O��*D	�)V*ԀA�A���9V"O�5�4$J)�t���#��)i^�h�"O$9##%���hѢ$w]��x"O���fG����e����&jF>I��'Y���}x0���of`I�	�'w��A� �("�0�E
�f��Z	�'�|��a�(�<��'i�1�� �ȓ�nQ:���<����cf�9uB�l�ȓG_~����Ҷ(�傰f�7�8��|��$���Y` ��elZ�i�b��ȓ
nN��l�"��B�`� g���ȓI�
�e
<d)��ۣ���G�n���H�����
���"C�>���ȓG����ͣD���P�i�
����ȓ0� �r�(>v,	�*U�̕��q�f�V&@���A�"7#6Ї�Py04�@Gڝa�)�f�[	pGbхȓ.�l`�'K̗G����≞9"�,�ȓ>U"���<RH�d��f�:����m�SNV`4~�h�/�{ �t���,�����vRD`pWlFݤхȓ0��a��BۘL(��C&ɡT��D�ȓo"����I�6�B�K�O@nt^��V,��� �/{�. ��'D\��Ʌ���X�B�ֵ��5��b\�`*P��sd�X��ʕ#!��12�<J$@��݊Q��L�1��ȹ�Ҹ<�8���N:����ɨ+p��E��:GV݇�g�����(�`����8T�����$��� Z�]^]�UC64���ȓ=��𫐂7T#\u)RK�2Z:��ȓ\D���$
w8�h��6O~\D�ȓ�:����v(p��b�4+�"���N���+�5a�p��C�3!�hU�ȓH��ЃA�L�*�.�0�산V�$�ȓ$�96�?e�d��N�CX�1�ȓ-疘����G�L ��W�'�\��_����5�Ewn����+G��伅ȓ�JXf���p�T�Ä��Y�`d�ȓ2��4���b=�FD"DɄȓW�FI�Ł1GC�����e��`��Ez�d��'��kgf�˵��:H 4��$�=���ʟo�洐�eї9��Ň�r���Lߝwb��Q��.�(���S�? �i��*��R�J����-��Qy�"O�lɧ,���D�}����"O��P���2lJ����2����"O�yR&k�>?�{�!�-H���W��/LOʥiAdϒA��Q�@%&{�@��"O�l�Ӏ�9h��R�0(�,)4�$0VCՌ)�M�]��)!��>����ڿ��'�^ QHF8v2La��c���4(��'@б�R�}/�ɹra�*{�H�cM<I�O�����.@��HB�A�AE�M�")H's�!�dT���D�iM:Ҁ��!-�F)��8�DIzp�O�Zd�Rr͍�k����O�r��uPKL�Yfp,a���B?�Ls�'�0TX�aY�~^�4� '@�f;��ҍ��)�4�VW6�%�&��zA&� Ƨ�=�y"知@�4y�*@l���ؕ����hO&���+Vfla���"��h��޳_�!�[-^H�DE�;�Z����\7n�!�D��8���oߩVyN�����J�ȓ:3\} ��;u�t�Y"/�+H5�ȓ+B8�#���_��� �$h,Լ��R�D�*���~��]�T��}�T��L�/EUT��W�܀��(��hO?KDb��v=s�
k��= �o/D�h�IV�7�h�(E�U��Q��g.D���T�>o ��+��cSc94�軣/��s���b��J��ȕx�<i�-.�}�2l^c���1GVj��q���O��ր�5b`Na�%X�HE��'el0 �cA�z&�+��7tU6u�4/��'��I}�'�����	�1a��+�`pa��'�����M�yK���I�ʥ)��.D�HЉ���h:3�O�_$�� �9�ɚ�HO�O�z ��[�ʮ��6n�/����
�'� i��A�n�q0���.!�M0���<A���3T��1�j�7c�I�#փ5�!�ԍf��T̑�y��t�у�-y�!򄊷@��<(�ǒ91����<,!�OJ((��ICI��ek=n	��Bx��C>��8�2��#;��Ja D���G��v��(�p�i�Di� ?D��aצ��)^L��@�Ը_>x*�8D�\C�T��M��+�3j��TK  6D��
�)C.)XL4��ӉR6�@�uG5D���'� ϲ�H`iPW^�� �3D�ٕ)�=m��iA��(O�����ǯ<
�fS�Q��,n��$H�Tu��!���D~E��;�C���:ul��Вe]'�y��÷%t�İ@Qn(2t�WV�y�J�A������.4�@͹!Y��y�g�[6��R$@I��&�A�yR�)��O?�o*��ea��Y�Z��=w�I�<�C͝�w����]�A�>�0QMB���d&�S�g�w���U{8����
	|�&��AOP�u�0�keB\.(� p':?�����'��O ��m�^̔D��J
,4����|b�|��kV�)����<�N�sj7b�˓�0?���5 �v푲�� <Q,���f�'ޢ<1�Q>��劖����1.�O=���1D���`mG �2��@늾|S�=UbN� ��O ���i����я*m"l#�D�a{��d��r����N5]�R�J����~�!�Z�#fA�A�V�F �+��\�!��
\�M�OٞJ��%�l��5�!�� 8x�d�08�����m�[���#��'Zў|4ę!|n8F"��s>)�a�,D����N��i��`	�'�
Rxq�e7ʓ�hO��>J�4�)@�,`��/�J��d!?�qfG e��Y"��R=�ֱ��ڦ�	�'�qO?7�V�2�Z���0l¢����2OўȄ�S9�~x("G��L٘e�@c�?�LʓF��}��=[���@HVO��)�J��HO���	*�X�[����H��(�?u!�䞟�Z����A�k��"C샌a�!���(#^�A�s
��T��hr�kS�!�$��w�į�h��Ͱ F%P�!��
�,�Z�Nτ������$e��D{��0ɓu��\Ȉ�f�[��azg"O4���̣8�|�El]�Zf�t�iў"~n��VD|)�M��ke���bO�.�C�	�U4�S0��"^�z(X�G�%����HO�>��!�J����(�[~��j��>D�H0􁘒���&ƞo�U��O����'��h��"����k�
�`'��"��;D�$�����f�򢃃�W���ɴ�3D��ksk�h����ނq-t��2T�z�c�D�BP/�8V��L 7"Ohl�G�+��(1A@�8�DpR�"O�	2��%0����e�5 �f��"O�L��C��P ©�v��>|4�"O�a���DVf��׬��;V��kT"O�	�dlʕK�\0��lW,J=��"O�=�r�G!N�D� u,<��6"O���T�����U�"t'�EZf"O����f&v�d�J���������	G-HAr�E�
Y���@�&f���v������v�K +�ԛ�gS8q������<�S��yi�+���E/?,�Da�$��$7�O"�t�Z�'>NX����!��òi���$M�a�6�����*"x�}#�灄^�!�D��)N��ۧK(WF)� �ax��I�7����ܺ��3`�Z�h�z��p?1�&�N~!��$�d����Tml~��)§e͘h��Ȟb�8TO�J����ȓN>�BWM]�@F6�CWG߻H��9'�؇�ɉ^����矮Y��y��Nͺp����	k�I5-_<H
׬I�T4�P!Ƶr��������K�24np�5o��e ���d� g�!�d_-?v	s�[�\鎨�cdV�N!��A����5����\dj��U !񤜪$J	��O�G3��c.�X����o��9"gc::��	�k��zmЄȓ����S�4Iw��<i��,�ȓk�A�d��,Y��e1�̑85� �'�@���A��|&�d�G*�I��ړHǾ���Q//$�pK��ʺD�p�	O@�a�Z=�g;��'��{BI^'c���f��%=x����5�yB���1ж�i�/�=nİ F!�DO�~' �'.��~!�	vN�� 1qOF(�뉝+t��q�!��l`B �6P�[��C��:,-�R�N��>��"��1@X�"O�#A5W
Y����]rt��"OP4��←7�P�%��3n���"O�����]f��#�"R"PH�"O��`!��y����.gK��ha"O� ��n7\����\mAj=�"O�q���1X�亴�8)��i	�"O��'�*����� |����P"O� ������?~ƹ�q ]:�ܑ"O��RE�If�~�����;�ޥA�"O�Yj��_�DRC�	t|�aB�"O�E�"t�HC$�l�<1w"O�	�u/0(<EA��h�Y��"O�5x�"�(a�x�q"�	�J�%j�"O���Gw�Heq�hǎ%�����"O�MI��W��,	��ا	�
��"O�0�. _�L���֍S�����"O`+�e7-�^�j�!�5;lزW"Of�k1�]A�:(Xs�� b�ԁ""O�$q`ؙB�P����EU~XXW"OB�x1d4+�u;�>nKbl��"O�����	�ă�fU�.ZUj�"Oz �%�̲"lF�@�eł45���"O�Xp��On�7�O�,���+�"O.�2��*h��<�6�[�'m�i�r"OH��эT�.a��Ŏ�u�2�J7"OЁ��!N ��(��d�Z���k�"O.�`r�38��	*�_�h���"OfD��GB�-�n�3��</w�!yD"Or��B�:s �rV	88�k�"OB�@���Ǯi��Ҍo#��6"O�槝�;ܽK�F�ə�"O IBTޕ|�2��'���J �l��"O���!��E�>mkd�1���P"O2�b�O0F;0��-����D"Oz$���%Zi���QI��E�"O��[��p��(��"T��]R�"O��TL�X����0#�K�PS�"O©��BC�p�Q�B9]��d*O�t�Ƭׯ'M�H��Μ#Z�M��'�r �o)7�*	����wsڨb�'b��"%�QHrax ��\��q{	�'�"l��TBL��L� S��r	�'���y�n�6R4~��t@m$���'͂t�@C�b��]�R)�5k"��'Ī�G��7�l�3��4�����'j$�(��))kd�1�J�YN��:�'�}"r�Q�M��(rs,Ҹ*��e�
�'MB�k钍%�L9e�<8�9Y
�'��c�B�n:8��V	��a
�'�ɪ��-i(Ⅎ�*!�� R�'͈�P��"<�����L8��'	r=�Gn����i�Yc�TZ�'�,Y�`���nDJ��]�4J�'�d1;P�.���7$�
O���z�'W��H��HH䑑�._�9��T��'֬q V@Ϯ|À�!���+30�'pr�c@DL1@��ظPH�]�|P;�'��H�fΧ�⧤9X���a�'��I�5�۽�D)WkC\w��s	�'� ���P�'��|0d��d�"d��'�dU�dG�:7BѻB`Jfgn��'#B<X���%Q!��V�� �Ȃ�'�xh���5�����:6�%��'�&]P�� L�pJ�)�16�)Z�'�nܢ�Oܷt�V���5/���'�2@������p���#}(�[	�',�������(	�CE:��S�' U˦a��<�U8�b�WKVı�'���Te��YQ�NF�I����D�A#�JNI��DH�>�5�ȓhi޽�qΗ�t��A���D�\�t��S�? ��cg\�,��t��(�P���@g"Ob�h�J³^w�tJ��/`�����O`�x��'P@�(��dg�(0��)�ə	�'�j}��K$M�84!�۸1d����$L�,�>���<�S�rj���vG�aW�MzׇR�!ChB�Ɍ*X��G��xi�BJҬi�t�<>hP���P�dӧH�jeQ($�� �i۽�N���"O��BaF�M��hǧ��T�py��+}�ς����#��D\تa�C��"Df����� a��@�
������J���a��ǿ__� iuc�;e��i���":��LaQ���;�*�B�MqlF#?�'���l{�9�.���j��|yAf&�F�8�o�<v�!�DJ�CZ��IV��za�a�����2x`\�k�ɺw��S�O��x2��14EP���ɑv��m��'1 uy1��)J�%ɲ��$`�`L�6�>YҥSLʈ���}2N�:^�89 o��/XȱE�֙ܰ?1���,s�uB&`�_��1#��>S�Ĩ��ئf ���d��`��`<4�����(D�
�џ�#I�Z����|���Q1��rw��DNG�A	�Ņȓe���n�\�U�B�L�=����'���6��Y�S�O�&�A6���޵)�L2>IDe�
�'+��G���r�6����A94J����'g\����Z�ze����6r!��'i�c� �I��a�2�B�t��e��'���Ѱ@��1�¤[�$݊ț�'��M�e$�3L&�"R�]8v�:�S	�'�p�g�;Ʊ�� N�)$���']�}����J,�A1��E�s
�'��E��O�
�^��0	԰�(��	�'�~9��fQX�����l���TX�'�z1�v͝!E��0g��}�����ņ<�؅�
# �K�W��S��:3�X)EZV�l!�`
��OK��)�&	��������	�'����c\�>�2�HV�n<l=�O8�q��31x�'i���!�_�OO�q�@M�"�$a���u� �c�'i��2dF8CGL�1GXjm|�h��i�ȀW�H�b6�,��팭�O�h�QN<)�L	�'BL���yY!4L�|؟ �'��(�B ��kG�	��:�O+6V�ij'lőN��bbª~F��f�+@D�"���OR��Q7=-�LJ~�Ԁ�-� m��+�P6�H��/UD�<�V�s�d]��IƏ9�84K�B�G}K�J>f�Y��j��S"C���s�녽m92�&�)�<C�-���PD	
�<|�`��4l�ѦOFiȒ��+lи&>c�H;�0f|d��h(�s�"�O�X���sǎ@q�ƴr�ft�㡍4T�` L����?�q�X�9X|�#׃[>+����ME�'��\�Q��8\v���~�'�8�BOL%W�RM5
�7������
��*�L�υL��;`*�*b����2���=�^�)��<!��1x��̡���{Nt2p�q�<â��o�x�ꄣD(U�� ��

(1-�q���/L=B�B5X��S/�4�A�>�S�Y�( ����4���*LA*��$G?x� �')��$��n:Y����rJ�)js��A��I,��H�N�#4#޴���ԃ�;D��'���D�N�]�\��S(ӡ'1��K������@HlDyT�_��إ��̘2�π�%�L/2��[�H}�q�d�)mz$��v�`\�slK	%����N��,!ǉ$H���(��X��A��ϱu�@nڴ�H�+^8�N�	���R}��?QZ% 1b�$�8�jͫL)��Pe�D��d�5��X�qPtG��+d<�cׯ�"	˼,ٍ{��~2T�P�
3��O\<�SR�	()�&ώ*�dh�t��5!"0t�Ț�<R�l��SM��΄�%1R҃��3g�^Ec��U�2�E 8s&�ԇ4a�T��|R  �r�:O�,Z'�˅D�䕳�)WQ�9�v^�h�'�;T�Hu)&8>�ڝ�b�~��,�uw�+рU�
�\�!Ǖ"�]!e�\\���#?��p��K�+�ayb�A�@���AGD�6�������R,
t;t��uE���26�̠��JD�n���;�P?�'�]V:S�Վ,8�A��Y_m�'ĕ�1��~���R7v�
���S�X���'�2断EX$�1�,��0�f5�OvK-�)+� �h���CZ����ߌ,D�P�a�I�Ai�O}6�1*���4+D3�&4��kC�Gn�\1O@<3q삒�>�ZĦ�<�'	On��H>�!�ÆKO�!�a�_^4=�A��|yZ�0���+'%?�8��򩎳x9 x�pLҷ~�htp��F8o�UH�͚���q�>,���'�"�hs«S�I��B&
G�U�М|��B�B�E����ybW04�q; �M=j�m	@*���Px�k��2�:t*�퐿e����� W�L:��g<�5N��l�����5%rHL`Qf�<���G9n^	z "Mx�<) p�E]�<1s,��i�n�C�œ�b�V�<�5�ۗ^. ��ɊA�`!C�K�<�t��iH�3UK�PN>����W�<	Cg׻I�YAR�U%=H�����W�<�oF2-Y�ɻ0��|��؄mQ�<A�i�:Y:H�+^�*�h��V[�<yA�ݲi�b�Z5Dי}Pup�k��.3�>����'�D5��FP*���P�~ݘ	�[�j���A5�5�7���"0 G��*�
�с>��
 AU c�D]���+�"��e@0ғ�B	�ઐ0I�(Ԙ`">�陕o��|2 ď5P-<��Q�.1�!�ē�t	`u�a��N���ƵJ�<�Z�`V�C&$�t!�-olX�)�矴)���?���QH�6��0�n/D���
�5MDF$��Ȯk�h���Ȋ8�?�t�D�y6���K�*[���3�S�6M�ю��
:�Q2H �5=ڵ��ɒ@��١���[�6u[FA�6AN�����H�xj����f�dt�'!~�h���(��H�S��)��]Ȉ�$޺	N��A�3X\��B'\��ӸW�:�bdM, �0@��d7-��C�I s��-j$��F�pIB5#�('H�B�-"�-
S�(@[B=ڧ�yr &V@ D�ÁRӮ���+���y��)%�j�P�FN�} `!��?�J�J�(�Ff��ǀ�z��`���%�ўTp���r���X%�h�± 	+|O����	5��` &M�a��(C�>+�����>=`�I&�L�Gf��
�Q��P�g��O���x��V�M|��?A���.�n��R�O?�-�Qf
�g��'V(  q ���WB ���oԶ7ڂa�ȓ/�<of�hXpĒ8{�N\��!	4�p!F)� M8�ӗ�E4-Q>Yϻ<{�M�&���a0�#e�I��A�ȓ&���L)y��1���$�@�"�K <�ƌҷK�1&=B��L��?���Ʉ61K�+K�h �KTp���S��8:'"���T��姜'G����`F�>�  �g�.��P��!�/SS����AsҀ�B�'�2�"f�b�����0I��Qj��`ӊ�0X�lh��)��qSR�",v�資�R�u�w�"M�D`� ;�,|"R�!M��u�	�'�ԄC2�U7�����^7������&�X���ti�c	��քKNՀ4����1'�~�]QΤ�4h�#r�4\(�iU�D�Ṗ�I��F�$D=S�V��'��qBf������9#0PX`"a�%`�AP1. H�p���hO���h��I�4XXU`Z�A�j,����fN-P���	��@ C6��q%`�G�H���_K�P����ָ>���GD�>B����7������Κk� �`v���Zc,	/D������ ��F<U��yC-�����S��'��#���`�fX0.�o�<�V�6i\�����	�D<�H��h��%��+^(��m$}rmˠ0T�\`�;�ɕ�Y�f|��6$�jD��h�Z�{�-ƕ����5A��}X���b�4,ڒNX)�Z&�=��0
+P�)ϓ<����I�G�NaI5�ߚD�@��?Q����>~����2�'{��k�E�1)f��A��u�><��!�\L��" #�p@���:NR��BN�.
8I>E��'�N�(�B�t
8���N1i����
�'�F(�3,��͐ �KC�X�]��'�HUx�D�d���f/�.vk8�02g��j�  'D����@%�D]
���|8D�P�
/D��X�d�	���b���5����`9D���J�6vHE$T,g4�V��h�<U�	�x=Hы�(�ƀ�$�g�<�����^��t�'�.5���{�gZ{�<i��-�@Y�̀*i����Iv�<�f��9s�8)�ħҧOS�\�T�r�<� ����0�ȡ"��sE���1"OP�0�Յ5L�����!�XQ�"OV���E2i� G�f:�A��"OD�!��V-��ѣ	�4v�1�C"O =�B�R,�����,	RuC"Ota�s�֨~D�Pq�Rm@��"O|0�$���[V�\�C�;*���KA"O��C�M1>m �ac�2I����"O�uۖ���)��
%aމs�~�2�"OJ4J%j�qv��	 �ښl�=��"O=��� �D�R��Hń��"O��5�� T͋8���Z�"O�j�ņtF~��ϼ�T p"O�%xBEC���h�7��,�� bF"O(�k�@�^1T�'�L;;w��"O6x�/��
)��F��Q�2"O\�P� ����#�F =T\�0"O�����N<ԘH`V��2NCDy�"OT��Aυ�3T��P0�xt�g"Oj	�&�nlL�hU"�`h �Q"O�,�eL^�V8���
q��m�"OP��圫~�*�*$�`p�A��"O���JY,�B$F��Bidi"O"�� �I�f]�,��L+Kc��HV"OrY�tI����ap�Q5d��1�"O��J�	�ltU�ԛf"H�H�"Ox�)pa�}�$��fC�O, Ca"O��8��. �Ҙs@�Sw�՛�"O���G��gjv�7iK� �X�"Op�@kMҴ팬Z�4-8�"O��C7�\ѡP�&0�⌸q"O�@�Րpn4��L�0�4m0"OV� a#�>���3��<�Ƒxa"Oj(k�;h(��/���.��S"OH=;�̜�VX�KGo�(��0��"OL�c�N�[�Ή����r����"O�)6/X.���ȵM�d��"O`�a@D\"~=��e	=a�$���"O�k���E@� !״6x-��"O�ԫb'F( p.�7E�&�"O��*QGS�p`>��fl�/%�d�a�"Ov@q��O�U*l�q�ñ?�J��$"O��3S͊0b7��}�� �$"O����/m�`"'�P�G'���6"O^8� [�R��hac� �A�؂ "Obuk�k|hBb���Vd��"O�Slr�n���ˡ�\��$"O�P	�$ �`h	$EQ4��qQ"Oj�87	ʊ]���K��E�"�0��"O,��`�|)���@��yJ&UJ"Oh��.��A�`H�H�5s#�e�"O��BP.A�̶��r͏%��x��"O���
�{I�6�ؔ@��lU"O: !�*ĦZ��c,�	f��"OZ�B��;,x���$9n8t�G"Oݺ�C�+pr����֞ tb��R"O �B�-�&�h�I7�  ��jf"OpQ)�r�20��C#�2]�e"O��ŠX�,�kԉ�0[���!#"O���Ü�mv�	Q!�*B�tmJ�"Ol�ڠOʛ3}؅�% V(Fql��"O����M�~�"4oߩ�}�#"O��!d��M,d��/L�o��Q�U"O�y���<>k�H[��ĚX��"O� MYҨ�:�$�pS�-!(Y1"O�dID�Ӝ�8	S�,�����"O��zŧ���c��]!%��]��"O�LH��) �%��
n�j���"OPq1�����x"M$V�N�ڃ"O>I+ҧԓ; 8�L�%0�hI��O<A;�'͂�,��M�;,P��)��.��$	�'�H�!TK ���8!j�(E�Ja����-w����$�ӎb# ���e�z�d���ZK�hC�ɜ-z������qPy�2a��X%~�u^���*�NҧH���X#��W��\С$��:�+g"O�9�^U���Y""��9�HQ��)>}���y&��v�3����$�55Ѫ��/�O�<1zB�'M��TDT�]ٶ�� �Չ��A�QC*�$����x��<�7H�5s�t��!��t;�R �;�pE���$�������*�uAҩCDB��²U�"O�����T;.�L�R��7|��d0�P��X&��dY����>E�tJIb�^�i��N9Z2�L
�����y��e�(p�#O4J�8��DKU=}��i�ZQhCɗ�y����'F¥8%Ah�yQѠ�0Ne
T��JՆ�sJ
���뇳 ��c�1���:d���Ä���O�=0H˶g��_rNUd]x0�	ָ�q��\̧n�仐���'��9%���h��
��e��!��GnXM��E�:����'�ظ����|�S�O�����R5"T��QB]>Z�b���'<���ϡ6��}���P'.c��
�'�xQ��G/J�)�!�@#SP,�x	�'�!2�Ά�*�x��	LVCJ�
�'�6iB'F�s�ё%P�W2�'�\q�_:>0d�y�ǕC˴��'ǆ0
� S�t���NN�0��5��'������F�v���iO�5���	�'0b���h;&��ŉ ��ب�'�:i��-@*�hQR/[�SVhi��'�>a��mY7-�b���ΤNc�ܹt"�
Qْq��;&�P�q��OfPi�!L^����FR��=j6�Q��	�b��@r#dD�l�=J���$�!��܍#�^���77�j�h� �L��I 6���9'�2!�S�O�L���J�[^��6E��!�J�H	�'mPQ���'��)u��6h��aX�>	*��h�
%����}���*?�8Q@G�!�n= VOD/��?���T�Y�%�5��� �hcn�K����ހXv~���B/O�X�9?��D!���a��p�C��#��噦���_�b�t=� ��Z`�����G?�y2�G�5t���v#��R���#!J���DE7�l���^��)�'E�I ��<�.`����("�e��D�ld��ƥe� �!��M�U�\�SL��#J�����O|�>�ǭ��<��PZ �I/���"x؟�GO��Jj�{B	��r��#�J*j���0צ�&��B��4^^��Ҫ�1B�*,B�B�(O"L�f�Q�^V�ڂ*W�O�I��iU�ܛ��=I�'�RT�5g�E�$�DIJ��T�FnE�^v��@��N��`�S��y��K7$��x�C-;��`��`_��y��E�{-z1�bI*9����W�[�^ܩ�"�B-����<�']H�`��.}�'ee��3&�0P��� oP�G�����I�z�\��hL!G�p9;۴2r�p��
;D��5�v��YΓg����0�X�S&�h/O�i�a3L�O��[E'�^QJf�I:��Ä�>�����t�zT�'�P�p��u�L?�b��#c�Zc��ٺq�,� �B�]�ƙ`�27��d��2���Un�3��<��C�Lx(�����&�������-z5��D�SۛƄյ8V<��/�4��p�qP����O�����T55Mlx[c܃^�F��$+�p?A�ꎂP����hT���?	n����*�I��z���5��AǮ��Z� *�>)�xu�O�C�ƄF��ĩ�H�8 �":�[s
����`��"�X�ѩ�����L؟t�P�&���,3��k��D)��+.v�&�xz�OM�/L,��a�#���P/�<�4n[�d�X��n�?3�P�{��+����m$���� ��#��?`vH9�a�A`y^�+ԥ�x?�* z(��>,O� b�'Q0w�h�fIL���ƃ�"RzS�`m�(#I��h1D�Πe����'����O��u���Ѽ[
���c�(S���9�I8�O
m*v!"��|{�ِF���FI("��0A򯎶61�A�
A�~�I���ɑ���':�J![E$�k�+@�fE:1�h�\�'����͔C��䤯|��m�Sa4D����Ņ��}�$�1#�UC��J^^���|��Q>��T?*U��oX y]�MG��m2bT�' �a�F��$3���A�ӌWV��D��B���#����1��4�a0�a��y`/"LO�xୄ� �n$Ze��P�dY�l-�$@�R�py���$��D�J�,�e�t@c��_����"V-H쓗�5"�f��5�P�7��ܻ��D��x2�P��a�
HP���q��^N�`@��+\ψ���ا�D�ȓd%|�A���_=@�� _�#L��n�`XE���ī^�c��݅�,�RIH��(m���hV��o_�C�>}4,ݹ��ɀ6f�yZ��@�|C�I ��Z�	��HP��q��C��/Wӊ��A�_�T�rg�
H�4C�	o[@ݐ#H�0�b(��:sq C�3��$�W@Ȁ�.����v�C��H*�k�M����Kx)�򄈁B.-��Κ�^�������j`!��B>|��1!	_�Q\��s"�R9b!���<�Ah+Q�[Bv4���lB!�Y.U��q2�D�$M��,@,<M!�W<7|D=`'�+�x�>B�!�$�/����(�qR|���
'!�N^
-��L���x��E���!�$K`�0j��WgHl�X'�\��!�d,`9r�T$[>6�
��uM!��ZU`�L£�9#�Z��/ɻ;EqOe���]�0|AB�=נ�{R.��O�v$Ig��j�<��!�0`�1kt�$;q�(�)����B�JUF��O�UQC���p���T�\:N��9zO����F��#���&�O0
�>Aa%��>i�%BL���>!ASð� ��] �#'A5LOL��A|ҁ��O��Qf�']]��AU�zj�I��"O��q��G�<-z���Gn����|�`VBb����LLa�O=��rө�%Q��W�]p"Ii�'T����Y����6`]�9�"�X�eN9/J\�'qY
q��>�@�UEAd��U�״PR ���`�Z�'���`�A�O��T��QK!�1��r� x�
�J	d�J�D�bX���,��Y}�IQ�Ve�)�LZ]Ę����Q�|�#�E�
^L���D�>Y��D���AI_����w�)�yR�R�`�1K�}G�U�3�
6�?��2����w�ܔ8t�xw�2}�Hx��k����64̹�7�P=o�~�����|K��&+��M�e#H#7b�9$���;(MHW]3�<zK>A6�L���DZ/��LH�'[��M���3�O�9�ㇷX�����I9Q�T����33��\�$Q�7T�� i�a~R��=[Tq���������p��ӵ�Ԓ4���'�>�I�r������l�B�2���2�C��+V�f�0��=pIvL��K�O���$��	&�c7�����=iwb��o���p-�R�r�����L��� %.ƹ9Ul�HW�i|ƭ�bŨr�f��A��1��=�'W\�v��5�x$�d5n�a ����3砤�Rs�O
���'�Ō3��zI@;z&lL0�'�\0P� ]�RU���1vn�i֏��%:E�|��9OJM���HL���X� !��"O� ����7NX��nY,A֜� p�O~ܨQ�Z��0>��[42R@r0�Y�w|�����h�<aP�ӄDQ|��hɳE}��dh�<!$���w�1�7_�U��8�.�S�<)0��I� �5Gb �@�v�<� �l�e�N�[�����W4@��d"O��Xs"Y�xr �e��SjZ-�D"O�9i���y�<�`�g�t"��d"OH @��hI�hIe S�]�0p�"O,Ak�hq,��CM�7��"O�ѩ'-թ��R��E?#n2�"Oq�S�[��-���1.���"O"��0�|�7H��"�-"D�|�ϘI���)����F\(��gG#D����)�")�x8�d���u6l���m D�\[SL��,���a��$��H�tn>D�t�R+�4�iq��Z$V�XQr`K9D�L�F�O�B XDa��ٽ:�L�Id+D�l
�LD�R/����Ŗ�$�#$�:D�Tu���A�l��i�'�#�<D��b�H �P��c�ܫ&<$Б@6D��F�J�\�Hm	`M�d
8`2��8D��3�)؍tTp�'#Hg�A�&�4D���Ȟ�U-z����	:-2
M��(D�X(��E�'()1bb��k�#*D��kRD�>~>֬�½cj��B2 ?D��6@��a�]<a9��Ȅ�;0�!��`��藅�2A4\]9D�[�%!�J*��U�՘o�����/w�!�DܹQ���S�U�R�:�s�O�$4�!�$
O�i��6
�`{Š�P�!���*�b,�լ��+�Dh����r�!����v�2"�'��=�&.�1$!�ӗ]�@0F�E2������"X,!�$�
-ʰ
���.pF:��p^�F!�d@:39^��fa�oGθXV�!��\�G�4����5vYD��6k�!�$��^y�91%�*��8�,��a!�$�|K�4k�J]�j-�bˌ�Z�!�$H JġZ�P���9�KՇ	 !�R�\�t�H�� �|�S$)�#�!��+�r`�V#S�|�|�""B
k)!򄚪5=�3��5=��"�b�3?!� "���j׉J�65c��M�-�!�"@KK q�d�P"A_���s�'��31'��w��L�1*ԙ-p0LY�'ώa�v
˒[)JY1L�,U!
�'�&�#� G�(�Xp*V�ʀ#�'o�ᘁ*�¸�����:>hTZ�'�jܺ�'�$���'\5*j��)�'�zX�G�GUY�3�(�-ceZІȓdM�+/��H[%�Φ����ȓ9��(�#�P$~�t��n	.����9'��!愉S��`��݁_ʚ��ȓ/'��4����b��T杦R�D��Y0PJ�f�63�TՊ��D�M����	+x�f�l�px��V�E�~^}
%ӱ�h㞀���I�S�ӄ`Z�)g�ѿ^��	�'�Sc�'������D����K�Nȃ	6��N��<�B)�=d�8�ON�DP*ȸ�ħ2��9�BA�i�pL Q��%T�Ұ%���I!K�Q��fy3U�M���rB)�T�xf�x���x���Oz��rG�Kx�.�1OZ7n�dEP�O��C��铲iR��rA��-s$`r�Y��6mJ��'ˤ#:w�;��lK�*�p�:!�&�M��'Ҧ��	�'5 
5K���,f�:���jT�	p��<��J0����Ow���΍����2�cH�Z�vL1�'��H���^�C:�OQ>�HB%�K������k��+P��O ȸTLޞ~��H�zvv %>I���~���H?6��V�B��u��(�����C� 
n�!��i�4�
U�>�͟剞v%J�hlܷ�����A"�&�V�����o�)�g�? 
)J���[ư5ʂ��>�3��"4�"}:7�6Ԡ3ȃ
3�ms@m�![�aۇ�d�l�����S�U��0�5�Ӕ<�vY�U$N�o��O�������O]��s�M�-<H��T=�Y[�Onm��aڏ��	M�泟�O_�:u��֠Q�b9s@k����`={P��I��X/�aY秈m,8��s@ҧ�!��Vm�S03d,+�B�f�!��$E���ڴ,� �i�]�?�!�D��c�����˜q�J�+"�ݓ|!�ٕ��b�	',��tX�n�:e!�W yxXyt��q�dX���	Q~!�Ĝ�B���1��:O߼탗!]�+g!�$���\D &l��/�ȩ��=Wq!�DK�D�Z��Sb�P��ј���6�!�$ֺP:��p��z�\B��V�?U!�DݹF�l��e�@ ?�f�S.�p>!�dK$OXi8�`P��=h ̓�I2!���.oh� �/`)�}ˢ�D'�!�dI�{vT`�ȗ�q��%]�!�D͵:)�����OJj^tQebP��!���B���˶�S�i`� �B��!��:���Ճ�	C������!�d�3P�Zcc��c<R��0���J����Sf�W����clΜs{J���^�y��.��y���aI4DR��ȓN6���H�M�� 0��N�v����A�訕bM�"8S�	/f��q��=�$]pa��?ƸZ7��.`����<ငq1/H9{; ��q��h0��~\0�6�20 ĩ��;o��Q��X�<��EY�T96 ����vU,|�ȓ|��P�e@�$�2A$ϵ�ć�#��㗉ה;���ɦEƸ!�Q�ȓh�x���׊7rZuyd��7JJ(���С*�)X����~h��&�rx%�B1f�T�J����I�z� 
R'7oB٘��_v^���� �yQAU�/����G8d�4�ȓi�C�R��� ���'C䰆�<7�+��M�f4hF�I�P�ņȓ�T���D͝E��s�$�sX���0B\t�E	^�lZd��� ��t�ȓ<l�U��j�o�f�s�j�xv�����4�u�ѝwڼ�y�cD�M�����Q��M3��|vr<�� ��d�� �ȓg�&�I"�ÚC�`� ��A`��ȓ1��F�/x̓5そ6����ȓs�Lh`a/@wf4�Qd��-N��ȓ�F�k69]�̅R���,,����O^	���2�0���$b5��N�\����%�<:c��!a� �ȓ.�^��K�-���Q��Šyx΁��ضL���>>�zy���b�.�ȓ;P.9��"T!OvT��p,	-,-���ȓwҦQ��N�NR��R&�'09.ȅ�&$i�@Ň�q���'-Z�6��ȓe�v�@¯K���(���t��$��G�F�8wh��[��� �H�5W\ل�1�J̢�Ɨ�|Z �Y�,�A�� ��E��	s��@32�4-	�ݫP����ȓW	֥��"�9_&���"�zE�ȓpV��və�!�FM��Ģ%d���m}ƹ�t*ӕx�B��M��1� E�ȓX��� ��7eB�sC�xҚM��S�? ���.ݗ� ��'n�>PqJ��q"O���P�֍x(����n��O��*D"OL�Pꇢg�}A�ؙaM��("O�X�������KG�TBa"O�Y���X8v��2�&0���"OjI�c��M%6�1�i?"�yU"OR3Q��+}r��N04�(�C�"O^�2BM3jq�=�0�5�\�"O�M�6B�4(���@�a�2iC"O�	�D����v&�b�Ma "O�mR��Z����v��6e6j"OHL�+¬^5C�ն,��X"O���	L�	H�p`�1]�^9��"O�C#�V^�&�K%d*nʆ<�5"O����Ӊ#H-���јx��"O~li�mL�5>n�ht"ژ`RP��s"O��xB# ,"ƌ�AA�$)؁�"O 8' ' y����[)^�	g"O�T��m��z�",�q(nɑ�"OZ��ĩ�G��(���<�C"O63VA)0ݚ}Q���.Qi��pG"OV$E�	�:AL��7�;tV����"Op�CÓK�-0t%
6׆�r6"Oj��WEY��"ah�U�#�}�1"O���"HCO��� ��ȗ ܌��"O��+S�q��#Bm`pR��u"O^�� �z����F�r�<��'�0��/��x$6��B*�r��'��A�+N�r�-�p`��-#B+�'��}��`��hj�Q���BrS�Z�'�	i��$)��
0�i~P��'r�=�!߬p]��X��՗t�y0�'�4��R��;���F��m�����'��8*���n��< ㇎4b�2�'����G�Zo���7̄1W𾝑�'2<� (T��5���5ID����'a �q�͵"2���(J H����'���S'AU�6�S5��B���9�'�~�S�M�,y��# G�(>ᄉ��'-D����)B�\e��!
�d!lA��'B�x���X��i��ᏽ`���K�'� 9Yp�,��E��	�Ē��p�<A���3(�����(ڟ3ef���O�i�<yMË?`�yш�3�>\���c�<� ��
;QR���/?0�5�l�[�<yBO�}z�����6/�D])�U�<�q�C�RJQ��1}���І��R�<YV�M�?8�Wj	�u`�I�d\G�<Ѳ�A(F���I��,�yK䣃F�<q�hƄ�Vف�\�wIkō@�<aa�Je0���'���R��t�<YB�;M�v=�p��1�*�Â�s�<�3�B##r��0*�+B�z�ʦE�r�<��f��S[��HW��r=��I6c�j�<�!	'��Hj��ܬI�4̑ �]e�<�VJ��<���M�B�M�t�]�<qD�B��e��
�1�<<�'�X�<y6���_�⁉�l����RᢍV�<�УH�����C�@),?�ͺ�.�O�<��I�&`!�)��`�
���-�J�<�C�4bF�`Ô�ͤKi���RD�<IW��B���Q ��KFm�~�<��Ӱa}���ѥS)�I;�|�<ٲ%�+Ql�5�v�ןO���r'B�o�<� nL)h�[�dM���~�^A��"O�T��+�&-��J]G�`�P1"O�PB#>h��@��D�^�v�z"O�� #](��:�N�7+!Ԕ��"O�YٰGG:@2f0�M�'���F"O�l����8E�L<0�KՏ����"O���fū*�#ª��+��`S�"Oj�h3��lF<�`�+H�a:�x� "O��Q�<V�:'H@�Q(�!�%"O`Mq���,Z��ec��H���K�"O�hd��>F�y��倄D� ��"O���1,F°أ��M�,���"O��C�IȐ1��k��z�v-��"O*�AgA��TN��w�>Ji�ع�"O(�6�ގl�t��� �Tl�M"�"O�L�R�V&?�(�j7� � 5:�"Ol�ч�U<9!\+ƪ��Ҁ�C�"O ����%.��В
�%�j�J"O�0Xgٱ=�T����9v�B�I�"O:q�(�G󨑊��̡H����"O�|�5a�%f����j��Z���"O~5��CS��؋���4A|���*O��q�O�C���
���,T�'),�zg��%�A�w(9��'e���,Q�rE��b��D� �+�'O�-� ��31��z�kH0��'Дx���%I�h<��L�W��yr�' � ��E�v��� �����'qڕ�#Y7;�Q!��֖���{
�'���*s��C�f�ҴI�6w�,Hc	�'9p�)E�J�u&F탡�6Z�E��'X�0$	7/� �Ca$b)�q�'ڜ���g�hS�e�E �O�����'�n��eXZ��}�%�E�Es����'��PJr�OB�c��	c�]��'.F�x��)t��Q@�+��	�'���@2��/`� 쪠$�+w��i�'��)�d�ʔ12xH7mUw�F�q�'"��s)B
R�@]xQ䝩g̮��	�')��˦g[&->�0�u�C�YL.H�	�'�\�� 0=3&8@��g���Z�'� ��B�{���e��tǔLR	�'\h�1�Ęb ��#g��X��'L$e�&�ʈl���Q��X�f��d�
�'�*������Jٚ��GB�n�.	S	�'��1J�ʵ�I {d�UK�%��y��
q��0��#�J4rb��5�y��(A��DzJ�#u,������yR��P�� i�㊜h�!)�̓(�y򎌞!�v8Y�ډS#�s!+H��y��KR��Y�=3P��0�yO�;j�Ā����1SN�݁��؆�ye�8 .1�UNS�O�4A JN,�y��L�r��i���7G� ��d���yR�_']4@&@͑E,$���3�y�<?��]C��R�6��-�"�0�ybI�
	�M�m�*0������yR��,j��8u�V�/��p%�Py⎙����ym�(Ѭ���Cn�<`�).$��)2t�"l a�<q�ʀ�P
 b�P?o`����QB�<�%Ƅ7�f�Ö��;X���Sa�d�<A@�B�b� �*A�\����RM�w�<���G$+��U�"�Ȱe�xGq�<� D�2t�T3A�IR`���I� e�"O�Y0i˗tk@equ(�P�4ly�"O4P˵*J /��Z7���.�>�"O2��t����Q�D���r"O.�9R�g��H�Ҍ>%*�"O����k��9�rI�@$�& "�"�"OL9��k^3�\��"i=%Ƚ�r"O�X��[ʀ\mܕ\J,b��2D�y�"�0`	s�b��=���I/D�����'q��Yk����:w�,IƧ,D���    ��   �  m  �  K  �%  b.  �4  �:  ?A  �G  �M  T  IZ  �`  �f  m  Us  �y  �  �  \�  ��  �  #�  f�  y�  `�  L�  �  :�  }�  �  I�  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(�'j6�!�j�Sy���(�GD�A�'�l�`���!AnU1�V�GH���'8 81����u���Q�J�5o|��'�QIE
�8��Ё�۵4jxq��'��aj֕yn~,�0�]*� ����$�O�}jǪ�/G
xs����r�h'�h�<a�IQ#gq�Ї�5^����D`�d)�S��4x�H����V������[��p��!jN}z�ۘ.�K"�ۚ-�H��'9�}bmQ�4�R�YP�Lx�����=��#��F/X��e�%��.)�$�7&٢-�!�р=�D`K����А&%���E{ʟ��ߩ+8�����+|i��pF�*D�� S�+Ī�ɴf�=/��ۅ�#D�p:6���PY�f��n�Yä� D��J��]�k�FX���6���c�K+D�P�Ro�#�X5J�Iu�h	`�=LO�� �6�_4U�4	K�#�&�,�9��'D�@�&o�Hy �� �(]y��1�y
� X��,�	��̒��P�$�Z�`""OlD��+R�..��ǯF��6"O��{���6W���"I�)m�t"O��91)׀bP�̑@��<w���AJ-4���4��.m^��	��Ūm���[�@1D��ڕ��9�4(d�^�2��q�v�#D��+�dE�G��q� ����HE� �ɻ:�Q�b>Ar���}��Z�o�5^��{��1D��8�Ӑ|r�3�	صV9d|&.���]�㉣X+����o��)>(Y��DQ.C䉍>��d�v�	4iP'�7
��B䉣4>��2�-*�ˀ��@<�B��;�hT�uK�#]W�� ����]CfB䉗z���bJ�K����7c�B���qà�$xצ1�"�\$C�ɺ�8���&��-B�u2q-�B�i%�	�E�Vǜ�aEBت�r<S�'���h��� J%�^���R5oK�y"�N������\=����.ֈ�y����8,42�I>� �d���yk�QЀI��#S�B�$$�y��	(�v8��g!}O��8S����yba��'LAs��[o��e{��K;�yb�w!XB�6���@L��yRτ?~'xu���ވK�̘�a��y��l�,#gE���̒�M�ӈOZ��E$���Kdǅ*5wt��^|�<����9�n	�I�� � `���J��H�>���g��Ѓ���V�����-E����]$���N	"}�Թ`�,��=�ȓ``5pcF��bq��u�J(MƆ)�ȓm��HZ���;��un@�7�zԇ�kÌxаjȾKwα�q�ɑ)*�l�ē�����92yK�o1b�؀[@"O��R��*k�pI��M�f�HA'=�ļ>����O�A!%��[.�P����.6��qR"O�$�OG�M�2���� |�|� "O��p%�1fU"%M.tV����'��'�:�jW�@)��\�jJ�!�����4<O��� �F�GoP�c���sBl0��'�Q����)`@ݙ����P�$D�p ���5��y8f�Ůb�U��7D�t�4�F2`1�	Ĭ2��X�A�1D��x��D�����< ���+�d1��n���ӌ� '�-Y�_�i�ł��0D�LhUDI5D�VHh0���v��1�f/D�� G.6-N cuc�;Y򒙀3�9D��ä]�&'�qFQ�HmLY�a):D��I�8r�R��
f$E�"@*�h���OdD̀���ػ��ч,���	�'n�t�g&�Z9:�����rzvR	�'b��5��0YP�x�S�'B�I� �20�!A*j�H��'H��y� e��y8A�$_�ݨ*W��y��y�!J�Oj�����F#�y�h$4��۹@�,+d#���'Kўb>�	����a�yR0h�'���-*D�T+g&��u�L=��ϓ(��K��&D��lObi��b�#M7���ذM%$��ӏQ fnM!�@��$G�T��b��y�E�*qZ�h��FE"Z�P��K��y����
��q���;��HI@�U��yR�Q�O:F�����51VX��/Z��y"D3g=BI� "�H�K%A+�y
� ������H�$��G��&O�(��"OT�r��צ!����'�<�T��eOޠbI��(N�Ya�'�V��x0:D�ۦ헣X2�q�˘�+�@� 5�8D�<2Qo��{^����8~F�{��5D����i�)W@�厇�A9���9�@���O#|���Nd��@̎�(��'%��X��E�k��@rRD�?s0�u��'�t��o�# H,���Y��x�h�'�6|�V�q���&�ř�Lŋ�'V�������f�ԗ �<=[ϓ�OQy�#԰~��8�,]4�] �"O
���b�/H ����( ^�z��|��)��j�N̘B��8�P)9H�'KXB�ɪ�B���OE2J��H����f�C�I�U�@��E��Ph!�c�y�C�	�"w��&�H�s�z�XVDj�B�ɝ]9〈sl�
$�
�(�
��Hy�B�I�7U@8��E+G"��h�XNB�I3A�({"h�*M����#\�4�XC�	��"��4�áAJH���&_�B䉺j��,ZW�	�2�T��E]#�B�I�I��iǂ��]�`���5t�6B䉸B����ɑO
�i@��z��C�Ɉ`�xlt$в'3؝���3��C�I� T�vm� v�Z��;%�C�6-ƞ���(�2V_^�J�JK.�C���8����ۢK�h���/�x��C�-n��p��숱OQ|��'��w��C�ɺ]h�sgF^�@.RU�&(E�sZ�C�63��:D��?�0�ٖ
�}�zC�I%X��sg

QR�L6y��B�I���-��E�c����2�P)�B�	�.���Y`��3J. y�!�elC�I(�H��%�������c����hC�	$Ş�+3�Ǝ6���p�#�B䉱~*�����Y�|��%�r���w9�C�ɥ]���fd�?nv�!�pÌ'غC��'6"���r�Z�0���!�!X���C�I�_��mS��#8��EI�"W�,�*B䉳Y���T�P��
e�eMPB� Ĩ�Ѐ
^�Zjq��n̩=RC䉖��D���г	��k���X"C�	~�z��F�F����f޽FC��$����W�^'�\{��/h�HC�I�+
�ϤE� ���O��C�I<R��k� � ]N�����O�2B�	4k@,�C.؝&]�3Ċ�B�#XNԒ�S��j��Q���!���$ZND�h��/Č	��F�e�!�G9i�^yP���6�"�A��v�!�$ؠB�ڤPtJ�9��x��;"�!�DЎQ��@��a66�ɤ�@�3!�->���P	n{`�9N�+Q!���m\5���C�2]���mJ�Y!����+5�Ҟ5F����mɽf!��R�Lx���g^�B�m�4J!��Џd�����3B4}�ek4�!�$
��8у�͋i����1HO 7�!���7N���B�J�M���
\�9z�'���3#��x�.�%��3C��Q�'�н�R���V����EK/=9@��'r�a8��O���dT�/�X\��'㞤#5M�ښ��P?%x�:
��� z�f��5R$9B��^�(��R"O��K��"9@lAAh'u���"OJ}A�#�9�͈4gHsj@�c"O��/*�8P'�pm���7"O��ڰ��p� 1�f��_ObHYu�'���'"�'�B�'�b�'P��'�z�(dMKo��I)�l��(K���D�'�"�'���')R�'��'N��'׬�d��d��sN�W
���'��'���'���'[��'aR�'*a"�b��}�ش�S�çR��"A�'1R�'~B�'�B�'�2�'��'?�ðK�!Y8�10�i�
$�� ���'�R�'��'x�'N��'�R�'��hz0�Y�t����"ql�4�'L��'���'d��'���'��'B�X�����AA��\7����'B�'�"�'JB�'�"�'=r�'	��E9��qC�80�}�W�'�B�'+��'�R�'/b�'���'���f�c%�(�aC�Js(Ju�'���'�b�'���'��'y��'��P�Ad-������33��TZ��'�'���'�b�';��'��'��▃8M�r���l+)��=$�'R�'���'�2�'���'���'�i3Î-K�����G�J�,�w�',b�'#�'���']��'���'"=�Ea�mh�kwƒ�

�Y���'kR�'��'���'���rӔ���OR�ԥւ7� ��� XAd)�ay��'b�)�3?�T�i)5�7�U(I�z�kP�N��X��2��D�䦵�?��<	��G�P�ǅ�#��tP�&�!6-ZHy���?�����M#�O��S"�O?I�Ys�d4�6�̽v��9�b+·Ԙ'�r[�$F�H�2S�t����'?3B	`R%�y��6m�9L�1O �?�C����6�'x|*���C��d�ڭɅ�ނ�?���y�Z�b>]���馡�I��:Ǣ�M��M�ĉ�ZwJLϓ�y��O�Y���4�&�����E�*��a�ܘtK��Z�'���Q򉩿M���N�:��s`�׎Y^�� �OP�%�0�����>q���?��'�I�_�>m����A��F��<LP�?!O6i4�,�|"o�O�,B��[e�����R�%���3��u�-O�ʓ�?E��'��A��R f���'(d):Ha�'D�7��7����M+��O?X)�rL� @�2#ˈO�
ਜ'��'�rE<Q�F����'9���J)D�|��	W�K�ht�vG�^`�C�ɅY��<����d�!8�
I)(��C�IR0z�CU�Z�2P4x�ę(av�p�#=Sj�q�3ā�_��a��]/:`Sd�!wd�81Ɯ<Ip�4 �0M�S�`m��jߏx��xу�ݹa��`�J/v�΍h��7|�-+��L5��hڅl�����
r�@���v�yr�P=X��S@F�A ��@x��@1�D_�~?��9�P(1�e0Î<D�H�S����+G�3cY1 ���rC,i� I�;F��h�V��qH�F����m���9wqR��q��n{\�:���S���3��'�t�0E��y;đY�;��P��DYE\I�v����P���3�$�F��e�)�d�\6V���c��ȟ?dȶ狚(u?:�v�-OX;׉�������h�	�u��'���8lގP�I�p���Kv�$�~� D�\-�����)`h���dT�:��Z#�'���*�o����d�n�b�h%�ӹJ��؅�I�!|p��V	��%�QW/�(5����ɭl� d����M뷶��,O^���<ª��iuZP�#@(2�|A��T�<� �"�2ɖk� ,�U���va��I "���T�i�9��@�2;b��3���U���2�#D� �(�^m$u{�E�EQ�0���"D����c!� ���ؓ#x�H	6D��)�/ժt�r��7W�'(�0��n D���Сb�\Eh�UVi�H�+=D�`i����g�d,���/H�z ��;D� �&,�07v�)�(�+;�Z<��`4D����=8D�S�j �l�X��qn3D�0"Whʝ�<Yr��H�����,D� ��I<�e��fR�>��I�$7D��نBV)"xB��4��g�&��A4D�ↈ����!3��
긅�g/3D��b4��:>Q��*R'Z�[��-D�̈�M܉,U��s�(a2�y�9D��c��D#".=�w�B4h����5D��
�T2�P�i�����s�.D�4�f����ՙ3�8���Q�D.D��	`�4<oZ� ����@��,D��re �)��!{7�I�f�X)��.D�X⶯�K(����<gN4Q��H8D�� ����<I�Xc�9 4
�"OVp�r��5Vv��$ቐ\�&y�!"O�xcՋJ�=z�͛Q �c�"OؔC�+�`�Q�թy�\K�"Of�O,S e���"Xcx�8F"O�  >L���̝Jb�5j�"O����~�$�/�q]XE��"O
-Q��
KrU0�Z.=C��a"O��0�)bJdTy�/F�ӼeB�"O0D�#�O�"�ȁn�*Y�vI#�"O �� ��zR�HP���0K���$��5\O��B�һ`#��@�+ɺg��h��';��F�S*MÐ�D�n��q�m٩6�:B��A��󏛆<]�ast�>��#?��ؿ?\4��~��+|�.��.p�.X��)�S�<��W�`�D�G.ĦK�B$�A{?!#�N2�6�Zvh�b��2��m:���2��xM�i���ǣ�	��l`D���3"�@PŊL<'֎Y�N��^�&H>H*X�������ቇa�f��E��;i� �#c�-�X��䆠 �<�1k�c���K!���	f�)�'��8 F�3���T���͖U����.��;��͎f��1D|��ɒJ���c׍�9gR������4��,?@���)X�m�>���K�1�y2aբ��oJ�I���0����Gk��
gZʂI��CM0��6ił�h���c�*SX��Ë
�u�ұ�d�'D� {�(+-��] ЋDw���Z�E�'��޴K�z�
�O�K�i�O�"<�s��V�,���N%C��!��XX��JLq�N�ue�F1̴9׈�1F9���A`�v}c�\�3�-�.r�f�$?#�9��)C��uE{ҍ��8a�غ�ߨ/�(�G�������L)oW�i���Ӝ8�\t:#l�9�y"�"���v,�<8k�b�@��y�f� *G́��f�D`[% *�#��5PT�R0)���UNȦf�,��
����a��+��L��#�Q0��dÚ�[&���̻)Ur�'"���ቒO�z�q���ef`�5�O�	X���$�$l\�}��9 hX�g*^��&91�B�x�0���:&ℇ�	�Bt���GƂ�OS~�c���HN$#>AV�3w}�Y��aڏ1��Q?���	�.7���3hСKĎԫb0D�l�"ӿ8��{��K�r�zx�@�l����"��w��u+���H�m����$"��NR;I�y��S�b!��$Y4\�g&�d��9A@O[�`�0M�AI�O� Kr��3Dt�t2�?#<YuFGET�DvjX�-� YQ#�2�O��g�Ҋs�:=��ՐLl�%g��`Bĉq#$�3 ?\B�	�|i��ɢ��:0�D�!-Z1t"=aԈV�tI�eS�b8��O��d3�8F�(�x�N��\Xn��
�'A�'��C�:]XP�����شvq�Qt FG�S��Mk��W��+S�_�@�Q��@�<�"�ۜ |)jEM4!��kqNw}�CA*��Ih��ڕ��4ApLe풦?ɜ���������G7"xᓭEe�����Ͻ��C��CM��z̬$�i��e[��#=i�e��f�?ݱ`��dD90m�D�:L��-D���c���?&�cB��~�L��Mx�,�����$������f���~�����	�l,�W��y��ϯ/�| ���.az$1��aϦ��� Tv�'�'�$���NA(h���2f�a�Z��
�mB��7���Zr��!P�򱙔��7N���"O� {�&��$�����d�k��ɫ��."[p>E��C��i)&��IF�9t���wF%D�H��F�Se�}��<���ەH�>)��˿o�`����/}*��'媉�␾D|*$Ӑ�i��Q��'e����-L0Ry�ك�@���,�����J\��e�X*v�'��y��ϧE|~�	��P�aB�2�-�>,����0 �7a��m��#h��� ũU;�M*�'A�M����Kcj��5��b�֙��O�՘�c�S~2�R�,"|ڒh�Va�yRr�!P{���X�<� �u���.c�����o��-;`I9E�Op��Ĵ?��m�C�<�Ϙ'�v���E�2#�����0#s��Q�'Av��e�8���KT�_87�����ך'v~�h�n��'�'��P`h��z��5��h�EӐ�:�#\�a����8�L E<!�%.Q(j�^D�$'�;<���b���	�q����J�0z��f˯��^��H5��djrG
�u�'F��N=����4�4�a�v����'j�
���3	h��Ye�F�B�L��TŜHBWG�>1!�٢���
+�x���P#�Ҳ`-��9�&�)�\�ٶO�Q!�gN�{~�@S A�#>�@��a��t�v�_2(� Iz���S!2Ms�&Ӽ���	%"}8�+��ʹB�l������?�`��jg
�Ě3�XQ�G�X?��49��A����c!?�5�C�^�s[��E�@9�0>	FE���i�D��10y�Y��W}E�rd���ߴU`�|BM�:H�I�y�O���#�ö�X�(w�Q2}H$	�'袕@�1q� ���Z�W�.�р&J9A��� ?��9O��?nϪy1�r���6�~13��? ������6/����D��I�L� �G	��-6ㇹ+�L ���V2@��� �~��&��YLn$��K,Dx"��` �3D��.�|p�E���O&�͈�<yc�mJ�ϓ!�����.`26I�u��/(��ُ{k��"k�T�C�#_\Pu�%��o��HI7�>ᆢK�h��DZ�y�����~"�i��4��њ�A�6���䀈&<]Dxp"O�\j�)Ź|�4[d;tʞ��$�܅fR�͓��A�4O��T?�O�K�0���p�� �ΔPc%Ű?��@�p�H�Js�U�j2�t�OC3�|apQ:OX�DYW��LUd#<�-��=t$)Ո�0O��I���l�'��7(Y�|�yx�Gҵ��iD�H�t`���3�dK��Z)p�g�f��$P�c�0��(<.y�YB�o�d��<q�p�W�"?��" '��O�)��4J�	Wެ#�/!��Z�*�jL�A@E#Y����닢 ��Īv���<���!l9�)����g��K���(
G����C��B�@��p؟�����djF��0*�|y�� �̅Iu'P�&�S�
:�(O��!AV6t��Q�e�+C&��q��	,I2��a ��S�X0%�~�1�ͽl��Q3Wg�L���Ñ�j�<ї�t��Aq��x�A����fy�}���a�-�6�ɋ��L�N�$�P���wK�|!C��E2!�v@��Cf��	BFl,A��c��`F� %��a��Y�8�tJ�5�Թ��"U�\p#C�<D�8�1��5z<�p�٨y��9�U%�O(=3T��M����� k'k�;V4Ĕ��G#^��0��IHq~5�aG�<�'H�K�hQ�D=װ��Oj�<aU��*���@��N�!Cj�|�S�ȑ�"�E�:�?�ib�0D\��*ܤl6�Lb=D�h�2� �?Ǧ�2���7q��j�a�mcQ�wd:�D�x�����  �d	E���ݳQI
�6�!���[�ƉD*&Bɺs�O��HX� H��d�'�u��@�% ��b��p��=��i`�y�5O1���$X�.�i��V:s٦0K�"O|A��l�`yh]�R�^��P��I7T> �q���י0D�Yrs@�o��<��.-!�d�@�n�`�D��'�F@��ՠQ�@�-VL�c�"~n�.{���`h�G�̬A��Ż[&�C䉙30�"�	Ym	>](T	G<04�H�iH��'|f�i���:E�h��AC^+=�ڑy��B� ���O\xB�]�7I�,��']vk��b�"O$���F�R]��X��T��&Ô�	�\�H�p%a:�'=b �
�CC�CM�8ɢ	ۯ/��d���V	�G�Y8)T��39�l�
a9h���/;�)��RE+��<�2�,�3p=$4rd&D���c#
}����ˏ�s� 3��>��)��=�����/(�a� Iυ��|�'-��R�a}�GBae��	�]�8���1yh���,ת'fC�I�[>}*W�W��F�|"=��/ӺM?�eΜ3J�\��@,PI@��� 9D�`bf�F7aIiƄ�/@av��@uӬ�� `S�S��M� T�jd�B��-�Տ)����"O(!蝏E��C$
]8���UX��n�0>�$��m��� $�֢���#��fX��1�K���y�m߅0*���X�C��x��V�yC>Qt�� AOAh>-��j��hO��Ӈ�Ӧ-}�!
J�n���#&Zt'�B䉿��@���a��Ա���sGXB䉮,�z�L�
Y�|��L�e`C䉖Z���L؝p�d|�RMޣmʀB�I)���:�e��}~��e��5�dB�B�6)��-�U�t ���+�C��9�j�@K�\F��6Y�BC�	21�~��&)��d� `bsC32�lC�IvѸu�*ơc��!K�D�4C䉋X���k��C$rO��3�#�L��B�I
�D�Z�̒�\�\��$��$yI C�I�|��À�9y�y�'uJ>B�I1X"@K��� Wq��	@c�C�:t��+�R�?n��P��ނ,i�C�ɸX_F�0'�=ۂĚ��X�.��C�I��}8�`A�c5 ��7�E�C�	1z�lI�٬�q���T=3��B�I�F���+���t��#�E�<�B䉳 ��ā&\�.��XQF V�B䉠5<@��ᢍs�����&:�,B�ɁyT\q�_�&�4cU�X�B�7u�\!�E
�)�24K�0�FC�	��Z,��+9U|q�K�6!(DC�I�K�|���Q'<�͔+�C�	�(J���Q   |8� ����eB�I�pt��$i�
O�L؊�IO�)��C�	:51F�s'�.h!­Q�rA�C��!v�̐)�P%\��"f��q��C䉃6ʸ����Z�8	­H��
-9l�C�I	P>��)�OI�4j�D���=i�C�	�eZ������J:JH�ԉ�1j>B�Ɋ+�⡒6 �UB$LX7�Q�B䉣��� ����/4�"`ʇ�B�	�dI�%�	L�-Y��.�C�	�1��#�!ȏdV���@D�!"�C�I2[�4��*46+!��XVC�0&�l����Cs=4�
��9�|B�I$?&�I�V-H/3m���¯N4li|B�I�oX��`�A�;R�Y�C�2N;!��Z�6�4I���zN �zG!-Z"!��ڑ1�%�B㗕C��kD�[��!�g�����Ϝ*�p{���8p�!��H���ˇ�5"�{4����C�	F��5E���<�1G,O�#WC䉞)��� B$!&�{cHF�B�	�p��H�@�w�H!)�=CD>B�	�w�L�c灥<"�2��M H�B䉷P�p����{wF=�1·o|�C�I(��@�oV8I�4� ֏�M�C�ɨB����dIȶgVI2�IK�K4�C��=1�j�Ss��2S��k�����nC�ɆSMl�`QlK�UwĤK���R�B�I�cȤ�;$m]�_ߒ��"HT3>2�C�ɟ<w^��4%I�a�d@T/F1M7rC�+%��C� rBQ���C}�4C�	�S��*���6 2 ���4-2C�Ɋ(�>�sDI�~�"��>y�<B䉴�%Kۅni �1�	�4%�N5	%"O��1*'�� ΚU�7*D�� >�鐻4E|����	>����"O��a��I�:Z2쀆t�dA� "O�%�r�G6GG��;��E�q��"O���
�p�0) �hܲ)v��7"O,;��IQ�q��
�B\�8a"O��+��K��\Ҵ��_|m*�"O&��d(�;T|�"��e[�	9�"OV���֪)L�,{�5g��y�"O�q�v���Q9��y�㎟q���"O�̙���`�����jn��"O��������Vo���1��'���
�dƖlz�ӺI����	�'6H��$��^)1W�P\x]�'���5"R�k�t�qK��M(�y�'�v���k��R�����R�Do.Ű�'�����X�~�1q0C��B��:�'Ơ�ZN�/d�(YՇ������'� hFՐOw�x��
V��r�'�������?Fb`)��&$~d��'��(����L�z�C7���y�jÁD�� �эS�>�R�0$¦�y���:CI�MGLX�P�,?�y�L�:2k�؈6��C	���n�6�y@���[�M�<�֝�am^�y�c� e��cϥg@�ifJ� �yR���gƐ� ��Žf�e�Ug�yb?9I���F��)Y�D���
4�y�$�� .��uj�@����f
��y"�O�spV)����&:_�X�lD��yb�ݽ��pXG��;3P¨!E�4�yB�9>�K�m; 8��d.���ȓF<�+����M�"h�pծE��W�0��Z�0Su�ߝ2@8�ȓfL�ӇH'9�]��N�KEfA�ȓ<ZЛ�b�(�"RB [����ȓ�h|���;DT���`m�Kj�ȓ\�q�bė/l%�p̘�? f���FT�ydE [�m����$Z� ��>����e���<�c`�K�'�����o\u:��G��G#N<�1��g�"��a���bPcW&�n�48�ȓp D�"&��2f0��Jrc����ȓPd�2a���mB:���k��Sz�9�ȓ �nl�Bh"s`�\Z��K�b� ]��J3Z��%H�m���g0u2�4�ȓ�:�r�XZ�6��׉�+ �J��ȓG�P�I���5J*������EuDцȓ��[��R���5+�����a�������`�%���2���Q����j9D��xҡF$Zu���'B��P�F4D�(��*D�R�2@��ϲvK�y��,D�P�3�ʕ�z�zQI��y�֐���*D�T� �4]l�$1��5���*O`e���
+**t3�FRx�D�� "OR]���O�|�R���˒s8�\Z�"O�k������ҫ��a`p"O�����7 � T:uC(^d�"O�I��%��qi*8:F��d���v"O�x���� `�y�O�fHЀ"O2�3�ϋmb�	����3a�H��"Oڸ�#.�BU`�.�Ih, S"O��8$��tf�)C �*�n�ib"Of\F�X�9\J@�f�.q؆ݘ�"O� ��(Ҽxj��y�$E�j�@	�"O� ��R/X�0%�31���,	)6"OND�a��dJd���&��%�T��"O�k��9�0��E�P6d��4�"O�t����?,c>9S"�"4���9�"O���Ɓ�Xl��7e���a��"O���p�\d�L� �X�E��"O����WK@����-�|9Pp"O*1��m�,OP���#ah*�S"O�z1��l������Y5pe��yv"O�1�ѩ�_FHUH��MIY��X�"O*�����?O��Á�vN0`T"O�����=s|�ms㆘)}\��"O^��SOAQ��0�$���}��"O�h�â�ZÎ=�ge��~��m�"OT���T���Ȕ�Oڢ�����yr
�N��Z��:H/v����y2��?,�V���-EZ����܄�y2�
h	t-�� �V\P��D��y�\�'<���p��`ryj�h�/�y�l��()D�acLM3�!*t�+�Py�g�~1�p$=2��a!�]e�<I��-� Q��%��4���/`�<y�)wj�|A'Ǟ�d�$P��,^�<y�c�7	*��b��z��؊1D�U�<�%΢�*��T�O:8-*l�S@KK�<�b�Χa��]���Ӱ|�@0�d!D�<$�:c�t�2A
�-�
�x�<�ҁ�.�ި�� ,��U�"�k�<A��ց[*(xI�k��.~�yI'!Gg�<Q�]$���F��p�4��@O�<Y��_���C&�K�=S���f�<1���m�������8% [��|�<Ab����9Ƃ�n2~�pCA2D�� ��r<4���@�wF�j�0D���#8'K�4h7k\� $D�	�,D�ġ�ƕ����,�1[��]��(D�����,(������34ʀ�a�&D�pJ��^�1A���B��r��a (D�xxsM�����B�B�0C�;D����d�:GĀ�JB�߳Q:yP��-D�(H��o��\Foܜ>2� r�>D�T!�	BU儔��-K�"D!0�=D��A��X71C^�!v!�8$L p�M0D����H��|0ܑ��]��Q�A!D��B�,�̫@HP:^r�i��?D�p����#
�و�'�43���3D=D�D�蝹z!���2ݝZ�V�k��9D�P��[-xrZ��BKի)?V�B� 6D��+Q��`�~�S��ҮWWJ�I��4D�<�"�v[��8����h�Dp�fM2D��2J�e4��:��Κ+�*�@4D���"hE�QN	�b��mdD��2)-D�[V���ΰ�;&!��2�xY0��,D����TXL�m�掏�G�,�Qe7D��beC�A�T�S6�v�4X�u�?D���E��H��=iT�������=D�Xpo׷f\q�@H�}���h"&D�4�0��	Z}�Y�U.E�$�dٚ@
7D���(��S-��Ag�A>>LH���L:D�@�r��52�
���ŝ;	�.%�Q�8D�LA�nR�"$R��q�\���x�b+D��c�*X�r ��Si���l��d4D�Ը�-�&!��jS��-�n4[�(D�h��ϻ7��U���?pA��f%D�� 4����P5+v��v����yZ1"O�P��ҷX�hɠ
�>5��@�"O M:��6'����(��LΨ�r�"O�X���m��h6H��m,�A�"O,���Δb�c�fX>�JyJ�"O��0�aS
�B�k����!�"O���kR)>���R#P�4 ����y�l�K��h���< 1��
�y�K.�ֹjǭ�μ��`W�y��RI)p�0Q��5x�8�1vF���y2B@� K6�a�'���r٣Pϕ:�y#D Mհqpd�= >��z π�y��4�p5�tKA�{��1�@�H��yR$͹+H�h:��1 �ع ����y�� r2!أ�ߴ��t�r�1�y2*��p"�A�M�I舠Ҭ�0�y��	�I�p��H��{�
K��y�R�L{D�L�x�\����H��y�cQ$��m+d�[�[���N��y��HD:���J�X��٣ӣԇ�yB-�"J�`�B肳HX���o�+�y�e��z�Jb�m�p9 ����6�yr�@'r�fU ���`�l��G��y�H�v�d�1F떬���D�yRC��G�"��VJ�;l0` "�yJ̦	���� �43l ����y���ę�Ae��<�@���݊�y���dbdHGù9/�Eɇ��+�yrfZ�% J��e��35�|U��,��yr�Տ4gN�U�91�b3�k�*�yrgR�b�*�!t׼"X��֨��yb���
TLE�ɉ�/�p 2�&ג�yB���o�Pq�0�ӏR���+B���y2�<v�b0q�/.J�<�(b���yBH#*�!�	<N��x� ���y&��)�0�%ҵ;d�r����y�a��N,:%� C"๋qǅ�yr���d�+�#��h��9 6�T�yb�F{�FRG �2D�+Rm��y�h�	U-�qJ��##�1��oL�ybJ�i�h������]c�A���yB�]u���A��>D��J��yℝ�&����U�XQ��S���8�y2�Sw�8p��'��|�9�G��yB�����B�ֲ+�� �����y�r�,���R�䠸 EO2E�C�	3v�:�j��)ŮT���:Q.B�ɐ��i�VCV.(W��S�a���jC䉇 Z�5�H��*�h�L��FC�I�s:��u(��������F
�C�I�B:�A�@Q�C����be��tC�It�F��P
�F'<t����;oC䉝h@(Тe��F��)a��0h�B�I;e�����b�6i����Ԇ��A��C�.<��I;F�ޠT�X��YU/6C��1zuD��	�}×��*sm�B�d_��˵�̞5R�M�W�
��B�	�V�F�q �L�A�����z�B�I�t����"�:��$%Z3X��B䉏d��)@���0�D�ڬ6��B�I�s������t���qB�����C�	}�9��m�=(=�pxR�©A�C�I�.Wܤ�``̱paVK��C�	�C^j��K�C��1R��'L?|C�)� ��:d+�%[�wy���>r<�A��,����NFN��Y�ٻG����ȓ^d�R�ǕIfȍ1���0 e�ȓ3��8�MP� �@|����_��<�ȓY���ʪoK�|��g�]�����䨔��-N=�й�G�|���ȓG`�D�#V0[����E�W�x��ȓP�~�F�����.]�,��Y��m\T�Q��T�
�Aǌ�=&��T�ȓ:���������$2$jG�u�!��g�&���-(��|�`+2�R$��SHֈ�a��MjX��&�P 1�<܇ȓs�L]�#ɕ�j$�1�o;�:)�ȓbDvQ��+U�4ܠ\�2�̵y����ȓd��ȢGr����ɳE���7��@���d��� ��հ�T���=,�х��*XhiPuo��"��ȓ~��)�7��Վ4 ��A�ט���p�D ����(O��1`��޺-��E�ȓ
J��	A�?����&O9l~�����p�ٵ�֮�f�1��L��4��m�ːK
 �n��K�\�tB�	6MztCV�LM���U��o��B䉤^:��4E��|�`4��l�0v�B�	x�=4�P�xO�Q��@���jB䉃z�ey��NYZ�zu%�1�fB�ɺS�B���Ȇ:�n��I��<e�C�	]4>��'�ݠB$P�Sv��U�vC�I�8���B ^'�����v[zC�	�|G�8#C����!��/u4C��.s6M�@��5U�X�y�H6�C�� )a�� �&B�$Z����C�	�k1nE���"K�eÅ�:U��C��6z�~��)	��"��,�zC�
r�� @'}�J���ŨHlC�ɥL��`�WI��w0q3Rg�)d��B�I/Θ	qM�hfnS���&P�B�ILD$H��j�/[�j4�#d�a�B��/n�<�;d �����*DF�C�ɣr�!�KW�32n�h��5<�C�	��UUi�*df9YEI�*P��A�'���p!��bJ�����6|A�eX
�'|6�1Ԋ�-@����GV�l��!3�'��@xf�	���a�P�A O��p�' �;���F!N��gቸ^�JEb�'0谂fO��5�W�[�Q!���'��y{�Ã�n5Z�A���=Pͮ�b�'��\�,Xs+X�s���*B�QY�'o|����Y���;ZQm2�!�K*D���A�#�|5)�e�5@�X�P��5D��d,�PY��2%
�^[6��S@!D�H���Қ#�(����J�n�2��"4D�Rq�����I��	NmH��7D��s�وB����Z9l)��s�+)D���V�*'?�]h�#X�L�� ��K%D��3V�BJ\9@6O��VȔ�a&"D�XI�IΫj^M�V�5A��ٷ"D�<kH�8J�X�����FdD��ue<D�xR���4��҆�i�\%8�k8D��R#���U����.��J���j�j5D��+��Y�z�hU��'ױ�M؆�1D� �u�l�x��c�Ƿ}S�����/D�h�è�(�ٔ��ɨ�9@k-D���FK�)�i��E"?\��#%+D�� 6�����8:v�;sb��(�|#u"O8��&� Ԝ8& �-��M*"O: a��5�A��Ё!�<�8�"O8�Pw�WP0x�*��lQT"O���.^!{^��KAoDQ�2��"O
�C��
#���v,�OV�	�"O�I:���"�9�k��x䞤 "O�]s��L�y~�l�u�ܟY�庵"O� n¸J�*E���h^�i�"O��Jc`yr��e!��~7���"O�1��Ʉa��L���2
��B�"Oր(P�ݔ6����2m��zm@E�&"O���2��e���u���p�D$q6"O*I��.�^�pj�I̚z
X�&"Ob5!�)e���ে�6>c>ͩ�"Op���M[-el�K���hS���"OL\�����&е9�Y_p��"Ob4SP@����}�2%[�-WD0c�"OD%�CZ�*���1�c_�Lb���R"OR�q&�Жe}���f��\Ɛ��"O�ՠ�d �[�gT8xC��[t"O��Q�d��
_�aYC%	,x*~E�"O����őR]��A$9-I��D"O��s���~K����B9?E��R"O,�e �%;�� �F��c����"O��G &9��Y�K�5aK�a˥"OB�@�"�aod�`��V�^J�Xr�"O�(��P�&hd+G��PN�A�"O����	��4�haI%h^�MD �C�"O�)�����f.��!*�I��"O�Ԃ�(Bn��Y8ǆ@�j@vy�2"O����H�C��eR� 2�hS"O(y����"��9��E��;'��0�"O�vc��+Ь�S�Q�9��('"O,ѰPI�t��x��eO0$Z=P�"OD��$�ʹ0MR}3v$���}3"O���才�^���0�,;2��9r"O�8Y�����x9y��cw E��"Od�k�I	e�5�cbu�%b�"O�t�!Ęm���t�ͼ	Q�p��"O�T)��ƒ̉CO�l(@=� "O�Y3��
-&��1ar�
2T��"O��2���O�^�9&�W��>��"O�A�q��
}�t�X��-?�2� "O�ӵ��,3�:�8�K]�3���	F"ORh�DMP�i��F녚d��T)w"Obx8�ߧ���dcQ
v���Ie"OF�SD	!c׀%���Õ �0���"O���q��=b]RD��eH In�@"O��Ԅ@@ò�0uC� 5��!�"O�x��̄�{�|�*TC��Ij�*�"O�hr Ǌ`!Q����m2���"O��J�'�6KghT	�gĖ|K�%�$"O�Jv�҈P.�b�dT�8��yu"Ob��� ��6@])f� h!n�҅"O��8F�X���	Ӆ
�Fy�Ԫ�"O h�V(�G�$���C!kV6���"O앰B"�D�|p�1O'S�	��"O����X�0�~�����ON�ܒ@"O8�q#��j����b$I�52Z%"O�����!6�����B�} ��{�"O� �pDC.T\���!!F`�*8�"O��'�zkt���/Za焥��"O�mz��ėeI���$��4���`�"O� L��꟭I��8�'#I�G�.�8�"OB�f-��D �%&�\/`���"O��K�
 �E*P�ч��`P�Cv"O��J���N�Ȉ�!Js:(#"ONĲ5�΄\�4��o��qmZT��"ObP3��ߩ�-1h��4|p���"O��b�n۔Jv�|�2���fR�	�"O@ �A�.Hzj,�&�&(W��p"O��A얰wJ���%g?�%"O �&M���,(W��8�Pp�D*O���H�b�)A1G����'"ы���'
f�҂
ͱ7�<y�'���Y`���!i괚Q6e�! �'l�-�(Z����o�7{U���F`$D�Dagd�)~A@�/ ���ɡ�� D������'q3�Dj� �!5��њW  D�`0�ƮY`��6\�
�b?D��!$�sͼH1��޷[�*�Z+3D��a��С/��c0��
`��M ��#D�H�Q�öP���aW.5���D7D����Μ#�@�z�ր/	 �`, D���t���s�lЀ7�H8E��!HrB D�,�W��+�T�)q@S�)�p�C;D�\���-g�>\�B���bhYc;D�,�sM�&j�xU�(�K��@J:D�������F
� "� �,����:D������n��Qc"�p$:D�0Z#L)8�*a8��_�W�x��9D��H5�@8($x7`?\אy�:D��h���W,6��GI�8i��7D�h ��)�Ȑr�>\{�`tC4D���f�q�X��f�U�X(f`�c.D�����xb��	�~��k-D��Xr�����%IU�4v㨽q�)D���3�ʻ��i��c�7{��z�J3D��ۆ&[�G3�KW��]X���),D�� E�_�K&@���*n�Xq1��)D���0Kϵb�&����A�ص#�2D�g�U�>��HxÁC�˪�a��0D�x �Y�0 B��#ύ	4j�{F�/D�T ���5h�BX��G�8��%`"D�0��J�Iv�k�l��b8 Q�l>D�dS�`�G��@���ɑy��š'@/D��1r�T�TT!*�
ڋ]F�ܠ�G0D�\VC��d(�Ps�%�kGP�h��,D�X��G |︸�Q��.�����+D�����Wa`ȂR)ŪFߚL!RJ>D��At̛�y�U0o�=BΈ1s/<D�0 p�g��p� 
C��)��9D�x�ᐫ>�$�4��x�{��8D��d�9'��H�=��a1�8D�p�ƆD�g
��hY�Vu���K;D���B�:0��z�I�8L�L5�9D��X�H�A�@h��υ+t�> �Qa5D�h��GS�(��7w�6�A�0D� {���,eФ1�C(хy�쐠��,D�X�F�/e����gMZ ���)D��������1@���u����h*D��K����;��ܑ�"��uS����-D��
%����h@B�9<��))Q�)D�$�"�J��
�IR &O|Y렄+D��j���=ol�SM�<EAtg*D����/��g� !q�� 7�Q�@�5D��!�h(N)(t��
�>#��Ѡ�O5D�� ����J@ܨ��%��$	`"O!�6��'V��yS��ʷ-�.��"O.ª�:��5��ԐX�bPQ"O��+�'�39�r4C�`S��0a�"Ol!Rd'N�y��d��N@�m�"Ot�Hd�]�*ޜ	�Ů*)�Uۄ"Ox���̧" P�F���I�C"O��@�r!xe�� R ;�Z�1�"O�E#��ݭ(�P�aFH�P�*�"O�Ժ�/��%�")�˕3>�� �"O@CC"���.���<%�"�*�"O~��H8+�����ٌ1k����"Op�����*V<��ӆ�lp欣�"O1�%��(Z{L�5Ywh��{�"O�q+�#2��y8�+��Y`i�F"O�dr���&�hEJ %����s"OX|;��3,�IFiK�v��E��"Ob\XB/X�p�X�*�'��CݮX�"O�eBTNP*v�(�Q�j*���"ODDj�fʭf��=82a�	���P"O��C_-c�FA�K�{��TX�"O>y#C�݅����	1� ��"O��"��/<p���hI��x�@"OjQ��
J?o��5Sm(/Z,�"O�i��6$��5z乓"O��X� �8"XۅI�lxe�"O�]�B̐P��E��bޓVL�k "O�є̐�i/|ܒP���L
�ly�"O
��֫ſe���Y�I�Y*�"O�=����Ψ��4/��:�U�@"O$#Ѕ;L��0�͖/f� �Y�"O��3߰D�d��So4�d��"O�]��ʇQѺ�b3d 3Sz�c"Ov�9c���!�� "v��> C �X�"O�qK�31����˂;5���"O����I(�ι���_#F(��p"O���g�#p7�< ��ñ7^��F"O8���Nl��J�(�g	��"O�,�"%�;����$U
�IP"OJx�����VA� 27�řfנ�7"O�9 c�٣ L��4&�
o��Ih�"On}���L�<��5ر��"q�Ơ�"O*�*s�TYb�9W웗zf�)a�"O���fLW�z<(��S-V�Ia"O�)0@�9� R���;UW,ؔ"O��ɒB�	1�T�v�E�VH����"O��I�*F	~Pcul��zF��"O���G	�p�" ��C;��s�"OtH�RF�C�.;7�B�Cz�؃"O�q�a���d!6��@�H�X-`z�"O��8cP.-T����I�L5��"O6mD�ΔS���uO �mb�Xq"O��BE�+C�Pc����ՉT"O�rf&�v���Ⲍ�'a���"On���I����*�BE�D�Lò"O�t@��)}�UQdc�ʤ"O����^!IЀ���-���"OBxy��?d(R�xѡVc�4xa""O�DX#Ů!�VPu �!R�b���"O p�@��L�=���?�:���"OT�B¯U��	0���qѠDQ�"O���k�s5�l� �U�2d\I�T"O��vצφh��A� v�"OVm�$D:&U��9�DY�3M�m9!"O� 6S�\�0t�5�%��q=,��g"O,�i��:�읣�R�'�2��"O�0��`�^��y!���Z���A"O$i��&W�!��$���RmZ���"O�ɘ���?�]p��:{�Ly!"Oʥbո�(u1G�>�i�"Op�"X387v)�������%"O|��Â�&G��X��V�i	�bw"O�t��L(X��P���!"O�])S�C<0Z�Ԣ���&B����"O��Q4�(��4�6.ƺb����"O�P��.��Z{P����k5.�+"O���6�9y���xfK@�~@���"O蹣t�ރT�6� ak^`0�"Ob,�B��1b|ɸ��ː6)�c�"O��y���1���	0%%�U��"O��g��4�S4*�$L�8(T"O�|;do��X�|IČm�ʔ
�"O�-��0D~�z6�_�`4�Y� "O.���i��w	D����T%�H3�"O8a#���
��Hi`�%-E���W"O�{�Eח`D�e*�D�%"6NMs�"O���T��?��ñ#,\2�ܛ�"O�$Zc�V|�����Ŕf&^)P�"Op�YaK���XP'�:K��"OH�J`Z9�nH�g� �U�Q"O���ɔkX ��G��3�B�"Op���#�)�.��g�e�>uG"O��$Ε�d0|!A�]� ��"O,ز6�-5�D� .��?lV�!�"O�����ĥ ��ࡡ�x�xY"O��ˑ.7X�G�����<�"OJe�J�/I��5��˖�n���� "O`����)h(dX`�Q�B�"�"O������F1��U�
�v\	h"O~�w�J�^;$(��4M"P�)"O��Ccg��`�5ۆb�X�
H�@"O�	:&��>J�<�!�\��̂E"O�4y��^(�0x٥�;ݺ1�"O\
&�GZ=C�%��)Ѕ�q"O d; �
D{iI�c�6ȓ#"O
����8c � ,��1a�!"O� hLKC-�`Q�K"��E"O&5��Qy�="R��K6ph�"O��iu�ŴKV�y+�M=a�H�"O��yW-�w%�a�5�ݤ��؆"O(���Lm�D\c��$�����"O<lsŮ�y�� Kޒd�0� �"O(�H��LAB��	w+;a}>���"O�,zB��Kݐ���9vNݰD"O��9��72]��Hj����"O�1P�F�]�@�� .����"O�q1E��?ؘ��瘤2�Z�ZB"O���W��Y���ޚW��uq"O&��U����磁L�+G"O��!s)�&g���l�.3��Z�"O�XZ5/[�3N:8���[9����"O85[����h;D!*	�8w^j���"O�� ʡv�H٠RA�#b����"O��P  U�C��=R���~5� �"Oܸ�e)Z������P,4H�z!"O���$�Y\բ`���` �eC�"O��(�J��h�bM�� 7	VY�"O�	2Ag��h�*�8�![�z��5zs"O� �q���g�p�wn�Q�.y3"O(0���<�<�C�F�2�s"O|�`D&��)K����w�\�zd"O~�80g9f��5�S��=��@"O�����@ߨM �g)%��q"OI��%�'u>�cg&�`��X��"O����()B��h�GB�o�ȕ��"O��N�p���$�f�P��"OB]��
Z���&��
T�:L�"O� �G��6t� ��KO���v"O���&9�"-���,'@&��c"O���1o��q�tn��P��J "O~5�B�T�W4��5n'V6�z"O8�"�[�T���L�3>�9�"O��I�̋*^IF$i!b�}��ذF"O )�u��#d<~M�M��"Q�R"O6�X$� q�6�a�K
�V�S�"O�]�tE���9��V1Ft��Cs"Ot�KK�)`� �dC,ZF��3q"Ol��V��t�H���Z�0�|11"O�����	%	4Mh�E*R20\0�"O��@�F�H�yK$Y�g&�Q�G"O�ie�Z�%�d$��P�fD�"O�l��FF��t
��ͺ��MЀ"O��� �N�Yj�#ب:
d�ؑ"O��k��p:dɢ�� %\>}��%1D����@(g܀Hps� 6i�n}
��-D���AEQ��p�P1�/@Y:Ç0D���T�X>Uxl�Y��:g�<��Ch$D�r��()lh���/(U6)���6D�|��-�}�1b�֛S8&{%�?D�4k�K�D�T$֍�!hA ��p�2D�\3�# �갸���7f��ܫ� /D���F��.k� �K�3� .!X!�!KX�)�Y)��2�c�l"!����R)j��́0$P��eDO5E!��%f<p�$j߳O�x�ڧŚ��!�N��d����B#�{T �S�!�䄱jO�(���S?z���G�Ǣq�!�$;�&�!��a:���F�t^!�D�0[���pG�ֆq#�e%M]�3!�d*Q�@u 2b2~(�q2d&ϵg����,||��_qaDz��R>RB�I�v+��Xč\��(�3�f�-:)�B�I�sʶᓵ��\��%pe�G"��B�3b@k�����=S$.��cl�B�	V�X���ԯJ6�Yir��zR$C�Xlp���#_@�+UdS�hZB䉤f����$�P�"� \���s6*B��@�t�Tc��<��#d
S�Jc(B�	�	n��I$!E�r�fp�S ]3�^C�IB�>AHΣq�P�
E�Y�C6�B�2,��i��F(pNdˑK#o��B�	Ts��{�jZ3�I k5-3\C��>�dID ��}�`���ό�� C�ɬ$�P�f.Q� ���!FʮLL.B���2E�gk^+Q��Y�ˤ;"B�I��ĩh"�8�Αq0O��2l*B�	m��8)�W�}��F۶n�C䉁Y�� ""��Q�TL��)�[�B�	�J]t�{� �:�\�@
,sU C��.�P�*�[�)q4��� 	��B� 4��`Ү	I��а0n,M��C�	�7�܊H $����(U��C�)� tY�`��jn0�y3G^%�Y��"O�S'�]�p�f�*p�"O����b�F< ���[-�L)��"O܈kt���7.F<p*(��L�!"O�-��')��M-!3���.Ƚ�yB�L���`(�#*�J 8#�_��yR�I�w~d��A�NҴ
��y������6AB�	�j���!�yB�R ڄͳBΓ�n�IR��G:�y2���6^0�c'ʇ�b=�PV舌�yr�@�? ��!�V��a���"�y����� ˾M�VH�s`�#�yb|(H��d�D��ҭC�yRHB�*��W)ٲ8$�e����y�jS;9\��FG�}�x��R�y�`O`�ۦ畀v�⃦��y�
���i���| r�jF5�y���V���*�`Q�vM&�P�L$�y2�G��|�E�;j)"�>�y2�͊/���鶥�4��Q��G��y�$۳f���zPF�9t�P���)O��yo!���e�� K#�yRE�EuN��珎<_Z�:��C��ybBU�u~���4�Ί.n����4�y�a��Q�'A�N�(5��Ļ�y�K��.��ј��D]�����y�HX�*�
�'� 4��;���y"�Q�21a��'��0�Tn���y��!cx����P�D1�sឳ�y�.E�6���O��F�Y��jP��y�LZ7	��X�!�$QΖ�w���y�dųN�xK�G�Nn$�V@���yRH�-Ur�ʑcW%M	B����K%�y¬��u�DY�s�?T�4bb ��yR�A�",D��nP��~��Q�0�y��ڪ	e��ђ��SPa
1�	8�y򋑝|6l�p��׬rq�졀ň�y2�8oV��6*�5n�ĩi�H�y�����`r�ޅg�:!O͛�y��с
�°����ZK�0 0&ݛ�y�UB$��Z?|�������y�ϔ���ݑ�c��Aj.�;���<�yR��]�H�@�B��3���GL���y�&�X� �y�Z7W��� ׊ߑ�y���+|#�C��WB�k'�yBCݧ$ ��&K����IZ1�yZ�0���?T��Y���?:���'s<h��D�����go�=��9��'��9��͔h��8��'�eU�Z�'BH�s�4�C�dܑF�V�'sZP���:��T1#c�o���'�T��1a�?��}h�k�"���'�V`R׊E�$�Ł0&�p�� C
�'fVY��DU�1��ܺ�l�a�N�

�'�}dL:T���qG�K|�aI�'�h�u��49�L��%��&E਀�':ഹ� ^�z�sb�����'<RЊ�"�_�Z�P��$
�R��'�
x�ϝ�D_]y!F�Se�a��'9���@71#8]�� ޛN����' i8�I@9QO��K���ZuP
�'J�A�/�(3��y$���V-
�'�x�ÇZ�<��y��=Ӿ�	�'�2@@�oRc"TACHOQ�B
��� Ё��>Ԃ{c�}�b�9�"O�` ��
�6���S�P|��"O�(C怿EJ�����|�b!C"O(�KG��#j-\4���Q�%�1� "O����N
�9T�Q��2����"O�� �JɥJ<BԻ%'=y����t"O�z��l8	ֿyX��R3I9�!��I�:�)F��M$BmW�a�!��<.e��!6+�91�V0r���:p!���"p4��A&Ɍ\�P�q���H!�Q�~�1A.�.���
�f:.�!��c��@R��<@�>��ڻR�!�dE�`$��NYG}�h�R���!���h�&�QpJJ�Y�LΥ!�!�$��	����`C�T��\��J�m�!�6C��q6��z��Q��W�!���5����LM�'_����F
�!�!�d܉a�@-
7�
=QT���?|�!�$�<T�1BQ`�3c��d+ĞW�!�dԷ?N�XpM$bYթ��+����3f,�Q��0'	�Y�'��y�&�?G> K�@�'"��0�
�*�y��ef�<C򋌏V�C�e�y�k��ylXt Λ�~Z��T���y���xgeX���'�ԳvL�/�y"��&)^���!���6�:f�\��y"��������f �𩘁�y��N+,tp�z�jM�8�"E�g@G�y�E"~��"�>)}2� ��7�yr�U��ڐ`�#.xf�"�mʝ�yR�A�LH�d�;)b�8樍�y���<�s���?-���B`�K�y��� !^���%�O���M[<�y���/MI��o��:��5  ��y��8��(yQ�R�HyB���J��yB�݉NF>tk
�9�������:�yr[�E%<D���[����ԅ�y�k�p�;E�4Vo.���N�9�yrOO&fA��s��!H0���Y&�y�1Ut�Ƴ;PހЄ�0�y��ܜ:��xB�ǁ-���W� )�y���"ܒp�©$Y��G�.�y�,�)nWP���*���d8w��	�y� �1k���� .�
� Y�C�0�y��u������ ���Ce���y">J��-�
��th+��T&H�ȓ0��u:Q�L�%��1�ַ	
�ԆȓbU\ #�
�Z�l���<#�	�ȓ�Ha aL�blt����6MP�}�ȓN���@�e��(Z1���2sf`��&^�� G��xj`	��Ey����p�>�	U���%r�B����$��gv,! �^��-�-��m<��ȓH��B'�7O�ɂ��11���ȓ;�Ta��"PoԸ5�"��*B���ȓm�J����5(Ȑ=x���CJ�l�ȓKP �# ��i(�H�3Ⰶ�<t�Y�ő1��� �*^=Ԇ�f�ȭ���U�k<L�D!��{(L��D�x���į8���AfO N�ȓ+���Pm
 N�Qp�Լg !��m͚�T�׶= TԘ#C����l��ty֧�}�2�#��"xrA����o��I�h�Ă֝F�����l<D�� �a� ���6@�d
Tg~_�D�&"Of� `D�	�]y� �B�E�"O< 0�l�is(M���!?ja"O�tÉޭ0���� �/��R�"O��"�)��PU�g)��E�t��"O�P����X���gƓȖ�bf"O���4b׺j�ze����(�b�"O�	(֡܇���2�4?�,탔"O�i��OJ
EW��s�(D�+��uyt"O�����I���#�!�k�T��`"OD%`���%q:�ur`'	5���k�"O�Qx�E�Y��@!4�{ߜ�+"O"�JF���%e9T�l�3��?�y��D�!
����t�XZc�Ŗ�y�����V�)�g�l)Н�����y�$�]�:�ge��5ȑ�@�yn ���qC�G�X�2�9a�#�y�L���x���ؤQ��ܳ��M�yBI,~��T���d(�y���L,I�V-X&z*�X!I��y��� ܤQ@��_��Ű�e^�y���>n��hyB�z�tqP�盖�y�*J%Z0���c� ��G�ٍ�yR,�bU��8�C���1��M�y�F?LRDB'��Ͱ=Qܐ�y��6e�>Xx�iZ����6#+!�� �e��� �'i��dB��7�!�Ę	N����D��5�f݂D"OZ\#`�+4�t\R"'@�^%$�QV"O���vl�����ҋ"��A��"O��H���j��|�j�5�F-"�"O*eR�i�1>4)3��I�h0�G"OB�+'�HNo�TJՀ#���"*O�%І��HaLjH�<e(��x�'��0�۹k�
=J��ڔFg���'�XH��Ѱ]W�#i��9R*���'˜Q1�▟�n�x�Ã �`�@�':vL�7DҔm/z�1��K�M��
�'T){�� 9����񠚚rG���
�'{�5��̌\�Ȑф�[�fT��'9$�H	�"m��I9���@a|���'�r�#$��t�,���L5�J ��'-�,���N�h0�(Фy�@���'���薬��|�䙠���r�1�'�� ꁧ�����du��s�'�x�k�E�&�,�`R�b��P�'W����'@� ���"TEr�{�'#��d&�� �C�p���'P�B���&y�
� �������'���ƃLudt�j�j�rP��'�� X���	]Vx��B�0-]
x�'�Ź�I�7Z�X&KD�V�����'�D�h���H�F�z�-�#P�x͒�'����j�v�0]ZT��O9zp��'F$��e�#X��)B�/
�v��X�
�'��h������Ԁpm�g%N1�
�'$��{ N��U�B.�X1�9a
�'}��3�hHF��� ��T(U?�s	�'#<�Q���p�"��$dL�A���'px(a�V�ln8,K�@·+�L�	�'�.�{�B�A��YƄ��mh�d�	�'�ح#Gd9@-��s�蝨_�N�	�'�@�s����e*AJ�e��^(��)�'�&d� �/f�$ɥB�:N$��)��� ��z��މb�\�2d�>��!�U"O�����ޱ_䔅ɰ�<�9r"O�a[�A�IH�17#j��"O$��`C�R���S��	$\	�u�"O&�8�Jʿ99���[i:���m�!�D��e��\�W�?XƲL�D+G<(�!�t�$��u��;=U"��ӫ_�!�!�B,%@���g ۉp�B��W$�-N�!�DϢ�b���������#�	�!���A��PIB���B��5�W[a!�d�g�"i�fH�N@B0���5D9!�D˪ ������+��!��$�"���I� ��Iu�̉s�!�$�/6��:�-Ǫ6뢌��I# �!��V�2�0�ܽ��� \i����>b�,J��JMr�g��p���ȓ�F��%��Z^l跠R���X��K�z���	<�� ���OW��c�����ŉ<�L(ÖK�7 �h�ȓY#�ذRd�^fr�j�dɥ2���ȓB����-O	A���n� h����ȓJ=�t�OY�[��*�k�=�Մ�BsKʿ0y�!����,�� �%?D��+g�U&>�Qy��J�;l�Pԋ:D�0ar��oS��C�K�)ax�(�6D�<��N��?�Hqs���;q~l��6D�a��LBj�ݣT��sp��e�3D��C&⌳=�L|�SC;|.���0D�X��� <1��#�ī+	�h�ǩ3D���7.�'D:��d���h�Р<D���En�$6�$ڲ�8&��T3h9D��c�ꓲU.�(�q��'cBEk�	$D��;B�b���㒈�=(���C#D���p�M�
�$)��͌T�e�+,D��&�Sh�y�sH�
P��rJ/D��Iǎ���9��&��7�iPI-D����̖`�  Zv,D�DOf�t?D��G�V��8��-(r6 �=D����^-��*���
��h`#h:D�P�T��lJvm��\P��YBI;D�\�"̌�/2t�`��dX>�Z�.:D�d�� �J�<��bG��io2�+6o6D�4#�dO.jP���)F��St�4D��s�Z�ZC �r�鞝u�`��10D��d��
b��d@3n�w$𳢇-D�T�R��	r��ń�d18����?D����ʮe��ʃ^8��m<D��ɰn�"Fm��D=�6ъS/-D�� �� $$�\��.�/X�*�ِN,D��"Qi�&L� a�	A�4�	Ȧ�*D��Ȗ����LI2�Y�#�$D�X��nϴ=���SWꊻM`>�� !D��q�S�PBQ	���w��� D��r1Kξ�$8ٴ�?^g��82�+D�(ᕀ�w�P��@ E�:��4�(D�(���8-1b%[�9�
���d,D���!A�(x�ł�
@p�?D�h��Q5R�f���a�@o<D�L��e�/xk��	���#=�"�hb�8D� ��D�0.�J�3�<je� !�#8D� �d��r�>�ӕK�������7D�<
�	�e�D b�`�,��5�*D�d�kщ0�s�Ȉ",�}�R�-D�4#!�����Ē|�x�@��>D�� ���G�M7���C ]4z��Y[�"O��3$Ȁ<�"���f� ]��"O�!�"B�M}�L{U�B�h��T��"O�B�O�8R�l��̂�||��"O~q�p�S7:
]���șy��)�"O���q�H�8!(�����xd��[�"OP�ㄪho�����&a^��r"O������
�������&.Snq �"O��b�L4V�RC!S5JNUi�"O:L�;�UZ7�ǩp�[�"O0ijA#�.9��XP.ϩR����A"O\qkрR�I�P��m�H��/�M�<�SH֠8_�q��+�~P ��a�`�<��?c湲�L�]�9��YV�<	�ѽZF0�`���m�,�C� w�<a���_�N�B���V.Ƹj�/�N�<������H0vt�I�&HJ�<��F�a�J����N�Y7����^�<1�G��N 
d��{�P�	s��S�<��k̻���ւ)��X�e�LO�<����X�Ĕc+��i�Z�NB�	�f֭��-&E<�2�Q�csDB�"�(��	�&`vA��j��B䉊mඬҷ�ݹL�j�7��6$C�	������Ā}/I#_��B�I%!����¤[�z�Q7G-S�B�I��4��S"����Z��*��B�W����Ǜ�JM��^�eU�B�GHDȓ�Iܰ@Pν���$QږB䉽z�~�	��̑9��SuY�C�B�I�}�"xzP:j��0�3�
!�vB�	�z"�`���ɤ*DÐ�R,��C�2Y��Z�B�6_�Xs@@�%B����O�{�fM�#�˟�@Y��.W>t1!�������R&�ƬY�Áy0!�D@+"mEZu�Bhj5Q�,�X!�$٬}g"�"N~�![��v!�D�2��\#w�LT������+b!�Ą4>���e�(x����+��PM!�Jg���Sb�Z�*����K9�!��	�<g<���!���;��&3�!�V
$���s�[ t���c�!�$��h��(�蝱D۾��mQ�X!�D��C�2�H�d��.�y��#8<!�$ ��졕 �>��8�dN�x�!�7Yv4q�����9�R I�P��!�O4bz8<y�/�;�LL�@�K+T�!�Ę	&e&a�g�S�WO����b"w2!�$R�u�2��cNӚX#(�с�X�fJ!��B����7F��֝��@6�!�dҤu��0�ؕ0H���]�!�D��4��#g��8Z�Iv�#�!�d�a|v��s �
]n|���7)�!�:�@�:�nN�|U؉��F��w�!�$�.y�A#�f;FEx9[�KK�#�!�$�"8s4 ���)��}�Ʉ@�!��G]���Q�Z���v��<�!�$ш3lQba�B�1嫜?X�!�d�?#�����N6���3ʋW�!�A�*E�ѭ�%"#t�!��'93!��L��m�BJ�9st$E��I�T!���\z�4�刕�
��%h��?�!�$W>]��Xs��6�~�Kf �sg!��9R�Q�2�]����! ��!�� 2I7%G,tc&��O�^Xw"O��ҭ�e#�C�&�N��ӧ"O�$
�H�z!��ȱ�	�T�2�"O�Q���1D�S���
c$��%"O T˱i�D�x����Lr�=��"O�ȉ5�S0:$ţ`����i��"O����O�x�銐8R �"OV�yU%V�&��0M P	☓d"O�H�f�
�Z`��2ThdĂQ"O�A�����H@��N�7`Z��3"O��*!n_"P\|:�B�)r`r���"O(���D�*%��pb�ͶXV��"O,��V,.���H���/���+�P�<��S� �T�0櫍�K`<����N�<C��R������F�XP��N�<q%A�[ ��fI��H$��s�<��,R�1hq�qeŝ.�5�Ӎ�J�<Q���9I�Ԭ����>@��
�^�<A�K����К��9���F�[�<`#R��4Bv��^ 䳃�Y�<��dT&3?�Q�BhVi�> �D�o�<y0�Җ>�Лa.�._ډ`��i�<� ɝ�>�
=��}��Ȇ)�_�<ϳIzz�R ��w��h�7ϟc�<��>�L-�fD�0]ɠ����^�<y�g�s6ht�����lƌ���NVW�<�ucУR���aD��Y_���R��x�<ir��5g� h�U�WV��(���s�<QsP0Y"Dٲ�c��x��1�w��D�<Q�+��|�
��͊�(�d�iZZ�<�	3v�I��]���CC�R�<���
*/��� �V�_nډ[�F�v�<��i�>r ���!`�sq�y��n�<�@�R"�ٗ��\/�݉#�i�<) ����DB��ɋ?I��Y1��}�<���g�~И��zl0���
o�<�բ�6f����
O�0]X�K!cLn�<��u�t��cۑ*�P%K@�<�ׂ�t���A�BK�H�X�e�V�<aE.Q�n[���ώ����xg�U�<Y@b�5(��`A�I����h�ʞP�<A�lķ$�����l~x��p��Wa�<q�ƾ=�h�ZWÔ>�|��M�_�<A�ȑ�bh�m�E`D��$��^�<���̇{��H��Dń2�����E]�<��� [�D�b K��ytܘ�Tk�[�<��OL�%aba���P�������B��;�ڕ��f�=��Y�pc��B�	P��BSH���¹!#k�)36�B�Y7��e@6����C�n�dC䉐A�V!`�"ڶ�x=a���,\�bC�+������m'Z)*�&Y�~�,C��1ZHBa#6t2i4�Q? bC�	�j��x$��l��O�.nC�I/Hf	2@eA*%��;`$�!vTC�P	��+��1,���m��&��B�I?E@��:�,@#0�����ϖC�	�}�)9��ǥW�xA �I֢\�xC�ɴ
s�4�0�ۂ'�F��O@�U�vC�l:�j�싿�ک�RoH�/k�B�	�_��R��֞h��d�`�PR�B�	?|�P=X���*:�i�`a�'p�C�Iy.~�s%m�7A��Eҵ��\��C�I�a-R-X"���v���C~vC�)� ��s��R5�M����4	is"O����E���5!!�7>dAA"O�pK2�H?4�ޝ�%��-g�HH%"O���A�]�hp��!���d"O�Ը�cͧ
�RU"֍72Y�w"Onp�S+�5�� ��Y�P,�!��"O�Ě�`��l���+�6�i�"O��9�ׁb�ƌY3��Ꚍ�&"O (!Sb�A�F�p�cR�ް�%"O� w�K�
�]�E��(�`A"O�0��,K(L=�ᱣ_�O���"O\D�Bȏ=Z�@=�u�A �.d�"O`�Ye� �;Zq�Wˑ� ��h@f"O���i�6w$|�bj]�)�`'"Oб��N�-7���5�����%�"O9�C+��jM>�P˔�H�2��"ORY�@k-F�Ah��V��{7"ORء�hA��*��מ'sNhf"O�Ĺ"K�U'fÇ��Aa���T"Ob�*�I؃]���v��4z*q�"O��t�׮�^�!``^S�Ą�&"O��҅.I�\�]�a��W�h��"O�h� �N�]Z�M��Đ��e�"O� M16h(9Q����� [�"O�p�_�15f��֭T�V׆�e"O��4DH)tt3l�T�`�A"On��bGJ��ӷ�Q�t�N�I�"O�ؑ��v�Qp���]f�0�"O�p-t}�$�+qu��T/�8HL!�?ֈ�)�㉋U�,�b$_!���/���UG��T���$$!�6	�t��u ��A�
�ʦ�	?Z!��ES���F�z&�Ͱ�� !򄐿"���i��|�
ӆ���!�SiB�Q��+f�@��C�\�!�ބ2�`1mP���qr㐄�!�DٴBԢ�JOK�d��Ѣ�5�Pyҥո9�QrGȞN�� @���y�ίn���s�mF.v���!l6�y2�5XZ��H�o`�m��EL��yRa�7�	�R�	t�Q)#O��y���,�m��Ҟdx8�t�@8�yb�{�^a�V�גtQl��R�T��y�E�zM�;գ�k:������yBȂ�-��Pصj�"o�Б��(ǔ�y���֑+`��ֈ���mH$O:C�	4��qp��sf-��)��XC�	Q0u3e�	Cl
6D�0#XC�ɕV(�sB�;X�P��W �.UtC�I'{�h!�OT�F�DX1�J]<As�C䉼6��p�F	R=�ly�b(Y��C�	\Ǝ�1�W�2��0�è�9�*B�	
�ȘV-^'x,���蛅{ofB��/n�(�sK�^�z�C����8`B�I�]�x�ҰIS
b�X���*�H^
B��$f|�92�C�+�R狝�MB�ɰS�Z�sƚ� �3g�� �C䉔h$���L�b��� ����XɪC�I/7�܂�f��B��!�ŲBǈC�Ip�8��� ,��-{fC��|C�	Lr�0� ..Pd�P@� �#�fC�	�T�D�S�KG�|�B�2 ��9A��C䉾+o�ĸ���	,�����'"C�� d�Z����qsءto�Li�B�)� ����ͯ
�J��z�r���"O(�Ve�#nL���$�z��8`"O���k��V�&��̩���9$"O�0p掔���� ��gHn���"O�0I��:V��Y���,V>eK""O������`��@��
IE(�1�"O
L�b�/b � � ϗ�3%tlXr"O��xu���#Q��)Ch�!M!��"�"O��� ���5z�H�����S�"O��aB�`�Y@���k�ܰ�r"Oz�s�o�*��䨥�y��y�"O�*_#̈�1e�V��9�0"O���N�!\�=�"%��a�T"O
�[ǊJ� ��h3���!()h"O@25�r��X�C�2h�(�"O�4Sp��<{������z0IA"O��Pî���ęҏ؀n&��i�"O�xk�FE��pQ��O�$n���"O|�9�H�&P9Z(�q(�*W^�5ce"OxҴ#�49�+d�2KxT�Y"O@��B$M�~4|�!RAL�'sĈ!�"O�U��I'�dms�Fr�9��"O�h.\�E�BZ�ڔQ���)(�!�\�I�p�z�n� Y����Jtx!�䝬� ,��膧c�<#��	H!�ċ""`��	+�9*�,ǯu!���-	LX`t *L���t�G�L�!�G�x�H��#�8y�D���)�,|9!�$ݲ$�(�!P�_�Y �LQ��\�!��ݚ\f̻�$P3i���Z���n�!�DR	�A����1�5�a�D��PyJ�/�mS��ƣ�<e��Ҽ�y��r���@�O��&��&��y�� ��,%+�/
�� C��y�A��7{t��*W�^=��KD��y���@�"�G��P��T�y�G="E����N�WnF��D#I��y��w��؆���T?�TKS � �y蝝X�Ի�lL���br�\$�yb�I� � mk��ԠL���Bb_��y�d ���@YF�OJΈ��G�?�yb��EAp5��ӭBWR�')���yb�S*[�*������?c��Ƅ	8�y�A�H���D(��C�P��	���y�HV�\'P��E7;Fh�"���y�$\ �@�I |E�Ր�H��y�!�	d��H����1v1�`s�"*�y2&P��	�#`V7Q~9:�
I��yr�N&*��qh���*/�<���C��y�E�x^d�R�*�2+.�P
>�y�,٠<,��2>.����[��y�fN6Wj���B�D�4�V&��Py�j�9Z	�]�AO�r�vuːiRc�<�U^��|t�F�ЖuG.��Gt�<Q�cYw��rQ!ڪg�6qAs�<Q�"J��28��JQ�@��whLo�<A`E�W�HE[��"ݤ�"���l�<1���1c~�g͝"dԾ8�`JN@�<G-�ib�E����I�4��R}�<�U�4�J����=�� ��r�<)Ջ�	� B�S�O"��I�f�j�<����d��8�d�:6IJ�)�hh�<G�ßGopT��R�+?���z�<���U´Y;p^����0db�<� �����3r���¤�U���"O��x��B�q���p"CD=79�"Or<(��C0UV��r��!�0��"O&�����m���)�f��M�"OH�L,OS$MYL,@�(`ӆ"O�� )��j�HYwoF����"O� *�	ղ/�%�b�Ǽ(���"O�9�Ј�5R	��֥
5[f�!�"O�����͊:RBK�Oe��S�"O�(S0-Ą#����K�1�"O|�$�Я�U肇�;sG���@"OF���	�G�|�bF��Y3��"O�ݓt���N�d��TI<K0,��F"O�$���*F��u�(�2l ��"O��R��jf<�@��P�*���P"Op��4q���e� �p1�"OjѺ���6A�T��B���F�r�z�"O~hS�*}�k�+L�>Qr"Oz�#I�Rw>��5k��q�0��!"O�����cB��t�۠ �؜�e"OȜH�+۬I�h1��Z�̬�A"O�!YU�śHx*�i�L� Ty"O���r��w�(�R��$�t��D"OV��� y�&u������Pz�"O�mH�H�`$���J�E<,K "O�q��`K�5�^Jé\�&b�b#"O���! ��Ud��QbD"Zj��%"O����]�A��yQ�둋"^�6"O��bàI�E��8��	�7ZF��"Ot���c��\zW�Q�W� ;C"O�ĸ��9x6F9zC�����f"O�;��@���S�e���p"�"O֐X�'Rʸ\
��±�c"O4�K3�#}��c�ĿV��"O��Yn</|h=x�f�$P��Ac"O|��B�U��zJ�fCDf��R"O�h���1	h�0*��%�r]0'"O���&e�K�Z$%�:�e�3"O"q�Ԏ740 �r���I�-��"OdIc�-H�fS���6�е=�i��"O�@�̓
Gn����ɻ.�*���"O�p�a*K/f�.�3W����L�`"O."�H�;��i��lT=0*�"Oz�It%Q��ҥɃ"c.�K�"ODL��o�8,M0��	qְ��"Op9(]��h��<�6���"O4�B�Ä�}��3�N��r�P(��"O�!@r�Љ~s���χ�x \��V"O:�3���;�1� �	�e�2"O�+���-O�U�+�0� ��0"O$�(�D����+E�!�Z��s"O�9��{B��*Uɀ��"O�J&�h�a:@�6��""OtE��E+$��U�w�/o�H�"OD����5�2PB���@\��0"O��0F�;��Ԣۭx��=9 ��d�<AW �~I�u��-C"0��S�Z�<���!(�޸2��C'91���`�X�<Ɂ�ӧ= ����o��� OB\�<�􈑲aB�(��B�F�&Nt��	ux ���%o���;��յx@*���b���l�n���{q)��;)��l@�; %�>"�z���-�r�X����
TS�iN�Z����Ȓ j� ��S�? H��� G�..��CDV�/�B"O��RwH�.y���W���:�p(&"O�H�� ;:d��kW�[����"O�8R��>w����
V� �)$"O@xL�	l��Q��F��-��"O�ء���-G�D`@�au&)��"O�������w�Q�F#�cDؠ�"OZT��̓_<8=ڥ�]D���26�'zp%�"Bh-�)P �,5����!Q�I�	�'��ZQ)Ag��Y��kAT6�\
	�'#���#�� \�x��I�R�Y"�'���@��Wvv)J�)ː[#�1��'��9�A¯������T]՞-��'P]��Ô'cZ*!X_�K�z1c�'W� �޸-tP�P�j�3��0�'jR!��G)S�z�r�$�����'�r`�* &78<aƪ&q��Ai�'sJd1�EClꅎ���Y�'+�t��)�?8O55��W3N�
�'�6��hW��\��Ԅ��L=��K
�'sh(8gJ��j��vΝD�P�	�'m\M��l�0�@���W� �)�'��h����\fxPG�RT�h�'V,a��J�M� 
S!+f���'���#r��H��iD���a�V<��'�X-��e��R�erD�V�U�&���',t�(��U3���a�W[8u�	�'U������P'p�� ���H-�%��'�� ��f�xQ�ç������'E���p�:Q�����/1�t��'$$9I%���'K��AD�Ѭ8h
�'V� �tF�*K܆�����)#DEMR���!3��L�:w�A��L�o�}�<d��c($�r���#[��(:h��ƙC�/�h�,�%	O��0?��hR6/��:v��b�t��gbFQ8���cHXC�5�N�<!5aL�t��g�σ2[���Z�<YE�[2�(�f$M7\F�����V~��H�m���a�/��"�2�I�gM��U��|:�
0HU�<�����M؊���"T~���x��Y(K��q���x�`��KN�3⊡&?����K�<"
D�qb�eN���D<�O����K�<6��!���2D�L\ 	��V�x�;�h� }�r5[��'r�p�DLM�0��c���l#�tQ��d՜,�2c#�����[�-_�I=E 4t�t&P�D�� �։m�!�D�7O��4
�`>'�a#$I3B��I��D�\�סj��1ֈm��>��yZ�1��۔���&H4�C�I�ʞ�h3�M��ɇ�S+m�d��1��5"��
ڑ�(��V��?����L%YYA�'�/�n! ����6Ma|Rk�~K��QFR-(�4�0W��hl
=�*Qt,M���t~8��&Ps8���l[����>ۊyc�f �	�n(�X���O9�	�7��0{;�	�~�����X�(t��!?]+��ڒ"OV	b$Å-n��T�g�Zm-�EH� աE:H��6��'{ݺ!�&�� Zr��	a��p�O��5>�U'��u��P��!D���n_�`����W3h��i8r�ޚE��.�遇�E�n��]P�E���:�	?/�^Lbq�ݜ\�,�s�ǳ`���^{��� F���yQ�����$���w�܋3Y�4�O�y�N�#"	Hs����� T����т;;��B1�X�~6qOb�8�Y����&/�K��I�eW�����,��u#��B8�1p�n�1�ȓX1M�J�^�D5�tn�9$(�X����n�*q�%�� O�إ+"��[5
c?�h31�Lầ#�7G�$��>�,�"O�m���߀
Dd#Ԏ�<��]����>��9��$ �E�f��H �e��.��(O�cQ���4�Z1�� ˺Q���'�4B���1i[�1D/&g�Ĉ��-[@�6�YP˕�m�pev�͛lӠ	04-#�O����*-�ɒU�]&&�����dEN���0�0;V.��r��Cn�EL���'uРm3�@T?;IL�	W��0S��]��S�? &��ԡ>D$���9
���(→#dV)��ēU�X��0�J#n.���#ڼK�����Xv��C�v��eU�<ك�V6f: �aMG-l�Z�>nfaCCQ=e��(t�*fW�ٓ��e2��@���:<�D�V�B�6^<#��(\O�Y�pC��h��˥"�1P�"27j�ʠ�2 5�m�Fb�.�1kC�'��z�瓥0��_l�t���}2g�'�(e�C
�L��Th(�~r��'F�2���� +w�,���M���x��LT��(�e �d���$iI#WC�u����aX
HxvNJ�N��<b%��g��~⤉�)aЕ㕬¼o�R��Ǐ�yBƟ c#��$�_(Z{ڈ`0DV�yBȡIV���M�0=��@�	ZV��KR�+q�mr�APJ8�p�I@+:-d"K�Rp�IR�E0��5p�H�*{!�\�
�Q%�"M�����e �r!�D�>rD(���"-2A�c�!�d���	s�aѴ�v�OH.r�!򤁗H��b�-ڞrJpJ���!��8T�-3�H�\&l��-��&�!�D��qʴL��`;���r�ġh�!�dZ�<�Rd�w'� }Ӵ��a*Z�!򄉺}�P�&�l�Z$�B�ɔ�!�@(E � V-Y�2�X��b��Z�!��ڈq�H��WZ�2�h���{y!��g5"�& �l�Z���AN�mJ!�d��(��������A�z4!�W��t�;5)�7y��$�!�$�<�X`�#���b��:!�$�x*�q"��63�R���(	!�d�*E��3��6���K�g�T�!��^�C+���6jJR�rD ��{I!�$��A����=t� pCG_!��t E�r��6{@H4ǜ7�!��
Lj,9
��)N��@
a�!�DH���1`T:m'40H�f�D�!�d��m���wn���BяK�:O!�D�dc�Aw/��O������Ɩ"'!�U-��mW�0���2���n !�Ě�_�>e���H�7�����!��[�!�d�2��`Tn�,תd�s�U'X3!��ؽ?�ؙ8�B�\�bt��$:!��K�"
�X�V�mu"FL�b!�)r��2�ȅ{��s��z�!��H����H��_�������~�!�D�3z�  ��d{�(��M� �!�Ē�(�B����Wi��;��C2~�!���[�*j��I+6K�<Iq.^9A�!�D��zI�Hj�f��|N� ��O���!�$P4��P���B̖���MP�2�!�D�=�:9ш�,]�N��`�;Z�!�D]8p�ށqQ-��9�\�aug��!�$Z� �(�#"#�	�ћ�&�-`!�+s��y(�-�(��
v#R�l\!�D� kXTظT���-���q��'V!�$�!f/�MKqA@�w�is�ʾF!�䂗tޠ�zW �l@�1g�:n!�D ?���K���B��X�	7!�U&�������&�(L�tG	w&!���(T"8gi��l�C�ɋV<!�D�"f%�E�v��&͐�� I�J!�d^�x��1H�%-G�I��VS!��.v|�\�UCڝJK���� �zc!���[F~ �"�����Q��ϛ R!��D�\z�����H:r���� �R#QN!�ȅh��iAA �3d|��#�,	V�!�dՋ���Kpe��Lx���d�<G�!�� �,;�Hgм���*�U��"O�:��������K٢B�a�"O��Pa�)@���*Di̜)���ل"O.�8��(�0��7u�rej2"O��	S�00F���Sَʹ��"O ��e��G���*[δ )�"O�AkH;e�C�	�U�|�0�"OB�.ܢ}��#P�K����"O&@���Q!O����EL�v���w�'��$�YpX�hJp&
�E��/�z�jZ5�2\O���1Ş*[�RE��'�0�B� G��1�D�:޸�Q�'�]Ҕ��(}��j�ū(Q��CJ>a�+)U��c��%L�^"}RትOlF�A�+J��$A(��Ue�<��LI#xj��	!��T8V��#,ɞ �W!�1JS���b�P,�~&���ao.|r%�f�E���=��G.$���d��t"P��A)_�rP�7f�<be{G╛��A�q@GE��(�ŦR��������![:�]z�-O:�g�?`�|��	��4�d���*��S�60�aɛ�P&D��V�yR���,vlAg�Q�P�5	�n��I#U�S��\$?
x��e�,�>p�	# ��}�oFwǲu9�$"D��)��ܺ���+G2d���pw�'�ޅ�am]��v$S�+ُt�,b>!'��"v�I2<@�Тrb��H#��:6AݵH��5����0�H#4�$�E�Į�1~��i���@7���ɊL@�BL^�G�ج�bCު)�����`���v��Na��'"�q���U(�˖�G�*�
��G�04�L���C-9��QT��
^�iC�=?��(΂y �h3fI�? Q�u�^���O=� ��	 $���k'%�0�A��'�^����D4�dX3)F=y��a�H�	&l�4�N4�dĻkO���O��'.Q)-Q&� �qf��=w1d�k�'(AVk�Zd��)"�O�c t(����86������ɟ$��yf��y�o	2�(���_D�9
�!���0<��&�v�(�r"���	xdy�g愋h�<��n�;��@����VҪd��'���]q�Hg�ظ� J��a�nT0r\���4b�|������,b�O
��Es�߫FYzB�I�cY,�#�C9>*BXv	8e�`5ze��;6���TeU��{�6�3�䈑'b��6X��8�!�L!��I�*����E!+���$*,��Aٺ^z�B�s����D^)/2���A�|�f����ay�OC� �@�h��_�v/T�;�E��^6$�В#¼�p�@OP%F`B�	�|1��E��vk.��*�KV.�O,��J�IR&��'#^ �H�4�%�A.V��r⟴�N���"O|��G�45��1�� >ArT�����]{�DCs�>�Co �gyEʑ�l��ʎ�q̜y�V*D�y�'m����K�jC� �E��?�F���&����+B�0���6�P5����o�!���uV��� �\T�� �&a�!�D�L�ҡ�uU��3�o�B�!�䐒)�`�ӄ�Ì6H}YсK!��u��)3.'a#����!�!��f��uS"��|`�X&�L�!򤓸,��� $9}����0�>E�!���>C�p�Pr�>d�<����a�!�Y�ڕ�E�D�`��mJ���C�!�	Q�H�IA��
� ���U�!�dļ`�0HFH�d�ؕ��	�!�d@�H$��G�ڟ��}�W�Y!��̓}���s�v�B�P�8X!��=�4��'������w'Z-#M!�!�V��U�׎ ����F\4V�!�WRJn c�gY+Z��Q���t!�$�'HP�GUZ��獓Ge!�����q*��U"W����F��-o!�E*khN��@ �P1s���>�!�d�8<F���#SҊ����.�!�� b�����\8x�у�H��p�"O���qj�W�x�3B
���"O^�S6�[0�&���� n��t"O6D��n�:	V.�:p�cS 1�r"Od<� ��?g� p6��DqQ"O���CˬP
�z4�K�}5p��R"O�a���C�U: `a16�W"O�A���Q�3z�h�Eg�G?zI�b"O�a9���;'I<]�ch� a�yn!�� ��`����:v(����:}E!�DC�v�Jт �r��i��K!�d�a����!GH78q��$@	M!�2��� 	&�x��!]�6؇ȓ<q̰�"BW�]`��4c_T��I��6ATP�b-^V�ir���yu.���Uİ%��/s{�i�r*��l�ȓa@h8�*opp�$DOYFB]�ȓ3h��'�N�ԐA�b���1İ���0n��b��++hfS'���z����"��5��+Ng���d�:;�"��� f� �D��ja�ʆō�T�"��xޘ���H�m�r�V��C~����2i���F�˚U4�	f�d�i�ȓ1�4�pa�ƣT�8����u��~@h`k�\�A���1�\:	��2 jxgΕ6�w(�N����b6(�{��Xx��0a K�oDDQ�ȓ0>r�q֎�|�H���~ߤ��ȓ3�@�r���AZlݩ�\�{Xa�ȓT�n`�Uđ��*ـ& �-��e�ȓG0`��3ı������bJ4���O^���fǘq����0��.�~|��O�#r���)+nT�)]X\��NO���p�N���P�7Y�H��ȓ+5H���W::|$p���ѷd�$��ȓ&���)/V)��f��5K�{2,(��5I���O4*E�Ywa<ݸ�e�<c���B�ON]2E�X�	b4ч���L
��abڀR���� A�S�� �v����dRH	W������ O L�É�!"Vq[g_���%ЛZ�f�bEI��gN��q�?D��R��S7Q���ʒ�	�u�Zl�@a<?ѥ�M�e�N��pA�9T��?	X�]�p�6���EI�#wR,�0$/D�U
M�<Eʥ�F�ya|)�QׂT�ܔ�C4Oh<�w&� b��qO&i3
�,��"��3:�h�E�'E }3�,G�G���@��4f ��a!�8f�!�(��@k��&�N�/��[R���&ɴ=D{�G�H����rk�)��"UfI3��Ĩ�+>���C��H#nRnD��N��y�*��}����E�n����'���MÂO�t�P�P-��Q��[�#U?�h�k��Vg�`�d8���Pt	��\�!�$_���8F�)R��q`��:z���9�Yc��%%���ۗܟrGy���,±̀&����/�0>yDؑ�rŲp.��"�MA�"��U�>������D./�q)E�V�:���8��D�#��F�a�ؼW��O|��Jկ?y�u�$g�~�6�aR ��{���ʐ1%<X{����U|4��G"�x!�X:Z��aK�L�'@"�#D�ӝtT����	�4!�UZDG��E�&�'�X;�����v���1���^Fȹa@Z�TC䉘� �A'  VZ ��U��k�0��u"- u���^��Y�6���qW�	�ٺ��b�A;L�4��u�ة	����DP�q�@4c���:�I9�,�,c��M` G�r���R�)L�|�Zfitt��d8.e�|�� i����`ҹ"mqO��*P	\2 �MQc��7>t�%,-����B~��s�#�@Lz5��:F��Ї�L̜�2�R�儑fJ�1����'b�flq��H�r2�ϰ"����2��O����;sTڕ�v(��o��EJ�ć; �E��#vJ|1��܃0�Jvk @�p[���#������"c��<x��3#tBd	r�=�S�? N��U��'Z��=С�t�����'|���!]�A1���-d�h���B�.杲��#��8!/�9l'B����^i8�d�P+?8�^�b�j��.��xI�%��KM��"T]���F�ՁSr]��d�*��t
��Fa�#�%��v.8���k���yr��8b8&Qb`�Z�}:y M��E�ʠCV�S� ��AA�҅��[4�x�' ��NʢWwJIIA �R%�,p��ʹ4t!��C��1��֧+$,��e��&�f����1N�~Q���:Z�ftJ ���B��Gz�/^x0�e�=7����F!�p=DO�.dx�u@�d��@LqA#ǵ`�M�rMB�*h��P2~D#��\Tx���'�_�s�: �Ь�C����V�1���0���AD&_|f�I�@B�4v
M˟��2V�Q.�(�`�ǱD\�
�"O̭+�
�:�A���M�V&|�6��; ��Ⱥ��X[��yE"�hA�>�ɢg&a��C�KtD�����ۼC�I'�l�QD =+�li#�Ƞ	F��	�D��O��S=����
/o�rA�/��xƌ(��0��|�$T�
I�L���-5��c�B�2���*���6FI��a���4]�th�Ab��3N����H3V)�4oܜG@����'_����`��`2 �*{ ��h�m��
���!��xA�k�o���Ȓ�Q�l'$�ȓ']�u��kV,��x��-y�\��ȓZ2��{t�/�l��hɮ1�ȇ�?��0d9��3�Ǩ>�$��ȓNv�q�!�ݡ:h�A�񫒳%�J��ĸa��(��:=�QBQ��*�)��B�HX��
�zɮ1ڴ- �8�$�ȓl;�x�� #Z��ˏ3*B�ȓ>߂t���χmEVU�NB.s$܄ȓ�`�{�S�eZ��(�'}�I��۬�G�&Z���煘m�p}��9L,��O���� �T�ZX$���@;(�r��$@�X���:+Ҩ��wY�l@��՗z�2\�E�M�`z8L��$k�		�*.CD	�S���<Ԇ�G��S7FA(as<t�5(K%`%N$�ȓ �@�zcD�G2FA`A�P!m?.��ȓ�^銃��h�{����>���"�^���LL�NZ�E�$�ݒ5( ؄�m�@ c$��5�2��E��pp��?H1`F�6<���I�!́GN܅��ΠP��է-l��F��{E
e�ȓ*S�P"��8_�)�tCǻk�͇��ְ���)��4�Eh�)f�t�ȓJ�6�V��4�RA��(a�<Q�ȓq��ᙐ�V,u�@պK�&f���ȓ@�x��G�|�qS�'~i�̇ȓZ�:��fDǂ%�t���鑶t?��ȓ@J*��d((8��WL�7_�R��p�zt��	Z�"(�e��/{G�,�ȓ4`�B�A �@�wiك8�T�ȓ7�x�zӬ2�@�K��I?Z� !��o~v��nܷy��}���/.�r��ȓE8��Ҥ,�\6p��{"��ȓsݔ���5�r� �x��ȓt╉ؠB���%j���<)�ȓ �v�C�C[��@d��)�Ni��(�!���HNȘ�I�0��`��e`�Q�o�,tr�X�`½b	�͆�(��(�j¡�0d���7�����(��j��u,�xF��	ò��Y9�L(�J�2gހ�pb�*�����
Y�ӵ�]��,IhR.L�71z�ȓp!T���W�yHA�H�1�����k�ҹ�tИpx~�0Ҋ#w����S�? �u�ud�^�Pq���F����E"O���I9i�(t�P��H�ؤ*�"OP�٥`�%b�*A׭� ?���b*O!#f�*v�2E�V����'"(�83Eƨ*{P�$$�9�`�i�'hl�˒�3�ڱJ$�ֵ	��R�'��=S�C[=,���!L���{
�'{�[A�D�Ś���}�X���'®��Cݬ�NT9���N4��'�Z0���[�f��<JVB��(�"с�'J�9�mP-�H ��3\b����'��i[�ȬzҀ�CW��9A�����'�tU�pdT����{�D�QM����'��Ps7lQ�5�9���Hq����'}��e��,4�E)�h4G�j�:
�'�$���m�H�qq	�%9�^D
�'�x��u��59$�� ��.߰$��'��=���0������p�1@	�'@����1�`�f�!Gn��'90��4ǂ��~�Q6kK�A��2�'��v��!Ό��`�ތTR�'�r) 9#c`�8R Z9`-��'M���B�`���J���ҡ��'xօC&lы8�2Qu����v!��'
^d21���:�V��v����'�^ț1��7RC4h G�a��0��'ה���A$x��Q*�$�;dP��'��Q��� ?��)��n�2w�^A�<��Y�Q���1GΎ�[@�Aª�|�<ǥԚ.*n�i�T;y��(�%�A�<9�$�A�<�P�܏?֐ЗG�<�X+M+��� 	�.9`mh�I�y�<��͉�z �q���]�w����H|�<if�[������W� �����}�<���.U��(�&��;��C���}�<�S"�K�D��Z�56|�B�Cf�<����ZT�X3����1�e�UO�<A�"?Ox�0��){ɹ4BGs�<��@�8@�´Ȇ+��m�f	P�i�d�<��@�'>�x��D*l~Q��.[[�<�g�����Qר :=�J�!(NX�<�⮘�ݜ�[���0y����n�T�<�SO�G�a:dG20�B� ��h�<df�á)�(Q��@���]�<��]� ��KK�&=+��S�<�E�W *f��˳�H�9����a�QL�<a��Ęt���{Fǔ�b��9�'PJ�<Q�F��h��Ñx	�H:q��c�<�Ac��d1,����J�mc�$rGB�c�<�1O� L�� OW 2�u��X�<�P�J,Yz�"G� a�B0K�ʆW�<6	�EKxi ���[r�!�N�<i�.U1 �̀Z�F��)g��2�L�H�<�ČX��8�S偁�}!*��nb�<���I�
�J�h��ݦ{)�Yҧ\�<Y��Z�����"hT5Y�*�[�<�BV(��Ȁ ^4Wz��`4�X�<���B�Ohj�����;�����W�<!�_4Djb���F
?R�E5��k�<��@\Z$�\�Ҝ⠝)���]�<�DM_�y��h 7�ӑmʶ�����Y�<ia!8�*��s�O�P�P��l�T�<���ël��á� -S$H�a�n�<� � �d���F�X8���"�n�<� �-�v)#
H!��ǭF�n�"O��i�)�K��TGF��2���s"O��Q��F������-D���#�"O�K�J�^���bR�I3(�@��"Oh�Ѳ	��(@<̨��L��Z�"O���Q�X�����#��&HSܩ��"OJ����P>q�	�s��wV&��"O������"�|8sp�P6���@g"O4U�䔍T}�m��X[���"OD��I�$AR՛aĐ�lKm	�"O����28���$LY�"OA��ʃ�Y���@c%a�3"O��: ����uj"e�&FI&��"O.�#f�:
�3�ՒN��l�c"O(SoI�1*�Љ�؁2�N�@"O�㧈ڑ%bu�4��Q�I5�'V��b�ټB�t�9�͘�h,�� jW�W�B���i���'���۱=�>m9s���!E��HIt~�Z���3v�l'�����Qy짺��w_�h9��G3q�>�	 �ԙ.���p�Oy�`�)3\<-���v�xi�U���=\�����0b<t���t�s+D�zӧ�gy�)��xU ���Z=4���1I���?�G%��A|��Kӛx����5��4�T�ٵh1tD9C�9�X�Rc�	#IĚY�N��x��1O�,A���Q�8cP�ˢ�Z#F�4c�,�ƨ�d��|�'͘�"�oú#m�\��c�X��O<��������OW i�!$5��C�^.�<�vEA�?�A�I����4��S�go���I\�U�h��dD�B(����(q���'�RL�ᓤ.T<aF�5�x�y���M�R�Ñ`��#�|6��|r��AwP��$f�="�N��C��}gxeɦ��W$��9}�����,��!#$j��3UXse)�pذ�'X�Ixb���k�.��.[a#���)�*K��XZ�M��D}N���!x� ��d�%5ٶ}I��*[��nz>��g}J?}�拊7=]���R��9�N9�󉒇h��|�'�b�mڳ=�*��ɏ-du�=� 32�<
 �����?q`��#&�Oͱ��LR���DPA�+�BV��C���CT��>�|܉4C�0�4�AV�z�h�`�@�D�(�f��?i��&&�4 !$B
�Nاľ>9��AI��H��$f��G4x�s'���e8rm�оi��+���ӰS���c,ϢL�кC���F\	3��d��Gx��~�ڕ�`Yg�0s�`����}��O<��1�)�$	Ϸ/��'�X�Z�HH��y/�L���!�K�U[�a�^$�yb$�3h�^-���γE%5#��9�yRl�<3��E��@3���0E��(�y�ȓ)���CQ�H��4�Ф� �yb���(������K��f�jTb��y")�mz9�Vi�}H�@S��y���s���ҏ[
+�R��cI�y"��[��B��I�$�E����,�yrE$ja��H��H0F ��y��V8h=���Ɩ:����M��w:�4љZ�P�`m�?Z;2���F�x��e�#9�@��Å:�Q�ȓAm`P����R�lA���(�}��X��MQ��#k��]�s�_�W����r�8��
�"M ]�U�C�`ޤ��{��K�˺z\`��J������{14��Нs���9��� ,@؅ȓD�	/�M�)���"#o&�ȓ7�Q�b��m�a���
��i�ȓz��]���^���P��㜛E�لȓ���B�+�F� �ł�i�<Q�ȓ-�[4ehD*GKR8�Y�ȓ5�X SG_9W���!fʌ�KIt���f>ʽ�$�@������'9�@��ZBP� .W�a"�38Sre��S�? ��dh3~�P���()�1�&"O�T 3�8p�:P#/͗:�А��"O@�B��(<�a�6N��B��`(�"O�1�nN�.N��3��J�����"O�݈a�21
6��i�3}�$��"O��P��bBP6��2&�,T��"O ���N7s�hlB`ǥP����"O8#u�ޅp�T�-� @v(E�"O��a K!^d`���"+_����"O����HG)��=��a�wr���w"O�0IҢ[ 	J��NpZ��+"O����8#�ఠ�3-b��*3"O�T���Z4\L���Ň�dM���e"O6����`��K۱zYJ�h!"O�ɚע�:j/bлQk�A>�ř�"O(���)g��$�H�6"�1(�"O\(i�(�,z�б3�l	���"O�̃�l�
m����@�t�-��"OĠ2щ�7L���1�ؐ5�ts"O��Җ)�>��Eb�`�
��!{�"Oruj�N��H�z$�@�\򢍩D"O�52O����/ӣ�$�4"OFq�0'�3
��m���	���'"O��ܩA�|�*�M�pdTi�"O*�K�dۄ+��р��R��A�"O�Pxem�5u�N�"���8QےP��"O��ϰ��h���
Y����W"O.Kg��1�"܂
�`����$"Ox����@7s͒yS�h��\- "O^�:u(Md�!Q��*}O~5{�"OzP�a�P�H^$0�m�r��	�b"O�\������V:/�p��$"O
�Y"mH",�,@XS*f�.�I"O�e���ףm�>�[���cq��I�"O��bhO-I��XH�
M�I����"O��1�+Z�FɊM���.C�8��R"O֘��L�u~qadfeʂ�9"O�I��Ǘ�Qx�ͫC'�sV�d��"O��A�CJ�}I���!AY�b�(�p�"Oj8u&�\�Љ���~ƔT�a"O��(Ї-N�&�:c��.���f"O��`���"�T�D�-n
�=C"Oj�#k�1Y[zlB�*^�C��`�"O����eګ����Hـ-W�{'"O�\ 3eV<`��qB��c-���'"O:	���W)AKxxIDO�����4"O^�)�JO�?�H�PtMZ���x��"O�я�	S�^��6N�I�J=)"O�(���u�r-!.��B�j�+U"OrŪ�hřVҘP��ӟ�,�p�"O�U��̫y<H�3�� N�����"O�9�Mދ%e����BWS�vQ�%"O� f��?K8��`dCQ3R���X�"O�8�V� $:L�����?x�^�i3"O�0���iW�A!cM8�R��g"O���D��$�T�L�85� d"O�i�������k⁈�s��h��"Oj�(kN�)��:!�,�L�#d"O@4�S�Q>h`0��tP�"OB	�T��_�@�Pl�5qN ��"O^y�L���0�2�^9o0-��"O���FIm�h��*�"]���"O|,��
!!�� P�^4`}*!"O����&B�H����c
��3�"O� �H�gG�M�H����d�#"OQK���#���f�{��31"O<�2g�յ}�r�Y�Cլ#~� ��"O>ăc�(�(�C�CW.=ӆ�:�"O�ҕ��fD� 1B,��V(-C�"O��!����v�&P��i��8~4y�"O�q���2��	��
ǜB�A"Oj!�u,�=���'�V"On4�U-6=ݸY��Z9th��'�l�5�Q�   P� �ܥO��K�'��5�ė ���C�M��q	�'�dI�Pn�O+�d#g�K�Ir�8
�'i���ϝ��IG�Wc��-�	�'� A�,Qm~��u���Z7A�	�']�A�>J4�YU�X��e��'��!�g�T�hKt|A5o�M��!�'��+ՆN3$�p��٤S4���'}J�
��3Hr숁Ɇ>��ɛ�'TP��l�Gy���@W���h�'�Z j���'i��m���h^Q�ʓb�l����B�p��U�!��?z� �ȓ3?Z���8<��`��B҈!�ȓ,�L՛pJ�XS���لZ���XB\�B�=>�T�a�c	\�ȓ���b�E\�t�ӥZ7�z��9.�p`C�v?d��KPf�ȓl)���U�ڥ=n�����
~�jM�ȓc�dC5KOю���c+]�Y�ȓ�(���+��  ����+5׬5�ȓR��hp nD*K帘� �)4T�ȅȓE�Ū�$��~~�넡Ү\������)���!x��{��B'� a��b7PtZŦٷ�֨�$�A?6<������,�|y�4*Q�Øgq��ȓ iT��P���I�,΋T&�͇ȓ@���PE�0da��LXs ��
I�\c�(�;>ObAWL�3�p��ȓ$���c������%� ��ȓ3o4K�%�?=w^�cɝM����T,X�!J�A��D���Gk��Ʉȓ0FD�+�^(��������U�ȓZє�W�'Bmh�@�Ȅȓ}�ph`��U�
��#P&	�f�x���v��	$�ש;Ez=��j>T��4w�-�A�ߎZ�\���lۇb8@�ȓ��<1�IC�0l4)��	�p�|��ȓ���.$`����8�^L ���~�<��I�42�n/ĸ��߉K>(���'\r��N����s��4E�*��'∡:R�F�g�"� "E�5�n�*�' ��9����1h��/P�	�'�l�;4A�����]�q��|	�'?�D �Fͪ1���!*�j��p��'!Z��T&�
����O�`��,�''��)��ST��+� [N$p��'�T�z�o��N�9��Z7TOd�
�'p��b�):?��BRB9����'�*US�	N�A$4���l�90�zy��'F��CW*]N����.\�a`�'���:�HY�B� Mٱ
�'�����	��O��!5�R�c.,i
�'�,I��oӿhԸaC�
d�8�	�'P��p.ȱ^��m��aɸ.wtH�'TI�3�X��,ł�O�J�2��� b0�Bh�jh�b��A5@H0r"O�!q2 �^��^t ���"O��A��`��9 ��#C[�li�"O� ;1/J5g ��s���0KEr��"O�f��t�jȈ�$��Q&K3�yB��Ɋz��ݎi�b�#pND�"�\B�#)�,�� ���Zm��hÌ�C�I�>x��;#��W6�� ��+R��B�I�ͺP���6u��Qq#J�m�tB�*7��hz�C �2q@�hfB��%�z�s�'�>T�"P�X�2��C�;9ވ�hҡ7���"�6^p�C䉢J�pmcæ]�`���ڂ�3IjXC�>j� ��k���A���	��|C�'Є�h[�1�ĩc���7[|C�	�q�"L8�&�7QJ�q���̢ErC�I)1O,�k���6�4X�U�ɠ$�XC�	

x�0�G=�i��h:sPxC��$U�Ƶ���K�\�}�WTKPPC䉢킅8W��B�] !猿3�&C�	�Da>��� $��q "@]�-�C��,R�M�e�ۗ6BH����F 5�B�I�;�8��p�F��[�B�x��B�	_m��+��_��rHZu���FA�B�	��Zɲ#�X�V��\��	<MzB䉀�(4q�kK9(��[&�G�bB��;9���[���2v�z���M�6A| C䉎o<j� ��\$����'�U�fF�B�I���T˘(��1CD&��B�	�:>i���k��+GgS6R��D�(H5Ƽ�mF(e*1���N�Ts!�ę�u� eQ��:4T�x�g��!�J+8��T*?R�5�g�;!�DE�AG.d�!녫[bN�
R��T!�ШdLv��Ǳ\&@9dO�9Q!�dЍyOdpz���U�1Q�h�2+!�O�>d�<��b�T3<�!*�,r!�;^XZ�pׂ��W$���g��j!�$��E�Pp��X�6����'�tW!�DV�)g� �2!���1k�(1W!��Q9M�ة � ������Z!�$�7��ĐC�[�-��Ez���V!�dS�^�V�3e[�!�*��%��c!�d��r��ś5�	6��%�c�V�-Z!��	�P8��S�쐘^{�@�G+=!��0;� �  ��   �    j    �)  z3  �9  @  �F  M  HS  �Y  �_  f  ]l  �r  y  n  ��  �  a�  ��  �  -�  n�  ��  ��  ��   �  ��  )�  ��  �  ��  ��  &�  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k��'�O�����;-픬�ª�O;v�92"OL�p&�V�Ae�Uk��K20)�"Ol�:��a޸q�JA>W�(I�"O���*�'SCF���� k����"OZɪ���w�f1b#�?��
B"O"�S/���p���{���3"O���S��J��:�oBXY�I��"O�iq�,Ц^\l��Ψ���P�"OT,��˓>{��x!)D
z�^	(�"O��B�=2t��g��?͢-Q�"O�|�� �Cʤ�A$�z�j}�6�	Dx��"g����ب���_�b~N	S��(D��aĮ96`�+#���0� �D'(D���d/�g�ޤiՎ�?>x*C�&D����S)*��C��Hg�a�O:D��t�Z�}�T��l��1PQ*2N9D�X�rدr^��0��R��L�`	"D�L(C���O;>�"\���$��>D���`g7?�Z1#���Ĝ�zp!<D�H  닗W���uiX( \jAXE`4D��cbB�*0L�AALպ"RQ�4D��W�8=�T�+�(��m�����<D�\*sœ qt�w�Z$��!A$'D��y��_7F6��u�׆J����'D�и6藡u[0�r!�W7WԕR��?D�8y�拁&4�A"[3���#�=D�<c%�ǖ-�@�q�E�Y�v�Xb�9D�qc��G��H�ƭY���5D�(ّ-�"�4�+�صWC�}���3D��`1��Z��s�*�!l�M��G2D�Rcb1"��Hu���G�����3D���Ȃ~`�Y�����i��#D�Pp��`ɨGǋ��M��6D�L1s*�9nޭS��G(�l-�Vk/D���'#�#�h��Bj��iq5ԥ-D��c@��.�"\��f��A�=s�L6D�H*aKO�j�Jt"W�ٗB6vm҄6D��{dE�${�u�&#�}�7�1D�H�˚�/��S��S�p"�����$D�t�2�=�\�j��VN�v��E$D����#r��x�+�tAn�Z��#D�t"���g6���g��CX`���#D��J�5��cMw�V����4D��I���-!|hŮ�_�2Pp%�8D��U�F�G;DqI��
4zoH��ԅ4D�H�����2�t�c�I0.�}{��2D���7mF�@��d(��G�k���@r�2D�PpR��U����CX=�\ٱ�.D�La⠕;o����+V䒘J�.?D� k�ev���X�'RP>����>D��e%��@kdـrCE&��b D����I�]2�*֍�<&1ޤY�l<D�{�W�,ّ�L�b�h��A7D�� �0�/G0q1��hv%͒S�`�"O�=B�ᐺfPLd	���|4�"O�4�g�6��I�$��/���#�"OR\8�d�kC.��"H�|Vn�A4"O !R$��(au����I�@�CD�'Hr�'��'C��'|r�'���'F�<Bt��Udē�A�<���'H��' ��'X��'C��'R�'F�陥k�c�Ty�A�� 8�A�'�r�''R�'v��'�B�'*��'�
9(&�J8"Z-X�ˀ(�I��'��'�"�'V��'4��'���'F��f��|>ě�Ԩh���2�'y�'+��'��'
b�'���'w� JW�֕3yM�ŨK�M{���'JB�'���'���'o��'q��'D|���¾g�J�ʦ�k�T0'�'���'���'���'���'a��'��zЫG�Y��8qH
X+]�!�'���'���'Ur�'��'!��'��xc䖺6"|,���W�D�"�R��'���'���'���'���'�"�'��dA棋�@��^}b� ��'!2�'{��',B�'b�'w�'/)h�M��>�Tr�GܨC���
"�'�b�'C��'e�'=��'���'�B��C�q��W��[5�V�?)��?i��?Y��?	��?	��?Y��B�:��P�"A{��m�9�?Q��?���?)���?���z��'c�l��F���o�x)����KI8Ud��?�*O1��I��M�#�/��� `MP�7�*�&�B�g����'�B��<y�	|�K��B�\�@���A�y������?Yp�ń�M��O`�;�jH?�9�瘯gJ�q��[ -�)�r`#�	��,�'��>%�kV�I���J�%�� }����5�M�"��^���Om�w�Xa�@�\/b�֭���F<��ɀt�'t<On�S�'Jy
���4�y"&\���+u"2(<��#!���y�?Op$��<Cў��؟T	�E-fT�*F@�'R8P�V.d���'��'6���1O��3B�@[B�a OJ9��`�@/�IVyb�'�r4O
���-a$��,�;�˰3�Y�';rE��wkdc��te�ܟ`c��'��!���tP8%#'Ąr?f���Y�D�'>��9OD����Q&C�S����8O�mڌb�f��?���O�%a7)\�e��)j�o�I�,���'�r�'�B���f���ϧJ�������j ڴ�[�/�MP5��V��'�H�����'�R�'@R�'ih�CɃ7F2�hibCO=+�z̻�W����4'�]���?������<���!��qa��mͲ�@Տ���QͦEr۴�y��8H� ��T�$��4hu)��|�B=�"/�1Or<�O	L�{�M��?��8�[y���I��f�p؇�Bh�pX`�'���'�����t[��j۴_�4(���8�J�c`K�:�`6��#R^�"�'���<A�i�X6��O�  �7|�����C�f��=�K��u|6����9��3+��@�'��'I�� �17�h�	w��H�<x�ql�9|�b-��?����?����?i���O�<�xU�_�F���f*�Cq�'B�'XJ7M�.d)�I�O ��+�
�r�^h���iܮ�01�F2��%���ٴ
��O<z�a�5�,?��&
��-����1#:�$7#B,4�y��n�O�;J>�(O���O����O�tS���%��(l���\���O���<�@�i4P���'���'�ӭ@V⑈��WqX�w%+\�����O7��t�|��� Pq����ƕ<7��d�JF��4���tkt!��4�	ş�B�|R 
0���I���!�����!#�',R�' ���Y�l�۴3�\���~�ՠ-	*78Ʊ�3m՚�?����?9��Ho��Y�t,#��]��2�*I�T�ݴa��nU�|ԛ֘� 3��]�~��d�~ZP�\���4��8�.��`��<�/O����OV���On���O`ʧR2^�Z�#V�nj��K�;Ec����i���b�]��Ih�'�?ͻ@6쁡�*C�E[���쟹S�@�	��?��x���,��V���<O�t��`��(�4xV'R�F��+"=O�Y��b��?�`�;��<�'�?	�!(
���ō9��@�ևݨ�?���?����dMӦш��F՟����|�ꓤ"2�i{�D�(�6E����v����D�Ot���T�ɱH5��3�)��O6���%c��<��l8WO��A���|�w��O�1�L�<p������J���� ����?!���?���h�6��U'�Z!X� �[��w	ߖrH�D�֦1�c@���������?ͻe7�4s���h��h� �Hh��?��5����8=ޛv���a�o!�䧙&@�����B�Z�f��N�z�l&�������'5R�'��'?�tٔ��[�nxAu�̚D�N��RQ�L#۴[� ���?)��䧋?�s �4<Ȋ	���xzX`gL<�����E:�4rs���O�J�1D�M��7�E�<5hE&��Bؔ��O�y��*O9�?�A� ���<�a*Vv��8�F@�%���������?)���?Q��?ͧ�����Y�L̟8���T��0� �(�%�1�S��ß���O�����O��� ��%Bs���c+�̸3�ҳ8߆�J֢
!]��o{~�+Y�*�Ԉ��Kܧƿ� �����#�z|
��M).�� �q6Ob���O���O��$�O(�?}�V�K�X����hxNI�aן|�Iɟ�ܴ/h<h�*O�D<�$�o�������h��%z#Ĕ6gQ�A$����ɟ�Ӽ#���nJ~"N�#o��S�+�u���:t��P����Qg�|�]��ٟ�I��xk��>03$	�5
P	U�#&����d��{y�rӆ0kRH�O����O��'1�&���c�*��)�$�]qX�'��֟����S���Q+l�$[5F�Ay�1�@{;���A�@zt��O���?!�c"��+FG������>o!.�
��K'Z���D�O4��O���	�<���'��Y�&	�Gk(�c� �(`,�qS�M�5�?q��?9�T����4s��$��l 5Ny`���%=�8M��i�7m *p+l7�e���I�g� ����O�,�5��q ��$���"`��R�y�0�'��'��'2�'�<7�*��`_�Y����0�?RD����B‾�?1��?�O~��?ͻl_�Q �И
��3���[Xx�˦�'�61OX�S�S7m�n��<ٵb�by�Ԁw��f� 8�.\�<a���`���� ����4�X��k`��`���FA(�Ȟ�"?���O~���O�˓\��v��A�R�'�b��v��X�ef�1m2pȣHP3�ODʓt�f.y��l$��J�f�S�"Q����\p�Qk�e(?�2c�"�B� I~�'&���K��?I���%`��Bwj5��	�f����?q��?���?����OX5)��޹8�rha�E��T�UCA�O��nZ�'���	���Iz�Ӽ+���Xy��q��
�Di��@�<���i*7� ¦1�5���E�'T�B���?�XC	/EL8�L�#dnH���D�M��'j�i>��I����ߟ����3�Va��H+Ch��P/+y.ɗ'[
6�x ^��?��Ԉ�$@<���w�1K�8�I5��.J%��������S�'H���Z%̔H듩��]�TrԊ��w����'*�x���Uҟ@{ё|�Y�pbńS�#�"�;VDO�G&�@�@����$��ݟ�Siyr�{ӌ�q���OF �Bʕu���뤌Z"t���4O��*�IiyB�'x�Ba�(�H�i���Yp�9f|HX�`�x7&?�!aC;@*X�I'���	���dARÖ�5l��;���:G^��	������������f����s�E_�C<XQ�An��:�N���?a����雨r!��˟�$����%�-r!ntӗ�?
�2�[7�۫���?���|*#ߏ�M;�OH�Kh�6W�h��Y�\î��'<&��d[�T\��O���|����?i��B���Kc�ܺ4�m�gl�1Zy����?�*O�Xmھ{_�!��ן��	Z�4'�
²q�1�^��6�ʱ��$��d�<Yu�i�6M�v�)
ԎcD, �!��B՜1a1R�(���*ݓ����Df���$!A�|R�P.@�0��U'�&	������\>b�2�'VR�'z��dX��޴��x��+ͺ/��@�3��.RX���η��D�O��ȕ'[£Q2e��I��M[7,`R�H��&���}��9CBh���L�DB���p�O�f��$G��:�2%hKɢv>\��'v�I쟀�	�����柜�IP��j�xQ�	���"V��3#�ϥ��6��"���O���4�9O��4��ҴHK�k�~lpTm�=h�R���
�@mڍ���?��?�����6� L����L���(Z�yq�=���<@�N�O�œO>a,O�	�O��JW�șN$�c ��VD�m��O����OR�d�<�C�iO %���'�2�'��l��$ղ;1�غ���:�p�$5?A���M;f�xRGF @�4��`ßQ l��i�5�y��';6���H���H��Op�	A�?�&��O���&�3y~lKש�:b����"�O��d�O*�$�O��}����l��(٢q�fJ�؍����6ޛ6F�@J�I䟤�?ͻWz
�ȤU0Tz8���� �A͓|(�Icӌ�ldQ�(n��<A��<:P�����"�`��͜%p�F
��i&�`��#
�����4�����O��D�O��d�.J7R8!P���1��BF+**�ʓ9u��gK�2���'%r���'����[�n�}���ǜ/i40�[����4n<�#��)�"H�J J���H��x�D�1k#
��pb �~4��$bbF`��'�hX&�p�'ؒ$8A�@-._�ܱ�hM�H�{��'�b�'����dZ���4f�9���o�N�
��� �r@EZ*a0�%���?1��^�8��ПX��4Q	�K�b�j���#�(/���{B�*�M#�O���������w��b�4|T����݈X�l��'0��'�2�'��'E��9�Hۀx���%��^�b8hdl�O��D�O�]mZ4B���'��|Bc�;`I��iӄg"���o�a2�d�<a��M�'7g�=�ݴ���ǄV�@�K�e8���0̄�Y�^�Ӧl��?�#(�$�<ͧ�?���?�N�C�$�wgSl.x�	���?������ç�Ɵ �	���O���Sk�b�D�l�'{��K�O���?I۴�y���<\�(�s� �R���ct-N|��E�h3^�h����)�RjQ�	��<YE�9W� �FV	|����ß��	Ɵ��)�Vy�Co� ���B\��"7����c'�],��O��?��iy�'���K!aET����G�u��@�'R6�P�\H�6*?ɐ��F���,�� �x�&d��X�"�1�$�$㔱��2O���?����?y��?A���򉅞��)q��&Q5Г�ڹ>&d�l�K�����p�IJ�s���i�-j���$�s)=.�t�@#,�ʟ8��;��Ş7!0TCش�y2�֕+;���@�X���t	�7�y��ڿ��!�	O��'��i>=�	�"(Ш��Br]`ph�H�{=4)��͟��	����'(6�X),1���O����w�x��a;��'P�kw^⟤�'���'��O�0� �,8�8�1j8����0?O��Ą�2�xq0���I�I�?��0�'��I�  >��KÔq�L�R��Ps�Q�I��8����T��b�O�2�"/ҍ�Q"�Xl��j��j�bCw�r�h���<������yW$�6��)��~(��[�⇶�yb�'�r�i��\��	m�B�	쟌p�j����c�;X��[E�
'o��=b�����%�,���D�'�r�'��'%D�8��Z�cs29��G�	k�`�yV��Q�43�F\���?����'�?�u��"`D ��5���ʒ�)��$�O|�$�Z�)�Sn)��k2J�^<r�%�"4*T"԰&���uE�T� �OƩcM>�(O���M2H#�a��,��X��Y2@F�Od�d�Ox���O�	�<պi��5(��'X`��ާd��IȰ
#b�|x��'�B���<Y!�i'x6̀˦�Z1iUp�446�2������X��Ymh~�B�^d�S}�'ݿ+gf��9�ġi�ʗ�9> �/�<���?����?i���?)���l�S�z��c�Ӓ7��*"!\��R�'*«a�TQR���<q����R$eȃ�G4)�L�ya��'y�� ae�|R�'Λ�O��!K&�i��I(&2��VBQ�@��-� V�q  �h/)��T���BAn���i�����b���?�c�	��@b�K�	N��E7�E�TϨ}���?�'��R��M�<����?���i
�OW��a�Ў��B� 3Ė�7���r��MЇ�'���'����?q�I؟@���xP�H3Jm4�P�.`��`@�z���A�4?)��T���-��2_�Ԡ�ᐳE� �����Z�&C�ɵ|�~A9�h��c�A��L�"&M���$J1D��;�-C�b�	�غe�����Ӽ �t�戊(���F�n�P+��I�z����j�-t�xA&�ت$xr	d��2?�~	S�A�Rƌ�;%��5W4�D��;�8EEϱM�ƍӄ��\��P3D�L���Q�zh˟2J�QH��VZ7m�;�����-#��ѱWǐ�,$!�0X#H#k�bE�$&t9��y���%3�$���V�IhT�)w
/��5�r��h��BQaN�Ax,����B���+�c#�5��A�΅�! �+�Q��N���A�hR$n����lj0�ҷ��
i�\ai��pT!�E'g7�o���a�`�EQI|DedC�LԀRϒڢ�x$#ȼJ���q�D�/t��Y��ߘd�.�h&C��?���?ɶ	o�
s'�z��T�O��.���ן� �gȋI>�]��"�]ر��ɪ4PŅE�YvHًT�\9���'�X|�U�&)��]v8q��~�r�yb�ɝ%v��$%ڧH�f�+��[{ܜD���&pI�݇�S��tbr��$a+hM�J=�]��I/��_}DɁ`�"q��s�.K�"�f�<y
�	$~��P�;�����E̛H�ȓ3�x��'��T�];f�.�@e��6hQXU��'*7z��5�y��ȓ=��e� �-t�$�"OKP&��ȓG�.�
@��6��Q�}�DP��IM�	���N�8���C:�`�ȓG/�mXE��| ueK�G����ȓO��4�[
,�2xu��3~(�u��-d����({4��D�M6!�ч�;j]���0�"����Q����ȓuoV��E��3p����Bo�7���ȓ:��)SrF�/0���2��.Q����eR����T��Ub��.!�	��:�	�<�t�S�J+�P�ȓ"�T��"��?
~}B��x�^%��G�1��O�Yx�"���#lv��ȓ���J3L�l��q�:E@rه���8�(ȉ�� �gy�����"鑳�/_ނ%	���f�A���-pq�5��� W�>� A�ȓ9�D��&)x��;��AWkP��ȓ[�V`q�@�!���#��ӊ$�8��[�t� �+B�i�S�R�KTчȓ��l���T��J�00뺵��#��!ʦ��;�nY"GKa����p:DLp���4Q�t(�A)L����S�? pT�'�U�g��L{r+C����"O
H�3Ɲ�b���Ã
�6� �A"O�|z��D1�0�3�4��0`�"O<�R╞YR��3ҋ�"��m�Q"O�ၐ@��Dd툧
rp�A�"O�a�6�ʫdrX9�E�[
!d<HKG"O~i���գش��W:MG8!�"O�������H�H�*N���"O��l�6W�<��2#�2/��Bd"OZ��ሟ,np�H�(�]�a�"O̔C��[�*���΂�Z2�Q�"O�@E�4W�������:'VjY`"O�љ�DW.C\�Q���hL�#�"OV�!B#̰r�*�� ݭ`b}��"O4�@F��!G�"����\�6��"Ozg�N6��Pzg�?+ʵ9"OS�h6�6ظsA�%�q�"O���C.�6ŰPy�M>i��Q��"O��uH�\���I��:�
�t"O����Ȍ�}L���PÉ�N2�8�"O�ʄ&��q*\����5n��s"O����,X�n�f�RA�#�9'"O�!��-	g�Ȫ�j�5Y���P3"Oz)4!�`}.l�E
�,|m�"O8�Ks��C��[�T�p�9�"O�L��Ee@��A��	;l 1�g"O8D��n�Q���r��MDZzqx�"O�yQ��)Q��ʵJ��}@�p)@"Ob�+��h5t�0ѦO<X*�"O.�p�?<�:	�GkS�,=�i�"O���B�d�f�z��]�����"O2�CW�|t���jj�<���"OTй�K�42r�H�Y��P�"O�t�eM�r���tbȐA�hx�"OL�I�'��aP��4�Y	F.(!@"O �W�?J����;S����"ON����>~�6�T*�:�R�"O|�ӕ���:�!6�A
r�PA"O�1C�'�Y�Æ�l���Pt"OLq����;E�xp"��#���C"O�;�J���(���חƽIp"O�<i��4� �hW'Qt���v"O )ޏQ�h�!�V�0�i��"O6ԡ'�	�a�Ѝ����� X<8�`"O��sЊC�bL�#� lJ�L��"O.�:�O�X%�`&$� 2D "O����H�+�jѻ�Ś68X�@�"Oؕ���K�����8MJ�0�$"O�i��MA'5	X�H��Y�FԊ1Qp"Ob��0h�(g|�S���d�qz�"Ot��5�����A�M�O�PU"O̵q�7a8�@�a��.�l컆"Ob�r�i�V` "�&\hiBv"O����5n�`�ϔ7%�*�iw"Op4´�F�r����M�h�vyc�"O�E��G0 cԢ�ŕp�٘E"O�����W�xD�Ts�+VC�@<�a"O��G�+P�X@̎�@���)G"O�@��AB�fz��#&��sw"OqP6ˊ&Z`Q�DАX�X�F"O��ɕ/g�\,����Mp�}��"O�\:�/��9[N�!�7U\�\�v"O(��qKJ#P2��M�d& T�"O$Ũd"J1]՘pI�,ˇ\����G"O� ~m�hѨ1V��G�Q;[�X�q�"O��V�A�(:���1��H%f芔"O~��u��]�č�g��-�$ip"O	3�c��Jq �Hf��I�b��C"O�� ��!I��D�c��	C��x�p"O���lX�qz����J�"�x<�"O���Wʌ>+��-2��[H��1"O�A V��A�f���[� �l6"O��"��3x�Ԙ��FW�"o2���"O~IGAY����7�� �p�F"O�YK��M�N�2|c �	�^jRHjc"O��0f�T�^�~(��@�v;��""O�U2��!m�����m�0*f��"O,�2��9�|%���ژ���"O�	H&j�+}+�),�t��3"OBH�B;$�@��?o��$"O0�� �G�X�(��ή*%"O��g!v�N�
��!�"OE�3D\��PMdmS� ��
O!���.2"��T�%g�.2�!8nM!��,��
�=��P����1�!�
�j3����C\�hH����)1&!�Dѓ�C�+[>\x���/;!�dB�2Ɯ�2�=u���c�V�	&!�$��ʈrQeT ����+��K�!��14�FyCࡂ:9(Xj�5�!��^�0p�����3��ڹg�!�$�p��IW�ȇ- ��rD�A�M�!��
,�R%�q�K<l(���D���w�!��e���k�(�*�Э�5�E�<�!򄕵L� MX�ɲ��<Z��V>V�!�DšE;��j%@�6�� [��R+j!� Jq]��K��*�xS�蚔*g!򤍛ޚໂ�L�9Zs�P�,}!�d�Nj�w�@�x �����
�Oc!�d�+f>$w���vIPY��"�M!�d��rH:��Sϙh��X���ϰC>!�$	2�N(���M�Yi$Y����m<ў�JF�ӷǀ��#,Ľ4#Ψf�SnB�	/2�L?{��M�i�%(&��$S :���"~���c��9�G�A��)R�k ��y�f���tX�oDT��$:P)����Ӫ>������0}XX�vI$O��p@F̶k���Dܖ]���I_Jq�6Aѱu�����LxrB䉡C#����lT�"��5�
Z�=ie�ȸֈ�>$�7!�	u&�$�Nު<JV��#"O<�@W0o����:16�ܚ�'�t�p@(�)�M@�CA��T(�w*����'��pB���*4��@Ax_�X��OpD�P�Yg�a{��19�A�W����-�7�Ս��>Y�gT�{����N�H��<B@�ǐA.Z����ϒU�!�$�&��BÇQ9�eQ�ߐKF��\0�l�������!�0}v��4k]�9GdM:d"O�u
�$�N���1�ă6A.�`��i�����/�)��9ǋЍe ��Sæ����C�'D� (Vǔ�S�*���l�B�"����>�R�ħ�p>�b\�VcB��F�G�<1X@�a
�pX�����2�y҅  w�@���l���8�#�yRBS�o�­ìȐ\�"�X6f֭�HO�rZ�|D��C�3hrY;�AL�h*Ĕ����y�k	�U��*e�e�*��J��M����>�O?7	:>j8�Y��1�
UȣI�r8!�$�}��M#Ԧ��9�:8�cKI�3�I-��|2��o��KcA�M�L0���W��y
� <��cٚ)L�	7	��H &}��"O�g��	Zz�8jQ�n�h�"O8DK�.<��(�-\���IJz�<��gZ8q;|صD��dڒ�x �Q�<��J�2��0����OVv��T@�H�<)�L�J\��ҢT3h�@�%n A�<I$hYp�x�%�PWv��Ю}�<�iF��j��+�"J3)9��Iy�<iw��_�� &�$�I��Wt�<��4"�^Y5O���`[ �
p�<�`��1�Ό�a��n-SU�Zo�<�k�_��1oT~�
4� �j�<����qdx�)�&_�(�a2p��h�<�"?��Հw�]I��Ċ]�<�O�j?��X�풭CD��q�X�<�l^t�l����/|5x���j�<y6H�%Vϐ��e�(!ZB��3g�<�f� i���xq�G�Mzt��
B`�<��5Jr�D��B�v���!�G�<�Xfa f�'��ivfD�<�	�o�6Pk�+V3Jq�9t�Bj�<ɄL��V՚��P�{\*E��)Th�<Ѧ6T��E���ͅ<�Qr��l�<�e� �|��4�� (Y�IRɆ^�<�b"��	�v���F<�`�`4W�<��	;1\�t���8^��t0Ӣ�V�<�3�YG����&�6-���II�<iDK�hn��E�ƍ4j�*�$�M�<aM�!�����JZ�d܆��3NI�<"�G��<v� O=
P3�H�<9��_23[4�ѱOtxD�G�TV�<���v��H��;h��sČCS�<�b("J�p5H6Ċ�}�]sT�<��)I�K&2 X��P�eU��#� T�<! ,E<&��)���)p?#��]P�<�A*�,>����H��`9F�N�<)���-��iy!b��B�0����n�<�&�l�� 3bȠ ����G�Fg�<!Dl	3~t`(0��h�:u��Od�<q�S�vw��⠉��5�Bȕx�<���'�P��w��	(�Ae.{�<)@N�,NW:l��(���`9��Ds�<���G�$��\%���J-�m�6K[X�<AP�ޥ=֠��.�wE�`!�_�<B�D�r��`��		��pvF\�<AgC�c+����-b0���dK}�<�C��Z�(I�GގXƒA�1�S�<�#e�
�ه�ۊ3~CC�s�<9�(�)�� �K
}��5��r�<Qϝ}�D	!'�V/*"�d�z�<I�m]2�؝���Ǎw��Q��Ot�<��lD)Y�H�s1��0!d�Y�$o�<!���8)��[s�� ^�L؆�m�<�F��"���pF��� �l�<���O,M�` '��C�����@�<&�'RW�!ЬYh�aH�n�z�<�S�	�x�A�ͱ?�dL�F�A�<�7hɢk�����,:{�L+@�Gy�<�p����-b��B(t�[�R\�<���(/��I���$w�x2'nKN�<9�ӷrG��K�"�+l��9
�'��၁IS��*����ڔ?^����'��|�$ᖤ~:��q��=c����'�@*�H�;q��hJ��05�Ő��� f @2X/JYL	���:NV���"O� S�ծ9Y
aq��-K^^\� "O��f��b�8U�K�c� 4��"O�A5F'</pP(��g�Hѳu"O��� ��
R�A!U�Y�lpjg"OBx[C���JIz@1A��B4"OJ@3�>y^��⏆�ؾ��U"O.0��e\YZq�	X*���"O�"�m�df<�P��W���r�"OB�R���]Hlm�
W	M6M�5"O���)��uؒm�HV�gC�(�D"OJ�c��\<Pْ������B��*#"O�����Sm�x�g%� :x��"O�I�E�X=�R��7Dܥ��"O�yW���_�.���%z�P�K�"O�����/"����d�h "�"O=�cj��x�&�H���#m�ق"O�=�2�)h��X�DBE�|P���a"OF؈��T�؂�����,}`B|�f"O2� �C�,P��y�!�
N�53�"O���3ߖ!`��&M��5:"Onqⶍ�(3��,{Rˏ� (ɠ"O~qR>-`�x1ݟC;p)�"O.x�%��;�D�5*�%1r	�g"O�3��Z�'[Xt9�iҨG�(`9�"O^����UH`v@[�H�gZ����"O�PÒ�&@��	r�,E��b'"O�4(T0J�R1;CoX�r�8�"Od�@�#�(Ժ��c�SÚ��"O0|���2a�t��QT#�<���"O:���^R�4oC=_I�q��"O��qHTQC��#�ԐD"Oޥ��ş1�h0B��݄a}8<�q"O�0#�� j�d�F���UPv"O��aa 9����`r2!s�"O`�����|$� ���J#L��h�"OXuBu)� .t�q����8� �"O�4�b� ���JӬ��<���0�"OJ���lƻ>���0�ʻ[ؔ(�D"O�]�e=n�n�"��Ù�Ɖ��"O��Y�MJ�hh����Y�)��2d"OFu/ٚH�L�q��D,w�yX$"O�x���f�|�!d��2���"Or�8ƉjW���f��l��p��"O��Xrfɜƪ �ȯΘ���"OD���&[� �氻6��;`��A�'"O�� �iض��Ss�\A����"O����/��0���.�:���"OZMb1�)~B>II�+�����T"O�e�C�EY�0�`�6>�Μag"Ob�۱ƛ�;�8�VkI�I~"	[F"O�]`��H.Y��U�gպ[b�U�`"Oj�"�I
j�X��E]@�`i�"Or�q#G�c`���s$Ͱt5�L�S"OPp#1��j��E��iNa7�t��"O8Lڃ�h�H�P0��n$B���"Ohg$ܧ����`�@:?��5a�"OVܩ$P("�t����jJ��"O�����@�B8�`B$��4B "O�Rc�UH�fJ��c�X3�"O���Uf�".�9(C/�5HS"OȰ�O�N�~pBZ��(ݩ7"O�t���1. >��C+��'ͬx�"O�y{C/�i;�3���9;��A"O� �ȡv� \/�œS��jD�;�"Ol(�k�f�{���&;��Q��"O�d[�b��s�\��!-&p�*QI�"O<�x�#�8�\�ENV�|�����"O�A���L���X׬+F�H��"OZ�д|oΕ22�N�:�8�3"O�Px�J�0xr��0%�n�r"O�X@��%:��%s����K֭�yR�λF�X�	��V�6����N�y`̱z�Jł�%Q\Qԩ �X��y�O+��a�s��* 
F��1�,D��KGd��k��`FSw�p�:0G'T�0`a��/è���)�i N��"O@�bp��(B��"��2@	Ze"Oȥ�u:C����� G".Ļ�"ODU�E�I�&q*� �╇O�XY�"O�x���TF�[⠃�]�X�
�"O��H� Q����F�����'�\X���d��9�eJG&J���'��}�R!Uey����ε�	�'�|DY���T����"���^´���'þ�	Q�X�V%��Q׎��u�H��'��x8��D.�֍I�KSY0��'�>���ǐ�����U�~�|H�'u$=s�AϹR�"�ئ���A
8���'0V0Ä�K�Dgz8�q�%���'���2�kȃ(:��d��%=T 	�'��u�
G
w�����QI@0B�'88{p�ٝT-����2,W��q�'�t"�a��Q�<Q%Ǉ�(N<4��'��L�C-�&��2%/ޜ
�" ��'bxӗ�2ބ(�D(���:	�'���[Ç'r-Ơh�f΃|�w�y��O;D��r6k�42�� �dҊ�yb$H	c\����&����f ��yB%1��� B�"�b��v�=�yk�/o�]�7���Q�#J��yg�u����rD[�!�0��B"��y��	�F��_�f�&i��8�y���0^3�H$t��=Z҆_�y��������f�:�@��ya�$vL�;��Ip%Q��L�y�J`2��j��L�=��i{c�K��y��Y�l5"� �NK�#Jb� ��y�մ"��!	C�\9LN\�D��y"/ӊ9�$0��؈N y��,�y�H=;��:VE	1��ٙgn��y2�%�RԨ�N�� �t��_��yB�?�,���z`��ec���y"�8*�\8�liD
�iD��y�@N0����/~`y�0��,�?����C�T��冲$㺌p0�E?X�ȓp�theA.:���A�- �cs����x�V�9cK��g�`���)M�9�*���2� l���ө1��@�g�|�
C創~�pH#�CNHd�c#�@�B�I�	��K��?k�`��] x�C�
10Rh���E.?t��x��.O�C�0hu�E�WG�l�����Nu�C�		1�M�1�m�a� e�':DrC��#hb�(��o}� 0eL1b��C䉚\]>9�%�(_�N�����Xl�C�I #��h�c�׳<������B-)O�B�ɬ0O�����r�������,+a�B�)� *|BMS�Sd}�s䔯���;�"O�`�T����z�yщ���2�"OCu�V�(���&�L�O��"O��v#�kF�:GT	vhf�i�"O�|⣦�5>��b�썝2�
�SW"O9	q/��.�"�Z�+�4P�H�P"O����G5l�<ٻ�����$l�a"O0�A�
Q�l�,q⒄ڎl�rܣ�"O �.C�d)����j�4�"O�е�Z,��٠�(��$�1"O( ��up��7NGc����"O�$���>����ȪQJ�8�"O�9b	M��8�1��@�C����"O� R!�(ʊd�#˦M��1�"O�az�LO'�)��C�f��iA�"Ov�hW��n��lH#a�|��"O�SӤ�94��f�ȨY}p�Xq"O��ӣk�PȈ��T�S� �V"Oġ��Y�n��� �L�K\�p�"O�m��cP�q�h�1�ɡk_�u �"O��a�U��s��B���3�"O�Ё�݃h�ޠA�"÷k�����"O�@ �,Y�E�Z�<�([�"O� 4�M[��|@ �Ⱦw�D��"O�LA.Ð���W-E6d،��"O�xSŎ	
�ڑ2gM_���x�"O�p� [�b�pa�6/�����"O]��`@4f�q.O=�t1�"Oڠ��m�O�\ ��;
o�k"Oj)P.0tD���C�8m��:�"OԈԤīN��Q�q���{U�pP"Ol�E%7�(�&��6k�����"O�؆�L�x,���J�O©�"ON8�D�.k�Ye�To��Qj@"O
�b쒧bi���`E*���{S"O���P���FX( ���C#:���"O4��M[�g[�m�d�,2d�$��"O�pr֞ڮآ�އ\Z�8	�"OUh%o�6fX)��oY�-B���T"O��s�.A,4>�����>�|8"O:� �j����O���2xJ1"O���*����ݲI��a"O�P��/�?�ni@ڈ2� "�"O�u3��G�Q���"�.�h���#"ONBb.n��4ˠZ�yz�1a"O��zd�MC'���=xL���"OP�l���9�#�ǘ(��`�"O^=��/N6|B�A�6��9G8���"O++�%#U+7�˓@�@���c�<� �ǆ[��M���r5k5lc�<��L�4aP�Z I�)�D�C�z�<�q��@U�0*ab�+bh���H�x�<y�,\❸!CL�<�R��'�u�<�A,�:e�1Y��B&8�p��2�W�<9r�	�4��ub��h �9�S�<�l�.Ge`���f��2�~m���ZU�<Qǯ6sΘ�Zgď�/ (����N�<��!Ѕp ҈r$��8��r�RK�<�g�al��RӢ�	�Jň� �I�<	�)R�wXкA�Q+�bpp��JI�<�6��5
�mq�ܩL�T@4�DF�<A3���*���a%b�.N�h��g�<�֣��t	ʄ�UO��<(����`�<Y�/C�I%�RE@��
D��X�<� ���ЁGg�.4�4�/����2"O���6�H�Nh:�����n�t��G"O���d敂E\����`ڼlݖ�`�"O�ܹ$�'O�����Ϛ�6Q�"OnM�Ќ�XK��ל]Ê$�f"O*�	02F�<0�.�h��ɳu"O�q75~A␁!�Ѝ*|P�t"OH�� �<<�~}p�fڵhQ��P�"OL�#�"N,����˼3d��bP"O����E^�gߤ�@��]�<r@"O \����.m���'	�	�,˔"O�]7	��H����eQ�p��"O}B�D�(�8��Z�"t��w"O�h��x �qE�E�dVԍE"O�I�`����ŝq:>�+�"O�d�����>:���A��$XM~�t"O���4��u�g8I@ɰ�"O�\Ä�N�R�J}z��!EHq�"O
�1�4��d�g��BG�|p�"O�@7.�&J�:lZ��~Z��'"O��+e�F":���ՄF�!�LU[�"O��cٍt���1�9d�@Y��"O:d[Pؖv'���֧�uвY��"Oĕ���>���sUFU9N����"O���w΄�Wd쳗��<v�i"OZ����Z�2�°g9�E1�"O���e��&��Z��� ;�9*O.ȒƧ�e�&����.+҅3�'�ԴaA�_�B�BC/�8ohF�H
�'��"�$Ӥ=I�� q��Di	�'� �G�̊n����OV�5�~��'b��r�T?F�v�!%+U�-�J��'����g�O!Ӟ���)x����'	f���d��"E����Ɠ����'q��R���q���3��Ӣ#+.tZ�'�v1V�ʨW�DQ@�'�N%0�'[�,��D�F;6e���F�(��'M���^��vmBJC���'�p�;�I� ��H�0�+ ���yB�p=��#S�Z�nʺ��K�yb��6�n�(B@ l��hW���yB��K��2�
c�P�kZ�y I ���"ɦZw�(�dȏ�y�_=<����RK�cUc �y"��a���r`�4L��1cR.�y�M�)�h,�`L2E� � �#X�y�@�~��-Ku+((涤Bp��;�yҏ�wF��bed�<I�8�@�y�j��.��@ĢSP^�lQ�c�yң�Ja��h�fM�W~����
�yrj_�!;6�V�W�Nގ	�����y⮛�*���E�)wC~�u ��yr>cm���-L�t�J�9�M��y2�R,�ؽCa	@r�a㣛 �ybM��H������iF�4!�숕�y2��9yb�2B�ɤ,Ӝpz�!�!�y�͎�q�X8ee��"�%�f�"�y��2W��ق�ʝJ�qo��y�ѯ/��c�+�3xt �5@���y2m2"Rj��D�±~7>}" hI;�y2�Ή(���K�{�]{WE��yR���$��A�5��3f�PM�E�+�yb��"/�H�i5�@5Z^|J�H�7�y�D۟-'Čzg�������]/�y
� ЙQ���u��]�c@�t9��Ȃ"O�Q��)X�C�b���׎@�ժ�"O�mH�D
0��qA�%}�А"O�l�$C�?3Ԍ���G� m:�h�"O�͓�g�q6�����'}�P��"O"���0�`�Ǡ<o�|{�"O���)N7��+ �"ac��K�"Or��&!q}n|`��ۺ&Q&��"O
mȑ�S�������	%��I�"Oĩ!4��M�-Y��Ɩ`� ��#"O^�`�79�J�=_����@"O4���E�qҤ	���{�"Y�&"O�9q���ޞ4p�d�3p���"O��Ѓyg�0��e�*G�lZ"O�;���aX��5ʗ�{��X�"O���M�2u���0@Ƽw�e*�"OҴp׀B�W���?j�P�d"O6��!@�E3Qd&ǧS��A��"O���E)
4��P0+�d���D"O=�"��tq^��E�ҩ$�"��"O H�N�D]�����&�� w"OH��5Z11REْ�U�}%r5"O�)3V�4
��*qM�&��qs "O���F�>(h���S֗o�}c�"O�4(BfA	
k�	��d�����P4"O��s��:
��S��0�o=8�!�D+�K�惋v.DI3n��Aj!�߷�%� ˠS<�I���k[!���3�<��g�p��`أ�P�N�!�$��,g^�*W�a�� 
#GԻ>!�s�8�e̯�@�1����(!��\ɶ��'S��&�(!��,j&����P�
ڬ��7�/z�!��R�Z�l���'�6g�ݐ��Pjq!�D
;Y��CR�[
w~�!(6HU!��ڧ#��]a	w�J�`��N�!�D��¸�&��:X�����G!�MKn]���BY��I�G !��&lȌ��- ��B�Ӝ(�!��A�!ӫ�?)T���A0w-�لȓGt^i*�ïj�����琑Z�ن�n�r��dm�%���w隋od���J|��
`. F�ֹʳ��?�ֵ�ȓ)ո�`tC�*ikL)�'�	� \�ȓb�릈Sj��*�"ޝ^��U�ȓ.�61#�L�A�깂pC�>�(�ȓk(\M:t%I+��rf��H���ȓo��C�G�#�X�U�֖̀Նȓz���H�k�,���iݒ>���ȓs�^��U�̍7�Z�0#mմG�	��e�F�p��bzdx8�	�6wpD�ȓ 66��Ra��>���Z�n��!��cr%��Fᗸ!2�x���H�;�!��-oS�mj҂��d�	����.�!���I<hgCe_�J���m�!�n�y�1Β�FX�p��M�!�!�$�&ez�{V兿l�䃧�D!���a����$0}1�*!��+BkB8�B@�E(d��$.� !�d�(C �8g�� ����v��L]!�d� ��|s�M5i����BT~�!��].&7F�B���K������!�dť%��᪂���|�*"��e�!��B�~\�A�_,�ָ{�N-Y�!�� ����3'&s�Ն���ң"O�d����B�f1DMZ�m
љ�"O�9gŅ�X��sk��U�p��"O��˲�95-Pd+` ܥY�^�x�"O���A�E�.W^ �ӮV�%�����"O����24D�CW��m����%"O�H9�G�C+�Z1���?xf��"O�19��/��"S搟cg�9("O69�*�}.$0��´�3�!��kͼ�H��Q\�1��nJ�z�!��"f���u��cn�"�.ɲ^
!��0��hiԫ�jMb]�s���f�!�$L�+�K�?>�sPD��r�!�,>ZX�!u�:~�k6F�)P!�$]-f��OE�w"i2� ܭa�!�D��l�����3,`����F�,?�!�$�k�~��W	�
y��A�E�P��}�$ �+�&(P.�a��H�U�A0�.ړ�0<qFoβ�LLH�\iZ�	��+�W�<�� D�J� ��Sj��dx�Qh��O�<1AD��`�U�ٻ-h��!�GO�<9ArHEC�9g4xp�`�<��N�}��Av#�A���˓)_�<� �#S�RxJ��C^a���U�<�U�֗Z��h���	4�Z#���S�<��g�.L�Z��15l�,��f�<�v�5�V��1z�~ �bi\[�<9��Ԏ[���0TcR0Kt!!��Pp�<1��D�m=�P���ԮK�ɰc�`�<y�`�3q$�Y
��҅і���l�_�<���i�P�D�O�9 , 5�QC�<��.ĺ#�02��P��T�-B�<�CaԕRp|P9�J�pz�V|�<1���>aPb��JP�+��{�<aQĎ���\I�����*��1�Oo�<�W"=?세+�w7����%�a�<�쁖sM�h�3Å�2,���Y�<�b���HI�Y	�*��m=.QRc�Y�<�D�A(hI��ʕE߰#�$-xS�}�<�p�%,t� ����Q�v(HF�}�<�G��9 �yS�Ё47�a���s�<�fŉ�rg���A�Gx
l0� �Y�<ᰄ�H``��
��$��}	�F�W�<��I��ݨ	^�	�zLA!΃U�<ѵ�G�\�>P�%�_�'�ܰ�sBT�<�CĞI�&���gu�t����O�<��̊�t��p�J r�dQ�'@��ȓ���S��,u2p�>;�h)��C\�0��B!`���	f��h�2u��s�r�!��[�U>���o��U�����]� Y�2ID�H3ܩA1j�-	�b��V�z0.Y���zTH��7l�ĢE�2D�pɉ�F�� 셅t��@�N1D�4�����qȀ�§0#t�P�!4D�$�dO�
]�e��>H>���0D��q�F�:=��S�u�Pi.D��W�E0��hԍMQ۶����*D���p��3	▅�B�Q�bh-D�q��h��BC�X�fފ�9��8D���!��i���fK�>�r9��l3��o���@�nN J��%O8�.eB<D�pb5#��F�(}�*25D���3*R#f^�ӧlW9?z�C¯.D�<�sH��Pl)q��տ~Pi�F!'D�� l�����>��D�Uh��a�,,q�"Of�R�딱v�N�q�Eۻߺ�Ã"O* �S�$+���W�nx��"O�0��]63߁/�ܑx"O��pw`#`z��� ��i+�"On�sqC9�`�d�8��!bg"O�h�Ԏ�}ֱ��&A1B�p(��"O�a��6R2T���V�DIC�"OԈ�-\_6�1;�X@3!�'W���B�|�Ps%H7y (9���`�!�$	%;�vha,��;�ɲ���if!�$6|Ԗ�� (9��)����?T\!��U#G�~}�Ū�1E� �*bP\!�$�=\@'	֑R�X|z�b�H.!�+nw`4�`aРI�h ����M!��KY��͖������Hџ,������|Zp�Ҏr�b�
��])]LX��N�<9 �}�8�q�ҤC3�Ec``K�<0K�c�h���Y6&$(#w��b�<q�G�5z�>����d�4D¥N�r�<!��R�+�y��Q�fCu�<���7KAܴ��-�2ao4��w�K�<i�/�$�Eb�̌�N�	��E�<y�&U�|*�eëG�֑���X�<�6i��8΀a0��~� 0"�^�<2F�S�����s��	åe[[�<�� � .�r+c�P��2��S�Tl�<yQ/��n�t)�G�j� �nVh�<��R+rjL��0�D�$��L�<��E�����&]id�
��W~�<y���I�
ģrm݅_�hiBa�ET�<�dJ�f<@�⢇�N�P٩a��T�<1��	w&L)y�B�v�<���^i�<�#�Y U4&�+�F�6�hH���f�<i�#��"�,���jβHXөS^�<
��P4C�m_�wA��dv�<2���G�lLp1��qH���'�s�<D��0�*-��i��kf�s�<�c�7���cf/�ETT��#� i�<�paF�QP �JPN�iD������e�<A��L�$;�`�9A��skTx�<�u�� �Q��	2~V��۴�L`�<���C�wk�1قN\�t{$��F�<���ͣ}:鈷鉑 ��e�6 �Y�<� &��C�n|ʑ�H6�eQ�n�<a�ޟJ�ȶH�8(,��jHi�<��O�]��R�C��j��H���e�<�rG$BB61:G�q�$1�.�]�<1��7)��`@��,F�oh�B�	6hCR]���߃W� ʓ97~B�&\Ƅ�������8d,��&ѦB�	�chV����S�Y�T͘���2504C�	�w����(��IE��(�4B�Ih��i��ͅr��\x� :
��B�	 `!���w�����ϝ�5K�B�ɳ\6H�'��1)���*6�� 4�B䉢I�H�"  ОWp�|�4斔,�B�I�9Q�Y u�	�czhZrJ�uJ�C�I�`�hy�N��Q�\�!d
'Fp�C䉵�(�@��U��QQ�C�ɫ�>X��O�!'���0$��2s\C�ɵjZT��$a�)I���A�G,C�	�J�!���	3<7Hb@�B�N�C�I�zI
��B�(a2|s�eK*X�B�)� X(�b*�@��m�]5T���"O\� �R� 6�A���<!;L��"O�X��2��)�#j�t��"OJD��ċ�3��x4��4�u�"O��:����1#��8/�6`�V*�"Oh�p1�� �ȧ��aĪ �e"O0}Bt�Ipr�� N�p�{"O��[�J�g��;DB��A!p���T�L��J�S�O+FEʦ�*�n�R�#Ѡ�n\k	�'�n�q��S/]~�X`�&
u:T��'�|�Aq�ގ_�	zd%		���'/�2�A�
r����lE�y��k	�'�,!Ya��,�2EX�JZ�t�Vii	�'�5"%�\���V0+��٢���y"�MJ� mˆH#3gj�(wC������O�⟢|R��*
�<maR&@�&�R�2A��f�<�`ۯN|�U"a@/��	+c�a�<QG�
)�09�cK�@���*�T�<i�)Ծ+#^`q�D�&��I��k�<i"<bQ`�� �޻3���f�<�u!V�̓Wd�#xm��8�K�<��Iׄ�p�C��b�A��p�<�4)�$t�t���aP�,`�"���n�<����VX��e�L�4�8d:�f�<I2`��_n@��ΐ�vV<��Eo	|�<�P�֚`|�S�%~́EIy�<�R!O� ��E��̚?mU��{���t�<Qdd�?d܀D����%�<�SQ�Ok�<y�G_�+�hU�-P�G��{�"�L�<9�I��
����(�4#�>�R��r�<7lB0|
 �A�T�zS��r�Z�<�TlO-&��+O��t��X�<�b�Z	�y���0L[$(Mk�<��'�*o�軓�Μf����r�~�<��E�&h����\�|S@3t��z�<1�Ѥd�R��ת�D�n�Hb�t�<�)˫���"v�Nr����l�<�0�B�h �M�ыÞ}�2����C�<����8$g��3��(���Y@�<��I}���j E�pZ����_f�<)�	A� r�Y	a�RF1�D$�f�<�"�A,?o
��C�Rv^Q�Պ`�<�)ə;V�����9��p��_�<9��� ��C�DՆK8��d�<1wGڊ&}05��E��(�(ã�I�<�3&T-/!PH���=k^��@ �F�<��+[3�L;!������L�<)%a�b8 1� �-rT��&�D�<Y��T�[`%`@�z���u�T}�<!�H�(AW^x�ǋ�xAؼS�D�<�&g�i먩[#ٶ.�D��z�<���4Eelٰ!n��<:"��ѣ�m�<�&�Ô2�Vm�g��fW����i�i�<Q��<'b*S�DM�8̺��Gz�<IS)Ч*��IF�Mx�����[�<AT�A�]��5���:=)
v��Y�<yF+߶
pb-(&�YL�-*�(^W�<�$��]���r7u�`�W*I�<���*"ڬ��	����95�n�<�Dڗ
�Ւ��7m��H�V��O�<N�+$$3��Q�SʒIhc��B�<)���
	.� T�9J@ֽ�wH|�<C�^�`�2�C�O����x��vx���'��][��I�_p�H`ŀ�I�F\��� ���9�b1��$�&^�h A"O`�`��C4"V��у�'Y��x�"O�(sr�[��(�Lּ!K�A��"O�u�e�����d�.5���"OPc	�c�-eި_�@5��"O
��Ġ��dP�z��[�ڡ�Q�'"1O�%Q����Qj�sq��M����W"OZ�ths��|s��O����"Ol���wZ���A�${��"O@P�� ��-��C��>iC��b"O��)��֔P.�� �C��%�!���T
Apa��A�I�D��n�!�dC6z���;eL��77�4�'b��F��}���a�셙o��!��n��54x�P�5D�(��R�1�9�Ӡ{�<��-?D����O�)�:��saTv�"�>D�tjsIֆ�j��p.Q
&-^��S�:D���"̭�\�YB���1vH��$.D��*�ҳYɺ��P ǿs�$���8D���E'�$��!1J_<&}���*D�d;P'�2켄�DK�$-�s�)D�tz@A7N�����$�:�g�"D�*�"�z�T��G�#N��8�� ,D�|����8�q�d�Ju��n.D�*��$1����%�eRm���&D���KI87m��'�X�@�Z�/D������G�uӀi�3�l���b D��R F��(ٹc�ˑI�xMy7�=D�4�D^lS�W�� `Tp���9��O~��I�$1He��8r�[��]8I��򄀹4Ă�����|�"!�Ң��yr/[���֣צ>)ބ�B�6�y2H+|_Ș·�*>x�
R��y�F��bdZ!₆Щ$r������yR/Gze<�� �S:Eh3c(��O�#~
G)�_~rAa�
|�~��D�b���0=qb��4�LĆT�XH�7�
G�<i�F����3����e4T�t��@�<�W��z*��ǍZ�daZ�C�}�<)�jEdX�I[�&�R���F�w�<��/�)\P�C���Q�А����W�<��
�S����)qe���I��NP�O�$)���C���0g}�Y�%��	3(��f"OR�P���V�lA�d�8s-���c"O
ݱ��K�7z�<�T�W G���d"O�e#�?�J�b�"� �tIB2"O:���-�O x�:1�W^��CS"O��W�T&�	Q�NW8����'�1O��,Q6�V�\���T#��Iu�O�2d$r7�ᚱ S?K8��
�'`���M�0���xA�,>�~��
�'�Z䁥M!k�`�[T���gJ,�:�'#Ta0��?A�!�ca�4]�`���'u6�R�G��]�>��#�]�\�b��'�� K���2ZJl	���@�^�R���*�'yAz�B���^�^�֡�12vE{��'e�4��E�zfz)���M��Y
�'%L�c4	P:;����È���V�a	�'�$�p��9s���ŭ,���'���#�8�BT`��:,�0z�'V�pa砋�E��}�C�t/j���'�X-��A�y�F�j�"٭[g�ϓ�Ot}�vk� �>5 ��ڋj�`��3"Oj��e�`�$�X�h�)�^�{�|�)�3� ��ڦ���녧Q��"O����N �;�<�фE(���J"OL�r�H�����P⒩6$>��"O�9�F)�-rN�EɆA��Og���g"O�A{�+E��I���TBp(S"O<�&�;�Z�� X'0`m�"O�!��5xj�8��F3Ј�W"O�e��0��	�Ӗ�`	"O&-8�J��m�\R���;j��ؙ�"OH�2�=U8��	�k�D"O��H�厷A�p�B�ܫO�4UA"O�ir'^�Gj^�g��[����}!�ݱ!�t �U\@0�g�7f!��D�.�z�ZB�fHހH�i�>8J!��]����A�W&<G�!�rɟ�L�!�W/c}�}!�$ -r��d�݄K�!�D�L�N�W����ӁЩ�!�$�5`;|0��h�$U��g
	��!���P0m3a��9lٸsn:�!�;p� @�cN�t-~$q�c�_�!�d�	/T� �
�b L���ɡ&!��J<��W(p�����U�&!�䁙`X��K�LɁH�4��R��[�!�䈺/�a+��D��P�b@�y!���lXr4J�A�,Rq�8�F]�h!�d�#�E�����``�a�TE�G`!��Õ\)�P�F��op�љ���E!��!\�Q��kVR��A��45�'vў�>qт`��v���g�2�8���d!D���Y!oo��g����lp��>D�K��*v��cX�p��q')D��5P�C�����Z�H�����"D�d�3��2U�p9�e�XA����!D����e�6gJ�)�5�&{�D��k D��a���� c�T�n���# D�@:�O���0I�N�_�Ԑ�F?D���G�9:��ɓ�@����G�/D�tY5�^*x��!�Ci��v_��B�9D��E�=�
�R��?���[%�8D��K���E��I[����> ��(D��*ʃ[�^���"s�ءK�"&D�Щ�a�.&T�T��S<��h�/)D���s�D�pɊ�q�(�7Tf�qU)D�����2-����#	E�s��(�n'D����L� &N�\����	 �<��0D�y��x?���2%Buq �1
$D�<������虢�
��cE�!�OX�	7|G���#�B5~yb�F@��C�I���	�F�X@Ԁc� J�jB�+/�T��O�t��D��$ܳ#�VB��.<r�ha��ۗGu����/4tC����r�&�������H�T�C�ɶH�|d��Hۻ�D�G[bC�Ɇ,l�i O�}�FLR���X���t��;��2�����s�T�#Ƨ,D�8�iR>[Pi�a�)u�"�u-*D�\q��W�=f��$��Dd�;D�P�Q�4pZ�)_ 5j�+b�;D� �e(�	o�~�Y6� 3amL=���9D�� K��>�t	�/�O.4I�7D��ҵG��wk�}�
X�+r�0Z�6D�$�DN��P8&akWl����A�8��O�����	>;������ih�D�/<!��C�cd�U�G�M�F�V٩Å�+�!�� ���u&V�v�j�UCR05"Of	��`�$q@��ҫ[�X�"O���&៖q���1U���*�!�"OL�1���i�` r�=ur�lj�"O=���(%t�٢���jJ@�Đ|��'LazҊI%?ʆ ���Q3Tؾ$S���y��P��5���E�S�d�S�֎�yrψ�dCH��uK�O�N@�rk�(�yrkS�"�q��#]�R�〬��y2m��*����b�_fI�f��yr"A%3��R��KR��B��
�yr����0���>F�)�\�y�HY}���� �<=��A#���yr��#:���Ѷ(#�IԎ���yB�4Y�8� K��$}BE�$ ��yr$�%@yv8�OH#29�����y"C�����s�L:-�H1�@���y�!�3�eQ��7%�>9�C��yB�O%'�h��sE�3�,j6BW�y�!�F��9Y�藢1���@G$ș�y�➶cD��U #D�`&�2�yr�I9�U��.$�=�$Ι��y2i�y)6�� a͖���1��Y��ybi�/<�v`��d5���2�ʔ�y�hR�)z>ds%�5QP����y"�ʓ�8д�1Y�0
�㕡�yLC�SݰUI��+�X��Bd]��y�/��Y%��C�cv�	[B �6�y��.���
��˦k[�u�A��y��Y�x�<*�EݧU��\�d˙�y��<yb"�)�̷<�l$���-�y2�؞�m��M%i変(!+R��y��U�GUZ ��'g��tX�o��y�ʇp�P���Y#`	0���y2J�<W�D��A5h�Z����y��-g=^�Re��^���#7H��yR,N�G��Qb(� +,�0FA��yRc�
P���O	'v��"�h�y���X�[��]�u�P<Q�n^��yb�1
��Y�v@�V�f��ѥȯ���hOq���2Sa�����r���'$�\�G"O���d�C�en�R6CƇ6n�"OL�C3*кvL����\�l!��`�"O�u)!B�����rwc�x��lq�"O�!I��8/�,��b�]��CF"O�Xveٷ�b��Q���+3"O��T;Ԯ%�T�L�$���s6"O2p���fz	X��\��&"O\e	��A�R@��
�.X�u�$"O,�QW�����7e�дp2"O�A��jؽ7v� 9���e�����"O$�#�^������+��qD"O0���
(9�L���dÔ8���1"O��b�N �B���"���X��"O�@% #�^����ʶV�*s"O�D�U�̧"-����D>4F�-�6"O
x�7GWlP�G]"h�e"O`�s��C�D[�F�-���G"O���❱MW��F�?�d �"O�1����A��EQ%�>1y~Esd"O6�-Ye��W"��[s�ȳ�"O��N������ŢK
���"O�|�tıJ�,))D+�sU,8�t"O
�:s��M2�|�v��-eLj�3�"O� T���6E��>�ti§"O(��צ*��[���-21�Њ5"O�Z��ʐ([t�p���;���Q"O��r�dFW����?�P��"O�,�CR�	QA-�3WNI U"O��ڢ.}����l�&J���S"O��b)8)^�sB�XO>qѱ"O��u��iNJ8Ҥ��+
���"O�u�AE�&��i��U�T����"O�Ԉ�C��t��A�`�"8q�Q�e"ORt�@��5*�@��2"��GL:`�"O��AA�H�Te�1(4�:I0�8�"O�)k5&7��A ���PTb!"O�QP�K2}DTt"v�=rp�"OFE*3��-0�m��f�"S`�@A&"O*�X&k�<�v5 ���-UJ��g"O29�F�O�{Nxt� 7?FyY%"O"u�73P��A��-��	A"O�i��@>lL4-�������"OTe�g�Ơ^TD f撁'�@y�E"O�z�B�#Oވ��Q�\�P�"O(H1	��d���e�*�
���"O*����Q+����,P���;�"O���1$4�9 êV�4
,�+`"OhU3b�Bg=`Q�Wj�	?���B�"Oj8��^Q�T����^��"O"�	@�, A �N=)G�l�"O���҅L�b�p��י=4y��"Op��P�TE�@ڥ�A?Q HMS�"O���!
B�^��X����-洉0"O",!���E�}
��D���r`"O�#7@V�l�f	�E�u�@i����
`�b>ej�CF�/-�]�l'�b�Z�&&D������;
"����A��Y�ظ�)D�VQ�d�mYq'1����D4�yr�Ph�pc�&Ӧ5wXyYF�	4�y#�!?���g�,*\@�����
�y�U�؈�����QX�%�����y�kF2d-0Yi��N���������$�\K�"|��'^�#�����J������u�<�p���(< �#G�E�Z�JSp��t�<�p�ؼA�j����Q
���*r�<ItS����c�솇i;|Y��B�l�<�G�3�l�A �C<��`a��7D�T��Q�)2e"�kW����)D��7.�Ĝ,3Q��V��|h��,D�\걆ך:��釩L�&ބ�1�)D�(�`�Q9z ���Dǋ�\r`�ů*D�,���ʿJ����� ,X|�w�)D��*�+`��u٣B��Z8�w�=D���dG��HY�����(.8��G�:D��c��;4��QIRN<!�p@2�8D��Z��\^�0���<!��A{"�8D�\�O�3��)���v�I�/1D�����͍c#*	wL��%m`�	�G/D�� W�M���qjbF,���h?D��i�aW9\�����F!v��R�H<D����N��A���G���x�R)>D�����HR��0d�(�|��Q�9D���b)�b1~����V�[�3B�<D�4�7,��
Y��x�K��䤀�<D���"/[*�ND:�N�5)� ��8D�`;2�!stIc�V�%Z��P�5D�Й���\��YrvI��Rdh�5D�!�� j���h��y+8ڷ�̱J�*�4"O��ueĵ������]�1����T"O��G�Ѹ �|tA�JO�����"Ox�SW��(y�[� �ehp�YF"O.�b`��	�Z�V�`XZŲ�"O�$#X��ay��_�2;t���"O�Ux��5%�J�Ia��"#%T�@"Opإ��bs�U�D"*�B�"O@���JE���a���s&��[@"OZ0��͐�c��e���z3�9��"O��!Ak��m�2�!�	J-���g"O�����P��8r�βq�$Y�d"O��[��]r�k%a�;�R�Sv"O~K7.(Dʢ����S=�"M)"OF|����7D3v%#�@(d��Y�"O2(�c�( �)�e�+M�`a"O��%o�4X,$c��
�(1�"O���͍ZLR��f,�b�Hx�"OiQU��;M��KT,� |���""O���M�.	rV�rb+�&Sy�m�c"O������.nj���ɞ�_`�tq�"O���chӚuZ9�2"�<n��9��"O���Ei�����[�t\��"O�Ъ�FM:� �h�1x�9p"O�8I�I�����1�.ukB��"OV%(,��\����:eil)�B"O�����=f��xa��MgD��S"O(-��O	V�EbT��Rg�ti�"O\��$K�_�$-�$�#Y4-9$"OBu1�� ��'@�S`��Ѓ"O6]8�ýR{n�a爂�E�u�w"Oj(���#:�����V#Y;��PA"O}pG,ҟ ��a4e�'"�5��"O����ę�:^X�s�ጜ7	RQ�"O�X���I5�d7�J�ޭ§"OVl��#�0��]�4�	���`�"Oj �%o̵.������%L�����"O4���ۖӀu�ql�ty�Ț�"O<�w��-��\�@�ޫ�p ��"O����5~XQw�]�z}�j�"O��[��?�:<��I�3Tڈ�۠"O�$�B�ܯbMD���H�$%���"O�y�t���B��=��W.0	�hX�"O�Q�A��;R*��a�%�j�ya"O<ř�bفQV�;"!8��J"O�ɐbҋ*�Β�I�� �"ObPRK�8%.��TGѪ|&Nm�"Od4��"AliZIaP� l�(�"Oވ��%� * wD�5tUs"Ob<�%�u�>�C�#�,�$CW"O�����}������ٿO�F5�B"OzE�P`NNG���!�ʭ%�*�J7"O�aC��
#��{�ϓ6���'"O\�ʷ*����W�fT�"O��p� ��p����[�ȁH%"O�������� 0��E J�A�"O\�6G�0#8Y��!^>��1�3"O
x) @
<
p��ef@c�0��"O*�1dB	 
�������/E�e��"OB��̖�$�&x��M���	�"OjeD��!x0�4
F���Ҥ"O.A�!�'�4�d�b�(�"O|T	/�.[Rت�6'#T-r�"O�T��ܫ�((%M��\G"O� �Q�&�D	!�ph36�ؕJyle�W"Ol D@L�J�"ܫ�+�#DwF�� "O��QA��4$�pF(��8a�]��"O���E$�(y����yD���"O^�#2ထ]#����EI��6��C"O�L;�+΀=DE�d�jx���Q"OԌ� ��;FzD0#Dx�)cr"O,Y٠��;�VŸU`C�(��b"O��20`@b�x1*��N���C"O�P���s4��#�qh&�0"Oz���L,[�!@Ԭ�(Pa���"O��`KX8]�0��B��"LO	��"O�t8R.Y�� �`����I;x]��"O8���"-c"|�7ƅ!Q?z�(`"O�'�Z<8�21�Yc$"O��u��g�Z��3�W<k�ИI�"O��H��^����1���HPh�"O��	�����7�D�*�y�G"Ov����P;2����aG�+M2="q"O�4�e�Bn8q��K��3މAQ"OD()�G�J���3�+-.�9ZS"O�H����/�fy �	-F�N���"O� iР�u�$�k�KN�Nq�V"O����U�%|�9y�Ǻc�6���"O:Eb���3B�r'ʳ縭��"Oz��(\�mqfE�E���:�"Ox̰���k+���E�vȌ] �"O�X��Ey�H�a%
رS�P���"O>�`�X�<�����)I�.�� ��"O2-�
�;����p��y�"O����Q�4��+�K.~İ�"OjU�N�z(;�i�,j�"O�ق% %Px�L`P�Ŋ#�$��"O�=��"K�kn`�3��V��K"O	䠝�<Z4h�I/����"O�qXr�!
ȥA��
0l��"O:�s��� �,=� �޽XuH]�f"O�`5�^�!NR��U�ZxW�t��"O�`��G3�@"s��kP ��"O�aH�o�+U���A�H[�l]~eiu"O����ǃ�S� ���/!;ƙ0�"O������(\�H!#u�$-��B"O�!4@/i�� x���<d���"O�4s�ƧWyh5Z���7�>H�"Oʅ3�۔L�DY[u�J'hĻR"O�|�h��Du3f���p�r"O��Y ���Y�5��G��P "On��n��B>|��i�v�8lA�"O2e�fL�e]l!�d煈t'�p�"O����%1���f�[�Ҥ��"O&����2)4 B�e܂����"O�X�u��&2>D�cd��vL���"OD�3��Պ�ڭ��b��Q��`XT"OP9rE�Ծ1$|-ȶ��5����"O� @��F�t�H�&�,ytBUأ"OL���b��J�Z�"���C��!�$M�'I
�[!���e�`�s�E��V;!�۸V�&ȫ��;
��P���!򤏿?�8�ڲ�^�"��s���P!�DT�r@��O������g��wf!�dV�8^4�8p�0K�X��g /3�!�D\x�`��MU!Y�G�!�$DC�rD�Dk�#�� ���D�!�ė	j��Pc�a�<�����"A�!�� ]�U��D�r�It�׏N��U"A"O��Ђ��	f��hC��E�>����"O
�R�ޜ6VdS�-�_�~Չt"O���b˂%x�;�,�K��e)�"O^�Y�� h$\A4J�2K{�Q�#"O4$:u��!Q� Y���t[�D�5"ON�9g��:��x�-�(H���"O���ӠM�=���R��ߗVC�kF"O �x������u��甲4'��"O񣔤�c)(�p�� �<��"O������8d�\c`ú~�S�"OJ� $��b-�5�T%rrI+"OV�*b�����!Ꝑu̎�y�"O)���`%�лI	
D���"O(������H�j��@/,���"OtA�@ �6f�n�����pp�"O����ЬF�T�����U�0p"O`��%��[(���a��,�B�("O���ӌJ&j��DYPaj�he��"O*��E�]�Ǹ��bT�d@���w"Op��DFWp4@I3�ÁY�U d"O�IR6ő�c+�0Q�͌,lSZ�@"O��Z��;���F/ �:1�p"O&��􈄰��H�T�j�~�+q"O���v��+$��hC&�	ۈi@4"O:���,��HJ��W":�=˥"O��ڐO�o�49Z����0��"O�l�u�I5aRl�:Ď��F"O,t�E$-Bj��읗  ��2"O^�W�?	��D�V	le#�"Oj=����
(BL���a�� ��؊�"O*@���=�h:#G�%���2�"O�h4lA��ܐS���!>t 8�"O0a�U�N����5��?B �e"O�ez�a�'1�=���\	�� ��"O��1!Om_H��O��ᩅ"O�p����W�rx�Q�߉X����"O�3�
��"���r��Q:܍�C"O�!��P���쩥h�x)$䒇"Or)X�M�HϞ0�FL,u��ɓ�"O�8R`�ڼ���;L���Q{G"O�!��`�*��1#!ۦ�h}J�"O�,"WA�E��"�@�y1�xzS"O�
A�8� �-(�`�p"O�mR�$ŗj�8d��oЮ 7�q"�"O�Ea���a�`͂��SC6�1�"Ol�E�NDU�+��KR"O����A�WB�:uQrY<�j "O�����{.F�	e�� C�ۗ"O��V큁w?6�S"hUq6Vq��"O�� �B]	,�Ԁ�S�A?S�f\1�"O��@�_*�
�� �H'NW�e��"O���	-�.qHͯv@��"Oi8��ш @� FM[�(D��"OL�I0G��7������0h ��"Oj�*�M׍�.%���Va1���q"O���((��}b�V�D�V 9��2D��S&�^Z
	�Ц�m^ ��2c6D�\1FoA5%tZ�k�փc0Hd8r%!D�X�P�C-X��@LP�kt�I#T�>D�9D$�2(����3G�1���!D����$2nŻ�NA�8ۀ�>D�����]梡�D�^�����J/D������xa6f��:��F� D�� ��D�߄_@d��ynP��S"O��d��'"�ĠRl-rO�P�"O����V;yd��`�K�UF��"O���C�PMP�퀱G����d�g�<YVF�3��]+E��THgo~�<aF&V+A�����VQ.�;g �e�<a霛v:�RӆΪI�̌�u��b�<� �-b��Yt�����Ð`�<����.P/)�v̭T΢D��]�<�A)D�GЦh���,/���C']�<i��¾Y�jC+ў5��Uk0c�<Y�F�4��$��͝[u΍e��H�<�w�� *�ޝPpMV z�d�w�FC�<!6�Q�8� ȲQ�B�2Q�T`��<��L!!x�&LSb�JDB|�<iDӴP�d��i�
6�a�"U�<I1b�GK���E�=+��y�<�4�C�PŒp@rN��m��=�w��q�<A �|��|��f
�W��顦p�<�$ǂ~3^�H��!r��'͘w�<	6,F�,�z��GN��5W}�<Y��W�ֲ�A�)L:v���	�@�<�'��8��h9��:(��x��{�<�!�P�zl�!@+J_:eh$��v�<� K�
��	p�����Qek�u�<�@��S�	ʅ����FV�<��Z�Xu+��>&�9ӑ�i�<Y�b�N3f���Eӷnp���\c�<Ѳ��&n���S�K�s�^Q0���]�<�!�ņLzY���b��:E��[�<1��1V>��`�X�JCЧU:~�!�.`f� �;R,��g�N!�ˀbA|��w�1P@����/W!�U
�Y*&�Z;m09�夕�	�!���O����T�pLA0�� q�!�d�G��,�f�υ%�,pNP�j1!��W�*M`"�0 "�l�L�R"!�Ĕ('ఐ�KгO����2!�Dݓ�&)��J���D�L5l!�$Q�����RNF�&;�}���4�!��B5�!Ϫ`�l�l��s�!�����K ���͉����}�!�I�'Ul����@��:�Y��!��Sy��Q�"M�B-R�P4�!�$Z�Y8ht�f���(ph��g�ΨK�!�d�)Q���5�:SUdɱ�J�)~�!��}y�-��Z)9ڌS�U
:q!��?�z�acM�5\��
+k!���Ҡ�Я6�����S1�4�+�'z�Tp�Ѫ>kΝ�`��/"�	�'h��F!1��X0��'��<��'�lQ� F�x�Ⰰ�"� �j�'UR�+��̼\��a�Jٍ0t{�'����r��6S�i�E.�)�Y�'늈�ǯ��P�lŁuiJҶ��
�'���hl�y�TZB%֫3c��
�'��X��Ӊ���z�葍U4<��'��R�rI ��R.T�f��'f0�;��ƶAB���m�Q����'=|ݚf�&{�ȨQAقA-"��'XM���=�hi�bV�f��= �'�,zG�q�Ȕ�ï�q�N�#�'��X@�I
�*D��㣒�f5D(��'����dK�/�
��o�>X$x]���� �9cAW�Sj�T����{0�Q�"O|��d��D�D]�
ГG��I1"OP�2��S��KH��V$r"O~�!u启3�p�gǒ4	ޠ�"O�az��Ş/B�% V�e���`"OdL�Q�ԲDP��!ʵ1��}:2"O>x������@����w�9�"O@!���Դ��L�֪J����"O*��1Y�4�6|H�Xh�t(1�"O&D�	˔Z�S��8���"O~���'�b�� ����$"�$�G"Op�K�$��� s�h	-lX��c�"O�]�vi+9:p��F�>w7
���"O(�F��`s�-�3Ô
	%tpp"Ob�(��ɣZt�RQ�ɆEi:��"Ozh8���;s�M�a	�#)2@���"OV�(#�_���x�G(���0P"O��WKN�Hn,}!�N/6r�"O���&�o�
����I����"O^�[jN'T�҄�09�ൡv"O`�9R+Z�2D�f�	 S@�t��"O���l��/r��M�<F%����"O){�� 	��k�d t"O��PO3���I������"O@�e���a��My���9U��Tq�"O��x� 4&��)@ݸ=xA"ODL��,X�]c�`�3�ЅD�콘�"O䠃g'Q�"Y��Y��(��"O"�M�/$�>T��H)u�"p�&"O����݃'��l���ħY�ȀP"O�	C4�rO�U���-v�4d�"O�ԡ�g7�ڠA�V's�>�h�"O�y[�k��AB0@j��]�#�
��C"Ol	�����`�I$P�j ��"O���Y�+�JZE�J5T�6�g"O@��&�p�����(��ᣲ"O͘�Ì$}�y��gE:T��Y�"Ot(�'�	v�ε�a��l��8��"O�TJ
�����u�H�C���Y�"O�Iʄ�D�#��P�@j�;
"X�&"O�s���x��y9E�)�b���"O��3���iel��C�cp䜑P"O �js�*��y�,� U�=�"O@�6�=}}�X9s��<JVI�3"OP�Qf��DnX�`#l�>����4"O�i��,Y��H׷W�f��S"O�T�m�,1��h���B"Of���e�}x����݈Np����"O�Ik�cE�e�6�3U cq,;�"O�[@��'1\�R@D�Uchl�Q"O,��ԫR�$�\ɰ��)HJ�Q"O�aREY4X�\����ߍ78PK�"O(��)��96�I��_6?ֆ-�Q"O^�sw�0Y����(kǆ|�"O,�{c�0=�r̩2A�@�t�Ђ"O��ㆢU9��0����3J��e"O��Ð>Uj����.HD"OV1ည#<�� =j6HȔ"O ����x�hT�#o��v����"O�0�#�b_p
 �0J�(��"O���`�%UM�0`S��"��L�"O�`�Ƨ��x�V�^&5Ӹ��B"O&T��X���1b�-,⌈�"OEJ��+��P+w�"pI���$"O� F���ǌ�D�64��0_*�$ �"OTy+7�P G��9��n߳<j�"O��P�R%5F�5�q����m
"O��;���l�d�Ӏ��i0.0"O� �Հf����S�`�f�A"O��bUcQ�S׸��$�CN����"O��Ѳ�� P� Qz���ib�x�s"OnD�t#;��1��̮xY`�"O�  M&Z`p`3��<X,�s"OJ<�B*X�34*0P��8?>��"O*$[7蛭ye4D�6(N����0"O(���$۔f�xx@І΍Fi�(��"O6e�߆$laH��ܪPֵ9�"O]��j_E���E�*d1R	�"Od	���Ť�HEQ�ā�}�hAD"OT첔��Yc����Q�p��:"O�=�m�#U"�h�BϫP|��I"Or�2���]�5�$Ǜ9lv�;�"O�`�eF���Cm��e� A�"O�Q�_�\84M�)up�"O��40�źQ���s��\��"O���3K�R3D�@N F��"O���
�>=���7���w��9�5"Oڤ
��pĒ&8?�d���"Oj`0��O"X��c��w��*�"O���V��d�:��T�I�;p=21"O|�yQf���V\��g��+PR$��"Oʑ"�@�,�vѠ0AF3���"O�p��9��FY�Tz����"Oޕ�6��p��m �Νlt\���"O�X��V�{�hd�A˜no��k�"OT,��g�r���	���d>q��"O��@�Խb����AçJ$���"Ov��6e��͂X�FU@�@܉a"O�$X"iͯ;(�|B�G^Z�X�"O�1�e�2Y���*,����"O�|�wB(:�"��g��D�"O 5�ǧ�7`Oz�{6+�t���	�"OP��n��|����i����ȓw"O��3)ʷ8�^h�h "I}�:�"OBY�#�:p��%��>2��#"O�A��m�8~F�ź��Ŗo��աp"Ot�z�"�$���c�d�RM��"O�Uf5o85��)2{��j"O ��E�}�fiQ8\R� �"O���fJA�aAzܡ��E=P%�K7"O��#�A{Q<���G�U�Vmy�"OR�{u�+~FRiZp�Z��W"O"!�2�Z�Q�� z d�0���Ѣ"O�z2�ԣK*���A�`�Cu"Or�3��љHrD��%�n��2�"O4T
"J�	fnfQc��Z�r����A"O�� �߯��1�d��>h� "O������i<Lɴ�۶8�8��"OL���f^��(�ҁ L�҇"O��5�Ė�neӆ!�	AO��"Od͐�$�O����jլ`.L���"O�e���B��гj�"v��T1'"Ox�$�G���a���Q���"O*��׀<9���.�/p ��"Oڵp�G"m܎x��c2��y��"O�XX�HҧP���B%�9ؐ�X�"OB��sC�'G2�1��	�@ў<��"Ox+0�Z)[J�4� ��>Î�0"O� �`Q���%WN)�#���C�J�s�"O��{�����4	&d_1 z���8O�2�	�gM�){R��>���T�I%\J5�"��"=<,��v�M�t�B�	;(.�`]x)�(׽w���"O�u�w/Z�~��EK4���xcRL��"O�4�뗓4Nj%�"��fv�[3"O`�!	# ��?7h��"OF+a�O�u�D���$�XE"O��z�R�[������Y�Z��I"O�9ZA�(U�H����Q!&�(�2d"O#��I!g.�Ҋ�$���"O���V��.;dܥj#(�0D����F"O<���`U�!.x)�`&�e��I�"O�e�u�/q8BC���R.�c"O����Ꭿ���˥#S���)Ѓ"Of�����)�~5�B�G�$pP�"O>���cŠMf��` ��JTJ�"O���%�g0�3ƅǙ]��QP"O���M�{~��J�d�<�$���"O00pq/M p�8�0`�.�����"OٱP��N �B+�f���D"Otd�g�Y+ �X��` W��TI�"O��$K?U�����I+\����"O�xr��q��2��`q�1s�"O(����`xR�����"3ݲ����'yP𩦏����I<�M3��A�_~��{���>��C����D&ǈt}\�I6H��E��O��0��/�NA��S#5�\0��՗P{�P���eK�C䉀LBb��o�8�8�#��.�dDl~JG�n�E�}&�P��ŗ�J}�r�I��J���-�X��HŤa�@)�թ�m�w
5P�P"�*�QWR��	�~$���7>ӊ��V��nD�)E�`�E��hc�Z�8�Y�O��0����s��y�t����d)�'���c4���{4Jݲz^�	.OvT��P�p��Uq��ئg�Q?������Ҵ� �M�;�ԍ��2D��KQ>!�X��L�ww��B�됒��3R��\@�(b��g�'��Pz��*��q���\�8��
�� a����I��u�G�ۙZTt���J^��lS�ey릱�5�G*�p>i"�ru��z��_�hM6�k�(d�'��PBB΂�qs��"ge�*nF$�[�h�?���Äjj�ه�A,1}�]X�-3D���p�	����Wl�U����N8S�(!J���}2�Q�k(┋P�sމBO�=���fW6٢'�1D��g"����0��� �D�ĥ�{/>\��K�G�:�H�m��GS��	C�	�Q�$S�`C����B�^�,��٥i-|O�9�"X��U �b�j�ƽS��!��D_�Is������(C�n�%�'�>����&�PK���M*�@ی�Ʌ�k��Mru)F'K1�i�f���H�X`��O�@� �B˹f�����'Lێ���'��!�����H���5:c���t�P�v��L� �Cfa��f�O�����9�N0,u��@`�ITP*f"OVM��� R$D�R��@Pb���T&T�p�� �(�0�r���6�VI
�	�(O��+U��)�5��hK�ء��'Lv(�C�ӵs����sO��b�n �@Y�U8v9Cae�1��Q6��6��j�#7�O֜�sL�6��}�mӐs�81Se�$ȸA���RdF�dM��1�Z�h����	j���7��� '�1>ʐ95ÖX�<�Aa��8�1�V(]РȪ@ʘ�0i��I��t��խ˯�!�N!��9*e�.L�})�@�U�C3�����
n!���w��{��V�E�4bG��*z�W��b�t���1%}��灋u�
�#��$��Ր�8�P��ӖR���	;L*ͣt�xt�m�eN�"��<33���D0��_ad�]iB�α0�`�H	�ў,�e��
GKUh��]�]�=aҧA�*�T�F.-Z$b�H�2%x����`�	#.Ti9�4;��I^�tUz�"O`���N���Ф�1�j$x���iY8�q��8	K&�+�mF:d#|B� g�Ŋd���wb�lb�d>��pYA�)D�,��S,#�:���PEV����.�?�2��HC0iN )hE�h�J��͈O� %�tċ�!|��s�բNV��j�'(V=��ݯU1�D�σ����Q�_/ (��",��48p��9�p?�3n^٠!�@J�,��ibV�I]�'ά1���! ��M��iЎod�U���X�D�Mc�I
Mn!�$�<��q�6	�ǐ�7*Ѽ���3ϝ7i�t�RH<E��co��a	�4�����?@�T̄ȓC�F=" b�^�d���k��l��+І��3�	"�NY"�&�%�U��͚�PV��wx��LL��ȓyy��^�qN�˓�0}��Ͷ�`�&�'d�ȑ���AEv`�ȓJ��I���@���!C4-cr��ȓ����d^�f
�\2��1}���ȓtx��sS���a
ء0�ųv"x��5L�Q� ��)�̉+ʪ}��7�F؃��dM ̣�Ů<����ȓn���B��N�J%G��Bu�`�ȓJ5t`{�)�{�h�P�#�<)��?Аp8"�!�H�m5>r�ȅȓKg�� /mYj٫���t)!�ȓHyL��"���H�.�'��tU���I�0p��G�3#N`� �fp:P�� 5ʽpbbD"'o~(�i�=b����Oj�3�K�?H�@� &;���ȓk�PM�u�BX�� � `v	���<�b��%{D��A�C��y���� �`9cB�4�l��@G���a�ȓ8�,�X�%�%mAԽ��O(-���ȓU�*%Cbf�`����!�!�T�ȓ�(�p!#٦
���8��V~I85�ȓsP�ł�I����"��-��|Hh��`�v�pJ���,o�������i�72J,:��/!JU�ȓ�栈�#Q!��Щ�a�%f> �ȓm��0��'	�c�:���6h@ܱ��h�~��-N7S504�È��:���ȓT%>l��@�xH֌�V�Lv�@��ȓc΄���7����P�u:���f�`��+��vRjEC�)a���ȓ&fND	V�U��<$
�	C�M+�ԄȓQ�4UIM�0`�����>���ȓT�ƴ"G"ݡRc��K���(�}�ȓ>��;�h .�̡�h�&����_M�G��u\�4n�=s�]��K��s���M�� D 	5b����ȓ:JR���X<K_�Fg�,|�Շ���' L6}@�գӬ��(��ȓV\�#AD��Nᴨ�t�x���t(UA�&҇h*��8��Q=z�<��a^�;�F_����H�8J&`�ȓ[MDq 怼mH�*� C�M&���Wf��pB*B0Q ��
�+@�g����33���C*j�t˵�V�>ن�+\�o�9�h�Rs��[JC�I?|Bvm��/ԝf�$��ī|p(C䉨1�@��C/2�Ԝ���h^�B䉱g����(,�!��N��B��U`��4�͚;i�A��44H�B�ɩcn�0"#���������B�>W>@)81c��|F�@��$*�B�ɜ[M�B�L �gv��E��� b B�	`��ѱcǆ(� )�¢��/w�B�I�L��@��	/�8 ��w!�B�I>2K��"b��#��ăd��5��C�)� P� �)�0�����o�-�.�ja"O���k����S�R�����R P���Y-#�ؼR�&� |�rݚu����!��=-��bDyƜl�s�+l ���B�*)G�W�D�|�',6@��
鈠�eO�N4��	�'�$B�&ʟ��U
]%+=�����%m��ɡ���P��Q��/h(�S$D˲��"5�E^���ddHZ�Z
"���%��6@����*$��T����V� �ȓ5RvȪ�%x��qh�-j4�`&�$�c�-X�f$�Ԇ�[��D�t��=�&��r�P��(�(���y�78�t��c�@��D���;�A�H��I0&(�	K B���L>i��',3��U۬a	,l�DK(<�LӒ\��Ms��?P� m��f�#|x9��n�6�j�C%Ȑ�Jh���ۋ<����P!o���h�H�+_ax�F�E�YkDυ�@�L)��M�Y���R�P�C���C#�[�u�Nyx7O��)V��A `�b��H��[p�� �e����yv`�1̚e�rhB�'q�iy@��~[� ѥ�~�b�ȓl�}�,F�K�<�B�,D�u�����v��TO,$�ڵy4.�U̧��J������=9����a�?B��d���J���B�� (g��k�OW�>��s1�|���`�0Xx��+�z}����	�B�X�S�&S�Ws@�
�]+FP��D\�4�D�ʳ�;1�B��h�\/`u���� ��YpR��ފ��'64�H���_5	�I[e��1���P�#?��J^hk^9#� ӄUd�������O���нXh���܁V���`A�<�`N�9
FF̊u��$	d(���� ����d�[��A� ���-�|JJ>q�ID�xs���')ɟ9���X��CC(<�����I��2��ES!�֙ZJ=j5���I��{ï6eb����0LO�Ic��>Cx�I�h���Qf�'���]�m���q7�ټl�\�GC�<� 
K����i�+�{�<i�!a�:lC�e�(&����Yq�PHѓ��3a+6�B`�G�O`$����H� 1�O&�I��'%�#�N���kd�����<w��� ���Q!����ē_��YunR1q9Q3%f���#�:I�t��O!�	�Wi���İ��S�K� ��T[z�d�������#''Y�t�" ����zR�ɖ&ްX�.�<a��~-�j�eq���7(T��[4ʋ�z�Zd�Ѝ(����n-�ɷ}ܩ���Ӗm),��ӴH	�����
_1xC䉯#x-�դ��yDbaQ��2"fB�F�6�s�� �7$X �@^8�"B�	ZeހZ7�N�Kr8��O�<B�4"Pl���:6b|��.@�C�I�� CS�F��Ll9��5�C�ɵ�,��N(�h�Rޜ��C�ɦ.@��''�<�P%�	pxC�	H��h#�K�/c���a��%"s|C��v�0�l�_��v�� ��C�)�ʤ;�L��qe�	"kb&B�I,�4�⫟4s: ��D�DXB��\\ ��k��'�� ���P�NB�>n\~�p �i{��rV �	lT0B�	�l�Z�H�#V�
� j�\�4B��$Me������1~���p�o�"3��C�4F&�`2�`���x9D-܈��C�I�R�<1���N��0���k|}���'b����&Z"��A$�^�i��)�'�8�#�$�L�n�R��A�I��5�'��H�U�y"H�8�*�Nd\@�
�'���bAH:T)�9��ñEd��	�'3-�ph@� �J�h���1�'i�(��@L�9@�ۋXa"���'%t�(FP�[����T���Y��'\�Ѻ��P�T�d9�S��${��5x�'�Bm"$�d:�$�L��tV`:
��� r���ܵ��RӎM�e؜��"O|��h_2Q����( ��5s$"O��	Y!KV��c�h��- "OTI��`��I.��B� @����A"O�a�-�k��x��[�It�41D"O�
�'ʤJ�8�Zs/�k^��F"OF���1^��r1��=@��"OB12��E�_:.�A���7:����"O�8!�B�<Q�U�K[�l&p��"O���ۏTR>���Ӡ	���Q"O���#�UM��Q[g���zP��"OJ({2㗌E�0�6&V�
.�y�ϛ7�` ��,fK�B�y�� �2�y��������һ�y"@�&i��i
�Z��8J���y�+:�DiRS�U�T��1H�N�y�Ə;t�!�MO@[��so�=�yB@�T֠L\&Kk���E$�y�.�.>���e̮Mx|��.��y�A�'М���`	�:�
HPG��!�y��Mb��%�P�>��(�l��y�6(o�A"�i�8�sv���y��%Z����O��>K`0�ef݃�y(�|��H5B[2�R��,�3�y�}=����Ҭ~2aY7�+�yR��Y_@��MϩFH�b�Ѝ�yBC�)=6IK�&�H��%Xt�K�y�A;X����}���@����yB'M�8|p���'[� �pV�Z!��<y��'Z�"��O� 9!a]��x�:�!3��(�W"O>���Ōd+X���	,p�N=Hf�x���Z��b��.�|�V�E�w���"��t� }�"O�)R�cL�a��`!��o�r�s��#G8��!���(�3���] Z(d@V�W���a��*4o!��_�IP��2.�ia��rJm�V�\�f���VX���G{c��JS(G&g���+�J,��|7�qV
#��i22��j���73�9jB��Z��Ԡ�M�W�<92&�!~�6��1O^�Hq �Ly�˚�=�(UPBD�D4��A���
�b��!	 ×&1�R\��O�f!��N�'l�%"ժ乐L?L*��� F1[�(Rq-���ītR>�<)���2d�T��*H@��a3�EX��	���>	��!��T57���9�f\�l�Vm�zDTi��J0i�m��	V�ِr�-K`Ŧ*츣<��[	U����ϑ"0��E�(���I.�qSBC�)��Taua�Zm!�dS�0� �@��+~�Mȴ<[29�새C�ăZ=��.�`D��w�<��
ʕ"�~�q�B{��	��'Q4�dh'p\�q�@'s�Jl��%��I�v`z��D�3�Tz����T�f�'�*9�2G�	q��ya��
�m�>�@ߓ6���6���1�<�R���u�F!tf�ҷ�֩=����\�
An�a�'WtȐ�I�| v�j�۫I��j�)�=C��@��~��%��5S�6��O�R̳����j��L�'Zf�\:�'�J���l�?�hqfMًRx���eo*ǜ�ch��`ي�PUg�\�B����;�U*�X?URj1@eD�j�b��"O�Yb��ͦ"SVjŤ�/��̰��'s��`z�#QC���2��<��]z�
��(O��D�+�8ӕN�0]o�m�0�'�r���sV8��Y�72
����P|q�܍!E"��C��Y��(�O Y���/-��1Y��6�(Hs��If����	9(�`U�5m	/킐i&�S�4 QT�+6�]�	L�|�2�PV�<q	̋�7�����ڞ^���H�i� �dC��z´ى��Ld��b?A{�3�ٲab�OIE�儉{�ə�"O�Hq��͌3��ٙ��W-I��q��a)��hSn_N0f��tO�R�@Q���(O�� P�A>�*)�A�ĐLV�K��'HdH�D� S�HիB��A�M�ɷn�F�	TCZ3`��S� ��u��d�fM4�O��4KO8-�앪�ǝ��֙���d�P��m
� &\q�I9O��=�zm���~� `���b��ZT$�x㑰�4��"OD�w�V-4�8IA��:��(�&���~�
����WGL���L�jE@#|Z�h��s��vk�h8��.ڦ�K  8D�H9 L�=-�d�3��Ažxc������b���;�)4l�6D�&���O�]۔$İ#�H���ᖡGDb���'h	R$��Z~�I�����H��'n�8?W��DFnn �����p?�G*W�DIh��:\�<�p�OFx�',��('T'�^����ɗV��-Rd��P{��0��n?!�d�(Tw��D-��F}鑦B1 �f�JU��L�6UI<E��FX�d��釽'�z�c��b��Ԇ�1a$01  !�(��o�pT<h�� �����Uc�I���y(��1�.!��{ D[���-�����:L"P�ѥY�p}[��Po4���ȓ5��-�Q._�2i��MH�kE�M�ȓ��b�FK!M�dE��H=�0��[�C6��,lm�C#J�&�hd��V�r�d��_�$y�Ҥ�M�L��ȓO! ��B��t��j'[3e���S�:9��/�&$ԅ��tO�m��Z��[���
�W&L���0D�$(d��K�¬:�I'�8��tc.D�LP �A8
�&���ȅ,)DܻqG,D���0�Վ9	���"h�Ь*D�26��(�a�v�$aO2�f,D�t����W|tD+a�Y t��;SB(D��z�V&�8��wBU�.8��d�3D��(WB�8�FT�SJ(��͹%.D�����~���&�h�"����0D�:a%;w��|	֬�LS$4�$J/D�x
R�0����
�����IcbC�		k_$]`��ܼ+�k���6C剋=P.��ǋ��>k�����!򄏑*�t����+2nٺX)�ࠇ�B|{�������?}����ȓ434�;v�+�|0���y�虆�X�*�[�&��~!�)��^�Q�ćȓh��p"/�z^�҅O�<ל͇�j����W� ��j��=Jn��ȓ��ѳ�N� �>�!"�VXr%�ȓ7?j0�2Fؿ/��XrB��q��[�	H�ܷ%�H$�\>% ��ȓH�@1���:�j�;G��4>��,��gܜ���k��˕ŏ>:H�<�ȓH�`�p��V.}~� 3G�"�-�ȓZ��:�'�/i/B�k��*!֒��ȓk&�I�שQ�u����s��:�L��ȓ����@/�ڠ���O�����ȓ7��D��(��A{�F�"Z�h�ȓH#@D(�� )N(��X�����ȓ`Ĭ�`�4@>��bݗtF`t�ȓP.:*�/�2i]��i�LM�X��^�q{��}CH	�s���Y�����YJ�eeā+�|4���7=�����|��i葥E9jrѻ���1`bv��ȓ.f`t#�jN��b��a�A�8AV���cH~�)�I]�+�4�@)�O����Qf(�j�9�Ȁ��CMOt-�ȓ��)�cŊ5lh��s6�
�c�Tx�ȓfo�(���;e|��%�v����U�*�󓏋�[>uۅ�
�8& A��{��yÅ�S0��ǥy��ȓ8v�� OK��~d�`'��P�X���i`�V��_)�)����i�����S�? �M�� ��I��`�g�P�d-Щ	�"OT���̢Z��ĸ C�6���"OИ"��E�	����磗6L]�9��"Od-&K^�L�� 0�kA@P��"O&���P4I�dA���:;��T;""O|E����;`4���\+�H���"O� ����8u��<8�M�z�x��"O����պ:�F$@e%Z `���"O8��r�њ�~pA�N�O����"O��bVe�#i����Ղ�5�$XF"OJęC� �6���H������4"Ov�@��O�1�[#��1�"OM"d ��/��:��
�w �k"O�:5$�=���3 ^=KGP-"O %�rJ�p�4����T�QK"}��"O*	s��(؜����w7&���"O.<� �9K�hZC�Z�>&t�w"Os�-��c��MXT�@�t�r�"O�|:w$N)
t������dRm�"O���G�$md*��g�ܙ�"O�(�-��Jw����f�k�
]��"O8�!�O� Q� ��ƝNp@)5"O�[$�չc�Eb�G��pX{`"O�):
��ܙ`t���0��|��"O��r��]Oi�i�w�
�� �Ƀ"O�] %j%?���ք��c�,E	�"O"+�� �vZVhcUȚUr�p"O*��� �f����O�B�Q`�"O��Y�#W�8��su��3����"O�z���v?�`�re�b=���"OZ�F��$`�t����` �:W"O��s���5)�2��@�Ch��c"O 5�a���9�,8�P�V�v~��1@"Oq
�ڥa������]�%J<�R"OFH�4#�Zm�D���x���1s"O�uf�һ3N�聠0;��{�"O<Ԋ�Ć�h��u�2f��	�"Oz�ӂk��M��5�RװYq ��"O@4bL=<8,�2�,�D���"O�uK�ýN>� &�Lmb���"O�3�6_MX�#ӊL	���Z�"O�A�َ$��Q��S�q�B�*�"Of=�q�Yq�"[� Pq"O��z�GJ�q�j�3b�$��"O$d���N�LDRT ���kꜽPr"Ot��OΘ@�n��Џ"�r`"O
cf�P���4��i	�q����"O
b�b�=��0�J�U��Q"Od�����o/��Re��)犄`T"O�ܪ�儺C�A�t��.y#^X�C"O^=AAJ�z�n`!T��<^$�"OF�j�Ğx�Y����/L� !�"O0�s�܋3KH�rF�6v��J0"OX4p6�6~�Dd
R#�= �<��"OZIr��5E�8\Y��4���+�"OND�2I?�ݘl<>�P�p�"Or�ѵ���E����˟�,_���"O��j�#U�MX��0��"R�9@"O�1ᐄ[�N��;�	���4�"O�`��)I�w�:�hW~4��"Ot$iP�'{�u*T͋�(��"�"O�t���B�l�
��L�K�2t��"O�	�AB;H��C�_ x�~E�G"O	��-N	A׀|��o\�J����"O� 8 �mҒ6~"z�Ο�X� A`�"O��a�߰Z�!bv,�K!�ya"O"�Kr#�
U�T� ӂ_��"O�)�ʟ�{NY1ԪB���A�"O0S��S�s�J!0�+OU��yA"O��{LC3����+ȑ6��� "O�}� -�hT�y�T���k"O�Uم��8�jt9Щ����"O�h�hG��t=� ���Vr�"O��K#'ц_|D�PD�kjTah�5OQ�5�ՉbO
��V��QQ��3��I�u!νSŐ�k�H��aɲ(urB�f��j��P�e���B���N�4B�ɒ"�@0ū���L�Vi�;$��B�I>�N���[	���Y'݌Y����$=?�v�Q%l�L�fEg1�����<1U)̭�X�h�Lߌ�Dtm_R�<9�iQ0
��Y��A!c!�*&HPQ�<A��R,p*���I�>r�Jb�s�<!��-��`��
ٻX�`h*��k�<���5��h ���3^��H �h�<9F��e��x�cŋ�e��8���n�<)�$4�r 0�O�>���A�O�<����*�X�YfRi�6���m�H�<IӈT�\��	VbP��r"�i�<�4a�`��$Dċ>�i(E�Q�~!�����H�&C<y8����%\�dv!�d��?� �C�!T@�D��"eM���P�x��]�ïIS,�¨R;c}4�Gy�gS:�ȟF�{4�ɦv���b�D<g{�ls��%����s?ѴgF�y�D���菷l|�I�c≟o���?�~2�	
'��+$�;{�4P]}���O�>�h�,�I/b�2�'%�J�����Op�����S.P�(�2BՇA~*���@�U�8ͅȓ>��ȷ������c��1>IU��\�܉�K���ԃPzb֔��8�"��C�N	��@ϕNL╇�srL���gֶO�ܳ�D�&��ȓ �n��v�����B�-@>c8,��2
��G�]�z��!�"i���ȓ'�*�# �k�^����[6X���ȓ �v���dJ�N-��Q�	�?g�L�ȓq��,��Aϡ~����S�\9Fຸ�ȓ&��`i��<}��T��5+�H\�ȓ��HӀ.0o#R���'�4=$�ȓ�
��c��:X�n!xPl_O9hц�?4�mh����ko�$�0Qk�2��ȓc�$!Qf�"����6���2�J4D���%��,��LaE�&*vH3j1D�P��^�S��v@Y�u��8�ua%D�<�g�U�y+���� (_��0`��#D�t	�߫bB�x��?L� K"f D���7,�RXB�ܰC��L��(D��Z�	]�o�z6��qQb��f�&D�������2e�f	U��ps�#D�t�  ]�~���{vG� ^��1B�,D�����ב�T�� Iu��Ġ��)D� ��H"0�z��ui\-dF�@c�&D��)����=}���喴M �b4a?D��ð	�	�����.�:bV�!�%>D�LX��� ! ,Ƞg*ԟC["x�ũ:D��p��� .�`�G
@�����4D��x0*�>�.4�CH0=А�f1D��C7.8AB�E_�j��7�3D���C&JK�L��	��b����'&D�� *Y�Fh��������e(Q�"O�E�>bp�D2u�N#U�	�r"O�q �D�*u���'D�1���"O܄�T@�3q�I2��! ���yc"O��R�6J�#�3;g�Kw"O4l���˱8�pœQ���t�8+d"OL�{A�3w`N�� 
�=v��U�W"Ox԰�� 6̺)9Djx���"OZ#Ǖp�T@��.[�*���"O���S(Qc�Q�m�/�R���"O:��TfàkJ����%j�F)R2"O��`-��P#�|
F+�[��X9�"O�u�&�+F$�*g��;vR��x""O2`
V�@�/��#5�֑R;�`��"O(����(|@���	><?���q"O Qp4�N�7-B���>�"])F"O�xZ%*K��.%F�N�$uڂ"O^��B��?�R�ݭ�d���"O�x����><�Đ �E>�^5�"O��5�C���Y�(<8De��"O�b��U�j�a��H��Q��"O�p���'�(Q�GL���"O����W"�vXh��I/����7"Oʤ1ch�(�,���$]r�AF"OZ�r!j6��T[ƀ��@@tq "O�E۶�S�bJ�銶o�H�����"OjV�ߞ�Ъ�LC%abT�"O�IK"c��ܬ���@�1J8[R"O0�%�$#�nAηh��y�"O�܃��ۂ4	�ԩw@�-sp˓"Oh;F� 5�
�aT�P(��3D"O�,� 	��j��ى*@z�h�*Ov�r&�u�@�y�ƚ�i_"���'$2��p͌*A�HU!�q�F��	�'�<0@șv�j����i�*Ʉʓ+�zTӲ	��P�~})��T&���ȓ���dg��\�ty�#W�W_�<�ȓ<����`��e��A�6c�@���p���Oܡ ��5�&A�V��Նȓl���	���\�ʕ��SM���ȓ���&��Sb�mj�l��xՅȓ`gl �7�9u|��5i2kҜ��ȓ9��\%�ߴq'}IVǓ�Jl�ȓQ`d��rE�7���E�.v%�݆������C"R2�����&-A���ȓ��ؠC,?*�;$"S|�`��jTj�`D�4H������	A�"21�P�UA]��3��A�[���Rv�qH��	�v�L8`A^�&�E��/NP�� �O�G���:�)ټ^[譅ȓ"7pRopܼjucC��a��Q��!��C7l��aҠI�/'��مȓp��Ⱥt섭,Y`��mHS+b�����`*�_cV�X��(X�MX�]�ȓh<�1$eӘ:��!�6`aeڠ�ȓZ!J0iԎזNH(С� `�}��p��P�#d�?HZ���M:����ȓ�T��j�6.$�Y'NI�Y+q�ȓe0||iV�S1x�`'J� C�I7��H�D �)SiFSULT��B�I�!!�,*���-�H9��U?Xt�C�I�A�jXS�n��W����˕N�C�	�(��)�)�Yșj��ɵ`~C��/h�V
U�E����9Roȷc4xC�)� �9�W�gx �q�+ē)L��"OJh�����k�*��0�1"O� Y�Bį���E��8�H�"OtJs�ݒH0Tq���L�V��"O�R��:8����D�W#�a��"OTu15#O�k����ViH�h��XQ"O"m�b*��0�%�׆@��1"O�mR։[�)\�[1f�6&�!ˢ"O�4�#��U��]��dN�F�x��"O`����K{$e���ڑx���"O4*
�MkĠ	d�ѦbnV�"OȀ��Y� jàB	 ^B��D"OB�"�>��s0Ӏ	Q��j"O\�y3F�t��B�++h�T�s"O�yx���u[R��!F�/h���"Od�,ԛub��Iޡh@�"O��!4*\�'$��"J��?��<`�"O6�ӣ
 �/��-Y�'� c��"O`]	aN�1R��6��<#2���C"O�yWj�
&�5�f%O�!-l(�"O�2�A�^#�����ֻ-�Q��"O��Q�K�L��Cpc�3%���h�"O~���X�`7٨���$u��"O�}kW�׆>IF-KQ�¤v��Dڒ"O.����ZYʍ�$��?)P��"On!�`Z�ihyA�A\<f;�W"Ox����¢a��|�� ��#��"OjY��Փ.qN�JV�}�r0�D"O�u���1,�n�{#	��� ��"OR�Zj�X2�gR�q�L��"O����	\�,��Y�q�51�
�za"O"���O�vM� FD�i��"O�9��%Gl*���Aa\袷"O�)H�k
�s
�%���|g���"O2!C`'%	�@�i�#�[�j"O��7�F�u�()����	~�Duڴ"O���'�PL2ʴ�C�>�@dZU"Ò���A��������v���"O�ɋ6��68t�k�)*�n�cD"O�x Q,F3m�L���*Q�X�"OSVC��{��Y!�fյ*5��t"Ofi �
h�|�p�]�fä�1�"O�P���%^�Y��	�n���B"O8���(�=a5v�HrV�O�� ��"O�9�@�G�]D	��M�V=x�c"O�؊@&�3|�ؼcr�Ҥ"L���#"O�����+G���r/�-X�����"OB�+������pB.��\��4"O����E�r�Z���ݥN���i�"O|� E��5�H�8S��=v��l��"OЅ���* ����uΜ�m�>x�*OLd�0��DN�E��>R^ԙH�'À��W
a��$ ��^-Ch�H	�'?��K���Ү��k-�y#	�'5�V��`�F��V ʧ�.�H�'m��U��-�<;�M���Ը*�'2�LÓd>-��,kS�M�W80�'�I�d�JQ�ޤA��+8��)��'�~!R �Q%�T���;4|NE��'�zxT��?@5X� li�'�1#wiI�`l�0��� �Ab�'v�p�[�^�*]��/$�ܬy
�'PB<��J��j�:�eQ)�Y�	�'��+��O�0"�S��L|O\��	��� � ��ȭn��H[S�_�j��'"O00(Uqz�����t��IX�"OX��F�@h�!�B��ҵ p"OrYb �
K,юͭr��с�"O�=��J1fQ���m=� ���"O\�Bb-ȯXr���b�
t��5r�"O�i���!]�����)c5��A"OzyѰ�E	+1������\�PB�"O]��n�'��� ���bdʔ"O�x@E�[�<f�f
P	�Rp"O��"��%I�$��qD� K�\�ȣ"O�͋B�цdf>�Y�cL�L��"O��br��Mx'lF�iϚ1jg"ON��̂�e]�-��+���lK�"O@�ɗH_�B4*�4r!vx�5"OĄ g�U9��d�wD�J"8"O<� 0/\�*��x�'n�<�V}[q"O��B悜a=��e�/��|Ѣ"O�8��O}ȈĻơ��6�d�"O�A�6���5�Hf�!�.��c"O\�k�痞W�UB�ϥ(̔(�&"O����l��̡��J�	ێ9�$"Oڦ���j�P�ʘ�W��c�"O��CF�Ôh���*�q��"O�4cV`�48��u�a�#@�ppc�"O�mZ0M�y[��8���1��d)�"O�[��.������E-�6"O���ӌ��'т9J�"D:Oy*0h"O�٣����(�X���
NP�IU"Of���/�0a�$c��N�Z�E"O�h�4ϔ'[�&�i�`h� � "O�Q����%oن!*��^.l���"O� ��7���Y���4y5��ڳ��B�<�1n�8 (�X;��8g�Ps�Ș�<iP���w�RA��(C*.��i0!t�<9�㌈z{�M ��N��t�W�s�<9��ԭ.e>��&O�{m4@&�s�<����jJ��{1Ɣj5��Ѳ��C�<��֔Sٲ��ԯؒIV
�Q�ID�<�&��"   ��   #  �  �  :  +  �6  KB  �M  �Y  Ue  �p  h{  Q�  `�  {�  Ν  !�  e�  ��  �  ?�  ��  �  ��  ��  [�  ��  *�  w�  ��  �  � s
 � w �! �' �. �6 �> .E rK �Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*hEz"�~���n.�h򂅵,�lq�Q�<&��;
��ʰf��-ꤡ�A
L�< !�6I���JŢðP�65��K�<�)@�,N��d-�*��F.r�<��펄o5>e0���2h%��
c�Kp���'h\�I�Ažc].ekeI\�P�E��'}|����Vw&5[E�ғv���'��8�'�H�aj�أG����'���Y����Z�,�A�:\D��'z�Ѳ�*%M<�hq�ū7��a�
�'x��YGd�1+�-0�V"+��A�y��r���[��̧
ǀ!1��A�DJ�d%D�hy����1�R��`��=jT*ԥ$D�4�Ġ��e�P��FG�	Q��*D6D��:��2%P� ����"l !�䆳M�`����7H|ٙ�D�
G�!�Dg�
D��NЈ�$2�̅�!�YJ< �Uo�G!)Qb�l��ɧY!�}�°>�#a���DT���>!�O��S1ʋz���`�����c>O����V�Oh]� �0�<�SŎ�
gkў����i�{*
��T�Q�B�X�� �u!�D�M��PĊj��.M�6���)��1�'o�$^A�hZ3���B���@��=D�$�wC�M�VM��m�@`J��D#1D�d�� �h�b�wh�1�"RU�.D� ��ˇC��Sgٛ �M���+D��IsቁC�|�`�p�Kw�)��hO��SŌ<"��L7a�)@�P2qK&D��C�� T�E�B��24�ZW |�����D�"�B�8fBB-i<z`G�ܕ�!�D�O���`�l9ܱ�tO/]g��.�p?1!�W	}_�[t��>G2��!.�`8��&�� @鶃��o|t�勆��� "OJ�`�,ς-)����V�5��e2�"O`q20���O����b�H���c�"O�ڴ��;x���G
Ǫ��p�"O���W�V�C��5Rb+O�ZnY�"O"�h^�^��0�⬒�hG�\s"O"|�bM/12Mу��$>@��
�"OV�c 
XR��L�0L�T?I��"O�t�RŊ�k��j`��b�3���^�OCD�t(-�H=r�}�lX��'Xx̀���,��e#%��:n*�T��'�tp�L��0S���N�Z�'�-�n�*��MӃ�& Z-Op��b�Z�[f�ÓPQX�ˇ�כP�x���IB~r/9:h��J3�v���9�Y��y�$�!��4"F���n��ATI��hOh��)��?5L��%-D�q�Qc�T=y!�Ď�z.zݑх�49�L b�mL^��)�'U���IHj/� �իe4����'���A�ã�$��#ʗ�b0�'<\HYDkTq��|�"�1	WF���'��5sJN�HL)	����	��''d`�0!Q�JCN�Q1�Ő4p8���$�m�O�\M���[�B�ւ��.I��'3�]�F��+F��`:�F*?\l˝'"ў"~��L9fac+j����B�<YtG�A�*xA�Ų?j��PC��U~r�'#|��ƃy���E�_�g)6Ib
�'�>=�d �<vB��:ŮU5u< x	�'��CQn�� g�� ����0����	BY�T�2/J�����\��C䉓F,��暼~�|�� ��fV�>y�����3�H �(^<.�8��Q�I!�D�&P�,8��XV�tS�eU�]�!��([��u���j�X�R'��!�J�F�aG�Rd�4�����~�!��$��H���r�@A���[�=!�Γl
�`wW�Mǒ �rJ��!�d�>!�u��J�t��((q�V�g!�d��h8P,a��E�
�e��!�đ*؀�Q��D�2����Љ]�!��)W�J02�I�$�fX��o����~
���?�a�Ȑgj��(׬
�}�'�f�<9P�Q�R�A�.�Qb�%��[x�'$�?�Ys��&æŲ�B�-l$�(�:D�(V*��U�H���J�yT�2�g3D���`Q>����9 u�SB�2D� �6C��E^\Yؠ�A�c���j�"/D�$���M$R�$TH�
��XA��,D�`S�&:n�J,;�CU�R�b�+D�0�H�.�dZrd
�g)��G�'D���w�Ӧ8s�����L��\�	+D�dzC��r"ջS�� �֨A��)D��rg [H�B]�G�6Z�l$��,D�XS�B��Ak&iJƤ��G�vY�e�)D�p�(�=�(h)v��O�F]q3�&D���T
�9=��y!)��=1G�"D���rc��iQ���,��d�1�"D�<Ǐ�y��ā�i�
��@ C,D����]�Je�m:�*R)e�p��7i(D��9W�ʑ�d�c��P�^��"*D�pb׋!�RU/����M{�>��0<Q��E�(��L��̢��tF�L��\Γf]R�a���D2�uʒ�yw����S�? Ƙ��B�)k��h��ބ=9��3�"Oi;m'_D<��UNa{�"O$4�E��
S�p3K�8"��a"OHl t��.B]��Whҝ 8��"O���Bʪ-�|��fUC+D #ґ|R�)�H���/��U��p@� B�	�|�`�pF�	�K��y��G\�k�C�I�-=�S"䇅Wu�[��؀K�C�G�dyX�e��P.6y��&֒SZjB�ə�M��K36������>Y��C�	�c�j� 6C�n�(
����B�ɵ@�=)' �Y�8�y�H�'d&C�	�6:ة1�A�%ư��ʌ9z��B�	��~���Z�5͘�A!��m��B��6�:��1G 8mgpx��$Xn��Tw̓#��a�	-j�~� u/ձH�}��%t� {�,X�� 0�M�q= t��$���2�G�4��<:D�ۼN�x=�ȓ�@��Kɻ`�D0RRe�����ȓ����H��X8R=�TC�+�\9��U����Q�N�X;N=�|�ȓN���C��D��ٚk�����m�,4k�EǸ7�6�իצ!�B�ȓOla%��:`ƌ̛Rd�#IF<��w�Ha��Iǰ=;�NDS�̄ȓ#���Q�M-0���+���=1�<!�ȓQ��d{G�mJJx��H�a�t���
���S��b��=���7}�V|�ȓZ\����Ç��Ke&4�P}��+s�b���b3���E�T�$�(<��ZG��B�C��({�H��+δ���ȓ$a�Mq0o� ��)��ڨ*���ȓ$���	�(;�R�P��j�t��F'ܐ���2k�����O��ȓ-alt��(��(�^��c��T�K:D�xY��D0���BDO�4�����>D��#k "|�K�dA�j�|H"�H7D�� #�)8�p��ݮWtV��%6D�8�����p���!�b�J�*O���P��]0��I����%�ʁ�1"O�[`��)[���O6%à�ۅ"O�I1���Cc9��̋/zZFy��"O��"'��XG��#e�\�RQJu"O����H�����}�Е��"O�pp$��*�������t$���"O�M�V�g��I��A��j� "OR���I��5D|�ʖ��<+n��v"OX�CeF6�U��#el��V"Ol�pE,�<�@��9����"Ox)S0o{�b���p�8��"O��(p�ǵ �(���K�=�b�:"O�{3�Mu�l�ʴ���o�<-�"O��[4��Ub8!(��0äACQ"O,q���B�X�Z��B�;Z��I�r"O(U�e��@2��ƺE�T�H&"O:$��/K�,	��Un �Xt"O�|��oZ0���g &�j!!C"O �� �(#��;A/�=Y��i�S"O�<���x����@���I��"O�B��
	[�	
w�-��\�"O挡���0�`����,��a��"O ����
��`²�[�xA�K�"OP�4) ;��l��@�Q.4l�"Oz�y��OT��h����	�$(0"O� T��dK��4�1�tN�3~����"O�}1�dA�=�r��L�jx*�c�"O�P��O��_�k�Bl��3�"O�}cs������h\��9�"O�c�@��+�8i8R��'(H Pc��'y��'���'8��'�"�'BR�'w�hIeA�=gD��C��N�84+�'	��'o"�'V��'R"�'���'v� Tb��$&(�%�E�����'�b�',"�'���'��'�r�'�&i�#B�-L	��
wň�OT�p+$�'�R�'Y��'e��'���'�2�'�V%N�vo�8��aO=�(5R��'Y��'��'�Z�M���?9���?1dK_4f?�!�Q��bj�I+I �?���?����?���?q���?��?�Faٓ(@�8��8xZ���bC�?q��?I��?���?���?y���?�4㉷F�=S0n�w���Z�)�-�?y���?���?y���?)��?Y���?��FM�Gj�!p�"T�.�8�A���?����?Q��?Y��?���?���?Y� ë>�ʩ+��+GԈ�0EH]=�?����?���?I���?����?����?�(��f��v&�A���st�O�?����?����?9��?!���?��?��)ùG1Z<�a"����k���?����?Y��?����?A��?I���?�#�&hjH4�$��&(�S�BH��?y���?���?���?a��C���'��FSg�y�"�Ǩ)U��k�d�6��?),O1�����M�w�P�:C<h1��N�rr�$b��/bV1�'��6�-�i>�	��A�
�U y�)]�f���Ѷ�PΟ���K�x�m�D~b2�l��l��N�",|1�IV>n��A�F3]I1O��d�<�����K��ar�	9bJx��J�:D�	m�l@c�T�Rq��y�
�X��dJ��$ ((FC����'��Ĳ>�|
�#ŧ�M��'�` 8���lj|˒f��h˚' ����i�i>�ɞQ�t� �C�
y��)U�2���	`y�|��e��Q���Zg@�a1J�����K:⟼	�O��D�O���X}��׫o�,�6,��6!ڭ�	�����O�Уq)�1��ԫ���d�//p�c�W)�#T�Ҏ\�ʓ����O?牋ZE�]���R�\Z&�3����M�B��R~2�t���S>?�F�ل�[
$�|�P�N�W���˟���ʟ#��)�'&��?-�`H=[?��\�!&�a�I4�' �i>5�I˟H�Iџ��	�A�a�W� �q�@] �ݕ' �7�LT����O&��/�9Ox�j!�(y���vG՜/� \�p,l}� o�ԕm��S�'9h`ڔȍ�4�rX:����`^P�Cc�P.T�������9�ł>8O$�
]w���'�ŕ'����T�bz8��-
�m��P���'�b�'������\��z۴C���3���g�߲�k�����1�v�0`�4��'q��e��&g��l�<#+.���^C���Uj&�<�����}��[�Ƅa���",�$�~�D'���/[�P�lHҡĳV�
ْ�N�<���?���?����?ш� ��4^�)S�Ш]侴�B��.?��'W�+l���:��<	!�i��'�`1r�g�8Q���")�D�[�'�B���D���;m�V��0�u�$Yd��h4��;�)�r�Ӎ9�� �5�'�(d�'3�6-�<�'�?���?AӒxqX��EI�/�J������?�����ͦ��H	��	՟��O�nE�6��"�f �"�wQ��	^~�+�>���i�h7mM�)J$ϛ�+0Fp�5�͋D�P����F�x��jO@3��'��ם�U|��by�w(<�3�\*g�Mj!mQ4L�<�2�'Q��'���O��I�M{�*¼Vt`��@n��}����ϑ�}��s-O�nZ�x��I�AJg�#3~hhk�ߋF��y�s���M3T�i{n��i��ɠ2�hs��O��'�,���g֢+h-1�G�8^Ԓ!�i����\�I؟��	����I]�t��!�@�[DE!~�\k�Ğ�L?7�ΡvJ��$�O���-�i�Ol�oz��D�[���� ����;锽Q�C� �M�W�i<�O1�~ +�j���IOf���;Ғ=a�-R�y��	�n���S�'�"��'p�7��<ͧ�?Q��ѳS���3�j�.�zJ9�?���?a����Y�� �l�۟��I���['IēC�F�xUlD5f
9��Yy������M���iݞO&�J%9+]&L�^�U#pX����X��-F7S��V+6?� ����_�$���;�<L�u⑩g(6�ضgcmy���?���?����h����^"_]摠v��74"�0xхD�'���$�Ʀ��Gg[y�hs�V���#x��M�ѧ��0���H�L����4�M���i�&6MI�[��7�7?�7���\���R5=4x�(�o*ܹ�5a�1Zt�+O��lZoy�O���'�2�'JRb�P�����Ĥ?� �U�	q�I*�M�`c�-�?����?�O~��aߎ��ghJ)&d�����)��Q��\�0;�4J���C1��IA�I�����
�6%�.lK񏙜��m�2"�=��I�9���â�':�E�'��6M�<�%@ӲcX�Y;�.����{��C�?q���?����?�'��DL����D�$��- l����9��u�Ƥ��hPٴ��'gp�d����O$6mϢ(���#��G��R�lĂl �|R�e`�6�P��X�
@AI$��E�r�)����� ¼q	C,BV>豳LU��F� �>O2�d�O6���O����O\�?E��/�**�B�Ca���m�:��Z����	��d+�4}�Uϧ�?q��i��'����g`���u��@�$[�(0��ݦ!���?��p˝�)�'�I�Ul��J.Bh�2��J�t0�EV�]�`��	�(:�	��M{.Ov�d�O��d�O�4�DR�� �8)]n�Y��Op�Ĺ<yG�iC��{�S�0�	o��Ļ]���%I�:�L�o�n��I�����٦*���S��+Ѥm��\"��P6jyX�$Y?R���&�{��H�W��B\w�� �	�d7�i���E"ejD� H�CC8��!�����	˟�����b>y�'��6�ͫq�5�T&�3,��M�&�_)f���g�Ot�U���?�6]��l�4[�N<�g5T(P`'��/���4z{�TR��6O���ٞ%˼��'=d�3��}I���h�K�-�<H[c�i�	����֟@�Iʟ���Z�t�7��)2�	�x�[���&_��6�?D���O�d6���O�nz�)��5��
ɂD�"�(��4J��x�O���OF�e*v�i1��I��sS ��V� �mӯpF�0*0<9�g٤˓4Û�Q�L�I��V�";�� ��yӼ�Q䋆ҟD�	���Py�i�0�qu��O��$�O��2�XQ\�� �5?��h�0������O��iՉ'L|4zcgG,w�]@��(i�]��O��k���%}�V9봃�<�c���Q���K;���)������K1�}2B��r*���O����O�$�'�?�!�fɘ��eNآL�@b��?�t�i��S��'.�b�(��]̲�"s�(�x	t�9%E���ٟ����-w�ɦ��'\�B�.��?����M��!iŢ3��\@0�
�Wg�I'�M�.O��$�Od�$�O��D�O�иT�̩=_�h���'U<�!�	�<1��i�\$���'Z��'��OY���M;�$ش,=#<J1�B��(�,�@�Ə�O�O�i�D���>ڎ�Z�,Ҕ0������}�U�A���p��˓m�u�g��Oօ�,O�lZy�}'B-�\�(���#5�(���'��'�����S�$
�47�T��;{�@��V�a��!@ւ�]I@��3�v�dKH}��e�� �	ަ�s(%;U6��Ĭ��3���Ѳ�|o��<	�!!:�j�lZ-O�l�;����@� `~��REgՀ��MZ&e��<	��?����?���?�����_����cd�w�\Y���^���ҟ|��4"����O=�6��O�����!��-j�8�oAQ���r��|��i�j7�ퟜ��E�|Ӡ�蟔ذ)��$H�
Y ���cL-;bq��'��&����4�'���'���A* �3$��O��'^��q��'��W��۴MU�����?�������<���$~pp�$��I0��$�O$��9��O��T��	,��WIT���}�`�t�0�x>D��U����x�D�E��0|�L����dE�8���Imޝ�Iɟ ����)�Gy��x���O���@1�����a$I0�F��O�mZ_�8o�I*�M�1f��%bŢ�DH=aо1"���ob�6�dӞTc��q���&r���d韠1B-O��G��1�h���c<\x 4O���?����?���?����	ʾt]6�5 �<+�d	��o�b����������?i�O�R�h�󎄣c^QjFFV-�FY`��Zyz�0n�;�M�%�x�O���O��-���i�D;� 9�B+�6r�t1YV�[�@��Đ.�Hyk�bU$�OD˓�?!��
����*g���1F� ����?	���?�+O�oZ(z�J	��ܟ��	6�����':���Ƌ��?��R����47,�Vh&����k3�C�E���£.E\/��O���	_	��e$�<��'m!^���?񥣕�Z��� P�4�8�rw���?����?���?���	�ORc�ְ@� J�F�'L��ł�F�O��oڣS5ބ����P��4���y�A�3{�xU���etv�9����yr�w�Xnڏ�MC�jA�M��'Q�'��CB �S1{�n@3!�,-P�*Wf�6D�}9��|BV��S�����П��	���
7�� )�d�[�&[� � �%�~y��z��4A�O��$�O��?�붨��H��'o]�_$.�������D�����4\���O2� hŞ=����Y��0�, ��t��"�D~�&|+H���	��'*�ɤgA�a"�͓�$8<��U�s"�����0����i>��'�7�S0 ��K��F���ŏ��:��%_n������?A�^���4��Veu��d�S��z�Q5�t�Dy������6M-?9�m05���i'�����C��q��0��Y�h{����c�L��ßx��ӟ��ݟ��2ģB2fG�� -Z��x�!DH��?i��?!��iH�x�cX��޴��IC��ç�M(;�c��I�����x�`z���n�?!�Ӧ�Γ�?�4D�=9��4@J�[84@a-��E����O�T@H>�(O��O��D�O��is�C�}�4�8��^�(zp�a�-�Op�D�<ǵi-��1��'���'�哊,��`�Κ�Tl����&���}��	��MS��i>O�i�b)�(H����T�̐L֭�+�4���+��L�	�?	i'�'�8�%�T�o����i(�D�IwP��A�ܟ���ϟ��	Οb>��'6�,��0���I)t5|����[���!�j�O��I��u�?�1^�0�4_�|�ƈ��]m�}�*��.Tb�i�7�J�	w�7Ml���I6GG�r��O��S�? 6��QIߨD#�[
��x���x�>O�˓�?	��?1���?�����)ͥzY{O^���Q�C�]0�b�nZ�x����I�����Z�s�H������d�J�p��/��%��Y3#ݱ}O�Fu�0�'�b>�h��Z���ΓY�.iP߀F d��8g�6�5�Q��Ol�{N>)O�I�Oܑ���i���H����M͠Y$�O<���O��$�<1F�i�^�H�'���',�qq�h,<��1���Y�)���čp}r)l�|�IU�	�2��|4�,#�Ǆ�rr�XJ2
{����&"@L��V&�$�b��'��D/�۟����'��QµJ�v"���)�t�|�d�'���'���'��>e�ɄU�v�9��0�8���&(�a����M�_�?��7��6�4��ŀS�P��Y��3X����0O��o��MsԼi�b�1�ie�d�O~5��e��J��B?m�p�W�I��p�$�V�"�Ot��?1��?!��?�dr�lۄ�X7x�)�)N�c��,OP�lZ�	wx�'�����'A�yz ��a���1`�E>#�`!�c�>1Եi�X�.�4�T�)⟈9;F���6�;���&� }#@B�*vD�'h�<���y��ğ ����P,0��*�* j��ԡ�����'Rb�'�����$V�0{�47�D�1�:*0`��ǥ}��Ike�V�uX��ޛ���syr�'t��g�r	xq�A� 
��Ş�wH������6-l�X�I4sP���O����;�츋D�ǹi�89�i�r���?���?����?����Oh4�*��̪G�V�b�k?ZP]�V������M�aRh�d,g�ȓO2��(�{qz�b��
6�`��u.Rn�I�����?�Z��@��Y��?Ѵ�] u�Y
��&,8֜�aŶ��B.��?Iǁ)��<ͧ�?��?�&(K�P���S���8%@v�J�:�?9���$N���*U����IП��O+��x���	L�<�/��
ri��Ob4�'�"�i�ȓO���O)*�Xt"-g����v�ƩQ9��8��ҫE"4�Wo�����$HP���OZ�2��ƹI9�`�
�f�5J�O�)n�/k�2A $�O�k^��+�)�Dxh8�f�ğ��	��Mˉ���>qw�i�������sȮ�!�`ч{V�
��n�DtnZ���4o��<	��4�(�[7�� ��(O���e#�!p�Y�]B��Pq:O�ʓ��=1r��Z�SSB�*X0]1T"�=�V��cib�'��i�ͦ��4~�"18��߽gh���ɻ\�|���4vƛV�?�4������}K��eӮ�ɑw��d;�ဗO�^�(���'��ɷ��D�'�n'���'�前p
pU�B�, ǚa�ǋȉ0D���	�	���֟���Ο R')��<� 
����x��A�Ŗc�����MC�i��OEࣄ��f+���� 	:��!ez���	&�P���Ù]t�'����ҟHѕ�'�l����@\<R��C~VU��'�-��DJ9xaLQ'O�V}2��'�6-%fk����O9oZE�Ӽ3,�"8�.,j���C�|MYt��<���?i��if�r��i��e>��7E����Ռa ��zeǙ!k�(h��h�Q�'��	ԟ��I˟ ������	�	-�L��K�	i�ذeS�q�"<�'�7�X+�����O0���Z���ykw��++d�)2�fܾWw��+�as}��'R�?�4���d����ڑ�\�ر
�EQ�xRp��`I�>H|酘�� ��A�kx�Q{��Wy���*��;�.�%�����!22�'�r�'D�O���/�MCB
��?�a���qɌ)��ґ�`��pD3�?���i��O�%�'Y$7��џ�ozᦩ u8� �+07���6��[�f�nZ�<��k�������p�+O��)��U��/M���� ��[5r+�LV;O����O���OR�D�O��?������a~Y�C�K(d�$0�&�Ο��Iן���4jk���'�?����'�p�+��,�A�Wh�y�Ļ�`����MKe�iH��A�g���5O��Ā@iX�U�B>[1��ʶg�"Ee��F� �?�#5�Ĥ<A���?9��?�Tl���AA3Iɗ9��CcP�?����$�¦�q�g�Ɵ��˟ԕO���$rg��W)�7Vv�!�O4L�'�D�V���$��S�?��T�?V8����Dݰ(Ej�SrB��L��2�*س?C-�'<�d��$$�|Be�Nm|��Q� �1p��Ä)
�f2�'���'��O��A �O@�	��M#v��*3�<��e��q�ce�M �����?�¾i}�'�̽>�ôi�=� ӄ{iےdl�*H�'Jqӌdn��Zm$���y��'2�h��?���Y��1%���Vu�s�k�1x&�}�H�'o2�'7��'��'F�ӛu�����0V ��Ь���ݨ�4�0.O���-���Oz�lz޽A�"x@� �["ٙTً�M�S�'���T�O����۹qߛ:O��U��d��#.��w��kE;O�]�G��?qG!�$�<Y��?��K 	{�E3�mJ<\����e]��?��?a����OѦ��a�kyB�'w>`���_$v�S')X
.Și���]}�"�$uo�&��RP�QK�>�:�:Q�_��0�'{Ή��,�&r()���d��&q�T���n<�:e�1斞T����m���=�Iß������ş�2�	�I�4�'�g��'6	�u��a< ����'�6�����O���O���O�EnZ�|| ����%������WtZu��n�� �4S��u����LbӾ����`��u�����?ۀ �e�J�K�<��	ϽD�����#4�D�<���?����?����?�TkԖ#V�;Feطn��q	���ڦ�bs�͟D�	ӟ�rPᆋ;�Č�v#E5VS��&�G�9��%�Mc'�'�����O��4�:���\�m��(f*F2�����*ؚ4�	���R���K��'�zmә'�Z�M��*�=3�0sѩ�5�ؼi C �?	��?���?�'�������.�͟���j��Hb��-I�y�Yy��|�OO剰�M�µio�6��)k�r�ʇ@Q��JXj@�$rf�1��f����ݟԁ���4Q�ju�e�ry"�O���Q�z��|)@σ ��ї톚�y�'���'�b�'���)�r���2t��0�BA��]*�����O��D��qr'�z>}�I �M�O>A��T�UkR
R�m�h�Q���0d:�'��7���m��V��o�<Q�e;8�(�ʔ$g��th��ͩ�B��� �6�X�DJ�䓷��O$���O��$A�*p��A��(�h�Q/��|yx�d�O�˓4x���؉"�'�S>-��̪ev\`ZEP��Q�3�:?)�_���im�r�|�L�`}�:���_Ԕ=Ô�
�,���f�J8lz�/O�IZ�?�Q�7�ā<K�ݘ�Þ�c���p��Pz(��O��d�O���ɨ<�¼i�\}��^����*R**К0�р}�剷�Mӎ2*�<Y�4R�	X� �1!�ֹ�v�ЍY�<��i#6� M��6�+?1�`±-����1�$#�:Q&�Q���>q Z�b�g��yRP����ٟX��ǟ0��Ο`�OiPx�g�@�\�$���E�3~rX �b�$�ȆK�O����O���d�ʦ�ݲ>Y�f�W�2||���_2!;��A�4;қ��,��	�2��6�u�Py���H�(���hS}N�Iӧv�$�4��BD�t�I_y�OH��9��S���J�����ҌR�"�'"�'�剪�M+hL��?����?�jÀcP��5H[�W$�+g��#��'���3Q�&@p�2T%��I�@�$�ҸY�#���jհf�.?Y��T"^Zrcd��G�'RY|�Đ��?£�%]��u�-:@M$RD,t�������8��Y�OA2@�":�R���#>�A��gd�@��Ǵ<��iz�O��;
y	a"^uʦy�B%B��צE`۴m��V�S�9,�&��x�ļK���g�-A�]HF'y9jA��D)tD�$�T���Ϙ'�b(���#&5��H2ݮ6�|j�O��o�.m0��������IO�'��}���nP���
�mZ�Yc_���	Ο�`K<�'�?�'e��$aˬX�>T�FY�d/���MӖ_�,{qd@�9��6���<�Q�27����,�u�Kk��?a���?a��?ͧ���Ҧуb,G̟tӣ��W���"&'^QojQC�`r����4��'\�6��F�qӪ��I�$��ѐ�*�_ڄ�G߆TRq���bӆ��Q�P#�z�JN~"��FO�h�R/u@�!���&����?��?����?1���O�P�ڷ�ڂt�.]-�%8ҕQG�'B�'��7m�6w���OJn��'Ŭ�(шO�	�̱ ��]�9T`�*w�*��O����0is�y���	�|�����B�Àb�r����5��&_^ڝp�O��OF��?���?��	�X؆�B�A��hĎIl҉����?I(O�Im��..(�'�Y>�p�ᙈc�^`Pg�	��\X���:?)�_�X�ٴ3훦�8�?EXQ�ܸ
ߊ}ʕ���O#�0@���z��V�\v:�������ɟ���|b��,ek�xȱD���,�'�¢_�B�'_��'���dZ��K�4!8�(CX�UX��N>z��2��β�������?�^����4p�,\�]�Q�*o�	�Pk��V�y�6�ZP�s�V�	�n\9�柒	�*O��-Շ6;<�s`��+��52OZ��?���?���?)����jGv���.M��؃�O��e`�f0�N�O����O쒟�d����ݿ0`(���"0�Q@�
d���)�404�h"��F���7f���b���q�B��*���b�Ol�����-�"˚|�Py2�'�r�G�5�T����tS�PQvDҎW�2�'�b�'Z�ɒ�M3�,��?����?�� �7���0��9:��z�i���'��������H<�gJ�0	��P���9VҺY�ȏi~҆�s��D%Q�g��O����g�b�Ǹ*����b	
lM�5K�kya��?����?���h���D��`�� '����6i���$�ɦ�8���П\��!�M���w��p���4
��` V�1���(�'L�7M�ߦj�4]�D��ٴ��$PcL���'NP��Ҟ)�N=��*��y���u�,��<!����ې慗sB�U����)D�Iу��Z�4���[��?���O��y+O(,8��ô+1iu`�<����M�3�|J~�d�X�`n١��@n�r�e	�L	>)*@ �����!i|5���[j�Ot����bĈ&6���@�G������?����?���|�,O��oZ9?����+pr�H�fBb��x�RD/J��	9�M�����>�i��6�����X�g�q/n0Zp��'���,��<�0K�7�+?������	���'��c��O�q8&�ѓHP�q��;1�D�<��� Ū�$N+fl���1�N�_1�h����?��5]��HF���)�ߦ�%����D��b0����R�nX��e ��W��f�~��iO�b5�7�)?!0/
I�? ���B��A���SAJ6d! �
�DL
�?a��"�Ĭ<����?q���?b*�:Zat��ˁ��|�����?	����զ�8�C���	̟��O��q�e.�5�4|��,��Q�jX��O:!�'�b6���SH<�O�H쒲����eJc�(u���ҏ)�0��"��% v�i>����'� �$�,���އU��
t"]w��L�VJ>�LzشK��Ȕ�߮�Ӂ���-:%�ۛ�?�����dOG}r`� #�	��� F�۴P��q��)�4pB�!��4���ɀ	رH�'WTʓ��Ź�.����3��:-i~������O��$�O4���O���|�$� �J8��k�mP8.2ε��g\�uN��'����'��6=�r�5&Y����a��Q�ܙ�$�Φ%ܴ,v���d�O�t�Ȝ~��f2O�$[��
 ^�hQ�������D9O� :��Յ�?��	1���<ͧ�?�-B��(�%�G�(����%f��?����?�����ɦ�RYޟ��ߟ�1��ݿ� d��Ŋ,�TZrO�[�tY�ɗ�M�'�iXO.d�%���a��Q�gE.HJ��+22O0��55f�9�3غ'J�	�?�k@�'E�X��p�� y��Q�f�Z�;�v	�V�'~2�'���'�>��	�)���T����5�KJ�u�X�ʵ�'L7Ml-����?i�i�O�Λ�{�����Di;�n������%1ش|؛���}_�6?O���6n�5b��~����a�`��L��H>=�$����(�d�<�'�?���?9���?���G�K�z�CϨ����3�����ř��ȟ�	矨%?�	�Q�2�3feǫ�4����W�^@LU��O=lZ�M�x����ՠF�!:�D��$U���� A���5�-������h�DN��O�� ��I���ƭrY4�+s�E�G�l�R��?����?���|�/O.�m�n�N�ɘX�ؤ;gHY97C�up��˥0�b��ɧ�M#�"�>�Ǵiw�6-���X� �f�hRv�ܲ��lb!�W�+�Lm�M~�E^,9�[�'���f� i���L@4G���GL�<Y���?����?1��?A���#��83�7-�<�k�!�.>"�'X�	d�4�j�5�`�ąئa&���%�5w3���E	�d�C�I?���?���|"v@Z��M�O�yC��]���A�$N�l��%���̱��m��-@��O���|����?�t�.xh��U$]
�f�ׁh�|03���?�,O�n��i�>D�I�<��u�D�6�L}P�%�*}߮��Zg���k�Iҟ�	���S���	1���!r�ñu+� ��E�b���Cѹ-қ&h�<�'4����J�	mv���B��D ��6̎�%ˈ��	ڟ������)�Sy�|���!�>u�\� ��BF�왗䋶^C����O(Xo�Q��4����Q^X=	I�V�m��A��֟ �ݴ ����ٴ�y20�b�Y�Ev�)O�N��iQ�kȑCB��
AթeB�<����?a��?y��?1,����B�ߗJnn�	@䆣p%d�j��@զh���̟���ϟl%?��ɓ�MϻWC�����0	YR��N&jez��?�x�O���O���ɱ�i���&Sf�����=�`�J�[��$� Oo@��'��'�䟨��:;8�ਰM��,c\��l��*dz��ȟ��Iܟ\�'zV6��t/��D�O��(�e�f�		D���wiʨ�d⟸��O����O��'�@ːH�� 0����?"2� c�@c���	�XY����Ҧ��,O����(�~�'q���6nQ�m�<�aW�ېE4�`�'���'v"�'B�>��ɽJ٪1H�e@�c�� �"���ɗ�Md��?A�E��F�4�^EQ�	m�H��4�
�O�v A�>O��l��M��i�Tٵ�i��	�`>� �O,j%�AC�(h��-�<[�`H|!'�̔'�r�'Ob�'���'�H���J�hm`��ql�6Z��}�uZ��pش3�������?Q����<a�ԁ,�0�H�B�f᳥�ڡhk����M+�i�rO1�z�ʶ�� *g�ugF\ 	�~��L���|��@�<���C3t.r���������
�1Ƅ��+S��@X��
A����Or�$�O��4��ʓ.�D٩vT�@�ؤ\�$�A�2���§_�%
�
h�t�L��O��o��M�i) =Y��Ag��R�nY�'z���d��Y�v���yR-�BG�d��S�߭C瀤v$�X�6�?I�|�A� q�L��ҟ���ܟ����@�z�C�"C`bԺ����-�q���?��?�ӻi8�Ms�\���޴��(��=#�� �c�̓")��A��x�n{�d�	��$a��?�����X���-R�B�k�A4`�x�äf�(xj���'�@&���'�"�'��'����`G_��h�ei��&|�}���'gB[����4<�&} ���?�������&��AQ��0rӺ�#uM\}�	 ��D�Ѧy�ܴbS����?Uc� ��L]�6uZR��
5��ڴv�,�%�C[y�O_�1�I,�'/��$�� +#�ɠc�$5�����'4�'2�O(���?q��Ɍ8�|�1��A H���G�
h����ݟ��4��'� �U,�(\(b�&��p�� Æi�g�	�x �7�� �"�Ħ}�'� ��?U�gX�$h��	Go
�I8�A��I{���'8"�'+"�'���'�哝f:&��V�$8Ֆ��b�
y����4H5 }����?�����?)r��y���=�N}�vD�>`�$���F�>_h�7��=�N<�|±
��M���� )q�L�%�i�U��P}��5O¤�V"��?mm8���<��?A7/V
WР���D�A�UH��ب�?����?��������K%��䟨��🰘q�5LQ �)�.�&W"��Z�f�I�a�	�Mv�i�ZO��2���S:��@׈�)��LSÞ�Tq�Q3	��U�V�B�5���Pҟl�f�=А-��"N����h�N͟ �I���	��<E���'���Y�'�,��,{�'.���R$�'-�7-� n��$�O]mZH�Ӽ�"�M-��q��"�k1�U[����<���?��i�d��i���5���k4ٟ�A���6M#�eP�m��uӴ��"�ģ<����?Q��?I���?q��V��" Aн{P�|�˖��˦}C������	�$?����9fH1ƀ#���@eғo�L	�O��$�O��'��ޟp��di̅覃��lю��'c�i�
my����Ւ,O�H�V���~��|"T��������yC�b�%ee�����������۟�Ty2�~��Ԓ�i�Ov�Z2�=ڤ�FK��*P(�O�am�U��IJ�	��8���M����0��xC,��XG�Z?�P���4�y��'��I
��Yi:)Op����$����U�`M���Y	c��i�1O����O6���O���O��?���H�$��P�gG��}�� ������	��L)޴��'�?IU�iR�'�R���E)CW�	8� �Cº@˳	5���O��4�$��kxӜ�M�X�`#��G�A�w,Uy�!����;Q���n�I]y��'���'`BgʐU��䄏u�����X�'e�I�McĈ��?��?�)���e'ju��BG#ҵ*��<�N���-O��DgӢY$���򟖵�m�.CT\��
�')����Q+Iۤ�T#������?	��'4��%��R�����3G�TC�(�q�Z������ ��ٟb>��'��6Z���X�'#�2> ���C̗�z�����<1G�ik|�ɼ>���,0�� ���!bF���&Q��z(b��r�V�D�+��6O2�d�s��Y0�'F	�	�&���8dݢC,,C��Jc���Ny��'RR�'-b�'��V>�T�GK,�u�geK�*�m�f��M�dE2�?���?)J~��3ϛ�w����	��p�����,܉w����'�(=�4������ps
nӸ�ɀ*�܉�砊�8�\VRrF>A�'��y��gN�  w�|�W��џ\@�O���� 1���$*B��<�I��$��}yrt��aV��O����O6�[#P�T������J�@ᔯ#���O�T�'�6mɟ�&��{qcD�X)#��PP�I��he�T�I5"$a�o�"����'������0�'
�)�	�/� ���Z�����'��'3b�'�O4B�A�3�-�0[ι��h;B���0��D�r {��AQW��O�D�$� �i�ɩSI�,����PMG
t��k����Mð�iF�R��i���Ol�S�J>���营)"P�!��/i���#��f4��O�˓�?����?���?���Q���� ѕ��)�/ ��,O� nZ	���	����@�s�P���ARt�@.C�B������R����ǦU	ܴT񉧘O�
D96�l���P�,˿k�a��C%�D�e]�����նdZ�!�e��wy̈́�q��<���6�Bm*�.��A�2�'	�'��O��	��M��j���?�e%9b.��J���,������<�ųi��O���'�^6m����ڴeC�|��=+g��8�KԒ���Q����M�'&��0Վ��8z�	�?5���n"4%B�M��H +�K�:@���	����`�	�����Y��I�i;��ݽ8=�!����������?���?c�&�	��	��M�K>��AH>H0-cC*��c�RLrFf��H�''�7F٦]�8	���o��<q��J�����2�R�w�I�V% ��E
��!�����OF���O��Sq�*���!�B9.�)%FE%)����Oh�9��Aʯ�e�i���',�:�;S�	�A�
m�6&� in�@��� �Mcg�i��O�i���]�K<FD ˷"r6Z&�u N����Gm(�����O��J>'�A%d�T-�4�*�����?���?a���?�|�*Ovqo�:zP+�D&K�,)Bo�s0�i�3�^�>?2�'�B6m'�	���dJ��a��H�!]����� ~�-W�W��M���ib~�kQ�i���O�0'5����<���VX�l�R�Qk�Z}Y�	��<�-O��$�O����O>���O��'c�`@�2�߈�` Z�,t� q�ԼiR�a��'-2�'��O/R)w����4@{"3�Ŕ0%S�����}�]oZ��Ms�x�O��D�O'ډ�i�3h/��6G�)L\5�v�	t�d؍s ���k'��O˓�?��'�Fl�ӹ+À�P0d\�d"|\q��?����?,Otxm�/�\��	��	&�tq�sB&<52�GH_"`���?�']��۴<z�֠?��*k�L����\"�)��/2%�d�Oju�%��.v��Zä�<��'�����?qq��r�a2U�?��Pe���?!���?y���?���9�}*���+a�|%y��u�~��O�EnڡT*��'�7��O�O�N�$"xa�	́&� +�48�Dk�vlڿ�M��߃�Mc�'h�:Yw���ӑ��Uh ��}j$��Bf^'K���I��|V���I��IܟX�I����/J�EW�����3����CKy�e�Lh�OV�D�O���R��$kR2� ΋�\�F�� mY ��>�i�7-LZ�)��?��� ���q��?\d\�BG�ZН2c��)� ˓v��7��ObxN>�/O "�1F�DuM��̤#��O����O��O�I�<�&�i�l����'�P�)E'ےFA|II�{�Q0�'�7M�O��O�d�'ir�'�T7mɕ�n��l�u'�X��K�2�Di�`lc�P�	ԟ�UCҗ*<��%8?9����c"ΎS
RL a�I�DM~�B��@�<9��?)��?���?A��ġ�7MЂcV�>uD  K��@oB�'���e�t�c�=�����q$�8�$-Y'�TF�q6N��#���ᛖLg��	P1eqD7�%?I2�E2'�Z��1B�`���+f\�R��O>�L>�*O�$�OX���O��%/�!n�6\�ǃĖP�P���m�O��$�<�3�iÆ��g�'%��'+�Ud�iNЕ�\�K5e��)������MS��iFO�I�\��[�Kߴ�Z5g�H��P�&Ƶ|�JQ���/R�˓�i�OViPL>���=�ڍiE�&7��=6gΑ�?���?���?�|�+O��l�8�V\#�,ߗ&&.�
c!Z�ΤrA���t�ɲ�M��b+�>��fe������V�P�:0	G,�O��m�Iz^!m��<i�O~69y@��?U�'�z��5�F#\D=Ƞ�F@��;�i
�j�@d� �ׄ�Ȝ��&�e���G�C)t��!�Zx��k�~i��H!GȞԅK�\z��V,��C*NB�m��b��ç<��6V�E'�1���)\� *3�)cG8�9�@�	Jdl"�ƭ(7t!R�Q�Y��q`ń�HV�(��
o���.��'���C�85�)I0G�;j��y3���d��h� ��G��g-%�Kᤚm@�JS+��� �A�59v�b�ˮ=�`=�ٴ�?���?���<�Igy�)��zJv�2SO����q�zm>7-_�/p�$����:;`M�઄� <��g�5#����i,2�'�bQ9X
f�����OR�	l\mA�!�e¹�0,�}d6�<���1��$>U��˟��IW�X�'>�]��[�kXl�۴�?����o9��Wy��'�ɧ5&&BH��ؓ%�
��8�c��	�t\��O��O��<� ;޽(��.8�4q�-�#x�ʥq�S�ԕ'qҞ|��'pb�ˬ\*�`ŌQ�X�!U?}�8H��|��'<"�'��I�]���+�O��q�b�&:Xx�	�i��L8�޴���Ov�O2�$�Op��d��d8�CNM�d1����%n,��d�>����?�����lp���OH�CN'O�� #6�^$������z[6��O`�O����OB!U�$�I�u!��;��Vta���W��7��O��$�<i厒�dM�Sǟ`�I�?p�.Ŋ'/6H���*c޶@���	�ē�?���������䓒����-w�t��g�(c��@�eϔ��M�-OdQ�Ĥ��Y��쟼���?���Ok,R"��AiツBΔPZ���%�6�'l�NѪS.2�|rX>�L>��!�D8�J!����b��mڃ_,��Sش�?���?y��	�	Uy�U�xœ�Bۍh/T����J#6�t6m�.�R�<����*qٰoT�x�,e�PGٮ}Nv�ۃ�i R�'����s����D�O ���V$& ���	R��z%��*T��b�`:"/�a�؟��	󟔘`$S�Ϝ�aE�5A���� �Mc��k���PQ��'V�|Zc�X�2AK�N�>�ڗ/�5_Z�;�Ov����4���O��D�O��;H>�4�8U�P0jL+,�8�D;$��	jy2�'k�'Y"�'� <c��/a?�hJ!�ק�������=��'���'��S����G�(��􊗟1���R��	� 5&\XŠ"�M�+O��&���O ��
����an�k�
�-���*�����l��?����?Q,O�R�EBz���'o���N�'H�^�be�܁zg^A��x����>�d�O���;4��OZ���F�/?�D.� J���0#�i��'���.���KK|������`Ӑ�;Cl�%�F�"��$�(�'Tn�F�'��O���W��ܫP��S�i"g�A���	ş�K'lS��d�Iǟ`���?q��u��՗r�ڤA��\�y���M���?92���0�&��<�~:�n��vB�[��8Q`�l��,VԦ-�#nH��Iݟ����?���I��}��X4����(E�a���l��J��)+��=�)§�?�`�W�?9~H��ȝZ�2隵�U6���'�B�'��|�!�&�4���$��L��?^n�1�2OT#�T�{�Ge�J��-�ĊJ��O�D��$`Qߤf�H�R7j_�q,�A*x����طX�D�_���a�2��y�q��>m:�A9DVly��x��]���'\BU�8�	F8�f��C�|px��u���� �`yb�'��$�OP��je�L��gڰF��B��0+��t�4ybs��l����@�	_y�Y1VJ�?=�Չ���=k5l����-@\���?����?�*O���|���|�!s*X���rQ�ڋt0SV���	ğ��'eN�[/����9�#��O\fH;$d����gnV�M��B�'r�I�tvOR��u�8��(r��_��~�7�i���'�剬5(�|!�����Ot���)O���"s��#� ����>T���'�'q��R3�y��'�I~�EU5�:qz���^����c/����'$��
��u��d�O8��埊�֧u�,	)yR4���,Ӯ �HS��)�M+��?����<!����7�*{��{c���Z�X0��듋2�p7��sn��l����I��0�S���ķ<iu� �ܣ%��6���Y��B���d�i����'��'��J�d��[&i���B:p���3HɡW���o��|��ҟ��J&���<���~2'�57{�MZ�K.
1FԂu���M����$C3*��?�I��h��
�<L	V�G4�����j�-4�n�m�ǟ�H4@�+���<������Ok,ȊINH�)�Dqs�i�Y��2W�8�	۟����X��˟��'��,+5�Yz�D�2�_3:h[�(�2R������O�˓�?����?Y�#Ǎ- ta)K
�
4r�@��c�͓�?9���?a��?!.O�L����|ʲ��4T)r"I.E�Hp� W¦Օ'(rS���I៤�I���i �0I�Fs}�ej��|�NPش�?���?����$P�:�R��OZcO�(���
�p�LD�G,�s�Bpش�?�.OJ���O��Ĕ���O>�$̤HnF���㌂�<L��a] i.��o�����GybOD�7K��'�?Q����&��J�H}����fŮ���@!
����0�I�4���i���O-rџ(�Ȣ�N�^ZE�לEm ӾiX�>v��,q۴�?����?���Ym�i��%�C9U�:	�7�Q�d���1e!y�f���O����8O$$��y��I�i�P���7T�8��#�D:���J�j��6��O����O��I�W}BW��H�ϔ,=&��f���EA������M���Y�'a����8��-�"�8z�dԫn�do���$�Iݟ����%��$�<Q���~�E�V2��˕��>'��]���¦�M����$U�?������V4l@Ǆ�o��BKA�@�4�?!sh�7	B��LyR�'�̟�
?���*�0�
"䀊X�2�bA��?)��?����?)*O��p�fL+�P,��K,O.ꔐp��7k6��'T�	�� �'UB�'�P_��]�
�t%N�0� Z�f�q�'�B�'wB�'��Z��h����t����81�jJ�D
( �-݀�M#-Ox�$�<)���?���.��MΓS9��I�Ƈ7�ib���+݆4��R�T����P�	yr�ϢM���?AI؈C5�e��*ޓ)$�����[�f�'�����������@E�b��OH�Z��Z{_�9� a�+/$4���i=B�'��a�b�㪟6���O�i�w�%i� �A�dءk��U�Q�'�2�'JB�_�y��'���uRS��qe�?q!�Y��
�q�'FL���r�,���O���韆Y֧u�)�b���T-ȗv�2�KE��%�M���?���<����?i���OA��Sů�9�P���#M�C)�0Z�4X����i|R�'���O��ꓮ�$��31D�׍�&�0�!o iz�	o��a�H��F�Ih�'�?i����c� :��B�ao��3K۫Uϛ&�'�"�'r�ms5��>9.O&������n/9�Tͣ1#)2���>.O\x������I���ۗB.�,m�g`�Ur-rf�)�M���I�(1�R���'�RY���i��c�c��D��0�#<�P��&`�b��ޚ*g���O����O����O�˓+[n�0���d��8�>���#��O���{yB�'������Iş�(7
գ`�M٦���c,Ԑk���/��Iԟ��I��,����@�'���+��k>��  V�UC`De��HJ�`g�Pʓ�?�.OR���O��DG�\��$�5̞-�ƛ�XKV����
�AjD�'Tb�'nrP�$�Jɐ��'g����t)�U����t��3!�n��W�i��[�������ɫV),e�	P�d sdH5��r��u�ǧ&�f�'�B^�D@�"���ħ�?I�'{d����͕3r>t�""M��ic��ŜxR�'�������Oj�ӵX���h���7��g��bu�7��<Q���"��v��~��������@�iJ9�
���[L��Z%br�>�D�ObYR�O�OJ�O��>)n#��U���g͠}��эtӪ���Iğd�I�?�L<���Xċ�� b����H%E���"��iyh��V�'U�'p���B�(���2u�=ȃ� 	���mZ�$�	�s& ���'���O$h��˟22J�� BO�#�J���i�'��5)�):�	�OH��O&�R'�O"N�|+��\=��brk����	�HU�}Ћ}��'ɧ5���;sR�$�p-&i�d�"����'=�2�O���O��d�<y�A�v��IɆ��\ڶ�_�91�V�x��'|��'��
�
��6cN�`/Ph`я0e�h#�'5������	�Д'�Y֧a>Ɂ6��8e�^�'���l���>�d�O��O��D�O�@{4*���9.ҽl4��{�Ag��3�G�>���?y����4��'>���B���t!%m�$%2W�Q��M����?��-Ǧب����F�J|�r@�w�n�1����3�.7��OL���<��&^#=&�O]��O�JTR�/9:����f�y&<�%	%���O��dP�0���9�d�?��I[���Qcm�6 �,��d`� �x˸�!�iV�'�?��'g��>���&���uv�<�Α0��7��O����7����5��.���������V,���iL+L/�7A]��oٟh��˟ �ӎ��'�ܔ�5*Q�9�v�{ƅ;TbH� �xӎ骵��OȒOD�?��	�D,��@�#�_��D�3㇠/��@�4�?����?Q�B��g�'���'��䕣B:��iE(̃:6�Y�J�f�|��M���|��Of����s@���Q�s�҉�4�ߍ}��UlZȟ0��W���'e�|Z� l���mI(FB���GC C^9`�P�lb�'�؟X�����'Z�J6��
 �ذ�D�%��8Fܑd{\O���4��?i�}~��we�)�a÷��0Zk�Q���?���?I���?�.Op��6��|"�'�:?�P�cF�h�s�MZ}��'rў��I$A���I�u��M��	�4'�:P�a�3G���O��ON�d�O$�Dۛj�'�?���	�,���.Q��0�SƐ�?����'��'~��'x2�}b͎6Y���O��u*�M����-_��Z����h���M�^���i�L�Vͪ��p+*�!�W�&�e)PgI&Q��4`����5n~�� b]�TzŬN��9��gU<����J�AತH�h��!F.U�����(.���
^�y�Tݣ�2V��+�Eү��9���&l�Vx�����F��S�U��b��8B �k �q>��"ǖ��rF�ż|�K3��
�1)R��/^�z���O��$�OD���O੭�w�&d��Ǜ��0�&*^�Y�]
�iO~9+�ӷT���Ѧm�-��O�<�'��,{m�Ai�`3�CՀ)�y[���:1�j�t 6a9*	����ոO��������o�$At�`�`dҢt#�p�3ϑ柀�'�@����|���DT.0a�;j��w���=�!�D�>'g
�Q��υ4�j<�P�E.m�� �HO��OhʓJL�q�펠Z��b��Ѻr�V@�#LF�I�	*���?���?���h���O�瓤.��� i^�
(�8�@m��B�D����7<�8=�&��:�Z�)��'�.���h�g$ϟ��8a��
����C'*Xx"��V8��@��`�(q��v�Zm�Ď�3B����O�=a���M�T�؄`�5q��8I��׉�0>�N>�.:r�&	(��Er�i�"J̓���'�IZEP`X���Ā"xI���1�K�4�#���>:�N���O:�Ci�O���h>��r�����I"s�B�
�R�o"�j�pա�1���K0D/n�z��ğ�H(�3�͘O�du�efd�t���B�&;���VE�8I�桋�D#_M깻��I:
����O�˓N:�܁�<�%�]�'$t����2��P���T��w5[B��hb\e��N2�hO��Jߦ�$��4lP���o؜�(UmX��?i-Od���
Ԧ���O�U� �'Ǣ�т`�V8���D����v�'h"aO�WH>aK���H�~)ԧ�ɲ|.���)u��wnfИ�ϡorX�'����t�����=�M��i��1�����&\�p�Oa�q�'���S��Y��+��a��E,�l��,"D�h����(��DP��7m~��b:OR�FzbN	a�`�#d[�6���Pb��5�7��O����OR)#�Ʌg���d�O��$�O�NقI$<�G�I��xb��
p�HWI�?V���SB����G���O|@�'&���׏5�txg!�m
���d$[���Y���A��JB@�O��',�@�*G�>���f�dY��'��	�36^�4�N�=�� X	d����"�+���w�<�H/<Z 	I���� ���<I�;�����Ο�'���aO�.��9�$�=}�
p�WBߚ",.m���'b�'5Bo�~�����J�	^���qb *�0�`Ňel�AQ��$'��ó�0=A��O!��\�D	�`a�y����T��@���
w��� 7#��fH��ǽ7�J�<qé,n,��Dk�x�0�F�ilv��I��,�	Ο��'�b��-u��� �s}�X
�BP,g,a|b�|��H|���i�"Z2@������R.Ø'\7��O8ʓ,м(z"�if��'�8��š� ��  h��m@B�'�N�����'��I ��(!"�"�$�	o�R4��I���EQ���gE�x��<3��`Ç�ȝ[B��W�ײmf�}�[U�z0�D(�h "�V@�'#jY����w`�qB�؜��s���7\�8]��im�ȑ�Ki1Xy�GD�> +��������N����Gۼ>0�|	��O�cA�b� ��k�#�Ms��?�.��Ta��O:1Æ�E� �c����e`Q �O���˰	���`k�L���A�ʟ�'��i(y�f�`�^5Ucv���P	7��K�hK�/Һ!N(�3vI]�H�2��c
�:l��.t�Rȑ��>@U��Il�H�Ӳ)�X���׺[��("^�F�tc�0��`x�h�@�q��� Ü2���ё�!O@uDz��A37VQ�d���r�U���%�6�O�d�O
�f�1n�d�O����O�C6g	>����Gd���VH��]*����2��$��{li;��|RG&k~�H�! i���(غ<`� Q}�%ķd��}&��k$O�3�0,h@�C�p{�Yp ���M�P�iB��h<��,O��d �l�R����_R�3�����	�'��`C��ջX���І�?OM�T��O�Fz2R>!�'֊�2�5
xT �;F�<(�	�'��V ��*�귀07�f�@	��� ���򈅘C�mjd.K,$��J"O�59�-˨� �f*�1.D|�"O���kÕY�a
�J]V{@"Of��@BQ�d�tQ2�'�C}���"O��jGR�6�\��am�*N_4��"OxQ��݊OC�(STnI�R�qY�"O����I�ԝ�㞷5.�(�"OT	����,�0�d@;<��aW"O�Rc�a�b@1a �e'ȼ�"OZ���B6N��C���W�M�2"OFU���1!v��`A�8	v,��"O�����A0���`�)>���#b"O(�y��Z /=||����#���z�"O���!�פv,͠`O�-o�i5"O��!T
J�Y�̤����Ga��3"O��+�kϛ����7yC��`"O���v��3m��|R�M��6���"O����mq� ˣ-�(�$���"OH��/�g��`)�#�|�!"O$ձL�.w�X�ꑃK�<��S"O�@��g�;qpdفvI?}��ԑW"O"8��#J�><y�ATu�R��"O�U���O��D �M&H�����"O���Q`�5E��R�._�r�LY��"O���bO�="�U[�M��� �"O���Ӥ��_��L�@)�k$@��"O`%BjO�f&Xt�`�K�d�z��'ML��@�޷V���Q�*�D�H��n��qq��-3��x�
�>��x���1Q��$#'!GIS����	�$��9R'�8""�$�6M�q�ӶWKZ`���Vh{� �b�E�-�B�ɬi�80z¨ܠ"�B����ȟ.� ̘���g�(�#�ly��ԉ˱ݮ@�t���ũ�<��c�P� �T�.S y5"��3G4GK�(��L��ȩ	�yڠ8X�N�$jJ
�!0ړX=fD��nJ�EE�k�!�!!6J(��I�i��w����*� F�Y�,w�սe���SQK�%k���5m�20WZ�Y£*�O�m��șcyp({��S�0��c�>Q�B�����&�M�� ;w$n~*�>e�Ӎ�&?+ҕi`��Iۮ���"OҹQ�V�n��P�C��*���-�;upl����K(���S�'L�TTB�k޵�R����<��L�a�:����6�T����z��� ��:�����+Q6�d�D'��3�L�]\���a��ў�I���#�*b�J�=-Lq��I9O��TD��j9��2�%N%��ac���O�b��K��ځ���)G��  jJ�����?X�p@��G$�.m�2��/F���D\��m��&��#.H���&��*Nl�BlO7(R��r�B�I)V
��
_�d�P�bF�\�T��`�@,/�dHR%��~2����4)���;n�H �_0=�����0W�̅�K�n��wd�R��u�U�� 
^��ucy��F�� )z��� ���(O��i`����4@2A*E&�Ls��'D�슣��y�R(0�n����52�Fðm8<�A'̗0�����o��p�4�ԎӣY��}��T��}YC�ʈ>����i� �
%ߕ1,���Wg��N����r��2�\Ǌ:�ԟ�a0��ϧ3�\-:�/!@�=;"�'�^EAEK	R~�,݂Hw:����S�;l�8Rꎌ	I�,�p��9x�>D�O<%>�S��X�{�&�b^ޡRU �D<�,�w�42K���A�!�?�#��M73�<��b�q� �.���WK،t��7p8r1��9A��=��R1��d�N�vFDB���j$0c�ȣ�6�L�TH��{��s�z기�PD(D0���M�<I��P���\��@ +9Y������a	����Z�#-�U���jj8Y�,xͬT;��K�~ �򩖳%���Ӕ>�O\�sunŞ��q�P��&1@��ד~T.4p%�>�#ٚ?��ԃ�@�[� 9[7팑.����W#YhAŦO�O7� p�f�9�yw��3Y�l���K1Y� <b��֓��'����(��|:�6�pӁ_7e,����Ψ1+T���N|�+g	��F�[��� [��G{�RC6�m�0�+���CBC�g�8�>�P�x>ٲ�	�0/|��)I��D��� �߆|*Cɑ>e�TL��Q�J�$1;�e؇r��I�}*�8�iϾo0<�֢�!��t�'��j�����	�+�*-�^�9���"a?}*�� ���"�/�r ��ϐ>4 �(�'�0�s$,}�ȖJ#f���gȕp�
�ȣi��elآ0jF)m��]C�@j?�}*�*��qʖ�	�C���
�` Fx��^:�8�(���ا�'od$h)��3(�Z�ztM�xҒI�BN��b��1���W$��N� �εa5��;!3ڱ8,�8r��I�}���]��獰�m��B�{���WJ�N��ւ�E�nUQ`	љ1�4�2��'��=ҧEƿR�0s#���w��}����!yRt��1eT�qC�k��s@�4]w������D���`݉{�A�w��>~��!jb�'��}94�>}R��;d� J����(	�A�9%��AЀ$��9o!��T>p��|"t���<�uD�i]F��3	ChA�՘ńEl�q=������IC�@��*D%t4\�TQ�(JX<�:�����J��	������UM~��! ~B�(��Iv�)�d�,��<iU`K�`lj P��9���1 ��}%�m{qT*O���A� 8�S
˖W@d���'x��QD�'c֌���״r���rC��19�h��Ol[��,�r)�dgܺQ����R��Op����,�$>��ؖ��\T�`�-�*k�!���=�^�*��B�&���HҌG<RTH��w�ŋ�,5k����&x(RDZɚ��C�zޙc�$� UP�Z���)U*6�4��a�,W�b�REB�Ԯz��:#�]�i�8�'���qN��rS�pJU�F�H�h�؉�"z����6(j)p����0<�G�ĵg�@�TC�;'���J��(�0�Q�,1(t�b�ēDK���� �<5Lb�VHG��=9�d���C��B'�iB��:�Z�N�рX/jt�A6om�C��2�韲����IR̪"D:ۺ�;s"O����J ��4bܡT��1��~������b�����g�m�!��ǒ+f�T�RM��lE)r�-$���퉡T�����b�m �d�%����4[@Y˔CZT�<3�b��R�V���t�I�BQ��f�x�@�6�����'���T.+#
X��X6?XB��Qx[b�9BN�.`?�j�/�10�ó-ֽcd$��' p<��	(DQ�CͥF�ّ@-�>tI<O�ݱ'�J�=h�y � �5!(¡����J<X?��0��D��9��̗�|J���Q� ��I#m��f�7pHt<���	^< 5��H l�x�L�����	��{�h���w�2\J��a��C�*|,(�x	�'�ڌk1,C�b��ȗ)��{d�Ia"�|�!��;��h#��ܚVC2�)r۬��D3��6�¬~�Ȥy��%4�zT�����y��tzU��	�R4.��S"I�]��AT �P:e�fD�V��ś�A>���C���$��#=��
	7qk��mނa�̥�i���!=̤�a�;5Z �"f]9y-&�֝�}�.�qr�Ðk2��φj�B�o�|��	Җ1E��3a=�A��+�@��%e	3�>q8N�X�O�O/4��w�0� .Ȋ"�إ @a��'rH��'�0�cV�5�谹�Ɩ���ٰ�>aw��a�.,+�i&2L
ѢI}�-�y�Џ��	Y�Q�`��b�牟I٨	S�h�;Nb��6I�d��yJ�F�1�,�R�M�u(��BR���@bp�gÂN����Fy��U�^(��r���jH֬�"��U��[�mU*H�2���պ��Q�O�	�"~#�rB�#�����k�I��؇�	�Ȭ}# HSm*M��Q
 ¡i���B42Ѯ���T>�	�Ca����;�|�ʛcDX�u�*Gs����a_�S��_sd ��k:v�u���Or�!�X����½�Ĭ�Ǽ��A��Ҙ�~�+�jEg'��+q8lȂ��!g���2�'��qڔ��NX@�mP#'�Lh:����"�z��gCC�2���@Ɋ�c���h������O&
�4X��\1	��3?���W�H`��W�`�-��˚U�ɏ@��iY���k��u@��	)��P���h�0HY��h����%����'F	��i½v�L��gER����d��pX$�Ucp��q��/���:�U�����(7< �}�-�"I.��A��!�p��\: ol[J<a�%�"'�e�ȓ|0Hۇ��-'S΅PG�F�u���3	��=�h�p6�L(U��X�B@�\S�Hڅ�����q�~�(W��a�F�h��;��C���['�V-te�`��9Za�W��J"C�=7�$��"�\Ő�@r+Y��~B(�ui��)���;	b$�>a�j +�R��bj�:�����̓R̓z����ă2F/��'l&ց��n�-�u+K)z�!{���7
� �ծD�p䑄��#2�n��K�F$;P�ςÀ= ��?oغ�j@*�C����?�	�$�U� ��yG%�-Kr(�1�:���2���yb����B���iã�	x�jس+O6���'p�ձe�H�Ch�]��c�x�1�C-;���D�3Q�:l�%H
d�~��w.[�KC�y"@/$.~��s&K��4=AD^�!Z'ܶr�����%�Gڛ��Z"k��R�'s��C�@�N<,$D{"�Z�0~�Q%�J�vq�I1� 9��m��f�26�QI
�v*�O��4��s���"\/ڱ��
_�2�ib$��g.,-�	�S�? |���Ȓhw�ZeMO�;ĊB��(��-�roI�V�ӧ�L>��|�E�'o	�3�h����L�$X�iB�-$��YfA�Vi�1�RߍV3�IX�AS!�~��rx�'���H�'�Z�"i�&�X�I^�^PP�I�B_�4�c�h�f��D�$��5�k�$( f�����!v�A�t`�A��q��A�P� �	4�&���
�d��6��">W�@+Ōx�0�
�::Ӆ�|�	0D,:	8׍�1��VĘ�K��㞤R��P�Q��UCvn:��$�W'\
�
�����*���y�JUTq(�	�e̪=��	��`�7,T�B�¼�ƣ<�ӊ}N��ݰ�vt�J�~��tJu��!v��C��#ʽ����^���J��Y�h��<Gx�Ȼ'�F�y�)ޡS=ܜ��$���$��US�`�UNQ>�z��c�k�a{��H�`�g�LW+��b`�[�q���R+D�B�K��.V�y��	
�;:,�@�%D�T:��D���=6l�{� �
�Rqz�Gե��'����p��)T�l�*��!n�\��H��9�圱cr�=�@튂=�}���U��������RE	�2�8��c�Z7�fYi&E�p�� E��y��t5c�u�S���\�ph��΃�h��h4��pafy�ȓA�y��O�N���F��f�K�лg��O�̰+�Bt�Cd�-p�D	�'����g�Q��E�/ �B�t��
�,��m;��ؾ
H�������0ZeC�9Z�1���>��qKU&����I	���O�ӠGD�
~�- ӍQT]2Y���ɂ;��jV��E�0ȇ�[Kw��	���AL <��P���G*q^4�s�eM`���i k]��a�/9V�����X�Ʈ8�|ȳfč�P�
�<�|bP&W�,�6�RFD�W .���_l�<�AN�2e�Z� ��-po���� ��iX�DLU ��4pt�rM?��C,��kOJ(�%G3(�X9�9%��2�>+��l�� TS�
�#Q�U'�fq��'ߖ�?1�PR5Xt�b&<Oġ���+��5��!  ;{j�1���
N�����@�O�����?1�B���f�t�F%єD�44�	"�N��xC
�g��	%i�>p�A��B���ɘ=��I�T��zb�����(P2��ͼc�:A�@A�"���%"O
<���^)n-����E���r���R6��<�"�X,5��;z2�kV�OX�<Y��n#�8�N���&M�3N�W�<	C@"�|X�gI$|�L	�`�W�<�&�\�zsМC���-1�	�rM^o�<��)�#F;J|�ă"�"�AM�k�<�%
�
D~ � �
i��i�<�Fmԧa����@P�Q�a���h�<)Q85�Q d+ۙ-i��J��d�<A�!�� ���gJ[�#�c�<�ŋBic�qK �@]�ҩ+��]�<�g�>G��}H�AAڠ<��B^�<!�l�/�p`�	)T~~͚�O�<!u���4�ㅫLp���TS�<ل@O1iFtڦf;����_P�<٤锪9���	�q
��Df�<I�F��!E��Ф�!	д9���K�<Y�h�xd�F�:M�q����<��٧H��3�Y�SԤ��N�<�$K��=�XU���z��Q�4g�~�<���;��\�㉈u�z����a�<Q��Ѹ\�M;���!�H��%�Y`�<Q�)Κ~���U.Yr��X� S�<���?Fg���G����4u�<��O5<(���[#{k�8��͑G�<��k�<}l��x��5����ɝB�<AVH��	0�T��`��u_9�'j-T�����Y#
��)��+ˢ|&%SB/"D���R�P� �`�bA�^�d^�q�
<D��hB@P���E_��qH�:D�ti��I�N�|	3��(���aaC:D��x��@?on��q���2B�Q!&:D��R�oK�#��Sp`T�6���7D�x�3��	X�y�lG3@<,!1J6D�� ce`d$�q�e�ЕX����U"O� ч��7�
��WB�{wd�HD"O����)	��|hHѠتLe�u;�"OR�XTM�jx&�ڛ$O��E"O��"��$�R� 6��"�"O^�$(˙���P�����"Or�N�; �#��^� �m�'"O��p׭��7�b@Y���3L
���"O��I�̃R7��M2H��"OL��
}��gk�>e��5�S"O��9�k�//�h�b�*�Jt.��"O,4�C*D/p��4s��-�Z�;�"ON�����{�������	��]�A"O8L���
��c�����(�"OXU���
$�~|�᧛�"�2MK"ONt�`h>�Z�qQ$`94"O�(�`a
<�v��U(�t6
���"O�LP'�D2�Q{��շJ�\ :G"Oty���<|��ֆ �t��TÄ"OX�#i���F���DC7�$��"O�=y�;*�l�S lI8�"O����([)tܨő��'@� �1q"O��0���:~���:0��15�!��"O(��웜պ��bk=Uߒ`V"On�����!4�Z5��?Tۆ�!0"O�t��L��t��]�La�"O�\�&��q�|�yr�nT�}rg"OT���)`̘���-L�49�]`"O��KH�n��	�c4@I����"OR1�vd+IG>L�v"�8_@�D"OXHHV�M�@8f1S�P1"ODc��*_a�{ա����-8"O$�as��k@� �B��g��܃S"O��r�K3�$)VN׎�����"O@i��H2��"���=r{��!A�'Yў"~
�"ۮ^�x����= 
Ԥ��y���F�0W�ءಠ�&g�<�y2��<P 0a�c�i��-G��p>�O<�b螐qP`,0��xT�)��	Oc�<qr
S.:R�q���*��H�Ec�<�B�5Gt��@�L;ZV�s�(�I�<�����~E~a�	#C���D��i�<iT��^��T"�!;�`��Bp�<��O�:
>6���CQ ����2*NS�<9D*^��tz��Y�2'��G��S�<є'Xx����.)��	S�G9�yr�]-����䐏a�n�P�",�y.LM�A����a!:%bV) �y���( /�� %Z�f�čÐb�%�yA]�.��pMߖ2b�I�#Ļ�y�g�&���A�-��D��� ��yrk�n�VYCЫ�%��0o���y�B�?"��5 ���_-�y��6	�$�aeJ� �^��$�yB@�s˂�H�mT�'�Œ�
̈�y�IHԂ���p�D����Ȳ�y���`	�}�"��a�:1²����y� ��.JYx�E,
=�\���J-�y����b�$	�Ĭ���ɲ�y��Ay�8��:����˻�yB ���b9i�&��tb���O��=�OwV,��CF3#&B�P&hъ?X����'k��d�L� nh�2Ȅ�5�F���0O��;Z��$z�C	���8��"O� ��k K��s$�-�փ�|��9�"O�4PV���?�����*F�ٔ"OR����2lFx��GάB~��"O��2ڞ/� c�4F�=j#"OT�BcC��t"�%(��1��(�"O���r��*�� �Lޚr��5S�"O@�r]�K IV�M'�͑�ʔ�yr�ŝ!ʤђ�G59�Ds$I��y"`!f�4 (v�^�2HР��L�9�y�
5��y��*�="�zL �!�R�<�R"Z� @,����2��iR�[H�<�UDB.k,��	D�ګ=���� �B�<�Y'��1#�D�0d���y�Ђ �>�[���r���.���O�*����qFx �v�K�Kt�k�)�f�<��">;���r(�;+�4�+�JHz�<qA�^�`'�.:Z��X�B�w�<iWL��	�2C�� ��l�U��l�<Q���7i�*R$��Se����\`�<����r���rE��'P�,��`�<��-/:�*�Y%�����M[�<�FG�蜝� �h���ʕY�<�
΂#��i�7�X�V�hYrԢ�K�<Y�� 2��Y#M]O�)j�cR�<q��N�8Q�a`�	�H�iCJZQ�<ٵ��>O�Z}a�!A*V���B�<�����p����Lp�5 t�]{�<QCae�BH�Q'C?(�10��Pu�<A�
+� :6E�2*�܁����o�<1V��� dq�E�U,V���S+_k�<��ƏT�V���F�x��Î�q�<I�%S]��E1p
Έu��hbD�E�<�'��!X}zV�X-!R�a��JC�<��_�~p-��DЅYliyU�<ɶ,!/"ڐJ��_ csjѩ��}�<Q��0u ���Ij�"yI���x�<���/	3@�* ��P��)YE��M�<9TbG�C���X�I�!_�*��~�<���^"(�@�(��S�>���}�<�!�$MJ�b��K�Έ�+�'�N�<i6��3_:�V.�}�,m�L�H�<��J	�K5059Iʺ�~ +ʓ\�<�'Eѥ}���Z��N5!\����W�<9�A�Er��Z0g<�Ƀ!V�<��ΈS+
�е.ʖv�Ydd�P��2�O�Q*ٻ!�~�t%X;~l��ф"Od"��	�d]�t�_c^��"Oܘs�I'�:M�3�ۘ ���J �O~�=E�$��lU����܂Z��ip�E'�y"��N@Ԁ�@�Zu�r��L6�y�̙�S��V,�h݆�P���y��@��jvO��`�(]Sʐ��y��?F ����ϖ�0�v�#��0�O��"�^�|��mՀ#*�6�b�"O�})������H]'2�,hRt"O���e��>C�@��ӧ��=��|��"O��r����|y�Lp�)�dm0�8�"O,L;P��}�d�B#�ٌ4`�A�"O�,Zfe����#��\�.J�1�"O��i �EU��a�o��W.��q[�PE{���ӃU�a1��-\���'�NdK!�D#k�dS �X���C��O.!�Ė�U*ȍQǈ�
6l�{Bi��*!�D��j�x��$�C�f�{R�� [!�� �h�v#	$��	��gJZe�%b"O@��g��1TPb$Ϣ>~���"O�M�C��8�ת۶@Gz�H�"O�|c�o8W�:5��M�M ��3�"Of��%��g��䳕(Ӹf	JIf"OP����9ր��'8�(�"OTl@�MA*{�KY3hJ� 7A�6�y�mB�
�)��[&8�Ca�ǥ�yB��8q�&`ZGƃ({��[�̕�y�Q�#8R�wbY�$���y�G
�yRL�	k�q��n������y2�n���*�ʅ�5 B0�$�yR+D�C���$�.R�(s���yc���vLU8����&�D6�yRX�|x<Q��X"2�(���U��y2�?"̅��=v����ujV�y"-�=0�X�J�(['@�`��d̄�y�L�P-8؃��țK�*ň���?�y�Ť]*�#�*G[�i�fϏ��y�@�-�6�Z���)>h���@�y2'۩b�n@�BD�~�ڱ�
�y"�P��N�
$H^�u��x��]�yrnO�X2Tl9�#	�E�4{Pȃ�yr��4���s�*�`P���W���yrL7EV��[b�*�JdBD`��y©ѿn��{c&Y�F���ĈU5�y�Ȇ�B�6�0�K��n�ԍG�y�(�0T�v���f�>	c�HrVm<�y����J�$���Y�-T�k#V��y��"7����\/rBH��K2�y��Hyp�	a���TAV��Tm��yr��C��i��	�!Ki����y���{�`�B��o�:��E
!�yR��<5J~�b��&(�!����y���d\�����	�\!ҲcY,�y"�]u������~�0��q��'�yR�˨F��4Rw��:,߸0KfF��yb'A�*I<)1R�R�Y�Q�5���y��O_��D�E�C&��`U�-�yRk�*$�*�����ZA��6�y"鄒5DP��g
��y��D�k��y�
�Ѭx%&K��>�Q$��3�yb���$��]��G�w��X��ރ�y���Qr*t���٦p���Ai���yB&�#�X��ffΓa�� ��=�y�A�<G�e8�&�D�X i�
�yr$�[�
��Ԇ�{(ѡ�e��y򪆤f�X�H�g޺y��xc-��y��h?f�	��ԩ#x @%�y�(\0v�~5��/Ý7��B���yb��<-BX���_%!����!�[��y�GH=S�Ѐ��Yِ1cA��yR,Q�\�FQQ��_�}�f�h��ǖ�yr��&j�P!�d-Bݖ ���%�ybI�1���Ը<��� u���y�@� l1����
ڣ>����
9�y����T�(�Ka���3���`���y��|D����.�zek�'�y��3b�i�K��$�*�k����yR��]X��	$K<y&<� �N�y���u�`�qC�~�����J��y��!~��3���:n��0�ɵ�yB�V�)Z Uak��hC�\�&�'�y�ƕZ����IL#_�X�0����y
� @��1b��5����WY*9|=a0"O}:'�Y5J�K�,��Р*Ol�Q��?o"y����%��'Ǵ�2�<=��a0����jp�'lH����5���&#ku��(�'e��J$nH ִ@��OJ�^�b�'����چ?* �(Z%h�����'kX���\���Q��G�6rq�'���5$I,
I��敉DP����'!8�Ȗ�-�`�a�K�9\���'D���聙?!D��!�U6)��L��'YH������M���<��'/8�s�e̶@����w�؇f�� �'$�TI1E�C�9�m�R�c�<�
ӡd��IĬl�na�r!c�<A�k]�y������휟^!�d��f����(G�	=�Ļ��R�6U!�N���!�%M.��hicM՛F�!�D��!��S�&Z�f���(�&S��!�$�f�RD�N*g��yAsD1J!�$U7S;ʱ����M�n$Q&݁y1!򄚊m(�pAKH�Ep�i����')!��O�=k���=R4D]�"�s!�dR������TL�0���Q� d!��T.��z�<d�*�!���!�D�,-�&k�C\�0��T�����u�!�хa���bL�8T���2��&k�!�K6H�*�F��-$�m�C�(r!��U�D�����[3,y��(N��!�DQ$�ѡ#B�B.聲aܮ�!��(^X:��Y�c(\����LX!��L�%Z���aDA�O���6
�:5�!�Q|Bt� �%�P�iոp�!��M�j��lX��'\�pA��� {!�DZ"����Rǖ
�f�uNީ`!��T�8b0�<O����U�!�O��515(�� �N��[s!�d�N�� �%�셹5�NgS!�řH�쳢�A�P�݉��E�+I!�_���xq�[A�T�q4��:!�Dݠ\t��rǇ��|+�^�s'!��0��Y���~�ɺWMD*Y"!�ā�u��i�eHO�ʪi!��S�h!�$% H�K�̈́\x�b���o2!�U�I>nuX%�ѡ�PA��E�&B!�dW�%�I���SE%��nT�M�!���%I���#jV/6a⠢�͚�Z!�ЈE� �I����L8ʕBBl�1$!�$�|#Z1�g���i%�5��N!"f!�$�N?�Yk�e�02����7i!��8�
G-��
���'�=O>!�$P=��v�T�.	\0�2&J&6!�$�?�1��H|�d�Gj�t$!�X�
]�,R�A.Z�*��/��ko!�D4W�*u�qg��\�x�u�V�0V!��f�8�7���>L���F�!!�[�{��r���Z�{s�D�s�!�� �!N����zmB}0p!L�!�ڵk?�S4�HT�Q�/_�}�!�D�ݸh��L��2��1�!��:�p�����ΤPQ��)�!��,w��.�	q�4��4��_�!� xu2����u�����@�!��]�u\�� jX�^N9�QCQ:F�!�� �L3��B1���!�&NrL���f"O�Y3��S2 ��36��O74���"Ov�4�����8��! �"OV5�u��a~�!�^����"O�Q����\M�d� ��2t�zYz@"O�9x�&�?:00���̢H�5�f"O��!A"�f�q�B���f"OZ�J4��oT��� $~hx��"O��Ѱk@0����	!
9s "O`�)G��)8��M�'�&�rU"OD�j���+%���B��. ���w"O�|�3��:����M��@��"O�E�c��z3ޝ!�֣��A�q"O2�(Q�z%�����^z(�	�"O��C�,��z��=�1Q�XW"(��"O��P@�ǖ���6'TQ��y�"Oe@�ԕ5�᳃��661�"O>0zf��bP��J����r=3�"O��#&�V!s���b��j┥�4"Oq��O!w휅�ӆD-E�F�*�"O��k` ��;�8��Œ�kG,u�"Oh1e G� �cd�%I*\d�F"OƝ;�/�,f�4�e唯=���6"O�l�fc�62��9U坯z�NIq "OP���fؕQN�00�i��2pp
F"O�<Q�	�O��#HU�;�>y�$"Ov���쑑}���G�(���"O4������@d�M�ef�zn"��U"O`+� S>%I*�#�V/`h
T�R"O��&�A.�z�a�$�Pe�"OJ�ْ���l����Ά2��)��"Ol��ׅ�� �*%x�V�J�E�"O
=��!�;n�%kM0<|�s"O:��A�����!9W�H�"O�Cdትf0X�e��x�\��"O�q�A�[�j�T����|8M�D"O��E,J&z7� �$�ҷZk�ia�"Op��c������c bF�D"Ox��'�ޔn�����
Zn�BT"O���u��A�P(Z���Z$�Z1"O4�z����2d
A��O��[�"O���`�(Y�n|R�
�:(�y9�"O0)��9/F�X��A�Q�^�;$"OV���>t>����ߌ3�
P	�"OΘp�ą#9l��CA�l��l"O��P&O�8f,E3E"��+��0(b"O��oԎyq��y1�>	u(�"OB!����+F���*I�B�A9�"O�I�uD�7����$L2�h4 �"O�Q���.����2<��jt"O:���Y>m?V�*4��x�@ �d"O�uR�$���dQ�	J�� ��t"Oȁ�0]6sSXe���۞Kj�!��<}v�*�-r�*ٲ�E�.>�!��#�D���
��f���0��L!�� Q5
hSߧrа⃁\�=�!�ā,����t
� [�=YcǛ2M>!�dԼ*,9�vb�k=r8C2F>
!��!Q#����0I�
���K
5�!�$$uy�I#Ўߥw��ؒ��H�!�^�|:��%[����M4 �!�T7XnP}��k���H�kDY?�!�dZY�����@��f�l8��:R�!��*�h�� �S�kn�R�.�1
�!�� ���`/T�3����˗�?ٸx("O���oةr8��I�$^�"["Od5��@@y��锟Y��r�"O�L�C��)�Z����hPy�7"O��Y̸t�\a3�A�7��3""O��1`��'t(h""�� 쪅�C"O��AW�I4 �t\b�炥b����O����M�>��R�9i����-�!��
�3����M�bJ���� ?����9�g?���"�(d:��O'2��TI�<Ya�[%]��M�ej�'3ŐMc�A�<��X=�F�z�
�.T}QrW�F�<���_
1b����,N0*�ɣ�I F�<a��޼d	��RO��A*P���Yz�'�ax�!�6PV��1g�eዛ�yRl̖~�vp��(�)d�"a� ����y�C��+��4�&�h⼨�[-�yR��R��:�̠{��m15�1�yR� 5tG.���M�<+�|������y���tVa� [;�6��RD��yROC�~I��d7�ʰX�끬�y§�G�f$��+B`�(V�Y;�y�H�x��� 6:��5e]�yR����!1P]�hgXh�d ��y���B���5ش]�X��t�@��y2�ۉ�0�hs $�0�D�͉�y��ȭ9u�	���C|�X!z��y�+�=�>	�"�HK6���IB��y�C
.V�1@�g=1��� ���y��K�Se&X8$X�vO�4���y"d��Q����#�0$6���F�0�yb��>c��M�a"_�w|��	���y�,�(K\���  �aD�Г���y�d��ިK2�`v��h7#F)�y��G�)��Q6A	�V�u�uF�=�ybe�{�`i l	eJ�<�wHI�y�i�
&]8������k$,y�GHN��y�S�[�6��`� `��A�7��;�y�a<3�BP*�\�R]����
֞�y��G %v���7L�� ���V8�y�Ț39�b-h���D^�̢��Y�y�˫T$e���8gl�����y������g�C�]�u��gN
�y2�;=���9���ר�"��#�y����v�P��EU�C�\���!��yR.<�}��'���^aC�����yD�>������R���NX�y"��>h�����æ�V�C�Ց�yr��J<%�� �x�.����y��T��LxR4!ƀ}�p����yb���)�Ai҂
# ET ��-���y�o7Ki��1����qCp�@G�D��yBLM;j��847`��SV��y��G�=1t4 �0]p]���y2�6{Ô�0a��!x����	��yB�ڕ.D���6�N<?��wd5�y2Æ�3c4�bSÊ�d�ē6�ڍ�yH�,)��ڣ)�i�&�ۅ���yC�P4�[�a?x�H��1�y҂V�IdE�vKD�"���j�m�y�mІ+����B��"�튵�D��y2�܋C`jm�wɊ
���[=�y2�ذ-b<�7�L< vD+���y�!��N�� ��	�j�fV��y
� ����G+l��Xj��J�_M�	"OV�A��; P��� S�qEH��"OH�ڢ/Q:��<�P/ι.[H��"O��cS�B��r(;��{;�mR�"O@�5.Y2|~>(!���O;-��"O� A�
��w�ZY�����`��"O���ޒn����a���I�<�ʵ"O�J@.O[�Y7Iΐr�: @�"Op��rFC�Pj�V��:���T"OREJ�bē��I����T8�"O6����j/&Lr�v��b"O潀Ơ�Dͺ�S�#��)^�܃T"O��#A��@՛U��Gѐ�"Ozp�ƉB$�,,J�&r�B"OT4���[+*:���	��a��"O�0�I&�JI(C*lxy�"O6p(�,R�dB�zc�_[����"O���^�^�Z��6A��O\�AZ�"O��@�W��:`��1e?��"O$��#� 2pNJʖ�#L����"O��#p#�-.�йP �E䅻�"O��EÔ*.
a��!*mH�"O��KdB����ƌ�h���:�"Oȯ"Oc�i��f�b]�����TS�<���,���Iv䗐sv�a��g�<)�%٘~���b�H�N� �K�$I��G{��iL�m�|�1mZզ�A�+�t',C�Ƀm;^����٥àT��F]�l�C�(o9�iwb�\2x��"�Pʣ�9D��"�&P����K�,(�,2D�$p��ޢզ����B<R�;q&0D���G/��](�U�mk���@�,D���%`٭i٬eňۉ$����@�O���(�$�|Fy2�6P�`�a MPy�d��y����#ƨt����#j��H�M�y�ą1J餬p���*h �h/	��y���=w�eJ�"!-j1�͍�y�j�3$���)�┻g ��QF�/�yr	.��M��B4Ȯ�0(���yb��C��Ѡ��Fw�9Ë���?����0<i��"9�zո@�X>WH�i���L�<�֋D�G���B���96���dɊI�<Y#(vY���@��cdjl�<ic��iD�`���8Z�q��6D�����)Ɔݓ�Q-��+ŏ/D� �� ľP�ХB�a��yCd(D����!�
�Dm�t��#5�Hho%�Ip�'���G��:E��K�� '�ԩ]C�	�BD�k3��Q��$��˒�WB�I�<���ꐋ��"����4y��C�� )�2���%J�7R�PrJ�$�C䉺~F��re�M�<l3���$#�C�	�^�@}3�fF	�6��7�Gq��B�I�z]��	��$y6��*E�Q���O���U�c&�vՠ�s��H�"/ڽ�ȓ�8���%�4����Ջ�/A��D��ai���B ����G��(>#�@��Q�֍5'�2�t���C�,H�t\�ȓx�����N6Y��A D��)V}��ȓ&�H��	Ə�$�`���%(b
܄�O��D���RHp
pG�U�,$���x~@�
�^i���ރu�p9BeG���y�%����ma��;<�C�E�y)Ġ"0]���/�.�꒢/�y
� 4��7�A���k5��97"O�I�q.�,�fd�у�,F�Ӓ"O�Ȋ4�=;�U ��:_74�s"O� 1+�F�<�Z�RJN����]��?y���?)*O��ӑY�X@�OG<�� �̆%h�~C�Ɇu�J:%m�Q��b���
PC�	3Y#�)�)0q,���o�oQ�C䉀6h �$ �%��ђ�B�>bt�C�ET4b�,M>tڽ�O$żC�	#4+��C�	+��¸M/�C�I��l!�Fl�S��ue��?��I�hR1�2��&`�f�L.@+!�d�l頱{�V?5�(=���|�!�dX�w��!@��
_?�	��ԬK!��?f|�2х��O�y�)<% !���d=��2a72Dc�(�:q!�R li\��+�r� ����o�!��X��ęź0�0i��l�{��'Ra|��a��r ��R;��Kv'��y"��]��e�i[\*�{M֐�yR�0[8X�õ{C�@A��yB��0Ѳ���V��������yBԤy�h��Ń�#��iʂ����y�#��Z �9�Y+/�&E�vbĤ�y)V9	|r��b�D�*���3��<�yrm�"Y<�����W�#������y���Q�r�30�Z�K��5YA׳�yKV�7�`��6��t�N�i�%V&�y���%�"Đ��=n9� �h�-�y�'O) e���ǬR�{�x�S6��5�y∆�s�"e�gb�m���U-�y���*����+"n�Mi�ǒ4��=�$6O�m�℈�t����L�%:wVlqc"O@A)��UO@<h�dJ͑g`�A��"O���UE��n˧SyN� ��ǚ�PyB��g�-�h�#R(�����d�<IծY�����ץll`j+�E�<�r���P�5��d�8�h�ɀ��X�<�q�߉;�*�[�Ө\N��T�<a�o��2\��nQ�z�-�!��S�<ᦋU8���ߟw��p�J�<y���$��|���S�sRU��C�<��D�Y{��Q��O^n�pc�|�<i���>\����E,"hU�P��N�<�U'�&$��D�4F��98��b�< %��9���Q�)���F��`�<)�G�S�q*�KV�)�!9@$BY�<q���b��E���ۣF����R�<��FW�+���j��
�
r�@2��X�<��f��(�U��ɔ�}����i�<���\� �Q��	V|x�B��M�<Qd�\�1�(uf隄hB��I�^�<�!�#�h�y���E]v�I�I�s�'���>�ƽ�*�!%�e�&�x�nC�I�2Pr���' j-I���,�HC�	�Q[�x��1D��1��)]�*C䉝%fuzW�B�;�^-��d\-m�B��1
.�<��i\�hF�C��z�B�ɠ	@>��ŋ�;�4%ȱ��v�DC�	�i�D��Q4*C�@@Y�~J�;�I��p��}�'Q��P;�EQ3����.G`[��0�'��1w�xLa���$P�����'���D� 
�"�	�����z
�'�i���ۃ�~��p႔(���x�<� ,E8��R.r��E+uŎ+c�R�Ц"O*0���&3gđ�g��px�"Oqs㦟��Xyb%�� 2���6�'�\���ȟ�'?)�OnRxCE��J�l\Ӱ���o�@
p"O �i3 E�U<��{���0F�a�"Oz,qݧ}�L��R�۶5Q��`�"OZQXJ �M8J%��|H=)3"O�5�RG@���d��ש}0��s"OP�iP�س36���(M��@w"Oh��+�
e�DEt�g���1#�'��'�2�,8RJ�Z�l\0	UP�9Sg\?6L���e�ީ��EE�hƭ��?&���&�\P�/��X�`�	�[-���ȓ] �"`�޵{�fE!�g�6_�q��@�D�X2h��^p�%�7XHM��aV�:P-�0p�T�s��/\��ȓ0O �u*�~���X#c�$��Iϟ��<��p�X�P%�2N�d����[�<A���x���~�V�� jYQ�<y����V��XR����r��S�<�ei.)o2���*N�@.���Ij�<������H�xw+-��)�d�AB�<�W�E�Nu.92A=L�9"�Ȇz�<Y&�I�F5�����j��yx�x��T̓v���RlM0"�Ƶ�Ŏ�$� ��|���ևW�1X�a42��M�ȓad�cS˕+	�:�)T�Aقe��ck��a�UO�2D�@�Q�P8��%Ȯ��B�ԔKYB�)�懗��ȓe(�Z�-�{��ei�P5���ȓ���ȴEZ-)l�:��{E~!���韠�<�4%B��c	�
�8��Nh�<QJ��O�`kŁR	'�XR �QN�<)��C�W�p�E� ��xL:sAR�<)H�R�R1� +޿	��4���D�<A�������c ��bL9ˁ��x�<�PmJN}x#�)˵n] p���~�<��-M��q�p"=�X�`�)�bx�H�	y̓L8"L��f��l����qoZ��ȓ-�0���JX�R��h{2�>7`���ȓz�tE�1�0��0ӳM�3{��Є�}�D�kQ�G-n���a�(L�qh��ȓmN�و1�߁}�Jܻ��̰G4h�ȓ
����) ��Th�26��ȓe�-����'b�4ků�	?��4���M~�+��$��咫[L���H�#�y��n�<�.S��qkɅ�y����n��=���@j�������!�yB���..�) ğL���X���?.O�O?uIԇ���(;1��"k
���NL~�<ђE\�k�
��� M�`��	�6�
_�<1a_�	�>��B��i��Y����X�<��i߯Sa<mQ�ƛ�cǈd!�X�<��
�hrʹ�,�v�y�Ҋ�[�<qbÇ�C� ؤ���(�փc�<I2i�l*>�!6��a�i����D�<	��F�aĐ؋g*	S�0�2�C�<!�eИZ�T��NAXb���M}�<��}�rp��� `���1�z�<a��.��T�� F>?~�����k�'���'�>�p��<�,q�W,Ҽ.f���(7D�|{R$�,F����:$ �U5D���A9l��Ph�\�_	�5��'Dў�>�S�2c  �Jc�*%.��D<D�� ���󂌐E��)@�(vid��"O�)H�-�"h���̃�na ���"O���+S�(eD���g}�=16�������J̧bC+#؁j��� ��vf�0 "O|��E�Dv�Vճ3I*6L�3�"O�	�ԥ�1N08�摪W�A�0"O^xⲠ
"��K����V���+�"O�8�փ��JF� ��O�fI��"O$�YtK��\h(�0vl]�z ���"O���")%H<A�#(YPGT����I�M�d�g!Y�Qb(�h�C߀%�C�=��� u�E�-=@�i^v�2C�I����v*#2�r$B#K�#D����hOQ>���Y"!_N12U2zW�}Y�8D�`q�$�-(�b]Ç)��PW���W""D�l��#�!9��A����tn�iw� D�Ҳ�3[���j�� F�
��>D���䏒yf@8�~cحpA?D����,6d�Ԣ�,]{Pz�/��C�	yR�%8��B��bP"�F @��C�	�P��}��O	*��<��%�#0��C�{�!��jU"F9ZP��E� G�B�	!�`�B���R�d�W$D�E:B�	�i�N0��C\�Q.�3BW���hOQ>�p2f7?���� �#c�f���9D�@�� Ĳ�ޠ�U��&}�bB�$#D�4hd
)�$m!��A)4e�a
#D�D�@9p�b�ؼ �lA�a'#D� cp�S�i�-k@f�kJP=�2"D���W��xI���d �
�I�>D���7&�XE��ʖ�1���VJ'D�+Ĉ� >��丠#�3y�Q*�� D��j�Z�~Ѓ�d�	Kp D����k�65|v��2�8/���Q�(#D��� �Y�Υ���S7s�`p�e� D���q������0�((,,Ĩ�D4D�0��,��؁!�,�;9]�s�K1D���#ɔ<K�Z�*)�%lj�L�Pm/D�����
S���!�S�Y� !R..D��yeMΣ5����o�,-}&eSAA6D��@B�$K�j�R
"�$��%�3D��GnT�K�$��,YX�RT�/5D���'oW#.(�SO�;x���2D�<���D432 1X�T 3���Sc2|O�c�����X�~�[ �^�F.�@�E2D��b[B��Z�CɈF(�F;D�1�ۂO	sUo

e�x0�7D������j��$�e	�Im�Ec�*7D�|{⨔55J��M�<x��h�M3D��A�̄I� QQq��$[\����5D��[ʍ���uH�Ѩ*d0%p�&5D�pbë�~�X.��Y� q:�.D���t���vQҤѰ��Ӹ�a�%-D� ����4*L@�b��+^�Zi,D�(��h鄀CR�� <��a+D�$���hl��7	[#4�85Z+'D��6���tD|uX��>/}x@C&%'D���2�H�q� �i%�|���hG
$D��kc)!V���AF+b���@/$D��2�@�����rF�n�|#f�'D����A�n��}�V%R�,�vT�%+1D���t�A�#6V@Ĝ	lRh� �/D�ԺS�գV�>�yR��9�<q�,D�H�q`�;�%�c�?Gp�8aM&D�� �dF(��Ud�H�#�"��#f"O���Bh�C<>��fl=_�صK7�'���_����#�)1�0�:��$D�L ���)
�|���\0TSh ҖM!D��b���r��"M]6"� �+D���v�� ����g�]>z��&�4D���a �YR%1��B;6�8v(1D���T�͋{uz��$/�60�0%D�tȗA��9��b��C�U�a�Q�#�����z�k��N�°2��'���"O6���h�9yu0�"��@�[�|�`"Ox��R�U�d�$z��4{�R�!�"O>���k�mgJy��C5<ta�"O�d��k��{�<�;LZ��"Ovb@�ʾ$J���KΪeH�!"Oz�#�b)U���s
�p�1q"O���%ć]>��Z�ō�:b����"O�Q��#��I�6��X ��v"O���"��?%�4�@w�4+��[�"Oi�Bg�<5�P�bA	 u�"OJ���ܠ[e8��b�O�p�H�"OPђE���42�Uw��(�W��!��10<�,��
��p�- �!�5y��!U,�9AF�Dq��]>#�!��)}�좥b������s�VQ�!�䆳
�$�k�Wx���	ɖd�!�
�شpA��-g��QTG��!�dG��e8M���M�ѥ�z�!�׼h��"�S��P����S�!򤚮ca�m�3���/���q�JҎ=�!��_Y|c��A�:�����!�$�vzI��O	"��ă֨�T�!��5n�x ���V�YSЫ�&�,E�!�D\�np( ⷠ�+&b�9��*޼	�!�$P:����%ӒV&��`�#�!�dТ@:�Xȁ�O�R�52��4X�!��N�%	���E��Ā�d�s!�č�)�z���Aȍ�p�+�b�p!�d�)�,�(qċ&@jL��a3J�!��cB�\br"C<q�����	�!�D�x|H��gۃUs>ũ��X�p�!�խ �.��uZ���i^�"�!���X��d�"%�p�FgC��!�&>0�0seLʹ4������X�!��ۣ0�X�6�]h�����׉[�!�dR�k{�A�ElWlZ�h85 ]�!򄔻 -�д����F�Pᥚ<I�!�D�m3.�RɝH�ച�T:!�dT1KN:��g�/���[�H]�!�d��N�Ѝ���!��愷��{�󄁴n�`�8��٘q\�[�̵2�_��%�"~��\$=v}�҂(83&1�`���y���1^L���.���dD�B	��y�F�3ht�he�٢��}�*��O��!E�'���!����d�����-oTL��'�T�qU�<<f!�ǀJ*�ź�'I�Hx�d���5�Ǒ�H��{�'�̑*�C׀4�p�����	�nY�����'
�>��v/4��̣?&�� q�f���#D��/9͌dZ�
ւe?��!�U!�4l6�Fɚ$EX���aa�[1O6#��'�<���5.P4:�◅`���'Ѐ]!�nي7�Tm�@?h(�i��'%
b`��"dQ�7�d���y
� j��Ă�� ��Q�PEV�l��c�'ў"~bQ���r9>
�iΠ"��3PO��yR�W0�l��#ҿ(P�� ��;�y���Wwhb��#S�,�H��Q��yr C���<�'b�+Qn���̖-�y"h�5� �ZR�mℇ�i��ȓkJLuH��T��!�JC������ǟX���'�d���Qؽ9���rq��rjfz�* T ��1%�CJ�ZT������􄎰C�	f�j��ȓ`2��b�i!L(��cGbȅ��I+�
��D;�!�0��qA���ȓ�d�f���C,a��O���ȓ}�Ubc�5"Uzx+R �@�.�Ɠp���&c�F�ZEhF�*j�\���'��Cw"ά��#�Z�P�'&\Q"��u#lXTI�_���'"�B .� w5rӁ��}�:�'������M� ����r�,ElJف�'�����ÝLq�u�1D��&\6���'!TT�\M�5s���f��'�
���j�3�&1��Er"�' �E!�O,6q�c�	����=��'k��ɒđ$�`
�
�5Z����'�0���a�3W��逵�� )�S�'r�qQ$��-��}�NI�}Wz� �'����b�G��� ��q�2D��'�Ĩs�m�T:����	.dY���'�,�8���<R�>P2s��q t���)�t��/2DˆFJ(���{��N�y�OSτYc��W�*U�i�g��y�hG�8����Y#mxi� ܸ�yr�E�x��f)�*`��V�y��b�� hSP���A�D���yr�>�j�(�@^�;�L0���ܵ�y�Kŝ.��C�+قK�л�I����?���(0��a��C�n^4�Їȓb���ĕ2W�����n8��/�Ġ a����fTU�H�ȓ�� @ޖTr�H��nٜeLh����L@,$��0�ˋ����ȓ'��D�!ɚJT�i�������m����*[&_��$�,g��ȓ8D�b2��H�7��U-�%���	.�<�3	П	cT9�b,"�B��=�I�uA0|.�J�L��L����0?ѧ�ߧPN��rj��QX)i�G�<�n���PaC2���J�0�ĊGn�<��C�X��P�&.4���;�Hl�<��e�p���3���/�3�"O��
�
,!����5*�r�k�"O�	����<0>�0��D茀"O�)YR �1Dd�a�kC�U�h��'n�	
ׇ�L�� �d�q��'q�Xb�BX2,d����KӜC\�H�' LIe+ǭ3���Q�[n��x�'��]
��?%h�C��Xv~]��'L�jv��	._� RC��:h��x�'�xu��g��x�j�Xb*�5=���'�䕫EƧwy�%���[����'�<a���^���a�Y.���'ch�kC�X+D�|�#h��S�'m�!{R
S� ��S��ZC֨�
�'��m��A�i� �#aS%P��a���hO?��  a�`Şu���0�!(~�� "O�sa�2d�d�sǏlԩI�"O��#ULZ8<��jd�K�6�:iZS"O�|�e�R�A�bS�O =�"��1"O6�*`O�z*�y���5-�\"O�=�Q��+Q�ej�ɞzqA�"O|��EêI�� A��ik��0�"O�ŸP-UD֔Y�wO8X\��'�|��'l@�[�G��٠gIƤ�
��'^�;Q�Ŵf>��@7&ӥCqp

�'����½{;��c�;`n�	�'��xK2��; 1�Ia3Q�@�2`�'g��ڲ̓�;i ؓs'E��J���'E\a���_R����m���h��yRϋ+L��a�סޤ����/����O~�d6LO�����S�Sq��.a� ��"O>5�@�މ_E�T@G������"O�����b����&E֙2�x9I"Ov@i�lP%�>�9oM�c/�)T"O8zc�ČA������_�H��"O�E0��<{���WbG���J��'\�'mTI(G��f<R�+�PRX�*�'��t���$5�H;i���x
�%?D�8���F�K�2+@�O�|�N�Y�1D��j���2��0X��ȃ|h�Y��`.D�<��ɏn�.i�#GF����P�H9D�\��A 2|t��Ą .����@�7D�xك'�h��}��@��m� ����*�O�I�/�Iz�	 ,0?�(��N�=]���O��d+�O`̚����^9�'
�"Ơ2�"O���G�J�1+��'�Cy�"O"}jtE��j퉑�*G�V	&"OV1x��W� �#� *��4X�"O��Ҷ	z�^2�� 6S�`���"OX|�q�G��I�ʚ��1��"O���ũ֙C��,�&N��ɀTQ�W���Ia���EF��3�J�O'Rmp��+D�A�]�X�}��XKd��i*D��
���k�D{0'̴t~8A:@�)D�@�S�� ]���Sd�e[ܼQ	(D��p'ō�:��Ahs��/V��9D��[�hV:ttx���աZ��ჭ8D�l$��Y�0Y6�V:i���p�$D�� �����7�S}H�q$D�x@I?Ct�0"&!ǆza��1>D�`�6�O$!H2�F�51:J��`G<D�DqC��+Z#u�R�\��A���&D�0z�!n�6ې1��c�F7�q
�'��<��HL�(㠒�D��	�'6��B� +=dr��� �O\`��'W�h�`ց44��$&�3�`��	�'�p�Yq�9̲�����!���X�'����3� �,vЩ�#��<B����
�'���9"-��_���g�?�I
�'?n�Q��8/��Q0�֘=�N� �'� b�n
���[���0��
�'ގɂ��7n�ҤHqk�61)ְ
�'>�( R�'g�L �G+A뤑��'��8�6h[|��J�#S	wR�)�'M\a ��^gw�h���P�y��Xk�'��D)�
k$��i�*�x��i��'�$�p#ѐa�
�Jf�����=��'T,���U$2Y��i��T�v�P�'�F�h�O���@�+�I{���� �P�A���"`����`"O�ɤ�E�)s�����9}@���"O�$�Љ�T؁�S��4U�t�"O��R��<�1F��&_$�P!"O@���NS�;%��B�ןN�H��"O��^�N2n�� �'U��|{�"O�Y�Ӧ!K�f=2�)L�'�,��w�|��)�ӿ&�\�3�ΪQ����3R)�C�I�X�>zT����ڀ��l�%"$nC�I�F���	��ͯg��tH��L��B�	�n$f�@��	�
P�qQ� xC�I1�:```�%`�*��7����B� ���R�U-d��BmD"$�C�I�_O���Ń�&^�v�E��;Cy���hOQ> �ӊU�H�D�	*�{�$D���7
�<7HL=�v&�-V��h�3�%D����
�Sܢ�A� Ў
'� D��Z�E��t�'%[�����)D����̲9Z�b���<V���l'D�L �)���ꝑ�!/`\��0D���!��/����!��BD�1�)3D� Raֳy��u�R��Td~�{��0D�`+�V)�l�p$���D�´�#D��Ȅ(�?f琸�P�_�B�ó.?D��@��E�W:y��N5CW
$��=D�@�M��%���[֯�7(������1D�X�`[V���w���}ȵK�*D�$ �eZ<A 9ې�S�B~����)D�Ъi�7�(��'G�,�P�'D�p��`X��a&��[EfͲ�A$D�S�@�'5���-ƗZ���q(8D�ث� -�҃äZV��7m D��j�JH�+���Ȁ����� �#D�@A�/��*��TҀ��-#�r���#D�Xq�I�%�b�'aY g
*���!D�����P�OphB�=5�J��QF D� �����lڦ���DƴQN��*�,*D�Pȣ��(wx"���(
F���J��)D��0Q�E��hYSQcH����	U�'D��ǄD|����3�r=�gK&D� A .R(A���� lL
��U�")/D�� w�_�SxL�"G�h���d�9D��3Ŝ�\k��U�e�o:D��2]�ThT�!���:X��*t'7D��1�ޥYr��t��S�R!k�+D�lh/*r��c�U3m��t�;D�02V� �v���#����&ak��;D�H(�Ĝ�"��83/����rA:D�����I��*؊�Β%<��j#D�`���4L�&`p�D�Ǧ�iӧ5D�8�գ�-�j6I��"���@�3D�����:4�h�q���;��ق�h0D��H#�R:L>ܩp��}\��D.D�{@��8pJI�#f��i�l � "7D����մO����&W�R*@B!D�����PP� �\�6�z��?D�$b"g#
;�:�g�Z��7<D���CH�3C�@��꛽e�
��;D�(���Ё$7a0'��]4��RC�8D��sT�E_"#��9���#	l�<)d���!T�DP���%[��RpAd�<��VP����ơm�0����`�<Y�GW�<�|�:�C�6����e	[�<�%��(=pB�AGK�D�V����Y�<� ��h�ƶ~^Y�f_,�
}*�"O�4��٣t:���U�z�\u��"O@���k�|��oɞA�q"O�YYa�I!<Z`��'霸��i	v"O���N�>(��qt�0�����"O�ĲB,Xe���K�I���6�
&"O����ѿn?nT��ȁ-7��:d"OĄa��H T�Bǚ�x+`�S"O��h���F��H��/��L���b"O�ڰ��f�F��גC���a"O�����Q#O�V)XS�Ց3�\�C"OY� )̱K�)�Skڅ #�$ �"O�I)c�V�g�jp�D�TΉ��"O��@�.\3y��w�t��1�"O�=)��̯eu��C�N�;�zQ�"O�xuC��~_\-zs���|�*"O�h#)Lq���P≇>S��4� "O��XQ�)+ٴ\H�i�:M��|0d"OT�p�ڱ_��(@���F�
y&"ON�T�� �x���UjԼA;v"O�<+M��C��y	g�� )�r"Or�p`K>e~TQ��D��X`��a"Ob(
�E��f����Ӂ R��	U"OFud�!#p���P3�(��U"O�A�GPpm�<㐭?Y�H��"O�-���?;�,l��L�+ns�"O�@��+�&Q��8��J�X��U�"O@L9�� ����*��-�m�c"O4�St��CfQ1�^�(�@;"OnAC K�{���S�"[���
�"O\\Kǌ	�p��V"�g��4k"OM��h�2D��+��l{���v"O �K%dȂ>�t�&g��{`�,0f"OBP	�_;#�<$��bVZQH�"O���@j�./��X�Be[��ڦ�Hm�<��/S�/�`Ȼ1hP�$�L4���Vh�<!@�W�?������P� �ɀ@��e�<1���E�������"9r�*\e�<����l=,�F	_/%���E-d�<q+R��n}�s��;O�<Pbm�G�<�������1&��}t��b�TK�<�īYVP�Ъz��[�	RK�<�P/�aA�`ڥGU$~�mC!b�<���x���f�K����r0�ME�<��)�T��#�)s�`z���C�<���Ȑ$%����	��}�y� B��<��C�O�V�ٲ�Q�LA&��2(�z�<�,
Nh�9��H
@\yCd��M�<�Պ��8�BH��j`�AP��J�<�&� VYJ�����7a��^�<��/�*M��S3g��sdT�R5"R]�<�� ǉs^F���0yBuB�Ϙq�<�'�G�7�Y7@Q�:di�eG�o�<�g�$6^���S���*l2�P�a�h�<y�jX�!)5��T&d:�0�(�d�<9W	��?=��	dmZ:��#Ą�`�<��j.
Q|�r�j�&�tAh\\�<���R�G*p��CA�%bxm��"Tn�<� �G#o��5c� ���59���s�<�Ш
.S�� &�9.���Fn�<p��+-8�@�Q	�ƨ�^�<�F��zO��:��ܤ9�%
Ċ�T�<�`�]1?b���v�O%u;&m�EUS�<Q5b�\^�Z�Bׇ0�~�C! RS�<� ���%N�	Mv%�T�	9��<�%"O����K�g[ m���C��!�"OB�2�.�#uBԥ*q�Q�f��"O���F��7]_l�S��q�"O� IT'��H��c��*^����a"O��8W�V�w��� e�Z�a:����"O�s4��$��b�
�Z&���"Oz�r�dGh�~�S��R�	�q��"O����`��=�iSp�з%����"O��#��(MlxQlӄ7�&4"�"O޵0eFдRDH�+��r_�(k"O�@9�'Θe�>1��")vPu�'�J�x�����O�'���Z�'l���d&�3d�j)�N&���"�'mT13��-��UH��#�HX	�'�Թ@ǥ}r�q�e���^Mb
�'|>�2d+��Q���A��=���S	�'ʂ,�a ՃW�85yGK�0��ձ	�'�����g�K,��A�/��"�y �'� p�2�B�uU��ꕋ)6nI��'F��5F�� C Ihv�K���'wbXy���Gn�!��ˆs��=�	�'~�@�׃�9t�Z��� �$�}��'� ��-R.(��A�;涨��'�$�p�Ñ'2$8(��.�=Fq�Us�'�ҠPflٳ\��av� /�Ru��'�<EIUNX�v��h5�����B�'��W'jR����膐s<�`�'�(�Os*)�%�O.or!Q�'gfR�FYad�b���d ���'8�F��z�.��V|����'5����n� |y^���.[�@��,��'_�ի���4J���$,x�2
�'��  �,�HH�2�X!#Xՙ
�'`�IJ��^X��s�L[3M\ �
�'\���jY�i��8B��?�R��'k�9�7D�bƌJB"ĵ1��x[�'�H��]�u�N�2�W�y��j�'7(��s����Z�`��"m�����'�aZ���8#x���cGf
�'���ᖡ�9p�x��lڰ�b�ȓBG�\A���5h�Dɣ�b3q�ȑ���8�A���t��x�"�-Nfz}�ȓjN�%���+p�L�5��5z��ATȔ{r��	uӮH�#([�6RD��ȓM|�e�ġt:�8
&�Y򈥄�K�:0��ϸY^���Vv@Q��g6L����8�bl1"M� L����ȓpU$,���H6����h<!��ȓϘ	R��?��җh��!�P@��*+D	�Ծ`g��Z�g�3ck�)�ȓf�`:fe����O%k{x��5���!��.��M	�:A�H���F!��ǭH̔���)	�6GBԇ�E��4���3B��P�ѥ2�$���|���:��  Q�0��J 2�H���^�ܱ�I
+x��i1�E�gz$o�a(<�`�1x53�+���PӅ�S؞P�=�'E����K�z�0�ӣ��D�<Itm�{����ř*S��0rN�i�<iB�`:x0�E��Lk� �t��d�<	��0l�d�9chH�ޤ2��K]�<��ƥjZ"q��Ɯ�J٦8�f(X���"�O����>L;��I�N1�2"O� 
x��oܤNPL�r� p�����w�O�z8jo�+Nf���"���C=�1�'����Q6y�E!"J�+H�d��.O,�=�O��'l>�+�G�'���� �r��H@�'��Hh�B�+Y�H���b,��A�'��l��g�RQ��]?ֈ9�'iV��e��,4�J!c;[<qC�'a�ս"��ؒE��uؔ��ĢJ��p>�M<	"j
	�B�"U0;|�!
��Vj�<��ɁZe��$G�B�@�3��i�<�w뒠^�(�3���&���#��f?�G����'<T�	�]��(
�����
�~��nQ�9���8U�%��Abڡ�>�%�)�I�hdxp���7�i����!���8\<�0V
[S ��2��	:>B!��13X6M	�!�l�Z���텻}!�$*<���� KCOl��,Ω?�a|�|�DX"\�l�s�Ço�=���W �M;�'��Ѓ�S��ՃcF�k�@���'����h����鱢��]DF(�'ǚ0���>@��q�A��B����'�j��6Gt�Ш���8U ���'�2hy3h=�r���Z�b�(�Q�'ex�!B���D-dяT4Vz�Z�OP��dՁ`L�5E� �}d�#�(�8��v
O���3hY�`}$��!��y�-���'���\q��v�\�f����!�<D������?���y�Bäa]��6D��Y�E�j A��y�TР��5D�\��.��Z�JN��8��fL?D�� +P�8Ƞ�Si�=L D�J �?�O&|�Q��9]��s%
v�Ɂ�'S ��C�X��؀"�(�s��2n~�C�	.G�*��G�#�
�� ���0���$Ie�'� �B{U���3��O�&���'��6+�	�(����WiJ�rpfJ,B�PB��G{���"ZB����&���8`s[*.���?��Q�!PeȈ����
3HƷ#��ȇ�_�!�4�:i��e�ef��[6*A�ȓ��4M��-!#�Z�Bh��?�����8>܉o�8={t ��)� B�f^���e��#�J��R�y�B�{'��Q�0V���'�D�">	�{"�~Br�ByT(@��iݢ�kF�U[�<A��H�T�����ב<���(���S�<O�`T:���B�)0�X�pS�X�<�I	�,i�ScJ+�ph����<q���hO>u�q@	Ef鈓���He���*D�����J 3֘$�`Q�I�2K*��G��H��m�4��q(�ܴ~��5!�A)}�)��$:�P�+I�������цB�I
/�Ĉ�Db�'6Qf%H��X�i�B��!a���%�Y��#��}���k�� R�Z��Y2� �6Mj)r�5D��	Gȃ#� �2� (/)@t�-D�p��w*�v`jxB$��Bl�:�=E�ܴ!x���7酣��p:�q;$�O��=�|:�4~ݜu��	z0dlj��@����'��~��O�;�8}[�j�I�=1��y��d�>���S�g�ي�e5*`�qcE9Q �~�V��q���8S�
p�v����v�3��1D��d�ɻ�x(e J�}#bH#�/��ȟ��� %.�@��UM�*s�U
R"O����Z����@��5�� �$7�S��ހ ���rlB4S�����ۈ����"O$)DI ��J$��:xPM��	ux�|9�(H�&��l��t32 1D�hQ�H��c��	  fؤU�,	@��/����%2����r&�ݪr�ld�@"O�)�mV`H�e��V�t�#�?O��=E�4`��W�=��ۻQ�n��Ԋǎ�O��=�O"1���(t6<��ģ���\���'6ꠣd�E�,�B���;w~��'�\} ��E�'�0�P�H4RH�	�'W�����§C���0 H��~`/ؼ�E{���iE��Ǭ�H�©Ȳ͋�u�:8��'� ��fi�!�r1Y�DpJ�R�Ovi���=D�Dp{3�"<�tNځ����9�DԱN���	�i�t�"�T�(R�!��A8'f�#&	u�6|:�H�h�!�D��H�0������!8Od!�d�S�z=�Qh�6c���!Y�8�!�N��J�P�(�TK�=���C�i�!�$ٮh$���"�O�E:x�)�@t!�䐍�P��k�:u,�AgI�}c!�dR�0��{�f�b����%)��s���4��d�'��[�.��\(pǈ�981���(�S���q��u�q�M�VК����y��,�rS��¤(�o֯�M��}�=O?7-%� ajb�1�zR���!��!N0p����a��}Ӷh�%�!�dS#~����/�PO�h�' �e�!�d5��XT�;o?����T*e�!�$[�j�\b�+��Y!Z��lM#�!�@Vr�͆z�03C��.	Q!��P�E|ur���������՛��)���x�B�S����N��<n�!�M,D�0�bG@*4ͼP$�߾]#Rm��*�>���3��j�$�9o��˴���Gj���3��rT�V�0H�g�3'�]��?K�y�AA�&�R4���'fb<��Z%��e��LT�=�4A
�1�h��;*V�JS�4g�j��S�" ��'�����pE;�@�_At�u銠!"�C�	%j�r�H.Ș(6P�j�g�'HO�C�I�r�$������9r���+�$Ϣ�>��8�h&���K��x�@�_��O.��d�G�P��)۱!�a�&������N�Q�������C�<S��P(��;W��d��EྌI���>�)��Q�8$� '��F{�����K�J�Т��z,�7 ��y�n�5lJ嫶f�z���M��=�S�O��u��l��)��UlY`��'p�$�1`11�ɓ�ia����y2�'o$H�f�3h�����05�|���'�z��C��J�RE0��>�2mY�'�t�B��[B
AiG��=�yb�)�S�2���Q��u*w�b1�B�	(s���
�������ɏ(��B�	3a�N�HV�����A ��1N�^B�7g_R���Q+=fl	rC6�:B�	�"��Rfm�R�cM�$92�C�I�����F�f�0� �����B��!w����,V8�R�XF��6
lB䉌?VVa�w&N�}��A8���zjB��6WT(`��2K�jbll B��j�b�`�����H�0.��k��C��*���$˓RP
���	#i;�`���� nQY�!�+��)`��A!}Ð�H�"O6Ps�$�FO��A7a�[��ty�"OxB���V���a���̔��"O�ӵdժr`0�9�$<@"O�C�F�:Wp�)v�]�M�"O�1"ȏ�f7hh #H#)��	�"O��˱m:d��1Ѷdԛ	)�"O��x����V���C�P>]_ �@r"O�h��#ղ%kzM ���i��"O�I��(��_ʪmk�� �\�y�"O����d��B3|�
�'R%	bDa�"OJ�)DA�c7"js�$G:��"OTY��?�x�W˦&76��S"O6�bb�UN�Y��I�x��"O"T!d!�u_�قq���d7p�X&"O���v��@�$<���@#|��"O��e/�;A �y��G�?y���E"O}� ђJ�]R1&�G���&"O:����X}8��qd[7v���"O>T)�k�R©����+*��L
'"O�aJ����A�	0"�^�4�k�"O4�I�c�n� ��_�_PZ$�f"Oz�sR�U3M8XIc��d:,���"O6�q���c��SEf(��"Ob|�FI�4L����$���j�"O���aJ)<������<p� ���"O�XS���0�zP���p$@�"O`]ۥj�;�r�L��uŘ���"O�)ae��b],�V���{����"O,q�#)��w�ni@ֈ��5���s7"O2AX��^�^���A^��1��"O�jA�ՈB5ʵq�	LbDf���"O��+ �$a�nY{�W#��:�"O�<1â�HF�b�m҅gd���"O|4aV��1XMP4�VW��t)R"OT�x6�>O���0B)�:�D���"O2�"�oL�B�Q<C�
)�ܙ'q��D�3_�T���"H��P&�W4�yb�0#�~d��N��y��ygR��yB�SN��G�6f����R��y�oU�%�>ɦ	[7H8��IW��yR%�q�"E�Tb�9O��%Cbb��y��,yx^�&J�ļ����y2�_�]OB��) �K���UB���yoƫ	r�� 6iM�L��z�@��y���oP�	觉_��� ��%�=�y����Aǲd:�`ۖ��a�D��y��?��{B� ,�� ��yR��2N����� }�*a0�	��y2H�/���!ADT�\����" $�y"�Z�`L �)T�\�_t�������y�f+9�Вs�E�����)�yҀ�<�⁹����,������y�Ŋ�Z��XGɛ�-�ZycB���y"��N��Eq��%�$�i"����yo�"������R�`R"���P�y�-���ЭH<~]p��̏�y�F�9fÖ���iȖ�Lp��$�yB���7���l2�~�`M*�y��B�L�<a1���ph�`(��y���Up�a��Վ��p���J#�y��e˺ՙ��>=��ږ�ߦ�y��f� �
!�7 ��IC���yb��T8�p�%S*�>�r�D�6�y
� �I���<���C���%"�"OtȲ�P�f`̸���q���`�"O>y(G�'��1���*}̐{ "O�eQcm�)���Y�W��W"O��[��Q�u����&Y�X�i`"Oڰ�S�1K���@eآh�`�"O�����9B<�̃�M�d�rp�"O�����64q�����Q��@��"O��[5]�D0:���(7aI��"Ol�l@�k��B ��.eJȩ�"O�0�a�S����o�0@�dQ "O�m@��)���B��K.&�[�"O�S��\*�yP�a.8i��"O��S&�TV����B��]5��)�"OΡ�å��wE����7P^2� �"O�h;@�%^�܉��]�bG����"Oh�Ç+�Y�R����c/d�c "O`�;���*�� D�-1uZ�"O|IK��pK������$9�d�"OH�*C��=p~�I�Z�#�d�&"O2q	��+�8k�J0G�(j"O�La"T'�|T@���� P��"O�A��Ɍj����kW'�Z�@@"O>����;���i��^H�"O&�"��y@JЫM�?U�(8�v"O����D#�m�C�ˊ"u�A{@"O�a����;!W�~Y8���"O����A�n~�8�!�I�G� R"O��ʓM�f��HHu�bL�b"O������n�6 �_(C� �� "Oƅ��*K�r�0M�U�n����"OT����_Y`PG�'���:�"O�8Js�X#�ι)eۑ��1�"O@�酀%V|�f�59�8 [F"OV�3���D4	���$�ı@��IeZR�#��S�Q��(с��0y���G��j�B�I q�]��U�%?ޝIB=]���Qg�4	MT�&�"~���H�4B�.2I�2Ǖ�R�ȓ6`\���.S�|�3�׀T�J���%d��
E΁�<ba{2#M�U�(e�H��=�f(i�[�ʰ=��gP!�\�4��ڦ�p�E�I������J�W/��7�0D���b-]�s�P٧�"������+�I�J@�Q en�X�G��cW��ظӊQ8W���pq���y2&!
҅b�MM�M� Q�U☪k6�xR�ܪe��ʓb�V�|�'^��JU�@�	����-��_�^T�����V�"}�a��qsPѺ�	�N`��@bBdBJ���m�t����'�~�P�� n�����܈P���I���s��ԟ��2C�V�<�b�����4	��a*�*u��O¨���'�FThя��8�PQJ]�*M�La�O0m��ջR����q1C�<i��~�ҧE�]]���k�
�TI���Y��4���=)���ɾU��H��3r�L����Y#?Q��k%(�t~��r���J�5�����>Z�jQh�8��XR��Q>�B%�~�\�'
݅F谉R�T �h�W-;r����$(6.0���*�E�~ě��~+4�D�;)�lUJ�{����Aφ�x�`�	3|�A���[^\=�D��,B0��aX	N�"~�	�>>$���j��wخ`2�� ��I��U�tƑ D��=��l�SфE#?��M��0ev�8z��'L\<��n�<�T��ɘ�^Yi�G��z�(��
9H|���dD�<�9��x`Z�r$ҋjEK4醆:6������'�y� �1��L0�O1���2QN���1���:1Λ�|
3#�2or)/��  A�!҃w�}1��ׅ,�t���J�)�mƭ%��ɵ��t٢bś��n�b�Y�_�V���'W�y:�-�m�g~��U�� ���������������O:tx�Hʓ^���I~Z��D�-]��Q"�KO6�9A.I6��ŀPL�s�f��� ��{�b�!���V.�ҩ�P�O
9� �5�~��O���G����q�:4�N���r�ޚ*�	vaOR��98�O��Y$�T�_EB��䏽K~�;a�>!�퉝��h���:�V�r��(Cۚ��W�Hr"���?~*q9�!Z"�|@����6'���D�&i����`�5A�� �G,N�:�������OLdcT�̠y��,����-m��q�t��4��'���y?����,L
v s���0A:�>��]L�ڌXW� ��� nH��+70�]`���2Ck�+` ���
Ds���9��1O`�� l�rѐј"ΜA�8b�Oʀ��Gt���H��)'�Y*���q! p�t��Pl±��|��B�p߄ �e�j�.S	�'5�,�q�=t|��3��j��1M�|S_����a��U;��ъɼvx��v.�l��9�OFj	���ģtLr=S��E7(�p
�L��:M+6�FT�H޲�B4I�,Ѭjޑ2��Ek������$�ٚ������'��	!ꖥ��B6��#.I=G&�?Q�bO�c6
c��KƤŬ	hNi+���D�8Y� �DOPԢ �4g�j	��
w
$���I9f�P�����/A�Iٱ&���>���H/C�U�!f�z�.�SֈՈ>1$�p�R(ho�#A#0�N���'��p�bIB�� �U���d�PM���֝b�4�C0E�70̬p�吮����V��R�[�$A�\k�nV$ؤ�K�<�Ԁ��`�\1j��6G�]�d�U�O	���d��m{��K5T��� �?b�T9b.���/dφ���-������H\8k��/�����ܸ��ɄdJT�(��jXIG��8��DP��P�p$9�Uu֘��$D$ˎ�f�
�MN�iU
_x�'OF�)�J�~JL�'4<!A'U(~q�1)��a��̨��� i������rFF��F8�p��	=�� ;vX&5t pD#�6}�Mm�d��ho?��'���� 9�t�&�
�=Dir�e�hu�̑PO� S!�Urf 7.܌!9����iC3BMI��F��@IA�&�9�\:�KD�m"b �
���N����#o%v(`2J_/����B��(ѧS6.4
9��M�	b�C�	��H��s�S�Y`���+$ܒO��BX.,аى�i�2~Xq�6�MjtX��̞b[!�d^-���+Gm!��1J�d��bp+�a�D�V� �?�'��y'IB0O�E��$$dπE��'P"�a��k��aÍ��+��8e$�&����'{�x3�FK�~~��#F��$��	�.�C!'?9#��=j����@ȕG�u��O�<I��$}#��Zny�X���K�<���ޔS��HА�6)�ժ�*�y�<y�M�;T��xS��`Sȱ��jo�<ҋ4d��%���[ 9l�sB�Q�<y���H�&�3@�!jC�H�<yV��a��);��&tTZpYN�'n��c��R�g��mc��($tP�WdZ=m�ȓ@�|�3��[�s@�a��=" D8�'���+�	
]�a�)�g~@N�g'�сdBR��~b�����x��]L,-ۓz��ݣ���#W�Y�$a@8�W��i�"�!b�'՜�pQ�a��)S��Z�\/��R
ϓ`�����O��bҍNB����,dw���T��:��\ra��+�x���#�X�w�~�� 3�_��y��xC+�O�(��D"|P����bE1G�0�Xwd����3HM��y��ya�ʀs��y��ا9ԠM����O�g�^�}��i�3M��Op�	���g�d5� 
_4F�X�B=4�(��I�7i6��*0Cºh�z|��k�^�j`�F�'1.��V,�n��Ą�����.�vX�fm�:J�x����u8��%a:�p���L�:0Z��+���Xb�"��Od�D��hq�MsU� �|D6"0�	6O1Le�f��5Vt1�8 ����!M,�9H,;����"OX��g؆=���f�@�:�BذfP��Qt�U�1 ��%�"}Z���;��U{1��j�60S��Tf�<���2X�d�[D��P\p(�t��y�I�Q^t �d�'�5[w/�H,�$k���L<��	�'qvU��ŝ�"Q�,��N�5��H
�'�E��EWz�kd���	4q2	�'n����ޚ9l$�BFM�+m*��'�x�� ͂4O����"�95"Ts��� P���su�8ؠ	ڈkN=  "O@tv��3/]��SF()����b"O��1�^���1iP�0�C�"O �(d��`��tbC�I�/�ĕ@E"O�8�GƔf݆�R�˞Vے�y"O6 �"�"jhX����,�>$�d"O��5㏶�L��C����x�x�"OB�(� �a�[D->v;(��S"OLH1��>R�h��L\1����"O$�q�)� ��XGJ[&Aʄ
�"OT���O�1>��xƩ�x�ؗ"O�HS�@@�pRP8!� �	o�xʷ"O�$��(� �:�#ń5+N�!q%"O\��gcV=*O�����_+Q"�M�c"O4 $�N�(�U�&D:b+�찆"O"��^�9����7}-05"�31�!�D�(0��Qʀ"�:| �($��x�!�D�$�h�C���J������?FV!�$�1SE�X��Le���#A�F�]�!�d����DeK�s�4���T8)K!��{:<Ź��О��Q�D
�yS!��C��Z@�A��� ej�0�!�Lc`8ap�.�
U&�db@��4 �!�D�2a�P���HR*S��}��(ʣC0!�D��A��ԡ��}�v�
S�T�#"!��R	�|��	_:�p2��U2g!�D�+BL��jթҬ,a��	��P�!��IW�-2����gg.�+�/��_!�d/JH�"��?MC���TN5-:!�D4;�8�e�@6�)�n"'H!��[��`-�l�ڑ� F�r�!�<t�l�Š�"=f�y��I�!�+�2��G��/g*�SW#��=�!�D�p�^@���[,
X�kS�BU!���'f:y��	��B�(��%:6!���L�8\��SB�!�5�	y*!��
�S!��JDA��9�@�s�E̟%!�d�1���!8�x09���t'!�Ă�wN.�z��� �����PyүI!{����ņAHbX2S м�y��$[:a�f�RR#b���yR��lJ�R��P�(Yp����yb�F�&
t�KP�K�Ls���,L��y�E�cuܐ��<wEZ���b�;�yRe	_� y�'�&�$�8ǈ���y2ȋ�{vh����\�
h1 Ƭ��y�L�;��Tre��>k�v����	�yr��cZT=+�Mոbb�4�1��<�yb	�/�tB���;41L\j"�)�y��&�v%��!�y����L��yB��&C_2H�&��CU����y"GE�Ks����Êg�<m ��ܤ�yR��:Z6	�k$�B�B�)��y�O�z�@�kΔ{<�h�#h���y��|@��!B	j��|�B��4�yr(�.kx�`M��D��!�<�y���r�L<�����$�a�4Hδ�yҮ�(�T=��I���Q��kׄ�y�aQ�tx��V0�T�A���y��Z�$d�/ {
�4�ʐ��y"�\���إdн#@LCᥟ4�y�,ݛ:/�4|=Ь�dK�j ���l�j��L�F<A��_�)�!�ȓ/�Z�@���1F�P��	J����S�? p�"�]��&�N�23�<	3"O�2%��:.!��z�gU�~%�Y�"O�L�DCO!>|�ۡH�m��M(�"O4�Q/̎n�Ԁ�D�ːmLrp�"O�8��˒?I6�A��8؈��"O<�� ��v��ŚS��N'�82p"O��)@#S�2�Z�KL���Jv"OԌ�s�S�u�2��`6o�t��7"O�B'ʑ=�X���+P���D"O�`�'%��W�8�i`�
��|*�"O�!��ͮZ������Q�p|��"O\�!��PBȌ����G�lXZ�"OF���P9b]�ĢT,�c���"O0��V(	�b6�a���:���`Q"O�ق�P:[GnuB"�0b�h0�"O��᳤�So6�3G#M8Z��࣒"OR�K��G:S�B�����sǔQC�"O
�ۅG�Y���Q�ѱ/�$7"O��㗭ʹ4!���	"u�^5x�"O�q�rEγ:�b��FG�=qe��a"Ol���� �>�X:Æ]�|tT�j�"O,t�u�r����d��.�$P1�"ORdk�gI�8W4�B�fT�(p���"OvD8a L�4�,�%�Q�옫5"O����$�~�a�5g�h�:�"O��`�͂gߐ�W�.~��$"OH���,����5�Ci�� ��"O� ��<�����R<	�u�"O� /�8n�`jUf�)��ms�"OXD�n�;��m����=ބ1�"Oެ;t�Q�PP��w��5�@�і"O^@`�1N�p�rP�H.�a�"O2-�Y�xJ��bO�7��R�"O"�9���a��En]�!L��j�"O�� SeŒJ�v�i�ā(+~e�"O�$g�S�u�>q9�i/�`@A�"O2���LXH|��!ɕ;��c�"O����F�8 �����b�b�2"OP�ă@;rʤ����9Z�j��� M�T����bj��k�IB�qX�$��ꂮúB�I�n
���ͣS���Ŋ^,ZM���&  �+;�8&�"~�w�r0����2��i�E#y�N�ȓAr �j6��Q?r�ys�@�U�>����g&V, ��W�6�a{�#�%P�����/�)H��P$�����=	���x��B�Φu)��9��!�+^��h �'Ĺ�yR	��DĠ��hUډ�G�L�'�@� 惷L��9� ��	ɴ	GŲ>Y��+qI��z�XC�I"-�ׅqIP��+)���qr=|W�5/O�����Y�4�1��]��(���8:��sD+=D�d
ӈK*&�䂖d��=�vD]�1������M-nCİ	ۓ����iH�
�⹢h�F�m��I2z��1���x�2Ho��t#��J��;s^H�B�l\�C�I&X��т�E�j<�A�1���qO�� �B�\�<�"&�6ҧ��C��"��䠞�7�p��pU�h���)|	"�i�*<~�2A�E	�����O�u��Y�Т���8�Hi!.˂uY�� �d"D� ����ci��#LJu�h���"�D�	�&J�2����d��0�ȤKB��QN�)�b�Ra{Rcʈ0 T|`��O��Yш9yX�[t�_$l� ��"O`,s�"ۤZi@1���K�n�h���^-���P����8.��Y"��D� ��CN�Z!�d˅��M�p��t��P� �F&K!��w��lA!��?R���F^!�$S�L�R�A�ۦV��U�D'�0]J�'��]�dg�pX�� ��('EϪs �i�a/��FW����'�ܣzJJ�pQ��%$�aKF�Dv|���
O�z��E%}�l�#�'��+�$!�ɪfRH���=#1��1c�)Q�p�j���ƃ0��9D"O$���ªEa�Pu�3<��t�OR=:S��6����L��}z�̮��,��M=�QA�M�X�<!�ƥF�A�C�>ԉ��^Y��'jMȳg���0<9�	G�[���Sׁ4S�T�F)|��Xbs���ʸ8` �w\#eM)B�1���M
!��ͮk��0�'�!��*����6�Q����uv� ��� F��jJ�ۤP��l��"q!��J�sZ`�Hq��%���Jӊ�)���E�P.D�NW���)�'nI$�� �,���z@A �D��!��"af��g�N��:�Mг=��O:$X[!d}�u�	ÓY�܀r��
�jK� "���Lyt����.���)Uʉ�T��4Ƀ�ǎ2�Z U��������@�l=��A�>1pʁcޅD�DAL ��~J�,j��QA�
�uж+6�D�<a�hRvx�łY*0��(��et�<1��L�x��䧁�%ေ#b��s�<��	�bwJ����)D{�t˵-��i�ą�=Ѷ�7�gy��Q T���Q���AǶ`� �[��y��[�;�u���Gw@�Q�gS��Փ�Yh�}�ȋ�}�J��UB_�F
�y��W��<�u�� E�Q�Ʒ>q�&��m�z���/FG�4�y�C�<1��١�8��mY�M)�)a���ey5)� 8�?�`G눤0���ɉ�&x�m.D�J��&0����sk��1KD�(⪋�b��uK���!�TT�g�d�yJhb�c�l�T)�Һ>,���G�}��'\
!왠�N�"Q�j�Ah�*�1�(�O�Xhd�����ӯO1��Hr�'���/N2��@�'캨2�	ʥ[U�P�S�F�Gd�$��'��w��W�(K�I�=�F��K>YS@I�8�R���1�'|i��a�	-
����*�ْҬ/D�Tth�1'N����ǍLt`�ѧ��B��{J���Bc�l�g�dfG��� �\;M��UK��APZ!���<���cQ��P֜����mA�����Y=����R�	�hYXUGV�f����Q%/[�z$D��$�'�X�Q C�Q��R �JА0�	�'p���A�
�Dx����ftC	�'�,J�&=���i��V�����	�'d�8��ˍ.y8�D�UF�y?�Li�'�T��튓�  ȖF�4X��'�~�')G��T��2��tٖ��'9tj 'ܘpڋgH���O�
������OB�@a��&r����kˋ��s�'r�� �T#wu�$���݅3��I��O��S�A��,�O�>�S!"6�p��7��--� ���,D�L�T�ڭ)�5�Y.�`��Ԫ+}+�_DݲS�W�8�� �'6,�{$��|W���)�Oz�Bb,R�6q)w��_"P` K�� �ڱ���x�D��j��y��Ɋ�f-0���O0��&�M�a���(��To�*�Tt� �kh�U계���y���h���Սd��u��0�~b��Z�ps�h�n�퓂+��I��7 7 �
�放kV�B��.-j�
#�ˠ{p��1L����'���e(NY��ɦZpt,�V�3FU�,�U��#�����	&�~��F��ed��9��^
)�dl��ʄgX�H�'Wqb���O���0q+3~�|���d��t�6����X���O���)d��	*9:1�ʹt�jЁ�'i�tp�׀[��(�p�[�nq���O�R�呇I�ȒO�>A{�(�%���a"��G�nQQ�e?D�x�E�Îy����C��Z9"�E;�d���^1*
˓aN���חb�|!�#إx�Ҕ��S�? ��JI�G�ժ@�R;
Uq"O��s	��g���&�ݦ4�� ɦ"O��� ���{a݃,�h�
p"Oz؂D�܏Q�,dZF��usHPSf"OPY��ͱ�2Ǩy���"O.y�d�ۛs)�|��C�� 1sQ"O����ʝ(&Z�HcbO1
݌�5"O�Q1P�lR4�G���,բa	e"O���h�=��G ѕN��䢲"O��
�pi�!��!#��s7"O���fh��hƔyS��"+�F�6"O�T�1���2"T�c��8[&x�8�"O\]�RF%S� [�Q�B����"O��� ��B��pS���	_B��"OL �6��$-<�c��4�f��G"O��6�D,;'�ċa�¯C~B��V"O�!p"�]:;���K�YkH�[�"O������GPp��-�QQ,,5"O ���K��P-�g�Ϟd@V�h�"O IA+Z�1kp��� !��U"O��b���?��՚S囀m�TĐ�"OD�+�/��Pf(��b�E龵��"OR���I�M�B|pӁ�"��"O ��C$�):�x5oZ'h�H�"OH�+��/'�hb�>$le`�"O�1�ՉZP2�p�T-��%(t=3�"O�=ۤ @�� ��֫O̰�"O:��T$B /`D%z"bQ��:�"O��c��M.Խ�B���� �"O�Q3�m�5M4%ȠKS�y;�s�"O� r��>]/���I�)�`Ȳ"O�A�ŋF8���W��:��"O�" ��5N�H�@��=w�T�"O:�Ж&.E�X7�Q�D҂"b�3D��1�[�,�|I����.��iY�'\����^��z�E��0|" C�;�ݸd��&�u(��1Vx��'��0�eτ-C����	���𠸧k�*]M1%d�E�b��{�ĭ��e��SC��XD�O�$�	F�[�P}��	Y���ـ�4<�
qC�bC2%C�T�<E��%�.n#F�����" �D��Q�ɿ^�����>,
�md��#	�'y��� `釱�&�p��	��,�w�_��|��'~L�uF!�R�S�D
B�ӄ$ߪ50\kRQ*-�!B� ��<Q� �5&4���>�D��%�;	I��	�OƓ`ЊE nd�����0�f8��"�����~"gF�gN1�7�!qev@s�S=ordPQa�T�|R2GFG�gL���̺��_3ۤ|�Q�\��4������9�m���ȡÐ;O��~�L?I�u��*+�zњ���+w�~���ƄYv�����W-y��ר�h��i�n� 0��g�V�5�8<�$�&�@��y2ME�P��Չ�S>qG���A$7�|X����a�&�H�%��;@z��j�\�VO$[�\�	�'C����v�]�4Xl�za)|3l!�=ތ��&˭\..�c��Vr}��)ЯT���V�I�Ġ@޴]��䌼a���HiL
��I�5�)%�	�{HFI��`J�|�!`���H<RD��D�4o҇Y��~
ç!��Q[Q�W� �Q��2
P")Y5�~�� !��T� �"���r�],�8���\�;��J�']���IciR}y�83a��ދhqz����	X�Ĝ���Z�����G�?��D��o��^	�������`����bX!u
��G�T=[ V�x8�ƕR�}q�i�3q�>ŉ�'f�Pd0 �c���;ċ̾<ziv+�1��8��I<C��6�/�(�z�/�X�Q3"ES��]�5a^h����E�5"P�9E鸟�R�$��se�����iuC\�K��y�p���W�ޤ��'�Y���[��O�1��٫�X���D�A��Wvl%��'P���"����s����)��[6(Ԡ�Ϸ9�j0!w�"fb�B�IH����ע{6�]a2(Õ<�B䉆+�.-���Q>4����wa��H�C䉅�� ����m�zt�b��Y@�C�	�+@:�*60������6K��C䉈wͮ����g�2T��5y��B�)� \�a� �Bx�`��@�;�T�J5"OZ�Cq�IJ��a`Iy���J�"O
u;v��S�&�H�����-sS"O� G`��W�Z�Qt�i��b"O�93�_2˅ 2f�Xr�۵w!�Dյh0<hE�Іs9�����!��-��\�n��*U�� �� Y�!�$B��t���(�2��ܴ`g!��=b�0Ak�	'l l@���76�!�d�7��t+`,�)����6�ʿU�!�$GBx#�f�#4���v�_<�!��y��ǡw
�ȑ�&��h�!򤀚PR�UIQ��*$Z�z��M��!��0V}������#"���$ț�UY!�d�-a���f*Ȯo/P��U�SS!�$60m|�l�Y&ډ���m�!���FhA� �{�%�s���J#!�$�T��E�a$G�3hl�Iٮp�!�$��-%����6L�F+��N�!��ة-7�-�bX�\�d�SIƀ7�!�$�)F���(ٍ�
,(2g�;�!�d��;�pX�@͞�S=�jb�ٿ[-!�$ý=�ŋ!*B�E�4�;�!3�!�$�7p:t�Aw�V?q�i�uA��Bo!����h��㙰!�H�s�J/e�!��<<�#���pn��"@�,$!�P$Jx�H���7DP8E�c�S)c�!�$��F�P슉'5t q�i��~�!��N�>��
�2����h�]N!�D_�+3��ÄŚ�P�,��5G%,�!�d֒u�^�@OϾ'�l�BR� �!�2��I9c)N�BƲ�'��!�K�<@Y`�ձ���!�!򤈑�8$�B�2�j�b����R�!�D��?�BA�`��)U+�c!�W�dvL����M�⤴z�CM�H2!��"}!B�2��³�*� 4�]�f%!�D�",>(xT�ª#.���)!��_��z��N�*NȀ'aM7!����s"OF�	�ɐ�ܟz�!��<�$�k� ���u���ę$8!��T�4k&]�g� (�t��#�/W!���r�h�̷f{����ǖ�!�A�q`%�$eTt����?�!�dH��|\��E��f�@��F�	f�!�K 'X������%&ar!��²'�xI��ڸ�<��vB�YX!�$G50�q�&n���Q���*!�!�Ď�5Ӝ�w.�-��$���B�)r!�ď�����%�P�����+}0�14"Op������\SNx��I�#bH��W"Od� �t9�!�B	-M�$�1"O�	����P����BbǰQ�"ݳp"O���e���k!�Q@��j,u��"O^1C�ɳt�2��3L6{[J�I"O�5q�#�d��\P0��yY�xS"O��F��Y��)e.�-9��#�"O��ié�W�\ ���ߞt����"O�h���ΐv�r���M�%f�0
q"O��ԳR�
� ����H�U`"ON@���0x��gG���5"Or���G?_\�rV�J�Dڔ9;�"O�P�S�V�3��ـ�C1 ��Ƀt"OZ�2u��#|�l��+ -G昀"O� *�t�G7��u-Q�RBL 3�"O�,��n��{����3>B��b�"O���Gc3��e��ݬ�
�p�"O�p�8�j�blӿ����2"O:�!ų Sv�@�;m�J�"O�x D��k[*Lk&��,kGPl�3"O�m#�'�P<�-S4�81)�]�"O|Ĉg�P��<�fH);�:e�"Oi�N�-v�H�rƂ�%W�0"Om�TE]�PK�+�S`�c�"O�����˯��Q�JtL�<��"O�,i�N�3 ����"TEC�M��"Oڱ�E�G�P��\Is"�w#��(A"O�%L��bސm�E�� pJ��b"O�P@�h��HP�hݫ����"O �x��<f�1q�M��[a�iB�"O�1P ��-����b�~�4���"O0��5c
1���qB� ���Q�"O*�`Gݻt)"5����!�̀��"O�ev늌,~}����"���b"Oԙ�,ނ�a�a�z�8���"O
�HĆ��3�Z��K��\��4Ѕ"O,D!)�9i�`�f�$4S���4�y�F% �>Rk��C�̫�T�y�6�tD���w��y;����y2��'#Y��#c�� G�̀���ޏ�y�I3��@�$L�2�Ys�@��y��iɬ��G5z?Ԩ�I��y��#����f#�)H�����Y��y�lM�]Z�m�����2�y��]��X����*#� ��/�!�y��Zl
���hӳ"���t�T��yr�3b���Q��#!B¡HE,ˌ�y��ݽ� E
��j�� fO� �yj�!�9��|�v*�y2�K�}�ӑ�4GRyk��C��y��O"Y��X�ƀ�*}�ѓE�D�y�!�0BRaI����Q���4EP&�yR�yؑ O'%��%B�&Y<�y��	�{�t}��;T,������y��>n \c���j�E��o��y����p.6�"�Ύz����!�ݰ�y��3T3X�9S��qK���p���y�@|lF�2v*!��U��F��y�Z DՋ `� +�n1�)B"�y��L��$�����0�Ū�*T�y"�*�j5xPZ�|1v=�7�ʆ�y�@ލ4�ܬ;��H�";� 3���yRn�=QB�,���bU�B�ۨ�y�P�f����Ϛ#T�����yr��:V�4b�nCPP���7�<�y��ټf���Ha�"\��-h�!��yR�ĳ2����,ʊc��su��8�y��b����9Fw�) 2	A�y'M)2|IA��LA @����?�y��O8h/j�#���<Վ`�`ꃸ�yr��(��y��N2@���è_��yR��2Vt�6��#a�dqb�GT�yB	�!{��ԁU�Zn��󍔿�y��59s �a�$U�`X
m�yb�Ljl�8v��M�� ��
��yr��^�^|���1N&��`\$�y2�1����^�dQ��K��y�� V��O�5P���iD� �y
� ~%�d����Ɇ�G�Ԩ��"O�=��-O~qr�X�b��Aj�"O��yG)W 1�$�'��
C	�.�y�/L�'�ʜ:���,u�^T��5�y�f��R�x37*�
o�"����Š�y��J:5����dӴif8A����y���9R��  "m:_/�<)�U)�y�	8|)�q��$� ���A��y�G�j �PɥIC�(����� ���y���� #G.�Z<l!d�Ӵ>!򤅪��tA�.ZC�I,I�!�ˠ��bE���t!^�qr��9J�!�Ă+U�5���Dn"I�wo��@�!�d�G��#v�N
'u0BQ)�P�!�$�֐���x5��{��W�h�!��� QX#��������@`R!��Ȩ.Gz4��E�tl�e�c��'qF!�[r��Hh5�̋ e�8�H!�!�dY?v��dػJ؅r�&A7)!�ǣXvĺ�C <l�h�o�9!��E;+wְ����0eG-y�nɪWY!�D�800"eH��=Q�N�G!���a����t��1Qd�6�Ԫ!�!�$W%'���aj����x��Q3F1!���`�����F^�6�nH	���U(!��a��AS��'n���F&�?5!��ԬA�����E�L����d�T|F!��P�Ȝ*�K�Fȇ(u4!��t�
�3�H-8ۢ\I#�Q	n�!򄘰'�b����+�� .X J}!��5)LZ�ɀ�,�b	H�#��}@!��]Q>�I�!�5�4CE�t!�dҪ�")QƘ�[����fϐ3&!�D��zD� ����%����Va���!�DӳHy*�!���av<����p�!�d�!Y[d�@��W:����M�b�!���(��h����%m�:T���Y�!�dV�3"���Ɵn�p�:���:M�!��bcd1�&/@�{rN�ض�ޗC�!�@	ad��AU�@lp���>�!��J�=��cw�?&=l̪���`�!�-v���-����\�GG�!��&�PŐv͆�-�f��R,?�!�V�Jz�Ё�,�/�Z��ǔY�!�dj�@|�"h\!/��pj���'v!���	|��=���q�2�qq�5�!�DE&a]�\3�Գ~'��5%	�[�!�D�9v<�0UDdIJ��ÙN$��'WPT�%��27n����7Jr���'��QbD+_%S
��X��Ɂv�dJ�'Z�=;6�؂	y�@	g�;t�<�
�'��4#sFо5��,���Y����*
�']VE=X6�ٻ��-m�1��n1D������11!.5j��=E$D9X��.D�8j��p��\8�C��B����g(D����� ^2Y�%��_��Xb&D�|�W*��/N�@��O2�"L�D%D�x�!
iw�8�B�EҁY�(D�� f%�\�Kׄ^�9�A�8D��C.� {B<�X�o�l�VE9D�ty���"4���Ab"@fx�'�#D�t�`�M�=���3�@>v����%D�x�aHZ���E�'K�\��5D�P�r    ��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   ��   *  �  _  �  �+  �7  �B  eN  �Y  >d  9l  �x  ��  ;�  ��  ��  7�  {�  ��  ��  >�  ��  ��  `�  ��  ��  B�  ��  ��  i�  T�  ��  W	 � �! �- = G �N U J[ B^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�?��+�сg��:�h(+a��Un$��F� U��yz�rMY(P.؁�'2Q�@BۓRLx�b54�n��'�Л�O��@k�b�P4ir��g;D���HB �𸡆㎨5�6���:D�ĉv�%ΤqQ�-׻q�頑�$D����-:*��Yg�к/F�`BR!�II���'\+��0�e�=��d{f��S%��ȓnydP��La�Fe��6E����ȓ�u��
O* ��1��@��Z���z�	�F�^ #���L��"O˭o��x޴��?a0�W}����(Y�J�65	f\�<A��%9Љ(Q�ˋS�X��"�T[�<�/P�	U-zQ��'�>�J�,US��>`Dx��$�ߦr���(�Cu�ځ�yR/�2���"P��9s��i���\�y2�֓zwB#4��4�驴M��y�)��GX�@��9c�}z�2��#�O\������j��<P׊�$Jl k �'4���y�zm��f�"� ����ݼB��	t��JA�Ȋ5be��>[�>��U�"}�'�O�	/?o�*ny G²M#�)����9���D��/r���8zn���	J�2�qO��	8��D/�T?��ӊYʊ<yF�֤f~(�*�K"�dm�H��HAUĘ�^�nQ���Ή.�C��/�f]c`�?4LY�RoH�U=�C�)� ���iP�7�e�diE;٪̰�"O����m�$����>A�<	Y"O$}@'bU�TV�ȅ�ݠ?��m��"O�K�M|��	��P%.�y����f��i��ʍ��.F�:�<Q�����<��`5 ���N����z��:o����ej��4/M�t�4���� ox�<��	c�oPL�QgA&0RdIg�J̇ȓ��i��۵O��(s�\�9D'�r��X�S�'q����g�����dXU��ȓ0���1ed�xZجX�$�f����?	�BJo���I�12u�匔�cDԻq��XZ!�Y�� C�[$�LeH��� lH\����s�����J������ځnw��Z�,D���햨J��	�k���$xP%~� ���>2`$���f_>c�`��QGzB�~r�_.�����q�T� �v�<�NP+$����5��!E�\:%�s�<q�^C;x�ʠ�� }g�z�"�e�<9��]2��<�QDTLz�$ٖ�c?I�:�؈c��@*,���5�Ǣ`�~مȓ3�^��[48E��B'�ꐅȓǫ�b�ɾhE^�X�"ܱ�X��ȓl
Y��)Y��艈AD/y����ȓ>h9bWOQ�W*��n��_�@y���+�S���ٹ_s��AvK_{�D�e�\��y�i�7Ze������ i���U�A<^�Q?i(O?��?51Ȑո2�˷�U3W�����'�p�㣋7on�Y�g� �N=��3�yB',lOޥK�Kʊn��� �n�$��O��>/&1 F�:~�������v�!�$���|DCAj�(yq�4۔#VnџxG�k�O�0J%J,��X�N^��y���!�\�����hXW�T���"�S�O��Q��wp�tB�d�>��]��'��Ȣ	�uL0Q8�e�J���	�'�R����"Kp�% ��u����'����y*�;&.ֵs7�d+듹�󌱃��$S2��3w$4$e�#>���I��*����kGm\��V-X38+!��rH	��H0.l�ы�-5$+!�Ӿn|Ω��0\Q|x�-̝�!����*P�F��U��W��hʉ'gb�Γ[��xr	F�x�1�[%fc��h��,��d'O ��y���fh��D�
T��a:f�>)9n�M؟؃��E#�\�A��T����8�ə�HO��2�7@�r{��f+,r?`цȓ3��Y�«٬/SD���D1�Fz�'�0�Y�M#�骤��~8����'��U��@����P�fO5%���y��?lO��p�≒�TYJ%D.k�h@ "O����nL�>�0�kt��=-^!x�"Ot}Q�N�EYΩq �т'J����S�On�M���R	V$���v�ٷ����'�<�e��*; ��"�}��b�'e�#B���8:��"I�̉�'�
��� ��Bc
ι
p���y"�'`����1�6�bFP�
��	�'�*嚅.�K�b����8%����' L����Do��C�>�$�Q	�'�"!���*p��Y�/УF��ո�'9p���hT 5(���Ԧ�m]�q�	�'�(��(Ǟ��=%�j��0�	�'אYд.� "�Ԅ�kՖZ74 ��}���� ���ʟ-'~��{4эB�MCp�'�'fą� Cb�����&��b��	�'/�ծS-�&Y+R ׫`6) �4�Px�L+*��P�+��_�4�&)���=эyB�T�������mB����H�oDL�<���Od%�%���9�R�U1�2#�"OpXsD�A�41���޶lʑ"O�X�P,�����"ēc��Q�K4}��>%?)�<�_rƖ��4�A���X��''"4��Hլ0.�����}���m��I�O��IM̓ڸ'�,
)]�^l�U��87��3��y%ъk�h�q��� B��(RcK#-�qO^�GzJ|�u���D
V����B��=z'�Y�ȓ0�\5�I�H6 QB����\����'��x"E�Y&���F����X?�y��F���m����*ϴ,7F��yZy��[dԷ_�b �ƿBB�C�����͑�<8,ۆ���8��C�I�#�q�hʝ;�2��`�	>ϤC�I"I�H�ѶGƌD4��z�C�.{�C�/yQl�����s܊e�&jZ�C�Ɇ,�qG��'%XL�����0~C�ɇ��}�L=!���R���C�
1�䤁6+��O����"_45iz�'�ў�?������	M�1��$uTr���H7D���sח9��B��<*5�%1D��8���i��A��&�����)D��y%�����B�+Z�s����;D���Vŝ S)e�7I׆n�~L�a�:D��"�����b��3W�-b.�`:D�dB7� �9�5/�"3g�w�8D�09$䎐_R�w�K�(;C�*D��x�'���4�`�4>o�dR�'D�����6��RHR}-���*D�T���E �mYc�Z�:64L��n(D�����X2EQ8���N��b�ap�%D��;n^�>�s�=v���A��(D�x�E��?�X��E�V�'۸�pFj<D�(�F%�r�H�vē�H�~m�G�<D� {��D!��`�GǅJ(ZU�f�;D�\��+H�G0+�LFN�*�x �$D��q��T"J���E7���!D� Ac��.f���F)¥G��$��O+D�P� °i!���#�3.�<ɡ@*D�|q����
���pE9R�t�`&-D���d���Y���2�E� ����(D�0c��FE4\� A)C�Bs��SE$D��Ҿb�m
�a8QV�ɻh=�yl�Vz���ү�8�$�:��J��y�%Ya�Aq#���J��̍��y� F�ҴBVn��1�4� �nT��yrj҇U84-)��y�����y�Ɯc�l(ʀ�M�7V�=�+Π�yRN
-��qR׃�2�>��7f���y�ḭ{��X���0�t Q����yB��U`�!� zi��'C���ybm��z�����x�BL�3�6؆� �Qk��O���'ZD���ȓ �Z��NA�I%t��*�7�b�ȓEw�$��ڷQ����󃟇8\����n�ƕ���):hЁ��e��.��ȓ+W2����0ބ�d��4�2̄ȓ�����	�%24i''D�(B&���y-�����x��*�;k�Q��S�? ��TdM�+�=�BP�(����"OL�q�O7![��Ƈ�&FB��j�"OT�ؤ��yL����P5IU"O���1��-���C哒0�2��&"Ov)�U;�@��ݏ�J��U�'�B�'(b�'/��'���'`���U�nЬr`͛��шC��Y�K�՟��������ğ��I̟�����	��H�	99�(9�WeUa�`�R��ϟ��	��Iݟ$�I�h�	����T�#מ2=�T:t�X�I�^e�3hJ͟��	����D��������$�Iٟ|����N�r��sIα���Rş����	П��Iޟ��I韘�����W�@�v05$ڊQ�е1u�ܟ���ٟ���ȟ�I����	����֟l 7EA.Qq�@�j
03T fK���X�	Ο��I֟����� �I�l�I��K���-���0"I@E����W����Iџ��	����	����	ן����D��%�&Ex�8c���൓!�
��X��՟|����	�H���H����t	sM=fE6�cƈ��~��3������՟|�I͟P��џ �Iݟ������k��J�(*~ ��P;�:�C�$�����I����I���������˟��I���.8�г@&@=U��� �!��A��������I͟��	���������Iȟ��I�v��u��+U��h��R
�u4�$���0�	џ���㟜��ß ��4�?A�0Y����R�{��0��+�R�|�q�U�l�	ny���O<m���ZD��l��x�@��=�n��a�)?AԴi��O�9O��W����; �3qB���uL��i"��D�O\T���g������l��|�O�>E��hO������-\z�qX�y��'{��c�O!d]�֢ç;���&[I�5�r�u�:!�d�$�ӧ�M�;` �x�OF!}|�`�p(V�� ���?y�'E�)擦%��YoZ�<7@�4UYn K H��(�$�,��<1�'���DN��hO�I�O$����a@(�����lnj�٧;OZ˓��}�F
�'��ѻ��@���
�O֥1x�{��YS}��'��>O��z��H@/�:+��E�ʗ����?��K=<�|����O>i�ol�����ؚ1�0H�l	�Sɘ�.O���?E��'m
� ���*$�⊓F)�'V�7m�&\��.�M���O��С3a�{��8�'gN�I�"��'S"�'gҢF�<қV����'	o�T��n<���'E�_������e_pu$����Ϙ'U<�` ��8)j��q�����Oxmړ�8�'����ȼ<FV�3�/
�g $��&�M� � 	�'�7M
˦��N<�|1��0�������#V; T����}��(�X���D��F^����dQ��O\�g�ɋ�a
��|k`�B�,�����ɖ�M��A���?'`��&�EAы�05�����<�t�i,�O�X�'�6���47�̋b��7g��<X��K]�x���"�Ms�O<u9�)E����M0�i��Dc��	�Q�:��-�09O��OT���O���O��?��� �9Zh�� 9[o�{�/���<�����Jݴc� �ϧ�?Q��i�b\�ĐD>.�0,�m<+�B�Z�G����HR���y��	� �7Mg�<�	Ip9뵆Б'�X���.Pf*����Ի_b2��x�I{y"�'r2�'�RK&��m�Ԉ��6o�(P(�F�r�'���4�M���Z�<���?y,���;�n l��fV?.��I���`�*O(�d�0c��'��!�"O�f��%��:|�(i0G��P ��3��4�TxҰi���&�D[Q�kX���@X>l�z��������Iԟ����b>E�'�h6�	u�v�R���I��	1� :���On�dU٦1�IZy��'����M+�n�9`S�<��l�h��*��F�c�`Tk�Jy�T�Iٟ��P�����gSty��:QU&؁��4"4�s���yBU�t�����	؟0�IʟH�O`����[�|��M�e�ݾe�{`�xӰ๖o�O*�d�OВ�(������]<F���Yï˴�T���C-;��EpܴIi��&����Qnݩ�4O����:ϒ���Λ=(�z?O� 9���?�� ;�D�<���?A���*Y�*���C��^����U��?a���?I����D���ma��������""B�AX�	F���d����S�j��	�oZw�I'g��/eL0<jc�#p؄ꦛ�Lx4�آs�<�5lAG�q�6���?�0� ] XѲ�n�1���#dѽ�?	��?��?����O:9���ٙ=u�0iRKK�o���C'��O8�m�)v�je��ӟ,�۴���y��4[uإ2P�VM�8[��Ų�yR/}Ӫ�n���M��%H>ݦ�'G�pJ�ƅ�?q�E�(#y���@	�\[r���
WX�'Y�	ǟ`�I�������I.f��Ӱ<h!isB�(<��'<�6�45��O��-�9O
:r��7��%GA�ԭ mJ|}�lp�2�lZ~�)�S%RP��'��(NxƠ	�a����"
Z�y�z�'7�;F����M��+?�Ģ<a�K^RȨQ��)*��q�o�*�?����?!��?����DJͦy�Eu��{�K�	��çnlv@Z�����T�ٴ���|jQS�0��48n��'<��$�K @��!�(��L
�XR��޶VD�3O�!;�)I�FH��Y�O�`�d���$��*��� �KA��^�� �� jD�	#:O����O*���O���O��$��.�aμ��'eRJ�p�fM~�����O<��ɦ�
�r�t�I:�M����򄝑_*�G��vH��� k��O�pl���M�*�0�B�4�yr�Q7z���dN';�L����#�v���gϊ{b�Dz�4>��ʓ8zV�+O��$�O����O|��h��h���Wb��+nk#��&NrnDrA��<	��iQ��`t�O�b�'3�T�wF��R 
�;�	#ъ" �H��'�ȼ>Y�i��7�6�4��SH��P�V��[�|�`�K8�:����� %|�@§>���f�}Y��g�l��-O,�:e% ܫ��є�l�d' "M����O����Ol�4�����OH�/��v�I�f1����ݽ~�p�4c�%c�c�'^�l�r�O�)Zy��i�bQ�E:\4qc�u����Tow��d�#E�R7mk������pP�~�IP7S�$��H�'��dڧ�[$r��D��C!�M)O ���O����O����O �'v�ڥ$b�76�͸�#��[��$ҥ�i"<���R�����?�s����3�Mϻr����� (����Ղ_e��)'�'���O����'!��HS�i����<@�� �T/��X!/W\��
 �%�¿i<��'[6��<���?���?P|�S���>��0�u ��?��L5~�B���d�ئ��`k����ɟl�R�`��1��$ɇ7ߪ�⧇d�	ǟ���O�,o��MCH>�D)�0K� ��V#��k�	��#_�<��O5Nerd�*?��(O2Ѭ;Rb��nZ>b��:]`6x5�^(r/�KPET�TO�'��' ����O�n���j�QD��;����"A�)�l�ݦ��r�w� �I��MO>��3�/P�TX�8�@\.c<tĸ7`�\?�ڴ%>���'8��2��i���O��#�ہ;k��S�/~�[�nO�d�.L��!� � ��.O�1n�]y��'j��'W2�'�"��6��0��
ܚ?R0���J�ɾ�M�T!�Y~��'�񟎘a��6s*�Es�&��Uq*�E}��zӒ$nZE�)�:ZΝ����$�3��I>x4��.�=HXЗ'V|��q�8�M��.���< �P"�D����������?!���?Y�t�@�� �������a'�k�U����,�l�
Fҿ}���0#�՟�ڴ���|
�U���ߴj��'8q�ʁ�2�S�A�xE�V�	3��9O �$�� $P���2�`*O������%̐4����`(�j��9Q�h��<��?A��?����?Y��Tc&$��t�P�-z�v�j��C<`6r�'��d���z <�Z���ڦ�'��)�o�/g�b��Z�e��r����ēD2�vluӈ�	��S6�l���	�b��$���E8�5�Cܥ`͈l�BD$:h� ���r�'j��ܟL��ğ��	�_�ĸ�c��S@Z���Z�a����	ܟ̖'c�7��c���O����|:R��<pZ�
 ˏ#3�ۡ�_~rm�<����M��y*���QB,V���*@��ʈ7����L]�F��|*�+��M� �|���1]eP�ɲ�э�C�%���'uR�'����R��
�4(l��bG�}Q�tK�&���P�	 �?�����V�|��'�n�E��� �4"�1b)C&鶹��NT�&��6-��!��Nצϓ�?A�̓�Zh�)���	gm��G��PI �뵅��o���<	���?���?���?�.�>�ӵk5*�I��=Q��5�`(����������I��d&?��M�;?rV0@GU�A)���gA+@	}�e�i��6�J�)�.eB��e�l�G���QS�������uJ�Ir����r�t�IVy�'I�d�*���#�����Dٔ.2�')B�'�I�Mkq 	�?���?)U�G��H}��W�'�R��SIY��䓦?�V]���ܴi���|2�M4]���`�k\H����y��'J��� "�#��!83Z���~�6���?�J�w�L����b�J��S�G,�?���?����?Ɋ���O��ȇ��D>4�r�ݭ��!��J�O�Em��c��TW�6�4�μ���W�_ޤ��3��Q�9O��n��M���n���b�f�F~��O� 40\wMVe���}LXX�jK�=����`V�	vy���$N^XU��νu��Q@W�M��X�P����7��	ǟ���iǪ+��}� ��t� �B��4��I&�MKc�ik�O1��Q� O ?Lq	0��h6r��&	P�.��H�<���$Qf�ć�����D�1XC���s�Ƭ��K$�p�[���?���?���|�*Ot�oZ�)F���ɮ\�h"B � |�H��%��ZI��I��MS�2��>�ǻi,`7��}�u#R%���:��o�굈�	��#�~lZp~B"F3<x��78��O׊P�vM^��ׁ	�F�2�Tj��y��'-��'�2�'|2�i���5Kf�[2y�x�+���b�����O�����q��|y� w�ԓON��5��8~�A��M��	q��Ї�K��M�Q�i���-�,b��6O��U�v�j���l@,~v(�ҥ�JPj-&�:�?���.�Ģ<���?Q���?�Ƌ����֋]���@��R�?����[��k������<�O�0��@U�W���`�D�F���"�O}�'�6��Ʀ%HM<ͧ��'� ,�l�&�����	u9Tx����'��T(O���ڟ�?�S�)�dA�x�n0��F ���m�r��O���O��	�<�b�i̽!�I=QB���Ʀډj�����H$r�2�'�H7�O֒O�T�'��6�H�ZH�cg��Cd�@�.�7�0�o��M��g��M˚'���/z8��)t�)� � ���'/L\���S���9U>Oh˓�?���?	���?a���	�|ה]*��[)]Od#2L0LŬ=n����t�'#R�O��S������"/R�D�Hz$f�	OAԙ��d����.c��%����?��S�X��)oZ�<�r�Éj�%�ѯ�c���+����<�� �2���>����$�O��d��Z��b�%R!��Y�cүG���OH���OT�0r��E:�y��'�rkD���MÖ'��~RTӠ$�,��O8��'�b�im�'��#�
ĈtMf�S�hY�X��!z�O��Е ������ �i�����_ោ����J���X��y���w�Ǒ�?1���?���?Ɍ�9�:Y��"��:㴀�n��c�,�S�O<Do�>nZ��%���4���cF��I�DuI�/D�@ܶP��O��Dk�d�䄟 ���s������(�b�]3��Rj�2撝�'b��hܶ��|2R�`D�%�$@m� F�A֔p�ٚ���F�}Y���@y��'f���3K��>0
���F�:���SƔl}Rjt��o��Ş[�u��m/&]QI��#�x`P�nR/c?v��,O��s�aU;�?��O;�$�<�k�&�Z4kM���$Z)�?Y��?����?�'������xӉt���a�7��\���͊P@Q@�p���4��'��e��F�y�.�$��.͈��G%8O�\
&�{�yC�)��x���9�>d���qݽ����4�w��@J_+xE ���)��q��'�'��'���'�I�p��-iybɓ� ^; ;z�9O����OZ�oZ�-8�3��f�|ҍQ2,� ���)Y�O}�����#C�1O��D��	ÓZf&!咟Xcth��YwZ�f`��L0=�&}�ڬ���v�0�[K>Q/O��D�O����OnM:hs"X�"��$e�)�O���<�ipfdT�'���'v���Okp8���S96�YS@m-t�t���'��>��i�z6-�g�i>��s��c�?� �镋HL�JeR���,A:�p�Yʓ�F��Oz!(J>�Tb
%+=؝Q@��4E{����?I��?���?�|b(O��lZ�:[��DM�2nA�A�ب']�!�VJ�џ �	(�M3����4�2��'i�7�_*C~L�׮�.�dЁkU9y6�n��M���\��M�'�� ��w�re�ӗX��ɰn��"��I<E�ֈ��e��+�N��jy2�'J��'���'U>a�fI	%�Т2(M�M�&Ei�叓�MÇ	M�<A��?�H~ΓCܛ�w�^�P�$����0G�=���Z(�*}ӆ�O1��(��j��~G���,�hu�#h�fm{!N�LU��)xV�@ѼiQ"�'���'���'�
hV�ma�5k�40g>����'���'��U�x�4<�~����?��v�r��%��X��tŎ B�A�����O��'�6-B��m�H<Y�
P�p0 �� t:�Ðe��<q�l�Hp�jZ?UYh�9,O���*�?�1G�OX �J�8|-��rWOFd�(�`E�O0���O���O,�}B�"R
�����X���k��@�Z�$�J�u��B���D�Ȧ��?�;3 t(�c"�zN�`��A�Sr>��.!�F-iӔ�䁃|քб��	YFٙ���H(���E����s���4��`q薰�䓗�D�Ol�$�O�d�O��$�8ٌ����)���Ќ0K6�X}��� f�y���'NR�Oj�$�'r�B�R����T�܍�� X4Z&��M�u�i1O�D�O!#�e�|���"� Vu-�nO1y-��XpǇ"�򤓺=��a���'�ı$�h�')���P�.�}l +5�"!���O����O�d�O�I�<�6�i�jy�'<`9�0͛� �J�X���_��3�'^7�6��7��dIަaJڴ�?I��S$�*�Ñ.�:��*�@�z��5!��Q~���8!�AbXw���&?%�.M�L��H��MS�};t�_�Lr� E�4$�,8��ٺYS��(��G�d��#�K��Qk��{��Z�XZT�ۂ@�ezx�[�A� I�l��F�o�L�fԻ_
l��]/,m.��8t�!Ĭ�
�@��C�� �n!SG@k^Mzt�L �X`W���ȩug֣M�A�Š�l���y`�5KC���P�� ֋	�	��bݵa���Z8h��PΠ�kb�#t��uAҧv�a �J��1��-,nᘥ!%�#�Kd�2��Ƀ�H�	
�(�����x8j 
�E3Bdz޴�?����?ٱ��0̉'���'r��NSr�����E�v���3rEߺ��'�"�'���vA=���O��D�ON�a4�Ȩx`L,yO�1���/�7�O0�S��y�i>e�I韼�'EFEiWI�Jl�%�5�A����ae�.���?�1O~�D�O��d�<��Dƈf�*hZ"�Q�J�I#���c���(��x��'�r�'j��ڟ�I�q�ak�Jږ2���*�&F9GԘ)���<�� ����h�'�`j&�>]wC[M6�8 ��w�XU�@��>����?Q�����O��C ���Ɏ������.��XH6��?y��?I*O�$�ca E�S�# Xq��/�p�� �<^����ش�?����$�O���ԋo1��x���3�P�����I6�U
��S¦���ğ��'\܍�š9�I�O���ư�x4���P���0ዐV��y:ҵi��	ğ��ɛ,ߘb>��I�?7M ꔘ@0���$�b��'8]�P�0����Mc�U?)�	�?I��Of([3��2��\:B�W-7>����ij����S�D���43�ʬ��V�O`�pa
��R�dn�)F�]��4�?	��?y�������d͵���*��D>D}��!0)\�e��7M�%�V��?A���<	�e���;F>lM<��'�ڂA�0��E�i���'��BRnO�I�O��DQl�? �]r��r ��4�˾M,41��_����䟐�3�(�	����ߟ�TI�v��U�MO�L'�]Bs��%�M���>�8�顙x�O<��'���v�&�Q'
3'-@�i���W�1�4�?W�_e̓�?������O�w+Ɉ'���ie���X�̔:7�P�^��ʓ�?	��?A�R�'Q�񰆞?�
DX��P2c�2�)�ҷ�8�OP���O ˓�?�uK����h^�!f��f�)����)	�Mc��?)���'��iZ�q���aشiĘ��%�>~2}pd�-o�Bl�'���'��Iӟ��f���'I� (����#R�����`�����y�V�D(���d�@��}�O������L�#`\G�$��iB"S�<�	�?�X]�Oh�	�?X���B��)���[6L���q(T���'`bG�S��\ �y��vi�R���b����g�03`��7U��I�v�:U����X���4�QyZw�4|��	M�V:zePC.�h��4q�OH���GW>�������~��H��l�l��%-/�6�ۊ)S��'�2�'��$T���֟H�� 0̈́8�sM��)��I�H�&�M��F��P��<E�D�'B�ԩ���T"!MåH�:ѡ��t�����O��$�">���|���?��'u��!�MCR��Yck��;@%��4��=UF�H|���?��' �E��e�8}^��j�aٚ9�jZ޴�?Y�&@���O��D�OT�<:dK�8���/_w�-8�E,[�ɦS���CT�>?����?�.O��Ē�:�q��	�r(Z������ ��<���?!����'����/-c���&&pr��BD�l�2Ԃ�����$�O��$�<��2�.`c�O�؁Aqk����'ڼ(�����MK���?����'���+���شD�yӌӖ�%0E-�7��(�'�b�'_��ȟiңBr��'!�'
Z�n�����,44z�F`ӆ�$"����DC0�LO�"Ej�b�-
�j?�t���i�"^����4%��O���'��D��9X,�#�4b.y���Z���b����
JJ�F� �~�D�E�X>x����X#]N�i�u�b}��'�F�{��'R�':��O��i���7��g�Աa���=\�XlˇD�>i�UN��k0��A�S��s\X9�C�!Q}r�$��0��7-
�$1���Ov���O"���<�'�?����(T�6��D��?O��ʶ္E��ɚ%�"<�|:��H�<�چ(���r�-��=�"��E�i�"�'�2K�3��i>�������R��-��)ҴY�h�`�2d�j����U=���&>��	����#Zv��o�;[� �rj�R .�n�����Z`y��'���'�qO�A�p��(N}*!�ĥ\6%0q7T�Hi�F�Q���?������OR$1WFۜQZ� ���X�S��}���BКZ.O����O��d;��ݟtX��n�t�����=��i��8*�Z���8?���?9.O��DȈS����#Z�t�r�h� a��|�vkA�|.�6��O���ON����E�gi�l��B��j��`;�!JedNc�\�������'XB�׏l��Sɟt!® 8���c�IG
'"�(g��,�M���'��&���asO<Awhȱ&�¨9S	P�j4��'�֦��IUyB�'Ś�2$T>%�'�4�ش{�l�Q��!��l[��U;�db���ɀ5��YhE*9�~J�S���:�ߖG	��'O}��'|�AC@�'EB�'^B�OE�i�aITMN���x�g�Ia*達�>���^L�ꧦ�[�S�k��L�Ɖɕ\-v�ЖkJ�}�F�l��:��Ißh��ʟ���Zy�O"�d� \E
9��E�4^�4���mY,6�ёtCBub1���ݟ�)TBK�1pYav�ݼdNj@) Ɉ��M{���?��t0�/O�I�O�佟9qO\�Qؐ�B�V�7l�(��%�.�'O�m�!�3�i�O���d� �߀'U\�ل`��B��;p8 7��O
 �)�<����?!����'}��3ÂѪD�艒�(f�,���O�ݑ���+;�������Iny��'̐(�V�
;���U�ـ1��X��j��	ןT�	��?I��xɼ��Q��!u�^�C�	K��Кq�_)a*b��'���'��Iڟ8�e��Lڔ&�"i�R�3v���{��4r@&^妡��Ꟑ��\���?�� j�Xn�XX��9��z$���$C,��?)����$�O�E"P��|:�/�hQu��F�k2��s�I�Ѹi���D�Or���H7=��'Τ��!U%eS��(N+�����4�?Q-O���̣dS��'�?����EC"�(�V*-����JƖ[V�O(��ȑ]��r�T?��e*�#u6I�qI߾l�L�pǣ>��M�a���?y-O��I�<��`~�UZV�V�8��ǫ
�@Y�'�R�%Jb��k�y����H�r�l�2�Q�3��e%֦�Ms�,ڍ�?i���?����)O�I�O��#pb)^~�(���O�VZ��#����-�����e�c�"|��c��)�F��l�KC�
�Tq��i�r�'l��A���i>�����+)����tD�jրѣmi"�Je�Ěg�m%>9�I�����2����.C�[����ՉA��8m�џD���Ty2�'N�'BqO|���L��?�0�� H<,�83�Y��G8x���?9�����O�s�kD�o����US�r����I�d��?����?��'�(� � x�'Җ?���� ӄb8�a�d�Th�ܐ�'�"�'��IߟԳP*[fZ֫=oE�x��^�g)"Qr�)U��Q�	؟T�I`��?��4+
hm� :,La:  Uw�ziI#�к��7��OZ���O6���<�a����?����~�ϣU��� ��	x��cH͈�Ms����'�R�̥���O<����
a�h���
����,˦���Oy��'������O��ꟸ��4eC� >n�ɔ�-V�8aC���D��?���ErJ|�<�OLJ	SW�W�Ǵ,�TdE5-V( `�O`����*����O����/O��D�d�����e��|�A���I�Y��I⧯#j��b�b?Ӧ&W�1��@A�M�P�BXs�'{��\� ��O&��<)�'��4����H.K���RfX?\�l}�w��5�0o�����p� �)§�?�7D^�(�P���Wl>��0c4Y��'���'O:܈vR��럸��M?ل!&M_���c�mG�L����/2�1O�X��GP������	g?�v��<WE�P��J֟h�.��,�I}rj�U��	��p�����=	���g�(�� ��"��9Au�F}R�5=����O��$�O���?�&-�`5*g��Urr���d�|�ꉉ.OF���O0�$8�I��s�l��FE�D�r��`��MiBn[�lhՓ��3?����?)-O2�d�\�(���)�� u�Àh��)qm71#�7��O��d�O�㟈�	�1Y�p+P�u�ȝ�JP���%��@D�T�-(�]�|�	���'#��O-d��㟀`��`��+��ݩ��H���	��M+���'$B��iX�=`L<I�
T�|�pؑ�G[�L����Q�Q��[y��'{~aZ>M�I���J��l�Ǽξ���\^g�H�D'��ٟ( ��3Hb��'L��GnZ�[ ؊�Ҍ}�8�l�iy��	pj`6�O^�D�O��I�L}Zw�TDx@A\�O��������X��4�?!�!2͓O��۟��}bG+� U{�|����F ��G�: �G�?=�87-�O����O��i�g}"]���,Xr� �l"YH�Hcᚹ�M�4'��<����D"���� �O�&@@
�����YRd��M���?��c�E�\�@�'G2�Ox���_�Y��a�F/"/�^H��i�"[��3B,k��'�?����?��R�+8�3���}�$�*B֭Wɛ&�'� ��6 �>!-O���<)����d64���I��iG�$YPLn}�ǆ�y��'��'��'o�ɀ#�L2��İDv��"�dVF��a'͚����<Q����Ob�d�O䈠���&cz#AM�.̬��e�)�d�<y��?����Đ�RYv1�'/¹���
sg\�B�[��$mZzy��'�	����	۟��dx��s���dOĄ���R�l�0PI�	��d�O��D�Oz�-�X�]?��I�dN�!���C��������L�9ٴ�?*Oj���OP��Ҏt��D�|nڮ4��b�Ze]�x�҄�?��7M�O���<Y����՟0���?�C��3d����Ìt��hT �����Od�$�O�-a�6O��<)�O.-ل"�s����Aܾ@�����4���8+�n�����ڟ��������Zy���[�0H� �G�0�8�;»i��'���;�'N�	ß�}*��8P+�����@xLh� c���Y�NE��Mc���?����A^�Д'Ođ��*��R�8:�&̪7�d���t�L	�?OڒOX�?��I�|�bE�C�ʁTR�1k��tv����4�?y���?`3*���Ay�'G��T�AN�����S���)Oܡ	��F�'w�I$���)J��?��AN���N�5? )�B�FQJ�R�i�,��e�듯���OR��?�1X5@l&�%)D����@�?=%�'eŨ�'b�'�'�2P����=�
iPd�ƪ0���E"A�r~���O@��?+OB�D�O���:5����.X�̌+�^-���0O����O����Of��<Acm	 Ni�	)$G��+@�E��r���{��6T���Ioy"�'��'�����'G������;G�Rl�C�)K��&�v�����O��d�O�ʓ*����E]?-��>Bo����� v�-#C�*';�}��4�?�*OT���O�$F�Y�1����ʬWj��)&�I5=�N��B坾�MK��?�.O��aek���'$�O�^�!�I�k��L5����7@�>Q���?	���^u�'P�	@RӂǠq���q�/h$H@�\���'DZ-Hc,b�x���O�����|Hԧu�D�p�p�X7�DEˆ
���Ms��?�7���<Q+O���/��a�d�"�_wpt���ؒt�7�8&X�8l�˟����S�����<	� �/p��HceG�A�D�@A_�6S��B��yr�' ��x�'�?��*Fp��@&l�"2���q��@�PG���'��'V��+��(��On���d0�&2����Mو/j�hrqb�ޒOh ���O.��Ok�] h��qҥN$�}�9u"�F�'�^)��L9�$�Op�d;���zs)�][�E)��^)�\�!_��q�a��ʟ��	��'��|@��� �`�O��^u0�&8$��O��D�O$�O��d�OJ�1�#�T�`��$^�2В5�؎]����<����?9���$��&�X�̧�  �.� T|���#V���%�|�	hy�'���'sFI�O�ۥ�=~�� 
��
L�4��5]���I�����oyB M(@	��t�2u.�L�̓AX�db���A��p�IßD��z��	V�� <�0ChV)�r����K)Q-�W�iB��'8�ɨppp8:L|����C舢fx̐�M��M��躢��C��'�b�'t@
�'��'��I-~�6�o�#4�����Y5Gw��_���e�@��MkuW?���?UC�Op,��`(lh=h�̈#����i���'���YC�'Z�'lq��$�><���Sk.{�Q�ǵi�:��'�q�L���O�����0&���I�,��R"��L�^�8�kA�z�@�k�4������Z>��'�HɁ<P5�&2sI6�����,6-�O���OR���EB��?��'��<cVdZ�Ԝ�U���@�(���4�����C���'��'Θ�;�U�Y�%p�"�H�c�&t�j��F�"ϲ�'���I՟ %��/��E� �ð<��U�����.�o�����d�O���O��pV��Ñ�$�h���\��-�u瀕�}��'t�'k��'� DC�"j�6�zBn�pcd�bK�H3�_���I�����y2���VX��S6C�>m��B�@�b�b�c��듆?������?��\t$���D�i �{r��:�H�06G@U:@^� �Iɟ���Ayb��%\��� �D�Ǥ'}޹bsH"?���������E{��'T�\r%�'��i��0"�F"���b%�	|p=o�֟��I]y�,&|��v��kLɹO�W�
�G}���T�?zb�O*���8�b��5�T?9�V D&t��1�@��'uϴ�;��g���O�l����O,�$�OZ��㟌���Okl�uJ����á? 6���	Gn����'���#��3�y��4L��P �!-����NZ�H����4�  �]�ŉ��?A����X��OBB���ޢXSn�@��Ѵ
w�1� m��Q*0+(���?I%��	{@N��$J�{����&�"Iw�9�ߴ�?����?G,�<�?!����)�O��	�J�$,5�Q�D��ݰTM���jwN-�ɯ���H|���?���c^e��Ս>��1u�����ֿi\R!ߝ1��I�����OH�O�����L5��:����/�u�5�Sx}2�OT��ك�O���O��d�<q��T�{tP����z�٤$C<|(���P�������	ǟ��?Y��[�h��<"��W�F�(�!�C��gl8JN>i��?����?a�fo�;�OϪ����B`��^��A(�Ϗ)�M#/O�� �$�O��d�mv�����iT�q+fH�.�j�`�I�"��Z�O���O@˓�?���?Q��?�V��l�2l{��MޒR`��0z��'��'���'(�l�P/�-�ēl#`��0\�֨Y2蓿!��o�ݟ$��Zyb�G%��:����@�F�mD%���;%��#De�R��͟t�	�Xj�"<�O�*����J�观�?a2�;�4���'"�o����	�O��i�p~��dm�� w��DI���ReE�M���?�R��M���OKxHȇ��KΎl�S'�#�v�Pߴ#���T�i���' ��On,ON��E�0,|bR0��!h2S��mx]�#<E�t�'%>���	�&æ)&#I@,ѡe��$�O>�$�;�˓��	�O��I�l����dDˆb�h��W�W���c�L��#'�	�(�I蟘�WV�lO���SA�!M<���!E�2�M��.-&���?y�Y?��	a�	�l1dP(�l�7���T.M�J�S�O��0�ǐ���ʟt�I���'L��ZA�\�L���7-˶W*t��c_;�O����O�D#�	OZ ia*���^����`t��`8�ğ�I۟,�	�l��*�w҂�@�КLZf��1#@�{2-_Ŧ�	ҟ��	l�Iҟܔ'ԕ��4T8�7=a:pA`�#��"B�\�'�R�'aW�`��j��ħ�qS��-�D��O
�5k�1�U�i+|��'*Bf  ��'5���S��
s�\��f�z��(ڴ�?����D�-z<�%>a���?���8.�$9Y�j�$C���C�S����?q�K���Gx��"@�F�S��`�IkwVةd�i��	������4V��Sǟ��S���F�H5�:��9�K�FC�o���'����O��, S�C�lTL��lU� EX@���iH����j� ��O��蟬Q%���I�J����� 03> �E���eb� #�42Ͼ�Ex��	�OZA,��mX"�ķ1c~���;^�n�����	ϟ`{d�ˠ���?����~��B����A>E���a����'1�Y�y��'��'C��y�B=g���`�G%Hp�c��l�8��ͮ$|�$�x��ß�&��X
e�X1���O��P�ޞ?��ST0u�=)�BG��Ja"]p"t��X�$����@yp�I���\t�	��BD�E���KUj����Ϙk	Z�:`�]PQ��tŖ**��6�D-��ňu�
?AC�(��?k�f�k�m��2��u��x� Aӧ샻<�^Y��@�W3���4�)G��H*`k�+�����D�(�q� 
�H�.Qz���%u��!��E�9�t��נ,�,����I��-"ǃ;f���s�MͼG��x�o�KQ�x��!�9�	��\�q<�1����E�t����@����=�r�a����X��4I�1��ɀ�4���7�W�)�&8��3�Q�B��M�Hhx�������9���/����D�#�`s��"G�J�K"��X�Q��5n�Op��!���y	6�sdGA"[lD��q�B�mc��I|����	�%4�P%i$-�����>�OB $�� �z���5͜X����j����=O�QFI`}��'J�;]=6��	ҟH�ɥ&�&H�B_i�h��˒]�`��̎갽�ՍϢ��q��S���'��	  ��(��)�1vK�x�oW+;kN@!MΒ%��*Tb�O?�D k0q��i����X����8����?I������|�cܩl���F��w���F��:�y�� }F�OI�g.|J��$�Ob]Fzʟ�8*��	&ĕbF�ݤ9`\m���O���W'G�8r��O���OZ�d�ĺ{��?�p�Q�
��Zre��[���DfU�; ��28:	æN��x
�U�g�'���"+'0���'\�/��t��OṚ �+Y5�P�ܓ����$�	a�%���'f��c0����ٿG��'�ўԖ'�$����Z�#ꪐ�t�sK���'0V	��6lE��n��qP���*�S��R�d�'n��M���Ŷh�Bژ3~`�rG���?1���?��o�������?9�O,�}�eh�+�L���	C[����J� ���ۀim$4A��'HtA+f�^dȡ���^��d鈀���B$MX .���A��'���
���?Q�eL5w�8�s1�H�|T�&f_��䓆?��������ȃ��8���:iɲ�Z���#�!�$8$Rڽa��)?�fa�!��Y6�Dd}�X���e�Ɔ�M����?9,�35�;mfh!����{?���P��/$���O����=J�����&�� QF*OL��'-��8 ��	���������dѐl(��a�Q��N�q�k^���)�);�p�Bnģ`v�K��
�Q�x����OR���Ot�$�|j���#!�=Bc-߅9��Eyh]��?���9OZ����,F�nq���W�uH��:��'BDO��дl��,����G��#;d}�E4O@U;��[}��'��S� 
���I͟|�ɹS��! ��i�V�`u�ثL4t�+J�r>�X1�툐c�T)S�%ɽ���.����4���^o������Ër�αb��#�:Ո��/)w�a�JзbS�F���V4]`�K�T�`M��%��p�i5 ��?iӼix��S��?�'�|Ar�G� ��h���?�m�
�'�20`��-v<ܸ�$�D�])��H�'�7��O��{1`T�+ީDj�(yP�c���O��UB��"���O,�d�O|����K���?�"�sBY2'�F�a��0gĊ��VhH��D>��b�fOD H����HO`���B�;��m�AkN7n)������$6FJ���ԍ+�8���2m��!ғ:$8��X�"��LR�J/�����c���Ɇ�M� �i�O�OW��$j̵Chjɲc�,V1����' ���×�O�04��zBf#�o&� ��I`y�Y�d�7m��݈YJ�k� ��`�[�H�\���O����O0�JSM�O��p>]y������jA	U�=J���Ǩ�oЭ�CK�R���H��ՕD�tD��Ò���J�$��n��J��ɿxR�l���;�j�@ƶVxX���	>NJ2���¦���[C�J�iŖ�IY|�huJ��M�"�"��<��Ҕ�T�����1�x���QW�<�2�^b�B��3�J?^~<Hx�L�<١S���'�F�#�e���D�O4�'kz��S��joj-�	�?m�xM���C��?����?Qv��)M�����POD����K�u3$x��c��p9�/P�1�Q���KFBUdX�qE��?m��$>)���Bu*nJ4��3l]4Jѡ3ʓ:��I��M+��i��Y>�j�@ #�$��]XH�#�$-�-��L�S��y⎁�r�ڰ	F� ������$6��|���x2�ü0�ܸ9wO9��6�,�yB��'X˶��?�-�������O��d�O6� f�91��DCc�R�P����W`�F��B)Z�E�k��M�Ou1�2L'&S�A �E�� �˅��)+CD�kq�p#�����\O%�1��>T�9���;.�<��K4���:�o�(0R7�ۧ��Cp���o�؟PE���i��t�Gg����Ya$NڨI���̓�?�	�^�2�� Y�,��@U�!,�Dx�k:�-,ҵ��Kc��ڡ!�<"�E�Q�������?�%�ML�Y��?����?�A���$�O0���h@��n%{�G�S*,`i��O�hA�����*�'��I�`�Z'l��S�H@�x���'�(� pbي{gzxϓ.k�M�D�M�V��`CĄ� �n���N�؄��?��S�'��X�pJr(�Y��At�Ո4�hpP�&D��kDn��Vd�xh֮V7�"A� 'F�HO�i�O��(9Ɯ!Ǹi��1�G��V���;MƼu�P�[��'92�'�"&���D�'�󉎤Cҥ!��'����`��u'���dNU>}ʼI�	�v�,���C��d� l�%nT��A��O�3�{�-&�O�8H��'c�+�F�u���/�0`[���E��' �I�D�?�Oe��)7�%b#D�D�;C�@a�'��袀`Q�P�s�g�8瀬3�'������M,,3��mZş��	j�� �#V�Y:^
H��̈�n�c������$�OL��� �h9�`L�lf��S�4��"�J�@ȑ�(�<xJ+�(Ob��	0ߘp����0�P���m��^�q��7 �Q�t���O��$+�	�O�� �@�;~��B�H�!��I���O��"~�Q~8��"蝄:MP��'��H]��񉁶ēB>F�{/ڒ\}�Hb0ڋ7�t�ΓR�dEXŷi
2�'���G�$��ʟ��I�Mre;��0  5� �/ZXFq0�Z�IĒ,	!�������|ZK~Γ�����O�FDjc��>Z������K����	>����B)�4"}���?��&Eπ��RfR�c5�Xb��H�,�i閧
���'�4���)u��:�*L�@�骚'���!ړA9�S�A@�Z��1(�#�.�
Ex2�z�f�lZj�O
����AӮY��ݹ�&�.��#���?CL�F�Bp����?���?�ն���Oh�(LHRX0�c,r�4�b�O�ԛ���Z����`�',O ���	�$R�r(\�V���G�Oఘ�/Z�z�h}�'�>,O�����ڈ����C� \���O��p�'�D6��U������Gy��-v0d��|Hčb�b[!�yr)�3Z�<,z�-�1v]�07�jh|#=�O��I	`nqڴ0�BvbQ��v��b�k�>Xx���?A���?q�����?�������=H��"�X9��l�.>8��*�r�6���	9wP���d�O�H�c!Ά]�L� ���;��aQ�'��l���?	�,ūDlm�ͭ*  ��
��?������O0��'1H��ku)��7��Xc�*>HWb\��^�@֥K� 7T��@U�	R�����	~y��1<F��П���W�d�Q�%:R��U�=R"�hB�Ѕ?V�)[b�'�"�'0����:O��O哵"B��Z�,Y�7�.E�n�T��<٧삮b-s��V�@k"T*0���~셈GA7D�Q�xK$��O�$�O���|���A���3b�v�������?	���9O��;���$?�����#Iߪd!D�'��O�����3[�d�5��}2BX���	Wx�x����1T.�5 GҀ'E.��� %D�d���o10�zBQ)T��x2�=D�,��݌E�p �d,Z �	&F!D� �v)�'f��z�J��2��`%D�����n��0:���*x�)A	"D��k7��m�Dٴ�D�c}(a�?D�|���կ<��u����4W��b:D��yw�57�
��`�k����c9D�*֪Z�{�%��H�Θ�0"�<D�軄��5'xe�p�I�W�p�*��:D�8�A`I&
�L����9*P�h=D�pq�`��#����%E�E�4���.<D��0��������3Lu��;D�h3�)�_��cv`�TU�;�a5D���ti��1�ܷ��(�4$9D�	��ѕHێ�J�\�hZ$�9D����ǽ�j(S3��F�r���(2D��[#�[�PfDP1�+�j3w�"D���N�L|X�׆��W�drdN4D����cL���l΄dw\=P�1D��b��_�w��[�7��y�`�$D����B=t��Y�CJe���j��=D��8�c�C̀��`B[�L1p=`c	 D�t0�[w�0��F.��'�>5��(<D��ȗ界b��T]HE�d�9D��`�Z|�b:�  3���W�6D� ��*\%��xQӣ���"�/D���Gd�a9��"T�ܫ"'�k�I0D��8���va $�!�ƁCL|�I��+D��1�K��P�.Q+|�QV7D�0�@/+] ��EA�fThDB4D�t*&�	�/��U�C�_�Lw0�1��2D��85J˾`�Q��[�O���@$D���Ǎ��+��@���m��¦ D�\Qw��k��E(�*�1W��("&<O����̊4F\�x���>� ���G�8F(��{A�Ą8�S"O�A��D����}C�T����Ց���(�a)��SãSH�Q?e�bb'r�u�D-@�d�vU�#k!D�ʃ.ӢG%� ;�F�
M��mҁ|h2,xP��C��b��'U��%87��ļ�W+���P
�K��q���'V<�S#��2g��+2�˱-R�����$l2Jt&������,�Ju(w�ܟb��&M+�In�Y�6G��ZDl�z���|��Ě�yZ��`�kő-u���'��9F�h�8@�D�����%؄�3���V����@D!��X�_ ,Y�K(�<9Ȓ�'`-ڐ�'��xp-�
HJ�#��%ck�}��'��<� ���!3��uEFx����&v�蔹�]q�<�l�U��JP��%�|"���
I)S�#��D5l�?�'e|`3�����|� c �M�;�\�s��fy�� V��Q�v)�i�'�UơU0��y4�C�9{��1����y���	5��,|�J�B')��<���0���A�T4���y�E���#�>C�:�
��h�'��R���6�0�1����`��x��[����JŠ܎�0�Jf�
���i%�P��	̟����S�6�B�՞SE0���h�$�!q�t�²i��+�l0��肁m�K�8�d� -D�; �*���{
�k1�X8Xb`� ��1��nZ���B&��d��)���	�X��4�J�ls�'��`%t,� *l:�\9�%���y
RJ�����
,��}y'%��Ms&#�=5�,`�D� j�h� �!'���2�4	�`���e���>��~����go���b��V�a�`�'��`��F�!`���/��x��	�D������V S�8Y��+I�/H̒�ݗ�� #��u�'>��6����|�)K(p¸Y�f�$vnUkW�%?9�Պa��!6~@���W�r- �I͟pd�4-6�UjU�5��Ԥ�A���b��]�֎��'Vm�v������9K�"����aHx��Q$!�	~�\ �,_;"a��Ѣ�O!x���l��k��h�(�-4�( �G0��'?�i�O��1��ߏ_��Հ��[�<�Aq�<����&L-���	cY �s��, М�O���2�!Ϝ�U���p�*i0���?�5��&�<\a��6�Og��<HK��C2��9#�e�NB�A�x��4�X~?5%0��-�@C.��D��$X���,h���N��eS��)%��+G������(ѨOt	[2m���.�v��K|�PQF�KV�����7�6����@��D��P`�o'XX��l�*%k#F��"cp|:�ƒ�-�\]�O���D���U=�%V�U:8I�ј�(x b[�`+tq�ԫ��6�UQ0���(��H6B�~B�L^"阇���8�x�H�z��5�c,��Y�܋����q$q�R?�A��F<�<��O��ʷ��X��2D
9s��Rb��<+����	��q�3� �/-��S�D����=R!�2o:wP�	A
�0��'�h3v�p��pd0���I-4R %�Y*��JT(��+D#� TaA�`8����RU�R����8,�ꨣ�ƙ4n8|+V���t	a�\1��C�L(�A��'N��ũ�)סO� ]2��7@��I�J�].�>�r���psV)F�n��a ���iE�D�5.����+�!�����5�/�1ю�Q�OM��1��֎I�"�ŗ�Y�y#��^��)��*I��|��'�`��KP>�"�[w3�,�B�Wx5���>�ȝ7됡[1�B�6���be`T-aO��{�	�U.ekG
�F���dE%G��#�U+	2=���9�0���P&Z� �(Ó\N0x���: ����
K_.TuĈ\�|��	L'[�N���鉇k��z�D#��#)��v�,{�i�j�)���3��'���X�dZ�忣'%I3�ԙ�N�-R�lp��酭����q�~����ԟH���郇W6&IK��W�^^��Q�W3#c�P����-#L#<Ѥm��^=�!ç
�&�����a~��
$V*�`@*v�RQ��#�?��P䦅��V�?�T]�@�ZC�)AfJH�ɔ<�@�h��];b{��!N�3J2�L˗D�v;ܴ!���[b=� �>O8MyR̈����vNʏ���p�ôgU����ݍ,g���5��IX��3�N;{���/�)����oEj�O���g5�Ӻϻ0�� C4)̖ê��dm�5���+; ����@87��"Uc�"��*�HL����R�&#=�;�D�Q
�z^��g���!��ܙ|��I�OZ����t� #N�Gf[�sy����H����'�B!v��7m�x�D��'wo,L��O �k��C2�<�ygi��	!��>�e�ݪ������gh,�ץ�-6ܬ���K?k�Ru���<���̈L���N?�K4�A�Dd�dH�ꏘq�t`��f�c�K@Y�D+���4�j�3��Ȭ �`d�0&�/J�<�e0O��HdWD?q�Q��>�a��C�n	��.�$[�PP0�5l)&1�R�'�$�����)g�`I5�ٵB7�CS�B���rť��Y��r�fZ�g%�	�6jv���'OJU
�镒.��S����MI�Og.IQ'�	��hl��n��|�O���b��"��� ��ij�8cQ���ЛK��|n)j]J0@%��y� �����M���� C��� (����0�	*��i8�		h.�93� B�C֭�@���,m|��b��'�0�8�iͺI��ɈR�+l&�s��O֭�'��H=3� ��M�ș�R�<d�QX֋As���Ѐ�)k��y�wy:h�aaJ6nU��ɓ@��k�r� ���_��$]��M��V�x���,�Ӻ�A\�
R~Pɂ��
{x4p��->i��@�d6OT�����<7|�	�N#��d��	]��l3�,(C.\]���=���D�Ob�p`��7�?٧]�Ql1�$*G&L}��M�� p&�X�Lʄ����ŢxŮ,(U������A��}Ъ�"�T6-��r� N��~Zw��!�p�Ѕ q$���y>,!�	�H\
�O����iI�g�I�1���A�A���x�烸J2�ZC
0��ɡq�>���(RI?��y��ü�w�[?�V�Ul+#\��n4w��qDd�E&�0�m�	OiF`B��4�4�F��f�3�I2|�xm0uCR	�t�	���DB"Iid��uh-~;�%�#��&��)DK�`\�RE�		����g���B峀6���U�fJ�$f�X`a�P�;���%Q�x��?>��i��C~2D>��$���9F'|<� ����^y�7�M;y�bP�ǐ2*Q�|c����*���%Ԣ���h�o}&�k#��?��?%E Բ%3�	�CZeC"���"[��B,Y6�)}R-UV�$�B,)��� Z�`�r%�
�06B�%4]�� 5o�h�B���� #�dX@�M_,s�b>�)�fN
/R[x�	�d��f�5`~]3#��m4��36�9m)��(t7��=ͻ�x��k�X�4�UjW40�H����8=�Љ�E��%vD�S�Y�L=��+@(VҰI�'�	��QNaX��"�P�R">1��!p
�H�&�1B�^�!B�0��ٺ�A�G	��uI��4才�T�s���d`��G�7tF���@I�9���%?�s�A4�$�#���Hݫ�(!D��9�j˾��X��C�(�e�#'��it$�U���xԎC�Q��'K"�t�u������
qb�H�'J2����(Z7[ma~���vVA"c
�I(j`r�T�b��@�!0�a����XDk �+0y\�S�I�'6�*�������p�T�8)~#>I���E��$�q���h�/ԍ@�|P�Z�f�:� 2pXb��Q���h
�����$��T�ds,�[�(����"U ��3PGFgAR��a��ٟ(P�G�t53�$�N8����$'���T��!<9<�Ӕ��2�HO�����U�ʪ̃Q� ���'Y�����@�d�K���"�Zu�A(�/Xqu
�߸ ����EG����5�^���>a��֚
�$q��O� f����k�Ʀ�XW)�nU�H��ȃ3���	�U�����8=`�X���d�yir��$'����w֮A��|2A��bϜl0� *�K�*hR���3%���p"�A�BL��'�l�+,�S�|	 j�2�4�������"t)6x`�I��YO��8����B���<Y�h�q�h�����_�t�vAv��7P����h;�tZf�U��*�s� �>m����I�%V\d)���3@ɓv�,��O�t��E����8V��'6����ԥ4��L�&��Nr�H~�UN��!)�0���/�(!��ed	Y�˘Y�Z�#��|�ho��?�'��1��Ϳu�.�k��T8�*�o�b�<����ą9�֕(�O����t�ك��A7jk�����%̘�c%N/��p���XȨhF�"}����D}? 
s��,%*�����6Q���I�+�d(S������!���_� ��i>m��a��Z�%�ּ8t�ӦΗoN}J�iUS8��KVX؞��e�}`�H���J��m�� \ *�b���	ܣT��0�'�Mԧ�Ob�����|�E��'s�́"*�,JΑC�̛}�'=���l^�y�D$y�M�2��x��'��M���%g�q�bKC�dTyb�'50-�'I�-��E�)����n�lhJ�g}�V4H"�]_
���I��yb�P�db���h���z�9����6��K�C�{B��rCDT����	�T :5y�/�(n�D5C�A�k���d�5�f�(D�ϔ8v(i`��� YQ�`6}��NMy2#UB��eµ�?�zm����4�]�`uJ(ON���	�/ד(#����Ú0~�×��B���b�|���$����f�>Q��>7#_r`>Ib��Eg���Hˌ"�@��	�NW@)8W�̟ �f�jp$�:'��\�T�৮J%D���p�cV�32^�'2�'xrhP���j�'H�1K �-m�&\��S��*M�L�tV	r����Q&�`����"�I�#��QЄAI�g�dI��
�e�"�O�� ��5K�y�`��L�0t��(k�]Pg������V�V,����V1+e�q��?��gy��"Ad��S<_� 8$@Wf�< �~ʒdۓ���\14t�!F� �l�$Y�}����KS'\��	��fħyF�(<)���k��H����4�xN�|�����Hf6�mQ��#�4���ɈO���Ė�m����N�(�!ŕ�
]n��"AĊE�����6O�U�v��5I�VE*6,��F7�n�50���<����$�^�@�:�X��A>g<j�zq�'���L��}Fv�	��>>�1�O��0�M8}�|}g���\s����I+'�K����f�P�5&ƕ������PxR	3��$�4�� ��<˔JF1��2�@_��bޓ)d�O�`�L��]�9~�PJ�������A�?�C�I�D�~H;@�6��#Cg*]N<�P����C�D�':��'X����)(�O�2�;cH�O�`(9�k	���H�`>Ā��؎�$�*q�4�6 I�9�d8(#���LWu�@b=}RN�A�9��'gܤ�(Yǐ����Քj�Z��'��1Y� 
�\�V(�[%x�'�hh&�(� �EC��Qvޡ��'఑yu�ӻr�@���aY�P�8��
��� hm�ъ�_��:�X�+�@ ��"O:�Ѫ�#y�l�Pkҿ7|��Y�"O�b�0�p��C	
xRN r "O&!���9r���pf��C�$"O��4"�/���A����(��ܨ�"O�a��_�T`V}`��~�ָQ�"OB�y��, \���m/2�K�"OP]�ԉ�!�`�P]%I�X\27"O~���[�B�̈́z�	e�V-!���Z�LQ�P�
t���y���%!��WZ1�B�@�T6`}3�M�,�!�F�(�T% � P��r���!��"a�lYQ��<3��z%m ]�!�V�@��p���� ��V `�!�E�����+ >�HڢOJ�R!�I�Z �������\�=��߆x�!�d�!X��c��.���խ�9h�!��AM�$yq W�b��L6�!�$Ռp��2��5��!�wK5�!�J�LQ��"0�^��c�I6k�!�D�y6y�f /"���CQ���!�D�ZbXD tc�=�4B��.t�!�Y
}���r�J&{ʎ�1��<1S!�0^����L�.��\��"��7P!��UNu�������#�"X�
H!�w�2 k�"Y�\��<���ƥa��DH�6����/��g���y"���o�\�0��>4��:�<�y�DQ�~���E 1<�(�A��y�畔Qd�뗆O/wb 
�Ҟ�yc:A_��X��J4&�E� !C��y�n�8J_Xuc�!���hЍG��yK?_載Xv�Ω$��Xxfg$�ybf��1���1Rl��dXU�S��y�g��Uh�5�4����z`	���yB��V����+�.��=��@��yB�P3S� K�m_nf�`�E摿�y���)3�b�z�':ˬ���Bٜ�y!��C%$=�kQ>���a2�[*�y�Q���䠑��8����cM8�y" ����Å� 1���-��y�C�%��1�`L	5����cL$�y���7Xƴ��� �,xff؋�yR�R�02F�����wH>��1�y�@�0h>����M�v�ґp���y2S4a%��%�)8��SUC��y�-�.O�X�%��,o��tγ�yR����<�;���&]��"7����y��T�K@���re�n=�h�����yR*�*�<�ٱ͇�m�p�f�đ�y��ϭLM�q#�Cm� ���/9�y2�Ҩ�n!x��.QjuP��[��yB���!"߻;H�[GGV3�y"! �E��m0H�1�H);g"���y��:V��'�0�!a�ɗ��y"4rM�w�ړ}I.�穕�y�X�k��*wb��#� [���yb��'�
08U&�"n`��!�yE�u��@Y�j؇-�d�;�oҨ�yK޺6k�1��-/�\1q�`��y�i��o%�48��+&K-"��'�y�[pQ����LH[�K:�y�AʢO��5s�b7<��xQ
���y��J"Z�x9��!.��0��ƾ�y
� 
���z`d:q.0B��0"Or�A�&ťMl�cB���$9d}��"O�Ձ�ȁ�!��a餀HG�.6"O����@ʨ�� j��y��*�"O�`�t��.��������t�q�"O��JE��j�=ªY�'] ɢ3"O�@�!�g�t�r�
�j|�@�"O�`J҈�{FМaP��?k�4�"O�a1Ҫ�k`rXq�)D�?K��Rg"O��"���7Z�꩙��	|5|��"O�����I�NXؑ�fH#M��+�"O��d���B$�9�ͮ~�r��""O�����S2l�A�@�O��Hi�"O4��Բ�X|s3OA8	���Bd�I�<Q� �+s��j�%��#��9I��UG�<�F��Z�(+F#�+Dx*qAJGH<acA��2	y������k�Ɛ�(!��2iƄ�d��Y�B0��U�"!�dұsC�ܫBf�j�Z!��(E!�#I�ddb0Ϛ�}bm����`,!�Ȉ�$��Q��3^R�,�P(ѯB%!��X�0�t����-$����	�U!��H�{��
���$`9��Gs !��7r��(�F�D�>���(ʴ!�d�[��� �:*F�(��D��{!��_�s'��Bk�ACHp���*�!� (=p�P�L�M/�С"Y�{x!��A7p��tT)�,)f! �|q!�d�M�V !Ӌ�0l���`!��RX!����>��0EW�	j��2©�<Q!�D�%@�0űA!�V���	�	�,�!�W�d~f,R�L֟-w�)Fִ=!�����@\j^v9+��/z8!�J0P��x�6E7�p$`���!�D��~�ҩU��6B�=aC�	��*�S�Ot�Pc�i��Ӧ�衤
�����' J�Y�Z TԒ�i�<T�����'#�ps��(&��␎�$5��r�'sў"~"7䏿R��� =#�.(�'QF�<9 I�����bO:r��@!�	Nz�<�E^�$d*��'�8pb�ط�^<���R��<�Ԥ�.�FE��d�
x��<q�-\O��Bb�]3Tn<����&.-�s"O�ZD�_��>ũ&$^Y�P�s"O�`�儼zW
 0�āh d"���I�O���K� )u2�!1�]�rj���'Ȫ�NF����p�GlT����'Jr��W牖!;���W�S�1I
�'e�X�R�V ~�bɇ�߼o���}��'��kF�_8Vݦ����';V���'r6�2��5�d��	܆A1��'��ݱ�@ȸlF �b�Xo8�ݲ�Oڢ=E��gN�L���ʕ 
�(pz%91�(�y¬[�}br�D2�t[�oͽ�yG��%@�YB�W	���ˍ�y�N�J�T��!�ƔA,p�$�ؚ�y��SZ�ty��%�0R�4��0�y�cZ'()�F�Z��Pi҃��yB�M��,�W�ɺVtDEP�̆(�yr≍B��3�h�yjш�X	�y� �<�r9���	:��`@啡�yB�Q&.�n!�5���H`��y�e��G Z�ڐD�"���7h�4�M����s�\Q���B���W���r̘"O� Zd3�]�S�8���: �F�q�"OR��L�*J�����΃,�h�"OZՊ��*sˌ|P�螪*D��O^�B�'�=Dl�AMO��2���9D��ș5l�J٫F�=x���E8D�ԑ��Z�9)�i��`��r�Hm��G4D�d��N�/(t�
6P���2s`3D��d(��*��E
g���;�`��9�!�dTRu��3$�X�g�~4	� ��QH!�D'A���A���0֨P����|!��\�$����ײ0�r "��ͅ)!�dD�mr��P�<{��my@`_${��6O��۠���U	Lh6�F1�ر�"O�HTe�F�0�݋��Y)��'2�DС+��QAf�a��Vxt}����v�E�0��a[K��F�^-�)p;�O�O�%$�98��y��C liR��2"Oxp	D˝%�fD�Ǉ�X$I�"O>�)�n�u�ě%L�c���"On��s`�*y���K���q�"Ov%h� G������] �"OE3�lŘVf�@��L�,��"OXI����1U$�,��
����"Op��s�޻DWZ���(Crh؝	e"O�$A�!ڔ&��M�#(�:{���'"O囃�>���Ц6����"O�)Y0/A�P-2L�l݈j�x��f"O���@�`�¹�7��36��`T"O�(����#tlJ��D�grꄡA"OL̰��J�u]��p!DMx���r"O* 1	B*?�0��I#g X�"O��	Q�^�R]�-�����r�"O܈�%c��S$��iD_<���H�"O�u���Z�t@�E��`�9�"O���K�� ����㌫-%�UA�"Oj��� M����W�R�N	ƙ��"OV���/[V��$fT����A"On�s�dеz
�o�S�L�
A��"O�0�v\D�3#�R��H���B�O5��"R.�)h�@P0�%JG>|���'�8���OۥI�T0¨T�)�(��'�rT����5�D���H9)���Y�'��Ճ���b��Y�I8.�J�'�P��#	 �Ի�K�O_zX������G�\A���6�0#a���B�!��+A��a�H�?E�N��Ao�,�!�$Y�xj�,��O��a�#p�!���)(ݪaꟴe�XUi�k��=�!��ه^��9"C�0+z�d�����!��G�|Qg�I��l�uK�}�!��B�=���q��4����d
�*�!�3SE(X���\2f��]�i�!�&I��]����x��b��-V�!�Ău��4�֏Γ ��@�^�F*!��=ּ��֙E�y��k�!��PeTX
f��a 8��!���sJ!�H�}�̉!�j�����Z&#�36!��A�z1{�E$+*2m����_7!��{�&=B�U$2�u���V�!��QƁ�w�J��"�Q�{�!�D���D��dLy�x�RU#A�#�!�d�6"�h �A�u�@p��/�me!�D՗VV�@K4K�?�������0l0!�$ق]���{򂀈EYh�"��B�0�!�� ���Çэh[����K}pT�2"O��0��Fi \h� ^�T\��"O��Hڴ��!	�(��G"O@�#��׸���aƁ΂: �QX4"O� ��*Cb�Hh3�J/e�h�G"O*Iq�D� ��b�kda��"OhS�(�'~�J�i!M�N\Y�6"O2U�ƊR	v���b�2�"O�8Xp���>�(�0�b��;���s`"O��Y���;MX�!*�`G�]��5�"Ox�0�NV8/e�T��n�� ���"O̸(wA�9�D��6�<W��lJ�"O�(&#�:�̚��­c�P��y�W2���K��^)!�fAM�y�EĶU�ܡ�%��>&P��r�N\?�yB쌥5�x 굢R1�"�0�
��yR@!	���Pe�����K�yRc�0�aRs�W��B��j�&�y�ƀH���A�.�V�����C��y'u)���P�G��r	� �L�y���5��}!��.�d��h��yr�؝G� pA%�df� S����yB��,L6X��l�O����#�y2��L^�����F�W���y2�T�f�Z
��@�� ����yr��!����H�, 2�{#�Ԗ�y�CC�S>�Z��!3�aK25���'�z%R�%�<[lU��J�2�*�y�'��U`�<��f����@�
�'�>|9@+�So�1�d(�)
e��'���`秙u�����ߓ�&���'��)���:���zt�2̌,��'����Gݭ~;�)S!���֜H�'�p��e�H�&9Z��`�$K>mj�'�d�H��ن"�5���}F|�q�'���	r��0�����Y6x��d��'���8S	�m  ���̀�:#���'찑M�)h�h���H�I-�,H	�'�Ԩ$��D<FP���
�w���:�'}"�x��Ҳr�E�F�U�m|��'�!�G@_0J���G��m���'xf��%i�~�bA����s�Bx�'�H���@ (fSE|�z��'��@p �>71�p#d�V�`bu�'����F�J�F�#����_܊���'�H��%F�8,�\�B�n�� 8䴪�'j�u����xo�Q:r�δ/V��2	�'�l��!�2���(��2=���'����Ƃ@�U�d�N���'o�D�U�/HS���6!A%v,Y�'ܜu�N =����D�D���:D���#O�&.��@u+�P�7D���u�сqiz%h¨��0ּ5crn3D�󗈔	Q"d9s�Tȼik�-%D��:�.� :H����Z�zĹ�P#D��po	6]�΄`�E(~R�)�!D����j�\h�b�;Th8�@ D�г�����
���g 7L�:�3D����'�&�ѡ�
A
�e�%D���Ge�/�>dsf�H�_�� /D���o36@@��F�q���Ҍ.D�H�!$�-X�xpZD��Z/`k��,D���<�x��m�'#�ăf�+D�l�Շ�g�R�{� m�ّ�'D�� ���񅟑abjM� �+�l�Qg"O�Ya&��z�p�
qF#]}Č+�"O�l1��?2�}k3�ta<Ъe"OX}�v!�2Mi��T�oHR=HC"OT�Hă��W��q�RfɪZ� ́ "O���"��zA鑯ǆ2�J}
�"Oj��4�¥H�<��ڶ<Qx�6"O�@����#ZpV́�&Ѭ?�Dz5"O�P�Avl�8JхŌ(%�8��"O��#���9��R҃v���""O��a��N�o�( Ѷ"ԪL�d�y�"O���"��߸�RQ��X;�AZC"OH�c"�AZR ���pʐ"O�@�F�����@�4&Ҝ< u"O�a�w�51и�T�U�G��U"O�ݫ��G ���(0�D�b�6���"OPx+��3X�D��҅� Hlp�as"OԬ���ߩ��I���v�t8�"O8�@��L��Ik�*C)���T"O�DpwN׵#t\B�	M��iE"Ox���@a�
ѹ�G�%rtT�y "O&��R�Z[E�H�s�]i`���"O��1oc�.�bD�>%I ��"OV�%솼T^�
�c	�a����"OHD3�=5��hā�+i�򨀂"O(�J�`�$]��,�᠌jN(�"OT�*�j�	YrDl#� ܎UA� 
�"O`Q�u#��Z@c�oT�w���2"O:0��J�M�d���8j�ɨC"O�(�!}Y�1GjìU�e�g"O\�q�	�v "��a)T<U>�ْ"O�ɹU,��4M�D�چI7�-B�"O ���*R	mۢ��c�){�]�C"O I ��G�	lHD	�"�:r�@0"O��!��^����� K���u"O���Qh%6Υ�� �䦉�"O�J쀿_��y���]69�"Op��G�n�0#�"����"O�I�b��aT�b�^�xt2�#�"O�G+@UU��p��ɼDs��Kt"O���*��+ ��c�
"U��S�"OE���X�7Oq���0M<�k"O��G�G*Pm2@��)X�0Q��A"O��!Υ<$�}[��­^���X�"O���E�͕��9A",G�<�H2"O�a2��TXؑ #D�}L}�"O�M�ƋP�Y"u�#a��W ��X�"O��	�H��K�擇'����a"O�hs'�ÿ1Y�ȁ�� �$�$l��"O�ݸv��
gr╱v/Ɇ���9A"O>M�䭀? 7�	*Ĥ�J���"O�LH�LQ1�aZ�D����k�"Ot K4fԫ+�VȘ
��! �"O��u���L�1�&{�(�z'"O*�q! !Tw�mi�+�dL���Q"O~���G��h�@�T*wE����"O�LbPc��J�Z�g���Y:U"O(�
���7A�?8\p!#"O&̚#��u,Ȕi�.��W���!"O��(Vn�=}�z���L���U"O�c� ���q�"S�""��P"OE��(����cU>c�qJe"O�5�s�լ�XS����wqV��"OF50PԨWh��0� �\�.e��"O� �Ԋ�	�5YhHA7��^�8Q)0"O�Xxbǽw�iق���u�]�""O�56
�$\B6���wBRp�A"O��H��	ۨ4��M�8[F���"OlHR�Ԑz���cӞY��X��"O��rAg�@���c"�&�9�"O��C�J#��p�fW?Q�Z���"O�P�4�Ų;�$���G���M�"OD�3�PL.�K�-�'Ԃec�"O�h���AE(Q��īV��p""OnM��T�J�N�@���P�@���"O��0&�\K̦P�ak�z!��Ӌ}��2��DSǸ�:��\h!�	3l�D���Ū8�X-bIE+�!��U�E�J�qg�	%�N��/�!�d]8]�<�ċ;q����0��>u�!�䑠k0�׋+g*�����ua!�ړJ�B���
D�C�0e�Wf^�o�!�DLv���K�ʗ	y�������tG!�$	�
QD�ӧ-	9l��x��ňt�!�D�Lg�K׬%h���L��Ds!�\=e� 0���=+2��bfI�'j��b�Cdޕ
���Z#���'�J4AC�<K�q�P"J�!�'����d�2u$pX�K>?H4�j�'Ӹ�I�'�� �P�P0�@�'V���>�a`�R|�L�A�'�bٙ��G?�01 C��T��
�'����&�ƞB�����>�Ty�
�'X8H��e]�F�=�6��*5&��
�'�l�µI�J������Ď2�RYP	�'���iЉPH>�����u���	�'^D䫗-Tu�dz���u�)�	�'��}�&N��3��0�u���s9bTQ	�')8%���J�R=�$��3�,\+	�'b 9���qp\���נ&�����'��@���Inl�󏉯*��EP�'�>�@D/�#ɶE�܍%4y��'�*�	P%#���u��,$4�i��'ZB�8Ҫ��Z�$e3$$ƫ)Xİ���UV�{�zL�hį�%C̪ j!�$w��	�R�O(�����҅Y!�̔*� �;�@]0ZO6�×�T�no!�$�!:
��26,u#�A�EV!�$
��*ɑ'��32�!�fֻ/.!򤋪`֍� G׊R �=�veE
`!�d�2>��1�f�>jo�%Q E�#.�!�Dռ'�v�AueYXv�3��:�!�D$N�����;>#�L#�ĉ��!�d�8~6���!A�t�"U��)�!�I�9��,J���\�2|����w!�dI&
�B�Y$�U�D>FI+!Fק!�!�<W}�p��Z44%�DH�k
�*c!�߂Y���u�8�QajِH!�D�,|��C�TP���)\6XG!�$ٰP����[���d �A�48!�dPB��q�)�N��q��EE�DT!�����6�YֶEp2kG�?�!�d�=��&.�W�0�ɴ�9!�$y� ����3�t�!�.OB!��X,�Qi޷��LI��ݕD�!�D�C:\��Ň�b�J8�B)�
�!��[�X��R�	)Z�j*S��
!��՟T�a��8�ƔI�@7�!�� ҽ����8��yh �	�O�p8W"O|�'[�UpVX����B�����"O(Izu�ҀTI���q $o��-8�"O���*C�'s�%��T�y���"Ox��F�:Aq\��F��
\��:�"O:�" /Z<�TEa�N@#[F�aC�"O�#��R�#{���Ǡ:	�;`"Opl�2���u�,y�#�)��dZ�"Ot���ɮ@P�� ��^0�v��D"O��A��֕FYN�{&�&;f,��"O0 ����� B�@[�
t���"O���r�L &�>�0��Wl	W"O�=x�'������ Ŗ>N�x�q"O
�5���q��|H�
82�9�"OF�{��h60��Cݛv�e;�"O� 1��"n���3��21��xs�"O��2sBZ+|��x�7��r���8F"O2�8�nϻ5Y�D+%�KWS�e�%"O���b�{��/Q 
2d��"OP�H�CM3�Ȁ��oy{�]#2"O��7@�(q�ޠ��+��y�h���"O~�S3!�Rx}S	�$�TLؗ"OP�̶ jιsq���"�N�sp"O Y �I�`4T%+A�[e2B4"O��S�!�,V���K�A�*fS4� �"O:��E��;J���\�$@A"OfP�o>��$ĥI����"O���d.	wOn�p �.��0"ObA�$�Si<�u"MD�lȎ�x�"O����,ٝC����wkR�@�=Q�"O�58��|I�!�	4rC��1�"O*�zH�-\Z�`��G��o?����"O�i����O�:� p��&yH|�"O�Y"�N�"i�@���1��p�"O"�
� ϑ<^�� S/��p""Oj��#��&4�0y�R��1q��ҡ"O �9����A	�l��s����"O�9��ʨ6��<�f��"#z�"OZ�)��uv���h� 0	>(�W"O|!�l�KL��th��|�j�r�"OXY˧AV� �����0Ϥ`;�"O@q�ƪռmt����;~Ä���"Ot��WE�tYr��X���r"O����,�lzU�T��iH�"O"8!`��Q�1���_�ا"O�y3d�n�Vtٳ.ӸSF�0;"OHa�DꌿL�BDpG�ÚUdе3�"O�M�ğ_F298�ɬ��|K"O6� 	�j��D!S�� F��ȕ"O-�1�Ĥx�����Ά5��!"OZU�P�M���1���`q8��"OX�ס�����(f�l�s"O�� �=�Z�	QFU� ]�= �"Ot��t�UY���[Uo��t���z*O�p�!iLq7jx�f��l9z�'F��+��М�HQoW���@	�'�0�BeS�J`�؉@s
$A�'3F�SFF�>��O[�Z���	�'?x�9��
4X*L�4����Q	�'��bg��,�Ȁģ4+F��'�r��h��y�q(Z�#.���E�<�#]�YT�α~��Z姊I�<�R�M8�De:���-7�6���L�<���P �Z��@I�J6�r��LI�<� D�Z�gF�W�"xb����gj�,I�"O��Z��ݹ��hqKY��<���"O>��B��
�(�ɦ���N��@"ORLsCCܺ}���*=�����"O�7�S�a����=s��"Ox�vY��a@��H>cr d�"O<�b��F;i�=���I����E"O(��T�	~,�Y|<�]��"O���1-/�6�!'��?,��{5"On�)�mè+��h�dh�$= l(sV"O:��.W�TАY�T�X�/���"�"O �	r�o�z(����s����"O4�;f�:5�1��'~��"O����g��A8W�]$k_��`"ON��g��̀b͸M��Hk�"O4aDʂ8F7"����	W��8""O�t�6O��,-ٳJN�����R"OVu5I��Ӷi*A�~���"OD�"��
4]\��qkW�bBL� r"O�uk�|�l��Ӏ� O[N9�q"O��2VnK*) �*��f>�1["O U�ƅ"&���Oٷ!'Z�BQ"O��Jchźo�ڌ(Q�W6 !hX"�"O4�r�Ɛ�F���bT���2��!"O� �A<=����G�3�(-��"O�Ţ��<k�e:�ǝ�S�|���"O��򍛻�+���{q���6f�Q�<��j��)��U��$.g�J��N�<�P�C�.~E�e�
���b�N�A�<A��ZQ#�&�/�-BR��H�<��d�5El=��àg�����|�<��f$B��j��x5���WIy�<IV��&X�KGɍ
/=�a�a�s�<�� �)j4���gK�2���H�W�<���¼hG�A�^�Y���2�(D�����_�9(�5
�� �����/,D��R���JH�!�A��J-|�{wo(D�l[�j�$4�B�CJ[:r�R��U*Ohah���3T�Փ��S>R��w"O<MH�PM!�-+0l0Ӥ��"Oh̛VÅ)D��kҐ"�l�Ä"O��k��� 1�B$R�L�W@9h2"Oڽ��kڛs,N�i �@��%�"O�ՙf�+Ɔ��CI��w� mir"O�9��o��l�4�����|Cb�#F"O�� �'È�zM��>)D%�"OΤ����E���XF/�=c,N!��"O<p�s̔	�,4���L+&�q:�"O�E#T`E��D駃��T�ra�""O��h����B&���$#	�t}�8�F"O`!��Δ�H3���gb�=:0�`"O�x��E�m�� ��#��Q�"O�|X	�RՆ�{�N���8�y�H�K�\�c�ɞ!����%�y2!'PN�Ih�U��l�!cA&�y��-W[�L��͠����Cv4C�	�0�~�hE�K�:�"�P��B�	sR�I&I�P�h���B�	�h�ryi��	=��0�QKA��C�	>��PAs.�!a��|�PkR�H�pC䉠+�R1����:pThqvfO�,�C�I�'(N=���2x1zw�K��C�ɳn�f��T�d��K��SR|q�w"O�{��!�7	�*
;����"O� �jQ�E�P�H�HЧD.S%^��"O@%�eMCWĸ�$i�/D�#"OX<5J8oFt����_�Z; ��"O��R��EKN���C�?ޠru"OD�pA���f����C�L�^ib"OF�D��G��z)���$�b"O���W�TRT�j2�N�1:ZT$"O�,�5���9|��ps�$Z�
�"O�T2$�[4@�:y�(Q���"O.����3p��P7G�\P�"Op��W� (m'd���~��%`�"Op��F�x9֍h�N�Y��Rr"O~��qF���/

����"O����g�KB�r�օ^�8��3"Oh�v��(mu�9�����EB�"OzE���n������CM�0�*O8ݹ�;S��2anĕG-�]��'#��rd��9��R��1�'2t�[���"nj��G�*>��ț�'�<T�TGI>ό��c���0�l�H�'�)*��pJ�@F��.���C�'����Ύ��)C�]*vd�q�'@�p1�3�5���8#�l���'�b����r���B�.L��S�'w�i�3�U�0���Z���hL��c�'�R��� lDn]�ACPҶuz�'cd����9Hk"h٠*�;w�|ah
�'�5@�CL8�����rF@�
	�'�� ��W=���O�V�ġ��'%�U(��$�S�#��F�h���'���!��)w�4ͻD��:C0ɘ�'PU�Wg_�Y�&����CH���'X�`@%A�==��S��&�p��'�t�cԆG:6�8���C�
��!�' ���K̸hX��RE�#X�v��'����� �@���Ҳ�(��'��&ʷ�f PA�U'����'����@.ɸ.=>�Y!$F�U��'C�0Pkδ^�ⱂ�܈n���@�'��� ����9HKS��R�2<h�'+@1�t��h�4��%�L`2�p
�'d�!�f�L�B!�1!!in�
��	�'l\\�!�˨<~��j�E0g��$�	�'Ev�#�c�=_��D@�����N8D�xӑ�Ы�R���l]-�^9aǆ3D��:U�-�2�15I p7���1D��k�H�(W2�ШS��J��A�+0D�<��G�t�93�jӘf���H3�ON���<����re��8����k	��<�V�����);H�D���
%�ȓ/����m߈b}���*��/��ȓkp�)R)ϸ[�N����:_����g�6	[ �-h�lk�&�4f�l��+�� ���$CW֑��O�::D�ȓV�б!r�B=>�`UҳM@�S�z%��}v����N9l©	���U�I����Yk���0��2+�2E����H
E	i*��	����	q�Ѕ�ȓCk�щ�g����S�N 6$��Htp��K�P�Τ���Gv^�ȓ7<u�4�d;��3���f��ȅȓ� �զ7gvHH��@�g��m�ȓ. YBJ oרh9��gU��ȓr�Be�e��"��ĠsO�Yü���S�?  ,�'�2� U��D��z��}��"O�L8��f��Y�� ��B�S�"O ���vrd Fe�2;�h��"O�P�4��m��HG�/sm�<
�"Oh�Jҧ�!����)����Xg"O�u����$쉐��>+G����"Oh���+� �ɰ�˺:ĕ�S"OZQ
�['"�ƹC7w���@"OU{��D5s�3�FN!BdbIJ�"OD��o�F{�p8���%���{�"OH=Xc��d�ؘ1T��)K��u�f"OT�F�6*�%�!;S�hLRQ"O�� ��_����U`��(��=�"OT]k� 	�dϤDIt��M���å"O �0��?"�������)7bI7"O"0w-
�V:D��"��4�bt"O֌�� �j(�Ikv+,P�c2"O�9	5'�=w*���)�n���p"O��	tnЃU4�������c6|�u"O����'�1sl��UR8��"OH�Dc�4��5�4�J) J`�""O��
v�B*��uҴl��=O(��"O:M�-1:�t=[�˙h�H�t"O��P�٢8�ie�)Z�p��b"O��j0σ���B�Ƀ�Y��@�g"O �1�
��d�ӈD<o��%!�"O��Iw	V��@]��|�J��G�IG�O�@���MQ�y���zK�/�(Hq�'���*CȘ,U�p@�C #��d��'����%�D�o_�`3&ñw��P
�'񂈫E�'�J�L|^�T 
�'�n�
�A)>*艣
�~ʭH�'��5 ��@�Q�ܼB��V��'�N��E%�@^\�u"��)�<��'&B$�Vg]�9l1�d�"i�y��'��� ��*a�ABt� M���'�(LɢA�׌�g�Ի����'*`9S�͟7r�h�	��U��'[���E�\�tL����,�"yj�J�'�h� b�����
��`�X���'�>�I1[�jA/Q�q�TE����"O~ y��<��!� D��S�,@��"O�A�Vk�X0q�Q�ny��"ObxE�&i'޸��ʂ7_4E�#"Oh	�P�"P7p`*���CL����"O-+�`@)�DT��(�2/�"O�e�9y�R}�0GG_Pvm�!V�0&�ȗ'��k�@�0��+��s�K8D�l����a `#s�� �JZ�G"D�$�!M��4 �̑rLA<xk>�@�n5D�@�]\A��7�fq��{��5D����T�Z��U�A�F7o��y�6 )D����@JT�>8rd�C	cʸ|
�&D��Hwe։�����A�1$`(aW�/���OF��>��N�@����@+ �V��P..�d1�Sܧ<�ŏS+��d�r��l���ȓ
�����Y+Y��,����>�����A��2�Y�h����g�K� ���|%��Nٕ ���M�TO���y�Ҵ"4�2����FN�%[s`ȅƓh��ۃo� �:2h��@��H#���<ړ�y"�.���v'�!x(�2�f���y�K:W�
��]�W����L��yB /P���+�Ώ:YbT8�瘟�y
� �������1,�!�А��9�"O|��׆�2��}�dT�3�6�˃"OZ�P%�
=iɰ����:t�j��5"O8\�'V�G�XxC��!�(�cQQ�4�IW�����U�Ü�"h0QkA)�2���i&�$!ړ��dS�G�!H�Μ�Ĉ�E��q=!��@=~�L�����Ox�х�01�'ha|���k�"P�Ʃ٬,���!@)�&�yU�9_��H�.�v�*���y��(@Q{ �׼�X|�]��y""q�P�2k��f�$�֥���yB��dC ����`�ĕ��J#�hOh�����xu
�HGNƪ=�>,A�hV�W"!�4��� �,��
����!��I��8�F���O
8�H�C!�$ݢU����ᏮAV����'Ɓ�!�� ~��c`��-���Ԇ��!�D�4<��v��e��T"�/� e�!򄀥U���s�G�@X�@� ��'���'���6�U�CA78���4E[=kx*T�ȓUr��8�D�:
�J& �H�,D��E�`��#h̀4�0n֠A�����A#J�,���'��_N�!��M���չ Jei�%�j��Ƥ�RdA�ƖUs �[�}�����0�tm�@ňtdq#�͊%ݖ�'<ў�|BV�F([Sļ�f�-u0= ��[{�<�G��HIR���P� 5��k���n�<����n �X�t��-"i�0�i�<!�\J��"ǖ���t0�Ge�<1�BK*0^��`�\��ݒ3l�b�<AdÑ3��-�0�����
xy�Z��'��F��/G�s2�� ȥ �v��Dl���䓐?�M>���͔/7F	{2K��`�r|r�f�!�D�`�PХ�#�H��M �2�!�� %�1�a�:
�vh���2N'!�D͈a��1���#� vʗ�!���:cd� 8 I�C�V��+ �Py�J2{��)`P��XZp�i�=�yr͕%���8��B����MX��y"��,B��9��Z�������y�L�apP,1#N3�&�#�L� �yb�Z d�&�IQN�&E(�{��Í�y��ߙ�0�˔�K�%^x�kE	�yR�Q5>͜U�P��Q���dnH��yreK�B��a
�MG8�J�qQ��7�y�j5L���e��2� e�'ұ�y"���*Ȭi;�쁗"Bl�3f�N4�y�M��
�p��"�3�B�	��D�y��V��X)J�`T�`
�HR5�۫�y�b�Ne0u�P��Hy��(��y� ^0	$� Ƃ�BV�+���*�y�[2�z$kAhP,~b�`�C��yb�Ĕ@|E�c�Y5& eC͍-�y�g��d��� !����(@��y�猼F��<���#�BH���X��y�oԯ� ��(U�ܮ���c��y�@ڬxx����Ix�>)2F���y",ƺYkfMB#�I6*�����W!�y�Q-G.���c�hH��B��y�
<d3rQ��aƑ~?H����yi����9����y��-)%����y�f�+5�0��C(��z��+�y2�S3f�^ճ4 I5 ɶ�r��<�y
�  7�*��$��*J 1@"O�(%�ӳd��+qBZ$/	��*�"O��Sħ
/�����[�X���۠"O�KU�$)4�C�F!�r�q"O.I��ط/V}����G��y���y��8`&\�B.l1�'�y2� ,>�VhY4�$�����y"ŏ�)z�D�5kv���V�J+�y��EP����g�Thq�H��yb���;\�ʲ��	��X��y� ����.�x�(�7����'f8�Sb��z�R�dC)�|1��'=��J�8�L�+D�0|��'D�(̴D7�@`��([V<(�'(�y*u`�4֤lk���E����'wh��"˺vLdze��0��#�'3❃f�8wT%	 ��9�Q	�'��U��NW����*~��j	�'���4mX�.B��u"�
&���p�'��������%#�	M4��'���BD(��;�zPkTA���l��'��PG�]=-	��ؐ��(=��'F��h%6DȘЀ�Q,y�n!:�'2͡�&߳qh�	Y�nw��x��'�i�喯f�J�h�X�n�B���'��ᷩ)t��(�K�c�9s�'.�����$!x�p��6Wmڨ��'m�r.�>:^�!�s�TJ�d�r�'�z����F sz��aQ0L, �'�����.@H��D&�"\�r�'��	�j��Lz���c�ͽQϠ�J�'�֔2V�Lk�v��g&K����'��r��\�`�씫THÊ+��Q�'��M��kGcK2m�CAz�a�'����'ʝ�H:��& W#_�h��'���P�ļ6�^�iE'�[�����'�"�*f�B����Ͻ���	�'_�Y��R�} ���f��O�a�	�'�̥*�f��^�Ș0ᐨ@����'"�a`�,{��� `E�-N^�)�
�'�T8g�V:S9$�S�@կEUX\�	�'~&0���V-#u)sM��'���
�'s�P�D��.��1�g�)Y�Q�'�xU�0�i��{�GW�� ��	�'���P �
-j�c�):�pQC�'����G/��ꬊ�I��hx�'���s�l�9i�`[����}��tJ�'�0z$�|X�� $>|&�d��'�n�;"���|_p�p�C�oeX��'��{��ɩ,�^��Wfǉ[�l��
�'*,8"��X�84
�
���$���8
�'��DP�ɑ)<բ݉3ΫM��E
�'
��ʐS 20���S�G�t�	�'G
 ��fC�"�K2�D:����	�'�(H����ݫ���:g��y�.�x X� �,#��xS���yb��S0ڹ�bN���>}z2�M��y+�7[�����N��a ��y�!��B7�փ	>����ƒ�y�)�&,�J����!y�J��g�1�yB�цg~������tn�a�7��y�41ER�h�Y``�І@���y2�R	:&�A�sI
e��	V��y2�Բ0��mӱL�Ej�����ߗ�y
� �� ��L�g�.|�`����HHa"O�Q	Q�J;�,ST/΍Bf)#�"O��;c,�v���Z�t/~�1"O�q0U)��)7��K笏}#x�6"O��0ChN=M2�uz�"
9*�"O�Qq2��b�� -��(��QS�"OxUs��ԑ��µ�!�Eф"O`L�$aN'��$��j,LF�<�B"O��3!Dҭ�1�	��B���W"O�,�%Aэ4B(+Q�{ѴeXU"O�p���Ӈf$<�qE�P�7_��""OR(z3+֩D,4E�������y���bE�f��3�����Z�y�EHz��(S��(2z��bF�y�͚2c�����Aq2�DX�g־�y��=F���]$n�ڈ�"b�;�y��6r��;e�
i����ņ�y��ӭW$���K�aՎ�"����yc8��@�5fO�R��4����>a�Oe�g�� qLƭ�5̛�#��Q[!"O��s��vŁ5K]��v�X�"O��Q!�G�P���ߌ+���Q�"O"�P���)q�^ YU���f)s"O,q�ү�W�t�c�Q�a
PT!f"O.i���+���;VO�!,\��!"OxE#"�Z6Kh^|{�Q"YVX��'|���<'���gk�&�fa�d�i!�dQ�4��+��g�0<#�-��Y]!�dʡm!6���ʘ�Ҫ����\!�$�8X��iU���}r�+�Pv!��3F�r�T��:-�~�+Uj��J_!���-?[� *D��=ʦTz�HʢG\!�[(2�>�T�� �0���gO:Y�yr_���'�T�`g��"oP��D�)c��q�	�'� �9��$o��8�K?���	�'�����Q5d(Lm[�㈟P>4u{	�'��`p4g�n8�9��<;%,A;
�'��9�GLC.hx��#��tg9D���e���k<�P *4N�x��$D��5N�J�R�2���&�6u��/.<Ot�D4�I*74>�xc� 2�^���
�V�B�ɕX�2�Rab�d�h໴"M�b�B��8|U�A�@��k*�$����`C��p8UU�٭Y	�A�%�9`�C�I�'b	
Uϙ� �O�lZ^C�I�o� ؀#�D�����L8s[C䉆A���AgɟT5� Ap!���T�F{J?}����`�0H1p�N���.D�ܘS��"el�8!RF�����
(D��E�$i�p`����N�lA�l;D��0�9T�M�Q���	Tn8�@�:D���K �i�:D���?<�&����9D��� �l \Mi���7.�Xi�V�;D�����]���N.(�.�xA$:D�X[ĈS�T��(��(�O�Ꙓc$D�y��O%
O�SV�D��aK�m"D��ٲ�L�<abǬ��u� ��5D� ���),�رʴ�+%��$*��0D��z��ʿr�]��	�6��ѐ�0D���w�1�*�b��]�UZӍ(D�pKA��t��s���b�~��J+D��	Q�Q�7���2��7~YxUD(D��St �!pj�36�^�E�'D��!����:0\j�����t�h�O3D�� ��)�ؖ\m����?D����"O��٣I܏�Wl�_�4�"O�L�Q&H�o�5����$��- �"O>�0A��o�$�q�2"��u��"O ��u�_&�Pqb�GPAP���"O~� �b!�F�C���[�"O��# �L�D~*G�֭k�h8�R"O�ѪcT�[D��{����&NhPx�"O�m����
��E����v� �S"O\��GE�v�!�φw4\��"O^l)t�^ Z`,
��_S�T#�"O�4 D/��&���2� Q:Ұ�"O����'B-9�`��`�ORƸ�d"O �"�/�� ��b�שX��� "O�@q�I>2�8e��	�\av0I`"O^9R�E

p�#�^�ݘ�"Ot(SpŅW��Uc��U*0�� "Ojy���4�A�b��< �9"O���M(h�(IH��Y
H ��ҳ"O	)�їj�0d �X�*�s�"Ofi�-�6$fĥ���C���"O�|��P+3�z��c���N��8�"OX\򦇉�&��k�.ALl�"O�� J�5:�PRB)�O$����"O�� =*;�Y+�
D� B�S`"O<�pK�"���gN***�ݐ"O�ha�!�'5��3���uyh�y�"On4j$�X}MVx�R�؉7b�T33"O���A�;r����فUY��Jg"O0)�'JR�m�8A�Wdlwd`�$"O(�T'�4�x����(RX���R"O2="'oW*Z�FU0����@<K�"O�8�����*�+�%6���C"O\ n��/4�92���?N�E��"O����'ZX���e�|%q�"O��J6F����qç���y��"O��2m
�&%��r�%��@�q+U"O����cPN�!pWjۉe��x��"O"ݪ��zۆ�S�E1?���	"O���'H X_�9�æ˺e�s'"O� ������0��"Z�!F"O���u�K�L�f(	�B�4;8c"O�8�qA�-y��}h �Ã_�B"Od��'���1���e���g�j�C"OLab�k�O�:pj5l΋$�R4�"OX�PR�
 � Υ/���"O���S��T��U��:�V=�"O�-��ު1p�!�7��N���"�"OfM��Ƈ�j��ɒ�m������"O���H�
��� CRu�r@QF"O~l���%WI�a�� �(8r@�j"O�ѳ���$\<�%0 /��ae�"OV���Ò�qJ���+R���S"O4`��"J�2���p��0�G"O�誷��;}q�D�5KL{	f�V"O�<�௅K;(\���~����"O&q8�J�H�p���P�c�R���"OT�cCJ�z�(��xzh�;2"Oʘ���X�l"��T�M$z<��"OMq�Ӷt�����OZjgV�"�"O"-��
��y��"��uyJf"O�ܠ��VX��4 L9Nr$��"O6� "D��8~$-ە@L�: zA�d"ON!��Nj ��X(?��#"O� �h�t�D�
B���s��)��y9�"O���pmߚA��H��(�|k��A`"O�|�b/mqĄa���P-
��w"O�)���Ǆ���jG�_�s"�؀b"O@�Q�o+$�j	�%ə�w�i�"O^!�@ �j�$:T�G�z`~h�e"O�UXPI�'Z~�yv@�b<���"O<���+�]�p�&�ɧA^Yp�"O�H)ed�"��x��CD??�ل"O��#�2ZJ���-4���'"O"Y�GÙ�lH�S��6}��"O$x��=[�}˳�X.3g8�a"O�l��C��g2<�� (S\���"O�lc�O�/V�PL�殒]RR��d"O��24�>�4�yum�TA�e�q"O��:��؆x�Ta!�Z�`0aa1"OlT"v�����@�f؅^7)X"O�ܢ��@�lR`�e��3F*�t��"O�`��(g��d�SFR�zyF���"Or]b�Ĕ zyH���ER�) ���"OR��A�>L�<a'$ל��mr"O��A�Mo��qд�@�|���sV"O�+#b�5>��P
�d�
��P�7"Ov����y3v qe�m}�""O�Cu��N�,*A�F*��P�"Ojhb���J��2�	"]�����"O2��D��~�f�(��T�s�B8"O�a01g�}}U���,R��mX"Ob�3u��"��%��a�~�H�"OD̝�k���� /+����"O(@�&N���H@�O5{����"O8��sM�2�lN��;���s"O��q�(�'��A�MQ�g{�I��"OlawhN�s������YAr75D��{��O��x�P'ï0&f�!#�1D��P@)Y��&���݄q�j�r�&.D�Xx�H�~�l�'�*sr� ��1D����PW�t(A�)C*V�rn.D�2�͔Z<��{�&V�om$EX`�+D�D㤁@�0� 9�������*D�����]~�a��̓��0�[w�'D���B�1�u#�a3^��x��#$D�T ��]awR91 g��Oh� *O���E@�t]���@oQ�!���ɐ"O%��Kع��-'[��� "OrQ
�l
�<m��ĉ ��	1"O��6��+R#n�{���z�"�a�"O�@�L�u���(Q�ɘ]���"O(1sT! ��@� ���Ըw"O�iC��T;�3Qƈ9&y4Ģ�"Of�h�dҩ&�$�e�[aJ(a�"O��R�#ãB���)*j2�� "OR��U��E@`�PN���1W"O�@;�X4E�F��,��|����Q"O
�z���7�tąH6��ݚ�"O��qF���\o�1�$D$M�<i9�"O�͑W�˘p������B�'"O@Ԙŕ�N�HzR�Y*O�4`�"O��A�cFY�,q��w|�F"O.@��
�w�`l@'Dg��	�"O<� b�\=t��ms�I�'vN4b�"O���e%Yi��hA63s6�3Q"O����Ԓ@m��bEN�V�m�S"O ���-O�xB"�	�D>"��d˒"O� ������iPDV�55�3"O�q��+�5|�P��B��R�W"O��� I�"r��5�N�BP��!C"O�0��g�b��zƯR�8f��"O�E�@H�(]�٩�,�i&p]��"O,%;��ٰY�v<[U+q��`�v"O��"%T�jC�@��T�B	ê;%!�D��Ot�!�P!�:Y�&LX���'3>!�WCY����D�9+��"�>3!�H$���0�A� ���0� ϑ9&!�d�f�q Z%o�يA�O�4!��0")�2�ν9�(��#�s�!�dЇo��X��Mњ8�r��v��~�!���bp8(s�"1�>M��*a�!����9f�Ö,�|}!���!��&9�x�����`�U�*+@!���4���⅍�)&L�v��/!��/j�lxx��݅qN�i�e�8!�d
�Yw�Dcb˒�.i��i g�Ud!�ɗdY
��ߡkeZ1����+rZ!�1xD����<|@�"�<T!�>��4Zu��63Į���٬ A!�'x�&q�G�	o,4؁!�
�R�!�U�+�D<�s�\}&��$�A*�!��h�0q��XN%Х(5CJ#G�!�d^�>�R��!g��MR����!��VHe��a^6�,�3�7[�!�Ď�)M&�ڑz���I�"��{!�D<
��ycOX
9�F��g�{!��бo����ƀ��`�3ÂӟD!�d��H
�}a���g����a��?�!��74x������3�	�woE�3�!�X�H�ꨛ�"B,oz��U�Z�2@!���S�P!��$�/3���CV	�jE!��_�Vp�1��vjY��G.5!��h���fnEaB�iCf�XL!�Ě���X2ϝQqv�
����~�!�dC��@3�2h��R�R�@F!���>�����9�ĘsC݀!�D@�,�z5�F�8P�=�p	�^!���s�����>L>�U;s�M`�!�D��R�2���5<7P�� �X9�!�X`�Q{!�$}�l�T�� !�d�9h���N>uz�L���ڛH�!�U��ta,ӂ�
$b���V!�?�N|��25������ՒBY!�dG*F��+��ǯ|?.�	R-W)@!�d
1W��!0�G���t�1�vY!�$J�?=�(���Q�v����n!�ER,�����|H��ڒtg!��^8W�ݩ%-�5b�р0L;]�!� *_��@ǲQ��XǀH!�dӓW� ��O	^�|i�e�7�!�S�
�TZ0��p_r02�O1#�!��͠�$���&K�$Y���c[?by!�DW��D�p���5ڪ�󑌛�e!��K���O?+���k��3N!��3K �d�%X�щ%lY�NZ!�dV2i�p��s�	�lK�xh���\`!�F�Ԩ[qʈ�+��P׈� 7_!�	�0�<�i&�W�z�V�Ȥh��_!�DU�d�+��2�>��*W�JB!���(zLPp��R�F1󆯒c�!�$�%x�
�! E�j�L�ʧ�>B�!�� �,��ݬk�\Ç�6ID�8�"O��h�O�~�%c�E�� c�|��"O��y �?s�&�X��=;t��"OQx�ߙ �ȵ!��ؚ2/"�!q"O�����k����N��U��"O^���M��Pٔ ���>~�fX13"OJ�H��Y1�B`jAi��+)N�X�"O��f�>����e�S$�ј�"O]	�S�w�2�B�g,Km��"O@t�V�G�4�t-h1��1rTNI��"O�5IW�a�Vu��1|��R"O*|;�/��/˒	�e��9�!��"O��Z1�l��{������"OVP[P(��RXQ`1+o�����"O�)I7�!���)��1~.��&"Ob�Ԏ]�7T&�1E��57g� ��"O��҆E�I�qcv(W��.;�"O��i%���T]�Ӧ��"��ts"O	�Ui�b3�4�'��<���"O�0�vG�v�A0�h�Z�P])�"O�@R���ЀhB�Zö$YD"O`�"B�F�li�5)�d�]���"O��9�)��bWd��@ռ/�t�#"Ofp�R�U�|�v���H-b��-K�'��'�剦G�� ��%P��v�(yTB�ɨ��Ͱ$`U�^��q�P�,B�I./��M+��sϲt��u�B�	
�6�{a���������B�	,_�l(�ĝ�+
�;P-M�+�B�	�q�VQ��N�2ij�(���1ۮB�	Q]~ɊR���Zà����J#T~B䉥L+dxҕ@���91��3m�B䉹 �Y ⊔���)�S�ɨ���\aG�)�iW3�Ĵ�@�^l��W$�!�D+u�D���շp�H���!�Dў\]�t�G=U����;N�1O���dQ4f����HL�5�� bA %�ك1�����g̓4���9��E?� �w"��(W�؄�mEH����&+�ā*��ʄ.p���{&��͚4�,Պ�P�&ܾy�ȓ>�����(�DH�kѦ2n �ȓR{Xx��|?d���"��<�l�=QK>���*>��tj!O��{&,:q��%!��^&K��@2�b�+_��R��(�'ha|V/�0P�TI�*	$���T��y��5���0W9[�qѧ-����D.�(O>u"+PJ�q��!��yS�a*D���w�r�ԽA�D5i����!;D���dG�2�hk!�h�i��F8�O0�	r��+b U�1���p���|-0B�I�`�+�O�X8�9�a�/'�nx@5���G{��)2B���J�
�/g�v�K'
�3�ay�(\@��h?p�C�.K�i��!��\Lv��I^�wUp�£)�w5,y�Ea_��	&�X�:�Hc��>I�JP�t�x-��N�D�8<ré.D�k�b�ٳ�����c�5ac���d*}�HB06̐8�=.�m�ClO��(O ���Ɔuxɺ"Jæ,^�,[��ׅ7�!�䓈Z�(b6��LI��)S����!��K�a_�;���C8��Calт
2��E�$�;�0��	N
�I�����y�	ե��Q�2"�/��Ip���� ˄�<��y2c�1J ��R�!Ș,��������>�O�4@M"n�- b�]��A�%�c��B�)� ����X�[!n�#d�q�	�5�'��OH��N�7k'*��@�_�&�x����y"�U�W��Y �j��Q�`��bJ�&��Ӑ��'�Z�)�ӶB����Tc�F�����*pW ��2ړ �.��A���Nո]Z�bQ�@���'��}nB�S&��y� ,�y�2o�_'�h2\�y�JA�1w��k����|%s�@�e¡�[+?����
\,Rja񄒫aġ�ğ*nD�@�A��~k�]�A��y"��[ȼ����l�\��va�8�(Of��dVTY��Ņ!)|࠳O�D!�My�R�Y���3m��0�Y!D�!�dӘ c@�S�[�(�$}	��� m����F{��������(q����ІF+�t1�%C�Ty��'׈�2pf��>N� �!*ϊ,�x��'L����G�l*��kȩ tf�3�'�DaJg���0!����"#�qДxR�7�� �3T�i�䢈�KO�lQ2����|�	���D��TmҼ�Ƣ�� �&)�Qa[4�!���T�YA����Z<Q4Aj�ay��ɾ=�&5�o]-2df����)�DC�wL�(�r�?Y�f����l�*ɉ'�*���aT%Rj
d��n~`-Jd�0�O��D�>�� �(޼a�˥r�<��D#�W�<��� ~Fl ���=�z��AS��?�
�'t$�R7DĘ8����$"�@�ȓ�|!⯘�n#"A�W{;O��0�y���'I0��1L�@
7��J\4�3&�'��r,ٳ%�X�W+\�i�L����A��yb(�$c�`�0@�v1�)k�#ٻ��>��ά<�q��S�Nj��D�9��=q��<�O�|F{J|�PҺv���sa��\Z��a�p�<іe�UF���N ;��q�r�\r�<)��h�UkNDr��拙d��,�'�tP�1A߳-��탴�"^?�ai�'����D}-��p����T�\1ܴ��X�d(�3�\([�*��N��j�`X"%����ȓU����wJ��2��G��o�����djܸ���
Y�J��W(��S~�ȓ_uP��Յ�.�߲^F��ȓ��}k�D4R8hTK�"Ֆ7& ���n����#%�ͩ�#��U=P���+��
�d��K�����8^[��ȓoP�Z�E��
���e��.��Ɏ]P�g\?�dh2Մ2�LK��J���	e���O���[$�W)`��h0%��Ya�8H�'�.�c���p��񷭒1L����'�u�B. �\%Y�@"s����'1��c0��Ng1`��Хk��t �'�l{��4o:��P�ϸ9��RH<��|8���!\=	@T�� ��m�l�ȓZ�(���K��=�Jp�q	J�P�H�IM<�$�ѵM#ܫF���@��6IWl�'S�?����zT�1IL�J��mZ�J2D����囅
VFq1��D���!q�<i���6i��(K7fԍ|���F��,>�B�I�o7<����.O<���	�N��B�>e�Z��\5)�L�����*V&���ċ�?�ѣ_�`��d�d�	0fJ�
BLIѦ��fV葐a�Ϋ����
�q���b��%�<�A�HG�$L!��"5<���"ظN�(}��H1HH!���X�F�@Ϝ.=���
��ӗE���r�H�C/�:p$�;��E�eHY��xX�����j�� �4{����׆�O�=E��� �H���D�ˊt[R�Ǜ.���u"O�:f-^"n�p��~� �մi�ў"~nZ���؃�P�#肰k�'{�fB� "g����K^5_U�2j��j��B�Ɇ�*�J��.<�y�p咽UH���2� mۤ�!��H������\ծB䉆 �0����؉*� H���P^�B�I�t��)�w�A�~�^��a�/c|B�I�lӔ����G�y�$�S�FFJ���7�	84�����bΖy�����m�B䉭m�X<e,�3
�A��D�M���'Jў�?�;S-�&x~��J#�X�5~`i���?O��IB�J��}�jB"j>�J�	�%ZO2 �ȓ6V���;2�:4�%	͝omN��?Y���~:��E�r� �{F`��	 ��y�`�m�<��Ӿ*b1��Y�(RT?�HO��}�8����	�%)$�I��I����ȓL�ݚw�	C��Pr�îI$�q�ȓDf�x0�l�(jP�R)Ln��ȓ,��\R��%a�>�I	��Նȓ�N�	���]A*�K��ehņȓ?���@R+S���'*�"�2���7�
��a�J}Dx�㜅duTi��Y���P�Eз;�aC$�PS�`Ԇ��$Ē���:���ׄ�`���?�bM"�m��*�v����>ͅȓ"�&����	G�@ J@�c�0��;P��D_�# ��0S㚟U�N9�ȓ��!Ɓ�;;�R�2�[���ȓd8\��"���.�b�2���%�ȓmð�#�D�G� �I��鞹��zξ�ځ�߳P�f���Ɛ3n���gpr��� �2-D���_0.�h�ȓ�`a7KK(���d2ʲH��rZ���.7'�U��'W�:�Ԅ�5����]>{�ܹ"�$� \�4��ȓp��lr!fQ�Nm�Egw�`��ȓ�d� B�Z �$Q�Q�%�, �ȓ[St
�(�* Jw�m��-��]��=����!��ԙ�Aږ~(�9��:^Ɯ��U�Mt-� �%sн�ȓqJ�(�d�
83Fr'Fٳ�A�ȓi�2أg8��R��/\�:t�ȓ6(�S��3�b�`n��
��ȓ1�)C�ŧS��!s�MG�,p���dL{S)�0�a��4�&��ȓ~�0A�-Spu25�Ţ�.n����yc4 �)Ű 伀@��� C��Ą�MΡ"!�^.Q/��s(��-���ȓx7����S��e"L
_h�ȓnw�x`0��+L�v�8�a�y!hф�	�Jp��jə(�8��YT��,�ȓP�hPy��F6�]P�O�������0����]j�f�kq��nl�ȓ'a$�էkG�EA0#ٚ��ه�51L(8T�!ƴ�G1��,����9��`̴J��Q�C+V>��̓�p��A3:&������G|��01�J`�P���`g$�k����y"mݮU^Y����6Ad��ǅ(�y�a�b�k���%��)���H��y/�3�*I��"i��,���y������H�CK8`$5x�����y�D�r��T�İa��IS��
�y��ˬLJ@���X:e��!pL�;�y
� �����^6�8��J�"AR��Q"O��x	 �衂�`?HCFE�t"O$����86��!�0\=&�x0"O<ȥ$�&<�DX�'�TAaqV"O@$��o�g}�@p��	�.6<�"OFE;�/���
�0���Y��Q��"Op�;�!V�8ИZ5�΋#�61"O�QeGֳ]���D|�n�""OY(�dӾ}-�p��\�wX��r�"OI�mI�Z�������Ip�("Oz\(���/�T�Z NP<��"OV�p����i`��D�8����$"Od�#�k\W NQp +�ip��c"O�Ա�	�@���!�A1i�H���'� r+�Ǧ3���<ɂ�P�_2x�T�\2��
be@x�<ـ�K�9 �.�?nӦ(RJty�@:Q��A��(��)�0lↁ�v�O����D�j`n1��"K��58�'M�5��h���3
�>�Nt�ߖ�Sp|��hY?"�����O���'��'K�P�3i�R�4���؃>�
��d�<�"�O3	�~y�g�\�&=���J6T� (��W�|���P��^1A���"8�&)���9c�0���Y3pQ� ��R#0�s&�xI�CG@��9�vݙ�LTuPS���jE�m*�"OnyYf�ʗV�DD�!�;*��>O�tIժD�(�A��8L�zQ�a��T�F�?�ke����y��Å[��e㐎;D�<[��I)h��y��Ls��Ғ��0P҈T�"��K䝉�G٩(È�?��3K>ym�!G��0X�:c"m�$�zc�ҍ��L	�N�#3ቨr��ș�J�8��%�7*F;^���r�-�,������f"=	��/\AX��f�H�g�Jq$@%m�<h���"=�w��R�@� ӵd �W�G~CH1#���3EΗ7h�5�P�Ģ,U�GyB�A9"����`��6iq�P��L nlZ���-�$��d>O�ʶ�T#+$��z��9J�dB4䍡lo^�?�Ȃ:�ṕB���]x��] �*�K���+�6L�w���"~��!h��U$}��FI�jm�Y���"x�La�aZ�Ed�\�V j�7�U�|�!YT&Hog���[���Uo����@�� b���I.{o�t�GM�R T �4��
a����e,�\���w!�:;`�e�b$�+r*�%	�~0�����/C�*�'Y�
���aS8>i�}�b��vt6ט�F_e��$B]6[���x`RAy�eQ=N �$��Ʌ�\pv�@-4�Є��#x0u�P�V�(V����,��?�� !,ӗsfͻ2���Z��<��/��"Y��W>.X���?���C�C��|���ZDBl 6�O+C�*(v�p?)20kxN)B��A�F��M3�(]�##4����v�<{�x���a�ǝ�fLR5CA++ψ<�F�]�ap��ǧR<��LH�h�څ�!�G�u'	U���0;ҠZ1�~�'X#9�a�CNfPk��N�Lt���e�ТE>��t�x�kE"C;�l���L�cE�����4�p����;g�j��M^�A.�)��@����[���M��{D�^3\� x���D� -7��h��F5_zh@P�:7�d�`$��`L�e Ƅ ���C�`OC �`�Xxt@@h�:6�L�����jd��� ޤy��Y!�Ҕ�^`A�sN�!�"<1��7(^)ăܚ�Jq�1J��K���
S�lt��-�-S��@ӄ�м��|���r%j�4F��K�aP�2�'��T���Mt��*��N��hK�q��O�PW�b�>-����>��D�95��,K7i@<@n5�5*V`ϊh�v#���`�e Ǹ^�d�!FI�n3�y#���!��*[x�1���l����� �x�DW3T�b��בݴYrA��/��2W�r�5O�QR��+�zU`�吩@Wl=�-��Q���ϖ6]���$��?8���3SWD!�p�M˶���{H.!�J��!ޡ�	P�'��0�s��D���c���Z��p����MsF�X�w�,9:�+Lw-30'%b���Q�̓�W�d�٤��w:]��*s��qHr��!&1vs�GFb�
����OV]��DȰ@Kl�2��F	��6Mӝfj&��C�Uu����%3=>�!fS~9�8yU��U��s��cc�����$՝e)�7��5��O�M �������-3���'$����]^n��C=(��qAb�i�/�	�����E��S�%T7"CKC�iRZ�mڐ�Mc���)mE�����W|��Z"�	p�����$I`��Aq�4:�Щʥ��"3�А'/��t���M(X�9�(�p�*Lrw+38�މ�%�Р0�܌J��C&q��	�M�(
� `���?hp�P:FO$u`b�:@`�.��v�M�f��m
�F(�h����8`QAc�9X��aT ��FW�1���5iؓ�M3� �g˜̂�֠r�:k(� yf�I��5�-�>RP����A��h!�)��⒞'ӈ�{�eZ`c�`�Ʀ]��Pw ʉNr�X;B�u����I?K�������"%�h���	=����t�^�>�)b�)�k4��ӱ�H=N���QC�!$�d��v3��Err!UX���Ɓ��էO�W~R�������^�)�6��J�l��>P]�IjBA�8mf	*�(�U�T��^:I�Q�C�עf��8X�
�l��y�[�,�9��2AR�ҷ��B�,�AZ�M�I.���J���R�5
�6�p"�@�J=&t�t+�< 6�M�p�Ϻ[��S�� ͚���v� 4�pc	&����L�Fo�E���n��!��/̂@h�F�S�tX�ƌ;~�Ȓ��O���lA'����H�6+��+�S�Gl`!bnX=?�`8��>�.�&�����3/��+1�S2Ei@�13��L� ��L�`�c��S*S��uY��ʰ�T�2.@:��%�K�^����,;�P@��V)1�
f�E�i�j�IrG�r�~�2q��+c�R���nF�!}Dp�LV�;�RƮDj�f�	�7�� �d����gP"AA����'��,��>���ǺbG�����԰��Td7���HE��U�P��ǈ�P������L�Rk0�H�ō�?���.����操P�@��q�	�T������l�B �v��C�qB���l�`����n���Q��۶�V�m��d�ߩA�er��Z�i�x��V��k���0𢅙;O��MR�#�ڍQ��]+R���Č�o�0�s2��!���p�b%�T�[s�J(�LQ0� ٗS>)z���7"�@�)�c�e�A%#tZ��SS"-�Rm@&@XV2	2w�	;2(�T�VJ1+�D�A���ecZ�rv�Gk�H�B�t�`P�e�#Z�����ŬZ�@�X�b8UnZ,�u _9I~��'�G,��{�FE [�Ӕ@�/��"I�ScL���8It���'��D*��c %#��M���5V\���2�IGy"��A�Tm����5%DA�ȶyPBi(T�u>Ic�!��0eJApǃN$F���Iާa"��F�Tq2�p�A�\��Ij^J�Ts�J�|,��P��H�*!{Qd	u?I�i߱l�Y�UFv8����p��Ӧ ��7�T�Qt�C;j��aI�	��o �ӏTCz��{�\%�!�P
\��a�CF��0�
Փ�g1���E�4=i.�R����zB�<���T���� uh'�Vq��X#&�X�&EI�U�4�X��ia�2�)��h^�)ƐC��L�l��O��p�R(BQ����lV�{V��e�Z�K�4E ��K8�Q�����V9@��ł[�H�2U��J:����T �}��y�/�VyF��AY,Lsa'��P��Iŧ����ڴ!��{��A�/
PtX���X�H�|u���$� ���!a�¥�O���P��"@=۶.�R������	�
Lb���0i��a0e�,3N6,���7��4�d@����C+}��qC�ȑOH0�L��5C, ��2�� ��I$[�)zW"Æ��FB�a�t�U!�#up�p��Ywo <+�f�$Y�	:�A�
$ʔ�`ϟ"��&�m�4)vJ�0)I��릅�o�Th��	 e��<�2��m_.�EzR)�6l"��q��GVf����T�}�"��c��*�Ra��W�(bJ�7�B�9$
�*�zYSj�>�u�'��P$ �J�N�aT�xa�Q�$�@�swI�>'U�lDzR�1)qJ���ҐU�୓TH�,y(X��jV�D�ႂ:f�SF�'�d����ڭ/��S�1ev]����;M��2h��j�1���&�v٘e��.��i�O�����$�>� G�mp̸�-Q%�d�
�J�	��G _��(2���u�B�����*���Rv�R�[��P���ũ-|���k_)e2��J�7tT��b'�
)����S?_��	�@<�����&X�1`�T�PX�ćO�JI1���L}hP@C4�4�T�%P�)
p+U �@l��^�L%��C�>:�z`��NR$j�,����U�04���5i�6e�V�K�'-n!K�I&"X�D�`Ӱ�@��/s��1���6\L�!F-�u�f�R�@H�#*d�-��i���\ '{�����C*Nو�BW�.WQ��8D` �^.>�F|���I7ʖ�-TH<j��[�B=��[X������3	XU��y����5K�N"&e ��$(��X��i*Q)B��>m��=BЪݐ��̖X�|	�kV�8�n%ٰ���8r`V�!{��
"!·�,���˝�%b7=XL8L��[}\Ź������4Sw*8F���g@��]Y�6-\f�Lu;G�Y���3�˜8αA�w��8 r<���]:�L�K�LE��S�G���đ�a�U9c��T9d
9#u,��`��;�B�#V퍕B��+RGM�f����c���țk<Qa����Z1�DR����+�B�G"�Û	����bZN�$� �_�G�$yـ.,�U���g���R��ۅL���9NP*�C�‰<���0""��n�4��5K� �����a��Փ�
�R�l�6]Q��LØNa��{P�=?��E��%�$|�8���F�?����'Qi�7�BJi��S �ڼ=��]�qeP�?�DQ��L�A}t9%ˈ�?mh��<)kH�;g~��3��r�@Yt'FU���C�W=�H�bh�k�� ,ю!�,���lȑ+�^P���"��X�m�Xǒ0�R�o�$ʈ"��0��A�e�üb�(��?$z��Xc)޶Y"�{F��{}��ǝ�3��I�E��=a���GP="z��(�N�*B�x��">C:Jx�&Ɲ*�j�bD�V�}.��#�'����ģ����i��,[Cb�b�۝J>X���I�p����d��!����4cĝ���)W��/]Ht�q�
�zNpYg��I9f��[�q��I�EDB�Y j@}Q�	`ae�:�L�*_�1,,$��.b�
5�+}#J��T �<��� ����VȚ������I:�KIގq���!�:/�,7�2,�H�[��QE�g�н��HB���I��@�"v�I!�
\�i�&��H�+
�:��AZ�[j����+��PL�?J���5�H��J���+�0����D��@��h���Ґ%��8�؅���!��ϔ�4!���	p�u �i�C��`�YwAx� V�]d`JfGQ v���eo�)��tH�	+�vH+���Q��4���� ��3�K�o�2�	?W-�iK�I3!�� ���"�b�c��Y��� CR�Nn�-J1I�T*��rS��idfƶr�����|<J��$�7�ȃ�jG�/F*�H�f��'�,�Q@N� � ���	Ba�h©���$� �!�x�:�Df�4$� �qp��!��'��B�իa;��r ⁪w������$�v	U,L)R�fpCE@�Q�!!ւT���C�J�#� �f����Tyaf�.;6�� B�	�j��͐�Dc��F~�^ 6�
�X�c�jc'�^�(��Q12@�)]�sv��2p��ɂ�"<�"A�a�nKG��-��iQ�f
%��EB�` t��l�#*e�xr	�O�b�Ⱦ�0=ч$�
j�q�`�e��)3�*K�{C����ិ�b|9&��1T��@��$ˈo+�D3��6o��RW��["?��ɲ�:"2)�榟�G�T)Q��'l�iH�O�w����M5)�A�-ݑA<^�q��8��43��0�1��vz�AGf�¸����"'Ș�q�va��$�8#li�D'[���z�'$\���(�ɴt:T�b�ȍH�0��U��
4�Ls�	�+#s�(p��H�N�	����b�&�*2g�Y�ݘ$ITR)�")ҩ v�$h�%��K�@��'�~԰g�Vdep9֥:M(�녏x>|��f!eW��ca��>[�h�觃WY?�2�]	$�Պw���V�D�4kŗ/e^�$�}ƺP�ʁ�J�Pl�"�,E�0��'��@��Y��֎[&B��t��dj�1)��]� �p���bՈM��ɣy��0��k���LDJ�䘱2ʀ �M h�� gH� ڨ=��c���Ty�Jrs���$���|� ty��0b�u�[�oZ� �35��{Xz��
�6&��51BA�3Wߦ�Ї��H��a{�ې'�![��~Pj$�t �y�HP$��6I��ڤ���OP̙B끬4�n� (�<k�x�ad�D�-��z�� �E뵤݉y�T�� h۸7�`��S`ٷYF؝����	���;3G�= �q��\�|�F���Ț;1�t���'Dn���_�]T��pa��;^�DZW���j7�m�!T��h�C�&pHx��6�^W̓sIp��vG.N�h��2�T�*:����Ufy���(+[�R�:TQI�Gݯ̈Obx�D�E�_��APDdI.g� ����IL��I���y"�ɓ	�tP�� � [��A �D,a� ���ǄHpU
 ���Jv� ,ΣG@�z��$��B�D'O1`bց[�49��ǉN��؞�m����@�8~�$ɤ�ʏ y�4Ȧ�)H�����	�O
�� �O���T@�:zr���DE��f��ȍf��kρ��(O������h�0se��Sd/AkIZ����̵$.���q,�M���2���a	�l3"�����L���6���85�-�3韼T�f���`�f�[}��9Nǰ��XS㊗9�M����>B��Swv��Y�k�2xٲ�k�s<���G[R���g�i
pU`�`�M@�*_&{x�LE��5��d��?��A�7��T|Ex� .�I���ia.���:c��:3��̈$����!�ɋ�1 ��c�)��M��Q�ٝ���*C���0��ܨ�L_�q�Q�/����� �<9)�HsW!�z�L���'(�@cw�;qp(i���[�� �A/� 6����G"�f$�U����R,"ȑ8:w~4Yr�0Y��<�q�ţ3���3G�5��!fL]$IEnUIt�GF����"B:�(`",�so�P��İ ܸ��b���G���J���L�@#�͛-+����jʭN�|٤+D1۶��"�NF���Z�4�B����3N�3g��/=�F4�go/g���Y�C��a�<�nL,]��@��^�02xx�tM�w�*�3�d�)C��4@�F Nߨ�i��'OЌ�*΁1a2)�̟�O��s�ʆ�V�,h2�lH����y��_�U�|p1elåv�q(_6,��c��iO���
튍]N��ҤU�f�N��tAơYۺ� P��,OX��d%d"��t���g�&����ÔZ�d�Ab&B>N�h)��yV.T����oS�R���@�^��~Zc�H���U�Cg�рdCُ[�n��
��v���k�{��Z`f��3r�I����v�.�S9��@Ȍr�*��c�$�T�Y����"}2���:�k��Rj��DMH�'KҔ v���>	�[���M�'��SmJ��� � �&!e�� �qy��\���)G���{�唩PQ��@`�:@���FY�6^L�U��'�C���~���K麻	M���"��bS�d1��	Z��HKp  �O��Q���""F��0��ܥ%EpPAuQ�!�'Ɛ�$9	��JjyB�H�A�'�X!b\W���A�G/zx)��#�Oxp9�C�!�՛���~�(DB�*�9@�^$À��=�x��Z�u�my�lMe�|���A��O��ZpG���.˅S*��5�u�)g�x�Ѷ"OYja�@�"�n1��ǌD�2�b"O^�h���8^`œ$�68���"O$b�� f����L�;J���"O,�90n�=_��X��	2C�H�"O����	�\����^ p�
�"Of�za��c� 	�d��(|2�YE"O�dU���R��H���2gi���U"O܀8��i
D��O>:F"��"O���âX�0��*�!_����s"OL��� FI��!
�d���"O����y� E2��Ҝ$Nn�� "O������mj~P��5%���E"Oڈ �&	2 ��⡒�G���S"Or|�P����亷@N	�M�!"O\�H��\!����˶D�n<�v"O��H�!L�c��Ux�J,�!��"OBw�D�6İXcm�;:N�!3S"OE'�2X�xE��=i!����"O��P��:�	R�L�<��f"O�ū���]:��Q,�1c���"O��ui��%bqf�-9��8"O���V��B�\Ȣ�&�K�>Uʣ"O���H8�AX���1r�
U�"Ox�j�nN<.��C�i�!c�E�"O��&H�"������
��0g"O:��� ���Zu���J�hQ"O�H`v�� PH��P

�^-�c"Opy{�L�+�Vt+n�%�T]�"O`���� 1v��l�o١s`�Z�"Oʌ��@��%�P�e/��rGVU��"O ]�7��,V5p�I�8,DP3q"OV�8V*�3u��TC�&��c��,ȡ"O�H����CL�-�u�ۿy���B�"O� �����J/�A�
�|,ݢ�"Oꠈ�*#fB�A�jL#oF9�"O��b��̏*;�)Ӥ1YTqB�"Ob��t!V9�PY3	O���"O8\���+d<b�B`���4"O�m9�ۍ]T��uc�""�|��C"OX��ԪV�2tT�S�U=u�h���"O@����ґ�7#L��v�H�D^�<�q!�+0)R!T7��a���^�<W���x�qG�W�\�>U�K�Y�<�`�ύ*��u�1��5/�l�T��c�<YB�_z��	�7#ۍ>y�]c�(�\�<	��$aR������1�s��NG�<�1�ۭ#1�PK��D�X��P���C�<��K�昼3�Lx�x���"�[�<��B�
t?�	�@��T�v�L�<IVl�&\ Q3v�	T>�����L�<�F9�ҹ�6�ɢ]E��I�b8�C�fZ�'�r-@����8O�!�T#L$���H��P#mp9�"O �s]3,�pE��]:)P�Y�`���@q(x� ���R��S�Z�d�i�+O-UǨ��`O��94C�(�����A�3 f�����&���2�ܞ/��!"�^)�x�0)0�)$��>`�"١E&P�J�v1ƣ�%q���dɜ:��a��E@%y6i�������'��;\
|h�x�N1PmL�0=	UB0b;JH��%U���� �B�''�ƣ��o) |R�Eۻ218"��
�q4�L*0t�5ZԄ\S}�u�ȓE�y@��1�2E��F=d,ϓd�	���L�r���fA�@�Yx�,P���OZ��FU� �JE��I�W\���'*T�� �qn$�[���}� Q��×T�Pw��9'�y�� �����M$qL�O ���טN�h5`Tϒ�W����>a��%@��#> Ä/L4|�R"�C���� .A��B cs��.(45Q���	�| ��2�HO���e旗��4�I�O�h2e��508{b��#�HO�"�B%
]*�� �	QA��/2K�2��Kv�p('���Є��1ʓq���b!��Ir�x ��$� ��z�E۝H��*e(F��y���-tR��ᄋ�(T�x��Äɓ��b��I�"cR��(3<l�YP&*�d��9����-��Zd����OZ|A3'�����@�I*j�*�Zt!1x�e��(*��ԷU�`��K9àh ��U!E@yK�IV �y,Ӣx�(�� L��&ԥcf� ��~b)�ce|1 .�2 &]ExA�%)�"	��.Z�d�B�) b�> �]� ҇,�i16��)��[2�$a u�bnۗa�V�y�"�<$�]:� ��5fe�W��Y�ω#prYUӽE
�aXui�P�'�(�!��K��p�������R+�,�w"F�r4�q"K!�|͹2�A�y!n�CM�U%� :�(�/������u7D�O8�%7�3T	D�1}�3P����DR��O���s�]�'�8((4gS���D�Z>��hB+@u21�ش@�V�5f'�f���d�|�<����,Sf�X:a���C�����ꦹ�5*�޺[c��$Ў�c�Q�֑7*���p�cΣ�05ڔ% y�Xe��	�u;�<q�x�%R�~�Q�T�E��$J��֨mP�)!��.,G�e�� с@��t���ij��$�)hT��(Ӫ#=�v�Ɉ0&�u����= QD� ���?����܆Nn�k�e��f�i�c+K�e(�E�dA�� VD��ƚ�<���(�Lz�D��C�V�nѧ�O11���%'�I:ў� �GU>XB���L=m�F�I({�Vt�W�;��9J%�J�J�D��G��x�f����ܠP��$�$,�*}�Tt�7K�:��*���N�N��w/�|Kh9�&�l�� ә*p
�'���p�'1Q�
�_�hB��NL &���Q+zF~�U�*#�b��AW,l_�쀰�8U�\�jb�׾-p�&��^��C%nŪ"�hŋ��.iV����O�	���]-y��	��ո1��i�En^ ;�݂W9O\�;�O�_��)�Ac����1ċ�92��E�Ŏ_�1ȸ�`l��*�I���+j��u��͊	���	�hB�0�*��.h�ؠ�P�	�c^RP�g�@�*1�#�0Y�x�e�Hx�('A}�a(vK"̨��υ'�YRT'\`��Vd����i���Yo0܉�kY������eܺ�F�]�'��d�C+3;<\9)F�18˛v��7�3�+�*[*���vC̤Z�R ��@?g�(���"�=k<�P�En0�[F+�*Z&���I%�5� ��k�H��򮄥����H��N�'���32���'<v��-�?Y�S�G�����*O�r��eFA2 ���N[
�L��Ҫ:RbPy�����y�p�'��#5��6
���P���\����aݍ�^�����՗	0R�0�GT-�HěF יJGPi� U�S~L��b��nj��t��
6^�xeǕ�(�DثV �F1ꕱ)B�1<�;��v���c���Z���� >�1g�Z�B7������z`~A�V�J�>KVT���M��Z�`�V6h��X�c���M���F���m�Lx��Ȱ�W}>�І9���ؓC!aJtF�I�hq��9�
	Q�⑤@�jX��}IP9�6���d�	�$ t$��GRƌ�c��!|���̘>W
���͋:�9HB���o�k e �KR�qc's�ͣ�l>Q��wЭ b��m;���vh��}4 8�Or;��Q01 �\8�肸�J``H?�����u(N��C�9kZ�'���f����d��>�������{�ziCF��K�����m@5���ֵb����D�h>���͘$hZ��q7�S�U̪	�7oS�.֖e�&�؛v�<B�L�2{�,ם�c��a�&�"J�J�f�<O�t� �\�֎�-!\��c4J5�n|Y1�K�j�N�ҥ[�G�J@�L��T���ϸ'V,\SW Хg�����ُ]�x�2���9u"fn̼hՂ��e�)F���c@P�a��ثfM�_�|�"� [;
 ��~���E� -S^�Ԡ7h͎3��4�gk�;Uc�"�}�ՙ�X]���_�02�(:�Dޭ!A�0ER����Js�.��*�D@�Y6�Gj�7�4Q�R*��WE�:@E�z������-��b�w}�8��Z�8�����M�<�L�h5��*0�09$�N ��T�~�C��o��`�ֵ�hN]�M;���DϦo��P��=f����	�6J�h�V�lW��#��]�H1��(ӄ��mԛv��"�v�[��X�Q��H�h���9T����]�|��'"�p�s]x����\�`�L�'����</:\�be�F6O̬���i�S]������(S|~@�D��k�
�)��	!8�\�y$D˧�`�h�F��vⷬ�EG�h�`�ֈe�d��@���}�V�i�dJ%�~�8FI.�f0�,@NƼcp�[�HHE劉���6k�Aj9���$�	-&���0�*�$p��M��t	�P�g���B�ы\�u_"iRCVxb�$A�m��U1'�&2I~y��fO�V�)�K\wZ0I��{g�@�P�ÑoF�m�NO7yz�2��<���ӻ?��A��k�^,P�P�[iX<���=���UB�
��a��c��=��lx��<h�A�%��;l�S��F:P�sF��_��I�1��?��p84AC�:e�m�0�����M��0}����,C#�̞��H[�6d��P��00���`��6�&]�!W>�{#�\_��P�ݎ*��\r�N��#��Ue��&/��h*!NT7!�Ƣ<��Y]ưp!��<J�֐h��Zu�R�y3-�x��D�2��� ���6��)&^bV�!��9e���f���8�[��=6�e����n��6� >t�Q��[Gˋ*9<�UJ7���h��F�<p�(�qP��%{��e��12��� �aJ�2\��[p�R�.���\'}���N3?�9rU���\ʔ��L���UFT�N �Ojl����,7�x ��X$y
Q��$_�J�cjƃD$������$f�p!�¹%7����־S@�:F��q�&�S2ک6Ex�S�a�k�\qwC; :��n�}~R�F8���"�ä�[���ay|�ˑh�$k(h�*�3^�Pqafƹ���Q�F�&��v3��xrÀ�*���i��F�2$CG��!=0kq���N���!���uE���3�eeQ�هK�Z�ʃh7y�\�p��
H�A��K�:�lx��G�$�:��O�Z�t�<[�.�<�0	�"/�]x#jƵrq����3Q��t1��K�>�A�c��=Rr��$,�*Oa�$QU�1�|�G���Y��0� h�.P4y�+��v[�0������b�ZU�4�n�w�N�\��ʰh�� aI+j� 5����{v@�D됅D��=� ��0C�$_�8Tr'U�T�P�+�
3.q�Eh�&xLeՉ�;Y]:p�!�l
�`g�k���E��:�����N�~2c1�[9]Z0d��Xi �0S���h���*I��#�d��|ܪv���lf���O>W@Z9ЎG/n�z}��Ɓ�O��s5�D��f̊6,�Ԧ1�
�a���PeQ"�,�$�*I�@pXF��_ �x2H��mMT�F{�
R��}8w�	�����r#I�_� m�	݅v}�D���-0���U�S�'��]`���$��"I��T*�a� �f�Hթ�2�k�T�y���0� �#���$ Cq��:�o�V%طC0��(:0��8Dt��6Ɠ�v�4ӰJ�!n�m���Ɵoe<a�AG�~b�N'3�X{S�?c�yp���#N��Y��ȓ2m1������m��	'g�rdY�o�,�jY!t��zY6mg���5�ۭ*�,�EE EԡvƓ
Ak�k���T1��Ї�M3�iE!5�"S��,-9��@�40�^Bs�>����/��-��(w��$��JΠHN���n���8�L!j��4�qdU�+������t���F�ϠEP�BVF]�$m�T��������V{c��0_�D1�,�~Q!"���9<����K�&[ �J��*A�2EC�!ڛ;�N]�]@=�C�F�6M{��Z�:�JQ�UB�|���D�of�l	�ؾAI2:���om����˄V8� ��T����V�C�VTQbb����1��51�Z�!�H����1B���� �d8�YQ�N���5����!FC�)�`��'[�o8�AT�@��Uؒ��'�F���Azr��q1撲DP	Ya�^���G�=zY(�5O�<��mOVC`��D��%~�1�4k�"��PHE��N>|M�g�I��O����՜�Ԡ�����B�+4K�t��m�>D����Yo"�Rs$N�ט�3�������VB�3E�u0d��x��S�	$x'޽a�G�G^��˗Hݱ�a|��P3Z��!��-{��qӠ�Ӕ\����dsN��'Y��>E�U	��]���A6'�/~��Y�`�Y�
%���Fk����Ɉtfv��3GEL؞I�y�����H$��`��iͥCD���k�
c��s���n��D�p$�x�2�&@<ئt�V	�&NR����
b��[�ʷk��5�3,��!c�O���a�`�$Ϗz�U�%��=��I�E��y�����/�X��������%~�,�C�ɞ3�M��GE�\^t`�'�<���ZvZ@�Ł�'y�"=5�O-w��҂�@LF��A��)P���2P/+s@���;^L�R�l,u�ם�E-Y��R�P=���7"x�0ۣ��bЌ)� �4#�\P҇�3=Ka~�d3b
W�a�1�d��$D��y�ƀ!q>n\y6���WCK�d�6m4jw�e� au�\9��;s�1�|E���ʪOq�Q
�!�+�0>�,��	F]@&C�X"8C�iǎ �rr�m�7#Z�=@�ð�l�P`V"c��d;��^� P2���zb�-n��U���c��"\B:�0/
R����:�B?�A�Q��:C��\jb!�� ���5|��3OA7�E�r�-��$0�%:1��`à�.o�=��L� FS|��I�Enݢ�i�f�Ñ�;x��AB�!֯~� 1��K�?r���gJ�%GdɊ��S��n�ӡGM�|��i:t��=%b� `"��/qn��Ʀ�1(��B����?��F�lm���]�P�K��&S�hz�-Mh�	8q��<kpQBUa�%P�.0�&������@�[�TY��Ե(�y��E�rp��PG�Z�]=�hhflʬ��9�'Ġ�:A@�wy��)U�>�;�E�u����w'�5D�h�vV�$��=�T��pʟ(C�����[�^����
������q�����v�n�#�e��t��l*�z�/�;���稒.����n�7g(�qM���L�:� Đ_tΜ"�&@�լ��1�T�qN�u���2n4�1-Z��@���$?�"�.�*X�@A3(���J*��,1`����C���r�-!�6T��#�,�2�	M�~11e�
�`���[��xy�z@
�:����`������� ����� 4�KG$�,�ɗ��0�L9�!#R<!�f, �l�~R����)D��g��v���J�Ԩ)BԒ�O���]r��U�1��|���A,(��y��2��L�@@/-���bekG�FJ����	),1,�Q`hϯT�r0R��<r>�������ReKǣDM��kgcȪ*>6��hέP����B�٩�'T�@FI��D�k�68)7�I�'��MۃO�*6����C�qSV�&�0&z��H�.8�u�嫄Xl �"�!�N���%Z�L$��C2,h�Ar蕭>�U��'���*
�l��CK�=x[�����Z�����W?9����EY;O���Jm̓L��5!����V/��4C2B$��84� ��k���#ÄR#A��<��!�;��O�$� �A+z q�DL�K}pM��%I�
�haD���y�G�y[���hA�E%` ad�MrrM���	������h��y�0#\�\޶Y��g���M��?O����-
5;�����&��qC�§�h�͙XO�MI�.6�"p�1��Lۊ�ᵄ��'��y�O�X��͘]C�q!��&���k�f��d�ߏ�(O����K�jbp*�/.>�y4KS�|8d�BfɍOԢL1e��<�:���G/M^��Є�˗Q�T�c�x���,���g���,��i���)O�b.������4�6���Mcs��7М K��ܧa׬e��哟2�L,#��0�ER�-P"�m�; t�2G�1c�F� �=2J����*p�+�
6�W�N��<\���*ғd/�]C��C��X�l�=V��Q�B��W'��qD�كw���3��`'�E{�Ξ@��H�LνU��qv��G��Ԓ� A%^�b*A7z�<y�i�/�d	t�'�>q�Iͯ)֦��䝻5�t�{�׭s&p��-{!a�Ό��N�����٢@�V��p����.��Y�؉ �M
�h04���'�,���˵M�v�|I��'�j��eKb��A���Т
ԝp�a����CAH8R�9�P��F�����8`���#ځH��ߊ	���[&�|�c�3��ы��;и�pvB��O�M`�(G8a��÷��t�e�Lu�f�c��S��)�B��_��0�����e�����`M3
���Pq!;�?2�K�-�x	㡠��D'"�R��!ఘ�"�ֳ�����D�l@�hܧ7.!Wգ �<$�iν]a��!�a��_AjZ��B������}�����yOq񡨋;|<]�*� �*y�g$��]���@D���	رL��yN}�qh
9�~Zcٔ���/��MR}ȒnM�1\�8��tib�����i�Vy���@�H�
P�B��ev)3c�:{��$��.�P i�07����H���0�{ܘ\�pf�4(.����<��pt��۔L�P�)�'Lt�a��;l�,����81�u�TW�����V�`���$?��fk��P���dn�M2���
��`��H"U�Z�O��`�����}�%��hb���r���B4�>-���J�7��� ��OS<a����)4:8�m׸d�x�'.J���a�j��)��S�� �B�1�'3���ꅑ
e@����kQN�
	�kSJ��\�@�u`դ�2R�Y�,ĉDT�� �9$�4�b�NWr�a�Ƃ�j��Rv$%�-'��d7�'}n��"���&2F,@W�KNB8�ȓ�H)���p�q+Q�������H���4��^h\�b�\�6�X��!��|P��%I|��@���{�Ҁ�ȓ̆%����K�4]�"A��n�]�ȓ ��4C�/;w�&��uΎ�U|tL�ȓ]1܀��ܐ2p ��ˀ!�Fq��g����✣/o+�Iaѓ`c2D������!��1��![���r��0D��)�ŉkܺQ0�O�!~+��3'B/D��RMj�J�V"�)}���[��6D�@���	M�֌KAL��N�p�Y#2D��sb�T�p�;�P�WdI��C2D�k&!P9SF<�S@�&Lxx71D����c�=#��Xk�nA4T�B�	�}�����Ǘ�r��(�D[�kb�B�I���!�/m�,P��K�h�B�	�u�ЈE�܎  FAA� ӄB�	�# �P�3F��;-<`֕%��C�I:=�Yڵ�^�!+�5B�����C�	l�<C�y��0�THWIQ�y�	
�3��뗋иx�V���Jդ�y2䇳f)�i�vaª`lX�8���yr@&R5�C�B< }�5 �	՜�yr�˞}Sz4K֥ڛ|����Qb�!�y��@"X`��)��h������	��yr�#!'�(3��N�k�N�;��H(�y�ˌ
+$̈�T�Ew7�1T��y����h����kͦY�6(c2@/�y��/Y���*D�)V��� ���y
� j��G �?o��:�D�(�Z�2�3O�\��-$�^X�O�d2t����g5b��Dki���@هvJ��sFF�J�t5xI>���t��V2��ͧPp�]�G.K;X�� �g�nl����{尀��%\�by�t+��X>U���K�a��L�.F�T�mqR* ���D����@�g�$�,Z�(˅f�H�� 싌�	�4���?E��6B��1�f��x�00�JK��M�VHS����ȟڵHB��)���qg_�E~H� �K�'���Ʉ�I� ��	m���Ŏ�;��O&h����O��;��w+<]�.\�q��c6Jěm�bD%�hs�L�7�qO��<d�A��k�N1I��E=k�m�^�X�d�	n.qO�>�礑b8A�6܅L�l#P�tӞ0Z���S)!����Q	`�(uAY�r"�m9��ЋK>�b��9���O��M������ �.T�(������:�@I>�зit*��yJ|*�����JJR+K�oK���G��f.`�)O�)�w�_��1{�"���N~24$�.&:(��&[h�z�Q�N���?i�c`��`�OQ?	�+g��H���؟z5�z�C�/l\5x޴	U�'��u��S�Ha��s*����I �ƿ|����ۈ���*Q���0I �OP�$�!���9�yK�HK"�u�l��S�$h4����2]bJ�`�.h��˓;�v����㞐*  !���ó{f���'JR>E�P'��$��R�*M�{*���'t�Ё�N��D��fW	cāK��x�6��1d�S�I�.��N< �ĹT�W����9SY�a
�l�@�|�Ѯ�<���~nZ@2��-��e�Є����9CׄߜrI�C��&
L��߳tL��!�䐾T�a��JU�
�Ydh��%\\��Ү�	�?Q���E�(R�兎-츙�çw�B쉀I��ERH�HV�ژ6;�ys7��a2ߗ^�z��m��Hc`<��Ȑ!�y�a��sF�@�-�"D0�	L��y�C�c.>)����nT�Ԋ���<�y�iU��q���o��*U/�7�yRXe9�E��g�m�(��`G��yb� YH���12}��NЗ�y�P��xA�T�g��a�y2ƙ9+(����1f�$)%��yrNԛjg�⣭�95�"��"�y��L�$�p�F�A!4�4��ZQ�pB�	�qM�p)��8K�T	Q�+\3gB�I��n0C�L�C$L�#��,�C�	�~�@)�怑�e6�Zt�R�2�B�	6Hsjt���X�u7���p@P�f��B�ə}ް\�ԫ�,1O�)J�
D��B䉉=�!z�!-l�m bʌMhC�	*K0b\�Ə -��"��
� VC�I��!b��9�`�*�	��>C�T]r8IA �yt��k�5�C��>����.)+',�*�	�5V��C�I�o�8�q�ǔsL6q ԉ�<y��C�I�s�^` �AO,E:F肨	s�C�	�ne^��(���ɢÂA (ʮC䉱1�b��T��9��T��S�_�vC�	�c�z`�� E2�@1�)�d��C���PPe�0��<c��͐#a�C�I�qX�H�/ ����"eصRC�	�4?z�e,�I	������pw*C�I�><�H��'���9&�F�, C�ɪ_X5��
ˤt�����IO�lM�B��8�#�D:b]�y��P5�B�I�^}.I�7m�a���8��N�h�C�I�w����ܝ�b�N�zT�C�I�qf°��[7ߦm�)M><�C�I�BG���h��`�n�h	�j�C�I>b/@d"w�^;� 5����(�ZB�	�5�6�ӳ��\ΪЁ��ǋCK�C�I�+_<x8��V�!18�HC�I+)����ħϻP�4�-M"c0C�)� x�j�.�x�0�_<Y�\0�"O<�a+^�rE��(���|�0l��"O&��1��&y.< �B���a"OJ��g����G�G|(`"O���&d9��������ʖ"O�i`w��(6bH��!�ߥV�dA�""O��坭q�
�JSf�N&�yb�ƃG����j��BԬP�taB>�y"�ga�-R�z<pc"	)Wm�9
�'�6$[�'R��.8��m�#= �
�'TeYt T�V���FW�)��i�'b6MX$��M���G�wbi�'�:�����g�xJ�,P��
�'�>�E�����j�Xd\�
�'WV��p	��r�6L9�W	��Dz�'{���	F>���,����p��'��l�
v�� �W� �Y�0���'`�T���l˴�X�L�W	����'�2���>���	q�F!W�j1��'�P9�@�>�p��C�)SG�u�
�'�H��s(ȱ�Ɂr��2 :���
�'�蠉ET�r�Dۄ�į�JI�	�'�N�C�NF1m����ť�
4�D�1
�'ېY�E�Z2�%p5.�%,dPs�'ڨ5���a�&��J߀) ��
�'ľɐ��O
zF��d�L�<�I
�'@d���f�5�\�R#�֬܌�X	�'��USO�=��1��U��i!�'���)���B���s����J�'��]�Eg�:!���iDA	(I`%B�'@��qGK0����@R�5��
�'cP��Q�&�c��\�|p<�CO�<y���3.����	�F[�����N�<�"��.ri�O_�H�sk�H�<Y���h�a"K{"�;�b]�<yA�W��&`��ܔ\�p�{��a�<q�Zf`HhѶ!�����6�\�<i�>vQ��yS�� e��)C�A�<Y,R23� ���]R�$h".h�<acH;#�$����:X���1�d�<��̜�9V�.QѰ�2�*Ĳ(�B��-Ζ��4���WbNE���(cXC�	4Y/���D�P&| �Ec�b�(�2C�	����5B[���jD�M��C�	<��L!R�'|����͋*a{C�I�����t'O��$Jz�B�	u�} re,|-��u�ȌX�B�I� ��U��EF*g�( qkǒB�	;"i�R�đ"+��T�X?4C�I�Yysϝ�5�����bT�9�C�|����QC��E�n�6���B�	�O]N���#���ʃ�˹i�C�ɝ\�ԡ�@ZZ�N�iv/Ƚo�C�#e�fy
���>�L\Z5�.QΎC�	�UG����V�@,�uO��?��C�*����'obԓg��W�rC�	8k��0���`Ll:�%��zC�2�rš�dن.J��W�!B�I�S�:, �L�Z%&Ia!�9��C�{-8$B���7fi�5�0��C�Z��%�7��&vRq� �=O��C�I�~2�:�՗Tz�C �"��C�	�)�Vh#����Oqd����ӴC��8�&�%%ڃ_��e6�P�Lh�C�)� p ��C�Fڴ��U�Ī{mz 
�"ON�JVn	2f�M���+~N����"OH@XD
�#R�BMH@�P(;g��c"O0Q13M�Φ<З�R_�:�B"O�Ma��[��VcY�=�ԛb"O �pacF:;>0p��OB����hE"O茱 J�ttr��V/�X�}��"OvL��c9P&=�n�SAfD�R"O���1��[�h*�F�n�"�� "O"�`�.�4��a�	^���H�"O$��E�I>, ��⎥~����"Ov��eI��8y�
�2p8Q�"OX��G�ƥzr��blii0"O4��N\86I)r�
�5]�$"O��8U`��>���Y,rV:C"O���S�}j�B��X���9#a"O�ș�չ3��|Xѭ�h�����"O�D�4e�1��Ta$b��
�0x��"O2ku��J�L�a���UcReq0"O�(�Q��Ō���.V�,��Ԙ�"Ob�����YB(�&��./	�`�g"O���٦dC���ɢ/�4e��"O> � /o�p�QfS,1��X��"O���@Y���3 eΧ�~�i#"OZٱFe	�n� �;2��z̴h2"O Q2I���<3(�
R�\H��"OAr�S�O����c(���q��"O�a@ɜ0"�d��F
���"O�I��E*+Gt��6e�l̄��"O��:�Ǉ F�l`�!�8C(��"O���e��,��������£"O����iRp���ԪaJ��"O~����#r�(rD��3-�P�"O �� �@+w�D�#ϐ��Eza"O��j�$Ɠ����U��!.	�i�'"Oz��aӕI�I�0#Y^�T��"O�-�C��J�4����	�X���"OT�85��>x���q���FB1[$"O���B%S�X�ŏ̴P;� u"O`���8:zp���OÖr)���c"O�$s
͸/� @� F�n�9B"O�"SO�+f@�İGE%u��a{�"O@���4NU88P�"�+��`��"O,��3p��h�!�p~��c�"O�� '�u��)�ª�/b����"O��+p��6��Ȓ%7Jj4�"O �j#"ݧ$�J��X�Yڠ��"O�=P�G�ڸ�&��&uk���"Ot�!ŋ.I5:�0a�Ak,I!�"O����l(|7���E�e.�dCA"O��s���.�T��P�O�q�B�#V"O� ����=~��2���dM
��"O��P�XH��b��a*`;�"O��)i��LI���,K�E�5"OH�Pe�
����M{~�;�"O�,j��'B�(4���. rqQ�"O���%�,&qr���U88��yA"O�t��}���6 AF-^��"OJ�s�A�2)�9v�X},F��'�bGQFt��c��=<+�'I�$XEB̥%���L�qݤ���'M�tɌ�0������fi���'@�B�/L�/v�z�. t`���'��Az s
��A��
�pt�
��� T���S)r��`@�W���p"OR�h�k��J,r��a-�r��}s"O�e��	��k'�� ���x�"O8TAp)���"&G�"��5h%"OVMje�k��E�G�j��C"O+�۸|��D�Rm��d܌{=!��M{f�Ir�G	�&Hh����7!�D�!J���#��q�lp%��!�$�g�b�q"��b(hyA�k�R�!�$�b��YD.��"d���O�U�!�DخpC��yW+����I�j��P1!�䐧#z�P3$�-0A�.�i"!��Vn؊��
_����� !�1�
�)�Ũ 
�BmN�I	!�Dǃf9��0y�|�F�֞_L!�d���L@"���`�(yCj�;!�@�tC�ᡑ%M�"�l��2'�%�!��#�6!�ć�l8��F��!��ο5��y
�虻\���9rf���Pyb-U \�St+�S|� [��y�E2yJ\%���E,���	�y��(���0��h��k�NЫ�y��]%Lq �ҵ��:�0@�3�ylƈnŴ�f���Q	wM[�y2����(5�N�+� �׿�yr�������6c� �dX7���y�,A��y��S,M4���.�y�Ԏp��eˎ6vV�Q-���y2��ML�l�%%�,m
<$٢��yңF<s�6eq� L�a�n��B&�y�ˇ 0  ��     �  �  �  t*  �5  4A  �L  �W  �b  �j  �u  �  �  d�  ��  �  5�  w�  �  ��  Ӹ  �  X�  ��  ��  A�  ��  ��  f�  �  q�    s
 � & ! L( �. 25 u; |<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��Inyr��-qd܋�FS$��Q��Ԝ�y��˪=7&}�)@
HZ����2߈O�}D�&D�=��|{�A���تI� �yr
��l����k��I�a@�e}��)�'s�T�:g,�(5(�K�
܀$�ȓJ�`�6 З`C��[��84��5��2��yr1�L�E�F�`F�D��݆�n�,m Gˌ�ZQ����<����>^�䨍��Yt!�:U�ȓ_��!���8%Kڀ� �>tp��ȓkb	�q�+�Y��K���@!��czT*��}M
� �+�ifN�ȓcA�|�ҏ>	W����g�n�|��X��B���n������01s���gE�j�:���A  8��K�N�2G�U,q�҈��˅�/�<��ȓ^&N�ypgR�[Ěq�Q�lg����T;4)����j<̛��)�LQ�ȓ44�����gP4�&H	/e*��ȓ�hY@�A:�����
�az(���2O��z�L@*_u�TA��3�2���S�I� p*���&oB�U���J�~B�	$1װԑ�H#If�O�9 ��"<@�)B"�@$a	F���f�©h#�^�<��f�([803"��(S�I8@b�H�ў"~�)� ��h�.ב9���i����<�Z�"O<�K%	��6��%�g��&r"@<"C"O�ёe�
�3c���w�"���"O��B�&�$�F��@΁��H1)R"O�h#���'������A�
�W"O�̡���9��f��������"Oj\j��O"� �Yqa &ct��"O�Ђg�pj'���-��`"O:��F��Jɷ��Q�����E�G�<!Rl^��-xAA�����4�M�<	���*��cfچ��;�d�<yb��
'~hU���9Q��ma�<�g�L�K챁���*2�6�;���^�<��KݻW��U��I�#?d޴ˣ�C]�<���#@����fJ�w�ΐ�aO�C�<!C�,?PnP��I'GAT���C�<���Gi(���G���5���:&�YW�<�2M|�1N�w���!*V�<�n	�h��#M�u����%�TH�<)V!Z>~�2��䅉7[ ����E�<a��ԭJ�,Qk�B�1eoܝ;0�V�<��f�o�zE��,&�h�q�SO�<��Wa.zT��Ä~{�xkp��P�<�d?^���Jt��>s��h�N�<�p�1P<Y�'Q9k$0m8���a,B��=q5�X�R��,[�!��mU?�z"=���T?����%�}��ԀH�P�*�&D�d�%��'m�<���"�rFL�7f%D�世a��p�z���Ј��"Q�7D�D����/Z�DS�	ΕQs���b�Т=E��4n9�$���[ {Ѵl�r�(n��	���l?ɷ���UIڐU������}}��'fT�!	�w�X�����P��4K�'�P(8���Ԉ0C�L�X�&,[�'Rh���R�Y��$�b��XeU#�'W�4s��L���#����!oT��y"ˋI�n<�e��� �L)�y""W�k.�uS!�I.g,+W �	�yR�	�e�TҧA�����/H��y�Y'7~E���	�T���d��yb��kc\P���Z=j�*��T�y⇒�Q�2�c'�/].x���K;�yR��3c���r/��+s��i�'��y�@3�vYA�"B3F=r��3肆��I�d�a|�L�z���ģSQNd�ï
��0?��+�?y��7?������@��%���h�<Ac�+\�(�ꐤ�`�Ȭ�gb�'�l����i"�h�D&R�lQ�u��x�!�$�gɠ�k/�� �A��8��299�⟢}�� j���≽>����ǎ@�<��,ɡa<���
�8hf�T��b�dQu8�@��E xJ���XǦ���*O<��W��?Q AŴI<�9�"O�QP&D�N��Ȳǂ�o<��y"O����K_a��ǂ�$i�(�4"O�`���M����a����"O
���DЖA3�L���ߒro�p��"O|		�*&Ơ����C7n�������(O�O�� ���|��=��Y)=�8�!�'����w�x�R�dL�<ŴL[�'�
���/dC�5�*��@(z����x;Q>��e�E	nG��Ǡ~���*P.8D��0gC��X�������H
�ن`3D��9�&��|Xc�dQ~w�iˡd#D�� $���bX;"�@���9R�:�`"O���CVkdYY�&[���"O0������t�E>(�H"O�A�I]�<WJ�Ãٳ�J|k""O��A���?�p�*r��G�X�W"O��Pg%Z��X����&'2đ��&�S�	^�Gd	k4�N��ڃ��*Y!�dD� �����vw��[�8<đ�h2	�QڈY�T1�j��P*���L��I-5��9��� 3|���Z<y7(��tp���2�H�fHn�<�A�Qu��e��X�L"8��on�<�5JAY�0�C/� ,Hb�ѴɞS�<�� W�|�v��2;�^h�g@L�<�&c��TV�M���.u��ma�}�<S���!��djbL�n�\�C�z�<�!�L�^fĐ���Y�W����k�퟈�D�)�0p���҃0�,q�4�F(��m����y�ڎ`� գC�F��`����GX����l��ͺGLp�ѡ�1��>���1�y�/�E�0�b�%9d�X��H���yB��+1��Aa�	F���C._��~��'���+}��IQ�gX�4bÇ	�V���p�#C%�!�$�#C�ԥCfG�q'���h��B�Q�,Ǔ1N�YE�"�y��S�D�څ�ƓG_�<+ЌS @/z ��U�<�T} ���A(<&P����jvyH:S�r�<ɦ�(~F-*��J4�����*�o�<��J	.U��4��CP�+�\$bŏIk�<����N�f�

ן]�ZC��i�<q�%�G�Z�a�ph�l_h�<�!)��gOX��цНEKzi�2/�y�<7�3v�E�1+"�J��v�P�<���y�� �-U{��LZr�<� \�c���H��חGjv���An�<��J*p�،3�O�~�US�Nb�<)aFD����O��G�hК�IHH�<���%��=鵬�?�*�� i�x�<Q���G!�5�4�Y�%4�t.n�<	�%_�i��p'��79��ԡ��UO�<i���3��[Ã��VEB���P�<y1�\.z�X5�3������dFv�<�����6�![��0�{� ^l�<�4�J�Q_v�+Q!F_�-AA�O�<Y�%
�ł�ş�F�x�dFu�<A�SK^�zDl8�j�H�u�<�C��4GD���##	�
e��[p�<�'"�tt:��-�3D�6��.Zl�<)��3�0)(��P�6�Xcc�Kj�<���D>2^B�H�&;IH;5`If�<��Q�΢�b#�ڶ ��lÑ�_�<q@ˏ�QRry(
;(F=�G�^�<���k4rpr5H�`����T�<��C8[����F�����fRP�<�d�L�	#��
8�xԺu`R�<���P=�|�R�M��@X���O�<�6bV	w������Vjx�p�#�I�<�%��S��D� �_6zTPp��N�<���n��%�D��4���q2M@N�<ѡg�l�&X���]16��Q.�J�<��E��P�Z�I�Ҧ�)1&�a�<�'��������n�x��ZY�<QA�07bF�R"�C�RS����LX�<���4����bX�V�:RF�
l�<� l��J�&X�tȒŜ(pN�a�"O�MR6�T� Y�!2d��>d2��`"O<Y"��Ħ<����ab�$(l�$Z�"OI��!I!#lXZP4y x�c�"Ov�
v� �Y��(�6F��t�P7�'T��'Q��'���'42�'p��'6�}�fM�AX<�bugҺ� �"�'/��'GB�'���'Y�'���'B6m���N���b1�Id�V���'���'���'y�'�R�'���'_�$��̚.UJ9�j��nPJ���'�b�'\��'���'�B�'���'t�y[��LY��AGżG������'f��'
B�'���'�r�'�b�'�x�
��@U�戩�c���8���'�2�'�B�'MB�'�B�'���'��C���3yk�X�rf�8�4��'���'��'�R�'r�'���'�P��NƜ	6��s��GZ�@Ɉ�'���'>r�'�B�'*B�'�r�'����ӣ�(9��҅�ɃO�Љw�']b�'z��'���'��'�2�'|HZ�X�c֐YS�%�j�&�Cp�'���'CB�'���'e"�'���'�\,I`��Q,0ВG�DaNE���'9�'"B�'���'��'kB�'7����� p%l������*��	��'���'���'���'3��'2�'�X��)
Cǈ��&���tr�0��'���'	r�'��'yҌr�d��OL� �2Q�}j���E��)!�Ky��'�)�3?�մiЎI���E�$��Lp��|v�I��͕��d�Ʀ��?��<���<��� D<^�&�
�d
������?�Ǉ��M�O�>��J?Ͱ��><�vD�C�_�>�\�b�*�	��X�'��>s�Ğ|��z�߹U��mz�*"�M�����O��7=�.Q�F�Z^|��oţO�
H���O��$b�4֧�OI�'�i��$ςA�������0&��52���~���n�k���\�=�'�?��@_4v^Ԩ£>\�����N��<�(Or�O� mZJ`�c����`�x����%ێ��A㣄�x�Nk��ן���<I�O�]k�U���A!�K+@�ĥA������cG�iK��7�"cF�����K3NK�J� �zWIH!gId����{y�Z���)��<a
�6`�Ru�7��5�bh��<a��i����O��nZc��|����Rs�|�C�5�TI�ĉ�<)��?���
E$x�4��dn>5y�'G��}���E�i,,��a�'I^��� >��<�'�?����?i���?�)%h��ą� ��\���P3��$�؟�H`E�Ox���O*�����7�Μr�A���������P�'B�7������J<�|�� P"ԈcϛBQ|l��,@8��� ��Q~��Y�p>P��I�#p�':��>��%(`+�0!�8(#�m'8���ԟ0��Ɵ��i>q�'V�6�6���g�li�`��,k$�S@��e��$Ӧ�?�U�H�ߴW�6+f��E� �.kV�$+$�)]�t�Y��]7�7�$?���f� @��pܧ���@
S� ��X�e��Ki�-��<��?����?����?i��t�3s�|��,+6R=���L�I���ܴyˠdΧ�?��i{�'��V	I�>���B�KZ�6/�!��( ���=x��|r��M��O	H�ōD8L�#D����ˁ	[/� ��:B��O��?y��?���CNzY��T����v�\�gˀy���?9+O�oڱ2�����ٟh�Ir�d��� �E�N8^<r�OM<�y��'y���?�����S�T��M�#]<Q�D�Ӄ�8��p�t��;3��탒Q��82�
T�I<<�Q��!W�X-"��V+S> <����ğ��I����)�ny�x�$��"/]$L�t!��ěPF�4���$�O��lZC�i>���O�LoZ�%Wִ��6Aq�8s��\�bx�Pڴ �&�. �v��� !��>Cx��\@y�O�>n{z��&��-�<H ƤZ��y�W����ID�� c��O��⧠C����4h�rC.Oj�$.�S=�Mϻu|Υ�c��;(	LQbBz#&�X��?���x��$�J�6��5O68�D���	w�I�W�H-S���`�1O^rw�E��'��'������ɕw���q���%���;J��W����	ԟ���🀕'`7�9fP����O���� �@������/Z;T�Z�tүOj%m��M3�x�h�*8605#�>uҀ�;b`�1����?x� V�� d����`K��c���׺W��-{�,��j�����ݍn�!��R�����k�D4�*�(ޜ����'�6�2x�Z˓m.���4�o��j��@ e�U�<�пi8�7MŦ-p�L��	�'6( !ҫ�?�wjEsb$M2%��lh"��4j��'��������ޟP��ʟ���� �j�p���B�E��(ɂ�'mv7-�pAL���Oh��$���O ��E�Z�n��*��L�\5[G��k}2wӎ�m+��S�'i��TH�%Q��R+U8Y(��gyRH�HTRY����'V�	;4Ц�"�I?`�Ε��%h������yڧ*����q���T���P�.9sV�;B�y���4��'�R��?1���?�����S0������@�;�S,.��E��4���a��(Y�'I�c>�� ���cT�T�\"��5	�q��:OD���Oj��O��d�O��?MI"Aݢ	�Rxc2�T|�Yy&�Aԟ4�����p�4�4�*O$mmO��,aKU� �$���`�ETH�I<��i�7=�2e� ,x���i;2XBiJɪ*6C�=�MQAm/���$X!����4���$�O���׃oB5Ɇ�H1KM&�Rd�F:���O��#`���Ķ!�b�'2P>-Cd�٘������6k��yĄ>?1Z�|��Ꞔ%��' �@QC�.��cڼlb��*��� N�Ƕpx��J:��4�4��/隓O"a��H�dD(��Mݔ3���O��d�O:��O1�`�nf�&G�'�fH����;l�(��'��d��y��'�Bj`Ӫ⟠��O$�$�G���8�G�[� p��C���D�˦Q�C����-�'�\{R�B",O���J٨}��qT˂S}�Q�0O�˓�?q��?����?i���iD�HQ�	�!�/��#B�y9���Ӧ RFCǟ������$?�����MϻL3483�M(�pM�J�!������?�H>�|���:�M3�'�6���-S 
�����CG�Mʙ'�2mc�a�ߟ0/������O���U�?��((3j�*X���`⇋6-4�$�OJ���O��*4�VAL�^�'�2+\5dƼ���"f���Q.�+g��OX��'���'��OTD��Mb���@eP�d?��R��4�w��>`9�o�-��'r�x��ʟ8�ޘ%%���G��$���O4D� 9���q0�{"��9l��ٳ�ӟ,��4~h� Q*O@n�c�Ӽ��&E�9Њ�� ��=�sl��<���?���i	��xS�i/����!�П�\�O�d� yA�i;K\	��%��<y���?����?9��?����CK�� $��MS��xg�K2��Ӧ}˥����|���&?u�	f�2�0*]=[$b�s�)9L��ٮO��n6�M35�x���.����EIO;%ĦU
QER)[����FN=e��IIml�c��'�U&���'�>��6I��(R���e�J��L;��'��'�����$Z�h�ߴ\�0z��u|`�r0/�(�)f�b�͓����d�u}�q�HoZ
�M#�S"lg�U� 2#��V�
��J۴���XZX4�����O���?adY��*�ׂE�d�1�y�'�"�'��'+���pj���Ua^��2I�Y���D�O\�d\Ц��s�|>��ɛ�MO>���J8�ᄪ��X�b�(� T<���?)��|j� I	�M��O�N4"t���!����NZh������O8@SH>�)O��O����Oʨ"�-of`�X���ܩU��OJ�D�<���i���'���'~哀k�	�S�LY�tx��l��W>�����֟�	P�)�b���dI�R�U;l�P�So_�/v�i�䁃e�L]�)O���?au�.�Ć���k@�Q���,�"@�m����Ox�D�OB���<�÷i2�Eұ��f@�qʳn]%K�>c&#��Y��*�MC�rn�>���i��H��/4����߹H�p5;���zm����n�x~�ˈ 4�����|�I�8v�z9�6,�TG�dcQG�w���<����?���?�Ȧٕ�����80��������
�%;f�R6mX�H��O���:�9O*8mz�5Zq�lq�r�дM�!bs(E˟��w�)��n"	l��<�$$K�x�ɑE�9�����<��n�"R*�� ������Ov��ɤ8ʄA�w.12
�щK����$�O����O��V��	����'b҃K�i����G��Z�,0
�*;B;�O�y�';�'��'���sRe�_�Bd�D���Jz���'n*�M�f%q`���"���?i���'h���iO4H�v���ӕ9Tx8��+_���'Xr�'������7�ɟ9g���+�C��!�ß�h�4Gi��9��?y¾i2�O�nR�3�*�{��QvR|H�$���z]����=[�4�����!���4i�!w���FtD-1Q*=ឌsC)Ԍ!Ԫ�$���'(��'�"�'��'����h�2xmB��`�I	J`����X����4O��T���?!����<9����4��:-@�J��A�K�%?�ɉ�M���i�O1�"]R�(�'.DHa �[H�K�E=�|����DD� �t��\�O�`!��5�D��Ǜp�P5�Vh��������@�	ڟ��fy��{Ӑ�P�o�O�$;`P�WhY8�D�+2l)�=O�9n`�F��	��Mˑ�i_�7��5������(���b�Byc�Hx�JvӔ�Z<�9pb���L~*�;^�pm�勊�9����'b<�`��?����?����?����OV�� �ЕW������;{��zTU���I��M[�˟�|���}��|2�V�m�B�je��0��4��#>QjO�,lZ��M#�'u����4�y2�'Ul�Ж�V���9�w)�(jvtyb5.fQ�I}��'
����<�Iϟ��	���a�K,�����>i$�5��'��Z��Q޴0�����?9���'i���C���& W.��u��/^�P�'��.��&�v�-$��S�?I���*vtȔ;�e����R�);�~�k���T��'��t-���lI��|�IB��Xa�I�!60�Xx*׆=���'���'���Q�Pcٴ)��}P O@�Dz8�t�)2΄�Ya�����̦��?�tR�, ش[|��R<�QJ`���^g.���i��7m�	
ݾ6�1?�%�-��I�����  ����8����b���Z�6O(˓�?9��?����?�����K�2�4-p�K�&�� @j2
[ <m��{�~���ß��IV��ß�����k���!s#,0��M��hC�蒧ɛV�f&d�||'��S�?����"�(lZ�<qW�	�h?" h�Q,Y��e�2jB�<��#C�&|��[�����D�OL��X�(~��#��!�0�I3 M5y��d�O8��O��gܛF(��JT����`��Π(8��V��%�wh�-8[�O���'�v6���i�O<�� �/Ld �LG%-�Z�cYl~�G��J��,b7ㇳa��O���ɲa����4|�FԢ�n�;p��<��#a��'�r�'������UA�#6�YB�DX�^r)�5�ޟ���4�����?��i-�O��đ+
�Ųa`�/X5��C>4����즭��4W̛F�S��4��D�-:8��')
�p �Z��R�K�J2w+2�p7�#�Ī<����?����?1���?���Ǎ
��eC�S��ȹV�&��¦�@0d�ty��'��O
�!$x-�V�z�u�R%�z-��x���pӮ�$�b>�RŉǞ$t�<�G��S!�E�7O�q��H��QyRM�5�-�	�'6剀{� 
�Ιe�L� G�N�-�	����Iܟ��i>=�'<T6Mޝi���3 �(��'�F3oDHiS%ۇ�����ܦ��?�PV���ڴ�F�yӎM�A�C���F��G)|y07��7�6�n�@��;.fe��O�'��D�w����XX�hq2��b�\�ڛ'��'=b�'�'�����kf��@	��9��t�bF�O,�$�ON�oZc��'HJ7�4�D�&jXs4��!�~�{ÎтK��$�|��4V	��OE攡��i���#�.�P�d���(C�/D:K����'	 �dB�I�`�Oy"�'��'B��x?`!��$��� �K���%x���'S���M�eM�<����?�)�%f��9򸲡�؛]Lڼ1土�ȭOZ���O��O�S�~��"X�6yd��u푦;�Y��᝖p��lp~�O��������R�%>V:����\ɚp��?y���?�S�'��dM�]�⇕=����Eń�B��E����c||�i��&�'3�'�
��?YDF=AK�t�@�&F�ѕ�T�?��)�j���4�y��'����� g�9O����^�-w�0�EM��]<I0O�˓�?����?����?�����tu>���Zw� pbV�ǿ�tlڠ9���Iğ��	D�s��A���K�m�3����\y�ȥሼ�?1�����|���?a
��M�'�����K�<BF���
�>�Fe��'��Q"4�l?�L>)+O��O��Al� 6���d�5	.��b��O.���O>�d�<�ֻiyfxa�'�b�'��yjV��~��X���x ��%��IZ}R�'7��|�S�p�)��FM�sQ�PXu�҉������fY��n��b>I�0�O����;���� �8\ɳ���6S����O����O:�D9�'�?!�H̞B�.P�����a����$���?v�i��,v�'��&sӐ���?6j\X�-��X����Sl�6���������	Ê�ݦ�u�i�1�ģF�#�FL[�摨�\Ł�f�C�t�$���'%��'���'t��'�]8v�ЉZ.��1f�=RKF�KU�xIٴ}Xp�B*O���"�I�O(�s����=*�B�C_?zxN� �~}R!t���oZ)��S�'g���@S��n��1)��Szi<`�wo�S�9�,O䥱���<�?)�;�D�<)�jR�@�Ze�B딌C�X$��̅�?���?����?ͧ��D�����%�B���c�C�h�v���Ï�"�������9޴���?�]�������k�4F� �a�7c|R��LD�^��HA	���Mk�O~��P���������w�z�Ëڤ=�H��u���"�����'�"�'`�'�B�'��j��R�H1,����(�X�C��O����O,n5>��џ�ش��& ����(Nɀ�R��i��غQ�x��i�� nz>(T�Tզ-�'3L �QN؎:n&`ҡ\�Q����`ZŌ��	&P�'��Iԟ��	ȟ�	7��H�b����Icg˲v������'�"6T�{x����O���|p��4��QȄ��(.a	E�v~R�>	Q�i�6Mo�):e/[�sjpء�'#��9VI˰Q�"��DV*Ĺs(O����?9��(��ЅtjdQPqIN����'��3r�!�$Yʦ� $*߳,�͹��ͦr�>(x��A�4��-�'��7 �������ڦ��-�"F&�{��3W2p��c ��M�G�i��ưik��?"�&�ct�OR2P�'
>M���Βax$��I���ࠜ'��If�����A��qz�
�JK�	��ê�M�t�K�����O��?9����S��PC~(P����!"��;w�i�O�O��3�i,��1��Q��AG8%�dM�p7zX�'�(eڠ��П����|�Q��'T:�3��F�|m��'�"�ٰ	Ó[�v슉l}�I֟t�ŌHu� c�&%\dIp��E��
�	���m��ēc��˕f�Y�k���V�f��'� x6��h�٠���Ƀҟ̠`�'@ )YN�H��P�&O��X��'H��z���2T��]���]����R�'��7-Z�I���כf�4��5p#Ȁ(j���!�Ě�g�6i��9OL���O��d�u�d6>?��J�a��'2�� �:f��2��	�CS���Y6�d�<����?y��?���?A��'QV�0� .���4�4��d]̦Y�VH�柴��럈�2�Bj�$A!�AG�x� �34�	�MsE�i&O1���7A��)���V�vر���XR�!3#�<�a�C�r�������D0AO\u)`Ƌ� �E[�Л[�$�d�O��D�OR�4��˓k��0V�R����8���D;@y���V�UGb�l� �(��Ov���O�plZl�Z�q"�Ō>f���B�Mj�qC�E�}�'|4� @d�i�K~���v|����eP���n�Hy�d��<����?���?a��?�������d��c�1�P���O�`2�'7�h�D�,�<�óiU�'��HG�CM����G�G��m�Қ|B�'L��'������i��$�OV`�n� ��ل,�V]���(JM)�	���H���O���|���?9�x�  � (�)�41C�[xG�����?�(Oz�m�
r[�1�Iş���~�DL��)��d��U7�(% M����Mn}"�'�|�O�R���-� F�e�j�"t&@�a�x񅙤K9P	��O^��I��?A�+5�$��j`��	���2�D
\����O6���O��)�<��iU�M�E�O45zT9k�фMl��!"Y��#�M;�"��>���Q�<�7�¶1,
�qQD˝h3�ph��?�f��M+�O�1��N��J?A��ĵ(��He�� ��p� a�H�'u��'4R�'"�'8� �r�v�6�,�K�N	A�����4B�ش���?�����<�S��y��S?X�\;��Ǫ}vЫ�J��JN��'ɧ�O����p�i��䎭�v�!���T�a�A��4�$�:�r]`�C֒Ox��|z��"� Ppu�Ԫw@*��Eȉ0��?a���?)(Ov�l#�@��I����I2iX4��O�%�"����hd�?a3R���	��<a�
�-`�i�� ۩>�@TR�.?�taK�r���)�J�@�'{���� �?YPaTq�D�n7h�I0�H��?��?����?Q��	�O�q�Vkޔ~~�4���߿�h��qN�Ov�m+E��'��7�7�i�i�F+� W�%��,!.��1kz��I���4f���[ݴ���(����O$ha��
�`����axӖ|�V����韼��ɟ���ȟt�$b��k�8M�VD� D �3`Yy��|��`0��O��d�O�����č�O*�\JV\P���|�D4�' ��'�ɧ���'�2��<���P*4<H!������E'�@�	#RRlܢ��'by%�Ԗ'Gd�`�C $�a�6m��4v�'�B�'�B���DZ�8+�4:L�v�n!����fIH]�SB �gv�r��
��$@}��'�w�~<
2�9fU*�
��0G,��kR�X0�M��'�x@���Ss���?Y�]�Q5:m�s�YI�Z�R3��x���Ɵ�����l��,��D�'m��<2���{��3�h6~F����?��5��ƭʉ��$�'� 7m-�$Ϭ����	�w�T)�b��`���O��D�Ot�䖨=�H6-y�t��1��H3d̺O�������k�F�[�
��?���2�$�<����?!��?�:Q� ��U� .E�Hh��
�����OJʓ6�& ^�v��'(R>�:&D3��sF�6T�r=a�k/?a�]��p�4mś��,�4�����9�"0rׅS�H�����lb�C�n� V��D)�<��'iJ�$%��Gb��;@Fٺ/(���Ћ��Ԣ��?q��?��Ş��Dצ�%�U8	d-I��kz�Yg��D6X��'w�7(����D�O��k��ߎ)��pY���;uإ�g��O���?&�&6� ?����xa��>uH��6}�-Rs}�����A1��$Γ���Oh���O����OT�D�|��I�?y۰9�"֭�2��IЖ����۠�"�'P���'7=�D��Sa�� 8�(Ӄ�:�hI�D�O��3��_3D)h6�g�\� �N#���Wg��D}��(�Ni�<R���~pr�I��_y�O�BN�<g�qH�'�-�q	F`��2��'Q2�'/�	��M�쒖�?i���?IS���#mT�b��,+���Z�H@!��'�:��?����=�T��ƤS�c,��I�iT�q�';���Q�O��ps����ƟXs��'��i�5�հX���������\$�r�'���'���'��>�I�1�L�'iH�%t�C�ń6$����	��MK����ݦ9�?�;���X5 Ry3d��-���̓�?����?Y����M�O����� ��'�M�m�<܊�\�g�$����':-ܒO.��|"���?i��?���{�LX���=P`Zc�CD��.O��lڤAF�������I@�s��UmP��U┿�p���Պ���O|�d'���Ů�8��	�dV����d 8HB���#��	5�@4���'2�&� �'�¼!�(�5vf�T��'�z�xz�'���'%"���D]����4UA��K�z���@"�߳4���S%�i�r��՛����p}R�'R�'�8m�e�.z8A`gӰ'�v=��N�x �撟���M��N����I��ؐH׮	�lXp!�.��0�`>O��$�Ob���OH�$�O��?E���P�Xi�hG��9�r�`�i�ty��'r�6mA�h���M�K>�DMB�N#�`��h�DZ��L�NՉ'P:7m�Φ�S�y7��lC~҉��� �@�HM%fbB�h��2t�D-b���?�&$��<ͧ�?Q��?�c˸V�txt���:h"4��?�����$Yߦ�FA\Wyr�'���*naz�Ye %)�
���n��h�	ܟ�*�OLAoڊ�M���xʟ���D;b�40��C�Q��+�L�O��1�!S�D���|�S��O!�H>��4Rr˅D�=4����fÁ�?�Ʀ��	Ɵ\�)�SNy�`�RPX��ǚf�8��`�S}����.�+���M�"b�>���$�.�8d*�>b�����48�	J��?Y�K���Mk�O�:B���O~������$�4X�����K�'�����8��̟��I���O���G�,p(�өF�>B�=�0��(,�6�)Kz��O���7�9O^mnz�mf*�
l���"��lT�q A*�����I\�)�S3'}t�m��<1�Ɍ�
Z���`�ͤ_M 	���<���
���Ip�	My�O�rc6Vފ �2�����J�r�'��'��im9�4�?��B��KE�T0��B,H�nd�mʉ��'����?1����D bx��OQ�U��77Z� �'�����^�&�酳�~��'F`#֪9���xU%ܧW�4+��'���'s�'!�>�	�v�N0���.��|`3��.K�X��	�M��\~�Nӂ�杕'F��dS0/H�h��g�L�*�	˟�I䟌�R����E�'��a�s
�z�� .^� L��iY+v�@ի3�D�����4�����Oj�D�O����5Nn2e3F�Id�L�5.�$W�� O�櫗>q��I�$%?M��5��t"�F�Hd5�(�,e��{�O>EnZ��M���x���Ұ@- (B$-��\�ש�pK�)	��!5��ɦr�7c�O�YL>A+O�8��#;x"��5�ۛC�(` �'��6-N����<8q޽��a�fzMq�f�;-�������?�^�t��ԟ�I*S8B��$�Y'-	�x���
 @��Ȇ�Mۦ��'(�h(׋��?�pV����w��!��DN@$�B��AN�
�'�r�'r�')��'c�0�{w�T�;`x2�˃J����OL���O*�l�C�@a�'|7M"�D	�R���r�	+�B)�uOW�p��4&����ޟ�ӭ)
 �o�x~��Q�L�,C$ß�����"�3u��4��s?�M>�*Ob�d�O���O��쏙c"%�$�@
b�� ��O\���<aB�i ��a�'���'	��:D��:�'ٿ;�8=�4&�g��Y`�	�,��j�)��@)&���3��8'�Tت��Z�o8���'�<�M��O�)ӟ�~�|2@t2�Q⥖'>��0���Q�j;R�'f��''��$\�8!ߴS����GE��h$ !��CA�-���zu�O.��d�ʦ}�?��S��1ڴP��y�e*Ƞ=;���-�	�9	S�i�N7mF1Tq06�*?�u*Ѡ28����	��Č7
���!Y�<���� `���BƝ�k�fmr�IFP0aǯ�7P��[7��+M�L@5�|�B`���2Kè�$��c܌�t �/�!��)���1׬�%G��I���7�
Ԛ�	y�B)��-��c|��)F���pqV��/S�Z���+�Zt�0��4���y�b�6(���i n�.Gn�(p��1�c�oN�̞X�����9Q`�<<վ4��m� [FDQh�˙�p���AO�;�F�B3��*&f!�F�׽`��f�'lB�'�����>I+O��V&C��LZ���$,/�M�ԯ�����c�Z���O]�%��%~^�
���n�x��W�Gg�7��O����O�m���U}}�^���	c?qA�X-"������0�(����y�J�!�H>9���?��b� �Wf�Z�����ڤ ;ά꥽i�Rn�	B�����O�OklȆ$��%�4Ӿι�E�Z�E��	�O7��$���	����ny��H�l��Z�I�@�I#7�� %����>�/OH�d#�D�OJ���g�,X;a��}h}����WO� T��O����O�˓V��9��<��Q�G"6�q��R)9�*��6�i���ӟD%����ӟ�٣nv?9R(�,g.n�rR�"FPpZ���j}r�'���'���L��1�����,4��T�����*�DK��%m��n��ؖ'���'�Y�C*�>��'��Ah����J#_��]ۀG����Iڟ̖'B�$�*�~����?���4�����K2����E�R�V�"�x"�'�b
*'�r�|rП�aʚ�^Z�<�pe�WH�8ⴿi0�I�Y RTXڴ�?���?I��nH�i�2 �Thm�4�:�0;�l~�f�$�O��!���O��O��>y9 i� 3lX����P)����h��|�r�릉�I˟��	�?A`�OPʓP;�x���!s����U*VX�u�A�i�9��'5�'a��$K'rJ8&�:EC��*) B�n���������r� D:��ļ<1��~ҁ�n�f��!M`��@����'��4��|R�'���'�����F�oA&j2�'|�~�p��l���$�nL���'��	䟠%��؋7.aB6/ˉttų�b��~��	'(����Iiyr�'���'��ɹ9���qrg�rVD�̅�,<:�P�/N���$�<�����?��鶴��DR�v��K�AuK~�;U@����?Y���?a/O��hT��|ʢ!+"��<*�.�l��!�3��d}r�'�2^� �O��ʟ�`�Ɛ.��+1��5҄u�v�ș���O(���O�ʓ4_�����B&[�0)Ǎ�G� ,��fZ�`�*6M�O��O|��|����3� ���E��~%��"���d�"���i��\� ���Z�O>2�'��\c���3� �8F����G"bB��&���	by� S��O��K�H;F���ӀO��FM	#p8������A��@�������?]��ulV�D>�9�&��;��Q����M#����dc��P�B��q=�i�� ̇*Ɍi+��ix2�I��'&��'`��O��)J�&DO�9��bչ`� 4�c&��փH(�Q��y��I�FRPAQgGR�VP&	���l�䟄�'蠤1�^����	Ib��s���(A�����R4�|k�y�BƓ":�c?a��_?�VX=�)T��"��̸����I��x�'n��'��'���X�oM��)����$Cz���>��
�����'�B�'I"T�\�\S�;rmކm4��ӖB+n�4��.��O����O���?��eM��G�%\;�pBb�:�F%��"	�?�L>���?�,O2����|��aS��V���,��"E:1��j�A}��'�|�Z� ����ɟ�j���M�cD�' +j��`*�2����O���O��'�L��3��TaS��1���=dv�a�3��W�7m�O~�O�˓Ƕ�����S,\a����W�j��uI �2Sw7��O��$�<�oP�D��O!b��5��z�"$
ԭɂ+�4$`"�P��M�(O��OL��F�OD������ ,�T׿<F� 2D_�h�l=�&�i��I�l�����4�?���?��'j��i�	 �,�� NR@HtkZ3!y<�1�	gӜ���O�5�#0O,��O�B���v�VHBL�U�P@�W��V'�V��Iu�7m�O����Oj��p}�_�Pk��/V�±1�F?p���	X��MKG���<�����7�៨b�g����{Q��Z� 2&�Ѳ�M;���?�� \�0��Q��'!�O]:uO�0V��oS�/@ q�i��Z����m���?!��?1uς?j����Ň-|�T��t,���'3(��0j�>/O���<	��S�h}��Ż��O�I8����K}"����y��'r"�'���'���]h\�����D; ߞ1�� �p����$�<	�����O���O�;7�ʳtG���nA�&�֭�A��?f	���O�$�O��D�O�ʓ����?��8P�F��H�f�;���H�d� ��i��ٟ�'��'gR���yB�d^r��po\`J l� ����?���?q-O�(Y�PK�d�'_r�j��V=�6��� �3L�j%�~��D�<i���?Y��y�����i�B���^�O��i"E+�xa�pB޴�?)���򤀔L 0��O�"�'��fT+�n�k�bN(l���j�i�y��?����?�G�T��<��O��y;	�	�^4���\�,��I[ٴ�� �rhmZ�\��ɟP�S�����VA��Գ
|�je�΍ LXP�i��'ײ���?���?q����&XL�T�_H��z@�	�M�JJW����'��'��dE�>�-OF� A�8i�Ω�C�M� �;jǦ=* {���I���I\�'�?93�-j�@���H%]�{EgA41.��'�2�'o�����>�,O�$��(��1q*���/I�˦}��bӸ�O0)��;O���8�	d+�¥2� +��R�i ���M�����uZ��'i�Z���i�m��ڑ1��6`�y*f5����>�5H��<q���?I��?!����N�n`�অ�L(*�q�"
�n����V}�Y���	wy��'Pb�'Р P磅]�BEB�,0nQ�t��yr�'���'���'��I�JM>=1�O]��Kڜ�$����D��X8 ۴����O��?����?�'�[�<�&�L V{B}pSd��U�+�mY&H��ڟ`��֟̔'t��5d!��Oۖ��C�]	`�:�S ˝"'�m���'������3�ǟ��OxIK���e����.K.�9��i_2�'��	0֦��O|���ʀ���cBB��͍_غM��Li�'��'6:칛'��'���U3���/NS6�q[�dF�U�vV�LK��[��MPU?]���?�`�O>q��hF�( ��3π�`�i6���ud(��OU� `��`��r�%��^>b\ܴ8{ؘ+%�i�2�'S�O]bO�� /xyZg�ҘY�R�r�E*l>@(m�T��IK�Io���?���ոp��,9ql��B�T阵�6)B���'&�'�(=ʦ*(��O��d������הW턹��M���(��e&���7�:p%���Iޟ$��*_<|��ُD3l�@�>m��۴�?9FGʭ=c�OL�D�<1��+ KM�^�[��W�i��U�^}�B��~��V�x�	ǟ$��[y�=TGzA s�Y�
�^Y�5j��qJ&XJ��7��ʟ�&����ʟ��f��MS��U�F)R����C(7lD$���������Lyr��H擝Mˌ�i��R?���C ��(7�O��$"��O����Aj�$��.B@LR�)�2xU Zf _yy:��'���'��Y��q�ʸ�ħ��x��"I67�i�폶fv��ɷ�iv�|��'w�N�6>�>qA�ՠ 4�h��Z=
�$�RF�˦!��ߟ\�'�@#e0�i�O^�������K�]2�gJ6qx���d�Ox����O|��<�O��Ѣvn_+���P6��{���iٴ��$W�V���o������O����}~�Y��~� �ʂ
V6�Z�Nߡ����O^x�G!�O`�O��� $�a�!?m}��pI���j���iv����oӮ�D�O��$����%��.��Q���,"^���F�ox���42�P�!���S�O��o���a#�TZ��yVn	�C��7��O��OZ+s(�<q(���$��t{��F�\����6L2`�"Y@G����'�j!�H9��O���O2�p&DC=4�*�)��O1�@Z3���y�I?��2N<ͧ�?�����I#?�t�1៿7`��)�T+r�O�BD�<	��?���?Q�4�
��"�=P�-�E!s�2�+T�_<����O����O �O����O��"4�ǄI�|T
� 
�t=s�§��cӒ���	Ο���Oy���l�8�'~`�	�M�2�!��>NQ4��?-�M�J>���?���Co}f�%Wεa6�S�/z1���!����O�$�O˓n�"tj��d�@� �r7��3(=X1�Rd	"V�6�O��O��$�O�Y`���T��)*�l�t�a�&��(R���'B�Iß(i���A���'"�O�wD_%d �U� /�R̪��Qk+�$�O����o�pPs�T?5� )�i�H93t&C#q�Д-bL�Y���n\��M�T?y���?�B�O(�Y��<��e�2�V
U^�(���ij��'����d*��?���5�;<�y�*	8\6M7K��mZ֟��I���"���?`�R�y���s2�@�pR|C�B̭I�����O��?i���X)�yx%���
����@%\�`ߴ�?���?a���+���|j��~��0�r̓B@I�+֝�g�Ă>?tb���� =�ħ�?����?9&;Ue|dAU"U):Q�ᄆf���'ZtC$F�>9�W>�$�O~�'�>��6�F�Hb�۠	�?$n�@�O�Tآ��O���O��$�O
Xٰ#Z9,0H�6a��A5��X���(q;�˓����O��O����OܬYclRg$���
�8U�	Kc��$V���q�>�E�ʧtՠm ��JC`c?y�B��&{F9��@�!�,Պ/D�Pt�-_�dx��䓕I!�|A�A)�I9����Ā ~�b�#�-����	,P4XҀ��x�n5���:N��0�c#
�!�D�)'nT�?&��C$��Zzи��
�L���Z ��$r���$���Ph�H[y6ڽp�H�i��a��Y0B��H7"�8���1�O�F�x���P�ITX-Y�N܅]��rc��*�$K�k���CO�}��� �U6w�����O�a� :`��rf��*�}��|z-���`p"�;z|H�K��ޫR.�3�>Ae&�'`��e.�(`��H��[���DğTe6��b�pp�<����I䟸G���'���
 aD�3�nI� lIHr�M�<9��\D�QZ�o�YELe���H�ٍ��#c �(s�@�V�� � d�9l�ڟ8�	�,����	; ��Iß�����] I�>���"��h#q��<,Ƚ��L
	��	,4݀C �3�䍉1MX�$���G�L�  Z�pM�'T�,���m�g�!M9�9�/���ɪĩ�d�&��	o~"�S;�?�'�hO�!hӈB:ge64��F�$��Y�"O^�����|�.$H�+ˉY��E������4���d�<���oI��^,��.ëK�,0�ဏ�?Y���?9��n��.�O���y>qʃCH}/8��&Ӭ.�d�+b�Q�/�V����
;$�u�a��`x��ط'ߤs(R�@%�	��xKqN�+��%B��D|����B�����DQ��S���&%��T�� 5C�p(1@׮MǴ���Oh�=��b��2#N�p�. 1�T�GG ��0>�H>9r��.��衡^�dʠL
0@Rc�5��'^剱`!~ȫ������7h���k�Fl�������0�����Oi	a �Op��w>� �'`��e!��䢭n��A�(�������%�T����d�31}vlC�N���*i'�~��]��N���&
���+^��r�'�@*��;l���>qB�5���U�;�D��� x��?1ϓ_��â���d���R2"|�� 蛶
���ց9�-�*N)�Q�n���y�\�h���_��MS���?!/�⸙V��O$L�$j�.R��
���F�R���O���_<"u��L!��|�'��-yT���VM@���+�![d�QI��9a�z��Pӂ�,�=���i?_*�-�S�=ZTX%�b��2{�d�	���4�?I���NH+B
�x�"�-v�)2�AӘ'~2�'K�hP��G	p80��Q-V ���y��|RcӴel�v�I<,�� �,��:��C��qN��[�4�?����?	w�`بU���?����?ͻ?�L���A8as�X+W(ϰN�����H��?H�	5��i���/�3��G+Z����ܔ{��/8Q�<�cSF�Ty�O�Z��	�}&��DH)*� �R.I�;�(�QLI̟��'t�Q��S�������h��,�/y@�G��g���çQh<A�N_�}�)x��
4�2��!�@~�"��|J���Ć�Pe>ѳg�]94��4. 1k��W� V��d�O:�$�O:կ;�?	�����H�	'��I�Cbґ_�dD�Q*%��S�K[� K�N���0=�W�ͲsS��#�Y���j�({� p;'aL#�Zq����0/��,��iΫss"�<w'"� �1I���0C�(�$�6W9n�aF�O���$�!N4�An��\�`����ĽOSa|�|��M u���袌�'@��hZԧ��Ϙ'T7�/�D��=��n�ޟ��	�VY^aX�"]�u4q�W�O�E>Q�	D�!Lԟ@�	�|B�$s�D%���Tqr.�0$�� ����j$OBM8ߴVpv�Q� ��gW��Rl�b�d�P�~�@�� <��x�Ò-�?�����D��#|�8;�k�F�,��Q �{	��O��$3�)§l��se�N �耪�`G�R^4���~�����V�ڥ�s�xgI9�yB�)�UU�P�Q�Ժ�F]�3�P6Ypl�ȓ;,>�pK�o��2�(�*�楅ȓ4������~���&�_.	|9��z{$1�G�Tu:Yb��:t�^����V�.���a�%�o��ʠ"O2M�ա�w�"��G�dN9�5"O�l����<B$t�[��4\�4
p"O*�3��	e1���' �oT��*�"O�1��+ɣY8������	J��H"O�y��h��LCIM�xz4�R�<q�*5�[�-Q�`sf�ق�M�<��<ћjP'	!\ 	E�OL�<9�垬/~�<sAk�"3���`�EH�<Vҟ0e�-���B�}���U��B�<�1D�3(��a#�p��Pq�t�<y��X 9�m��ōe#��[E�m�<��O
��"T��a�H�@�<q�W0J���Ë-qj	�*�|�<aBM������	m�����t�<�����bf
M)dFAW2M���p�<�R-�.Œd���V41��l�dBX�<)�{���F��0�@Ws�C䉓c|h��HO�1?�\+Bd�vC�	��LВܥ}4��p�g	'��B䉺$-L4s��[�A��X;b.�9UlB䉤�2L�qc��t�p���n�|�@B�	(��t��_�P_b=���;E��B�ɿ;�v�J��
4��W�C*t���L�O)�\����&X5.�>%��=r1��:$$�aJ0$��k�.(j���32�Juf )����M\��I��3�|lA��mpȣD���9;�B�	%f���#
�+��R�.��bP`�I�|�ѻ��Ek��s�4ӗ��+H�W�ޙ{� ѓ�	"D��1CR"Y�f�t6����0�a�$�!f֯ 7�cW�[:L��x"�«+�]�� _8ȢX�R�p=��
�h�y�����K/>��uH�`�S���h�j�'�����/^�3�O0d1,-f˓�m�1O,,bÃ�-v�����E�qs�A��dD�3x�J2��(oB��T�R+�yB�Q+s�@�zG��u�l�:c	G6n�0SĉW���Y��v�,����3?���$?����V���&�T���e�L�<Y�E�Z����&�!��[�˒�e��8��@�;)�P�u�;\OЉ�#ʇ�9z����N�|�vUy��'���i#��&;��ۄF�?QZ I'�#(6��3dW�v=���'�
���o�'dn��Gϣ?�Ь�y�O߃ЭS���=}xD�Dn�1S�ؚÆߟ�|��L��yRO�,�"���9}9P�Ѓ�I���0� Bؙ�\�ʼF��O�p�-�Q�Ҍ����O\�e	�"O,��!=O���˖(R�A�H��f	Ѳ���񐥏�,	"�ד0���#kH�S+`���E�(�1��ɉU��H�&�O�Oq�3�H�
fN=��NV�H`�݀P�>R�C�IX�n��HM�0�nL3p(�� a|c�L1t Ц`�|����F� Q>�B���/Ȉ�� G!zɂ!���3D�(㵠�Kw����,�1*��ɸ/��
�p/Ȝ��D֕8�>�'�Eh�,Ϯ+�\����#dt<��8R��$�]���y"��&ܾ!+������ ��!�*K*gr@�F՝;In��2�'��y��޽d�F�1о(�Rg�$%:4)yw�[�k����ȓ)��H�B�[^��gf=��u�<cn2}@�t�v�.�b�U�p\���QH�+�6`�ȓ~�e�2L��|��=g+؊(�A��H6lC��'�64���,B�'�0�h5q 5s*h�a� D���p��+`ЀKga�`��L���]*K7�����4�1O�иX��' ��p���%�ӫ�7m����)7��Qe��v����4�>q{V�=�¡Kğ�\��I�3d�J�&�d�b��#K��
"e���<�<	&m	�P;�=c��=����!��f��l֨�9�>8�CKð(m���?7�I# �]�G<A��Q4��wK�B��f��XSf�2���x�;]'Hi���aX���⬒�`�]�ȓH^�X�`�K��xxC'����P�Ů������>�ɬ��л��g������ț$
���[�0=	C��R��e�ե�|;�FHZ$D��9ض�J%2�L#���'��d�.�,��	�;���v(_6sAȼ� �D��b����-l�ѹW���-��ȍ����:q�2�G=)�� B���D�PB"O��h׊ԕ��X�P�L�PdR���6-H\���$�*�(�� �ay�c��o�@	2��e� C�	�O�aB$�'E�ѲO2l'���:f�2|P �Kq�z��$�L=:�i�6�xu��9�Ms˓aZA�uhĥCg��;������4��(p�D��<︱�E�
�����4��0;b>-j5B	�h#J�	w�M9g�i��4�IT�h� �Ă��Q�2���0����~���Y�6�H�i���>n�
!�N�<i��ľV���n^�����*�5(DÝ�s$x�G�<.gn����H���x8C�ǐ>�N��6�'8���	2W�t��B�0S��� ED�q�D q�O���C��h���a"�?#<��I><�>����&|*}�	�ʟ��僿��i�į§/@���A6�|� �$J�U�V�\�r ��$OQ�8�H��Ju�'��+�ݐr��w�p�1uo �:�l0ZU�Z<+�N�0�kFN�2�8i�	��i�pwh��P��\GF�;�yR� ��F�9����� s��;Ϙ'�l�JG
P�	°��̕%b]
݂��D��iH 4�R8����@�[�0�J�n�4��� U���Պb�!8�u�B��P(EM�hVaz2ɴ�b���@7��C$_��yb FY�z}p+�d��+2ٔֈO��3�۾0����sfH;S<��kG"O���V/¶�`NS����J��J)/u"mEi!ړE<��P!14��̻d�:�I��V�]��.����Db"��{��	Ij%!��\�&Bx��T#�;?�:���J��U7*b����B���KK3a<Fy��Í�1OEIE*�9m���"� ٓ$N�����OLijdJ�&�ʓh)HD0����%y���V�ɑ~�������o����C ?~�냧��|����n�)����䔂6�p K'�f,z��2S��#9�h9�1oɓ^����tBQ$K�ў��!���I��Lc�����BҦ"�O,�CТ��?�i���2Z�L�p�gW�^@�Mk�DQ�V�()�Ŕn�':�����!S�0SP�
� I9��A�f���Q@�1L�9ӎ�Ĕ#M��I8��I�F�J�PD�O�8Ѣ��S���R��уŴm�t�����yr��5D����BOE�<�TD�6��'�P�F�x��}J�ǔ%�4��� u)��e�Է$��LX�M�O�R�N�/8V�|H�״e4���aӪ�:�ӒQ�ڍxi��<�ܥ� �Z�#!>,��ͨvy���'��B)���Ƶ���O0-H�`Q�=!Բ�7cD+)�|Єh>v���F%+ғ?|	�Y�X01�dW�>"d<�q�+�Oj�#癞���'(?�B�����0(@,�[�I��2��$�hMEzZwЀY���Y�>d�%�Y�������L�.8���B�4=��PI��O�>a�=c�;S�p]q��պ��W��J�%�l�Th�<i�T�ʐ�d�)jT�Ȕ�@�T�� �(ؖ1O��:GMƱ(hui��Vp��0F�S�����r�v��b.c��YG2�D�Ņ}�2Y�A��(}0�6!>�.4�� ���O9�(��,.�aY�k��ׯ,LO�I�"e��M�����B�P�$AѰ����!�X�0tˑ��H�ִ��M��HO��""l�;$�ܤ������( i@�'Bf�A��]*+�ɧ��'L�ܪC@V��1PT�!v�f��V��r�N��#��=Z%aab����#=�;�k 2�иC��#c�x�AqL�
r~V�9�B�*a�D$��R���>��O4��aak�clt��;Ox�Cu��X?��8�H�%x���憌+U�1O��⎜z񫌮C
�X�C�'n��,P����ͨEcr:W۫$κ���+?�Z�[6"߱S%0�K��'$���݈�r8SˋdN�� ٴz0���ɞd׀�C�F�*����	����Kr�!}l5��b�q����<|<��7B�#T�D�I�HQ�:z��ٴz��Mq�!Q��ְ>������64X����}��� )rH~h�#y(�'$� ���t�ɧ��{Q�����U�R[��S=L�xQ2B�N$R��1��	�=<(#v/I�? N����E(��p�N�4s�XZ�;O\eℚ|�ㄺ_��)G��H2�i���~r%I�|;4��7���[��HO
t���[�]ZH�����?��U��c ��2⤈$"@q���O��"G)^�x�� @� �O��!���,v��	#\��@v���jjb-���̦�x���P&ȝ�ڴ%7��Ћ�S��������?!s����nP+��IO����aAY�]IP�}�t�d�W��*�'E�P)��Y&����d�10�e1�#�1b^�=�g�֜u.����^���N��FK6�~���5�q�w�� !����[�t�V��l՜�@�Rh��wX�Hk��	t�'ΠTq�
��v�HD�!(��D�@ѵ�X�6�X%�p��>)����ʕ�F*Ȧ="��KKB��i�^��DKA,�@�����7 ���j�Ɂ�#�Dz��� �ls���$�`����~:�+��'��xr҄�S%���B	�:�zƦ�g��(3Q��<U#�7MF W�Ȕ�H>�q�O�T�D�H� .�آ��1r$�\��4����¬mz�!C*�(CTG}�fR�&��Ezk��hf/�+bpJ����	'�`��".���#��?��D�9ph��"
K�6n,��S�֬O��ۇ��<��{2E�ve󩒍�b��[�j&���-�TA�4$ ��DF'R���T?a*]_�T9����G�XйT*�pc(���	e̓tk8�A��a�����+zJdCf%v �<�p�'5
�Y���*�1B�^,l.��{�/4E�U@ݚX5n�bQa�1Jvb`�t���[���A���9�I�-�����r� 7m �e��p�dۈd�h0�0d	 VNў�XAƜ�7-�Y�ec�V���3f@�l�x�*���vPi�K'��ZE^���=��_��5�v�J��k��_J�-���M���>)���/X5� G�-~�FXd�F�B���i؞���@�W,0aAG� a)����~`����'7,�����>:n|hČ=iJ��U��'�|��j��<�XD}��T��LrF�Їk)��ׅ�!�?a�W�i#�4���D�N�9�i�^�W`^T�#7O��
� ޯ&�(8I?�Sb��>zN黐�w���ڴ&����wBϥl��Aeǆua�+��8�}/�tڶCG#_��3TGǈ[L��O�![c���Q7�	���[v�j@���Cup�A����^�\����8&Z@:P>4(m����p!B��`Λ>xۖ�+�)^�E.�*��Of�聳e	�b�:T�2ړ�y�$Յ&���xE'��Q�bw���Px��R�>�8U�6�\+op̸���
�C���ER�ˬ3-��3��Rk��p������pJX�9�jq�ƫ�U��@H��'B���P�]4�ȱR:7K^i:q N:8��S�Dϗ���!�ݕ��D3}��HG ��6����F�:qQ�`(�E]��^�ar,O�#�R� Ł??A��H�,�4��E�Le��)���k�'L�P�@E�J�����$HCV-*�Q�T5����j8�H�/X�+�0ڰƃL?�� '+��z�Ժ��M�`��$~��G���a��D�@=D �Ŭ;��׷\�T\
"G�>��U �χ��D�?Qu!�<]��iS	�_>j9�%Օ@�~��� c�q�I���%O^�IPE1X�����D�,E��-�.�?	5���n�4	6��CS��剚q(�%�p�,����GR�9���<w� 2TX���]V���P�a�I��U�z,2H㥊ӊS`nB�B+R�OtAQ�m�/a=��4�F|!PfA4]���+	��p>��ק#�{���PVl!,�`�z|�5
ϛG��y�h�&QBB�FzZ�yg��th)3�DיQ+2諀-ֹ�y�ΤL�j���Cԡ}�5!�W��M����j���Kā=i�4)�"�yg�A�'�8�eL��F����&	\)�y��R�u�ճ6R/(!|�N���y�ǝ�p��pQ��'ְ�e���y�n7;�-���6Sq��و�y2E_=����C�9� �J5Ξ8�yb�X!^(��#�ۏD�zQ��b���yR%A.e
�zV�M��d��L��yb��..�f��
��t�����y"���g��!O�5>ݘ�`���y�O���v�T.,.D���i��y��W�4d.0�mS�,�dPW��y�t�BqB�'ءmH�`��î�y"�H
IR�"M۳tK&)��y2���2E��]�l�$�i���=�yR�ޓxEi2a�Tar��A��y�^5�0A���� ��T�T��y��1xz��]�t|B�z�U9�y���,�>͋��l6�4	��3�y�픮aϠP�̪H��p�L!�y�.'t
�1y�l��9�ҝi�c���y¡}"�m�*�2�6Y�c�F��y
� 
	ĀB�`A�M���#^4�c3"O���0��k)�XV��'����Q"O4h�&P�XI �PC�-�p��T"O�� �Y�0m �b�vdi�"O�\��d��$x�(��
��qj��S"O�Dk4B�
 �M���V�pc�"O��; ��p
�(���|V\E�"O��qgm�: ���@�ZIH�aG"O�m�B�۳|�����Q��"O2����v4.���]�O<p,��"O�����j�čB�F�fC�Z�"O��.\�h%�F�8�l8`"OI{���%0���:��ڟ>�h�i�"O�qqPa��jb�9�䞰&�r!s�"OXuAa�ѴY�`�&ɠ��8�s"O��(a�"q��5�4��;b�~��v"O�jc#\�y�X�ŮP��"O*4���ەETL�	$�4h��{6"O(1Y7��z�V�2�]�M�Ī�"O����e]�V��i�[�JF�UZ�"O:�rS'��;渄)"I�m�>,00"O8t����p����`�|z�eD"Ol�
P��
�����m�>��3"O�
�,���{f�L9(�P#!"OtM�ԢY-Tx=)F R�)P�"O����P�n�&��,�٪ "O��������[�/\		eN ��"O�jB�ҷ'�-[��9eZ�dX"O��04��.�����';F>$u`"O*SE�(S���Q�"+3J��E"Ox,1���F�bLs�!��c"ORE�S X2s���'!�,fF��D"OL�(��g��xBPn��3e`1�#"O��ע��W`:�N�$qq-c "O�}k񈊻R��1�&M�$s��[�"O� y Cg�kVe�A_�&"O�d�f�%krD�a�
�S!j0��"O����!8z����Qju�"O��c#�DNN�P�R(ti�d�"O��#K��N|����sd:���"O4|9�bG	�D�A�0_AB�"O\y���K�dh�[�JJ#i����"O�}�����iC�}���[	��}�"O�ᐤF�J�ڌ��GC�m�0p�"O�pkڝa���ڃI�Uj8K&"O P�EC1��	d�FeB�!A�"O&��kA X�L�e��v-�=�"O�1���pL���D jKҹ�"O�+^1)/¨3B�X"q/~u��"O6�:䄈�(�rՋv�ʨ(�Qkv"Od@P�E�o��pc ��%o"�)��"OL$9V�_=@��P� !��=x "O��	��U+[��( ֦\�����"O"T���K�05p�A��!p��R"O��(P-I��`Q ��+HH�9�"O�4�0�U ����6`�g:�9t"O8�rGdʮ\VrK�푈#����"O�� �n�/A猜{�m̄{����'x�z���C`T��R����H�'u~:K�!��D�6qQ��# ��yB�S�U�6�P���EpI�����yrK��B(@G�ٝK^u��ć��y�&�^[������!=".��6� ��y
X�Icƅ�F��=68�!!���$�y
� DZ�d��0�~�QY�e`e3"O���O��R~ m��'�O;Je�#"O>��7ńG�0�b�D~)�y+�"O���2ˊA��M��j�2��"O�E#aHQ;w<q
��m��4i�"O	I�e�9��Q�a*�<��q��"O��B�6k'��xWI���t�""O�h�EM�8WkR�)&�܆��c"O�1	��Ǐ|p$�$��/e*D"O�;��M��4�8R��I�"OjX���	%�<h�bpEd��"O�%P�h؋Y���Q%!L7/��'�'�:� �`�4��o\6E8��'�ք��bHr�0�zteZ-x{@ �	�'�P��r�1_j�2���%�݃�'&έ:� (}4�"t��	���
�'?H3c�B�I"����*FI����'��Ј��J6�����"v`���'<�h���;k�9 R�r�x�
�'m$P������V�)Q�-s��E]�<Q��I�S���0��I�=P��Xtk�\�<a��ynxl�'z}�c��m�<� P+'.�[0AK?\�b�r���t�<QC�Ƴb�P���M8!-��CCEK�<��l�/_F�$���&X�5���W{�<9�剗��J�ʘ�_��5��t�<���6����>>�|("�s�<�g�$�~(�A��?Z�zPOF�<�2�ݒ]8!j5�C:����TE�<����3�"�i׍@'Ad�1���U�<�U�! 6��`��`� a�XY�<�@��S�R�+��Ĺ%�����i�<�rG����A���=_�$�
�<Q��� �na�ъ���ȳ�s�<y�R<� �c$_�2pA�_f�<���//�5�sFP�)䘜# KPG�<�RP���E�&B/.��=�&�j�<�4�V�v���#@�D.	�z�"2�i�<��ʂ7M
$�d�n �m
Θp�<���^� �ڭ�c*t� R��B�<i �A�p�`�S�),q�(�@�<1�$�0��(Z������!F�S}�<�%�ʝ	 >hb�ƍ
l!��z֢�w�<�E�#E����.C=��dRE�Ji�<Q%��:8s ��Q�75m<t�oe�<Q�m�/8	�<�Ѵ=��L���g�<ђ ч$��� ��LD���k�<��@�7�>�h�G��3S�`�g��O�<��NNIl���ہs��h�ʂI�<Q�Q�K������>���#��E�<�emX�nX��t�;	Tܙq���<���{*�<�Ў]�YZ4�PE�P�<� @�rCfQ����Llj�zbFAO�<a�/��j�k�2=�j0◇�f�<YĦT)2T�z P!G�|*���}�<�d#
!>0x�͊+���	7�C|�'R?m����7��[�n��}{jd��M;D�(�Gҏ lI�MLU|J�Ю9?y���+
2t��q�J\��0Fߋx֢=�ÓB&�l��j��o�t��ċ�अ�c�UBw���x�(gJ'm5����IR}�'&rvv�kT�I�a��AC%e��y�O����\�D'U�x$j�m
�y��T�'���+re��N��s"F��y
� 8t�q�7+�B4��SY�Y�&"O�l��#ָ}�d�Rq��uVv�X�"O|Y"G��g�0u�f�ǩ>�x�w"OJp�cҠf�]`bפg V��f"ORt@ƌ׺mI�������/�����"Ol=u��.�l���R7	���"O��@tA�bW��#�h��~<�a:�"O��KabD���D#��2'�4� "O �C!�,69�x1�I�5�8�5"O�x�/���N+����)�"O<�AQ-Y�Yh�դ0.�X�)&
O&6mQ�E[��"� T�.6L�f�ʄN�!��/�L<�f�&$IP�ȓFV%�!�đ=Wi����8D�l�$FM�A�!�d���P��7��C+��kTE�<|!��խ�༠`�$)��x��#��|!�DЋy�0c�`Q">|��"W&c!�dZ�D�J,��C	3
@�ԋ�
t9!�&;hH8���C?$#�m��JG<,�!�D��*�5-��knГ��&�!�$H!A�ddS�H˂"W�Ł6�V4%�!��Z{�p 8�Eô08��P�Fאd!�ȸ,�c�R7^��m��o�SF�	Z����I߀k(\�٢/�:V�WJ(��p<��D�8B�d}��&'��5�lJ�<�P�W�j����G�>$"��a�C�<�&�ʨppk� 2�v�Ɇ,H}�<�5�g~r1�i�X��CDw�<�ck�"U���2�@ J,��1J[s�<��C܅�\��k]�K.�����F�<)Ӄ����|{���
��&�}�<a��	�5�,���J�Z�b5 ��y�<�g��/Q�"�ȏ�zI�d�w�<�uk����X2*οo�^�%�)T�0�K�.z�b`���]t�!�l)D�(���U]$M�b]��B�z�&D���Cd�;�҈:3�-C��1�J#D�S���9�>����t�ʅc��&D���V�_�q�8���J�LTTc�7D�ೳ��-"�la�H��ab��y�!򄉎u�(����3�4X�aҁ�!�d�?3�E���lJ ��i��!�N x^Z "��A�vN�H��2m!򄀾o�T@ �-e�leR��U�!��iD��� �@�k����E��	M!�7^�f�"����<i2 "�z6!��Ձ&9FȡR�GQ�0U��!ʲ";!��O)"��-<܊�HqFF�w�!�D�"y~(Kg�Q�(zt��gŶ|P!�]$�Uy�I� �ᓭU% !�d�~)Z��E�=�6T��� J!�D�;M(�Z���u�.���k��!�� 
�܍`�̑0,�D��g*A�!�Dܠf]BD0��[�l��a7jP�!�dB�� hBE��P���çn���9E�d���GG��m���%,�6��ȓE�Z���f
��F�i���=y���id���S{^4X&�V�J1���W���+� �a�J��Tœ!)��͇��V�6' j�H�U��y?�l�ȓ7*�qC�I5z���2p�_�'�8��ȓ*�\����ͫ`y���M�oN69��r���k�O�*!B���Ɔʺ`�乆������#3м��6@kb���S�? �ݒV��/X��K�F�]�V"Od��R2%�,d��	�&��`R6"O��yT��J|��s��$p�4��"O��1��li�	+%�Թ+�>�A"O2�k�F@�5���1�%B?(�<*�"OH�����)"d��\� (��"Ox9�`� S�� �Їv���YV"O�	r''Q$c8�B#☪#�!�E"OR���
,�8��Aȴ�"O����Ą�	D|� ԏ*Y�B��s"Oh,�V��?J��Ah�e�hu��"O�H�����ӬR8�|Ũ�"O� �g@�^"J�
c�ݠW�Z �1"OT ( �=q� ر΋��f̳�"On��t���L�Xȁ���X��"O,�3��[6nz�M�U
¡b;��Z�"O��Z�I^46% ���ꄀ"9�0�"O�x`���>/�p@�S�?@ �"O���"�X�7�,#���[4Pr�"Oxm�a��ExN���3u����"O�`�Η+,�т5e͍�ݐ%"O�ˢ�/+Y�M�f�Z:j���@"O* �E��'Z��CO�݃!"O�yb-��RB� ��6"O��%5W�4 �K�c��)�"OL���-W	tD^<��;[���"O�}ٲ�J�h���pǂ�Ϝ%�"O֌��c��u�R1��&��d���
�"Op�#���Fc�Qb君���C"OVHb����j�LM����~��Q�p"O�|���Y 5A��P�"GJ�8�D"OZQr�B�?~����G��	����"OtT�EH�;o��Z�C�e�<�"O�}�R��5� �Ӕe�Ow\�5"O�����ϴz��4�Wc�� u`��U"OH��ŏ+zi2���ǚ'����"O �q$���nM���	1H����"OX�kaF=����.���a"O���"DQ�<S"o�N�,("O��p����1���Q5�
0,��Y
"Oڰ��/R�y��&/��*	��"O�91�8¨����&df,eKs"Ohx@��cp:�PAˋc`���%"O^eQ���"���
�b$�}K�"Oz�
c@�t.X���H|Z�P"O�0�$(9gx�� �_�8I�"O���ȹ{t� �QN��d��5"Oxe�S�X�tt)+矅.̖�J�"OܡCSGA؈��L�6�
�""Of�)��S�	.N`
�"RA�b "O�s�N N%��$�*0V|yT"Obxa�dX>+��PE����H�w"O���׌��Q����ëJ�C�v�Q"O��zG��f쐁b�U"jߌ��5"O�pC��^Z� �IϜ2���xB"O�B�m��%�xI�T(Ɨ��Q�"O���C@�0S���,�����"O6x��F&g8����#�V$)�"O @0���$YL�2�C�y�0H3�"OT�Pe�&y�A	��Qdw���"O,@�A�y��0�c��+v"O�-� ٕ}���3���;�� ��"On��TK	$%@��_,�д"O�L�WT�C�̑��.� r���"O� |���?(�!�3$�-S��j�"O�`*MZ$'V^�k�#�6Q�tY��'�����@en=#4�	�;#J��'�6����ɖx��e$�5�`{�'C�mS�Zg����/&�A�
�'@ �9����@b�B(z
�'<��2CCC)bL��L̚w(,��'|,��g޾Tc�a��*.�ؼ�'��)г��o�Bt�叫.פa�'��xCr��jr��D�Q"q��'����M�G+Z��vf�L��M��'������Cu���K{K<�b�'}��
0��d�<= T�� � ��'�tJ��*7�4��ά!��� �'����i{6�06�I��r��'��� �B�<�68�u�� ����' ;a��O֡z��#S����'`�-`�E<)/�KU��NR�,��'����mћJ"I���Ƴp�Z��
�'I|�;D�U�l�L���l�5�
�'XX�JR
�<8��%Q`h��MH
�'�Y�e�>=c��f�$�!�	�'\ZċP��+0��p3��
m&	�'sn���FĢ]V�j�k��g� �	�'Dn���*8��sO6jL=��'=j���� 
�4�
��h`���'����I�f�$�ƨ�\�<��'-�`�i��M��p�ٗ �V�H�'!!��n@u	 EA�a/���'n�вD������6Iݡ[��Ic�'�&p���ٜ3�����hɺ؁�'���o�#0�(`�d�)=0в�'���A#H�t��A���ژq�U�'pŏ�<䞸��H�j�fi�
�'��1��1�<��K�`��)
�'H���ə�.Nu��%W���2	�'��D+� ߝv�}��c�O�����'��D�1+�z]�$KdEF:�Y�'E�hZ��Q�:���f`í<�B���'�`�Xu-ћ1!��9a��7��(�'a�l*#f@p�hL"�h5���S�'Z��#`��k舍�0��/�$�(�'�lAñ� :lM���'�&d��'�a�k�L�Q��$�ٛ�'1hD���:׎ѩ�E;P�T��	�'>iI�S'� ���E���9�'�n�1�О?Qp���F8'�����'�h����0�D�e鉥w~�{�'��H��ǈ�{��iZ� ?k:p#�'P��X�i4oI�̻���_��`�'�`���B��3��%BQ��z�'ž9�fR�N��U�C��&4�<(��'������7T�C�\�+�v P�'�l�A�ϥ`E�"�Y�S�$b�'���H�#_�&v=�@��$I��;�'@�̱��D%i��;pfPPC�Q��'!��rű�xZ H��V�E�:$Q�'f��L�7�p�#�P�F'5K�'�8"�?V�$�` ��'Y���'y�i���Pne���ǅ���"%Y�'6D�0a�AF�� 1��`e���'OD�S'F��>ԆM�TFC6#~�Q�'@��0�)�&���i,�#�и@�'��D@e��b�I�T�݆ ��	��� �qsB�X�G!D)`�H�4�Uc@"O��j!�ْ;����0��h+*��6"O<E2��ț%oV�A�$^�]2�E �"Oƥ���L\�0�A`��*/Ĥ��"Oibueêapld�ٽ,4J�"O���1�,�HeN��"R��w"Ox��u�I�|���#�0��"O�P��@P<j��R�H� ��"Ol%	$(�.,L��� 4�H8'"O��p�*������i�7 �0��"O�`F��#\�Nl�R���K����"O��#��5o<rx���9@Ҙ�"O��q5i 8^����/�&�1�"O�;%�ߠ#�����j�RX""O Ԣ�k_ST�PdV9?�p�c@"O�$	�Fö]�Xp����>~0�2"OR]ӑbK�eV�jSdŇi����"OR	���d�|u��a�|V����"O$��e�ު8ڹ�bkB;F󨀉 "O$L9T�ԩY���Z<+;�)��"Oz��`��<'���⃉U���aV"O���f��&���#��;o�dg"O$䒧	��*��d��d�v��:w"O$�#NJ'=�TT���Ӧ9���pC"OXTBC醠8��R!O[�HY`58R"O�T�D�Ծ(j$Q�E�ӒB��(q"Ov��1�΄L�����[��@g"O�G	tL��&�O�3=( �"OU�aD�]fX��&鉌V��1C"O`$��>U�����N�&/m@"O.y��A��Ff��Ƀ)"�1(E"OT�+�fK�8h��)���?؀"O�1�O�M
jYp�W�4�vРp"O��J�/܊$��6h߆�~ �6$D�(�&�8l�̄#*�:O"� ��=D��!�C�.&�QaE�AT����	7D�����&��2�A)4МKg�0D�hT˛�a'V��01v�t0e-D��9��ƁX2AQ�끮u�v���&*D���uLU�2�I��F��m)D��آ�L�S���QŁ^9�4pc.*D��p%�v?�U�5��w�� �;D����m۹m\~��k�s
��[�>D�X(��#��A�Ӳk�z� ��2D����u(E��"r������+C�	�Q�$�s�@�h!<�Wדe�B�	>�ȉbf^ h�ؐ*�'�B��1c� �����7��03�e��[�<C��;��`�5GQ��� �I��(C�	i���IUZ����э��n�B䉏�"-*��S�9Z&��hB�hoB���ʴ&��"A�(,B��8 �,	��'!Y@�r��42W.B䉄eF���P˛�Q�xt�p�syB�əL@0������d3q"�Q;B����!��X��rp�&'̵}FB�I�xƹS3H�'1o@��!^I6�C�y�0���>0nn�a �g�C�	�D�b9��E��4����u�C�I2c���8�!��#V=�W,C80\C�I� X8�!a��+�b#�fV(6�xB�I��Ve���#b:\�U
�,c0dB䉍�uys��8N捙���670B�	=){ʉ)vA73�ˇ]�ZfB�)� ��@@,FaYv@�O"4C=�!"O�e@a�݆VHFAZ��B�5@N�5"O��9DK	/K�0*C;Xn�� "Ohl���!q��"�\31��� C"O2La����=�TI�b�5T�lD"�"O�`���@fQ	����H��
"O �a��0+Q ���Ϫ~2A.�yB	�8hКa���1��8`�[��y2��4
���	�;,W�����>Q��y2D�)<��ePeU-r~`)�� �y�%� �ꃅD;4lR���
�yh
�~D8a�Y�t�cҦ\�y�dY<{]���#����a�����y�˔�2t�P��L��u��q��yR�1:�%k�J��f0b8)ABƥ�y���P��Zc�F��
�"�� ��=�����ˏ3�$P�%˙	 a��P+�!��
VϚ	�0��yk��0���8v�O���dR�ZҮa�$�X�Jh~���S2?b!�$�nL�V#�6�:�"�O��DF!�$](cT()V�&\:���\D!�� u픸	pdY?5��!ю��!�$��4���+s�6Z@��C.]-c�!�d���8�#/��b��t�!��A��X9�MC���]���1�!�^�a��p�ҢA�x|ląȓt��w�ʉO�,��*�$gl~���2Q�z�N�1�A�w`�n��ȓ7�vA��*�5A�P��NB99���ȓ ��X{Vaہl�D=����/iv��˟x�'.M��ףMT�	��<T���'#�t9�K��p�^�h��{e&�
�'�0]�to��eILk#�I	�
�'AB�fe�x	� ΃G��P
�'��@�m�~��r��ٸ:C �b�'�(�qm�.~<�Kщ,w��q�'80xSF&�� �� ���ߓ��'�<ण�R�Y+z��(E��i�<A�m��N�!��AɿG�4��LGK�<�!�,s�&}�"tߢX�3��\���#�v)3&�G�<����
�;.
�A��Uz��B��?u�
&`�/l=C�I-hpQ�*@+z�z1ǘ
)��B䉚Y��B�n�3]���Ћք_Z�C�ɃK-v�QO�j�p���\�B�I�0A�Q�3�х!h8��#���B㉺]�4�Z&�L�.Ĵ;0��6w����'�a~�.�~t*|��D�+��y�
���y��J/3H��c�q�pەe�9�y�FR�d� -�Ҁ:-R��e�y���&��tI��;>�0Z0%��yR��Xa���@ٻt�T�$ȓ��y��	�@e�ϭn:t;4A[��yRɘaQR�!vy�r���	��?	�'�dJ�O��'�"�J�f�:4Nu{�'an���͐Z�6t DE�=+�2��'S,�P��3�9�[����3�' $�)u	;p�*!�c��*<N%#��$�<���)�V��'��f��AW�ߺ	�ў���J�O�Z�kue]��ҷ�G1kG�[���.O@�+���C���S�n�r��M�U�']!�dӴ:0�΍��l9�J
? ��w��yT��^h:�S��7#P��N<D����`C3��Y�I\�@Qjt D�� X�2�K�S�̨�挝�}���C��I�G�D욛�����-o�j-�T�����'�R�O�~IP"��qv�����8nT4��'�9{fOB%d�1�l[�cY�a��'��j�]�	�l:7��,Ԍ����x2�:��!��m�\TZ7�H��y&N*mI�6&�6Z���f�1�y"���-��X��2U�e���É�hO����N6(xz�����(`�PMݿu�!�x�hpZ�g� ;$��64��O���:�����}
DőF�Er�igO,\�Bi��ORp��t�E��)g�O`B�ɨI�^���%>JEt�yՏ�
 FB�I/�T���ؑUR ��P�A�"B�I;5��m�'b�(�(k�OY�l��C�IPL�!Y�l�0"Ǐ��Vt��鉲E�H X#�պU%8�)�'��pG{J?M3E��g�̹�mA�#�N�<4��I��͌j��,��'�5��jeK�w�<qU��/O|� c�	
M�B���Mu�<HI�8�l�A�n������q�<iV�_�uB(�a��34��-	��DA�<1�Gō�(���O�](�̠����<�`@ XTJqIVK�)-�8�ё��}�In���O���b�ײ�b�{w�U��t����'i>������xPg>-0�
�'@|��q���V�1=�*�{	�'��,�Ťa&��8�a
0)�q��'
=�!��2`�͵!��J�'�*���y�L[��
En��'�����X�y�LX+Ĩ3�ܘ��'��l�R#��[��e+"���$x��'� 8���m�>�fE�p �9���x�O2�~ؐBɅ�*��{q����y�ڢdp���C���$�Xeya�� �y��ӛB���R�[�#'l9�7,���xbaW�7c��w�F�,��m�*L��tx�l�'�Z��,9=�J-I���*X� H��'2�%)��ߥ5��́χ>G�MsM>i��?����	�k�╸�k"��d3�G8P��0?I�G��?��0a�bf�щ��c�<yV��y�p�0��R�J2�0��W�<��̓����6i�v`��	�k�<	���4�]C�
V/j�����'�g�<��B�'qL��G��"
v	K���?IK>���~�@��W^A�lƕ}U�q�R�J���͓@���h
=�����Q����C�I@����o
7!&���IE1$���bT�6D��x�+�n�i�#ą�Y��6D��fm��h���f났ni<�2D�2D�Ĉ ǃy���4�� `��.D��	�d�9��<�C&�B0V�)�	П���ӹL)�t#0�j�ĸW�-�f���O����y��M;�4�*��9��%�O&Ջ5`%��y0!ך>d���V"OB�c���N]�-�5��,�(M��"O1� �6Qi �� �>J��a"O�@���Me�����f���p"O��K�J��#�68R�%*�"O4x�&�K'@��5`���7|K
�bP"O����FU�<�vY��C�,3:"O��J3��5]u����
- �"O�|	5�Y6^��P�V�^|d��"O�;tO����r�m��#U~Z�"O� >�P&d�0F:�ub1�D
)I>Q	�"O p�qM��=Y�5"�ηk>6�q�"O�q��_`0�*�S�'NPG"O ��&B׀��m�Oʔ7�6�w"O����"��D?*z�� rԢ"Oz�EE��L)(D)�n��
v"O%�ô�´Rt��!9���Q"O���B��󅅌[ކ��"O��]�sO���1%�o0@���"O}��W<C�́��CJ��f`&"O"4+ G�;J�q毑�N$# "O"���Ըeخ|9�.�L���u"O�pk�'N�+ ���E21℅q"O2��EOL�Q
W.�VU��"O���CޣȬq!��,�xl�%"O���ω�|!J��J /�,�r"O�	��IH3x�b��E�EW�NI#$"Od���.��3���dGY�z0a�f�'���'��E#���# ��#�G�a����'Y��[���!���{�B2
��(�'d�����Z; �0���BV4e>Y)�'!n�@ƼaX��0)���H�'�`4���Ԡ.�<�8cE��0��'���F)�=0-�B$��Nd%�'I� CGm�0z��BD�;��i��?��i+��b#�@?'Gd1�á=p�5�ȓIu�I�
�qל0�'J7h��ȓ9Y�<S��v#�lܙB"�CK�<��/֦]
��ׅSء��Nl�<��'�"\����d
�m��ْf�~�<�����a�rd[+rl��Ĉu�<���\w,xT���Q7XdPyp� �G�<��"�5� �:�g�T�~�5�G�<�5��&@P�	��E�+:��!gz�<)��Zb!F8���P�M��s�Rr�<��kC�NZ������	Q^��珌r�<�
Z;f���މ=�捲B�Ue�<4�ӣA���q2'aܸ����K�<���:\�M��I�3�ր"*�L�<�`��p�I�k��:Q��OI�<i�b�=).M�5�l
���KC�<%�E.8��
S��SZ�LkEAt�<��^oƴ\skf���r��Vo�<� *0 q�����΁kR�����n�<��D�#KI.dqC��<�laz7d�Q�<���ߢ3Z� ����n�ؑ)���t�<�SH��P*��OE$B�.]��jCk�<��3�az��F���� �d�<Qp��&��X&��b�d�Ҕ�J�<q��9N�0����
�*�<	�w�C�<�r���H�:(��N�~�ܑS g�<����8�P1�@�S�Q�H@���}�<� �E�.U�}���R>������c�<a�	����5��#�tsB��e�<�A�L^c���f���=���Eh�d�<�B�)o<ڍȑBU�&昘Yǉx�<�hD�N����!ֶ\I�i O�u�<QV��@�6Q�ah�lF�xH�% q�<� ,�2eBsb̰�2�	��SD�<�e0p��AbS�mX�9(���T�<�g�h�4���KгW$�4����h�<���ʕ�� ����XEt��Qb�f�<���[�(�v�J�R,tiH��H�<ɐ,��/1�LC��9`<��ө�B�<� �#��(pLe�ч����{�"O��p�ĈfO��w�%_�HU�"O�J��Rk���r&�Q�T}�W"O&�F��W�Z�@e�D�����"O�)���Y9�
R��:�X� �"Od�2'A+�R�GP�!QT�[a"OP 1�C�����-_~ͱ"O�9�JK���Z7M�G���	�"O1I�
 SR���͟'̲�؁"O�Us�K��b5S��q�4P�b"Oj3��?q&Xt�3�V��f99f"OFE���UTC�,T-�r�B�"O�%Ђ*�5~��@3恌K���"O��K�S j~E�S������2"O�y��i�fL��M�	�px�7"O���gM�8�4b�,�	Vؽ��"O8����'m�v@�t� N8J�h�"OX)#p�]P�n<A��~����"OE!LE@c0�PV�<!�t"O��Gح.l|0�Gᅣ�""Ov���&Gp��0��I0Y=�m��"OΘ�T�C�>��=���y"O�y8�F�9g�v����
tX]qc*Op�!�g����]�4��&6�N�
�'���ö-	�u��ȑ�T��*uZ
�'1���c!�@n�8�al,A4ݩ	�'MR�GT��Fe�3��F�����'�h�r`�·B�D���KͲQ�ʓ}VX�b�	�&���Ƀ�E���m�ȓ�v<*ǩ
��5�P���!1숆ȓO�\��a{�	��!I�k�R	�ȓ_�D�ʓ��i-���o�Y�v]�ȓ0(��K��-%s,(�!�#p
�U��0@-�'-Z|�� �%����T��W�]��J 2�&QJ�e�_�d��A�xl���� Ib�
@mE��bu�ȓ'�r�&c�>�����H�G�`8��J2��1
��^�`����X�`�΅�����IW���h�<Liu �5>���ȓG�|тg��8>p��֩͜9�Ha���pD�5쇖,w�	8����vy ��ȓ.�XA�-�!h=昃w"4wc�܅ȓzM��y�9D�z���E��X�rP��w�4��c�Б"Ar��߄�����
0ٻ�@�6�A�k%��u�ȓ9���s��P{b:����(J����{Y��0.=v�F�0�)�~��e�ȓ)����v�	��KQΏP��
�'���Jb,�g���9�N�Oc�E�'�1�Ti�
r�|h�40y& ��'R���DD�4�v�ِ��04I�yJ�'q|42��n�����ƺ0����'�2��
*fid�)�+#���)
�'��XѢ�"AMb5���N"bU`�'����ǉ^4���&'KL�1�'�U "ǣ|���U�T�KNN��'�8TwfK�t�@���%�G��)q�'|L��T��3+~N����G�\+�'D��9�O�{'B7oE�l��'drC���f$P��2�R�2�'Ѽ���h#i����E�,v^- 	�'WzD��� <�2���M�0�h�*�'(屷�*i[�l�������(�'��XC��$Fh���:�z,b	��� :��j#\�l�2G�Tnt��"O�1 5�:{�(FD�x_��"OF��� <�\4��MCh���"O8�ږ �"��U�Ԑ<Ԍ8A"Oͫ�!�Rl⍀����#Ġl)�"O�)�ϕ�<h��yB�=w�"T��"O��%ϒ*>�>�!����2"O�I������mB�J02\��"O��;���	�n�Pw�=m�Ұ��"O2 ��d@����7-۞M��1"O�B�E��k�@����U�Ĩ<�Q"O"�	ҡI�i��H��L��:�"O�I��${a-��S�S����"O2�*У���CDll��M	�"Ol��
�"�$�Sg�
 �"O,��@ ,�����$��1ZG"O*�8t���q�.���CT2Du&��u"O��(g�:��|��˶rv��$"O���O�|�L�a��5
t�x��"OR�vmԜz2D��"jyV\��"O�l��A�خq9 :@q�̂T"O�1Ӫ��[x�𥬞6Q@�a�"O�1;����@e:�kZ�]���"OzH�N��J9H2��|�J�2�"O�x��	�4:t�	;��+ڐa�"O�A0G�/Ȋ�zEMx쬌BU"O�x&끑s�P��"� C��d�"OT�Ɯ7�tI��A�SSnp�a"O�aP��4<��p�N�B`,]��"O�%ɲ�$��g.��L0��"O�xH�"�5��t���X�P�T�s#"O�X��"[}@
�a�9}Z��F"Oȝ�5��m��)��YjeXii�"O`��A�8%`a��,��*��P�"Ox1T��'��%[�$E�L���"OV-1M	�u�`��>D�Jp�q"O��p��?e��90��B�!�1"O��0��%JO���j�#���b4"Oa;��\���C4* +��ew"O��� Ğ���5�7�$!9�"OM P��]���	����"O���jK4	~�S�pF��"Oҡr�I�pG���FĚ�Al8�"O�-���U�F��X��Bsd�'"O`QP��2Ӛ��7�D-]q��cc"ON��"\�`�-��`G�+� ���"Oаx����YRo�g��٘�"O��0�\pعb �'f^�ۇ"O��G���z�����o^9��"O\�%�PPp)-�
mP.���"O)�6#٪e����"YrBb�Z�"Oxue�^�J9��L�N�`ɑP"OYs�l��J���'�D�||��"O�U@&!	GR��u��\s���"O���5�ـH.^4g�=BU�I�"O�����O�T�"��ɜ_"e8a"Ö�����b�b�$\ 
4B$"O0-#Ԍ����ժclUQ�"O���6J�~_�X��A5�����"O��ysD�*���q�.�*��{D"O��;��2KQh(�R�ܘ]�tpR�"O�Bチ0F�f����*� e��"Ojp��іr���s-�./��IxD"O�,��MOۂL��:��h��"O� �y��ӴW�{D)pU�؊�'%�'�a|�h�#~�l��D�H\�2�o-�y��
$�܀�&�RzD��� �y�Z�m̻�Z�5�����`2�y�f�s6�cCE�>E�P��B+�yR	G�~}R0����D�D��R�y���%;q�L�L�8h�kV�T��yRJ�?��٨���x~���"5�?9/O���d��g`4�R��XI�D�E	M�$!��͡tS|XȠ�XC.�aA(�)p�!�>��0B�`F��U3gF�m�!��[C�\E�"E���P�f��-�!���(X��p8S��0���q��	R!�J�`�4QR7�#s�����CF��)�C��Ĳևݓ ������\����?���0>����~z�Ib�ί
��ڵ��m�<�w�B,`�J!���mJ1) �m�<�a)`�t`S�ǥ`B0	ti�R�<��Ɲո�0�C�Df<+�j�<�%@��3�[�)F�t?��2'(Ei�<�`c
���aF���F`p�j�'�a��dEX�Mrt���
p����y��|�$궫S��A�W㍥�yBg̕d��Ta"��JK��A)�,�yR(�=��Բc���/j0L�G���y2�(u��U�%f�Pj�	���߸�y"��3q�i�@���Hs��@Á��yRCK�SF�8��33���:C�ѕ�y2L�\>\����;wX�����yr����#`+��hV�M�y�ō+E�}9��װv#�R���y��#)�fa�⡑�A9�9C�υ�yb�3z^����I�P�ƀ��y�W�9�h��ɻG�2q1B��yR�͟i���G�:�t��E���y�F<R��;ED����$;�y�c�h�Q�����-�c���y� ��h�	��`#��M��y"H��sH�5Z�B�Y�X`�tLG�y2�R%`�4�HU ]*J�-��ǘ��y�Ęb�4bԧ<����e��yb�S9m�`�2e�B�j�������+�y��c5��$,�
A)�8�y���9%H"E{奞�Q��X���@��y2J��1��<ya�J �MIG)�,�y�'ٗ�5�vhڱE�(��6�G��y�ƭ�����4sr8l�2�I��y��~��y���dDθ{rh�yR��$je�ĽR�pxB����'�l<��/���L�IȫPl8�'g�-s�!ϥ��̸�LI(}E�Ej�'x��#�OL,Z�|I��ꆦ,�������˄g�X��h�z���M!�DW�v����2L.":�,�≁�U6!�đ$`�@ɱ,�,H
V,�"I.3!�D��`�0���̫�����
̘
#!�$/K���qDJ!t�ND����*l!�ވeՂ��A��*"�I"�\�X�!��Q �)��O��t4��$A�G�!��T  YLϕ%L�m��c٪�!��]V�1{��E	,���qD�т�!�D)Y8Y �i5ӺU�/G (�!��W�����N���:�n�y!�d�8;�>)���Ir��S�.R�!�� �I��V�T0���@�J�U:�"O�H�Uʉ�8�2��i�
(&"P�s"OИc���*@r�880)={��9F"O��*၃�UE��"��� �M��"Of��'��cX4�haF��r^�I��"O6����}s�5���$w�`V(�yB
��EO���Ӫ&At��EN��y��Q�WA���I��HF�K��y⭍
 8@Q��+a,��H�y�G�t,A`Uǹ�HI���&�y"�@�"DHSD�_0I�f,��Mq�<�0%E�+خ�{�ČnL-�^`�<1'�_;Vm�x�q"�$���w�<�r�B�?�=r"/j�.ȓ#�s�<ɰB��Ss���m�"C��m�2#q�<	�&LG�}�`0�6=Y�H	I�<2�9�ld��Y��`5B]�<���
u�6  G���soH��� X�<�%JM6,8V��R�S�l!&�����W�<a�Q�u�B��'FN�� �k�<��&��Q�t�zE�ԔRhDhh�L�o�<9��M��1v��2o>((�MOS�<Ie@֐Q���F���;O���gUM�<!󋉷\f���`^<ysx���AGM�<���5(j@YPF�7<~%�W�}�<q�	&~k��f�1�Cl�n�<��σ�ޘaBϋ~�ܱ2Il�<ɵ�'$%����.J����ff�O�<��ب+�l-�Ѐ�lxR䱱�Bw�<�QH�|��p�e�z@�LS2iQL�<q��8��w�F:O)T��g�F�<a��h��@P"��)�*lj&�D�<��ሇ.{�LA���{s����eRL�<��b�m�^E+�c�1���bHG�<鰇�w��&� �i_��x�y�<2�ޑ>q���Ѐ��)��@��w�<�Rm�|�#	�R��Db���t�<�#
�8*���H�)�y�&8��t�<�m�:7�S�Ɵ�DAk��Rq�<	/�X,�l�4.^�Tj*���Xk�<ѣ���g� )�쟺k���$�e�<����*!�����<RjL���\`�<��	�(�jȋv���@�"ׁ
`�<��aA�MPVӰ�4f>YR-�_�<I�Fɢn��]c ��3_�� Wi�\�<)7��
|����"Ζx�� ��T�<IM�_4H ���=L!�`�?T��ۗȄ���U��0<��]�wf%D��Rf��%$^1c!@�!p�/D���ѯ�) j�A@��K<^и��,D���Y�
DHqW�]� �j�g&,D�J7�L�ub:�3G�(�L����)D��h��T�4P0Qi���k $�7�'D��A��ڎc���T�hq���C2D�����z�S��\%`��)�;D�`BcU#`�R8�
��<�����9D�D0�l�f���IK�A
`�8D��n�	`�2��k uj�6D�@z� 	lA>8�e`ŷ ��N D����/��aIn-+e��h��a- D�t� l �#,��8h�����V�)D��p0Џh�^�y�R.�Q)��(D�8�%(O��4q�O��|���x �:D��
%��,dÊQ#��V�̠���:D�� P�83�ڴA݀��� J�y0<}2�"O"��b��=?z����M1%��P"O��c�KA$�]�g�s���"O��+pD��l+��u��T�@��"O�p���E��}�B$��m��4"O�@��CѸ-k��d"��*	��"O�K�Nɶk��,�,"��e"O�y��(��W��$SV�"۶0�w"OZ�x��ōlO�l�v/�l�2Ő'"O4t�s	�08�O;(��C"O�i�mŗ�Pp��.�_��1�C"O|��E�GeX��FY��ɸ�"O�-��B�>o{�x��V�V��<ۧ"O�-���V��G�K� ����"O���t����(�S��"O�Bh�w�j(���B"�>iz�"Obd�1ȟ=K�"�{U��o�*q��"OUA3�1u�05y�@,8tR�"O�L� �@G�,�z �Ұ-�X���"Oja�/TaAx��a��,g$�I�"OnՐ����;�LIZ $1_d�y"O�� �JW�)���k�G6Ova��"O@�B �\'����R�(��Y�"O��83#&tx9b�ƣ?+$=��"O�e AC�`0�����VDI�"OBB����0U�D�9��5��"O�=j���2sXذr�� �\i	Q"O�������&,��2@L��PU"O�[�g��d&t@��)�@���"O��Q��˿q��p8�b.'�"I"O`��B��5gcfD��C�[|��j�"O��{�
]�(�bbΗu��H�"O�� Î�:d6\%�� ��'g���"O���"gX�]�L@�o�'d|�A"O&���T�i��m"T�Ѿ@X,��V"O����œ(����̜NHȲf"O`mRQ�Y)t8RY�M�JQ�=!�"Oj\��Y��H�&�=.f<��c"O�s.\��8��^�k=@}�"O�Y��J�s7J�3�:/�1`�"O���m!��rTBׂ*vx-��"O�4��L�i{��["��6���9Q"O(���A0K�f�I�_7T@@)"O@�EP��hb�Me7tق�"O����A(<厱Hf$�,Q%�eE"O��mȠ9v������8$ay%"O�qx���Q�!� �%AV�Ѡ�"O��@�eaȐ02ŌJ�6oj��"O��b�D���4KL�6�`B�"O�|1���$)TYH�'�+ &N%#P"O�HRpc�,��+R���F0Y��"O Ę.Ŷ*>}�P��2GR��"O�AK��^Q�PF	?^�2U�D"O��GH�x8��wT�|��੥"O,j`ܻ6LrA��@P�i 4�C"O��(��T��5��a?J��"Ou{�f��
r�+��O2TJl���"Oj@����O4���PE���I��"O1
�� _CR�aց[2-�TTh"OT��'X4X�8��*<~t,�"O�pK��j����^^�MrP"O�x&��~�
yP�K�[{���g"O�E���W7T%*�˂K�xD��:p"O��9p�O�T$J|ё`�'��Hp"O� �5�WI�"X������v��ub"O�R�BՊ ����(4�tZ!"Of5��D̿l�ޱ��m@H!�	a"O���!"	6R�.�(Q��E�0��"O�� ��M�-��	iŌ��!���"S"O�@�g��0���ǐDK�"O@���!̠���� G��S¼���"O������>	��8���:5"OX�`R�!�Ix��L�c�&��$"O��� �w���\ }j0�iE"O�݁B<A1�\��Ɗ�_��Ӣ"O@�dԪ^9���E�yve(�"O�!�@�5
&�Y��-�b�k!"O�т�(�3 0>Y��U�N�ta�'`�h�G� }N�3Ԋ��v�{�' ��T%�5-i����.
�`�����'-J@��]��z�I��G��N4*�'G���5s�����-	�5�T 1�'/��s�;hZ�)Z�F�%?J���
�'��9ō

x��򩌅:-�`"
�'�"�����+b��!m��-i
�'�<D�Sŋ�e��ȫqmڴFx�C
�'�b���[�&��pBM��C)fh��'��T�±*��`���R�p�'�� �$��'C���EUFƨ9�'k��2�����%j*�Q�y9�'Ij�X�N�r���C7�ʶH�H���'I��@D[s��`��E���'\@l1բߝ��ȥ#��ްj�'F��a�C"pa��ŏ��`)J�'�~@2�Ƶ(���b�H	(���K�'��l�B&]>l�6z��Pu`�'Z=�+��w��أ��*}��%��'�2Er �۞{�{����ѻ��C�	��4�&.�1w���xW���C�	9n�&�h`�K	 ������j�C�I�1�0]��KȞR�.)s$/[;-K�C�	(zj6Г�%V�p��U��O\hrC�+St����SɊT�/΋NԮC�	��
��W�0�6114�� ��C�IH,�B��V-C&���n�K�HC䉈738Q��凍W�m��C5B�B�E�����LϦ���t��C�	��\hJ'\�2���"��C�ɫ`d񓔧@��ٴ�ؼ(��C�	q*U"��� ��4 2��;l�C�	#�q4�ðB�q,Դq�*B�	6{���d�݊ ��@P	R�0�(B�+i�d)i3L>�ڕ�a#w�B��9]*�wcϟ�9��MH�&s�C�	/ Y�3�"Ü��@Ƃ4��B�ɟm�l��U�X�8���2�C�I�P���#����n��)�}> B�ɉZ���w�V��DX�fi@�K�\C��)5��@�b��!�P�0�#L"I�nC�ɔ)�8�B��^�n���DK�X_\C��fk<Q�k͚�"���n!!k.D��i�g��H
�xҏE�՜�¥.0D��"`�+$�b�Άʬ����#D�|	 �#86�d�ףM;iˊ��� D�Đbi[�r�:i�E(͓`��@�W�#D�@OY"�� �
M�@�R����"D�<�1�N R����h��I�����?D���F�h��d����8��*D�� NY�� Z�0��钸Az�t"O ���D>,:�3dJ�	 � ��"O����Ճw�2���i��5�^��3"O,�y��
Cm������o���"OX���E���:�؅:��e�G"Oʽ�Q\[D��	�)�yL@kt"Oҹ���/���[p�]�'F�@z�"O\u��KW-G�N@R2$!�jL
u"ON�`��
��c�I�X}ٷ"O�S��;v��a��T��q�	�'�&L�E�N�o�e9��8!M���'�� ��c
i��&�B�Rs�'�t�)B�Se=i��Q-�䑢�'��T���ѱ/����$�୉
�'{*yʇ�(|d�v)�"خ)h�'ǔ���D��z~���@��@��'$�YB��H':\P��14D�t;�'2ڱ���^,M�T�M3]�0T)�'��4�pC�/"z��T��*�Y�'1�h� 9��]s��%{�ڥp
�'Y ��5p����a��"	�'l��s!��p������^��	�'��īW�=	n��BeY�CD����'Of�+"olHHD3ej\c�'9��jу�t��m"q�ڀ�`�'��@���)y�Ų�K���^(��'v�Hx�&M�G LȻw�ܶg���'sN��jE`P��jG�w�,��'Q�s"�@�h�1۱̏�>]PZ�'�B�P��/[B�I;�g�73�h� �'a
���Oܤp̬���+�C	�'����b��:�<a�oϩ#<ҹ��'�4��J%B�N(&C��I�x+�'��T�����iRBl-G{�г�'�h𘔥�#7�j,�ƭY�<I"�	�'�RE+ńZ9޸mIuN��B���'��KJ5%N�!3�\����'O�q:��&e�0�'��zV���'/n�tE_)���f���mj�'(���DZ��xم�&��'>���D�H[����߳L��j�'���*�	?�L�!	�8Ly$X��'�b���L��2�&e��NU�K��9��'^��k#O�2�D���ۇA�����'��I�Þ�&�N#�M�=�H�h�'L��M@�.2�|���MMBn�����Y�,w���Z#O.��
� Y��y"G��Q��!ᒌGjEJ�7�y�,��'r�ajU)�":������!�y��>_I�[�.�*������5�y�oM�nҙ�QMՀ�N˒�yr�}��	��/ڂ���h�jS �y��ar�LA�.�tl_5�yb`���6t�w��1��(P� �5�y2�s�0Ը���$���T1�y���0���!�ar�(A��y��
bzr�Jp�	�+H �!��yB�����d�`0 d��F8�y��2H!6�˂��h�٘���y�@:�X��\�r����ybh'S(��b�$[�
�̸�y2`�$V��!a�@��T�$��֢�y�kʅ7,����[u$)C���y���0Ip���!ì P��� �y
� ��!aQ�U|�8� ���B|h��"O�<����_���Rǹv�dw"O��#�N[�V��l��[?n�v I�"O�С�Z>tG��g��7:�~�9�'7L�!Bύ�z�ظ�Rg�C`�X��'�
�Q�E��j{4)��I\'f�^L��'�~1���{���k�
ܷ9t�0�'ܥ��H!8X:v�\�Z{�'�v�˰e�-"%X8P|8��'��A�!�@I�]�Deʸ>3^���'w�� ��&\h��'ô5�,(����v� q��5U$��8 E�i���Ez"�'{T�
�l
�.X�!N&U>�䨋�)�S��mF<�L���E("�q���;�Mk�'��(9�L�Se�0 %
�D.�X��'H��&�(��;D"��h���!�'�6(S��.bL4MbS�^�Z����'¶�0��;P�h"*{���
�'	�ّ�ģ<�����V�dh@�	�'?��� �ph4P;c�G�Jq�0y
�':���%&��_D��z�j�;����	�'c����&t�d9�H �,�v=�	���'�����"5�4Z�8M�L
	�'�v]����!'�VUS�d)/�,�{�T_���'dv0rQ�	�Z�v\��[<C�ܐ���̴D�1#�ٺ��"oO�����JZ��ϟP����pG�lf�e�ȓo�Aұ�X3t��Hڢ�ږk(�L��HhV���T25�
T�D��
k+��ȓ)@�z�j�Iw���t�τZ��}��S�4���ϻa(�+���,�T�Γ6Fb�<E�$�D�2aA�(�n�$]I揕��yRW�-�l"��"d�6�˔����yr\� =L�6���1��{� D���'�ў�zD$��K#�큂*Zj!�B���TY�� �����'�O��HX8g���`'�<B�C�idўb?Y�'���(R��8�Px	b��)� �'؎���� �r�4m��OӉi:"���O����T�v=qv��,�h(�w�K#�a}��>a��J�T�� ��"�H�8�X7Cg�<VFӤr�b��`��+&�"h�|�'�#=�Op>\h��A)%�(�9�C��!7��I���!O��B���2M�H򠮁jH$R�"O*�Q���x�SN��/>N�b�"O�Y���5�>4��M�
�d1Qf"O�-�b㖯5���c�� �xA��"O�����~S88���,{�)
f"O�EKUC.Zu��;bK��$c^��f"O�1	�kB w���!@�a][#"O!��-F45>*�����"��qSq"O*% �aL:E�2�6'J�@�5"O�\�Ѐ5@X����� �0��`s"O\ kr�؃X��j m��u��"OZ�Č֕Ub��:㬟�F�����O�=��V�>�"F8 �L���F�#U�����z����>�偍%Y��0`ʁ2��4B\�db��D{J|��ފU
�� !OK�4%�`��I�<�u���K��͒3È�c92TK���ɦ!F{���i��XR�H��60��
��d�t�p�'�0У�Ǧ4v�mчE��a����'�:�)�o˯sp8w��Y�쌐�'!�y{���iEu(s.,S��Ds	�'��a�H�ו���
FE]�#>D��R��(Z
��!M;!��V<�O��$�>� :0�P��d�ɰ1��'t_P2^�4E{��	{��P�poK0%��M��d�0K'�	ɸ'Kў��х2=��h5�&O��i�sjQ0 �|"�"}���{P�I�G�(1�H�X�/���p<!�O��'d|�qFEȽ
|f�#��:�"D����]���iV6ey����M\�أ��>v!�Dŏɚ`��F�'�a8�	@!�XI���e՞Р,�Ï�-Y��	6,#Q�"}z�݊!S��b4d� �^(*aL�a�<�&nP66NA#G�_&b�1��M[���=Y�\4
��kdF��1��b�<1 I9T��(&�U�l}�	Kw+�W�<�rO�Kl8����X^U;b�{�<�g�J,UY�`[�
�&%�P�!�A�<i�n	d"FP���	8x��KY�<y�����%AMн
�`q���E�<����>)�Y�^r���4��Z�P}�5�U���Iqy��I!H.1i؁g����mM��y���#.�X�U��=Yڍ�2�L!�y��&���
��%Z��B��<�y�.��Z�E�E���j�!E���yR�ĉ,8lTz�C i�6�ܳ�y"�̺�<����ԏO>i05nN��O�=�O���3�� �}����.�}�ĨJ�'-R�W�j��
�ܐ,t P!���7$F|MFx����Dn�)`��ƍN=�:y���"O2�=!T`�i�`�
����Av���D�I�'L�?MC�,(a�F�q��0f���:��-|O
b���2Ȍ' ���qE�0j�\Hj��/D��W��g� �T�r��Z�'-D� �t��=X T�# �gif�@��>��4��>�E� B�̙�ա�>4O�i��ANx�<a�*�>D@�4a�#	jqb/�p�<I���;�	���>DKk횢>����X3�\Y�B�эZ�L��GڣZ!�䚏]b葴� ��)��%u�!��G}0�E��I�c�(\H�V�����N`���چ��*V��ybK�7Y¸��'�3D��P&)��}c���?E��r�0D� �ec�]�h�%g�%<�ZIP�/ғ��'��'(�P�����A���"��{i��6N��pƉ�Z���)�� 5l���+�RL�S&�n�։���/{*P��ȓ6���2%D<�\	����H��Ć�Ld�Pǩ��Y��ɠƦ��i�N���M��e�$��+9�5Y�d�rՅȓ ��Qӡ�/.@������,3��ܭ!$hΛܬ#͖cc`Fy"�'2F���2:�3`h  A�'�0���v��`͆+,2�m�#�<$��P�/7K����!���r� #D���6ͽ"�6=14�݋mtr� �"D�H1d��X�r� F%��f��C�!���<ᓬ�e����T��^axeEP{�hF{�K[���$J_vv��B�T�j�n� ��I�l,���)�E�� �5G�\?�C�	4��������XZ�^�C�I~���FF�sq\\x��l��C�I#!ziZ����<d�jSXB�	�R��=h)���M���w�����\�k��%T͌U�R�^�u�!�_�`ܶ0Q��
�Xhl#$��T��)�'n'*Љ���9�p P3�S1%�V�;�'Yd�RQ��N��(`2�D��LI��� �)�1~�apQC��f
��8"O:�z����i�4�B"i���"O�5�����d��"��j�v�9�"O���g釉�l�#����M��(��"O����`�L3)1C�]�O�zX��"O|���vRr���k�?J�09Zf"Oz�X�cF�%��	^k`���"O�q
2OǭFGfe"rc>��D�8D�@9�+D;n�6MY�O�#m�r �56D�����Z
C��b��mP���5D���T*[�#P� B��a����4D��
`�N3���/J�{��M��N1D��;�Y�ƘX�+M�(S2d@�-"D�� d۠j� �i � ��)B�%"D�����i�x��Ȝ�b���B�:D���R8��8 p�M>�9�f!-D�l�`�����۝:u"�z�	\�7F!��pL�����Fr�L0&�I�B!���+X��;�-��c��8�R�B�o;!�d�48��d�$I�aA��3v�?2!�{r�j�`ϣ5�i�"јJ!�@W������,.!6L8b�M"s!򄟭\�4��X_�vCTAێ4�!��%R2�͊��H�9:#���!���(J@B#P5V�8IRdӄ>�!�D*�F�k�����.H��� h!�䘩w�����9�DcK _!�E�t]pI#;ˤ,pT�-S!��	y�EZ�MK�l�+��c7!�dD'��@�
ڛ!�(xR)D;5T!�D��KNt��e�(�I��QP!�CSduj@EƸ~��(�&Ρ)�!�$�1\�A�53fX�D(�#\�!��܀B��b�Č�:��@\B@���'�L!w�/L�0(��8n��	�'�)��� �#���Ca�~L@PS�'�fT�PK�O>�t�fڀxR���y�]��zF��&�ZĈ�4ؘ'P>�y�� t'T��� �u���+�'�<e���%C��!�M̆RU���'H�P�-�+�p�EA\O�8A9�'�<��Ǣ�|�t�i��A�r��8j�'F�=j�QJo�Xw���A�'�h'C�P��!+"�L<;g����'�̸�E�6?\Q����=2�m
�'�.�:DF�4_�n呀�7�l�C�'Z���WO�
Ŗ��fF�#p$���'���[
�o�lA���$	z�"�'
x�9�N�m.��z�ķruU�'�2ջG� �,��}�뚉�(���'זQ9�&Q#h�m�����Y�'<�S�?v�i7�	y�� ��'��a�^
$�Q���C?s��Di�'� ta�i�(P-�� �z)^���'r�u�A�ؠb
��U.��Y�,��' j�a G�'W<�T�ґz���{�'u �h��a��ã�#�0̨
�'���h�=1�(Y��ژ�Vp
�'YH!�5枛;� ��勇 x�A:	�'�j���JT�	,�]�E�Q5w�J1z	�'��<[6�L<TrTl����=_��'"�!��]147zQХM�ް
�'�L��W_M6$�hT��+�us�'�L��n�tԩ�C��;~w�Z�'�( �C[b�*���b-l���
��� ��B[�kB��E����6�8�"Oܨh�N�vH��U2�LqI"O8��1�N�j�=!B�����c�"O�ka�]4JK&� A�5G���e"O⁡���4PP[s ǜm�f)0g"O��#�N�
��yb�ښ0<�W"Oz�q���<��P �,2s"Oh9��.��I��<)(�5Z�"OLЄkP�Q�T����{�� �"O���CAR�j�@�`!e	O��ˑ"O�|�u�^�gaH�H0��Jݹ"O��{�l�6)�2]+��^�Y|�t�"O��֌@>]F,
 �G�#XTp�2"O�8�&��#5�v�s��%�d��""O,��E�"Pⰲ1L�:��Ts�"O CB�z`V,qU�B>KV�i��"OJ��X�#&HaBˋwJ��ZS"Oj�x�,�C:X��)��
��Ai�"O<�3��>{Q��js�6f����"Of�I5�ީ�>��G,ؚ'FŲ"O�����10�xtS)�X ���"OF �D�N6�y��Ѷ_(�$�"OЌ(��N����P�x'v��&"OJ��#M0�����'��I)�`�g"O�p�U�0O\*����ڲ1���g"O2A�7���vS�`� Y���ɥ~*6I��FD�O�| ���\ ��!��B ����'�}���� �ԽЄo�*Ȑ5+sܶ|�<"R�K��s���3�(|�\��+Ԛm6����+D�0��f¤���@�"'9�����O$D�!	ˏ7),i�c�>LO��S�fÞq#��kԨ��V&b��'�2���%�"s���s�ƀ�,�|=�%��hd���E�Ј%�!��X��A�X�KI�EP��ן`��O�³��" �-��/-§9h���jXI���*ZX��ȓG��M�0�)D�T��B��� RD�އ�.���hy����p
T��H�鵏	�W^x�qV+.D���r	�$f��&�Q1��U��O$p��mn�(i?LOr]Q����)d��TH�3c1�D���'�$s�#�?ebEq�kX�v�v��AaT�; �/
^!�ď*�xu{q�Q9
ST�+um��a�O���S�B�V�����&�'`�b��4DD>R��D�P�*�����Jv����1;�*���kZ�`�&0�Dg02X��C�"}��9Ol�hKH "��m�p��u�q"OD����Qp���y�oƉG��HѶ�O���ŅL�}1L����2g� I��-KR����2*_!�D�&L|�@�r��O
pQ��fJ�!�L9P�d�I�b\�1�إ���м\s!�$MZ��r"o�4'�P��l�lk!�dc�|�If�Љ<����q	�'\��$1jU�m[�G�%l���LA3�ޑr�^6uz PҶ�,�Ox���jߦ��3�I>Q�� ��'1$E�feT� K0�"�F`?t�%6���H\	[w ��aρ[�<�6JEI+�`�>Pd��\lyr�	�v\�զ֡s���BA��0f*:��6�,/Kj����ȽS��C��/@�By�d�	9��পI�UIn�R$mՓO��I	m��\
$6�����0$�|P�m��g����Em("U�rH�5(vE¦�\�j:25�J"7�� �V'iM��fc���a|R����AA���%IEm���OB§��dZ��g��7R�B�S:�`����E�r��aaG��2<8B�ɵe��vo�/~_H˥BN)_�˓��Uq��:�d`׍Y�)E�#}��"Κz���r�̽t�+���	!��+v.yz��@�,�.=A�%�����&uY��lR PFʰ���{��[����\���������?�#�$����4 �\����}�9��6+�RY3P�
{߆ Ё��c��� $�0"�4W���Ʉ�ğ l��e�Iࠩ���N'm!�QS/�.�A!b�r�(������JB�qjf�M"�yb!�8@%29��ƢOނ�ൣ���yBbZj ��m��^9����;F/<-����J�7��Y2���	~pV� a�ٿ]!�>p��J�"�
�.4j����X��pG��c!RЛ iB�dk�0�q^?!k1b�ɘ'h�D9���L���p �-,�[����;�Q�#TD�k�k�SR�����Fj���iS��p�+ue�h��0Y�f+LO`���ݟx���$d�|�ٙF��h�h��b{� ��dU~����W+��y"�,Z������MZc"O���7k�;���i��@Th�p�٭~�� �����R8D��@$6����+K�9�1�� ������9��Ug��	PF!�;6�����
Q��m\=JZ�K#���r�@F�f��X��N����dπ�"j�x�y%��-@ֱ�G��D���x�F�,��=AD�ˈTi4�"�ET�(0���H</F:%c⏀{��ģ�C�/�"���$R1 �̠��ĉ<H:�7�O=p�kB��Zܠ�+'";x��?�t�G.u��K�ϑ�8���WMLb�rQg9`O�͠��$XdC�cC�@'�`;���I0S�H���iC�i�*a���+# �"r'É>0����S�)��b/&p8�С��.j�&q����3���
b��T���Zq пL�6��1O>��-���������`<	@���Bz��X:	�����U�j��\Pd� "�� �>P���{�L���P��*�G��}�$�]��D�3���۠	���-�O ��灓&s$#��8W���G� 'I��-Q�n��#%O\�r7l b�d
 ��Oh3E ܨx�ʀK�ܤV}fuH�cMb�A!�)L9&<�Eb�OƘ��S�tCd���N.
�vx �il�Ӝw`��;u��%D�J���f��7�,5ˋ�D�v������Ɂ�:{b������a�|�q@��YW���m��P���BJ��u���;~n���,��`���<Y���@Y�W���,VP�X$�S?�"������t
�(\D�D��<1�"�D/V ��n�����(5Pa*6AA�ők�f�H���VD��'E,^��¯֊9?���P��e�	p*����'��h�C�
{�\��'�) �F��z��Ř&�������ܭ��j��>W��@��3~@\P�=��P	޴m�*�`�m
XtX;�O�MjP�&M	S�l��O�̸�m�$���r���i����ɍ*޸QB��:NT�![��ɩ
���	[9��Oqa�i
9�(�4 �Go�&:>z勣cT6�z�KWDÀz�4I�sC־8=L�x#�W�wM  ��$=2n����~po$��,ٻ$�����#9�I��a�8NȄ�s<O^9�n8����~
�2d�\�<!�LS-S��q (_�jr�l��@�C�:�ReH�5���f��'^н�O���|���i�H��
C�_�� �CO�=��0�&-/^�4H��܂>���#/��i�@�'(x����^�gբ��2�>+��I��۟o�+ �i�&I��C��� ��o��'��$��|�v��5j�>e������	RH��U���D�]���	�(��!��'����&{�7�'"*�(��*=dB,b2m�0z�����_�C���v��-��	�6� X�3��_|�!Ư� �(��8#G??2���h��1y��'s`��a�z}�I
J]���cC�_��?�I"��iڠ��޼H�:!)%��"��)��Z��?�dO��TN��>�O�����3>�m���yb<]�#dO�YI�%�lP���)�'�u�d� q�����fK1@�|	���"8j�Ɉ�=o����4r� ��qL�0�QCP�G	��I�q�J�KǉO��s�^�+�G���H4�'Q������&y��ܣ���D���K��\����OX p��&L�" ��g4��>9  +54�8��
�ȟЉ`Q��:m@ ��	#j�d�!"O
��+��
�M��쉰fX�X��H�=��ݔ'Þu1�b�g�#aYի:vǌ�g��6N�C�	�Fj�%xL�.�(�����+�5a�F%�����'�Ɣ����?b�beK����ϓb�fm[ҩ���$�	%�xaP1a�G ⤂�/�E!�d�U)$59�Œ�Ę+���e�!�$E1z�朡P��
�21[Vl�3�!򤂞v>l� ΂%k�:�jv�X�R�!�d��F����f��I��顲��2!�d�7Ly�y*f�S�y�x	����6!�D�;C|h��ǥ ���Ӑ�ݦik!���gǢ1J#�3R�������Y^!�d��W���iA�6"��"��&2�!�d�-]�0�IǀQ�a �ћ�ż"�!�ą�%���8E%D+nט��&:Z�!��({ߜ��,2 � ���q�!�dF�%�|�z����/qD��S1M!��%LgҸ3���� Eĕq�b�>!�D%��UQ�ች����K!�� �I!�I�t��"�Ι�{ X���"O�l�3DP*b(�y48 P�5D�0zȏ�"��)�(hs0����&D�����:zk�=� �F�+�>�+�d"D�`AI��p��E��)��`t:D��{�JE�0d��!�+|���Q�8D�8Ѷ��V�h��SM m:f�q%�7D�����6@�.EZ��LX{� /D��˖���X�1i
|	�e�S�,D�,���� /4l�&\f]�H'D��W��(0)@)��l֦O��؀�c&D���RkSd���0��=���ei0D�h�u�"�p�n����2�I3D����A؍L���rЪ% ����.D��q�O�C�h�9V���Bm4�20*Od5�t���?��(�@ΣT�`,B#"O�|�7Ě�P��jO�.,s���"O(a�YD��;�a�&���w"Oδ�E�'o��ź׮Ml$X��"O��@���<� �OU��"	�'"O�L�0+
�^���׮��<���"O�Ճ��&$� r�oš 
�2�"Opl��#D42�Ē��$��a�g"OE;� VD��5��:�.$�"O�e�W�����UAňEZ
� E"O$��@
0m�$ȇ�F�5�V�!"O�a�*��ȔJ�$T*��3�"O)��:��8Ji���R�"O��YąE�T����+`%>=�"O.�:�ӓ	_�IZ'�DO��u"O����3@z8�gh_ R�*3�"O<X��(Ԭ)h��(�� ��Q3"O(41���p�t���.�=����%"O��*�a�9*C4x
��Ѽg��R�"OD-���ӊ}`�F MQ��2"Ob�!��B�\\�󅏕|6 d"O�x fΛ^|��Ӯ�|�����"OL�
��%4��`(G�����b'"O~��I��h���[1���<=h\��"O"I�s,L3V1�!e�H@�IA"O��u/��l,�0G[B��5	$"O���!*�\��iH�R�P5�T"ObiK��ښ~ٴt��)�&��"Ou#֥�2�lTK^�z��p�"OJl��,�;M���94�W�Ľc�"O,��!�_&��ـv�UD�Α�`"Or��#[�lo����J�l��1�"OF�����Wpx���hŦR��
�"O�� ���?����g�X����"OJ=[��v9��QC�N�ri@���"O~�V]H��"�Y�QM*�"�"OL5��]���b��0J)�a+v"O!ၩ��i�*��Xz�ir�"OD�iF�ߚ"�2���.̛0m��Y"O`x�`R�D	Z���C<��"Ov�)��ֆ_�^2	�E$�4x"O�%��;�"��҉&-�&"O�\0��F:(�<�E�U�Xe&�@c"O��)/���� A�yH�"OKI[�1�F+K~b�B���ybo��%Ę��"��z��I@˅&�y�C�1rqCp.J-V�E:����y��N8W�V�8��[0o�"ya
�y� Ý13@&CZ@�p1� ��y
� �}�7f0�ҦJ�)JHK6"OD���  )΀��#��E
l�pD"O<�@�Gͬ���H�:>4+""OB�0t���b.����&Ï���+B"On	����W�\<�3�רmH�C�"O� ��+KNx8`&)�7T!���P"Oh��2Ϝ+5d���DK�)����"O�0ƅS�<1�#�͜v��(�"O�99�H��,B�4KQ? T��"O� S7@x � �B�|b�=#"O  su�@�,�2R�W-UjR�[E"OB�
�3Nmi�ǝ�`���@"O0I���$�8`�B�i;�)�"Oj\�.X�pƑ���8;#�]ې"O�P�)��T{V�&y�1��q�<��R�e�I9�,��6LX�h�I�<�M�]�\a坁:֦@Y��I�<I���W���fL�'T}�pp�AS�<�/�CYD ����\$�����q�<��^�d��` �͎c�&P��P`�<�F �0`N�8R�G̼����Y�<�Un�0�ƀ[��L Z��{3�JB�<@b^�&�h=��jǥlG�Ek'�C�<AӡCq3�!� ,ωm�zYK��Jd�<�1@�VƄR��,w���ĈD�<I�G�8W�N��dٮM߈��d�
x�<���46�`�vM��W���32��u�<���V�<hl���b y+f(�[�<Ѱn�rhvq���#$5�,#���R�<�q��.2UR�Xu�ӗem>Y�J�'����Q�U.3T�>��H'"s��q41�T��C/D�,94��L R��¦g�<�Y�&��Bgy�T D�S��yB�Dw��B�B����G��y2a�*-�����,���E�?�)H�s�.�poB��0=1�i>]�}3�F�H0�:�/
k��<���&�r��>6c�� ����Ĭ���W$rk$��bs�	@A�y��P�
D!R�n��?9
P/7��ls ����؉SC�Ha�l���_X�X3"ORab�̒N����쐜O�c��'%��� ��m��	U��~@K�K�5�gD�Q�@�{�$���y�H �lqw`;x�r1YpÇ:�?Q�Mq�����W��0=pk	4O�(f�:
�h����R��������.*	A뉴8X�"�nO:(��d���E0#;���ȓTuR8�֯��a3�X1�CG9�d�?!g����H�߿��4d�" �!�x�a$D�HvƁ��"O�}*��Ɯ#w�`闣�3!ˢ��v)X� �f�"���)��<I"�S4=s��ɴ�\��ک2e�WT�<qp��.�������|J�#�V?iP��-&�"(�ۓCV���ЩQ���`��-P�Nd�ȓo���zu�:"�f�3'�;}RɅȓ;��l▣�<ZH��&��2[�`�ȓ�db㦁$ÚP�щ�@�^,��l�걑�!ݤ-�� ��]�IZ��l������;M_��@�+G�k!~<[��?�L��ԅȈ��>qeʉ5�T�8U�݈H�Y0�ICl���䊇(�BTm�(N�d�$q\���@���VEG+	�!�ě6ވ���2�����7�剖.�XHf�L�Y�X����E�O4riA�'1p�8ԃC��pnR���':���d	�#�� �N1wK��Z#��#{G� (�� �X0#d_���g�7)<DP��O;.����$jl�I��	�5.(t��� }��i��6T� X�o�mP����C.i���+Mm`y���d��Z'�W�L��?�U��TT ���\;Y7<5H�O e:��}488�������
�'��y@�^��Q��v�`*Oh���F�}<VP���&uX���� ΍˓��3_�@y��2D
��I"O|�@�,�? � a�$_�vq���	1��pأ���b�Q��/�;�ϸ'�.܊c���R>�|J0��kX*�X	��$Ĳ�:�X�I�:
�0Q��Y�YHtЉ�j�G+��� ���0=�Fb�#_At���+���
Db	h��� C�*�|L���T"ATiq�QZh(}XC���.|���N�@B�Ieq:��v&ؼSB8�v�Q�EL^�'"��`v�ȣ+����b�O���G�D���x��Dru�^�$�mz4���yB��h���؅L����b��p�|e���^�[�Z%�H�"~���nV4:¬��` K"fe�C�ɰ]0伲@�5C��I��*	;��	�e�)���T[azb�#1<B89D���w<��huMV��p>��b�7\'�y@��4t����ɞ4]��s�^4S�C�I�SP!�ץP�Z��mC�	�pz�<�AׂU\	��0�'kxHt��`I(A0�D�3A
�p��\���:�9����p���B�,�CpS��pi1 �w���O|�:S�P$l��4L{I��J��y��[/������ [~lD�D���~b'�% :���g��@��/�p$U"�,�aE?�O�@�LxX���Wm8JY���Ԫ0-:ج�0/��y2e�j*d��L1.���h���(Ot��Q��i l����A�H�X3-اo��
d��h,!�Ė2q���$�jq:����AK�6nQ�Q���RG�|���i>��#�lΊ���f�̓w�̍�����xE��h��TP��GO<l(�
�I����d�=�5��'��!7c�� ��l�vaĳ4I�1!"�p1��O�E��O0�v%A��ͱ�g��}��)�//D���f@�Q�� �����4�[x��S
X�ه�ɽ0=4 `���5��y�2�Uϔ��M�b���Ň�2�y��RC����� ^?��C���M�B(�2ހ�"~n�x�ڭyEˇ:�0����PN➄H��_+!��������yt��8K����.�R<��A�O�Q����6rc����,i;n�"�G�H~b��"����v��,��E	�c>�8d�G�F쩋5m�kN���-B�����8s�|��U���BG�p�ϊ/|�,Se�]�(,lDAp��<�'�0P��%���&}ʟ�q�CT�Z�"P&N%+��ZRdF>�'��Jr�~�`L�O\6H�դh���%�(v�\8!���!�u˳�ЙRY��a
��S��M���P8)c� Z��֧fN\�˄ojd ��b�K��j特M��M�6�P�*g�S�ӑw�yЇ�C88�jX� ع[��	��.��S�G�b�'�IX�G+�+g[�,�����3��*,a0��r.�#+\*iH��|bn,�S�.f$���.#+[ �K倓�O��J��;`v}s��+}���}�ĪFnLv��?=
��G��ҥ�n�H �hP/�O~�*�i�*��DF�y�
-�s�W��)�Vcܨ,A�� ���F�@�Fҝm9ґ�2T��*�G"N{q��'��qc�K042 ���7Êa0sO�41�s�aCP����K�eR#v��TI�	6�2�*�$T�5T>	�� �K�@�� �A�0�
�DY�/z���'��)9�%A8��'��5iS�@>�~��S_������50�|���#T��
0�2�O�D�5 �%�?�Ջ!�&�.%��p�e�:ep�'ij����3q0������ɾ��S���"�r4"�i*K�,C�	2��� ��0,&�8����p��<��(�9���ؾ0L̑Ӌ�L>1v�eM��#��ׇ]Ӥ��DaXH<!&�����1�F8O���� �}�QaJ0�j����?F|����4?��X[W
 �S�y��Z4>��PKG����nD9_�����
s�<Fi;D�(��	?���k�d(���U`"D�t��aĽT[��DmȖJnh
2D��9G�^�g~*��3vd�4m'D�08�`YQB�)�O ��ծ0D���֬�GY�<�p�����+D��;0+��zDf�+CYfU$L$D����TU���z���LW� ¦�?D����bS�C���@�DCĮ�!;D��AVlK�V����$I�g�@M�EO4D�h�ԋ�!pO�D%�#�J%2�/D�� @�;S�H9YzZA&"�?[a��b"O�4��ƒ�6��BBCi�lµ"O2Es��?h�J������12"OD���Ͼ��3��[�Dm��"OL�K��&�ڔ.^�=�*1"OnY��%��8���-sZ͙�"OΨ2@Aۗk�(��1&se�U"On���p��t �.{��(�"O��.YC,�A�WcRl�s"O@4 `HQ;B&��QF-�
Y����G"O����X��1k�ѹa�P�"O���T�b�dؓ���
�v!��'��0�Ń�z'p�yu��6KJh��'6�U����s�>]�a��!s�		�'�� � U�B����adȬ��'x*��Y�i+j�ᅣ�N`z��'�mS�F1ej*X�9��Y�yƝ!�Pt���x��U3%](�yB$��&�������y�����)�y�F�sz IIw�?vGF����D�yR���	�~q�5+o�l�8p���ybN�"�~��K��gTN� B1�yr#&j��<����Q�`����yBϔ5���:����i�'�S��yB�q�İ5$�"���ԅ�y�-@�YZ���M'$*t9��
�y�FÜo�� ύ,&˚�iB���y�`νB���a���hk����y�	C9I�uQ�R�"Li;ӄ
�y��N��@��$BX�	v�s���y�H	2� =q"��
+q1�J��y�g�H�雳��H3 yP�\��yҧ�7!N��ئNވD����oZ��yb��BV�TС��O��Qy���y2bωbF�8F)]+@�����Ǣ�y2J	_?N�!��E h�B3�[�y���_���,��M%$���O��y��K/7'a(���Hz
�C⬅��yB���sS�HSj̀3CP9��h��y���V���׌C�6䘅)��� �yB'RZK	�#T�E�R�qwV��<}r��"�ȋՆ�8�g�	�]�ȓV�f�#� i�Ж��?	%�Ȅ�+�� t�*��PжdZ:�t ��8�V� ���E�1���ǰW���<�b#F�P���c��=]�U#d�ـ/7`0Eo�?��� � |�Z����z5��'�
�� �m�b��x�)§/ra�W�\�L���@jJ�.��|t�����0��S�O�
aY��͈n�l�Ն�
�&D��PU�ވ��y
�'kZ���
�kw&�8u�P���Q@̓u�T��(`���`)�5"��0x����@A<c�4p����ا�Od`�(Q ��Xn�M�B��V���O޴��'JD�S�ORr�ۥ��$6!�Dzc#u���'��Ij�
$�������Z� _� <�s��36��h���)%1��e�?Ep��0擆N�֙2ǋ	:���{�˙.�m�4]���'K�8̟JЩ��d	RS�p�2$�(�����\*��D�Q�"|�\�5��(J~j���k�<a@�Xq��h��4����%lc|��D;n'�(���:Q��壛W�D+֬IG(�1�F�E�'`�Y����:Lᥡ�%S�H�� K�I��a��)��Y�q��Ax��ϖ]w���P�R�F�-��<��TE�(u�P��s��M��u��Y@?y�b%��?�1�}� ��?�R< �
�*sF�q�[)Nm��
�>� ���<E��i��	_�vP���_�=��`Pg�Δ!����'�(��$ú{t�q]w(Q? ��9t�eA�"@�ew���e��̩�K2 �(�äE�(�a�� ��bU"2���Zq�=��M�bnۮV$�(s��/��L��O?�� �a�"삯5
��S�&� jς�Q!]�.�,�R�`��Tsç5�(�I�P�I|��@�FN��R3�Rd�
��'4Xt� 6�,J���q��sU�K,�bE�s�"D�L��+r]�dI�0|���@}�I#r��<������G�>��e��ݴ"FN����ٟ�|����2Foz��Uh�\cT�����3�B�	3)�	2eȕT�HIF��,)��B��3n�n,���2W�L�I��P5�dB䉴����q����E�O�8�FB䉠lE a��p'BL��iφt]B�ɦtd�XГ�٨c��k�k��v�C�I,h�|)�Q���v�u�,u�ȓ]Nd�DH	xŻ��ǜL���mGZu���͡Z�����)�>~��u�ȓq|�x��jX�A#|��,<*iM�ȓ	,#�,Y�Bq���� }�8Ʌȓ��{�̍�C�6m@ƂY�p��0�ȓ��Q�튿!HV�c���5R�:�ȓB��9��+lV��I6b4CEa�ȓ|ڲ��@��[r�) E��2M}��ȓ}�p�c�ِ]C��Pdȱu����ȓ\P��V,��k�n囤�-7��$�ȓV�zQ P�ْY�lc���&w?�̅ȓ]���w��y[��B��#*�V��z�@��k�mf u�E I�u�R���y�D��唞z��Z�l��`��.����rD"�Z���}��5�����B��b1�3��1_o�)��?ʜ�/z�2���oX�(��Їȓ VZ����0%�84�b­?+����j\LVb��qLH-�$�V��V��ȓn��e�hӹ&`x�*
�w�䉆ȓm�,(� bX��b�(	�p��@��'� 2C-�NGM`�LI&�Ԑ�ȓIن5�d�_����`pB��$�V��ȓ/?�gg�#����lǭsb��ȓ|��h�0	�*���h�(`����*�l\Ձ "%���r� wx� �ȓ#R���$�@3+X�ʒq�@\�ȓw^�L���1�t�y���Y{�-�ȓ'He��_.+5j4�vO:l8���b��m�AJ��w����G�=v��Ї�!� �Q.-|��f˂�.�`��oZ�x�R�0�S���4$����3&�|��hJf��@��3b�����c
H��!��g�\�3�#&F(���hf��"m�P��,C%��q̀D��Ig6	V$���������^؆ȓ7 ��xc!э64���Ϝ%�B���z��|(  �a���"�kܖj5�Q�ȓ]��h����~A��[ MP'��h�ȓ�lL���,c�h�;PM�YF���xy��	�!Qv=���^B:r��@��%�&��m�f�&�4Q��k�t���˓7��Q4M��r��ȓ�N��� RG,l�"h	��jI�ȓ)pz�������όR�P1��g�j���Ř
Fٰa��jZp�ȓ5:�5�Ce_	.��p��?zч�0� ��LŒvK�8�!�7[<���ȓ\��h:t�8p��͢r�X�� �ȓ{�,�h�bּa
�D�����%�b�r�C��H2���y|�����$hդ����ա���y�Ơ��S�? �D	N�%���! M�H8�AB�"OJt���L�A�'�M�&1��#�"O��2L�9  I֡�'"O�=�6A�5�dH�u�H9D
�Ъ�"O0�� #A�c,pA"�e¨[�0�*�"O�y��I�FG&L�5���UB��V"O�]��/�K�t�c��4�$�h$"O.	���C#)ux���
l�I�"O����$H�<Xc��%���{1"OD�qw�^"":��!� � �H阕"O,��i�6����Y�"���� "O2�ZPd%j>�չ"K�I����"O� ��葵P��(�@�K (���B"O�I�d� �����˽zc�8�"O"��`ʭIԁ��EJ�W8��'�^�ka�N�"����"$-cz]��'�\���i��Zcf�
k�o�K�'�nHx�.T�w�2���z�r�'�(〩�({��%�P�M��E��'� 1C���_�\3�K�J6�1�'R؈���qA����I��?8�:�'H��@�C� u�^�l]�h:���'����1��[-����[a$dz�'�hl3FׯRd�{%DA�O���b�'E�1��B� ����FS���'REX�+ P%~`Q�"I73p�b�'�T넉5�$�`3-�%0�@��'J����V�W"j|�C�(CAk
�'5�	�aF�7>p���F�N�ܨ��'���SD,ޒ�H��$�̀D�A��'�BȊs�	5$ЎF�&���'TA*�Ɂ$X�4�hƣԣ6���'w0����|?�!�������'��=�D��%:���3���Ƹ�'M�t�2U�^5�	! Oؿw��i��'6~�+��aa�Q���^uk��	�'45��.T�ܤ�pw��"@��L��'�j�I�H0��)���;���
�'a �����>^r)�c�18Wx	
�'��U[mՂ-y\�c AӮ: PY(	�'�*EZ�掻"hܹ�Y_FV�	�'k��c�MR�A��lZ�d�=I�� P	�'�`��ț Y��ҦNBI�v:�'�8"S�m��옶�M�G��'e�Bc�J�{�6�zv�D+Е��'
vɡ�H+ayvd�/ �4�z�
�'?�ԛ" 4djFX���Eф��	�'�F��Æ�M�p����R.}�	�'5x@7�܊sV��+cÝ�~�\��'�*��`�=l��3̓�D���'��x'�%fN� )���'C��#�'����	W:�5#���>8�X0��'/d��DFAxv�uA��2S�d2�'.F��! !u�	�$G(p@�	�'ެ	���
����O�q�r�i	�'r>h��U7,�x�5I�m`	�'Q�x���߲����
�X(x�'����h�*����UJ˩�M��'"u"q\�+*���ui@�x�`��'V<��"�/E�&��U�8e;���
�'��bI�.Vf���s'�X����'o���̚~��TT���H�'���E1pp�Q�T�Ē1��X��'�$��aa�1Kr0��c��	Ag0dX
��� H��/ء]��P�Lo\&8��"O�0�����aR,�Y8X)�"O�@�E�F�G������?���R�"Oҙ�#��nͨъC����y"O�t�` �0�h{���B���J@"ONe��Đi\�x�|i�"OؼB���56��Hc0�\���i�""O$������B�н�(U�d��!�Yk��=X��`�8�`u�ѯw�!�d��A��|��K�5z�D��@��%�!���z�ً�F�a��)��/N�!�8J��]�sHNOȬX/4�D�"O�y2��.�|ǅ��W-��1G"OWg�5H�\T��(�0!"ONq�0�I� t�vC�'"����"OX�΀�A�B9�T$-f"�=�%"O���g6�*�L� >E�"O�����"�&h�'�+p@LP"OdAӢl��0 ��P�#�h�~��f"O�-ivB�?	�����?��]ʑ"O�dhWd��CdM"S�^!j�IqQ"OX*q�٬���˲Ϙ�zg�(@�"O��[t����
W�/a.0	�"O��c��2g�`A0�P&
�R�[�"O��h'�	�h���`�����h��"O> Q��FkQ�P�g�t��\J�"Oz<Yf���.Isb&Q��Dp�"O�	��J'D�|B��&ȝ �"O�T�E
�g)Z�aD�j��"OTD��iڢ�R7�L&+�찳"O�=�6.�3[�Jڶ(`��=x�"O}���۽ns��37Ҿ���Y%"Oڽ�e�)E@��Ҥ�+ D�R"O�Dsp'C

�:Ux#Λ6O��9!2"O��gg
�:T���ZNz��a�"Oش�DM�3�2e�qk�=ex��"O��+deU>=��DS6��`���"O8���'H�2+��q�`I:�p˦"OF���dS8Q8�x� <0���t"O�}ؓ�Ay���qᡍ;d��c"O2<+ä܌Hs|!�Ca��tWN��0"ON�@��H����	�sL^-�g"Ot�c�k���[�FHl,�"O�3�O3C:�� ̏�.3����"O]�"�ҰiN��9ǁ@�e����"O`Q�q����f�A̰!�,��"O����hMt���L�q��A
r"O
8!э��Lr4C���n����e"OD���Ƴ?Lع[$�<H���R"O�Q�C[�0Ⱘ�ׯK!$���"O��;��������m=^��=x�"O����@Cc{@�
��^;q۠U�f"O(��DC�D�l��î�"	�����"O(�k�g��q�s�ݨ�M�"OșQ����5~���g��l���"O���_���]�K:H���1�"O�k$Β{�d`P��:Ƅ���"Or�"��f�N�
+ŌV�`Bg"O4�XF�+��y����<V���"O�u�% �$7�U˃�Z�1�X�3g"O�%�ˀ�:��M�6��ʐ�`"O��)+l�X,ʧ$O��"O�i���9	v�|J#�^
k��a:U"O�KgH����h��À=t���"O� �x��F�9S|�c���:<HM��"O��.A+�4���D�A��i%"O8�)�b�h�Jܘ�)ߚMk�ȉU"O�=���5j��5�rJ� hF�b"Onͪ�G�
\�d��ލ-?)b "O `jqN89
����� "TI�A"O,UA�N�I�b9j���>TSV"O>}!���k�D��D,h��)'"O�)f��T* CV�0X6|��"Oba҇,i�Vq�T�Z)[���e"O�P�	   ��   �  >  �  �  �*  �6  eB   N  �Y  �e  eq  �|  �  ��  $�  ˝  �  g�  ��  �  <�  ��  &�  ��  <�  ��  ��  :�  ��  ��  �  � j
 � n u! �( �. �7 |> gE �K �Q �U  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01�m�{�0Rda�#��i$��� NMӠNF�<(�������zVޙ@��	L���)��uv�8��� �	�"�Z?�!�d�2DT�З�J��93g�D�$�qO��'�?�p���ZD��+v� $�����=�騟�2��ӬCp�����k:�1�>O��C�)�x��a�W�	�	��
��NB��	�'���p���e,���T�L��M١�:}B�(�O�iR�F:+-��K��-9`�|�	q̓��U���T�o`�@�(÷k��ȓoδ�v�F|c*@�n�r ���?�ӓ@���[PfN86Rt�� �/$��}��ɭ�?馕����I.Ŕ�hD>�T���(-D��#��S��x!b΅3�F�і/+������}J~JE@�.+�Fm{��q�V1���R�<�0H��g���B�듽[ZR��'�FR�<i�#�?���5�7z�P���s�<1`�%JH��'���Iʖ.Qy�<9c�3}�\y�A+Q+G�f�PE�]����?���FE��Ă�a�)e�a(��Q�<�u#A����U��N0��;h@d�<�Ã	!=���A�g��-OTm�2kMd�<a�C�kE���¯ �`S�b�<y���8���sǮ~��%s�O�^�<��N١,�*!�_��X���PZ�<����}
B�+��6E�⬸�U�<���2@o����:W�VDVE!� J��źqoƨ5��@� �G�!+!��
�2���ŉ�����=1.!�dK�2z䱵��4��"	� 0'!�D�TӞ��D���C$BY(��!�č�u�L��䅮	�Ex7�:1�!��˫!Ɛ��#�6]Vj��L�	r!��DU]ph���>A�*�7!���6}�PI/�
7�5�R�Z�(!�$��E�x�f���g"l�P� $>$!�D��M��;S�юg�9�ӂ�>�!�4oBX�����l�Dx3�؂~?!���,ԃ5W�}�a���N10!�DP�g&��s��G/0
���b��x!�2GԆ`�w� �$z�����b!򄕊#������ ��XIүD(!��F��� ��R���	5�!���T|Q��P�*�jE*��W�!�D��l4aC��[�/���hB��!�!򄀑I�&�ؗ��V (�D�U0X�!�Ğ�3�b	��JI:(C4x䅘�N�!�d�+V�IS�F�\@:m�FC�L�!���(wp�j�N��E�a�qe���!�$6zĶ�k���~
p���"�!�䟃Um ��J�XGT�����I:!��+��ŋg-�=IFj$�`��/�!�@*����O��>Ľ��I��!�F0cUĵ�E��(OZ��:���/�!��)Q&1�զ
ih� �`��By!�DA�Xb�Å�id@xi�`gk!�$��vt��4H��0`V��"[�}�!�DU�z4:�ŏ��;��TC����^D!�F�W6�8��C�e I£]qE!��6x6ܐ&�V	!���hA!�P��޽Q�P	v&��R@��l=!��j����� X�l��4�C��Q#!��lkL�)��	Ґ�YԀ�?�!��K� �攚B��n�"YԢG!�%&^�	��ҳp��e)�$R!�� �)���]�Zy�]Y��Ɍ�M�c"O�Q:�(��t�����{�tuS�"Oh8���%q!�@#do�"_x
*"O(Y���X�7�`��ܗ-x=zS"O���B���2���H��v�']��'��'P��'�r�'��'SN�P2H�PTp@ �9E����'���'�'W��'"�'���'��l�`&Q2h@tYP��� ������'Y2�'���'���'�b�'r�'W��G��b��P!3��3&f�=��'��'�2�'��'�R�'l"�'���y�N�T���[ a )�|��'G��'���'�"�'���'�'IE�iU�U�0���윅=�����'���'��'���'��'"�'�Esi�qFȐ[2��+-֌�q�'�B�'���'0��'�R�''��'������{�F0x&KT@�`a�'72�'�R�'1"�'�B�'���'�`aQ⡌�d���j�$.:��p:�'-��'NB�'�2�'kB�'0��'��ʀN�7�,`�0�ȁ=Z�`��'���'�2�'U��'12�'�B�'R�|�`	۔H�@�C�P/�vIc��'wB�'o��'���'"�'r��'��hk7F��P����S�V}d��#�'|R�'
��'���'�r�'w��'r �F��e�Z1��T�t�j����'r�'d��'�b�'t*t�P�D�O����-/�����F�J@E��Ny��'8�)�3?q��i��`&�6����N�<,y�����N٦Q�?��<��Q�@Q�����$2�-\�y4����?b�>�M��Of�S��O?Q�cC�zD�#F�͈6t�!{�� �ȟ$�'X�>y����MY���(?rDh:�A��M�1��q̓��O�6=�` ۤnH�#f��S��%f����O��j�P֧�O�$�z��i��"!���a��ɇ�
`ĂG���|�x��A,z�=ͧ�?y�C65�.p�T$\&O��I#aL�<Y+O>�O~lnڷv�0c�P�Rm E�� pBU�+��쒢�LU�]�	ϟ �	�<��O.E�@�,C��-;q�K�z@� 򵛟��ɼD�� �K5��<E�K��|�V�K
|.z�qA��:e�����wyrW���)��<�쁽:�Q凃#k`��)�N�<!�i�ey�O9oZH��|'aD. t� �֏\4X�p�IW��<���?)�M��|X�4��$u>���'���9NS��tCRj7JY�"��:��|�,O䓟��J!���Hk֐pi��5S|dr��0ݴ!&\H�<Q�����z�<����L�:�f%����7f��?����y��$�'0"hY�t͒,K0��*�j@��Y-9V]Hs(�2��dÿ�bͱ���O�aL��Y���!nFJd{�k�6�<p�,L꟤�'�	j���M;b��<�qs�¬�O��Aad�[�<ɓ�i�O�9O����OB�$��m��4�&�X�5=&�t*LU3�1{�f�&�	�~�NI�I���i�?!��צ���ư�;�lM�ޕa��!��Ȋ5O��Ľ<	+O?�K��oÜ(�5�/%<l����4�I:�M�u��i~R�w�ГO���-ʊ*�]�!"[�����	m���'���';�RΛ63Ol��)�OT�C��,1&1h�]q��yc/ ��?YC2}r�>?ͧ���Oٸ�L�|2&%��iM9d��P
G?OOBXoZ0O�b�ЕO7�Hs+\�Gix��d�C�T���O���'[r�'��$&�i�Or-7(U;M,���iW��&���g�O�0z 
�����i��'�&�,�0*�:m�̀��]�p�&����Οh�IDy�Oy�ɗ�M��18/2����4q��V��2P��+O�kӠ㟨��O tl�31�z��ٴJ@��!8��� ۴�?��o��M�'(��A�g�&1����Öߖ��6)кێ���B*[��<1��?y���?���?	)�ȉaE
 V���#�� @zj�ȦA�6�qy��'��O=��|��@��u!��?�L%�%A�1��m��M�O>ͧ���Qe0�4�y"c(��u�P��9n���+�ybʟ	�����1��'��i>�	9��ܓ �[&;�>]#%�J�b�D��	��	���'��6m�!����O��DCA���K'	�Rg p�T�Cg0���O��o��MH>�B��>�4� �7��@�X�<���*�H��#T��'_�4�Ɵ#��'O�P�ɞ3�l��Å\�<�B�'���'�r�'}�>%�I:�t��pWw#0�R�柗?Hn��I��M��U��?��;���4�N���&®z��p	� V沙��1O��nڟ�M{�b���ߴ�y"�'�]#��?A�@�.����'�B�w��-+�%4�'��i>���şx�	۟�����ɉ�$��DEhp��[�vM�'2�7�� {�*���O��D,�9OJ�G/� rL����I�"�L��O�|}B�|��mZC�i>M��̟4C֎�ga���7Ɔ�R�R<ч�S!x)�yfe/?)�o@'X�J�$̞����D��`N�A�ĥ�V=b9�2�Vmz��?1���?�'��DӦ�Y�M��TB��0�����Ž09��ڰ�Jɟ$p۴��'���+b�� c�ZTn��$���?NS$t!U*ӓ|~A1h�Ԧ�̓#�Re�3��o/����y���u�C��� R|�J�s
2XS��+��i��2O��$�O����O<�$�O\�?eir�5	��	�DL	D�c��֟P�����4u�x5ϧ�?� �ip�'����A�2d��1�!�\�����l.�d�ƦA�޴�:�C��M��'�2N�*(+���\�����ļV� �.��h��|�^����쟼�	��\X�$�:���
 ���78Պ�Lȟ��	eyn~�@
���O"�D�Oz˧p�x|�j�4_��i���z%� �'���
&�`t�<�&���?Up1�Pav����ɓt� p�e-����SC
4�<�'U�BOΟ���|��� ������)�ҩ�g�\(W���' B�'���$^����4(���Qc ,KN�;rcY�F�`���d���?��j8���d�M}Ii�V��"���|�ʔ2�ĤM ��Q�'����4%=��۴�y��'��'��?	�R�T;�Ο;k�$�B�$b��s��m���'��'�b�'���'���:wO�-������n�� �Z]��bݴ��1I���?A����<٢��yGE@�T��C�L��U0�I! �g���i:�7�X~�i>�S�?#�+Gɦ��Xތd��*OR��c�����k�%A���O��#K>Q*O����O�0D _+��+jG?{�J]
-�O��D�O�Ĳ<���i�X� E�'�R�'�"���b�Y��;�#�(���a��DV}� l��=l��ē�B�Zw&�݌5�G�U�'�HQϓ�?q��]��X�P�W���$�L�{�R���B�-�*�*$%z���*�R�D�O����O��d$ڧ�?Y�ș�jȌ�$?+u&T��nJ��?id�i1u�W�'B�p��杲<zt�BdH����1�#ȏI&��;�M��iQ�7BM%&7mu���	�r!�����Oct�"�ҫ{�I�G�;jIV��K@�I{y�'�B�'���'7rl���1L�X`���V��Ux���[8?��ß�'?���e]��R�L�t=4q'�2Y��*�Ob�o��M�x�O���O�찠WJs?�`˱aS-C�Ч�B�"����_y��X�} d�	�{>�'�	:$F�Q̷ �,9 ���U��@�'�b�'�O@��M����?�F`(Gv��Q�{���a#�¥�?�0�i:�O1�'v7����];شeĘ)v��.�x8t�>�v�2E'
�M��'���(X����ۊ�'<���w��!�'ń��Ǎ�� ��5K�'���'���'���'��h���:8�� B'��S)�As�c�O���O��lZ�#x�ßx;ܴ�?�(O��F ��Tpb�
R�`s-�H�Ɂ�MA�iO�$iK��v=O&��AbhL��%����$ ɕŵ�?���9�D�<q���?���?A�@��_�B�*Ы��k�h УE+�?)������ߦ�:�c�ay��'
��Os�e�w�٭@��X���J����O6��'6m^���kN<�'�"�	�i�mwn���F���B���"0��#^�,x+O�	ñ�?���%�d�2g��}��_���|���3l����O����O���i�<9��i����,ש����_�m��!��B��,���'��7��O\�OJ��'6�ƤD�>Z*p��n��}���$B6��Ŧ�r�f�)��?�b��/2��Ц�������A���.��Ġ$�����<A��?���?���?�(��QCrFA�B���O�}��)�f���z��ȟ��I�D��B��'^�7=��icVDUV��`"U{~��zЮJ��)��4>[�����O2�4ˍ����?Oj�E��6�i�&@~U�E�F4O�0�#���?)W�0�D�<1��?����r�]ء X�_w$ј2&��?����?�����즭ֈP`yB�'	N�pc��9��<R�)�{o��)��'W�'��ʓ�?IڴH��'���p�nȸT:f���Į|�$]@�'��g�7*�:�z�J����	�?i� �'2��ɜ�z�ғ��q�����N#w2��矴������R�Or���S������.����Ε7~32�q��]H�e�<��i�O�8v�M�LG@�i�ꛏ��䦝��4Ta�恖7|������
SU0�T/ݭr�D�kDKڟpr�����bR��'�̕'���'F��'���'��`�ƛ=H�Fy�P�$E��T�V^�ߴr��-r-O��$3���Oj��PF��WH�/5�2� �얉m�����sӌ�&�b>�KrG�o�̘�j� W�2�`W�2�d��yy��]U�D�	�;��'W剣"��O�33�8H0��9�ܖ'�r�'��O��ɘ�M�5,���?�,� 2|<"u�ɦ5^ev�_��?�ճi��OPȔ']B�iw�7͙b�4�a��Y41T��1+͛f��d")o���7o�U�&����aL~b�;"2��0c�&����aB�w����?���?����?�����O����o�%eD@a4mZA{�qa��'���'�"7m��MT�}-�v�|"-�7p�`�sQ�B�J��OY�l�4Ox�l� �M+���d��4�y��'�2=y�W�t�:EB��I.�!룅��x��	"t��'��I����؟���<ddk��vI�%���c�&,�I��l�'z7m�������O��D䟔�)�NO�5	��R� ���J�$��	�����ON7-�S���I��wf������R�z�ȱc4Gzɹw��=.��,���<���<���8��5l,����$~I�"ʗK��p���?���?y�Ş����ݦAI��}v8%z� �į�Q�����,��4��'��0���*��cC�ǂ7��iQ$!+4f6����H�m�'���k�N��?Q$U�� �%�a♧C�B��U��81�9�5O���?y���?���?I����I1��x�T�֯a�-�3�I5_1<�lډK�H���� �Is��iڛ�w�r@�T�G�X誥��dC/g"��D=�Vig��Y'���?���t��mZ�<ɐ��i�6pB�A;��-H�<��o@�;���)����D�OB�$"D�
Dhd�b�@"��/޺���O��$�O^˓4S��τ& R��'�B��x�̕�$���*�~���[*h��O@]�'5�7M�����I<	�jџ^���ҡO"�$*��<��Π,�d��
�3!��m*����)�Rڜ!��M B'�!Z�.@!n�pS�.�Xa��'���'���ܟ�ぉ�.S�mx�Eב]i̭v"���#��(v�������4���ygAT��`�Y�����q�4�'��6M���=�ݴ��u��4�y��'�x����?͚�Ɉ�i�r�Z&iJ�@�z1��)קy��'��	��|�	�h�I���ɽV�*i��+C	%t�!�T2^���'q6-#)�����O��D$�9O4�J�G��v5J��3��ɗ�Pl}�q�Nq�	Q�)�S:?\&H
�(S�V8�hC��[	X+ ����U�`���'!`���ٟ$B��|�W��Y��	1�ۣ헆Y�(���ϔӟX������I֟��yy�&~��Y�u
�O�1D
�	$A;@M�,X���O��oZe��-�����Mk7�'A����B��i`
Sl^~�J�+�:��Y&�i=�ɮD��@��OX�'?���'.��b"�O�S�d��1	�Nh���	��x�I۟���� ���i�0�KSf��	�p��@@	��?y��?2�i@�%��ObOmӎ�O���"�0+�J �r��|�%�T�MO≇�M����o��M3�O���&�9;�ȥ5���9��v,�R�*���WC:�O,��?	���?��z��}���M�ȱ�d�����y���?	-O�nڻ*�<�	�h�	H�����	�����O�,�!�E�X"��X\}BNx�t�mZ����|��'18�)�O�.��q	���%,��iۂ���C��܊�I[��d�B���bM��OȠ��_�o��a�d܈�L�+$��O����O����O1�����e���p ��%+�<��Ȭx�4\�P�'���n��㟀��OT`l�%��q�$ɚx�8�r"e�5M��J���M+�늘�MS�O�UB�D����<�ѕ����OP�`��@�`��<�)O���O���O�D�OV�'.M��AMP0U����![m�)C�i�@�'v��'X�Ow�Bl��n�R�&�%�ǜmzD:�gC�S�v$m��?�K<�|�Ɵ��M[�'7,���� ��[sG[ot]a�'��pRmA����֓|r]���Iş��� � �:E[�aW1��(��Q�I֟���џ̗'6M (�����O���֣}��3��Q����G$`�x����O�o��M��x�-Ԉ��㯘�^z��]���$_13���{���;�������̖��`2� t���@�ڤ��,��B���D�O����O��$6�'�?��DFAb\��!��T̀��4��?�ƵiW����'���hӬ��<DԌ5�-� Tę �'7��I��M�2�i.6�ϜD&.6�:?I1  j�����6�	��<Č#��G,�2J>1*O����OT�D�O<�d�O�)��EG����Sѭ�3S���b4J�<��iE
��4�'�b�'R�O����qC½xR��5Qj�!	��43�:X��B��1&���?��Ӡ J��[#��=A� �h �.%���%��5�ؖ''������ԟ�cp�|�_�t	v���X�������C�Ɵ��I͟ ��͟�RyB�n�,$�3��O��h�Έ�R<��`� �6#�2�X%��O��o�y�%��I"�M�V�ibt6-6$�r� �XhJ�c�DKD�W�Ӏ�	͟� *��nG�'�Qy�O*���"�ܜQ됪+f:hB����yb�'�B�'/��'�r��;+˖Y!�C�e06)be��W
��OL���Y�Tnc>%�I��M{N>��#�cs�A�4䓊*l<�7#�]>�'u�6-�ͦ��Ә'���o��<���[=BD���
6(f!�E�<C lmb�T*q�d�������O��$�ON��E3 3b¡��s�jy�7Vg�:���O\�r�V�u��'��[>e ��ɐ ��p�s@�z���� ?2W��ڴL��vD(�4���M7��������y���*�ΕAe�41"�-�li��<��'f�B�d^<��`d�Pn�
J"�&�X�~
�����?����?��Ş��$�ȦY�U�Pa��Kd�U  ������1^
�	��Hzڴ��'��gg�6��NY�T�F�^+x{�)�s )��6m�ئ5^æ�͓�?�2�׷+�D�����K#|��0'J`�����L6�<Y���?q���?��?�*��tC4�q��QF�J��j��t��禕�ן@�I�0%?E����M�;�^푵�=~&V���5���!�i�>6_I�i>���?���]ަ�Γ$��);�#�6�H@�'��/H^�`Γ>"Yk�m�Ot��N>q*O����O�EpW�	i�R�S�M�:PA���O�d�O����<���i�j���'���'�Ι;%(�Vx���$���/$�@�\Gy��'�f�;��\�n1bĈ�#&Rp�Ĩ�'}9�D�O�`b$�5"�p"�´<��'Ӗ�D
�?)&c�+��$�JC�yB�7�ı�?q���?Q��?����Od��#k�!X��@A,� k?��`��OtoZ�F�M������ߴ���yw)�:�$���H�	��5��U��~r�i��6͘��0����?�䮄����]�? �u4L׺qYB����J�\x�0���<9���?����?���?��Ö�	�x�B��6L��B�(����$�զ��+��(����D%?-��*S"h����o}�4G�YB��H�O�loZ��MC�x�O~���O�jM�t�]�cgx¦��1���ÄZz5{7ʚIy"�u3`��I/kf�'0�	�#l�X�T+@/y� ��Wb�����ៜ�	ܟ��i>e�'$(�D�$qvr��9�d�ɂ�h�Xԑ原���w�&㟐�-OP���o�t��yG��&3Qz�P���[�1��/Pɦ��?��a�#�H�IY5�������3𾘚�Ȇd\���p��^���O�D�O����O*��+��*��y7�ޣT���@Ł�+hA-OJ�d�Ŧ=P��h>����M�J>yC��=;
n<��\�O� 9)Ìт5��'7���1_c�tn�<)��3�*�K��Կ	N�AG�K@����$�P�$�����$�O���O���E�5��Z�nW�l\�3ǜk�t���O^�Yp��
�Ot��'�"^>���ۛn�\`p���/Y��wc7?9X���	Ѧ��N>�S�?EY��U;k\\�v��&O�p��o֐U!X����h|h�'K���X՟�|��XHHE@ 	TCm�`� �����'}2�'r���O*���M{gd�ڄa��}8(��%J�S��\Y���?As�i��O���'�7��,	��F
�vZ���d�H�D���n3�M�$�W�M;�O�sV���rd��<q��<�
����8%�
�b���<�+O��$�O����O����O�ʧP���+'�H=�
Q�&*$�l���i��!���'�B�'���yr�z���,*�@�ň�$��'���S-��n�8�MsҒx���IZ�ZJ��3O�ŘV(�+�\,k��Ӊ?��K2O��!OƳ�?1��8��<1���?�7���l�k�c��B�;B�����?����?y(O�n�y�8�'���#^N.)�f�
)�X,�Ƃ� ��Ofm�'�(7͆�{I<�%cA7z8�RDk�P0�aZ@�p~҈־x�����i��Od����i�"GT�iqsb�L!ʶL���>d3��'W��'��s�=xb�� ���#@BֽwM���2e����ڴL��̢/O m�|�Ӽ��-$� t��Æ%?28k`��<AV�i�v6͎Ħ�j�����5�'q$x6A@�?A��)�V��ɡ}oh�C��&dT�N>�+O���O��$�OR�D�O��G�8OǌT"R͇�T�`Ѣ�<�p�iP�I��'IB�'C�OH2kC��n�B���*��TC��:,(����k��'����?-���kW�Ał��P�H�5 �	���Pr`�<)Z��A���O��M>Y+O�(s�R�/%伱�C�"k�\jo�O���O���O��<���'IL���r�|��D�oM�ip��9ɨ�+�"՛��d�v}ҊvӦ)oZ8�M����9ɚ���lK�	��sg!��\pɈ�4�y��'�,$�f!U�?M7W�����ߍ@�ۆw)��i���	R3|̹��f�h�I՟@��ןT��͟<�Җ�E=p/60*�C�e�Zy���?1���?���i���ʘO���s�>�O8X�K�md4鱤�]�]	Z0z�CE≃�M��i_�����0O�����k��yzB'F�
 �`�>T���@�&�&�?Y  "�D�<����?���?с���@8lp���xh3��+�?����$G��0�n���	����O�,�"���	Iȱ{��Ͽ~��܉�O��'��6�Ħi�I<�'�:P�O�M�:,�%	��$p��NA5��
���*W^���*Ol�ɜ�?I��#�E�n�܊����5�\Q�g'�����O��O��4����O�>+��N�5lT��B�'�N4\laB��E�4X�f�'v��eӈ�O�K}ic�X���Vs�@�DI��=K�tc��ZѦ���Wr��=Z��O(��%��4������J�a�8�2�$��~�^,)��m���'c��'a��'�bT��Sq� #&�;I�YA��'<�d�۴n�B P��?���䧨?	p��yÕ�q��H;7I�R��1ig�I�%PX7�ڟ�%�b>�3�*Цi͓U������]�j�˰�;R����l�Lq3�M�O��kO>-O��$�O�}��(C$Rd>͈4�޽�)$��Ov�$�O��d�<y3�i�&A�F�'���'�*�c!,P�12��ъ�3~��2�|B�'�z˓�?ߴ�?�,O�j�-�c�R5Ba���m�ȓ����j�� e�����)�S�d�"��؟��G��6-�%jd��X�p���ӟ<�	�4��ş�$?a��ş��	�yY�t�����铤�B�������M+�kZ�?9�g�&�'D�i>��8���k$酘�BЈ�'�Kޒ�����ش�?Q���3�MK�'b�#�(a� ,��\a#P�K��� �S-
XV�|_��Sޟ��������+ "
0|~\ t��3;C�	a �zy"�x�|�B �O����O����dR�P]�I�c��38�p��+̖Gv��'ݖ7�����J<�|R#�ɔ=I��R��:��q�œMǄ���$ʫ���Mv	k��'�V�Op�l=��3Q��7N��W���
��mA��?����?���|�+O����OZ��� \�r�"�aG�(�����
r�DE���?�%[���ަ�ܴ��(j�dx�T�1��T�����&�MK�OB%�������#6�	�� e(�c�*n�	��aU/V��@B?O����Oh���O���O��?�1�i^V%D��vą��eS1~����ON��D���:��o>Q�	�MsI>!�d��"xԈ��'>lj�]J��H�'�6-���S�-x�}lZz~�b��� Z�x���8MEn<c!��`52q���A�?!T�.�ġ<����?9���?9$J(n���u
F�?|��0�.ʖ�?����D��|� *�O^�d�O�˧8�h�1�ս j�͹��.����'���<���~�H &����?5�6Q�t���9���P�Nٚw�Rn�����c��D�'���Lԟh:�|�$�BҦsf��..��"OD��'��'4��$V�`�4��1�,@	�`X��KM� e��!�&T��?����F���o}BDm��aё��"�ךMX�(��P3>lmZ��MK@LX��M�O��b�˓�J��<	6��H"��S�Aw4�vR�<�/O��O���O&��O��'K�X��NK(𒀡#�3.	:ƴi�l %�'���'��lz�{��>�$�!A݃ �J�P��M�M۳�iI�P�b>9�a'B���/�0Je�F3y�,�J
l���V�D0�`�O��H>�.O�	�O��y#jS�CM��(F-؅1x�8��L�O�d�O��Ĩ<�v�i;D��'G"�'��};�lF-d�Tt���м!8!��d}�Df�Ȭl�ğ��'�����a^l᱕
N�xpy[�O��rsk��?��:��V��?��OD�d+S�?�B(3g�%U(n�Bj�O��O:���Ob�}2��O�"��b�	N��E����z�nh��)�6��' �7�:�i��" �D�\��M�R�A
�Eb��Rܴ���'^T�hq�i��ɗD����O�a2�cX�V&�(DG;jEaG#_f�I_y�O��'oR�'�R�lb$��=�ji�
�DA�'�M÷� ��?���?i��DE�#\��b1v!�d�	=˺��?�ݴ�?Q�O���O��G.A�p����H��u	⛦B^=3�J�����7F�d�J�.	ҒOlʓ{��p����#N�X%��-3f��L!��?I���?���|b.OrqnZ�/���Ʌ8����,}{ l�c�r�6X�I��M��J�>�շi��7-�ODĢ$�5
p\0M���֨,
�p��hn�6�՟4�d Y��B!?A����S�I��V��9�h�8��P�5��<a��?q���?����?���4l�9C����懎H/�	2�dվI���'qrgp�Z,�%9�Z��̦�%�T��d��5xd!�O�
}v��ڣi��\�'��7��ަ��	�j��qo��<q�H��H �j������L�'E�C�����<����4����O��dL�
/��*���)Zbx�S��f4��d�O�ʓp����!b�'�[>I��K�!�(h�͊�!�j�[�c/?�$X�lJ�495�&�'����W����ӥt)�y"\�q�uJ��
Y ����������c�	�%�l�0�،:|��"C�0t�~l��ޟ�������)��~y��m�VtСAQ9{�����7-gV��hȠ=�D�O�Mo�N�<��Ɉ�M;1�;~	0A��^7���t!؆#��6�'��@G�iV����"}�$�On�7p����X0<Pu͜sT����d�O|���O��D�O����|b2U���q�Â-Rh�2��B*Q��e�0l2�'"�)S���x����w�բ�)�KU� ���4B��F�'��)�W��lZ�<9�KL�?��s�薶D�P�27,��<���07�b�$֮�䓶�4���$��)�8��+�.(Z�BpED%�X�d�OX��Oʓ7L���̛���' r��0�lL�w��6�����n�f��O���'d6����e�N<�g�ZIߊdا	��[!zxg��t~2O(2ZZr�\2a��O{P)��5a���L+~�:�Q��2�$yqO�^B��'��'���Ɵ����h@-s	��ɾl���dKئ��IN�4����MÊ�w�T�U�2v���"�R���XB�'�v7��ئi��4�.�3�4�����np]��'�0i��TX�F��vO· ���ӥ-;��<���?Q���?��?���X
la�B�r������U ��@��|�Işh%?q�I<o�L�����?M�!��c��Sp����O��m�?)M<�|w��m���"�.ZB�9��(:ucF���H���Z�$��a�$餒O�˓[
�"�EM��[c��3e����?���?��|+O �m�0VǄ4��%S�<���(G�txS���][v�I(�M;��#�>�i�r��t�|Y��yV$㗃�iu�\�qC�'�|6� ?�sM֍SS>��߅��ݿ�'D�nȜ8��DJ&<��e��<���?	���?Q��?������5MT�{� ѭ�d��c����'��cӚ��1���D��M%��zOJ�X!�a d�A�!��&@��ēBA�Vh�O��fH�hƑ��z�GJ7Lu�% 4`өW�HI`F���<��'6�'��'��'Hr�'X�����>�&LK�G�q�ѣ�'��^�4Y�41�\T����?i����@	J$����9���`��Zv�ɤ����Ӧ�1�4Mo���)�=`�"	�2l�xY`@�o��y����VHH���@�d�<ͧ/f�$��|m8Ě�M&X�BD���P�4�`a��?!���?��Ş���˦51&����F}��;{m���QlEY� ��ן��ߴ��'��˓�M{fL�v�f��J�7UMl�Ƅ��Wd����ЅDlӔ��㟄����T��a�fy���W!��V+��m`RfiS,�y2R��	�Ißt��ʟ��O��H�)Ί)ud��Cу_s.�$x���2#��Oj���O��?�����+�]'V*�����3k�|<z�͘rK���`�n�%���?���b�Ao��<� ��q�� *�ʌ)DLOA�0�â>O��)ϙ�?ٔ(;�d�<����?�G���2D*�M-�20���?A���?����CӦ��p��Ey�'�� ��2?���0�2���;����w}҈{ӂ�mZ��ē�F�)��Ҋ)��=���n�q͓�?9�f9��A�&Z���������dM�d�%C�M��(��W`J����A�����Oj���O8�D-�'�?!d�Q�o,J�kC�I	Ck0۠L�#�?q�i�� QX�lH޴���ywFϋqTƴc �
#ĨHZ��G��yB�l�zEm��M㥭�6�M��'���"�t����q�$��$DZ�\�ȀcW����Y�D�|rP�T�	۟`�Iʟx�����2W�x���=f�	�,��n˓���	g�R�'���D�'�X���m�0S�E���*h$���Sg�>iA�i�7��P�i>��S�?�uJ��RV��bㄹg�E²C�=@")eF�Hyb	ˈ�=��b�'���5E36Q��F�7��mS,��:X���Iӟ��I��4�i>��'�P7�ï
u��DZ;~�rK4�W�9��Y��7"5�DE���?�e\����4dݛ��}�$Dk&��%�l@'
�?��e����iA�7m~���ɭ,��1��O�y�'��t�w�\Z#��
Q�y13(��l}��'s��'���'9b�'.�t!`"�Vfx�`cj�'R��e��O+x�n�$E���A��ny2�g�^�O���b!@�ex��x�OT�Ol��[���J≸�M[���:P��MS�O���fa�H���I��џq�p��%�;f�����3鈓O�ʓ�?��?���H߶��6�F%a֌g �K��Tr��?�+O��n��
�4�Iݟ��	d���#mТ�Q�e�;g�`ʔ]����a}��}��n6���|���]��!"��Dma�[�A^%K0@aS]�{C��f�������A�=��OU�lތi�\�S'��~�҄�1l�O����O����O1���k�&�Z�fA�A[?O~�����_�H�%�'�v���T��Od�n�;R�S�O�@�R�#Eޮ�Z]�شq���\5^K�6���K7nUB���D�~y��O_�1�v�Lڡ1���7�y�U�X�	ğ���џ\�	ß(�O��	� ̧ L
��恄���F�y�4����O����Ov��������]=^���)F.��m�az����������M�|J~��ǀ��Mۛ'd�"$+� a�\�'��=��و�'�"iƠ�Ɵ��#�|�P����П|�C�R�/������/*�h�lɟX���t�IYy"�j�<)[F+�O����O�Ȃ�P16�C�ʞ
P�ce�,�	�����=���&J�ICfۊnzT�@�Y#�0 �'��(�TH �>]�B�����Ɵ`���'��Hb1�]3L�=h$f�..�b�'�b�'{R�'��>���{l�IE	��n�V�[�}u�l����M�G���?��j��&�4���˳ B�\Ft!#=�r4O��n��M;�0�0��4�y��'�`�1���?�Y�)�2����+]tN��Z��U$��'J�i>�	Ꞔ��ş��	7SZ��P�BW�1^U	�L�/_n�'�6�ǟD�x���O^�d(��+^Ⱥ(�ANO!:8H�k'A��T�$Ę-O���}��&?��?y�I�o�h �/�R�����U)�r�*4,R�� R0�d��O�A	H>!,O��r��ʅx�m��jM�o����K�O��d�O����O�)�<���i����E�'*���ޜL�0Uل�	�s�����'��7�8�	��Ӧi��4�?���lH�@wG_�[�i���5g�bИ�4�y��'�"D��E�?��O��I���4*��]�VmL<*���\cv�t1O��D�O,���O��$�O~�?�	��֩�ʥZ"�O2A#�HrG��ߟ��I�|�45pʔͧ�?�A�i��'��H
�F �3KԞ�%;�'a���M'�i�)ȹ6B��6O��dCuӺh��$^��-0�,�,[`t�5oO&�?)E*>�į<�'�?����?Y���)Q��(�	�,|�
|p�hƶ�?�����D���VgADy2�'��ӘvBѱF�Fw$tpv��i����	3�M��'����O�F����̰S�K�;U6�˥I3m#BU&:�r�/O���[�?��o5�d�#^��Y:����(�D\�s�ޫ(�:�d�O����O���	�<yǼi����ӧ�1btNuYĜ�Uǎh!��=R�'��7�9�I���_����T#���)�0�|��H� �MC�/-Œ�4�yB�' x�Ç�C�?�k�O�I�rB,YU��u��,x^�|��5O�˓�?q��?I��?�������<�D��.T���:�fP*dX��nZ�'�ҍ�'�����'L7=�$5Q��j��R1@�/h�x��NӦ�ߴ�?�-O�)�b�$��F.�7���Ó䁜?b2��u�	�/�R�C`Jz���Cå^�R)E|��dy�O����6��-�&��� l�4]��'�"�'��I��M����$�Ov�ڒ�)qjD����١PY�5hV,7�I���O�7�O�ʓ^��1:��S�D�E�2�
�K<��̓�?	f�.1�:�#I~B�O{d��	�2��J�V0;C��!�DL@�5;��',��'r��sމ��ڸwj�$��n��Z�Cb����jݴp�\�j��?�s�i��O�\��ipԑ3��� sa_��Dm�lm�ڟ���j�禹��?a�C��l^�	ԿC�B䨧��b@��D�#E �2L>�,O�I�OX��O���O�I�$|�ޡq�m< ��tˀc���D[禁Y���Ɵ��	��(&?��	�)�� �B�V�}0��% Y-d��O��oZ�M��\�O��d�'��C� ���V ��g�h��%L�<�\�aMb�ɗ'n�����'�(@&���'����E�b��� �U�Pxh0�'���')2���T[��Y޴%�0�p�r�1�+atU�V)E�(��9����]@}B�f�Ԁ�������W"�@7�Ǉ#.-��
^-MeBIo��<I��v0N�C�g���);+O�����(��NH)�����d�0h�=O���O��$�Od���O��?I03��s7����i7�H�'.�ş|��ɟ�h�4i1B!�'�?�E�i+�'��U���B_^I�2Ȅ-x���/?�d ɦI@�4�Zuɘ��M[�'�o_�-�b�HPa^�n�^h��Iķ{?z)���ϟ��6�|�Z�����`�I矔xRn�5� 䋗,�ujҙ�����D�Iwy"�z�L2���O��d�O��'3���S�oх�$ R#�_�7md��'���'o�f��O�O�	�t��1�
�kؘ�3)�106H�5��XVH��*_�d��˓��q��O��L>�b�Q</�- G*���4�C��3�?����?���?�|�+OnZOkd�`�_��ၤ?N�Ԣbb�ɟ��ɺ�M�B�>��ip���gϘ�U[�W�ޞQA����i��o���m�l~���/UE�5���Q�� P�
�0u�U\��ǉS�v	��Ky"�'l��'c��'/�S>A�H�.}�<���U+t��Q�[�ME	F���O���X���˦�]�5�z%�­��W�,����πvd�A۴P���5����0h7md���2��S��EP���l,"����d�L8i^R#h��Cy�')$��V�L:3U/%hQ��D�	`��'c��'��	>�M�&��?Q��?�����/��$����7_�X��߼��'^��o���q�l�&���J�Kȴ�w,���I�Ш<?Q���x<2�R!�=��v8*����?	GC�s,�2��
12��Ġ�(�8�?9���?!���?	����O��Pw�0���V`ؘ ܘ�-�O@�m�v� ��۟�!ٴ���y�ʞT�����u�
}pp`���yb�iӲ�n3�M��*��M��O�:� ����
+�l��%^9�����w�O��?���?a���?���o��	Y!i	�a�>(hSH	N:v��/O.�nZ�'WJ|������	q���,aFƓ�y͠��6&�5��(to����O�6́a����	��ԧ��u퉦pH5�"C\�|1�AH��$�}�ՠ��-mn�O�˓F_8��'-��Ū�H&oef����?I���?9��|R-O�<oZVp�$��%9A�X��O��*��g,Ѕ�ZT�	��'�X�Igy��.}�	ܦq9��L�A609Ѕ��|�����̗�?��oZ�<��w���*"��%�r`2*O��)��\%�G\���P�f�-<y�9O��d�O��D�O��D�O\�?W[2K����#�v<�E1�+_�L]��'1��w�>�Ї)�<)e�ih�Y�l�Ì�~�Z{ ��F� AY���&��c���JeӲ���r��6-u����'>D�9iD�8���è,/֬�2��R�b�AX��Ey�'���'C�ݦN��m�P� �R��I�b �A��'V剔�M�E'�?���?q(�h8�rc�,f��yCJ��lq�="��H(+O���O`�O���O/�5jd�к1vӤ�> D�=C�A\�F����,\�E"�I�?�
`�'��%�x���㺉 e�U�ѭ�2���'��'"��$V�(ߴ�t!��
TWaVaz�
ߎsL�)� _���d�覍�?!�Z�xش
q�-�"5�L� H
>�pH� ��ܦ�B�4z�cߴ�yR�'�������?�W����OM�1W�σt�:EzeMq�@�'"�'!2�')��'���=������`q�M��MR��ٴb�zD���?����'�?	@��yg ��9�y3`�Zuܶ��e�<+��6M��P'����?M���R���o��<I�Dþ0&zP%��4	FBd(BI��<)c�[�&��E�����Ol�D��.]�Ԯ��]����Գ"����Oj���O�~����>PZ��'�bG�*�
����ͻչ�l���JN}�p�p`�Im��L�����,.\2ԵI׌Љ;���^�t�s�nĨ}w��K~���Oё��_x���@�P&��b  �)y~j9k���?����?��h��Ό�s�.i7g4B�<�:$	�������MʐlVgy��aӆ�杹9�p��T�u,�ɧ莍sͶ�	��M���iq�7�ɦ(�N6�-?��O���)�d�:P��N|,Ś��Y�x�luIL>�+O���O��d�O��D�O��y���=!��b�J4W �Qů�<�v�i�4�p�'���'���y���SB��4
�GC��C�!ݭe��ʓ�?qߴ�ɧ�'&��e�`�J�{�NG@��Hp�-4ZDX,O���C��?�a%8��<a �^�M3� 2���5ZxI�s�æ�?����?q��?ͧ��DƦ���E�P�2F?ri��퇼m�k�bΟpܴ��'��iٛf��O&6P�|S��baǴ	L�:g5~*)�g$e��z��8�D����X�K~��B��1{Uh��CY")��E�B���t��]���XU��ql̬�U��.V���k��_aR��G�VѢ���"^�fH�L�Xe��  B[�;~	;��'�e�Q@ɗ|�q�g0B��㬙�y��)�{P�C�ȼ*���x�I�ݲA��6"��j��]s�Dl��`C�R<��p"݃{9z$���۞wL>��4@�3�m�V!B90��=�gQ7lH�!ڍg
��3�ޔcdn�p�K
)�j����G�� �ɜT�<"޴�?a��?�Q�߇>ǱO��ĭ��;�KI%}��l@�F�%�l���tӌ��O����(�:�&>���˟��	.�� tis׆�=dC��bg�)b�p÷i����[~��'j�꧰?qK>y�Ƌ�:YN�"�V�H�"ٛ�o�Be�	�r����&!?��?���?)��n�2�U�9���ϮCjqB�0�?������Od�OH���O2e��V�A�Y����d/Yss��h�(�ß�p�����������Ɉ-�	��%�d�X ��A�L��wJҨ_�8p
�4����Of�Ol���O���f�'M��.��J�D{�'�w�z�Q�a["����O��O���O��ɢ|j�'B�p���:>����Ô,�qߴ�?!I>���?�P*��#��'� ���@����Eר,l�x��xӘ���O��D�O�)���|���?A�'e����6:�)��K�O�Ȱ��x�'=2��&X]��y��n�{&��7���@ L'�p]R��i���'�e
��'���'k��OH"��5IF9����`�� \���Ɉ<�M#���?1.��C����<�~r�Z�H��V)U�V�xy��ݦ�0$	��M���?�����b��Vx��1IW'.���`�+��m��n�#<����'O�s�E�*��D��Ǉ�fҥyEn�����O���=N0��'��	ݟ��Y�V��B�w�����$/����>I!̛>���?!���?QE�ބae6+��
�A�E�&�'] T��.�>y)O���9���ꀨb�B�r�E0e�G:s��rtZ���A*�h�Iٟ��I����'-�}b(�{����@G1�r��ϑ�I����OԒOt���O�Y�"�Ջ(Fb)!�3�54肯D]ܼHM>����?Q���Ğ')��x�'\�}b��-D����%`VN�YmwyB�'��'�R�'Z���@�'#�ldDCh� ; F	"n�� b��y��'K"�'#�0>�(ʨ�N��Fζ�Jt���qU�<���^n��m�֟<&�t��֟�*S*�Q�mC�A�@Fе�jy�,l���@��HyB�Bl��'�?���"�K 5r�H�AH
]��D��,@�	��'���'u�9�3�'��Ի�O �Ӯ)�p��Vf�ޔ(��{D
6��<$� ����'�B�'x����>��cS�a3���T���$O��\C��o�����*fT-�I�8X���OWzP��g@7VL�s`B�N��@��4N(|@ֶi���'�B�O ����\j���j��X��t�O�TA�D��Aq��Z�b!��y���?I�+�Eb]�v���x����כ��'��'�j�/n���ty��'��d/q�E���K5�X�MѱO�4���3�D�O��d�O�ı����o�%�!F�h� �o�٦��	�,8��+�O�ʓ�?�N>��:���x����u^��1R�Ϸc5�	�'���x��'�@�P�'���'@X���A�о^�=d�9+��A�gݨ���O���?�H>����?�A�=jb��"�DI6)��K('bH��N>��?a����$C�L�ͧ��L�&H["7��*����Bd�'���'=�'��I�5���i�A"BѼ<޸��d����C�O����O&��<YC�W�C��OD���[�l�B��`�����:r��'P�'�剑%E$P��z�INH/�iC�G
7���z@��-����'K�V�#0�ħ�?���C⤚�v�"U	*"fp�;�Sp�Ijy��H��b���ٟ����^-��9�T�B(C�Čs�i��I\v@!1ߴT���֟D����$\��!�v��v)QСj��w���[�H8u��ş�L|zO~nZ�o� UaO7� ��g�.xH6-�8,"r���O���O�	�<�O� �H�M��9@���i�	`�(#�g�6��2�ׇi�1O?=�sM�3:%n��S�\^p`���$�M��?��y���,O��l�d!|�̘�4
:������{����<g��*Y����Ĥ�Ps��m����Qy:ց3DDgӰ�D���x�/:��\�+����}(��өP(QܮP��T����+#1z�b����hy��'�PPtOE���}b���-.�|�3��E��П��	X���?	�l�|	Y��c/nQp0Ĝ�nQa�`Y:ò��<a�����OڈP�e�?�j!�^�Xʮ���,ѿ����~�P���O�����┩F@�7m�B)�]�BN��ar8r��Q&2���՟�������'�2��".��P�R9p!v��� /(�qq��
P7P�oZ��|�Iey��'�����ҕ~z�B	���(	f�Z�n�
0(�I��M�I˟\�'� �A!j!���O��ƌ�e
K	�B`x2dd�
e3��x�T��9�R�l$?��V`�a�c뾨x�(ܺbx�	n�jy��$EN�7�OD�D�O���z}Zw�6�B`��Iu�B�ƕ�j���0޴�?	��5N�y��?�-O~�>ar�*�����a �P��q �Dk�����Jئ���� �I�?��O>�JY"M��!	bxe�A�U+V��Y9#�i�p�'0�Z������ꠘ1f�cE�F@҉>���Ѹi��'�R�sQ��X��'���O�9	��a OX!^�=@S�i���'����/Ѧ�yʟl�)�O���\ -Z*����/�:aΛ<w�Hlş�ڵfU����<����$�Ok��U(��i���$���3�h�����a�H��������l��\��'CXض�C�`U���Y���𡎃m�<ꓜ�d�O���?���?Ѷ��	R��pC�d"����Ywt ��?���?A��?I+O�YB�C�|� F��0F�����h�����i����'���'��#��y҈O$�Z�`�3Fy2	A0L:7��O��O���<�	R�H���ß4j�"�tP\4*�-[)4+V���L��M����D�O����OP�Hs��x��'b򕲷MY�/U0�k�@	n&�,n����Ify��Ԅ1L��?Y���JWJ�Gjxʔ�R->R8V��rX��O0���O��dN�wt�|Γ����Y$�f���-2��!�KN��M�*O�,�v�ᦽ�	ԟ ���?� �O��Ս]ET!�$�
#�R8
�(�wW���'���%�y��|R�I�>i�`�0!ܿ{��ԘG�yH�6 ���7-�O��D�O��t}2U��{�E����єw�D!��M�׎��<�����)�Sß8@`,O�+n�x�Q����$q�͚��M��?)��`A]��V�x�'���O~5j6�%L�$\cI�p�y�T�i���'�4e���yʟ��i�O��� >2;'/i�T�q����S��mƟD���4���<�����$�Okl��.@<!h��)x�}hfDz�&��7X��s�'��	�?)��ܟ�'�jdG&܏;b�����©Ffp���B�q�����$�O��?9��?Q���
)��cG�
L�����)A ���'�b�'���'���%bL��OL��H�+{.:}J �O6��r�4����O�˓�?q���?i�#��<�G�A'Hf��t�� �4� ���'�R�']�R���7.^���)�Ok�'K�\�1�P�N��y	��J�T��v�'%�	П�����P��~���j?�e���vR|���K�ȀU����=�	ǟ0�'��;A��~"���?a�'n�ިjfm��~�v��_%$�y�R���	���	/t�
�N�	S�b��4}j5�5nϦ8BZ-0G	�Ϧ]�'�h� a�z���Oh�D��-ԧu�-��Fi�W��K#KS[B�`m�Пl�I�_[H�	��9O��>�b�cM�*�4��%��BA�&��6��0T�dn�ߟ�������S&��D�<1�F�|򺙫�IU,\ !*ubş|����Æ�y��'��~���?�%o)jd� S#R<#������ٟ<���'hr�'� .[���Xyr�'�� �5h���A �>7�ep�A�7>���|2�ݲ�yʟ����O��D�->0�iV�}�^y0���>�m�ǟ��@�ҕ����<Q����Ok��..,�!�(k��2��Gm�I�?����qyB�'�Ҙ�T+ {��a��ƞ�/;�U�Y� �g��>�)Op���<���?��R.�ꡊ	jT$$R�����������<���?���?1���$�C�r��'  �Qy���	�|9*aA@Z4^�nZuy��'�i�oZٟx��|�l�i�@'[�sA�4����4ӐCt���D�OP�D�OpʓM��A��R?��ɝl@�K���/(�j���i��,u�h�4�?a-O���O���k���O���#Ul=�VN�H"-�M������OH��<Q1@�*/L�O���O��8"���Z̙ �	_�+��!�d �$�O��6|��$+�ĩ?U�&�֫ֲ��t�	�I�a��qӦ�a1�I��i��?���"�I�:gĕ�'1�X�V*_�<n�6��O��W�e�H�D-�8�S�|Q���EgK*0y�_8"7�D�6��l�۟h�	ϟ��S/�ē�?�bH���d��$�Q�֌%�E����ƭ���y��|��)�OVp*���|Z ���B�2bv� �ۦ��I��X�Ɋ*h&�k�}��'��A�i:d۵��"T�i�*�<f��f�|2��j�\�����O��ӢRmx�) �^�89�%��g(�6��Od�����g쓩?�J>��Rg"��Y8H%, ���0ZNx�'�T)��'@�	�(��ן�'�|U S�'�쉣� ͚%��֟0�xc���	c�	ɟ��I.�t���@
�
)��Ax�:%�p�ԕ'��'�BW���"����D��(+Z\	��B�+��������D�O ��=�d�O��J3����Z�?P^��cV�c��3�VK��'���'�2V� ��*�+��'W�|�y�#0t�Ĩ1plR�R.��z��i���|��'��)��yB�>�H-.ո$[�?�~1���ؖ`#���'��W������ħ�?9�'@-�AR��4$����˄�!g�J0�x��'B!ͭ�y|�П�!��!��֍�}[��J��i��I�����ڴO���П��Ӱ��d�R����D�t���[6��F�'����Q��|B���	L�%Y��p�DP�+�oR����*$\�6��O����O���P�L2!CTA-"%&�)a� ���iV�ۂ�'��'��,�dUe!�,R��ș*�t*b�ʿI�mП����"I.�ē�?���~Re��8zzEk��R�,��x�g�(�M�M>��		�QB�O�b�'�r+��{<�h{p�5�p�+�,�	?jz6��O^	��ƻ<q�S?9��s�I&�\:FJ
Zޥ0���RV��J�O�8��Z&��	�t�I����'GPlp� �}O��3h�*(�"Q�&.�W��O`�D�O���)�	�\GB�co�#`oB���H�=�PŠ��$�I�T�I�8�I̟`�w�L⡂I���rL!^cWCA��!�'��|��'�Bk���D��4l7h��Wݱ9���1�D�	���'��'B\�@
�Ԏ�ħ[�>A�EJ1tzm@�	=D���i�"�|"�'��*��'A���v-�l~x9z�D��i�4�?��������h'>��I�?��� ���HC,�4�A�1��`��x��'�]�O��޽ ��>,�H���^��YK��y�9+�b�'?�@�+_�I�0��D�*&v�!)U*D��8��1β1y�!���ʸ�6��%�$��o˾�x�J�8Vy�;EGǙu>�	X�oM��\]���H�EX,���� w�"��A�]�甸�f�/����)XU�0ϋ`
X�Q��[��0��V�������9y�Oɧ�� ؔO�D���h�� �"�k�s���!+�8i0���O����O�Ȯ��?��_d0aS-�=��Pp�!��ZA����'�Q��+�P}����B_F{�� �tSj̱Q@��+�(�#�	���!l0�I^�Q<l���hO�t�&� �b�e��E���O��d�'���uyB� N���i\ hPQ:���9�yrM_9P�)�]�CǊ�af�)(
"=�'�?�*Od�#d�ަ)r�����<�E@*YԀ2gj�柈�	����	�=[&,��ܟ �'+6<��PcF99B}�ba�&t��y���=Z��DZ$��wF�{�r��#ǩW+W�Ș�cP�U���C*�iq�Lz��єNYma�jr���I؟�2�z밌��E�� �� ��f�g�'�џh�Q�S]��dDưo�����5O �=Y�JЋD�ɻ�䝐fJ���&a��<���i�B]���Ԧ���)�O�˧x����+8p�6�V�T��)Ȑ���?����?�u-�82qX�	�/E�p�F��򩕴����I�\bF|� OY"Q���f�X�4�(��m�lb���IlC��2��X�ip�!˗I�+s���/O:Q����O��2�Ӌ!�R�{0�L�BS�؛!	�pCJ�z��=������C+�MP�H�w��v����=�� @��aùV)��:V�����
]>�m�ڟP��R�4O�z��'��N,R�2mP�J��S�8��I
z�Nx���^�H	q#C�K}*�^c>�D
:o�0���Jʏ$�����g���(���zdI������O�< "��<l��,2`ᑨy�ΩJ�d�#��d�Oz�S�Sb�I��n���Ed.4�C�(-bB䉆i	&	���V�G�ʴ(�&�'}p,"<	S�i>m��=t� t���R)5�P�'X%j8�4�Iß�I��uˀu������I؟p�_w���'�r�3�!R�n�ȣ��ٔi ���VK$U��uG��gN��Ef[������i:�D&��aޥ�
�ʒ��5�ӿwڹH!� hh�!�ޟў��g&��kY@@sG��/
��I����X���O��D'�$�O��D�<)�� 
O�ʕB��;�lX�Үz�<q�Eݰ�B��@1�t3�,ǸH`�����⟀�'�� bf�s�0,�fE�j���:�Hc��xC$@�O����O��D�?<�D�O~擑V���������c�Κ�xF�Qie/F�$��(�tf2�O4L�`B�h�8�#��V�%Z�$�|WR� S�S�m��!M{X�����O$��V!^� ��#�@1)R�P�7�X�OD�$�Op���r�1@��/HZ�7%�8;1�����M
������|��_��IJ���O�r����K�A_Bm)�O�<(�<��'�"�ga	 ��l�t��5����'Q��c�X�Z0�uy$d�>=8��'��1��-5*вd4���H�'����HK�9(p!�Ħ�.5<1�'���JP��:R���pd�/>`��'���Z&�J〱��������'��]��ܟq8���v=�� �'��T��G�74�����l(!��'��$��I�A��sূl�,���'GT���BӪ$e0�b�Ԅa[]��' ���0���h�	XX��H�'�^� �խv��QD/	Q^����'�>�#wF�\FX����>M�z}�'� \�GAln��/��F5ڌ��'Р���Z�B[HEI���>dp�'�H�t�B����NE�1�\x��'���3U�U2\J١��,,i�
�'��hbȡBf%!S�)��h
�'@ ��#��rގIWjK/
��ٲ	�'�r`�g���<�M�uE4��'��RD�I}�(��5t���3�'2�Q
�����Qkөm� Ua�'��p�V��TA��O��I����� �4�w �>��E��·}^Y�"O^�b����>����1�z��`��"O�u ���5���0y��UH�"O��0�f��FBƍ���(��"O�u�7���RQ�M�5F؃r��y"O=y�j�0��}�5/͗ZS�1Y�"OP�� *�6w��H����O8>� �"O��Y��!mjT#���~��1�'"O�]:�"�Vxa@7�r���a%"O ����ˇHpN�b�뗽D�Ҹ "O&��,�+=�P]#���P���g"Od�Ui[�G�$�	)��Dӈq"O8����>r �I��!�1P"O�j�P&6���(��R���"�"O@�#�e�o�T�bh��v���g"O�!��璾i�4e��{����"O�t���$�P=p�J�d�l�"OiX��@��i�6���p�$�@"O����K��,a'��';�!�"O���!Ad����$�7�*�9�"OҐI�A$q�fT���t��XA "O�h�B����P0N��X��S"O|I�A,Vd���"őv��"O��1U�B��lP�S��$�(K4"O���CL��>�i�E ƅK8�!ir"O��� �	4�p���L,���"O4���J�7X:u�N�(-T]�U"O�ِ2`��lb��dҷ�j��@"O) �e�*?�݃�Y ��P"O�	ֈ��7J h�� F�u4��"O���j�8x�x��%M�aj@!W"O&pI��I�+/ź!dC�t\���"O�!0�)C�d,Ő�bL��J"O-@�D�-
��X�W��)��r�"O���A��*]�Y��ÝA� �q"O� ��F5��=�� �R��Q#�"ObU�-Pj.$s��3�H��"O���O�<u��k�z��E���O��Kg��n�S�O���ˀ
����*e*غFƶ�y�'�N�� �I�1�x@eb�09�DHH�t� ��$�p=y��ݞ��MY@آ�~��&�}��(���r{�	�c�"Z�f}�����:^�)"Or�nTxB�@�a��X+*���I3D�V����
�<4lgk�"(�
�j˵27!��]	9:
Ы�-Re1s� D)|��_�h���>E��E�k+�ƚt�۳�]5+�B�ɀ7���b١Hw~e	$����'��܊� )\O.�	֧ԝ@�� hS�i��1��'�J|Z��N�|��E#�	��M��u��чȓ>���b	?[�މ�����@��5�D�ZQ@F�(�8����H�V�!�ȓq
�y���*D�@�r2��9�� ��,�
�TDɇ�):W™&W `��V��z��9�zRr�5�v}�ȓY�bPy&��}�|�GjX�"F���'�܌����-�EB���M~�Յ�|�t8��DC��X� ��8Ԛt�ȓT���JR��1~�xr�\rW���r�t*��ȀVi����E�"�f���4?��K����9dV���!���y�ȓ,�t� �*\�褕(��g>p��D��eHN[�ɰx9f�[>	ҤK>qV�I����/Bx|��'+)D�Г�m��<8�,�-,y���?��Ɂ'ł�����K^�g�'��UaD���U��CцI:t-l��>�l�ծa�? LeC��9(�)z�FY�XҒ��5�U5l��ò�'��1�*O�p�r���wʆ�+��D6"
B�`�,WFJ�[a�?�c#NU�#�⩠P!ܟ\�2$�9D�T�t�Բz�BA�C��?q����#w���(=��݃��޸\0b����2����O�/�䰇/�a�!�$C-z����1��0`�T�%(N�k�"��w>O�,��&N7[��T���?#<y��"�K�AI!-�b�AQ��a���hC��9D5H��gF�>�d�s
�!���0�B9}nD���M'�O��y�gP�;�����/خP�D���ɝ1��,���6��%��
<��%7�ĸ��&V%]�v����g�<iC	?^�8�'�T E��"1�Y�<!a����X%�- -�����ӥS�ļ ���Bk �r@I�62C�ɉ7_���q&P�=(���"$�pT�8s�k����/J2 K�E/FxcՇfdF)P@��5�(Đ1#\��0?ّ�J0�.��Q�j��U���pi� ��G/nɊ���GK�B=0��򤗛L'��@�`�&<X�	&�Y0��2�� ��7���l�艓��1H��A�Ј�x�`e�'�@�*�O��:������j �БiXV�X�1O�A{��Ψ8=�eԋa1����i͹%���Z�#�"�pa��&J���ťG�R!�d���ƈIJ�@�ѽֱ��:OX��d�E D��x7l�X&1O �{10�z�
 
�&DL>�!c�3P���r�'�P|�SKD"�n��.
9�����������O?)�ӏy��W)_�r�Ћ�2 r)����S�
i�������� @!����B[#	���*��-��7K��@��&K��t�'�8X)�:�O2��dM
�h��JZ;�p�����i7���6�qO�#Nt�DjS�� 
P�+�Z(\^��@$C䉔"u�@�Ċ]��L�֋�,Ac�L�҃�l��lPn��O���|V�9��BS�$7��څ��M�'���؁���<��c�4��՞;�YѰiJ�6K�>*Vd��b��Y�4aSk�f(%��}
�C7E�n�ҡA��kL�"��� ��qQ�ݘ��M��h�5A���>v0ŦC,q Peb!.��b�-C&��|�\�?�KG;{�,[��P�Y��`���J��dɪ�~b��O*���N��?1l�����#9�|��seΆFR2�S�/��\Ȼԉ^�f�?ɤG	�x�~�q%�BZ�x�D��@#����ԽioV$@��R2c�`�3^�R��ɪDHp]Hb$�+��<�3"����|br��0�F4�!`\"o��Q���C�ɘ�ލ��A�G���i�x	�>	r����D�)"o5zj��\�`�
ْI���Q���>?9�)�x�䌠B'S���ܢ��Z$i�����=��Y0�K>� �"J���'ٱO*�X l�?�����~aE�)~�	�_����q�@��K�$_�Q�,Rk+=��%�
�)v�4����'�v�>�6��/�F���IiJ�q��[�8�T�_F�����I^��Q����#E���$M��� F>{�hH��.݅;<�G{"KۯMh��І�"�M{��R�]��h��U:V�`�`�j^�y�+>O�p���|9H�'����J>a1	�"����ץ"Hy��ޘ��7-�U�:T9R@<6-כ:��eاfO�J��i"%�7;�剛!�re�4 �v .)�`ـV����$GV?uAd�	�1����>9ԋ�	[�i����t�� BG�C=�ܓ���Z��I#�m�tE9����`�#���X[��@�1
ND@w�>Yf�4�0<Au�	�b���$Mի��pP���{Z��`'ܪRT�>��'U_��m���X�"=�d[�#��ؓ'xH��D�/ Ϟ�#�X�h�A��6>.u1��#S�`hI<�f
�Ǧ��jH�@؁���E��lm�c!Ԍ.b\��)�x1Gy�?Sll�g)Ĭn�\��	��JD:�o�?,�`H�`�A��U#Eр#z�����T�?c�S�M23ـ�F�h���ea�>qc��&L��D���@K��>	ǮBN瞬�㎌m�~A6mHp�	9sZ����'�.-2�l�4�"|J��)[ ͫ�����O����C�}�I�`Nռ����M�T;P�W�b��� �G�2<~�@CŐ��S>e[S!�Y�>���
?���6�7��Ip�~%eЏ,�*�%#ʇ=��|Q��/��mҀF^>Z+��rŮ��<q%�M���I>E�%V�T�H��'Ts�b�c��іE�b�I�I�H�B�2�$�<�}�È˃m� $��CQ'F������i������e��9�0<U���Z���҉?1��ɓ�ϷI �E�hA(��ˎ�|y�}� ��!\]1O���:�R�X�,�<"0]9"���4O���O�k��c�naTOL
$z�s�M�H9���a �F|�L�#�`�G�$�ԥ[���A0��_�����*[���u>����E�2����p�;�(���"'�M	�Ti�Z�v��"O� �X1��Ҁg�(I"Iʄl4����5s�,zr�<�BˀI���'���0f�-c�Q9�
�'��Y�(	�	�jɈ`ݢn�h�� ��~�A�d���Hf�,�
�O�j}� Жah
P�$��z��-��	�mC��VAXux�Y��'�x��(
U\�p�2j��tQ�'4d X�D�N.hS��;1�T��K<Ѣj�6⢨����,@k:�}:Q�)4E� ��4#B� ���P�<�t��<�.Q"b�� q�`!�UƋ��� �O��@���7����{\��UbѴ
���UM����t��y#2�A���c�G	`���Ǎbc���]&�MȖ"˻U}��d��5 9���g�-�BFޛ	G��A��3�\����0�r��
n!Z���Ԧx&-�ȓ�$x!�*_�{@��k�-E���ȓR����/�(lr���#��32��ͅ�JO��4AS%&����i:G��C�IxȀ*t	*~���G��B�	�l::���Ib�6��IW��B䉺K��ٸ�ʏ�zN��"'*�TB�	($_D�á���R!={-�%"O��) ��<�\�b
aI�=�w"OLq� �տ_\0x��K�1D��"O����<t�z��"��W1��"O�9"��H��z�Ȁ�C'|,��"O"(�k����y��g���� "ON5�Tm&d�>���$_n�@�t"O�L �DĈ����� ��j"O�y1�iJ���X���W�~�Hx#s"O�y8�û-�&ݐE!T8ը�0�"O�p#e�P"TM�&�����"O����#gl|x�'��mO��P�"O����q a˂��V <��"Or�u.�z�����"a�E&"Ov\��<h�t��McN��R"Or%��D�*}"A�l�0Wi~=c"O��
VH�$.Y0@��(`>0C�"Od�Ъ��q��k"埒FAnp��"O8]y&JKD@�]�!E���"O4K���/;� t�ך{�x�p@"ON9Z�(�%$�|���@G=s���"O�,bӅU�$@���A�%���Ї"O����
yv=h��A6����"O�X˳N!�T9�C�@=�x��c"OZ�*d
�3�tP	`M�	�r��"OR�B��L j���L^Xj��"O�����#bi��P��M�!�"O^��*
<q{�r�ɍ5V@���"Ot)�@΁�crF[���T�:\�q"O��[3 �_����'U�7f~�h1"O�xB�ia����q��~�R̋�"O4i�Ѭ�"hʔ��d���k�"O����R (������9�ڌR5"O���d$:*��K��6\N�Yx"OR��e	>W��SsH �AU�� "O�9鐎).��1�f��7V��E"O@X�/��m���0h\�_ �"O���s�L-�R�3��	���a"O:�H���#�򈉳!\�\�Ґ�"O"YA��,V��J�o��n���s"OqX�.�d��9@��m�� v"O҅RTŀ�^�&-�v,��:��w"O~3���-�=��J�f��$sS"O��hD醳PxY�A�tpm��"O�D�Sb�V�ڹ9���72�4@"O� ��p��A�la>�V��Oj�k"O�-q�mȻ(|���[��"i("O�p0ӮM4Z�Z�{v˝�+���ٱ"O6��EF�/1�pu���[�Q��4��"Od�0u��Xu��&��(h̀���"O�5��Z5;f"A�s�՜n�8Q�"O@=@S%J�8�4�0viP�w=�@"O�عW�2tF����K�o�8"O�lj�	F��l��M;�0���"O��F��$d��� Y�z����"O�%����&�&\YVE\[	��Js"OB�H֢����]3#��o�0���"OnH.w��*�c^5����"OB��"+H2q����f�A�6s��r"O��w�X�"RLx���=E�H$b "O�z�J���4����� IX5"O0��0͉e~,�&��e�FTq"O �Ȱ��:.TT�N��s���"O|�$i¯�h��'�V�=��"O���b�6���q��C�4�� "O���%N�<u��J�������G"O�B+o:��򗄙�r�Bp�P"O8��C�<����✨L��c7�#�S��yrN�,��"�_=Z���Q�fI��y���Б����Me>���N��yN@1)��"��ъQLRi��Jܑ�y��A�{��ȃ0B�Ok��bgL;�yrG�"�\cV�D�M�\Xc�FG��y�W	�ʀ�V��e	��@�y�h-_#��ig`#Q���HpgӁ�y��=B+�88נ�6��Rǉ���ydE�0`�C�2E,�`yAd��yr&C���H���!JKBy��fC��Py�~W-+kD 0���:Y��ѵ"OZ��c��a�t��.�/�(ur"O���*J������
A�] �xy�"O��Z@�� u�����n�r��CA"O�l2���)P�P�0fSd�HE"O�t��A�i% feV�fhX��y҆�:N�[f��;L�0�A5�y�	�o�-$'�74`t �΍�yrČ�c1��
3)D�h3����y��::(t2��(p�B��y�bP�S8���3�� +�\Ju)��yr���l`��B� �:u�'g�9�y"	�t����&����B�nL��y��ށM�J%���0�pb�nO��yBgB�8�b��45���%��3�yR�� ]������5d<a��L��y�*��H�2�s�^-4DX���
�y2̄!����HQ*-�vA�0m��y2����D�ų3�0�����y2%��)C(�A�.�='u5�u딭�yB�԰b���V� �P������y�c��|I�[ ��X�90����y�H�Q
ZMp#�N-�lY0A�A�yrj�	ĊUB�O]�>�2`h@��yR�Vg�R�R�G��[F<��!�6�y�!+W����A߶L.P}hv΁��y�H"hݨ�AoU�B��4��G�"<Q
�z�~ �Տ·aC�aå�%v�LQ�ȓeƦH	��3�~ �[�$X|�ȓ?�h����R��T�G�ߞj�̑��#���8%�Ӈ�����ǝ ����S�? �E��`S�g���ŮH�oe ���"O���� ,|d0�-�������"OX8��a�MnL��Q ㆌ{U"OX��SI[�T�䁛doE5K�A�2"Oz�Ф[�2�~��n�1 (i��"O����)�)l�F}��hTN�x�"O,�J ��m`�f�"���W"O�9s�Bfq�M����<��k�"Oҹ�ᗄph@��ph�2b�ܸ�D"O$ؚ�J�3q02,��˵K�Z\!%"O���L];U���\�9t�4��3�Ş	�&@�%e��$��pc ��1�h���`0�L�a�X�h��Sh���<��G����"��8h}ބQ1k��X���ȓW�y8��\�, 9��H�E`\�ȓw�8A� 5��(�" �1Q��hR9�`�Jz�0p@wn�a��H�'�ў"|�N������H��GGH:'!�d����F�աR� �c��  !�d�G���M�_zA�U��P�!�ĕ�n�JUH�E�5~��h+T� [!�d
|�X	3���h��(�Ӡ�H!��ڕ�bqQ�/�;�>����<*B!�!>�i�lؤ3�P�$T&y:!�;ubB�	�JWV��	T��hL!�$�*�ʔE�#2Q���S�Y�bE!��W�p�v��a��mH2�����9'3!�d	�x�
}`OM����3oGA�!��3�"��%Ժ4�����͍k�!���R���^u]R���N@�C�!��@.Ou��1�%0�%"E"Z��<��'�� �!��f	`����N$�uq�'�H,rs!�B����@E*��'M���Ū���dL�o\m��;�'�t��^�x�T���)Z�.�F,��'�.�Vg�=E��3qk�0��s�'�Z�	+ӗB������7�iA�'JJe	�������V2�N\��'ĨRbC5~�tT:��;V�@�(�'����"�S"��	*˘� ����'w�L@� ��+���.z�6Ĉ	�'��-yf��M�&�C�q�ҭ��'��rc�,ٹ�"R�eU@!��'��YDGۺ%���3��.ʚ���'X$,�ƒ=��8S�.�Ȉ�'ɆՓ�d��6� ��B�W�s=d���'w��"`�}P��ы߹j����'>Jh�k�h*˓�0`�,Y
�'�����H�F1�3CD-#�*�+
�'�)��J�;Z��L#bj�5!����'��`H�-�����A� e�|�
�'�~���K=sL�dS�f˔.��|�	�'u�E�l�1/-�I�P@R'y�l�	�'�.�n��91��Z�_�J��]�	�'��!��c�c��!h��
�<|��'Jў"~�� Q��|z�`	�T�̨��ld�<Y��)pkl�&��c
Ѐ�R��J��t8��QW��)	��Z�l��2�\�(�m!D�����O�6q[�+��Z�l8@�B!D�xRB͓PQu���!d(dy�<D�p�sA+H:Ry+� �W"4�k��7D�r�i��)P�8�Ċ'8l��5D��* -��7�@�&�ʞ=�h�A�4D��gdL�$�4�ۢ��6D�� ��YC��(u��	p�ײI<MJ�"OԱh�
`>�j�@ƺ��v"Oش�EC [jx���X�K�
�# "O����O(}�f��� ��D�v"O�`�p�dU���F��x�꠳�"OR�ЂBn�D����5%O���q"O��rd��~��9��閃75��s�"O$���AЂ�vc��/��r"O|��H֕+���〪j&��Pg"O��a1&�����θ�v�;�"O�K�Mɘ~:8��tG��"��l��"OF�A�K��<�b�Զ�����"O�q{3,K�ʨD2R ��t�̸�"O��PԤɂ�8YC��f�> �"Oz|9��-@2@0�''#��4��"O�ţ��1A=�=bǇ�h���"OĬB�d��O����&Y�l��"O��h�%��p�zM*]��aѧ"O��G녡8��%rc�δ]���)0"OV@P)^�5��3
̟^��Cv"O��� ��$A�ꬹ��<\��X$"O���v�L�z^r�����o���£"ON��/�D�x�*e
�/z �z�"O��p��A}�Pv	A,X ܈�"O@ș�OH��t�I!5P����"On�8B r%Cņ��Q^��R"O�����3qנt��03Z.��1"ON�I� \��ec�&wr�"O�a��k�7D��zf�Y�C*��V"O4H�f��:�mA�n� vS�m�Q"O(�ҁ ~[�09��*IA>�p�"ON4��Eo���.�
�Ș7#D���Q��78.��Ӂ�/^3�śq�&D�ЫeK�;sɲ�R2怞wVJL�T�&D�t���!>YʰX@gR-h��C.%D��t!�c��H�+�= 4�a�8D�t�5@X3!m�(�¬�~� ��!D��hs�Ut�H�� #�����J>D�����F��!� �l��x�$�<D�hS�ϖ�ȑX!�'j��ⶤ7D�\�#
�����Ō�f���`5D� b�@�����S�()��Æ5T�V�O��*T��.���!vWh�<�R�iNIj� V�2�̨)���O�<�A͜�a�4� ���P`�Qa���I�<�qė= B������\��D�Da�<��C�Z��r�n�3i ^!	3M�`�<��oG0t}�U�CД@�Hq�vi�P�<�H�M ����iQrB�l3�!TW�<���X�$�t�S�C�v�D�
��X{�<���4&��,;db����&�]v�<�B�+��t��&�5��%� �u�<)�#D;?���)I�22	�E��\�<q��
�A�܆IH�t��g�M�<��e˰L�<E��Q�2ɩ�m�M�<9A��+֖P��@�����TL�<y���)��Af�՘K�����'�K�<٤P�K{��S���U�ĀįGE�<QpJG0� C�L]��9��~�<�C��EQBԋ2W�8�°�s�<� iI`pTKp��Lh�l2�r�<)6͇���'
Tg���Iq�o�<�g�
�F��Y���9��(	A��u�<� �6^�����`ˌOi3�J�<� �Ź$�0(c�`�ˇ�5�8|YP"Oj�q¨]q���2b鐹֖�"O<�D�&ڮh�q蟣���"O�HA�ʖ��~}%�4�>��"O�P�� ��~j�g�`r��)"O�����#.H��kG�U	T�jH"Oș��`�&�.9S�b�<��P��"O�y	B-th$R�a�}9��`"O�;�@���
6Ɓ%�V��5"Oj��PM���ur�CQ�`�"Od J�+u�(��Ъb�UsT"O$\B�CI;b�e�&aO�S\U�g"O��7c�|�)�����y��%��"Oɓ0��:m��A� ��e���"O�m{�!��LPx}��Z����B�"O�v�L���3Pu�QR"OĀ��IϹ}�\�Y�$�	\;L�&"O:���[��������<Rv"O�z0�L
r�$s���.[P(�S�"Ox`��P ڑzd�K.���B"Or4����(7� 10�MD�(�q�f"O����m�1[^�����^T��"O�[�	�#*�0���[V-�d"O�=�"h��9x}����]����q"ODJ�O�?���)@m��hJ>��"O
�`�M�+}�ꭰ�,�� J�Āu"OĸҢ���(|�E�3� ->L�)�*O�3� 4�)�Pg�+)����'�&}�j��|z��K|���'��h�@����8�G̏:E�vs�']��_>M�bQz���?��5��'m:y[K��L>�E��
,3�ĭY�'C8͋��)c�ٜ)T��'����Oћf߈U��9&i����'�Nd �6an��r&ƚ9�1`	�'�l�h���P93r������'8�EZ��֭lҞk���)Q�x+
�'VR@�u_����po2P3 m�	�'��8z��?��y�A�\Tp��'��h �� QƲ4�l�<S�]0�'��c�;��[�YO	� B�'�j�;��$S��q��/�4H����'�8Aѐ���Z�F����:��0��'������)]N2y�ǀ�a<��'
dp�vH��ex��3 ʰ��Q��'�d�j�c�Bm��3�.Ԍ��'���8!�݁��X��&Y/�H��'�(��ve�8(�k&���Q�l܉�'�p�G�U���Չ�%Q����'Ϟ ���YS5H��LQIPP�r�'�
� �
�y�H��ė3-�(��'@��C��6r��#���2��c�'�D�I��ڂ&�|��WE�./?���
�'zz��6f�T�0��Y�.w敒�'.���� 6u�H; ���o@���'!��p�F8.�>���*T�fŜy
�'~T�0 o�m�$���E�b�0ez
�'j(4a�4s.�H��S�/����'I``���3n���3�]�#븬P�'	p��sH����ȕ��0OK�� �'(��Q��p�؁��LD��
�'5�D�q���|�c����x�@	
�'��{��P�f���CԊ�� E����'�z�1�����j�F!�8!���� Vt�c�;_�T�@C@"wK@1p"O�O����B�� �ș�"Ỏ�K�(6=X���95����"O8�d��jx`h��ؠi���3s"O(yHCO�/T��#��!C� YC"OpXK�D̠D:�2��N�$dau"O:l�O� W��!HCQ�Ig"Od̋@�_�"��{���<Fp�r"O
��Ae��A��a�E�RL�L3e"OP����	���T(�GT(*�"O�R��=�E9��,�j�"O��[�4W��&1C���0�"O2a3�2�����]�w=��rf"O����-��m5��2b�!�]K�"O򙠢��+NΖaBկ�����"O@,�Va�lC�U���D5-TH)�"OZ�@w�L&��DHũ3� � �"O��a��_�0�N[4I-'t�{�"O��h�c�Q����d8r�"O
|3���&�R��U�� ��%�"O�ذ�ׁw1�E`Á�k@�<� "O`@��#4�D}��!Y�}0̽˳"O"0['
"a8l�#Bwn%X�"O Y��ÖF,x��� ȴ�"Of����M�\�ɂ#E*+�R܂p"O�$sK?v"Fc��|:�1"O�3���n��fG]Rs����"O��j�a\
JK���Ui��X�0 �"OR4�u�M/;��᱁TB@՛�"O���OM$S=2�H�X�x̢l86"ONp�^=&�����
3�p��"On�avN����� "�n��"O�*�	�T&\���&V�nq�"O�%{���*�	�� ��Li��"Obd��А�
��υ���h�"OD���Ҷ8�Bh��� 5<�̪�"O����Q�5s��#U#S~���T"Oll���Ъ#b]��̚jD��4"O�b�Mgй*�.�9��"O�l�'�5E���b.�
6��t��'�1O�A�T���zL ��@-v �#"OD`��>����M?~ Py�"Ov�a�������bh> �$��2oI!�DQ���0�bG�J���S��@!��2at⁫� ?V��E�V�P@!�D�3Ы��!_9410Ǌ��y!�K#K�΍JĪE�d'�|�P�A� M�{��$P+04XȂ��-ii�H��L��7�!�W�|�a�iHzh&� ӥ�"/�!�ϙt�$�R�G*� I��

�!��*i��
����?6a3S��(!�$����t��%e�%h�Er�!�d�7̺�n���$�s��T@�"O`�	B�B&���[bʗ>^i����'���
���6`�]:@�G8��K��'D��Y�@OS��`A��aP�@�b�*D���bK�z��Q��)�P�Ԉ�gk$D�����ρ\V ���n��jB�#D�8���'�2͓v�
t����B�"D��f)Z�|�0A�,��<"�
?D�xr�����$r�b.°Ģ�	"|O�c��
g-_�r���O!+\� O?D�|���1B_��h!���cr+)D�l1�`Z�l�L`)�!�
]f �xe;D�� �H8go�������%��Y#"O �h撙F��D��5��eA�"Ov��v�Q.p�+�J̄_MF(C"O�RlO�c2F���.^:JP̂�'�	 hQ��!��M"V>ܹX�+���B�9'Y�m��ۣfʉʶ�Ds��C�	�3��HK�N[nЈ� w&æ&�B�I�C����ض !z9�b�E9uTB�Ɇ8X�p����e��H�㞽�|B䉐C���{��֔�c�[�.C�I"��ڐ
��8�h O�QG�C�I6R�F�3.��;6 �S�G�1��OF���U#=�b�o�46pm�G�H�!�Dؼ(Y��P&�5z��P�oTe�!��pU����.&�~��b.߀#�!�Y�,�%[0U��M��KB�L�!��&�x=C��pΙP�L�"�'%�Hc�PBn��i,F���p�'��	��!ךL�Q��=:�`��'}�M��iI��Q�`��* ��}z(O��=E�NʲlE��b؆{ �Whǐ�y��ד;�~p+�ϒ$" Q�����y�C��OW�\b�
��'�c�`���y�M=_�����J��0���^��y�c�u�Fr�k� �;����yA����=���юL��H���+�y2�˟,� }����u���#��8P�	ϟH��a�IV�'��gP:�P�s�M��:m�	�'��q;P�ܱA�L�������'�.�6	���0(E�(]�
�'�@P(�mE�]pXxs4iӴ;Z��	�'cΔ�b/D?�@t�Ķ[�xH	�'��	�(Nu�ec�bqb��'���g"̚i@6�p�gݛE[:�r��?�N>Q/Op#<i�  d��A�+��x��J�<��A�p'�K2�?��!�a/�����q�S�O�Z� �ᏎH2΍�Rhƺ#�F��T"O2$SM�f�ʍ˕�9�a��M7D��ʲ�W>J����L�I?�e���?D����U��4m��*sZ�]@ph?D�PKX�"�~�����t�Q�%M�<��
Į�p#�lD�8B��k��a��I�23�
ݗ5�2-�/�O޼�	����?E�$LPX��<Q3��3K�(YҮ)%�!��3�T�ZB�ɺ;]`�1�͗#U�!��&W�\\��瓪N�p���� �!�ēr �`��"��"u��7v�!���T�J`P�Ͼh� ���#\m�!�d��x�^��$ʁ�������$�!�Dǣ��)9��/'�ε���M��)�'S�n��5��pߴ�S�%A72�ڬ��'� ���@�8,y��H�zH��z�'��U��K� Wh��YW��<��0K�'K���Q;~�2�[�_�3=|��'ڐ�+/������H(P�8�'?��bT�'����F�N�
���	�'�����0D1pI8V�U#�F��'�9Y�b6
{ZX�Dc�tB��
�'���A��J)s�������qB �	�'��%�{����㊐�h�x ���'��:E"�>�ʭ�S�ȺP8vT"�'Jv�s!��j��}q"eǏt���c�'�޼;��C&U ��؂��r6&��'��(e@-qVʁ�FW�t�6%	��� ��b֛QAҴ�bۍS>�"O�j��t��QrL�(F�邱"O��2���/� y�2KŜ&4�i��"O�E�@��0u�X %�� ���g"O�D��͈W����Dب)k���V"O(xiƆD�iU����cF�Y��"O�@��(ħ7;v�r��Z $K�yѲ�D�O&����,"s��B@�_�&��L9f��=f!�D��S�A!�"p�Py4�9%\!�ĕ5���B�Z#'��}�&���>!�Jht��$��r9�} e#P*H!���8'���$�E�P)�5c�e!�Dʄg|I�5#_Iv��!�;BN!�ќ��0���[�Sc�X��BֲR��'��'�a��`A��J���X�w��@�e�2��'az"k@�R�=h��	|b���-͋�yb D�ِA��KYuݸ}�M��yr�[ZpQ� �	ss�� �I���y���47��#܈gc��k�	�ybE��I�$`
'�=`�A��ڗ�y���Դ)űPk��҃�F�����?�N>���h�.@r7��S���q��F,��҆9��:�O�ѡ��7K7�[#��,�D�CW"O��s�8a"X�q��Ի2���y�"O`9����i	��i�j�s�4p;"O:(2��R�s'�
fq��K�"O�E���K��|��ʔ�&��a�!"O0�:� Բ~������^�AkJ8p�\��%96���ܑ����#��<��LxF-�w��7z/R�pB̉�q�d���N&x{�V�,^���ņ�8��ȓM�8�uGN�z�������( }�ȓj�t�F��o�<���fL�Fr���9
TA��BˣA�:�惔SY�ȓu�iG.���]����>/E��J2��0�ʘc�J�Pg�;gEb����	�u�a������
��,ܜC�ɎZ�������D�҇�7�|C��/�@mH֩3������GJdC�	'4~L)*S�ѽ6��hh�%1&C��[�@5��M�Į�@�w��B䉱7� }����Y�8��dы��B�	=�Xi���p6V�Ѧf[�Z�B�Ii`daB2��30��x���Jf�C�<P�.cj��~�f��S�(Le��Ē�9g�qU̗!ZS:̢��[6!�#B����i�(h�tkZ�3!���=~�P�,�,�x+'��*�!�d�g+Ȇ�4
�(ɂɞ���	D�����  �!�����A$m��[R�,D�����78�(%!�NK i�H�j6D����F�'TJ��%FȞ9��='�3D�\���>{�����c.�Y*�*04�X��N0~��ě��D0=[��a�<�W&߸-?l�qK'o��<"Te�_�<�"�Ɓv��5�FV$'G$�I�@�w�<1qc�05_�`�U��`�.H+(	m�<���J���F�>e��X�q��M�<�1��Ǝ����6H �C!GL�<1f.وn*RI���г%:�����Hh<	$	R.N��l�͎&	�A0A�<��x2�͆U�V�Bң� ���S�!�;+;�1�Q`�?J�<aB�,�!�D��4�b6�+X�� �=�!�� L�s"!+mf\x�!���(���{7"O����H�I*�DO�rR8$��"O�z'Ś�$���ßG� ��O�Y��cND��&� ��&��W�����<�5�G.[�p͐)I�iҖj���D?�8��H����j�*x���g>D��s*J*��E;À�N���t�)D������"X��D��/�Q���(D�T�A�նY<쌉@S%��C�M%D��J�R��=#`n�?K�\fO&D��x�@w��RŊ��x`�P�*?���O���>��H� �,�t�H!D2PN>ړ�0|��P�;�h����T ��k��t�<��6D��=	(׉�jlk��z�<!R�ڙ�hi���;�Ȣ3(Z^�<�pbD�}r��q�Dػd��aJ��a�<)�K��x*F1�m^�\n��7Aa�<��C��R��EG�4���E��UyRW��$��|�珃�k���V�2&���Y�(�VyrY���	s>	z���v����?4��;�,D�\�H����Ms�"9���4W5RC��4+�2���n�y���6���K�HC�/���c��}0�Ё%�sW�C�	�#���ÀFAP���!�45�B��4�Z;��	�!������*B�ɩS}�hs�q�¡��b��v�x���8p	�@'Q|&�9��[39��ȓw�z���-رH� ��D��U�>L��{�,���P��{rAÅHR�X��l���5,ǯ�V�;���5j(�ȓA���r4��c�Z��'��Z�"��P-2����2��-� ʣ�ZD�ȓq�x����>���jp
!\�1��$�� Ō��7%����o"X�����| ��K�v��e��[�4t��ȓ\�z�ٰ+P�
T:�3���vu�ȓY!x����o2Q�fk ��lŇ���  �I�.��9���5Fd��A�`|	�fD?!W��L� �:��ȓ9_���(Ϗ5iJE�3�*m�M�ȓ@�رdo�)BB�r4��ȓ���R��W��NИy�a�ȓj�$�t�ҥ�.I1��D\�مȓep����[� Ӡ���b�o�\��ȓ+��	anX�AE"����Ȇe�Ѝ��I�<A��߳
��L���F=3F��8e�\e�<�jA� 6����V�0gfm(E��_�<Q�e�;�%�deډj2������W�<�`I�b�J8���ZWJ-�OAP�	S���Orް�G���l	!��S�s�iC	�'"�q��;Jdc���8M�xr�'Ɔ�"a�)
��1�Y���\+�'��q���3b�\�R6��_1�ńȓ:��K!/�"345ڰ��sV�͆ȓe���4+@1�třp
�=H�Ɇ�eg>ѱ�NE1���PfY�2W�ԆȓjT�֏��{����&�-Gl�h��#�
]R�f:
_ �pRi��sO��ȓd�E��F1�.��pÀ�7��x�ȓE� ����?.���K*p���ȓE�Su(N�>��@Q������ȓ"y��3��1�`a�S%T:'Y���ȓ+ĠMB���*,��,��VB���`3�U�0�[�=�L@��ɰ[p�l��S�? �<˳��S���K��{�h(K��'U�$(>}>�)aG��B� Y�4N�&m�{��$�;|KLx�H�V�V��!m�"Q.!��+ ]�H(P���^�r(PЬߟ3)!򤖤1v��[�,�0��؃Ҭ�8�!��8W�5�3� ~4Y���#�!�d�]�s�n�+u*�"����{�!�.z��e�P�*5��4�����!�����I>O�M���[T��01�Iٟ�IŞ[``9��L9��py�� ٞ	��	R�'D��thHl��xJ�+Ё)��N>�r�Ҡ[�)Y�p��P�ajPm�	��Ѕ�	����q�B��jj������18C�	\ �I�c
_4V���L�&/C�ɏ&�Zղ� V�Nٙ��ҏb.B�I�B@�V��oX"���-t�&���!?a#�k�$536��T#Τ�c�ux���'�fp{�刬}��)	�%)� �����hO?�`���*x-t(j�eH�I�fIŤ�pyR�'ʶ ��DG�^�ft%@J�M�HQ�
�'�����l�T�yt�Z36��R
�'�������K@���SL̤x 9a�'���Y& ��XsLR��D#� �8�'bJY(�F�'?�%��O�Q��'��:2��@�RS�A����?��y�OR
w�h '��:&��qp.��?��0?A��^�G�Ԉc&Dgp h��XU�<�Sd���x��G� �jٻ� FG�<i!�ѥP/X<��_2�XiAΐ{�<�v).�^=�pBΗSH8��k�z�<9�-��]��5��-�-sנ�q��X���O��T"$���]36�Jb瘿Z��l ���'>� �L7 fء��ZQ���'�|���O�u0i9DJT�M�F%�
�'�Pp�%�D=@**���6J0<���'"d��GJ�� ��7B��+,�@�'Fu`�o�?Y6z�Zddȵ(����'�6t����=�!h�Tv��(Oh�=E��ENZB��uD�5^L�Q���$��>���y��g���r)Г]�Te�#��y�A�n�.A�U�\�S�؀B�͟�y�̜>�	��,0w��f����y�[U�JdB�c:W�ƴ@e��(�y�^��V�1�#%NV�#����y"�E.���#�� ��P��%&���)�S�O��2�bE�t+�ɶ�F�1	�'�,��J".��#!��4x�eZ�'��쀕�˚�0e��ލ@T]�
�'Z�	dK�\6��`��e�‪�'�
�1�QllIk��\��H�
�'�
��`
������؀Y�QQ	�'�L`�iQ�k���
R��`�p�'#,��T�J��j�KI�4	f@���?A��?�����i�ODb��	�H��8 �\��B<��X���>D�0P�.ޣw���2,^��#ĥ2D��8�7K�Hԑ2=�/D�`�em���X�QE@-E�F�C�F+D��0�_�-�� �� �R���a.D�0a@3E���ؤu�����.+D��ȡ/��.`8��X	K�<���OP��O��$�O\�'�?��yR�99�y�hǹt������O9�y� \�!���Ch
�8!�/�$�y���F��<�&.ˆ(�R�O��y��!�j��7M6!C~����y
� �8��T�e��x#��s�6��2�'�1O�xwGDr1HQ�����Fex"OX	qWŘ�Aj-��[�y�� ��'ur�'�R�'��ݟ��<yen͒/�DKf���UHv�I�A�<i��˵�\��l�BK �c �2T�́wNޏ�J�)��TAQ���ph(D�ș��WN���t̑�^��"2�$�O�$�O6�ɇa��j���1N1�8B�'�h�S'�Y�B��"�:5�YH�g<D�L��Gԁ=ې�	��Z4H�r��8D�qbl
0`E�s��Q\��7D�Ȓ�+5�Vj�H��Fa�F�'D�T��F�V�h���g�C�PX{�$0D��
��7F�\dKu��%)�x�u/1�O�re �����`�D\hbi��|�B�I��(m��g�+;��T*�k7\����0?��Mԍnn�_{�t��J�M�<!aB u3r�3���[���HaEo�<!#��+5'lQ� �צa�� 8��Vi�<���I-f��2�K�-�mbGT}�<�C"ө�\$�5/���y��d�<��-^���A�����ND�I3*d�<y �=M�`��B��J*��ƖG�<�'%S�ZH���&��=���9b�L�	T���h�@��)��+G8������$D�h+F@�Iþ0�sHG�A�hSA�!D�к­�:�
LB��DG�aP�?D����G�,��Q�jͺH-� b�!9D�,p�A�)c�\#�e�L���ا`6D�<ʆ�@E���b H�)-���b� D�h �O�O��a��*�"�T�*Q�=D�C%�"Vȡ�MQ(�VEa�k=D�0��QR��e�7'�j-R6�8D�LK�BQ�EE>����S�tB��6D�\��KE��C���|zj�(��7D�@+���e:Ɛ3cH�6f�isD!D��1
['x�dQq7ʗw]�!0R�?D��5˃OW~�(w$�,��"�<T����KV�V��n��GCl`�"O�qz'ϛ3��
K��,�"ObU�"��f.�,��H+ԆM��"O�M0��<p~\`�@�h� lsC"O �0S�v���"i��M�<	zr�|"�'�az�ڬŊԠ1��lr�8:�΋-�ybh�F�
Tp�%c���ԅܱ�yr푌@T-�q�4\Z�)c� �yR̐�}u�)�bL�\k$u���T
�y���z��Ԓ�l�$c�4@���y����pB�����%/��yr�W�!g�L��3�`Y��hOL��ƅ+S��P�Sj#�4��$�!�8~��+Aj�N2��a��J\p!��\�b5,qcr�����eQ(i!�d�'yt8!��'\�6��,0%�G�`O!��?ʄV�Q|��;�Q	��q�ȓ_�(9��O�D�D���\+�	����1!ǜn�Xpy�R78֠�ȓ ӎ=K��tE��'��6�����Q.1��ç|ӰqR�쓨���~��ń�M0���V�I"G.���ȓF㢅3���X�ʼ�t��d<4Q���r���σI״5@QH_��̆�Z�rb��MQ�;��C8:���#� �N߯/��]����:r���S�? ��j�8O��Q��ә3)��x�"Ov����Uxp��,���x�7"O�I�N�/O���EK�1x��"OV�ڐ^�M>�J$�-U~�%"O�]���+5"���H�}��"O�ܘBeT�yKN��q�
�7��A�"O�p�D�A����`͵%&�*�"O�T#�@�t�B�k��C:�H�"OXt8у]<k���Ӗ��4)D1�"O���#�^���|�U�Ρu@�A�b"O�t2��]��V�� �աq'PH�"O�=�D�_�(t��ӝ5>�+�"O2�ZW%խm��ր	�=�ze�a"O���T,��6z	��A	�,�L�v"O�U���;m����Ca�f��%� "Op-����M�����`1K�f@��"OЌ20m�'4!�L�o��d��"O��B6�P�,�h��hD�s��01�"O|�P��R-*f���Ҵ�,�h�"O@Ԃ�o��.�R�ѧ�݁��$@�"O�ԛ��Sf�c����Ꝓ�"O�Z'AH�kn&��ĦG��p���"Op�xc�L�
D��ş�Y�jI"e"O�i`d��f{��d���""O�5aC$�4K�0�6�ÓM��b"O���ek̄:f��ъ'$�ik�"Ozm1�K� #/|-ZcӶO�q"OLh�&��D
��[���`�"O���0����b�x"O��7�՛@"O�Sv͒�n	��(�,�N'�8{v"Ò���J�  Y��\<��i�"O:1H�߷��Y㥋ҒK�x�`�"O�ѓr���e�d���B�X@���"O�����4-ȭ����!D��"O�ɚ0�[�fp���8�p�"O�`���Joh����.Ɇ_ДU"O�)���!*rM��ޛq�Rz�"O�[���| ��M�+z�ЕC�"O4��.�	@�qp�X3-�Ե2�"O0�8׬�d2�`�a�94˾���"O>A�Ee��z@���.R�V���Af"O �����,	�`���d�J���� "Oސ�ꏦ'���Av�H
H�X�9�"O�0z���)8rH��5�I�pr����"O�0��*�+8�j���H�-MR�4��"O�|Pť^�*8fDabn�l��l�g"OȄ!֭R(=?��ǍN�o:||��"O~�く\H֨��U�6�$��s"O����z�h�ȱ)B��8��$"O}�eK$+�1�N�^�@!�"OT��a�P�̒���,�6��"O�h`r��=I.�ER���i�h��t"O�ecã�y��6a�W[TtKs"O]�f?\��%@_�D��8"O���%���&�z�c�o(���"O�=�H����DX�@�%Z��0�"O�\�r��#&�Btxq�V/�$��#"O�p�&�����y�M\�`�@��w"O�¶�Gkp�c��`���2q"Ox����)o(	8F���v�����"O(uj��am����M�W�H��V"OZ�K��V7x���[wE�"����!"O�I��hŬ2�n�i���h:^="�"O|��G-�E0:����)l9�� �"O�  �������E�� -�Z"O�����
"�a{0f˕"�q�"O�(#��X!�@�6eLx���3"O|ADқR/aR�EZ����"O� re�I����:��֖�<ѻ�"O|�Y3�/pi�@
�cU	u�քy�"O��lÜ2�4�00��"[��A��"O��I9Y���b�0מ��%"O��+�i��>��@����
ϸt8Q"O�	j��8��ȅ��>�y��"O��裁��O�"�۱Ȍ�iT����"Ob��.� �f�%�'aK���$"O�I���زq�t'۸DD���"O����7fLL�匒:V$ x"O�a��6�<@���	���"O��PA�C�
ݜP�
�@<[�"O��$�[�YJ�څ	�69��"O�-�"�=�����\� xIc"O4}Ñ�� �q���0d��=�"O�4���ĄuX�)07D :XBqkW"OL�
�F�<^�]�4MG"{��M+�"O�%�d@	�9k�aۖ�M�M�"d��"OVrR�܎3~�uyï?<m��SW"O��Rw)I.0���ͻ2\�U��"O$w��1kJ�A�5'ݎXС"O�!��CV�"�P�U%C�f�8�"Ob�h`iD[�̔X�#�2D����"O*؋�	S��22m�T�i%"Ot��P�+@�"�������h}ڠ"O\P2T��
qC�0$���}��8F"O�9�!���N�h�e)W ^.�X�`"O�)q&`#2�L�'�^ez� 4"O6�K�e�Q0�-I���~� �q�"OD�p��	RD X�oӔu{̹��"O|��"!H�2A���T�8��,k"O*,��@�kt�� K��QyZ<��"O�$ᇇ�^{l@�ҙ|`��"5"O8����d|�pQ�ʓ87Ih���"O<UI̕��b������y?j��"O$��C�� �dP(e�NI>�02"O.e��.C<;ކ��VeC�i.��{�"O���ło: MI��E0 ҝP�"O*T�E�L�Y$��!@e�&��C�"O,�snߌ(`\�e�ו�
���"O��z@��d7����R����;��d8LO4��FC�U���Wc�%�$8��"Oj�(u3� E����<�R"O�i�0*��:�8l����*���"O.�PC�6P��[�◭N�j�G"O, bs�48/�0[T�C�*�:���"OXȡ���E�h��@�Q7�8\�%"O�a�E�#�ݡcb��,r,�"O��HN�7z�V�)@`ʑ(˸p��"O��'�b߸���.��-*A"O�4��R������P��%��"O.U���I�-��x� n�t���·"O �kV,Q?�#g���V���"O\��P�ƥ u���>"��A��'����i"��9��&`�sA�\�H�!�O' �[�͊��f��p.$=!�L�� H��"�@�p0�Wl�S!�d^,y�Td3��1��E�k�!I!�$&>T� �(�?:n�4ҁ�-Z�!�I�\�֨�4)^+wet�K /Wh%!�� �SpT�Zt�q��.قb"Oz�H6�MF؈��Cv!��"O $ӳl�6E�	1竃&a	�]�"O�<���Č'A��ࢭT�!�ʤ�5"O�M�e��<�<����@�(��'���~b��Y=N�Ӱ�֮���RtH �yrlj��BqKP�Q�C�y��x,)��m�5u�@hmS�y/�
6��*4��"l����5�y"d/s~�@�mǮh?�E�Eڒ�y��6v��a�VJQ�Z���ӱ���yrK�<��a+�ʙ?T�fբ�����=Y�y�Ő<��Y����S<����y��	!^�mxա@�Ihࠈ$葅�y�^�C	�J'
§8}Թ��	&��>1)O�YQ ��,�(5��?�d[C)=D��B�KaܒXh�b��ic�p�2h7D� ���8�X��AOR�3�O6D�d��CB����5fƎ2�V�p�C3D���� �$?�EjT���5�R��r.'D��9%��rTb$�bM��>V~lAsE*D��xT�N��I��խp���;U�;�ON�IP�tcÌ�n�z��%J Z�C�	�i4��Ή��&=��jB-s�|C�I�S�̔�Ҥn�P�q6#L'29jC�"0Ǩz�O?��9�v�KN��C�	yizݐ1���e΂TY&���{��C䉷���:��4}F8@�-(��C�	>:��u'D�'HD�(�&D��h��d+?�*]#J��T!֙i2V͂D�J�<)�$P?u�y�c��
F��l�B�ɚE̼)�AJ/�1���L4�JB䉸A� ͠������O�q6B�ɘf�"% �	�6"p��rk��$&�S�O�2���G^�2�����H&yJ�!q�"ON�C�o��p$fL>}>x��t"O��ٱ���C�tL��G��w��y8�"O��s��,Kg�ES���$���1"Or43K� 
(��Z���!pl��R"OdIBf"1_��Y���-[Rls"Ov����� M=���c+��DD(��a"O0ԙ�d�2�дK@�ەmC��(V"O
uۦ攏SQ<t�tʑ =8T��"O����J-f*U�C�BXi� "OP�� N�.�U�^'���*�"O�TJ��%�(����#GL$��"O }(�b5�j��2>�q�G&D���لl���'��4V8��$�$D�) Ǔ%~�Pc�o� <�fa��!D�,P%n���v��8CT|i� $D��A‒)���+	<Й��,D����A�[�P�`��D�R�`T�!�+D��Uk�2�
�{��
`H"u�4D����18$��e�@�[�"�k��4D�xB�)��;R���1��92xP��3D���T�J)?2�3u����X�7�>D�H`s��L��+�ᄌ`\��e<D�0���#6��`SJBɋ�Uk!��_��8(�2D�(	#��]i!�I�z��dJ��"2�d�ȃ"J9`!��G�C����(D�*�҅����!�DR>4����Ğ� ��b��$�!�$�Q%��6�I
4�*U{�R�P�!�ě!��̙�"�{* H��&Z�!�� (a�@(~r�2w�ݪ~�zXˀ"O܉��D�z&�a�떓=�A"O�E���ȭW��B��Ҏi�dܢ"O��ei�t�E�F�̂��]��"Ot% ��:*�XS����}����"O*�X��@WJr��HC$w��;"Op,Q�HN�.�������0�p��#"Ove��V�w:�%��!�2�Hٴ"O H#����%���M�U��a�f"O��x�'B�'J�ڡ�0����"Oެab'��+�50��Br0�C�"O�	�5���j �1��B���U"O,�(���)�
j�d�f.a��"O���4G�H��`xc>&-�X"O���-
����U�!.�"�3p"O� �$�2B�,�q��szܙ�"O����F0W�<seEǔT����"O��l�"ld��� �Ex��B"O�(��H�x�����:��	؇"O�P��%��|@�w�њZ���ڲ"O������Vj�i5�=a{f��B"Oܤ"ǀ�iR�԰$
V
M�����"O�h[�Y�s~��EC��zߔ@"O� Hf���*�ʡ:t�A̞K�"Or=�ԤÈ(�` 	���w��m�g"O� ���ђn������$v���g"O�q��mF��
!aFN28��X�"O��
�g�i=���g���0�"O�岀�A� <j!�#T6}��"O��륫C�@�f��"�;'�>Xp"O��RKӃn�Px��Ag����"O�H�w�#t�$|qj�9A�,}(Q"O�D���C�J�F)��ґ/�l�a�"Oʨ*բ�='�X�LڊU��Y�"O�x�r�C�2P�0��2�f�)�"O��F�ψ� J�mN�7�l���"O�@@CdX�A\���cO71�T�	�"O0@IP�=z��xQ���Ʊ
a6D����+Q�	S�$a���u����*3D� Z��B��8{�*��$�T�<D�(�7&�zp�I����q] � �	:D�L�	��:<��G�Rڬ��ǃ,D��87 ͛eWD�9�`^�]�꩒25D��薣ǡK�X�"W�r	�(Z"1D���b	8W��͊ւ��N�1%e-T��
օd��(g牘hTA��"O.�`�F�0�q6:RΙ&"O�8뢯A'FQ �aƦV�U����"O�t@�N__����N� i�ܱ�q"O�	Q��I( `���C��4����0"ONM2��Ӥ&�n�U뙐s[��`"O�Q�3-أp,x�i����L��X"O����`�?��Ёu
����p��"O>��C�.G�cL��m�8�k7"O����M�=,�R�ʗ�S�l"O�e�낚,�`���ۤ�|U#u"O�m����k�����(Ց]�2-c7"Ohy0F�2yQR���	̨Q��#"OLข�inP��h�2i|�)"O�	
_���S'ڒ#НK�@��yތ+ʂ,Y��\  � �22�#�yR�P%Ɯ�2f��@'��DÞ	�y�oBi�`)���51;���W᜹�y�ˌ=κ]��%֒)H�pS7�^?�y
� " �S'_� mYOp���R3"O�QX7eH�
�Q5h�g����q"O�9
2�wYD����\1� ɓ0"O��Y�GM ?`����@G��8��1"O�����h*)�P�]
8���"O���bU(h0� �<S7Y�f"OvQЗ�ͱC&����q�,X��"O��{R���H�,7eђ��Q"O�,"�f�,@%.��`퇂l��}�T"O�8)��P�y��8⡝-R�"OReI3��b�1h��'PBȹ�"O�a��:�БfaDW�H�"O�t��j˱�"٩��U�� 3�"O��XDꙮR9l�q�FZ,a�nub�"On���<uRp�i��"du��"O�4! 	'y���ɴ*�<V���2""O�4(�����X��IM�,��"OHM�Q���Jap�z���.�D���"O4�����`��M@�gմ�Lp�"OQ��wH�yhĴ*r�	�"O@%a���o^<Z�&Y�nn�|IW"O�j�c�5� \�`��?l��T"O��	�a�����X��|{a"Of{���s{.�ۑ��lפ}(�"O5R�Ա��Z%�� º��"O�� �!�f�`rd�HکB�"O���J�h�b9z�'䌚�"O�%"��S���b��?I�Ě"O" �� ^#B�
���(�~=�"O��1�N�-8���1���*~���@"O���`���Y�HL�d�2�"O>P��+�_z<A�̖6�8�ȕ"OT� �&2>�}��,%��b�"O��[%*̖1��Ƕ����"O�x�t�ի]�h<w�.m2y!S"Oʁ��X�"L0��7�˗(�f�"Oʠ��C	�]�V�WƘ��C"O�f��Gߤ��s��>�X"OZ���b�d����5$�p���"O��2���(R�� ���C)jP�"OE�B
�v1T|X1'؁�� ��"O�%��@ɢv��ge�o٬�K�"O�1q%�*p�pZ��;@�t=��"O�1�q�#��0���F�� ���"O����']�3'�yxr��f����s"O���&��+�ʵ��̘���"O�� P"�?u��q���?�rh�G"O�%�լ��������W�"�xU"O�9 �٤	&Hh�0��>z��Q�"Oڤ�U�_}�����[{��Q"ODu�4Ȃ�)��ݦ5��!�"O�l�3��B�%�$��_�xY�"Oty�ǂ	8��bB�+gtB"O����;~�$���ݨdY�lɗ"OD��
F�:��p& Ĵ!D�@X"O���h�
C��<�4��\Dn�Ps"Op���
ȓ>���D�W�>5�q�2"OxcAS1�.p�7�eI�-��"ONL�p��	��pˤ�ѿdH��q"O�=�7M��^�ܳE�]�c$��Yf"O��G�F79����Ug[3y���x�"O��贍ؗyR ÆWJ�N$��"Od�K�B9G�{�f��=�@h�"O$���[�����UO���("O� �S1 �)X�m}��E�3"O<i@�ӸJ�.0"k�N���{A"O��QɕLm��YF*�l�H���"O
l;EcЁ!�2���Ș�8�§"O����Ň�f��b�֠%zP{�"O���KN�m,zP�#��Dt �Rw"O�!#�d�'�Fh�cF�� �pY �"OD��Q�9߾�
Q썽N�<�*�"O���Ʃ	
�d��JKl� u:$"O�*2�M fY �	�ѻ?���"O��q�«R�>1��H�']�0�j�"O�)C� �5��iBɞ�[�p��C"Ofă��NY��ʷ&V)3X%��"O����x~r]X�˃�֭��"O4]��<L�n��D�P�<q�}�S"O��AH��D���iL�]vR���"O�ԱS���!Z�J�S�/Q��8�"O8��cƘ�gAL�V�Z-n��q�"O�D"c�9% i	dѵ"7�x�U"O��4��5$D(���5ʵa�"OM�#H�-!�Vp ᦉ�B1r��D"O4�R�%s4E�׫@�b�š�"O �a���2o-@[�T�^���"O޽a��1�|�[�K�H�(�h�"O�A����VU�5i��,�:�`"Of�Xs%�Q������$��B"O�1h@.U�.���T�orv@CV"O	����2(N����cK��pc"O���1�� ��M���
25�0��"O����䐏T�x�s��Y$S��[�"O�HسbB�>w����Tz$��`�"Oyz���!d�šQ��+�<1�"Oec���	w��W�?�&\YgGl]B�	�`��)˷&�hk�g�%^0C�?�����&�~�a$���[]HC�I�m�� �W
NBZ j�@:|C�I�u}8��'89�D��KQ.@�^C�ɞ#�l_���!ʂ[�rB�	]�0Mq3JғVw���boI*(�ZB�I�B4�聆�B����'�.Hw�B�	+-�Ȥ���	W��[�/��u�8C�	�(��C��6�H<�îK�y$C�	�=V�I�����Ҹs�bD�B�ɘRj�v�(1��xbt��0*аB��ąFf���ǩ�7'���Br#>D�L@A��;]��Y��q�Ir��:D������1=��|��*W(}y"��<D��&��2=hm�.߬Pi�Y3v�n�OZ�S��M[t'QGؑ��ٸ���'oIX�<�����,�
P�
�*+����s��Q�'�axɕ�;Hb`��/eF9S���*hz���>�I���X��J�hA놪ܫ	� �y�"<���Y
w�̋CmD_i0ۂC�9U�Oh�=%>K6F9rn�!Q�n�0�8 ��%�<ɛ'4l��Gx��#d�uȗ�^� 50`FS���O�#=	BY1T�1ٷ B�O�Q�v.�]b(�Ob��B��<��R�e�����E�T�x2��* ���+�_��Kg�	>
�C�60>��[����XW��2 �8C��<gPء�
�7����K�C�I�Yk�˃
�;*X����*A���I]y|ʟ1O*�#���@:�^�oR���Q� SA�)����b@W  �Zt������IxE�{�$��Zx�P�!�Ďg����,�(<j�X_���D!�� �|@6����Vd��ꃱz{HX��'�'wr��ɒ�F�i��_m��ݣ�фzlB�ɭo��Y��O�u&(��[�h!LB䉘XנL�.Є|�a����F(��=��"	�����q�b�Q��_3mK��%�lE{��4�܌6��d*��X��3+J�.�!�d��1��ÂݼnDv��a�F
��y��t� $�tn�;ZAd�����C䉨���j������ K�E� Ol�=�~�AF��}�TϠb(H���_�<����
?�^d EKV��0r"HY�<�1���h�'�
�iQ+����B�I�o�����IZK@����_�pB�	,}j�B�AŴG����m\!s�����O��	�<��sh�S�xQ4ۉAC�'cI�����[�r��ك�sO�C�I�nr>%*3n�/Z��$yTGR�hC�	�[� �.=v�b6���4z����'k��xr����BE�G��!h1�]����L��qTJ�=E��P�t���o���w��<l�v���ܰ?��j��`@v�2Ç#/$� ��m�=�y����5�f��vS
hj ��,�y�<	��E�#R���D�m������]�<vaT.A������$��nHX�<��-ж-@��r�N�t}r�L\�<IrG^ ;�P25/K"`�E
�*C@؞��=y��ݐG�n�z�bU�`a񆎏|�<1�d�j%Bͳ��iZ��#��z�<��E�S�"���A�V�L�`�jVz�<��G��^h|qvhMt��3&M�<�,S�IۆM��T�4.����
Jy��d��(��$���p�ǣ/9�t�P��ēr(�)���b��� $4�#u�F�HIec�F�>!��D4`E�I>!�}2�i6��Ce[�5j�1���8lغ�OzOԴG{"�'�P�hw/Ȫ<����j��#����p<a���'����a�-�"�Y�� �<D�V
O�Z�l�1bִ��B�{H���F"O�1�F��Q���x����B��;��T������TAD�0�b��3*l|�3- 5%!�Fb-�t t�\�+�J��D	ƅy�=E�DcŦ��y����$ ��t1�
��m��')�|ALφ1`��U�$��5 �zQ��� 
ˠX�,��S�N�؝�!6D��;���2�R]�$�E1�g
.�D?�S�'$�B��N398�ѓ�)(I^�ȓ�Mг�& nq��+�|e\y�ȓGFh47(ǫK�8�2���7�Zt��<5 P�8&1n�����6 ����ȓn�9[�/[/?�d<��A8�T���d0�؈�c�`���"`K2�X���T�f��u��-m��Jf��-f)Pa��r���i��hn�a�w@ͱK�ȓ#���+Ο$J���1GbǤu<=��A/��IC��z2x`�H#$}���ȓt�n$[ ��GO�e�j�xo!�ȓc�قȚ5,=�A���3^�d$np(<AS�S�hB}kr�ĩ2LX]��!�v�<��G�,"4�rQ.D��Yg	Eq�<��
�&S���ޫUC�1eHn�<q#��<Ap>ѓ�*�*2�&];$��N�<�4	Z�J-��e֤!�����N�<)UA]�iF��gG�]���4�]J�<! �H�a�0 cj\�N5��PG�']Q?l�
XH�MU��d���*�̘�W��B�)� B� ��P���h0w��w��5zR"O���G�m���c�ȹ��u;3Or�Ӈ۬n�B�g�]�"��`�;�#�S�;��`� ��/cX��	,���ȓXp����L�zf��oE�'r$��oz��'-پm5���%O�H����5[.ظ�Ԟ�����E��^�ȓ<�0�W�1����W��+P� �'B�}�`̑��rH[�T�iज़�yrG�<5�4���Pf�����	��� �S�Oi�ɩ�[$(�~�J��"OX�,�	�'�t�2���5}�Zph�B�M��<��'�$�����
7d��m�(ztL��'�����^�M	��*;�~�S�(&$��c�b�WO�a�W�÷)��l�E�'D���X�NM��f�RqZ�b�.;D��)D��0R;F5�c�%p&=�Q�9D������56R�ju�H&���a��8D��y#�H�B��Rj	,z�iw�4D�@t
Ј�̰�b'	a�ihf�/D���6�OPƌ�eɘ��lj��7D�$�o�	n��%�s@��ԡQ6."D�d#U�V6)��$
�	W��vl#LO���!W%P�R��C�(I���/ D�t����"Ӛ�j���95HX��=D��01���w�D �0��u�()j D��{s,gN��#�$�1c�0<R D��.�#%�"����� W�ash�VC�ɥ�v���&U�Qd�Z�(�>��B�I�yv}�#kF�U0�P��!ftTB�Ivͪa�V&N68���J�p=B��.�"y���M�2`����=Ĝ�<��H O�$�&*"��35!���M��"O�X��W���j���	�}K�"Ol\�ExV铡[�,T
4n��N�!�d"|����䆒âѐR�Z"X2!��7~|��UKG��h8�	B�!�DD�B���s`U��J�ZR��N!�C�C����иd����#�i!�D�+�j0������CA)���!�d�3eF ���T�"����
�!�$�-l
6.��(y0`�e`�!�Dї;&V8(���e�����]��!��_�vP�$ؗ	ӉK8��Tn~�!��;XK���Ae�<Fq�E-�j�!�$G�E�+�G�tfx���K�m�!�d�0�T-J&-U(Z�^1ӔM�� W!�$_>u��Q`$�c�z�PK
IS!�$N9G5�!�`�]0������_!��?s{�=���S�F�<K��*S(!��Y1JA	E��A^����CT#!��! �J����D/:<�`����!��V�a=������ZL��(���7�!�D^70АCg�
�4ЂK�1P�!�D�
� y�N.7�x�����(r!�C�R�,����);�$��K�@{!��*+#�(TID
��rf@`!�$F�`2��P�?�r�sd/�MO!��r�t��`�K�z�~ y��N(eW!�dۼH��V�DјD4O̐:E!�$ /��Ъ1a����}W@��1J!�$
����G%�78PL�!E��@i!��i��i.MB,	B&��!��
]��8`���`V@�*çM E�!�� NZ�g��T p� ��h���"O2Ţ!��F�3$R�IF4�"O���� ��DX���g��=	~�}��"O�Ѳ�,L-^���3k�=&�ۀ�ɴ]����#�9qxq�7��d.�I�b�`'��{�|�c6F�4!|B��.O��X�ƾ9A��kQlV WOVB�I	8�� )=x[�ɺ6�W�c�B�	�>4`c���zw��M�B�	�d��9���. ����R"v�B�ɇ����9��braQ5:l�B�I�	��Ys�ߋl٠<#3g��h��B�w]��� $���Dh
1�%�B�I �����Q�"0sS�/��C�ɨ:�E
6,�%_.�wB��i��B�)aީ󕥏�H����� --�B�	7:�.����/v�Ԙ!���vC�C�U�pZu� ��|"B/j�C䉒q�Ԙ���ݐH&��`�mӰe6B�#&��͒W�֖A�NjGg
�B�	,dޠP9�@E�����al�8A.C�	�h�䔋'.�F���a�G�I&C�ɮV�� � ���!��l�fB�C�I�k9BآE��4ڌ�@'
ėL��C�.hl�;GK
�'�J�z�W5paXB�	pR`�w�F�4�`�&FH���C�	�?��KVlńo�H���F�6H.NC䉠 ڬj ��e5J��
�]�vB�IE�|9��w �k��ߌc�B�Ɉ.�N��@ U���r�
��zB䉂Wb.t��/1��]#��X�C��.��#���k�"�41�B�ɗ�(�`f��[Fj�@@
�žC��G�n�aw�гSnQ(4�]!r^�C�	�]D�5��يf�.=���W�C��>(x}I�F�!	�:m�e�7Jv@B��4F0H�Q�喂'���1�Va�:B�	��P̚�E-ⴻ�A�w�TC�8n��!q��{"��5mW7`g�C�I}6�v�.)G��� ��9,�xB�� N��9D�~Mj5�a�}�C䉾A�,`Ʉ&3?VmJ���Kf�C�	�4��DS��"z�Zm�u���(s�B�	�i���@S-|�2e�@�B��B��C��{���D#^�2���C�'6�4�'gEP�i�
��aC���\
�ጇE+8�a!�	I�6B�	�kPP}s
�-@<�h��6@ B�ɛ"�� �� �k0�s�&B�ər)�ۧfە;����*N��B�	��@'쐙`���#'BLPRB�I1$y:0�u��R^0	4i�>B䉌;���%hÞl�هK/@��C�ɵp)��1�$).��C���
��C䉬i|`�P�_04Ct�� \�#�PB�	�3ڞ�9��X2&N2�L��C�ɺ'�������z�YC��R8C�I�9�HbGҮLlT��C ��=)�,9#������_�A�6�Ӣi0&�'�$&�!�����HZ1v�̠enγJ!�m�HF0!�d���S��M����;5��qaf
�	jT�<�bT�<i"K��i{��܀d��pJp�L]?�u�[��8{%�۰<U�!���_�sB��u"�L8��)��W�U8R�CHn8N4�ͭ"��T�e��-2l)�ēÆ��AW82��l:$�JSC�4Dyċ�Ϟ�����0���� P}y����q>�,�C�*͐8�f"O�M�RO�1� `)�dV=]�҈��]�+� �i��wNlݗ�����w� ��I�mN$�D����y��	��p��W:ct��b��~bG�9�ʹxc�ա1ay��9E�H�gI���؆�#�p>I ����ms�Qk�����ީ
F|�gK�OŠ�'4(�+Q�B3D D���!�c��d�D2&�!N1Fb?�9�nD�u�h0�ѯJ��o2D�,z��:��+Ѯ��[��mr�o~ӂYc��2 ��I�"~nڟH�T Q�d]j2���eh̢M���d�DL�-�C�ذ=9�L�(u�(y��׹,	*� �Fy��	�_�, 0��׹/

Р҇Q͖�Br�\�*�xc�혯ag��1 ��}�<�cfL�I�D��V�$/5X��ÃQ��yr��'-�΁�э�Oh���Ǉ����AU�g���S��T MU�1��g@��x�Ue����#�A3`�0d�� �=���P:\6�A��F�Arܼl���,5'�'�<�7i �gt��b�'<h�'�{�'e�y���J�hL$>9pd
��v�P)��J7@6� p�F�pWi��Ʋ<Hs��� լ��D��:=��M�JEzB�+f���$�z�鈜��Ӻ���իN@��5,�2���q�ON�I2pA�q)�>b�2�@t�W4��B�I.4���MF.M8Q��_&X�,�RK�x"�`�O���,2����ǬH8i`m^%^�"�%|iL�B!Fѐ5M�@��9�z���פcT�R ��S�n=2��^�/`�$�B �.��y�W!5����R�N�/ N�2�_���gy��
$ �h$�H�m�8�i6$�V�Xq�G I�p[���)�<~ѐ8B�fV��E�6t����w�I�2&Z}R�E�
_NttS�=E��Z��x��A�yD��'6�A�wF�&~��O����]@��¨��'UDuI�d>��Pq%	! �
��v�G�wObC�I�b��*a/A�"�	5�8nH<�H�@hC��r�6�x��1S�.�uSğ:�-Cȼ�Co��f.1�V�LQ"��ҧ-$!����7�a�!���sI���?���(�Q��Z�3�}4���I>E�įձYH�gL�m�"pA����	�߼U���>Q M1U�c���R.�Q�B���\UR`���>���TVh����=6��|���hH��KN j�2es�jX=�C��q3����,�B�v-Gc�%/�=�c�\j��3&�0�Ӣx�v��SA]!�^q�eN�a��B�I�M���;�MI�r ac0b����Dں׊��Gӷ��)�h^Lē��-�ڔ�$��awnM�
�'�ت3dvOdU!�'3N�I�*O�!ɥ��e�.ec˓$!��Y>KƁ��g�G`Bm��	Dk\AP�� vp� 3b�F�Z��8��E�%���YG�'���QWGO0x� ɳ� t��@@�1L��@E{2���.J��+���@�jS�y� �B0��W�T�U����>)���+6�E��݂zŤO��ܝ�D`�._|�h�,��`�N��%a�J�铘��ǉ�:��� A�{��Dq�ȏx����8b
l�W�O|����'(����K�A0�8��A�U3d�Ol:A��V�b�X�!��(�	<W�0�I��&XP�}����Ú9�'h�<��VwZ�yȱ �"�џh�t��7&�{p��.CZR��e'}Z5h5����O�
yi�k��>Ő��pYꀮ\XT���	u�p�q�'��[��V�Z�
�vgH&.p��{�S��xp ��0J���"���D�Ă-�̤S4r���:����r��_	��$������ �K���!@01���kͿE8�ĉ
|3�z�������'IX$0D���r=	�fY�:��d���t5�=�@a�
er���شaÖ�ip˙*�ٰ �G�{ǜaC�,������;��OJ��AOM��q����i8�h2��'��I�UFH�j�rSß<���zV�M����3i[��]����)f��~�D�3"��p�FOX���e���'�tQ���אÒ��m�9&j��C�~r�+�W�"�0�),Chh$Jo�<I�LRM���Y��Y	L����w냨F�*Հ���"�������x�>�F���O�a�E�X���fa&�`��"O�X&,I�:�^���I,l��)��e��P���?�����q�\w�Q���0�ƐF�b��
Z�E/T���%lOPMk�(�(����!�Fyp`�c��RRg�$P(�a�%��d�1��tp���T��B�Ϋ5�O�ᛣ���%�@dbb�L$f)\�"`+=��.R	bt,����/%��� ���;�yB�[�Ξ�C��E�A�xj�+P=.'����H>!�Hb6��5��W��~
� U�A/'��ա'!x�<��"OP@Ae�A�?�zg�o�D�aVMETX؃m��Tx�����d�����\�cMСY&��On1��B+l�a|r��,bVyk�nX�#�`ŠEm�\�^�@��\���9��V�[���J�*�m�C��!N��kuKM:�Ol�Q7$աhR\�2Ǚ�A�����ق�%���c�Nü?*Pk�"O9P.ΜF�����z4�@�1b����A��x����g�O?���n]���F�cD �7�^b!���h�~�ĄݷhVƘ��W��IwݨEI��A�j`V!��ɼJ)�/ۖ���.i�Hӂ^�l�R"VP8�@��n_ �la��e�,s�V��e_Z���͗l]a{b���q����	�S�T�� BPp$U��L�`�>1��"H6
$%'��-�0K�>�@� g�]�iP#=Q�*NL���}�w��b�~��ak�)�r�Ӊ�`}�c׎Y�Z\1��|����3P>�Ȗ-�~�r��d�[�}�F
�Ҽ��=E��4n���S�`��.�-Ҳ�Q���&�(�ѯ�ayBێoM��{�ܫ ��)E-���d�B�J�ߓ"�%�t�$s�މ�����R�zq��ɑW�n����'f�i㆘���X��C7gT4L�	�'���2��Ȕn�4�;���,��D���Ă&c�"~2t�ȫi���fSy�}�C�[_�<�ᇍi�	P�bƔ_�����Bg�<�5i�	y���CeJ�v�>��%�[�<i��\�.��y%cn����S�<�c,�,Do�eh�'O�uH��A	�N�<1�f�
{�("�%�;��h3@�H�<�B��!T`�p$��#Q��a���F�<��[���q���j�$P1�B�G�<�"�Y�n�^�!C�A�@Ú-!�D�<��X	��G�=[An($d�B�<i��3�l��BI28������g�<�E�n}�d�e%����ScNZ�<�櫐�5y��+�|lp�!D[�<�$�.~�Q:�l������l�<Q5ΐ*=_��� !�,�XZ��Zl�<��ˆwՊ0��nJ���<�#�E�<�C��v]��d�"0L��i�(�[�<�i�+X8�#���mgX��gGT�<�Ń�_�T���V5|��YV�<q�۸��Mjr��]dd%� hDW�<1v'N2%���ChB0Rn͈Gm�I�<	&F�$v����<���i�<����k�Pq�FǺ�5�B�i�<14)A�B���N
�v�yЭMk�<!�GM�>ҵ�1�Ҋ@bL�lRy�<�3��.`BmQ���pB<2��H�<i"�Kv�ޭ��i�#d�%�gF�H�<yk��T�"�P�<|�C2��F�<Y���@��b)<4섻�J��<��*)�u˦�ՠv�~h�fl�x�<A�����l�D�M)�pCeGz�<���b��1�t�3c�����r�<��/
,3EL���)�*��hg�MJ�<a��6��Ti6���\�FH�h�<9Q��=|v 9�H�
4�`ːD�_�<�t��1w���3�ØO��1V�<)a�ǪLET���.��i����%�N�<��*n�Sl�	(��ȧ-Ep�<2�� !>r3C���>Ȭ��Cj�o�<�BF�!��d�5���b�hB��e�<i�l�!%n����O��t�a![\�<Q��$�qd��v��1�ȇE�<�pgT�Q���
��٘^a2���L�C�<y�;.��"�cCE��f��}�<� ��򰉌�
��*Ed�$�*Las"O�����t�ܜQ�A	�qq*�;S"O��Wʄ1�ཀ�o�U���Q"O� Xah�2�܌v��YH��d"O��Q�Ո�t���+]-�t"O��G'	`�Ls��G(�d�J�"O�m!�	�f�-AS���V޴sd"O�8h�C�L| �O�X�y²"OLy`#O9�%�5o>T�b`�t"OhD8V/������:>�J�V"Ox �E����ĭ1M���r�"O�ċ���< _ܰ���T�VQ9�"OT�E(�Z������Ӽ�zV"O<�����y�  U�!hҜ�7"O���.��~��Q��@�5Úp&"O(��� y܆53d��M"l�"O����(�?���M 	~$��!�"Ov�KR�ǚUъ$�wKݥ&/�k4"O��PǓ)�^@2��W 81ʵ0�"O�&�f�X�����KݪL�a"O|KW!�p8L�����(�"Ol���+�$��Z�lW��ۑ"O4��w͙�W���C,T
g�(D�@"O�*���;�\�:6a�0%N��%"OJ�1��25n���.�m����"O�a��[��$Q�tN�ot��"O�D@�\<q�B��E�[�1 �ݺ�"Oh0�O%o�4�� ��9$��DKW"O�1Z�m�`��� f���X���"O�<���;�<�c��?�zI�6"O,�`"��rǠ�`��ފA�쁱�"OR!0���-q鎕1pBƄ|*"O|��I��i�4PKr�H)k����@"O�1P%��7�4�1�/^�i�����"O�h�,�%'��C�ᆏ(�PQ�T"O�Ai��\ +> ��a	�f��AC"O��"�G:c=R�0���P�\�"O�����(���K�o�0a	.��e"O��g� "�\��Q]P��S"Oޙ�q��6pu4��6�<~Cdm2�"Ot������K��qZ���"nM2��"O�h��"K��S ��1,%	�"O$��R#��,�D[�`b�Q"O	��C�Z���C��xw&A(�"O���p�E�?s��K册8t���x�"O~�م�Դr����Eă�l�AU"O��JEA�)0zl�E�H�OQ>qC�"O�Myq%4mQ�t���<����T"O4T#�O��H�dр#��I�h�ء"O�#3f)��"���}��|B"O p`���	=�l4 �#��+[���0"OKٳ�����R.�zhG�U/�y�K
Jhmj0�@� bkw���yR��@RBDA�D�q�!��	��y��A�]1��#i�M�A��oW�yB�7�h�����BA���� �y�s����T�0�
�bDlV7�y�L��L��w�F�7j��R�,�y�+R�5��,[rJ4+x�B�'C�!��+�����7E>v�1�!��G	Z:����Ǜ%d�Ԭ��Mgў���Oq|�D���£Z��ӶEG�A�l|Ѣ
<�y��U"�����i����RR�F4�M�cھ3<9��A0}���i�VQ��	��Q���< �"	��� �,[6�GJ߶t윸Q(Tu�F�O�X��%!`�ʕj��;,O|� K�_e���g ��`�'��$BZ�"P��ǖf%z��SJ��(�
T�҇�6/!�$̄;A�4H�j
;J+bȩB)�7L�Q�t��l͇=M��ʊ{�'An\D1��&>��2�Brn]��3�L]Y�G�-i���uTy��3�j� v
����[��)�矔;s��"2�Y��|�سg�4D�hP`ֺdvE�w�R!��ۄJ����k[����Z�e]fX���5
�g� ���4ӎD���7�O�\��F�Z�h�rp�U>_٦��LU'm-N��aJ@R\C�ɳ.eXXbw)�3��)�A��/�g�<%�"fE�u�H������^8@)֜P��L4*�6��W*Ǉ�yf��Qy2E%-�>x�vC��M[�,�(J�����6}���i�`HhѬ[=)Va�q�Re~����Ͼ݃B!��%*��D^0Z��L	D���*:�2M(f��I�o4
��P��t�*6 �r�]�d���ek�rl�q@�hR���i�b^�!��S>x2�`�
>p�����Բ��O6�rf�����d�D�A��?ia�c
�;�$�a��N7b�1�L�$
=stO&�A��ў`�l�6e�s|������E��y��G�dY���gZ�M��Ȟ"?�&��|�'��С�S&@���#cȒĮ����d�M��K���ħ5��ur�a[�[�u鴆�8�X�[��&R�5ꥀ\�Kl�1�sɕ~�`�$�����Ƶ#��M[���<�W��ݚ��w-)}Zw`<��d�lG� ���Ȫ)��:W�Wq\�!y2�q�(d�R Mo<YDCE�0�������7R�}��;G6�n���/��s�p�h��ڽ0�����
�i�ZYZ�w����̐=d�bQ�t��,c����l�
��B#�+0�R5{&	�(6pt�NӆZ3�j+Աb�ȵ��� \�0}����3�V���1n��ݑ`LL�fv�D�Ă�#�?9'�37���YC�3�	�4!���*�'E�]Ð
�d�L�n��^�I"D�6
�T�c6�'_�t�"�թ	���R��x� ��,O"x
�/�=L��	�X<�{V��+i�q�a�Љv�4�Q�i]�:���k�������i������d�!�d])	��Ƙ>b�I�Q>5���N�"���?U��#�y7�#������t)4#��]��x"Cޟ!��)ǋ�X��ɦ 
LZՂ����s��Y��m�n�4$�"}���X��T��R��ũ5a�F�䜓1���K��* (R9&b1O��������%$�!N8Ց|2dE!	JDzr� (ipݠ 㗷�LD��fK9����G�9)2��$�	1��I�ꖗj2E�F>eEў��.�hpƩ�����8Т%��jъ��k���<�!�� ��X���#]�rM
�@Ѐu��)����d��S�f���{v,�k�p��f�$;�� ���*�CbjZ���#@@}�*��'H��N�6����ɁiO6�B��Հ�(ER"@�v����	y ��9L.���ɏ� ��Xwg!����'�� ��"� ����'Ȝ��a#��䀧>��EF+��O�����9W��<���]�e ȋ�'[���W�c�jD��ĳJ�b��y~��M�Jҧ��4H��f">�N�yI�DiJ�p�<D�8�-K�ΰÂ�)W��؅;?q��R�L)�	ϓ1��d�B&V'���V�^Z���ȓwe�5 T�ϋR�̹Q�@�;W�<A�ȓt<l�33�a����'/�j��ȓW�"�1�D�q.�X9"�>� Q�ȓOTl4ҥ��b<.���"��}j\0�ȓ>�\Xwo0+0@}@�&�SVZ���C�m;4�,=,J�����4`��ȓo��,��C�B���B �Tf5���N��H�ҴP@<��LR�O��ņȓ]�D�qRl���A������ȓ2J:h���ؓN��9��
Ǿ'@��ȓc|�J�� �&�	R�Ղe�
��иqS&�ΛɊAШ��$��ȓ*��)1 ��4@��ar�u�Ȅ�PjEbg�"� !��I4]���T�Y&$U=~�R���Y�$�t���S�? B| ��N�����g������"O��j�c�,���%|�<�D�I�<�����C c��bD�[�4�$y�QmL�?!�Dߺ�����������W�r�Ʉ6kl�8�`�}�)ҧWo������L%����#e4�ȓ/��)�ĀR�,Hش���@�O�Q�Љ��)#8�
�Y�ʄp@�X�o+
ɋt(�r8���C�ta{��ˤL*���&�ޙɰ��T�OF}b���a0`�#��
QMN���O:%{֋�3
����d�ݴL᪏�
��apE<�y��v�f�� I���\��璷�~cGM6��DT��Ӄ\j޵)���Q�����C�	%V1��E@6?���34�ת@���'|
	��O�P�����I4e�M�$m�r..aP�.�183���D΍aـ!+�+������0�N�wk�]�֠�	�'R�=@��5{�!i�et�p�Z��$X�6�05iӧ���O� E� �����ta �����'g��Ƥ�6$NJl�鉅@��0�O�)Q�JM.�O�>9���R�]kHx������aH>D�����?�`�{�� m��!�g�>�� l����<i�E	/���� `*� @�}�<��e�*� $6�̳\m�T��*�t�<!�(��kF }���,f*��F�H�<��G�8)DF�IG '}^���b^K�<1ӮP
 z��Y��P$Ȧ͹�[S�<�2���f�qdS:�VU�4
�H�<�a`�DhB8 1��24K  (NC~�<�AQ�`*� U�ߨl�ʅ�PÍ{�<)�o-v��Z�B�=/���C�*�i�<��O[?\l��BVRv4����}�<���a¼E:�χ!�F�򳄔z�<�q��FK��%Y ��j���S�<��ǈE��ԅ;V$�2��RC�<I��~,����Ϝ}b*!Į�~�<�f(�\�6�sV���P�W `RB��5s��#p`��AZt �i�b�C�I'3' l�Q+؎(�Y������C�	4P����*�-lHI�s"�7n��B䉟*�@�Q�J��w���HGkI���B�	**&<��WhW�<��x	��YψB䉅hۄ4@D� v `t�E�T �B�ɭ9 A!�/�V�:({�ߐ2�lB�ɍty�����ծ	@@�r��!lrtB�͊�%�NxAT�H8B�pB䉇V���̍�
��4�WB�*:l4B�I�1�00�ì��
� ��ԆJ�X��C�	�y�h8��*#�P:�l��%@�B�ɷ[�$�{v�V=���t�խ�ZC�ɍ-�`��
>&�+�l�d6$C�	�x�)(v!�	EF(�#�b����B䉪
�������VD$�>Hu�B�	�aB��0E�1qx�vF����B�k�E�M����B�LB�B������(W��Mې���c�B䉢p�\�ҍ���BÇ��\�^C�IK888�d����_8�:C�ɔ2D*t�Z9t�Ia��C�ɏ�M��,�<]`8��.G����8�d(�$X2|l�Z"I��N�V̅ȓ!Ø� BY+�y��
��6�~���z�.|���ſ A��h���z"|�ȓ,�y���<8���u�XX�ȓ)���d�Ԓl@�30!�͇ȓ(��<[B�S!zS�9��`�/!�Ї�S�? �HǤ�'(H*�+� ���qY'"O���*�Y��(� 䆶q���۶"O\a��ӧ1���)�B�}�$��g"O��{��yŊ�ȶ#R�jD2T"O�)�@]�[B�Ő��l��);e"O�M8G�G$e�<m�D�țP� d@�"O��qv,�
|�ܴp)�s�$!��"O���1��l�<����Νsƅ&"Oj���	�Jl�!��D�[u>��@"O�ti�LO��X򤄗��H�4"O|+
�&�!����k�p�'܊�`pX%���z�K+v���H��d��P<�P$�;\�bu5�����
@�b�����(>Ь��+Jk�!�$
�O6�4e^2%�M��L�_�!�$C#1>4���"H2 �k�!�D׃`�,�1�Ç<t��/2]&!�DI�b:�$��M�)O̠�qE)ؾt�!�$Ƣ}��I�g��C��y�a	S�h!�D�0 ������?p�)�q�N�#�!�$�4|�[ÅR�BW ����^3!����=�� ϶;.T�!6cǶ>!��O�����fNN
��K'�]%`!��F�Ot)kg)�!I�Q�C!�[ |�V!L'|�48�ᡀ�AW!�d `�fm���#�:�p���;\!�D���`��^?Y)5y"ϒ>$I�O�]ڏ��)�T�f�}zs& �8Y(ׄǹ�L� #�u�Is1���~*&J(�D�)p�sD�Q�G�(b�6���i؟�9Wd��%~։����T��� ���&��aif���j�6NU��'��Ȕ����W����1����
>�������P��(O�O|�ɀA>ձŅ��u�
�p��� ;A�����(OQ?�S4��2U�)X�A�g�q�Ǽ�(Ox�}�O��Q�o<�CHL#B��'>���?�a�P�1K��x�x���)	rI��OS�hhFLO�b��Ң�� ��'�"�eo>��I
S��8W�T*T��:d��`��*	><���%��Ʉ��|y&'�b?��nW�
\�eCP�杖9cD�>aG�Z�� �"}r�(��Q�q�$��2HT��PR�<�B�/b�	1Iַ+0��"*D��SF�n���TAS� ��#�d(D�l����qK��qT��^4b��8D�<pu���81���YJ�"A.+D�< Q�S���Ň�P�8@��l'D�������*ό!�"���?��L�%D����S�4%�`��	�l����$D��b�@���h�揱�2&D�\x�ǘK�h���H.0(����$D����� ��L{P�F/(�2m@r!D�t�5�C�Oo�@H�X5��3D�l��eȹ~D0@���V����1D�d����&JJ�8ኤA �d�c<D�L3a�<yFJPQDF�ojI�p�;D��v�B(<B�d���\��&D��P
W�S*��f:@}�8(0�8D��5bW
;N�J���ʨ�x�%7D�l�AS�'C*�Pb�K�h�#	5D�\�O��Y�hdIU/W�k�D�� �-D�l!�nK�6�f�
B䀦}4T�$� D�Tjf��>�R�	�)�#R X�T@>D���u�v��@�L���i{a`<D��*�5i���0ROJ�:� %R+;D�D�!mS2o<P�hLˍf�H���>D��(�\4��]j&�
28�V�I$,<D�X�s�NxT�*����ؠ�'D�����f� r�Ƃ�M�=sV�#D�� ��K0k��ze0 ���^�~툜�q"OvAbS$��o�h8kF�Ԩ~��	�"OT��djP� kBp�E7;�X&"O�uXÍԍA��je��mF
��"Ǫ:�n�*c?�PS�$\GX��"O��0%�ܗHuL���F	g4�LS�"O6l���=�j�Sb�Q��h�"O` �b�C�%�
|#��?m�@���"O����U�3U.���BK-�xZc"O4ᑄ�ϲ^���v�<	�$��"O*��æ�6��-�"V�w�͋"O�k�A&Jb����&Ώ(����b"O�|Z(ޱF�HeI�����18�"O2��B�! �vd�B�<1Z0��"O��AB�ִ$A��2qJ�l(�L��"O0���[���� eB�,�h7"O2�(rFS.8���"�H�J���R"O8I�1$�(�t�G?,��@�p"Oh�K���%�<"��P��L�
�yR-��@��cve���XđV _��y�'
��(�9%�7d$0����yR^�bB~�Y��R�|x~�P&L�y2"��`Sg�>c	<�`l��y���+u�I�e�S-d� ����y",�(`��`��爗G:��p�K�y"Q1w�L�z��M�P8��V�y2'Y>L��iȏ�H���(@�=�yV�4@R�@[�,�4bD��y� \@ٻ5"�"3�		�%ה�y�eG�<�[��Y/�z���lV=�yR�O,����lS��:�3���y�RJ��@8�&)�X�ҥȝ�yr�����aAc�����d��y�̛T�*�qvmO<� {�$�y"H�7I`U�@G-��%���y� L�_bts��R<;x�A��F��y�bB���⁕�3( ��y���C�E�F�*��3�B�yR��]�d�@��޺����"D��y���8>yDB%E�U:���.��y�f�"�F�)WE�O�Ȱ��˾�y�
�`���: "#E�t�����yb�ߍm tp�&M�:o�x��
�y��B�44d�
#$Ř+nZ��/U(�y��JRI��	���vi�xi��ā�y��S�}��u8�f_�m�
�x"�V-�y�(ˣ/�5�p0�M�Qi�y"�"=;�H`@&<�@a�I�y��n  xZ��c�^yQA���y��N�w�ĉ&�ޱ�%F01UZM��c�����"�^+�h��Aݥ
}�`�ȓqxi��'I�������P%��@tA�Ѫ�>N����Ha  �ȓv����R�-U.�
D�uo�y�ȓ2X\�hj<8����	-�.H��:!�y���Q���!�V��}���ȓ)�� 9E�I;vk���6�8�pI��/uTirV�](�;V�ݢn��Ʌȓ٤ՋD�U$@��I7��i&��ȓh�^u�Td�iQ:�DLO4���9���τN^I���:��D�ȓ`�*Ց����~��H�]9u�C�Inp�IQM�q/fD;uq�TC䉓w�̄Ý4Bu���T-~@C�)�  ]+��3w��I���SR��4�A"OF���m��kG�ՈpA�r�p��"O�$�uEݨSʐ�F�d��qXp"O�ɨQ�P"~�a� F�\��<��"O��'��;d�)��Ć��� "O$��W�)���1�BɯG���"O6� �:O�&y�OY95����"O���]�O�m�T�?�-��"Op��dZ�m��#ܥ&��e"O�����O�N��p��Ќ9����"O��:�'v/��[���9�r"O��Y�·2���y���!	���	�"O" **1���S��jT�d"O|�p�LߺVH�q; ��p6u�S"O�)�P�1P�{7��d!te�3"O�|8��M'���q3�#6a��"O*�a�2��ʲ+R�0h�"ON�v�ŏRpHE*�J��XI7"O�Is֦�$Y�j<p�HS�"O���P�(�@�����"_��(i�"O�X�nΰP���J�"D`*R�"O������4#dR��va¤o!&�G"O�ip�Y�4�����	
�NJ��"ON�Y���,ihdEAfHR8*�#�"O�T�!���a��<_p(0"O�͡��G�}���qV����!��"Or}�v
�a̖����U�#���J�"O�)�F��m\`�$�[�p�(9��"O����0n��r�J��r"On��4���v��+�!o�f}��"O�"��ʠ669�EJ#|aJ!
�"O�ip�D҈X`�hX,Y�\�9�"O�qѦ�#x� ��G.?�:�"O�5҅#"����W�φB��!(v"O�(@&K�0�	�#P�~�"�"OB���lH�kvN��r�*�ڭ�"O��)֦�4tyZ����.B�H���"O�$��a�d�J�S`'F)DsF���"O\��"PY"X�v��4�*`�"Oʭ⑍�%mS8��eKԋ�VH�"O�E� L'"�fH`Uh�3k҅�"O�@!�Z�O�N�rt�L#ꪘ!�"O�}�`Q&�ݪ�#� t�|T�"O6��� �([u�IQD��r���Qs"O�P��&�j����ծJKF��"O�!��-��)3����N;x�"Oƹ�S`�v.��0�̽9�6)B&"OH1B�"��kb����A3�"��'"O�d�b,��1ʨ���jY?,�FE	�"Ou��C-b�L�C��	6�� 0v"O(� &oE��hb�Ĉ'E�p<jR"O�S�J4`��ӣ͝sd�QP0"O�U��N�9��A���5��p �"O�A8���7x�zq�	Ӎb�4��"O����E^3o<)`r(�Y�r�9D"O�L[���Di
����Z$�8�KW"O�T��E�|�e����V"O���&��?�x�qb�T��z!Q"O0:��Ņd�Xy bI*�d���"Op��'�؍�傑�I�$Ϟ	�5"OzB3��#j\����u���"O���Ta�60����2��y��y#7"Oh�� S��<Q�n��4�|2�"Oژ[�*�v��e ��{j��S"O� )�t��5����H}jZ�*e"O8���m	)����@��/]p�bb"O�
f%�K�8�En[�U��[�"OJ��U曰	b6�q�� V׶e�"O�b���u����8<�\%�!"O� ���(-<�{��8�B�H�"O��)���*`r1�Q�:Ɔ��E"Of�b ��/$��*$Ǎ~��A�Q"Ot-i�o�(H���W0mP�IQ"O ��/���j��0%��J�xI��"O�P�J�t��4k�C�Yaz��"O0�1�8�J���@M�� �"O�-��ƈ�^�P���g� :�"O\�P�,]�]�Ea��=x�*pJ#"Oԕ��׈#,zaxG�^b��t"OP���@oܘ��'�1![��"O�y2T�Y��!A�õ9Hvp�&"OlԸ'K�'�
=�a�N9��;�"OB��f�9Z�z�=|MI�"O�A���;D
�H`ꑾM[z��A"O
8[aC
�]�F0I0 ��
H�U�"Otq0�aj`�P��P<Z����"O�𖉚0��<���a:Fp�!"Od0h���)i͂��臊$��Y�"O"Ab2]��0�e�����*O� fD�� ����B��	�'��m���nm�͌;��	�'i�@�wb��pI~-Z0�V�I�Z���'��@2c�?gv|�J7�:OQ~�A�'��<���[<�I�J�7T��)�'W��LѨ9��!8�i�=4�p�	�':���WǙR,T����15��h	�'�p�V'�	��ku%��u�xE��'�v�s�kE&[�6Cf(�1<e��1�'֔ �O$Ema5g��0��2�'�V�k�X=A���%D�*���b�'{>Eb �T!�1y0��5�t2�'/��+֧1�$ @P*��N���'j�Њ��=�V=��������'E�p�����p�Jp���� ��'���9
]&��!k��h�'��%�  ��