MPQ    �    h�  h                                                                                 	lC=������K�9�1gbB�wv*�+*�J�0*�\ژrs̈́��i;��
i��x��Xp0�Z��0IE0��o1�\rD��e�ɠy��XZ�!�˔�#Y��5��4��Hzh^�L䎄�Ozs�?r�)D:<�V�Aw6�w.�3U7�9���f4����!^7�N1V6�J�
��S�p��p��5�~R䔏H��O�g1��A�4�S+ o�r,L@���տ&_�2��vVA�#�P��UDf�P	(���`�#�����v?/�٠\�p��32>���-�� �"� ���/�{�0i_3Ed��W�X~7�֠�fn��t0�I�������2ί�ZC�@dI��/e'�5�,y�̃������K��u#q7g�HE:tg�����؍DҬ�O�.�#!�0g���`TFa�Do�{�`��X���:͍�( �<�~/����J���g�N\L���a��"��)�iRf���'$��O3�}�ת�F]i+����h�:e�R=�HA��S��1���d~������`��Cɉ�{����t�2r�������I)��j[�����pݨp/�*w��45���O0.�C�^�P��6�/��ա+�������Vh;�E&�C@)n{�ʡЌ��J�L ��J���b��?����s��s\�8�΀�75XߎZ�b��y����qYv6B3��-�k��Fd�#�_8��.��l
�u���oFO!�yT��+��$ei"�A�:�Ϙ|�p,o���K/�y���Xl�0���2�G��IL��������|5�,oh{ ���<7�U��fD>���YU+=zQv�m]}k��1���P�f�TK�G��#cq�r��/0�#�a��
<4ƽ��aYY|�hK��Q��~3�d@]�w��@�09�hMD�Wt�Æ���)���E�h��F��Һ�J�)�,������F>JE#��7��-�{�se���15�@�੾�oVB��G���6�_��#�#�3�$LW������<���Ta���p�Ҽ�̰�v{��B���"(\�!�j�����omri8	ݺ<E����f.Y}w�8��c>dп'Ԏ��:�QE$$0I��J٪�b�"ک�H'ʂ򻘚��ܔ���Xc�.~���LZ�Ñ-��#��K�E�Ŷ᪥���c@n%��x��2��;s���B�f���w�����~��C�!I��t�5\է�ZN�r
k��x��P�����ҙ)	�m�h�o�j�`����]�^F�Fѽޞ��4����o�>�\S|��H���V�Љ�ط���4j�2J}J5�X��@��\I[�l�pV�h��@�-�B�����B�^
���^��醶�s�x>����ɎG�+__�)Tۡ��67.���a'�d}0���w
��"hUmd&��W�{�3B#�Okk@ـb���#V�m#�iD� x�E�@�.��=PP�g�AE;���A,�,`����9��~U��K����ft���;<�X(/+y��Z6 �����_����  aA2#xPA�a��fC�(jT����5��`��,z_k\�0��)��M'0-4,�X���	5��/zZ�9��I�!�~2%�7�d��ȧ��Z$k}���(�2(��u��&�>�ZZ �Ws�Q��~���,�ܬ[�4�*q�M4������[����Y�{�0�'��ė��me��M


9�6�㠴y��\�U>�f�%�: ��u~���L�ص��KX�~��v�����B�yN���&l��lʥ�j�
o����ĭ�[�M���!b�����>�x�Yz�>	-��+���k��V�	�/d��_#��(��8N6�`K��'f�߂�A޳���&D��BBZ��1�cE現��k�u;�!4�x�c�P�;&Rjdg��(�9q?�4�.ds�Ǝ99�!��9�W��)&(�Dd�z_�7-�>�(q���#h�\uGy̿2A��t!	�g76:CA x�01aP�(�k**e\�V�yO�w��PP ���c�`c�5Ӷc�/��?�:�$<4�E�`/>-�}I��e��y�0����A,
���L�C?�ߋ���jG>�(β� 8f��ث� �Qm&s`����CD�vd&�8����;}P�GW�UJ%�@Xl����xMj!~�=_ؠ���`:H���$��?A���Bf� �0�l�k��Wa��Xa)���8��۶?��N����-�����$��x���' D�E;�̪�L�	ڠ��#���MO��cs���Y���^�,�1��I�ɥ���_��y�e�����B��y�CQ5&Z��X��[]>`�%-_���)ĭ����(w�#e��,7|��zhŒ���h
[�j`������+��,���y֔=�������+�fOJ������UU3�Տ]�n^�3�;S�S#v�J�����thiT�{R�%uj�>T�N�U���{�0�������`;��ba�uۧ�4m����>cZ��o ��$���g��6�ft��̤|N����da�6%�,��*�sB:��<9�w�i�S`�â18!`���8��I:Q���_�<�z�Θ������jp��8�K�#?�7�T=|Lo����Zz&lf?Y�<u ��c0��)�\2�Oe\+,/�zx�8!xo�՘I?-�R1�a�~�p�`��҆�mPH�׻ ��5�p�kq$�(|^Gt���v1��'Mҁ�������w+40�'ku �R�:=K?n�Q�p�Hx��M�9��H�����^L�� ��䓽hO3�����T��E�k�z	Δ�%�Q�������:<�"��654����ۣ�*(��|��� ��P�^uPw|� �̞a�6��?��k��&��%��L�]�x!�,8�����r��D�����]@�?�բ�l��C��ק$X���S}}����͘3IÚ`�M[�>�����v>����Э�CO}�T�n�n��6��P
��ι�le�w,
d9�4b��Vz�0p�Y��x��4���=��ځp���rx�c%nm��O>��N�ެ�p��G�]$�wĻDF=����r�1e�^'�D�����ig�<f].:ǵ�RS�4�w~G�QVc�C��R�;pBv=H5�&J�Js�����Śݨ?�u&�/��7�߀�I� \QO<�s���\ʌ����6�"�i�o�cKW��%�g*̑l��D_2x�;��ߊ�ݸH�B^ ��`"�r�ի��qClM�x���!Xi���X�"��}�'�]���4��=�K8)w��A@��]eph�ׅ[�n�U��MD���7����ebH� �׉�V/����^�֌I�J�X��#�}�"n�8�0E �����Co
Ί`=~sd�&�*��o�z5on��EX�N����ww�Ƹ몪�:���Oέ����'�Y�	jj!Wή0�m�፫F��W���{ǯS�����O��c�2<��Ⱦ��^��݋�i��6	��Oe�>��"|þ��^F�й�����1�gM�]Dd���Su2�M�
������S�� �k~����Qb�.ݖ�w���u��U!t�1r&�܊��̄�l���*��Q�+>��E]߂��D5��ъ$�૾.^�?����Ҹ�o�+�iA��eVC��GD���&"nv��+�˽�n3LO�J��b��O��ɗ<�s���	����kX�5#Z����L�0'ݸg6=��ΈD~�\��ֵ�_��S.��lE�ėݴFJ<�yz�����$��"b�:��a|(�o*dK*���:��X'RY0��2W���$'���.��u(�-���?th6�u��k7c���DKϜX��&��Q���m����oM�%���bT�4/G8��#^�;r�̗0�|%�
��6���Y��Fh�N�L�Y~��@,�$����C��Y"t!m��	��)0g1ERpU�a���5���[,�y�Y����HJ��KC�N�Hlb��)���21R��@_`޾�4V�m�͘�,v���^m��B��nNPL�u���ߜ������޸�M�G§�qZ(������˧"_P���ڸ]U���zmMG�	TE��Ԗ|��.�Ѕ��cY����h׎���̌�c$�t��� P��#G�c��m`�������kϲ��)�?�%�!�~f���q�;E�����_��heVn ����~���;�H)�r}If�4^��q����~���|H�/{B\��vZ���r�ҴMH���Z~�}�@��SA�(~�hߜ�j��L;~���h����F�S���&��u�� oJ5>_��|�~�Ԕ�3V��#��Xw���Y4�r2�q>JG��1�,u�[�="��Oh��@�BA���k
��O�����:�(J�x�:t���G*(�:6FT����%�.���a��I}�z"â
�҄"C�Yda�Wu�q3=������@�8:������H�i�3x3
��;�}�_�wP5��\�h�{���,T�?�~�j	(B92\UU���Ɗ��<���}�x<��/�s���Z��GV�����5s����YAma�Pܗ��>{f�x(%8F��E��"�K��5\�&�$}t�*�-Ǣ��s���>���h[�,B�\���2��o�����4���x}v��cN�(�#���@�>� G�,sn���RB���q���24��ŶH��FK3Aד�(���x�����::w��3����
w� �񓡠�k�}�UU���`0m FE�~���4'�p��Ks�B��!�v�i��=T8�5}�t����+%����l�m�j,�w�^����Lŷ��C�s��u�̠�y�x�|z-Uw-�7�f����V{�C�j���g�#�d�$'N��������D�f��k��d��L�D��]B��Z�����Y�"k��l�|��x�@UP�7R�[�w�g�t3[�Ϫ�._������~2�TcWW�:&~dH˼ҡn>䇼qS�"��Zkw���Y�2�t\�zg��C<�%��c�P��(&�*�=a�1�]y�����K�W�P��`���у/)!g�O0<o�Ô��y(00I>ex#j�K���c��
��L"�}?S �-�j��(��n S\�m�h���OQ�*D`y���>C	v�l8hHf�V^IL��0�U�O�l,�?�s�!�F=��(���ۉ��$�����{/�B�'� ��h؇���<�ȍ�B�)ν;8Z���:72N6x��*�����p
��Sa��b7�De}\���e����į���z�[~Z�t���Ž��l�'�蝽؄���0����e��i�ՔC��>2&������[x�����y�~p���+����#��~p��u�	|�#z�%��;Oԣf��D����������	Ƙ��2+=m�f�11�3z7fJl��;O��u�{3:͏؟k^��Ĝv�����uv�7��]1��/�BT�wRs�j�����<���6{���M�����`V�b�C�P�	�o�9�,�]>^ݜ���r���H��:g��6�it�%�?wN�
��DrR��ݗ,�x*�B	/�w׉wOϙS[�ʢ�p`�-8�>�:̿��:��,!�-�+z�.�aIpQ~��fQ(?`�)/�BL�G'���J&gY3��u�T���n�>��m�\mϠO Ə+'�z��Y8�\R$�>(�- aI�p6r��d� R�H�=� �&��yO$P`�|�����1*ԤM�|6����R���RF4k�H'�R5���R"u����l����XR�(zr9Y�HG6��ɪ�^�] M�ߓؐ���5�̸���}�Tb���f/L	)%�%g킴�Ų���*�q6��y�����*y��7�N��i�˥u+h���� `�+��g+6V���֗�k���g2��'�bԳ8=,Ө��nm�/V��H?�/1��������~�Y�B�i��y�ع��q�'�NV�۽�M6�}��$��x�v94 a�hb�Cj�~���Ln�Ϭq(:L����Ee�>���2
:dTY`bz/�zkxռ�1��m���2��>�i��C%p�r�8�%I`�����Щ&:N}����W���?�w?�F��8�7������^"K�U�)�$�W<��9:B��R.n��⩇�A�c�����Sp�]HP�GJ���c�'� 
��R8&�Y̾�쑀�*I��CO���h�\b�UA�6��it��k��ףz�*��l؀�_ͤS;�a��$��HO�- ��%";�]Ն��q~���>�㚖a�1XNX�� k�'7����4�%H��:�rC�A���] 1t��]����T�(D��7�-/�b�r �#<�q���j�ҭ��I��XT�1�x��n8��0 �O������e���Ydj��%f6�3�5*���7�t��P�ڦ�<�p�tb�,�:*ʒ�
�u�vgҢ�υ�`�!���0��=���~F���>�{�}�N��� 䞺�< h����� �<�Ӝ��4���\���,�y�9�Jùh�����tK��T��5P]�+�'����׆Hy[���{'S����>�~�$ ��`��˔����?{�U��t�,8r�sǊtA�̿r������S��O�d��l��`c�*{�5b�[��8��FZ�^�N���5�E)_+�Z���;V4���c��y-snq�R���x�w��L6+�J�=NbgJP�Cӗ��s����M��`��X��ZzK1��/�k\����68�w�㳰��@�g1_.�U.���l�[��2%�FEwpy�hT����$���"���:bO{|c�^o��K%�#���{X��u0�xh2�>���!����1���.��/Ih������7���lGMD����J�!U�Q,�m�j����:�e��T��^G��#Y�rD�0l'L�n
2��Z�%Y�J�h����G	~�@Ӵĳ"X0�2�{g���t�6,��,)��E���|��Ұ�F�o�T,'d�������J����|��cv���ʬ1�E=@��ʾ۪�V�_��
��Gk��U�����(����L����=���OƆ���D��ca6���H�4����"��0��[͸8(��	ۑm(E�	S�{��w{�.D4�q6ct�ٿ���.��ǭW$f����x��`�������~I���$����
;.�M�ʫ$r���ɸ9[��1��J�E��l� :����n�.�Ȩ�;��ԗ��cfg�ä�V��F�.~�z��g���s\L�Zy|r��E��8~��R�x�[�O����wh��jՊ~���cȔ�F�	��T�u��Ң�0�o�p>:��|���/��V�ss�V���DG�4�82@�J�YŌC�ǭ[ԉ��&�jh�N@�)LB�K��l���"Ǡ-��{�*��@�x����*�ZG�D��2TQ�� 4m.�c�a��}�i�=�5
x:t"�5d��kWO�38T���@O�s���#i�[x���6ti��T�PƗ��w�>����e,���<vk�9l�yU����/�װ�X(<2�D/aε��fZ�z#���_��M����A��Pw�����f�p�(�;z�����|�e��
��\2��!)N"-�1c��j���gқ��Р��ç�^�2�)h����݅�P��}Q���͛((����z�>@-� �s)���t0��i�"P�4#���Cb��z�ДCﵒO����F��u�j�Ǚ����
҈�ȬN���}'���U�΂��� ��2~�4�!��+�xK��m�t�"v�`�x��4Hǎo�)�HQ>�}��l V�j��l�9P?�#���pؓ����/w����x���z���-�	�ɡ`�ء}�Vvݚ���0�]N�#�"�|�AN�][���P�L��f�M���
o��GD�6B�nZ�u������W�k�y��׶.xh=�PD�R`sSR薡�k�jԲ.Z��D�����o�DW�S�&���d<5K�m6�>߯�q��W��mE�)�og2�N�t��Egm�C7插�qPR2(AB�* 62�NyŇ�;��F\���>�`ٿ����*/�dz���<�뵔���#��Im�e3���fƞ��>
btcL]�K?�@�ӁUj���(D� nr��kQ���SQ�N�`4��9bhv�8#	�q_ �p��V �lǼ<�nN!48�=�aA�C�R�V�0��}�$+�Swr��v�JB|� >��آl�ڷ����L')	8�l�5�$N���u�.��L�����.^읇�D �5�� j�B���(^���1�O�� ��B��"��Cs��?�I��ȴ����em��7<[�˧�9�*&�����[�$�ڠ�Y&��#�OA�}����ٛ��0:�|�lz^W��Ҝ����ǠGˣ�^+�qB|�I<��$��o�=H���l�����fE�"��в�0��30~-�Sg�^�ZF��W��@v�Dϩ�݌��T
��R�*�j]�ܬ���A#{��}ʨ��[b�`q�bW�r+՛�����[�>Y���%奘�5���7g�O-6�J�tGO��ڑ�N�x߁������,��*��B�k�����w�TLSV΢��u`u��8�:G�!��6����ȼ�u���pm2�U?�*�
��L�u�3�R&b�*Y�y\uv���!&���\��0O��+"C�z.��8�a�#�?^��/Pa>3Mpѣ���v�[V�H��N�6��+���T�<$�U^|�`c��I1�BMH�y�����WL�-�4���'TZ���OR}�-�jq���>Yv��9���H⨡��p`^� �>�����$��s��8��T�tq�a�	��&%"���-��}G��ؐ��W��Vf��;(*Ծ��D6��<9�F��uy � �cÞ���6��%��iXk��:��^��D7��o�,n���`�ኇ%��͌J%f�5z���~�����6M3��,���i�p�V�M���W9V�mv4��h�K�#�8C��(�J�/ne������ �����������doTb��_zF���ϔ`��7H��PFڙm��n�,p� rnܐ%$s������D\kNx�`�&������Z
Tw�x�FИ@�r^��g��^�����B�߄�<�)m:��R	zW��f���M�c�!�],p��AHk:�J�3R�>�m�;��u�R&ģ5��u$�_�,�6ԝO2~OCM$\@�7��"f6�,�i����٪�����u*�bl&,_h�;�A;�|�H
�! ��"�o�a�'q����LU�������X	���x.'�����}m4ᦌ�]�m��A��]���VK�d�?��rDAj=7Q���H�b�c\ d�r������2S����I?�XX�}W�s��n�/(0�ͧ��v�9r?�@����d��� =�%��5�Q��R���D-�ځ/�w��BCd���:��B���!�)�����w�!͒�08����G�Fr��u�~{��.�ɐ��˲R�ٷ2<�ľ�O��[T~�@��j%�,j\�d	$����:!�ôk���/�d��x>�]>�]�D�b���JU�CG�Y���6`�S�oW�a�<~^糼�~�d�D���Tɚƺ��
t�gGr��O����D��;�з�ꪺ�����{�+��d5=�� m����^�}N�G�X� �+�k9�^V�����-�Tnl� ����2�LQ'�J�.bB�@�H�їD?�s�J��I�����X0��Z����"���u�B�63���>C��V�:e_��.�|\l��u�͌gF@��y0#�\�=$�@�"j:=��|�R�oU��K �B��iX�S�0� �2M����<ˁT�)��nN�復=@�h���� r�7Y�GD�aĜ��cQ�=�m���"L��|s@YT�,BGn�\#T��r�y�0'YA�צ
�y��5�?Y
�-h,��B[>~DD@�qA�=�DW���A��,�tW 3���)� E��ԗ���+���J�,b�F�I����2JVyk�Od�~�(�\����V1��*@��o��]�VSrWxh��b���Я������䴣L(�T��cMB�
������Cgg�]��Ѐ����b��=�"[�R�D�S��)�mc/	���T�r�v.jׂ�ipWc����{b�w�����$,,��W+ٻ\k�S΄�
v�c	��x��E*(��{�I�ۨQ��o�0�X��y�Ev�/�[4���n�����c!O;�V�hR
fB�9�(\���:>~�B�2�<ͥ��\&��Z�>�r�i��H��!jn�s�2Ҫr���<hWj|���1��/n�F��=ޯ14�e4��o@��>]R|V�'��oWV�����v��E4�{�2���J��ӌIt�b�[��⪁�&hPt�@X�B5�s���_��IDv.W��Vwxo���E�,G ����T�o��b�.�e�a8,�}a�0X�0
���"�Yd�D�W��33!�`P"@
��b��m���(Zi�k�xi�H�1��LP�dÒs�	B��2h,�8����9���9ǖ�U˒������2@��3��<mR�/������ZGh_������+�ϥ��A�=P���+fT��(�_2��[S����ƽ�Z�4\�����^�-=�t�����z�=�v:.5oU�*��}26� �J������ˁ9},�>�l(�����l>��A �E�sDR��񉞰8��]��4��׶>CE�����V�^6 �ʭ�����찄rߵ#�����
-x��g)����s\xU��X�֐n |�%~��e�;^��d�K�
a��yv�鎴����z�j�������8��l^�j"�M��A�^���e����+���AQ_xӃz#�w-z/I��Af�<�Vq��@��Uq#q�F�N�.v������f�4�R���~D��&B���Zo�ߜ�W��6&k�+�2�Nx#Z�P7��R۪k-���o�7.U��Ɵ.p�R������W�&��!dwB߼�>���q	���T�C����Լ2�ˑt��Dg5�C2���A(ZP�((\�~*�N���*�y �J���A:���`���$�/�y��ԗ<��1��b�IȮ�e�����Y�}
=�uL��?��?��*jX�n(�n� ���cef��Q�`��9�4�vu!�8��o���D?����e'[Νlb��iJ!��`=��g�^�G�ш����$f>�)�q�BBw�~ ���ؽc��2�<�uv�)Dh�8�yڶ0W�N�X0 �/^�f5�	�f����D�L�ƽ�*�]Q:�i�C+��Q?պ*���;�!�$)��D�h���'������
L�eH�#ry3�4�&k�X��[��c���ӆ4�4�^.^�S^�{��4�����|0�z٨*����w�;k<�����̸İ~�?�ϊ�K<=#Қ٧9��iwXf@���qM��[u3K����N�^g1���	H�$��v}qq��tťT%Ri]�j8d9���ߟ��{����yG�E�`�Ab��^��e�b+�>TCր�U����g�6�"_t�"��u̫N�����T�g��,"�*�"B��s�w���SQn͢BA``0�8�o:�\�����+߂�c��p%Ǯ-�p�{%���?V���g�L w��m�&]�zY�G�u1h�'w�5fU\㭔O6s�+��z��i8R�(>�s��b��]�ay=�pl���N���z'HA}��Q.u��/�:$�j|/?��n�1�R�M���3��H-m�0M4��l'����R�I|0Y袙��yf�޹
9�YH};aƿV^]�� �?�A������N��s��T�r��\q�	ߥ&%݄�H)(����ʳ��m�����̷�*/� 譫��{1����u� -	 �7���Ճ6�8�L[�k�Ͱ�]������)��,	]��rw���:����e9��F�f�B��y�x����������瘄���b
M��+钦�����v/d/�CV��g�C�lz��#�n@�����&�o@�|ȹ�ը%fd��bp �z!h��
�I"ϋ�����j�)u�pt�r韉%���� ���߱�Ns���!��x�?u�w5��F�v؄��p�G�^ӌ�?���C{<���:8bjR��(��"y�c���c��ps��H��bJ	�3�⃙vH��`�&���H�����Q@`O�m_,2\{[��$g6�a�i*�F��
�e8��*�	�lN�_^P;�AS��{�HŢ9 U�"1�,�<�q�|O�I$$�Y2�շX�#,�6��'-o1��]D4Q�Y���hO�AQE�]���(n�����-D|PI7�hH��LbY�� -���
�`�߭gΧIz��X����n�n��N0v䣣#|���#���/�Cd�Q��4����5��B�mp�¿)��\�����1�뛐{:�������D�*ҘR ����!��0�NF��ԙF��0�a{]h�D#k�������<V�%�קY�c�EМ����G�?�K��	8��Pï��om����������f�]�J����,$媆>5��6���S�ޯ��~9�׼�Z��얛B����z�ˠ�t�^r����*=�5�6��]ݛ�;���l�\*���ύ� n�5;��;�B�|�^�����;���,+���|c�V��=���쯚ng�J�<2s���LlC�J�\{bH!���×��s�/¤6��ֶ(XK�yZp 1c&��&���6.3�Ι�u���',A_$�].wa�l�;3�h�F;M�y�����$��"���:O�|���o��K>�Ko�XX�0�u2ȵ��w����F��� ��pshg/[�;%�7��Q"�tD���)�w��Q��mI�E�=�����,�T7��G		�#OM"r��P0���`�
(&P��)YE�_h��7�=ͺ~��N@IN��X ��N���(K
�9t�)���q)A�hE�GsԲ@�Ҧs�%�,��=*�����J��+tB%�����~�s$11�L@0�̾�0�V��j3�8�}�*�K�x���n���L��x��Y��ŷ<�/�����Y�8<�o��RY��Φ�"p��c@�n�����mޠL	����Ḗm�^.Ŋq�$�c�|��5�R��=�[$����V��;������딂���S#x܀9�σr�����6�����y�K��w�tEQ��N:�9*in�V��;�ė��<f���c�;�|�~֢ ��
�`�A\ApfZ$�rv����x֧��z�n����j�Y�Fh0�Tj�k�ݢ�l�����F��]�
�R� t)-o�G�>�G2|���e}�V���������4�ޅ26e�J�er���8�~&[ʁ��Âh�d@�<BK�N΂�J�Ӡc-0q���9��x*��`�FG��˙|T�~��V�.��a��9}cbsϓ
ni�"��d�WF��3.��ܴ@��rX`���j�i0��x��,��p��P<�Uím��F'��,�"�O;��P�9"yuU����x���8<��/����9/Z�u�������>�lK�A܅P�h&��)}f��\(V�n��rƘq:KP\P��������-��*�Ėe����Q�F������2�&��P�G��v�F6�}�,U(^�ߦ�N`>�� x*�s_�H�j�O��'3ܘ�!4Y���9���W�
r�T�y�ҒE����Z���Y��P�.����
���"$�� R���U�8_�q= ��~��mEvaء�	K�G�jc�v����Rj��e&�������l6��j����e�ęϺ����f�0L���[x5�z�X
-Uu*�Cp�׮]Vl5��<~��{�#1��r�N�A�L��䂟 f�;����*�}�xD��wB���ZJ��O�z�*5�k��)���Nxޖ�PR��RV�Vš%:g���3.P'.��j-�vT��@�W�x�&���d�o�����>�_!qdc"��e�]	e¾2�h�t*xg�tRC-,�����Pȹc(wL*�8��ry;��q�F<8��a��`Oq��"�9/�Ke����< h�����+0I#�
e��T��|��Ի
�L�>�?$"ɉj�˒(��u ��m�~���clQY��`J���/ �v�_u8����������Y��=]l�I?�d5�!��=Kkr�yݤ�L8�⊛K$��8��$�l��B҄q ��+��z�ڭ�H�P�-)��8+�_�+�NGV��ʿ�41���zK��ߟ��%D6�Ƹ����^��4�^����D�#�v/��='r�2��}Yص��Y���'oe#!)�hD���/&�n�DY�[Ɋʷ��Xę� w,W�g�яRX��Y|K�wzT����w�T;��֮�̬��'OͰ�� �Z1W�e�=�m�� �&�f;��L3���HH3ff&�IV�^B(�'�����>vx���n�\�`��T@|�R䯵j��:t��w�{��;�^����G`���bM��NP� NQ��`>O&���I̘1�\�g� �6}Rt��'<N�:�UZf�"�(,=�&*|(�B��*�(r�w ��SL�Ȣ���`븯8�/�:=ۀ��Kq�f葘���ki��r�p����'?ѝ��`�L[$-�i	&X�YD6�u�!�Bh_�A��\��O�y;+סz���8˃Y�75��ž��a�g�pg������H�Lֻl�t!�
�
�H$��|�����ދ1;��M�,l�N����":��Ը4M'����vR3�7��6b�4�"��	O9
d'H��ƺ\�^�M� ~�)�)�4�xž]IL�� _T3�}�WB�	:��%��p�c�e�sԢʎ�7"���JG���S=*����h2��*�Q�<�u���hu� 1+���<�6g4�mk�o��I��Q�d>�,�d �㤆�@J0�y�0��m,�+�C�AH��/�Y��n��7�.����M��?�Le�M����3��Q��v*,!�ЙC�vt�@q�n�-�"�k�w���Ov��ccbd�ؓb똘z��E�!��,.�����O�-��=hpT�rd�n%���;7��z'�Nn���iר3Q>���w���F�t �谘ܝ'�^Ǉ�f�U�U"<�uL:��dR��:�c�	���c�(��yp.]VH�\\J��a��5j������&������ը��l̊O(}��*0\�5��&F�6��bi����O�X�N�)�*��sl��c_��;�a�5��H��u .�e"�H��g4q/m�����D��r�X���Q�'�_:�s]k4��`���clA���]Q3��C���Z�]�WD�V�7�6��*�b��� ��k�����x�B$QI��lX%���i_�nI�01D�>���/�$����j�FdP�Z�K3۶q5[��Ĉi{�:Fr�7g���x@p�ro:;�B�;A&�_�(����u�!C׾0n�~�́�F(L�eH{3,*׿�f���&�O�<�����#im���վ��"E`�C��*R��p�êя�oХ�ڨ�k�S�Y]��d�����؆9Cvy�1S0pN�W�~�k�=o�܌����P��冤t*>~r�ϊ���p�v�q�*����`�`����5����5��v5���^�;���
߸v:+5�Q��׆V��F�3���Jwnb�С�����A�L�ZJ
4b��񤾁��z��s�4���ڊ���oXf�Z�
>q9��^�xH6)����H��B>�_�)d.Rf�l1�$���F6��y�����$�<"
$I:���|�!o��'Ki����X�#0#��2C�l��Ձ�G���IU�1�����h"�Z�V��7O&���`D7�	�Ĥ|�Q=�m�V�X��_���Tr�%G�\�#J�rU��0�x�	�
����O�Y�pehR���8_�~��9@K�s��fSޯ/�E��t�S���pM)���E>���Ϳ�!e�� c�,�nH�R+��ΌJ�/U
�T��
��N�;1>΢@˞��#�V	������
��ƀ�j���Z�GL^`u������-�J�Ϊ9�7��kF}c��.���/�"�10�����I��z& m���	�0L"5�hc. ^ ��ͅcŒ����-�D�x�k$7c��uC�q9��Ɋe�����Y2�.ףܻh���z�������j�Ɛf����8jE,`��шI�ԫ_n��?m�����;���^��f��U��ƒ��%~�"^����f�\\2�Z�)arQ���9�P�W�>�iG�`=����hK�ajrf�=���n�e�F��Y�e�Ѡ��7��o6�>�R�|�WV� �[VնJ�g�v�u
A4�aG2�K�J|���6>��[�-�7�~hƁ�@8�B�F��)/��7h��0Tl�c���x�T�{G�GZ����T����.�ɰa��}�x�_
�0�"��kdMIZW�{x3)��G@�W�-�G�r�ʹ�8ik�Ix�\_�'�Ԏ�z�P�k�ȇ�����,�,@i�������9}{SUA��2���(q����<��/2����]Z���B�u�)�e�!���G��AY�kPH����b�f
r(/�����Xz�s���\�A���x�-�����\��p�2�,����l�v��k�2������.9���
�}�kOp(�}V���>QY� 3/Lsz�����f6��ӮY4��ɶ4�鲜R-V���$-��b[�w�&O���<]����
�`��>�;tc�i�KU����Lq@ ��3~��1�Ф�\��Kߤ���c�va�ܴ)�@��`���Y��ݮ�lQ�0jDԂ� ������T�f��2���v����xP�z�-0ۛ�Rd�r��Vg�H�����±#L���Nd0������S�f�bg��(�8�7D�Bx�Z%I��r��S�k��˺��.x��Pm��R�y��ġ`|S�;�.K�3�U���]���>W�:�&o�d�C�>��>��%q�귍�e��'��l2�%AtH��g>ԤC(6��l�P���(�t*��mݝ��yvQш��7V{��v `
���=D�/�<��ڿ<[�D�g��I~�
ed�U����O��
�MKL�.?����=*j�V(u�� �tY��`̀Q�{�`����*�v+��8T/���"�5�@֜m9���l��D�_V!Et�= a̔)j��9�eZ�$�R�H���gæB-9d o
u��P�(���+*�)���8��|�&��N�5~����OSf�\�'����N8�DћƳ�����FD�y%��G�����������I����T�M�pɍ�0Q�� #%e����.g�2�*V�&!u����[�m9��M^���԰7%h�s���݉�a��|f�9zϫ��c�ԏ�qǣǃ����za��u�&���}=ى������f64���#�aU�3�
���}�^?l�b�}�Z�qvs+*�ɢD��T[�R_"dj��"�uq���x{��ʹ���j�`�b�y���r�[V���*�>J)��6�����.&��g	�6X2�t�(�̫��N߂����ם� �,X%1*�{�B�T	�c��w��4SG������`�|�8k[:�yB�f��5��N�f�Ϯ��p=����)�?L�H�y>L�X��ż&S�Y�D�u��E]y��P��g\Y�Ol��+Ѻz?��8�/�t�c�|Mř�a�p����l#bH�< ���������f$<��|e����n1�Q�My��i�u�>8��T4W}a'%1f�x#R��w����������y�9E�IH��hƵ�
^3� 9A��Dq2��w�8dT��jT����R3k	���%S�r�~/���ʚ�i�.]{x���\���*��#���EW�·�^u�k�6 �>۞���6��k	�u�S���7�ԟ��,?���������4r������������j��׮t`��-fD��]����D�Ǉ�M����b��
�v%�y���T��C֠����n���]I��Χ�rQ���Z���d���bfQgz�׋��~��We��jڪ�٘�&�p7T[r߆?%�k�v����NiQ�7Ҭ�����k�w+sFa���#�T�8( ^۞��EO�!/<�K�:.u�R�t4���<�X0�c�^��86p��H��J����ϩ ��-�F�&�A�������0�xO����I\�/q����6�+|i�օ
*�"t���%*e}l��_9��;��W���0H;�� I9�"'����qj}U�3��O��͉>X:o��l_�'#p�N}�4�һ�R�p^��AP+]t��^����u�8��D�|�7"$B��}bE ��.��>;�V����I� �X�'Z�d�(n��|0�q��Y�k���������
�d�����6��5��ģ��µ�R�3�(A�oz�t�:�����~�zƎҎA�P|�!~)�0	b/��N�F����]3{Nt�:��\���oI<����ͷb�l��(+]��皝bd��+�e���å4%�w�`���h����]�m��Zzކ4q7j�_�g��SK ���La~��o�x��5"%��Cɫ�z�A��tE٥r����z̫�K��������$���g#�̻ʂ�5��ѱɅ�$^��.�XyB�1P+P_J�rl�V� �n ���(n]0���D�c�L��SJ��Xb�Ų��+����s�Y��Z�}�L6�X�Y\Zf5a�\�Wq��6$�"�O�����]p�_�.-��ll�JĞ��F1�byA���}$8�"��j:��|OT�o&�4K�Ț��X���0>�#2���kM�d�|�����N1�h���q�s7�|���Dr�
�_��IQ��>m���s�i�� $�k�T��%G?Ь#E�=r�l�0X���)
�ݽ��nY�g?h�g�3�~U�@�g��h���6ފV���ct(����)��8E�vF��^�Ҝ����4,|g`,���Jg����޾�d�)�u1y�,@f����6VdiQ�A�����A�|�E�����L��I��� ^��;)��eYͪ�1������T��$���ؚ"&�����ø��{���gm�|7	?2�ɖc��.{Q/�,�c��Ϳ	~�$̳�/$�.j�д)��W5��tׄ����v��	�����Ϲ����	��$*�%n����@�m��E���L�oM�n�!��Ȕ�&;�ӗفFf�����+��� �~��7�C%���\w�Z�N�r,���t9���p��d� һ�Ϫ&hf^6j��{��˹�:� �qF�!2�������@RQ(o��)>�}B|�ԛ��Vз��º��06�42,R�JW�_����3Х[��V��:h�8@S��Bu����C��Ӱ��T�g�D��Yx�C���SG�����T=�j����.�+�aI��}��q�w�
dk"�~d���W|u�3$Hl�qU�@;��H��͏N�i�C�x:���"�0�&r}P�b����&y!��cY�,{1������9؝qU�{��M�9����\<lo/��1�5hZX�S��[�D�
��"1�A�x�P�Y��fe�(̊s�8��h���N����\����o�-n����B���M��e���&��Z�2G���Ʒ��I
��<��}��)�
_(�d%���[>�R
 �S�s��m�`P �Ae���4�4w�/r�����ꔯ��;풪R�*�ad߆�#�M�
>�Șys�V��|7U`"��w M�N~���J(�V�K�!�`�Fv<��d���`�[����&d�i �ll6�j��y��������ۓ�G�<�!�r��xklLz��S-a�ɍ�@�`:Vb�QL�I)H#g["h�dN?a��4]�&>f��|�c���D1�B�,�Z %ߜ�p=�`��k�ʺC<�xTp`P�ԨRL=�C����3�ֺ�.F��ưC���e*��LWx�&JՏd(*����>ˏ�q�m�����[��2c�t��zg�S�C#�R?�P>ե(�֚*Xo�xb/y����sR2�*�t�`Ţ�X�/�� �\�<�d�Q.rI�Ǌe���Ҳ�ʸ<
�+LIQM?Z���TjiR�(0K� �
����;UEQ��`�"��%>v�<<8y=�ݣ��B��w�z|Xl3W��Z�f!�=��3̯���B��@9�$�㸄�b�B�W *j��	Jڣ���t)�W8a_2�!�N�4Aa��j����e���)��qDls�Ʈ���n+;k����Rt��P����������s���>���+�l�Ki@�{>�e��#�J¥�%��&|��P�[�p������=Q���=��
�2�E�[���|��#zJ]�>`�������z�����5����>�[�=���X��:�f1���^���3�ο�?Ű^�u������Mvn�@�$�,��ֽTv�]Rڴ�jɩ������m�{~Fj���G�%`ݯbCWE�Hű�~e�3Z�>EL�֑.󘆬�AF�g1�63j(t3\��F<�N�p�����Y�,s�#*r�B\7X����wV��SB9��Sj `a`�82��:38�G��Zl�4��aQ��(�p�g���o�?ǐ�v�uLѬ�����&N`�Y�rub��x�������\�k�O�+�/z�U8������+e�t��a*�p=����ǧ�HrLn���{����$wj�| c��?1� �M4B�܄��ڹm��~ 4���'�����R�x�A�����*���o	�9�Z�HN��ư�P^n8� ��_9�n�����$-�Ti+j�MD)	��&%�������i��Dh������4۽��*@l�ޟ<�`�
�2M�ur�!ޭX grS��jK6!��}��k$	���P<�ns��ڌ�,ځO��h�������N$��5��!�����0�`��I~ʳ�j��#�g&�գ-�B�[M}��C����_v ���6���C��`�6lun����!�S��m$_����>'d�"�b�)z�����a3��t�� �#�Z/4pRt�rZ��%��f���=аr�Ndt��Z��X��v�w�rmF<� �^����Ho^	ґ���?�<B�:�.�Ru]ޔٷ#��oc�]^�tp��{H��'Jz����=��'����-&�t�Y�/�K��DO����\,J�\�:6��i;�����=+y>#*@g�l���_�c@;}D��9�H�"Z d��"��m��pq��&�k��z��(�X�D�ˇ�;'����)��4k��'Y�eAb�]�Ԍ�yv�P�$u�D-�%7�1���bj% P~u���_�ьͭ�/TI+R�X[���_W~n���0��p�tc�%��ά��fid�����]��5ј�ľ�=�0�~���c�����댖k:�p���:�Е�\�	�s�+�!��0�X��;�F��au"{i*F׵��7�:���#<'�۾�o���q���Y��x��������B�禟à�D�����`�:M��I�\]f���N"s�t��/������"� Sf��M �~�2伳7�Ї���-�����t`��r�������)���o������)��6��a���J�5��	��}5�MD�^�y���f�쩠+k���� �VeGɔ��{�.2nX��M����rL�W�J ��b��c�4�S��ŧs���µ�p��
X���Z�K􄐩�F���!�6�Ϊ������x��_�4u.� l�|��9knF,~�y�L:�H{$"u�" �X:���|�?�o�9K�X�\?PX���0YW29ذ�F蠁@���<��Z����h���ی�n7E�E�d�D�������A#Q�j`mz�d������a�\�T��G�c�#@&rS�0`���
����g�Y�~�h�f��.�X~���@z���<����e�)���t� ��z)R�E�>��c��P�&�,N������{~WJ�V,��@�ꈖ� R���1��@�3��i=V��$d>����Ѱ� ���<L������B�wv��<��ٳ�/���ɴ	����#:�ӿ��"���>�K����p��mo	z���v�^�.�d��U�Dc����!���Z���b�$m��L�'���?~�O��O�u��k�1'Y�TS���G�2�������w�E�}��G]D�
�n���u.�O�v;0�'�T|f����}�M-n~ǂ����2͑��\�?Zw��r}X���᧍��_=���Ԑ���h�K�jhg�]]X�,[ț��F�w����QVbm)�o,z�>��r|B�U�6f@V��Ɖ�v��M4'��2�x�J2箌5yΨ�[�嵪�Wh<�@nP�B�	���P,�����4�DbJa�J��x[���YFG�\Txt�']z.׭?a�q
}M�O��-
�w"eu�d�ͽW�L3�Ղ�Am@�&�c_����j�Wi� Mx�E���(���xPme��E����>��,�ۄ �x�93��U�	��hI	�"����z<Y_L/hS���NZ�]����_������aA�v�P~Y���4\f�*(�.<�S���5o�)�:�$\!���5V���-)�$�I��f���]��:��h��hq2�����q�d��ʷ!}���)"(/kL��|c>l ��4s����ۯ*��e�I�4*���*��h���:�ʒz���V�-�c윙Z�!ւ�z��
�uQ�S�	�q�~�_r�U;ǒ���� �"~��V����;�K������vik��7b;��V����]�$�l��Ij;�����Jrŷ��H��xX◡L�-�jx���z|
-�/��ب��V]���.����#����\N�����S1f�Ι�*e���DLdBn�Z� � �܏��Nk�3$����xP�+R���ꓡ�`�q��.A����e�>����=�W�!&%'*dc���t�I>�WquYC�@��@�J�2>��t��Jgt�qC����1}P��(�ˉ*��<�S
�y�w��B~�-�r��`�k��s�/���7`�<�>���:
FI4�e�9���}P�E��
�)aL�
 ?�c���j�ſ(�)B ���O�s���Q
��`n�� ��v��?8�⴫�D&+��R��GK�l�X�Us�!��=|����!-ʽ[�8�$R�6~���]M�B�J ���)���1���]0)0=38���NXT$�(����R�u~k���dDk>Ʃw���u	&R/�����=A\����'�p��]�	�
~V��꯰f���yUe���^	�� 8�&ו��u��[�/��:���%�J�aHvҞ�ѠT���o|��5z�.q�a��0wǧ92���p�8�g���눫������=���ٓT���f,���]7y���3��(��,6^���������@vieөő��T���RUgej��L���[�HR�{y���o�H��`�i�b�Thr�G���=�Ω�>@�����f�A��\��g�y76�tn�����N�~6�fb۝S�>,�%�*�LB7:��,xw��RS=���b`d8MAh:���\���7��O\�H����p��Z�֎?B�`Q]L!��:��&I�YU�bu������Ҥ�\��mO�M +	%z��
8>Y��������OY�ae��p�{U����"L�H-|���
���=�@�$���|�O����1L�5M���ܟ���4é�t�4͝&'[`�ݎ�RDs�h�����; �J��9��H���ƫ.s^�] ����z!���s������_��T���Hu�	K''%�3���N����n������$۸�*��虆X�{��­ΓuM��z/ ���16x��8bYk?�Z�I��Iϐ�d4,u@������Q^Q��Kt���⊜�Ţ�����B��䧬���8��6���"�,�MX�I�~�z�"�vD�/!����CUS���n�X=��r��h_�`Ք��d�w�b\"iz��Ǽ�d:��\�����`�R�X0pm�ur��%k�8��F�KH�N_����بdR�hw!tF.ل����n��^c!�w�"��~s<#X�:$]RPf8�ܾ��goc||S���p_Z4H���J��������bE��|� &�����#�G��0{O�k����\g����j6�u#i�3g���DX����*q�l:@�_oPk;x�̊F�AH�� ��"��ը%0q��+�����2����X�:�ˢ��'���4=in���uT�A��]�U���ˌ��xDh)7X_|m�b�%r �@�%��Ls����If�aX�8�Z�nZ�*0b���t���)�·f��d!���PM�Y�5��N��«[���*�/<I,���s:L���l��а.�҄�r�ʝ!�-N0?����H�F9��{�Y��0���\�� �<�#���G��"I:��z�&�����p��	�����AO8ÛZ9۶I��=
�UR���H�]Ajn���2��r�*-N ,N��[�S�����~��ȼ��dk>��fy�a@{�o�t{or�
E��� �!�B`����'�q��H%I�(���&5�^��'R��蟨^�HF��I��#�+���h�~V@�B��!���nSD�������L��~J{�b���o��K��s����c��5^X�G_Z\���>ԩ�;S�I��63!����y�9�4B_�.�4bl�|2��r�F'y�y��(��4$=Ү"{�:�Υ|�J�o\��K[Ě��4XDW0tIr2�#5�!���{*z��������r�hS^qۧ1r7����ʅD��Ȝ��QNF"m53b���������mzT#�AGuP#;)JrfYt0�1�9��
��|#�Y1�oh#�K�)�E~�:@5��0�xlA�@T�7^t^�_��G�)�M	Eo&*��SҒL]�8A,�������v�J�l`M��S�{_Z��W{1�v�@�]q���&V�8ȋ�ɠ�7*���y��e�L/`{��aUX�Z��y���X[¤� �g���o�Ӻ�z"�����W�ڊ���mJ�b	���:�Y�.1�m�J�c����Z����)��$&��ƒ�ق������ ���_�����l�w��C�N��������9�cG�E�<��/��n��P*��
 �;K*�ϖ�f�yx�OV��yv~�b���À�Lf�\�8�Z��Rr���y��(�܃Z�k�q�͐E6h�X8j��85�X���6۱F��v�v���7��!�o�u?>\3|}J���V���x[����4B��2"��J���pJ�i��[��0�H14h�D@��Bk�\��ő6l^���]!����8x'����G���7��T�[���+R.�Oa�R}�ߟ1
ZG�"@�d���W��j3��'N @���~�E�i}�E��i�xp�u�伎���P(����o|u�
,�!ք�����9�BnUr�-䃮��*��z��<�r}/� ��Z�,s�S�z`�3�ؖkA
��P?m��͞f�(B�nC|�^���i[75R\�5����%��-�)k�0o��� �ҽv�2�/\I����2����<K���2H�}sW� i�(ʑ˦�v�>b�� d�~s˲3�V/���"�܄-�4�7:�%����i+^ŏ��ym�1b�������߼�y�uM�
���OĠ����ڇU�Y��1� �z�~|v����؍A]K0|ڧV%!v��*�ڢ�W>�Q���jѷ��!�l�f�j�戂[�ą�[�%���ie�����wx�r�z�r�-��P��a�C�wVXe��j���Va#�7a^NN�"N�8-���-\f��[����i�Dg͌B�%�Z�<�;P��o5k��ں�>x�ɡP�\RB�:t�c�Ѱn�.<�-�f�#����} WnB& ��d�d�RX>�?�q�@9��}X4FMQ�2�t�JNg��C8z�D�P�p�(��@*���.Ҁy';��ݨ�(p���`;T9ӎ�8/��L���<��8\?��I�xe��q�i���5�
�GDL��F?�d���jYd(�(y ���$e����QEȮ`��l���v<�8�l����*�-im�:�li�e�P�!V��=7�����*�86��V$��s��X�_B>= ��i�D�ڙ��'�)kBx8��e�W�N��'׵���y����ŮP�d���D��hƤ���$����Q��Q��q���b�V�q���ekء+W���v�q��e����A��}u�ٮ&2V��0��[5׶�����{	�ą�T��+� W��?��b�|��oz@ ��O�@l��B�����2��p������F�Q:�=j����]��p �f'�^��xt��;}3Ҷ��5�'^�C�e��+a�vd2�ڇ��L��T�x?R�9�j���&)���V'{tV	��-����`Db9r7M���/J�iu>;��G�����w��gu�6�9?t�"��|��NЬB��Om�k,���*h6eB]F���w��S8��	{v`ׇ�8h��:)��7ç�RM��j fW����=�pn���#\�?�/,��LG��շ&D^�Y�/qu�H��l<�S��\
��O=Ԝ+.zPh�8���6X!���*(�a�Papsmp�z��};H����Q��f�v�!$��|6�s���b1���M��ܺ�Bگ8'�O�H4^�'�'��I�R��#���)��� ��%��9�ЩH���Ʀ�q^$�� j����)��d��t���ET�F7�Cƙ	���%����Ϩ��_n����s�_���,۳�*����T����d�(ppu(~STf� �9���6Ӎ����kZ{9��	`�$KF�P[�,��Ϭ\�O��eh���}���s��#+�E	����D�U�I�����<�8�NM3��鹨$��Ȟv��hmЅ%�C'��,�n�բ�2��ͧ�c*��U�O��d�tb�:�zh�]�1���P�����ڻ=�Р�p��rPQ;%F�z�'0���=�NZ��H�-��`��Qw���F�A��� �	�U^�֌�ҿ��A݋<>��:�R+�B�O �)3�cw���*3pD�H!Jp��`�$�����1,&��;�N����9��<FO�ef�\��?��v6�J�i񧯅;ɛs��o��*��Wlu��_
].;s!�X�Hl� ��"��Ճ��qne�P:���/��ވ�XkP�˽f�'�aW�ߜ(4x�Ō#ͼO�AШ]=������FH ɪcD��R7�}wn*b F] Ƶ��.����yS����I�T�X��5�U�}n�r06.����{�b�V\d��&��xG�j5G���� �&��ڣVu�֙亩�:�:����'���˒1���݅�e!/�0����u�F��B�{���׫�Φ�ݏ�;G<]����?��}@�Ys��A璚{y��6������Ö�6�Б���pw'�?�]Bg�ĨF+� �%��{yU��T~S���C'�~��)�I�����ɼ���r�)t�jMr�h��q�K�\�A��pR�����̮r�4R�ӂ�}�5_7S�bF����^�7,�i��b�+�r���iV/������MnN���ѷ���L�J�YPbd򕤪�͗�H`sֈ`�k�V�}�X��Z�t��(�Q"��zQ6�
�`?��4׶��f_��6.���l���o��F"��yR!W��n2$XOe"��:_��| vio�>mKA�jyX�W00��u2/����},��`��M��5�_Bh:��}7;@%iP�D#	��0���,Q�A�m����[���ab��T^^G��#6p�r��0�#T�5
�dm�W��Yl�h��l�$�~f%�@�}��DI�i��n1��t�97��$�)�qE*.��9���/��lj�,�c=1��q��Jx���� =>�����4F1*�@7�f��/�Vu���:���2粢}���F�L�J���O[oR�l�۬�99�%���g2���Y��ӵ�d"7��%��5'�f��m%�P	�^�d�T��.��|���c1+�z�&��L��d��$�Q���1E��r����ń;1i�E���sܧejϊ#�������V���pђ�6yE�uά�@��n�����i��#;f�h�J�ofdO������~�bm�T���Q�\�zmZm�r�ư�%JC�×��U����&� �uh��ej^��a�����F�����Q���7��9�o"��>7�#|�0%�l�V�z3���w�ayj4]��2�%�J�2���;��[�Ȫ�ܰh�V@�TB�LO����qhàjXO� }lx��u���G�xoT�b۬]�.�?aZT�}���c�
Վ�"�d9��WM"3���z�@lv���Uv��� ��iW;�x���<�7�P��+�40z�Y�����,,J�V���9��LU-���3R�S"�U�<ϥ/�h,���Zi��.Qf��j��>��y�AEӋP�D��׆�fv��(��Y���i�ْ����r~\W����-�ť-��U�K��\
.Ҙ�)mN��$�����2X�5��DyȚ=�ʭ��}N;f;�$(eآ����>��� ��s��2��΃�ұ�ܿ��4`�O� ����s�� �蒬L���;�dG�W��p�
O����颠�|:�U�U�pP�8�U �~w�z3�HgKKY~�ѥ@v�h:�.qJq�LD���qݚңl�.j��6L���~f��_��zn�M�"���x�%^z��-���>)P��Y:VSA�b�1�z�#��<ٯ�Nг��s�I�a�f�>%�t��$)�D�VFBdҚZ�x/�v6��1tk���T�px��P��gR���O�#�Lō��w+.7$��xሴ<��,ܦW�y&�*�d�1�����>�GQq+HO��p/O��E�2�X�t4#�g��C	�cvPo�(��*}�<�	��ybЈx�#a�(,�`�\�ө=/����eQ<G���< �7I� ePA��#t��;�h
_��L��!?+�2�Mzjz�(aGT +�Eނ�̯�Q�� `Qe���v�w�8@�.��!����I�l���K��!�ٲ=�2� ��ʳ�-�ѕ$����}�SW@B�J0 [I��_�f�F����)�g�82e���N�J� #��X�H�R�+���:9�D=�JƟ��jf��*��k�3�h�L"�����D���������\�b��q��P6ejw�ԇ{�ю��&�6Z��[P:F�x��V�~��5�~G�����VK��Mٱ|��z�1����}�{ȯ���}��1��:�f���7�̖�=Ey��	� �o�f"�U��O�M��3��2��[�^���N�Z���v_m�5����TǇ|RK,�jZ��a��~{<{o��%�	�x5�`.>b���(�ݱG�����>6u%֢u���V��g�j�6���t䵦�̷N��*�]_��#B,ĥk*�	jB��OIw'|QS3$x�d�a`��!8���:�3���݉������R�2�9��p)tN�>�?8m)<L�iI�p�&?IY�?u��.����bq��\EISO�z�+���z�!�8���$��4��a��p�u�����H�;q��m���QT�$(�|�(����^1�Me�B��'��*�P�*�4C>�'��$2R��[�r^�D(g��ŝ yV91�HK�ơZL^ %�̓�Q:�ߪ{����կ!T:��>7L	(�%?K���������٪I��Q�Lۮ?�*Q>���|���M£1yuot�r� 8���06.tn����kud`�?d����ԋr�,�[��~8�a� ���R���>���j��Vg�[ٳ����]�I^��&���Q�M�������X�"v����8�@x�CB�0���8nbr8�Ij�$�^]����
xMd,��bRs�zC7D�l�D��A��~���K��	Up��0r�Լ%!w,�b~�ЁS�NUo[棳����XCw~�F�I:�/ܤj�^�j�-�v��[H<Y�8:�R�������cr�qp�M�H(bvJ�R��;��������&�)*�j���|PZ��hyO���@8\�X´-�G6�?�iL<���������d*��8l�*�_���;n᱊��H'ÿ ���"d��^�qV�Ҁ�������9sMX&�u��S�'�\��<�4�q����Js�As�]����ʞ���#����D�U7��r��b{�� �c�I���B�(���I�?X,��P�'nY0��Ű9���f�=�)�;�dW������f�5^��'~¡���~����i�}��:U������8�z�����!j��0u���F�r��|{���&2���R�v$,<�뾹W���Wfv(�\A��.�a�+�Q��w�Ñ W��L9)�������[]�9������$g� i����Sm�S� ��Z�~[��dҢ�x7�}8��Q|�-��t���ry�ϊL0̗�f�x����#�'r���b��8&�Gb5:0�ѝZ}��^�FN��rQ�w�+�c��^��V�ҥ�Z���Q�_nI�ա^�e�OYL�JJq�%b?A��y���ps�-���I�8�X�ZRS���C��W�6�λ�Ȑ�1X�x3_��.�^�lX���
�F�y��ŕyTt$s��"q&�::N�|;�Mo���K�F0�m/X��m0�9a2���x��`��\�z��2�h�5����7��D�nD^jל����ZQ]�m� I��>R�x�#=��T��.G���#1�Fr�0D5io7�

ъ�2��Y���hY"��4~���@����x6n����1yl)t����!�)cf�E�U�T�҈1�G��,��� �lvJ�LN֒��;G�q�P��1A1e�^@�|���-V�r �x�����-;����􁋡LeU�ȭ1�o<'����ت��d�ZM?m����:�Ӱ�J"�[��oy��ƺ���m ��	+W�SE�O�.�^,���1cL�C��-��t��̟OJ$>�Φ���8o�p[H�V�8���ܚu:���41�%�,��A��X��������ђYF�Es�������:n�:�Ȁ�;��T��+�f?�5�� u�sO~������|��[\�� Z�$�r���`:§^�ރP���'q���Ah��Zj��.��޹ν��l�RF�9,�,��X �q o��>i�|�6��o\V��c�.|��%�4xш2�,JÈ���L���[�i{����hmS@��Ban�p����ܠ#RS/ �[s`x������G}�����T)����(
.���a�u�}~OBHq
P�#"��dt�W�3<����&@'N��l�����i�xix��}������*P�-��O�eW���L5,g�h��8���9DgkU�r��آ⏛��0g�<
��/9#0|�+Z�e�����`��"6��|�A�1�POja��_fѳ^(�ٮ��_�Tq9ƺ�L��j\�6�������-Z'�fN��3��s<��6� ���U_2�/�^�ȵ�b�(.})?�vGd( ?Ҧ�ʣ>xW �&�s��L�Ҟ�`	��!�4��ݶ��y���F���'Wꪾ�o�M����+0�k�,
���Ȅ�������U�uw�sR] ���~r�gt���KfV�LF,v���P�f]|�G��� ���U�l�<j�H�����4�[�`��s�2Π^3x��z��w-w�D�y���yBVN=G�@i�5#ӓ@T1JN�du�����$�Zf{+�Ͻ`�ߚoD��GBߞ�Zl�?������
k{�[����x@�sP�d"R8��*�ӡ��>�B��.2u��u��o��G[�Wd�w&��Yd�E[=>�obq�o��q�*j�_G��2ϵAto�gE�
C�S��ȸP*�[(k*�yn���y�!b�^�̀30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4�y^�*г�j���&|f~o,KN��xslЗH�S��ޣaQ(��OU8p��ӳ�ę^�|�ΡZ���%C�A�R�n�X���<���.���R��_@n^��g���+�¦���,t�_�_��t��T�(�gџ�l�0����G�KA�����tf,�8��'��J}����/rĞA�ɢ��`��F�qX�ߌ�����a����:��дd��-��q��!���7'c����~ZX�ox���\b� ���y�1Mfߖ�E2Gb.�S��^'��I�d�0�s�fz�={���|Y@�.����su@��_7ᢈ^.�)W�{p� �H�>��~νU��M�ز�����
�y�Q��]�����U�-j|@�'[vv&&�/&��΂|�S8G}(;�^f�&�<4�~]��X/�\�4�Iށέm�<�	�▴�����G������X͎0	��h�ٺ)��An�l�jǲz0��{Ո�᫶��S�� �� 9D�1A؋=��c�lR����U<��-�e�
��Im�g95K�^���(��jc��K����52�� n��e����z�1��8K|�j�|��;s|/�������`�D��K	�p+	�THˀ`�o�FRD+'��
8i��1V��05�Q��wExu��O��VGc�Y��leykD9|l��[���0^�mO��x���I�k�����T��ݺ|Eo�E0~���x�;H�WH
��i��������EC��
����v��(d�i������F�7$�z�$��Iy�,��;M=<� ;�$��qGU���n�L� �μ;,���ѧⰾ�]���t��[���1����>V`��y�J�^�}^�����e�kbt��'����ඟ>�u��>٤X^8%H
��ɭ����]�&�4�,Ԙ�r��p�$�:��$ˮ����r�� c}~9�Ǉ���c:2��|�Ll���[r˔�����٫،���,}܃�a�%"�5l�f9܃�&�%
���AO&�la	-�8��3�D�5�;;'�<���1<��rV )4���\H�i��y Z;І��ڽn���L�e�D�V;�H4]m����)�9˯բm�a����R�sd��J����p�\֢�h�E�r�A�Sނ���-F���">��_�A^vӀ���W��36���sM��H��~Cmh1)V��%��w�ɮ����Hqw�nۣ@m�7rVE0�;��h�zF�饋�U��Q���ѥ�(	�������.�.}@V�2{5��X��B4S��/
Q��T�}/B~4
O��NRjWף�ؤ{�
Yg�o}�?�����J�d#�	�r�KWܑ�\j*���4h1��D�^�d喂	�����	N�6��L=��C�1�3�vM	�XYg��X�ʖ�����ᩣ�w�г�s��\M�˹��GC�k����]���J��%�&�2��==�ժl�Q	hr��SZ������둷i������F@�r�st�%C��<�)#3j��������G����N5C�P=~�"lIZXM�|o�q�^�e8=u�&X��?�әI�t�0�k�f��*Ms��t��&���De#8!4VW�����H�!'�s$����~��v�O%lM{�Ǝ���ұ��%I�6��q^���gԻE�\Mk�*?���+6�'�!S���?-�?>2 �a����4�ǜU#>'��-,��y�n�=��0!���4����E�$3��#l]����'N?��F"/���9RGt�,N�ܪpE��s����朿8���(y�떦�u�`4�:-�W�Ƶ@�_�9�`���56zo��ĸ�B���#�G�ûDz=�ԇH�,���>��Z�@�B[4����T����G/���> ��k��UI��gl�˅� �&i���*=����hAr=y.gB)���wzW���i��6�4�	;&r�S�C�D������T�sLS�'3��P�ݞ���C7�"t���\T0�Uv��^f�P��}u�*��2A��>k���/�������_�2��f�|ex�q���(���P�� +[���}%��A�!��c0TI?c����"њ�L����y��F��w�hu���^�!�H�^�yc�2����"���O��'�d^6�*C�tp	я�j���Y�v˫h�e0���'���ە�{'�n;�` 2�z�nJ2���7R� �v�(�n�pJBT�W��V84i_~�e�,n*⪣w'd$r���l�;L���_j�dzб">�����9��e��T)l:h��d�H��������A�'�ۭ9�~�w%5���<�b	������Rq�%��6���w�� �H9�ػj
��Ơe�|�$����0��.1�0 p%qEw0���e���z�JQ[g��k����߿�4������n�H˩zMZb�� ��WG,+�+��b�����df-� ��v��X�Y��ųxb\���,�y?	2f�W9E=�.!��)�y�t���(s����~{2�|d��.���,@�0�_���I>�)]d{g� ��ͩ��I��U��ؖcL���O�����-y��j������,�U�<�5�'F�|&qY�/ѭ����1�(וGHI��h2��R�<�u]�8/.�e4�f�9l����D	��FE9<9e��ci2�;�E�s��A��A�<	�WNާf��Z�ް����*x���!{��X���;�|�)�P�>�Q㜑Eh<"�5%���1i�������d��?)��I��B�T�J,�[+�ؽ�����u���5��">�X_�Jt�d� M�\re�#V}��@�ŕ�Ηgcќ]-��l��(p�7q�2�(Ѥ�!I��P6]R(jr����_��1q/p�� �CC�]��a�KՖLa�3����&��_../��iX��y��_�K��R�Zܤ��\�$N%��f�X>��}�����I[ʲ����#H%x�3s�d˟�i��ƀF��/��)<eħ��c���1-�Vy���4��Q��������k����G��7���}(�Lfsw����S�4���5⫒�*N�G�N����f��Kl�xLK�AQ#���ca��߳�	8�u9lY.�R[o���0Κ�V��Z��N�RAN����@Ck4��0ʍ��;R�-�_�^K/g��褒�[^/��,M�J�Xt���>�g*�~lzT�#>�� �xA[�i��t�q�P�*�V���n�!/+�\A�] ��o$�x��	8e�i���W���A�K�(����h0��h�玀m7�X,����+��6��e(M�AM�Vx��[I�����c�����T=��O��Cp��"M4϶�Psk��P8���:�b�Z3�!ܼ�5�:��ϳɽ�0]o!�)!`�2��X�jP�7�v`c�U��na}�M���6��b��ǩ�r��!�{�x�vi|���߄���6N	�$Hw�~�6a���u�&x�ͅ:��9�h>��1 �y�u��:��hGDAGF3>�O�*#У�7��g���;�����\=�K}�$�OT5|T�<��g�(����)9�l�@C\w"�f�����%Ƴ��T1a)�Ҳn���as}z��2[�U��`���W���>���u$#�ވ��U������AYx`ދ}!35"���ĘK��4j�c�K
<�l4C����&���֦���W8�ZjB��ϒfP|H_#�ļ�~�7�b�M�߼��	[�ZH"�#��euR[w*��٤i�r8Vc�54� ��9=�E����c�/d�C�_k�h5lK���s�0��O��Hxh0��Ek��)�d�`�^^@|���Eg�׆2b�x���.p�
^�i��p�m�f�
~EEz� 
��/�a��r�j���?ҽ�M7{6��=,�`�b,���Mm���"$��kq�4���E���Ϻ���,�ƞ�~�o��p5��[Y�A�Z�T]��
9>m�a�p�_J���48�Ա�����k���BO��`�୦'�L�$��y�X�S%z�{�$p�� I�t}q�+���eYrgALѻBJ:q�h{+����r�Z�p~���[��:��ԟ��^L�B�rk�� c�`^ˇ��b��0�ّk[3�>a��"�UW���m9�&v�������O}<�a@C>�O�3�8��!�;�h<���Z��� `����HŚP�PPl;��!�q_T�t�L��V'�dH+L*m�.l��'�9b�2��*h�[�u��]ڊ �AX=��4^���p=Lb�K����xB�S�e��J�����~��RA��w���Ɏ���J@����g�W4X���$m�n7V(u��wr�����J�?�.�A}������VwV���;J�:h�`� ��L�AQ�ʆ����(�H�� ������}w�Y�I�����F��jB�視x�]
Ȓ��Hf}B�ZB�ڭO�S/N)��W�&Y�;U�
�s|o�J��2��d;�I��W��\�ɩ�1��7�1�=��$R�d��	l&�H���7B��W_�R1���vd$EOׯ��� �n	��?�?�^�:H'��u��D#R����t��>q�]l�"^���\��&ܛ�z�=��"�#9@	�1�r�9Sl�t�}?�|'�`$ݶ݄���F�@�}�r���|H��s~�#J!-��p���板�:��W�E� �P���YcSZo+��s�q�{^Z I= �&�'��~F���Aޖ5sk����sz��t�O�&3����8X�=WŸj����!�I�s� ��Ly,�GɁ���0M����T ��gV����Yq�����X���|MM~:����j���'�����e�ڶ�?����,�"B4�\U�e�'V��,c�y?�̸�i�g���)lD4{h���Ԣ�ۗå�g��J��~�vrEF9�ӽ6R�Wm��y��AƎ��sk�*�5E�O�]��2�,ޯ`� �-�@��^'��w9��P����v�Lz&Д�[��B�#=���x:zT���?Ɔ��bՏ��W׬[BҾ����T.���^���x,�n�_�-�T���B�� T�i��]*T�%��AI��.� ����5�W�si�e��K~R;nh�*�C��BDH���i�۫��,['J�6P�����V�C�Yȹ���N�BT�C��^3�P���u�^���]PA2�Ѫ���M�����V�o��3��x���]ݭ�a�3�d[�tx�ۉWo�)�.1�e�[�]�P�tC��D����ϸ-��/�iPI'�1�P0�����C�S��_+F����T�H��>^�sPf1u�Vⵊ�Aص����s׼�<���9�８�����C�x;�����<w����[���޹B%�R������I�O���ѷ�䒔\�@f�C�&��u1�^�x����*і�t�M�R��"�����(�d*K^��C�Rp&�Y�Z=��jY�H���h0�5|��ɼEda�8d�+�3��w�J�=۩̸/v��󘿅�.�J�\�WD#�V5`(_�
�i�d��!w�FP$�A��G}lMi����_�b�d�`���(�[�9ث��7/l��A�Rn������M��b�'��9܎�~f����+�9�N�K��� ᫢v��Sq��4p2 �V�՛2�������e{�$N{B�Mh.��q ͆�Et���X��ձ�z��[�����Ჩ��;��ߚǌ��HWrz*���|���tG�+l
z�,~������-)�=*GS��Xw��� b��^�cy<��f'k�Ez��.�Y������B�����sAQ���M�{�.}|�e+.��3.@�_jވ���)ZR�{�� �7͆Hތ�-U��� ÈL�N��E'R(�y���D�U�=}�Y'���&n��/n�%� ��z�G����6��n�%<|��]��/��44�{����L�	 ��DJ<�;��`~�؝�X-/������0S	���N�u�`��Z�-	�h�gz��}>�{3k
����9�R�y��N��9Ghy!5g	����ȷ����;=��A҂����kjJ	�+�V�ӛ^�Ns*�z?�2G���S�(�JQ���}Y�\��7��u��;X�Œ���ƞ���o�I}2(���q�~�2^���=�gI�<[6�������_Gf�qL�ֶ�̣C����^A�Kr�	L�^D�����6i|1V/d5�X%���i�K+�ЗY��=\�i%.�|fՎX���}	Q�ꔘ�I��ܘk�U�%!���Ht���#��fp2���V��p3����Vd��Q�c�^�k]W-�gK����q�VQ�����-'���(�MU*7�����7u}e��fPЧ�Kw��h��8H�@��z������J3�Ȭwl���!8N/��P?�BC�~���zY^��F�m%��0Tk%o�2ہ� m��yS��z���K[!�\��� 
��$�� 6c?i�?h��	<X[��F���	"l��5�j�v�#hR����O�Y��������5�;r�m����L�!��=i��j�'W#Bԗ�Ls�YB�R=hF���G�81a�t���b��`��m�I<<��� ��v_z��"<v?����r�D��.��N��e�:$�����ġ�v�p[e�y�l5x�c����aqpi�×<H�>�X7D���@��5����Ё����b��h����*?<�!ǝ��b86�o�#3nlw���n�*g2i�O܇<��I۪���A��T�w7R|Tt��?%����Q�����#H�)������@2�ޚ��?��Q���gc�#��P���+0p,�x�6A�����)���'h8�GC���+��s��-�}��<Y7k�H�F��8!�]K9���})���R�
s�g�os�r���'��ֈ�C�ޣ�`�|��b�O���8�Cͤ��d��W���F�j�1#��p����z\�z�	��3~��[]?�PFf?�Y)�_��Y�v��,
�����Ք�!�F�ئ+6SzXW��w��\����A)�.�j�,�|��;u�as�m������00��G��2�"&��J`���?�wY@m��v2NO?8�>m\GPD��;+E��	_����؉�_�:T�~ju}��GE�CL񹶙vTد�M!���7hTB�������ݍŭo������\�!k�f�*Z�er�����x�T잮�����%��U�#ϩ���{�e���M*Q�J��V̰����T-��⚕� ����b�@=Cض���К7�ɧ�R���w@�1�%0J��b�Y#���tM�*b�ߝ	ݹ�E�(��!:�@�br�#�Jw�9�y,�a��N�U�-��IM�[wһډ:�]Ύ�[�	Hڵ�c�xd�� �Ƒg(�G��p����P�c���謸p���Mt�]�=L<�~�"4p��㕐aZ��laE�y�,������=�+-��^����9���9���/�RY��I{��$�b�Ef�H��N=�im�����Х��Ѽ�$!�6�H�����ڪ~h,.�Z���X�6����S�mB2ϡ˵۱�Q��~��c7���璘׳�UhyS{��*P��.����L����_��g���s���j����K��2 �k��$�j�i�w��)v���D�� ���2��l��tDH2��O2��lR��c��J��$������|Y����Z��8%/1M)OyW��w���!GS\Y�	��%#+S�M�[�3/��4��i�^��~�lg�r)�@�}j�ژ�3P+A�Y�^��cD����rNK�@�F�e�}��!W11�ҚC.�{�S8�=n�&W.�\b��^�!�u�'h�.��Y6�Q����b�K	�@�m\)G]�
�1�j�]9$��x��{����_����!��fT�Pe�e��	N���=��Jl��R����{Zn���0N���3h%�`���|�ШG��I�G�!}k X~��o	�;�u��*�=����.��8�:�w��Gl�b��@umo:lUG��Fs7aOL^��+0wagZk}���q�\}�*}^�O��dT!������)y $�l�\�se�G��b[�e�=�Z���J�)0�n8�����zGm-r<��'�N�1�(\ȗC�������nuc�N��)U���{�݁��ǂ�25b���h��j�KJaݬ5��KH��x��OB�(ub8"w�j�����|����&��k��wH�����G�		��Hb4���;R� ���i�kV��5tj6����������:�Pc�@-�3Kk;ʇl�n���Y�10��6OᶉxF���>vk�i𤔔��O�|�E�9��r�Uxܰ:�n)�
�}ti�zҭ䐳J׵E�7�
�#3S�k/���a]��57����}폃�q,��GMT�I��$�C�q�印2z���楺%k,��Ѿs5�����$b���|�v"�J��>�&-˰"�J0M�t2��}�E�]k�_����;
���w}���4�5��X�^F%�c��d�Z�<�fg�k��nr����˒:�q���7er0�����~P+S����[U�3WM����hyH�D���N᫜��
�x�ѹ}3��ɳ�Тn���χK:�3�&�����2W��x�r�tn��5ST��:�L��9V�?��i�o����@ܮ�����'���\hq��Ц�%b���1Z{��LJ�"���Zᕿ.8Z�c6g� �f��^oר� p"�������4��ӟk}|��g*otA�t͹��� n�aIi^u
u�)|/�!"1@�{�i���� 7 �HI@���LUe:%֚�#���$��_���������ǽ�+K0�֜я@#�m�
'u�.�4�ڮ��R`>�	s0���U>��d�!c�1��;k6��L�¿,��p��!ר�^X��7��DZ��2����;�,4�����-�\���)�Th�����JrO���VJv�6�7vc_�U8 �>~M��(Z��U!�><�I&���D�f��o�(>z�d#ŗ�PŶ�o�c���_9t�G��r�޾�&�`�h��e�����ߘt��
.K*�w����U����e�"p*:�l7۪�6��?�U+�p����W��Ζ��D�L�	Km0��?W�sDB���.��v4n%ڙ��L�;y���t��vw:���_�zY�E�^A^5��L�jL��*����A�ms��%>m�2)���#� &�P��)r����x�u6ES���������O �Jk%G ͒�/3���Z��;'�B�'S͒$p��8�̶ʧ���(���Zq<���'�l�A��TH��)�<�S������y�9�N�~zʁ`6C?�����ucF���x�kЃ�l�Z^�)U���0�cO���x�� �k�����X�s�;|Q�*E��Q�'��x1��c�T
3��i���҂a��E�=�
�T�x�5w?4�}��Ҕ�70�%�8��U�,A0�MI�b���$��q�l�������v�ڮz,K�ѳ�t���˝'
��VuM�	}�_��>b�����J%���	q3�&渚Kknu���ܷ�f��Bk���0��ʷ�X(�%�������Q!��i����, �!r<���0�.:��0�
�L��r��D��~E�|�0b�$�:� ����L�l��g�Ɣ�y��䣇e�K��٦A��J�a&Ψ"��ʔ�aT9���&K4������O2�)a�w��D�35�R�Aq#;��g<�h���~~K �t���%HZ����;\-���5j�wL��WQ�VٺH�sAm�Hhڵ�79�s���C��:���N	��D�����]dp�l��z1QY�͊BS�	�o�R���H��A�Sƀ����~��?���I7L��}ˎ|Umt١V=.���R!�:#w��S�� �����a�Cf�Vѥ#;���hB�n�������"Q�݇�]�(���Ə�:]�}�*��>᭰/���(�=B�n���D
���`�H}���B��]O.��N^xrWc��ذS�
�@ko���2	��H�d��$�~=�Whd�\vN֩�Cf踋�1)���dq"�	��6����B�!�خ'��%1P8vY���G�ʡ�V���ƾTã�f�?k���� ��YA�����]����"�MI&�`{�=��i���a	tir0�5S!���d|ݪf���L���w���E@Zr ��1݄�F#?0|�^^���쿑���p���1PI�ݙ�lgZd_]��4q%��^/�;=�&+&�f�K2��V�ދ��kc���6'�sO4�t �&H�:P�8�̛W�6��@4�!3�s�������\H��[(wMZ2�����^ip�1�u�^�qj����QڏM����l�-1�7+�'V�����˖|?J���ǋ14~)U'dT'+`,�yT;o�Iz���1�~w4���8�ưa�/lQ�_U�3� �<F.U��R!�R #۸H]ܶ����s }C��Gy�D���������`@Oe-�]��������EF���$ަ�z��(�М�B']�#�^��O�zI���*ц�Yl�w��LE�B�ea���T���S�&�Vͽ�t��4������W�% ��Ki9@�*I�꜇�jA~��.�pN���JA�W��i00��@��;�!G�_,�C�ޜD�A�~<��`)N�{�'?�~P_Y.�+�CÞi�.ԕ�c�T<a\��^(�PM�eu�N�TKA��+�ʘy��mf��������������x
j~�r"w��S����[3�;%�X����Q�ot�I�(����&���qyo%өR00�a�u�U�^�7��T���+���裁'�"�ƫەz�3��^��C��p�	돩¸L�Y�+,���0�y��Pb��6"��7?�z�.��/+݆��J�������󂊵��Q�JN��Ws�8VD��_
���8.nl�w3W*$�c;�(�l|㪍�_�$1d�N������&9����톦l�ۢ�����
���9j�q��'�f�9K�~����Ҏ�H����>?�uxR�1�����}� >T
��8]��/�[�!e*n$���)�.=� ��*E����GP��-(za[sq���g��RB�j�R�(�#�{%qH�1�z�������c�+����[r��H���v�dL�X�`��Q��bh��ԍgpyK�uf��EI=�.�;�5��� ]p�Ztsp�����{��J|p]�.����2�@`��_α����)i�?{�M` �_b�5yt�UtyUB%~�o*K�{�ۭ�;RA�_yʼ��T|���c�UeU�_�'�g�&}6�/],���2�(�GT���8M���v<�&]�8�/��44�ŉz�ۖA	��J�R�<�h��o����ҙ�' J�X+`�M�m	&�WN�Jۏ�gZ���Wĺ�6��,��{�LJ�mZǈM��$�]>�(@-hH��5�H�=��7ʙ�n��j�t����Q�`[FJ���+��B�ق����,ĎA������dw�J ����o\��(�/���j@_š�O��up�i�w���/(|X�q<��2��=�lI�6�0�v"#�s�]_��q��`�,�oC�*�mm�KaA�Lm�3�/���2���>/���XT-���4�KD�f$����@\���%���f$)[X���}�\�D�Ig�x���c����%�����$��ƈ�uy�o�܀R�~����5O��3\%c�F���-�t��~!@�IQ��E��Es�Y��w%��K���z`y}4Df��Y��m�����虪��f�E�|�Q�#J�|�F(+4�tX��w&j�0}�A'�ړ(�U>��\̏�_,�m�޺�_�n0,�E��2Z*đJ���~�u0]mJ�.2���?]�>k6�G*�ȹ�r�W�_����m����T�:�u{�G��Hf�jm����#z:�gL6���(�DDMN2źs�1Q�ۂ��*c�����/f��$�|�{�{qo�/�3P
����u��[P�340'��\���XW�,�m�Ʉ"!`D9`ʤשQd�jiK�ܯ/����n���M��66�����?��f�v{q���h؃
���='96���HpH�g�*��G1ܪE�{}&���+��]گ��ߐ5����S"�����O���j]�"]�ۢ"4��/��. �F7AS�J�꺘O����"�f��Du�:e F�7&}�<�~҉S���*�n�-҃B�D
_��8ֻ����n�a�$��|�V�u��iP�b2��әa�31����n�!A���'�ə��>�`� ~��,��pͷ2=��O�$�������N*�T���(��6n��m	;Rf]r3g�Œ����/��T;�����Pg ��YR6����ud��	�n�d��ܦ����������f0���y�:�����QǴ�>tZ��3�g��y�zi�,�K)�|ʸN�SLT�*��������[Pk7$0K`�Z��{SN	�E%���d���-��n-&`�G�s���?��Q����ip��z-���������Xn�_��Ѻ!�3\���;�k\;�}5)&i��A�Y����;�������6�k��B���2�	�nu�����ء�&�9�X�12�^ۻ�_�p��n��3S�	��xjF���q�i�Ȼ�X�@�ј~3y̥w������B�����_��Z��'�J��"�d�ȕ��Z���gz�bf-t*o O�;"}�և$��4�	ӝ�|�s��B�o��tJ{�Ͱ� �vI�� 
sT=|�Y!��v ��gc֠��7�'I~�a�J?��Nښa�#�t�$�k�ִY�R����')S�0����#�G��uy��4i���>�/z0S��U��X¢j4!a�7��% k�:�Z�½p��Ѯ��q]���1�X��i�H���\���V�#;���҆[���k����A�)��=h*h�ԑCrM)��ʮ��i�v��SU6oB><|f��`>���5b��'����;��9pJ���I����1@���>MF�vX��r������%�-P<횱�Z�JW.b�f�Ct���&���E��&�]�j�M�0�g�b���t�tiH������i�Uꫯ*�T����V��@|��?��J_�����aP(�N�X)-(D�i��wn9�V�!�*V[����Q�c�r�d�(�����b�(~!GI�p��>�c���H�µ���t^��=h%~R/lp���,�юa����H��D�W=�p}^�#z�g"B���Ϙd�����/-@=�.l�{pƎ$��=Eo�d����i�l�Yd��Ųm]�$=����&"��)-�v9H~��%������6mLQ�o AB�����b����~�άc�?����s�$��y�B��
Pg,���!ܶ�ӥ��d=�a;�x�j�6b���2M��M$�@u�jXz w���vV8	`i S��2̳��U�4Dd���R<����~��dB-�����,P-��Y
%�8#H�Tx1�pk�G�4.��sG���Y��ʏ+o4O����3K��4�z��3D�˳'���D�T@��v��3l6L��`˅��D;(��N�b�@�6 e5q��=��1^Z��_̢{5�������x����Q=瑷�h�}��SI��/l�	T�K��8�$���&�v�G9@H�x�$���f�rPK�����]��l�7ec©N5��W3��f�B���->�y�4�����N�M3��`��a��c��I�ۛ=�f �5��ٝ����u�%���?Ϩ)���aT1:�"�D��)��U��u+*4:�̱G���F/XO374�z��A^g����g�\���}�1`O�ݑT��š�.J���)�u����\ӟ�B����|��r�v|�0h)L�n�� ���z���;a1
��j�ݛ��ȳp7�[�+�ܱoփ*�b�eU�`Q�ݝ��<t��r5�*@� ����j6�K��+��Т��˯7��o�D�h8��j���nG|�����@�d4�Dɷ�=��O�	�r-H��Q��[R7a��:��i�CV��R5I$R��x��������xc�X���kW�_l'yf.a�|0�<�O}��xb����k0�@{���	�|x�E��5���x���
��
�\�ia�����߳��E�D	
�<*?�7����J�l K���7W���VV�<��,�LM���w$z�_q���J�߫a����,���Zs&����{�����0��f��>Ik����J�(gӐh"ԍ�w�a@�k��^�����*��	���(�	�QFfX�m'%�E�� չ�X���Pc&��D�2�ré�ї�v:ͯ#W��SHr̯��ϋ~�{����Rq:ǟ�آL���N���g�#�<c���A���ܟ��a�	a-�"��2�Y��9�&�&�s}�L�X��OYkYa�M��+^�3�IF��]�;:A<d����ӥf� �a��m�H!H*�,�{;�E�M_��aoL�/s^U�V^�H��ms�D�<8�9>��@�T�7g�A���f�~�=���[���p��`~#x���Լ�S�+�6�o��q�5&���I0A1����ik��Ǯ�&"��޿�3�����m�ިV�����M��A�~H���~u&�S-����V� ;&�.hI�҇����9�Q�˰���(|��\&	�aƣ}Ӹ�%0R�����χ1B&�(�T��
$���s<}�[�Bq,�O���N��W�z��5�
,Oo��TÅ�dvd��%P�W��Q\ݦ��䨾�ߙ	1�� �zd8�	H�4����թO��k��+�1W"�v@�{�8��q"�ݖra�;�2����Fl��� 繅��V9q���]�
o:8��ec&�y��'=�p��F	۝�rwYSHˑ�k����uķ�Y��e��+C�@��rg-z�X7���H�#&7��%B���1�ә�3�� %Pp�>����ZK]u��}Lq̔�^�T-=�M&+�ۇr�`��ʠ�r��k*����as�Svt�+I&��w��8�W7W�"���r!ښ�s7m��(qsţ����%M����ڗ�%����*�I��q�	C�:jz�x�M�T��F��Go��'ݜg�d�c��?q81��l���a4EtU�
�'���,���y��y�p&�п�F�4�}6�����7t��������K�ZZ��(F$��lR�4z�?���}���[sG�Ҡ�\�+ë��N����Lۈ�`��-����:.�����,����<�)�z��z�7e@Bn2##ݑ�V��z0?��Kކr���'���sB.���4�T���: \��M��Je������0���� ᮙi@��*06d�NsA%:�.)�J����W��zi7��'s;yǜ���C�D$�]��m?ۇ�%��'&K�P&�����CJi�ȕ�'���Tc��	e^cP<�u�D�+��AP��xڋ)�1t3������=�voS����xqs���X�������[헵Ի>%7��4q����I�ǈ�L4�-����6���![����uCM�^��{���=��;�H�"Ô��bSi���^	'KC8e�p�2{��ZW���Yw�;�{q�0�����ℼ����wO�a�F���K�-��JE�/�Tj�%���ʅ�IJ5&wW:"V�N�_�R���M��wZ�&$����PlC�C��4�_><d�^���b��P9�~9�Ԭql���>�"�[�F�A��Ƹ��'�#9RK�~����<���CV��v�Ƽ�E�X����Cv�j�� ������)��kWeq
$-�����.$�� �d�E*Z����?T�z��N[��6���;��T��1�����2MH>��z .��2O���[o+����"���_�U�w�>�sxI��X�*	�X�bOs��TTy�;�f��LE��^.��\ ס����@+s7�Y�B {E��|�_�.�ѵ�jh@g�;_��/����)��{.�� �c�|��|�UIyq�V���Ba����x��[y1�M�y���	Ul�]�*'���&$�E/��ΰL|���|�G{y�?�'����<r&_]�QL/A�4j�9�5<��8	�1$�9��<�_6����N���U_��- �t>.	-�!N�fJ�Vg]Z�&���[�xǖs�{���t�:�o�
��?�[A�2�h��5��9�d��>������1#�P�K���4g���[�X7r����� o�e8;2�oK�����O%�X��)�]�h;�d���r<3�����c�`v0><U��9>�K��ᵱ�����dH��*Z�������[�>�N�#r|�P1�o�'�KF>9�l��w(�/�3�5ie�e�s.��7~�*�k+�V��b�ӣ�#e7��*'�O7hf6��?�(���x�ң�W4{����߰LQ�m]�?$L�D�-.��	���q��jچ��L{q����9�A�?��ݱ����N0D(��^.3��U��jy~~��s$�M��zdP��PU����ܕ� �wv���M� 2x$E(^���Y	3v�� Q7Z%t~��Ts��L��Z&"@;��L�t�����	ޞ��hw�(`�DZ~d�LQl@�}����pzq�i%���I��u����<8�M��X�BAǙ��&�Y�S�F���%�����o6���x�����SE��Us[K�\�M5�w
��Q ]R?gK	h��	�-[���5�ZU�l�5��v�hȍ ����<�Y����Y��tg5"�/�k�!G�!��������E�r='�"��գ.s��x xm=��$����^@a�Z�<�����k�W��|�@M�����fv�b�׎p邈�.������m:����$Mğ��v�(D[����>��a����q���Ն=H������>n��T\���CI�?4��<<b7g���"�*����6ޝ?~�b6��o^0�n��wIG�l�8*%n}�͏#<ۯ[ۨG�����W�w@�|RN��>�Q�|Sy˄�f)� ���>*l�X��?W �QX�N�e*#t�¢^ �+nR�,����ÓR�g�/��8��Vْ�8+�{��a�}A�6<�b���F�8�:�]����P��)�ќ�2sѻ�ha�p߆���(�E��<`��Œ ���58��PeC����n��/N��)���hM�1� �pm
�Ve"zmw�8���Y��~��]=m�F$;R�������W���/
�҅�'J����F��+��%X�Q�w�Xޠ��A�fz�����dA��"4��R.m�ή�ӱ�����	2�`PQ���Q��֊m�,2#/?ݬ�>��G����9O����x_��6d$�]�&TN��u�WwG�΍L��?�4��-{/!$��H�T ђ�N��(6Uū�q�_�8��!S��f�Y�b��r'x��P�;�Rj���+�D�2q���k�Hݩ+v�������f�M�l�XކՔ�8[nx�-2�1��o4��>8b�:CV���7jΚ5��D�ۦ?8ѯof�0H��bg1A�V�_t�L`�<��$��7֯L3Ĵ��B�\h@^��a�Ju�B�7��a2.N��-��I�wPǮ�x(�Ό�[�L��3��c��td_���D;V(@��G���pO� ��c;$G�$�cDkt@�I=�sT~�A�p]�~�8U=`�aC<�����&�'=�G�@87L�=���R�ʲ"//��P�L{�\Z$]|E�%�Y8L�;i+�~��������5'$�f9�Ɵ^������r�~&�*��Ց��6�f��g�B�������O��~b�c��Ր��W��h��ƩPy�?n�,�aP��OI2ܘG��`����ؼ���Z�=jҷ�I�'2�8�g�j�b��j�Z^wc��v8�`�N �32n!)�7�ED�Y��^b��[�� */�H�"d]����GY,���Ό���1ˍ!�m���汌1G�kY���p�+�Q��]�3m7^4��-��7	˕�(��� p��@���X9]3��/�W�#��_Dae��7�NI�
@���e�u�_e�1��՚�h{�� ;��$������^9�`;hԯ������݇�+�IKX��+�����Hj�h�9�C�x��`��LI��@{�}��?ᆎ��e�?N����9e������Q����g�ӛVV�~~N��y3��`n�z���fI�B�_a� V��u[����u
���;���4)�C+H:���� �,��7 uM�.:���GB�F���OU���ӵ5Ǜg�
A�t���{\;(�}���OҔyT���e6����)����~0\u�[$������cs_�$&�)n_}n6�!�_z��5����)��Ӟ���q���i��[� ��Qw��ء��I�U��DB�Oݿ!��${�5����Bpw�L�j�K�ʅ��j�IU���$G�u���fI�8 ��j@���P��|�c���ĺ�>��*&�� �Ew�	Y��H�%��$�R�i����ix��V��5r�0�&Zbʑ�$B�8c��(�R�ky�ol�$o�,�#]0��O�;6x��v�WkR��h׽\��|Z�TE�tǆpn�x����샦
�'=i��W�k-��@�E��
M~�jdF���qһ"�79׊�䫃�P�,��>M�<5NK���j�r����%�1��D��Խa�p,�#Q��u�tM[0��!Dg���l�f��T���FA��F��tx��R�!t��'n�M	/�K;AJ<І�"�����J�cؓ��k�ΚZ��
.�I����m�(�Qa�n�a�;��1�m׈,+x��ˣ�6-zb(�6�M�q|����X�_��c4cI3����p�u��V���y�V&pPN}���R�iכ���3���\=���E�Sx����U!G �`��M����j��������mn��M� �6zYV���)�/��'��{�?%�C�1�y�D��6�/����H�gf��n�1#�������)M�����E@]�&��S��<µ1-"����C�z�ٶ�],	E"���/{)v.G-�7h���Q�T�'O�x����ϛ� =D�D�eG=$7M]�<�c��:	���%fɛ�
SD~+��I�P��'6���p�U3f���4���V*�����bS������:D���By�����Tٞ�P������Gz��S:ep��=�Bg��n�ŦrIb$���'�>|��]*#�tJ�RM��3�^�98J�u����Q��;Vc��C�  5RU��U�d}58�����"�#�l��#-������0��&yC��:�߬U�Q�>4�N"P��z_g�+WyJh��]cK�7�����S4��T����2����s7��]`M4��bSu���"���C�dt��-<(�n�� `K�]����f��Q�]D�P9��J�u-�@Y�y��nv��"�ۜԈ�p���#}����k���+D5p&��k��:tYq����m�����f��k�B�ڦ�s���n\�(��K���&����'2���AP�w�`n���S���ܟu���di���r�@��e2N�lS��A��V,�J.A�T_Z��Q��"�Z+�����`Z:tqg�!fft2�o<�|��"d؂��A�4��d�$1o|�{+�,X�o��9t
�l���� ���INK
��|T��!�`'���n�2և�h7e_�I%�"�фs_E����h#��W$�T֛+��`謥F�/�0�K��T&?#hO��4u`��4�N��O?>y�10���U����!hr����?k{�D�^�D{��8
)θ%���X���/n��#�����;07�9Y�Y�fג�m��N&)hS�hӔ��{U�r�a��{
���Dv��U=��>#!��m�R�:g�����nD���������t.Y>t�#
U�P��oZ����w�99�9�yo������W��%�e�?��'��JE����*#{����W��;�qeϲ�*�iB7 �U6m��?OP�����jW̛]�;ףy�4L�{�m�U?���DG`ӑ���cU-(���{L����8�{(L�.^�怛�7^�	��hj[��y�����d�j�߸��t�� K9�����Z(x���E���w���8�T �%�m�����D�Z�|;l\�aܒ��`�7�B��6� /�(�k�Zb<���l�d�L�	���bs�U��f�� 8dᓁ&4�B���H�Yt��F[�?%*]��(�oΚ ��k_�h?ES�R��킓[��\1@#v���:Ɇ �&?��^h"0	R��[�2��:�ح�l��5��zv�U�h�|q��n��%l�YKŰ�񔟣��5��}�C&�e"?�F���1 �'mc��m�s���'=~�_HqD��a" �����v��A�����1�L��H�v� P�&�\�.{�S�<��::�ü��7�vI��[{$�B������i�Qq���m.H)Y@��������bj���-���Eub�&��!��*����I5b���o�Ayn*Uw� ����*����e`�<s�>�@ֆ���7�j�8wظz|�0�ɕt���Q�xL���yR�)�������$�����?� �Q������#�|����+r�,�Tތ|�+k)���d�18!>=�*_�+��İ��T}�C�<o���'�F�v@8w�z]a�����)hz��ǒs��eĢ����}�/֞�ߴsq`3G������͘i���bCc�3�=��:���
�� �?1y��p�0���z�k��W���~�]��bF���'���5�@��,N�K��
#��!���iF@��+L=�X-�w>��H��A?���@z V(�t0�w�m��F�w$�����]N'2r@ב#5�+��ۍ��mb�2��j?uހ>��G&�8��9\�#�_����g@��5�T� u��GޱL�����k�Ń`!�"G�"�3T�2������]��C�ܮ�XP��c!��	fR ?��0�r�$�����꜀�c����:��ʼ;߈*)�$��:��Q
����M�

�.��,3���k"-ʿҚk���D��b�C�PS��������ܼ���,q��l0�b�����;�t#�e����5�d��!���ܴ}�o�B'@�h����J�&�ς+a�9�Nr��-"���F�w�wE���$�[V����c��Id�ڋ��2���(إFGC5�p����Vc�^�B���q�t؅�="gE~L��p�({�����_�a�.�ʂ0���?=��^X�0����^YU�^]��J��/��~���!{j��$��(E|�A���	Oi�l����9�2K�g�$w�!�^TW���p�~~��*�p��[6g-5é �BH�6ˋY�HMu����o�8��)��M,�i�p6��y(�z�M�5��]3{[��mc,q4���%����r�%F���P6*���v�LHL�Ex�3^U��_'a�=p�����.~!�3
`t�Ʃ;�lj����:�X��n�U�M��6�_�����r���ʯ�{����y���I��g�g6q	����HZN�g	�A�q�U1���eh`�eՕ;收�#]��i�2U���r(��#/"��ف�!��<�A˼&z]ou�"^�1/~�'.�֓7+��tt��$z�O���ʺ����D� Se���7F�<e���.R����[�ҭ-�D�Z$��֥#o��lɞ�+���{��V�����jab����m�]+5�4��1�����������m��w*��A&�V�$ά�#g�n�qϟᲓ&gM��o�2o:D��������n�Sl"��R���5s�W��i3䷻���@�u��Z)�?�ʕt����c9�=X�����Z���d��"7����K��V�Z͎VgԎ�f�=6o���`"׆����W4�ӷ.C|�+�mo�M9t\[�'� ���I���
��|G�t!:�����|���78"IX���dH�R{M���r#��$�q��#f���"��EEC�c0�Ĵѧ�U#��8�"~Nu�h�4�W���r�>-�0�E�UVX��|��!{���c�kN#��4����n�+	������X�?������ߚ�0�;���,��]U�E�,�0�)�VBh���:rg���n� �Nv{�RUP�>��K�@7ѱm�#�&���a-�lD�32���ն>���#�UP�μo�~̘ւ29�:��,����>�u�� �e�6v��mE����"�*��!��mg����ek:*R(�7�XK6�K,?��,����mW��"�v@�(�L�O@mH�R?o(�DZ�0��$	�6��L��ڱ�L��ҷ�ތ�����h���V��5�U^Yq�����jd��,�X���q��5ҋ=C�J����o >�?���B���x��E�C�$/�$����. ��2%_i����|���Z1��;?,��?+��<���*�䷊��ڷ(��Z��X���il�n�Ǻ�����T�/��K� &���(87���YuBl���Y�o�F�Q%=E��o���辈����S�>~�@�[��\D��j,�%� (�?�f�h_�	��'[_�F�M��e#ul�d�5�Rv՝h����&Y^���dȯ��1�5�����W��y������Y��¤�3'@(�ԠV�s!��	�=їv	uW�a���������� ���(��n�+�>��Vލ[v�������Mq1.�W�/ :��6�or��J�v�=[NRR�u�b���0�\�#q�ţ� �GH<Y?!��ԩ_{�{���;u��1H�'�Fb����48*e7�b,�
8�ba�co鈜n}z�wf���Z*0&�8��<����m���N`��|rw���|�Y���H���Q�l1bu�lM) j�a������c�X?��Q#����#�i�I��+�J�,��~��M���j��2���8���}�+R�O���:}L�\<B�mŤ�FH�W8jZv]�:ʛ�@){�Β~sp_J���ʛ���pn��s�gU�`F_�+���Ƥ\LC��M��X��-�t��;�1�×p��!��z;8��öx�D�~2�K]��4F/����;e�h28���6�>��
v�`�r�P���uF�;[+�X`�w���;zA�͓�g�i�!��V �J�m�7��
���y�Űt^2%1�1*������`��m�*�2F�?hI�>�JhG��G��I����_y���7��q�T��1u�@sG��L��ٙ?e�ؘ�{!�:����T�#�����sW��V��j���U!��f�\��d�r�d������/��֦���x���Z�,�����
-����M��a���_��=���۪-�����W��b�k#C�:��
�`�e�Ϲ�*�m����0�ǣbr=H��HHtV��F~�(>�"`ͯ�ۤ���8D@ɘ�,�;J�:����aN%�4-5?�w��"�C��η�[��r�c5�zdĿ�j/���y (��G�k&p��c���U+��n�t�u=U�~���p�t^��n%�t�a��=��=ϫ�Y�=��뻎�_,�(.mɘqk�ʽP/z���9{���$�XE�҆ѣ��zi6 �i�d��nֲ���$j�lɱ�F$l���f~1��C;����6��>ÜX�B�@@�>z���~mu�c ������ Э�Q�=yo�wB�Pt�TZ��#K������=C�Gs��E9�ja�
��h�2ɭ���r�-��j��w��Bv#��k `.�2yq ���DQج�߶���J��8�z���ٮ��9PzI�Y��L��茁�/1�W�t��A��漒G<G�Yޥ�����+������3�Y_4��R���� �W�u��ۄ@9u��Cy�3���������D̢��"7Nt�#@w�e��Ҫ��1kG��[:{����|�O;ߥ�z��J���bh��Ś�?��:�����?K2������x2��s�h�9�x��f������y)�̈J@|�5n��p��Vu#�?���4�hc+�J���k�l��!L�}�r'0���O�9�x���rhik������ؾ�|VnEa_p�l��x-E��,�
X�i��b��풳��EtwE
 ��]IKfI*d�I�ʅ��7�a75ڐ�7Gr��1,&|'M�]��6$�� q8#߰�^9�}Z;��,0b��8 ������6�����5��N_>�kA��5J��K�.����ֿ�+�ks���<-�5���'�����X��%�ns��!W����_J���e��ra�1����:�j5Q����r**�ԕ�~�$ՇU�O��T:#���!JL�yT묁Y���_��c�����ӝ�v�ca˯�"��w@E9m��&p`a�B�v�AO7��a:.��R�3ʒ���a;�@t<¸�"H�Ӄ�� Z � �yH?��
+;����О�?L�p���:VaN�H���mQ#��ڳ�9���^�f��B�����8�w��C����pw�ˢ~�uV� �r�S/��TDE�+�����T5�AO����fɈ^���E�.�"�wm���m9H�V�u��φ~���z�0Λ�rZS���Ȥ��V6�g;&Ph��:~��kQA.���!(�UW�z7�?��}q����T�խ�=Bėá�d�
B!�e��}<�BώO�	N�E�W�(��u��
Jܛo���:λ!fd�PN�� W�7d��������(c � �	R&�[�gB�:����'El��_5�v5v���h�q���T�%��YK�d��	Σ��5����ҧ�8h&)�"t`�FUw�1u�'mx4�m��s�5��=~6V_}HD�Pa"u'�����ߪ ��wM�����L�S�H�Bv��m�&�(��h.{Ay�<�g::S�ü��7U�vIs�[{9�B���K��i�Fq�{-�mcH).�y��#���,�b����"�����b�[O�!��*��'���2b�6�o�6�n*�4w�U��i�*� T�eu�<sH!�@+������jIw��|��ɕ�,��?Q�-�<��yG)����/O������Z�?��Q�J����#�*��A�+��,��9ތ��+������d �8!3�*�+��(��a?}ٸ�<o����IF�ˍ8w�r]aE����)h�i��<}s�.-ey����}�L֞�Sߴ��`3���l�ͭ�荣Cc��2���s��?� �91y[2p���=z�����L~��C@~�]��aF��q�'���5^K��K�e
#����.��cmF@ME+LR�X-w>��H��A?0��@��V�0�t��w(@m�]�wo���ը�]�2ru���B�+"xۍĄmb�H2��Z?u�{>�lG&���o�#`|_�� �߫��8T� u�i*G�L�����j~�Ř�!����",.T�'��w����Q�C�������	!�rfRU���%Or��������q��c&��O���q�߈-������.�Q?4����M��C��,���J��-�T�kv�Dv�beSC�e��Ϛ ��Q�ܱ\���h�#W0��Cb�s���PRt#�b�+�5�b�϶ɯ�,�}a���@�}���b�J?��wNa��NrΕ-"q���Iw茉����$ �[K��˂�c�cd����m��	(�Z�GC��p����rbc�@��B�\���tؚl="�~L��p���9�Ք�a��ʂ�����R=���X]����P�Y�T�^2��J��/�����|{jH�$�{E|W��R�ޢi��Ĩ����犲g9�$w�"�^�v��;�p��~����p+e�66g��é��BHˋ�a�缛~��>cMM�U�m���^P�y�V��SYPa)|�{��0�,�����^'8�T�h��1rj��~��@�2V���J>��!3jR��w��Mv�by�{ M� 2�@��aID�;�L�)�$J;�����u���(�f���Y�[2Č��r1cg�%z��.��I+Gie�Y�����+�ł�4OQ3\Q4�9��m�W�-�L�BY�V�@F=&��B�3&��y%�BޚD�zl] �N�h@$��e������1X����){��e�KҼ�߲K�t�"�K�Kh��͚1���g#$�önK�c�����%����� (*9zN5x'�T�Q]ɂld��iՙ��z�&*�e]C�NE�ׯ���� �a<���[G�����
���źNQ�>3~x`���WV��_�I5���-� �I+��Z�1D&u��Ķ�ak�c���]:��ߙ>IIM�H���cu�:�HeGځ�F���O���ych�I�gp����a��\�6}!nrOj��T�3Y���E��u)O����\Ϡ�������2����J�+�)n�uv��Uz]��H;?+/���:�>���m�"�?�eWα頡95�\9 UI�����W
�6�p�5x�բ��U�T�jpiK`�݂�!��hM�q����K��՟8��j��,��8�|^|*����R��卜��c���ݮ(	�Hx���8�R1�j�t��iv]Vy^�5
��i���?�[mj��u�cGV���k�:l!��h�Qo�z0�%�Ow�ux���Bk����:�V���|�E}�݆��x2�N��U
t,�i[����ѳ`E�a�
��y*�N��4�f!�S�?7��0�S��6�,B�oMj>o͂�$t9�qT���H-����[����,L�����$��"���P]�ׇ��ߖ� L�>C-`��+JFQ!�J�!ԇ^��NJk��X���F��CG�������X���%���z�:�:a�Jِ��y��r}gё��:�я���r�e��~fQŇq�E��:?��)<wL��$�H�7��B��󔇦�^�zs3�'	h��a�y�"�M��9	�s&�ثw��
OӂiaVTŦ%<h36�5�b�h;�S<^��>���X v����H[��ǰ;�3��G�����Ls���\V���H�f m���?98ݢz�U����`�Z�רw�:�����p݌���S�&˴�+�S�q1�p�5s\���a/���Ak�Y�9�ɤP֊ ¨�J}졭�t���m��V���k�2��%�xBk�շ��F���I�VR��;��2h�X��k��iQ���@(v������ۭ�}��޾޸�0 �I��B�K5�N�T
^L��5�}XL�Bk4O/�PN��W�82���
fc�o*-'��һ��d�{���W���\�uߩW��Y�1� ����dr	�9�^�գx��Y�mt{,1a�v:�����E���[R̾������ �$�93ڏp���_��w]�1�;��rص&�Cy1�=�k�9٧	��r��	S¨D�%8�噤�����3p3��w@��sr�����E����# �}�_
�;�b��F��-~�Bj�P��o��ZE5�	UtqFS�^p�=�&e�0��R�����l��kd�	�W��s���t�ʟ&ɑ��'O8nL�W����A��!T�s�.�"j��ԡ��DRM�
q�����_N�Rw���q�\��t>��
Mc}vІ>.��XA�'��Z�^B��L�?��쮯���yU4��UH?'l�K,���y՚����}-���9�4��:p���"��0��hH���]��EFb��S��R4���5��RT�,
s��C�K퇿%k���>�&�BP`���-)�3�i���^�&�?�j���z<���1�B��"#��z��z*����&���(����MYBhz��s$vTD� �4֑�â�ā�u1��*�}�؈� [x�i��**F����A�0.�j��Q��7[W-��i��G�!�9;�p0��[�C��D����#����G<' ;P`s�L��Cc�ȏ ���X�T�I�ë�^	�KPN�u������A��Kb=���.�^��v)��{���c�I��xkX2��ܨlؼ�I[�iU��%�������3oIL��;2��h����p�O�s4=�D�u=�\^'�Ͽ������T��ꣂ	"=����Ȭ��^CyxC��pV�E��:{���Y�Q׫5�0�J������4 ����X�1A[*AN>��c��ZEv��+e��g�� �{-��A��ܒ��w��b��t�h�q�5��	����I��e���>+g �D�~��>BJ�;`+�	p�����-�}D���������n�JԼ~�`�N\�f���Τ>�f���L��f���W��Z(Ј�q��2H�@��IX�6��f�A��G��_*'.q����R�C�ȗ���K5Z�L��G�-s�*����/��X(�r���K��кk"�p	6\�m%q��fx��X��}l1��W�JI��_��8k%dIA���b��V���d�C����h���/��&�{�cf�nn�-��p��2�Qp�B����-С��2�X��\�N�N]�}��/f�r�"*8ٔ�h3�}���*��г����g�fw�Kg3�x��	��p����a�i:�O�8IE��Ĳ���F����DE�m[�(&=R���1 �����2�!,�RVS_|�z^n�Lgu���"�ى!n�,�X1˸B�t��g�i`l��e����`�A���tߜ$ѕ�Pv��.����/�h�A
��Uo8b��
a��4~��Z�@���L�	���z&(g���. S!��G�.m���,�P���(6�FL(�� MUn�Z_`�V(�c	���N�0o�ǣ{�Ƃę�{�P�:��V��)�L��3{l[�"�����/Ԑ�!E`Q����*}j��*��+����n���MU� 6:^�c����E���`�{A���� ���A,�ݼ6��x��H��g&lS�.�1�Y��b����<��b4]Aۖ�O�z�\!���6"�ҁn���yG�˙�g]�}�"{�-/;Φ.j�7(љ�S��a,�O���G𘛭�,D���e::7�<��C���{ȱak&�����mD>PU�	��֢|��c幞����lE�V�ic�͖bT�������n�q�x��ҁ�N���A�e�T����up�N=~G����f��"�r�{���x����4w	R�3�b���,��5)ݗBvH��͟��E �
R��M��rd=��P)�����$'�v87�M��]T�0��Qyk^:U(4���Q�Ir>����,a�gd��y
Lw�\*YKP�Dʿ�MS�x�Ta�Z����HI|�7k��`Y�׎S5B����5��ȸd4�G-��ndٗ`}��z{��&Qk
�~k�
��-w���_������__H�q*����ȴ��[̢-�kb���50#P �Tg�Y1x���R}�P���OX�]���bʦ��܅г�nT8ό4K�?=�&?B}���2ܔ׻�V��7��nH�OSY�D��|��5�-�$��i�[��FX@�|Y%7O�,� ���
���fQ�Z��q�"��s����d��Z� �g�FTf4�Ro����l�n"$]u��^4xZ��}�|�`R��Ԧo��t�yB�t�W s��I���   �  �  �  )  p*  �5  @A  �L  6X  �c  �m  �t  �~  `�  ��  �  P�  ��  զ  N�  ��  '�  |�  ��  1�  x�  ��  �  L�  ��  e�  '�  �   K � (  �( 0 �6 /= pC �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'���%u&q+G���'��Y0��'���'oB�'���'c"�'�"�'�z9Yq��*g�Hr�F�A�^�ʕ�'(��'WB�'�B�'h��'�2�'b��yQ�H.&�*`�`�I=�\��'���'!��'���'��'���'�>9Q�� ���g���l���'z��'��'���'���'�B�'t�H�r�P�7 ˔�G�VC
�a�',�'}�'�r�'B�'��'F��s���L
p���M�,\���'/��'�2�'���'��'���'Z��ql
�lr��D�":��I1��'���'-B�'�R�'a��'�b�'���a˖�c��X{����TJ:X���'I��'!��'���'b��'@"�'G�@u���\H93B�p?����'X��'8��'H��'�R�'5R�'V�H5�-r�,�C�$Xd0���'l��'��'x��'D��'RR�'b<$� '�<3�)�� H8mxv�'m��'��'��'���'B��'c���Č��Z�b䡈5'�iCu�'�2�'e"�'�b�'p�hӮ���O�x`E@�a��B@���EЀ��Gy��'w�)�3?�B�i�!�B#�g�̥�T���$����?��<��mA����4�B��m�����?5"���M[�O瓩�jH?�0��[��<`����B�^%�2"/�I̟ �'��>�"6��Q�
%�QI��/�T-Cr�Z<�MC�a̓��O
�6=���#J=Lkܽ@t��=�J|�@��Od�d�Pէ�O�1 w�i{��ܒبg��
`.U�p���[�h������=ͧ�?I��)X%8dyKT �Q�"i�<�-OR�O��m�N� b���W9�A��>e�x���'Q��T}�I�@�I�<��O�9#"�%%�|SG��j��Щ�����	�i�,�C�:�6i�R�Z��(BU�D(����/�l������ry"^� �)��<� ���u�"L�MZd"%ώ�<�S�i�ށ��O��n^�S�;eպ|H�bk��vR`%:� n�����|�ɾ���lm~2=��,�S�U�H9'!��jX�ђ6ƷVjڠk"�'�<TS�' �i>y�ڟ���֟��I�f8l|�Gꐝd���vL�$[|*5�'3�6��U�~���O��$�|����?)�ɐ��h�.)�T�ZG��#��IӟH��x�i>}�	��,��aó$.���4eЁ25�c�P>?4�hoZ^~�`�B�����?�����<�/O\1�R�@�c�  
R�̴yIrd�ҋ�O,�D�Oj�d�O ���<���i������'O���O%�Pȫ������ti��'Zr�|��'���ҟ���џ� ���`P��d�M���g�zF�lZ�<���_�p:`?��'����w�����E
&O�-�bM�:7����'\�'�b�'�2�'g�>���%Ƒ&��|*U�ߦ}k`�B�e�Ol�D�O~ow���͟��ܴ��)�$����d��Yk�f��f}+I>i���?�'{(�1�޴����2$Y�Fß7���h�2Tk�Sq���-o:����䓯���Oh���O���A�r�>�Y�S2� ���ӄr��9� ��"A\�mK�f%�3g���'���O:���c�t�eӎG�|��%���yB�'�:��?��O{���,Z�N�!�F��^����-e<H���ýjw���I�?�� �':(�I�[Ij扂�<�Y�K��7�&�[B&7W� t��͟�����d�i>u�I꟤�'O�6-����yHcG�^� ���}�(}*RI�<���?�,Ot��<��.:aK�l�>}kҠ{1��:�����?Y��#�M��'hNY}�Ԩ���Մ
5k�*�N��"�M	c���<Y���?���?���?�*��HRwm̆B�� [��Ú@��U��򦭉b�ڟp�I�%?�	�M�;:0��KNn�� ���	�4]#��?�I>�|r���MC�'<*���e.�(0��;AQ9�'\6 ��������|�Y��ȟ�YV�PT���IF���D}�U��؟���ߟx�	Cy�~Ӽez�M�O��O� b���C�i0Lu 9h�(�I���OZ����Gy��m�E�T*�FL"��&?ѰK�)Y7�AD�׊��\5���
�?�@��W��d�S"�$2μ�1�$���?���?���?!����O�]���Αf;�\�q��6)���r��Ov|lڭJU1��ԟ���4���y׉¡ ��"C�_�;���Q��_��y�'d��'׼i��i�iݱP���?5Z��o���À�0Il�������'M�I�(�	ӟ���ӟ��ɷ`<0�kZ�HK���%�wJ`�'�7� �8H����O���t�	�O:��>	8��0D�B4[ΚDZ�陸m�<��'���4���$�OR@��B�nl�A��hH)"�XP�h����6��<iA� )�����?�eW�<�*O�ۗ,��e9�i�EMZ4y@w��O4�D�O>�D�O�x `#�<�V�i(�28�>�Z�V�(����UFUh�U��'�d7�1�d�Ob��'���'2 ���z���@a,V!�U�-/.��i���O�5Т����s������ 5��;B@�8�㤍�o�,�'5O.��O���OV�$�O��?yS�'���&"��F�*�t)
t��������\h�4iÊ��'�?9��i�'��]c1iL4���[4�S�M>j��3�|2�'��O:J!s¼i��i�5b��
 	�P��^'?� ��k��0:����d�'8�Iٟt�IꟌ�Ɂ}:0ٹ&�Αo��h�2"O--F�D�I۟\�'�6-�6����O,��|z��}�Bh���k�kCM�z~b)�>i���?�O>�O
.|W��?�@nFe&� ���#qQ�MrĲ��4��X���`��O�A�1���Lc���$m�x�i���O8���O
���O1�:�EH�fLӸ�b,���6�j!zv!R���'M�`w�D� ��O��$׆l4�؞�|��U	�UYr�d�O�����c��Ӻ�6Z��U	�<� o�r�a1�d�)+�
	R��</O����O���O���O~˧b44IWc�G���u��'m�b��iq��h��'�2�'(��mz�a{ �K$9,�K儇K��8�m֟��I|�)擊�6]l�<� .J~?"a�i+�^D����<���&���D4����4��&�%���S3��a!��Nv�D�O���O|˓G����J9~��'7��.wTH��`�z`�
���O2Y�'���'r�'-��Z��@:7�8y@���Y"���O�9��Z:?�pD�%�:�?�%��OM��Er
�)��?~mB�OF�d�O�d�OJ�}z�ZG���S����(�&�y���=�6�޵>���'u�6-'�iށ����>"�xb�I�k�2�B��{�P��ߟ��I�c�LnZ|~B��L�R|��w���%�3�T`Q��688y��|�^�����p�	��	��\{OJ�18������Z��-��xy��t������O��D�Oj�?��KEk�,A� �V��
���%ȟ���OJ������	/HcJ`���R̔���ȟ�3�ԲףG�����'7Έs��Ο�Ӗ�|�[�l�h���`�<��e�ҟx�����	$���By�d��ԣ���O����o�<Yy�����ۘ@y��Od��O���|�)O����O���1u�:lJ�k��1Ϥ���#��@��kr�@�	ǟ, ���c�TU�4��Vy��Or��?�la�P+��[ڬ9U%Ǵ�y��'�r�'i��'����ǚz����b��tÌ\1u���P�p��?�i!<):�OO"|��OR��*�gx<(@+�L>)���$�O��+�x��ش��8T�|���P�y�Zˀd/�%CG�@��?1��(�Ġ<1��ɮ;3����K�Ha�5�ML+�O(�lZ8������	v�D�U)D�p�1]2<�Cċ���EB}B�'�b�|ʟ葑��:����W#�Ce>H��TzHP2E遯y*���|�a)�O�I>��i�`q�\+Q�P�k��I�`/���?���?���?�|j,O�oڂ$�9Ŏ�E,���cX��8dޟ�����M#�rd�>Y��M��3ꖙ�\lI򄅐L1ֈ���?q���M��O �:g悯�2I?I��Eށu��Bh?KH��#�k��'���'�2�'O��'�哢O�a�œ�]Yz��O�<��4m��)O �$��8F�O��d��]	
�lM�5�Қk����VNR}����쟤%��S��L�	��~�lZ�<����7s/�z�dH�C�*����<9�A |I���z��~y��'��"v|Xe�j��~����kN)k8r�'��'���M�q�?�?a���?�v�H
}ˎ�Іm��z	�ѣQoU���'����?�����z#$,XU�E��bx���4[�'�}���@�t�����~B�'�00�� �z�,FE�m�e Z�<���R:|! =��R(�< Cp�A�?���i���U�'
��n�z��]�D�f,��+H�62��UMב3�\����Iݟ���d�ɦ��'t~U�5��a��lݎJIjl��∞%��T�	�?QcK�<)O��������O����O��!`��9���G@�,�&pHv�<��i��՘�S���u���'�R�B�Hxt�U�_}�(���0y�I����P�i>��	 �Gh�7}��l*PA�+n��(@Т�U���o�[~� ��"iV���䓶�d$4����ʂ8d�*q��C�Ah$���O���O��4�,˓@����4���¨��ـ�@F�HoR�1r�xӞ⟘B�O��$�<��H�R�V IEG������V�3B�	Qܴ���[	P:�8:�'@���n�+��̲�L^�HN�I����2���+�OX�	���,I�2)�FȾ�(`(�Oz�D�O�Imڿ +�+\�Ɯ|"��.)p�I�A�U8����(J�'X����� }c�V��L��O�=oR�<���;9d��YPz�G�oV��4�D�<1��?����?9�-	��4!��_�>5����?�����D^֦A��Lğh��ğ��O���QA
�4�ҁ�ӌP�C��U��O���'���'�ɧ�I �%�R=c����0j����=D� ��-�7Wv8[S���ӹo��|�	�P��x7N��G�9��'սC�^��Iϟ�������)�FyR/m�������p��L���ِ|�0
��Q޼�$�O4mZ�aC�Iݟ ���Y�d��A3��֎#�;�ȟ��I�I��)lZZ~�#�#w��=�SJ�� <�*�+T;0���ZR4M�%��7O@˓�?���?i���?����)�)����f_0fn{6d7ElH@lZ#���I͟X��Z�͟h�������5?���:3-
TNd�SĎ�?�����Ş&�}�ش�yR#L	e�Ό(G�\�]��A0�Y��y�L�r��)��Z�'���֟���b�&HQ�/\v�J`8��;L���П���?�@D�'�6M/U$���O��䍤G�FqZ�OV`�����i���D�<���(����H�?q��Ҥnk���I)�}Q"! �<���HшѩF�<|3.O<���'�?	���O����|NT�ǯ�S�"�Ba�៼������	��G�t�'��`D��1O��}QE��V�ѹ�'�(7�"�n����4���ɝ�w���S��3C��(�?O\���O���;N��7M0?i�LV((��)C'�y��7RVJUrF�H$<$LT�H>i.O�)�Ov���O��$�O� ����
?�USɋ�uZ~�2a�<!ּi~���'Zr�'��O[�N͡I�F���iY�I�"��c��/)*���?���ŞM�zJ�}��ՙ��P�T�w^�M[�OB	"T ���~��|R_��Q$M*;�0Q5�@�~;0e�t�����I՟��ҟ�dyr�t��c�!�O*kP/�S!�t����R�@���O�$mZY�QG��ݟ$�'��-�j �C���`懀��`P$�+Ư��������}N��Px���eာ>� � �G�CB�2�`����ǟ��Ißd�	���2�f�9oI�`jD�g��;�Α����O}m�,�����0Qܴ��`�Ũ��-;d���f#�|�t1JN>����?�'#.i�4���3P1̈�EH	[\���ٺ)W�kU��(�~�|�V�����,��ПH*a����l	���@�Լb���d��Zy��n�6@Ԉ�<1����ɑ>��)HV����AwE
,/��I���D�O��<��?Ś�JĘZg�͓����r�����i�D���w��%ʥ<ͧC>��Y�?˘A��E�9b(Y�f��%��D�	����I˟��i>A�Iןh�'L6�"\m�pK2/��v���S"�wC0�����O`��Ȧ�$�������O�5�s���F<��@�]���Ps��O���@4/�07u� �Ie�x$9�ܟtʓ7����Ď�5I-N[F��(0#��Γ��D�Od���O��$�O0�d�|�g�H�D�T)YW�+�t�rV��;_���%�B�'���d�'�7=��� H��m�@"�	�K&���Od�D$��	��nR7�e��!èΥ8�<�᠏"""d*�g�T�s�	�!t��Ey�'M�� 7M�
w#`�K�!$Q��'���'{剏�MC2Ȃ��?���?����o"(�Q��`m<E������'U���?������̙�$��hoM�RV��'<@��D����Ȅ�~��'�5��Y$e|�1jҨ|�L���'�6�z�cC�
>��œrN�!�b�'q�6Mv�j���O�TlZ_�Ӽ��È�L�Z�ɂ*F?:A���	�<Q���?q�6��Xܴ���яn�uQ�O_�hŋ�4C̊�Yo�x� ��E�cyr��(P�X�Ba"���S�
��jy����,	������	_�'6-�w�	� tJHؤ�����	9�S���Ɵd$�b>u�ėNK��g(�5�e��n�b�lZ���S�WCa0�' �'��IupR��֜~��� �^���I�x��̟"eߦ
��L�'w�6�@;C�����3Yؔ�B��@{�:���-A��DZ����Icy��'g�듖?1*OP�iۣV�h�Z��(��ғM�`��7|���ɝPL�9���O���'v��wz|�x�f���4�L�e���6Dz���I��(��埤��П��:t�N j�91D�ǘ�(����?��?q#�i����ȟ��o�X�	�@�8��¹(w�H�e�Q3T�'����ş�S�J`oZQ~/Гl6�mZD)�-R<\
��(���"�g?�J>)O����O����O~�#��� Ls�ib�B�(��)e�O��d�<���'Uf`���?������xdTp�Hʀ�8P�Y�<i�ɤ����O���&��?���f�`)SC� |*��f��X8X!���2?���|�M�Oj���n/R�Γ]@�Ȑ,�HW|(C��_�o|��@��?��?��S�$U���?�M�G���(=��QҪ1�f�@���Q���*O>�$ �d�Orʓ�?y�-��X�P�ߡR��#�a��?���%Dm#�4�y��'S	����9O�Z�N�{f�!��fM S�$�v>O�d�O����Ob���OV���O@ʧ
ծT�f|6Be�� E�-�M�Ҹi�HJ�!�3�b�'���O�'J�wb0���P�\��s&��2,���'X���i>M�	��%���� W\U{���5R�)���B�̓f�8���O�@`N>�+O���O��+@	
.(����a \�T����`�O0���OP�$�<��i��X8�Z����1%ؘ�9��=z��]���J.<�?Q�Y�h���T&�sDQlW�x�d`+uh>,��!?���ȲlD�8@ڴ��OȊP���?!Ъ��Z!�4�ϪsK�l�%�=�?���?����?���I�O��r���GNU�� r^�HWM�ON�nڵ\�I�| ݴ���yG���H��	�м�!^2�y��'�"�'�vIPE�i*��4/G���ܟ� 2eab�D�:`�* _�`Uj�:�$�<����?	��?!��?!"��7/[ }���X�KyJ��i�0��D��M�q�F��P��ԟ�'?U�IB�R�q�*�7kHQ8f2�!R�O|���O��O1�bt1���W�(�&�ϗg�qP�K� Ak.� �!�<�J�J
�ĕ�����19 aJ`GX	,\^U���N�h��?Y���?ͧ���Yæ=A����p��K�h�p����0r�����+Y���޴��'v���?����?��n��xݞ͋�T� o�Ueh �r�L��4��D��\4�������P�s�痎Y�bD\�.]�髒7O|���O����O�$�O.�?1)��\Q�5AU��l��i����ӟ���џ��4�@yͧ�?ad�iv�'k�ઁ�QB%T��$+H6f��i:2�|"�'��O���$�i���+�j�A��U\r��(S5c�%J��$���6���<�'�?���?�����	>�$J�-G�2IZ$�[ �?����ę�əńןD��˟8�OA �@i_�v�ToZC(��y�O���'H�'�ɧ��@�C 4A�LY7bu TH4��~���&�N�x�us�����*�BLM@�h��h�'�*���Q���=�� ��͟��	��0�)�wy�%q��5� "d��]��$����IĘ��z�*؛���u}b�'6�PI�#bNT�r�(Y%Z����b�'=�.�������������<��e�� m��(A�z����i��<�(O����O��d�O����OH�'�2]�!u<!3 Ϡ5��
��'��dA��?Y��䧁?1���yǕ�v�x��@�6-��"��z���'ɧ�OV�y���i��F�vF2�I^�E���Z���X��t�̟xqB�|b^���؟hS���8-���a�GQ_Z;'D���	۟��JcyRO`�x�!�C���Ofayd�1Ht��aD�r�"��O
˓�?�+O����O��O�uA�LA��<SA��z���2O��$�1(zP$W:2$˓�Ba��O|���9�XĨ�G!�n<���ι6��dP��?���?����h���_�U@<@���d��=qbm t�������
S��d�I��M+��w������R�Dl�xQ�x$�s�'	��'C�=˛v���ݮl ��SLRQ�B�]�Xz PJ	�>�蒕|BZ�`�I��<�I��|�Ip�"�9k�(� �-�5x���sy��i� ayR/�O����O�����dV`���"]�H鰁��
m��\�'i��'Vɧ�O�b<�g�6��ġErR�iH�L��C�J��c]�@�$�64�Bf�g�wyN�xà=B@.��e`����EY7h��'�b�'�O��� �M{�n^��?	�L�_�N����81�7N��?�c�i�Od��'�r�'����$��} ���yC��z��0ۈ�(�i��ɦ#�l|�tٟ�����"��M�TW�9���ω�|�D�O���O��d�O��d3���[��Jtj݉(��i��@ϸ|�8��I៰�ɕ�M��*_�|2�s_���|"+[er����S�dQ���@!��'�V�؉�A�æ��'��=P6��:V�T��FD�Vy���K	;����	�Q�'���şl���x�ə����2�K;|%��#,Դ�����'� 6mCw���O����|�,حm�� u�2�	��ZI~R&�>���?�N>�O�@x�d��}�@����+�.���
O<�|���G��i>����'�&�x�Ŧ�.@^��$���G�B�S`�Пp�I؟@���b>ݕ'�7�M\�PA�p��`z������M}!�F��O���V��9�?��_���	�=�p�y�'=��� /�!l�����؟T��		ئ9�uw"<���/�syb�A;u�Ii����2�L��l���y_�x�����	�������O���+<���'Y"M�<LP�KjӚ5ӑ��O���O������Ħ�ݏE�:�rdȲ+b�av	F(��	�$'�b>e��Ǐ��y�:Ī��`کE�R ��J݄qߜ�Γ!
&��䫥��&�|�'���':a�%WY� ��D�_~� �`��'B�'=b^�H	�4\S�Q���?�Rf��@*��Tc�J�m޻��b���>����?YM>�f
��F&赛��"�
�Qp�e~��?�(�ّ� �E��O�,��A��I�	�N�`�q���!�$m����'l�]��ɟ���0�	E�Ӷ4��П �����H7�`��Hl�%N��J�4PV�Xp��?���?	-O�9�����@	���Y��Ԭb��jW4O��d�O��$E4�6�b�p��O��R��}2���3@��r
��"�Q�� :�$�<���?����?Y���?i����(�L�b���.��"�!���$�1�E"؟$�	ן�$?!��F��r@�=|�)�Qo�d�T��Oh�D�O��O1�qq1���wҩR��a��hiW�˪��	�&�<9��V�$�L�d�����S9_�,���)U��LM�4"�#pTv�D�O`�d�O��4�d�c˛Fd�*�h�T�D�S̷3����W���y��h�㟤[�O|���O���H
NT(f��4Iv@�)ʂ>EΑئ�iӲ�(�	 b2ʧ��;&K�'.�t��Cō1��K����<����?)��?	��?!�����X���?���K�%ſBEb�'�Os�
(�F8�$��ަ�'���K�d���c�	J�^`Vy���@�I����i>5��A��=�'�D�
� ~�($j
�k���RK,V�e�aՋ�~�|�Z�D��۟X�	�ɷAk�N��b�8REZE�T֟���LyB�|��u���<A�����yR���O�Tr� ��8t�I���O|�$,��?Y�W�c�����9*�ʬKȥ~�H�q��������t��o?1O>��h�bB�AaTAT*z��$1Ш��?)���?���?�|�.On@oڿ*�L��������l�;
J��!�Dܟ�	(�Mc���>�OF}Y�����p'�"Ob�����?!�́��M��ODe�J��O{�q��g��n�f�J��c#.�x�'R�'��5H6��'���'��O���7L�e>jֈL�Z����N`�V��l�O�D�OT�'�?Y���?ͻ9	,�+�̺ p��r�..6��<����?IJ>ͧ�?i��9ɐ���4�y2N�0�;���+w"���ɖ�y"��C�ȴ�����4����A ,;acɏ���c&�ۍ[����O���O��5���C�Xu��'�b���̩�aM�S4p����¦U�O�h�'I��'6�'32�҄��v�`Px�.3e����O^���fޜW��7-�^�S89��D�O♚���)LR����dR�i�^]T�I�����OB���Ox��?��b��<��%|�(�"�n�|d��Y	s�i�I;�MV)���d����'���i�55�Kw��ɰ�If6�)��|�����4�	�	lEn��<y�>��+6a�Rp��CO9o��,��%WO`L37oJ�����4�
�D�O����OV�d�
x�^� ��c�H�x$m��[�˓\��#�i �������mH�h�t���p��oW�?�������	}�)擷MO�����W�8]*�ݽRv�S���b��{�r욷��O�YM>�/OH��sD�/מ�
�MM�R�z�)�O ��On�D�O�)�<�S�iJ��'����{�<� C�R  ך!T�'��6�3������O.���O�� �f�x
�KEN2��H׳x`��ݴ���"�M�qџ�����nC�更�TJ�.9i�5�� ���d�O�id��O�$�O���O1�(H�jS�E���*m��T���O4��O�o�6.p�����X�	`�?dL�˵��(��Ȓu�N�{��H$���	Пd�	�W�h�lZ�<�����Jjܼ;8���#��/vF�!a�K�a���������9OۢQ���E&�h^8����MsE���?����?)�b���̄ |�,�U���7�`(枟\[�OB�$�OH�O�ӧ0P`"��2��m�ȏv	nyZ �;\P�n���4�����'�'DLɓ�n�b��kp'HA����'��'r���O)�I �M��X�2��tp�O�D��@A�^(9�����?᧴i/�Oz�'��I�9��y�T	V�5��(ʿF���'$��A�i�I&i޴
֟��9��`�ELJ%w�F=���	΢a��M�kЌ�g�פk��� !���< Z�NO/c������ҁ�QO '5��q�s D���,�dP�,�O�`-��!ǀV�rGÌ
������3��@D���ܢ=ظp�f�R�����Ak��b��]:C�cr�)��Χ�H�W�٨)��Y��U�����i�!}-�D���14"�1a�ău=�q�$�D �������`�8a
Qu���š��%r-���Íi���&�.O�4�΄3�tt �&��sZ�)	C߄/��5o�ß�������S���<�ӌ�'(5p�K
���4Bڑ֛�Vc��|2U>�?qR�^6xܶ��!�I9Y#pH�S̈T��'=2�'{6,X&�>�)O��d��XCMT%�*�x"l���Za91�1�Ɂ	{t%����ϟ��I5Q*�$I��Z��x 0�D28q �h�4�?��.
k��Ly��'�ɧ5(�5^ �Հa�.&��b�ʞ���ď)x��O����OR�d�<�"� ���Ԓ6�3]
�q��W *5��Zv]���'���|��'�"`˛+��$��Z/�dͳ���Z�2)�y�'�b�'��I�U7h�ИO
V���!��hi�y��J�8�4$��4����O��Of���O��$���ز*�)�h�A�=ʠ�)�Ⱦ>���?)���Ą:�̌�O��*�#0.��v��Z�+S*X�]��7��O(�Oh���Ot�3EI1�I�	�DL����-3$�c��6V�6M�O��D�<qG�:!��͟`���?��ˊ	S򢌪��(Gex�j%D�3�ē�?q�X ��x�����d�������[�8%R��G��	�M�)O�B��N����I̟�I�?��Ok�s�����׻v��vL4V�v�'|�o
�B�|b��[�9��ȋ���<#V��e웶�ċy5D7m�O��D�O���_h}R\�ٗ.�m4�H����'?�ER^hX�4j䤨�2���OFm��Jw�4P#�����5�E��-��ǟ ��_����O6ʓ�?1�'�xҗ�Y��rebG8i��8X�}R���'�2�'�I�n���Je���t�\)$0L=�6-�O<)9�n�B}�S�|�	P�i��{r��\��%@��N �>��U8�䓫?����?�-O�a�Ε.PX�L:���̩�D��y����'!����%��������s�]��12C,� X��E�3�H�:ł,$���	����Icy���7#-���>���;ƢY:In8���i��6��<y��䓖?q��:d�'G��ʥ�k�j�@4�ڰr��٘�O����O���<���l���̟���Ϡg����&�L�f �� ȗ�M���䓿?��M[���{
�  �{%��=d|��LB!���i���'��	�{Y��L|r���1#��11͖,Q%��@e��'���'R��'���yZw\^%�A��� ���U�[Cђ`*�4��d��nZ���i�Ov�)�a~��҇_Z|����QT�y�I���M�(O����OR�%>�%?7-�	�bTʁ,��J9 �#�=w�6� J��7M�O
�d�O��)r�i>�h�B� |!<���Ŷ4�@X�Q�-�M��?�����S��'��_�O��ˀ�B�&���$MV�7-�O��d�OF J��q�i>��Io?)�$� +
�T��,��G��u+������\�I-������Ia?��hՇ-\�{�č��@Q�ɂƦ���5:*���'4���'�>��U��j5J��"���$"�$�5b�1OP�$�<i��P*6�Z��V$8�j$�M�Z�@DϏ)���Ot�$9��Ο �7�p���`�Ud�H$��1p��o�1��c���I}y2�'4��՟2�&dٵK?�d��&B�$6F��վi�R�'P�O�$�<)"�Lަ��Gb7휘q� <Snm��<���O�ʓ�?��l�����Ox�ڐ��G��D�cW
p�V�kۦ��?����䈵�'��tq��55���P�^,+���4�?1���DEsj5%>]���?ט�U��]�c�O�j�T��0!Jf(O�˓�?�����<��>8��χ�\�f�q�<Ǆ4�'?���(�B�'�2�'��X���4?�NY��V]w��BdF�8_�6��O�˓L�:ExJ|�^uV�1д���đ�@�4k��ƌڢ��'�'4�d\��:V��tM ,26���L�,�;�]�\kFN:�S�'�?^0
��%O*d��,��mږK�>�nϟ��I֟,��,߽���|R���?��#
�I���3�"I��P�.�P����'s2Y�0ʯ��ʧ�?��'T��5��Wk��X��Z�h~�� �4�?�������A�����|����5k5j�H0��a���'��:f�=?A��?�����D�'QQ�ڄE5S?p��@��\�R8��a�	���j�IryZw��� ��ה%�ͳ�"�JdI�4�?�+O����O���<����X*�ə ~Q�QbZx��x�"DPi�������ןL�'�[>��I�(���c��ޔ�@�7#������O����O��?QWKV��i���Rt�C*aD���Uo�T���w�L� ��IyB����Q�Nဉܽi�� 	#-Ʉ��8n�����	QyB�ؤAO��'�?A���5dC�c�&tI���:n�xr��<I��	�t��ӟ��f
l�,'�D��
�rw$k�X��'�+�<�mnyb<Y�6�Of��O��)�P}Zw��f�ԋ'��uzu"�&I��4�?q��Z���ϓ��ϸO����7'ӂ-HiEa�{�R�[۴��`R��iZB�'���OR����đ?P�]�4���Ղ���!�r�m��*�I�Ж'�� �Dص?����Řd�4��G�ӪR��l�ݟ8��ƟxGi����ĸ<����~"`ұ7�lx�B*I|��c�̓��M3�����سt��?E�I�`��h��1��B�K
r��1h���o���X��BI��d�<����D�Ok�C�Ә|��Ժ7�1��+O"O �I�6$(�I��|�	ȟ��	ܟЗ'�4�rf�� a�t#sE���0$F&��gNN듯��O���?9��?�pC�e�����|dhQᛀL�͓���O��D�Oh�r\��S0����ڂ2,!��4
t��r�i\�	ȟ�']R�'!Ҫ�0�y�%(	A�u�3iX�(%<��n�-s�7m�OT���O��D�<����f���ޟ�7��}ͦ|	g�OD�t!� !�Mk���$�O*���O�X����sӤu����\)X�Mǂ|]�\ˤ�iLB�'��	���믟���O������%^�T�85�jJ0�X���Y}��'R��'�l,�'�U����0(8��ň.�:tq ��5�֩nZeyB�p�7��O:���O����u}Zw�X���'<}�!1��:\$|��۴�?��)%Q�}�s��}Jq"�%[�D�uKƞ:d"'+¦A�v���M����?A��R\�t�'q,��� �X8"b��d&���Et��0��2ON���<I��T�'>�%3���^�Hࢋ?5��Hq@dӞ���O^�dʋ1���'^�̟|��,m˄iP�3�TY��N�2 "Xl�cyr�'D��yʟ��D�O��ж�H<arm�I���CYl�LlZɟ̨!���$�<������Ok�/;i��q���[�@Tk��ɧ~����{y��'��'��5���^^u ��P�d��<1�	�Jvvu�'��Iʟ��'�2�'(�[�@4P|��`�o��I�
�dr:���'	�I���Iş �'@<�A��s>=�`,38��S�+'�HdR�sӜ��?!/O��$�OJ���2��Y4m�Y��*L/(�tͺ�A-@\Jn�`��㟴�	Iy�^�MR`�'�?����m��ĸt�vD#�bK�9Ϟ�mZ�Ԕ'Z��'�rJH��y�U>7������EY`g��[r�;i]���'O\�,��%�8��)�O��d�6ԪC,�H���Dh�f��i�� �P}��'Rb�'s2qٝ'��s����;�=@�"�#oo����a�J�2�l`y2�����6��O��O&�I�S}Zw�X����Hn��Pd�5w^�޴�?��0�����?/Oz�>� ��D��
� |�0�S�T�u b�izpR�}�@�$�O��D�����'���.:�(�!�ˆ0�VA��͞^��(b޴*b�͓�?�+O�?���ü�6�Z�kБ��W3}��H�ݴ�?����?i0+5��Imy��'y����/����Ӝ<��,S�"6z��f�'�"�'�*����	�O�d�O��� �]�vab�c�&G ݈y��k�馽�I�^���O���?�.O����N�Z�� #lDt8�LK$U?���RW�
��c����՟�������ky�.B��Y�<=*�(��f�`qp�>)O���<���?1��'�N��$�̛`O��`΋93&��Z�K�<.O���O�d�<1��ܩ1����
Â`�Q)�|r08`�@G Z���Q�d��Oy��'?��'�$�'�}�aNQ>P����W`�O���SQ�s�����OX���O��.�<�k�[?��I9E��z%aC4o�,���-q)9��4�?.Oj���O��$�R��$�|n�����xg�*~�FГ�EܷYnD7��O��d�<�������l���?=㳈U�*�ԑG"�
<Q��L	����O����Ov��A8O���<1�O}�̉�(�:"x`)p��3$�]k�4��$35�m���������S ����X!֌�!??pt{Q��g�:�ط�i���'b��'�r\���}B�ؗv�Rt@En�#�0�qA�ަia*�:�M���?�����Q�,�'����S�4��H��˯^�|� -x���
W4O����<�����'Z:M�g�,	5 ΤZ�r��'I��'�#��'v<�����O��	��yqG�[M#$�V�L]@6��O��$�O�p	�:O��ݟ���ٟ|�W%ʛ=ň���az-J2����Ms�����a\�@�'N�U�D�i���e�
"d^鰧�h�6���>Q����<����?����?	����Ċ6 �>�%K�,x�p��;Q�Z���^�Iן0��]�	ן4�I)y�@��%k��5���)A���Y�p	��$������Iڟ��'�z ˱Jt>e�$N�9�M��m�M�6KD��>a���?M>i��?� ���~f�%���'h��D-��K�������O��$�O��\z��0���4��2��])֬��KXP�ԭ��:�6m�O��Ov�D�O�]C�;O��'F�mB��̚B�-p�N�%M��#�4�?�������,%>M�	�?-B�#2ĨX�R,"��x�bK�ē�?��x �������4��!=�D]#&倥D��e�/��M;,O����Y��)A����d��n��'ĔKPb�5z�%�֏�p��!��4�?��q�Z(�����OP�����
0%F�ӥm}pqP�43���a�i�b�'b�O�*b���Qǐ�{�5s7���.�������M���W�<�J>َ�D�'�����N'�p�눣0�:��b�q�����Op��XS<=&���I��<��4���t�^ }_>
d\��-�ڦ�'�41��~��?A��?����K�0�ׁ�}!�6TP�6�'���4�#���O6�D"��ƪ b���{�tY����wLӨ���m\�<Q��?1O~��kO�on$D�Rć�e�@0xf�ɪG�\P8іx��'�b�|��'�B��T�F�X3 �<w���1c��[��Qڥ�' �I͟D����'KDm�e�~>q#&�G�}T���H�4*VT8	�c�>����?9J>���?Y����<��C�$>�V�!�훹+�f�����I3��ȟ���H�'��:�:�Ϭ	��y벦�5y����*7?��`l��'�l�����D�ß�O<��qEM�a6��gŀFq�l�B�i��'��IfG�@�J|r����1$��J�iBh8��R>��>�+Ob��6�i݁跨��v	��b���opr ��e���O�9���O(���O�蟔��á��L�N��.ϻ#DxAr�L�9��Iy2$�-�O�O����VB}�vH���jZҼ)�4�&DP��iw��'nb�O�����Z�q�Dh��i�S�$�{g��4�@�lZȟdE{��|��'���OԪ;ߞe�G���`C�!qӶ�D�O"��3C)�����O:�əw2��G懫i>,�fۚg�`Ҏ��d��ߟ��	����Ҝ������ک|6v�(Ea
��M���8~bX�-OP��OR�|"gG����BV�ϔt����k�*s\�O�`B���l�	ß��	ny��-[%`����Xt �;�jC�����m6���O����O����5K����X3�C�#�>�{p�!Yxc��������I˟@���f����0�|��pm�-ALQ��� �4��m��@���\$�D��qy� �'�M�@�'ҠLsG�0YV�
�&�X}�'���'h�	�ȕN|ڃ!ԃ����+�mS@�a��3����'��'g��'9�ˊ}�,1%^�C�%O?k�H�	�LA��M����?�/O�M����D�۟��5e �j��//`�
�+ي��݀J<���?�%N[C�'4��X�'H���0���Sd4�S���hO��T���Ŭ�0�MK�T?A�I�?�(�O2��,L�;:̨PD��q�8'�i�"�'s�����"�S'ㄵ�M�)�6� c끉/�p6m��	�V�m����	������?]Jl9�&$ Q0�+Z���ٴ5���Gx���O��1�,]�Ę2���^ː=i'������؟��	�S$P�L<9���?!�'��J�g�C\�M�7f�,z44��}�`���'�b�'1�+=� H=�H�.�p�+uMJQ T�i�r�\���c���	}�i��Kg�ħ(/�P��.6�(���>i�	�b��?���?/O�8�5��u�&�`�S�`��a�e�C
!3ް�>�����?��T.�]B�iL�M�$��a��vA�����\yܓ7�$���/v�k��	�5ڰT��i�p�4,�+Zh!��m��1c�2_�<�%$VqO����R(� L��@�P�i2d��`�I-
ǆI ģFF��C�^�+<Cp|PB������ 4{���G@	:*]��s�4m8G�&w����H-T��=8���4vF@Q[���1D�ڄ��j����'�X	v�0���-C�d���O��B,��2r-P� ����kP����zDV,��������O��C�x����%[P�����tS>�y)ǎy�X����;�����e7}r��R��q�	��7mZ�'N����A+G����s��"E�>�<�a� ��O��hem3}�BA��?���h���d̦0���Bq��2�$K��\
S~!�d�~�b�21��"$��ʀ⋸Mfax�)ғ�0�#��'c.���گ/�|y Q�D��ȟ S���(Ko����џ@�	����65�����W��!�
�U� �b�Ŗ~殍a�
�t!��v�g� s쨴L�HA��Y#LS�:�j�3%�zl�����q� �2�3�d@"/ yK�ȏ��p��M�.1�b�D6?!֩����`�'���҇T�MA��Y&!��m
����'���ز�Κ�hb��axp)��O��Gzʟ��ں}hVNءM���"2�!9(��+Kj�~Z���?���?aV��4�$�O��;E�y���Ӷ^����#Ԛn�E�W�S�>�7	�� Ta{��=���S�t���$�AY��p���N�ID�=lO�����Ŧ%*�1��t
t�c�+�+r�'�ў��?�&��,��I � �
�v�K$�^�<)q�Z�� �jÏo؜�w��C�}��	OyrČ�,� ��?��m�b�p!ԯ��B������?)�Nk����?Y�O2��G��9m�h#����q�0������O���� ?��x���*G�hqѳg�n{>�	�TҪ�e�,;���y�gI�l�j�񄀔�r�'��A����4��%c�+m��5hc���I0}>���_!���h3�S�BNC����M�6II/)�ty&��$���'fQ�<9*O��3�i���u������O���I�'D<�8�.�(E��[�Ék����'�B�ӧOV6�5���|�'P�Mx��S�2rl
�d�g��qO�Ы� D ��F8>���t�6pN���t�Z���A���.�)ŗ>�4��֟�I,�M�����O �X���:;!Fa;�$Q�6��'���֟ ����+�dE:a�R�S��ѱL<�1� �%c�x�i��7��O��mZʟ�{r- �-z�ԈV�O�4i����<�M���?��)�b�s�D �?A���?����DI�!!����B�Әc�Nh����8͘'���
ϓeJ�bff�F(��d�� F�4�=	��[x���ԅm��ݨ�O��ܩ@����L����)�3�	1VS���7��������H�!��TU�4'�Tʎ乇)̗E�����HO��(���{���pէ�+È��Ĉ�A��e�r���,}����O0�d�O�����?�����H�3d9�qȑ<��9J�g��9��EksD.��}BAߘM��hɓ���<Eɠ��`զ�JgO
��}Bo
U�|�	��u�P��V<)��Q���?y���?�*O&�$2��N�x���Ϸ�
��었�C�I4J4��Q�ޱ}��<Rf+�JFzb����O������CS��I
(�vՑ��<�T�Q�JY�8QZ��Iٟ��UCUٟ�	�|7���j[-`���0�$�A�l��X�t��� A���x2I!V&��LƗ����0F��Ç'B;	��rѮˬCrT���ߞ�2�'��I,$#2��''Ƚ�L9�@`
�I�c� ��	*Q �(٢�<r١�+�\�vC�ɕ�M�1i�0����B�^�:$ Z�M��<9*O��"�/�v}��'n��.:k���	>m���0��%7l�@`�β!�>���ɟ��`¯7*��*���&^�8$��S��\>��g�%Z�R�`�mN.J��	�<�'�r��oߐHu�]�B�|ۑ>��gH�;&b����NM0o��`�%1}e��?���h�X���=�pu�Q헓^v~���fN���C�I�eyV�ۣJC>JMp��.fSaxBM ғ2>��c/_-_���HCHv�n�!òiv�'_�E�(�:y(p�'���'�R�e�Q��ʖ����@�݉NdP����GE�m�H��	%	J��C>��2⎨~b�\`��8<O��K�F�6Y������G�M�ua=�����|�Њ	�^��7垏g)��Чe[��y
� << ��D�jK���,l��� 7��ؙ���ӮG�n�I��:V��{�dE�a����m5���	꟤��̟�A_w�R�'���:(�L��*I+!�)�0���0O&�sħD6
4HЦ�y|tа�ȧo!���6
]�1C�#B.�h@���
 n 3��'�B�|��'�����:=H^����V�V�IQ��I�Y!�d�
[%�1��.j��H+��"]1O@��'e��
��b�O�D�,��=3 �E���)I
ɄE���D�Oj�2��O��db>}JC�0T�F�H�.G�~⪍�F�h��r�&rjXด�د�p<!׬�A��P�A2U���҆8�
%R�ǹ\�3T�i �x�(��?����D��ҝ�Ć��1�JA�kݴXd1OF���R�KtN�8`Ӑ;�2Cv�T�*G!�d����I�C�0�0P�wjH%َ}�W�b��E{��)@�u8�x���\=�9�tk�")�!��0h�F̓���b�H�sDJ��zx!�d@�WĒ�qˈ�H�h�����5ht!��3z (�+�J&RuԴ��$�(_y!�ĐY�y��3V�:�E�Oj!򄈨;��0 ��g2�r�b�4*�!򤝀7�8� �d��q`K^�!��ņ	�.8��`Ӕ*t�Р4`X�3�!�Ě�-�ӗ��nj�0���T]!�dS18��m��_�s�@i����-	G!�dϩ7L���+��R�㗆A�B!��*u��t�k��zW�:!�D�*MC���� �b/��r����!��K�Y�rq7�o�,EbA��;y�!�]�}�dX˒l�0)��,8����!򄄁p�\ي�W�O��<b�$�!�dA�AV$i�I,EU��)_	_�!�[Ze�i�E�m�8{�V��!�
� ��aK�'Ez9�FiϔO�!��ٽ&�^e�b܉}T
�Q�+D�!��/���80���@�)�F�.q�!�"T��8J�IM�I)65˱@̷�!�۹]��i���Q�P|���d�U!�ܩu���f��<Q�(XP�I.x!�]�2}���̋�C�6�"��Y!�!L� �7�C(i�4�3.�Y!�dZ�lr���E?l�p�d�Z	E!�D̘z�;�޽oTp�i& T��!�䓣GN ��䊟5|�@B�R�!��1�|a)��Q-(�v�h�(:BO!�/�tų�aY�g���SH�9k!��N�8K ��[N�"p&� �!���3����NN�ut���増�=!�D�W!��J�ƣd҈+�L�-s�!���:U��5 �H�98g�X��(L
!!�� *=:��H�n��p��U|w!�$�P�̸��	+�y)T CbU!�dO$�*�[hZ-�,A��1'�!�Ăk�x�)�o�<֌�VPc�!��NPցXE�رE�z�mߐ�!�$�{����/ldp�o�F�!� �~���͖*Q\�0�!/�)�!�ʜu7���ŠM�\���.�	(�!�d
��9��G�2p �gٲ\!��,x�ʤ� nO�N������ȥ6Z!��.Vڒ`�Bgߵ#���a��A!�ӲnĦ�����$�h��5�!��P��h�ٍW��ړ�Y�F�!�M� �@B� ޓ��9An!�$*]�99��Y�q�VŅf!��=&<-B��&��̣�c��^P!�� H�! d�� w�hk��^Ej(��"O��Q-̾�$���-*�E��"O�y)��R:ʢ��#j��;"O�E�f�K�7]v(����C�� JT"O`a���أR	� ��U�<��ܨa"Ov����Н�h�*FHē�R��e"O�h��H�}5�л&�݁S����U"OZ!QU ə�d���K�/[�|��s"Oh�ab 30�x��w�ޤM�%�F"O�%HҩFt*��Й��Q"OΝ[W�W�L��(6j�'X.�C�"O��ɤ
��D�� z�	���`Ad"O�MA"+�A]��b�B�C�K�"OT�##-&#М����{���&�'��i{�収m���Y�j� ��]y��W�B��4^������]E��)��	�C�`��&C��>���^�&G�px���T�>a3�
N'V����V*������:��g"r��:s�܌@���4�Q��/Ĺ�ff��S���Y��Pp��g$�e�e
�7��B��λ_�z��ȓR���g�����ZB͝T7���O|�5��?�~dW�G�`,$��E�6TF'͡MZ����6���	t2��-��3\ԡ��C�$"��X
ci׀.88�M�z�dI f��E~���i4j��%+�1�b�:� �r�t���
]��Z3+�gi0���5+�FI�>@��8p��!XX��Y��v�աk����v8����o�Dr��(a�^�af8�)�>ѓMG/�*,sC�YL9���q0B.U�L��/��P
r��$,U6O��E��0H|���DH�,8���M���䞮&Wܐ��V<W�(  6.H���	�Q�l����B��@����$���~��;:�a���$���c��5y���D�^!1O���@�0��L�!/
_���Z�����'�ܭa��6#.����J�o����b�A�?G$�(�\�K�υ�a^�'�}��N�x��Kd���x����ϗMn����B��fX؋�����O�pC�_\���ϫ �6���D<s<d�PCc�?	�a�9̄�1�K-u�Fa2���K�'����ƈ�{rH�aŊM�/`�c��n쌙�����K�j�a��]�f����(�$MY`�R� n��">i�$@�@d��!̼��~�<ݘD� �%���C`�|��Z%gL*Z�� �@璮#��(�f� LLĻ3�d� �Ź7k�K�.�86a��2�1O( ��ML��Pa��>ga u��-�)bք�*3��8	��0:�B�
�-ڄP��+��b-� ��f*xt��ئE5?�(Ҋ�0=�0n�6m��v��_���e�n?c ��3|4��ROU�mKvh�D�V�'Tآ�7*�����:y����'�@ʖ�;�P�.p��e�(��D�{@�DxܓO�Z 8m�Fx�;F�@��T̼a���H�#W� �B%��I��A�,z��J�' �=�"#h$�c�<�&+,(��$`��W�.T}  !�I9w-��*�dM?R 4I���Ģ>1S�J�F���!AP�tll�DI\7��h���1�Jq{�.�i�������(o��D��i�Y���8LOfY��EK�-���2�N�:���@�OLo7�ꅩ7�?J�fX��M[�m}��0�J��h``���=H�S�J�S!�DR�",����ʙ���㠊�+�$d(�J��਽	�Z;
�1O���JJ"xͲf2�<�TK�:5��� �Wx�b��';�\��KA1����$�B,�6 *� ��\��<�<)�(��v�=7A�(�,5�6g@�1�k"&TZbh�bǒ�F�x�F}2���b�RĢQ(��k�,�i��q!�A�K>���Aŋq��93@�;B�t���S��T��gA}��� ��Cȕ���T��a�a���ZƦ?R.B)
Sm�L��TҁӪadJ�ce�dI9X�B�Bpns�R��gE>q!�{󄜈%=th�A�?:�Z�s�̘�L�ȈZ�K��Yt^��C�T>#�1O^��G�DcG�� 1�H�`�ß� �����:�����'qbb�h�;f�1b.�1G�n�;p)իMZ��<9t!ŋ�Z�c"E Fa2q��\̓A���(6�ܰ28i�lb�(|G}�'�&��X�8h�d+"H(}@'�qH�Se�4`�j +DK�t�Ji���u��Lb��4T���	{���� �=9�F�K����z牍Z����7dU�d����3;#����yKFc���dX�O:��tg_,�.P�\ �dH�P�:�"~F���P��AOM>Ĵ`�S��8`�t�ORH���Y�H�RI���9O��;?�X{����L��"�^��L�'�1�2�'�&m���&s����%��:ƜS� ���'�ƝQ�(�F�Hl0�g�a��S�:Id���D�TK�[����J��8��L{����L���Y����
p��3� e*2�7���Q`,&���2#�A�b�Z�s�;P���`B
.s"��T?��$�E�D���Qi�">��%q�s�������*�R�O�D�x��Q?��?!���$�.��������k�In���ڠ)d����	O$�Z�UI�5V����м]�E0%�� ���ɬG��CD��k]v(Q�F�L�">��@�3<��u�ۮC�j�ju����r@X�8(�����!�hxE�B�<A���c���RV* K�r�YP� �<9Bf]%%� ��"W�E�
qA����h��HJ�L�\��08 ��!'d�i#W"O ��C<S�l��5�S �(��#
i0�11�F;C:2u�B<��g���6,�G�_�
��|��,�L�\͆ȓj�QŏfA�B�� �3q�EѦ-����$���{�,�_�"!"b��rU�l�E�3�hO`!Ip��Hƈ��b�L5j�v`´�JB�X�YҸ�*�ѷiF��j��B�<���+��1�M��oX���6��Ħ�g��fB�H���ZYFp�$��OQ>ט!E�z��Ǎ�e�mˤ�#�$B�	�)�,aP���0c�䩁��3.5ܐ�v�&�?1�C�:8��<�V˽~J�E(�I�R[H�P�[9��0��=�����7E� 	Vb�W�L��`��3v�B�҇�E��zA�DL��<a%T��=�S�ѭ/��. �I������ܓ�`�
g��n|sf��0�0M�*#��͖���؂2�2����~�<!�"H�&���,�QaFm�Nr�� �d�OI"�n�f����)��y'n�4-`��ːoV�/��aW����y�Lȴ��t�h��;�(1˂&ʓ���5�hP`�]�g���ҩ�C⟠���<�1�a�<cLx%KV�/LO�2f�f<$)��]8n9�D�?�u���4H|����冣�4��tKI5>)H��DY�jHu�\��#�X"\I1O��'�H����D`q���A�Z~��DX�s���:2��Sg50X�Q�daKO�<��E�T��4c���]7r�1�i�.��!I3$_F�na�q+8w�Vy�bM�PˉOf2���w�h(�v�X`p��I�%����
�'�be���W�^4�ą�=W�&0�6!W
�>�9��T#�H�q�b.�bd���7^c�Xa�7&��`� =�:\:�<lO ���C���Ѡ{ր��G�	�lzV�Կ%��I�}\��Ѱ��d؞p�'��uh� S��	�H��H9�ɴ�XpK���L�O���R#�	_�$$�4K>���'�跖�1$�L��'�
qF(�[d��p	��OQI��3?��ӛCR:�Y�/��6�[���P�<��,$C�0�ԡ�(�ܑ+V$Fh�aq��!�:��1(�&����!;=��4��H�az򃈭z�X�A�ST?!6$��Ԡ2�M��ԡ3��^�<!���>C���x�&ͣL�L	c@$�A̓�( �(�3b��~%���p&քYذ�bQm�D�<9��Wy�$���<��LH�73�@s��0}�#������/_2�1�D[�~q�%i#L�&7��B�ɡw�D8{�׵Ey��P��B�y�C��B�\X��'��`ѫU�w� i�ՀU�B���ӓP��i�&V��hK~�s���,.8+��ξ��C��-a�x4�aE�n�|�ʍ3mrb�|�ƕ)S�����7Cj��adHKx�Y�3�ʜ7��C�	XXJ�F�Y�ʡ�R�[�6"����L��T?����F��O����9"��Y�S�{��ء�"O`Ȼ���4�2E����/gP�����;�<`J�&KDX�P� �Jg$���	0e��X�d,D�<Z��x�D3 �Q,%�J�F�)D�X�ˑ*)0:Т�Хd�z�qU�$D���Cl�T�Vĩ�s_��(U>D�x��@Z�q~HJ��O6G8|+�:D�h �
�(Wƽcb���d����3D�8�6͎1W<�{`K1�xxE3D�X����	&�8�r0�
0r���Pa$D��؅PWƶ���ʏ7����#D��B&N��y�}�pM�r�~(� =D��9gKO�z%��/G7\��c�O D�H�s(9x���beGk�J��5#D�hS�G�2q��A�=N�J�cL!D�� ��sB�^���yDU� '��s�"O(�,A��h�4��@�d@2"O�3+)u`�Pᣃ��Ҵ:""Onq��L�;RY����Y�"հs"O �6-�6u�Pp���_��:4��"OIcэ�6_�B�"�mɑClB-@"O����u&���vW7Ee�E�"O�(�V��h�@a0�x}ztp$"Od��$Ř�G�f('�\�YX�a9r"O~��Q+K�&�z�Yģ�)/G��e"OZ�Q���U!����@�3V�kA"O<(˶�Xx!��ă��*�t�"O<�.�4k=�`	P�Q0g`2*Of=Jf)�Y�vug)3T�U��'��*@��$?�T�Wj�R���q�'_�H�eD�<��ř4J��I{U��'񐕛u)�?���{d���O��Y��'�M�*��F¬��sa��^*�*�'+ u&����y�DV4��5�
�'��1��)иKj�"���>����	�'{T(Ar�:><�F�K9�Y��'Jia��B�z���:�/��$��'�<�X��S�NA�0�(U����'��d���G�[��E�2#OH�m��'�z5����?5��j�ŰA�r�Q�'M�P�N̪v���f$:��p�',�T�6`��3��!�v�:�͸�'U���,G��Y#�� 6�����'QZ!���D�4<�(����-K����'@��v��"z� fR-9�~�Y�'�jqj�G;L0�����"O���
�'&=��M�wzb��P����R
�'R$�6_Eb63��Fˢl�	�'��Hb"O(nlhzU�Q+�lI	�'�pe�v�IU� <D��ya���'��쩐r^��b�^����c�'�*%5JT���N&r����� &�yb��w�-Xq��h�D�1���yN��W�1�O��bZ%���ybJߨ����& �r4HIK&L[��y���^������bły�%�˱�yŗ�C$�,i�/��% �ÈA/�yr@�c;��I��&�"${#���y���sN�۷�J0tD�r @��y2邇�,k��+|m*�
���y⯍+|
�Bi��"�i�ѢG��y�'Ȩ�t`�@�r{İ�m���yRn2ŀ�a��Z2j�z%��(�y" �b96E �닼c3P��tǌ��y���&8���6�73�Z`($E*�yr�6U&�y�n��(��=+FŇ���>��OL �xC2Q�3ժ7N��蓨.D��PoFP�Jf��/!�pY�(D� �wM�3ˈ�0mʘy�d]`*$D�l('_�\���F���R�骁�#D��H��U������Zw��ӵb?D��ȰgO'���&�L�+���Q`<D�x�U���ITDX���n͢1�u�9D�8A�)� g�p�@
Ji����6D���D-}�|�)�k�F��De�2D�#F�Ϩ
l�5S�AR�2 (�5D�<���**
Z)c[�W�ؽ�`�>D�(Z`I�j�v�Ȧ*�?���2�:D��(A�v݂PZ7꟪!������6D�� � ��<|��%.�2C��\�"O��)Q
�l5��p�ź����F"O������JB]hS���ԬѴ"O�I�#BJ�d���9vYX$"OH	H���%� �����$&z��"O�J�J�[|DL���Y���"O4e:�+���Qz���(l�ly�"OxY	tn�A�a�1�T;di9b�"OXi�e����A�F	f���V"O�mqf��,�p6��
0RLyq�"O�-cE�?rf9pk��c?�@�"O>�At�	�4 �Y	£�28�nm)#"O�J�.��L�q�O��dX�H5"O� ��ƭo�0m�C�C"Rt�L�"Od؂�5{�a�d¦9n$��v"O2Y�!##�\)@�B�kU���p"O�$�Ζ8t.�i��ӁtCN�qA"O�a(�)�!=f�]�5�Op��k�"OJ�b�ˈ���7�4c$l;!"O�at�B�F��	��/\�OHZ�J�N���������E����/'#&�i���yR&H�+"�BeCL� x�B"ˁ�y�b�!T��욤�����Q[�Py"kĎG$���s��%5�{�Nz�<Y"���-�r%8��Z�u�h�ꤤnx� Dxb�00R���DG��e�"5�yr&ĿK:3`ݢRT�iC�c��y��G'[�j�j���L�ym�&�y��'�NL� +��A�<��'�0�y��O�+�Vl�k�Ks�9ar�M!�y�@��|��o�x�N��P�ִ�y��A�KN��� \��W��y�ؙ2(<S�"	fZ^<*'�֏�M��'�3`o��oQ�����+��m1�'�i{3���%d�
E�
����'~N�0qL�0A�!��@�'ln��	�'q�eY��W�*��dPq��W�`	�'��8���S�LR\0�D-V�.8�'Ѧe��3GP"�f�S�6ʺ�[�'��`�qɄ�R�F] �ě)q�|��'7,4	�HҫA��q��⇿ P(p�'e�����'>��L�a��8$>�\x�'T�3&Ǜ%�hhI��!��d��'���Q��N��'.��m��'����gJk\�a�/�z�P	�'�idh\�x�ĭȆ��@հ�'z�Q"@�H� X���e�B ��'�z]�!]H�	2��!V�̀��'�@ 0��E�F���釠b ����x��I�(�����YZ,�u����y"E��y+ܔê�5K��|h�����y�,~�����Z]�x������'�ў�O�����Lf��a
��P�b�4�P�'��(�ZM�����Bhc�'H�ظrJ˴|�	"��˸c�,qj��:O
��գ�:���$g3,�4j�"O|e��nKiʚ=�;I��� U"O�Q�@�V;&dxxY������'l��`��H�6&��1�/W	i	�DzB�'_�ܨ5�A�b�;4B��T�{���2��e��i� ��"���L��`"O���c�& ��P m�Kv�
�"O�8���." �8�E�>]k^Lt"ODa�ȃDy8�q1�X,Q:-i"O� �����M&~�NLR�)�,O2}	#*O�x�W��j�αP�!Up\I)�'٢`j��4�+T�O!Q���		�'u`1�Ck�8F�.�8Fl�D*�Z��6�S����j�\���߫T�t�Rӌ�
�yb	D�j��!F��S��r��ɬ�y���#�l���M�x}�ħߠ�y�F�{&�d�Gi[KAB���D��y�3h���'oA�J�<�bް�yR��"^��xǖ�G�ly��˽�y�NQ�:�p�ch�%=��ݻA�̤�y�/&-��`�`N�@��xpm���yB��0���!O�1����*��y�+��r�P�!����%��h����y2� d��T[R���$��DC ��yR	�#+��h �-�� *�i%┷�yo�x鸠�ri^�L4�G�.�y�f\t��F�9|N����AZ��y���MCt��Ȍ{�Ne!��R��y҄�|D����J�i���5�U8�y�O�\X%�b�17@�a��yB���L�)�f��2���	�y�H�o������6�)��P��y⡂ryXi&���4�d$��Y��y��JC�D�IfգyF�($IL-�yB���r��3�[>�$ЖN��y������ۢh��F��Qp�Ț/�y�DD�JITp�������y%�Ǘ�y2%<L�J)���I2b�'�y��ԣg���R��-)7� �����0?�*O���g��@R�H /=Qot�"OZ�Y�ҹ�����ɱY�`(!w"O�a�e�Qݕ��P�{��83&�G�<Y�dξ���� �X� ���[�͐E�<���	0)v����A,S�ċP-�j�<��?��PW��lܬ���GL�<�1	ߴ$.P�DO0hb|��*X_�<�����ZvD�Q3���.� �U�<��+K�iߎ�x�e �w��!�ɖE�<Y��ڒk��m{�oޟU��d��u�<!
��V���!�J�z�h�#��Y�<Qa �9&b���λ_�d���V�<鑋E�n�x�q�K�%���0��	R�<����o*��5�ȅKn8ѱMR�<�'nƉJ␩��|�b�)��r�<9��D�Z�KcBżFތ)���t�<��M�v	4�b�B�D�rQieMMv�<��M�=����nB�vu���Ee�r�<AdC�~�h\H�"�4��8��En�< )�$:�E�ĨWZPxK��B^�<!�3�Z���%{Y��2G*A�<QtD[��DT�N�h>�S�X|�<���X��6�ܘ4� �3#��{�<�jF�1��p��P9#�
_�<!���T�9A"�7Bz$� V��A�<���Flᮨk2N�f]�P0f��h�<)��5\�j {�S�fm2Q��fCf�<��ݸ<2�9��.D(.(��X�L�c�<���P�pxE�٫g�B�В�`�<�⫝��@ź�Kר-t"�!%�^g�<9큮!��Ja�էB�\)�`�<�J%1�0)rM��U?z�Іs�<15�s�q��'�X�
c�<��:~���j�UIj��uU[�<� ��@�����2�(�W����"Odѱ�l�4u��A"'E�E�¸G"Ox��DF�3d�0�£]<	 �xC"Of�y�c�:,Y����$�	i�T�be"O��X��4���â�(�(�
"Oڬ��ˋy�nl1�/�S�F�p"Oje�a,��U����JB���#"O>�bF��G��+�B�+aƼ1�"O�Q1�&AnZM��V�]�A"O�$JքؽP���a�@��s�&h��"O�E��KS�L���eo�-�D0C�"Oj	࢟�T��ʦD�/x�2"OB��T��7U�]�$�<x}�"O�� �X�W�D���t��'"On��O�pO�t�UI��%�[�V"Of0 �XO�"�G�K�0�F*O��q�逑z��X ���4Y���'<�4�!�%h�Z4;�L�<WَL�'e�QA�녋b͘�`�Y+S��ē�'R`LP��è%�V���f�=q
�'(����hL�zuv��V����`��	�'8�8�oM8n��tk��T69��
�'���z�H�4H&4h���K+)����'���B�f� ���i� \ĸs�'�����˄!Ξ���Z�$��
�'E�Qdq!Dh�G"
fdQ
�'k&IJ��ܢ+��<�d;��]s�' :�P�E��v�����@oM�5r�'��sD�#/pds#�/c+�	+�'��Q�m� cH���bE�$-���'R�*F��GR�����0d��'v6��0莥-���@"��w����'m*��O�=-�xA�A�h����'!`p�v�U((��%Hg Q178����'*�X8�Ƅ?a�`��F�/6�`(�	�'F2�c�͛7�*1Z�	����	�'HL-0�Nٙ]�Le�o�i4m�	�'�L��֪�4~�nu"r♐��r	�'8,��c��4{<�����A[	�'^@,�B�F�"����@����x*�'�����ĢPb^�٠f��h��1�'O�#R�2@{��k𡏳�*�P�'��U�fN� ����j=u:����'vz����p�P]��M�?x��c�'�I�&A�=�8�I��5��(�'wX�dl��n̜ Ǧ�}´��'�d1��`
�̌�F*݄p~�i�
�'u�r���)jdc�o�|F�	�'`��陾Db6��5��ml����'iV�R��ܚljpň�âW��I�'�$�;Alݴw4�G� b�9P�'Uzq�M_4)j��vG4i+����' ��TO�0B&Y�����e����'m�u�u.��_,��h�pَM��'���r�+�G-:�O��9�p���'ppQ�k�[b�	�MZ�r�'UȔRh��d�$M��b��v$��'%��g[�j�rIP K
����'f�[�_�G6��"7Ϧ(&���'�Xq��T�`���v-�--.p�'U��DN����3/�O_�i;�'�~�ض�yZ��I�c�22@�t�'�4���;u�h��+�!0nf�'�x��LܝL� �H��$�"�K��� �qY!��!.6��]%J��""O��)rF��8@h����Ϣ��� �"OX �����Yd���	�/��ѓ"On	C�su��U�7}m�"OҤ,וl�F�!���W�L��e"O�A�iX��[��R�Xk�}�<�1���EG(\���̓<�TE���U{�<	�(��e�ƴk�G�8j�p�F�t�<�#隿q�h���u���Ze@Np�<n�%^y���C�N*���AF�
B�<�Q/^&	� �Y��$�\U�Zv�<i�T�g ��:���#IoZ}�"K�p�<��iQ�=Y0���>��Q��Gp�<�A��j>�����Q42�Fa
 B�T�<�"�J<��{/B�U8��ׇS�<Q��0X=�S0+�*�+��N�<��l2[$�n�-"�B�Ka��M�<�cGУE۔$�TL�d�tHs��
H�<�v	��<��Ţ���O�6�� �G}�<���57,D��G�`V�mj"��|�<դצsm���AO�og�,*�D�q�<���&Zm��X�Á�>���+�A�R�<�d�72��u(��_e�e�P��P�<a���~�hڇ�@� 0�]#�I�<9�mZ1j6Q`��_�H��ʅ��@�<��bͪh�⭸� :càQ�Q��S�<QK#,/�� �B�55��D��	O�<YQ�C�VT��!dgX�XS���K�<IFˆ�@ۚY�p-8[�� I�<�ǏڂZ���i��Y�U��P�c^P�<�C/�&4���
�Vy2Uz�s�<���VZl8��_0���S�<Y5e�
&)B�.�5{9��\N�<�B���T]*�S���u�TB���s�<�c�۱a�p��&EV�[H�����u�<�U�_����
n�(S��E���Wu�<)Ef�?��5������ ��q�<��LX�\�V	d��
Plxs��x�<�qj�.I�D�,�2W��u �Gu�<!�m	2�X�1sk۰�2�+�WG�<�N#�F913��Yw ��w��y�<�r��oު�ґk\ P,mzծu�<Y��h>����Y�r}"�bKo�<�O_tA8�K1�߿a&�tҕO�A�<�f�9k��JǊ�"Y��Y���U�<�Ќ�;b�[&�.��T���l�<�E�	��|H���U�&�a�#�T�<��K8M$�h1mȗn� ��u�<�6���'�L$�1
)v��u*�o�<)3n�W��:ňM�A��k��s�<YV�BК�j &A����R$�n�<a��2&�%k� ٧���P�L�g�<iCl�,-sb���^%YjY�ï�}�<a�)�Onu"Vk]�UP��2hu�<a��K�|T�� Sֈ-�7%�m�<�e��!�h��Tۗ*Ɍi{#o�`�<�JQ�*=��@R�ks��jS�B�<��BŲBT�:���A�X��J�}�<3�C�.1�� iD'��E�w�<E,�G�@�wLJ$SĘx*#GJ�<iԩ[�t0ѹ�׹o��mr��[�<q�,�p���g�2.\�n]�<!͞	;I�|@T7%}��a��<�GK��)��y+��C�����R�<� :��榆�;�jHÀB�&��lI�"O���m�uz��"�"(��H�"O�h)1��G@ ���A©A�6�B"O]bb�,{l�	[���¹	�"O^��7��qB*9)�/�%(+�I�"O�M��ʊ�d\9��Pp�d��"O��$-Εi������H^��C"O�Ԑ%NQ��@�CeRL�j�"OB�8�/�Cpz�K����2�{�"O�@���&�X�r`f[�|�x�P�"Oz�1bi�Oo��ðĊ���e:�"O����]�|�҂�?�2�2#"Oft�P���Z�Q��Z<�(�b�"O�,
�j�|*@y��J�qg8q"O ��$�?�\��hMOt	7"O.�hHm��:�i�{C��"Oji��%ӞF��t�ӛ13���"O@!���?[2p��@��Jx�"O4P�c X+��;�٘d�̐�"O���B-^b��̓V&1\L�"O��c�ł�2��� `jmZ�̂�"O�q(���hS��s�	�n2Ir&"O�0Z�%
�z�jϐ�6O���W"O�� f�5�P��ş�(<P%X�"OP�SS&�4b]bѫcW�5<�dI�"O��p� �d ]�B!��p+Vmj'"O���錵|�8rb`&��c�"O���3��73���`M�33S�)YS�'�ў"~�e-=OUn5���9g��=�!#���D'�S�O�<����f��%!ƍΙ!��r���'����łA�fP����>9��)
�'e&�F�:Q��Q�$���h�	�'i��ˁ&Q!Ox�%�F*��kR�,A
�'��<��OU�f!��k�@�1��I��'�H� �&x�V�֗��L>I����> Z���K0�4LC���,�!��S(��95�x���k#N݅K!��\��h�������mÑ��O"i �*NC���YƎY�x�̭�G"O2H�Q�:���[g#ü[���0 "O>���7
�樘4�ώ�0���"O�Aё@N�l�Z��v-�J(-J�"Op��NU� Zn��"�_�<�`��"O�͡à�mˌ-xc�S�L��ɠ�'0!�ĝ�H�*�ŕ�L4j�-� q�'�ў�>�scS)��q´��%�i���,D���סI(,��{7�֙K j	˔,D�L�S"�6uL@��@ur@��-D��%�>x�q��Њ�<���`7��c��@hs��
M#�����	M�R+2#6��]���¢U�<@�0��/8.�A�/D�@�2���V{��?53�	�C�Od�=E��4Ojq��� ����ـ�*#��lX�"O��(�d?ތh�JxizW"O�c�H����Uj
وv���R"O����%	���p4�Ս3�ZH��Y��F{��IF l�<L�g"��:K�ܻW���da!��8�N��j�
6�8�F�](>!�ݺK�JՋD���*<$������]�z���$��B�`���>{��a�ڝ�y⭍ 
)�Qɓ�\��t���yr(� 0�v����B�7�y���l�P�c���Vi��
bF���yr��� �eFU�\AqKH��x� |ɉ5�I�ba�zI�6>���"O����'@�!,���'�l( &"O�A:wn�2I�*��0��$������!LO���Nڍ2M��7�(Nh�y�"O����蝆iP"��8dŢ�"O4��)X8�ZV�X)I
��Q�'�I�w3�1rԠ�P���FǄ�p�B�	\,�}X���<$�}���҈U�y�ɇebb��J�l��@��߅=eh�O��=�y�L݊6�J��1�*�>��G��yB���"̎� Bϊ>"FL�����yr £@%���v�oi< ��y.@P�Ȑc[5e�X5�f���yRLW#\���AP �Y����k��x�'An�H���Ϫ�`��0�؅h!�דc@ +3jB�y���pr(,,�!�GEQ�l*�"�F���42�!�$ƳpC��I󡔃n qd�M0F�!��N�d�:xe+����+�h�G�!�Na�����X�P�ʃ ĀY�!�DL t���#��4X��z� ��$���;O�zU��EL��g�2���Y&"O��c̔�e�ڬ�&L=,B�4�$�<YO>�˟v�b-< ��+4h�J_��C6"O�$���
+1��D�7��Vb��"O�)rŊ��-�8���G�h ��"O`u���g�*-0�HU�xfI�"O� G��$ꤔH�GZ$eP�1"O����n+V��zT�:X&]���	J�0、�zVE��%�"n�⼘5�8D��0g�3L��%�G�d��e��!��������F#(xa"h���'�P-0�f��q�kЧ8Qo���'�X���a�#6Tp�fTB�t	��x��'7&��qB�ѓp2|��Z �yLK�%6�|[�
L<kXZ�@�h��yb�рa8�����0�h�S�yR�>z�.i"i��u�|��C���y�I��AJ:pRr��Q���y掅7�NU��gQj�8<�^.�yRş�^ώ��@AE�f�<��(��y�,n9�����,Q����!���xBI�(���S5�@9i��� �N�'&�!��"N���D;���� NG�!�$_�l|����LZ�+c�=`��@��u�`��7E9B��Bֹ͚��ȓU�\�W�sC���c�m����'nd�[�'�rQ��쒎g�����'�!a�O0�|�c�G/[�9��"�'.�e�r ��t%��,��D�s���'@��&�Asq!�f��
2�	���?��*��.uX���O���"O8:g�܀� ���+��1�h�"O�U�7O��JܮLZW�B���"O�᧧I��qv��8�r� "O��ʁ���T��WiȍQ͎� ��0LO��:��k��!s��>M�j$c'"O��qK�����C�D�<{x���"O�����ػ8�H��އ%pX$r"O<��A�1�
1�l��XQ���"O6�J3/Iej�8��Қ#?��u"O����mΛ�)���� ��"O���R�O�@�6<����
>	�a�"O,xyAk�2��v��)!��}� "O� xɳ׮�͖ш0o	�F8�"O����
O��f��V.��lX�҃"O��BQa��HHb�,{��x;�"O��{Ӆ��wz�[��f[�D�"O(k��"òHC`�=����"O �r��(K���Q4Ꚓ!�N�Ӵ"ORM{�eҌ ��8'�D�X $��"O��:A�^�X�\9�߄aj�80e"O�j���D��a�ӦH�H�ޱR�"O�\!c蛂Aj��y�F�"�	�t"O���C!"����F �)�\"O��/3f�r@��΄��č��"O���hV�k�H�RX�v��� �|b�|r�7o�,�J%�ђL�-��Ȟ�BC�	�<��)�F�V�A��Pj�C�yY���4 \\|p !�@�!�B�1bsR��A�KMD�����n�B䉲���qR��h�L�=1(P���d�������=b6���V��ъ!,0|Otʓ�y�OӦ/F�:q�E�I-�Ȣ��&�y���}P��2R�
�A�4�04����y���(��H�AU�<�>�TE0�yBa6]��}PL�7Uu�O���y�MÖioT�5/;Q��yiJ8�yҀ��]C�i����7���*,O��y�J ����ߜn�q0�jд��3�S�O,�lނ��� ��v���'�b�AT3+È�aգ�����'�)�A��'`��B~�BA�
�'�(�C����)��p`�	�
�'�%!���.G�1`�K�b"��`�'���C�O1w$$�����8Y�*y`�'DB�aV��	�l�gϖ�>��99�'�B�{�ʟ{�D�&��5BCX� O>����iý,��æ[*9���#��.e!򄂯ń#sA�#�%b��!`�'+ў�>�! iD,k7���eM��cQA�@%4D����K�\�f�I�@�s;�C�$D����`�'^2��j@��s���"D��H�C�t�`�
�E��|�0XB��O��=E���E�Z��l��j�V'�u���:�!���.N�(�3��>���"0`��W�!�D�&r�� �J	)����sM��P�!�S3Jgz鐀&x�(�/U�1x!�d��Fؼ�Q�ߡI�*�����/{t!�dN�Cl��BD�$9~t�!�i-m!��*(�,�#f��Ja��C�_3:Y!�Ӄ+
H�A�BԿ!�D� ���WS!�\�+Zp2�l,v�z+�n�2$�!��$(�B�RSLΝs�Q7䁀��'�ў�>�8&/�2+�Liਖ਼3^�$u3��4D��[p&ٞn#ny��-�5T$u�f(D��#� E2�J��t���)�Y�(<D��V�[�ie�l�,R�AE2QJ�=D�TWiEff��zE�]�C�0��<�	d��k�ƟO�6S�ɝ�xK�![��9D�0���ɯh�#M����Ҫd�!��20�pgc��*C��$	�!�!�¤=��8 '
8l�13W��J!��?D�%#�oX	!$�82�Ζ<�!��,����$��Ya썡'S!���/C�,�'��'`I�'�иM#!�D/p�3 ��"3�j��tm��
!�o2��r�j${�6�D��u!�� =������!��@[��B���"LO���՚n2�lD�ҶXs�4� "O@{�@yrܥQ,ɺWkt)�"O�!#���8(BA�U
n��#��'_�d��Zy&�Y�(�P��dB��FS�!�dK�=�BP�'�@;_����*9S�!�D�+lT�"df��$xbń�!�W�	�T	J%J<"4x��,�k&!�$@�3�6H֏�� 2��`,#Vk!�ʃp;H�Pr�`S Z&�ջ5!�dH�H`�2��?4AP k&��3!�D�>���hׂv-.e�l�3!��'x���p���#z�jVAҎg`!�$�;1�R�����X��!p��M�9]ў��S3�2$)���Y�r]{1�$m~�B䉬~T(P��5L��`�FwhB��6?�~���ǾQЈ4#p�"�R�=9�'�d��C��,w�8S`�]�v�`M�ȓR����F�]NX�bVoߋ=y@u��y���B	Ӯ)�lt�F/PS�tX�ȓ�e %'�<tb��2�֊��Ą�,4ƭ��E��N�'iT
?BNԇ�>�����`R���h!m�Nz���?�zĭ�w��L�MU�^H���j Ys"�c0bѡf(ӕ"�؆�IH���́f��@9 G� ȓM�
��T�J��
A�ʛ�T0���s����R+�mD�
o��ȓ|��զ�!�h�G��z�5��3�&,�DJ�B@��� ���iO�	2L�S�,���cX�S�̇ȓrb"�T'a��\b��0#�~t��6<�(Qc�)G�j�I�k�� ��1���Kм	�q)�#;|��|%}�4�$̲a��ND�@���wp�y(�֊s���H
0���ȓ02�x�I��y�g�J_l�ȓK�`��ƀu�0���%$݇ȓGT��*JДI3iP3�`@��t_J�7�
�d�:�ǎ�{�bA�ȓ2��s4M��i�8eK�/���ȓ$�,��nW9 �����#�0���G{"�']JH���(��A��/"�&�)
�'�Ą8Bm#*p$-C��ճq2nb
�'��{狏W!��zD,jQ:r�'�vb,� b��4�V�c	���'lX�ȓ���P��3X䈰�'��p��b��(�q�ٛS�R���'h> "�>$��|��j�EP���'���`TfD�O	�A);	��'$D@���'�� ���7E�,r�'�f�Zh��7�����N�+*Nȝ��'����@��:�Dѓ�HYWδ1��'پh�(B�L���S�FwV���'T���'1Cc�0Y�IԞ)��F{��O ̹H�H�%fK�J�K:�P��'3����2`�d�lR�[�@Ap�'����7!���d*۹W��(�	�'5t���G%E{�a�@Ã:����'XB�;�C��`P���N�2�T���'=X{�BL�::�R3h2uz��
�'"���%"C̀ �����V�P�P
�'6�q0�d�JU��kD�� �v@a	�'��9�I�#}�>Dz�O�F{p8���� ^�1@�Q/w
@��7:9�6\4"O���AH�%;v�R�Y lێ�a6"O~�0i�	J�����f�2T�$�{q"OB�
�*�- �vP�(1�� I�"OT� �JҵZ!P(�B!ۻa��ٰ�"O�5��D�)*������!*�y
T�|��),6"�p��� .�q .�K�B��%Gc(���L� J��u�A+�6oÊC䉍d��������J⣖�vw�C�'�H�a)	�.���Z���h���=��PF]�"!+{H��۷GD��j��ȓiŲ�����K��H;*f䕅ȓ*�~�f��7;�@[e�j�ֱ��:h;�I�M�`[q-�h�}F{��'9V�q�dE7%"�"�)�?.T�H�'DP���̗n��(�5�C$�p9�':�ia̚�g��H�ݠ|+�Ku"O�����N0��B��<E3���'"O�T(e��3�f��*[�&D��"Ot����Hk���K�A��u�'�ў"~j��#jkʼg�S�T��ȡ�(��?9-O����g��j#�9�|,S�I�`����^��͢e�ĸ�F� ��ϕX��ȓeN�� %��, 8���܌��A��Q>��wK	w��U��dB��B��ȓ4�|۰+Zu��ݺP�åY��h�ʓ7�!�Ǫ�\�lQ �a];�@B�ɺU�L �ˑ7�2�a��5;'B���Y����&��`���᦯˚I��� D�2D�@.e���;R �?��)�6��	!�$�:ab�pW�6�]`Ձ�=m�!�]++��
C�Įn�<{&@ěo�!�d9=� D�&CM4)m���άg�!���@=Z���EU�A�F�t�!�$�	�Х(�!K�DOj�#�L�9�!�D�iPx͒�nթ1�	C��v�!��E�i���a�����YG�!�$KtN��V�O9#cfI��%��6�!�Č�o�:��%��78FJ\�é�!l�!���/3�	��_�T⭨�'��I !�B&k��	���2Y:�9gǞ!�D�q��Zw��'%�Z��e)V�!�D�7Q��À��'����EA�V�!�_�" ��)!JQ>S� %��F��/�!�F����U���R�kRN�!�ԛF��a勅�x?�U
��<�!�$	�J�;%���h���(X��ȓW��P�����-�*��cb�.�6��ȓp�IC��*&W\��ON�O��܄ȓ]��1�%�P#�x7bK8/6&X���R��Fġ�ihm�>4
�D{��O�mp3N2.�z�8'c|!�A	�'�HQ�6&8,ap�VCC�CfP���'��(���C� t"�h�;S�T��'Ħ�{�㉄Y|Ja{GC�Pw���'M��A䀨^/*13Ðys�eJ�'j��5�	347��;2J�5����'@"#��؈w��gJ,O,�p�'�]�S��>~���� ��XY���'���ɇl�?t$I��RJJ���'8�Ekf	�B�إCC?4o2���'݆�X�f�1��#5iC!+���
�'����n� |JI��苶�28�
�'M�*�&Ƕ�>ɑ3��0h���	��� �����_�In�����^)ON�R"O��`�N�5u�nE���J�0IZHAd"O��S�,�N<Y��C���04"O��������iӃč,%��9�"O4�ɗ��#6��K�bEY<�6�?D�D{���7 N��s�Re�Q�&�>D��*��5�I�oߝy�r���/D���D�'_�(�v�ް,�P���$,D�H��c� {�@<!��@�^�� ��>D�Th�ϖ0BZp�t��8 ����l)D�̡`i؈d�B�ײNhD��p�'D� K����@�z��H׹z%<9(5F$D�d�'.H�r�)3�U�1�i� D�0rd�1[w������M�f=D��Ge�Pr~��'�ĩGґ"ō/D��0��O/��a��-GB���� D��9#0e��c�nA�	$��/;D����L�:?� iV"8��Ex��8D�8�`N#2&�$[��I{�����4D�`��D�L)��@�C�NS��8f�8D�L�ᔂmz�l	V M�����;D��be$�����.F
d���1��;D��9v�S�+Dy`VK�!%z@�D�7�O`�.��q���P�I�$�@��Y|\)�w!w���J�cg&(�ȓ{6�<	3��`M�8K&`�,B������G��l��y2�	1u��Ȅ�mΰ�ϸv( ���+9�$��ȓb����� �%�x�x$ӤZ�f<�ȓN�� ��ͳ(^�Ю@�r��]��06"�@�.	��x�R�@��h�ȓc�f�!�*ߙi+��%�L#zP)�ȓ}+rX*��/)���H�'�d��ȓt>}����4����o�<rv���,0X���V��q�# <f����P���0n̍O����!޺9�0$�ȓ[?�LZcbT:WE|MsVF^�
5"%��9^��׃M6R7���p�h���a��q���_	D+��C��J=]����ȓb����OҊx�*dk׎=��E�_�,�|�H�9{�z�N(��x�F�N�<a��ͬ� ���ʮ>m(��Xt�<��\�>��!	 #�y�C�[�<��G�SވHkWił�쐺6��X�<I���<�=��cؾ�n3�`�S�<q*�m�~,3B�ٽ4�b�"\g�<Yd.G�G��+w�Y4
�\)H6Ϟax��GxaH;6����щ*/��u��,��y�%.m�<,ĉ��+P$�/@/�yroB"V��Ҧ��*�Z�����#�y�g4)?��Ʌ*�.)����0J��y
YTY�����8!4��g*��y�&��
�� �%7��a�F�D>�y����Up��o��{ޱ�s����>Q�Oj����Ʉ*����_dV���"OV`�%\G銌��/��Ye�B"O6�rwb�;�f8�(�S��d34"O����d�U������3c��iH�"O<lH��Xn�Q�,��-��9y'"O4<Y���9�U��_�b:����X}�<�a�B�������)Ų]�ŇƓR��0#`��Ӽ4@�@\(Q�*��'/�Ek�*e0�Yj��ˋBK����'4�Psd��<vX�G%�)@�~l���� hhSO�$��ЮM/
���"O���듅c�����ʁ�%"Oکע�<J��\*�����1Cv"Op5�6`]���C�� D�~�"O��Q�2�hI�A�e�F	 "O�`���B�d�sK�2|��y��"O��A�ʑr�q�$��	L*��"O�Xj�܀1���V=����"O�cS��%��|���&�x˧"OP,p���
�긪g�Z��~abC"O�y���e򐈠SLZ�3�:Р�"O
a�i�u���y�Ȏ���S"O>�A�_[4��S��=���T"O��;aH�h�|��eZ<��%"O��a�Nϥi� �3Q%�%D�D�)#"OD9Yq�':RAqVK�6��!`"O�e��K_ƄՓT)�*u�H�"O�s��I)�2�!J��^�(j�"O.M�R��/Q��հh�*~O,A{"O���p�@�K@�<��T�`��"O찠����6*��2���	7��)�"O� ���/��,.��E�!"O�8��ҼqN�	�r瀫:Il�1�"O���F
۶7,l�擽s70�"Ox�9�瘝' ak@f2'�)�2"Oڑ�U�%@�&�$5*4ݡ�"O y�SlӘx�N�S���P�"O�!�c�Ø9��"�l�,�|���"O<��6�m����JĨR�j�{#"Ot���[
O3�E�RDܛ-�F(Q�"O��LV+reH<H��Qخ�J�"O.	���
�`r��,VvR��"O� ��o4T�p�!ɺO��m� "OV�aUjHD��eF��$��$��"O8�"-�04��-��L�h��y��"O�k���q,`�U�H}
���"O�Հ�
��=Vj%�q		�
d~U�G"O�HБK�4�T��K�A�X@�3"O�A���˛@��e����/^��RD"O�d�����%�ebw#��Ĭ�b"Od�j%��KTذ����!H���ۄ"O@���"�@pV���S�4��|�R"O�$s�P���j�W����s "O\�:d��rȾx�1E@blLI؁"O|Bŧ��'��c�mQt�"OZM�&h�@<-2W�W�\BhiH#"Ol\�҉ƙ-��Ur��1�U�"O������x��1�c@�9Q(�\��"O��q�G�-x䐑H��<h�"O�5x�X"w��lS4�ֽj(�X�"Oh��o�%EU�I�&A�_�.lq�"Oذs��	ra�ǣ�>1v��6"O
I1�!��Y����a�� ,�4�x>��rM�P���A{�F���&.D�<B�H@M*$�D-��o}�)��.,D����=}���E�r���j�8D�̐�`Z�S�nt`C� �=dB$�QL5D���C�՞c��	0�ę�=4�y�%5D�##4G,X�h� "�mY� 4D��ʒD�R�<"��gb���/3D��pkT9/�D�2��k��9zF1D� �!eȿe�j%I��1Tku���.D�H17L�U^0�2B��0�4�㴧(D�L2#��$2��x���U�4�vB�)� �� h0@����A&�
AT���"O��Pf	ʏk.���  
0+944ɂ"OpK7*�sT�ѱq̐�.(�$��'!�ܐ��ݷPvh����<	f��U	%D�X��<��r`Y�]du���#D�\�lINz5���9��H�j"D�� �!�%�����!.$0���;D�p�E瓬/���:��X�"b���),D���lX�^��'�&#�&�:��5D��"�kɯ0&����#�8b>�Z�9<OD�$?�	n�Ȱ���S7�iC�(L,)�hC��sY��`�ʡk���0��
��B�I'4S�-�dg� T{\Z�̆8	<�B䉨t�<��f��y�1|2�C䉎p涰K���<}�A���A�C�C� t�H�����6At�p���^�C��,5gPhC�ϩ|�p5a�
.8��![E�=� 
/%d�3�Ԍ1k}�?Q
�
�N$��'ҍ[��)��A\��u��SO�`r7�	��fR�)P�0|���!�l�i�)���	��c�bą�C��膊�b(^hI4��]�ȓ(<�x�*A%�*`�HIi��y��-�QibE 
Ʃ	�
���Q�BѢ��4lZa
�#A���܅���L�T�,m����.�r��ȓk����S�385S�-:X/N��� -"�%��1e^i��%�f�* �ȓ<*( ��׎/W��(�Ɣ�2Pи�ȓ*�&0�	�s�x���G��t�8��2d.-�SW{�j�c턚WWj���f=`�@%T�[�>���VC'���Et��KB�za�H�h�4����ȓDqju�dNa�-4��\S&�ȓN�4q��
�w~�P�0퉓�l ��4�����'B�sd����ʊЄȓQ�h��B*���i�K�+T�Նȓq����U�Y�x)WNI�0.���ȓiB�X0����U��c�|�j|�ȓU�T�yp(Ҵ��l�"ɔzv��� ��신��1<�>��r�?�Z��ȓ.�,��dn�.��,y@�[.|͆ȓ�=��n��!�c��	�ȓJ�a�WY�rɁA,�S�6Y�ȓ$w������n����I�i�l�ȓ9Z�a��Iօ)\��BbfN�4����E�@��d�N.T:�}�E��$�^��ȓsv��I1��1Y��������ȓ,��m(s��.:��>��P��n��8��^,�4�rLޤb�ZB��t��9� V��x�Ɇ�n�B�2a¾YӔ��CY��ѢG$b�B�I�t� �C��W�ș�&H8=�HC�ɹ ФM�3�C+=���@�J�6��C�	�f��0v�ҏg�E�a���C�	=n �XR�똞]G�R�*N;�C�I'U�V!��CAY�D�
��L�hz�C�	 GS�LҰ�S�@���(p��0P6zC�I6F�fPB��2B��A1\$h�bC䉗�\�(�3}���E�)[�2C�ɾ�M����\��fH�)��Մ�g�x�@�[8w��E���
>f|�M��L���Q�&�)��1�-�>9'6݅ȓ/+�`�+����Hr��?� ���S�? 6m��Ç�^�H�R 	�k�Ҁ�d"O����<]q���qǈ�>�^��"O*	AԀ�4D�,Sл�����"O�]&��4����&d	�����"O�B��)H6��#��Цv�CC"O\��f���a�	����6"O�	P ע4z�𮊝)�}I"O`L;V�9{L�!�L�A0�"O�Hs Z10�� KULɏ7�ira"O�M��Ĭz���@ߴG"�p�"O"�铈ݟ��E�E[�k�@@�F"O6%bE*5R��ip
_��v�k"O�=����mw|(�(��^\���"O2��s�/t@B��?BE�1`�"O��hq�Bxu�#����~ pR"OiK�����:�e�L�F�S2"O8E�W�o(H%['�J�4oJ<��"Oz�A hG'��<#�%c��a�"O�4ˇ���*n�
�SJ�}:6"Ox5y��K9���QC�6P�	0�"O��*4$ZN"\�$ �b�	0�"OԈ���"�0��e\-Q0D�G"OD��O��T���"c]2W䶴�%"OԃK�$�\��!�>@��i/�y� ��LSB$84�����6�y"l�1�V�1�ɰ)���w�E��y�3iB<k��Ŭ)D�!ҵ((�yrς,\��y���� ��a5K���y��Ӎ9N�A FˈK<$��$	���yR��8V9��G�=�r����N��y���#QB��D�_�4�:P�-�yr  /�(��F L�3G~Xhb���y���fO�CR�^71�ʌ�$�$�y���
��Iq0��.�@ ��޵�yr �Nwl��G�)m��L�y�Z��T�7�O�(��C���yh�ȞT�غl~��A�ퟣ�y��ӱ=��@��=N8�t(UIH$�y�LG
�Zq��z��J����y2n�	o�Ŋ�����i����%�yB�ޒ98,y�kǰOݤ)"�%Ƥ�yr��v-�n߇`4\3Rm�*�y��	y�!r��^�!�ݢQ߸�yr]2}���T�Ķn4��@Q`�;�y�	O�"�����c}A�6�y��ߨsq��#�Y? d�1�M�y�)V�Dg��*�X� ���p�i�=�y���w_:8Q����u�B`�C���y2�q;����s-Xm�c���y�͖	���Jg喞:������Y�y�`�2J�.�*ƊV�,�\lI�&�y� CTTL��D��W%X:��Ά�y�披a����3�+K����գڪ�y�G-Q�x�ө�.?�\��W�y�H�	,&!єa 40�\���'��y�M�/{�0���A"8��˱���y��$w�ܸ�lP�P�N��O	��yA[誰�E�*E�P�!<�"C��-i�ȸ3�V i,Qo�"+��B�ɸ;�dp�͜��qsTF�+��B�I�g���A���0�����G�!�B�k�8	3�.Q�p���R��b�B�ɷ4����d/�EeN���&bB�	>Y�@3���B�>�'j��(B�)� rԩ����QsP���p�""O�!Y� K�c{`�U$�
�t��p"OJ$�R���Xt B ƽ�
e*f"O$Ejg�A��@9H��L(d)�4��"Oj�s�� '�F���ǁS��=@�"O,,�兊/�jI�@TTux�0"O��!th�a  0Q@�]Y]�"O"D:b$�lŦX �oR&WRD@"O0�P���z��0I�+NjH���"O.�a@h!�ܕ B�	e0`���"O�X�솤>J��W�ܠf:����"O����IW���8!p�Ϟ!-�9��"O�i�O�&
B� �'Y"����d"O.rc��!WÞ-���<1��j"OxDS��N���	GD���Z�q"O����j޿Q�$����=N�PY
�"Ot$2.Z�4��Az��;O�`AF"O`HqEoM�U�H亠�)!8T1�"O.�iJ�?�0�)sE�9 <�;�"O�`(ժˏ�T� &<� �S�"O�h�Q��	N�-U���;$�7�yrjڝ�6��Ȍl�8��l���y��a�ŋ�+��b킅��E��y��iM��*���G�DPQP��y�&ɘZ��z�L�*���ρ�y����^}[�慮W�"�H��yb�A7�*�:$k7S`$$`���#�yr!M�*:i&E�@����	-�y��P�_"�U�7��@����#��y��	N<�����5M���ŉ��y�V+Ჴb d�;/��H�BRG�<���J�G\:�cs L�t��P��^�<�B ��2�T�@+�ţ�'_2;�C�ɩ�ځz�m�
 Dy���۞.VlC�ɜyv2aH�i_4iG<mJ"��9Y�C�I�,��|q��%��R�"�8�/D��!r ӏZ�t����e2�k+D��H�E����̼*z�X$O&D��"����4���L�3G�*'%D�� �ҕN���Q�cݳ�r���>D�� D�FP!p��B1``i�>D�dI�e��.
J����%P����)D�d�T� �RJ��ア�2�����+D�,+B�@�%���T�W9^�<<��)D�`��˫x�(��dԗ��5q�()D�8X��L�_� ��EqA�dв(D�l��6M���Q�m������$D�4bB&��G���	�8��8�,$D�8H6aE�*,S�ș=�@�S�!D��b��B�kl���m��W���"G?D���5�ʞ-��MX%L� \:P���=D��S#bE�6
�� �%�� ��C�7D�4	EK�,ip�H9��Vi�pd�)D����'@:	q#��T�-q��Sw�(D���uF�-R-x�W�&��ts�'D��K�Ɏ�.tHզ�3�TI�m2T�Pq�AT�)�$��(G;C#���e"O��[���<N��ggH���̀"Oj�:����{��ग़�p�҂"O� ����T>��rař���{�"O���c�3UXn�w[*[)dEr�"OR<�C!O�3v-(4�Y7y|�)�"O0t9��M�K�NG:Q{�i"O�]Z��S�l�*�.�>�4�b"O� .����*��@ N�=K>��7"Ov�0r������^�1��"O�u[�J�G'���R�Ȧgs� �"O��3�Oѷ�~! f
T`�Es"O���s�(5���ֺ$��xr�"Ozx�բ@�HT9KU�F�D�"O����2!����/���X1"O"BC��r:}�P�Cd�|R"O���߃b��ɉ^�4�v�rs"O\�R(�"-���`նq��Q��"Ole�%��� �K��'&J�{7"Ojh�Pl�;-��%S -¯�`��"O(�@��<=��2�+�-E
u��"OX��i��"�C�̓#��H�"O`4�1���L�ʗ�[4X4@�3"O&}bj�5a p�#B�qɌ�� #!D�ȱ�Gz���I7t�4��D2D�\�G�<v,=8s�E9�
�Z1�1D�!��]�>s��Hv�e��$D� E�߷0�djLY�kڌ��e$D�@(Bh��X8�#�*����ad#D�,�a��*J]`�Hւ,Y���7�?D��S�On���c�Α]7腡�� D�lh��F���كN�=c���`"�#D���T�;W�\Q+�@fۤT���'D��@@+�'�^Y����#Dy�u;�9D�<�UCV�s�9`ү��N+�8@Ӡ,D�$ccG�'��`�SI�vК3,D��JK�#�(i�*K�~nV��@(D�hapϝ�D��µ	�+fN`��F�%D�x�`�^&v�Жj���Zk��"D�pR�h�
=|0���Y��a��=D��(�`}_�=H�'@(2 h��;D��۠?j��2b���%D�H�6ǂ	d�6��oB�Z#0U�W�%D�I5$�=>��<I3�_	ac��18D��h���)G�}���&k �5D�A�e �J��e�o��Q�� D��5�E*\��U+T�'. �)�=D���v�W�J��C`b��a�h=D��h�/
�t����)�Z���R֭<D�$��]�k�H��׍ߤ?���AE+9D�dI]rF�4��Y<d���O��!�D��Q|<���#W�bXi)VhͯH�!���&��9Y�!�Ա0˸o�!��ƄG��<����;:�E�I�T8!�k4� z���1B5��d&�o�!�!;'0�j@��5'�`Q�E�:B�!�dϯ#S���'�$>{�ݐb%2!z!��
��1H�FF�B`�,[&#� �!�ƨM����M��b�ys�S`!���i�:����#��j���!=I!�$Z-��d �w�\�����%�!�$�>S�%�C^��Ġ�!MP�K~!���S>�(��R���+"���#!�ă9!����� I�eeDY�7�!�d�j�K�g��(;���b�,�!��T�-�����_+��A	��!�$ݍ{�t��"厫aJ�Dł�9�!���&%�����_�|]l5��Lx�!�1A������S tH���N.�!�+|�hIH_�Op�hYv�n�!��ɲc��ݰ�Nވ.I�,�r!R�q!�$�n��Q�i\%�28�p#�=!�� hի4��7�x8Ã*=x"OT��e�>hتi�$Yx*�C�"O\��s�p�(���:�H(�"O��R�
�[��S��V�"O�PR�O��Lz�dh�	594$��"Or�c���,<H�E:w�۪$`a�"ONx��f��6lP`���()�|ف"O���(�;0�m1��	'<:��)"_�����<�2B-9���s����e���V�OX��O�����2:����eo_�T��2�"O��ી�I���s�X��tڦ�,\Ob|�t�T�)(�)���R"JDQ!�'ɱO�8rA�9H�����	Ϻ@�M"O�٢���o���x�h��*�<�b"O\}ؒ��l�Q��}���A"OP\��H�9.ѳ��H�C�| ��Ii�O��ed��[L\�M�@�x�	�'�8��wC��,�dE3DX�2'�Th
�'44׀A�>�(�n�A��0
�'��4��J��n�J�O�?�6�Y	�'�Z��AfZk��Xz�GL�Y����#OMA�n��ՙ���=�2�)�Z�X��I�80E��-��j�B��R����.lO��'��5"V���X��I]�V*4�
듍�����,T�A��+�L�"���|��1}J|�OT$ap �8��Ȑ�kD.X|�0Y��Iw���ɓ�~w�� ��^�x�f�h����M�����,�����!J�]مF	� ~�  �¥W����G{�x�l���[+R����s���-�X��=D���c��.�H����C���m���6F隍"G}��5�Aլ���)��:��-zE�-�p>�ܴ��dǪ\�L4���D
νȴ+�m��D�O���$� ?�ҝ������J�iX�qa|��|b��8���kP
­l��Z�o[(�y⫚�Z�=*�M	�8�r aZ-�y2�5K���xC�D��q1�
�y2�>/��	��Ɩ����ّ�yr��n��|��C&N*ƵZ"����?�" �OdU�C� �ɀ#⍍s7�9�"O.̚��N$.�b� ߪ'8A�&Z�|D{��i��!���V���CEC^4A�!�V8o��h��4��aR�a��:��d���=���ٟ- XI����c(6D�� N9T�!�d�.�%9d��!V�T�� �!���P���NآB\��E�j�axґ�$'���_�^�ha�i�<kk����j(D����'��� @��ϛ�6�����)D�l j�. P��#�m��(�R��(D���C8u�<@��eD< ����� 4���� a}*�hLW�6m  ����~�<����h#�q���[�eGt���C�S��i�0��h{*l{��{���8 �6�6"O�WN˔w��!CH�
�D�в��G���O���8�

'߮��CAؗ?�M�	�'��H� ��P� ��Fʚ+�Z	�'t}� ݼWw���ա�N���	�'j�8��U�K���˧�0`�@�'�T2� �E� ���n)C����L�R}�_��S�'~d4��\.Hq!V��!J�h�rs� "Ar�C�^C@���R�w2F���L�-���C؟̣�
X��6�e��<^��D�=LOV��$I'w�)�2�?T� <Q2�<Q�	p�'2�P�H�<.�l��c�.. l[�'�J%���j��Ӗ�O������� Xr��.C��{�bE�	��e�b�|�~zǥ~�����߭iY��'�ě /��;D�@���GEJ��&��n$#�8�	X?	���O��P1$���y��1*Z�����'�X����$�,�%��O/NY��'{$�Dy���S�w*��p�;Y��t�\��yRb�1��H�a�N��y�Sj���y2�\ 0�q5��d{�����	�8�1O�t��'i,-@��vt$�C �<?����\�$�8.\��aK@�3c���S�; x��^��$}J|�'N�dp0ۖ!���a��<rZI���HOډKtM}0�!�@X�Z� R!X�(���)�' ��9z�ƛW�Ti�	�i���z�r,:d�ЇW�0pjS7y�
����M#𧒟*�<#���,W��+4�TC�'�Q�$j��'v0�!��ҖmS����ʳ>34����D�O�#}2񏗙0�=�ē��H�1/����D#��?#<9E�Ѱe6��kL(|����Bk���'��Q� G �
�:e`D�`(Ru�dO��xr�6)뀵3$�M�t\�կ�%�0=�شj��'�P�N1`RHXE�ٰ �.W<D�4aѩQ$Bht�U��.?X��� 2LO(�(C���~�8�8Q&}��_�<Q��	!+v}{K�Is�M("�X̓�hO1�d��!���>y�3�\�⩺�"O<�A�i�f�Ң�l�0U� "O1B�m��;e$TZ �5_��T�"Ol����	�����_'q�q�"Ohx�À_�)Sɠ U�Bn"\)C"O4�;�]��0����>?���3 "O6�� &ʹ���3Ɲ�5NĈ"Olɒ5 �
���B�%�r4��JP"O��26�3\�b�.C�B$,���"O��pDO��	��Ś4��;n��Ɂ"OD�	AfO�h
�`�
���I�"O4�xA�ʔk�͚`ϗS�\��"O���J>Q������R*F��IS"O
��E�A�ay��Q�ϣd'�|d"O�ur�B���(�
5�@�1"Oܝ��n�ex�@+�bP5c<TA��"O^���ܼf�¤��A�" &�"O�\g�'D=ZQ��O�V�dH �[����ɸG�1R���< Y���g��}|>C䉳	d���
"w�
��7��C�	�<�r1 �O�_��y1�e�B�#<я��?�I��¹G��	�+�&_֕x0%3D�p���d��іǖ�B��L�X��I5�hO�>�ï�e}�U�bJ�i��()�@;�O��y�m}�]���5"GRX�cIP�y��* o���$j�m�Si ���<!���� (�r��L���sd!���^��d�e�۵V v}ӵe�ab!�D�9w^�4 �+7|!�FK��#1!򄀝#� �.��N����J
+��Ic��x�c(�)(<Txa	G.s�	P
3D�䩡�J�R4�ّ%_'K�b��@�1D�@�l��.H�C: �P`�C�9D��05ir
��� ��[���#D�k���xP*�� �M�eR�h��"D��a>{ڌ
�C
`�D�BD`!D��X�ɝ�u��$-�=�8��3D��*�*2���a�K�e��ٱi1D�03�)\02���o�%� 4S �.D�`Q�d�,���Kp��������!D�� f9���]�x�>x�"^!"MZ�Y""O�u@¯@�U	�j�lW?$��b�"OȍD��]�v����X7p�k�"O ����e���z8���"OԴu4w�z�A$A�Dl�0"v"O�������| 3F;@2=�#"O���i��_��a+q�5C�*t!��I����N4�yq��X4��Q��2y!���{�R���2^0c����!�7m�޼3f�	�:i�I�c!�$�!HW�D hH \��́g�̅L�!�DC�?/�����'.x��h�>�!�_�^��Ib�+���b��҃zz!��ՁAv�TAƆ;v��ӵ�6>�!�	��a7m"j~e��[�fT!�޲N�|QZuPF4`� ���K�!�Z��A�S  
T<H\���	u�!�Ų%�F���K�O<�e�`��8�!���L�� e�!-7Tq(v,�g�!򤍥lj�CK���08���z�!��]".צ��KZt����JY�!�Oj-�L2��3	/(�����A!�� r!,��w߾V�J'�< !�ē7�H�!T"}�"(ZE	%�!�dq+R��LS�LƐ$��Es!�ė�2Ӧ��C�����0mF�?e!�$�)�zx2�&�PQ��A�>{]!�$ߗ�T�r��\t�=c6ʑ�P*!��T9��� ߉~~�hr��2�!�d�S���(��gb�a��	^k!򄂆#��H ��V��88�E(@h!�d�.�X�� ���{¦M�eL!�D�/]�
q����9@�� G�L�n�!��^��\A�K��W�N1C�;�!��Ƃv���Ad��B�]Hu�Ѝx!��MY��6��+T9��ܐs^!���}>J�i�'n��u1��45@!�DS�|�R<1�ʆ�z��m�Q(!��4�r�ɵ�'j�4����.A!�_�8���YTD)J���a�;E'!��%�������i[�23���?�1O�J�kZ+8�V�"��XF&��F�'K����27�H;�̆�F!�$N�P�dD�d�D
��h)�D�!�d1+� Dk0*�|B�had�)�!�Dז��ʷ�X�0=�5SQ���|!�DʡTH�-�L[�n�lYы^�N`!�$1\�,l�`K;G� 1#��j�!�D^.(o�����V�#��}�&C� N!����~���6G�8��d����!���=�lJ&J��?u�h�d�K�;�!�$T�!D.]{�K�x(�9RM��!�Ï��Q��e�;gǲ��c� �!��+ai捻��ȞT�&]�ç�	
�!��(��m��G�6B� `�݅4�!���;,�F8��+����d�Y�!� �"x�u)��D�4�#��Ĺ�!�y�JI��&N+}���D�߇�!�ųjz (�,�u�٢��c!�N�\hD�B��.b�l�5�W� k!�dP	s;b��҉D�u���m߁SG!�$ټ7���Au��>���+� '!�D�0sdhz�D�B�rIy��Y#�!��ޑ4����V�Ð1��;�o�)|M!�ĕ1%k[�2T�l��V�ݠl�!�� �se��0�B� pJ�^����"OVH��)�"�X�c��_ �8}��"O�����b�f �g�0�"O�Y�'��0�s��1A��9��"O:,pEk�>b��X�4�U�.��"O���-��C��s�a�`��9�"O<m��h6.?����W�H* �%"OP����6R�$[bݦ
nʥ�r"Oh\��$��2 �nH�%G�� "O��Q1�K,h����clO�=D���"OZ� �` fI^��ЎR1orH,2r"O�@���'x�=���J�~z��ô"O�x��8>&�Y�j�Lo��"OV�X�`
����9�}!"OJ�1f�S�z�N|��
��K@iX�"O��@��Ѷ�׉S/KIX�yV"O�%��kHg�2h�h�XPҶ"O�p�䅧-�qI��H�Y�<5cu"OF��Q+O$z��`��{��P'"O�Pp�OC1���q+�,@�"O�U��BQ�JY�-XU�Ȋy��"Oj�"¼Ee ���I8\�H1 "OH�	V*
n�P����?gDT`�A"O@	�傅
�lIhp;QH�
""O����.�;�r�c���D(��"O$��	J�y��!�'e�	y$�EQ"O�	�*E�v���z����9��U"OJ�w�\�Va,�P�#�^f�5�"OxP����m���� /n��d"O���Ւ.	�C�`�0_�I�"O&��u�SS�����@�D�1�%"OJM�aR�p�\m��uaR%I5�%D�@��NԮI8�,I�N� �%D��� N<)9��9�VpI�d�<)� ʔ2@��S	ӓS��x���u�,;��N�a��e��ɝU�)�$jR�~�y��p�b]�U,ĤK3|a�Ovŉ[�#��x.�&C4
��,/Q�,٢��+g��b(�g�FjT���	d-�$B'p�U�ȓC5���$���G���;5O��!�\8t�	,K��*$�J�Q��)���F�_&8"~dr�/ܧA�,�a=D��;`
��4�1/)� ���⤟�`e�@��`y)t��]X�(�#X
�ā��+�`3�9�O�+� +a��;
5Ӱ�2R���3�.h��Џ^�tC�	aB��ᔬ�?6��dZ`"�T�.�<Y�	�gN���4L�>��O�j����шw��{���u�ԍ�'�"!ခ��o����d>d]1i,�QX}^��S��?�"�<���nΞV�*q��.�A�<A���3׮���F���EȡN}?�V�6}ش�%��<�®�"Bl�K���>]��C"OVX�@�'.R�H4�K$.��6G�*;�DͺG
�_�B�	�u���#kU���ԗ ��=Ib�ĝ��pȌ�iҗc�B�p�kf��A�#���B'!�dû'�l��f��J�Ti��i�r�Q��k��	l�>�X�M�)���h�d�y��h*�<�V⑒p����$V t��@�d]�K���13��Fq��I�Q�d�-���t&�$#����n�^���y$�D(`颅дb�CC�I�H�6xrŭ�UΥ��M��B^���.C'W�^Q@U�[�:��q�;�>lZ�m�D�I�?qbխB���M� R�"ljP�#��+�ax/��`qC�i ���ï�l�aE$�t��eJ����X&N��4B�TB��8�j�榵�'q���v��qj��֓4�$���$�U2��M �	�f\�h'	��7�@��d�-O ��E	t���P#�ȅ[N�n��m떝�$͜�(�	�@˥O���ܧj�Š����0=�"��;��R!�H�
ߠ8���V4-��I��M�~������.�hu��ʘ�	9�i]�m]Ma5k�R�$���ȏd���IN;,�THo$�OB��B!	=h��(�"?ڼ�����#dҌ��V�� &D�!�M
�OR-Bvm�<h��8��\���D�2i��q{�� �Q��-d�E�F�C�bMd:�ɟ��=��)ڐ/�=��*{^h�)�I��\ڲi���K�`CkܼQ�(�u-;Tl=��Z���$		�nӬ��"�)�	c,��"4mD�2�	󄪋�g��˓����L�(-o��;�d��>�U3�M��i�2��bfX�pI�ם�36�b*
�)v䄈����-�牬$������	*�x���9;�����)�n�@+�e���o��B��e���,�p]Ҡ�v~��)�O�b�8��g����ӬW�Z+���P��9u���`�`�U�x��DU.W�N@�ƇI�J&��7J�rĘX�����mp�̂❱{� q0g�	�9�ם������ś�%*&�C�.�B}�%��C�9��+��D�;���6`���'(�&1�%M5Y8xI��->�>�����'P�h�u�{��i>��ڭ����N<QQ�U�ʥu$��!�T9�b�ry���������H�T?�B�`ވh���5/#����%Տ>��r�a؞���>TJ͈���/���I�pɢ�)����>���#@�&d�$�O���'���H��Q&?��g@���c��^�aV`���"G0P�5�u��F�T`��X��<�U��m.�$��5]���'4bV���
�As�'	���[w]<��/�/��O�Z��@JO�>Q��	͸F��-(A�$A�p��c?����I^V��1aӢ�,J�\9��I+,��0�i����O�qr�"8uNduQ��N����W�0��ME2S.�#��>E��J<6J�*�&�/V��g/̾��D�54Y@��N=z`ayR��#�^#��ܦ|B��*۱Tp:�'�(�T�f���~B�Z�Up4��+��x(���<
߶#p��$N����I>Q��0DUGD�Ii���I�h��O@iYd�ĉ(,������<d�>āH̥E&�Jr~Jџ`�p�"4�%�@���Ї 鲉�"]_�X�2�	�y��Pê��v�5��
��<��$[�aB�h�?��)�'

�1[ %�8<Z$j�X�Ct�!��xT�Y1r�Y�����'�[ rċO>	�^Y%z��|�<y֌��Iܲ	��Y���u�v��{(<a�U�Q��i*��T�
Sry�L�,lF%�?���e�'-hF�9���,8�P�b!D�<Q��:P4|��K��R�$��!D�H���+άdO#f�v�1��-D��s��QB��h��]�ipH�5f(D� �u/�)N� I�B'e!Ftеd'D�̳�b��$�"1Q	[�X�*����0D����͑R�T��UiR�X�RL���/D��Bg�Q�
S�\*�e���:̚'�+D��{O��s�dda���39uؔц*<D�d(砏�i�Դco��;h�zV:D��Y�"L�|��L!FAX }i6��t"D�$A$@�6�D��$�8���dI%D���� �:�����Sߌ ���$D�옔�\�%o�0[�K�|��@�@A!D��ңaP�f� ��UH5[�xs>D�P����*pjx��/�l�+7?D��ҲlĽ&�H5��}�\ɸT�.D����n�,��4��EĦL����#,D��(�,^1`�h�AMI���"9D����b!���"@I��ِ�4D�4�U�&~���S��-����&D�(k��
8s-Xe�Ic�q�5�&D�h�Å7`��`E@75�Fu*1#vӺ�I�&8��>�b��J*���낹9jj$���B���U��46�A��O�|9t�P�A|�L�3LM�o] �)s"O�e��E�(�TB��f9����x�(�#�z)%��6MZ�D�Dgjam�O&��zI�$�q��'?�s��#V� Q�௛�/��@٥��e͔=z�*�O�!���H߸��C|�"^$(U.ػ��Ć>N�VΊzy��P� <�r!���c㠤���K�7��	�DJ�Vg)�Q��, 9㶼P��4O 0S�-�f��Y7G�!��"SN�Y7 G�9���S靲k�!�D�/8���Y�#/���ό-����GZ(�k^<t)�e�5=�Q>{��*^�x�K"�T�q���k 8D����0��pP�L�?�ukW�<U5��K��H�D��̢�#��r�ʓ��b�����N�~X^@�an�o)|���=�O����.� ��
� ��Vظ�f�A���vJ̯
�z�*ď?l�h��'H�T�c� b���Ň6[H����dNz�2T�U�E%�@q��^� ��\�U�~�f����	�A�r��(D����\
O0��s� ��S������<YO]+zZ�Z�N�-��	�Bӌ���{�n��~}D��ë�(�ɉ�"O*����T����0��˛`�j�ax�Z=)�ʛ�H��!&��s��OI1O��*/K�y�X��m�;h���;A�'e��s�X'Zi�A�`�e�hT�4K�8\o�Q�%��b��,F�N�az�a�0?�j�;3K�2I�D�����O�гE/-a4\��E��>�d  �O _����I&{F<�0�P�F4�B�I�[���nV�"X�#	L� _~�iF�7&S�Y��8�U z�ģ|B���/Wh}����Kx9;@C	C�<it�i��PJg���1V:0�Bl��C;���vl
$ut*�C��-�8��|�<��&Z)�T�q&�6~<1k��E(<a#-T�/&�:�[�=��A9���ur�r��¨@�u�S����=�F�q��]
G�K,(����K|8� �GI<,8��0��-�D�mZ�'߆9�$"^*vV4�8�ϑ=��B�	�c{�T0�i�pUv����j��O���U!=���F,��h�@�Y�����ĚS�2@O�hJ�"O24*�b��R���WhK�q"�(��G�##/�"M��AF�/�g~��P-bѐ��X�F��}�Pꚭ�y�)�8A>�����">
�{3�S��M+ �'0����K:w�̴��.A�	����dV4z�!�D����m�.��"�cB��!򤒋z�m+�j��D�����NJ!�D/j�PIr�ةc������p6!�4(np�q�B20U�5�w�D!��2�8�a�͎eM��!��z�!�D�8;r����(��a`B��!���-	������3�����B?b!�d˓I�`pJ�M�'�4ȒLܹ`f!�D�>=�͡���ktp������cu!�"��p����g �Pf �]�!�d��c��E����*�"��p�i�!�$�`y^��$
�s��#t�HZ�!��ȫg��ce_ݖpU�Ʈm!��hѲB#�,R�0x�3+�!�Ğ%���fHժT� ��BA�m�!��
?+h� 㪔�R6�6!H�!�$ϼA��w璅�lE0�a_�!�$Q�ir����R
H���#၅��!���|瞤( �DX7��G�+�!�¤>� ЗEW7_5.!
V�ۗT�!�$�2z��;��E���
HH�c�!�D!n&5R�'�i�g��!���r��
��G�n��y�À�!���c::���^�'�t�@��	|�!�d�/S�f����l�"�����(�!�Dz��XJ�d�8j��U��e��a�!��"'-�A��K���0V�U�*_!��)�����ŉ
.�$�3���!��K�dSB4�ӏ�w�&���b֧9!���V\�P+�)ŋRt�V��_%!�*x��5S�g�~K*%Rנh!�D��^>���:�$�� �$�!�ʔ��r��	:�B���� �!��I�e� ԑ��G�Xu�k�+�!�D���z}Zӫ��H�XA!��ҞnJ!�DO�'�5�DF�O���`@(0u\!�"[�2`�7^���a凁5&!��A�I}@�Z��*[�`<s`Ǉt&!�D�� ��p�/��]��ijd��4<�!�US�,�1�����遵�N�Mr!�� 3���&�q$�(�nCT
!�� ��1��Ύw�b��QFD5s�B���"O>Q���o�yqW�Ŀ�>l"O((�����˗OŜB��A��"OFe˒��*v�<�8,�.���g"Ot[�6Tj��e&Q�xɊP�0"O`|B���><��V5-D`��"O�p��A�2AA2����A6a��ۢ"O�� �`� O@�
D��;:�b��"Ot��,@�3kP���jZ��B"O��`��F��L  ��)~�;4"O�EꂉJ�M��&LA�!��#�"O�L�%�_wנ%����F��<"�"O��+�X!M���K��P�d���"ON]�e��4u2�q�G�ٰd��xY�"O&��׊L*C>�mA�(w��1R�"O���(݄}0�Ͳ�%M�/�v��"O0�{��T
T�$hU�.$�V�a�"O"�j�+I�8r�8Y����J�z�1�"O���e� 15����
�r"O���+\�\�(��Q2I��yz"O�8K�D�2f� q��J�D��"O���o�<���(��سB��""O��������΋�S�=K4"O^��7�}�]�E-Պ$*\�	q"O�!�3N��"4��C�J�!b�$b"O,X��#Iy��È�$mW�%CC"Od�B��Z��麴$A%J$ �c�"O��̔�M���Q�Mח/L0�P#"ODؙq&�D��D3��HM��!"Oġ��i��QG �ӅT9 *Y:2"OK������7k�X�`'��yB��8�r����D��`� ���yB��+�����ٔ
j���g��-�yRo��26~��FH�	�� b����yb�-V*8؉2+\������/�y�*��W������֭L聑 ��	�y���Evi� ��*
B�@ ���y�jɨ&�*h�C����+PGY1���H`T�� LOZI�l�\|	�c�P�9�|�;��'rT�h'J*#��� �f�f��T�h�:=v�+�`�Mh<9 �=�T�$���*�"_]�'.��	Pc׊:�@�4�	X�j��R�<>�j�z� ̕$~!�DA��HݲŢ���t�Wa��f���A�U/^&�u��+�wy���'�����¡[�F1�EHQ"�-r�'��c�ɇY�a��ǅ|�V�'<N�:@�	(82:�+��'�V�I�gdQ̤Z%C	vxHM[�$E��A����a\��(�//D��t�Y153�Q9�`��x"�[6C�,��4v��l���aZQ�$8��j��iz�Z�9 :�F!O$`����gI^979��ȓn�|���o\<+�$XT�O�3�<�L�l���s�˃GW�)����L��i]�pCD�����:D�\#G�)�n�S�Q6o�-(a���HQ$�\e��e�5(IX��a��J�R�J��H,{�괠UD �On�I�2��0{���98�\qp�����i���<��x�"�nf��s��ۮ�!A�˒��hO4��R�g�^"|��*ۃM欤	p��*ֶ���kb�<�G�	3։)��P ��\D�'e�#�X�O�"y�AQ�%TH��2������(O�X1�KK�=�nǼ2B�Xդ&Nn�8�HT�<!��WHBi�L>%>� 1��)���'/��d�������a�^� �C�	(�E�h��1��YccFE�~ވs4`��l�r��45aZh�G��8F
Q�f��N���?M�hZ��L���
:f\�2���  axrj��]Pr�!�i&A� ۤ�~�i�jp0�" ��#R��i��d���������'`���hu:� �Dʹv���r� ;8\|S�f��zy剁A��H��՛ ����\�1J� `�N�X�!@o(��� ��)�*W�-�墧��OPv���O�xa�>��i�
ӓ\� �ˆ1�f����#���᥉�x(+-_����\�V��1۟N������~�؂D�F��8A��2pzP� �h���֒E��!���w���c�V(� ���a��w�l� �nκ=�v�����*i\�!��V�u��˫OTAې��R��=	)��e� Y�v��@&�L����$>M��z�����HSMӼfE�]b���"G� �s����F6PI�-]85�

 �tҴ=ADS��QV�"U
��)�	�=�	@)۔M�l� U� �8&˓mV8)�����X��υk
H�E0&N=I���F]���lB:�[�F����j�N�6�^��>7�t�[)t�&���(������WI(�0+��у9�؄n�>V��c	e�0瓘T \U��O*�<S�@��;�ޘb�J�e�$���J1�"2o��4d���Č3�tU0c!@/��	�C�^�(�y�GȆ7L�RL02 ��U�y������A��L���M?)�~�C�����Q@���5����!����'tM:��Y���M�@
R�0<]P�D�"UA��S0Nݕ��i>�r��t�d M<��LX*����xȜ��&FyB#�9g��p�F[�T?)0S.F�1��!4�:4q�@C�d�X�F�B�����D,)�	�j�"L��	�I��1�Ѵ^6$��#����!�L�@ЇA�4j	$�'?A�ǁ����dn�'lJ���cE���q�A5y��\[R�\��eg�!���P�ҐuR[�, E(Q*b�	40�'A�D�\w�P�������O+�]����d 	�鑍Q�Z)R��ңzL�q 䈧�ħg�f��f��>��Hc�&@�E{v/V�o����c�52��)��L�WbҢX���#�XH�0B�ʵ<��6ea8��H9}��)�*o � '�R׋��S�`�ѫOʁ��C�1��B�'��ȪP� �dSv��M����I.}�L�2�x�kg���'�ܥ����az�;1���Ӟ�"u��0�����'���з��.�QY�%�$~3r��baԻI�@M����U�	T4���L+�'i���`!�B��&�E��F҇�LF~ �X�S ZS����?5�P\q5�ժ�^C�I��x��R� ����D x�˓Kc���!�ӧ(�p%P�ɑ/e�v�T��-@H�p"O0��rJڃp4��2�&�$�f&#���&
�.�0F��dA��`D!Tk��p���
x��q��;U����Sg�oԄU@�,��x2%�	h���jS�H$[K�%�b���y���/"��eːQ+�
3%Ɍ�y2 �/t�̻�AQJ��8@4M
)�y� 3�,�l��Fa�0XNX	�'�<!k�C��!�5�I  ��]��'2��ǀK�V��{&��7$���	�'(8y��E3 ��a�`[	
�u
�'���+3V�����&0tb�y �']:Đ!��=~��I@��k�� 
�'��z�������b 
pl��':�@*LZ@is���
�n��'���[�n�,LV|\QdE�vȸ��'�:@��bԭy���s�ƤXY( �'z����*�<d�&��C�Q+dP<P
�'�~X#�׌U�:��FF� e���	�'E0�sN�h���S�L�a�'dv�Itn�v��P����2�%
�'�H�xA��\�	�q%Bq�	�'�T=�s�]�e�<�a�(1��-�'�4�e��R>��M�-�|Z�'S�F��b��h�F&_A�� �'iF]r��{�"��UM^�'��<��'u�8Xs ��cP�͹�hޞ��)��'���{�� =W�L���&E% fV[�'����ƿ?6� �M��.̉�'g��[� �)}���8�:4P���'�r��\,��V��~xj���4�y�&��;p@i�C&.G��}�Q��y��M�s�j��<�����޾�y�/��jlxZ�T�,�`o�y��?f�]��!q�
	��V��y���4N`��B�.Z�rB,��܄�y
� PtH��ӈEZ:��l t�J*O��B�ټ.����Y������'�]R�h�I��	�������'��(��E[D�n���cV��T��'C��q��59bJh93��VIn���'rep��(��A%KI����Qb\���>��:=�6�k���P��ȩT�[I�<��i�5B�Vk4g
��"���/�E�kv�c#a'���v���8.<���H�)S�	8E"O 8� �s��j'�;(M����@�gb}p �>	@?�gy�H�I�FI���)~Z��k��y��ńW�2ų�,�X����M;c�X\H�n�>ƾ���uf`ɡC�)�����ƴ�뉻g<	�DcD:3/��(��Hw捋"�tLi#"4"!򄊆5���8�d۟kˎEѵ����qO����C�	K^:���iT�
��s�XG�vY���E�w�!�$Ѽll��b� 8A����*���F��"�U�T�|�'sn��T%�h'T(2UA�b�옣�'"�  �N}�#�Vd�,��aZXJ�!Ԇ�0>iw���_1���ɑ1mT�Y�G\��xb4��sQ>�7O�rg��R��a���p0n��"O�e�u* ����a��@����C���=����%6�bF
�+��ɻ�n�K3J��@�ȓJ|x0�D�͠��ț��t�B)��ǇHEqO�}���&�9�F�$S$��5��7��ȓ4�ެTI����cf"Q��}��&�L��տ^�9�BAO�mB&�ȓo�H8J��@?v2�r@FCx�PԇȓsHȍ	��0%��A��,�v�B)��t̠�E���~���M_0Xl�����8Ӏ�/-Z>�*�bW�⨇��0-8&n��V�0,�l�R�Q�ȓ.UB�(Y�O(��A)�Y�ȓE��y ���%H�\�*T��p��ȓ;�1���@>@v�B���Z<�ȓ�� ���S�|�b���69������F�.j��0*��(T:���P�0��"6���9���u�hM��i���t)�����Ղժ3!�4���2�*��
�H�yBB@� /�|��;K�ɪ���}�\�@!`����0~����L�A�l[�m�%s|��ȓlWb�S�A\�t�kFNݕ	����s��} �f6�[%/�	���ȓ�n�x KڢE�As7��uL���!�H���-z<~p4�ZѤd�ȓF��t��lǇ����<y:p)��2�l��U$Y�yzT���{8�H��1}(��y�f�����VY�Q�<�	 �QV�mh#gS�z�n,�w�{̓l�H��Ө�t�LH�s.ҳ �D��ȓa{�:��ǟC�H��(�65&���/o��в�ӂ�A�3E5�6ń�NaTt�T�udX9"5��H�R�<�v��<Oڮ��`��(�8���C�<�,[�
P�l��"º.�v����x�<��$�cܪ\����6%}F����L�=mK�"<�'��	�T2R�2q��7kפ��^h�@T.�>����5k���I"rq����B�ɟ��$�L��<)LԬGM���W��2Ph@�d㓌B��I��)�&_�S�O+�jS�K;wn]����;�\D*�O�زD�)§r/�����56H���pc��I�dH�P��<E���\M��;�/dw�Y�1�ʛ{*M��ө_k�l����d̂1ؕLE�b&֣<!vB=�b� 6�RU^�2�j'��Ѡ�$��(O�Op�<���Q��h�d��~3�xH>�y��3� ZE!��*o�i�FT�p4p" ��>I�O�Y�S�dl�(6�6mC�aXA)��X@@M��"��`y�hTaA&
M�ĂM���6��L�����|j7) m�N<�� c&Z0��LR}b���o�;��4g됢�@B�		��) ���O�� �͔�%������1���t`��<�	�'(�QQ�..'n,�e@LW�d��@�r��b�f���de
v>M��隍�U���7ETtL��䏱WҼp�v���,��C�$~���'�H��t("c43�2�����	Z��rZ���0.�#�qOQ>řB��06J����8� ����OL�s���ڸ���"0�.��Z
�xIF)�\J�(&B�?ᰝ�=��'E�ɳ'�0E����iCt�Y4��4!���?�'�NA�`G(B~<e�V��a�&�	�'�<\�@��'|̠$H�ٗ`Q x	�'�N\i�+�4�&�����R�� ��'��D�߻�<����{�=Z�'�X�14��.4�<YR�N0+r�A��'�h���L�.I��A���D�'�R���'k8р�G�/�8)����A[�'m��G*��R@�!��J-{�'�!�b�כg�h���ƋS�H�	�'�[ H��5�9y��	4&�|z	�'�P����#�\����
&�֥K	�'r>�J��N�:���A ���h�	�';j�@!,D&���:AoG�Z����'N���pi��4���O��U���'��h���Mf4�⤭�8bT�S�'�~䉳��1n.n��$�`�.-j�'�x�c?$��@�ӈ�,U�t(c�'t���8n�Na�#�P�EO���
�'%(�;�H8�����
b���
�'����ɱ#�cw�݌X:Q8
�'�ܵÑ`�#g�4yuC��s�q�
�'�P���<X��9�D
��<�	�'�����N�"�b���@ ���(�'S�X§0R�9(�k	 k�i��'[((�2�kn������W,����'邼�7A��@c𕰥�Q�DXָR�'�Ab�M4�L�z�8g28�
�'V��� O5' h����X,4�@�2�'�xU����5#2HJ�㌈Zj��'��i�F�Vږ�JW"2�8%P�'�@��ǃ9W��ɶ��h��|�
�'z�M�dH@�}=�x�%ُY����	�'������=����e�T��D 	�'hyk�NY�hlT�!�D�IJ���'��	��J�)� 8˲	�{�$�'�>0vL� Q�H�Bu�
�zf:p �'"�0��\���h�$pJ�Y�'������T1��;���7V�i��'����+�n����͌��y��'v$���T�����~`�E
�'9>L�P�.z�E�����BDٺ�yB��|μA�嬜�� ��,F�yb�%-2���aE֣N�;�H��yD�n4~����?9:ԫ���y�-��{��4�
m��-��y�㐡16ʁ�æ0�U�����yr�-@����z����(F��yRř�B{�r#��&L\d�V�3�yB�ޝ)A���u��-�QxsI*�y�B���ҹ� I�\�<%c�!D��y�j�8@���a���\��A`dĽ�y��T�	t��{�ЄUy���Ǥ8�y�%,O�����I��L�7��'�y�N�8�B�"U���8H� ��V"�y
� xh�g�Xi����Pc���"O
�d	5E[ e�ý!O2P��"Olٰ��Y}ŋ��L�,���"O��spI�c�(��fD��
�(�8B"O�`�����N3NECp�ō1�
,��"O�i�uO��]zJC'��"]d=�"O8�8�œ���I��C b�ʝ�!"O(5��+> I�b[�
�*�p�"O����H�-s�mT�Hs���"OD���ʟ"A@ٔ��i,�z"O�A���0���'2\�Dإ"O�M�P(S���C�W�?�>��"O��� ��c��y$�<@v� [�"OqW�5^͢����QZj!��"OJ�ȳb�?�x�BB0{E�"O
�I%���.����5X�8�"O���C.H��Z��1 ޚw��1��"O$�(%���C���)��d���
3"O�,�s& +����9U�ܖ(�y҅ҏk%�D�dNI�SSJ��0�ȱ�y"l�2	mڄ�V_d �� �y��I+��b���h@�wD��y��^	@p��ғ� ���7�y(�@�R�"Ӣ!vp@��fJ��y�$ђ'�4�c �WŤXzk�y"L�G0���)�:��i�����y�NԤ7�{�i��d����0�՝�yB��:zX�xA��Zהa�P�$�yr�܆��)q��JY{�I��m
��y�D!2�̤��N=z`C֯K��yr�Z��y鐉9[��kUEM$�ybI�[�����;4*.�E��0�y�#�hy��s׀U���`� -�y2B�83���P"k�J��$z��A��y��'	�lې���@�l�����y�lх&��S�̅�2�ڤa��y��(X��[Y�����O�m��s׆(��̘(`��q'�SX���ȓ8�԰���f���n4�8p�ȓA�
H�enk[�(�eoO�[�乆��d��P �=Rݸ�g)V  en���x�U�"��	#�q�*=b� �ȓ�D�`�(ٌk��X1NB;d�ņ�Wb��E/��?�n!B�*I5�$!��H�r�%U!�:��α�Pu�ȓ1�H괉S�v&�,��	*-JY�ȓ1-X5IF�ې�pJl��k V�<q �Cu�r�:f��+O����S�<��,I#�r'��*SP\��PP�<QVLS�B�D����Nؠ����r�<q��ߜ*&��R��
�'z\y�/g�<!��۵�4 2��n4�Bq��h�<�RUX'ܽ30i�VO��ҡ{�<����*DZ��3�&�6���C'�\�<IQ�ܕn1* hfL�cَ����r�<��ܕjXTQU�ۃx&t�jŀ^Y�<���j���*Z�(�2h^�<���-�:�:��Q=jt�RR�[�<i�FՃ%�X�tn�?YD��b�AM�<�À�9wc�j"�B�.,N�:���E�<i MP�'��t�ufK+GX쐂,�A�<�tEҡ �4$��l�}l\���G�<V�߻��]�CBN�V�%ip��@�<9D#�9M'�q��'}`��7 �z�<� H C%�W3?rF���Q�l|#f"Ot��H�4z�
�ɐ��42pf���"O>4�%�ȅk��4Qt	D*��D�"O����^��!*� �3L�%+s"O\��*��)��Q*qIQ<q"O0�Ѐ�g`�Z���YKn��S"Oz���
.cв��@�C$/�=P�"O�qBuI�<&�N�)���o��\�p"O
�F � �Db׉�&�����"Oʜ�QC�#P���V.K5b�l@��"Oĵ��EC�E���΅,1p&�"O�e�v��.s
��rPǀ,"Tj�Q5"O5�C^� ��q34��2io�չ�"O��D �/��i'���M{���@*Oƭ�-�*�&a
W�!<��k�'�8e0�(ձB� ��f��	���'�yae�[�1X��T�X�4��')"%IT�Y��;SK�C�'���q�B�0I<�bsF	1}��+�'�>�Ɇ�A'/���P �кv�R��'�&��bMe:iÚhxq�	�'o�9Ҳ+L;$)6����޷b&�%�	�'���Ä�L�:+�x���ĕ`���"�'�t���c��k���UZ�n8��'�8����B�uI�|	 iU)&�\���'B�Dcg�4%z3R��qT|��'*]�Ao��8�����h�3K��h��'�̉����YC���B��DLRE �'��`h1��7��x"A�̊C&�s�'�� y�
[+C&�������U��'��I�AeɭH���J���
�T��'����������烽�p��yz���C7:R��@��ɀ����T|���t�a#B^�PM¦�}�<I"%[%G�:5jԋ��}���jM�<��$�	>^��8�D�K�b��3��K�<��+E��� t��&pJiyB��~�<9�Ꮢ=�� ���# �|���͟N�<Q$"IH�	�J�1�D�#��@�<��(\�'��Q�"О9Ĭ�r`Fs�<9�J`�����d�ht@'Fs�<aU$P �v��s/�H� �ekf�<�K��1S��s�Ǝq��Y��Mj�<����s���r��%^>𰙇��h�<���:�&�0�	 w��q	&E�d�<�Í�fq�]�� �V�Z,�3�G�<ar���&����������!��7�yRd��d��%��5`��y�G��p�`P9V�S�<�����y2��L
)�fJF�FZ�L��Q��y�{�\�T�R�@(���%�Y��y�k�,P���bI�g	2d�-��y�$Xk]$� �܅XA���U�J��y�S��mB�+L�M:屵���y"��u���a�E�	G�����Ґ�y��ۦ
;�P��N� #K��y�Ʉ*<�f�"A/\)CV�]��y�թh]%�"|�V��ugP �yr�t���'��u��PiԷ�y�n�4x���i�
~S�ukd)@>�yr�ԗe.��oޥs��٘���yBM̭����N��8t�#6	O��y2��� C��2.t$������yr�W� ��"�dA%����@��y
� ��fi�N�N��r�<d�a�B"O��r���'���E��VN "O��#�X�Y�`�!E�?YM`"�"OR�z��]�2
T{U#92,ؐ�"O|0�aJ"\�^ )���"w��"O��; �(@�Ax�A�"��tr�"O���ȅ�"R2nYJ"O�%�@Fޔ[�x�����l�,t��"OXt�"Ƃ�F��Cw��G��w"O&��PK� A^0I�A�)^x��"O�=9�-�	���v��{	F�S�"O�T�0f��D�d��O�"^&<r�"O<��/@7�P��5�;�݃"O��G]W�����.9M��M"�"Ol���   ��     K  �    �*  �5  _A  OM  �X  2d  Bo  
{  �  ��  �  �  ��  0�  F�  ��  ��  �  [�  ��  �  ��  
�  ��    x � [ �   U& q- >4 �: YC �L XS X[ �c 	k Uq �w �} d~  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR��D�J���ӳ] �K��F/]$	����kϊB��.p2:d�a�,��������=QÓh�D}*���\�<�{ĥ��1	bq�� U&�2�A˼m2��v��$&����
rdk�A�)!��T��ΣT�8��re�q���W4O ��Z���+�'�δ+Rh��Zc�,��D ��2�S��f��zA�QW1�ɢ�݈�yB�S��n�A��M)3|��
I�v6�=E��ULD�S��"�l�B�C�tgZH�ȓp�(8�6̎��.��7�(1�І�_�%�l�-�w�K����ȓ{��4���`��n+h,�ȓd�Y9`X�^�zQ0QN�GU�ȓP~�����+���
u����5)�ذ���
T
���A�N+���F���c�H�h�>�Io:[�M�ȓ���G���,�+�T�g�0��ȓvU�M	���}0�P;�/a�f��ȓi����P�C*r���� T/jt��ȓ7��0�R�#!�X\�4�c*)�ȓ#���H��&l��:�"?r�����na��جT�0��j3R��܇�Z�ڜ�B ��w7��1��X2���ȓY���K�K<�fX�&�VL	�ȓe˜,�ӨN�Tu2tX��ĭ[NrP�ȓ�x�1m�(H��dϰ:�����4x�M*O�����,�\��>�8� 'ְ%?�8�3��t�$(�ȓy_��Q`&��fut�@d@Ϊ>�-��qXXգ�
�?Q�����'����Q�հ <A\ ��j��#o�0��Z����-�;�`��q��-/ y��g�&]6HK�Q �/I�����"D����@�,c�vh��F�<��"�g3D����l�Z3���^2CG0D���Р� 'Ava���ƴ�V�1��/D��A��� &C�5��gļTzJ�7l-D���rF�+%�(:��_�Tl��7D�`)���6 e��@����B����+D���a"ϑ"���b�C[t�$��s�*D�pڳ�& �*��e�لF]y�U�&D�d1�-q���/�rߖ �&D����oH�B����w��JAn`�.(D��:�`
q~��Kq�^>2\��!T�XCe]��H�Z�@5h���2"O�M��4l�d�
׃��8�ndñ"O�1b�b4��-	c�σc�4��"OH�y���ov�y���D�s�jU�"O0<"�*��0@p��-b�
��"O>`��7`��ܱ� ˅8:3"O��S��=ǰ�Y%-��N���"O� &��'��=y�~���L����2@"OT�	���Q'�Q0JI)RXIw"O��KD�5�F��(N;( R"O��#R��39���(ٯi�4A�"Or�PVꜴ-c��e�؞
�����'B�'}B�'��'o�'���'
&p�k��8�5i��3O�AP3�'�R�'U��'�"�'.��'E��'�Ќ
a��R�`A!�D�K�^���')��'�"�'���'�r�'���''�y3���o��@3����3��'��'�b�'�"�'�b�'�b�'Bh�CQ�S��)en���K�'A��'+R�'�B�'�b�'���'ONI�GXt�"�J%Cۓ�8���'o�')��'D��'�B�'���'aV [c�]�DJ�)�����bD�'���'�R�'���'2��'���'��$��D��ߠ��4*Ol!6�'Q"�'�B�'�B�'�R�'���'_�	��e�,y5���U������'���'�"�'*"�'�2�'r�'������ė/*��;�)��c�u���'r�'���'\�'<��'�'�3P�)-X(�q�fA�����'��'�B�'���'n��'��'Ԕ9y�HG�<�����dݷ6�bLH��'��'WR�'2�'���'�2�'�F���+��: 4��e�e�~ ���'���'$"�'[B�'�NvӮ���O��	U�wY����^�!�Ȭ��xyB�'h�)�3?�i^�ik��M-gYV���#M�+g�����"����ڦ��?��<q�zXU�C��W>�B�b�7A�����?yt`E��Mk�O��S��J?�7�7eD�G���^�,ٕ�-��ş(�'��>-�C���
�o؄p�!u��M;�A���O$L7=�28�jS�	Y�lN1fXp��r#�O��D{�ק�O���ºiE�����\#�Q�I>)�PdN x&�$m����E�=�'�? 
�(��e$(���׎��<!(O��O�@mZ�?�"c��9��]�bKB陁*$��`��X���I���I�<�O�`e���̞���Q��٩2&�,��O��K�rf@Q���?Y�b�OTx��ꖂ��#���(:�|�q�a�<Q*O~��s�,�wfP�<\��o Ԁ!R�c��ڴ�b��'��7�&�i>9��ƚ�L>j$���S�����l���I�d��!\�`oi~R5�da�Sk���P#C
5i�E���&n��ꢘ|�U��ʟ��	Пh���|��� =!nJP�VkW� t�ەIAyrA�O.���'��'V��y��;���x�`H�IW��+����_I��DX�v�x�*�$���?��SgT8��	�^u�#C`�H�IS.�����542���7�2	��f'�'!��0�ڵ��$N0KWxAx`JVU6����?I��?���|j,O�n�<vHR��I,
�<��*̫4��+0ρ�C,,��	�MC�2�>�#�iN 7M�Ŧ�+@LAzGX�5N�i@�����+F�l��<!m��u��8g ������z���������"d�4�Y�E�0�%� ��<I���?���?i���?����,߬��dJ �L{k�p�4F[�5���'���f��1�6�t�d٦�$�({%��,OE�����&O�8�3
2�䓈?���|�E+���M��O��]wx�b!N)˦�����=�F� �G�O�t�*O��n�iy�OC�'���(M)�]�2(��J�&q ���"�'�剂�M��e~	�I�$��P���O;d�&�b�̡���.6����Y}
l��m�"���|b�'f�j�q۝��,�$�^R��|ɗ�.ъ`��ML~~�}�y��'h�i�'�wH�z�(�W#E�	�h�Iրt���'��'���tR��ݴ!�H���"e���C�
KI����i��?Y���F�'�'oh��?��o�g�����Aպ'x��""<�?A��i;z��D�iC�c>}��f͆�����j稄�I�|��e ��^@:P�)�M#*O��$�Op���Ol���O˧n��ӐgF�fC�
'K�'���ĵiʂ����'�"�'��O�ҡr��2�{%,J���c��0�� Cv�'P�fi;���(�D}��;OzaׇG ��ٸ7K��I�A�P2Ov 0R���?��Ĺ<��i��i>�I�iH��x�M�QyP!�r��>�*��	��D�I���'G:6-��f�$�O���ƣw��t��)=N� CӉ4h�,+�O�qm�M+��x��
�\�x�h˞]�l�M����іͫA�����I"�u�I̟����'���$Bڭ9\���G���].����'<r�'R�'	�>�]�d�p�����?ZZ\z��U�s���I������*���OL,oO�Ӽ#SG\�B�`���8qx8Y�R�<)���?��i�x���i���=�,1C�O��ףJ@5�����^�1㐅Py��oӲ��|*��?)���?��#���d�[=��P[�-A�it\��*Or o�2Z�E��֟\��_��֟�#�ڋx��R��)'�.�@E�[/���O���j�i>=�	�?"�O��>DaG��mdQ+ԧ\82�����-?�F�E�{e���^���Z�՗'�H��W�V��4�3�K�dY��S��',R�'�B���S��c�46�F����-@"mx1�+k6�����8I�D���8ћ6�d�ty��'���ehӒ	D��.-�`�ǣ�F�[F�Y*)�7�r���ɥw�(ut�O%��H����� �!��a<{�4��DL������7O����O����O��d�O��?�r#�T����憭V/��ٟ��	���ߴ7~��O�67�>��S�*��𢁓b��,9ԏU��2�O�4m��M�'�
�`ٴ�y���n��$Z�BT�r�L�R�^�A�|�7�X&H�)�u�O:��'�r�'�r�'̜u�c��2k�\�sgϝlE�U���'Q�T��ܴZr���?����i �W���z�l��̕Cv��;6�	����O��D,��?I�g Y�VQP�	!$ �q�LТ"EX�{`���4�֦���ĀSA?	O>	`k�	2���̰,�����)�?I��?	���?�|Z+O��o#��|� W#l�j�)\���a�GmN������MӎҪ�>���nm��*3M�~�x��*�m����?q����M��O�LS����zI?I�ê�(.��82� M|�5��k���'�'���'%��'�S��4��2(МE�`�f��'ވY۴M+z���
ش�?9H~ΓM��w44ѵF��]n��w��*n}|����'+Җ|���e��EY�4Or%�F��5d��wm��0,��1O�p:S#�.�~�|�[�@���kFD�QlΉ�!��EӠY/�۟��I��8�IPyB*~ӒaBG�O����O�P���.�(0��'���xrO1�������O��d%������Đ&��#Qꩩ�(_�V��I�(�``����+K~��`�������l�GM^#St�+6bϡe��9�I������IT��yg�W	t�� �	Q84Ś�Ķ[���f�zH�5#�O�������?�;�����üT�x�ʳ���p�r��Nӛ��s�b�oڄFz^�l��<I�:���������'ϫ~"����*'����t�K�����4���D�O����O��W�)�fŊg�r$�B�!&˓Yb�*�P�'�����'�riS���5>��i�dh�
F���h�>���?�H>ͧ�?�����	j��q�pi�:�֘;��A
@�X�'v"�0����R�|2]�H������L�{�RR�܅�@��������I���@y2�~�R�:��O�)c��Ĉ/YB�@�c�&l���O��l���$���O��d�O����,Pg~4;�� ��
œ�v�Y1G�?��3O����B+�*��L���?i���a�5N�6/Bif�!�H����|����x�I퟈�IO���D���8Yk�E*ƍU1b���?��G��f�X���$\ڦ&�� &�Ns����mO
D�&����I�I����i>E���Xʦ%�'.���K�CM\萗���4���O�X�������4� �d�O�$�`�4\�@2*d�2g%�O��d�O,�u������_O������O�rH@��b�Vy�Ř�'���j�Oĥ�'HR�'�ɧ���'���au
51���(��m�e��ϝVȌ}���i�rʓ�.�:�	\�	��`��=]zPY����"��I�L�	���)�S}y�moӮ+D�-z��tCݡ8^�h�2�хp@�	��M��2�>y��#�dls�l�,O
.�h7�Ԗv��(9���?9v	��MK�O� +%�ׂ��O:�ٚ�G�
�b��b�'����'~��˟�Iڟl���(�	l�4jͦ�����*ʹ^�����̑%�r6-&*U�����T��y�ǜ4�$�˧����:�s��&�b�'Qɧ�D�'b�䊥.$�f4O|�C�I��c���m��#�2O6�JJ8�~�|U����Q
�=�ʙ�s�EX���9���������4��Xy�e�&�����O��D�O!�Sd����q�c�SJD��0�����d¦���4J�'m���1 ?:p�� J\+�>�ڟ'J� G	,���������Hh�V����ҷ2 �E��lT�KNMXBИ'tF���O,�d�On�D1�'�?q�(ю��Qc3��"� ���]�?�ÿi�6|�g�'�ңq����1*%>h (��S��U��^�u��.�M�P�il�7MS.9/�7�m�8�	q��z��O1>�3��ѿ�ֱjp�D�)C��}�Ey�O�r�'#�'���̆-�*�I�gW���a��cД@�	��M+����?��?�K~
�	8 j-[Y֨[DRsO&u��P���ڴuB��)�4������X��t($�"X"@�Zv���(�a�R���c�Kt[��D�IQyR΋�\�p v�ͶIߪ���m�s���'�'��O�剨�MCBω��?�m�>l&�P!C�V�+�D� 4�Z��?D�ib�O���'7B�'~��Ob����C�x�@h=1���0%�i��ɡ-�� �ҟ䒟��/YV��1���9#�� ��6��d�O��$�O[l�ܟ<�	}���0Lbfd�>`8h6�ņo\fLB���?Y��C��6�����'�t6�1���X��X�V���1�]� A�F|ܹ%�`�ش��F�Oa��{�i}�D�OƱQ��9�CLׁ<�}�oD�X�,(;��'�t$�<����'��'r2�iW�ٜ�T0�GUc8���'{"R����4w�v�����?�����IU2v=|�Sbn\�����¸d��	���Z���Y�4����)J�����!+�˂��|T���5�JT��h �j�3��i>�0�'l��%� AF�����U�����.]ܟ���ПH���b>��'47-ц:z�b�N�(t���˅�r٪1���x�ߴ��'��듪?��ic}Dr�����^	�� ����?�e�ܗ�M��O��!֣B<��π �Y0�@_9B�&`7�&F����R1O���?���?A���?A����I=F-p[Ч��@���t-��o��n6Y5����ן��	S�Sן������e��#�6����@?)8�U����%�?������|
��?�6I�5�M+�'W�X��$ɒ;����"Ot��j�'K�����Xi?�I>�(Ox�D�O����-HrIn���(�g�O��d�O\���<d�i�x�	��'b"�'k: �`RM�9Q�A��9���'�'��듵?	���$.4��"�al�颥n
�6����?��旮f��-�ڴ$C�I�?#4�O���u��9a!�����]+׎��2@����O����O��;�'�?����jh	Q�ʪP-�YC '�?���i2�QU�')��s�.��]�W_h���+�-�}��=9��	ʟ��	ǟ@�!��٦�uwW�9�ɐ-�h�%`��mrr!a%!�|���Oz��?���?a��?��P|�!�0��P���`�ת��",O�l� �T=�I�P�IE�s�P�rN�8+�!��-�*=�*U�߁���OV��"��ɔ�7�(1t�4h>�vfI�*��]�U�n��0�'H��D��m?)N>.O԰[K��[D��R�PMrY�L�OH���O��D�O�	�<�t�iJd�@��'l,u#b�TB������,@p���'7-(�ɗ����O����O8��X9ci�-p�/�J��� ��/{�7mc�x�	>U}�!xڟ>˓���W���X�,�e�bYx���>��?!��?y��?)���O����/�\GZ�	Wl��b}�=��P�8�ɡ�MK�*N�|��
��f�|�4��\�Rm�k��i%��3]+�'�"�����38�F���4	�4�R+K�kYR��E��+!��H%��c?�H>1(O"���OT���Oܐ��`�:�0F��$k�C�����O�˓<��o�0<r�'d�S>���L7O��YY'�Բ4�H:2�:?)�^�H����|'���CD���$�r*�!�V�bo�=D���Y����Mr.O����"�~r�|�/�$*�`eH���
޸�@/2&�2�'�B�'����T����4qsz�a�#M8����M�Nb�(�`���D��Q�?�\���I ����4��*gr���	֟�q������Γ����4�	�<q�g*6�hD�	8! kW��<A+Oz���Of�D�OD���O�˧%_�M���ʀf�x�M�/K�d@аi挤��'1��'M��yR|���#
L޸�ъˢM�b�_� h.���O��O1��(�+x�4扁o��")��m�a�F V-OA��*�"�҆�O��OJ˓�?i��sH�+ѡ�B��ʅ��<��� ��?1��?Y+O�<m��(�h�Iڟ��'lHI!E�'42��h�c��n0�?Y�P�H�	ǟ�$�����T\�ą���+��M�Մ&?3C��3r�s�4��Od���?�D�5����+H�H�pM�,,��d�OP�$�O��2ڧ�?��P�|�@���G�}��`���׊�?�]8��������4���ygo�:XRQc�v�kWL� �yR�'���'�S��i���O9���,�����	-�}"u��r��C��(	��'��i>�������џ�I���`�&IT�]���J�|�ĕ'ـ7��"bU���O��3��1Z>�b�K�O�N�ѷiӊ��P��O�xn��M1�x�Of���ON���̘V�(�Fi��6Lv���\;,Τ��O���o�9�?�0�İ<�A��bA�G�2ʚ-��F�?9��?����?ͧ��d�]�w��͟ p$0q�e!�By*fM������4�?�J>�V�d�ߴ	��&�yӸ|��� �e�B�H�#���:u.�MӚ'V���E���8��dퟲ�.�5G��|x�oR���(���'X��'1��'�2�'�����Ӭ,*(\ahN�r�0��c�O<���OjLm�<�b�#՛�|�L�4҈;j�8=��Cw�ѩa��O�Yo�-�M�'�vLߴ��$��i��5
�<6�Ph0v� "o�uP���?1�/%��<ͧ�?���?Q�7?T�K�&�;��0%ꗧ�?I��������b��Jy��'���?#=�U���6v��v��&,t2�9n��֟��IT�)� K�3z��a�����"<�m:c��
��<S��*\�l����-�ȟ��A�|���M�T��ERĽ���24L�'#��'���T�d(޴h5�	r�T�%&bh�U��7V	��K0n�`~2�p�T��*�OR�䝖
� M�b*T�ʤ����8��O��Gi�P��ӟ`�D��T���<��G�YE2@��oXi��(�1��<�-O��$�O��D�O,���O4ʧi��cmC7Y�r���OV�|��i⵳i� ��'��'���y�Jr��Q�F|z��lS.<
Y�K�m�����O �O���O��DZc��7�{����%�+*_�,��`�$x�����%g������[��,��<ͧ�?Q�gW7F�~�R�C���LR� ��?���?�����$���	Bg�e���۟���e�A��E`���q��a��s?��ܟ���E�x�D�bM
�RGFxVa�4�ŗ��)b����\nZq�'[6���ş�2T��[�tиC��6'���[�@U埴��H�����G���'K~<k�M�J�VU���O5p?*�t�'��7��]^���O0�l�g�Ӽ۳�m�tP�I_�@���*��E�<���iT:7W��! cn^Ϧ���?a�-�*~H��B�? �H�"b�7q�敊�+ �1��*���<ͧ�?���?9���?�U(�zr*�Å���۶��K��d�Ʀ�@�wy��'��O����58��@�r��i�E+�33L�
]�v��x�$���?�Ӿ���B.l��-�ǣػ8=�O� =��u3Bq�tG�OR��M>�,O�ȉ�ڻ���Q�k,:��i"�"�OZ���OJ�d�O�I�<1'�iӤ,K�7� V`�s��X���@��KC�'Z�6�;�I���D��A��4n��6���2TO��x�̙�&�ԑa��i��I3gj��¥�O�q�N�N	%��tp7M��i�� �F+��}��$�Od���O���O���+��	~J(�����F�ǧO�r �	��l����M��f��$�ͦ�&��rb+X ���������u��#Zm�֟��i>���fB�Y�u�-X>0�@ňC�./� ��ÁGf���O�O���?����?I��2Z�L�[6�m�&Am���?,O2-oڬN������h��w��\w�R��D�Ng�$X@��"���R]}B�'�|ʟ��"EŬ?�NY�Ѭ�^h��xg*.RȠ� �}�~5����&MD?!L>ID�"�����⇯+b��A���(�?9��?	���?�|(OTMlZ�U&��I�#�\Mp���8$ㆁ[Xy��y�8�hp�O���<5k&AST��i����E��{���D�O�B�Ma����K"WM]����P����KC&�Ze#B+.HԵ�7�y�`�'���'���'���'N�ӟl�<�#v�\�=XH��G"[�,#v�X�48������?!���O~�6=���c,C�W�ذ)rG��	�P4QU�O2��-��I8O��6�~���� t�T��>6�z�{�p������A��d6�Ĵ<���?Ѧ"H�r$��h@H�}F �ɰ�?���?����ݦ)��K�ԟ��	��@�N�?(�H�P$I� 6����`�T��q���� ��l�	P��uS-D07ߠ���2Q���	���s�-s��n������z���'12O��nH�s��(�Ց 땩\�r�'"�'������R�eՓxJ	��"Skd�qh��$�438XH��?���i�O�!L����F�+����f!�C������ش+����$u��F��H����}��$�ު<�Z�bB��R٩��>a��&�̕����']B�'3��'Ė�� E�i���%jH�N��P�_�\��4=�h�h��?����?��C�2=�`0��NJ��ݡ�g�C���	�M���i\�O1�Z`QA��K�&�Ԁ�	_^`��J5[jI�䜟����Y)mrəD�	Sy�/g���h�"DU�Tը��Q�0��'2�' �O��	 �M�W��?Q�>�|�����$~���L��?!q�i��O��'��6M�Φ�8ڴT�Nh�׈�u{��A@&eZ��f����Ms�O��;X�@��6�S�ߙi��I?Qn�y!����crL%�'�|����ҟd�I���	����B蜑-�Ȕ�U���X�T���G8�?���?�G�iN
�O\b�|��O���nͮO��`�j��9�E�v�9�d�O����OD�QpӾ�Id� .�+��<+� {a�h��
��)pj��~�|�_�D�I��	��<#�T�th����/X��m:'�۟���_y��v�hmh���O����O$�'?�D�� n�x:|�1M����'�>�]���%~�(�'��=\� Ţ+��XӔjDv~)�У��N�D]*�i~�O�����R��'7@���J�?�ΘV��> �� ��'���'�"���O��	�M#A@�����,K�B� �7��*��5���?�Ƹi��O9�'�<7-96�݂��
�y�ȍ�W�Y�)�ҕoڷ�M�v�Ĥ�M;�O��Z���
��O?	��Z�\} �}���s�z�H�'yB�'���'3R�'��S�J�&���S�x���o�3�~�:޴_S�p�-O��$=�	�OJ�mz����-(�Q�Ņ�i�Hlx��6�M��irPO���i�%4�6�x��`�k�;lE�!J©���в'"v����ۤ&�B�Am�Idy�ObKJ�xh�5ɂ�N�EB�L��ÃK�B�'��'(�Ʌ�M;�L�"�?a���?a�,ɼ@�D��W�"M>�� �J���'\듀?����'�Йtn��ѥ��$z9`�' H�c��M�r踋���������'��"0�P(e:����m�j49"�'�b�'�2�'��>����a?dA�����k�FA0�z8�I��MCvkW��?��h��6�4�B��u���2Hr���@��
�4O���O��Ĉ 8O�6�b�8��
'���E�O���w��"I?�8��yɸ��ӗ56�O���|���?����?���,�� Q+7�8���o��\�~� )OZ�n�&�&��IȟT��X��J���)��<��y�C�C6/X�0�[�������$�b>�qqN$���0a�%S�ju�@%�h��SQ)5?���@,,���S*����!X<Q��R�����#IG�}BV��O\���O�4���rs��j̧�y�&��f��&E�E_6MK� _��y�)v� �8��O����O��d
�C �p1i<ul�ĪG@�o�^I�i����ş��;��*0��'��T�w��p�wOܾ�R�rǜ�}����'��'O2�'���'���Q�KЄ=�IUd\�BE"�S"��,����Mˡ��\~�h�@�O�$)�HD1rƸ=��A	���#H+���O��d�O��pӐ���HI2�1� ���g�	��䁡#��~�c���~"�|W��ğ�	Ο,��'�2b"�5���|��Pu�����	}yRӴ��������H��N�0B$5
$i	�1d�h�����$XR}��'O��|ʟ,D�E9�r��r��!�f�s��B�md*�"7jlӪ��|��J���'���&�K5
D�Q�G�q#>	�֬П �Iџ����b>q�',7���X�1qVG]U7��3��x5K���\�ߴ��'����?��H�5H�m��	C}�`U�M��?��Sip ��4��d�K[ry����őY�
����wH�w-!�y2X�������� ��ٟ��O�N%���'�J��d��'���+W�~�|����O����O|��|j�{K��w��Hj��K�(�F����V�p��ȳ��n��ymZ����|Z�'��eH[��M#�'�8�HA�W�!ʺ���hՍ=&��ɝ'�~�b�K����s�|2]���)���`%[��I�O��0�@�ߟ��	��L�I]ybnӠD)��O����O��"J�6H쐖$� T�q�.�I���D����ٴA�'*��f�Q( A�PN]�,C�'��҂�̅���R3����3��czV�$�*=�'G6^�:Al��qՀ�D�OP���O�$-ڧ�?�t�69h��A��8p���zA����?���i;��7�'.�zӦ�杹h$��i,��I S�gh��9�M�°i*�6���u�p7l�@��1^*�a��Ob$�1�@�ePj҃/�h{�mC�nL}�IRy�OLR�'l��'�b�~�@�fF�\�T�5NZ�)R�	��M���,�?���?QK~��N�<�A�mL�^l�! �B�>�x^�<�ڴ;���5��i_� T(���)�F����
�����o	�[��I2�0eie�'�ڡ'�l�'�li0j��.��p�ǋ̕R�N-xG�'���'�����Y�8�ٴ7��;�'Kb9�솂GCpI�*ܥauA{�\Λ��ds}��'c��'�nl��[� )f")Ee
9)��H�4�F<O�$J!e����'?����?]�ݮKAN��1�Q�E�j�'�3TZ��	���	ҟ �	⟬��Q�'M�� �� 8� T���,��}����?�����F�M)����'#X7�#��]�V��C�)��1��� ��M&�`�4^M�f�O/\���i���O�E���`��	d��1K� ���8��E�r�O���|���?��88�SMns��C��
�����?I/O��o�A��������ID�4��:F{�H
��ae�!��C���D�r}�|��mڜ���|��'<�^d�4\0Sq� �;���	��V�m��qRS��o~B�OǺ���_+�'N�}!�ƵG�6d!�*� )@P���'a"�'���O��I�M[���RdD�He�W��D�[��1t�2���?���ii�O ��'Kf6͏�o�6H�f�B��T �@�U���d�J@n���J�l��<����سt�����'<z|���O�DZ�Lz���(/zn���'������	۟��	S�4E+e��1�4Q'S��;B�K�0��6�ӝ/�����O��6���O�ymz�}���&yVٲgN�1&�n��G�ߟP��l�i>��I��{��AǦa�|�x�qf��7"k�T����[O0@�f6�|��&�O��M>�*O���OPLde�$v袭��f� _Gu����O����O�D�<� �i���r��'�2�'Q<�Pc-�9q5δBs�	����D�Z}b�'U2�|���X��W,Bv�ɀcL��y��'v~�#���s���O����?	��O�aCf�T!z\6|*�I�;K�X�i���O�����I��P�Ix��yG���$81V�4n� b�(�?bX�	h��ݨ���O���i�?ͻOC���たTx�����6��Γ�?9���?��#޾�M��'�ReYy6\�S$�	X�S�8w�ID,$@�l� U�|r\�����	�����şh3J�2!��;`'�[���p��gyB�j�l�!G'�O6���O���4�$>kp0�2��.A�P�@�P0����'�7����5�I<ͧ���'>O� ��N�5���8����W����a��A����'��eBRR���Z�	ȟ�}�T��7���(X���� �1�:Y	T�Oh��%���6�N*?���Or�I	�{ƌ�<��
�0:��!dO�)=�PI21k�6�?��?���?9A�A��e���h���`�ӗ1PEK��2�����5�����Γ�?!���<>b�2(�������
�Z097B� ?{~��-��0����O����O���O��d�O�Ygb[)O0L[��Ԋw`�����Y�saM�3���P��	�O��dX��%��e|�|
��n>1'�0�����`jb�T���=�C_v� �џT����0�	�|�t�l��<y��r�R0Ì�W���
�^*���&�Ȩ2�X����䓔?�O��'n�%�A�p�HV*�h�ڱʤ��3�|=��0��E�3�4�Dd[A����'WR	i� �Θ�C6����?�:���'��|����b�$�����r�y>��O�R���\8��gGs�0C��),d�`���ΑɛF�����:A�$:�dԁ'�bI���\��q�A#WT�.���O����O��	�<W�i���k�K��(���fM�����s��G46�r�'�7M?��6��d�Ϧiچ��\�	�&]�fl8勆�M���i%��z�iA��]E�m2��O��'p�ao��{*u JY��Γ���O��Oh���Oj�D�|B�DN9~Ar�ш�>N]C�K�E�F �%^#��'�����'�z7=�1#�@�:/������-�\������@ߴGo���O?�5�&�i��� ��c��8q� m���E�D��!7O�B�ї�?��h$�$�<ͧ�?)7�C���q(٥)��]����?���?����$Ѧ%���r�����hP"BF���(�W>s|�`�AOF�3n�I��(��|�=Xe�FmϫB��pQD�B�P�	�\*��#m�fDm�V~B�O�����?i0��m8�\�p�Z�L��?���?���?�����Ov�R
�-6�H�3� ��໅J�O�lZ7$�tv�6�4�L�	�N�

���#'^�O�����9O��$�O��D�%7�6m3?ɗ$� "~���z��C�c#�xs$�+ M'�`�����'[�'��<��\�퉌�`���jE�+���2�[�h۴U�ZX͓�?�����<6�c�n���V8���@ᕿIa����@�	E�i>U�i#����m�~�[ �-Hv���$>w�H�G�iY�I�����C�O�Ob�&565z�F�\I�V�_�( <����?��?a��|�(O
]o;et�2mQ$̚elƯ��0GK_�=1�I��M���k�>	���?	�o*t �l	%�*,��r0@����M3�O��p3��
�(���Μ�b����?H��X�W+V���O���O&���O��� ��=#`�9%üזA��G$~�~��ܟ��I�MK���O~*g�&�O�}� �Z
"U�x��N/"6P���?���O ���O�Ia�g�f������Y`*��8z\5W�=�h����On�Ov��|���?��!D`��٢_���W� {Ȭ�
���?�,OjinZ3I��	�����?���C��I' ��s�T1Q�\2�R�H��Iן��IF�i>��+Nv(����1���� ��EMzm���rߠ�m�g~��OI�e����n��`1-��9�&(R��k�H�����?����?��S�'���֦!����D�8 ���'EO�i��f�P���b�����b}��'g�A�b�9m��ku�ц%�ʼt�'hb풇Z���3O���ļ@�^��O?�	�J��@*v�S1&.-ʆI�/��	ey��'o��'���'��S>q0���wf�`�č�� ��|p����M�s	�?)��?�H~2�&���w���cu���N�)#�E� $��8	Q�'�|�Ozr�'�}øiS��]�K�0!�t�٩i�@4���3O6!�w����~2�|\�H�I���!��B��ẵ�m�~LW��П������IOyfh�n���%�Ot�$�O�	��Ǚ�dO�[A�E	r� X<����$�O�7��I�	$��;��L���;PH��4��������E̘DpmI�!?���?���d���?������0j�t��T��<�?A��?���?���9�>���ʌ'*܈ʒJ� c������OH0o�3Pe��ߟ0sݴ���y7�ԩ.(fxx�GGt^��'坯�~�i:r6�E��	�%PѦ���?�ЪD�%�r��U[���סR%�Z̨���h�fl�M>�(O�I�O�$�O����O��P�y"α �����(C��<!�i��Q!w�'���'��O�2�ώ#Ġ��$�ܧ���a
���	�6z�0D%��S�?��S0U�P��*� }�zaƆ�+h,42F/�8K�6�bW�Y�Tl�O^mL>�,O	b ☴K{�uo��3����Ak�O|�D�O��$�O�)�<��i�ց��'��b��E<x&�q�LB�BA �'�\6�/��<��$٦��4M �fOнF[�h1�ED�p�.��y����6�i_�	�X���O'q����xa��ônH����Ӌ~y�{�<O>�D�O���O����O��?�a"׏B��C#�J�Լz�J\۟�����|�ڴot��ϧ�?��i�'BL+.�� d0i�n\�Xea$���{ݴ�"d�W�M��'��!�r:�@���R�<�]�aBP�]���QeB�ş��c�|2R��ٟ �I؟,���Y�3����&c��-/lQZ�Ɵ���|yr-g�H����O����O$�'�T�*5��;½z�@�)j��P�'Xr�
���Nu�Z$��b��wfS�}�!�բP7�A �;j��Q3@Yk~�O�V��	�V:�'8���L�{j���Ș�S�81���'���'����O��ɞ�M3��D�4x�l<U{赢%(O7�� (���?���i��OB�'��f� �/���"�׶y��T��L�S&6�RЦ9�+���'��d����?}��6@����s�b=�7Ι{��|��9O�ʓ�?!��?!��?������׀;�P��	�@��|�q����EmZ�Mw�=��۟���m��79��w��Y�#?\r$:�)_�#
#��{�"�m���S�'9	:y��4�y2`C�_��Y���U`\��&�y�J]�I�Z��I'��'��i>��I�s��G"��*4�cX ���	П���ɟȔ'@7m_%`J���O����
PT��$> ��`�����c��4!�O\nZ�M���x��!�Vy8��K�Z��8����9��$�1��Īԫv61�$�9��s6���G(G����c�Cw�8d�'�*���O����Ox�D!ڧ�?�� �1��h{0,��W�:���ɛ7�?)�i�����'~"jb�@������p�53PHQV�]���I��M���iZ�7Y�[�7m>?��̝;�i^ �6y9d/;�h%P 1��l8I>q.O��O���OZ���OD��`C�q���jc�7�2|+%��<!�i��@���'"�'��O	r���_}����C�1
��$�[�-TJ��?Q����Ş	 � �vh�"E�H}���3S����~��͖']�$���WT?�O>�+OFysR�ѾZ �|҄����}k �Od���O
���O�)�<1��i��	�'ζ�e*P)b�x�ćW�b!�'�7�,�ɫ���O���O�쩂��1E7d� '��̨�k�._�W��6�(?��nź(z��|��;"��S �#fLJ�(Sg�%|IB�̓�?���?���?�����Ox0IّCL�J����A��R&*\˝'<B�'Q�6M��Y���+�M�J>��	�~���
�/t�M�@������?���|z�ʇ�M3�O��qA�/M��))�m�oq�t��G(�����'b�'s�i>��Iʟ�����za�A
!�P�$i�<5��I��P�'KV6���{���d�O��$�|b�ǂ+6M@�ꔥw.�R⡟_~���>Q��?IH>�O�~�cG��('�\� ��SE������)v.D �Q���4�x�(����O⽋��L+h��yx �N�S�P��1��Oz�$�O��D�O�ɗ�*2����<�ջiI �C���H���*b��::uF�X�䘥�y��'hҗ|�Oo�I��[�F��!���K�R� �@��H͟�����m��<��iCε!ɖ(��9O�Hr/��"���f�Dta54O.˓�?9��?����?�����iA� ��)�3�F�x�v�蓆;��o�.��ϟX���?іO=r��yǤS0?X'�	�k�����j�*,r�'�I՟�џ ���
Ml��<yc͎��"j��د*�,$k#��<a���!V+��	[�ky�O<��ʶT��u�r�^7Cb���Em�*$2�'��'��	��M#��ѡ�?���?�U�R�+���)ԍ�5�,�ȓ��'���?)����:@A��*���#��^�J �'&lT' �8𽐉�t@ҟ��1�'��H���p���L���yٓ�'T�'���'��>���w�pw�����ȿ.�d4V��ӟ�ݴm$�'�7� �i�U:%G�v�@R���o�&� �m����ȟ����7�pMl�R~���	Bi�''��g�KC��@e�}ߌ�{J>Q-O�)�O���O|���O\��s(П^���oQ�8g���ν<	��i[�0C�'���'���X>���|��`�����.��C K�/��ѯO��D�OƒO��OT����wa��aJ�?ĺ�ړ(�8L8�9�D�s���8q�p{$�'즍%� �'����Pg[4�A����6����'r�'R����U�L�޴*](t���Z�����љSU0��N�;�:��� ����'��'P드?!��?	�	�==(I�Ao�:�04�aaG4UkƬ��4�y��'q,��V�S�?y��O��i��NՓ����@��0�
�rᘱ+�6O�$�O ���O���O��?-�a��F��1aG�E������K�h�IӟH�޴8�>}ͧ�?�@�iUW��%H�%�8s�n�}9�IQ�	����	ßT ��W⦩ϓ�?�K��8�
�X�B	�2D�`B��i�`���O ��I>)+O���O����O�y�ǌ�]��Wg��
���s��O~���<I�i��1k��'0��'H�x���Y�fH&"֒�����5u��eF��͟���^�i>����*���z��5$r��f��|�����/Y�	�r�oڒ����LI��'F�'\�xO�4�U���J<M
t�'���'n����OX�ɇ�Jd̟�7��5!/?������O	���������۴��'����?9��JnU
�'��f�G���?���J��E9�4����Ur�g�?��'����2�<QB$9���wW�Dk�'��	��t�I�0��ޟh��[��lӺQإ���H�.nz�B,'f��7m�z���O���8���O$�nz�	��O��{l�	��HJ���@Ɨ8�M�b�i��O1�6�q KvӘ�E%!`��f������<O��r���?1�-���<ͧ�?yeB���@�R�]� L;1�B��?���?i����d��h1��ß�����(KR�� e�1��
S���)AL�p��'��8�Mc�i�rO���:�VD�&�ѓh-�Q�v�����FЇVG�ܡP�6擀TM��ן��D4\TvBN&��9f'���������	��`F���'�VA�'��wP�Ac��cښ�ˤ�';6��-w>�$�O@�n�N�Ӽs��ܫG�u
��C���B���<y���?)��O6� ܴ����B�:���?����5o�Bupv�B�/w�}h��	M�IGyR�'���'Q��'y��ƿ|�ܡ�H��h�@!�����3�MCtG
�?���?AL~��	]:0u��j�HD
�b�\�	�U�T�I��'�b>����ۭ?`���W� ��Yib �sT��l����J�'ƙ��'l�'��z \�AT��e��b�4I�d�	����ğ��i>-�'Q�6��Z���� ��ɁA�C+j�w�R�[���dZަ9�?�W���	ş�ݏw�(Т�D�p��T�R�C��:7��U�'v�
 �F]�H~��;����d��}�F�qcU5�J�ϓ�?a���?����?1���O"����F�r�H�hIъ3YR@��'���'հ7�J��i�Oęn�t�I<0\0:�Ř"�p�3�)<	9��'�,�	��S�'$vml�R~Zwz\�h�ϫJ�H��B( )4�x�c�F��D-�d�<Y��)o�mё��܀��b�-�OЄoZ��M��֟t��K��@1l�r�b�����8rM�����Ox}r�'��|ʟ� h�N��K��(���p7��pLP�1�qG
c�v�����H{?9I>q�a�=@ l���
�b�8BmWx<i��i|�ʀȝ!5��`�$�-�d`�(�$����5�4��'I��?1w�M�sn����̀�l�@���4�?!�5l���ݴ����P�{���?�'c9��R=��T �?��c�'��It�� 
�I�}#��
��T	���M36���?���?��d`l��>r(U�g��K�����.SN@���Of�O1�j\��be�x�	�+EI�@�l	��E�� �0DB�'����P?YL>)/O˓LԼ��(a^�C��8����	/�MS��>�?	��?�U��?7ɖ<�D�	��9�t����'�J��?������Bc\�H%��7#�22���ABH~�o�VQ,����iR<���\b�'���c*pdk�&�Q�ntxL۬�y��Qo���;񂗦UB�h�T��Y�Rls�N-#���O��d��?�;V�p9�ǪU2�cG��PQΓ�?!���?�D��?�Ms�O�J�T�ov�)Ŋ�V ���T�Q7%RZ�%���'xџ؛�J�	�r����$�Q�6?��i�椛p�'���'���=Ѷg��uZ1��i�6�&�9
VS}��'[�|��$�B&8��xG˓#VFt컑��?kH-��i���}U Y"(���&��'{�X�4��&`jl4s�n��`�j)��UY��Gb�+>m��S��/t(�aV`D#�rCz��⟐��Oh���O��ƞ؜���(� Y@��ŝ#Dl`�j���v� ���?E'?��]''z^9`���<��iׇ:_~6��C��DQQ
�j���j���%/R�q�cB՟����Dc�4*�H�O��6�:�d�L�}�ą�7�,��E��o�p�O����O�)ˀ39Z7-6?��{��-�C�&kU�9�6H�{}|�C�����~��|]����ǟd�	����f`@�M�L�M�Y�|�¤T�d�ILy�'b�Z�"@�Ol�D�Oxʧ1�+$ωΑIw�\�*��4�'n�:��6�}��%��'$���WM���,(���E�ehr�]� ��zŌ~~�O!���|��'�\%(���+�܍�w`/,�1��'Yr�'e��OV�I+�M��`ȲE6�yJ�eW<���S��<(C���?1ұip�O*|�'G(7혙07x�ISgLz{J��Ea��i��m-�M���C�M3�ObّWG����M?�1wCkn��b�͝Y>���`�s�$�'v�'O��'^r�'B�� �V��f(֖M3�ԃp�H�[QRa���V������?������?1W��yG��9�3��j��]B������7��֦��M<�|ଞ��M��'� �I��Q�pwjp"�`����t��'lY	������|�V����H��U�c��Z&JX�3dX��J���������jy��u�>]�7��OX�D�O���k�,O.(pe � �l��)�Ɏ��d��� ش��'���[0��<}�A��P�i�����O�d[@oS�����C���?�C��O�#���*_
�ٔ-\+��"��O���O����Oآ}��"q��s/�z�6Y�1#�@���x����O��k4�'�6m&�iީk�����[g�W0$L�=�gc�p��47ꛖLiӜ��n�L�fJ����/���P[s#�g~<�6m�74 L=����4�<�D�O����Ov��8':tє ��NVy
F��3���%�6� �0���'���'��QD/�+�P�80�M�wjP}�6�>���i#�6M�j�)�O59�ʂL|��� m�ڹh�@���N�ڬ�����O��PH>�)O�M�#&�.'�bݘwO3�ڕ{f��O8���OV�$�O�<Ac�iu�H���'���FRZ���lʤO0� p�'�h6+��8���AԦa�ش��$��n{R`˗R8W�tAQO=���P��i��	<Mo`��O�q����8����-p������Y-\����O����O��d�O��� ��Hx~�d��$&�
PD	=ߚ��I��P�ɻ�M�&�|"��K�V�|2�R5	�]���9dp��዇�X�(�Ot��g��i�'>�6- ?�e)�����l�oF	+�I\������O>��N>�)O�I�O����O�����X�ti��K��<">�3�`�O��Ľ<��iB@ӂ�'���'�S6F,� �K	'T'd2�aA21�.�g��I�Mˣ�i=�O�ӂx;�9I��+o�����Vb�9��ht�&1�f!4?�'-�0�D@(��q,H��P�� $O>u�(�X0����?I���?�Ş���ߦiWNK%G\�8�풒��ܓ�քʶX��ɟT��4��'Fb�i'�f�R7C.V$�"�՞y�1ǬXf(7�Dʦu*&�ݦ1�'#R����
�?)��<�"��Zª\�o#�P��9O��?����?���?i���	�}�� ��a�	(������M�~�Tm��@_>`��ڟ��	Q�Sڟ�X����Ū��t�t賑iM&��� CU��rݴT���c3��	ݦT(7�c���#��/0�)���?�B���"m��A���R([��Dy�O�
	e�Υ�.�g���S�/���'���'��	��Mc�γ�?����?��#L�G�^�j�mĶs+��c����'.��w��֌{�ޥ$�� ��"�T#ԡ�K�$���CQ뗐9\�8V	$��;�����C��?���p�8sP"�C׈�ϟl�I���	���E�D�'�:�Ꮾ;�z���A
�(>I0�'XZ6'�8���OX}l�T�Ӽ�n�WI$���T��p��â�<y��i�6m���Uc�)�ަY�'&�1�a��?�"Y�f���p�2Uߐ�y��J>�.O�i�O$���ON�$�O����(X�/��ŚW�Bk9B�!�<a5�ir��!�'.��'��X��勯��H�@S*�T�1�k}�r��,l����Ş5���C��;J "�,ɥ+,,-���hd�p�'RX�X��K�T�T�|�^�0�능R�������72̞i��H ş`����	ß�cyR�f�Y5��O
��p�ۆ|Yp����4W�V�ۆ��OelZO��h�	��M[Ծi�7��!H����1�ɣ'a"�#�D�3��E�|�"�ͦ	�6H�@�>9���;uvɁr���F�'��lrϓ�?)���?q���?!����O���ԑY���lW��X�e�'���'��7͙�|����O�5l�b�"T���.�K���6Q^y0J>Y��Mϧ=S\���4��dp
��p�H�TA!� .�*5�6��c���?��1�D�<�'�?���?)���l.����-
0��2��.�?����\릡��o|��Iǟ��Ox"�`B�݁-���I@.FZ���x�O���'|��'ɧ��	�/ =S�Ǐ�V�в�lř�����F�J�7�>?ͧ	�:��B�	�1�$	���#3&�a���{�R��ğ��Iݟ��)�SKyr+f�n$h��ްT_�E�0-2�L���ַT*���M���>���Zщ	��UD�!ke.��6���H��?A�Κ7�M��O�@�
Q�O��]��!�%fz!YE�
��	�'�I�L����Iϟ����I]AD���ΠR�bD�w��U�p7�B=����O\�3�9O��oz޵Q�]$5�f�Qa�o��
!�T�D�IZ�)�ӛR3:1l��<Y�ϖ�L�̃�o8]~�����<�@ż:����h��\y�O�rM��NcD,h�/e���X�h�1D���'UB�'��I�M����<����?�d�;y
���/1�ؐ0�Hǚ��'���?������D����Q�l�&��J����'���ؒ�8�f����~2�'��U��]"��a�J�M�L%q	�'�bܑ��c ة�/�-��ڕ�'�|7�&JB��D�OF�l�p�ӼSlS#I�Р�[=wU�e��<���?���6� ڴ�����U�uC�?�"��;z4�	6B�w%|�I�Yy��� !�z��uc�2����{�X�D^��Nؑ�I�����s�' ��u@T�V3K���c���
	��\���	��X$�b>�CDΈ��aFU�dt�93�"la�0n�*��)_�e�'�'���;#�l��LP�tr���e,%��������{�!����ޫ9�W+�9Qb!�#'����	��M��r�>A��?ͻ�0���U��(pÉ�~Oz�"�+��Mc�O�=��JG���4��4�wU����.�#{�|�PlK2��,iu�'���'���'��'!"���Mx&ђ�'�̘��P�>�X�� ď�&���#�'	��'X6���Iw��O��� ��øvXЁ˒hʆC�$tr�lr�t�p*�Sv^�D�O��d�O�\�d#|�L��꟨�@�k�8�Ώ/�tiWi�]|h������%��)���?I�&jl�@V	U�#	be��BW�{V)67j�x���N�����S)������?��)�f�wM��
�F>'nnm�J�PjZ<x�'�66M�@�D�O��$S���i�|J���uC"Nאu�B�G�g(03LS���]��4������'��'a�S!�-x��9VǄ�9�L�$�'���'l���T�'�2S����4[i��C��ݒ'EV8�Sˎ�R�����<i���?�I>ͧ��D�O�� <.0)��͟�fL\u��K�O����H�d7�g��I.8\�Z��[@��'�(\ˀ�V7J��y��BǨ�ja��'N�	ʟh���(�I�����q�4�$! |	�`�(-�*��q�ʍ�7MMS���O<����ʧ�?!�Ӽ�v�\cH�� s@�;>EMU4�?1������O��Ol��԰fv(6mt�s#�H� �ȹCNY"�Rlg{���g�;��D+�$�<ͧ�?����ms���(Nc�x0�b���?����?I����[Ȧq�A���������*�Ä$��IZA��R�>ɉ�Wi�	՟��'R"�'_�֟p��b�G��m�5/��R�:)��4���Z�b������)�'I��,�(d�����\�c����o�0h�|I�cO �i���*�?�N�#M�;&�l@9G�D��� [�m�:|�,���J�E���(3,���)rf��/E��Hɱ^
CP��cj�)q�&,����o�u��� �.��ɲ���%Qʨ�Ї�S!8��,y��-S��3~�<���q����9���!d怨�䇳Q�*4n�8�88���<&���RB�|�YR$��_�L����)7�̊4g�SN�`Z�͛!���93 ȧ^_�����	�K#��R� mr�c���c,p�# �&]�Ā�E*b�ZQ���Ŧ��K�h[�}r�'�ɧ5����2�a�c�� ��l�e���d��771O��D�O��D�<eK�;.�h婵hՖ>RΘ��he�����x2�'JB�|"U���`(�/{�8��L!	w�K4��n��b�@��埄��Cy��
h��S�|����d�)
�i�i&Tꓥ?�������^-p�)� x���@7
4�課�ׯS�� P����ӟT��Dy�lҁ]���~=�g�K�3��]X�F����c��u��z�xy2`ә��'>tu���E]��[�l��&̫�4�?�����d��-�jT%>����?����B :]BcGS�Y���arN������0	-��L������ȯS�P�B/��{��npy"�Z�z	j6-Nh�d�'���&?)e���1[�`"��C6%��ɨ'�ئ��'2\����I'H��p��A�� �!�����fo�N��7��O
�$�O�)|�G�Lh��\54S�`�폪-���ҷi�:�ȗ�4�1O����: � %��&@ ���h��wDPm��������,���8�ē�?Y��~2�	6�,��	=b0Y��lX��'n�J�yB�'��'�p��)HD��"�X*W�`K�
b�0�D#j��'�t�����'���}��fb��j6���$0���x�@��<I��?A����L�_����J�o�=��[�>�PgL�Q��?�L>I.O> 9�͞�#�Up�K���!�����h�1O����O��D�<i����rH�i[�X��@�*_�i�0(��+�=!0��ڟL��f�Zy�����$�6���˕��HO�L��X�+����(�	��X�'qK��)�i��}@hC�r�~���_�P�6<n�\&�h�'*V���}rL�=���p%�����@B$̑�MS���?9���?��$���I�OF��q���E�v��YU�8Ã�5v�'z��''�Z����	�	�xR�l�&�.5r���Qr�&�'RCD�F���'��'=�$�'�Zc��j��50��	�%�VF�۴�?��0*a8!%w�S�'t4@�Kf��6�����Y*��-m�'?L�Iß4���\�ş0�Ir�do�7���/ �4��2Ӻ?�J�ξ�Gx����'?��Iū|-�l�rK���t�!��m����Oj�D]H$����i�O��	�Orݒ��E�(-�4)�!۝[$X-��d�T�Sǟ ���D��H�3)<P	���%���*6�ʀ�M�} �T��'�2�|Zc�\pEʶ���DH2C�C�OUe���O ���O�˓c��Ivd\�Uy�ř=~�p �& @� $��jy��'"�'���'���r�[�5�T�Ƞ*��ݺaK��4�bY���	ߟ,��ey� �*����<��Q��>?�XDPB��p|�7M�<����䓧?���5��1��'v��h��^sy�4�@�C6Q��O����O����<i%M��r�Sԟ�hQ.�)XѰ<����&�"@���Z��M;����?1�D�zd����	' O6%3�ӦE40�8��%r>6��O����<���]�S��S̟����?�-&I�0����xo*��6F�;��1$�P��� �-�Z����%�R �#E(R, n��憶�M�)O��Hc�O�=��Ο��I�?�ҭOk�3=v%���[�#�jI�6K��_S�v�'�2���O��>����q�0	�/)�|�3�i�p�Q�	����	�����?ڮO�˓mh��3��3\����
3(���x²i��<����/��ߟ|��/��G�l�u����vI��a�Ms���?9���(��Q�h�'���OѱB*@vfUp�/8�t��U�dF'Ux�O|���OB��
)Mͤ���O�.if,�Yq�>�ʴn�ԟ�s����<��������'G5X3�}��g���Yr%Ob}�b�7��'	��'�B]��'aP%v�aj��_��Ha`�Cauy�O8ʓ�?�K>���?�'��=a���!��Z�H@�W�f��bI>��?����D"aJ�'�ZY�GfN�~fJ��#�=��0�'qR�'B�	�����4�'�,D���E�yc��@���w����>���?����dϫdh��%>uqqb�8��LGG$7!4U{v-��M������4�z��?��_�~��P�b��(��p�U��+�M����?�)Ol��ӯ��S矸�s���'A�jT�k��DqcrU9uE�>�����O|�D%�9O�n~��([���h �p�7�&N$��_�,�G�C �M�ER?%���?��O�)H�iؤ ~�c�X$U� �iH��ӟ��I�ħ�����ES�����^�d�c�tӊ����I�L�I�?�ZN<ͧ.��x`&	�F4@��D-X&_��a�G�i~j�0�'��[�$?�f��q�O�q|�1��k�%!&�L鷹ib��'D���)��)�L���7��D���)LW�H����0��'|ƔP'0�ҟl��#Q��AH�Q�Qy�kדM\�m��h����ayB�~ڌb�@�{鮍�P��RE�&�G"B��(5�4g��H̓�?i.O��$�?�"9s΁69�ty���
w�]:�
�<��?a���'�����b�
}��A;n�\Dy@d�	Em	0�B��'!rP���	�E��'v�"q��n��x�"�FA�:�m���I��?��O2|'iBЦ��c�#�H�U��MP4:rJ&���Ojʓ�?9�j�,���O�T"�Xl$
���S	F4�!�ʦ�?���?A��0���'��Yv� 2`\�(y��<ID%Ђ�b�V���<A�8�B(�,�L���O���Ɩ(Óa�<n���j�
�,�n��%�x��'X�A�g�̑k�y��� r�HCݛg����i�=Nځ��i�剓!��tk�4b@��X�S���A�H�I[��P�Fu���7)�Y����k�ޟ4HI|M~n,u��� A?ͤyS����<6�Y�d�OD��O��	�<�O���T,�	�N��T��8k0$HZ�dcӸ�sd�k1O>5�ɶq@�i� ��*Z�����4f]�%�۴�?9���?A��pw�����'��d�9
�H3��;S�q�?_��F�'h�I�
�������O��d�OB(�1=b�9#���E�r�s$�ަ���*	|ց�I<ͧ�?O>�����'\v~xД�LmPD�'��e�"�'O�	��X��ǟ8�'>�(�m�}n2#U���*V��w�߲5O���On��<Y���?1`c^�	a"$�v+F�[���бK��G�����d�O����<���qF���a2��PBE�u�Y�Ug��M����?����'r 4�"��޴g��;T �T��T#���7��X'�T��Xy��'����V>��	�v�va��M�B,Y��M�ai-�MˊR�'X�ȍ�7M� I<鄬T77�a2)��_��"u+����Ο@�' ��A��+�i�O���Ƅ��e��� ק/���j��x�]��Z�c�럔$?9��]7"`��Z\杘�*�j���m@y�n߲U�6�X��'��D�/?�c�W�z+B�rTf E��Z�Hmoy��"5[�B*�	+��i(T�NӞd|b&8 ��CڴG�0hB��i�'�r�O@�O��-�����G�NQ^4��"[�sò�l�&;Z�A����`�'���y��'�Z�A��+iRLI� �
l��&e�6�D�O0�$�q5
�$��S���K1�# A��+ܮ���ʛdn�nП̗'�t�3c��~��?����?Q�$W��u"`ʅ�8����B�P�6����'\�Xs��6�4�8�D3����eY%��*�$FDҗ�v]�X� � ��x�'��'��Q���V��2�0�gh�O��XP�P�˝Y��͟��Ik�MyB�[�oe�0��eN0�a�F'�e1�T���'u�ݟ���ğЕ'lZ�[�n>-і�e"X��ᎠWw�9c��>9���?�K>1+OΡ����O�0`ǉ(y����GjPb9.�*��n}�'���'V剒3H�QK|b"jX���qT��6�r�"���w:���'��'��I�f��	^�����z]jXP�̕Q�Ù�\0��'SZ� �O_<��)�O�����[`���C��}�ǂ�=�H�HE}"�'���'����O�˓��TM&�Z {¨�v�}�%fU��M�+O��cW���Iݟ$�I�?���O�.M�CGJ!�o�i/<l9�ٟY��f�'���y�[���It�'j��P̭	��Dh"ϼ6��]nZ�By�Ȣݴ�?���?��'%��	^y��&K*8%C���-��?6�6-S���O ˓��O"�3u��y��,J��Q�働.��6M�O����O�8xօ�]}�\�h��]?���L,zJ����b��4�\ۦ���iyr�ߕ�yʟD�d�O���L�lv����bD�z�B9j�Tm��Fo�6��$�<	�����Ok�J�9�meA�R��h�0�١��If��Ɵ���ҟ��I�l�'34a�-�Iv�M��CS%�����-V&����D�Ojʓ�?y���?QU��%#,�+ �n����\�c�`�ϓ�?	���?)��?�-O�x��E�|��F� W�$�0!dR�uͦ9;�����'�\����ğ���	>�P�A'��!�E1\�"m��M[s���4�?����?����P*�fM�O�Zc�eP�U9bѐ����$��4�?�/O���Or�$D3�<}�<�LQ��E�n��S��ʋ�M���?a/O�@�f@�H�D�'�b�O�@�C\���X�"ġ]��t��a�>����?)��q������9O2�#^��ei�
��݀�@K��7M�<y2�B
=ٛ��'���'��$H�>��O�r�{F�W -KD�JVA'=~t]nΟ��I�G6����$4�ӵp�pr
��e� ��P��0�7��%fN4l������X��8����<�aY�S�EBY(/��3A`��Eʛ���/�y��''�	i�'�?��g��U@��B;I�})TՔw%�F�'@��'�(E�r��>A*O����������o%�7�
1����@�h�<���<����<�O�b�' ���R8t��%d��d��Q�F�'���a C�>Y-O2�d�<Q���$(�jTu�$�D)D�Z9"�g�v}+Ҭ�y��'z�'��'��I�"���/ƍNCXx{�֮B�d�ea���ĺ<�������Ot��O�lC��I6mF����Cf���3��+0t��O>���O����O�ʓF�~�y�:��}�gM�h9���C�����i��	ޟ�'��'y�b�(�y�	N�6:�B��lF��連`Nt6m�Oz���OR��<!B/UB ��џ�X�x� uQ�eYW�8���蔞Q�86��O�ʓ�?q���?�����<I,��nQ�P@`�ʎ19D,�Ĉ6�M3��?�)OB5°�]N�$�'��Ot ���G�w^�Q��~5�Q����>���?���lny���9O��Ӟ e~-�Q�W��Hk��]�Pt�6��<�T�G� �V�'lB�'�����>��n���ɐ.|Xt�@�Ep0��m�ԟ4��81����^��Kܧ9�v���ձ�.����K�Aa8\m��7���!޴�?����?��L���Wy2�O�����dYP�R�3�
h�6��c��d�O����O�Rh:� |�{Mݳ4�q �		���0q��i�"�'R�ߕ&֒ꓴ��O���5���t�ƍU���Ԏx��6m�<9��N\��S���'�R�'��`;Aߟ�����$�����f� ���>#�n��'��	񟐖'�Zc[Ԥ���{�-[�\�v�(��OZ��>Oh���O���O6��<I��<%�T�R�� Lq^��mt\N̓�Y�@�'�Z�D��П ��n���ɳ�d�f²E3�z�r�t� �'\R�''�P���c����TE^�>5�ȱ�J�/ ���@��"�M�)O��Ĥ<����?���`�~`̓}����9Ak������L}��'���'!�0=(V�詟R��J&n[x0��A�5����ܗ$�lZןė'�2�'\��[ �y^>7�Ғ���k��� /��#!�H�6o���'8�U�P��fI0����OJ���r�SS��=��Xc�/�"�Q[c)�[}��'`��'�Z{�'L�'Z�i9�hq�����<[����+(e��6W� P� _��M����?���J�[�֝=[2��)��l���V!?�7M�O:��ѡ'��$�O�ʓ��ONDՋ��B{�~	cBn˿j����4F�X�W�i�r�'E��O����Y<K2�`s ��e7�R�­P�`o�o$�	cy��'e��$�V�Hj�엘*0UrV�,��hoП��I某�!�V���'��O`��  �==�b�bqG�	���:�i�'�D��)�O|�D�O8�d�٪d ��/ng ���ƦA�I�K$ޑ�M<���?�M>�10�b1��)�I��I�%΂N
���'E2�k&�|B�'
��'p�I<Ay`�s�	I .�Ԙ�v%Z���!����'�2Q���	ß(���7��C�I�6��}�&.+�,�w"`���'���'��O�-�2
~>!�jR�e^�XS��ݳ&�̩�3H�>����?9O>���?�U��?I5i�;a���I%,@/鰙����d��	�@�	� �'阄��L=��ا!�f�	[8b'��21!�Y�w�ŦI��E��L�	�JUHu�I|��:*�!��D�"��*���3ܛV�'BT���r%/��'�?�'"�Ј�'���R�kB�( ��������Op���O|xR0O.�O��|��y�⍙i�x��D�X��@7��<1���$OǛF�~J��2C���q�E%:xHe��K�N
�k��rӜ�$�O�Y =OX�O|�>MX"���ڴZ���ᅔ(m77���-+�m���|��̟��S����?��oX��s�R9iuHS���S�m��t�]��h�Ix���?��)��8Y�%�̓R��a�b��Pk�f�'��'�����-��O"���xa�/��a���Z��m �L)��=A�\0'���������.��&���)��=���W>TfE��4�?�P̒�[p�'/"�'�ɧ5���K~8S��U�> 6)���D
���H1t�P���<���?����
3�&���g0F�yQ�:go��:C��m��?iO>1���?�UcQ*e�>yIS
ЂGd��$���n�B����d�O`�d�O���Zȡ;�La(�BU�hrR� d˺[v̙SZ�P�IП�&�T�	П���~��C�.ʔ��Cf@��*!�Yx�EN ����O����O �L��I�b��%�/l��$B%{Uv೔��2RT�7�?���D�O��'@r�i�֏!�E�#d�4gx��H޴�?y���䍥_9,9'>A���?�؇{0���@&��Դ�xfc��'g����a
���᠅�4�䠸"�i��I�����49��S�� ��$��k.hQa��LX�MJ$g�Cz�	Hyr�'��O�O֞X8��,hi
�$O8�l9�ݴ!�jqBR�i��'2�O�LO�I�!R�f�kT�Q�i�p���)^��'�����O$���ǜh:�L���K8r�]Ѷ�<7M�O����O���OR}�V�T�	[?qEF��L�ls���{�@1A3mЦ��Iҟ��I�&��)����?���q�f��p.X�&��2P%��X-��1��i��Z�������O���?��4R�9	aL��a4,�kb��u����'�6�ɚ'�B�'���'��s�l��j��:��4j�Z;��(qN�pQ�)��O�ʓ�?�.O����O ��>�8�C�ػ<n�c���!s 8O���?����'lA4s�<��Ȋ�܋����Ee�4"���C�iZ�I���'[��'�B��y��"�|M�W�֚8�b�{U@O�8qX��?����?�+O
��g�L���'�|mHd*�^�`�q�C�a�ȤQҠvӎ��<q��?1��7����?q��!�X��4��4r�͐�fڥgW�2�i���'��I4X���������O2����FAqC �F�N0	 �Z�:��'b�'�RF���yRP>�	b�#�ܲ9 �U�5\�a�i�ߦ��']~l�B�l�f���O
��򟘐էu'\-N��L;��S��}�C�'�M���?1����	eyB�'rq���(�YK��`h`���zr^��P�i�����Es�H���O8���Ne�'��/�`JU�ܪK`�����?t:޴td4Γ�?(O�?��	�T��i)�-
�(0��b 
P�4�$�Cݴ�?���?��狄��	fyB�'�DC6,r����^9q�blb�n	0R����'A�	*0�^�)���?i��,r6���**�P��̕0Aư���i�B��=
`�듾��O���?�1!80��b�
i�h�0gǌ�ZC�p�'� 4��'e��'b�'�B�'IBg)� ���K��	ކ����a��������Ĥ<������?��'�VX")%���vOw��t�ܴ~4���'"�'�R�?������|JQ��qv��t��n�ԓv���A��֟��I՟��?���~r�K�Qx؀a�k����'����$�OZ��Ob��O,P2�O����O���A W��kVcI �<��M�����u�I۟��'�Ƶ�N<���5u���s&iZ;�X�@զ=����H�I�$���K��T������I�?���O��'�k�l���@[��ē�?�)OF����i��j 
Z�X�b��� H4e�cj�B˓/f�ɕ�ih���?9�� ��ɞ�`4JvM�-]f�k�O'd�OQsG"$�I�?O4N����)ď��'�ƕ��i�H�p@�'���'�2�O�S�$l,e���:2�����;W�օ�6�fa�uGx����'��A��J�@C��`I�:%�����o�Z�D�O.���)�*��>a��~�� )��8��x�"����8��'��Mq�y�'�r�'� ���%J�1��G��0��sMeӠ�D�y7��>�����k��Nyʐ�)�
;E~�q�Q}b�:��'4b�'�[��iW�ȅ~�6l2wG�:�
��#�K�����O<	��?�O>���?����k!đb�HX:�4���U&��<���?����D9H���̧Q��9�
��WZP�gL�<h����?I����?A��\�'}Hm�0
�8>�ME�vi��ɫOD�$�On�D�<�G	̢��OZ"`S�eA�g��D
�,*Uf$K Kb�~��;�$�O|���O���Ձa'p�E^�G^�c��iR�'��	q|��J|2����e�#:��Z�&Mwj P�c�.��'���'������T?cg�؞(x�u`�o��UT"��� q�N˓W�h�%�i[맽?��'-���/2��"�M�������rk>7m�OR���2}�b?A8"%X"�d[��4^u��n��G$Ӧ!��ן ���?�xJ<Q��	�L=J2��L*X��	��Ai�q��iQ�!C���S�$��ЂK)�xA�O�"�MocD�M���?���yb���tV�x�'�"�O�����%s��"��S�v�ⲵi���'�����yʟt���O
���jQ�5��i�:�$��D�v d�oZ���2�LG+��D�<Q���d�OkL�v�.0&뗏<���g��':�	Ӡ���0�I����	H��'��ቇ*E.5㰘V���Ԋ��w�F�xPT꓎���O���?����?���S1��qP7hT*�JY�g�S	W�vU̓�?���?i���?/O�kE��|:F�_�T:%?��9c��0�n�}yb�'����������B`��k���>�B���d`���E��	�M���?)���?1)O
�1���r���5�b�"6�����J;<T $�M������O��d�O��X0O8�wD��{��L?B���"CK���ir�'��I�w �j��|���O���;pllm���3�4L`��X5MUD�'Q��'�R
��yB�'�ICJ���7"��$�6f�
P�bKզ��'
,�[��x����O��D��קu��"6
R]�	�({4������M[��?�%���<�M>��$�χG�H� �³l0�f�[��MkĈY)qc�V�'l�'E���>9+OH<��i60j�����0^�P���O�����f�L%� D�d������cF�)c}� 9уɒ2Д]@(:D�l��b����$�CF�>�X�� *$�OƄ�傊+ʈ�u�!���f��7Z�\ #p#��Q��i���ΡwT�C4J?�hy���l����=N��@��&��}�����N�T0��ѲZ:��� \x��5�Jif�Kd ��!5h` ��R'��p�ԸN������X
9��l˧��7f���)%kzEd�2��'���'�҅���'��i�@4��0`	�>Z:�m����Q�Q	U�mE�Q��.9j�$��h�N�'F�bH�(�4� �<����LT�
z�l���SIu�7-ժ3pACag�U>�#� �� r2�'�D��/$n��ʵE�A����I{�'@V�ӷ/�}��D05�Q+Z�x��'�����#D��G�	K�m��'�V꓾򤊆8����'#�R>]�t���:���Va��&ű&a׍H@�Iڟ��IC}�y��E�	�1�G��?�Od��i�Î�$��ɚ��۷HF�\i���v	h�� �Hy�v&7�i�����M� ����S�Er,�GyR�Һ�?�����O��!rw�P��)�hq:"(��<!	�_�zHb��jlxC�P�1�rx���-�ēJq��q��#N�d�!�ܪb��H���W���Ip�D��3&��'��-$�xS�]8F�� /7ɒl�a�,5~,A���	h}*�"b>��
4��9�@��<M�Lœ�(��[� ��HV�=��T҅�ا����O���T�� 8�0 2��.l\�Mh�dٽOU��D�OL�S�D�	),�AC��� �#YIY� B
�'���s�	Y4"�\M u.X3+��0���HO���cAX���J�s���BJ#S;�����(��D�@פ���@�����[w�r�'�h�8�oXP����A��?�Q��'� �	�	&>�d���\M8��   ��A�"x�X�$׾*�H�f �*�@�r�C�6h�92cD�9U���=W�.��L�v�
���.����	-{�ԁ��ޟ���t�'i"Z�H�vMZ��&Ee�;�4Z�":O��=��(�'%��P�]])�9`G�"��&�'^ɧ�)$�I�`�iSi��u�8� �92�tC�	�GJh�r�g��1OjRsGQ7zB�I�b�`u�#��[m4�Ȇo�+�C�	��|��	� V�N;V��^�B��6�-P����a�2�j#UqpB�	H>FU8�3��&L��HB�ɬY{��
qNZ�$��A���c�C�ɘ_����"�?U���e��9BʄC䉳^������K�ѫ��XkbtC䉝#Ę��vU�:�b\yl"!6LC�I�EOz�1����:�L�Y��a>C�I�ua�p��7G�h P!H2݅>D�`Q���J�A��K+�6@��&D��ɗ��
�&L�0��>  ر�*O�a(�M<*�v	��
���B"O���p+��2�q�D�_�m�� �"O�����O"
eniA@���xp�"O�I;�a�+y��z����$@c"O��s��ʕ$X �����d �iɡ"ON���i
7-f��:%�4J�$	�s"O�e�%.��A�b��K�`�B��"O�͋��L�,�r�	
T2%���"O��H�[�C��يQh	y�ui�"OX��8]��	6�KEp��"O��'�з?`�k7�	2[��h 
�'��U")�5�.�;s�ռ{1���'{.9CĄF�w�hA�]8�<,h�'�M����q�d� )C4L�N\K�'���l�%�j �[�n{��	�'펬�G�z��@g�d��`��'��p����=3��< ��C&Eq�y��'�(q�%(�N��X��r�����'/J�J�	<+^&!��E,R�|���'�QP�N$&Q0`0�n�45�L�h�'9@��gJ&\��d��Dۆ;��1�'��#&	��<�0D�S��:SV1��'��h����Jj��2C�,�D��'�<�[4߇���s��W$��`	�'�z��pM��+�rI��MY��>m��'����Ά�m5�S��3xԀ�'�A� ���h���"�@�'�F�2b 8W�<5�Q*����'���&F�akb0BΝ��y��'��[G!R�>�1�*�
q��I��'7,4{�G�
G��*)�#�LJ�<9
U�|hN�9��	*� ���+�|�<�U��T��������]���Sz�<�����w��P�ӥ3�-q���y�<ɣ��2�1��	��֥Rv�<Q6��4����TUNk�1x�ct�<��M'>o4Ș3%ڕb1����+@q�<	'F	�`^`	� �D��*Q�j�<��#ȏZ�F�wgA�dFDKg�<�g�I,IjY#�n >�� ǈ�W�<q���\o�� ��F,ܽ����U�<����%x�*�q��`�h�k�<iF��3k�9;B��B�`Kt �e�<����{e�x�wIL�C$����ώe�<!��ƳH8�i# 7���
��NH�<	˞�Yɰ�0���i9:�0L�G�<� �����

ufpS�ȡ	j=�!"O��{2,O*h��q����3�l|��"O:��
��Ox��!R� �v<rQ�"OҐ�B� ю�"D$��v�$�"O�h[A�ԥ*�FQ�Q�_�I
���"O��IU�@�#�f��V:-�p-
�"OH�(��{�H{0A�Ɍ���"O���"D89v�	8�j�	���R�"Op�ЅbZ6k9�+���������
Y �E��i�d8|�2�#V��%��`���y��E�
����T@L���(�5�~�憤�D�=E��oY�{��I���>Z`y����yH�$�Qiȶ>�.�Ȅ���ɒiu�}��'�4�� ��@RC��D@5x�TU���
>g{d�	bH!:*xкTI����B䉆D^������`Jv�׽&i�"?arJ��#n>��&OȊHW�`H2���5Q�+.D�����ۚ@�\�R��J� ~<��uf,D�h�C�G�T�����FhP�d7D�h��N�/�lS�c�=�J�Q�,1D�(�J��N��a1�UH��{�%<D���F�:�Bd��a?E���ps�4D�t�g��1E�:ใ,.HB�Q
��.D� J�:M�2؉5B�.v�tI8b��O؁���)�'r`}�&��*$d�yZ U�OH��a���$A�x�(�
Q��8aZ�Q�J9[�h����?I�	�/�|���*޵��O��S&e�8u�Z
���i �:EM�`�6�G�D�t)�y�M�d�kL�`q<��P@�Q��l c��77>�K��C]�V-2��N���z�M���Ѵ�6\�u��D|�=qdĆ+v�(���MWh��Ua!�_!����0�Y(K� DJ���T�7aϱT�\a�*,�2�)�Ջb6\��?,��)j��'�L�h�iҷ{5�������:�?���Q0~�P �2kF�QB�ER�jދ@%�'��d�$�Ծ��Ϙ'k��פl�"L�6��j��N��<��+�(k�3d�V����d�4'��;Ì�'aq����Z�a�$�e�[�7�H\R��'�4��a�K�wD�Ay����K:r\��b��e�P��b�7��ٸ�򄝏2b|�qb��a��I����2�NQ/,R�fK��fV�=�)�##̡QЃ�TE�ؤ�����&�;M,8�@��[6��x0���<�7l7�Tp��@ ���2�Է[�h<�E�' ��@�� n�H|����3D�?!���W�q�8��Q?5LH���l��'b�(А
 �Ϙ'�D�iV����3�K�d����F)���y���;7?T�I�@N�*�3�I*Um����	ʕ=��`Y��Dd\L|��@���|��,<O\\�a�P�M�}�cF�>�1:��C0ML,H�A�P�f�w�I�z��zA�B2ID<�j�����?TVR��ʎ�I���G{��)g�~9j���T����O?�V언�p��Ӽ��U�C!=?1�l�}0딇Cx>PT�ۦ\h�c�&D����pf��O�M�e�Ff�B�IbI+'�|����&?�����|3��� ���y"���J��u �ڼ�@(���	$bx�	}���*J�8t�N!��(OBP�+DD��B�L��h#��ˆ�'+����(� E?�Y���xA��Z&s�@BF�G�t�X��'n*�H��͚N1p< �#�
n�����$��$�er��C,\�q��ɰ'�ӉSE:L���N�\q�"O��EI�Qu]�#�-3���x%�'��]P����Z�r�0�O?QR0�K�I�X�x���Re`�*�
�V�<	���%9�XRmV�w��貣-_Qy�AI�]%޸�Þ��p<q� `�=��m
�q��E�4<a~�A��P�_��p�ƃT�`�"�HR��5�4� ����*��r�ra��R&j6��	A,�ѓ�� 24����FK)�����F!���e��a�1�X!/����U��������
\i�ᓡH�Й�NG4u3�/@sȖB��1')��`���5DΐU��,�6�tb�T��$�Ye�x����G��,1�#�+6XhB��U��x�薔�����F��}4�$(!(� H�*�e�I(<��@IAA����o�ڳ��B��'�'�qO� f�E^�
�(q�r� 1zn�%R�"O6$#Viś��e�c(��֙�<*Ð7h�qO>�3g엏S�n�q��.|��0��,/D�tiA/�V�Q��`�l�\�#.�	�,q\��'j������ +��R���Ѻ
�'ꢰ���^�J�@��S搨�(�+!��S
OV0����}(D�����{���!c
x)�ՏR��OA�9HAl�\b��J'��	�',5�t���ORV���N�
��A��i�NPE�8}r��Z�O��)���q����'�?u7�a�M�2��OD9`�a�`����A�Ih��g��hǯ�>q���X�'e���,b4p�$l��m�d�q��A�Y.>I�!�E�}済 *��k�X׌#K��%qm�#b�"��Va�=y����-sp��'
@^IhJģj�Y�4�
�p�셔��<{����m�p�'�y�)�3n�lT��#�3GӲ�1��y�1�
A��#4���R��v��x磈 4ʨ1�Bg��L�
�i�O��SB��7z�d�'%N`�1����вgL�B�lC�rE��� ��;��=뇪M@:�Ի���!�x�����hZ��Z�{�,�f��X�,J�k�&s�
��q%��Q̤X�l7�{��3J�E�ջ�U�h�R-`�cA�kĥXҍ@4?nT�W�a\8)�"O*���j�K�*��������ҽmV����[Kj�9���*\*6��<��>�.�/CȨ���� �����L)az�'���dL+er��r��I�N�z�cuj�@5� �ͱ[�9��_)v�^��]h�Z��4���`sㅏyВO.�I��Dy�����
]������ڲ֢�H~��i�1�j�Ӄ��:��J��K
?�zqZ�ψ�C�]��
(�8��E��E{�Ii5��%QY���ψB��\�aP�`�d�AT�V��hkʧN%IF�Ob�1�d]8���s�$Q:rJ��"N#V5�1m�-�f��,�11�r�� HRd{f���X�gj~�@�A��(��d� ۰
&F� 5�P�A�C^v��C� ��	SE]�p���8�m�8@[�"N0�9�D���
�n8)`u�#h���L��'+�t��6��UK�~�1A<I;P1����e� B�e�5Y�����Gc��hYD4�X�')��Q2������-��} �Iώ;�5Ä��w�"E�R�����O �k�)+�R�N4ɒIS�Fu�P���ABÏ(r~�ŊqgL'j���B�8d��� ��'`����N�49 �ղJ�zE�FA�Y����$M�1 ZL�t�W�d������).Z48��ĐWjeK��Yn��ªʧQjd .T�QЀ���'/@C��S�qT(G��'^Mn �wB`�H�K���j���8�``�R���V����݀FbF�	��C(W�a�pN�>7~,C��
U�%IhQu�ʑ)CK�,>��SQ�K�t��S��V|��ǀQ�	�hA<(Z��<i挤:(��+˭N%�(�/�~x��B+ʯJ-�Ӑ#��2��i�p���w�<��B�/x�� ��/J�9�G�1#���R����!L֘�:�C3	 � �<��b9�	���ܴV=��ZS�P%`6!�'!��.c���`��#�*��*�U`.C�	�:ˮI�T�ת��N�6t� C�I-Vi`���~�Ybť_�R�C䉗@����hۨ)��8��"ڕ7�C��'*���3�_m��)ɇ�
#�C�	�q�8��\�y��MӲ
#J*�C�	J��l� ��-M��r�!Kg�C�"���׌W긨{7��$[o�C�(0�p-�Q쏿��HfDѩ%~C�	3��|����'.����b��5�C�I�WxrM�s��=n�6�����8y�>B�	�6�h���<�R���-Z/�B䉟M�����1|(�d�h�C�ɣ1T�(�i��L L�P0�Ӷ��C�ɄQ
J!z��O@�§��?�B������+s��� ��*^*C䉢8Gh�(B�
�NB�Do"(�X��zLD-;ɇ�f�y��q%�=�ȓO���W�X/1F"�0f�\��DՇȓz-ā��U����M%I΄�ȓ�0;�͟7&ʝ�g��z���:9�H��^�=?�1���P�a<�<��9�%1�-%wrBU�ӮB<O~����N��@��鏬#la�[h���̑@�<� n��Pu֩�5���E)%
e"O��������Ԥ�)@��C0"O�,�C59|�6��e�p%��"O4B�D4Co�œ�!�E�pŃ�"O"��3Μ�V ���/�{ 4ɠB"O�Ȣ�˩Qcb�X�#	1r�0�"O����/ ]����$�ψtR �c3"O������Rڨ���K�	C(��"Ox@Y7c5rJ(Y�VN�<r$� d"O�)���$R�����X8C����"O� pɎ+e	M�eYE`IS�"Od�:wꋁ-R%z 瞣?&�Щ"O!s��*g�"d@G�¢-"�( `"OV�8�HL!�j��6K
�Q�@2�"OX�"�aP�~,f��v	U����Q�"O`���	��pF��5�2î�h�"O�� ��צIVh)E)�
{�$�S"O@��"
ؠ	SL���%D�(��ɰ"Oj�����<�u�E�X��\�s0"O�K[�9��kY=3���6!�C_����`U�q�Fia�*Xu!� � ؎h���8A�������!򤑲qȆ�Q�A��"o�.I�!��٫6~����84�`.P5Y�!��їx���0)C/��Yyƍղf�!��=4Ӳ����+5��m1�,կdS!�ď�SSi�+�J%Ae��"?!�D��+%X�mͯZ4� fY6�!�D�,p|��k�+�(vˈ�+���4�!��<.@�Fm�P����r��fm!��M�!_����/-5��]���#Xb!�� '��p�����qk1�B� `!�d�6�r�FN�;sh�]!�D�%/�`��6��C��u�&��G�!�dL�+e�T��?J�� &A�k�!������cA � |�л�ŻGT!�$�#!��B�W�Byr�&��6N!�$GJ<��֢ėI��qD���_!�$�c��%qr`�!P6�,HV#
 G!�D@�yr��� N4g|q,�;>!�D�K܆��LV�/f8�MM# !�dԵ��p��.��XL�FA\�!�D��i�ٛ�$�)W�\b�\;V�!�dϻ �� 
6�N��8ɔ̜<p�!�dj����d�>H��\8憰An!�����%�UD��2���H�#"7�!򤑕&J	�֎��.t2ܐPI�#!�� Ű���UT��)�g�^�!�d����EPQ
�HRr��s�Rb�!�ГY�ݢ�'�l= <�ׯQ/@
!�� �,7�� &kѐ+=�󮀥y�!�$ԲR϶��엇{�8�% �CB!�d1�0E����i�x����:1!�$�{M��·"�?���a��/5/!��	�fa¤X��b�X�0)!��,����cȚ5�NLJFcgIc�'����p�|��&�^��ԑ�'� ���Y�p��FT-]��s�'�D����6P\P|�oŅO�  q�'���e(4��tī��IN��
�',e���X%���*�tR6Hr�'* �I#����oЃ?�<H2�'�Ƶ*6�T�G���^q���D�6D���u�ٶwg�1���2"z�Ѹ`�3D�� r������Sg*
�o��B�"Oģp���(
�b�n�s�4�(�"Orl@C�^�K-R3�䟴jʲ��"O�5h�'���ٲ��.㎜�R"OH-1��0_�X� �w��%;�"O|h�bN�$/�IG�W�W�j0"O:�A��Φ4�n�Y��O	1¡��"O�e��W=�Z�cw��6Q���J�"O����
�+F,XP�E��A�P`0"OVX�7.�*���*�(J\��u@�"OJ� ƯG�G?��D�t�9r3�
w�<iP�K�r���K�,ph���p�<�&�Pj\�l�S��c,�l�<�Ue�7g�je���C.r�y1`�c�<�bj�e,�`���N�=���H�Ʌbh<��kY�my�$ݰX�(��G��;�y�N�p�Tm�Ï�!S�&`�����yrd�D���H���@��3U��y�#_�pԜ��A��3�XM:�)���y��U9�.�#� H�����y"�ݱn(�Ϳb�>P{����yb���0��d�F���Y掔`�G�y���'1�� tIA�U�-X+��y`�m���
ef�8G��:ŉ"�y®X$9����ǍגKy0�������y��آ���`�W�B�V@*��]��yK�d��s�!ـfRx�����yr��Cw: �P�+r� ����y�o׾k���
��P)q�ļ[�M֑�y�^5;���r�N�b�T���ʔ �y�H���Ȝ���R%e�~D����yr�����D��7^[< ���S��y2L��
�+�>cɒ���^�y���G+P\�B��6+��A����y2 \�gn�E ࣓>*i܄�3EU��y���z�!d�6 ��pK���3�y�i�$����m��d�H-9!�8�y¬�3[���E;_Ρ0R�>�yR�6x���1�^U�<������y���&J�}�U�[,a�BA� T%�y�i߷;��`�-�}�Z��ͅ�Ps�%2k_�<��X)���|N���=�bT[�h)m���k4E��=��@-���Od�а�!mE�pH�ȓ\z��س��#���Hd�F�]�n��ȓ �jp���;JҪ����n���R��驢"J#Dm\Ѫl ^���ȓ!0Ty��R&�<���� lꡇȓ� �/�Sղ��aK�!�`�<)ŌCM)�<"��Yݴ�9#k�[�<�ƢNh.MC$�^,U[�H3�Wb�<yu�]�8HpTNB+- (�Z�W[�<�M݇X���r����s�8�
�*�P�<9��H���vO�J�q�	�I�<�s�K���@�K¬|"9� �M�<���%u�s����#�U�y�J�Vք��O[�A0�`�M�-�y���!F~�)#N�*=�Qr�n�y�K9{T
�b��O/"מ�6�J��yR"��F���a`hÍ)���%ۍ�y­;��Y�AG�x,�ٛ���y���]֪p��Y1XH' )�yM�<U	�#uJ�0M~�̀7�D��y�(7+������M�P窚�y
� �)���a�N83shQ�kܖ�c"O�y	3M٨9F��2H^�����"OxȊ��.�P���ݮ_ʰq[u"O�����E;�~��6�1`Ĳ�`"O <)��πa�p��!��o���#E"O�2Ǉ�gO��v
Jm1 �c�"OHɘtJE.% j���"K�|����"Op�R f�;S
�E:bб(��<��"O�xgP�7CJYA��ӄ>���hb"Oh\A�.V0{�E��${�}�u"O~9��(d�Тv!�U\ }8�"O�p�&��bS��4JR$O�xQ)f"O���#^-5�����<A��)�"O����55�������O>� �4"O�؄��[�
�D�ӟ.�E�"OZ��a�S���Bɛ�E9F	�S"O�`�
�?��[�"�-ú9�"Oz�ɇ16��u+�!i��}��"O��@oJi���%I�+8K&"O��P�I��8�$Jt�\�H�u��"OA��a��;ndx��L�{�v���"O���S�ߴA�ɢ�B (���"O�,:��׫-0���� �bw0�h�"O����#ߤW�h���\�Sp�1�"O��X�'��,����@��(n�q9�"O��G��
,P������sg�ظ3�'Mў��L��m�u�W�f0f�h��1D���0�&2DI3(�_�\PRa.򓞨��i���GR���$x%�B"OtӁl��zp���R����"O�p�)Y0 ���9)B��`"ON�
e�In���Y��ݥ3�HT��"O\�Xq`�. lh$�(T:/$��{p"O6�9���BN,�9�撾><�}X�"O���D��([����@%N\u*"O�2�D�)*9f�Z+Ysٰ�Ґ"O�����	}(`��u��r�Z6"O���"��'f*�#��_�{�굑"O��F��f�`-�X�4rp�ط�Ii�O�����
]j��ꢇ�5�$h��Ğ$S�ƞ%/猙���	?�]��!�"�i��
$#�H h�'9n����e��| [" j���1��
v�ن�D���e"�8rI��c/�L���Z'��z��ڈ>P:�j�j 9\l؇��8e�ТO4n|�������pϘ��ȓY�˥�L��z�	9pt�T�ȓl*����
�U7p}
%�� �4ч�H�@�`��2��9
��ExHԅ�l�f Wc�cd�E׊X�����]�>�X��
:�͒��M�D0�ȓPC�ԛ�cnX��D�99��ȓ%00�VO!w8E���+�+<D��;�+�*^��SC�}R Y��	3D��PD0�����(�+x� ���+$D��6
r�1��
N�Y4�6D�ؚQ�0Ȱ����3\rQЅ@4D��̚V�|5ْc�]\���'�1D�a�
�n���k"��+����0D��z0Z�6t�U{�bب 񆕱�3D���gH6�
��Ժ �'@0D�<��썄~~�X��CV~|��WD+D�$�R�
Aɮ�R�k�J�%D�Li4�	�X�R\�'�v��h�%D�� �,�����p��걧��}]f�K�"O�嬘`E	0�GY�H?���"Oh��Q�,5�����kO/��ҧ"O�l�a�I�2�d*1kԨ-���"OL|1T�ss�X��D-f����"O�3"eİ;����d��R�Ƶ�"O���5.؈��Z䌈ie$�A�"ORi�$Oے'İ�a�D�L�ʐ8�"O(L�Ś�%o�p���K.>��cG"O�)˕��kQ^�*�L�"��r@"O�̑fe����bs�@��L3�"OTI���<[N��a�CV& �F,�"O:y�Woݔ%��c����q)V"O8��nT�}�t{��_��"O�Jч'}�ƁK��#/��x��"O�����Z;d���Ϋg�1�!"ON�$	�C=�,���ϖ�a
"O��7e��61ްA��k�B�KC"Ov��� �̥K�H΂���!4"O�<��"��4ކ5.)c��=k "O�@�H�E�L���M� 9�fD"Oz-�� ]ar9�D̀)s�Ib�"O�����L.���!�����
F"Oʁ�#�L�
��)�	֍<�xm�!"O��B��̛Y�<D���D�H� �"O2)ЗIBZ������Ŕf�$��"O\aa�Gk���-�4Xޤbt"O�<(֫�	q(�%8�-� U�-J�"On<P�f�,H�jË.##�1i"O��',޴k�Dm�C��1�$�"O�MZ !��|<�PIE#e��*5"O��(`�?z4�d12jX%Q���"O>uY0�$�%p4ϝ�-�f�Q�"O-[��_;Y�dC%[- ���c�"O p9Q�Ft�]:7��Wmbt��"O�"��pt�x�����P8�H�"O�y�@ �0rTcֈ=Ldٔ"O̴�f�	,>��6�^���@��"O.�X�^u��P���*�(ti"O�X����)5Vd�q��t��X"O�9��ar�iGaV�f�z5�a"O(y��K}@��"cR{� ��"O6�ر��?+��k���;�B�X�"O����Z�/��)"��|�2H�C"OR��͇Nv��@J�|(d�"O.pq�����\-����Xf�i	S"O����)�(�T�`%
�]�U9u"O}Q0@�Hn9��@�<�N�YS"O��B���yE�+��(F�X0"O.�+�jD)x)oC>�X`+�"O,	�B�֧z�d K�Η�f��W"Ol@�����B��0��K�	�Pq"Oఠ��\$ � �k�r��"Oe�� �<K��y�b�E�-슸�2"O�QI��B�;�h��OP�K�,"�"Oحj4!L�O�����('�ْe"O����*Ю%K�gF<�ơZ�"O�	����i.H������z�ٖ"O�ʃJ��y �h��ڇ5-���#"Oz��ժ�y�8���2$�x��"Ox�H��A�?���y��Z0Z �P�"O�t�B&+T����Z���[�"OҨ+"��p���t)��J�"O���`h��W>��8AM��r$��"O� rP����\�Z�̃Y����%"O�m{4�Q�T|����^��i�e"OV���(�B�"i"W�ħ �~��"O�MJ�g�[ZQ���^Gb��"O"�acDۭY4�Q�+��vc��JF"O��ǆω^��B5@��GI��"Oh��E�LS�-��^$ �����"Odِ�M��+�8��6#ǽ]*����"Oک��N��Z�(�"3%�8"O|�شO[r��ٹW�Еd��[�"O�R֧B'D���d��ȸ"O~lb�G8X��!b@�0�.)`�"O�`ؕN۫Z���X� �~�n,xa"O���C'L��ɣe��\���"O�Œ,
"��Q�� ,�B�
�"OrpK�AC�&*ze1��W�~�PtR�"O���R㏡���C0$�+]@��""O���,	�*�PQש0d@PB�"Oh�S*�U�,�R�K�ifzx��"Or8���O1%�(�Y��	F_|��P"O
M��M��X�X�CG��#NF��"O����U�I�(���%N\��"O̪f�Z�su*�8ÃϡonL� "O�Y�A�	9Z8T�#��S��-{1"O� �nM2jW`�"�
q�#v"O$�5�[2w�%�k����Z�"O
٠�[9�JT9�oW�J�J��"O(��W��8�d����)O�~SQ"O���"Σ>�=����#��09r"O`Ȩ�eE0\�PE�����F"O�-��+ �.¸��c��E���:"O���	C�2����l��aq��b"OT�ʓ�
�Q:M��L�	"�"O:��������C�MԾ/�2��s"O�LJ�NW-#� �r�G&���97"O 鲨��m��ܸ��?:v�$��"Oa���Ѱ[�f`8�Na�K�"Of�3g.�?�����N�L��E"O�!�,��������9h1P"O4�Q�ǯyζ�s�iԕn�j��"O�u!1nN;����ȕ�L�u�G"Ot�Pd\�^�8���':~2�ݑq"O:E�B�uӂ�c	&��إ"O*�X��\^�D �͖.e���"O�d�����_�L�@����w+n,�"Ob��5�Җ����7޸0'�=:!"O8jC$I��8�ɛ�N�~��U"O��"W�Z<X��H7%�^)��"O�|�B&�Iֽ@d'�5��`#�"O6<���ڀ�^�a�TtB`��"O�Hh��6��Q ��tiF 9�"O@�B�Ȁ+8�A��Ҽ{Z��ye"O�T�Sg�?)�6�#�#����[�"OjD:c��W���%$O͖�ڥ"OJ+���e�4,)&D�(C(4��"O�Yh"f�R�f��䘟(��"O��{�L��*V��b�ħ�R�23"O̡3!�ُB�2]0s�]Fn��u"O�PgHA6F����',F�E�u"O�e�7�q���b� C%Uj�!g"O�Pb`�I?I�t�0��7QlHI��"O�����ڷ1x�!E�BR<̻�"O��d�_�k�<m�'��/?*��c"O����P\ެX�"_�Y6B}(�"O� 6�g�qRD����+��@"Onř���Xˡ/�K�8��"O���b��e�~�A"�
�K ��7"O���?/�9b�N�P1�p��'d%����r���Z�k0}�JH��'v��Qږ&�T ;󊛭g��'>"926oR�M�z�s�ꈵ_錥��'N�q�~ �|cC�PM,����'�`x8��7G�h��HN%He��r���hO?��O2u�T�R��W��9EOQw�<�r+� 0W�����\�:�<Z�e�G�<� +�(@��A��ȊE�D� w/�A�<��c���܋C��8N��Bb�z�<�@[�J��I%��D���"�x�<QR�P=	Ԑ�^+�z��B!�uy2�'����S�L1O���if�)G��}��"O`-�� ւC�h	����|��	ZT"O��C����r�)Ң� w���a"Ot��rd��)O$8���X��Tȡ"Op�c�ܠI&����T ��Xp�'�1O�̋��P:Uz�Yo1R�d�S$"O�d�'I�2|m��M�,N�D:%�'�!��r��
��$P��,�b�0&�!�1ajxc��Ǐf�jp1�K�w<!�DM*�r����t�<��@��M�!�DM�S�u�3�J�0` ����p�!�d �2y�d�-2L�������!�$Ԗ��8jB�Ⱦ?�ၥ�@�-��d��Vvd+b��7�M�����B��>v} ��Μi�~=;v�V�B�I:I88�M�g�|ي�eE�l��C�I�p�Z����<�*���cC�S�C�	 &��u���� Q�`�SI M@�B�I8 �p!a4���)��B����)�hC�x��(�z਱�E/˒ՄȓhJ4��J&�2t�F�(RBj���U��bM�*?����#c��Є�w_ �1b��:Yߊ �&��~V*0��A�����L��\����Kך'��(�ȓ	�0��N�-<wn�*��@���ȓ-��0� �05E��ʕ�^�=��p�ȓnC��L��Y`�?s)V0�ȓ7, �VA�*p�<ȕ�4_����	Z�'�lpkDU|l��f�*^��x�'[�ق�%��;�-3$V���Z�'��v�_'ikm!/��K��Ah�'�xd٣��*R�R�r�엪B� ��
�'�&<��m�C0���%��<�
�'J�-���!��`c�R�4�������*�'3�0�� '.B�@����ρE삭�ȓ1"�}�#�G�tDXqgB6g�Y�ȓE�"剧lE�Xt����Gb,ф�*�Vx(7C011��`���SYR��ȓB%D��BkU����4��`��eDLʔ.���j9��հ,��(��
@T�� ��ac̏4&��G�'>M��
 C]ȱyP�CU�� �:D���S/�z{HXrD�7mh�X�D&D�x6��`�N� �e��[K�%��e!D�t�H��#)I)ΑZ(���*D��Pd#�7Aa0����R� r�i3T���T͂�s�4]x�EO�sN�T9�"O�Ѣf��g���c�D:j����'�1O���܈d|�!�`�ua ��"O� �<��i��@ zQ-G;[����"OֵS�Ŗa��c��Z�8�2� "O��j�@�n���8�"WO�U�"OP�����6��ձ"���� g"O�����ȴ4s�;��D�C���"OA�ᝧ/�4�P`)��3""OTPٰȈ�4"NY�g�w{D1�"O��0�Z-[U�����"�0�"O*��R�9�rݫ��̊[�ċ�"O��{�r��r��[Mt���"O$�	R��J*b�� LV�#Ր��7"O����=FFp��=1N�B`"Oԉ0 �K*`����Q�CH���1��0LOԄȳ�^,�R胶�ğczT��`"O��X�@�~��9:��3�ؔ��"On0�
˜�:�Q�I�0'��% �"OL9�#(��l�ڝ��g�fY2�"O��ī��t% `�V�5�Ա��"O���W���)�!{��ĉjaT�a�"OT��t������U)�E��$?LOxY��S|�he��gFޑ+Q�'7!����#Z��Α>��y5"[�!�d�=B
8�qҏպ|���S���<�!�d���<��&ô0>Yk ��O�!��Ŀ��]� �΍ZZ֬�1��!�D�~�4���$B���w-u�!�\�XV��P�ʹ9)R%��.BS��'2�'[�	O�'��$���J���x��P�x(����h��ə"�xy	�ͭK���т�TC�I#����ɀ,u���%G�\JrB�I�>1���t�
�&h����
@�B�	%x����L-�&`j��^'�B�ɥj	��Y�PF�Ɇ�xLC�I�]�4��c	�I�`� �X�e4t�=�-Ox�?9�$ˋ�vD����[&|:��j���U�<I�L���HX�/���%�>m�nB�ɢV|����c�m(IL��C�I)o��jl�-���D
{��C䉋A�f��2�F9��p����C���1{é��=z��q2'��W��C�I"f�i�Cg�g��ٓG�60Z�O�d�OJ���O�#|��eL6"�0�l�_� ���_f�<��ٔ8�Q�4m�Z��KP�Ni�<��&O$a�ƹhdZ�?�����bK�<�WJ�{c������}&p�b�}�<Y�g�2ev%�rAS�0����|�<�c��YH����ק1g���	�|�<)c��V�UGS�{|���@T�x���O�bH����/��(��.
3����	�'>>�&J��z�脪Sg: K�k	�'�fU��+|CjXP 	eߦ1|B�	�v����Ԯwm���q �#l�C䉒|��k�ȍl�ذ󃟒��C�+[Έ���R<v����%K_�(��/�S�Og����a�m1z`�3�#B��Xqg"O̭҂W��L��c�B{j�2q"O��y$(���=�d�^(@^2�Z�V�F{��)C�r�����-�`E���ً@�!��òb���R��Hp%F J�O���!�D�ZY>hY�hא<��B<��'$a|"�DP�
)(F.�	\BP����'�ў`�'���R B�zZj #wO	Y��l��'K�h�҉�(�����bD"N�؝#�'�h(&��b:%�Ə��E������� �s�?>�����̄����e"O,uIE#������ۉA����"Oġ�Gm�! QQ�?GId��c"O�U��>?�TY���*�"hkq�d1�	ߟ��'�PaC���O,��a�h�Dl�
�'�x|�L�$�&)��ā�zm�u��'�|aSG��S����a�1<���[*O8���O���VA�uRL���yI�?�!�DE�{�4�t�Y�;|w(Ɋ�!�䎲i}�T ���2D)r	�+/>!�� o���Ȋ�����~�!�X����CpZ�5�$��X"D�!��ob�=Q�	|���6J�!�$��qr$�A`*5�ej/A�!�Ε*	��hç��,�̡�4��V!�$ۤ|�J}�3(�:y�=B�ه^!�ĎѨ�,Vm�.�"�11�O��d-���r��fz8� g 5�H���'�ўb>�'׸�R�)
:���L��h'(
�'�\u�1+Ģ;@��OY�Z����\�,%�T�'�9C�䎛i�b��q��
P��4"Ofx�HJ���A���ഴh&"OP�1��-cd��p�],��Ђ�"O��;�%I�)>h)6jE4d��@*s"O6p�3��+�b}T/�gs��3GOz�a��N�XA���^�S���9�	=D���Wk�Kv�L�h[/ ���9��hO��I;R�k��ūn�b:1� d�C�_rn����"F�z9�EfK0^�C�I���]��m��6��M��'��R ~C�?>��eB�ѰjS��	3�'C�ɒ&dR܊3o@1Q�����C�n���O������;$����q@)3�윰k�!��cy��A�-�5�)��*]��!�d�Pt����$Uz!rA��¸R�!�dۮ[p2%dB���x�� �!�ɧ<�$u���	6X4&+@0{!��V'!E�)�A��7c4�	��J J!��5/�;�c�� %xA��O��Y6!���!QVp���<����K'!�$؞jE~�q�ʷs3 ���C�n!�Ͻ-+�\�Bc�{��`��y�!��]%@��%@>h�ڜ[���"�!�d\2:v��&�H.C+X�Va���!�$��8*�Z���9�{���h�!�ׁ�0�H2&�F���1W�!�dK!`��A�DK�uѪ�a�nO-0*!�I-Fp�W���d��q�bcǓCm!��y�.� !i׹6�,\��!P�MY!��9�YJ3��-��fG�M!��Q/_��u���
0�x���:j7!��_�[��*��1r���rml�'�b�'2������;'+ �i:�L�
I��v�|͊T	T8gu�IU*D���ȓm����X�bQl�3��ղ%�(D�P�7劏�1vؘ���w�1D��Xp��"��p*�R$~kp��/D��YS"H-xh�����E�4%c�'D��[�G�0O��M���܍%��l�R�'��G����]�ܨ���H�\Q��͙\'nB�I�%�4�C�*ܿ,ؘm�P�M f�(��0?��l�5k
�z�!�o��19� _�<�S	ֻC��tY�oB�VB�sR��Dy��'w���'ܫ(7T@#Y=f&��x��� �U8�AŹ.�����A����"O:,H�(ԅ9��!��D�	���D�'��'�r�'�ў(����/z|JI��킛G��R&f�y�<� �� v�!�.�1��(2	~�<����U��4z��M�`�֌p᠐z�<0A�)"��2`��%; �ЅLv�<��'Q Y�p�˚%I@0=�G�s�<���ۯws ѐׄ_�!�a{��l�<1�,ĳG�D�C�A�q��E� B�]�'FaxR
Z�+e���@NԲD��y���,�yR���D����f�-{~��dA���'laz�a����ڷ��1!��l�S�
��y"�S0q�;���3l�1�#W:�yRHO���B1�î/���`R��y��9�J]����~���KC)��yR��6{Ӕ�)0/�I�h�R���y��X�in��U*�9����[5�y�M�/{�K������yRR26n�'��4�B屧�Y��y�ß7N�0yP�S=p�4Ӈ��y�ÊV�H�B��D���
g����y���0��9�M��C0�ҡ���yR�V�KmP�����:4Dj�Pb#���yRB>co�u˂�R�&(�0񢡃��yf
��.I��
�FY��C�(��<��D��t�\��r'[�N�����A�!�F�
�j,�GD�E��s%��9!��/:Pxm���K�f � V�Y�!���4.��j#H�q��5���GLg!���=Ǒ���/L�ճƍN>�Pyr�L3p�V���m��Jw�$� �y���E;2����J�F��T� ��<A��d]�<႔*B�P�h�����!�W.6��q��/$�
��@G� �!�䗾t�hz��W��J1`<2�!�dF�FX�g�"h��%��Ӑw!�D�	jeQ��I��"Y�sEY�n!� ��i����X9â�}P!�Es�T���Y\�� �"+s!���Wg�鈔��S������1c!��&B~!{Q�óQ8�����<!��	w�D�c�͆�*rP�s!��`�~��`ҜC)�����x�!��)=n!ҴnG�wo�]����<<�!��q�b����Mbnʸ�``ҼJ�'5a|��ǆ{>�$�V F�B ���,�y�D���������>o��jO�-��?i��:JŉŠޡ�Z��EなDL^���'�5�4'^4��p��LI�'(��'�J|Ka�0�����Q6u$��
�'-\���E|Xx𛖀�{05z�'��XA���bI��!.r��+�'��ڵ��?�
��Ua;jh��+�'+ܘ�@LۏJ�,��ANf���	���'p�>�I�t���s���2������X;9X�C䉺
4 �Х@�!��Y5��1_LC��v~��pt2F":��¼:LB�I�\�>�u�ӸGT��Kf�V&ʓ�hOQ>A3���ҕ  
�c"ΑKA6��+�S�'l�V�z�n��L����A�,�މF{��O-p	{��C�t�]�ѥË>���#���2OH��� nnZ����;�"OB%X5��T_��(����I�r%"O�P����h������xyr"O� �(tNB�VJ<Ӂ�F$j3�=1�"O0%����LӔY�N}��q�����O���*�'~%: (�ܵ1�H�ڧ��7T��UD{��OÎ���	�%T�1aɄ���0�'_����E&zJ�i�A��]��h�'t.8j�I�\ry���5Q�^� �'� �
 ��8;�^mkЬM�Ih��Q�'�y��K,�XA�n_�4�@� �'3�M��lL L�"��p�>.'����'�J9��'�x�k�fUxlN�*-O8�=�O��	�{�씨���*X&������B�	�
D^��X�M���`��� ӸB�	4$�Q���6Y�$��3R�*�~B�I.A^�s��@�J[��B�O�X�jB�I��ʹ��OK�|���QHdB�ɩ�6Az�d�(8B9��HU7Z�C�I�~_L�G(����*w֋�n���O��6��?E�<y"L(,~Ёakׄ�e�g�<	�ˋy�j@��C]�F�|ʄ��b�<ٗ�O
wi2XZpM�����΍a�<�wоZ���z�W�l;-LEh<��k�#E�$p�� WhHA�mP-�y�h�q�@�#l�S���U,^�yR�� ẽ��'6M8� �wh׊��'�az�f�c�B��Fg;I0��1a$����<�J>E��-�;vpQ����FQ��ٖ�y�̰B%H��W$�P��������y���;�L%�ƥ�K��(!M����x҃)g5�g;}���`� �vX�O�q���u�΅�v��B<b�'�ў�G|R��DD��!B	{aĎ��xX �c	�'�N��h_�Aj���cͅn���I����D>��ӧ8����Ӟ@�Pi2Q��3"�@�ȓj�,���U[��Ń,A� �ȓ��f�#'�2$��BH1µ��IR��+ԃG5L���hAf��ȓz���#g��a锱�W��,G��%�H�	D���'��P���6.p)B.����i�
�'4T��D�!�6A�h�L�"�'�<񡣢��M<b%As�0*Xe �' �ԛ6�T1d���A�M(T.>�#�'J�L��P!"�e�d焳yk����'_naaAbډX�P]#$��7D�-A�'���q�M1||ڳ�Ք'V޵X�'��5�
S���$���iIP�'�l�S5�		B����𦑍5F0���?1a�Y(Sr��D��W�iN��y�j��TB<��A���'
7jbj�ȓx<P����(���dԽi�L��ȓ!wj�b �X�!�j\����]0Z�GbZ���|z�F�"(������̏|�X����p�<�hO
)��L`���p���/�B�<��X)B��u��jܻr�ԙa�AB����
}�Ji�fM<^�$�b�<'fч�6X��c�<_�݋v뙒o0�ȓI>��#�A!"w
8r.�la�ȓjkԠp��T"��������]����P�k��^?i"(��� %l�"��+D�`��J�+P��4L���p�&7D�d���܄;`\l��K���) 6�'D�\k��R�t <h�$'Pb�mvA&D�����ԙ(O`X5��$��!c7D�d��� ��p"�/һ3�*e*!D���Ƈ��K�q��32��Y���<I���3� �I�� 	&J%��s�ݟP.�ѫC"Op��	8�`]K�&��5}��J�"O~��� ��:�dX�%�+Lֹ�"O�Ih�+̪3��D[ě:8r���"O�kK-_ 	���u-���!"OD"
���\q����7^Q�b"O��(J��I�<�b≲A��hr"O���I*#N8@"��1�[��"O��*��� e��u��,K�Te*1"OD�c)]<	���K�\v�س"Of�C�� l�#0/^�9jr8�"O �����(�FH���Y�����"O⥐�(��z�$��Y�G�0a5"Oҍ���2HZEpvL�~�hya"O��0��d�T��d��|���!�Z�����<Ȑ���זK��4a��݅5�>��0?yv�ox"80w�N���ㅂ��<�7k�?R8`eM�g�8HHs�g�<���ޕ&�N!�Aؖp�fP�g�<�ĬJ9>�<�הG��p����k�<��h�&������րy`��j�<1�,�!H��ȋ��e��^�<)�çj�f�I���!��XZb��o�<���AO��8��FThV\��h�<9p*ԤXgj��g��2.ҡ�,e�<�Ta�,<(1� �n����Ϗj�<aǃ_5phLrD)QtӌP�Ԥe�<Ѵ��?���
3�s$\j7�]`�<��-��.���_�|��IЁw�<�6M J�E��.J7tD�Q`q�<���/i����e����)adX�<i�o�>X�DPF�
&����TU�<բ�>0,)�f�	(�F!&bWw�<�P�յMք��p�z~P�0SMAw�<�J_65�
ic�*T1x�� �w��o�<�Į	N���h�N��)�ڑ���i�	hy�X�lD�d,FP��] ���$\�=X�З�y�!S��: �C�RN�L8���4�y2�B=��
�#�>ʅi �R��y���3��$4q($��oC$�y�-�Pf1�B�-�p����y��^j̖�q�������A�y�#O�V��Xr6W�%@CQJ����?����e�4 )JgA-n���g��y��s�N4�E�l� @9��Ƃ�yb�Ѓp����@g
j�n��CD��yB� 6����s`��y�t��C!K��y"� 06��W)�q�؍����yRN�3�BkCѰ��eO<�y"B٪ H�#3Ɋ�e���P$�]�y���>ltM�-V���s�ߢ�y�O̢O���P�S��ϡ�yK�i��q�F�\56}���S��.�y��d �(�R$)St�R�R�y��T"�x������\��y�޻0��1�6�Q�Npa j'�yR`	i��ȁ,%b8i��_��y��0�v�H`lV� ��sCG���=y�y��Z%�X��'k[�qQBtS�d_��y©$E�J�sa���A�&��y2ć�;�h�.�|(zY0�Cѧ�yb	S�*eʭsw��y�T�a��
�yb�пb��YO��oTrd�a���y��܎N�b�h���=f%���a�Ӳ��'!az
� �(Qq��5���WE��R���'`1OQ�q�֏z|�`��IQ�����"O<��U,�G���q#/�F��l�"OP�g6w1ܴЎ��|� j�"O�	;��I8x��xe�G9f���"O0I��$E�i�����G��ʟTF���ܫj����@f.9FL@��ˈ�y"���U�Bꞣ����uc��y�"�zk
�R�-�v�� ��y��= %p0Q�CA�iX��S�6�y�
6 xb�]	Z�A�R���y�dJ�"���q��V�f�I3�Ρ�y U�|��1�D��#��-[��K,��O�#~*�c���P�3� ������W�<�dO ]�\�ׁ� w(�A�FQx�|�'��Yk᠂3/ǖ(y̆2/.�B�',p�eD�U��c�&Dv{�@��'��0�2Ù"E(<=A�Àp�*��
�'C"P;�ҥa�ک9�
��B�	�'�8d�PC�Gv�z�f��G��A��'��u3���M-:(r�a
:+88�'�^e3ǭ�/)52�pgIZ2g%�
�'|��b���$	|�	��7m�B��
�'�p������Q)iֆrH���	�'6H��p*C	7�(p[�A�:d�d]�	�'J���F�P�,���!�I�T%�i�'�T��/�� �b�ү9z b��O�<��3�Z�3(�b ���"O�
�c܊X1�Q$G �aP"O(Qb`�/s�&8�E��[5�U["Ox����^%�0�cg��Ib�"O����bġvmvx�lD �b{"O� �SF��$����P	�v0ZH&"OTA���(/��m��C�B{F�1�"O���f)B6��dj�,�8n(�@�"O| H�E�p
�c�+^�H ��1�"O� s�f��a,b�B�,.A�<��"O�%I�)��%j��@�%�2$@�"O",�`�O��x�̉>&ՊQ��"O�xч��H�>�k]�#�n�3�"O � �%¯ex!��ĚX��9R�[��D{��ID#���Ȁ��l2T+�X�!�DW4��C&�./��w*?.�!��L$Z4j��Z�İ
I�G�!�D'y��q�d,GzD1�VH���!���t%��T]���R!�#b�!�D�v���a��J\qqO��v�!򤓋;�Sb"�\�䐨`��!��۫%Q�-�s��r�>��M-�!�DA�8�V�I�vnQ��Ã!��
c�p�@F�qY�%Ⱜѻ`�!�D��'Q�����c3����BVQh�C�ɺgE�`��
)X���F� 	tB�	�GZ*�� *��<n^E!צ��'�B�!A	�4���~�k��
5K�C�I.24-J�A��Z��x(��'D�8S�XctҡI���جc� D��4)���NM�5�VF��4��2D�P��i��Pq��΀�OJ�W w!�ãFB�@�2�"8�:�i�@V&J!�B,!U��
�"F�\��a����S�!�L6����Y��RI�`��!�d��B�*��2h�w�\فO��7�!�Dd�0ؑ�������o�3�!�� ��!.��(�8�G�}4��E"O��1���G"�P��D��Kq"O�a��C	!�.����&a9���v"ON���/e�t\��[�N��"O�u�䌓+�h��a�I=��c�"O2�i �
�d~�#Da��
�Lm	W"O��)�+��0�y��I�j
г��'�ў"~ҥ��A2����F�*	�A�����yR�M1-���2b���N;Q����y��� >leSWB��K��d�alP�y���-i�$����,K��!B��yR'�Yb�{�>0�I�)A�y�K��Z�:`�2B�8W;�IY�%�yB,�?_`"Ԡ���|;d�A���y�����6�2
Q�|h�)�)�y�	�
��U�E�6����W8�y�R45<�j�_(Xf|#a���yG�T���b��L y��M�ej
�yR@
3Nҝ�רW� Фux��	2�hOn���O�܄� w%���t�X�-�,�[%��2LO|=#�n�� S��Q�.A�k�\��"O�Mٴ���S?��)#^9x\�S"O`�Z��
bb|0�D֩~��P"O��	�;xf�Tz��Rf���h�"OV	{�#I TB&5�U	�.�7"O� �pፙ?�J��� � d�4"OĈ�RJ°�;���<�����"OFu��R?���fhva\ 2�"O�R��ˑm2��8���9`L�r"O,y"���X�q+T��<o58z�"O� L�ǌe��g�!B��)3"O���UBێ�^��"�Ȟ)@�
�"O�wݨ^
6؛�)�A���8��'���C�i>y���@�a�TXCᑿ>yR�'N��y� �b��p��GnS 5�v���y��U���]��.��l�&�Av(Z�yҥ#1?x�`2	&p��:FhJ��y���	�N}���G Y��bR��y��|���1�ou$r(�y�d��?�F�9R��z�d��ܣ��$:�S�On�K��;��-�g���K�M��'�<A�E<\���"�W�\���'UNe0)�'y�!�2B�'^x�b	�'bB9���B�v/>E��H��X�\H#�'Rz���hH0pn|a�!���Ȩ�'t��S�\'�q:D-�#"���
�'Θ4S4	#}r�y���;F�����hO?)R�$�B�CB"U&A�K��B�<�t)�[�b���^'k����X|y2�)�'�nu�cmH'8ߞ�a4�F�T�V4��C���k��58P`�I�S�,�P�ȓPB�DM&y���7�B�Ĕ��Bah-R5�Y�ArJɊsM�����ȓx�5����#p쬠�D�)�j���^)]�D��
$� ��4,̤Q֎=�ȓYK��I)�N~��/
;2�8��ȓ0%v��e�R�?���ㄟ+�P]��bF�qW傭vݴ!�7č?$&%��A{4\q��ڻO�Rp)�g�i�����&>|��G C��(�,�W|�a�ȓ%䵱Q=	
�(DoAC����,�\S�OtL�i��Ė����E���Â@�=~�Ad&Ȇk"X}&� F{��t鉑65�)KVi�S�aAEH�4Bh`����?)�Ʃ�?9��?a��z��y� ���c"�[����aΖ4A����"O0(�ee��BE�$ K.D?P�2"O�Y���όD8��(C��m͚8�w"O�8��$�s�Z���ٻ��`Rb"O~-2�(�9�yDC� @w� "O�;�o̗���jC@�nfV�b��'fў�|B�'Em���獜�$�ԮE7�d��۟L����->�m�I^~*���0�~��tH��!N<1�#���̙�ȓd:p�d���x��l�sx(���̚��T�QD!�� �wԎ}��:�¡:�FI�.�q$�� o=�<�ȓIٮ��	������ȓ�|���X�B?�d؆�HhĦ���_y"�|�����`E2�΅V�h�)�IEojC�I5��Jb/<;�CC�NP��C�ɫR�p�!%��!M�<��o`�~C�=���1�a�d��8�q�ZA$C�ɷ&�d�Hq��c��qCG�4<� C�I�I�Wj~$�`�զ�),�C�I�+�ƌ;a�
Ib<H��;Tm�C��o沠 ��!��[tc��2rXC�6󰐳v�Փs���颊�&�|C�I�'�@x�B��5��9���Z�d�B�I�v��D���h.ɣ%�6VoxB�I�*"D1��K�6�$I�P&�)AjhB�	�L�(����ò`����2�3~=tC�I��T�囅P����a��0~~B��j3���^yƤZ���$���	�'QR��&d�"�X�q,��2YD=y�'-�F�W%0���D(�}��:�'��J�
�1��QtKތ]>�R�'}�ะ�\�m�^a�3�K:�(	�'`<,y��I5xC(��"OH-r:X���'Y�M벥и�j�$�ҨV�NI0�'p6�(��PKd PC& H�z	�'�� I(Q����kw)? l@+�'>�Tac��*|P|��3)�5DX0���'�T�2�hުb|�&��H�>1��'f$��ӎU�%B"T�F���BF��'x}��ʷS��|k]�;I\��'g"1�G-�:\���O H
�'����E��?Va��S=,�L��	�'v6DIS���
�� ����(zc	�'||d�2�նh��k�L͏!����	�'�>�pk�K����Hgc��
�'����6�J�j�r�A�!�3�T	
�'�ıa3F�9�:9ZS:3~4[�'��r���|�bZ��	�|��'��2!��J��B�Ë�{s� ��'^d�H��ě0�hܪ���y��!��'���aD���,U���j�.} �'SX\ad&P4&�3��F�eن`�
�'�B(Ѵ��� ����7iA[N m�
�'���1a���E�>a�g��" dLe�
�'$ą�/��S�B�"7�pL��yr�ґe1dCC�.r�Х$A��y�L\�e!
�	\88���E�ϛ�y�aY��(U�Wa�:Aq0��@Ŕ�y�,�X�P�����8�x5	ѪK	�y���Q( ��Uj
���I����y��S[�2b�&`�T�4	
��y�%*y��s"Z�E�N�D%@��y҉ �����Q?=��Q"5����y�CN:n|	�eĭ!�P$Y��2�y
� &����Wj
����D�VQ	�"O��*�ˆhU^����	uO�<��"O�Y��(� `�U�h��04����"O��j$愗q�`9��V�(2�1�"O����/�0{Q�<��!`�����"O�S�/�%�Q	���l��"Ox�`�I�����JPs{�ݓ&"O6}c�oE�rDxr�߾}�&��"O�4��*�{��e�S(;�jP5"O�d� .�@�Bi选�.y�|��"O%��Ts��=���6Yv���"OrAEA�P�m�V�@�9rr�T"OjQxfLލ� �%�N�sbD� �"O>��	�8��H�������d"O���w�B�Č�D`��.ы"OR} �ڽV� ��O8-V�K�"O��T�<;Բ���dG�"O؈�cI^CZByJP$��b�@*#"O��a�ŋ<Vjz��Py|$pG"OR��u X�8}�Y�Ո�b����"O i��)�����IAF�R�j�"O>-�$��?6����Ɂ�g�BУ�"O��4� ?W�a�.w}lY
"O()�'ՎW��۶L�Rcp�е"OFmr�@F.ST���e�%U�|��"O���(W锨Ie��R�N��"O䌚�o^#��(*�㚜z�L9!"OD��D�P�V��%J�MR/�ޙ3"Ov��f�Ƽ4,��3��I���"O���SK�,F�!����g�
�YU"O���؋8��\A����5WrM#�"Oj���P;i HPJ7 .̥�6"O�y;��<e^���"��QT� �"OZ�8���W��\)ЎN,xP"O��rbo6wL�x���ҩ�0�Q�"O�tbV��^�f�Pc���f�J�XS"O
}3sNG�j������\���c�"O�ڱ�N	&i�4��U�{ҁʢ"O�����7N�v1�\�US�x�"Ox]P��H!7����:<�#�"O`Y�R�S�isz��υ���2�"OrdK`P2k�(8���q���r�"O@�+�hͳT�ik�.N����"O�A�pjԁc��k1̘�|x0���"O8-��
�p�0�j)0`�4r"O2mxRc�:#��QهG�+?a+�"O���K&\�8ڷՁ_#6�0B"O��6
�pP�E�L��Ho"O������MtVM����}��	�"O`���D�$��EF	�.p�@�"O&�h=ˈ�b%`G�
jH4%"O�� ��9\��If�Q1��P"O,4K�j�$�x|ӆ�,qE2hi�"Oj�0�����h}�"FS9���e"O.����ħO�B�����/}zr�"Ot�ȧ�F,^G���FA�-�e"O,ܑVI��F���zL�	�  AA"O�i��bT-8�J�ӡ�'�d�t"OV�+Ю�wZJ%P�i��M&�Hp"O���F����TbU.h��%"OFTb$</���a�F8R�
���"Of��Q1�Ȫ��3K��ҧ"O�	a��ф6Q�i�5)�8���"O^�BuC2'5llfW1H��s"O� Ԡ���ښE����N�0-&�"OTШ��#ZP�UB�ͪ 1�w"O(�{���t���'K�"�5;r"O̡��bG�d2�A
�9J��,:"O��z��0
����aJ�6&讌R�"O:��ӇE,ۣ"��p��\��"O��[�$l5FTPtc�g�¸;�"O(� ��h�Upb�[cz�j�"O,�¦�G�v�fx��YFDX "O�9b��\* X�F���T�H�"O�Diu�B�s �!�"�f��r"O�eH2l�*oY0]���QkP�j�"Of���PV�� �-vSX{t"O�%j�JI�Y.D��b_m6p9�d"O��BB�2[q�}�!��sDP!"O
�#NO���@Ѱ��9"���"O���m��3i0���E�� ,��"O���
�d��M��%W
�h�aD"ON(�RNV	H�ޙ�v�7�8�"Op0!��39�]P�D�*;�	XQ"Oll��ДvAf��A�G��Y�"O��e- /K�蚀���u�d�%"O�-�W!�z#�d�p�g!��\�z��m�2���l��&�!�D�p�j�C3K�-8�ޕ"!C�4�!���HN����`�;N�ީ��o2u!��̓7:ъ4	���
����A�*�!�$�f�ص@C� �phj�(�n�!��L6�J4��:&�]��]o�!�D��-1���2`�y���9E˿xt!�ą�QB��S�����`Q� *�!��Y#r��i��A
2�����ϔl!�$��D	Z��s.џ|�&�S�d��Bf!�ǭ\bb ����'t$���X$i�!��#sXm��)M�$"��d�� &!�V�]=�ēV�M�?"����
!�X-B��{E"͞���4	T�!��U�`�J�fű]8l�i�)�!��[Ha�@�T:b�Z����l�!���,\�p �U=1zX��B�;!��%��9į�Y@�c�C�;,!�M97Z�(8��4  �6��=%!��ώsed�*e�́{�@�QA`��J�!�$Y	q�� �9����G�ӥj!�ĝ�&�Z9�� ?Z�$�s�mO�!�d�� T�PiҧI�|��U��d�!�	�#lz$"5$�W||{g��6�!��Ds�D�3յ{X�h𗂄0$�!���.#>��"��BPG8��0�U3�!�$	�U�����(,4� ��\�m�!�Ւ}��Q�I�7l&̈�7�
6/!���)LBUǭX�/-�x�GG�c0!�DH��p�a��˛���V��f~!��׃�>ԣ�nD>@��vN!��G,C6�(�'K9O��D�P	!��D&RE����&�p�Y��T�i!�d�|A��5fI�1��ɐf��d�!���k}���b�/W��}�Ԏ�'=��Dy��'�������+5�mȱȕ[�ޱX	�'(��2O}��3V�_�S�4<3	�'��X�RS)B*E(1(Ԡ d�Y{�'aXp �Mܬ�a��A/0N9�
�'J�MD�X>_C�T�H4߶ Q�'00��f��0/�d���R���#���>ʓ��� `��B��)^�̴`���e4(�P�"Oڡ��ҁ[��l��²��X�pGyBj&�')K� q'Z�S��ŌLcH���(���jR)�sT��9"�A�4��4�ȓ�0qi�#�`S��[��*T�ȓ_�����DRTFX��{��pD{��'Tt�8Wl�6�X[p`F/�4��'�݁Ҍ�}��������?��*�QS�B��S͚�끠շ)st��'�ў"|*R��$���I�2@� �'��t�<�hʧb�H���?H�4[��px�Ex��� ���eϕ'e�E(e�x�#A
E^�A+�N�G�J�b�;�C䉎׊|���S�:S�k$ɖAS�#=Y��T?]Q�д=�vq��+^�/��Z@;D�x`��G�U�nآ���4.Q���E-c�b���S�L<q��!��h��,�>�li�,ȓ\L���	B}�IRrd��e�K���<�!
�3�yH��L�:���.�v}���\���O��~�Պ��A�d!�&�ܺL4�5��J�\�<1�
W�� �J��uB�D�2�U}��|B�*�g}"��,���z���j���i�>�yc�%xpI�F�6.X�D�'�M�	�'(���v��+�<oܭ|����"O&�2ǂѰg��bP�21{�I)�"O���v䓰i/\0dV2�,�h��I~�Ie��x�-�4���J�H��V���>XRC�	>;�� �d�A�'�0�	s��h��� 3m˄[ �� �'��0S�'Q��:A
��HҎ��RQ`}P�`�p�����>���9����#Lq����g�q�{�^�L�Po��9tH��P� B�΀�sY
=��I}�'�"����޷j�:53g��G�����>�#}�!�K&xpj�:��$4��0�JY��B8����eH8+A Ɇ�8�ژ�E��,��4����O=���U���0�M��a��@K���6�!�Q�r22͒ �ޅ4�Z�b��E��p�Ն�ɛNf����e����ِ�+7�C�	2poH���9q��uS҈3Z�yE{��9O�9����7:&`�n"c!����l7D��ڶE�b�:�
Q��XLn�lt�@���2Y5��9gG� |��y�ȅ6�
���<�� I����RŔ-I��H���ě��B�I,_뒰X��Y\��4�fg�&p~�B��g�i�/��l���q@e$2B�I�F�qC�/1�|��%Ԑ]�b�d��P�'��:�F�9���D�v�2@"�4Z��	W�'�iD�4�	IS��AeQ8E0��,���y��'Aܖ=��@��2eg������Bܓ���m��:}��q ��2s�igѩl\��0?����r�E�#A[�2c B��)��O|�[ v��&c]��@�υ�Y����I'��d�>Y��@�@����%Y��u��o[S�'���=�'C����H�*mL9i��!,:x�=������F��w�,	 � &
��Uoݞo\�0��-�q3,��L�c��0� Ȑ�y�?��9��V�<w>I��*t@�Xu ğ]�C��4R�� -��f����wǆ7��n��hO���D3��p!�;_�x���, �V���He����CCc��^!94�%:p1�>�����W��\�+r� G[�4!�K�1��'��3�)��U;�E�`ɃV-t�I��	j�!�$�.9�v9kC�H8	%f�bUo٨m��O�D2�`�IX5��J߂?�q�M�?)��B�)� Υ�&��+��94I�@��Q��"O@�Fa]�s�X���R.��$��"OF����KȾ�+�&�"u��tӂ�'����;#�.%�|Iۦˆ�ՀǦ!D�P�c�N�j�aaP�fF����G�>a���S3|.��*�/�$Q�0I�[6�"?)���PcR�mЀb�\� ��k\H�O���D�k���h%�9zl}���C!�D�;�V�[cFm䎑y��)!�D�i��@�˅>�x���N,xQ�`���/~B���v�ĉOIjA"C��f_��P���ȟ&�0���U��9�W ���v�Y��'�!��T�l�+�(�Y��r��+��D2��z��~��S;W�n)���O!m�	�E�A�ybM�V���2�E�gG��0%���yR�6g�YF'�-,�"iS��ީ�yBI�\�P�e@5&2\��0�y�h��ٓ�K�!�XTB�ᆫ�y2(��'\���"!���dH�$���w���O���CpD�ds�8�R�5<� ��'Y��z�A�\	��cl�N� 9�{2�>\Oxc%�B�#u�9��X�7J��G
O�7�I�(<���E_-xN�D�5���a�az�D��X�B<���tE0`˃���!�U�ØmAF��oB��"�!���2y���ʊA<�y�"�J�\�!���H�h�QV6o�n�	s���8�!�$U�9��xZS'�i�8���[�(�� ��ɔ���Fk2-(s�ŏe�t#�"O�i�� �+6��Ħ�%��Q0"O
�"��+^�*$�3l���"O� ��ː< ���#e� c��S�O��j���zJ�]r�g�?6���&-d�܆�ɲA��ā�τ8�tS�G#����$l��b�8с �7�
t��!^;+�jkfm?D�lH4�3k�i��iZ�#V�Sv�>D�T��+���U��&Z7Bf=[�<D���$B�~�<�$���p�H}K� :���<9�R�x\�,�!�� S^	:�G]x�'�Q?=� �Ӑ�P:��Β+�8�{��8D�ؠA��+'
d)pҁ�Y�>@X��<���'1����&N!g�r,A׍�8'`A���:lOFm��%W�r �)�u턣UQ����
OF6��7+�"�ؒ͛�=s��e�A`�!��M��� ����7o&�"!�Y5=��x��	�)*Ƞjv�	���Ό$O�>c�����)�ӇVz<ਖoE}��a$���2��B䉺2�@�"Jj��A��M-��+cDB�S����(q��H�g@�Җ�¡nB䉢'��d+l ��"H�s�K3=4z"
O���I$l<����[-lf8��'�:Da�S��y6���}��dX�'���R�2D�p�䢖1:��1#� R��!+1򓿨�>��V�Kň}���9Ex��Z�>O>��U��8 ��*��W�*j��z��Ëp���aAÐ8�P�*���p0��O����Ԟ!�0���"�<-��m8���fh���C䴟����'	�Sj�aʄƐ*6)�tJ�Y��B�I<'V����r( �(Eo].F���$?�S�O���:�I� (� ��(��
����4"O 8�ƩU7�L�����d��8s�"Op=pvMؑ*T�-�"f%w>���"O���V���_vVy�CE�9 �M!�"O�5����V:�;����$�4�qV"O� p���l͹l��y �M9���9�"O<U�� <&t����T�j�"O������}�e§�/x��0B�"Ov ��"�.<��V�G!>qqw"O�-"��|�P�0 �2X��"ObX�2�OȒ�;����#��,�"O:�"��8D|4����3����"O}����]���"ЧM�+�bғ"OZ	���ο~�J)pW���.��"O�0�d��W���rC��rx^��v"Oƨ�g�/,C����薓-Z��I�"O�\y�YmT B�	fQ��÷"O���j��8c( Bvd��q+R4rP"O(J�`����碚�U����"O��pSƊ7L���V;N��5�@"O8u�g��KΝ#",�:��3"O��-9O|L�qIC�R��]���yi�	���cQ>=�HXs")N��y҉��2̌�ό2�� �'���y�HܶK�̸#"O�-���kG��y�䎐o����6독 �R4� c?�y���-w`�J�[�Dը�E� �y"�#-�vE���*u������y���1�z���Je�2 �qʄ;�yR^�d2��p�T�VѪ�Dd�0�y�M�����+�%�A���y�h�%�����Y� �¡���R��y2H���SRbj��Ɵ��y�i	������J:�P��EV��yRj��h4<������p3 �5�y����F�`u�4�	���F���yR� �,N�4o
��H�/���0?��$�e�X��E	y�����a�	��,N�<N���8\��>:KP5�g��p�<���4� ���*�@�RӉm�<c��1E�h š�&Dʀ͢��Jj�<�t.�%0P~=��#(��E"ǆ�k�<�A.�f@�cBã>��k#�MH�<�0�٬���.ܳ>���I�b�<9��1BN��$�J�T��	���U�<i�� +���6��`�cT)e�<���I�d$I�h�I���02�Uf�<Q�X�,����'�(C�� �(P~�<A�	��J�Tn��+�)�m�t�<Yh�	[����%!�~�h�Bw�<9��\�;������X'��͒R�Pr�<��"k�H��ЭV�w��i��Zi�<�����@��%���=cX����VM�<9��Y4�I	c��X�\@�q�<I"���Fqaa��8� ���Vj�<ѡ3`5�T��__7���u&`�<qg�*Z	��"i�_7��S-�^�<!Ǎ��9טqh M��4S�g�Z�<a�jJ�:�V�§H�Xj|hH�kZW�<٧c�L���*�r6�-BL�<I�j� a&)�o{�4�D�a�<�C	��h�c�� o��`ƨu�<i�� U
h�[Q�L�h#D��1C
l�<�wƗ,�P���L���j�Ai�<yg�MH���	ط=����f�<Q�eڢ7���h�D��%ǖ��%(\a�<q��{�y1�$Z�@Z�zrC�k�<q%K�2|ؤp��&}��!�c�<iЮ3E$Q�q�*E�
yh��RE�<� J�uHb"�Q�ti�:+���"O��Q6��uN{&�%�M[�"On��!T.L���#5΃vz�т�"O����9c@	����'r�pz�"OL��B�G$<���#E�vǶ�ku"O��`�a��3�$yb�J���Y"O<)�)"uHvEbG(Z�v���"O�z�˙2��c��?,�Nm3c"O�4�RO�.Z���D�Xξ��"O�%h��ϴ[5��	��ɷ�B��"O�$�Aи?J,p�m̞m�F"O`X��D��'���5+�,~�J@�c"O�h1�DҚu���%�14�H���"Op�C"�ϗT�
���f�D���� "O8�ZN5��� ��Ir�"O~�;ꙻZ/���K6��Q'"O��07⎞U$=k�ˑ�k/F�c"O�� �B�:d�p���@(��'�\�a���8�Go�?w_�uzd�ӹ~d���-(D�����QP�<�0ҕ:���7L5�I�h��{����:�	@ /)n
���M2C�I�V=���*�7<`���D�@�1u�QܓU'�>�!�&t:�#Ǿ��K¡=`����ȓ�L9�-��Fiԙs�n�U�o��D��I��'H���ĎJN��W`�]#��(�<�����<�#��4f�*���»-#jXң �`�<1`��NZL�[����blF�
F�P����ׁ ��y9�A��6ml ����!KТ���xc	������%S+�~�N��w�@��h��D�;�z���K�7��i���:C!��B�&Y#e
R."����,N�_�!�ƳHu���N�	Ǥ�*"J� (!�ÁV*�Ȳ������jjqI	�'��Qc2(Ǖ��EVe�:]��A!�';��3l�	J:.�B�QWx��B�'s��XtdJ��#���v)��'�c�AK�O���8�Ǣ's����'���`$�L�\�N�0�lƦ68",*E)�G ���I�{��H�T�6\��`��,H{,���1n�>d��3}bBM�U�T��T��9������y2i'L�*$K�B.��� �~@�!X��$!��E	P�~�e/�JG����tiIȭq
bT`V���q6��ȓL�E(�gM w�T �a�>,�$]��'��<y�E:�䫒����9O�Tx�
�R�wG����ę�02��q�E �\��� �V��D�}0t͢c)G+:���hY�bX�#V�>�x��+O~ �%��[��p��4mbH�)��3>�
�� 	u��"=9E�75.μf��[	Ri���~2�k�Nx ���V)�@I80��Q�$K����i+�H̇�Iæ��&a�]j"萦O�G�h���,�8h�����h*���%�yh/6pL��#���Id˟)_�!"�K���BB��$MR�+vɔ;)\�܃g<d��%P�b�@��1T��D�A����(oV�0ż���ϣ}���  "U�Kz)��-@8�@��L�62�3(��ez���tG�A=�L�B��0��ּi2 թ��O����Ro���q	�E�N�1R4F��1��pS�X�+��Fy"MP/B��FA�4�����*)��ɑ���AQ��e^<PdF��\�Ⱥ��� "dl �e�A��xzǧ�4��(x�.��Q	 x����CA���'��.D�(҇�|���O:�n�G�oZ=�
�CD�ڧ7�(�`�����DQ�i��H�L<��~���"�F�T��LЗ#�>橙(+plt��H�}9VЙ����?��Q��T�ǃ��4��w(D�`�bBUkr��%oX� #�3�Ȁ�+>���Q*|V�\��i2B��a�:a%F
%�~U��X�=�JiC���]t�X�4�?�'ۨn��\-6\0���dTa�\H�ф�}�F��DM��w�'���z�	[�+✂q��
(:�4�O�����J�bΨ����7�Xk�
�A�"@�F�9G��yi���6k�d<%��I<7Ɛ��֊�;qQ���	��LL���)j���7e�̟$��̅hچ6�v�,��D������r-�П�CЉ�$��@��j�)f�)Z�7O�
rAƪ�ēO���0F��+�PH��M��\��,�v�I�`1��	�k��鳕��l����=�g�? "��"�A97FҨ��O�lh�@�x���%�1O��q��;��=�|�xdk��q�vM��G��7㦘�s���F��I<=��y���|�;n�ִ���W�R'�1�3"ڻ�Px��6��h*A�\	I&������D>>I�qn��Ɲ��	dR}@
Z�aC�|X%�2;���$��j��ٓ�$����;t�5�& ��/&8Y���R
�'_��D'˥u�8��'�[-d��Y�L<ѣϔ6X�>)�N>�~*� Q.�
L���b���ʧ%�i�<��CT�P �s�
�Kj݋b+Թy=qO�M�5�<�3}roF� Fꍣ!dO�x*�Q��R�ybK��P�F7y�L�3�"�/�y���^�p�����kt����AW8�y����8ۖ�!ŌX;aMZX�G�&�y��2}�����3����ƌ��y�� n����0�5��$�a)�yRF4Rr��B��˾-H����y���t'ް93�K�=�L�p���y
S���0��"%�4���F-�y��@, C
��Y"lR� d �-�yR��.YSL�����,P�hRAmM �yB�,=�0��#�M� ��%pāٔ�y2�M24%n��k�I��]4�M)�yH�g�}a��X8�� �$���I�r�����(pF�E� �(c��8�I�9O!�D0��HJ���[Z`$c�H� `2��Ob,C��!b01�1Of��g@$8MP���gA�ȫ��')b�t��A��;v��i<�����xU�t�aR@�(�Р��bުn����e����Ox�r�^�|���;J|�"�ٴ%1y�G�n�x�#l�A�<��H�+��=�V��qn�ReMQEy�`�����G�W��S�O����a+U!M�D���ĳ#��e�ǓU�<} 2e>͎��O�gt�P�lݞjF����I�<͘(�GH
�� ~�)��NQ�3�	6~�h��@�S�~\rdHI�hv�;�ဴhPM����oѭr��K|2�m� \�����2N'��@�'�.Kx����S����"9NV}�a���/u �H�f�M���r�i�b'	1c20p�OL^e����+s.��O�Ll��0�v����b�r��c5�OT] ��&n�7�>��y��Έ=��;BF��t�$�Ӡi*�<��<���'v[��� �>᥎΃z|��ƻ%.��#�u�'��!��ʶ���Ђ�9�v�����"?�1z'�¨;tzDZ��_I���8ⓟ���C>���GB�o�h��U�	�6.��S�g�����$��/\&���Ś6^�hQ���K�d�
�&r<�:1��I����.��N�6z��h�'�
9��g[j�'��Y��J�a~~�y�K��^�]3��� �|IF�V5�0��U�P���6�:��uZ��y7o�#��D�"�N�DBZ�E!?���,�4�
�J+}J~B�]�[����#�J�>Ԍ� �f
M&�	�_�Dع5ER�n�R�!�)��܎�;��	�:S\��g�.�L�E����I��<II��@�d�z�'V;����ņ'�h�AT*Ǩq��d9u��!C��l3�ݗ-1̉`4��m�b��,�O�m���!.�b�Ѯ�F���$�	4�0��n��(1��/\H؈x�@�!-�j�!��� N��M|�Y	h���"���`i��`�''�i"�I���B��I^FF�}���_J~�]���A�t�y!���}$���D�4?<���Z�=8��'�����DZ� $،�"Lސ
@s.O�X�.K3L285�9�'u���I��O�}�,�:��I%��}�&UJ�`᧍�5g��1N�jx�Y����+)@X��F\�N3�]�5�� �Τz�R���i֟x@��8y����.;�6�]�R @�")�d˟%eAx��)�)p�챰��R��p>��ެO2�Up��^��cb%5�Fa��R�\�`�'`��)V���(��G��,��=����jR�]�P��k�>��:��Otj!�B/�h���4��#[�z�H�������:`h@�C9����ՙ?�0MY0)����E��O�(c(ʫ
��q�5���	�t�����Ʀ1��>E���"4$�K͸a��]���8]q�(RS�B B�Ĭ[F�4B�$��������.և ��,��뚭7�z��I>��6�~��� ����5�p��Q�4� �+�.m��7O+Lo�t���i�!���sp�ā>=��Å�u^�O����NK���<�H�|xb>%�,^�f4	sg�.Ahhz�'D�0����V	���l��t�*qED[��I���)�p�R��O?�I*U�vP��7Q����%~�i���� h���;ɢD���/)��P)wY��X6E�a'zAɖ�'��0�RQd����P�*��4��QTi���~:.Ł�εd��Z�h��&��d�ȓB�Y��`"+�J��D�
�50Pd�ȓd���,�?}vD��p����2��x���/u�����M�}��-D�����F�\T$�Z:sa���/9�T�a.Ĵ9ӌXwE������/fI���(;��@�D1d{���a1R�K�ñS�} t�h� �ȓ ��� "�E��M �@''H��ȓr����4Cܻj$V�j��$L�p�ȓ8��ѥ�יn��Jr���x��]��J[��5��{�2X��i�.�a�ȓ*���0n҄KM^�$��~-�Іȓ&��Cä`p�QӨ��QP����䃗��l#���G��� �� ����("E�K�vm�����k�轅�ܮK�ΎJ� � D�V�[`������
�Ké[58���H0>e�̇ȓ��!�
�%`�i���&w�ܩ��*�`���*K�@�8��# I�6�z(��V]��¥�׵z�@��GְM�N���>ނ��o��I�G�)_-$��4D��r�� ���؄�ߊ�<`�'?D�غ�	S�j�!M��8�d�9D�|	rnU�Z�x0��n���1��7D�`(��'O�}�J%,qp�4D�,��!S�w2����'�,�BQ�7D���b��B�
Ѯ�#��B�2D���Ɛ�v���CH
s�́�f,$D�0�����l떼���r�X �.D�$Z��]�'~�4Yrᏽ�z�8S�8D�,��T:��Eq��Lz�:� '#2D�`He�B8tL`]`d�
;p�xp-0D����\��� ���Nx��@��*D�X���ߙQ/& ���2}d��'�$D���d�1	�cFM��d~�}SC#D�d"�G��\h��iQ�W�\<�f�#D�l�1Nɛ�8Dh0�O3"�
$�'!D����푕m��@��C&���;�!D��)��I ��B%@�;w�5�A?D������U4�Ņ�Z2�I��<D�$c0�X /Ц��.ņ5ԞY�Q,8D�|��J_���*׫��Z�`7D�"�×''�4u&ث"t��"��2D�lcB�D���������s�3D�T�@���i�	P�N�&	�3�1D���G�H�c��Gj�PI4�A�-D��ҳ��I�,Y�g$
���[%'D��a�d	�^+��R�&y�C��6D��IL0H$~ �t����a�$4D�|��FC6Br�i�c��6X(���ti8D�����ψ�D�"m�,9S�9�3�:D���0I�ny�Ú�K4��c�9D�p�4LN�(�:����_�o��pR!C6D��;s@\�=��QEʖٶă�+D�ܙ�
Q l����O�^�cf4D�P�t�Z@;��E^�#��)6D�Dȅ�K�qW����0��x��4D�ı2�v��9�b!S��p�&3D�$*d/�$D �%-$�� �1D�L�匈hT���K��P�h,D��z��.!FL�F��5f�x�!D�� &���ǆjS �˶��<�n�  "Ob��u�Z �L���?�6	�R"OX���aZ2vn��Sn�@Ű`q�"O
�!Q[�l_�t�Ƌ�ȔP��"O�XP�_�i�%#�EW��ya�"Ol�ѫd�@-p��ϙY�0���"OB\[�O䬐խ1k�ҩ��"O�R <{ذxYt�A���U"O����/�"(Cd��a�G<I"�1CU"Od�C�I�F�H��B(Y�ƍ��'D�×m�<>� ��LS�F��Db%D�(�֫���X�82"L+k9�3E$D�4��*�*Ar(;#�K ���k�O?D�0����[To��3�b�J�#/D��_{ 8��D��<��-D�,r�KY34��ʣ#
��͙��<D�h�0�B�BO𤫖��2V�~� G;D��p^�`P�"�퍼8tQg9D�0{��;X�v�Iq�I�xѳ�7D�xB�AуP�L��U�D&} ���#6D���Ԩ۱�����c��Dh�Ӈ6D��Ӥ��eF�PX�}�&�ʗ!��)y��h
�"��!(�!nB�!��{�pR�L�M�X� .J*s�!�F�w���=4��i�C팈"!�V#:4HQ�[��T�U��4[!�D\�)����M_���e��h!�	�sX��2��ǻ#H�]�ЌN!��]��.��+
 4JQ��F�g�!���3ld8Ec֯]2V=d�ZTk�0�!�0z�8 W�ǀ(%z�E��<H�!�DO�4Z���e'����Y%IS};!��ƪ>��R�K�2k(H��Ñ#I!�@aL@ �D� �z���P!�\#����\�d��ٛw�!�J�B�8�"�O�HOޭ �k�!�$T�$�9�!�J3s60R�MU�_�!�D��:�n�a��44<AA�N�+V�!򄚟4�Ј�V�M7�ˁ�,c�!���;^P9v�<XH���4:
!�$";<��}�Eb$0$Oz�(\�	f�BD��3����/��͒�*ѬуV:BP��,V:=Ȫ��I�u��8q�l��>^��
� \
B,� �dn+�!��1�Ɖ��F>9�l��ǔ� �d��6���K�6?���H?�#��+ox�*���ݰyc@9+�!�?/�B�	2%�t��σ��C ���qBc�	g��HQʁ����`�'Ur��'���"#���y'�_5�������&$�����>��K�M��MAĄ/��!�ªR(p�E�%U�|IZ���n#��D�V��9Q!��p�Q� �S��+���yp%��,ި���<���iw�LQ������mV��?�n�e�@9_S�ICvC_:".�)��-֒_���e���0>8uC2� ��W)z�T�8��E. �|�cGd6Eh��ԍv�P��ޟd�q�'���hŮ��k��4j��MCd% �	��-Ar��q�<�Ԉ�x�}�Q�2 �Fh���M+N��I9��Z���S�[��%�^?!�DW
+���9�w�e��m(?��90�'����P��!𝃃�׺@,uyRƝ��� �F��~��	Qw��6-@&<���I#&�ъ2�85<�i�BF-v��a��U�H�*@��(O�"䎇.p��1E S�`�@j�?�k��D>�-��h"wϾ��gթt���D���4bߓ[p�Eq�*�<%�%�f(��.и%����皳m�v�P��Yr�I�?aԻi� Ĩ��Z}q����Kaj8�%:n����at��xQș�(��4%%�6;[�@������RnO�WQPi�s%g~��hq8O�[E�շ9]�,̻g���<WUru�,9�|���v���˥"لFq�De;^;�k!g�$�z�+&a��UZ ���4�?���z�*�v�
�u�|�?A���E0d�1�L��q��@~�'[�1J�%�#3�qC� �<u�'7Z�� ����ͦ(�ű2�]�@u��0p�84�L�"�Q(w���DT�K
������D�3F���y��X?Z�H���8bV�Q��ן��:�⅁g(��2�=����8_ b�"RD+X4���`���yҏ�?�>�i��)i	�9��J���Q��!�fZ���1��>t�	��k�n	@@�H�[4�C�ɭ<G0�9𩂺 �"@q�@D�����#D���	�%v����|bOh�h9!���q�l��Sm �Px����uѮ퉀M	�O`� ��#�X���[�ޜ؇��)\��h1�Sa���!xD��E�M'�����ܰ���S6t&`+L����5����X�!�d�$2��� E�E2�6�p�)�6FƉ'�}���S?l�ɧ�O�h��`
UF�����:&�
�'�5;����>��t����9���0B�0`�z��OV��@gQ#ڑ�Q@Q�~^�{6"O�{���qb �Q�σud��ʳ"O���f%�L�����<[t�R0"O�$Zb�Ԏ����0g�+W(�3�"O�M��؃]:V ���� �d ,�y���7J�"��D%�U,ҽ0�͛�y��Ȯ\k2��!B�._s��h���y���e[��J�Y��飇D�y��M
'9ؤkAi@D��(��ʫ�yR���F�d̜L�4�����yR�]>	�����8ARȊ���<�y�[�5��,{0�^<k4ʙ���I�yr'�+M9��y�Oזcj�c#ȵ�y�ON;-��ԡ���]�~ Qb�
��I3���P���	(|�� G�5c�t��Ƥ�4R�!�+HSȀ��Ww�re�X)=�r�O�R5"(?�1�1O H�p'�S
1Hw�5,�}�s�'\� g�<C,Jv	
�L�PDȮT���Sa��`؟l��#	�Xe��S��>I��)ؗ�/��%<n�!��OE� ��U�3�'(���`��U�"{����"O�d��l�Zm�!	%Ʋ�V\��C��C�(��֓>E�dD��v����eN0ލ�g�nX���ի3h�O�x����	2��� �� Q��!���&��;=���Vl�3�3X($�Ck�l)��`7�I�N`,�"�\�Ñ�JM��PF�Di�-���M܇U]�*��Ύ	O������o��u���(k�줋��Q�]���!�� 1@�↨.?q3׋e����vWD��451�;'��HT��-Z-�0�VJ��Y��i#��0D�Y![M,����Y�V���r�Xoߌ=�%���Su��!(U��'>>}���)(�ǐ<jȲ4���6���H$n��D��=�ʟZ��tM�m?�yJsh� ji��%�DI"o}����d��j�̄�SOwC-"��*Y�F˓{�p<3tY�-�j�
���ɵE�Ȕ���@$�{�F_/ܶi��̩��O
�P� ]�Fi�O@a(���`��[���Nh9�2�T���$��E��4� ��
4n���Pw�E�y�^8���$k�I�!�� �K�H��S��*׬!c�Qu�)�g,נr�N�Ѣ�ʿ6�^L8u�'�<:Rm���-@#âێ*�*)RM@#��l=�T�Ԩ�D+��O�n�ƨ�N���$�yo�8rWΒ�&\`	iB�Y�����$�"8~+��@k�C9H��!C�2uG�A���Qg�&��'>I pe�:�>����¸�v4�a�*��\�n����� �ɟ8�A�l�*3�nԑ� ��!��#�$
�#�+1���JMж�3W�^�㒌Pʕ|^��-y��3�;-P�qE�D�4M!ФmCud)UF�:,�$��4�@<�JنE�~P
c��xUj)K �1+��e�'V�I�e� ���ϸ'�~���+Q��2��˱bX��X��t�r�H�E�t,��i�ҦaإpW N�vQ �G�L��0?a�F˿9��[A'�seIk��NO�'���2��	4�?	rD��VH����V�Ze��E>D�@QÉq<�����͚h��5�6�??��a�7��K�M&}��i�*DX��D�	��T����Ub�!�D�6y}��"���1�샧M< h'�蓇�>q��'�l�eΞ�ư���
.^R*�X	��� �<`�*LO�n�xU+�?r����"O�	"�h�T�h�0IT4��k�"O4<9�n�'�ФE�:��e"O"�`�3�Ȉ�s�Խ-^r=��y��w�H])G��&�N�A���3�yr��9W`��<�����Fِ�y�U�>NP��Cڑ	`f�1���y���&L��� 
Z�{�p-X�$2�y�)�q�-@d	'q�<�!k��y��8іL��ʬj�j�� ���Py�l��`��eívFe����[�<���hYp��Q��.jpt����_�<QRC��e�"ɒ&%ϨaRD�j�#RX�<��jڲ(}Z�)�_/D0�*4��@�<�ï�+%�\|рO����-k�Vp�ȓ!^\��wa�o�`�0+¯i��y��{D�*���3r�9p5JR!	*��ȓ@��-���F0�Ha�c�:�v���b �� g��I��\�f�K=rM e�ȓ&@$�VN�;F��p"A�]�U�ȓ#|�Hr� ����P�+�\y�)�ȓ��X�#W?!���ĆC%c܅�ȓVLx��'d?���%W�4�\���%֜��%�F�}�X ��Z��: �ȓq6X豄���;��r�.�U�zQ�ȓn(@�)�|�CW��!�� ��o@��8E��/tyX��|�����\���`U��IՀ!��B�t^ZL�ȓc��Q:e���$�������C�I�p�d(���vÂ8 �ɐZ�lB�I�D����Qb��L�H��$���9 C�ɵcʴC5
2?~< ��X�M]�B�	,F3��Q͍!#L�� ^C�G��	3Ռ˶j�M���5��B�	;���0p����0�
C�i�HB�I_������[����*ߑr�C�I($!H0��"7ӄxtΜ3�C䉹w���"�O��J(X�-�~C�� p/�1
���p��5�
�qHC�ɛ����f-w~�Ń&�ǰb�&����2@��� ��OFz�ceHݍvq>��!B�t-!�d[�:tЅ�T �oz�p;��Ɣt!�����dQg�bvH!��j_�^!��/! p@
�HQ-`jx��(�q�!�K�Xo�Y�ؚmhr�[Շ�=�!�$��DŴ a�&�GV���GGÙQ�!�D��x�a�!��#S�0��7�H�/!�(\��-�-�� ۣ(J:?%!�$�x�&p30-Sz^E�ΗK~!�$������U�e��VH�G�a{��!�;y��1��# �qJ�>+"��ɉ�P��Sl# ��-�"t�����K��5R���&"��ذ㞢2��.P�uPFjد�Q�b�ߟ����=9��/��U8��%dnh<1�A	"��������b>eq�J7j7�<05���QJ*}rJ��,���=�g�I�7�!��%IZ��8�.�z��I��,M�?E��dWbF�南�^�T��f��jIt�80F$�)��M	��K䩋<6��a�I�u���҄��6��O���'o9� @�,�v���TH�]e�=o���'B{B�"��h�p֝�(丄A���\�P�!�S8/��݂R���U��)՛�?�B	8�l��!ɬ/(�;W	B:.��A1�ƫ8�����<�bh���a������Դ���� D$l��c��6x�=p��O%*qǞ������'G� �Ò'�)����d&U��x�<�N�d�L�':2����O�"��i!N�Ь �����̬�ڴC�<i*�)]�4ҧȟ� ���a��O��a���}D�`w�ٝLD��'�J���s�p�B����w���r�'� �b��0h*H�P�`Y�`f��`�'+�lI�*Z�k��p�lZ$�qC�'�!�	:8�a�J��,��'>&刕*�3:X!s�ώ�%`(i�'�N�R�'E�D���8�ե�h�!�'��!K��W\*J�x�c��| ��'�0���W�����A|J�`[�'J<ꃏ�4��!�&,ɍt{(x��'�����gL�j�t�Pa�>MZ���'
���E�0K���gHח;�@��	�'9>[$�!�z,��hߏ0d�@	�'�28���'aK.�k ��Tu�9
�'!�h��Rk�0`0ϝ=E���	�'�\�:P�*�<�����l)�\��'D���ց�Mk��0�R�1˰x��'�|hb�o5��� � v�Ј��'�~�{'�q �@�cK1D���	�'��S�hA�-�"E���3>Ǽ���'�j�r�"���\�4�ې4m$y;�'��(�� I3z~����h̜{bN	��'�^1��@���>� ��ȏoM�,��'͢�� 	]������C��m���'��ĚQ�ӷD�LШ��'���'_<Y����A�p��A+C/@��'��l�7Dޞ�\�Sѣ^7/ҭ��']t�O�$M�|ʑ̄!�b���'�V�Z'�4u��q`%��rTr	�'�4��?LN�uY���^8�
�'k:�	&����uc׮�r��(	�'d��t�]
S8@3wF��5�n8h�'���tK�=f���Ӿ&�`���'6J��&��C�Б{����*��[�'~Ő�i�<���Ҕ�ܼӸ�Z�'+�٫`�ih�ys��:V�ȓ}��;W��L��E�#�E>�T���m�|8a���
�>�(����챇ȓ.����u)�E�Z<�rLZ2V)���Jm$�˧�	?�|y �Էz���ȓ<n6�Q�&�q��x r��6���ȓ
��X��DeS�]���T0!�����&� O_������+�ܥ��]�4@���6N.t�P��%zl��@�Hp��	 Lb�sd�E�w� ��(`�hBW��X�p%�b�إPx�U�ȓd���[ЁՄO��MSŅ�f ���8�\�����J�[pC�: �х�3�j5Q@�0jj�z1/]�k_&t�ȓfK��h�)I�|�
���.[�xЄȓ(ZF�2��KrмR"��6���~����h�{i�z�L��Ψ�ȓV{<���(,ty�q �ȓT`b��\���#`n�=Z��U��e�B\q�� �Z�ⱦ�5h+���ȓ{�Ʊ���f;�@�� 
��ȓc0$m�[Z<^�[�M�h�@��8��k���10�v)�w�� m�X�ȓ_���O�4��4GԒC��ȓ�z��PI<Q�t���p�ȓ*�m�鏲o���B���K�Pu�ȓIݼ��cl��Oe&aQ�Pr���ȓ0\�� @�Јdf�0�VΒ\xԆȓq)>)� �V<j�L)��(�5?h8��S�? �9�T�j�L�6�\t�:"O�	hޖ#��$95�9�Qq"O��(ek��3��@qmGf���"OL,B`C��l��$j�-��l��|1!"O"�!�(F�(/��xЁ�aۄ}��"O����DJ�THF�G1��]`"OԐjf�Y7:6j��g�g�и�"O`}���#��kUǈ,�\�#�"O�h�KܹD-������9~��T�"O��1R$�!_K ��"1��"O&=+L����d{bVb�,	�"O���완!'�y�#��%-(Juj�"OV�8�� O�x�H�@1W�|s%"O�x�%�&���I4��-E(R�d"Oj�8f.�(�VM�Y���3"O��X�L�1V�ք2�	ul.�"O�� 0�X�\�}RP'�����N�!�dA�~�1�I�c�|��u�E�X�!��4'P�9�ʜ�J�{�E_*Y!�D�������-��hjB.!���/�t�Brk�R �9'���FN!�$����áF���l�,۬a�!�Q9��U[d!C#�V�Q�=�!�DO�zC���FX�"2����D &B�!�DX�:�rl1�� ".(Z'iU�*�!��ӷ^/��K��3"
� �7r�!��{�� ���$ �����p�!�D��o�=��Ef')�f��O!�N
J�jTҷ��(ƀ1���&d3!�d]�
�%�w��((�sfeݼ]�!�DШ(�2�v�4	�!8F���"�!�đ9e�@���/bɺ�h@��!�$���P$P�g�f�*a�F�?5b!�ҡ.8pԺ�l�R����p��gF!�D�+�zٸ���:&��d `A-+!���EI�u7DN#��i�O",!�$� Rl� K�|w���
Y�K!���3����ǼcH�w��2�!��J��s楉,~oD�G)��f�!��*ArnXSpc�5~^��e\d!���="�����ޖ
�h� &I-oG!��ƚQ�}�$@��d�$� �P��ȓH�NM�rH= �
�F�ĂQ'�A��{8����m:=\���b� �tć�D9��4�G����=Ay�d��P����OE�51� RN'H �ȓ>�^��p+�'Y�!� ��"j�9�ȓ㺭�`,��b4���P�I�ح��=��I�NDa�yä��	HX=���42$_6#��@�� ��(�ȓQ��ċϖD�
4H!O۸Q�2��\!0�ɅO|��3A�ϝ!w��ȓ�Ɛ2��#鞜;g�E�2��0�ȓe>�UcuHA]���sҗ'�DЅȓ7ꔜ��	�dI�1���͐�lD�ȓwc2�����-){��D�<�X<�ȓ9��S1��V	���6L�VZ�	��,�����!XH��"/�:�6ȅȓ~]T����B�0cj� ����Nk�8��KP�2�V!k�ʚ3^���ȓS��9��M1$6b@�b��H}�H��o.^�8�I,]��s�&�����ȓ_��ӈ_�`��rV��P�t��+`P�ۦi�%d$��r��W�A'�Q��S�? ���N��6`��C��9]O��[�"O��: %��,�?Zq	V"O*uB)�#cy`P�ci���ӗ"OJ�ҷ��+���c��8���"O�v//R6��'Ƚ�� �"Ob���D]	Ն�!'L�^vLI#"OJ��%E�2+@1.�+����y*7����ŏ%���y�͘��y�#[2i)7K��R4r�*�(ɚ�y�v�(Q!V�^	?h�3�gƛ�yZ��	�BA13��rC���)
�'���d�8X�
��g�B�4�H�j	�'H`ěT�A�N�,@�7���,��'��|2p�C���H`��( �)��'�`�{��~f�A�ϸ O�y�'yT�k(����0P�f������'���q�U�6T0�@�{=�,A�'PL ���>hX��v�������'��T�Є�Z���;��C2QxHq
�'�-��i���}"��ǈ~!P0	�'F������Bl��#�?rԵ��'.����#r�E'2s�a(
�'�^���n�?"����$%$0S�'��%��E^����B	��'���C�Z���UO^���c	�'B~�)j�V:`{��P;�x��'l���W�!RPkO6G���'����(�<q��� ��QHL��'�&�b�%\�x�*�it�x	�'2R X�J@'�h0AB�:{�h��'����ga��s���x���#yM±��'��02���qc�	X���?T�'(<ЁgØ$�x�@��n��#�'i�����-�!��J�5D�X�Qbϗc��Q��2W�pa�4D���׃̓���g"��P��e�0D�)W/V�H��1��O6j�[@d/D��A'M���lb(O%a��i���/D��'T�q��yH����i�-D������t�쀑 �'i���6�7D�T����y��+1aZ\ИSr 5D���a�So4q��WD����*4D�H�d�X�Z�<��%,T(��	�dG$D����#	��X�0��.,�`#$D��B%h�P��L�$ʷ�!D���9_�Z�Pd��<Tu�m2�� D��k��.D~A�Bn�8�c9D�Q��� ���s�Ю`5�ZA�*D�x1F�>"�Y[Q`�	-8d��";D� �$�ͺYC*�蔧��ỳ.D��z�ȁ$fhD�A�c|�F�7D�\�������勝Y���3��5D�A0�D�9�"(+@�E(hf��`C�3D�@Z��Z"?�d����?afYY��-D�$��d�.I����4:�Har��,D��8��V첀�`��u��p�w�?D�Ȉ�Q�T����nJ� �wI3D����O���z�� ;���Ң�$D��9���[s�ÕOT"<�l��#c6D�T���Z�U��
�E��N.���7D�,¤��
"sl@�`�S�S��*:D�(B���7�Zhh¥,/���@/9D��� f4aJ�ӕa�z�ڑiB�6D�`륦ռ�6��m^�3U�9є3D�� ZX�A$Z�TA�!Ş"�^��"Obu��`�+3n���	�=/�|�*�"O�)����&��4��fR�\Pm�"OL�aF�[_�(5�@ ��V�\�"O���3�߷-���R"�E�b����"O�D�    ��   �  c  
  a  U+  �6  �B  �M  �Y  Je  �p  �{  ��  ��  5�  6�  ۧ  %�  ��  ��  8�  ��  �  ��  #�  w�  ��  �  R�  ��  �    � � $ 4" , [3 F:  C �I QQ �W �] �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z��Yb�с�5|O�"EG�;֊�R"�O�~Q:�F�'VP���Œ�'蠢DO�	J厈���4D��@Q�Ђ:�|@��Tfs���(D��`D�J�=Np�A��׭7����Q,%D��z�oV5H�r��.Q�����$D��p�L���Uk��B�����F"D����`���2����{�& �E�<D��PL��j���H�G��:f;$��S���T����t��n�����^�D��� �F��9^	�F�=[`�͆�Im�)H''��*-���t�S:E��ن�	�H���
�e�pڶ�3<K�̆�;�؄�c��v�`����֭wXވ���t~� �6XvD�e �8�HP��E��y�D�9;�px����|	J�fƈ�HO����"��aA'ݥtǽ�!:w*7�!�p��`�:�4E�*ɠ����Gu��E{���\�B��8�d
5s�.,�(�8zE!�$ǈ`VaR�킍wz�q2T�
�-!��QI�V}z�f=n�����,a~�V���J^X+ָ{�儏v(p�R��5D��)��?1� Zg#��o�2���(D�p���%HА�(��� ��Ȁ�"lO4➼�eO\;xz\���%$��1
!D�p
`f	 CHA�0���-ƵH%�<D�pZ��CX��wf �B4F<D�<��"J!���#����.�aDO-D�qU"Ո0<�i3K��$��X��0D�� @��#aǵu0�IՊ[�zl�s�Of�'�6�NQ���I�k0L�F�_3��݃�!X8Xaa}��i�d	x�Ա$o��\�j�� ��Vhm&H�(#<E��4'u��D��* a�<x��S�RU���Ms�B��D��<3�Z�V��#YRy��,�OҜh�k��Z�:i��m�N[S�'����O�4�V� �ń���/( H�"O:mKw����b�GF	ڷ"O$��$L�GE��;A��t�V"O�p�##�&6yK83�� ��ݬ�~��'�̀�=E��' �R�yB&Ӽ!s�$�DH�:�y�DކE����B�
}x�^��'J�{�A�^]~|ӄԅ<(��B'	I�yb�����1q�E�-����ȗ.|�B≎;삔t�+I'�h[���8E��B� :��)2��a�,���	�3HԮB�	�s@�@���d�j����P�B�	Z�
�"�7d|�b�KD]�B�ɝIhZ�q����*�y�JO�jC�I�ynD4�7@ɫ	�8��B->0�>��}b�f�qiA�'-P�i&�G�C�z���DI^�<�sh�E$4���(�D7�)Z`?1�]��m�|yr�S�\Ӥ�#��J>�+"
E�V��C�I7B�F�v/��q̚���2j��tE{J?�����3>k-���I���A(6D��u@I(S"���n�#^�u#S�y���>9��'��	�E�l���4�\#�4����'|��R��-Mu��;�!a*�e��'��D��EY�3�F�4���Q'��+��D �S��퇺V�N�ر�	�<y�0��+Z�yAP2ez�=Hb��##�А
��~�ў"~�Tӂ���`�[�$��iD�Rԭ��a�$��΅�U)�%a��.P�l��\�.��hǾ �8:�a_� �����B̓'@�1�F�z�BQ�M����ȓVN^��ؽ���Qp§ ���n� �EE�0��Qtn
&V��_�<�ەi�#G�L�f�I� 	�ȓ=�r!f�,`� �2�1�t��=fPH�bd�3!��,�
!H����l����JƑ@��\��OC�f�4 �� ��Q���
� ����[�����-��l@�m�!_~����$��2M�ȓ^`�ђ �8z�Qb�1n�Z���.�C���J�~4aC.$@�ȓp�D�z��

�V1�S)־�ȓM��%L��	B�� �
S"���|/���%�3-Yt��N׋]�����.�ѕ�Q�F&~���̈,M�]��t�����^�U�FӅ.��S2���i�{�J���?N䉇�����fE�,Mq�(�,D��Ѕȓ	� �� ɠ�:��Ơ��j��-�ȓjJ&]!g�B�x���blV�k��U�ȓ{R"q�N�!r$0QR�&z�}��T��a��W(x�]���"^���(�ڢFC=�8@��j�g�pQ��G�"�BG"f��lљr�4�ȓ�M�P/W>o���x5�ŕ"��
�''�#r?B��K���a���
�'\�P��mɀ)%�;���
�'�����X�v\�[4	=oH`	�'�����U(���i˺	0����'4Z��[1����p �YL����� E�����Y0�)�J�iw�!q"O�q�ʇ�gs܁�˓�*I!�"O�Y�6���I	@�R�`M�"O���# R	
R��0K�B���t"O:�!ck�a��L`Æ�'��xi��'��'&B�'�R�'r2�'��'u��W)��C�5@��J�L��'��'*��'���'�r�'���'���L�1d���XC��qՊH���'���'���':��'�"�'p��']�e���nA(\�ƪ�u��Y��'�"�'���'|R�'���'��'�����M�	`���r��k��y:E�'��'j��'���''��'��'h���@0
����V�V)qJ ��']R�'���'m��'rr�'z��'MD� �^9D��8R/�)'M���g�'4B�'�B�'|b�'"�'���'Q�����Eg�j��4@�(��4�'���'���'u��'$��'���'�ژ��-���J�_���ze�'��'���'M��'J��'��'�\];���u�eナ�'-����c�'u"�'�B�'/B�'�r�'�2�'��+I��``I ��7Ȱ5�#�'}��'��'��':b�'R�'�ʱSA��,ol`�2oH�=�����'�'�r�'Y��'zr�'�B�'�J�-9	⬱B�W&S���A��'�B�'�'K�'���w�
���O��[�G���"�|�2�:��ay��'~�)�3?A��i�BU�e���Z0d8!`%֘ Bh��������?��<A�M�	S^`aCN�#s�RI ��/�?��:u�\��4��dz>���'���5!]ZA�0��~���mS�`bc���	ly�
ff�ZF��Jo����&44,�ߴ>�*e�<I���'i����!T�(�+6��q�'�4s�n���Ox�g}���M��3W�V<O
P��dٳ2w6�a ��>
t�-�5O�牛�?�@':��|"�Ql�,°a��A���Bq� 5t0͓��$%��F˦M���7�I�(��9��������ߦP����?�X�������������glJ�
0�H\�Ũ'ʗ"h���l���^"#Exb>m���'Dx��	�Lxf��+P�N��dr�h\�$�Jt�'L�	��"~Γ��Gf��F.�9��f?i:�ϓjR��偫��$�ϦQ�?ͧL�|hh��v��$��hb�FAϓ�?i���?ib+���Ms�OB��+���L�f��:�=R�Uj�dKFUO���|z���?���?����t�'��)O�X���g ��(Ob�o�t�,�	������?}$?岁	G#��`d��]iH���KĖ���C���ݴ:������O;�$/C�Ty�����Ս@�`Ԡ�ݗ|\�h �ih�˓2�u 󊦟�&���'�]���ȈW���c��:��8�'���'�"���\���41
<��_P��n��m��Qt�!+=��������x}��p����IԦ�"Ջ�9؜sW�Lu�Ը��L&�oN~r㊍3�N���6��O�fT�E:<�$�N3�N]�����y�'�b�'��'V"�i\�j�0���I;t�:��b����O��d�즵`�gl>��I+�M�����6�3Q�\0j�.�n�:WN�$�� ڴz뛦�O�Θ��i��d�OB�w���V�`��$�[8��$��lP�`h>LH�'��'�	����t�	�]�D��P�f
!���<I��	ȟ��'�6-t#H�D�O����|���}*dt:u��'eP$`t.~~RĮ>ac�i��6-�J�)Rт	����kb�]�g��,#To�-<a/�?�MqX��xm��9�D�&6"q���39��°		9.���O
���O���ɷ<���ij���lѧ�r�˱��?��Hq!
.,�b�'�7M1�����$v�~��'-�Q����Ty�T�@����ܴ<,D8޴���H'D�U��O/�	�R�>���LD6I�бʗ�M��	Oy��'B�'}��'|bW>���h�=0�j��-j�~��o���M�kM��?����?1K~���w$�Ҥ	Ͽ5�`R�H?��<YFfoӴ�mڳ��S�''���ش�yR��7�!be+6Np��p���ybA�V�@q�����d�O��әBIL����i�������)K����O�$ca �O��m؛��?|��'��*
>?�J��>dд���ٯ��S�������ē��9k�4�?�)O���F�GuhB�f��,v~ũ�:O��D�&?h�0���LF����?�y��'��9���v���kD�)��Q��6Z�8�	����	ݟ\��J�O���<Ab�41f���i�w�����$l�I�c�<���iM�O��3BS,�����a:��3�N�&5�dxӔ m���MK�`ͅ�M;�'%�wk4��'-oj��BՏir��H�ќt�NԛH>i/O$�d�O �$�OT���O��$_�NB��!L@��t;dϲ<q �iA�M1K����'*��֟���'���e��N�Z��'c�@D�i��>Q��i��6��Oܝ&>��Sߟ�PcŅ�l,���B�zv�IR.Z�<Ϝ4�V ?y�d�z��������dV3oU�HH�`�	x�ܩ:LT��$�$�OPa{��G>�4������q�;k�Ԍ���4�d���D	�0pG)�!'`�Q�9A���X}��'���}��2�iϜw�v���.� �81G�Z,8�P7�u�h�	3�a 5֟���*�{�? ���gcD6I�HHI�I�*!�F7OD�$�O��d�O����OZ���$'�n��D�%-�(�x�M |m,�u��Oj��Ʀ�@B�MBy�'��'k�TF�U���Ր2���B�a���7��6�q��	M{(,6�}�$x�fK�0���ô"�x�&��&B!���)M�M�0T��N��h�Kj��?9��?���t�}��ÍEO�����A��q���?)-OX�n�%�<5��蟸�I�?���-$p�1���a{5��62�����D�'aҴi�D6*�S7Z^�@��Ɋg��4�CDN�;��`���Մd��y�&?�f��h(#0�m��`��?ͻ��ו�-Z@OC$|��x�&��Ɵ����8�I͟L{� p>-�	iy�p�]x�o2>�,�qT�I]����h��t�ܟ�����\�������[��a�f� ���-�b�EIXw2li�`m�Ϧmsܴ6I2D;�4��ě�&�&� ����SR�h8B�cY���Fȁ-iLz=)�4����O���O|�D�O����|ڠ�ܲ��圳M>I�sh��9�X��ݴW��e`!O��?Q��2U��?�'�?�;.	4������sw��	F��(�:aⰰi�26]ݦ����O�`�v�i���}��2Um@�EP�$�v�����,X�H�h�d�Z�c��R���۟��wC:x���,��.�qA����|��럄�I]y�x���d�O����O�p���:����-@�K^��f�O�˓�?��O��$h�lody��Ee�(Q��5��y"�����j���� G�F_����u�FM��P���'^�\��I�,�\],B��D�tg˝�?���?����?�����'\2�ޱc~���"H�#����@�+CREz�� �g��O���O���<��Cs�Jw j�y2BU	To���aT?ٴ �v�mӪ}�d����ӟ�j����Ĥ�nzd8�Յ�Npt���bJ�r�\$�'9<7�<ͧ�?���?���?yW"Q(�u�Ҋ�|��\i�m�����榡��ʃ���̟|�OB�'���CDX�A����!��)�1@X�X�4	w���~�
����	�B����T����Kw��j'�tSAaA��u�@��\�ƣ-2R��Py��{�P�1q�Q�K�;r���`,Ǖ9=�H���?i���?�$�VA�6�)(O4�o�:f���S�J"�"q�߻#�6�a$@M�:|�ɽ�M[����O`��'���i#.7m�	���fY�=��[G��#5E� q��r�t���$xćH����-?���n'֍Z�LNbi~%t��l@�D�O����O���O��+��H7�LI+bOF&<��geahj|	E�H����Or�l�j�'���'=�	�8[��*	U���h&�@ `� <�۴��$|�!Dx��R�6m"?)���:�����ag�`Dj�?��m���O�q.OT�n�Uyʟ���A�3�g2�!�B��"<Y2�i��Q���'v��'m�2Q����D!��At��<���G��̟(�I���S�D@��u��,ФE=
gIG�Z�lG)����<ͧk8��	O�	(��%�V��=hv�iѕ��q*N�������ß��)�SGy��c���1�πF+���WKR�b}��"������O� nZt��L���Ŧ1�!d�!u������C���"��?YߴI��t��4���к�����$v�˓l�,hs J�mi,�y��g�P�͓����O��d�Oj��O����|�q����`)Z�(Ҟ_U�h!!��a��䐧E���'/ғ��'�7=�8<B��M1K�P)�� E�m�ń��=!�����|�����5�Ɍ�MØ'2�LS�1��`�㚘z�Y�'���J�˟��1�|�Z����ß<qKS�t��	!F��L�:���NX�� �	ԟ���^y��{���Rf�O����O����P�?BP��%�/�X�>�I ���O���1�d�hb؝��-��M��a㎛ a���O.�Z��+(�&	@Vj�<���O���DX)�?�4�67��2�"�4/���C�/ɟ�?���?i��?Q��I�O���#X�$F��b��d˗��Ot4lڥ\�����ܟ� �4���y���x����ABJ�,
V<{5���~��i?�6m�ʦ��p �榑��?A��ޫLD��)	<
쀡�t��'
����R#$p���J>�.O����O|�d�O��$�O���BO�r���:��]�tw:�Iϼ<��i�ɲ��'�2�'t��yR$w���GF�¤������(��Fl�F�&���?����6}d��.��v	��D�	;��b��H��59(O�HH�W+�~�|�[���q��3`,��'��cC∫�ƚ�4�	����I��Siy,~�zةq��O��%l@�$d:�+N1�Q2T��O�Ql�F�5����M�Q�i�7��=�] �%ڪ$Gة �G�a�B��q��"$J5�?e&?��]91@Z�jr��
�]g((X�9O"���O��$�O����OL�?�fG߆|��+7�� YVџT���@��4<$Χ�?��iS�'��pf�0�`4�dC�1*d��.��Ʀݚٴ���NB��M{�'�b�N47�Y�����pȬ[3,ڣ��5M�T?�I>�.Op���O\���O)�GV��L�@lD�\�eJ�O*���<�i��*�'	��'�Sy��j!E��|��`�7� ���	)�M�5�i�XO���$2˔?_qR��W&�f�x��H�H��eF�o�b�'C�d�q?AN>9��t}���e�m\`	���`<A��i�l���k7%k �1�a�>IV���J=���'��7(�I���d�O��� ̝4h<!c&���BA��O��m����m�w~�N4��%����� �Z�H�SsRl�@��h �(9O�ʓ�?Y���?Q���?��򉃳t�JH+%�7"@%�q�L(�f�oZ��f�'j���ܦ�ݛX�N�SQh�1����E	ן+L=�	Ɵ�K<ͧ�?��'�>aK�4�ykT�$T(�X��%��	�����yb��ue�l������O��D�^�ʹ�RE
��r<���%hn2�$�O����Oj�C؛�hq�Iş8�ֆ�0/.t�RR�//\حhDO�'�$c�O���O|}%��Z�LL9s	BY0�Q�N
a�e�������jBwQR��<��'_nJ�I��b�
0Pj�K3�ϛN'n��A� ß<�����I��PE�T�'�0a�&��W�H��I�0f�|��'�7ٺt6�����4� ����A��I��	��U�77O����O��l��A�~ o�g~Ҥ��u���'`�	!cJ<)��	)�KN4��TIL>!-O���O����O,�d�O�!�ǋ.c<A�T�Aú�Rb��<�e�i@�X��'��'��:��C��):�q���p�4�82��B}��'6��&�󩘖b�qs�B�f_Z�:��č_�����v�z`�'%n�S��_l?�H>�*O����%[z@Q���	N�.�:`m�O`�$�O����O�ɱ<'�i��p���'�!�L3C�5�%�
C[|�W�'��6�(�	���DP����4�6�	g
U
�d� E����S���o?&�ZѳiU�D�OX���MS���tP���S��	��L�O����C��N��y���I��	����p��W��,`2�AB�ǙGO�`�E���$�OJ�m��I)\��֟�*�4��l��y�C@��aj�m!e@�R�&��V�xB�`�ʽnz>H! �=�'݈���]8� �YƍE3?�I3b�S0�ҥ�������OZ�D�O��DT"��Tif�ށ@��4�U�Rl���O�˓A��fL�d{�'��Z>�X�N�Y�9�Ck	j�!5�"?)eX��+�4Tꛖ�$�4�l�I�-�<A��2�VɁ��>}1<�A䎞�z(r7��xy��O�����[I�	Z��ހ.��[S+C�n9+��?!(OB��<���i��t��ʊ!Q��A���T�;w)���r�'k�6�;�I����즍�b�P*D��`�pX��DG��M���i�豓Ѽix�d�O^%bA�۬��dR���G�8�* [�$�=3@T��kx�T�'�B�'�B�'�r�' ��`���	I��bR�K�>� ش��A��?9����'�?aw��yעܦ(B<X�F�P4"�$�� J-���c�.&���ZM���Ӥ�	�F�3��N �G�)+��?�P(�$�OܓO�ʓ�?q���\-�q횁0P�vH�Wv�m@��?����?�-O��o�
pM*%�	��.U����j�#��)Dǆ�a� ��?�&^������!L<�Ѐ˶p��@���ϙ�V ��~~b�	�3�e�i�����	��'�W�+�|��M�b�N4��%�S���'��'�����3
�� ��H��)g|�#7��ȟ,�ٴyt��?A��i�"�|�w�.l�C����q�̍�b�YC�'26��ܦz�4�\:�4�y��'��p)f��tv��t�d�e�C>v��R�H߅�����OV��OX�d�O��\�x]�m���
����d!���P����)$w���,&?�I&c��ч!Fu�؁9"��~hn�I(O���h�"�'����lJD�>h'.� �D=r�FA�u�ԸO�6m�wyb
Қ��m�����D�>D��$-l��ى��?B�|���O��$�O*�4���C@�V�ǷS��/�p�r���<U�N�bd�Ü�y�&s���0�-OJ��c�:�lڥw0�x�fO~�\܁��P5k�BC������'0����M�J~��� ���V�R�&&+2
]R����?9��?���?!���OW��Iq��*a�NŃe���.�A�'#R�'�6�B"�)�OxnZ~�I�:oJ�(M��)K:P`�����]�I��@�i>�r�Ϧ-�'>��(e�_���J�哶M�-�#��������D\�'��i>1��ݟ��I�7�칷'	$Z5�*���40��Ο�'�R6ǇI~���O����|j��'�i��L|�9�V(K~���<!��?H>�O���J ^����ѓ72hx���>
�`	H0.Z	F��i>ћ��'/E'��0��6IK �J��L����!�ٟx�I������擖6���Iy��f�R�aU#���p�0#�&dQ�
I	@4f�$�O��l�Ɵ$�����>Is�i���F�7f�d�q���l�p8��yӦ�$�� *�6�q����]ȚA�Q�O���`ƹ�U�\:Rq���d�.�]͓����O����O����OJ�$�|:3��%P��LbD#'�2��$��DIN�ݘ��'��O����'C�$p���_2L��1��	B�a�kS
�5o�> o��M����4��	�OV4k�y���ɹ���P��#7�F9)0"Φ*��<bR��O�lI>i*O�	�O��/�P�)N6"]��zV�W<2����O����O0�LV�&�G.Q��'^��>=�8�3�M=y� }A�'޺��O4A�'�2�'�Ot� ���m�9Y"잩��cԝ��s�@-eK�lZ���'Vɜ�	���q�h�_�*��V�4P��r���ҟ��	�����4E���'ߔq����8ެ�U������1�'9�7��"?�����Oz�oZM�Ӽ�Ҡg\�}3�D
�VA"}8q���<q��?y�is��¸iH�I+ �>�  ӟ� f�U���
[�ѴK�D�gA?��<����?���?���?��hʨW1d�QD����Â�H��d�ܦ�h�ן�	��$?�	�{�Y'�+/y��T&���PX��O�}m���?I<�|:�!�1�`dD l�ޡ	&IͦFv���	���d�$(���E�8�O
ʓe�J=�U��W�<h9�O�&G���{���?q���?y��|�,O�=o�	��=�I*~���çV�P �l�wT6V���	�M��b�>����?Yտi�t�z��N�T� �ň�;�؄�E!� tϛ����cSf�����:����p�wIßWR⽐��ҍ1l4Ɋ�'��'�"�'2�'���ec��������m��@Q*�Ѐ	�<������^���d�'��6� ��_+xb��
�C�<8�<}�2n4:���&���ڴћ�O����b�i��I�V"���"斃2��]�7C�VeX͘�#�;-f��+���<����?!���?Dm£S�6��ro��F�����R��?�����$�צ̀����<����O����&j�
�(���6���Oj��'K46-��IkN<�O� ��c���*�n�{cC�9�Y���<v=� �i;���| k���$����cܤ��W�P��L�3�ޟ,��˟�����b>��' �7��
t7*�HA�g~��Qu�N:�\��e#�Ob��Ԧ��?m�>q��i���{w��/ ��Pˉ�$bEz�l~�HTm�z2�x���U� ����?��'�T�ץ�>b�ظ�0$�*��8Q�'Y�Пl�����I��p��d�$@ڶ����|a�� ��8-�7�K�A��d�O�D!�9O�nz�� [=9B��	ufް	2�RAɁ�?��4�?�O�O���Q�i�dO0_*S#�R+Ov��� �<^���1>�f���D��Ol��|��%�:x�w'�3*�j���y
����?���?�.O�m5H����I����ɇOk�
?���r�ݑ}U�����j}B�'���=�d7+�J�*r��9"����f��X��OF��j�vRQ��`�<	�':'��$�?���X7F���a�5�\��,@)�?���?�����l"!L�j�fa�a$�%�l[�ԟ��46N�����?�%�i��O��<k"����I�>h|� (Ѭ|��$��1����M�r����M��Ox�jh���&�W�05v-sC��s�e[��ȾN,�O�˓�?����?i���?��
�j\0�T�*��\��;s����DO��y���xy��'P��|ꂈ]�o)td UC�K�t���oy��'|J~�5 �"G��r�*�b\40`�4+�T��q�;���ş'в$�e�^�O��Z�f$ӃbJ `���W�js�a����?I��?���|�*O��n����'	ش#�/�]cࡑ���:�0��'�7-,�ɼ��$C������M��#]B�&T
�΁Z���5K ���4��$�.�.����UD���0�.�:��1�`H ~5�A����-e��O����O����O���-�ӰxV2�R�h]90_N���җD�f��韸��4�M[����|*��A��|��Ǯn;�8:���1a��XHtKB�	xO�im��MK�'+���4�yr�'z�`�B�ʌ�↏+R ��sG��I�('�'�ɟ���۟h���
���ŋ�=R9�׎N3B����̟��'�d7틵[n���O��d�|�ˇw��т�'s����~~�+�>���i^27�y�)���˃X�D���M43�̚�k��)?=��NV��M#�R��t���,�d���RX�U��$�Q1
�"sK����OV���O��i�<a�i3�Q���v�~Y�PJ��T�qH>{�"�'L�6�9��+����OD '�ߜg��M2�a�)-��S�b�O��mZ���oZQ~b/Χ}�"���W�	S--�tI���?O�2T0t@4 �$�<���?���?i��?�+�캥
���|I�����mE�a��Z�	ß<$?��I9�Mϻ��,�5m$l�����z{J�� �'қ�-��O����O��$�6�i:���`8�(�B-)f2�8�������&):غ�1騒O<��|���}?:�a���V)��AUc�q_�����?����?�/O` m�&#�P�������iʸ�wF�n���Ɗ&͆��?��Q�������L<a�j���m��,Y��S����-)p�U�[���|�P�O�h��krݙ'�҄)D	�qhZs��+��?��?9����zxx�¸U��;nr���`�������юH�y���M���3�?���?����4��N��Q�&<��V	p�n �1H8w��d^Ӧ8�4�?�B �<�M��'U�X	A�ơ���r���t��}�P�T�M�;��%ƙ|]��S��P����,���@��� ��� �.�.NCǃnyR�n�䨠�Ǽ<����3_�?���.��ZV�9:~�,ڲȕ63o�$�)O��m�>�MK���h�R���*
�5��EI<yP�!��fP��3����#�� ��f@�	Cy��)�^ų/�:��ƭ^M�R�'��'w�*�O�剿�M;ū�&�?9�\r��0a�EVb!�ٓ���?���?).OL��>?���MK�uPځ;'���-&�5�ė7p|@� \��M3�'���hȦ��S���������u�Cm�0Ud�ɧ������O��D�O����O��D3���T�,��@�t3@�'V:���j���I<�M#g@'��dR���Iyy�	DFN��e� �D
G���rT��A�4:��O�\	%�iU���0� �E���].%�LP�B�<Dݞ�)����?���$���<ͧ�?Q���?�2�Z���(���Ew衸!L�'�?Q���?I�h��tZ�tHB�?���?ֳ��4��-������fS���r#)��${}r�'�BJ?�4���d�� 4����o>Z	i���0&_��+@��/_�6MMyy�O�z����Z���hh�
KV�:p둿A��#��?)���?��S�'��D��y����H@bրX�m�8ڇ���]������ߴ��'��#���m0a�� �h���b�.P�6ML��dMRܦ��'g��#��T:+OXu#�l�AE�K�)�a��D��9O���?����?A��?I����i)pG��]F8�SB\3��mrFzӐaX���O@���O�����I���3lJ�xz�nB7:�ި+�� kU���4?n��.��Ɏ�o�6�k���G���.����W@&GnH4�d�d���'	~1�� �Ĭ<)��?�q�%SkX�%��L�&F�B��?���?	����$Zצ��$�\qy��';��څb�$��PC��H�L�X����a}�@q�p5m����a7�1���9�B�&V�_�|�'v���G�<Nw��D1����~2�'��"Td�"�a+�ߞ?���a�'R��'"�'��>U�ɎnK�8��EqOF���b�$��	��M+eh�(�?���l����4��i�E�8t��c�I\� 1�Z0=O^��O��n�[�T�m�<���t�"�HR��t��A��7;5ąR�#
M��R%�D.�䓈�4�~�d�O��d�O��d�vC������/!=��
��{T�q��vW��'�B���'Sޔ1B�ҏOv@9E�7 ��A�˩>���y�x��tb�<����M�`��@��i�b���*F)�]����'��%���'��I{3L06�ꉹ$��[߆�{
�f����/'��FS�b�p��Fe^�Ie.�9l�b�<�p��OJ���O�lnZ%._D-R�a�3miu���!>4*숡�\Ҧ�'������V:L~��;q,V%��E���id%�l ̓��?�� �P݌�9s��(�	2"�!�?��?�#�i6��������%���W#�"	���Rk��^e�<3s��?������l��i9�6�#?���\&􌀹�Ɏ?9���b� ES�չRO���$�T�'7�O����J7�1X1�\��RY���!�MóF��?����?-�v�ZQH�D�]�6`���P,h`�����O�)l��M�ґxʟLl׃�n�,�X +� ݖX�eĆ=���z��%����I�f?L>	4n��	�~x�f�4'�5��U<qU�iw\� �WT���R��.�^�q����b�'��7�6�	���}�j��q��%֦��F��E?�8����ڴjL�%�ش���ДL֔���O%�ɖK��Dd�w ���P�@�o���qy��',hHCW�őA{��Z�/N�ƨH6@`ӊ�� ��O����OJ�?=����!hC�����Ř"<��E.^���Kt�4�%�b>��D�Φ��>��Ö���"b�Q��K�73d�Γn��Xp1����$���''��'��DO�"A�T=��,)�Fu�5�'�r�'��X��cڴ3�FL,O�$"�e��)M(><��n��54⟤9�O@`nZ*�M����d��&V)1���8-�(�n:?\��O΍c�I8�j�;�����S�q>��ܟ�i�E�@�6��G�P�r�(D
џT���X��ş�E�D�'�.)��D� l	�184��/����f�'fh7-�!�"�2��&�4�iSte�e���q�F���$Q�<O�|mZ��Mk��)\�Ѫ۴�����(a��IW��#π'[�0mj�\�X�
(���<ͧ�?	���?���?�t葓�(I��m�(*�>9Cb�&��dO��135�<��ȟx%?�	�R舩Bl��9-
�p�L���p�O��m�3�M+���O}�T�'�4ER�
RL�0�#�/p�3��::p= �O0�F�ȝ�?� d*��<	��V%U[ذ�c':x6,�z�� �?���?	��?�'������
�,�П KtHI,N�����r(,Ui��K��y2�w��⟄�OPnZ�M;�Q�����ΌXg��H2�K�l��+2���M;�O��л�b��d�wm�@Rq�ÛGd�yP��s�x̋�'���'�r�'q��'�p郷*"r����C�
�"��0��O����Oj�nZ:i;d��'�87M&�dB�&���F�*{�Y�n�&Zv&0'�X�I�p���C��oZ�<�����H
BWܨ=KČ�~�R����'Gt���3�䓥�$�O����O����J��pK�d8�26M�5TT��O�ʓVY�&ň.`TR�'�BX>9$�$�KEj��VXXJwC8jO�I����O���~�i>q�	�}-h��/ޏ2�`�j��I��I�w��B��*3�Lyy�O���I62��'NJE ����G��y#�%�l�4pv�'�b�'k���Ot�I��M�i���@%�iQ�hk+[�Z�J{��?�6�ih�Ob��'��7�� x�tC�OR5���z0k؈q��	��m��!�ߦ��'z�IÇ��?��X���Iq�|\�UgM�e@!�wDj���'�"�']��'"�'W�+{�ra86�R��-���kR����4��Q����?����'�?���y�nJ))2a���Ue��Y�(X32
��'ETO1�8d�o`�`�)� ��zW�@=w�P��1
� &/t��v5O
��%�W>�?I�b7���<�'�?�rE��:�$���ab�HpC�ϖ�?���?���������g/Mϟ ��ݟ B�
D�8�2U�����&��e�D
a��]��I���	<��(�вg�&pzi�h-z��!͓�?� '_@�"��4��?mzF�O��d�#^#�T	��P�i1��Ir�@)	��$�O��D�O��4�'�?i�II)h@�ͪ���j�P[ ď=�?�g�i�X�R �'��w����]!�
�`2�˔ �>�{�B�+'�牖�M��i��6M��Z6-*?�熟�rVF�H�Z�qfa��كL��J�X%$�̕'��'��'[�'�h�RY�](�!`A����)6�前�M�3�'T�LB��?��'U3�ub���?a1e�7l$�e	�m4	��0�f��ZW�I �M�s�'������O�����$\m�K�鄉9���I��� ����>��	'qLl���'��x&�h�'��:����`���l�5�BL��]���I����i>e�'��6�\1C^����GŲ�KPƃ� O��aBoRJJ����e�?��^�<��ԟ��ش`Cv�3���B������N5*8h$)�I��M��O������Ĝ�4�wR�}�6��<�)�f�t��p �'2��'xR�'KR�'�,)���J�eI`�g�U6)�P��B�O��$�O �o�{�R�'ic��|�hW�J��Yp�(M1v�ۃ�tO��l��MϧCq�](�4��$ѮW�BDõ�")$��6Łm�T�j� 4�~��|�S�h��ϟ,�I`�D����<��%��	�NZ�	[y҂f���	d��O��d�O�	��T�X�GF.n�F<���XŐ��&��s�O��D�O`�&�������dʛ�[�m"�F��6�P!���U&M�=X%�æY�-O6����~�|"��R�H��/��a'
��T�_�x��b�6(��E�3a��Q����H���aM�P^����O�lm�b�_z��2�M;�o�L�ED�<s�����)ڌs���M~Ӥ,�¬d���l�MUİ?Q�'�����R-\D�a��+J�:"͇�O� �bćO�(q A�5��Z��W'thP�b��:D��ς�[�h,�PɊ*(J��g$�8;
�l�w�	9���"bE�/vR:�cȍk��(�
�%6qhiB�5!9��X��v��S��qo�=d�\$�GA49�"e� k�Y펍�FN@�l8,�3r�U��N�1�m�3x�,�j�B>-�r����4?&� ���"L)��$�n������6ዲA��a��A�>v]@1��>7<�P'�z<�=7�N�H%��B�O<��pdj�,N
$���y���ON�d��`4�'=� ;��Dk��AzF( ��^��)شNRXy������OCB�UF��l!��Zs*�eΘ�f�"7��O����O��R�l�d}�]���	B?1W�J���������ئe'�,3�l�ħ�?���?�R�Y�ک�`�R�lxzq
�B�,]��6�'jD�a�>�-O�D&���h ���ԋojfZ6�(m�4�FT��i4/��\�'��'�bU��p�H ]���D�#��ɀc�l�&��O2��?�L>!���?y2�E��8u��!`A��h��ɷC�X�<����?!�������ΧYX�I+�F��}��(aa�A��n�{yr�'��'#b�'Ĝ �%�O�TD�H)R�2�h�B�%|�z��X�P������TyBcX�EZꧫ?Dm�<$��]�a���9���	4i���'�'7��'�������
�W�X���'��X����r�Q�x���'z[��Z !�����O��$���3��S>j;D�U��m��D%�r�	۟\�	���q�?)�O֘�i�+M���q�+K��Hڴ���Ȕya�Qmɟ��I�\�ӂ���ƪ������>�$hx%�S�V�6��v�i���'�h�ß'��'��>���@3J00qMc8��I����TL���M���?Y����P�t�'��a��a
�+������7�"@YQm|��-�QE2��F���?)0
0n��}���R�ȡaG� fٛ�'tR�'�L@@�>�+O��䤟���JO�bE� �-g2�,��%:��7�Th%��������I�*���cH�5��¦
��dj޴�?i�'�5��	gy��'Hɧ5��_,�$��ɑd8L9%M��dS���O
���OJ�D�<)��A�dR$�I��
�V��Q�ֆ�"5�U���'�"�|b�'���$c�T����&`d���J{�d�u�|��'��'��2]�q��O�.ə@�_?�h��Y����O����O|�O��x��h��,Ԭ�G.�	{`Ґb�E<,�1P���	ޟ��IHy���2�J��+)S*>�>�3��צQڶ�j����e�	G�cyB ���b�~�ֻ���)� \`�:$h������ԟ �'��p��=�I�O����Br���7a�Ј�b���z���x_�p�	���'?�i��ːJU�lA�(��!ļJ8y@�v�P˓ZTQ��i`맡?�����I�ru��;�"��XXP1C�Х'�27��<���?і������4-!6�:Պ\Lx)ʤ���%n�,w�Xy1۴�?����?��'[e����&=���u��TD�S��6��L����O�����<y��$�NP:6��<��-K����X״i���'"m���O�I�O �	%�h�c-^�bt%ҧ��	�@7�O�˓<�iq���䓔?��9�������A"�byX�!�vӔ�D �I��L���P��`M���FS�f�T4¤FD�K�MC�Y��z�ܙJ��c���IRy��'��� 6�Zg�u���G��&U"��@H�(��D�O���+�I֟p�I#%����c���hTxn�%}<��FR3@).b�p�IyB�' Ƒ�Pڟ�$����	)��9���N�|�J�i���'�Ov���O���a��G6�6��	`�@�����U��Hbcj����?-OL��Ư`���'�?	��Vf�p*�Ƕ\H.]��G�WK�����O��DHH֌�B��x�e�@��񐲧��"Oʱ�$���M[����O4m @�|���?��[��;8lN=�"�W�Y�M�K�I��,�I�J2����h2�~2��Ec_�� 7�wD(���n�Ŧ��'���*��}�"Y�O���OA��C�l}Y���4v\$x�f�Ϝ_d%l�m~���?�������4F|<���ϫ1� �@ōDy�b�oڥ�VPcݴ�?)��?��'����\cNpu[BĲg²��3gՏ#H����4O�1���?����?��'�� Zb.�29�PE���Y� ��К��ǁ�MC��?��.-�x'�x�O��O��q&�P(������V���8`�i�rR��H�GHʟ<'���IX?A�M��;�f4�?W	X0��ͦ��ɪ2T��'l�'��'3�{A��kȼ�F)�J��e�$�d��L��	ğ���ϟ,�'��Z��|�҅+4��U1���7O���O�Ĳ<!����Į�.]*� bԨzL�-ڇ�P	�M������O���O\ʓ�Bj�0��)��O\�[��c���J��!P���Iß\��Hy��'��ßt�n��*
ι�r�����KD$������O��d�O��~�x�cR?��ɒ*����ׅHmH}p�#N&Ei�$��4�?!(O0��O��d�����3}�Ï&┓�(NLGV�@ ɝ�M���?�)O��r�G�S��':��Oj����M��t�r��Uw��q��>1��?��R		�����Tg��	��lڀM��j��RŬ�?�M[(O���Dꦉ����h���?aS�O�.�4CW���ФZ�`�f�/�v�'��G��y��|b��uQt���M����䬝�盶oFY�T7M�O(�D�Of��Aj}�Y�H���I�T 0ĊU�� ����M�g��<�����.��ȟ��jQ�s*����
#U���J�R���O����O��E�_f}�V�<��{?Q�꜄}��]�$ĕ�aGȁa�mQ䦑��}y2���yʟ.���O��Ĝ<�|Q; +�<p
v]��ɐ:Q���o���4k���$�<�����Ok�D6&����F�J|��1�AU�&�'�2��'6��'u��'�rS������o��F�1ke)4a���O˓�?�.O���O`������%��(P�1�&�&K����8O�ʓ�?���?+OR�(6@��|J�$�%\}��BO1�F�� ��I�'S�L�	ڟ`�ɥgrr��%K�\ѠE�3�bYn�JuP����i@r�'���'s��`�����$�����U�"��SB+Z-Zf�oZ���'�"�'����yb�'0�$��x� �@	8���4(�ܛ��'W���%�?��)�O*�$�7@�3���r�սwD�����l}��'���'�V���'��s���'S�b|���u&�'M�<o�mnLy��ΩiQ�7�Ov���O��)�|}Zw���E��#{Zͨ�OԨ7���4�?	��y��9ϓw��s���}*���b�����D�'��A������hfi�*�M���?����rX���'��DX��@�����tp��@�@��v���y�|��	�O���dʝ�~�f��$(�H@���U�E������ ��I�X��Of��?)�O�L�����A�c��?�8���4�?A+O�X��6O���� ��ݟH�r)�-5 ek����8�K��M��H��4��P��'�R\���i���#�)3������%jN.8���c�h��&Y��<���?Y���d�s�\���� ��$Sc���B��e��Jh}�V���IQy��'\"�'��p	���;_T�u�Ԁs3/�:W�D��?����?���?�*O�DR�Έ�|R�Cڼ$�NԀu�_'�P��sk@��i�'��S�l��ɟt�	M���	�y8 �zO��@D��	G�T�n���B޴�?9��?������Ҹ��O�Zc�b�{5����m*f,i5Px�ش�?a+Oj���O�D�<(�1��F3�U�߀g:x	*�o�<�M#��?(Ođ9�[G���'���O$<�a��3n�,9Z3L�<pbY��l�>���?���(�͓��$�O���'+�Y�I�>�j��rK82�7m�<Q"�M1�v�'���'���N�>�;n���ò�>S!J� R�n���x�ɕ_���	����O8�>}:��P�hʪ�Y���|�u��~Ӷ�3M���-�	ݟp���?)��O��9��({g$�5J�0Y`��"<�H��D�i?&L����=�S�h3��ӟ36\��D"�"߽�M����?���1#��{�R�\�'��O`�s'ƞ�(1���EDE�l��)�Ծi�2U��+��a��'�?���?y'f�:{�B=I7(=��d̾-����'�F����>�*O�$�<���[b���8����h�F-Y#��Q}r-��yRZ�T�I��L�	iyB �$s�$	elr����F�ŘB.I�h�>a,OF��<i���?��.���T�����+�/ `�����<!��?���?!����E�1-�xϧ7f��@@�'�T�2� 2,�o�Ny��'�Ο��ҟ�z��a��8�9	| 9���/Q�h<��b���$�O���O��0�ּ�Z?e��9�� � jՄC.0*���dA6o�"d�t�i�2W�|�I�4�ɀ_����v��K�[�pi����cL���$͎��'�BP���� �����O~��Nŋ#bݑi��"o�����u}��'���'Dhųʟ0����+��;���Ղ��H�*���M�.O44Y�EWȦ��������?	�O뎚�T��Q�ĭ�/B��j�ៀ����'��τ�yB�'���'q��=��%��-3z,����'$��F�i�ph�3f�����O������'%��;-�����=��K���6����4|��`��?�.O��?�Ipƌ ���/k��e�P�[��� 2۴�?���?	U�\8e��oy�'c��C�3x�f�A�$� ��Qd�"CR���|�(�yʟ���O����Uڨy��8Uj�{1� Q@(m۟ B �J3���<I���$�Ok,=�i�Ѧ��A��h �#�-�	~���	؟���ߟx�	Ꞔ�':�t��(�2 �@��VS�E?*s�O&���OĒO$���O�42��T�v�y�SY4�m)�g�J�L�O��d�O�Ĩ<�U��+�	�	�z8�/�t��\�KW:z���� ��a���$��y�p��Zh*B�ο\��:���U'���'r��'��]�܈�����ħ�\D�F�{�B%sPf�	"t$��i\r�|��']���yR�>1�ґ^^<��Y�J2�hXb�����I؟$�'�R �Շ(�	�O2���IR�%3�D����|��BT�*�Ĩ$�p��蟸Q�D���$���'H�J-1V��6	����2Ryliy��� j�7M�G���'��$I;?!�G@"d�� ��&J����,ɦ�I؟�u�ߟ�'���}rW����CsI�#��(�����R'��M��?�����xr�'��,����%,����#Y(��Ox��(�%6��F�'�?yPO�uKl��c�8B� i�rb��)ћ��'R�'�b�Q�J:�	����]�z �`��P��&���%�0��>���Qa��?���?� X	?\�{��'f�@��Њ	�ݛ��'O�8�D�4��˟��'8Zc��h�	X;�x���? �-��OQ�#��Ob�$�Oʓa{n�"�Y29��`�7e��Ey���Ƌ�]!�'�2�'��'�"�'+�-�W��Sq���1�~u��+ˊ�y�P���I���ICy'�XS��R�Yz@�оp"�c%n�"SӒO"�d>���O ��*!����8<����㊪/��!�r#�}����'P2�'��]���'C߉��'n���pd�α �|ס?ހ�Ҹi��|"�'����u��>�1͛b`y�.�*�����m��ş��'Q�U�f�(�)�O�ə�'��EؠQ��)�:
�=	�i;��O��������;���?sAb�1���1��MG�P�ՠm�Jʓ>7ȼ`��i8���?i�':i�I�kE��g�+Do�m��">z�6��O.�dҾ0P�/��-�S���"�_�l�"��S�P;N7
6G�kS��oZ��I͟@�S����|��	b�=2��n�R���[���N]<a��'��)�'�?�"�ׇ� D!��°�B�I�7AN���'���'���ꦦ)�4���'O8h c�d�zdA�@ѝ�ҥi�4�?�)O�e�ЈFS��۟0�	ßl �+����	S��R����Ѩ.�M�%�\���x�OkQ�P�3%�1Tt9��D�g���0��>��
<�?q��?1��?�����d�?;�8�i	/us�U8b$D�8i9�cSs�	ޟtG{��' ^l��I��:���cG <�b�8�G<���'��'�"�'���	_A��O�|��AɅ*p"�u&Ǒ+�A��O���(ړ�?Y�-б�?釣ÃYX�TC��wu��"R�I�����ꟴ���`hU$S����	ʟ��B,Q���1��3&�pK����M������?���)��m�1��q�4mMR�p�O*">�XT�3y�J6M�O��Ģ<��ڶR*�S����	�?�Ig�<Z����C_�Q�*х���M���lR�5��On���^	��7��Q��ZF�f]���i���'��`�'���'k2�O��i�q�T��hU���L�(趭S�j�H���O�<��	
51O���y෫�(^�,u��ǟ�Z`���iM| E�'u��'4��O�B�',��]��P���������
���P��4d�N�:��O�S�O��߄մuQW�2.$�������6��O���OTM`��BB�i>)�	����F"�1d�#���v���GM����'J��y2�'��'�V|2GC�<7|��W��#T���lp����ԮH�N�f�����&���P�T�}�(Q��A�>K4���,����Dr�Yv����	�����qy��_l��(Bâ	����D�ڕ�� ��g)���O���-���O���I�I3p��f4N,5#fO5j������O��D�OT�4�
a�5:�������t�hD���&�%����ē�?�N>A��?�2�L}�,����S(.x�Uf���$�O�$�O�˓H�yJ��TF&%&��4���)�:Y�	��u�\7��O �O����O樨��đ�}��@���24�e�ݔ)����' �P�X�m���'�?���u�Q�� �0$���b��nR����x��'����O�$���Ϻ@-2��ӣK.	��7��<���M�g^�6;~����ѕ�� �� 3�T~��kQ�(>�%�F�ia��'c\�ʌ��)�2h�.x�5�F3P��#�^.��h��G�7��O����O����|�H�(���e+, �8�d��q$�q�i��-���d.�S؟���AM:/w$�4G�8!����u�&�Mk��?��a���S�D�O����^6�=צ��4/\����% $c�dCU�#��۟��	���pgi1oZ��Q�_0��m�j���M+� -���Q�$�OT�Ok�$[� ���,G5!4�8���&���S1�c���I֟���ayb��/~*��$ �u�؂ G�49ָ�7�"�D�O��d<�d�O��$�- )X�ýB)�&�8��ԫ����'���'""[�h#�OP����$,��p���kS���o2��d�O�d*�D�O�җc��I+.���
z�x�D\?O28��?9���?�)O�ԘQ��\���'.���G�(��k1��>,s���E/vӾ��<����?���;p��?��'`8&H	�+A��r&L,si�Cڴ�?������ſ�\ �O>�'��dm���7��"=V�$f;kB��?����?�efD@~RU���86:p�s$Ftb4�Ii͵�J�oGy����HԨ7��O(��O����u}Zw%�,0''¬�ҥ��#@�][hEp�4�?��[�:1̓
.�s���}*�-�=K\\�C'K�:����G*����T�K��Mc���?A��j'^�L�'��iNڝQ�ˇJ�!Ȃy���hӴ@g8OR�$�<��D�'���$��1z ��+�+���Ƅe���D�Ox�d�R�h��'1�ğ��ZZ����]PN��"h��% \�>���ZS��?1���?�g�ȦJ� �b�/����Eʵf��F�'d>i��>�)O
���<�������Qh��A^,2���E�CO}������O����O���<a�%�oն���C[���H�^�H�1a]���'�RS���	�����kL���)J�:dG�Ύ�Ь�g�$�	Ɵ�IߟX�	By���4è�.?^l�s�ٿR�}��B�4I(�6��<�����O��D�O�٠�:O`�h�F�,+JH�5K��Y��&Sj}��'UB�'��I8�d�í� �d>?���Ђ�N�$�"�`���">��n�ʟ��'�'*r'Ʃ�yrP>7-Mg��xR� z�0���`+(D��fU���)T��I�@,X�#�Tu����%z��ɬf5btH�� ��TC�I g���c J.�R���_$�˗�QV�X]���u�X�E�GȂ�_J�A���N��!��V�d�T�[䇗#8pX����.�|���A�Hܠ�#@ ˲�B�I�f�<n��d*���9�|�`��B^#'I�\��Ic�b��H'�����#����8 �7E�Q�pP�Q� 0�,YB�c��
Sd��O����Oɬ;/�<��FS���\����*y(���GI�����Θ-��x�ba����O�f�'��q� -�NRQX��Z��Hұ�/+� ���4�����9�.��3J�|�0 X��4�ݴr��B ��1W����B:����a~b,��?�'�hOR�㧣�-Q�|�q��.o@�8A"O����������,X]r��<���?і'�,�Z����,Y6�ې́�{-��6Lٙas&mʒ�'�B�'���`�a������'Mn�2ӊ��W�|er���p��+����X�Hvl>`9@9ϓ,��$�e��d0q��"Q��x�V�X?V xC�	`�+�[<VP��m~�cA��-Jq��)��̟���r�'��O�%`�,ι(Tܰ�B׸X�0hA"O���sM3%B6�{3B'N�F��e}�_�tB�	����$�O����4��Ei₄0'�mz���O����1X.j�D�O�擠 ����`)7�V�s�'82�Q�j��H|�� ��ݕs|���	Ǔa��U0���DwTu���O��I�Aj��0�#Rȴ]���'%�!���?A/O��6�� 8D��r���&�4����'|OTmˤ쑖�XJ��<5�L��eO��lڗ@@�l2�F�V'����F`R �`y¯Z B���?�(��Xy��O��� ł
Mx|��",ߝ3
i���O����;� aH cX#hX��O�a��i�#_�Ԓt��*��� C����	�V!L]�BdY H�ra�Gn��?Y8���Qp\T��I;z;����>}�K��?���h� ��&BJdf�N�GK���Ь�:)�!���(<�H�+�:f����e���axR�5ғO?��ې�~�dq R�V��.���[�����<A��ˡT<�-�I����I͟�ݓn�b����(T � �3Wy����O%�I�2DL�@�)�3�$���`:��(%$�RS�|��Hq�=3}@�!q� 1E������]��剶H\���#��E�Ä8�̡��q~R���?�'�hON%�MX�G"�x��3 1��"O>LrwD�Ce0@�F���h�F<ّ���{���?�'����u��3�2苰�D�����/��~�� 2c�'���'��y���	��d�'�"J����n$Jt�@�$_��N׹4�����Ј
�H�Dy^}�Q,�w�
)�$�� �`����`X@7iÞJ�[t+T%jx�Q�ɘğd��)� ��)��E�vo�!�$�'[��$e"O}��M0I8�r��;B^�b�dD�]�,+�i�B�'�R��`�~'V���O�t�z�B�'�m��A �'��H��|r$Q�?RB�*T�T�	Ɗ�����p<1G-]D�YR��(���9���Z,xv���S�x1��[�	���bG�T�K����D��JC�I*�@k�Iy{�����$3�2C����M�"Q+� �$m͐l����,���VW���i��'�哐88��	 /���1DG�z��M��`ӟ|R�)�	ǟ<��ԍfvE�$�����|�+�A[����L�����1��>���NA�ab`�v����'I3$�Hf��s��$��ؠT���'�P1i�ɘ��O=�QT�(���#�B��U����'��@%����C��y���Ó�X��Wm���v(�x��릋��M��?��S!T�q怯�?���?��Ӽ�-�[rlV�r������+0z�
P�;O���Ӻ	������|�O�H��:d�ñDЪ%
��*�x����z���̶lƠ骋�L>�2b
�c8̝���ŠN���c�$��'���S�g�I�#4�� T4)/$Tp�A��8B�	/p*�s7��;9�X]�6B���@����"|2 O:NF�;B�Y?y�Bx��`�9�Ys'�;�?q���?��M���OH��v>1��R�O+ - N߶j�.�PĬ���C��'xGXD�q��MN��6dH�L#l*�)�X�q�]�}Рq"�ˠ9,��&݋<���(�O��8���:.���@ړP�Z-s�"O��P1�EL��b4H�Z��0�q�Ni�(}�C�ivB�'�ֈB풴	�>P���R5K�x�@�'���ոlw��'��	Z�?b�|�e�.mB���%�NQhG��p<1��O��FB!;c�?cY�9�&�ӓB�@�㉍����9�Dİ?�<����J��M!�>]�!�D:{\Pc1�ϸA�F,*���6!�!���q��M�<D�x}��O!9P��N&�I&l���4�?����)�2����"A0���Ơ�2�P�s�P2�d�O�%���O�b��g~"�UJ��qR2�ʮ���$呐��m{�"<����kLLc�{��yY��T�DF6a�'��O��O�ư@��^�p/�\A�%Ä9gTH2�y��'k�y��I�z�JQ�X
��Ց!���0<�!��c��@q��A�F�)�$"�z�8޴�?Y���?9R/��cv�I���?����?�;un)!�o�7<,�[��֓!TB�Z�y�ۈ��<	�l�r\䀐F�[!^R�b�fܓ)��9�牔1@"`:�m>�x3��[�(�0��<	��[��>�O��t'�'*�05�� ë)����"O��9����U8�i�¨_76d������(���Ӕn9��Z�)³g��MgƒM����޹8m"�	ʟ��I՟�R_w�R�' �i�L���Ѷ���C����D'@FHGL����$M�{ r�
$�V'Y�jCk��]��"�ɦa���䉦aEn��� `�:��B�T-~��Ȉ2�'���'�B[��	y�s����&C�?ynv\�'g�4�<���e���@%L"h�{k�3k���<��T� �'Uf�#V�iӺ���O���*3i�Ջ�#P6���h#E�O���Fc9�$�O$�ӻ�A���
&�pa�'
1q3i�y��h�`D `8��z
�z>5;����"�e�%�O��K4`��$R@���;�-@T�'�z�h����	Fd]��a>��L0�>����(?
� ���|�ԡ��ϒ)oYn����W���,U�@�j h��)�'ǘ'��\p�	zӎ�$�O�ʧ1a�82�"��7��Q��y�R�J>HI�����?�UL���?��y*��	0\��5���,���#Q�ܫW���'\�b���	\���B2d�c�����>1��A�S��_�<� D���4-��_�2ͬ ��X�{�!.N^�B�I��l+>Y��	<�HOf�Z��\���RC�1HR��a��Q�	ܟ��ɅA,(,���O՟ ��Ɵ�i�{Em^DJ4�R@�L�P��D����a.M�q1�$���;��L>���>;Jxp��N�U���Ş�g���PE��A�4XYEEöc] ��}&����Bҙ&$�G�C�[������g�X����)�3���	S�ap�a�F/:�q�n�!�� �m�ʮ����7d�	�ɲ��02��4�4�O*�ǧ�W�����D��� �+&A8v�ˢ��O����O2��ݺ3��?1�O��h8BEܕ^6�tpa��`=�T"��x2�ю�����R@`Kօ��`yT9�'��Z�OY.|%j�e��5�;�I���?��SDV���Cr�je���P/����ȓ3�N��`ۼ!�XMbD#07�b��<���DU��(oZٟT�I+q��(�AȤ5�aI#�$zd��Ɵ���%�ԟd�I�|ʳ�e57M*����BL�rD]qyq��*R�&�xB�
��'��ms�lX�<��R��%�����b��h�Iz�ɮ(� "S�[�d_��P�-�-?
B�	�I��fI7�fX3�舲u��C�� �M�qb�-h�x���@H�@5#�v̓;ݞl +O����|�5$�6�?�q���5P�1�P�ũ@i�%�W����?Y�g� S��ԋj]V���kEN?�O��s�E2��H�Yi8�ѧ��<?"�'��C @�,M1����`�O@�<���Z!����U�<��2�.}'�?9V�i��"}��'2�$49��� �pțE*U�1�'M����ő�}�呫;ռ�s	ÓPq��H�� $X�P�:Ec� iX΀�)��M����?��,lSa�&�?����?A�i��T��и���	��ᓠ��Jc���P&*<O0�2LC ���E�n0¨9B���,.�yR�_��Y���O�5��JO�/$1O�%�������6pȒ@�9`�*����(RrT�� V�X����'�P�i�؍{�8��'�<"=E���W{�l.��S*�5^a���p@V1u~���'�"�'�a�i�I��̧z��y��U�\�n�W�N�'m��g�@F<A3�?>����gO�M�i@����m���=���3$CR�t9P�R4�I)x�X}�A ��P��	/��8��L]:��Y�ćК��C��f���BGU)"�x#7K �bc��؈}�
L$O?46M�O������F�X�����A�(|�n���Ox4���O���j>���O�OH5��a�d��Ñ�׵o{n0���'[L[�B�?e�<c1FQ��*	�c@�
�p<�`��ٟ�&�$��X��0� 4A���r�3D�|��"\9J�P�{UNۥ!3D #e�0��ܴ%4�Q�L�'A\={�M� ��<7�@L����'*�\>�sc�џ`�4��1��@�(��f��]c�!Kş8�	�x��	
Ŋ����S�d]>�����"Y����҉�4l&}"�/Hf��P�|��4��t�j�N�d/���iԶ��ɾ���Oj���O��?�����bd��XDa�?l�1�C$�I�����I�aͰ���F	^���
���[�p���@a�'Ͼ�Ru锋@��I�%焬B>��(��{�$���OH��)�.4�J�O�D�O��4�L	����,�1s�� k6��#��4�	�QU(I
��'���&�?@I��1�L�"8� �{�ߑ))J͆�	�O�(�Z��NmaV��"U���IG~��3�?�}�I�����+�\Â�
�<qqd�/�>y��/�4;�HM�i����5e��H7�,�����D�O��<�r))�U��
�!��|蚈�4�'5���ת��as!��DkҵA���6���9���+�!�$+��DB��+�L�b��	~�!�D�?\|J��2�Th�B�ʢr�!�dJ�Iܱ�!
�����C�۳!��R	GN�$�R��6��@%��7r!��'ef�X�hj�j��K�ei!�d�q�T��oҠeV�{�˵sM!�D�K 2�B�����R%��,;!�d� A�Bd*C���W�,�+��Q�/!��J�xe��j��ǋ�\�Ze�BY!�(X��%aѓT���	�j�-�!�ܦb��t����&2`�z4$�{�!���tB�A�(�h���3����P�!��>6P��:��'9���Y� �<�!��̭;���+��[���a `�9u�!��  �+��/|	b�#��:����"O�h�Ă%LJ䫅��q�z��""O�IcT>S�hYu$����U+ "O�iS�#�����8S�T:v���"O ����:?��e� �O��8��"OLxq�K�+s�b�x#_���� c"O>��FC���ءe�W�P�\� �"OD<yū̾��83c�S I��3"Of�QdK<u��jS0l��7�3D��S�i�q�n̓w-X�t��X�n1D�� `$ݘRG�����5Ya��`Gi+D����Z}R%�4�ȕ^�ț�>D��e�ћI��0b��&Y�^��b�>D�@ E�=����V%�J�dd�ѧ'D��I��9ØL���_�-Lr�1�!;D�,ڳ��7`!ND�c+߂-�>0� �$D���,a�.�{���*�P���4D��k��C�D�씻��D��b��1D�����*u&�q!����n9�Ђ0B1D�8�c�,~�Ti�4KQ�`J�9˳l0D�h�·z�>t`��0�v�(�2D�ԣ�lıx���M�
��P�'<��.�&iR����.=e��T��kK �I����}�|�'̔kJ�� �i�@�'�w�T\�A
�(9�]��';����"C^�۱#_Z i����:3���w""�'/1�0�6E�A^r��^:0��ȓ5!0��u��>SRȹ�/�9.{\�X�X/�sU�|���'FL\�	��Wl6ɩ���/t��p�
�'t�)��˅Z�"�x�
L=��R�'W>�ڔ�ƩRha{bM͞Rr����K+$ȗ�7�p> ^�C�Ty۴S%V	����a( �A�ѷP�v�ȓm�\}�O
�P�
E���k�b�Fz�c״a�.}Ï��J�����/g��M��( �!�d�5a��`�R�ܤ#�T�����!�Z�A��ip2H�Edl����l�!�D�/.J�iTӸ_O�|ѧ�N"c}!�����aZ3u���s�IT�o!�d��$�A�(�����Ƣ�)>u!�ĿN/ұj+�%|����&:k!��	B���(_������-9P!�A"P� ٪ h�R����#jG9!�$"�YX&�=�~Ah�`�7?2l�O�ștC C���H?��P���U��uk��� q��Y:d!#�Oy� kC?�:M�b�I�����	�3��K@��: ����~�����$	�����ڇf�ҭG}bg�;�Zm� �P�]�O���íP�b%�dr�˗�}T���'/\�VH�cL�)�ҡ@�8��'R��X�NC�%JF�Gr>�3@�^�n��IX^2 �3	3D��Q��7(�y6��'z�:,���"��ɱ},��Ua@j��g���y��)� ^|B���+8bU��	�\�ZxRܘ@����b�-4�*�͒ 5h<(J䯚*)�~��ǒp��`��Dy�n4;�� ��y�&3� d�� @�L`Sc%'�y�`5kq�M��?-�r\��f���y�(F�EQ��e�P��=!���?�y"HТbi��HC�+F J�ˤ��/�y"Bʋ	�8����X�o���2U!���y�+	`@ݰkɞl��r�ߕ�yR�[_F%�č`�(���M�y2�����@RhɌD,B1��V�yr��5M@�� ��=5~pɐ�`��p<yp��t���!KR�	���jqE�
����f�6�\���)B�zBڠ��'��C�oB��w� Q�Qz���>)��C��q�f�L� �%ėB�ȓ�� J��
)���Nϼo+�|���^j�<� ��� � 1s�"�+ ������y2π
r��Ђ� )���r��	��Ɂ7,A�p���p��XҐ��/^���Ă�L����+vL6�;���&=�5�"��n�R �lۏ~Lmїi�>��"x�I3���J�4�2�s�����S��@��6�|�`4�	(e�����K�q9�A�k��`��
��^�4�*�A�'"�[S�&m,�ȩ�M�韰�u*R�u��x�i�r̒ ���J	LTb�l�0�"�$y�>�{G%��*L��'d��(�R�(pс q�D��v�١$ɒV�V��,gJ�At�4��0��/Mڼ��$H%w�,�1aJW>�,�#РŻ?Ts5Ί7���2��~���1�t�3���VX��H�� ؚq�ל!��|X"�B����1o�O�����C�����!H7j�8��>&��哇ƚ:��v��>Y &�x���Cc��{u^�g�j�����'�!s���:%�%I��W�~�*я{�R1U�p��;$���j�!Q2m��Q����2cbW�G,�}�4�C$2�u�c�G8w�fd{�
�%�8eC&�H7}Fz�3gjG�����q��7>����M�j}N��1��9��q���=0����>�8�r��~=���E�*�N��'�M��l�v4z\���(�قuȈ�N�] ǣ�'n�a}���	����!�
F�D:#bX���q��d�j]r�a��H�jeH�=��	�Ϣ�7 S2.�̚R��92��AjeT
���qo�m����J��\�XggR�7/�| @�#z�v	
��J #��0R��A9��m�p?it-��^���
&�	�,{�Xw-��F�B���z�v!��cF�+2�$Q�T�~i����O�Z��ۃ�B�y�>�HY�2Ez4{��¯H���/��$:���H�=�ņ�/x���T�C��@���4ر�I
��OȤ��T�O��0�
I�;(�娤�\�|P���r�	=#h����C�jJH���D�W�2�Y�{�����e�⌨}Ҭ�� �"J��s�J�!���G����>	��Uąy���yr��`���o��Vi��&O N=c(�?��H?9���hh۷�Awϔy�"F��Yt<|1e(|OD9�A��7q�iر�Y	z�Șk�*����*����Y(��-]$L�@����R&Z�Ia+�x���B!�R��B�tLɡ]�jȰik��
��O�\�s��7\(���E!�`���'�|�Îu���y�F��$1À")���u����2(�9FLH��iך k�#=Q�l�0H��U�I�l�$U��<O�� �ix�<����j��q���O��Q�Y�,^$T
Z���Q/��4�h��C;��	d�^u��I��6��|�D�E�>���`��J�LJ�����4�Z��c����iɴ4*��*�L;�I���;���rUO]�]m92u�,�,7�O`����;��k5̄(%�Ƹ*3L]4\�:����v������9ʤ�sQn��d�h��q@K/m�+W�ɞ[�>�����P�T����h����ė�����µ}�F���l�J`qǢ2`ȭ��$�j|����Oj!r��**�"A�¯�1A�`s��	�OQR8�K�&xԔi5m�T,��
��+�b�$F)X�c�!Z�@��}��Z̓h�QB@��;@*�  ��1(�	�n	D���"�O�!���P�� CMU[��*	�>��)mI�I��eQ�;��|�2����Υj��![6�J?C�d)�"O�T��.]/5�|��)�dm�I�R�L�'���O%m��P7�W-2�H�O�2iߒ&6d�r�5ȮpY�ܵS�,kfK6�̕����%+��\�ι~j��O? @����ǀ�05��IԎNw��A���;�io�Fq0��Q1��Gz��<�)��m�<	��q�w�]1�PM!��)X�ȑp�=���,�1O����콲�a�;K�T9�(N�����	_��Gz2�+*�D/�m?�"��;gh��jCHG&z�p@�C��iR(�q�'�1O������',����w��-��̇�tA�r�3E�2b�yr�_2`��r����b�fNEa"
%k����� ��h��	W(ڰԈ���3���|R��i����v!ƖB�|pBG�P_�̴(7��,/�bm+��4���)O��A}��AJ�	8>��aש
L�0�i�:I�3	�G8���pO���	��V� ��Qɨ<��4�n�c;6�є-ô31*h2�C��_zȷ�ծ�0=ѥM�J=���bG�,����c%[�FK��I�^��QT-Wn�Iʟ��'�l$�g�y;NA�9�Y�l�1%i� E	��}!kޱ:!1O�| %cΑz�Q�)�N�d ��R��̓A�T˄�H0袤��M�H�'��������M"�o F2�1��d۶��M��CYzx��d�5v�l�4g��0%�����	��|�'s�(9�`5j��$j� V0��N��sVQ�B�^��p>)c��� paϏ3{v}"#�Uy��i>��'��٢�����Pa�ўqҎ����-3az�`�)�h����Y�0��ᄒL8&�(���(��a��U9�<9U�=oШ���݋2L�Qp��{���E��,��e�H<c�1O�a�X#0���'j�d�H>���9CT�ӷ�-0�@%bFg���p@$`Bo�B�ܓ7LU=���=1@�������W�A���8C8Q�����t*��-(`c���a8�`@�fԌ`�lQxRA�X� -���&t�F�
b�'5
WaH�(
�d�%AS*
�֝aO>�!IC
��<	#˜�%��̀`�AS��1��&S��p=q��D�/��˨On�p��]t)���C�D(It(a��'����G�T	�)c��F/�� hUsa癘y���F�]�r���'�y��T�8�� K@��+{���Q��ۯ9̅0����17d��O>1����q�d���D�<U������LhܓN�2)��"buGj98��<	Cb	C���0!�� ����$*Fg�~]�t"R/V1nz٘���mbhH���Xbub�B���IaX���
N\2��C��
��"�I�I�����c�<��t���oB�y��8w�
P)V 5� ��G�Ɂ !��J-p߶h���6wHf4��HI5y{�y��7�f5��@Y9��� ���i����b/�%��eh��b�az���2c2�ks��)��L���1&�bY9��ۼ} ⫁���=�"棑�|�a&��y���=��
P���'��>�Q/Pp� N�� H�������xy �&�����ɾf�^� �c��U-�oy��i�E+r_:�3
�S.�����7%��D�����'�J%*D��&^�@�c������S�'b��@��ނ��Dpae�S�ć�0 MCUBÍ�D=�����1�J�'��4�z�@��h��y̧h��'re�ւ��z< ykCK-&>L��'�rd�f�6�h���@�Z�N@�#�%�mQU�(O�tآq�}rz1��I!\�^��@��4o~z�8D�^�n�t����%2ܤx�׃�w�t�� �/� ��Չ0G }�t�Оaޜ���A�Px�ϙ !����9o�x��A��dW3�ޕ1􄋣l,�8�dI ����Z�6���� M�TE�<+��Y�y"F�;H?L�s'Ó7O̺�J�Н+ⴼ����7�<x����$0ܻ��ԝxB����ܵbv��2�xa�ȇ�yRɍ�X�ȱ�V�[�I[vl���y�%��r�f�8!ȗDJ�5:���4�ybfW(L�-���7@������\��yRG��aN�`k �Qan�k��P��y�c)iL>X�gǎ>,��"�IH0�y�N�<�uZ��͚"<�W��	�yҪ��WX��3`�`Ț���y���Br�T+ËL�6ʣD���y��ݶkd��9�m^.c�$P#jG��y���L�,%y����pbc���y��-�T�&�)r	9�Dʻ�y�H:��@A� Rܰ�Ԧ���yR`"KtJ|�N�,!��D ���Py"�P4v�z\˴MԌCM����t�<qg(;M�����-�}���)��Sp�<���I	/oJ����	P����J�j�<فC��	�|�
��ẔjJ^�<�E�U|��9Z'�W�!g���"�GX�<y��G�n|c�I0A��<#unFZ�<�E4�ƀI���25}�X�f$�L�<��֔<�+��G$[pă0�	A�<����i��ԩJ�Y$Yۂ�r�<1U$�@�8�����
�.�y�<A��^g���E�Ջ?��}��'�N�<����L5�P��2_��0�jFH�<����R��
��
R�ޕ���]y�<��N�/y��Ȉ˄e��p �Xr�<i�!�3Z�d<c�a��(8%Ęj�<1�.�����f�C)��y+F�g�<�����p�3�Lu��ۤc�d�<���:M��}@�
�fC��b��d�<���F�@�&��Pxl� �X�<��d�ЭPu��c�ڌ���<��$���S�Hc�Ԩ%Ør�<�w�BR��tp¢GUTv�X5h�t�<�&��:�H��ED$R�U�3�j�<�S�/o���"$n� `]���b��f�<1S��6#��]�b��������N`�<��ܺ�6ݡDؾv�����\�<���1� JPO��e[|Ų�BIr�<I)<D|�M�r�Hv��ы,l�<�T
{L�edlԾy{�J�g�<� �#�,Po�|A�Ȟ&XިE�a"Ox���)G�%PGIׂlI�"OF�xf��'|��`0� �8;��Yk�"OԠ��	�ao��� %A�pM �"ONQ�V��Rb^��� S�ް-�"O�H�f
AwH0��$���*݉W"O��ٷ)�血���48����g"OLh�A˴z^�P���R� ~@<��"O�܀�&�.�D����R8STu��"OB�ȠJ, '*S�؜�I"O�����RY'XA�#�����"O8X�5j؋R������Wj��CU"O�m�R������ԤANn1s6"O�Ͳ2J� ��	G�õ��Bf"Oh��p�2l�T<yU`ƀd���e"O��{����z��/ȥ �-��"O"��u�N#�>���\�H �,�@"Ov��2c�=�ĥ��$LI�"OL�2"���~g�	� �V�٘�"O�8ʃ��`Bf��2/��2��%"O 0�Cy���A"N�,���"O��S�u�r��Pi�OU�˴"O:��U��wk�m ��7MB�)c�"O �R�eψp|b��g�s����"O��� Ũ~n �����V�4e2"O�qq�P�>/��A L�*i�U"Oh[��F-Nx���嘸A��ec�"O6I�a�6J�< rE�6�|�G"Od�����x羼`��K,v����"O8���l�7��0��L4�ࢄ"O�h@󋌓-�,���
���aY�"O�4�FiV$�骇c�G �hp"O6�i�+T�zU�Y¦Ȇ��ι�"O.��%��(N�*�*2H��y3"O���T)�%y*��v�8+��=p�"O��x!cC0h��3�ŋ�W��!��"O�0�q�H"$6x0��I������"O\��ċ�.�`bI�^�h"O`-�
F�5� 5�V��8��"O$�K��<I����cŒ�t0�"O�	i�̀�z��ݣr�E�@�(�"O6U�GZ�r<P�E-F���()�"O�y V��y3Ȅ1�L��q�@}�%"O�,y�mO_Wƕ�f+|��!"O���m�<�HYБ�� ��)Z�"O(تe��$PWt\B���8�0X0��'��'���h��Ö
��p��N�	^@@�'��8�A�F0�aT!�0 �����dԷk�����g��-[�?W�!�Ą1)���qEȖ%sDePeJ� �!��ӽh2��:��	7Y*|��	2�!��P	)8���X�J�
��%�9N!�O 8�>ڲɛ+m�\��AL��!�D�<2��`���_��h���D�!�D��O7j���D�,�P��2EX=�!�_�T�����C�`xR�ɸ�!��&lB̈w��4�J�ƭ�!��	�y�F䂕D�5$���0�ͻo!�E�n(�����K�����-]�6O!��.�BD�[1Et�TA���r>!��8kɒ�*���0n��Tؠ�!��%)4.T
��S#nW�t`&l��F`!򤝔:4 P���An���Л>9!�K� "���	k
�!S�-!�� 
�I%CI�
�yQB�=|*��"O�-�Ql̨*6D	�n�\^�R"O(1�3ǊC�ʁk+--���R"Ot](���+��ᑯ
6�8a�x"�'��	H���D�R@���q�
�'���FN19��P��9m�%��'���@���(8�҂�@-�İ	�'�
�@!��qM%b�  l�A�'��B���<P��*⮌�'}�b�'��BaD�j*$�@�IJ0m��=�
�'��LJ�O��{�/
_���j�',�@A@AJ΅���ۋJ[��;
�'�P�(�O�S|:��m_�FΊ���'�p&cЎ>��%�g͐I��'dzu�A�8|��Dg� a����'�v��#&�yK�_�K�.��ȓ3Q��pR�r�q+b*�-Նȓb5\h8E�!>���#��Ϥ	~����EȬ���2Z��Eb�o�LM�1�ȓt���Yg�9Fj������@��ȓӆPX�똏_qYIc�Cr'�ݤO�=�J���;q�,;�8�7�T�<qw��0zP�y��+J���y z�<q�c�W�b���'�?OB��Zv�\�<i�'�;f��	�#�T'Z[�x)5eTV�<Y��*r0̄�F���"l�r$Q�<���4<0��5lޅ#=(��aZO�<���_%f�x�e$��N�ػ �Nb�<ys�̼D��x���ۓ �y�C�S^�<�C��:zl��r���1�0˄�[�<�h^.�"��""�:ڎM(�F|�<y�MY���ۀ��K	��A�'�a�<�ҠY8�����.G	U��!����d�<�pG�R��8&�ZR��j1(�U�<1f&�?@�D�E�H���VF�R�<�w�J4��,�d��<	}(�`"$K�<�V��'%����[.SP0j�o��<I�G(z���ʥ�Ȕtt|�q��u�<!���.,�l"�!�%�_>-{�B�I�}�h=B�GѨa�R�Z�읓*U�B䉅LT����#1���්[[�B�	 q��p�Ƈ�5G�c�V��F{J?+��
4D^(*�<�D"&�!D�x���8m�m3�+U P�fT;�o�R"<���O����EU�e��IjęA1�|Q"O��Cʂ!K	z�x���&1�)��'ݛ..�O4�R�+�<���C���@��3"O0T�C&J-!x�)å�ۚq�E ��,�S��ɔ;��H�D��=%�T5����Zg!���c����ݠ$d��+eX3wd!��"a�ݣ�`��d�!4ʏ�C&!�D�=�z��D�=x�j$�4j�Oԣ=%>٘Ө�J��@�%ΑV��J�a?D�Phgɏ+1N]�Q�wF4}��!1D��0�@c�v剷�S�3�H#g0D�����6;����	>�Ȉ��*�>Q��'A�S� dպX�s��`�f��'4��{3�W�`8L P�кZ$ʰs�'���G!Ⱦ`AmCR&!P������D!�f��ĉ3�;^O�� GR����ȓ�j1���(�6ܐ -�$N~�H�<ы��	S���۔�!����X�!�!M>� e���
o���q'��fd1O~��C^<����A��jd���lJ!�� n�� ˔_O�miB�-�P�t"O4=�#k��hx<�c��8`���"O$E�%o(:¨ɡ� *�@i�"O^]I�J��O�/�&j)�"Oؙ�"k�qmj=��u�����'��	J�
풠�R�|t@ɢ��<��B�I�L��r�$�4ӆ BZ+Y"����7�Ʉm�.��I[#{�L��I�B�I�4�~%�bk�z��ۣ%��"?ٌ�)��$�4C3�D('�����!�Ą,�����"��~3���'��Kx�'_�i����'��41M�&3�F��	�24��
�'�6lC!�ǂ�6X"�D>/��
�'���a*��(�L@�c��+E�2ۓ޸'M�X���]|�H2C�F'$p~ i�'B"��ġ�pT�i��/��*��'����6|�Za�֩
�H���'��a#�\}���LM!	�n���'�ў"~
ceب �ֈ��D��KQ���a!�q�<ٗlwt��"�Hx83Wϔj�<b�W�!2��`7�ir�tK�a�g�<Q�'�"-Vmp��O�XƖ���eZ}�<���y������*Q��XF%Gx�<��� 0�( S���$7�:��5��s�<a�mB�+��a�kJ 
I��@�I�<�D��"K�=��͕CJ�xǧE�<A�h..�ŉrߛ�B�K���V�<9P���a.ap��TH\���dT�<y�H�r��Č`P�b� I�<1�-2-\}�ˋ�8Lؘ!�
G�<�
#y��dc�G���O^�<�ҍ�xvP]��e�M�,���%�W�<	�&�<b��U ���
c��@Rrk�z�<��+[�~j̃�K�-#U�����q�<�3�նj�5��N�P�v$��ny�<)��L�J,���ْ=������u�<r#Թ}�$(�7�B2�E�"Y�<Q0B4\��I�V�@�VF����.�o�<	�ڿ~��,�p�S_?~u�e��<q�7W�40�LZdFF�a!n�T�<i�F���7����RTq�u�<1���-�� ��Z#'�!�&q�<qү�9	U|$�g�J	gr!!MUi�<�Gj²�b�����T�8tNO�<!�FčG'`�2�I���]��$R�<�G,9N�h1��f�z�]��o�i�<�ΟZ�aҕ��g�n��R�h�<Q�`��Z��{j�M8�cWa�<	��	 �!�% �<�z�z�e�U�<Q@ϊF���p�c��͐ۀ$y�<ɡ�&jp.�A�!F @���7aK�<C��=�h�RA¤D��`�O�J�<���&$���	�7��mP,�F�<a�,�(Zh� �s�~�-�u��K�<�$A"kAF�0f� �,�:�S�IA�<	�O�W��U���k[�u��b	y�<r(��#`d��W,��f>�I��w�<)�� <^���K/2&7��/�yr� �̸�I��Z�����h�	�y�OT�xԫ#lZ�r��&�Ӷ�y2�M2>�V4#�T,8�(��J:�yҩ
�
�ii���2G��[A�D��yr#3.f&�#���r���I�y���j��mb�߀"��CW!�5�y
� �%�чI�W��e���K!���q"O��B��!��cQ�G�,q�"Of��b�?$���m܆��d�"OqR��S+g�Y�v�N��<�7"O6�x���"�xi�!�ī|
ɉ�"Oj݀C��7p��ʕ�*g� ��"O��
@Jβ50V5�e��TY��	 "O�< �<I����O�T�L�"O
r�V10�0}�E&I����"O$\�q��M��5cV�D+0���"O:X�d���������H�rh8%"OB	���0P;ȍAW���D��JW"OT�aM���xh�O�%�Y�a"O�riT5@ ��
w��w�nA�1"O}ǀ8!>R��#��,�4UBe"O�4:�O[v�p�J��H#dYl`�"O�e�7ɝ\�>�Sb	#���"O��ڴ,��fp��@�aP
gxQ��"O��`���	$<�E0�lJ6ɚ�"O��Ҥ��J�%Y��R�S)��2�"O1���4� ��d烟C�RE�"O�a�O�: R��(ӚQ�4�"O���L ��5?��h�c"O��[��V�Tc��s���	��i��"O.� 'oǒK�LPaȈl8�, �"O�}��:y�:�� :�0�"O�\���n�p��u�^>aa6"O���e��Y��,�M�5�܁ "O2�y�����.�[���i�"O����z�<��G�	� m�ى�"Ol����	J��C�O� i�ɚ3"OzU����1��r�+�C?`��"O��S��Gu(�35l��m1F<h""O��	�a��t�\��5d�8��r"OD �-\���B�Z
��ٱ"O�d�w���f����M��5�"OZ�$��&4l0EU'���"O�`iԁV5J/2=Cc\?x�
�"Ox�z�����.W��6��"Op]����8)4�3�O���>�s�"O��C��
��@��o.Iq`,ل"O:l:+Ng�5B�B�2�β�!��F#z� ���h�R�ȩ��	�Q�!�D��J�d�H%_�1s 1<.!�dq��y9qd��t�5�^�
)!���P��	� ���T���bm-!�:3����b�)\Q�Pm	!��Q��a��`V>H28��ˆQ�!�DM�Mt�đ4l@
�L  ��P7�!��i
 ���ܯD���� �#$7!�9o��Z¤ϸ~�~�:2���$.!�$ � �v�@��@�@��4��*!�� �N��e��Z
��3)�6	!��[�x���sk�]T�A�j��J!�D�8$�|Sv���I �$s C�
F!���C��e�*�!�z�Z"�
n9!��&<��x�`�S�S����i !�D�\I����� ޖ�Z�I:!��9/�
pIe	��T_���i�O!�d�9M���Z�cF(9�|m`�Z*!�D�7	`��� T��JP�]6!����e�7 ײS�"�<Y��C��n�f���^�>�`
ŤQ�C�I4��h��7�n0�Eŝ<��C�)� ���v��2��� �	G�P]�`"O�)Wg�&0�����%Ǆ>��,a�"O��r ���V!�Tb���ê�y�"O�e�u�́NU�	cmK�~��]��"Op�I
R=d4���-a�xAt"Ox�C��-vD�hE+%�"O� ��P���\�&��an`�"O�\Ó���8@�$K�XL�"O>!��<�b� �J7�(ux�"O
�SwB:7��M*U�Y�a�`�y"O4Y��Ag�k�AL'|u� �"O<aY��.T��d@��J75h�i�%"O,���./t��0@V:Y����"OL��g^�>>|��ӅVu7��K"O�JC���5���Yc �쑂"O�S���I�$���F�D ���"O4ͪ��R�r�%�V��]wT�#'"O�	�匄� (jթT�Μ.�`1�"OȔ8%}�1��Z�l�ڶ@�!��RA4�B0�)G4r�q"OB��`�܀e�<��%��R�"O�+@ �k�dys#���:�s�"O���񌘙 ,	����y��Ԁ�"OB�z�#�j�@ӧ�d�fx��"O���"K���<�j5(��T�`��"O�y�f��BUu
2*հdM���"O��â��(��D���)]����U"O�0�P�ոWN�]�`�[��~8"O�Z��FOx�ófHZI�%"Od�ӓ��&[�!�� Z/LIj"O:�k���:�ѐ���	<9{�"OL�+%I�<.[x����ǋ%�M�b"O�MZ��ԏbhf��e�#~��c"OнbP��ij���-2�0ZS"OpT�3���`��\:|PJ���"Oz<�Ve �><�mϡgEr�"O��j'�̑Df̠3@+�&Q*�� "O�J��Y�<�	%�w�"|Sa"O��q ��M�p��Q�
�u��#%"O8q�Խv�Τ1uhN�1��A�"O��i�*rA�@:ҦN)ar�h:�"O>=�����X�XRA�K��(�"O.S�FiR��U�j���"Oԩ�dO��[`#��:y���"Of�8v�3Id8��t<*�xA"O8��'�en �`�B73:}�"O���M��}&�A�$ߠ�h	t"OzѢ��W�V��Qj�����"O.t�q,X�����S�B�,�"O�vY|� �H$j�����4"OxE:�ϛ�Z���F���ad"Ox`k5 F�#��b5��r�p9
�"O.��1#D�X��=sf>Q�r�K�"O��k��A�2�<2��:�0�"ORUj��9:>�P�@�9S��d"OH�+$��y��y&�=>\��"O���U��bvtpQ�AY����'�B:OX\�e�Z(P�yPU��nk\���'"�T��(AKؐ��eI�~g܅���3D��b�N�?pˈ�;�낗EX����0D�P:@�'Q[6�Y�*!%h%;��,D��2An�(?8��!დ�My;7+��i��P�P�>䞝a�m�0�0�ҕ�+D��C�ϔ2D�����(>] I���(�O��)� ��K��;g���i���?d|J�3GT�F{R�'�1O��R3�wl��0]�K%"OBQ�`��$F24���6xUB(b"O��㵀��"��ԁQ���"�b�C'"Op�0ᇏTx���)ݟ5��0ئ�|B�'y~8yc�z62�1��D+,�C�'�b)�B�֧ ��qX�-#D�<es
�'���b��\|hxȇA�'I[��	ϓ�Ol�
��H�E��NK23�i"Ob,3F���i���E��t^�Ц"Oh� T��*���flZ6Z��"O����H�]¬�����2$A��:�Y�����)X()R������f`|!�B�Ib�K��0A`��� ��IG�C�	*9��݁(�J
���)��d�O�����BT~i����i���׬ΏP�!�Z1��0r宐�,�� ����\�!�߼Qۢ�1%:�Č�p�TX�!�dT�0і%�6[�`��
��r<O֔hse�[��lJãG$�z�"O(�۵�/�lQS����?���"O ��"	1!R���W�R�33>���"O� �1	��P��D2�F�I �p"O\q�Qj�q�N���d�F��P�""O�(�'�?�H��`톹S���7"O4�{�j�>f��a�R ;��b3"Ob��qL0(�8 �)3=�l�g"O*a2׉q��E�)��
�"D"O(Lx�N�6i+T��ǉ;aRL�T��3LO�����$��٢�DC�<����[�|�Iٟ��IIy�T��O?N*s�������J�T��'2�h��\�	p예4�Gxt�'WPEj$oU�NK����雙>ր��'"��G.W̤��&@7 5�'x.!�a�?c�b����W0 ļ;�'�������+x�h� LM�j��`���.OQ˵�	6LD�i�� �f!d���'��'��)�-
�k7��7/�� %�5xH��'�����L9_X�퀶A���
�'"R�R��'*� 1�2�L�db�0�
�'��\��ڲ]lmт3_��Q@�'1F@��Ez:P�Q�[_0�-O����O����_	c�8�* �T5M�IK�,Ȏ2�ўP��:0f�h9q%��Cĉ	� S:r�O�ʓ�0|b OUt�tl�sY+!{�`X�K�<Y���6+蝡E�V]m�\ؖfAI�<9&�M�IKh�w��/=�]�P$AG�<e�h�{�L��)���&F��<1�d	�r��]�ǢE>\�$���Ŗ~��b�ȠG��V-~Ȉ%�S;vᱬ*D��J0�"k�nu�̊-?�B0ð'*D����K�x� �r>��[p�&D��D��	�n�`�O�O�
��#d"D�0J T�q��y	�f��-+���l=D�tّ�YW`UӰMM�c�8�g7D��R�%�7���Qn��|?�x�6�O��DHsun�ѷ!O>m(�m���4o0�B�ɥW�(�#���D��A�,�j[�B�I�8u�dhSgԝ!(R��S'Z�>ئC�I�-f �P�ZiނZ�C�>V�C�I�&9ؠ��#��q_�q�V'!,�lC��B�%�V�L��v��e�0a��㟀F{J?��ж*>�Z�i
��5DG=�O0��$��i��l��r7��t�� ��S�? n�˴��&Cq �)Ȟƈ-i�"Ox�1�A0H�P�AI�s��iY�"O�i�ф�'UJ z�*3H���"O<͢v�:���i#y��!��"O��:��P~ڈ���A�o�ʥ�0�|2W�h��S�@��t
s��AhP{cϚ�z��B�	 O�9�3G��;Ц1Q��\7!�B䉻E X\IFG�R�.y���ع;)j�d*��r���]�(x���Q�CS*uj�,!D��R�ÔN���2caM8X�p%%D���O�=i��)&b��0ъdR �6D�p�$��;VM�S�̜']��J@7D��)d��2y����@��x��6�5D�T���$9���E*���+a3D��8��~�R�Y��
�&?�`bC�/D�lQ�H�����:h���) D� ���h@�ص,��%�"�!%=D�T�u�\<L�=�R�>"�
��9D���G�@"w��۔@;o�2��sB"D�D0%Mݑt�m���
�iE�w�?D�xZBN�$a4 ��U���g*OfM���e���3n�7N�D\`���z�O�����R /r��f�ȳb"|A�'ZLs4��e�2x�a* ��'�"H�+(y4�2�Q�RL�@��'t 3��Z����3�O�,��
�'�ܹ��f��E��2��-���'rtu����u�pK������,O:��dR�*��g��$,��hW�Qq`!���t\� b�l���fb� P!�$�v�� ��o�
3���bȬ,6!�ĝL�ɒd�j(s��;!�D��)Mօ(&#"���gH�eў��ቶ3��-�Zr�ݡAF��3����@_����I���{��J�zl�q�uI'U����O��$*�OPuBPEF@�D�s�i�~� 	��"OB�����z���7(�}��@Sb"Od��Y{n ���-L����"OH�`U�$1B�8�kڝu��O4T%�'8�Qaƈ�1*��&M<D���bΖZؑ�a,GTD�g�<D���cH��mAv���"Cz��@%�9��3�Ohܲ#�-�|=�UF�2gi
��B"O
���|S�Yb���UST��"O��В-;_� Q�c֮A�ГU"O�X"�����`!���9>2�� "Ol1���s�qA�N���ˀ,̊�?�O>!,O1��?V�B�Z*�����L�������<	U��yH0�1�)ѡ$`Z���C�<a�S�ɔ��e	N ~�v���$��<���%I�������|���q�<a7kU�S��\`�2�lt�w.�j�<e��,�T�p;W�L$�*MR�<Q���5b��s�V+�
T�ΑPy2�'�����BL�����ھ�k	�'{H��׸y'���� l҅b�'y�pAɈ83�L�*$ES!D<�
�'��Ax���6��<���ѡA���
�'9��E��h\ʭկĠ&�P�Q
�'/F�Jpc��Aj�����e�c��y��Y�~��W&��<�R%1VB���?����sS� ��jԾs|ءef�->�d�ȓnr!���<���G��D�ȓ%@�zU.��^�v����2d��̇�S�? B ړm�'�0y��:l�v���"Od@������eȉ+��Bp"O��!b*�a�8���V��}�D"O�e�g
$1G� S�Hڣ0$4��"O2]Q�Nٌ!�ޭHp
��$�K�"OT%���P�I���QU�,s�T(d"O�H�Tg�.�6!JJD&|lZ$��"OX�0b��#oӰiJ�揄KX�|�p"O�d�f�8<�D(�A-$W�9�"O*�ެ&�d��["9��w"O�RWDE6\$ܭà&ۡXW�) `"O�����Ӏ��0��d�'p|��1�'LO YcdH;O��t*�N/��2e"O���%.�S�D찆n[+k*�bQ"Ō������N�Sė�J?��re"O��a��3h����!�IK!N��2"O�Z�B M*MFiЕ-����"O�dKe���D]�ȋ� PLd@@��W>���
{�������D#�$7D��Cg��a�rZ6�A6kJ�y�U6D���4	٘B��[F͊�z���'M'�Ic�����m�줻��?����:D�����J�T�8�bd��C�Y�0a:D�$�C��Pl0�3��\_�	JbF>D�l�#Ù�s�p�G�:�<=A��<��0|��*]7J�us"�R�l���"PN~�'��Y���n���({��UY�x0�
ƣ�y"�� 2�C�g/�Sn���yR�B�v�����Ic\.���ކ�yb(�5Q��(0ħ˴r��bWH�8�y.�M�H<�g"��T�~�2�E��y�h�MA�Ib����c�f��v��?1�R��&C~rr"I�!�"���,ٲ���	� �'�Ш���B#�\
o]H@s�;Ҧ�B�%/D���&�լ��!�[��<Ɋg�-D�@S��ɄM�	#rJM3$����*D�lI1�\��`��U��I�(D�� �N��=.���L^�2��"D%D�L��A��6�@�4I��j�.�8t$!�Iʟ\D��'�lX�4��&0������������?����	A�g�dM/!�F�dc('��H�+ރP�!�����S�����xB�N�\�!���YB �)�,*�&�[Gޮ�!򤛙H����׍��J��!F313!��]����2/V�F]r�Oʅ!��]�J��̺���Y�ٳ�Nܢk�r�|]�"~�$$0w�4��/��{�b����y��>W�x���H8au�����yb+|<��AT���
R��b̓��yR��'����G$U� �l8��y���6�HB��U k1"���=�y���?V�X���wҀ��Ee_��yB��L$�-"�*>uʚ��w
��?�����t�t����Q�+���q��-_9�@�ȓ6+�M���9��R����vxȇȓ��A�m@mp�-����'Ŋ�ȓF�p�A�F\5΄��9#�@l�� ��|�����Y=4���6p�b��ȓAZ�K`�70��`��*EB�@���P��0��H� 9��i�!z�0���)]����J��|;��o:�,��fD����G�E��2�c�>O�̈́��x!R'X��@�r�O�i�(8����0u`I�z�: ;�E�4t�M��S�? �YpQ�kך!��H k(D�P�"O�i�L��-�ntBJO�P�7"OjU�&M8&� 03���*n?4�T"O����FIo����I��1( ��"O4�2'jC,.T �Rh3M/���"O:\�RaΨp?H!�Y�n��Y��'bў"~���Y+Ji �.S%(<�����[��y�n1��E��C])����"��y2DX$f��Q+��X�ZY������yr+^� ة�7l8\8\��ꄣ�yb�<U��l@rJ�X�v��,X�yrH��h?��HH�]�: �v���y�*6��л�Y�=I��6h�=�?���������8�C�_:6�R]c�lN&�85a��,D�P�"�:F� �q��{\l��A@+D� 6`�"<<*�
�j(��7D���4�F�*j�2�c�=i��A1�4D��k��x �$��8<m���-2D�����K����� �Юz�x��+D��ʴ�W�7�����n͊b˴�i��(ړ�0<�H�.6D�Jр����Jp�Kr�<s�.W�k���,�&����H�<�a��
�rѪ�/��yz5�SF�<�Nט��:�$�&,$�0�F�<�a�@+1��ј%JB	m+܅*�MC�<���Ųf����3��r���q��~�<�ȕ��q�G�=Ų=���x�<m�\NlR� 7X�r9���w�<9Fō<F���3�އ_�$A0��w�<)t�[�;�p��U�܀bX��2/�X�<�e�|.�B��^�4���Qz�<��؊���p�ŵ�Y�0�u�<)���F��)«�.A��`�U��e�<�Ӥ��oiV���˒T�zE�7nBy�<�䄋,�>tq�OF���}iӦ�z�<��ܡ}�f`���1�ZyId��`�<���$4,����v�r�a"�Z�<��(�\��ِA��  ����V�<Ia/�p+(\h���=��Q���T�<�� ��$b�����J�,�#���h�<�!�

F�xDs����80r��~�<!�	M,k��2��������Gv�<1@�Mm�.U
�&���m���Ug�<Y2L�Hw�L�&뛧�a�Ǟa�<�BlL�5x4��a�ڠͬI����h�<i!���5u��To�3ٜ����g�<�0&�Rߖ3g!�u�ѓ�I�<��)+��M0o����.;�C�I��)��l�%Nb<ْ$�(Wf�B�ɖN�L��5jJ:p�h�R�U��B�I�c�+%�Yd<�s��� �lC�ɜHܱ�a헤��i��j��B�I'g��P`0���4-�E�D
�� C�	�Z�A�U��5w��Ź0$�6C�	�aZT�֪I+[�mhp 65B�6�����P� ˠ�y��qd�C�ɻ=�4$�J9�Lqq�Հc��C䉬#@�W��4l��1Z`�-k�C��&
#xiI����7���w�F$K�B䉤2jv�I�MT��zո���$�<B�ɗK��+�>&
d%�Ձ��a
�C�:,�̌��!��FI��c��
��C�IU\���t�'8��U�P�Ň�6C�	 �d4�6$��h,� ��.]�C�)� �K�O�9a���`��Y�"O�l��Ϭ<df��0#�9�&�2"OV}{sŋ�4�B]�`H�%V��%"O�`�fԹY,��[�hϝ�� F"O����0��ehM�@i��{�"O�p���R0��ѩ'�u *!Z1"Oĥf	S�Sfk�L�9KJ�U"O��yP�B�+�R`��	52�ȃ"O��3
�#}�PӪ��5�E �"OPq�)�M��U��o˘mטy@s"O��'�UNZ�q����`�S�"O*`�TرU��(Y��2�6##"O�u�S�(!�SF��<���a�"O"�&Ǐ?�`���@ƽ8D"O �+����G�Z1�%lS�[��ؐ�"O.!rĈ��<�P�qa�C�1d�('"O�i�3�?=��adN�G�}�"O����憕SdN�zbN�[��t:e"Oj6�9$$3vF��6ps��<LO�H�秒�K�@��B�Ga���"O�Q��$
� �����gU4�+�"OL���pd5r M��1K��%R����	��p9��\���E:8B�B�2M�&�)І�g3.�h��&�B�8d�Ĺ��&[����ԂO�4)nB�I�:��eY�H�G�U"��w<B�� �r��P�Zj��ZE��w�B�	�zL�$��`
�>��D��޾�B䉼b=��G���%���ؐ`�=!:$C䉽V�<��6�	~�]��P�HC䉴I�%��П)�VT31��%GD�B�gh�]����0<�a�
�\�B�	)E����&"����f���|B�I3eB�Tb$��+�
���Q-83\B�I�"|�TGĹp0p���)@B�	:N��`����.>֕�4�O"_�C��	�r��6�ֈ!POM��B�	�X� ���0��,#" �8��B�Ƀs�аy'�Ƀ�@�̯8t�B䉩t��bf	R���X�"I{��C��)xv���Ū�?�@�ȇ�eB�C�	% �|� V���J�bd �)&��C�	��44�R�S��(H��F�]�fC�I�h^�|I�^�(
n��n�:g�*C��6j�V���@� b�ݽi
j��ȓa�Xؓ�.�(=i�͚���,��ąȓ�و&������ݶ9����)���"�M#;|�`����O���g�5[���i�A��#11�5�ȓV�p`�
�4�nUS�#[6b��X�ȓ9��3 A�aH4�u�D�=� ���B�z|��L�V��K�'?�Ąȓ�H�q��
,I4Z�r�P+{���ȓT�\0vnǙ)3�t�̇;ڤ��x�x�{`�BdT��k����+�p��ȓ	�l�Jfɋ�q L�S�z�����[��YK�
�XJB�X���9�����$�$�+V/_.v�`��"�:fHK2D�$I�fو9�thz��	������<D�\��ܻ9N�A�d���z�TW�8D�غ�ĩ$"ԌĄ»a���I1D����ǟ8jBfT:��@�%����3D����,B�BE�"!��}��P���5D���pf[�p6*�x��B�h�Ҋ/D�� .��&�B	n���"!(�6��"OZ �1O	�Wv���eo��G�Ȣ"O�%�4D��rP<(8e	ѣOҖ�h�"OLyp�[5P���N#t�ڤ�s"O����6+�~=ʡa,K�&��"O"�S%�,��h�`U�s����T"Oڭ�D&@�*�إ��7ҵr�"OR�(a�e�R0YĚ����$"O�`���C��h�#�Ɂ2�*	�"O�8:�'H���Ug٤	H*-�"O�q��)G�	�hy� �1%:� �"O����*�'?���V�L#6j��R�"Op}�$A�/W�h�Z�F[snL�"Oĸ����<}c��P��A8dC`T��"O��)��N/|�ݑ��n�ZH�'"O��3ALR&=�ȕ�pĘ�Q�hm4"O���r�Ф(i��9�c��i�`�*�"O��Ra�� ��u�P��� 0��4���O ���Ћp��2�KP�����'�0-�!�[�R���RЉ�"̲� b�È/!��Z*c^d�7��b)Ʌ.ͅH�!��,ޝ��	K	u��9@�#�36�!�dW-'�||{�E!_��UZdcD�W�!�J���������1�~�!�d��vl]�uj�������Ð���O2���0�Z�����O����T� �!��?R�8����I��@BB�uT!���#T6��3+Q�R0 컧���q�!�$�&ry~���
!.�`��H��5�!�D��<0��(A�&�ZéL��!��Ӫ*{N����wLx(Ƃ�{�!�$��j�-�Da	�e�\ =	��O����`$��pFN>G�6�7瘤u�!�$���Z+���9[����U��!�ěo�:M�a�V-$��#!H��!�$��W��1�'�@�S�d�$�!�ж[�ZMa�7L��@��#�!��ܗd��nM6R��8`v����!��N�(|��e,�(�EƜZt!�dͤe��H�mK���TD
`!�˴b�H4N� ͈ir�Ғd!򄑢3�<q����'#�"Q���.;(!�d�)��"Bj�(?4u�X�:s!�$?!�By�
Ϟ[0���럮x{!򄚖	�&���*�e�j� �
��n!�DB�n�@�E�W���H���u`!��[.~p����� I��� �T�S3!�Ė4��=k�AU���E*mR�{�!����JQi?!�q�MP�!�ݟe�F� �Y�<2����l ��!�Q;.d�!m��2��(ԫ;)�!���B��p[v��E���P�I�a�!�$�{�� D�B�tvfP�D�!�d�bL�pI�L�H&��!��S�n�1@F�+X˾q8pD
�F�!��ߥ~��9�B�{��S��͜l�!��\l
�K%��(u��h�Ə̩�!�K�B���P�e-�����H�!p!�$O�u��X&�V-[�(9#Ǯ�Y!��R�mEb2�f��|+8鴍�:=�!��G�V���r�k&�IeB��E�!�$$r)��Q��?Dd�e�7�!��J�v�N9�b��']$�5�U��I�!�0�� rThD�	(պWcP�B!�� �<��惥XS ��GŇ*(��"OR�P����bD3��8~x� �"O��X'�ܹJ^�
d��y�����"O>\�#�Y.g
�$۳�żH'v���"O�9#HJ�z�lYIA��q�"O�lUK�i�`9,	��9� C�yb��1x�ҕV��6sb�H�t
щ�y�� Ԩs�#W!iR�Ak��@�yR$a��{4�>]������
��y�d�d�)�f�Z'@�ҩ�T�� �yrj�Y�u��@�97FB�Dm_��y��Z5qL� `�֠���a6���y�㛊_`���B� FHH��ք)�yҢ�3m+�<a�@D��H��h�
�y�("t��)
�CP�4^���Ua��y��"fɼ����0��������y2�3h�E����)2H̑R�ڽ�yRk\�-`|�#gT+N�Ċ��/�yr*�Vn�:�ƙ���y�le�\�G�^|�*Ǡ�y�������[!z]�������yRBR�G(~��*��h68A����y�
tq��P*[�cS:�����y����.�����D*�rM�"�y�o�'D4ӠM�==H5
�$�y2��:���ۆK��
�Z�٪�y�	ьI:x!�G�U)q��A*v`���y�"Ь���g[�8�$L��y"N�E�:�s��6c=��4AS+�y�j�;j4x�c�`�ne�Fo��y��A/T����UJ�[9&y;�i��y��Q9$=��8U���W�JÕ]3�y2H߸�zl0�톭P�6�+����y��8-C��H	54�����jC䉅d#h ���
KB
]�񩂉?LC�I�C8����C�x��0Rm�]�FC�+=/n4ӔkC|��((��3��B�	�P[4L�G>�t����&n*�B�6]"���قl� <����Z�|C䉻d�%���ct�}�G��+HlC�	 }$8�b"�X��q9�G� LhC�I"/�� ��^���Ui�
ݍ�4C�ɯ+��1�В���i�Jۖj�C�I�*��(�!�?���C�3��B�	�A܄�I��X���. ��B�	V����L�GqN���㛂�B�ɪ����)�6uZ{0JZ�h;�C�ɵ�Rxb�� �qJl�R׀Y5ZVHC䉯�L0�0
Fj�`��@/�?t]C䉥=ʼ�N˔;�<)k��#I��B��3"�I�%,9�6{�'UB�	.M��5ۥ���'WNxT*3Z�6B�E>>�y��}�2������M,B�)S����U)	������KAO�C�I�U��J�J45N��G�,)8�B�	�<��Г3���8�@��x�BB�ɤ�P
mX�b����*-�nB�I���q�7H���FK�&�|C��.X��
>I�Ჴ��'
�\C�I� t�ic)ݣl��MQ�Ǡ��B䉎~dv��
�0>���7�ʽ|��B��%e�pI���n�&�H��	�N!xB�I�l%���@dB&X����a�2K�jB䉈N��B7@�ƶh�0�Y-zc�B�)� ���@AX�����cY�gz��A"O��q����|`�D� ���"Oڐ���:]X�#!�� pa��"Or-R"L��r����Օ��"OjP���"	��p�e�3G��J�"O4����ŢZ�X�� V�]!pekp"OT-Q6΃k��P� .S�v%ɳ"O��C ���3�:h""�V�Fk ���"O (�KN������hjA�3"O�t9���M��% �K�DU��E"O�uZ!$�$����*J�W>|q�"O�L���$h�N$�D/�"08*�Z�"O^1��H�4m.*���Ώ(v%8��"O�t��_z`;�mW� n5Ca"O��@Ӄ��+�j<��~:J��$�&��0|���A(p��ͱ��]�@e�}�<9!)T�5�M)S. ��&��f��A�<����:x�X�㰠�6e���cP�YS�<i�@D;t��lÝ߄�˅+�Y�<����oų$_�mz�D;�oAS�<	"R&f�z�㍰
ưk1 �M�<����M�*,آH+8�� �
K�<9�˟<h� � �+
�@M. �G�<��)Χ��4�%<k�!�%��E�<!rjP�Tf~�r��G��`aNZi�<іoηV����h��[��9���c�<)u��/+ �Cj������^�<�����*V����[.C�`�� �`�<�d`à1�ay����ы� Hq�<��ѽR��D�-�v�v���^Q�<с��OS��A�a�.=�q��W�<�r��1N��:C��nX��b�ƆS�<��!�0?�MyA��H���g��R�<�R)L5t�{b�W�an ��U	 N�<�g�����@��[�H���JV��_�<I�ρ3�(ٶIH+Fz����GC�<I�g[4IT,�u�٩W��8թY~�<�7+¼y�:��dBQ"J�:��B�<�s�i`|���Q�SV4�A �I|�<� ��:5�*�!R�7����A��x�<A��\D<T�4ǂ9?~:LyG%]q�<��*�9o�@�C��G0�h��g�<y6E��<�2����9��#�~�<��"�7Q�bܓ�Y�6|Q�+�N�<4B�_R�U�H�� _��"�I�<��ϟ;1=��i���H�����]�<�\�8h�2n�0�CUB�<�&�����Ɖ�yڑ�c�@~�<i�LǼUф��$';#FI�G%�b�<�Q'��z�x� ��F�rrX�:�
Z]�<�� ۗeq0���'T���^�<���K/%�b11�!Yh6�"��\�<�AV�]K J��"����1��_�<��G1��Qd��"}b��r�U�<�s�$��UR.��%�vm{�o�R�<�Fǿvf�t�J�!#H����XN�<1!�k����T��1/�]�g�Of�<y�hƟ%�lA��i@�"�vи�(VL�<�i�#�$@3c��,�F(�tD�N�<����Z<L�XǞ�O(|��c�<��ʛu]�
�䄽O�Μ�b��W�<`�OL��R��W5d���G�l�<��My�n�sEV�"<�x2�AC�<��=p0��#�0
L0T�<� �2��fW�Q��Ė|U�0I�"O$�
�J�a����uJ*Ѻ�"O�)�f"�E>��%��K9D���"O��#�V�_� ��!ێ�\ݻ�"Oj�-[�O��F�ב �p���"O�P�V(�M�Eڳ=E�J�94"Or���mC�)���7��=Hή�Ha"O`Y��E�3A�TNܲa�z�A0"OB�1�F��؋���U��:�"O���� �DtC��ƙ�B�"O��yS�}m��0�F����0;U"O�\`�[���[�M�P�B�"O����]Kߔ�@�D�ں�i!"O��3ϓU^����ү3ª�"O��"�GԔ�ce�%�a�"O޴)U���>�s�A���m�6"O�i�5+!TTq��Y`�d��!"O�����΅3#�=��C2�B�`"O^����3ʖ��6�J*�>H�t"O����Q�lH�1��܍W��I;"O�LR"C�v�z1[a	B�f�p"O,J�,V�#!�d��+���X���"O>듦 ?6M ���kU�C�����"OP��ą�2F��E�l��dՆ�P"OX��]�	��p����i�t5;Q"O��Iu�I�6�"Q(�KS���Ȋ�"ORe�4���x�H1k��Ez"O���H�7&�����#ޛZ���"O��׭Y�T�D���I�qmT�"O��6jF�"����.f氢�"Ol�e�P.�d!k�CϽ{]���"O��Ӕ�Ԑw/&X)�c�>)$�0b"OlH:q)הoR��D�S�4�rݸ%"O�5�!�I�+#�hi�֨R��H!�"O��a���-�= 6�28M��"O1��oS�P�.�"w�	�:�4�T"O
|2T`��I|�!�5J��6�+�"O$�;q�Ɩ(�����;����"O��R�N��n�؃q'��^�&tH�"O����Q��A(��Y/1��Y2"O�	i &+���߫>��ố"O\���l��M�XU8*��! �"O��)�*X�T��:]���`"ORq��l��=,0��Ŏb�z���"O@����"{�N��� W rH���"Ob9�r��^=6()�Bֹ&$	Ȓ"O4D��є$����+�
��H �"O�e��n	�K��:��3TLF� �"O�eq���=�K��̢heB�a�"O|a�3DQ�d�,9��#�� q���"O>(J��*IVĒ"Ɉ"p&8x�"O�=�EL��*�ʀ �k׼hܺD"O�5Yf�G$`N�p� A�v��l B"O����c��j/��X�/�1u�څ*&"O��qЭ/C��d�oĤv�A�p"O��y����v��5��YsJ�sb"O^@�/s���y1���<lĀ�"O�Ѹ0��&9�i���0�0\�e"O� �r�[�e�zY8s�̇����"Oa2�肨b�b���o�F(@�"Ofa���ߺ�����U>H/��a�"O��@/�y���@���66jq�S"O������V������5<�ᩃ"O��d�\9V��M��,Z)�h"O� n���Z
o�T؊ċ�/���"O(p!����)r�X.c��̐�"O�(��H�gDL1�I�%,��5�1"OL̊2� �DgԘDH�;`ą�"O�U@'��g�Y��T}�����"O`t�� =W��sqeP�[�$�h�"O^q�"��'U�0�*a�5��@P"O���5��)%cS![3,�d|B�"OfĂ�E��Ah�c���c%l)�"O}@�'M<��H�!oHO���P�"OTٲ�ϝ�I�0ٰC�Q�6D��"O�$���	�{eH$_��@!�"O�%	)�;?�p�ZR�S?lH��"O�	��	7������-I�-�f"O��H��UF��@�-M7X]�"O:y�b�@)~����C*7Ԕ �"O�q� `_"��ir��T��zɁ�"O�R�Z��t*�đ�@T&�"O&�Q!�D(0�N}C�c�u��U��"O0Q�O�6!_b@ʶ�̣	���$"O����Z �0}�G�Җv��P�"Oʌ���fU���Dgu�9X�"O8����U�MM�I��W�X���"O�|��쒶"evl�f� ��TQ#"O��CG��hs8H��%��<�0$P"O:a��gM���/�y���q"O�����G״����K4�P@�"O�}B�Z�RI!8E��R���5"O�ԲgO�	~]���(Xn����T"O��ZE�L	<
�`b�Y޵F"OH �FCߪ4�2e
dlP�C�"O��'�m��BLE�]16lV"O���cn�����5�}Ҁhu"O�e9�k�I`�
3@%P��y�"O|9�ꃏCb E�W`�4:򼵓"O`t`�IU�i$n[�tb�"Oġ�$n��=���J��Rp"O\����*��Y����p�@R�"O��
��~�2����P'���'8n���o6��@��?����'X,�!Ũ^�H��-�f�ɵ8VR�@�';t�`�y�^1c6N�.�l���'����qF��4��aV�̽0�pX�'�,�8cΞ�}c2)�V�%�f���'��h��h�Y:�������Hq�'Q�ɪ�d��{gJ��,��]���!
�'��Q���m��	j"��`�61�'�TEIR���E4X��'�W�F��'�ڠ�sB��3zIصč1K~Ց�'_��0
�/Z�vثŁ�4F��'��r!EQ&s��m�0��y��(	�'�h�hV+E�AD�]C e�*t���{�'�q�&F �D�GeB�eW���'(r��ŋ�|���S����`�j	��'�R���.H�4�b���I�U��j�'F�Ԋ��Ə)�Թp'I�LC�U��'?�tp���d[<����LÖ�8
�'���K�,L�y
q�L;r�l��	�'��l�l��FxHd��
)V]z��
�'��qH�̪Kxv�R��6b��"
�'�r1��f
pF�!kS��gf��
�'�~�Wn��w\��㮓*a�L���'$�8�����n�r��!,���'..�3KM+;���J�,�2f6���� �x�$I�@-���1CA�m�ID"O\���3���%� �:
օ`�"O ��ݿI"�i%��3	�(��"OBx)գN������NL'w�t�6"O$Z�99���J<V���"O~��B��Y�x�;Ak�T�4-�""On�/zY�f�V�r�R��G��$C!���]N��&�ǽ}w��q2��:�!�$�=,r$,�eǑ3V��H2nοx�!���m�4���Q��Qb�Z0"!��ŏ:����n���b�I!�	�!�\T���Ά�N<#k�)[ !��!i+�@����7��X0��K�% !��k��<+��A�W�������k�!��A&�uQ8�`�� hM�nG!�$d���4�
|�6�x"�I�!�ğ>-�u�S)��{�T�8*Ў9�!�$�A���ׄ˞<?<9��jW�!�D�j"$M�!(��e�,�*����!��ڝT�x�(��Bk��ǭ՞*!�d��8��%�ri^����E4!���Qǚ�{b���������;J�!�DѤE���wdٟ$�9y��Ff!�d_./��Aȁ,��M��� !�dN.zh2,(7���
A0K�:-�!��Հ|��M�gC����J���#|�!��P��x ��?�E1��0e!�ۭ�6dh�"��p�,Y�'�?N!���*wH����U�9����j3!�D�o4 ���>2���菀`�!�B�R��u�ܻ	C�Z�k�!��*f��4ab ź�
����Іd�!�d#!����Ɇ�`��̠'-�iX!��ȍ�"e;��u-�UZ@b8'!����"'M�0T�&$H��lv!���v�4�u˓|�`��B��l��Ox�=�������z�~��$
	0C���	D"O ٺ�O�t\��Z3q �!"Oؠ��ə�wEA����"\ܥ��"O���غM�J��b�X#t��"O�<cdA<4lM�gƇ&i�m
�'�����N0y�,S܄r���	�'�ĩy��Mb�9i�m�nҼZ�'��9&�ޜqH6�b*2�a��'����F�430�򂐋*@�i����6�o�	�e�H�0Ձ��j�N܉�"�(��>����,-D�L�t�~�Q�dН{�Op8�͈GNV1
7%�
M��u��O��X��R5'�ʖ�J�Q��y�n�,��'�ў�b�,'N_eY׌�m�h��C�'o2Q�&�/o
��X��9~x3�'��10H�،�u�,h9*�'�lL#&�%m" t�) Q��'��-q5��f�ry�Bi�6I}����'(֙����}�8B3O�C�e��'rҬC/;�Q˛	B>�9��[8�y�o_��`���aϬi��;)��O*�;��#}j �V�V�lZtl0/�N5��J�A�>�S�'FF�01$��2�Ԃ�A*	����/O�O?7�,�΁��[��,��W�U�����ޠ�F�ܫS7��sw'�"Ɣ�'�ўtGxrJ�O�^ܠ'��l���2�l[��y�Ի����h��\҅�ٸ'*ў������@1t�eS�7	|9p���.�S�� ъ�!<�p�kWJ�a��P"O� a��̵,�4��%�^I�� #�x�C�����Ҧ�Z;��
�g�����:$�Ȱ4ĕ/W�.DI����$.X��$�Q,\Ur��'�'o�)�s�x��NL��`�@��Z�7ݒIsA0�`bz�}bugK�a:d����G���jQ��f̓�hO1���h�hO�Z��u�3�H^�z�� �x�eB��Xe�=�~� �6��:F�M-�F�Z�'��y�K"C,�طI)+�:�2�ҙ�p<Y���
%�N�{�jQ�.�حIcE�L�p���'�J�d��iצ�
��<X
�'-nD����6��Ȋ!4����	�'��yXA'L�Őh !&�r��1	�'���p�$�~��0l�>�%%~̓�hO1�T� �o�����F9V���I"O�-�!�Cp]s���33˖�(S�Iox�p����6[�&H3��]ohѹ�o&<\���Q$�$L��O�YG|�q�"k1���Ӡ`+ ��'MZi��߫v�` ��	�<!���˛(���ɧ*Ϻ-�x�E�&)!�dM�z=��AU옃7�p!�#��g�'�ў�>���n	�N0D��ڠI��� L"D�t�$V78ܦ�`r!XN�(��!D�$k��ԏ|���>[P�0�:D�,��[+/h�M�E��7FΥR�	<LOz��J��%C�n\��˦5��Ҥ�V?�!��Q�� �̒)�Ji��*ξM�!�dؙ.�`m�F&L� ���ڡ�A1P�a~2�Ol�c��������3qx`�:2�
f�<C\�b<�(�%�2�$ �cm�m�<)��<Ȝ��2��;*�@��i�<��՟*'�Ii�b�B�I^�'��&��h��\��:���>{���b-D����E��w� !-8��y4
�i�O ��)�x��&%5�n)�Ə�|�bYq�'ғ������3���8v�|G�����-�#=i���O�,��L�G)2��d�D��4�'��OԢ}�A<%q�	��@�A�9\���ɕY��݅��a�f0H�� 48'���fڋo�C�Ʉ,c��(��8��3C�юC�I�Z>}Hf�s+�j!�R�D�.C䉴U�b1u�P�l�9׌C��C�	lL�`�
}tlzҀ@0q>�"�S�O&�!�"\�h��ke��Pq��'�qOn���i�HJ1ʵ�
�m����"O� i�)@6M�Ib0iL]�nԣA"O�!�	͘;�&�!'���S�2(bD�D �S�)B!G���g�i�����X�X��D{��v�!���:(fN0����*̪��{����>deh"�&9e5\yp��v��=E�ܴ�x���,̱L�����(c�rԆȓU��,hE��.�4x��/��DІ�(�$�1��e�(됎X*���)���;G(H�@2� �^R�8Ub#$��
���&x�"�D�Lc���C�#�~�'��)�Cۃ,�HX�R� "/�����(On���B 2��T���N,s<mH�"O���]�w��]�s�]/W#����'3!��_�7=t8AoB�>���`��H�!�D�$_��xmʠ3��y��l˿)q�}�������
�9���@�U�<�؜!�-D��a�%�|����+�n������7D������^L�(3䎁�z�Xa7D���
�R�$��kY�>GZ�;2 4D�� �BΜ7
ոu�FNJ�\�yP�"O6t
s&G�X��	Q4-X%S���P"O��[p���B��� Q���V�OH��D]2z���H�<Vre�e/	�!��ʦBo4qҷ��'����FB7{qO�����
n�:�#]�-�v(�SQ�!򤆪xIriYց��(�DXH�a����^x�������w���G�[@B�e8OPJ��dI�i�d��H�]p���\J�!��\�'����� �	��m��m�1O,�=�|⡁A�U����1��i<���'�I8��$���.ƅ;�,�ЦE�f&���#D��K��7
�y�s�a�0�F�!D��8�l�/
ր�W�K�b�&)A�	?D�Xr�
������$T�B�E����<��'�qO�2
��Q��ν:�>���Ġf���$1���  Q��q��r��i�@�R�9֬����<��OdU�'/@<��t�hPR��<��"O2�0@ I�+1�xcDHQ�:�P*a"O��!��ABtH��,**���!�'��'w�K�j�@��"���JA
�'P2ԑʙ' ����b���m 
�'a�A��E��S��s�hTBH8�
�'�0ɘed���h�'n�3��B�IX	�m�� z�:98RF��Ƥ�����	�Z����Ǖ�{����?q�E�IY�!���7g&�����D��&�����ʁl2��y��ڢ ��u�e;D��Xv�Q
_�|Z��F�QJ�y9ņ�>�I���O���$խ0�ġ�	u� �XPB@�r�!��[�n؎����O��t��#	+9v��:�O�ܨ�$H4}�4x�)ڃL0��� "O 9Q,��r*����&!S��c8��hR�9�vE��Ѻ/��K��!4�����& ,�c�"�e=~�r����x� �R�nQ�q��D��k�h���<a���$"L��1@�4+d�ȳ�ӹO�!��	4јP��B9oI�4����'�:�IR̓i���5�.Y����8d�0�ȓDIB�[�BV"+'n�H�	'V�j�IDO9k1F�,^<2i��KY�B7�4p�"Oր�6��0�R �b�S�����"Ob �M
�5��\HQL3R��U $"OH�0e��btF(��(Y: ��|�c"O��h�+�0/�Ѐ��%8Y�`]�"O�M��jƠ7�Z�S@��.��%A0"ObES�$ۖ O��БL��/�U� "O(�Kd�:R�#$L���,��s"Oʬ���C[���,]���@�"OR,P0)y5nU K�!=Խ�C"Op!S�(�Q��UA���~�#A"OdMh&fZ�$�8Ep��9��Ѻ�"O�}iѧ߽f�0� ��1N��ZD"O�a�7�Z�x���{�lM9�Y�"O<�Bu���"��|�P+X�4��1��"O�-˶���,(��#K�8"s.u�P"O��YG�D-T`J�j?*r����"OzI���ߦBwR���Hęo.���"Oxt�A��%HX�!0����Ya&��"O�r��΍0֒���@�s1�<0b"O�L�/ݶD�tY���^�@B"O�mqP`ŕ�~�	� �Lv�yP"O"Y��iʜ@�FJ�X�0�T"O  �&xY��߶�X}:�"O� ��U	�&1X`˗ǒ#M�v �"O88IS+��v>"�0�fI��,U0�"O�9"V��N��u)$Gº8�F$�V"OF 9�d�<v���@[:7�FY�"O 4*�+�1�2���ԕc_�4�"O�5 ��#?�:	��B�S*�Xq"O�%P�	�?`��(��A.�`۷"OZy)� �g�<�p��)`����!"O��J�D�.	��`A��5n[�="u"O���GU'xPV �B�W��"O�U"p��Rz8�H oRD��2�"Ol8��K
�A.��IQ�:r��A��"O��(����5S��D�t��|�"O�9)$A��0�b'I�p���{�"O0ђ�̐�M�<�l]�p�0"O��P��U�M�����+�����"O^�Ԩ�3<�hY�$(���Z�"OX�82%V��T�q�C�(���(D"O��G�5�%I�ȊY�v# "O�t�$�O�4�l��NI}��#"OFa�TO�@��DIc�+ `���"O�Z�  ��iU�b޶� f&�	\!�S�)r�� ���%�����>}!�d�2cA�T�%.�
C�B$�a�?!��Hm٦Lxp�<`�F�{���!�ד'"�PsH�Wݜ��b監Z�!�D��Ag� *  ������ �j !�$�y�tz�N8��Yo@š�1l�A��Ӹo8��(�n��y⡉9Y�y7YW�mѣ�yB�]B�L
�C��e�� �=�y"c12"h���0,,���e��y2a:7��ȹD��'9������y���m�8���-������yb&˽�jM5M�<1:��f���yb뉽^4��H]
,S.������y��7]��4��D�1^�Bh�P%�y�ET>-l,PȖÅQFI�g�G5�yro֪Z>����'I�z��ŉ�3�yr�ޣ.���l�%�� BE�E�y��.5lP�Ƈ��$�,��7�,QJ:�B�F����h��ߨ|��92�k� &�,�C�O�!�$K	F
�:lD�8����zH�ݴF���-�E�r��	$��ze`�!�`�	�f+JE�z�8r��J%�ƭ�~��Ԣ��F�(KalH��y�#����jg.�B�2��B2˸'��3�a�l�f铯6�`���oZ
]��$��bA�7��B�I�[��B �I�GD�h�!"6��څ��#ʒ k,O���Y�@��mµjI>��bd��%�&C)D�8�e��E�@q�ʧwFT�� �Y�D5 �D���hj�^�H�A��>�����¯*춱��*9�l��0+�h�r�oڻ������M'	�����z.�s�<��j�v���N���+���Kܓ{L���t��$Q���`���`�`r��1et��˦�T��!�d%+�4����&< :ʓi�]�L��� 9K�i�'er1G�,O����ƌ"�R�JЯS�����"O����H��fQ�14���P`���Q�i�9���J!��Q��I��(��Si�B��a�g@W�i���d��zp���&|�c������#"/�>i�)��O&D�,C�~��K%�Q�@�N��dj$D�� D�Ρ]Y���N�<���O�ʵeZ* �&�O?ա� �9E�����* �t�>Ա�O�h�<Q0d�#E�2l��>#><=H��l}�![�r��١�Bx���"��9���%�"����@.:�O���V+�8k>��� ���r�.W�j���O��R�8䀑�LlH<� !4���3�EIےiD�Xn�'ւ���@�#1�������(��L� � LQbhiWI�>�!��ȲHx�R1[�7<t�󓆗�;q�$��"��*���yy���'(MX�@E�+�,[@/kKX�<�j�`���DWN'(	��N?�ՠ�5!��LZ�H̰<A��44�峳�N�,5��� �HE8�܀b��$ȱ�S��%v��2��v��@�4�Y�ē�nDb��ݗ):��
!���m��EyB!���zl2�\�+8��M�,AU�آ�Y<|Xl1�"O�\1�R�[p��Cs���]R,��I,?�+��<E���)� $���4���5*��v�Ʌ�T���@c�[�Z�d���"���'�6Ųv˗�:`D���	?v]�H�e�5I3.�Bs�C���������s��m�`�ե֬U�N� ���Cf�C�	s�� �$�تښ9�� 8�C�I~��(P��}���вq�x�)܌�	�n���R�x��צ�F�ء��I�{j�B$\�غ�IV478�.U/aDN�Z�%D��Kg#G�rtP��(���9Ԧ �ɾ>��<���:z2�M3̟�v�)��.ɪ�t�^42���P*^X�H���$t~4�R�Y�bt~��6b@<��Qb�{r0�$���I��H�R��kM6�~bÒ[�Hl���[�"ʒ��l��y�e��Q����/��&tLx�ǠS<�?e�
+�n�Xg�6|6�[����?��O&vHp�瀳~z���
?��d��I�Au�͉�E�\��9�& M>���-�,��ÅT�"�x�R�|����N���� �o��4k$���>x����U��3�.'���K��P�l���E7$�`��h{��U(/8�5�t�Wyu�9�h 7}哌_I���̜����H1��^����X��؅�ahڎT�h���]�*��!��3D3b���C�m�<������Ǽn�2����.���A�B;jĻ�ꂘl�>東<^���%N�{��1°k^0F���Dކ1E�/Z�jQ"!�N�P���x#�U�l���S�@�$��8[EJ[�7�P��fOʺApQ:Q�'���(S�T�j�{�0��ʁ�H!`92M)���;庄����>�z�2ٌIY�(ДG:)��� S6�	�����H
��v��8��
i 1��O�-PW@[��6!���|�=�@]�	�����L�8U<������䦭{�z[��rg
F�7��T�� 8���ge�)��Iү�T���C��11���jZ1D��
g#�>N;�q!c��B����D�03,��J@(
���#/��a�sc�H��*M�P��6�Hza6���z ���`�O $�~�F�l}���t�S�Y2���u���p>YV+�$P㾈A���#j�
�)��x�\=i$�	;Jh�f���A��L��(�D�@������Ğ�UI�K"e���te��DM@1���J�J�4i��(O@Q&�� @GV�"�!N�F�*d��fS�<`�`î.Ghj'�w�����֖g2�o��,�u�F$4>�8A`I������#Xpxl#�����4��,n��(�U��$5?�Ͽ+�C�/����ҕD2flKAB�m�<Q�(Ʋs%��)��<0I�MK�N&�h<#W�Zp��[S�#�"H�'�HO��(7+[�z᳠(�38�2z�'��4� ��&x5��r�jȴ{�2�Hqj�4|ր�Gg\�!��d�����a}�6r
Kŗ%��d�C,hаEy�fr ���Д#��@�v��i�S I�����
a�ݪ"V�h��B䉊F�0�Y��Z�B�te�&�A�Z�֨`�h��ay4,�ik��
�h����5dA�s����P,jݸ�k�)�y��)y����'g6�؀Wꐃ4+j����ɑ1��aJ�}�p����@�q#�& t���,Ta���*B,+�OPA�$ؗk4~�8VH�#^�����C~��q��P��M�#DK�5�}�ș*gQD�1�Y +֐�T�+�hON,R�j��r�Xvh�4&5 �'W�����ݑJ����&ɜϒe��y|!��'�� �(5�$�_�B	�I"{� P*Mw�U�Qm�@�O�b�:0�!&���2I	�;�<�"w"O���/�)eڄ�;"h	=�H2�l
��~2�]�@p�X�!�R����� e�t쑁��?��J�ы.wl����@ɬ���������&)$	W蹹c(��/������6T�ܣM�
�hH���ax≚�m�T�=IP��;���Cޢ��}k���B�<�&h���t�Y��ܚ�r��J}�<ِ��e����T��:��8��+Tl�<A�k�Iy���b��!Mt����L�i�<� >DЂ�̤?=�@8����~�U"O�A��O���+��p<t1�AE�l�����Ox<rc��R�R� �҃yu�y3T"O"E���I�Ro�(+�*A��H�2�>O��	�&ϳp����B	z�z��� �U��d�E&)�{�,X�}"��ɦ�#A��Ayz�r %U�z�J�
,#D�``P�O!0q$���
 ,�$�!���G�4�`�Ϟ@b�>	Y@�I�I� �҆���Gf#���` ��i��@'ȭya��(�hA֍�x��Y�ݙB��O8�}�exz�i�F\")�d�E�Wc` x�G�TnqO�}��_ՠ����Z:Hq*ĩȯk�Ե���{<���e��&@�a{R��(TT�X`H�,��D��,�	�?Ye Č �>��8�����|Ӥ	���+ra���"F�W0�h��'fj����g}2�X
0�,��D���"��@������'2� �/G�fQD�$M�pZ���ń�/'�����!K���'Q8Lq��Zj�OVhYݥ!���Ao��W��+A%�V��E�1b=}B��PS/?�Zu`l��F�	�Ξ�6���È{B���MK3ym�EW�� t�fE��k�0����s�.	��I�e�H�P�R#62������Vn�	�.=�቗E��2`3O��u 
Q9��ƍA!�*1"O�IH�Bܙo-���"M�r�
��"O��h��4r)zU��E6��"O������P�9���P%ڭ�"Oh�adM�n�,k�KI�q3"Ot�k��2QT���U=.		P�"O�����Q�N��G�([�m8�"O:��虸Fш��ǂ�'����P"O�t�7EԾn����\"�� j�'@�����ff�Ɇe�j$��H�'*�t�1A]�l�^�)��?S����'0J���L�2��HF�e�����o�~�I<)���;g�	9 �iȘ:D�]�<�U �G<��$UlXb��XF�m] Zä8�)��\� P��aP?z0A��[	A�B�I�)�T�c�֪�0�sK�2���䍘Y>�S8,AD�Ǧ�:�����97��d1TvGζH�m`0$�;��ycf#�dp����Ťg��L�`��{�(����a�az�L?
f�O�e��g�^��"���jS�4ڠ"O�l�^�G���E
?G����DT�<@���{���'�k�f�Y2&E�$�i��յ�ycP#g�a����%&%��˞�}2�Ћ��<aUa�#S��3��5�{Pw�<y�i�)v\i��M�:K�V�p Z�<��c�VX�)�5T4���T�<vNf�A�ɰn8:qtcP�<�'nTL�Q؂	��v�Z��e$�Q�<�hΒ8F�D���	~B�XJu��W�<a��8|�0�8��w�:�BV M�<�FI�B��aB��tC�Uja�a�<���K�>��u�q*�)l��Ka��Z�<��n��a�P���)|]؜�e��M�<i���E>D<�2l�?��m�/]f�<�f��m���PT'W=9��*��k�<�" ����㦊F"28k�z�<��Ή"l(Z]Z���t��b�w�<���ɬj�J3�9ݐ=�4GH�<��j1>�=("�K�lp�KG�<9�n��H̰�O���kf$�A�<����/z�����1+e����}�<�	Y*�6�����6�5I�V�<�3	��Cp�(�Qۿ/���(�Sk�<���X�U��@�YW<��rN�~�<!�AM]wx��	ĨT
2`�R�<� ��Rqe¶��CN���@"O�0���1x &J��ڱ��"O�=X�`_�$H�+P��8�"O@iKw	D+;�4x�@
</�(YIp"O�A�C�9-�� 8!���
�+"Ob�aT@;ϐ9�s���P����"O��ʧBI+<DCU�MO$��b"O�q2�o��jH6 ۝`j�*�"O�z���7$��LcD��\	�V"O�!�!C t���⑳b$��"O&�y��#P�9���4���T"Oʄ��Q� Hs�Q&#�Ll"O�ؒb�]/P��h&1�B��"O��ɀ�j$l����A�Z�t"O"�9���/�M���F�c�$ٗ"O���0�!;I��3uJ�?]����"O���,��iX~���)8�Б"O��вj�R�(!⇇9H�3 "Oڌ�D��_�
��Vƅ��V<�7"Op�j�(I�!}�*%�B$l&�T��"O�����������l yط"O�xv- �m�ff�"'ŲW"O�$P����{F� ��Ä!�X�`"OdBv������^, r8f"O.L	��T��~�."Vv�XPS"O�X���2I�z�C7	b�|*�"OJ�X�dZ,b�:	ԍ� F�ѩ�"Ozi����^��iSmG�	���"O�ԙuj��V�t a��_&��3�"O�-��%:~�bq�T1<6f�"O�!��wY�Ͱ%'K�Zq�hK"O���A ��_���FT ��<��"O�Pj���.|R9�ৌӲ��`"O�AKv揯
����V#�VQ8a[r"Of����
�3�蹐���qW�<(�"Oڄ�F�msX����N���"O8E��O�\4R��,N����"Oj9�E�V��$�����<a�"OJ�J��}�	�0-�=˰�
f"O89�!��"3�]��T1cĜ�"O@�!��2G��H�6�\�$�:|��"O��1��ʑ<J�b�G�mf��@"O>L���DJP�5O̹\t� "O44��j՛X��1��eS�+L���"O����У2�)�r��3i����C
5:C�|����#Eȶ�b��ķH�l(0�$D�����*2�$����>~��9�RDl��trf�x:��ߓFu�u����:����۔Z�\��I,~0p��FEֵR�m�м3���rx����0��B�ɉPF�Т�努W��}��I�$��XI��y�Z�r��U�O�Z�O��Zae�S�^�C�'�P�C�1a�.is�i
~~i�S�D#?��8+���<���/�gy2$M$sn4E�D�0J�����#�5�yꄃ_�|�\�}�����Դn�J,��!40���J/lO� �"2!-��B�t�|����'�4�Ӑ�(� e"�i�E@�D�<���R�Ϗ�xthQ��'P����Uqm�4�]8dR�h�{®�6#v���`�=u��>Us�T�y�@i�$�'���	sm/D��y�.;|�� G�8����Am��̬��I� ��5�(���n`���AbĄp���0�W��dC�ɺR�p%�B�Km$�@�/P�*�6��*�D� )��=9��ȹ{�`|r����en��a�c�u��LH�f�W;�]�E��;�̐;T� 4�����4��Q�҄��"m�3&��й��S�? 1xu/4SNA�S.�
J8T2�'F��R���;�ɧ�����5(]��Hh2��21x:`�a9D�� �
�*Or]P҃ϓf<�%�G�>��k�y� �!1<O]i!��8x�ޠ�`�=�!���'c�3���DPVܠ�OW'b>43�N_�h���x�FU{�!�D�2klj� �/� a�=�Q��qM0	aD*���z�' ���&�[�yԚI�eN��c�v���*%�\��!�1,�%��[�:�P�rb�=�(� ��3N��)�������|O ��oE -��f%D���/�y�|�xD�G�z��奟����Š-0�Up�˟~X�����M���1#΅�anH3��5�ON���M�Q<���' L�HEUP3�����dM-&A��'��E�M�./���ꓨ��u1��X`��m�#�,,��b?��e�K�.Z$l2��Ϡ?���ӌ(D� �# �'�Y�L�޸Ã��< X�I⁎���2(O?�d�$^�ZH���=/h؅¯+A�!�d�ML�����3[DR�F������r��3i6�y2A�+"��L���<(M����W#��>����#u��*"�ώ&;����!��3%���y�݁<PA�JO�:�`D��y�D�}��A����To(Q5�ז�yrO�z����� e�P�e��y�I�o }�����d�+u�;�y"nI;K���*e"	��,�ٔl��Px��� ,n���;)D�Z����F�Fi⢆�Z����R�'A�"D[�e��}KD_N8�DXÓ ��9�o�"`��d����%
EU*�X��j�nc1s��*D�C�D	kT$8���-t*��5+,-B��ΟJ{pp�#IX'K��#������V���Ի1<�#׫�	=Aڕ��0>�Q��/F�(�i3J��i��]0� pp� �T*Y�Ne��_�������X����շk���g�~�hHtmG�U����F��$X�A�OtM�͌'I(����o�����p�����IJ�z,�b�a�T��RеG�<��F�ʓL*�p���)�����ʾtȅ)T#
#>YkAn��0� �ʅX�R���t���Oȴh�E�U $(a3ю����N�c=Z�⥈\H��:��8���34U���@L(����-�:�|;Nߑ�8u�2k^�K��3ǳ#��%�@,�ǟܐdm;�d kb�_�|2fNI�.��pqGˈ~�4[GUV�'_�\�cmE)%���Q^��+e��?ݪ}��"T9/�tʦ�I<Rm�S�[.ҢΦhP�qѤ#T=��3�	.Hzh�iH����@VF5˓ �DL(P��Zx� ���$Pz2H���)��,NthB�� 8��|@��C�7�dq�q�S�w�ȹ�HK�V<��D�i�����VS�� �jݠfqn�ѶHσk�~�`*Kf��=:f7��ؖHQ��(iV
\#�~R����*a-^�M>������?	m��^գ�K�$���	��O��je;GmԿY�>9s��s���j0LV6r�D˓sfȥ�c�A0X���(y�����K2N#����i��s���?��"-t�,�G�'{����f�^�}ڰ�2(�o��E�PE�4 s��R�M�A(<� ѭI�Z
�KM(hJ\Q1c�Ojy"hD/6��5A�́?�|	Xd+��W�F��~���:.7�����B�����.�Y�<�����P1K�N:b2n�䈂���b0f��U�g�v�
��JG�	�X��ԡ�� ��D��F���W���r����tm��u)*�XBh�,x�jC�	2R���c�m�#�-{'&S6�C�ɭ7�P���G:]��A����8n�C�2fĥ)v��;;jN���K!r԰B�	0,d 8 F%ܫc����6��1bZTB�	(W*�ѐ�B�P݌�7k�*d��C�I.yJ�A� �JPE���ğIcC䉐-�*X(�g@�%�6U��4��B��?��Ѣ�����R�^	��B�	%m4p�)���>c�ؑq�݁�LC��(K����!9?,�ZH��SdC�	1J��1+�1jw�\R�o���hC�	 �x���"�I��
�L�!��B�	�Z��2Gm�aF<4���=J�$B�I�c~X܃�Lz�B�b�
�W'6B�I�o=9᥎��t�K�
G���C�)� 6<iP��w|C鈷T5��i�"O���r�\7�6p8!)[=s86�Q%"O�áN�*,�T�ƏYC��"O�|+��R�RwH�QZ�C��c�"O\I	bR�&�6%���04�11"O"�b0��P��X�kǂB�]��)�)*�����O�]��j@v��Тi�!?��e��"O���Z�,�j	@�b��w��p�0O����V($���Z*�HػP%��PLjR&D�1��{bA��%bL�(3���8�i�<2�(�W��0u�Ҹ��g%D�����0f䮡`�����p� �ɗ@>90�,s��Ɂ?1^-��K"8�$�Q�N�j�!�ě�EBm��˾(S��Fb�:?��D�Յ(Z��Oz�}����X�`��r~�0u�I	O��ȓ,�f�{ЦاK�9x���d��I;j�M�tAXE�a{�lS�z�P-c�ρ���d�` ����=�`o�	
��P�,sӔ��U��U��ÕB?M�q�V"O��`�f#~}�3=�2��`�dY�0�A	�H��s0$	�bĥ�e���N�І"O>�
�HG?PN]�&b�y����C��z�P��U�$6�g?�5k�����Z����A�2x��Ke�<YINX�hbƭ��-�����<���ϧd����
�i�P��r( Z��X����*shh���>�ı�1O�!"�F��������R"Oz|� �V2Gw��1fɎ~�4� "O:\�C�O�d���5�[���`��"O>m���\�̚�(�Ă�1�9 S"Ofqha?[p4��"�{7dRR"OFMSEiӌ+��Țt��1A=��;�"O�����^3-��p�p@�+�0��F"O^���f��"q����Mѧ�y*�"O~�*Z
Ep� eW&H��"OF$ꃆ��06`�� �:_�& h�"Oʹ�ѡܳ]��8�.,[L��#"Ov��?�D�1e�<&1�q�"O C��B.�s���%_ͬ��"O�A�"n�.��i��54�V�I�"O�T��>�nܰSLGL �"O:ѓ�)P�i^Q��ɍ�9�v*�"O�`{S[�16��bF?����"O��8�J�6LH���	 �Ȁ:2"O��@�E6���g�݃/�jl��"O`Ĩ!��114������}��,h�"O���RP�*��)�!u�L�t"O�m�F̎0n<�uf�{kZ �"OvŻc�V6�\{f�����2W"O���M�>q�Y�b�ђ!�<��a"O(Xf�J9h��5�:�,3"O�5�u�	j�V)���)&:P%"O��`pfıE4dx���kϖ��&"O���dA�7���2�]0(�\�1w"O��v�h��Ѓ'#U��ҕ� "O�E��I�<{�)"U/-�TLs`"OP {���j��  `��Fp�9�"O,=�ׂϘ9�8xiW�@Bur���"O�d'��	ؖ�rP?Hij�b6"O�i�ᡃkW���2Ͷ��G"O�P	�N��N�t�q�W�I��h`"Of R��	�&z�	3��F�{�
��"O�aV�ɢ��PH� ���K�"O�E2CJW�>�xm���.Gw��"O����Fބ/���UIֲ1s\i��"O \ʔ	
^�n�CRj�j1"O�L��C"|��L��C�3Rnu�1"O� ,��i�=u�Z��B�=xZ*}H�"Ov���L��58ș�ƇoO>=�2"O��3T�Ќ5>J�#�)/%<���"O��aj��	�Ti�ǈȖN��<�"Od	b7�L,p"��ѧ�ܕtz �W"O�yђM�����c���+j�X�"O�����^&�`c��x0N�q@"O�5��B��Q< �Z&�ӅM"d�Z"O����+��\ǨtzV��/'*ijs"O��J�T�2'����^�!�xz1"O���̊�	�h�q���/P6Y�"O6aS1�Nm�&qw
ߑA\ђc"O2���:FܱahD�L0��"OMR��=k�܊6�J�j�v@�"O8M��,�p�5��E��"ɸ�"O�H���D�Ei�JG�.�be+Q"O���A�oi��e�N��`�
6"O�D��Ò��8I�C� eT	��"O�e����4��PbDl�sEnYbv"O�u�	O0Cz�|�%��'J�	(V"OH���[�m;��h�%L�Y8lЪ�"O�,!e��\����Ć/GZɹ"O�܈2��F�t�R�#;.��a�"O���!I��u�8���ßg/����"O��9� �\�L��O�)+,a "O� �p�p)H7I�m �:�"Ol2�GG�^2�Є�G���HC"O�lJ��I�8¬43���i����&�&$~���
�s~�$��(���Ӗ-&��8�]�䬐��ϱ:��i�r��c;���-O�<�O|"47O���Ov��D拪+�&|+td
>�&��AOe���')� �D�?��Ģ��Xv�k�c��)r�����ZA�u���s>	S'�D<5@����=d�nuѶK3}2iC#{ɠ��Mצ��H����Q3@�4�����B��@�O����G��T�>%?�'B$�F0f�1q�%D>?�$�b�4D��� �⌵&o���/O�?��R�A;��u��ػ^��<���/+d��`
����L&�)"ҧ`��M2Ԍ��+$ ��P-�;T�ulZ9I��$�O�����O��sӘ�6��(�VA��d���B��i�Y���(�TO�?�R��<�H�if��4j�B��J�+��I�s�$�ĕU>��QlY�G�- �G�����I��Ĕc�ā�i*�Zȹ��Nܪòh;H�x��V���5�p$��A�Z>FL��Ș���� <`���]�a��䜶n�#�H�a�+�kq�Qf"�"�4�HDK���y_�e'�(�Ak�D���çU�4�7.Ջ~�@U�擄jF�Xe 	3~�P���* m�)�' �~���Z��n�{���;
{L���ǘo��a�Y��9��OlZ��ԃ�u�x8�S��r�Y��'����d #y�{�&�
k��m �'�
q���[�Oʨ=a�� �f!j��
�'�F�j%�-�h���IQ�Q���y�'�" Z&�[?x@C�g�'z)�s�'�,���U�7�|\�L]/R�y�'y�4�"kCo6z�;�NM����'/���W����dAfE�0,��'jvP�,�0s�0qq��N�e8^H8�'�R��0}�~��g�ۼJ�p��'�: �%f�58<�a�O�T���r�'�����Ί�U�=Y�D�����'>��.�`�h�ɽ>��4Z	�'��ٙ��9��13��	8;���'�^0 �@�#����࡜8-��U*�'E�bH.)WΠ1�	�8M>��'gx�	Gn̶$V�i������Y�'�&t���͞E���dIΠ��A��'�,���ZFU:X��!̄����
�'On j$*!%4չ�N�LPҼ��� �� ��� _��*P�9{����"OP��3��Y�Z��f�U	z�� 0"OzM�4D��?8<�\T��*�"O��k6��`�MBc�ͅPJ�D�"OJq)��;=���/;p,�X�"O�!��7~hi3�n �yH�"Or�C� I����S.D�i�l��"O��Cfj�9_,ez��j�>���"O�jE��o�V�C�
K>�zS"O�ሃdȆ?��8�䘍Q��-i!"OBD���ߤP1��aj�-,~�HÓ"O޹�t�D>g����:zk�(0"O �2�Һ�&�P�oMV4|��"O�PD'ؒo�`@	�n��80�Z"O��B��Zm|x�!��#Н�"ORE�U�ћ1�ތ��J̲�6���"O"���h��k���:�L 5R���"O�A���w�A*�o=�0��"Odl�4`I}
��
��y(Z0��"O�1ˆ��`�����B	h22�z "OD�cu�ځ-��4 0aґJ<`�"OnY�D�/�V��בr
:D�`"O��X��\�	�ҁ���(p   �"O�-[`�݅a��2�J氨s"O���6��*c_��p5J�)���P"O����9�l q0jv]P�"O�5A��$JO�Iqc�!dZ���0"O�1¶Ҷbg�,��A�$\I�\ˤ"OD0�A�S��� ���]5��z�"O"ic�I�1 �Y�,�,�m�B"O���X�M��i��i�3av�4xf"O
����;@ob���G /l\ր��"O� *�d�Y��F���<��mQS"O��V$Z*��B���v@J�"O��!�Oӗr��������l3va� "O����Kb� @�ŉ�%yJ�� "O�,�PI����HՉ�EbXQ��"Oĭ�f/�6{��5s�Yd)N;�"O�|s�RI�R�P0A"��"OJ�9�&��P��4"Q�+ x3G"O�}k`�R�RU*�!�;���#Q"O�=�dC	_PT	S%;4����"O�$���١l
�%2�̿A&U��"O*d¶�Q3Ҕ�"`�>&�=IP"O�I{G�3�q��;! ��r�"Or��GHV:��B�Ǻ'��A�"O��5I8e�Z�3��~�,\�"Ol�� ���
\z���9���	�"O��!�ǹs�>�9w�H^J�Ū'"O��@ĳo#ؼ@�
^C�$��"O��b0�W;��p��w}.(�D"O@��"�ɒr��!��3_Z�M�C"O�`Y0�%[{����$o���Q@.D�p1��СM�|�a�C��b3����/D����A� Űg�B�I��{%c9D����ə!H/`��pg
$�DYa��8D�\ڳLE^
�|�tF�"E��
�*"D�d�2���7��$� )U����("D��Q�]?j!�WD"j�%x�.D���cc��h���Ui����d+��,D���gC�+y�4SA�v�[$,D� 0%ɟYApD���٭Bt2}�s/=D���5*�qy�Ī��53���*Ӂ(D�x�5��lp�MyЇ0M �ZW�8D�� ʥj���Eo.�s�%J�8<�"O<x���1"�aA�
��9��qpq"Oa�C˝�o�FD+�AR�"ܣ�"O��3�.N�Qp��� 6.$Ч"O>��lO�@���6 H��)�"O}6�Ia
��!��/�JA��"O�\�kɡkG��2ӦɴCKb�{s"O2]V���L���$UK��I "O�Ƅ�F������;e��}D"O��1�M5�*�Ǥ[m*]��"O>�h�ص?�X�9���!-x��h�"Of,I��@h����#-\L\��"O$��`�%E�@;��уpH�D�!"On,�UhZ�kC��H�ƕ�n6��"O�Hq ��;s,���E��k$�j�"O��[dC�ݠ,!�@\��r�"O�2$��eI���p�T�$��QCC"O��ҳ��*�͚wɔ�d4�<j�"O,�ZN*ea^a�����=��Q�"O�t�S�vyf��牖�{�V�C"OPPЇ��H���R/�v��"O�z���^�)�w�ǀf'��
"O�
�H*���c�b	z2��@"O�u!$��!g<���G��t��e"O��(T ^�t����o͉1��h�"O ̣��,�8$N׭&�H��t"O~��$E�-+��K��_�?�	��"O"�8�)�)8a�b7�΃p:�Q""O*�C�A�=�48�D�;B� �"Ox�J�B�2
�N����t��YC"OƐ�W?(@>\Z�ޤ�l��y�F�h�!�ԋYC:84
@�y���4?������W�MCS悫�yr	C�$��˴c����]��윸�y��'�d(���^��uz�ꇝ!�D�P��i�W��]Z~�(�	�!�$߂ �����D�##Q@��)_!�G�,U�]"t�D��l��EJ��T!�Q!���`ĩ��L�Ԥ�b.9�!�dڈ&)Hsҏ-I���;�&{�!�ː֘0r f�n&�%#�OD�!�$S$+��P��V�F|�5P�Ͽ8�!�$ƬJu��k���Q[��pD��9m�!�$�-�p] �HDZ��!��bH~P۳f�P1��8P  pg!��= 8ᓆ!�2� �R�"k!�$Z�f�%�N�g����Q��@	!�$���Ȅ�FªP�\�s&��76#!�$F�4�\[�ז����ԇS�!�$A�gL	�Iܩ/������G�{�!�ė
o&��s,h{��)b��!�d��S�F�b��`���d!�K����#jO���\�� �>y�!�Ě�O4�m�$u��hT
Ǭ$�!�H;Z�(�:�eA�-k���ܞ-�!���o���@T�oL�k� 
xq!��"Y��	�#��7����,f!�D5��q��D�H6�%�GW�N[!���5Wx�
�J1?lH�e�V!�V�'fڕ�,�=sPt��n�,�!�ǼD9,�AnR�7���g�>�!�Dڅ8-A
�Y�B��%��x�!�$�?j��I+���L�$�� �ݘfp!��ҺH>���C/z��ɕ�_k!�� ����ՆOJH�A���<OL �"OXZ�؍+�5�&T�#(���"O��z�`
�~#D�#�$�`¬�z "O�L�a��Ǣ<�g��d�ޙ
%"Oĵ�G����P�9�00��q��"O�hc6/�?1����J�Y�҅2�"Op]��/�0���#c)˶ELt�s"O8����ԉ|{b `��V�9S��Z�'�R���F��T�:Q1'L��$e(�
�'Y��z�/V!p�NT��hZ�!���'�DEbwV�4�H0��♺D�RD��'�����\�s�L���H� Dz�'��bQ,ע��1Q���x���x�'�h��(B���F�C��h0�'�6��REf���g/�k>��'��Ŋ϶D�� ���ҁw��@	�'���Ԃ	גYQ��Y/��T��'���Q�+=a��X�.W�+n��
�'Z�|sDf��s��hß.r*�	
�'�~��#ڸ57Fp��#� dR�X��'�%�&#�:27��S��_S�-��'O���n]��@j�!Ef)�"O>͋G�Dm�i��dM!p����'"OFL@�b�=B�`��f�� ~^�&"OLuHP�0���$Y�\�k�'r
����փ
�����(�	�'H�ܨ��E�#g8(Q�Mc�����'���-ـ_�Ѻc$mӪ��"O���ӥT6����D�{��("O�X��-Y�I����E�W� �H"O���a��C�4,ӃN�a��(u"O�(�@*�C'��z�L�HW�H��"O:�p�(U;nJzQ�֯�14Z�=�T"O�P����43�p:��/X����"OH�OH?CF�@9��O�VT. PS"O��s`�>U�ԣf�\�B�� �"O,�Su��=+̪�@�S��3!"OX���4p�T�Au 8Z͈�"O��aLQ�V�tYqM�=��R"OJ��K)�6Y!q��|�
1@�"O �I�P0H ,8;�Ӑ:S:M�"Oν0EN������^T�8��"O���A�'&!����i�9m`U"O�,�Ge�vH�����^�PȆ"O��Rg㗭����x�$�u"Oɱ֢�'H�4A�c�����"O"�A� �5 �*AH�ݖO���A�"O�I��͛hNx���K?���6"On]c�	   ��     K  �    +  �6  �B  N  ^Z  -f  �q  4}  e�  O�  ��  �  ׵  x�  ��  ��  !�  q�  ��  ��  ;�  ��  <�  �  : � ; � "! s' �- 4 ; �A H sR <\ b �k �t | B� �� S�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O��jg�=Pz�Aa`�#�h��!\��̇��#=B8#���fB8%pS��H�����fȉ'�$!q!c�	^+F b�ǂ!3�v|��'��EK%�ݵXF|ԲBER�/�f�ٌ��#�
ّ���5�`��'c�6vH��C$"Ox}e��N&}A�A�3Z`X�"OJi1�Hճ,U��I�	� 4Ft��"O�D�tkI:��͠�(A�Iddi��eOuH<YS@҂+2��p�T�w޵����h��\�>y���BdlcL
�g?x<����d�<7�5�)�늁yD	�`��J�<�"]2����ܿf:����G�q�<I&��d�ɓq�:Ρ����X�<񥮀�8TΩ���y\^P3�N_�<	BdJcV�����P2.�"�J�,�v�<i��1i��#P��,+=hR ]q�<���	4M\���#���:�����o�<i���3ZJ���5Y�%ԞU��g	h�<i�-
�Z����&��U@�ɱF�DM�<����+�|�h�O��i�ʤY�h�K�<����u�
� R?
Kv ça�<���.-���4��*��ZVŀY�<��ꈍ[����Se��e:��Q�<�%��$f��F�S�r��TeXX�<��(g��K�GįDlz�iU��P�<�w(]�>c�r!�*8`9K�"O���T�W���!G�Q�R-�"OHXB�X( �i#B��)^i"O"5K!h�5��В��+B
p�Ia"O��Y�Xr�-���,�ِQ"O���j�"�U��-�~��"O&���Ǚ7�l��t,�V (�"O�a 2]`��:G���ya]�&"O2K��ƹEέ�F�� F��QS"O�%�⋖�s�J�y"nԵ'��ۣ"O�Yk��z��i�`�@�p��"ODY�̙<RE��NK�l/2!��"OJ�jv�۽;�P;"�̼#j�P"O\I�/���Y�	I����q"O�D�$j�4F  �H1e��N@b�"O� ��
�/q:��W� �!��Ժ"O깚��
=%dU�f��3���7"Oba�6� "j0]H"�sΑJ�"O촁LTf�䍐ANL�r�4 T"O�LU�]�FP���2�xX�!"Ou���]�9��]ao��)��"O
�H3 ��Y��Qo�)I����"O�u�wƓ-r��@�7c��_���"Oz9T�ȧ&u�h�IK��< D"O��!�5�6���\�f�"�"O��k�eK-fCu����:���ar"O� >��sc���5S��	�C"O���I�8-��4�nO�G���"O��X �].8pw�R�u|�#"Ob�[h>S`�b��C"4]��!"O"-���[T�]!u�v%���Ĉ�?����?!��?����?1���?����?�C��J$d�bbT*v B��?���?���?��?���?y���?ٱ@�&i��(^@i���ز�?���?9��?���?��?����?i�f�	2J�x+�QEr�5����?���?���?���?���?���?���)rev\IQo�Z��=��2�?���?y���?y��?���?���?�� A�7{��9��+X,�ᑓ�?���?y��?����?���?I���?�jȍaBN��3�N����S��?����?���?Q���?����?����?��BL�`\��ߑ�v +p.���?���?Y��?���?)��?y���?��ᖚ͜�C�\�mHP�$�?���?��?����?Q���?y��?�U΋�@�Bi@rdݭn�����A��?���?1���?���?y���?����?���<��� ���m�BE�CG��?1���?���?����?����?����?AR ��d ʽ��  T�6��'f�+�?���?����?Y���?)��?���?�֋Z.1P�u�#PR��a���?����?����?���?��dQ�6�'
RgE/\\PC񋄇6\v�{�eN"�Tʓ�?�)O1�����M����]xb�� B�av@ ��ŕ�P8%�'2�6m&�i>�I��q���S� @p�f5�T���K�����	3�Pm�[~?�ڱ�S}��[�#�d�b��-�,��`�1O.�D�<���IĆz#B-��N�:%��y�D��b�&�lZU'�c������y�ǔ���1��D	7�����J ?2�'I�Ĭ>�|B�E���M#�']
��s�R�F�>e�㣕�m���'�����6�i>q�	�9k& �`��a�����+t�J�IByғ|��w�|�kv��n�����Nd18��U&���p��O���O6�|"�Z6D��ؠ�TU�#����Ot�����G�1�t���G�J�$�(w��x� $�<{�v=j���� ����O?��6fH�ً���y\�a����Z�牱�M�&��u~��yӎ��Ӱe�p,�'e�Np����42���ҟ���� Ӣ�
����'��i��?-��"M�SD�K�D�2T��h��?3*�'�i>)��ڟ<��ٟ��	G�9c��*H6��A�F�]��P�'�\7�g4����O��D4�9O�)��L�e�=�"�Hqǀ�<����?�ش2r��T�O!�t�ϸ!.�
�A�:_�:ӎ�) ��R��By�l�3��� AC�8/�Ɵx�!dʓ2�r��M�v�"$�O(
�����?���?���|�)OFqm�)z�r��	!��s�=|�j
�NC D�J��?�M����>9��i�7��O�uʒ V��q��o��5@�iM4x7�v�l�CԦ\8E��$A.�i�	�?Mj �S���nϨ{���h�A]�n���H��d����ȟ���˟ �I���Jg�̊&\�c��NF��5JE)��?A��?��i1���^���۴��S��2��	�0"cnL�c��b�yB�i�,6-�O���eӐ������ך���b�	B�+��@b��)r".ͱ��'� Ȕ'��7��<���?q���?��M��A�}p��Q�:�.L�֪���?	������ l�ȟ��IޟH�OpA������,ѢJ�j��ON<�'In7����%���?�8�h&�,5�N$yn�`C��3�I��N�?hl�'}�֝����dy��wa~����Co��!J�@ ̀��'?b�'���O��	��M#`o�S�k �%a�AXa��j*�+-O|�oZJ�g��	�MK�/M�vK6��T��:}#�< �B�I����'.��Y��iK�$�O�-	 ��1���@�<!��8]jV�����;��=@pE����[���	ğ��	�d��ϟ�Oz`%
C��t�<�:�"V�l|J��q�8����O^��O����|�4��w�����:V�\E�6	]�OS&�z"�O�6m<���I�O��6Mb��jP�sG4�"�J�d��#���I?��X#�'N��'P�6M�<a���?q1�����PCP�����K��?1��?������F�J��O�|���|*�I�q���kH-��2dK�C��$��	���o�L�ɞW���Ԧz�\8Zӈ$���I�h�7�Ŋ(.��AB�ULy��~�͐��'�X��I�F7d]1`H�U����T�G�=�e��Ɵ �	���Ic�O�R �OOz$��jS*�3��I�:��Z�Wo�I=�M��wLz���
(a7z�:�E��@J��'T���g���U6�c����q�"x1�O��̉�l�AP���tL�&N9FE�&l
Ny�s�:˓�?��?!���?��?*�6�o�Ā���ܫMr�)Oܙn;�\e��̟<�	w�s��kT���W[�����K��� �������ĝ䦅iٴ���|r�'�?Y _�(��G�;�dܡ��D�+���Ӈ!Q��򤖺_u��k�Fy��X뛖T���r΂;`��t�M0�݉�E[����ܟ��	ϟ�|yb�k��5K���OBl�&i��/�6	�/�9'� 0t6O�Qn�f����I �M���i*��⠴IQ�$���0��,ɶ8�q�im��ݜ�`�����B��e���MA[N�� �s� m��0⡈S)~v�h��4Ox�D�O����O����O�?]�it,��M�	�E�WcT՟����l�ش�Ĉ�*O��l�E�I|��@ o��Y.f���XZ���%��[ٴ@���Om3E�i��)L|��Scg�L �0��7	;\Y��j�0L��i�ЛÂ�'���'@"�'J��'�@e���R�fR�y��#R��S��'�Q��j�4�d����?9������C$�r��#|6݉ jH�W����'���w��v�a�T�O�"^�������T�k��C$
9�U��1�@}h���oyb�w�}��'����y��Y�><4
TD�[D��	�'���'B�'�bc�<����<�'��Zj��Mz<��'�[�7AYʅ�;]^�ʓ;�6�'��'�r�䛶�ͣ��D9��/'N�`�,̯e+�6��O�p��`ӎ�H\L�xd��r,OHx�#�F��Y #�������K�צ	�'�'h��'�2�'	哵u}B��j�.T�P$	���3����4_\����?���:.��A٦��:pz��%o\�;M���7�ˑu$�q����M+�yJ~R�"�M�',h�ٕ�-`��9  ��$#*���'��FPޟ�H"V���4��d�O���ۓ¼�����&�A�h�8���O���O4˓Z��G�����'��$� Y��L�I9���C�]Vk��|Bͽ<����M�I>�7��p&�d��I�����u�x~bMS�B|2����H)R�剷�u�E�ݟ�"�'F�ԁ߳~��HsǗ (`�4�'^"�'4"�'Z�>�]�q�Q�w�5Y ���Ь��5�����M�U�
��$Q����	m�i�iA,�J�2D ��;�4q@�H��tnڐ�M���q��ܴ�y�'q����c��?u˔-W<lN%d�݃x�\q��Ԇ��	6�M�+O2���O6���O���O
�3r�U-��9���L�q��L��B�<��i&����'F2�'���y���;x��s'��g�9g�@�wz*˓�?��4�����'�?���$�"�s���SV(�N=�V4 ��.��Dѻj��;��H���B�vP�3cƠV�j-!��:��b׀���'�R�'k�O��	��M[1�
�?	�F�CX�(ŅVyH0����<ѣ�i�R�|��<����M+�SS܄+�`Ʃ~n�^ x���R	�9�M�'��,B�{������S���1�u'�w�r�8Aj\G��hs���0�
��'�r�'K"�'���'��e���#=<� �g�^�R/D���.�O����O�MoڤJA�-�'�7��O$�*܌�wJ��tOT��ˊU=��aH>	C�ijj6=�@1"��t���*2��D% H�q�k�o�d�{�`��]W*������$¦��'N�'��'̒�Ӑ`@4T���C�m���P"�'6�W�Hr�4K�m��?i����	݈)��黦D	f2kMPX��Ot)�'�p6�̦�'����?�	&�@��)��
� �L�;�NQ� ���R��#a�"��	=2�����q�\�����k�A�A�XiS��E?v�>q *��?a���?���?�|�.O��l��8x��������ѓc,���3?��iI�OLL�'�6m(	�q�4��Q�Lsf_(Z�n�|ʑm�ݦ�̓�?	���!�V���Y~2���rD�۲�M>R�0�d��6m�<����?����?Y���?�+� ѐ�K?/��p@1�fK����/�¦� %�s�L��� &?牍�M�;d��ͨ�IȌb��6k��@��i547�9�4�N���O��@�goӊ�	$��SP�Z�&�(2"�9a*��I������',���'�6��<�'�?�����4��%���B	V��?���?A���d�5j��2?�����:A�x\�8�e�%��Mj��k�>9%�iq6�)�d��6�2�H�U�6��(ՙ=;��O6�r�ƈ@�����,B_wD$�ɞ?rb޹h�t�ȴ@�ԆhcՅǨ2��'B�'`r�ȟ؀��D5x¡��\������ϟ��ݴ&e�5�'Ƥ7�7�i�u�P��^m	��M�eki��㶟�n�M[�GV\�s�4�y��'���t/��?i⠥��2��	��� /T����JRS[�I��M�*O�i�O����O:���O.b��V�G7]R'f�!i��C��<���i��A�'���'���y�K����M߮{6@}ځj��FJ0�M��fgt�F�O�I�����= ����e��#`p�A����8@*E�s��k�I�M%��$�'�0��'z47�<��2&L�\#�K7.xޜ�ũ��?��?��?�'��D�Ѧ���i���`)�&2��d����32�>f��1�4��'���'`�6�|����$	��P⑬�.6@��1`N'NuN�0/f��:�˔�I�4�~"ù���NYIe�	��S%.��yj���OF���Ob�d�O���5���vx(�E�^�~��,�bϛ�#�������I?�MӦ��}~�����Ob�YP�X(MT����B�S����UO'���ŦѪ۴�?Y�n��M[�'�b�"h�d	ԈX%M�4R�nWZX�!��Nԟh��^�<1޴��4�����O��䚂6��h��' l���kQj��kG��$�Ox�YT��J��y��'��X>u ��V2*��}���_�V�E@%?�q}��tӺ�l�p�i>���y�*�ce�� [ K0hW�:�0���o�^Q�E�*?�"���|���T�˓��[�"�9ʂ�I �qeb�*⧟?�?i��?���?�|r.Ot\l�
�;�MO~��A�s��bD�Aqy� lӨ���OdhnZ�5o`�cWl�,FD�O�"�~Y��4P���f6O|�	#\�J�(�"�վw"��$��� �-�cg�^ۜy�gA��hĴit栗'+��'�b�'�R�'h�'@�N�eT�ٵꋄp.x4q�48Yٹ���?������<7��y�
�����D@'v�Za����6�ԦXK<�'�"�' 8zy"ܴ�y�˞(*h$�Ө�r��t�6(ъ�yҢF(:�`e�� k��I�Ms-O����O��2�
�A�ЍA�(�+�K�OR���Od�d�<�d�i��0��'
b�'@BM��`5���.V���2��'!�'y�˓�?�޴r�'�Sǀ�p�^yhw"_+pY<屚'2镍wRܨ5��	W��.�u'gM���p�'��ez��:jn 9*�g�N8��z5�'[�'\r�'��>��2[���,��'�ܭQcȖ�I��	&�M�ܻ��d�ɦM�?ͻ<T�%�,E�4XN����Vg�&`�̛��k��oZ6:�\�lZs~�ݧ'�.q�S�D��G�8W�X�cꍸi�R`DU�jٴ���O���O���O���:�
��	�qNV8���
"�VʓLe�6��L>��'	���'ʄ0��Z)�!B�������<9���Mc��|J~Q��!��A��fR�H���` �
#�(��i��$�ph����~Th˓�vS�����@�8k����_K��Z�kZџ�����������Dy)p��IZ'�O�!	�ϭA�����J�t�U�F;O�n_��8��I�M+ŵi˒6�C�<�����b�ZX�4@V"IPry�akh���ΟJ�Kʸ:����Gby�
q���Q�`�R�V�5Þ�P���!0��I柤�Iȟ(�	۟��I^��XF��IX���`�ƒQ�m����?y�؛���7-���4�MI>�w�>W���S ��!y&�L�zV�'�R6M����� $čl�g~��
#�T� �8����!�Z"�t䪴��֟0�C_����4���Of���O����'0���b��.3h(A�EI�&����O<ʓ=כV
 ����'8�T>��Æ�&�)��Fؼ7֞L!V�:?��]�8�	ݦ�hJ>���?�gQ��xW�]((~�H�"�p��X��^�wKV��'f��]'2ReKyb�w����D�E��@+"��E4n��4�'���'�b�O����Mk�B�)CP6��ߊ$H>��'ϩr�Ҝ",Oj)m�_��"H�I�Ic#�\+*�T�Q� W�����8�M�T�iJkG�i��D�OBUq�"ɫ����<Q��$-	�
�5�<��RE���R����ݟ���ٟT�Iٟ<�O
F��&��N� yȀ��C!6I���cӜ|��9O���O���$Z��]�$�mޓu������UX�41A�FD=��J�"6�w��#$���r�l8����-x����$�|��+g�)K1��	K��hy�O�� H�6�-Q�9�"(��A��?���?Q)O��n���	ʟ(��#?QL���O& <I�F�q�)�?1^� �ݴ\��i;�D� �`���E1�X�:�Fį+�I1$6�q�6��_
�b>���'����<!X��A���f��!b�G�]�����П���H�Ip��y�E,B�Vb�#�H�v���D٧QW��rӐ�p���B�4�?IN>�;|�0H��E	�i��$JS�ۇP���kX�6�r�b�mڜ<ln��<���2ty`��.Hಌ�'M�0m1t�מ��	�BJ��䓙�4����O����O6��, �M�'�yuJ�sE�s��L����2���'�����'1rD�2n�7���z����`	�S����4f�f�7�4�6���:��A�.D�xqA�ƴ�X1t
 b`�����<a`��)3��� �����G��%K����N�A$�
Ae���O`�D�O��4�d˓UM�fŞ,2=2 �Z���ڭ5�&h)��	��yr�q�|�`�O�HlZ2�M��i��|�q� ..�H���χ�4��a,�/R��1O���^" a���^\$����;S]�L(`C抍SU@к3����?���?��?����O1���<*�����L�^�ej7�'��'��6픔T�b�8�֚|ҍ��"��X��Ӑ]Qܸ��OB�q��O"�m��MK�'OZAQ۴�y��'��*b��;q�8�&�c�\�!�6p~>��ɒ&�'x��ɟ���˟���3<�0����( _�؂� 6�����T�'26�(C`���Op��|��H���zh���ukr�kCm�l~�J�<���M��|�'��S���/��i�`Rtڵ:#�ɢ�.ycq'��S	<0q/OB���?���4�D�w�Zr̓1Id=@i��8z����O��D�O���	�<���i V��$A�a�x,��i�1��|�^&^K�ə�Mۏri�>��iB�3 ��+v
�!Ǐ�2/�d�� t�r	mZ#N��Qn��<��rBH]Ac�y�-O��x&��G��i� �U�>y��as4O���?��?���?������O�48���L:�MZ�&���m�h�@1�Iȟx��u�s�������JS�6� v�
�͂Q�������`ӄU$��S�?i���#yv�o�<�I�o�0����4��
�<�VNн2��dL�������OT���ET�xՁ^�<n�@'kގE-&���O��d�O�˓+8�6���B�'��l���'^��=K5�;�Of��'�6-Y¦͛O<�ਘ1gR���񎉄*�4JϤI̓�?��p��2􌙕��u3�iV>�� �1N����A4��`@2���Or���OJ��'ڧ�?I��I�	.��� �R�@���H��?!�iJr�2@Q��H�4���y'狇[3��Ek��t�)�nJ��y2j�� lګ�M�TИ�M��'T�.�(ά���ۀ �ၧm��]� ��ٳ�ᐵ�1�d�<a��?9��?����?Ѳ.�:�xi�BȴR�.��� ���Ħ��@ܟ���̟�$?��4'4P:��:[��A��	�+0�r�P�OT�n��MS5�x�O��D�O�>�J�i�
g�0�r����b�����9���P[�x��"�1i��BQ|��py®]bV0�DlұUN�)��ĝ ���'��'m�OM�I��M���J�?��L�1��Q"TeĢ;k��!҇A�<�i��O���'W�6�Lަ�Q޴<_fAS��f��5��[�5a�	�1HO��M��'2B%̧Z���S���?����4!9�leYU��9������Пt��֟��Y���6�x�mE�8����2F�1K۾�k��?��4]����q�I �MsK>�p�#L�%PrM9Z��"g!Ѱŉ'46M�Ŧu��(2pt�l�<!����1�@���H��b�����\���H$GT�$9����d�OV��Oh��GwB����11�B$�DǞ��L���O�ʓc@�栕;���'-2_>E@g%v����Fό4��(���O�p�'�*6-N��ipO<ͧ�
�А"���&�Gh�k�I���:1`Ơon��*O��C��?	p�"�D��|2�a�@lOd�<J�$4����O��D�O`��<�i����N�ʔ�qW� 
̼�q�'�<!M�I�M{��Π>с�i����Έ�V�B *��"$쬰�ha�Zm0p���l��<���tD(��&��	p+O�ӓ��t�v$�5��+���3O���?Q��?����?����iX�4�DjQ���IJ ��ei��?��Ml�,%h<�I��\�	r�s������37�͝C$���
�B�5���33��v�`Ӌ#��ɞ4u�7q�7nJ�-,p��"F�%��3�
w��b��'Nb�	my��'���
��8:]����7�]�Z������?���?I-O��m�/x%�������bTN�Y��r�N��)L7{���?iA_�$@�42�6#�=BR�@�h�*qRmB`�!n��OI`�~1آ��<i��jXp�D���?�Gd���������4����?���?���?э�	�O&0���^���Q�gS����Kg��O��o�v��d�'�6�8�iޙ�VD[w1���r?�J�n��Rߴ ����|Ӧ��եj�<��.<x�$���hc���"@��1&M� �Byq�O�䓡��O����O�$�O���T�,��ъ�c(�2��0d��uh�	*��G�!�'���$�'_�� �R�7]�Y���H�����<)���M{%�|J~����N��j^�BL�9�l!���p�ʗ:��гU� H��S���O,ʓ#�����j-i%�Ò:h��?����?9��|R,Od�nډa-64��5Nl���� ��@R�D�"��I��MC���>���i�B6���q��8��T:G6h� ��CpmZO~2D�#���ӿ<%�Og��>��� g�Ӷmo*�0���y��'("�'=��'���)�-����p���I� C�3��D�O��$Ԧ��BFvy�v�ΓO�<(�×1���B�*	�MR��:caJC�I��M��i���~���>O��ʃ:tE["��P��L0SQ�yQ䴩B�4�?!�i#���<����?����?�kSS�]��GԊr�\uZ@MT��?Y���D����(�#O�t�I��8�O��@g��$�!�B��]�v���Ov4�'�t7���*K<ͧ���J�4�n��&K>�x�����a�3Ǜ�Tk�ԁ+O>�I��?�Rg'���O0�r&E�&�[� ��5(��$�ON�d�O����<�c�i&�̈�M�2��]�%ON]=�<��"h���MÉ�O�>qҽiV�ܠ�E>N�e��I�&� �9g�m�t�lZ�^BL�oB~"�E4O�Y�S&��ɣa�J`8���~d��1�ȧqTX��Fy"�'�r�'6��'�r\>���eųzD�� I�70�|8�f��M�ń��?���?�I~�?=��w���&��Z�{ .�*��i`�zӚ�nZ-���|B���j�͊��MK�'��97ɖ!Gj�(piڪ=La�'���	rϟ��3�|BV�����ĉ��)aFЉb0�\.&
��*�ɟ �I��\��Zy����d��O��D�O����?ݺ��̈�m�v����;��2��X�����4!��'�����mx�X&��gmP���O� Z��R�.�*��:��^��?����O `!��'���ʓ]���1���Ol�d�O��d�O��}λ��p	�͍)�12�"�S�B)K��k�6
��F��I=�M����Ӽ��/K���afK�kwB����<�q�i��6mݦ���M�����?�F'� O�����e�u����;���p� �|~�-�K>�(O���O����O����O�YZq��y���5EEaX8���<�g�iR�E���'���'���R>�,A���9S%^(w3rP�P)�E�R�O�o=�Mc��x��4��/mdZE�QCZ�2���$+�'U��*��Փ?t剮l�PmK��'Q��$�|�'�t��e'G+\;�eLR-x�|X!��'b��'�����R��bݴSV���A����E/[N( j�\.k�\�"���'��'���ӛf�|��o��{Ϟ�y��^�T��lr ֟SD���HC�����?�qjƾH���������l��?pa�Ɲ?M 9��	BS��$�Ot�d�O����O���5�S�h� 3`��iz{�ƙ=��}�����ɿ�M�6!����ʦ�'�r�׈9X��"��	�is*�z#C� ��0כ�imӚ�)�t�7a��I '�z� 8��TC&��D(���^���aRcG>�?���&��<����?��?q���{��	�&�/2�%zȝ�?!����ėǦC����	ڟ8�O�m"��%'|���A��<���r�O���'װ7m����M<�'��7G\-OgJ����Z�'_0�)�șYs*����/C��u{(Oh�	߇�?���)�䓯K����,<N��D���(k����OF�D�O���i�<q�i+V�z��;��K
: j̘ӳ��>w	�I�M��K�>��i�p���Ö:m܄���D���-X�cg���nZ`�>�lZ�<��:%pҦ��ص�.OJ؆�O��i$S<#<T��0O�ʓ�?����?I���?A����<*��sF�ֻd�D��$p�j4o�=F�K�OB���O���$�Ȧ�]?1�����7C��[�FU�u���	۴����0�4�*���܈Io�,���hL�WA�#$�r�C@��(j=��I�xb�Zr�'��'���'��'���U
��H1�4� G������'�2�'�2Y���ٴYY�PΓ�?!��E�L!��ϳ<���y�Onx y���>���i� 7��o≉;{�٢D��$|�@�D7���蟬@�N�Cn�sè#?a�'Q�$�dP��?�@�&Q����\n9��0s��8�?Y���?���?���9�����R�0T20�qC��R!�\33M�OX�mZ�Ssl��'~�6�4�i��bC~��E1O�;�.Y�r�p��4,&���nӜԺ��~�l�Iğ<���m��B޹N�4m!�fE�o2
l)`�K $��&�x�'�2�'#b�'���'�V s�ҝ>W|��g�ڒ'��Q�]���4w��8͓�?q�����<iDgE�_Cn�	��E o>L �g�H�>v�I �M��i��O1�t�I��
�b^�����4�sDO
<_�1S���8h�pRL�r��Uy�ДR+��C�&�wmɁ�$u���'q��'��O�ɟ�Mk ���<1��")���q���'(��	A�I�<Yſi��O���'�ҳi� 7m�>"�=��T X��Sa��&*�&� ��o�\�I��@��xu��L-?a�'���ݱ_���#�ė�47~�07�S�<���?���?���?����؄v�-�3��>�`@�^��yR�'���v�@�J���L��4��Y'� �oZ�,�*���C��$��e�xb!g�B�n��?��������?�u�F����`�4;&h8*'e�2���p/�OM�K>1(O��O����OV��ۿ-���PC��$�f��G�O>�d�<d�iJB5��O��D�|�h،B�)Ď0�r)j�E@~RI�<���Ms4�|�'�.Ll}:w�
H��r1�_!Șm�FC�'l8,y��i�p~��O�rx�	�a/�'S��(�*�Z��U2�I�A����P�'���'�B���O���M��V7
܈��)TQ��qyC�����a+O�n�Z�W��I �M˳䚡G_8�bCt�a��7J�F�k� ݱ4 l�8�I֟$�b�����my�!�/>z���$����q+C!��y�Q����֟��	ԟ��	韼�O16�;���V.h0�q�
'M�i�t�|`Њ�O��$�Od��������W�����$_.��&��)iv�@X��M�ě|�'����j�Z�xٴ�y�b�(V�Uk c��^������y���(���I�'�IƟ�I�fN��i�薏.�N��a/Q�P��	֟��	˟��'i�7���R&^ʓ�?ѣD��f�j``���E��h0Ц��'��V���x��'�\صfV6�H�jT�B�V���Y�y2�'���0�ܱweddtU����q�@�ş��!�7Tk�!)´q� �#ҏR�?���?Y��?��)�O`�)F��2�U4!ݏ+��9���O�o�=d�$��'@�6�;�i޽���߷dþJ�C�z����"l�|B޴t���~����r�d�t��🬻��M6o*���M�b�9/ٶ�a2ؽ'x�l$�x�'�'�R�'��'*��"���.j�M��
*Z�.�#Q�ly�4Z�0����?q�����<i��ߚ�$���Ǽ�ܠ
����nN���MK�iC4O�i��(�	K0q,eb5M����`9f��V{f��Ґ)�%��$�{V���V���OZ˓)�%��՘-4֭#��P�bx�J���?!��?���|*/O^�o�`�\E���_`�Qf��ԁ`��,)y�I��M�n�<i���M#ӻika�k�t�",P��1\�P[����=��:OH���'��4���N�˓�j��_�����E�}o<1:d���bo�D��?��?���?Y����O�<�@a�P-Qʱc4m	r�4� ��'���'��6I���˓P�&�|��G�?i`�(B�S�}�ëܯa�zO�n�+�M�'0_bQy�4�y��'�~<�3���yAp,�F�D���p�'Xi�����A"�'���ȟ0�IΟ ��,��)��EĂ)�E gN��jy��ǟ$�'�J6�-^�8���O:�d�|B��Á��u�P��1N��0c"Tn~r�<)��MKa�|�'�j @K�	֩�v/ǵk�9��H$-��c�^
/�@L�,O���-�?�1�:��O�=���*���yANH!����O�$�O���<q2�i�[��I:������B4?-ȱ34�4Eo�I��M[��<��4�B��5"��L��&�A�x�A��i�B6͒�[m�6�$?�b��O�������^u�`�4&p�Q0�E�_`�d�<����?���?���?�)��9(���+H�L��6v-捋�̦}BvL�������L'?�ɀ�M�;'�Եт�HO��9���%{��r��i�6Me�)擝Aڜho��<� ��*5`�7M��c���t�4�8O�xk�HJ:�?���$�Ī<9��?Qª� 7p�ke�/��vO�?���?����d�˦�sr�ܟ�	֟ s���x;G�F#+Qqi��Kr���O��l���MKD�x�c�A V�X��Nu|L@RI��y�'_A`��7�	Q�W�d��4��Eϟ�6m�KJ]�ס�UQ���W���	����I۟�G���'Dq��ʬ��jǌ
�a�2�I��'��6͏t�˓y����4��Ha��؜MH)��gQe�&���O�6�R¦Y۴d�r���4�yB�'������?U`¢ޣ;�~aţP�0�t��dAP�vm�'��	۟��ȟ\�I ���LP���t�G�Axʨ�a��ה��'�z7M�$#j ���O^��5�9Op	{b�W�|��̹v%�=�l5$	pyr�''�&�9��O��t�O�l�qSf]=ta��"���$�	��r�ֱcR���V#��U.R�X�y�hF�_�daS4�'���т�H>9���'=r�'F�O�剩�M����?Q��ۘ�:,���S��h�U�<9ָi��On<�'7��ܦ9kߴO��]2�eI%E����R�X|�0I�M]��M��'f�&�J����J���?u�]J�P���j��`;�-C�)��}���	ʟ��	����՟��I_��ܚ�{�n�{�d�1��	TU�}p)O��d�զ��U�#: �i��'�Фs��
���s���!̰���i-����1���|�r���M��O"���D�*C��a�K�Rd��֩_y|�R��Ox��?a��?���DR�}�-L,4�t���*�xlř���?�)ORm�_�����̟��	D���Xb,д1FIDT�Խ"AL�����H}B"v�>o���S����3����g
VZu�`�BOFJ�2��зMZ`���T���A���C�oD�`	$��F��	��N2Q;"!�	ğ0�	۟�)�SHy2.|Ӵ�U⋉���P�M��)��G΂s$��d�O�	m�|�@����M��eǅ�l���'r\���@[�fu�6-���o���ퟠ@A�%#�ĮXxy���H�����}�
Bt����y�\���I��X�	埸�����OÒA�k�:E�V���Cj��9"�~�T�b���O���O��?i������,��E`�u���mт�)0Mϛ�fl�T�$��S�?����E(pn�<Ir�ׅq tCF.]-�f	���<!7 7j���D�0�����O ��u��1�J�;S:��	�+F�V���OX���O��[B�ƫ ���Iß� '� ��y���ƹvŎ ��Z��x��	��M�c�i��OH����$��0�QBZ%ei6���8O@���$����!��������O~$+�o Q�BaD�jH]ef�*!�Xr��?���?a���h�*�d�%���{�K Zn�@ #�~���i'�My2�oӊ��]8X/8�Dc&R"�d��	����8�M{r�i�7m�u��6{����=A������O68��I�*f60��cг� AH�&@Q�IsyB�'���'�B�'�N�-A*��6Cɝ3��s�L�j�� �MC�.ֳ�?q���?�I~Γt���� T<hNP�/$%�4���\����4>�&�=�4���i����S�eP�B"�	i�<���V�]^�>��d��<Qv#�y`�������Ł\�f���FR�}��`��ZS��$�O@�$�OL�4���|�f�9).���*���p�*ަX�
�j�Q/�y"m�^�R�O\l��M�Ŷim�̚B:QyTY��
N 5�1e�|��f>Ob�d�27�x��'{�pʓ�r��Sxx�@`ƾrV����E9%���̓�?i��?��?����OL�9&	H�-&]�U��f(,�S�T� ����M��B��/r�h��<��JN(+��IU�E7}�`�GV=)��'��6��ަ��?���lZ�<a�/�����e�!N���xND&Ѣ�!_8�$ލ�䓚���O����O���@�y2�EX�MM3H>��H����:wd���O����&%	����'y�S>�ka�ٱ1�=3��L��O'?�!V����4i)�6,�4�f��=xW���X�M�/C�^$ʳ"=lU`<ʡ-ѴN��ʓ�����O��H>���W��E ��\+q�,�[�͊��?����?���?�|J-O��mZl*Ip�@Q:o�u���֫kP c�Dy�b�R�� �$�E}Rnl���1��d|��ԇ3d�֡jV���MK�4	����ڴ�yb�'�R�0��?Y��Z�䛒�K'35����,A<���p
p�x�'��'�r�'���'��z��:1�'i��Rq����hQ޴U� 8����?������<a���yG�̲E@�B�>'tfa��%�9~D�6���i�L<�'�J�'tq���4�y".�n���h��^%��|��)�y�.^��i�I�<~�'��ߟ�	J����R�k�(�zQ��#{u�Iǟ�����8�',�6�J���O��䎽" �S�_��Z����5_i��"��u}�xӸ�mZ���(�E��/ϡ$XL��P�N'b�ܕ̓�?��Ł�`�J42�^�����R�waB����$1R�̖($V�z��O�^���D�OR�d�O���'ڧ�?���3(r��@(�A؎0�녶�?�b�i9x�X X�޴���y�(4y��p�aj�~ڒI��d ��y��o� n"�M;��5�M��'&bM��No���3yU<�#/�Vʴ<C$)�8K^8�W�|Y�P�	��,���L�������J@�Q���P+"h���pyRBiӒ����O��D�O:���$��n� I��VT�h�PhI��!�'��6�Ǧ=�J<�'���'12z\� ��G����I&��Y����bʘ���6:41��.�O�
L>�/O�=@aL�4E�VDD�ְBdV8���OJ�D�OB�D�O�<�Կi�F<���'"T�
��ȋB<a��*]=4��ۙ'1�6�&�I���$E���Y�4�?����5�����P #��i�2	ʍTU�T�ܴ���$N6m��'��O�>�،#@�I�g��;v�=�!�
� �H��ԟ��I���Iڟ�	M��
\�����{P��$ڒE�t	����?���Ư6�a��M;M>�����4��&�a��@6���y�Z��(�4tW��Oe�A��i�ɵ�j�b_�*����"�^�(g�,#"`�\�Ily�O-"�'�b����qh�m�@�r<�#��CO��'�剂�M�2���?1��?�)���#&�A�k��K'N�fi~�ps��0�O��lZ��M;`�xʟ�hfhܭH� 81������e%O�j����3N��]|��|j7��O�u�K>��d 5\��D�����Y:����?��?	���?�|�+O��m���:P�.��4��k�4K��+�iycr�����O�l�k�0�:�G�8�d �5/�/$�|���4q囦��.�V3Ol�$U9M<~���'{q��{��u�@�+z�IwJ��.En-����O��d�O����O���|r$b�R��
�뀱iVT��tЁ_�V��9U���rS��y�S �<	�� S�����J{�27��Ǧ��K<�'����-$����4�yb�Hn�����܁T����2��y2��Jx���.)��'~�I�4�I�yva�׎��*�I���rK�M���d�Iޟ�'�7-X"�����O��D	)IL���m[*6|�y���-R]�⟴��O�m�>�M{r�x2�L�nO*�#Q%�e^$!�+�9��$J2Mˤ5 ѠBqlҒ��98��slD�D@�n�;�O9?[�!ʕ��. �0�$�O����OX��*�'�?A!O|*$0�0��R���?A�iV� h!V�`�ߴ���y�"��oLd=�gQ7�F8Q4���~2�'���*d��i�ҍp�6�V!�)�@ �}��K�;[�����
%g�P� '���'���'���'/�'ŘM!Ž1|l��Ǝ1�P�BY�� �4�L�	��?���j+��<]䚙`�f V��ф� O��'�7m�˦�SM<�'�J�'y��K1nԳS\P����y�I��O�B�L-j/O��"���?��4���<0G��/�@T�Ձ��1�����?����?��?ͧ��d��q�(��t���5ڽ�*�#cE�m�C�h��K�4�?yL>9�R�<޴m��%~��!�V�ۖ�D��ЁÏz&��t�i��6�w�H��t�h[@�O:���']���wS��9E�'L낌�@�
J�t�'���'"��'ER�'���:FB�1���d�F��$�3e��O����On�O��'��6��Oʓd�z=���P�n�����5\��xh�x��q�n�o�?��6��㦝��?y�K��@�so�E�>Pz�a����0�g�OԙYN>-O����On�D�OЬ;��ƿMt�6Қ!
"�� ��O�d�<E�i?��e�'o��'��S�(�y�t��c�����D_rd�p��I��M�#�i�,O���R	�?;�܉����f�YP�jȠ�d�*�-��2z˓���+�O�T�O>14�ֹ1^�����3�L���K֤�?���?����?�|j*On5nڶ2X�P���.
=�=D��٨�j�@^@y2Cp�|�d4�d`}2�a�̤� `Qc!2C��!b��{�l������4a:H�*�4�yb�'�,Tj��?usTZ����F�'b�a��U�41@���
t� �'<r�'2�'D��'��S�(z��q�5*��C��!����4)U�x`���?Y����<���yl�_�8GA�:;�8�W���7��A�I<�|Z��@.�M�'����@�/ >�y�A�m��2�'�P!��C؟4�֘|�U�0��쟸#���7,?t5��@V�X�x���@ퟸ��՟���Wy��l�,��2��O��$�O�42����B�CĀ[�F�0�.������զ��4�'����s��
R�Ju{v홮<m��1�'����*gl:m*�mXq��	�?-�t�'h�E�	;Aҥdm�0X%��H��:� ������ܟ`��J�OwaR�'6��Ԡ��l�	p��#;2�d�ʕJ���<	�i:�O�Nդkl��I�J&�p��e� vq�ݦ�ܴ@2��CB$��2O��D��d�x��B�БuUIs�č�(^�Zϟ���OV˓�?����?����?��l��0�mJ�)W��{ŋ�� ��/OĤmڧ	�U�I��<�	V�s��q�Hͮ3�|!�3%	10�P�S"��'��Mܦ�۴uH���T�O����C�5�1���M�����B�lEY�^%J��2,
���'�(u'��'�l=s�lH>�����O����'�"�'����^�8	�4/P����x�����'Z*lCf��w�!���}�����_}��z�F!lZ��M�Md�f��pF�IQn@S������۴�y2�'SJ��4���?���U�T��ߥ��T�&��a��E�;鲐��r���I؟���4��⟘�Zk�3R�Ҽ�'�� �E̚��?���?!�iHXڳ\� ݴ��s,D��
�O
�8��Y���L�|��'���O͂�J��iJ�I8Ubi# "�'E䌱�`,x
� ]�,��X{�I~y��'*�'�ҡ�SՎ��v���wS �£N	�?9r�'g��6�M�ӧΩ�?���?y/�6�h@�{��y6mvK�������*�O��n��M#E�xʟ� Ne:��˱)��]Ȳ� P��JV,T&8/��@U�� ���|Z���O�|�H>�k��3��w(Ld��#�,)�,���O���OL��<��i�fQ��9A����q��0cS�K���*��ɲ�Mˊ��>a�iQ�t��b�8`��-!�*F�+�"���n�Pm��3h�El�D~�"`��1��+��%k�0�1$�Ҏ�t��,H+ ��Zy�'��'Y"�'��R>�{�'�&p��s��,
蒰���?�&�hyb�'��O}�b����F�@�E�dx@�0�Z���Qm�M��x����Ǉ@i��<O����2@F�8�]�2�ꈳP5O>-��ǋ�?�s�&���<����?!@���Z]Z N_%xb�:�Y��?a��?�������p���ޟ��Iğ����Q�|#���J7
"	�#�Q[�yu�I�Mc�i�BO�H���˼B�T���}B������8�4

�w5�Iӂ�C��u9B��ӟ�#Wc[Yx� K ͅ�k��a��F��L������ݟ�G��wk�����[-?�� Ӑ ��6G\�p�'�7�#G���O6io�F�ӼkS��#�������@M,dY4JF�<��i��7-�Ӧe:����-�'��8�R��?�x�m�VZ�֬� ��ԁc�U-T��'��I矜�	�����㟰�ɹ0ˮ1������љ��<&\���'�N6�ɇkG����O��0�9O��� �A+[Y�$��Á/DxՊ��Uk}�Na�\�n-���|j���R"��$/q�-����.d�X�a
wehP�����Y)����wO��O���H`�СEDQ�x� jUo7XlP���?����?1��|Z)O(pn��mj4���.N
�����P-���_2*��7�M���>!ƹiIB6m��5Z7�/L��K!0%�͑6Q�кi��D�O�92�fһ��a*�<9��ǿs����f�L�T���/8t���?����?���?y���O�F=�<$��TC?B?��3t�'!��'L6�^&X�h�j��F�|���fN�!0�1j5�9�b�K�2�O��oZ��M��d6eh�4�yb�'=��bȂ���Qs�j�7_-���2G�,�$H�I3��'����p��˟��	^c�c��8����m�)]4vd�Iܟ��'�7-\�'���O���|�4�����Er%e
�J�}0��WG~��>1��iu�6u�)"�)M/`���3�Ɛ2Nn^u�엩1�z��Ƃ�j9����ǟrԙ|�dX!q�h��N�9V>��ǭ��r�'3b�'����Q����4E*Z)�'+�&AD&�c�+�;n��al�"����y�?�[��*޴1��!YS �s�'��!Ό��is$6���&6�/?�#!\�	����DȊm�8*�\
&�,k����d�<i���?���?���?�.����Rf���-S�4��N��:�E��L��ş(�RG��y7�����x��S/Wh�ي� �*�Dj�Hu&���t:E�z���	c|���(z�F�s��E�&�.�;l� A�'�'�\`'�H�'���'��D1u/�*@��������I��'�B�'�_�:�4R��TZ��?)��q(�(��"b�H�"U�PwXi!���<i���MSВx�Ǹ_��t�CF6�ʅLT����^̓φ(|��f��������'	�qv*��`8:���A����OF�D�O���/ڧ�?����e<hi)��T�u�q8�ˁ�?�'�iMD���^�,��4���yJ��%5Z%z�� c #;�yRG|���n �M��E�M{�O��րE5������P�5��!>᪜ �o��G�|rU���	ȟP��ğ��I��L�QG����0#�ćIq�E��Cy� k�n���N�O�D�Oz���$���څ��L�z�t0 �� +�B��'F�7M¦�L<�|��	� d�=@�o�>��7kG/ T�G�����ެx�0��wKҒO��5�l��Q 2}*AX%l�-������?����?	��|.O�oZ�@,^)�I�Y��xH��/g�4�!7�Q(5�X牸�Mˍ"!�>��i��6m�O��"g�p�N��R.\qJ�胉�g66�>?i�#V&4#��)9�Ӗ�5@Z9 ���`�	Cx��N��y"�'���'���'���	�!�b�����?V�$L`q�t���O�$D˦��b�ryB��F�O��
Ѩ\�pn�Y ���0�`D��{��'T�6����Z��Dl^~MU;F_�Y��o�8�I!��mMt���������|�V��S៤��ʟ�0F��&ٰ�����1&z�	ş`�	Eyc|ӈ��I�O,�d�O�'%If-*���:K���%�-"�i�'f&�2���i��$��'bu��¤� ��q���O-FxJ}Vg.XW� 9�����4�.Q��vt�OD@�d"�n�~��O�o�r�KG��O��$�OR���O1�˓	���i��lt
�h��غy+\h��&�E� �fW�\cٴ��''\�Qg�vML`��KSL�!<���1�O/?w�6�֦��$�����'b� Bc.��?��1Z�d@5'�0��q@j�0|$��zQ�o���'���'?R�'�r�'��;]�p͚$�*��xц��-��t#ܴ�
�H���?������<9���yW�B�<���7�#QQ ���mu$6-M����H<�|2��Ҏ�M��'h�)���'9�J��ǥGP}��'�j�����ٟ$qt�|�]�X��˟	���.1�B�(���R��nٟ�������tyaӜ ��O�O���O��%�\�k�>��� I�@�*�P�h.�I������k�4&���� 6�2�ٵlԸ�p @3	[�����h�	���P�q��V�ӏ�⏌Ɵ��V(Y�q8T���� -�t�	"������	ҟl��ԟ�D���'혅�$�,~���)f%A(�%�OBxo�2)�Q�'�7m$�iޕcEۊ=<b�Y���96���ȧ������Y��4s�ʡq�4������ �'-��X7��\�>�C�M9xu��Q%C(��<��?���?)��?񥡚�	��uAkҽ�%� �P
��$�㦭���Dy��'�x�ӂ
^���)GN߹&.Ѕ*��W}bAm�t�o���Şv�
I��"��Ү9���J�9����+�_/0�Z*O^���_��?	 J!��<�,��ZH$fu�j �7���?)���?����?�'����=ۓ-ȟD��ˋK��Y��݊c`�Bob���4��'6,�5Û��hӪamZ�NF(�c�n?� ��qP
���m�Ϧ!�'ĝ `ɓ�?b@���w� ���.h���'�Y�w��eȟ'�r�'�b�'���'��fmX�g��9�xA��Y'q�8�I�.�O���O�n� ��͖'L$7�?�$�&����TKK�&	���3��j�%����4^x��Ox���E�iM�ɭ;;1�'HғE��%���,~�)�	ъz�"�B��Ky��'���'7b�ȫy���c��*s�B	�͌D�'Y�	8�M�4�<�?���?�.���C���'�8$��́�}�X�[đ��[�OؼoZ��M�%�xʟ���nE�51��(͇��@g@ϬJ��l���3U�R��|z�%�Of-CK>a�lΖS6\����z$�0���?����?����?�|
/Oz�o�33I�13�+FP#VN�S�rs��sy��xӘ�`#�O5l�-ot����œ�1�l�+��@����޴3s��AJ>4�F������S50����{y�Q�ɀ�r�j���yA�,Ұ�y�\�\�I៌����`�	���OZ���CnB�|�3^��U��͂�5��pM�I�|�IW�s������cvl��o��I�A� �l��:věրm�x$�b>�i�C���Γ~���#�?v�>�	 ��`�ϓZ:*�#���OI>	.O��O �PA�֔�v�h�!E3.&���tL�O��$�O���<Qֶi}؄ј'\��'J&I��A�q5P�#g�В����r}�w�*lZ��}�D��7mK;z�Q���(P \�'�`��l�qr@���dNܟ4���'��NO�i��#�
r�`�'�B�'�B�'��>��?���Qq�ͳ�nZ�:�(�	�M��G�b~2�oӖ��ݨr�и�'���&�AW�&��牳�M�V�i�6-�>9��6�%?���@.$Lr��A`� �6��$R�!����-
PL>�.O���O ���O@�d�O����	b ��%�̲8���2��<	�i�,u��'A��'���y�IN�[9��R�f�wy��+�dl��di���|�
�'�b>�z�	X`et4 �]�D �aD�F\����/?�"R<=������䓿�D�� R*�H悆Bj��Д�[R�t��O���O��4��˓V�v���y�EC�r��yђK�;'�b��n�8�y@x�z���O��lZ��M���i�v`�ͷY�� �/N�^�ꍺ"'�9�v���w�J1P������h�I�0 �\���8%��)�&3O����Od���O����O��dI�ZV�9�<��A���.UfDE���#:ҥ�K�Of���O�mZ��tA�'R&6�-�D!%o�a���$.�NxZb钄@��&���4z���O��◺i����O���&[:0�a�	�&E��l��
'~ ��+��d�V�O���?!���?��8<�,��(ɟNN�Q,�$Qs���?�`:L0B�,�
w�(�,O�����瓰j�2A[�CP
�b�T�S$*Y~�t�I��MB�i�RO����@��.�<2YP���Rd9p�kge&�@9�d5Y��˓��դ�Onq�L>!S`�C���B+�#[?��x���S<���i����@ο:��u�vF�%	���+�$����&�Mˍ�F�>i �i�^А	�>?k
�ض��	e�0��eӒ�l�.�x�n��<I��O:���c��D�x)ODi��M������T!ztv5ʠ>O\ʓ��=�,���$�k#LK14:ZI9��K�$���ɀ�qo��ʟ������y�⌓jt�H��*gV�9���ZL�6�ѦM�N<�'�b��E�d��4�yb�Y�8��$rVLR����kRFǸ�y�/�g�"y�	�&.�'���Ky�̌q�,D`ê�#� 4WǕ5�0<���i,l�� [��	�a�:���d�(+b��&��?QFQ����4yQ�fl(�$_�NV�EIu��4^����	;m�$�O�)��e�'D�.���d�<���9��D��?�a@R�6�f=4�\^��d:��Wg�<)� �1)�>ɪ� P\�n�{�-���?1ÿi���b�[��{ش���y���{0��P`O�%P��y�D��yR"c���m��M�4�[�P#;OJ�Ċ6~�^����7���8�%��s/aK5���*�|��!�D�<I����*�,�:�*��(I )6%��	=�M[)G���D�O��?)k!�:���+���'�N�#������O�6m�I�韴����x"� z�%@۰d�@5I$��y8���c�<!�d��6q����䓵��>�H�92�z�AB��a|r�w� �H���O(u�� �Q�`}�Gl�0Zk����;O�IlZm����4�MCտi�>6� B���h2̊b�Xa����
N� ��7�k���		X�Z�"��O�2L�' �t�wrl:��l���cgɏ�&��(�'A�2��/�-+01t*P��Vɇ@�����x�ش2�^ �O�6m#�d� �]�S�*i�Mi.��Ro¹'�Hm���M���q&l��4�y�'��m����"m�����%J�gH �b��:p�5�I/�'v�IE�.�1��NW�]�$S7*C�$}Exr�rӸ�X׬�<1�����T ��M �HY�"��!X"
��ra�������O 6M\D����i�<�V��%�
A<q@�)�6Jx�c5��	7�Q��<���o$���D���U�N����ܸ~�DdsA�r�x���M�˱�p�3�L�g/��Zp:
�C Q�L��4��'#����Vl�/~H��(?v2��J0�:�6M	���
5N���5�'N���I��?�J�Q����F-�~ݐ��Z��srk�̖'=�{��_��ѥ�O��'Ţy��7�G;�p��?���$Be��>@Tc7n�.*DD�b$^	V�@�m(�MK��x���f֑ �6;O�ܒ��K,[��@0��h�4O���K��?)Ӡ7��<����?aB�A�}�z�{�.G-O���C���?����?�����礪���ty��'�(њ��

���� �Q�p����f�Mw}�/j�fo��ē6?Ԍ)_��pq��N�����;?���M�1Dl�(B�X&��"A�mZ�Ll���H�D��7BM�)��DZ,SJ���'0��'���S�$��֕��@	C!^v���П���4<p`�'��6�,�i�)�����RxBu�}�����l�Hj�4/��v�d���a'}�t� 'R���|ם ?M��3�@�5L�����&]j C|�R���͟���Ο��I֟r�ɄS�ܔ��E�u9Ī�hyBai��]��8OJ�D�ON�����Cԍa@�Z.]�����
M9Aθ�'�v7MP���!O<�|*�,;�r�"�Y�"gVA�&y6`���i~B�L�n��IRB�'��	�*�� ����x" ���ϟ#�`t�I���I��\�i>y�'��6m�~1󄌌&�2�B�l
��`8� 'W�H=��U�?�`[�4��尿��4ev"Ń��G4i��2���<�U���M��OxR��ܝ������wt�x�$Nٔo'zd�#�3��1��'�B�'�']�'�(�Lڄb
Ak���m/|�y�1O����OTm���>�:қV�|2d�a�@�ځe�Z6"�� BI�Ht�O$�$i�󩎪7|7>?!��0:c��{�� ,3`$Bk_>d�l��"��O�	�J>�*O���O����O����\h�� ��L�;7��x�n�O��D�<ц�i0@�'W2�'��S�?�RoB!u�:=����$
l�:�����M׷iȄO�SG�h���1�H����1r�Y`0!�j߮�<?�'xԮ�����J�0J@���NF�:"�G"����?����?��S�'��ݦ��$�~�t!�D������Ǐ)fc��A�&�D�A}b�y�Dp�wbFj��)��I*e�ftʢGT�� �4��2�4���@��i�����SԐ�f�9,x���c�6��Yy��'��'A��'
�P>�Cc�CǮL���Z"��ܘ�@�1�M��&��?����?�O~���c��w��:'��/}ء V�T�v�����z�D�nZ���Ş.o���ڴ�y��ƴN�pAH�+U�R���6B���y�	T�Z���mb�'���؟��	�rUĜR���"-�V���}\v�����,��럐�'�(6m¶^�Z�$�O���R>M؜���(T|~��P�ԥ�:�X��OܼmZ��M�A�x"�="d#j��i��d �hU?����:u�P�d��*rΤ��h	���~�&�-5����R"&5"F�J"*"���O��$�O��D3ڧ�?qc�>-`H|z�o	�[���;0m�
�?	�i7 4�A[�x�ܴ���y�n	4}�Ҽ#�+��X�\2�d@��yҥm�xtl�M�����M��O� yt�ʁ�J��֣0c��X��B�tX|�� :n��O\ʓ�?q��?a��?��I4i!3,E�^R���C��[@�-O�lڦh4&x�	�	n�s��s��>3֐j���?j6��v	����X���47Љ��OCF�"g�8,���;e��!g�DPs N�w�&���_����`:12�Co�IFybh�ZA\�ۥ	D=%p*h������'�B�''�O�I��M{�<�A`Ժʌ�Z�N�C�82�i��<a��iI�Ox(�'��6͈��(�4-���81M �	�%��ܤm�DZ�, �M��Ol����/�j����w�-���3��C+���a��<	��?Y���?i��?���� T	\:b�M�KW�	��X��y��'�"Fz�Bl�!�����4��1HZ4�$&3\3��s�#_�� I��x� g�<�oz>%���զ��'e��a���'�l�,� df�%���eRX�	�`��'T�)�s�H��J�(�xq򰢁2?���� �!�j%�&�X+W�񟀗OP�������T�br Y o����L}Kx� po���S���^�"$2`H �[��d
DgS�&=�=8am߄i���[��3|�b^|�䈸�������P��8B�ɕ�M��f��3� �*Cj�|�0Y���U7_�f)+O`o�v�z���'�M� ����	F���]�pb��U�Ϧu�ݴu����4��$�DF(�+�'rbDʓOb�0�I�0�0T�v,ڑ�z�Γ���OV���O���O���|�Q�=f�^h�ɍ����7�B�:��D�O���&�9O>�nz��3��?B��RqטrH4������?	�4�yb^����PXŁ���	�_y6ċ�k��^4p}����d���I�hq����'1*,$�������'Q�ES�%�`�R��$�:60����'L�'U�V��9�4������?)��8�Q�G�>&�P��1Hi=�%/�I����O`7�s�8�'�����k���r@G�*�q�O�ӵ��3��TТ�Ɏ2�?���On8����|���E%�M��� �O����O����Oޢ}��j��I��f��T	f�M�z~l���GP�6E *��		�MK��w)�ht,����8R
������'�J6��Ԧ����t� hoZr~�
�� ��ӃF��1 ��3{����8z��+��|T���P�I՟P�	����g.	�EID��7����U��ny�{� �'�Ot��O�����F
h���"G�E� ��ȉ�<Ҏ��'�7���!��H����P�?��U�5�6���Ǉ�%u��仢��
ǣ�-v��-d@ԣ�N����[�GQ"t×(څO|A+�V-趥�����[�"�$Q�a!�Ӆ`Gr�Y�JۥCG*!�Q/>���5���C�l�4%�9(�r-�2��h�cj���T�T&f�B�ѓ+K 2�.��m��I�@qRf/8��0P��h�Ը;$� k�z���Iң֢��e��Ԑ[�U�|�m*!��7$AnA� �c<��jtL߹,�r��Qc��'h$p���X�H�ܑ1F̔�2&΁�ƈ�,�R���`u�d9�#c�c�@�ҡ��/^��D�خD赎�6"����q�6�G�\"E�(v����5��^}��'v�|��'w�J^�$��!Q�Z1��S�h@L��%ài�6M�O��d�O6��O��`kC�O�������c� ./�̩�3� �0L5�'	k����>�d�O��H�RV���x ��]�Ȼɉ����%��MK���?9���?y��	$�?���?�����ͷDrr�!vl�#0�R疭6�'G��'���8f����������c��)G��8W��Сp�Z�X��f�'�c��:*��'��I�?������0��y����eR��4�67��O��D�[i���f��I͖+8@�f�<|�����8z����N�cr�'�	�?���џh�'p�Y�b6�u����e�,Tk�{�ˆ�B�n��y����O�=��T	�Ԙ���A�r2��J!�˦e��[y�_�)���Zy��'��D�U����SHD�}:�5ae�ͼb�*��<y��?��'�?���?QE,�Oꂝ���@+�ԋ�2;���'?$a�R��q����'�ē�?�I��+k�@�f-E:t1�'��.�^�H�O����O2��<ɦ"�\�H��B��FpR�*c��$ ؉�cX� �'�2�|B�'���ݪ,Y@ Vh��֠0ǁ�&�|��':��'��	~���K�O .U·�4jT��Hrb��b�x��4���O��O����Oz�9#����p��+$U4�ЄR�2�j�B�>)���?����^J]�O$�	�-BY1`K�>���� c�ws�6��O�O����O���>�I�@��ȡ՟$�
1-�@� 7��Oz�d�<)��ZT�����H�I�?��v�l���J�/�ưH׋߱�ē�?i���N���Bܟ�8�G��0���U� �2��i���
t
�L�޴�?���?��m��i���w�C(Ɉ�+G2h���J�z�,�D�ORd�,5�	nܧ X�@�$�9#`�hƠC0Tۮ oZfd\Zٴ�?���?���/(�	Gy6GJZ`��?VQtu�Ҧ+�T7M�e��$>�$)���h���e��lTB£cR8A��ʝ�M����?q�<��]��[�h�'���O�R�ς�m$��qC��saf�`��i��'K(b@L/���O����OV���Rg���b��B76�4u�$�TצE�ɸ�|q�OF��?�O>��+�R�cm(=���l�&Z���':`����'��IƟ0�	� �'�H���9 ����0��,x��Jq�ī�x�����Ob�O����O�p)UFͮR^e[F�"C�%��΃=_ВO��d�O��$�<�'�N�I�bڭ`�(ÖYtA�E�x��\���Ig�Iӟ��I1����4LX{����� �C���r��O����O0��<Aɏv��\{sdX�m��ܸ��Ǣ8m�Y��-ǂ�MC����?I�}A�Xq�{r [��"|�ũ����"�� �M���?y+O��R���K����s���M�xjq��a޲E��qÊ=��<���L��?1I~z�O�z��bE��*��D�p�L��޴���6;*�oڐ��i�O��x~��5��}pS��.%�v�����M�)O��`Ť�Oܠ&>�&?7�[1. ��8Ō�%y@�x[i�<nZ76zx޴�?q���?���v̉���@�}\� A!OZM��q)G�t 7�ҷd`��$�O,˓���<	��$S�1H���N��J$ȒD@2����i`��'���q�PO�	�O~�ɕ���Di���H��։cF���4�?I*O��p�J�}��'5�'!`�����#ϩX��x��^�v��7��OJ\P�L\�i>��IY�i݉ rG�h�r���Eʎ5���9�#�>3@��?M>i���$�O�i����2�i�e5�t�dj�-1�ʓ�?����'^��'e:5��N6Hdx0���Y;V�i4�GHf�x�y��'H�IʟLHƃ�X� �8�&Υ*5������hйi=r�'�O����O���CF�;ϛ�
�5	�N���������?.O.�D�^�r�'�?	X�ډjɂ$�����)R���nk��?i�d�:T���q�I�w��ժW�	�Vy�h��ұ��6�O*��?�E���i�OZ�D��klC�=K&8�%��wcN��aJ:7�'�R[���.6�Ӻ3'`�p1���� wx)�L}��'�I���'��'���O��i��Aw/���uy�7�0d~���D�<� Jz���'L ��a�Yj�|� c�	HL$�mڹ���	�	�<�S}yʟ��iqD[ 0�Ƭ�CΗ�H����\}J��O1�h�dP (�:	zr��=�T��b	��l�꟔��ӟLQ�dٛ���|���~�F��2��A�`M�>=�6�j���.�M[����$�S6(���y��'Y��'�ʄ��+0 IX#/�:+�4pf�vӰ���?j4h$��ڟd$��݈Z`|��	�x�lq��F�x�F����$�O����O��e�()wJ�X��	�O��&� �ےk����'L��'�'M�	)*��5s�@�	b-��P�B�XJ��d�Z��0�'"�'��P�0�������d�ƕCa.�#��,;� ���
�byr�'���|b_��2����9�%���lyF	<7ص*T�����$�OV�d�O>ʓ�,�Ж�A�5�Ι�$H�Ex���P�L�u�$6m�O�O ˓RV�в���(h�d*P���#@n��sǉ`$6��O��$�<���L@I�Ou"��5F-����0{g�۹d�&�QHR����O�˓}`��B����'���욿g���mݕ/:b�AGU�����O��HC�O.���O���⟶�Ӻ3u$�Y��&�=J�P\�)G���'Y��-u��y��Gӊ	�u�4�W?v^��;PL��Mg[!�?���?����
/O���	O�D�"�%bk�E(p�S3ga,|�ݴZyܝA���N�S�OW_��xJ���$uԅ��I�:|T7��Ob���O�����<�O��p�&!B4��+܈����f#(`���Hg'֝&>�	؟���$DLڸ�ЍC�N���#�#:���ܴ�?y���	dщ����'��QZA�O i����p�0Y��$�eL�j}b�]#QRT�������	Qyb��!z2$PE�V��B�ÀS�nY"I#�$�O��$2��<���9� 03�FΗHF`��B]�B��?Y)O����O�D�<i��+��	A�AF��C�H0 ��@�J֩*��I� ��J�	by"�hy��H`�Z�I#���)�����N8듅?����?q(O�ѹ#e��d�'�Z( �Ŗ�g�"�����cV�hV�e�p�Ĺ<���?���~�d\ϓ�?1�'���c�l��Lg�*:�XU�ߴ�?����֔i�^U�OZ��'�t�R�a� ��I4���Ef�����?y���yҊ�m��^��'"N�T�C��q�ܸ4
Ncu��l�_y��3Q�d6��O����O���DL}Zw�[!�� ���H�&(i�ش�?i�dK~H͓�?.OB�>ʂ���)����HB�M�Ԩ` a��08$e��������I�?�ʯO|�P�^���GĎ\�|0d �B�y9P�i�
�a�'��'��z����dQ���S�Ūbi���֊#���o����I�ԫ6D�����<����~BL�~<`����T:n���g_1�M���?���x�~5�S��'�r�'}�E�3�?�>��!�� �H��j��dS70���'����$�'�Zc�,1�O	�_�2]�b�[PK<t��O�`�e;O����O����OH�$�<��·RY2���g�,B�a�o�IF�x�U�D�'��T�@�I�����-4Ad8H�b��t�9�<�I�4�Iܟ��'|J��u�x>qh@a#p)�NT.���.v�8ʓ�?�)O:��O���U���
jx���(͘}�r����;rՔ��'���'f�\�PX&J^���i�Oz��6�H�p�<4#�Dj;����䦑�ICy"�'1R�'�^���'��7��4��N֏N�t}����F9D�m؟t��ny2D�D���?y���2�H,%�޴u'�-XUNGJ�"lu��������8§�q����ly�ݟ8!"�
�9���#��� q��2��i��	F�y�۴�?q��?!�'3q�i��#k߬� @掍	���ȓg�b���O���t3O��d�<9��$�W"���#�ɑ7�L	��k�MCCj5���'���'�����>.Ob1x��/
HUaQ���h�������R)h����џ,��B�'�?B� �Fn�֮X�i�&a���}I���'�"�'y��(5@�>�.O0����[E�Y3C�e ��
4��]�!�fӘ�D�OL�D��OM�?���ΟT�I1g�&��#�*��ϒ0P2��ش�?��.�A��Ly��'���̟�(3G(�a�ǚ����@�]�uD�`cb���?1��?I��?	*O>�b�OѵBע�bkROx�PrX��!��>�,OB�$�<���?����|Xg��%��`Ȱ �P�a�# V�<i*O0��O����<�C!ZL�i�| 섹��W�f���wJ�W�_����|y�'v��';��!�O���V%BXTE _�(�b����M���?��?�*O�����\����5��
�H`,����/�ހ�sBO��M����$�O���Of����?�q`d��j�w���`!]z�m�ş���Ay��Z8�4�'�?A���� ��k�(�-����4��28^8V�h�	䟐�	[��T���'���
�G�-KSe�&	�,܀w$Ρ`���X� �#�F�M����?A��JvT��ݪn�B�# '�}�\)�AH�d7��O���M�\��,�$7�Ӑ[t���d�*��DlF�7T7����.�nП0�	ğ��ӛ����<a��>C�� Y�%�4����h�t@�6$0�y��'@�Ia���?ae˄N�>�"�H�C��������P5�&�'Lb�'m�y1�Ŧ>!*O�D����GL�+=��Y�D
�n� �Bp�>�/O&�2����ݟ��	���]20�e1�N�#��L� l��MC��p�l�YUT���'��[���i�u��AU�RPBa����#k&�x�&�>���M�<q���?���?Y����d� zS"�q(�<U��Uȓ�ԫ>��dj%%�[}B^����^yR�'�"�'�q�� uZ0�X�gA�b7|]�E���y"U���	��TybĂ�Y��,P��5��(G��Έ�l� CE7M�<!���d�O���O<�(�:OL����:�����R�
1���Uܦ��Iܟ�������'���Q�G�~2��C�*�/XtUUC�'oI\ɱ�զ��Ijy��'���'Q�:�'�s�#��R|�T��)��O�&�i�B�'��M�α鮟6���O6���70��a�
eq�lҁ�Y,j̕�'Z��'�B�� ���<)�OҠ��� �i�m�3��&{
�*ش���BK���o������O|���}~`M�~˘�9se��4sJ�S���/�Mc���?�����<�M>َ��ۿQ��!���,7e�!� -��M����.��6�'���'��T�>�ɾQ�4�#@%�ts2���HRC��ٴ��͓����O�⌀�_k��wA�i�'�?L�l6��O,��O�R��BM��?1�'���$�)fB��LӄD�F�Aٴ��M��M�S���'���'�>!R��EN��店$:PI�ԙ��d�����<v�b)�>a�������7X�����>'��i9b�C}2͇�A�_��I���y¨��
��U�S��\p���Z��EQ�0�D�O���*�d�O���Q�/�ҁ:�EO
)��@�B�M�WpSU�O�ʓ�?����?�+OH�����|:OP!�&r�"��	� ����l�	��$�H�I���y��f�*cŚ���9�%�� ��b#b���$�O<���O�ʓ[�l x&�������y��E��~H�%,�
)��7��O��O>���O�uJ�c�O��'v$�$�5=v�1Q�&E��=�4�?9����$��4&>q�I�?��MܵZ ��(]tڸ������?!��&Ix�����䓂����
9N�X�E�G-s(�`��!ǻ�MS)O��	���Ŧ9���.�d���Q�'�� W GhBGÑ�1�}�ڴ�?��*h�����OH��"� Q�/���
�?)����42n�$��i�r�'0B�O�b��"��I%L�<4��G�&�EQa�-�M�%��?�L>����'�0�R���
u� ��h� Q<V�r�Is�����O��S�}/�d&� �I�����]՜�Q!�>tv�Ab��2aB&@ns�	;/����sy��'���5�Ԉs)3�Ё/*�l+�ğ��M;�r/�Ǖx"�'��|Zc,����.t^�1ՠ�7R�h=�O�E�3��O���?���?�.OR��ǂIx� ��H�$�`����6Z-H��>)���䓘?!�� �ڨ��d��S3�-b¢�eҵ�.�<-O|��OP�$�<��L$��3,��J��/'ԍ�uF��r1�	��xD{��'��@{�''X�"d@�W� ×�O��1�cӆ���O���O`ʓ5�6勵��d�)J��0 �ص�<$���1M�6M7ړ�?᧡L��?Q���~ªJ(vH1���(<��lʠ�M����?	+OLh�G%IB�ß��s���# 1N�
#���$�1׌=�I��l���Rǟd��ly��np�u�2<&X�S�L(�|pz��i���'����'��'z��O2��5&I߇[�Υ�@(�:d��H[��
��M���?A&�F�Ԏ��<�~Rg"O�8����Q��UD:���W�����X��M���?����J@�x�OG2096GJ�t�b�{�c�v�Dx�t&x�Jh��	>�	�?c����)�J����� '�Y#�ʰ8%z��ݴ�?	���?Y�#�?!����I�O��ɦJ��`�fʆp���G��*?ԐQ�yB'<;�*�`��O��D�`t�IA���RAP�ǅ�La�en��T�V���'t2�|Zc
��K�'�f\�Q�G�g,.�A�O.l���d�O����O"�S`�q�!M	y��m@�JTVn�� ��ē�?����?�dpaKe8_�,D�D���>�`��q��?q��?���?�o����œ �p�pg�*'ZL$�L��M[*O��d(�$�O���	U,��i����W�ˊ�����+�$�8�ЯO(���O���<�2��4�Op��E�5JH�1�@�����c!�}�H�d�O⟘�g�2�ӄ�liH���A�JT�F��(>	�7��O����O*���/˧���&��#��!0�0�BwNKZ�bQ��U��柰��t����i �~BAD�k3P�A��:����@Ц�'`*DZ�i�꧔?��i<���#ў ���ą���n�:7�O\�Ĕ�"9� �}bq��"��]	"d9'�R�Z�����c�զ)�	ʟ�	�?�J<1��r�� >���c[-0)C0 + �A��iv����ğL��D�='��r�}@�p�F���M����?q�~�,S����Or�	(O��gi�n	�!���H�b��5�9�Iҟl���d#���UzL$`��0jת8{��7�M���B�Q�q�x��'H��|Zc�z��q� ���Cq��>�A��O
����O2���OJʓ<�Љ��d��4MfͲC�įNc�`$�FN��_y��'���ߟp�	��;�I��� )��焗 -�QPEBo�@���|�I��	���'�hU�P�{>)Q�3t0�e� H&�t��+z��˓�?�)O��D�O|�DH@���I)K45y��A#��[f/U{}r�'�2�'��I?@lfȪ�F�K�%ij���Y�w|�ٳi�	^٨�m��l�'�R�'��K��yr�>y���80�vi+rj�y���T��ܦ������'�7�x��'L��Of��Sp(	�Nࠤ?e�:,����>1���?A��`��	̓�?I*O6�/���i�䍪sF�1��ÖaѾ7;<���%�V�'���'�4�>�;-�ʼ�e�ȁIӾY�#�V>Zt�1oٟ��,/�#<��d���}��Ayr*�7fJ*��U.�M�5�]�RL�V�'���'���>1,O��K�G%��uQ��A�>Y
o����St�4�'3��)�OLP2!�Z�� ��i���[ڦq���X��0���P�O˓�?��'e��Z��A��Mq!A�!?@<�2ڴ�?�*O<p�4O�ǟ,�	y���$�>�����1N��s�R�e�ɻoKPq�'�"�'�?yH>���I?H��nA(w��+3����I�fUbc�h�����	ٟ���9Q&���#
~�V` @���A�Ly2�'S��'#�'R��'G6p���w�ҼBBC�/"`�P!gJ�N�\��O<���O����<c��
MP���6 Yĭ��-�:ot|�!��&L=�f�'���'��D].<��ɭ,c�
�a�'���@�Q���?y��?���?�fFH��?a���?�
0�8� �02���i���C���'�'�P�lr"A1�$W.#�Xȣ����$ш��!��k��~"�ֽ)����%�4
�ƫ�y2�%@\&��m�{���! �X5tp�M2�e��M���w�KQV�G�#MG�{�l�j��Q�R?`X��r���DMle�k׭wdD�{�(�LvB|��CY9D̞���Q�z�i$�� p%���mܻ[<��t- �X^ܠF�[�5x�%��W�`7@�s~�`�aA#>�ʑC��Cư,�aӪ]6�$�OJ��Ov��;;6�0�؛67 �1S�̘	�Ę��fW�10R @�
�\������Oe�'Ő�ҶL�x76�+2�I;��Ҧ�U I��\ɔ�:`֠S�]�I�x=��+�|�E�%K���݉W���2⦋�W���G/!�U�Ie~b�^>�?�'�hOYPv��:)���s�㗶U��p�"Ob��V?M�(I+�!����|�����i���?�'�\5'��xה�W�C/-؜�f$��S�
��w�'�r�'Vr'p�Y�	㟜ͧi����N�~�#���~����`D���\8�V�R����ϓ&�l����ڇ'�`٪��$utt�# m���I��4
B��;
ϓn��(�����8���?�(țt(������o�'��Ol髧K� n�6YYg�
^QQ@"Oq�����Ii& Q�1˂��M}BY���������O��cegK�?D�fN�l	�7��O��D !��D�O��S֬Sb�|K�j��5�
T�OgF�8&'N�����b,6O�!���(V��u,�*l#����#>.i��C߳.��i7��>�p<���Ɵ�Ity�Yr�j�!��*�4ੵ*B#Ϙ'��{���O� �	mj�\9j	�xb	r��Px�Bǻl���嬂��xtC$8OD�B>��ڴ�?y����݌?�����gW���V��L�+�)��P&��Or��P/B�l�v@�7�~�[>��OG�l*׋^�+�:���;2�O�P����S[����L�~ŞU��ڼS�ҹa��?�ɱ'�.(�tj�퐈aN�A	(}��ۡ�?y��i�\6��O(�?90%�
&}Yd,a�T82h���p�H�'B�^��g�S���Th�OvP�鐄Z�;""��<Ɉy2�iv�6M�OV�lZ�4R��@ ѩ��ª3yD1AaT��M����?���cF6�FC��?����?���ҿ!�B!]L����V�x����N
'Dh ۶縟��׍� v�$?c�Z'׆z4����K@/�y�GչD�m�T\�s���s�̒Q[��>5 a�<ɖ��x��#ՌX�_dT��$�^��?��i�r��*���,O����5V�\iBA$	8W��i�.Z�����>y@�D9��ɒ5G\m`��c��B��q�X�m�]��h�DP� ȲB�0G��G�� )���� D��Ћ��u����f(�ZMD�>D��2tdѦd/�=k���%8V�"�7D�,�v�A1��t
&��2M|���:D�(q� K	i(���JJE�AKk9D��;EJ��N�$ܩ&����Y�c�6D�� $�WB����#��<�D���"O�i�M�
�!�`ԌE�~��"O$˃��L�ddO�mrx$"O��.CҶ��Ʈ* �����"O�1s  �&����N˨<˄��E"O�XQЌ�^)ld��k
;Pj2-;1"O䍨C��BI9��U�-N�T�D"O& "��_�9r�"�'"I�}*�"O��щϺCd
1��=v+�ѡ�"O �J�m�#Z�|���	]�vA��"O$��H�<P�P���nH>�X��"O�J���T�f�
Q�e����"OH�!b��kj�lZ�
���@r"O�-�q`�3�L�
��a�h�i�"O����]c�>�; �T�X~z%+�"O
I�G@���@��@�s�%��"OF]�0��=�(���A�"`[d1�"O�Z�GL�?�(��`�:n^2P�"OP�p�̓.hNt)���
��ґ�"O�ْ�5�u�MP���"�"O<(J&)�6N��Y�V��yS�"O|m(�"�'o�*�Ɔ���"O|EC���+�f5�Re&k�}CA"O<�i�>/Vt!�qi҈N�^�y"OR�Qd.��Hb��kt�<�dղ�"O.C�I�\���:���,�<9kS"O�4Y!G�.y%�Ī���-sBdؤ"O\�p�ۂ/�Q@�n�3Wp|�A"O�)��#r��! �ѫ"�f4� "O�=�R"�w����KƝl�\��"OP��Nٛdv`��Ȣ��#�"O��7��פ���F&$�J(kA"O�����#&��A�"�����c"O�A@��r��B���̌�R�"O�Y�%�5R2��넏C�<��"O�0a�_9G����G�#|<��\��s�j2�S�OU��+���H0̴��Ȑ�zR,���'�D ���F�/:�W*(-]>�I>Q�**�0=�գ%���kC�V8;�A�!��M����U��Un���ŉ�
TȽ�����n8��&u�u���Ca� ��v���u�ER��i>s�'�>׶<�p���y�6��� 9D���v�C�g���O�A�>!����<�Go>���(�xIT(�<W�
Y�R���y�$"O j�jӷ?B�R��E)r�n��2�|B�D+v�az���/W4j�S'�V�lh7�{����9�n�bc*�0���\�j�L�A�<Q�"5X���#��.Q�	Y7���'�pub6�S,u$.=���޴%�hI�N3�C�ɱ��@*�Fɠ"4<	�A̘
v<�!�����i=Q�p��F�K�%n�0�7f��x�!���pf�Q+I�,�f ��PXq�'�v � �'S�Y��(�x��&į�~I��'[�0����`y��,�.i�b@�ˎ�y2�"L�ű�l�rvl\�F�G�y����2^������,� f ��y�,[�x��q䝰ZL������y��t�~����C!? �A@Ȓ�y�H�(�B�k���\r�g�H��y�e�$N��	4��� ��H���y"Y�D�y�%Q
hݢ��Ѕ[!�y�+E�<l*=c�e|��A��R�y&/wU�t�AÝV}��'�R!��'�txjL<��T0�.�fY�W�O+.7��{WJ 	����S"O� ��qG�*$:E��i��\�tԁ1@���!�0���(���)^�6�yr�Z H�����h�DB䉱T�<,��F2V�0�O�}85�'d�'+����!���R7C�&X��Ub�4=<��C�;|Ofh�C�>եJ��M����UZ| u-PU�$�1��a}R�J'<'b!��i��\�j$a#���')|��L<e&������� �|ՠ)�J(Y	`"O�̱����u^|��.��R��Eo���' ��P3��H���]5��u@ӂ��c���hQ-\�"��C�I]6�iE�<F;��h���$�打R<������6ZX����Z�'񾠻冈�i}!�$O#R)� �@�7��-B��$~X!��[=��t;�V�yL�(�A*�!�$�(K}:="�%N@f	�e�N[�!��$s\�}������|℅�/�!�$ܽP�\s�JE��U����T�!�D���t�6��%�s���X�!򄊫U� ��V��c0J!�D -i�to��V��a�O�<<!�dO�e�5k�i��,��l'��6!�ϗD�:ibpE.2�<5!�e�72#!�P�;�`���20�B1�J����y��P 1O�a����RJF;E��)��"O ����k�x`�IO���z��>� ���X��x��$��y����ӳDLd����yr���qB��Q#��G�NP���0gxQY�<�r�����'?� c�Ο#�Z "��|�J]Q�� �O�!`���Z��A�Մ;�l�%"�:��3̓- �Lڵ�'и"A�=�aې�/9�"�{��� i�n�s�öd��bE��|:P�B�B����59�Փ��x�<�{/�Q+��7�����uyB�X&\��Q��3��B̮~���`��3"��(�.!W�&��UmN��!�D�k�3���(	���u�(K ���V#L<�n��~z^�Z�e;��ON�c�O֨)���1D�z�x�oז^D$�QOV�*�̇%-(�:�h��`rJ�e��V �Ԏ��J6�	 �D�y���8ŨO�)xH�7kIzQh��Pb1h�;��'�<XT�[�XE"�G��M���P�X<BH�'R�<�x�Sᗴ�?�E#�B��l�V_8�2KY�_a��b�o)?�Ei��twRɢ��ǢM
��F��}�f	Kq+-�d�J>i�dI �LG�HxZ`*H�y¤@(ּ̉���?��1Ҥ�̚z����g�Ӭ����7�-�N���4�iR���'<�!��,��X��T2[LD����u<� �[\p�A*�P+���`�X2	VRL��	ߎxd����W�K�$�d�i~(�����G�	����
`NI�S��X�ax�C�035 qCuF��n>���+��,��K��ِJ�yA�fޤt{��;u�/$�Ař?4RjdA�@J�����-4?Ʉ@��j��p �)B� �(9�NZ���O��9��b�m.���c 6e܄8�'Wf<�� m��prF�"G��(ui�YH��	��)Yb�P#req��'R��Xr�M�[8t�P��9��- M�'C��i�a*��~�d��r^:EI��s#L ��,�G^�J`�P�,ыz��zҮ��T�!tK�����΢���/9`2p8�{�.TѨ=(�ȭ�����ݶOR�tK���-�@�b⃏,�!�$�wo&�+�
u�jЩu��%��'�z����ERs�n��~҃O�_50�z���Qn9��p�4�F���5��I�~� ��3��,���ELi7��	���Z�A��J�/.���I�9~@"|
����?�Al�9n*�!�W&Q�7��C��Q�c1�4��"'NV�_�J�b�F��)ݸ1 �cG;"d��A��f���	:�ʐD{kH�>>A�w9����*�0=������A��Ò��m��[����R��cL�sì�<X_�����i��8��ɴ+/�M���R�2b Y�*\=8�O X�"Lx�M��jj��r�E9q����o��ih-�@m;�8y�  ��{�!�D��τkEx-�6���d��\Q�K߂Δ<+�x,�2���$�|K4?�OҮ�˙w���(��&F0��E��D��	�'���Tݒ(�@��&�ݤ8WTH�0�dB�k��x�D��h�E��Tm�'�T\�,]0F����a$9o�p��ۓ<��� �% �|��2� ��a�l�'u̦�bT _'<��!P)�;&IFxP�d�
��t�ī�{X���'�N�vr̈s%��'D�So/��)rT�ٗ�4z���3'ƅ�s�FO\��C��� Mc�eg�V�؇�`H<QSF�??�@�`$��-R�`1U��=u�����+��P�&�6UޓO駻y���.�Vز�oA�7�&��怽�y�o��
N��`��[�	Z��F[|&)%���NK6���L�*v���ɕ�5��d=��p�)n��D��F�|-���,�1 �cA#|IzY�4��+[D����Ȍy��3E����
��AO XH�͚HM_x��s��dY8���8�l���H8Y��#�'k#K��1�
��<���}�T\�/�,K�u��"@>g%F�a�'c�hǈ�jxB��`��c0�*1��6h��/�J�> ;kـR��)���E�#нp�8W�>�l�r1"O4=Jd��=�҅�wa�RuBUFÃt�&�KK�tj������i�4a��t�תX�L����ҏҧ-N�tf0�O�u� ܀NpZ�i]N��[��?<��{� M�t�@cˑE����	(\O��ʲ�J"Z��������1@�� L@d�T-X�L@Z.r��M<h|B�BF�#"��a #A��N]�ȓ4���b�J�W�����؜h|J���lF��{�b�!k��̋¯ľtv����94�-�"��$2햰#A�e��?�"��#8`�?mB��YP��2��0'������͔%^хE�
S)�q�9���'!#�O�� �
7�4�j����
�^��1�A���b��E��̬}��|��H�����0��	������9�x��X�0: )lOD
�KT�ì�w�T�J� �sp�'�TU���+�DD�1TT���[>Xe�D�9?T%��)+�Q�A)�Zg�;P�[1jU�@��I��5�.OD�8���h�P��խL�_UܽCcP�@��͎.�J��b�*V<;��'ҧs��#�H�	!�5�U���*4�?�pV�b�?�.%��0Z��X�4:y{"�ڟ	�~VG��,S:]
�<�U�ߤ��g�*�2x�d��:*���I^�d����+����'��>���#�7��H�ܮu�ޠ��C]u1�l�t���G��'�(7a{�*��}�19g�ؗW�쌳��D��y�i�w��#<!��O�/��Y�!�t�L�m�{���ST�
s�8�jSM�PټB�	�?���,��C64�:s�jM����׭<w��qf�S�|4L{�c]�b"��:��\T,C�	�i��@ ����6͘�bZ���6^f0��CFY�)��<c	]�Br�	�B�����U Y�<�v��-�!1r�L�<Szeʀ	]V�<I4�p��@�A�U3Ut�D��J�<!���  ���!Z.��|�T��A�<9�kA9g�J�s��(2@=ʣ��z�<)��?a�pX9 ��*U��!B[�<�v�A�<8��ZSG�.�ʘ����V�<�bE�#T�j���O�806L0���^R�<����`C�ţ�
�5�̠ä�B�<)�"��k�P�9�E��-�mpF@�<���X�N��� &ׄ�@(��Xb�<	�*&c���e&xP� �G�<� O[]+L�Bf V 8��3U��Z�<9���!������O��t�aZ~�<!�*�7h�4�g��dǲ��NA�<	Pi�j	LCe�YQ�%�H�@�<ArER�0t�ܡ�!@�.�m��z�<������nx�i�>�jTq��\t�<�R�2eC*�{�/�R=��X��n�<�'��WLy��=+
�1r "T��	BKɫe{�)���f�P{`�;D���F�fR��Ef9#��@�S�&D�����ۼ^��tqD��4V1A�2D��q�D]�Pyd˵$�+�B�:D�+D���!�@:��0��HT�0�H(D�P�c��P�N�*�Η�C��Qw�2D��J�#��rtQ�b�+OD�<a�:D�@2�D�C��#��G���B�,:D�@y#`��t>mh�gN�|���*ǎ9D�Ԩ6��!�4��JM���`�f9D�� �5�����QZ/݄DZ���"Opt�#�35��	w.ɔT-H r"O(�"$��	lL�$�[#H50$"O�	��W
7u@�3�kD�@�T"O2���"FS� ���@�dXQE"O !oU�D�'�Ⱦs��X* "OT�:Ff���ȉd����"O8T9@�� �ġa�"���"O����&��}���@�S�s�Z�s�"O1����.�q��E�F)J�"O&e��	�Z
�Q[£Ǐ?��1"Or����=$H�#����F�`%�t"OBeS��ӫ��8V�	�C�n�"O(Qh�1�~aS�+�$d�x���"Of	ɕ�̺h�dH��%f��"O�@ȁ����֨��CW+�L�"O�aG(T7n �K��àl��B "O��a -��8��q//r�V"O�l�c垞!zR�3�M�aՐ�"O�!� C��k�(�A�Q�&D�D"O��^ �j���^Yڰ�"O�!'B����Ȅ-S�K��A"O"�aaXU:���m��>��e"OD�bC��
���I��;_��"O�kg�
5&DP�I�8i�"O��J�f� "E:S������Y0"O��A�	�RW,�맩�1-�`�"O�`�FX2o�����gS�)��!�G"O�x�t�J1q��"��X�d���'��%��+�R�`QI���0�'x�"�ڥ4O�1,Ҿ>
ZE��'�.eZ�j&WnJ�9��/>�J���'yHl�#�L9b����Ŕ;<z��+�'�N��.VS�^��G�#9�V�I
�'�~���h7m��|q́�>�,�1�'��w�Qei�I���%1v����'-T���n;FKX<P�Z�R�Z�'# 10S(_*j�kWeW4NL���'.H�F�!h�pegn�?l`��'G
���I�m�F[Fl�*'��#�'Wb�%�߇S�T�dH
�i�"E:	�'kZ@rw�%��@D�C�s#����'���УO\�.�lx�Β9p��$��'d���.��	(x�`�G�=�
Ւ�'�\LQA��l��4"D�/:4�8��'^�@i'�N�/��%"��܇5�
@�'������Xb
})#N�3,��q�'R�bI�1XHi��]�.>�Ɉ�'��h�FH��?0���\�����'s~tQF�
&wiB	��m�$P�������*��)*m�o]*��p�P&.�!�D[�c����o�+G|�2#�5.�!���dHl��j��\��a�k̑IK!��&ytֵE�S�_�a�TDT$�!�DA��9��އ9k޹�q"�?&!��#�J�$��:HUX��b��V!�DL<�.������/�����i!��f��{7��@�de#'��5K�!��2D7�}�EC�&<�Z���E��~�!��<H��en�7��m�U�m!�ď&e�Qq�B�<T#�X��
�e!��HJ���F;zr�x�cP��!�$U5'�1� Jjo��ҩĭ)@!�$?[E�8��g��y�����N͝F!!�� 4�ʖ�
>m1
�x�J�,� �I�"O���j��J� �3�G�>�D�§"O�iҗ�X����G
1�`����Iu���	��&
�����W��ECb�V'!�d���Zx��dC�R����g(�!�d�
�4\s��M�4���fN/L�!�$بs�`�,�6�@Ec4�P�]�!�d��O��h& X�G��E���8/�!���ʪ0(0,��r���J��Ҥ�!�����'�
�V�z1`i�!5�!��s.����O%Y�F@���U�	�!�߻��x��ށz͜Yxa�R1k�!���B��h��ޯ,X���9k!�	4r��3G.�5j��	��!2{!���a��8c*��:YR q�
"Fl!��o>XT�T :��!+��W ^!� ,r쵚@�N�@��1dˏ_!��@&�`��n��1(ZA��h�=6X!�V aw(qc�,ԅ3q'��!�Ps��S���T���oZ	�!�d�Z�f'��!��aSU@�[�!�$�2>�P0�0�/N��A1ae!��O�E��B4̘,i� ^7(:����"O6������O�ب!�Yi,�$��"OL�!hG�k�n�yŨ̬w�D�:�"O���a�W�*HE��҄%"O Q{ӌى\�,$C�M9~�>ŘV"OrQ;W��*H~|��q�.-�-H"O"�1�&7O�PjU��%�6L�"O�Hy�%՟z��4	Rˊpڦ��"O�I�v�ڬA�&9��J^���"Ox�6��o�~e�b������F"O�9� b��F$0�U�2��\��"O4X"%E�lԮ�3.Ǝ�2�i�"O8ŋ��NG���GB4���"Ov�J'f�qnD�F����I�"O�z��´��`R=6����"O��0�;�|P9�[)",X��0"Om����tm��Ԭ�;��U+v"O�% "�˅��m�	��l�"OHM�懌(��j��FG�bF!��y!���w�l��7�=�a|��|�#yUD9�B�?q��-�`H�y"�бad�  k�,3�|]9ceˮ�y�ś%�p� ���(U��(�A%�y2��M�V� Aj��k��Uң���y�Ʈ��!%' i~��뒋6�y2�]nAi����c�N��b�U��yR��Y ��T̀?/��Xy��
+�y��M)&8�X��O4s�̈�y� �*;[|�0�U�n`bwo��yB�O�AȾ����T�
3Hy��+3�y2e_&i��8z`m\�{��)c���yb.�8]��Me��f�2�
SG���yR�\<}6�@��?6�y ��%�y��3����)��t  B��yBA�b�j�Cu*�4�S��N��y���[p�9�&��fP[�N���y�ǘ����(�a�H��:!��yr�Ɨv��� �;=8�}���V;�y��3��� �i�#,���˥+݁�ybA'=X��5@�=�8���G��yrj�	l&��&L+}s�y���yrui��w8��*V(���p?q�O� ���Z"kY��Y��дY��9�"OV�ڦ�͛?|Պ�C�
* ��"O.I���J�V�%C�#�>\��A�"O���k�,"�x� �$
X�+W"O�\�Ǣ\�3��tC���*ɜ}3a"OJ�;f��XJ���2D�ih��Q"OXq��f���p�A!r��Y�"O
T����"�N��$E�5a���"OT��P���z:(�I��QU�h��1"O8�`$��=i��\4u���"OL���艥L������^ ,�a;�"O>��p�L�\g�i����@�)�"O�	�g��Q�X�36�h�!p�"O� #^�ZG��3 y�b��"O����(Q!�`M`q�E�ش�`"O�$�'!�A���"�!~�y�"O��Xv˝Tb�`�p!�P��9#2"O�I�� �:>�,�!�	h��x��"O|H�*?B�p��b V�2�"O�Qs��!���V��!��Y "OQ�2��'�쭁 ��,_�� g"O��`�ǅ�0����A��&дx3Q"OĤ$�ׂ?�Lz�LQ�*����a"Ob� ��x��Tp���X;���"O<AY'�T3hX�dx$���f1�P3�"O�M�OM#��� �'��+ hi�&"O��!�FYF��;�E�.5ٖ"OT� �C�-����&W\��"O�CEj��T��j!/��@�D�3"O<qb��#LŦ�"�nC�v`��"O�h��^�N��B�]��� s"O�z�$�&GS&�Y�KށE��2�"OR 2󋈾`��d럊,}3�"Ov}�0K� En�x���{�xyYA"O��IwE�=D�,="�����E�!"O��iS�s%�� ��^,z�(�"O�3 h 0i�Д7cO���e�"O�ع@C)#0TŪUG��p��!"OP�٠�ы�HJ`F7n���;�"O��� ܛ$��$�T�Hx��!�"O�ݻ�C
,{��I��.�"i��m+�"O.)�t�s��(1G�?X�2��"O$��ɒhI��r�K �8� �p"O*lhe�͊Z��eH�o�
@�9��"O<��N9L���j6ُ@+&$�&"Oz�pl��n�Њ%�¹}6��"OX�2���Y ֌
siѰf����S"O�$
�Aڒ{��|0`"���"Oā�P\8j�	��ሏ�h0�d"O\�������n��$�s3"O�����D��\Y��NI��s"O¥��E���:��_�%���"OXDY�%�(:��-soO 9�T*4"O�5cK�H�Ҍ ����(�m3"O�嘕��?�^�tOګCfH5��"Oh���IC
W�1��@"d��"O�p5�T�/	l�:Ө�� �"O�Xf I}�<4	�g�O�2Yrd"O���DaB���z����C���!U"O�B�!'&�c��$z|1(B"O�l ���	ca�)r̊���T"O�I#W��9W�R�ӄ텃����"OF�1�l�T�n�%�����"Oj`IE���̼�X�BԨYz��"O� ������3z`�H�qcC	���"O.�aw�ʡ(�+���_� ��"O��FBL_��QP+ɰG��a��"O
 	�B?�ĐuiD�c�XI�"O4l�6�@�.Mx]X@/�=VI�@"O8�x2�P�F��!QM��Y� 5�"O�(���A���땟%̌Ej"O�0��<�9��,��ȯ�yD˄�`���MD�Y�h��I�#�y��I�E�~X�#�T��prД�y2��|q���T�4u9�t !�D��y�-L)Y&���e�7��m��W �y���Hk�uB^{���$	 �y�X:c`Бh�A-		6=q�F%�y�h�m՘<�R���-��l
d��y�"I��BU��9}\��*C��7�y�J���tEJ�(t�D#�I!�y�Nn��@ '�'rO:4�r
���y�3`
�L��Ϊf$s2
��yb��*;,��J �`"(B�i[��y�KA�J���V�b�����I�;�yrlҖ(�x|��ȋ9X봴����y2*6K|:���BM�?����,��yr��"{~(ەl=m�\�r*��y"+�,2 6� ���%c��QAG�y��A�:d�9��_�f!Ӂ����y«A ,(���*ǺP�ȴ:�a��y�CH;/��ق�Ԭ(`q��j��y�ǝ���Xw��#�XH[�����y��ϛar�����{ؼ���F��Py��Kԉ�W)դk�H��[�<i3�ч3�� e�J���E��S�<�eo�) �n	���L�T�@a?T�4�G�O"��8��)A��A��#!D�<�u�Z�疝pʅAФ�#!D��H&)FK�P��P V��"*D�*2���\U�$9PiΑiX�Cj)D����րd��� �o#7��Bֆ(D��(�6q����
�_��IQ�8D��B�� �f5 c>v�����i3D�h(�Rl�TP�ڪ	�8L�R$D�Hsg+&��$�e��1 ah�
G"D�`�����;�%�R 
Su�%k��?D��c#��6�����L�y��>D��swI ITZ�Mިa���i��&D��rŃ��Lp�Ы/A�5�`ш��$D�zD��K�Ⱥ�(�=:ƈ�;e -D�,��o�3, �H5��C~Z1��9D�(��h�%3�޵���<�4Qx��2D���rm�6����'kY;>i�/D���#�.&�HjS�-	Z���(D���SE_�X��dI�f V$�m�+4D�h`!�ߍ%�����2T+�ءF�3D�D�($�%�+ɺ?X�̸p5D��	���
�����Z-|��rU*3D�$��#��'�<%��D�.�D���n0D�$ke�ȽR�Fp�0��G����k.D���E�PTX �G���b����6�-D��A 	�?K0\ �(J�ts����c,D��	݊r���8��U?S)�m+b)D���B�^�:>��Ժ��	2�'D�����/5���k�0?cz�kF%D��T
T�<DM�VMʒjA8�3��8D��Ça�o~��1��A:�L�q�:D�� Z�� �_�i=ԁ�"!|T�Y�"O\	��?"�z25"]�fE
m�3"O�0p�&E�A}�1P��Ύ+�01"O�*R�M}0�j�!\�}� ��"OTdf�5AP@mR�ÈW�D=:�"O ����4�d�K%�<� b"O�`��Kґ!�$e���T$��x��"O��3*��H�h�A�	�H��Q�3"O��"��^-n���YOF-+�"O�,�bBW�N`񠮆�wK܈��"O6HksB��D���G�nCH�6"O���,�:<���l�*1U"O��v�K��J1�&�H��\��"O�ГaB3����I�%f6I�t"O�)0K�V(@�!���m�x01�"O�5;��R?�q�07��1�"OH��5N�'`V���;fj�,X
�'�� x��Bm��,9E؉+���
�'\h`�G�9Q^Y��c�3 � ��'�`��$D|U��(�C�J�'�<9�E�':F��+g�,��`�'�pؒF��-U�+�%�"#t0<��'#$QS��[&[�.)F�k�t�k�'8�E�U�U�tƊK�y���'&|��m�aI���X't�B���'v"$b�搭}~�Xv��v��	�']�ĻBn�	�¡�U���bVؑ��'::��AS�, jI%T&D�r�',ƭ�V��l-�Xu�N
PO����'Ր��#Ͼ�3b³O��<z	�'��m!�j9�
d��˳?�8�	�'^��[g�F�oF4l(wgҜv�~݆ȓp�P5C�%xB��#1���A��l��zh
]pl��lJF-���X��Ň�C�&�@AZ+�����.ɖk��B剤�n�F��4NSr=��m�.p�C�ɕy.��� gK�C,p����gP�C��!gjt�`A�&|heE��lC�I<<9���n�;�>�7�_�d�B䉓iP9xw�!��P0SG]d�B�	�+P�}�%�U�R�,�b��B�	�pԥ7,�96�\��V�e�B�+k��a�2���ep ������NB�I�U�.���P<Ҵ�H�f��+�$B�	����]�S��Uzd	�c6B�� 7��xc��^B�~�"Ƀ�cG�C���@��ym0�!G"_܂C䉇!~��oTv�Uf�ZH�C�I$C�J�;���@J���D�١5O�B�	�Ilp�g�2���e-�#;/
C�	�#��h���"*)���.�8�B䉭L��9���"_3`�ċR��B�	)��#�'ڬ%q2��Sa�)��B䉷�Ԉᷫ�*{��tHJQ+��B�	b�m�W��8��4�	ۯb�C�I.F9h�h���9��q�D��N��C��>x��$� -��*A�q�	�#s��C�I��(}[ī�]���T$�![(rC�	�(f,��|����/��wdB�I�t��ڡ(s��2Ӗ{��C�I,V�����8��Xp�O�J��C�	�^d�)U�#��"�� ]���0?фo�-פ���M���a�s��t�<���҈G�|�҅ܓ�0`�"�p�<� ��I$�ߚyw�4�D�&"22:�"O�%��ՠؐh�b
]�0"O��)���w�^�)f�\� Ӥ�8T"O��T�	�^T�9��"��{f�	�O���e�	#�였��ޠSf ���'�
��gS=X�(��`ьJ7�{�'7Ĝ�ӧ�(���i*+B)��'�4���9�x��)�$"�9	�'���3�۔H��!N_/	��p�	�'<&,ۓ�� �b�f%R��5��'^�U�aã.EbP�G3BXTq{�'E�T�JA1@�9 ���6��q�'�ΔȁHԭS Q�#�n[�'7dI���^hxs���P	�'�.�r� ɁXHT�+H��(L�h�'$�qYƬۢp�"�z��%���@�<�QG�	��<����j��Ԡ"�c�<��!$|��0�
�z�f�p7�]�<y��R�S�� 4��N�<���d\�<ËU�V`�#D@4Md nY�<Y��D���!��l{�] ��HX�<F�בt�����51�X�dQ�<���6x�M�uH)l�d��7��x�<�%J��>����ċ�;3�C
l�<���Y4z��Dn
�K���bD�Q��y"���%�z=��J��ɘM3t���y2%�:8��B o�s�UXI̐�yr�aBE��ā��4X�.��y�d�p��Y>�Y��W"F�=�ȓ&{� G�/dC�0S�lK)&�f���e�2��_��n��7m�
�p��,b�,٧N��f:�� NW�bX\��	ϟ�����C�}R�n��i���rrB_{��O��=�}��cw�p��Kp����!^|�<Y��0d�D�!��6H����I w�<��͕$�ڝږEK�G�By0p�[�<��N(f�>R�N#O��S��]~�<ٕ�ՐO�A+pKC�b�\�cWR�<!0�I�M�:��1���|�R͡a%��T��\����+?��I!)��Y�¥B�i��$�Ŭ�N�'a���94�˴&��w��8ǌ/�yBѽ'o<����A,ı*�,�9�y"%�O��(#��:ݺȁ�*�y2KN*\�~���%�*���p��yb���\���&���ġ*@'��x1x3>�9�늕	T,�҄�R[�0��*n��e�c"M�%��C������d5�S�O���05O��c����4M�7"O�����;}�4�0��6s���sF"O�� �#�?.H诏B0d
���U�<� �4$4Ѩ��7�Xr�,Gj�<)��Bl�*�!����D��`\p���hO�'ca\E�f�:n),1�ƩɸS��ؖ'o��'/��$+��a�.%���v(�:��zR��A�<�'�:A�@�9e�[#@�y���A�<1�b�<&lj�
#7���i�<��B��1�Nh���R
��%�d�<��O�� �B�Ύ�|0ش�%a�<�� �P��©��"�\�ro�^�'�?)YC�ŪTJ�<Qw�H,c�
hz��,�d�O���<�����k����J?i�1Qj9"��1;�D%D�0롂U�v��(��Y�e&�`�"D�t�aG�<4��h1j�w$Q�
<D�`Yh[�RDIQ��
!H���m%D�� @�����g�V�3t�Q>.� �"O4�:�oN�[D�I*!�XC���b��|��'�t���l@&1:�kIe���1�'����%��3K�2H�nFX��J
�'��9���S�n웅g�K�"�{�'T�H9�ƠK�d��%F��6��}A�'�Fј��>zƬh;U�9.���"�'D�<�rB��?SDT��G���Ti!
�'M��s�͏?������6ظpH�'5�k4��h��(��.ۋpA�P		�'O萲����ڪ�2�@�<i$��'t���E����2Cۚ1ܭ
�'"�����0 9TXA�+"����'R���sfЬrܱK'U���`i�'	2@�Pϝ=�B"a_!D�ȡ��'5�-����N+�̬f
�}�	�'��37�*x&��#�^4	��в	�'
|��f5X�"�xCX�z��'.�	���:Z���b��Cjt���'M4!I&cäu�DyҌ�=5���	�'cq(�*�0��P��у/�T���'jD�� �p���j:*G���'e4����:H�\��t��7%��`�/O�=q���z����H�}�ȺN�w�h0{�/D�8�B��izr5���KK\\��N-|O�c���D���+!vXٔ��=c%d��*D�h��k��j��B��3s&����)D��X�`�'!:0("�����Q)&D�SħS�S[��[4�N��!Yҏ6D���D�;<a� ��E�|#�=���OT�=����,7��'f�*P�:��th�Ȗ�L��l�*!���p���F�_.�0Q�!��!��5n�mbfK	��Hyr
��o�!�d F� �£�@$l�0�kb*V8Jk!��S�F�J������\�1p���ZZ!�Ƕ[���"�M�7s�b�@�ʊ8Z!���2�6�;kJ�V�ڴ��O��i���'�
uY��ɝhϠ��W��9����'z!�Ğ�W,�B�ˏ$/x����8!��0va"�J�ԇ]p8��+B�H!���.��U���>2��a���|5!�$ێ� ���_mҦ����O�!�� %�:�k��>�D�sr!�ב?���Jr�7�(��K!mM��P:!����7X�����^�WP��0?���׿d+@���A|
��6�Ay"�)�'E���R4+�	q%L��ES�:C��`��:�C&?�V��遌xc`T�ȓRsT� H!x͘���l�Z��D��IIZ�:G��jC�����F�DrN���e��=�5A�C�u��.K/�����.	Yש�3��0�%��:��(�'�ў�Fx�&c��ҡ�
�����K��yR�1���A@�<3B��v&���y���g����-
��Zf�
��y�-N�[l�;'/֛nG�)��'��y�`�F:N; A�<�p(+��-�yR��,70�j�W�;g��(�.ɿ�y���;U�ȍ���(. ɤ���y�>A��Ƀ��4�&���g��y"%�)I��37nH�1%��+��#�yR�¾�R@�5�W9S����'���y2S�0�ؕ��X$E����"���y��[�h<\U�$aX9>�x1K��y
� ��	�mW�Ex�Az X�
rZ��B�|�'az����`D㊛O܍���@��y�_�0�b6�$|��I҆���hOq�
(	Ƭ�%/T��O����=�"O@ݛ�'6�H�p��Lp~��"O�E{t�]�_��tҕ��-B](�r�"O2ap!Â-V�K3�VN$�+""O��X7A�lӀ��YB�-���|b�'���#5J���O�9����6͐��!�CoI fFw�`@�Q�߼ y��I��(�L�Q�/�(D���p"�y�"Op����_ ���JˑEW8̐�"O\Dk�iU�qz0<a&I8r���*�"O5�Ί�P@����ҁb���'�:����{�&�ZG�2]�B)C�'�2���N�Ԝ�f��7V����/O��=E�䀪�f\��MU.1F�P����?���?��<�š�&EvL\�p�F&'j�{i�Z�<A���iX<��FOА)��I��K�<�Ӛ34�J��V�fPb���E�<�D��$-\��D��xU��"�Ln���?��o\XGJm\�pV��1N��5��ئ�C�mצW��X��,+�PA�ȓW��	�茳3�% VD�Gt���ȓOT�!��*B�JaL���VNm^؄ȓ)'�P�sB�r�H����KѺ��K}T�Z(���Eg��~�21��Ӓ'*�<�x�J�+[%O�2t���O�=E���/U8L#��7D���'�өQ5�'ў�>}8p
�=l�!Э[b:H4�L7D�x���KB�Z8T-E,hFLs66D��DJQE<b�ȠJ�C�Zh��2D�`��e[&�p�d�U�^�)�,3D��!B�.tY���F��$A,D�p
�呠n���i��Yʨ��$��O|�O����O��=yd�P$O�B��4L^"��}h#���?i���'p��`��ǲ�̜�`�L"]�ȓe�n��#�,hkn4diE;1��ȅȓs�D�qp���L�.�{��S6���ȓ�|\�ĤٝZ�x\suK�1{ؑ��9�.�A�g;�<u�G�ǖW1>��P<��'��"֖}k2쐎n_>�ȓ�������B�Q�"�(�H��'*�':�\"��O�1�&����hR�'��Y�t^�0�4�#���"�
�'�P�0N��_(�٣�N��y��Az�i��t���F!!�y�Gb��å��
w���K���y��H:\Y�)R��'p_��TbL1�ynH�t;e�Y�dlL��!f���y"
P��YeÖ,XZ`�Å��y��!
�h�x1��Wդ�3B*ׯ�y�	W1�s� '^�^0�1E��y�@
tH�DلbU�XO<`Q�+�yb`���lp�G�D�U�`�����y"�ʭ%H��[�K�29G�9��F�7�y�l�f�N=�E�]?,�	q���y��'c\�8j��B�bF�S!=�y҈
fi�x���tI.(á�R�yr�˨@C�9u�<j��Z�"V�y�A].����2FJ�`�@1���yb셍c��P:�(��-6��HK��yr+�1�R�`����$*~�"L��y��D!2�]a!+�$0LHM"QJ�y
� ��I֏
��3G\� ~h�0��'��3)J�9���P��8�e��g��B��%k<(�14���壌7"�C�I���ۀ"A�a�
��d��7g�B�I�wj�J�<MµJ1,�7@�B�;�*�y��(@�U	D�)c�C䉵D�@��h`�!�ʈk���H��	�j�2����Bw�B�T�J� ��B�I�'�����bv�9x7K�,���ȓaF$��B��<r�S&��t��8���pQ�F�D�����'�ń�	;��+b�8g!�ӫ7/*U�ʓ*�‡G�F�8�ird�<D�jB�ɑ*R� � W�&+8�0��1�VB�	)o�U�!)]3K���	1GđQ�����O�a0��ׯ$ʆ)W'��X6 D��%/�*B���aL�;'Ф�;D�,I��Ʃy��"�F\o���b�i$D�a�N� s�����3W\ Z�K'D�(Zq��+R�` �B�6"#X��� D��%�3/"<�p7-��S��	)D��"�a��W�@1/I	����%�O��D�O���F�1/d���T�G6`n~���&!D�����$=Ob�hA��99�n���,?D�\˓B�M�� Q)��m$X4�w9D�,Q���T��]���V^F0�D�!D���o�`�v\�ec3r��*6� D� 	a#`���� Q)Y5p�`�D4D��P���"N����iХ9X���?�O��d�Z��	Y��^l�|+@(����C�	g��\�!_�0l.i���?P�C�ɤ��H�4��\���%��v��C�	�~�h��5,Y�A�ؘ�bB�+_�^B�ɑ�y�
��M~���j�*G	*B��$>�FMa2a��M�t�B6�*$*B�7L���O�U�&����
W����z�`;�!�(�h5k���+J��	�$=��K���T�'b�QV:qM���Ê�{5ja�u"OT=��݄>�Z4y�@�$t�:�"O����4gp"��n�E�H�"O<�*@�֨�ȑ	5M/.�6(��"OL� H�h�8��%�˃�ע$H!�$�T���7m��R�*H!�I��d�!�s���	�E,q��˦EL�N��Oz�=�+O4�jU�(�| +���80K�hs�@�OrC�		���P� ٣6kbБ�FǛb�.C�7@^6Lr!/�_�Z|�����C���̘���S�S�p�1G�Ήv�B�	�O�Lzi@:2*�8Y��L6HC�so>E����?�p�Ŋw�*C�ɥ�̔Q�G��l��T3A��=�H>����J9""��ۅ`�Z���8������$�Op��'gǚWB]q�u��C"O8�k ��g(M�sI�!j�|@�"O�I���Z�zU��)�Iy�@"Oƹ�BO�����лd
>��'Բ�s���:��L����v�1R
�'�0��Ņ�\FeP��\�h ����*��p�΄�N'2�a �@�z��'w!�d�DZ.�( I�q�9��]6W�!���9�����ƘV<��	C}!� �ᤅ[����S�^�Y���]m!�DS�L�zd��܎H���aţ o!�ʳ`�b=���'`4޸XPb�t^!�� F�J�l�]6���VO^2��9��IH>y��6L����D�Z���bv-:D�����r�ԭ��>c�ĩ�Q#;D�@3fðzD�h��K�Ab1*:D��� N�}��"�疓b좥�e�+|O��<?�4�/!(�'� ����'i�i�<a�J5�h�f"_�Nn�|�<I�ϋ"dڅ*R͟1�D��a'v�<Id�(S`��)E.��v�.}@R*�J���hO�-��̘��Ņ��YD(� ��ȓvH\m
���w�r;��QRч�Ej��y�i��֝:Ao�;Lr�1���v~b���n���G�NH@�1W��1�y��Z7f��Tb�?w>�`&.��yrO>s+j��昤8a4݋e�;�yR ��	�nX�F�ڠ[�����?���0|"�$֣z�tQh�" �@��5`�I�<Y�l���x�Z`JA�(:�M���Q�<ђ�29*F�[`eڜP��x#Du�<q�J \�\�yA OH��IS�z�<�#���D0.�HU��3A���f�u�<E�Ń>�	��%4��rA�^����?9���O��2S�8"��Y�H��y�J!�DL�@! D�|}̘�rmU}8!�$RSG�Yd�r
x<��L��x�!򤀉f!01� Eי#M�r��<(�!�D/�dH2MD&=��lS���Rv!�Q�2����J�*
,"�FО1S!�-}>�`K���u&
�Ge!��Iy�ԉ�� �M�BdΟ6!�d��zU��wD�ٔ��:�!�_I����ŕ���h� ٶX[!�$�+�p�	��Att0��
�8^!򄜚R�(=�Q��xT8��f���!�d�F��)�cO/-�� ��Zk�!��úq�>@a�	�	[�`:��*m����#?(��G��="��D��\f�B�ɉj�v�Z��[�sVD�T�,�B�ɟ\&}��.ٔT��Ce[V��$Åa�M!��)�¨�!fĀ:(�'vў�>y+�&Q&eF`k�ɚ�`�R8y�a#D��5D�Xb��T+��u���qN.D���C
Ō6�Z):F��&~�����L+D��+�]��D"�RYpƁ1�.D�����N�8o���ǐ�G>Hr��+D��H���5Zz,Z�jN�~wE��3D������s$e��J�@��q %��9�S�'A�荛aa\2R!8l�5H�2�̵��~8��(�(T��X]:R	�6B�ȓ�h�uʉ��n�(���*$fŇ�S��p׭�N�������7�ɇȓ.�⁹7�G�!�D�
��(��`��c��İg�F�.�t��˷Mg���ȓ;*i$����԰�C5'#'���IS�Sܧ=|��J�g�.����l��ȓU���0���+k�D�4��TqBh�ȓ	F��+/�<p���4"4~5�ȓ%�ؐ�g,�;^�$H҄%M%�����;1"���Z������T$\��h�ȓ;�Ȩ��KX��X�▥״st������Cɸz�@��!E��q29&��$�@��m�O�,;%��2�TAy��ջX_,��'0�1ѕ�C���3-9ϐm��'S`�i��S������!<ޖ�B
��� ����A�|����bT�
�3"O��A�ӤI>~���V�O�%�"O*X���3M���Q�^�Y4q�"O���6.��"rؔ�Cb]i�l��u��m�'���9g	߯@ޤ��C�����0��"OYx옲v��(X������q "O��Z�AA�h% -��쎜G�V ��"O��k�?,(��C�ۜl|�z�"OHa򧤃�t숍+���zV��"O���"�$�p(��+
/EH�Y�d"O�	9�i565�8�aɳvA:�@���S�'u�D�I�܉g��3 \���LoRO�`�ec�urqɔ���:S"O���4�����I��]�p�	q"O�A:P�ل�F%��I_�k���2�'�ў�I�<&�T��J�y��l��M�ul�-{`�Og�<	����(�� ����"^X�<Qo˿w��� 5a�!g�Q�<��i��}��Bh�c�\*6AhB�	�K�x}0Ī�)����P�%XBB�I�/��7GB�X���Uh_�3 |B�I��m�2-ۈz`H��Aʎg�0��d�<�O��e�D���Ub��"Ӫ�q"OB�˶*?� �['����i�"O�r#Q蜄�1�_�9���"O�"C�L8��`�8���y"OZ5*t��
�h3��?ﲔ�C"O x��K/΄I䀀>Z:��9"O2Up ���x|r�+K'rf� �E�|R�'.b�'��O���<J��湊6�*����B�4P�	�'�:x���1wO�p��ʊ!ON��C	�'*�"3��n���[�OF�K��p	�'�pD�)>�<E�CP�(L��'ָTx���$���*M��d�r�'("`M&qb���g��nL�'le�A�ʅ0e�؇�ܞx��S��?Y����OJ�S�'��x��!�4A�^xa�!��E)��	�'ڲ���쓊5t]�S�C�EI�'Vf��Ej	#}Lh�n��?V�@B�'�̝��ؼ��a�*=�2H@�'@��i��χ#���%���5�$���'�T��ԍ�w��M�+K�3��"Ov�Q%*  �xP�7B>Vn�H��D&�S�I�=�֌����5o��h�ԩ3�!���!Op(�Mx%.�&ɋ�B�!�dHR |�G 
6$����Y?3�!�$�7f݆a���U���"H�^!򤝖o�h�2'��[����i.cA!�u�mi��JN��\��
cC!�$�O���QW�wh�pZ�@Ɲt5ўX���e��<	t˒�D�h��'K_>�|B�I�,#hH�7�Ù,��U"��DB�I�Rw8�#�|r�_)O:4B�	J�0�;BbJ)�P�v ���2B�I*��u��C#�)�\>(�4C�I�{V���	W�r����L#9,C�I9H���V$�K��(I��O�d|6�?щ�IS+: z��O?D��H&f�j�!�D��5k���(��eƕ"�!�E�H8p`A���aŠJ�H9�C�;y��׭��_ ��
�BC�%aG�#�-G�f���#��-�fC�ɦ"�H<���[�� TC�I6o�p�UG�
�D��w�I�T�?��� ��W%B:A h�3��ݱyL�YAD"O�1�č,�V������3D��"OЅ`��ЕM�F-��@M=!����"Opl�C��ڲw>�!���7D�k�B9g���+��b��7D����gGK�[��l��P��7D�L�Df�(�J�٥�H�@E�x�v3D�tKפ��:�SB�k�t�"	6D�<db��A��݉Uk����(��g!D��b�K���|aJ�q�r���"D��Yj��GL�%A��B�!D����=jv��a'���l�`�S�2D����]<}�⸂�dƤFJ�g�-D��cPGC =� �0���.cd \��9D���C��9�����Y9���c �8D�`���+W���&B_���ɲi5D���P���ZyI�
ԇ{��1!�@>�Ȉ�n����VWz<܂s����u�0"Ox�?Cv-��Q�L��Q���y)˘��	0�
�	����gN�#�y�HV-;�r庥��Ut�e[��O�y"j��N��W���i�y�W!-�yB��`��Ly@FU!S�q�'��y�	�\"��EL>~�ά�6b�9��'���O
��D#Ҙb��8'���BP����yRjjcuyq��&fld�qЊ��yBh�>T�<����]f�!�d����y"���v8�9ӎA�Z)���g΢�y�.�UH9cS6{8�LK�F7�yb�Sd( ���y����Dm��yr[��pe���m~�Dh�&����?)���dL܄M��J�h߼[��K���?Y�'����U�)`�ɹ���.��-*�'0B�@�fAg�C��
���'nf ��V���1AdÇ �t��'ֲ�s�4g��	�3�C%O��Q��'2D	0DŖW 40A#����Y��'ͨ���Y	M!ތ��ˏS���+H>����?açQg�	��A���fȨ���E�L���I~"d�)9�\)c�%ʁ_J:m�C�D��y���'L�:���=Y�`i��$���yҧҸk �� s
��`d�!H&C���y�C��v�R�H�`���`���y��. !,���I��/�8qеJ���yboϣh�zA+�-�D4�u� ��d ��|b�y��L*�1���\�}1�yb�;)^M��`^]l(�x�����yB�I�X�S���bM��+=�y��� ��X7�f��TQ&���y���a�$P%g۫g��x2v#P��y��r�i#$Ğp�[FJqI�ȓɔT2��C�y�f��O�D����}�$d��)Ȧn�5
 �>�
��9�ecK�%oYp���J�8aC,|�ȓv��bs � I��]�d��"4��ȓqe�%����8wT8Q!�"B=FeP�ȓ���"��Y2R	!��t�]�ȓ@
��F�RKF���%R�m�h�ȓwD��{�^'8�� [V%��6r-��Y �y�ʴ��#rE {f��ȓ���e���A�4��Տ��̄�I�֩ڵ 5��9Bd�\�0��	�ȓNӂك��:V?�hZ�ϕ�DT��[�|��#Q*�i�MǘQ�*���S�? ��"�'D�@���BL�X�a"O�����6zW�Ȫ��޼D�N���"O6���ε%�u��kQ��N�!�"O�Qi ƕ5@�� �EQ$+��ٙ�"O���ÍH&qA(�U'�B�`pq�"O&9�$��w6c��F+��'"Old�%e "�9Q�qS"Op���g����$� �5�"O a��H���3�T�P$bq"OB���M�R��M
GZ�|�b `�"O��	�����,As�D�I5�"O���N+��#T�_�e��<��"Ov�{F�2"l6�;B)C�k�*m�T"O޴Ƞ�J�>ȕ@B*��D��#s"O��CP]:� 	��(�I�HI�"ON`!�ߊS��*���=�H��R"O��ŏ�;z��I$@��XӺ�
"O������/ +���0�$����"O�%���T7y�����fRfn~4��"O>�ʠEO��
�BƳC! a"O�8#'QbN9�jܡ!Ŵ��"O&�t����V��ɳ�"O:3�b=9��(��.B(vy�Ԫ��	ϟt�'�1��tF�q���c��BQjPHCt"Oĸ�'�/l��EDH���"O�QsS�
 ��eÃY�D���"O�P��2z��usT��B�j�"O��� ��E7@���3� 5��"O\���
$Gc�xb�Ԧ�
�P"OT�q��$��0� ]�
��ȵ�'���+�Տe2����	��1d�%9��$�O���B���IP�$S���$4W B�I�tW�1�'6�j�'F�
B�"B9'�
���7�[�O7�C�I�R��ĉg�/T~�%A�AFxXC�I�9��dZUf�'��1�����>��C�ɹ*����t�\�=10����Q�zB�	WR��ضM�N%"�i���#H�B��Dl�l������YWϠe[~�K3�'D�pQ���p9���L=}NL	f%:<O�"<q ����'�=g��MR�� [�<�B&��{��q!b�_���r�j�U�<��nY
��0CAM���@���y��V	,������4��T�"3�?����h����%��B�R/_�b�j&$�?4�}����a,��#�\��d�N"���C/D�$j�*�?�} �o
.�m8��2D�k�`�^�̨+YD��)Ƅ#D�h���֜ua4�Z��pI��;D��F�0x.^m����YY�U�d�8D���/_mj8&�	%��q��<YH>Q���O$��D�b (�'�An|����'R�I :���I"O�aG�m2EA�2EC�ɺ@x��������v� 2�?a����#;�H}Qg&$�i����I�!�䞨w��*'�<y�,L�Ҋ�q!�D�t��$�fc�9��ثA@�y4!��0��n�u��<���Μf�"�'/�'+�>���l�����W2r�\��@O�t�0B��Eh��5��I�)���:�*B�	�K��b� � 9�"${r.
�btz��8�I��G{2@ѓ.D��G�h�(�ZW�B:!�D�VG�,�G��$���� �-!�d��Q�����,xpnH3Chȅ�!�� �e��L�FҤ	�+�� Ja"O`�@��C�$���r���}�$i0#"O�qya��MR24k삠�(���'z��'N�ɱp�b����H߇T�#��',axb-��W�}�D�]�V�x���Z��y�����e;���P,d��g�ǭ�y���z^d��� ٿOZ����	D��y�lQ�!��b�K��5�j�a4��!�y2��[9�3�W��PTsc�+�y�Ѿ�s'�Q
�Ε�!����2�O���bQ�t�f�0��<(��Sc"O�C�i�!�h `Uм`�>�4"O��X�f�=�
$�0���	r�!HE"O���J�v�4rd�kLԺ%"O2�9��?�"͓"��Se�T�"Oxe'ǋ^�n���S/XyA�"OJi��&��T�f�t
��K"l@�X�D��	�8��B����x���qs�A�4�C�h|��� g���x�Ã�$C䉼qI�P����喍��CƶG|�B���YcGIP
�fq�5A��B�	"h���Em_�3�(�Z/�)�C�Y-���f��:8 c��-�vC�	2�(݂f*X5/�Ӆ��n�2B�ɎZ�h!c�:Mb�$+b�2"B�I ���+��ݾ��ISu�d�B�I�{IZ$1�&o]��{����C�%9���V�F��e�`"� \�zC�|�X Ggj�N5��۫+�PC�ɒP��C&��5�2M��Y��B�I���Y*�Ʌ�欣�?A�<B䉆c[x�e-���s6�¤	<B��6����G����C�E��tJC�	�#Gi'jbx�KEᐐ!e.C��	)V�XFX�Q��i�Ȑ�`,C��^�h@q�I!;�¬#W!ٴ}�C�I�>Nl	�`�4����LH��yb��#�.=A�$%{r�,��Cގ�y2���v��*m�>���ز�yr��WZ�A�b��3��(�0O�9�y�ŏ1-8j܊QȀ�Ɛ�5�א�yr%�T���K�h�՘d�Ϝ�y"�G�H� ���`+2�z�M�'�y�#��P[���F������"D����,PK4��q�qU�y��	�0(��h�-�&lxQ�N;�yRd�	#�9!�F.1RDp��5�y�II����j�n�'�e�p�˙�y�\�i�q�Ug֯z��X`�A��y�
�3{�iq�H�<	v�QcN���y��O��z)#>Tx]�rL�6�yB�Ha��݁5
�N����
��ybl~�8|�䌝�?C��	ՀE1�y�T�X\FՋc�PE�4�d����y���\G�@yu�?DL]����y�Jt��� ��.1�������ybnZ ]C�l;�Ӫ�΅:�.9�y��ΠQ��yw)�}�&���yraܙ%����c5���F��0�y"�ʌv�B�Kq����^i��ۍ�y�LQ����+Z�W�j=#�n+�y�B'OP"���m� WP�p5H-�y�B�q���E�pTX0��y"΋:Yj�D�Pl�(<����*��y
� �lz���/䀢�ŉ�T*"O�12�C&o�`��`c� w��YBT"O�4R�T�Z��uxw�ތth��&"O�x��]=Ib����֐����e�<����	5�a�e���Y(����y�<9��)+6�xa0%��k
J���c�l�<�F"(h��5� ���x5v���$i�<�@d��H��ܑF'�"�#։�M�<�[+0�4PBခƀpsEƖH�<�P`Ls�����ʢ�l�{ �D�<A��G)�%�AB��F��"�A�<Ѡ-C8U@y�q�ɾO�r !hM{�<���1��pa&Ȁ�1Й굋m�<�v�O*GV�;q��0r�
 ��M�<��?t0-����K��m�+W�<q��.- d��hȩ9��@��B�<!�A�>3���KA��jn��zpk��<�`�a5���W�ݧ"~�ҦD�|�<�Z$~:.���s&YBծ|�<Q��4�xe-N�
�|͢eLC�<�a@2�u�$ꍀg�,TzwB}�<��oB�:��Qi%-k�pb�Ey�<��U5!�d���S�{��i�C|�<��B� b9��Ν�At��F�^�<�4�@2V\��"Ӝa!Lh� g�E�<Ih2����G=�!6��D�<�5�R�A8��{���<N���PP��B�<��EB�A�7aҴY�^U�<�%�(%@��Hs.A63�>�H5�CP�<��>8'�� ��&t{ �H�L�<��a�NkH��h�"u�>�s��OE�<�Q��'vb���l�"	2ܓ��e�<)�� �?q���(A�րYa�[�<�`l��(ؾ5\4\Bth�Y�<1��K���RB�T�>�+���A�<�E��v��Qa.S5h�@H���]@�<I���1岬k�n5!
�|b4��~�<A5k�>nE�e��R1f��(:�~�<��-m�����F��-l�c�%u�<d@���r�C��TB�r��l�<q	�-oR:�A�酿c����@�e�<q�)�xFJ4R�� ��������`�<9Ԉ���	`P��F&��ֈ�E�<!#��$Q＄�c)��<� �h	@�<�rD��&#����;Ș���a�<q�A�L60PS⍞8��1��M�T�<�.�	�9 B/�;�ݫ�)�i�<��B�1�� � ��%"�+d�J�<�'c����2 �P,E��Y� ��]�<�V��(�e9 �ϼY��r�<���݃U攠#�KK�\��b���w�<qv��3^�\a�T��>�v� c��<)2O[�{�
abFďtr2��`Lt�<I��T/D�|��F�D�
�@�&�Y�<���"���H!k��U"�遅W�<�T�L ���ll��EלYlA�ȓ%ff�0�ߡ#��uq&�ʢh{�����(it��y�ެ:�ܵQ���ȓho慡"�"��� ��/?�����N�d�X���"����!�\���I����ւK��mK"�#VX�ȓPR����.��{��k��٠R�5�ȓ%���J��$%R��
�L�`�ȓW^(p�ѿel�ч���xP��S�? �@�iWrE���Ҝ1���`"O���O�4�xqC��L�HX"OV�����\x̹#Q�ܧ3�E��"O���f�#Z,�Р%�'�>�0q"OFB"/�5^�d�h�F�!z��E�""O����A8Jt�X��%�)|���x�"Oz����vZ,jQ�������"O����$J�2< ���V��"O�C"j�@�vQ���J0\a`"Oz�q��5}��!q��BA4Dc"O�0�(����i�ЍN�2F�s�"O�X�El���5fJ�'<�0"O
�8��H�^r�y�B�s)��'"O.�P�惙_���z�а��W"O���L(>p �B�%�|Ը�"O҄��/˘u2El1�䤀�"O �:�D+jԬ���d�� @�"O6I	�Ș]t\��$�łe�����"O��؄�Ѐb⦠K�CF;����"Oz�3D�D�)������"�x��t"O|��g���j�.�CU!T�`�"O�L)aAԸq��)�B_��(h"Oh`s��	*ot�09�O���Q��"OȀ8����1�fDa[�E�l�n"D�0��矄&��L:2A�`n�ͨ��8D�x��
Q�)��e��E䪕�D�5D�	Q�� �p�;p��	���x5O D�B�a;(�(�c�I$}JX�u�#D���E�(|D�c���C;2l�!D��ʗ��;9=d�@lA-P8P��>D� S�H۴_:�:�+��Uv���B-;D�Ȑ�N��L,�&��><��dm-T�����:$h�r�,O#2�dp4"OR�X�UF+ @���[�*B�Q؀"Oʴ����%gj��,A>���*O*aࢃ�ot�<[CG1n�%i
�'NJ��EOw�颓��\j�d
�'qb�{�������G��
�'�N�H�ʞ���X�BI:���Q�'�����i[�9��膋ƫV�Ex�'����!���s���2��#I h9	�'�:`HsbHɀ(	 nԕ?:����'*"�b���:s�h��º;vQJ�'`��X�,��2q�I�%ۈ��'�}�F+��C@\�k�@Z5#<�x�'�����mA��-�g�K�J�<x�'�2����������g˙L�Z�'��A �=\+D�Pf&�&	�Zx@�'������Gt\9v�	�|����'n1K eh~ĸ%1r	:�"�'�n�h� ϛn��H���k�4��''���tC_ 6���p� ܾgI�DS�'��as�C=:زlP�@	L\��
�'}椋Q-]��v@!�e��L�}�'(d@�.��t�ҡ!�d��K��}�'�BU��O�QmX����A�1	(ِ�'���Y���]�$��]��'�V�Ӯ�v�h� ��^4��e\���<����*H��� ���L���i�&G��}���������@��A��I+^ك�7D�HCD�\9kT�T&иul"I�i3}R�)��9v�LIq� �qWH��f��c�؄�I\�����q�ӥE�F�����a?)��P1��1�D
iC�W]�<� ��E�?W��R'��\0�!t�'>ў4�n3Wтl��N$5 ���!D�<��E�=z�t���b��I��"D��j�&B��ܨA�%%fN�x�G>�OP˓���1��_i���!��Q."(�'>R�'�x�(���*R����P���;���y�>�`�3$ -�D��?�y"퉲Dr��ᗉ	�(y�@��.���OD#~s��	#*�ؑ��,"�����D�<��eV#F�Q4g��f�+ph�}�<af�U fB�<۵�C"]�n�EX� �O>��Q�
o�Q�whۗ��݈[���� S�2e�����HP��I2���5���<�;�(�2u�$�I�e�`��&�-q85���:D�$"a��[\�E�a	�6@�8�9"�"D���@[�5��1��Y�\�ڡ��H D���gNY^����?�~T���3D�ԨQƁ#`����ޱ@�L|���0D���*W)H��)��
ۗ# ` �7
,D���ƙ.
�zE ��\��'+)D�\s�n�1g���t�V�
��*�"'D�����C� �l3C*�2 �:ykP�$��hO�S]�:�k1e�\-�8�ƊP�kb������`��J��\v�6� A-C|C"�n�ş(�?E��4q����7/�)a�����?�LFz��~�b�;mQ�Di�D�<H�
ف6�[?!P�O:��dOC��n�Ix��[E(5P��r��1O\��?���JA��P�%br��⤗pH<I$LV2?,(	�mB>� !J>.��	h��,��+����x��.&�S�A6LO�⟬z&�D�K���pL�Ȝ�S�N�>)�>ъ��wn�q� ���2[Q~���[j��&%^Ni�!�@���s��p�>�ۓ�����+��s��9K���,[�B�I'R�6�!4���{�\Q ���6Y�C�	?/����bED���$��eɘ�DUz���I$�I�n��E���4(�$��"^3�bB�I,$��I��ȞZ�K'��ŰS���4�L	Qr,@.��c�Ƚ8;f8��N?I���ϙU���� E�a��-�&�)���<)�d��NْC�L�I�.L� �d�''@8Fy�Q���F4�D$�7"�6����bO>��xB�. ]��ᇌ�S%��VA�$D��o�P��h��q����T
�+4D
=b� ��'�qO�"�O>�"�'��fȅ�t"O�Pc�	ͬ|׌ԁd�)~d���&�>ъ��)�	<����s#�'.��{���fF!�D�A5��5�Ȁuwe�592���)���`vn�*T`JD�L�~�p0/9D��`��_H��;��ؙ|�@���!x� �?1�ט'Z�S4K�:���@&�Z��ML2#���m�H&��ib�́53Xg��h#��!�v�8	1H�S�O����SnS%,��rO0uf.��'k<C�Ϲ��P� U,q�ZTA�'����Ȅ�V�Jm#�B�<��1�'�s��6�P)��A�
#|uy�'�����	 0uL
q�-o�{�����&eT-Oc4x�f	r ��#��y2荿~_nT�#%[oD���&����<�OR�Ђ�*I�����m�3.8D�(��	D���	K�1[��'�+�6ذvCN\$!�����+�C���� �0bA�1�k��ħ��I�"xRa`ff�;_�썀3'��Ɠ5*r�j� fPfru��Vٖ��	�<�5�)�~�H?��S�? h�ℏǣ\ŠMC7�C���S�'��̧>iCH�h��$�T�R� ћ�l�[y�'�Jy���'��5*膤XJ`�CU@�)b|����D#��?��ɷ1�rϒ`�$��S@�; )�U��!8���s�Ж*a\X���y��C� I�#N�E��ܐRLL���M�g�Z5���?NIt�Y�!Ewar�O�q�g���̦��Q��j���'ԛ���{���U`ި Y�yA�g�,sK�B�I"1��tS�&�)a�z8 ����G���<E��B2	 @L��ѱ`EN�T��y2�>x��sLŖ_��I`�lÌ��'�$܅�I<#�n}�fi�'	L%��e�5|ߐC�-)�H|ˇ���`�`���^%A�NC��uV�}'��9iE�� �Z�RC䉃B�ja��۝'��*v#�
yvC��3k�^tz�T+D��x2�LK���⟬E{J?����o�B�+k��^�(���:D�� d�!"�jLAS�R�J�X�{Q#7D�������J*`t ���t�v�	�A6D���U���x�TykR*�oF�tm(D�04E~�U����9XM�%D��@�e��Fpd3�eݣ{��l���"D�T��E#p��� �'r����,�$��1z�%�$��}0�Y�A�=H���p?!��܄mD��[�F%Rݓ�
y�<AA ��`� ��2k_R`��I�<9I��h�݃��	�@��(*���o�<�g 'i��xjgk�
{\z��Jk�<����(>��SSÔ��ZÔ@�<	Ď̂qp�أLN��X��c����?����:%T�a;��E�}}��3�O�X�<a�B�'6�L��gG<l����`̓ט'�0�|�JH�f�PdIp懸F��]9�/IY<��85�a�Q�p܀3cPD���'�ў"|*��-,AD��KF�΍0E��v��D{��� o������:�KebK���'���$�&
I\x��BMD�9�&O�GR!�4���2�*G*>�	i�M��!o!��ڶI7l��%�+g�RD��ƛ5���gy��'� �ca!���\��BL�4�
�'��d�`�ͪ�t|Yʈ)t�p�b��$<�S��b���&��Htb8 �jɛ�y"��]�@����%,�q���mZ�Q�Q�"~n�$2. I��ژ!�4���H�P��B�I*�v�jA�Z�rrE/��.�B�!�T��N��&��YS��h���	v؟�k�%�;9B�]��-��kM��#5D���1w��үO�=9�'�J�<��.�
"�9��K^j	.��#ꓢ蟂�3�@�$v����$9�(;�"O�l؅���.%.(z�OD�+�aЇ"ORT��oÞS;�uZP��fQ�"O� �[�v�`��P�Åh�au"Ox�Z�)ǈ{��K�%*�@}J"O���P��	4�H*����^`A�"O��GLΟAJa�s	; �h�"O�ț'30PTH%ŏy�nppE"O �qf �z,Ȅ��m_�N� �;�"O`\#�#X\4(P�ވ(b���"OR���������wϞ-T��"O�P�T�*8��i���8�<���"O�1Ɂ�7k�vd�qDH#h6bUc�"O�T�q,V���-�Y�
� �"O� �Q����4X�HJt��"3r0���"O0�pqBD�D2E�sѱII\�
�"O�L GlL�Y��M����RJ7"O��`�śH��Г�+�:^$��"O����Z�0�٠�, �2�"O��s���d� 0���(�n��"OmS�Z�&z:Uб��\~�\R�"OL���ώ�k�6	�ݳjl8��"O`�x5Ș'd��"dH�N��s�"O� K�G��d�"�� �k�V\@�"Oh��AN^��y8)^-1�<i��"O�A�a
�$��
"G��\�\H�"O�Y�W���]L	���U��P�"O�Q�EW|�P���!8,Y±"Ol:s��2_��d��I�%}���"O�Hb%*�>����e,z�x��"O�օ�Aײ�� ["l��p�"O�<���7Lr�m�`�,	�"�`�"O�	A	������Ώ�ʆ��`"Ot����DZf��\1���"O���uk�m�F���<d�p��4"O�E{�%F�Y�e��.C�f�(Ɂ"O H�#R�_u�d���ƉC�V`3�"O
���A'+���Y3$^H0��"O���gJ. ����~��Y�"O�L�"e�X��Q��F�-5bΔH�"Ozm��)VT�bd�3�W�Z	�p�"O ��Aǋ��4X�m��E�  *!"O�ya�/5$�p��6%��i����"O�=�`H�6ލ��ж�`�"O�I!`��5yC0$���Z�2���"O��b�S�)F=��I����9�"Ozi����S�ڕ*0j��A��Ը7"O� R¯ײU0��ɧI�E��tV"O��	001@�0���"2�X�"O>���Y�+�2� ��=g�T�"O�]���T6~l䱁�ѕ*{~(��"O� DȢ3fA Ӎ��`��!�"O4���D<Hf�a̙{�rܙ�"O8I�!͈�c�f���i��t�$)I�"O���c��_�����G�2p��"O&�s�B$_��=A��:X�ƕ0�"O�l�1"A�RXÀKL�[��|qu"O�4��I 4E2z��'I�����"Ot9Xc�T�s�,�y��6$�*���"O����/I�z�Icg��$���0""O���Ǚ�3 ���Gm!3*5D��;��l#��3W��v2��t�Nm�<�"M�A�"�QQ"PM����c�w�<��J"f��e�Ň�"4��x2�	Y�<�`C�8�J��U�E8�| "�c�V�<I��R�qf��IG?Pxyn_P�<�ևp�Lڦ�;?�B@[��N�<Yw.&bǘ��G��81'�L� j�R�<1�eD�GcX��%I0M)x�����A�<1((�~�S蛲�Z���&C�<9�$DOǠ*5aγ+�~a�''{�<鐏ߗa5nА��)�H��g��J�<Y�H�|,Lp$`�{�2�Q��\n�<u̖�3yl��т��T�1�G�<!��DNl�i�R��\|�<Ac�2|C�E%�	�ڨIIwL�}�<a�i �E��r�]�	i�U��";T�����Ԟ�&�q0k%c�ˤ�u��I1,B�qO?� t�9�aH:�d('��
޶��P"O�q�H�;l֌@��lJ�Q��X �Q�\#B%3+BY��Ʉg<p9@�գh�Q���P��N��$!@ȁ��,��!A��"7�s�Ԋ0���u
�'�mq�)_�y���k�͇8<�J�+���_�u�����Խ��OvĔ�K	"����s��3�����'O������9���F�� "U,���4:��B����lӧ�����UDX�z�	u�D����p<qQj]'��'#Mi$iJ�7�f�h5��\=X�OީI�ㄨ/����
ϓg�Dj�˂D�i�ᇏ�z�'�����CO�S��c��r��h�������n���x�"�=n��7H@h<��	L�q�����Y.�( !�B�W̓�<,q�b��ؘx�k�*��IN���۴H!�Qr�dH�hݤd����D<���x����ϨEMv�"w���Y�����iO�:$�:t��/��I^��M�p+ҭ���rƯ'�xy:ed������}�qO���/VU\�!���C.���c_�����4 R��'"e:�ΈO���AM��~ (�Ofe)PfÛ鸧�	ڎ|9[p�S�RO��`�*�2Mӄ�9��ʄBoRT �'&j��� O�������'j��0D�P㡎 N����5
Qt*P��p�g}�O�fI@�ƅQ-r�8cC�Lp�˓	�R��!fB�D+"�\"��$�۸D�� �R��RJ�ϓN���kĨ-�)�'$��YS �
Z�4l�J�qM���Oa�b�U��D{��;�c����#�����p�O$�3R��,�0=����T�upR�Դ!�����O&g�yiP�x�B$�;�q��N�L3������#_Z���-a����$�Ԋ�Px�@\��` �H� �X���n��<��i� �(!Ҝ|��@��8�=�S$FFykD�$���KEI�7����-+��7���2��_�ZT�Q!��5�L�#�N�.��)�θ�!�����S�O�Z�"rQ�`p�8Q���-In"�
I��YҬ
]��t�eB�k�OZ�]�W�C�p��܂�m˝Bd{L���u%9��8Ǔ2B��H5��E�
��SM�K=�lx�dڋV���5GT<٨2��l(�g}BaLn.�J�	��80�$ՁH^���됯%^���ɯ$	N1���s�0��4g��X�G`���t�䓻�ē�Mki֑K�6��D��z}���5{�B�+_2\��a����L2�p��	�e�h�Do�(��DO"S�@��%l�|����!e��O�1Mo�\¦��(5!v�	A"Ц�~RF�7`9\�Y���	���c�4q �W���S�ȁ�g~�O��C��	e|�	f�}YK�;&����&!a�:yh��	+D�a�D�I:I�e�IOw�����I�y��h�Hp2�S��ɪ��};�옮�P 2�)L?s�c�\�{q(�'23��Qt*�7{ڀc�����N�P!��C�+�8L�h]����(�)�F�"a�:��t,Vu���1Ï#y[L�S��M�N��,��쎳9��%Թ&Uƈ���H�<���q�!|QX�3�N�����|0��38�@fF�)RK��H��'	�``r�Z1 �(1���`͚���B�,�%S��S�v�Tc�L�/>(��%�� x���eʐȂC���TmD���x�A� �J(u��'���O�BEƎ�X �$��r�E3!�X���0�%�M
xs��ڑE��m��o�>!p@ۂNў�tl���$�n�,�����$�.Y�h��<���ޑ~�|I2�"PH�2��Kƥ(���O�q�!ݝ@N���/_ *�>���Oil��1� ;�a~���!��!��;����U��;_s��A��0�F�5�>=8�[?%��Ϟ8����O.�X��"MT�A�hD�[N�p�C�'�*�hr旇A�:��raĹl��X�pe(Tk.H��v��2�E�=�P�5���+]�E��k�Q�2�[�|yaxboZ�kZ<@Ҧ�v ޟ]�6�Q>?�B����@>Z�YV+Z��yRJޡRm&i$ğ;��e0p��1��$Ȉ>tZ=�P@�
f�R�k$
Md�O2\4���]s���9����r�� �'(�Q�%���]�������a��lyע�']� �㵨���1�Jȗ��g�O�<�aᏠ����'ʨ2����I g�:��Ab�V� �Щe0mXQ	̖�p�ɕU=�� �SF؞hR�M�Z."�Q��׿kNɻG�;�ش����F�t�f�~��yBYw6��t��9bJ�`����7���+�'�h�؀��B!8e �.�*�Y��'ٸm
DB��b`��Z�f���;ҧ'*Q(���Q�H��e�e��N���bÂH�� �?-\���O� )3$�رd�(3͠s�j���D��f)QԊܓL���'�N�:��}2�?8�Z�!V  2sh+2oG���kp��+B�<y��4!�,`��TH����7���� �x�}0AK�}ў�)AB�15H�� ��u�\��˃�'�� 4ږ#�"�"��'׽�<+QL�cH<9��� _>}B�x�2}�l���E�%.�����d�v��E�U(U#�;��Q�R��c���=�!M<+L���'�b�[քD؞$����AH�iZ�iC�E�� ".yX�h�����_�V*��'Dh��.[~�P� � �
H�������w|�����"�Rap�"�ZuH#J/D�܊F N4.϶I�Ն��i���Õċ�n�dۢ�[Xf���/��^O��҆��6��	>����S>Y�x ��� M՞�y��I��hO�%�ďV��R�$�7#l��BbX�L�z�h��.]HQ�&M0YI"�#҃Zd�<ɂ%D�k�0�'ʰ#}���rb昪� �r&>��CG&]��D){\%a��T2`@�5 �-qh�`�q%1��$�'탕{���m=Q���������@ݽn��j�'˴@�$��O�y�
�7 ��2���K��AȔa_71��T���΃��Ƀ?meZU��� Y�u���bMV�����-\U�T0� NIa~B��&�	+R�ɼ4�6�1�&��Y�����C������A"lY��05�pɽ6�4�I�h�OE0u�4gX-~����8v����$�Mw����MQ0o7���Pg�~�s�Y&K�ɠA�Y+co"�S�+�?e�� $Ҕ��O?���|Ν�����,�R��1��-<��Č/��q9�"�Xd�Q�#%��� C�!�, �%ʀ�A�v%h����}9��чnp��$�E�i�e�fm���R��-*�epA��4cCg���fA�L|Γ)n٪©�EBy��G��Yeq�3b�a*�m"�O@q��g-d�`�r�|r�`���+?F���R�Ȇ�M����n�?9�lN�3�^�{�	_\������_�r":}�
�֙��G�OF|�v`�*u�d���ʲ��4���{�(j `�8�8�1���p>��D�*޽�$iT�%��񃦚�'�@=	�GC�t�2M
��I"b��?�� ���Hs��!�n'N��4�b"Oj�YD�� �`2�
�R �!�'vD�H���$7��P.� Hz�yd�����Â�V'Ҝ��[?��\�ȓ$�p�F)�2W�tm���ָ�v�4j��)[�ֵ�~�S!̗a���I0h@\7���y�@��ƚ64�8�F��q�S�'j��D�䌛�Tͮ@+���h���"bJ����Q��J5q�T����,�0>��3Ŏ��F���f��L ,e�`#�kV�p�Np��ƙ�?a�p�W�.�� �O�t}[�dY�@�A��5=t��Rߓ(Dq�3��>����� :���0H�I��f����j�ቢv����*�,f20���j�O��X!`��.���c�@G�օ���;8�%���ɀx*��@a�Լ5���g�M	#� t��b��N�� ~�ؐ �^>�Gx%U������o��Xs GWF	j��.�Ic�O�a@T�U�n �3�ϳ?�@9SGH�R�\X�@8B��(ӓH�s8�P����3A"yҢ�V�Dn��d��OL�	c��&��8�H�C��On�XT��9���&8���t�M��|CH3]!a|��C��l���jJ:f�{5��,&�؉��E� �G�`�!g�����#-�^H��yB��$�>;V�ٟ?����S@0X��MC�b$�0�>�wt�n��`	�Q�7��S}�y��#��LhuO���%��7U
�0Ђ��oe,��׭���ft[�-� (@��Ų'������k<���I/%��IF���.���o�$$��g�=@�]�Df�6&C�	�s����Ce��XX�MJF�E�0|�,���Q8�ЬKv�^�O���5�ѕ�jQ�Ю�0V:l0
�'� u�W�߈r���GL���|�a����� qG�<��'�gy2��[x�{����ju!jq��y��J�b��y0M3:��P�\�h���	��O�\#�#lO��A!�ԱX�z��Ƭ�<���'$�)��gξ!����i-ҽ:P���
�L��b�.*�����'���P�b�{���җ��,/�ő�{B(֖��T�GDċ��>]IGh�/Ip:��%Dq|��w�-D���$A� D�1r�K�8�pH���N�Q@ Z��l���DɩIG�M�r�H�i@:03�P��!������j]:�Q:ǧ�6b��
)!�����'3�X���޳f���뀈Þc���b�'�P�aG%G%3�Se�!	]М��'��A�A�j�5�Tm�rؖI#�'w� ��s`�Sd��#cj�'l�@�0�����A��0E#
�'�(FY%G��=+2�
�|���Q
�'�`�I���}M`�J�M�z�1)&D�� b`��ȉ(p�V����ߎ�h42�"O �����n�qo�H��y`@"O�DB�fǧ�T�)�.WA�Xis"O ���U��Jݓ��
~DI�"O^��:��лC�08���"ONb���10�r��5n���ab"O��y��!g�nd����z�
q"O<�)��X��L�W�G"r����"OT��g>#1&�{W�Fd�1�"O�I��nE�i�������=�A`�"O���@�W����3\���Qs"O��Bc�1n��0��
x�2�"Op�d�Y'/�p��N�*>�����"Od+��c#ߡCϨ�q�j]!�](4�`��pF��2� =���W]!��'Q�ȣkC-{��H�"D�!��M�,
|| ��O>�e���7�!�d��-�d�$HԛB!b�צX��!���^CJ��u+U4
�-�t�.Q�!�P7JD������a�ٌ^�!�d�r�I1�ح&���r�� 0)�!�$S�6ư��P�
(`��ip!�ޡ!�ټE~�!���	~ö��EG�`]!�䙺HwB�;%�M��ơ҈&k'!�dтV�b<h'$6y���� k!��ޯ��Yb��%s�M�K\�	�!��
.C�B�k�(��01B2�D9!��X�&-��!�������,�=?.!�D�>>��xᤈ$~����+P�t
!��>�k��X�S$ԂT̗�!�$	�"��\y`��s0J-���8$!���A�pH+1·$)�d	Q�X �!�M�0,���EnA�5a��MV�!�$��F$�I@Jj��CVfLz�!�Ā7�^E8F�|i�1��Le!�$R�#t��C�"����ac���q�!��JqZ����:�%�M#�!�DN��J��s��+s�f�s�,$~p!�䃂8���0r�q��5iJ�`f!��}���s3k9D0��8ǊT�!���F����vK)>�rt��&�!�D��<��<a� O��0	�LBT�!��2I�yg�<5��yh d�.|�!�E�JO�Uh��� i�V�[�!�D�n�"pCp�6qdV��q�b�!�
8� ��.�C���'(d�!�DR>Mcp��dk@�[:2$��g*�!򤅘Q�dMHC�z��0�+Q=:{��������$͙�Fr�Y��	���A0-2���8u�1H�V�&�P��u�!S֭ـ8M���ʀ`�@���QP����v$�􂇸{�����\��D�R6�A��,�(��ȓ>�@R8 |%�T��Q�$q��cg�M�4��� ;�)� CR���Ɇ�锡`�H�"�4W�[|X��"J�Z`A�0+%�R�i[+����ȓYi� �	@��ԎL�<�,��ȓ^Ԑ횇�͠�5��@G7Ype���ԝ�VjR��qk�!E�"nЅ�U����,R:x�2�ô�Ɔ"Q�M��4��-�U!�$.EV��O(����pI�F�Ͼ�(A�(I-���ȓ��Pa&)�$Y�!䄊*e�FH��S�? �E�*���i��էP���{�"O�r�b^�I���s���=T�4�;�"O���CS�����e��}�n�q�"O@�7؆���j�P�jhAz4O�e�1�L-Ƹ�������A��zy���V>P::!"Od;�V�+�6%�&-S*A����^������5N�T ��ɓ85B����� �f���E
���2 0@rƨk�zM*4�1L-��H�$���'��9�"���=��m� 7H�0��D��h�EA���O�4�Z�n7b���#"ƓyֈD��'( ��MM�8�X��,]Pn�xشbж�I�ǖ�?g�ӧ����dۆV�����2��YQ���y"$��Y�,�Z��A5a��s����d�#U�5[���
��<1VnG9�����A,�
�r�vX�xE�U<j���Ṅ29����E^jtEԇ�!Z�񄔚b�<��.o��c�*L�,���l!5
L2kv���	3t��Q����A���rS�L�V�!�$�)��xP/S5D��R�O�wɛF�W �U����@��s� ��P$�?�>��HɀG�,8D"O⍚7�T��͊�g^�V�t��W���l�&;�����'�f��᫁8cS@(��L��!7�H�	�Adp���V�u8�1Q��]�A�>-H� %:L`PQ3�>$���a!�$������ɝ,+�,����f�Yb�x�ɏl�q"�S�)��:��ɘ��A�tT,__^��DE�3�ɫPi�(����^���[����R Iy7�d�+����{�����(�蔊��Ȉu�~ŠQ�"M$����1C �G�B8���I<jZ���$E�X��R Q�!�$�dr<��@R�B��Ö́"⦩;!�GsyB�?1���}&�,�$h�!1mL4�T*�vz��V"9�`:D� �R�3��X4��� ���ZȄ�h��9V\�M��ɠ�H��� �
	8��A�Mƒ��$T�\�@@J�`�`2�
_J�
3$�	G�i�̈́H�q�' I��	T�S�O<�Rv�	Ad̬�PP�=�
��I��q���.w�%�u�G�O��{�C����&�
7Rj�qN<4�k����p��1j��F�()\�z@(��-�LQ�꟢d�剡*T���E��I?�.�N�[���왁BW�r4�9�#��� y��>�O�Qp@�Q�f�hA�ߏl5�[���� �D �.�W�O6m95Dxɧ�[@��I�
��t��)��q�p�c��ҷx4�r7�'�p�@�ě$m�ld�.0�-�"и�aFؘQRF��QK° ��9��(l��)U���&�	oR� s,�hⓅy������V�V3c�FZ �OT#C��X"��A�IU)�10nx��!ł��M�� �#z��H�<�4���
�5��y���A�  b2���'f� C~���q�B�6%�(O�	CR'����i�4d��<�kH~���<Ĉxp�\ g*�l5��Bm����ʂ��-H��/�O<H�b�P,C,����H%iN��K�&+��"AdB�9M�L�FĞ� �<@���.I8��	�oF��wZ�Ċv	XL�L�����wxQ�0_�����֗����W%��R_,Mx	�*cvUA��Z�z_tm)Ӈa����'�N��ҋ�(-��O�~]�W�_	2�aфG�R݆����|/Ќ$��+pP]K�fK��u��q� �@�E�C�. �d��9� �O�%��'��$>c��Xrc�6ˠ4(�A�\�9���<�F�P�
8�K�g՘#��0�-��Ij��g�I�`�u���y��`��P |���AQMV_��T�5�.J�@���j��r�h��GP]y\���O�3���4���O�D�Ҡ���p��~
��#�� %Ǻ9Y���ob���	{���Գ,�)IP�Q�dQ��F<"�B)۱Xr�X�)kqO.�N|rD���Ua0��+!�*���:O<�S%�=@����D��.n��lZ�%�,�y���8A2�OB�6��C�8R9���s�8<9/�w�0�'��yhRD޼"�Q2���E�>����1H����&s�ԉs�O4D����˜�N�t$�m�s�P���>��u���#��L��~R	O (���C�D�t&��q�g��y�)U1\&�'\�m��u�7��?ё���*}�]�&�<lO"��B��0.;&����but ��'�x9j��*W*�lZ�z�1#��;h�6��P �m|�B䉈}X6	1� )��ƯڔpBV�P�B����x"�S�Z�l35b����qb��C�)� N	q�V'.�~�QqJ�7{�.5VȔ�"ba�"�'��s��c&a��<��E(ϒ�G�\ ���$D�x��.��$�ӏ�7j"�ٶ��p��dI���q#.<O��z�EM�$+4hg������'j8���~�8��Hҵ`���L�G[��O���R�1&�&�2W�F�V�ЈO����d�#�(�"��Dc^0n���80�ذ
���� ����@c�.��
ۓn�p�v���*"���q	|�i�6O�A��eȔ�x	<}J|�@�$m��z���3��݈�Qg4�R��nB!�� �@p�`���?`����[5��*|����-a�` �e�N�~�'�f� ���GE�	?k����2ֈ���ٌnKV��:���	�Jv��)S�+Լ��1�ȜU��IA�>y���O��:�m�Ê�
��� ��AE��:Y��
��3Q"q�(p��aǬ(�|�I�J�O��r��ObQFkN1Pxh�ӓ�xA�e��K���@DHŠ�`a̓[C䌂ꋏG�Pҧ����~��E���\RV����a1�� �L `�L�0"Oj��+�l��)N�\�M�%�>yӏ��3 �t�p�ί_Nf���B#}Q?Ys�MT�W=dl(�E	8������"D� �f�/�����%A:�,B���zd�؂���J�Zҧ���ǺY��$9���P�uP�.
<�y�B� >��`��n��_>�p����~bFt���aǓf��K��=~Ozh3� ��	��t�R�;�O�����c��������Q���YE��'��EQ!m�<�3o�R�P8�m��X��I1P�/<�ri;�'�21����T�'��P�x����3)�
�J! W[>'�a~�m��H�@�+w��O��\X����H���0�"J�C��E���n\<��I�|�$��q��.45.!�"���w��=9����
�rB�+�I��H��F���to�W� ��F^D8�(3����y��
+��h8r�^2E�
��ף��?�Bʊ�&=�c�y5>Pq!K
�h�����Z7��!��p��M ��%D���vB��}�,ъ� �6d@��DF�:n+�P�G�R,K�X#�D�@a:�'�O����ݳ6m��X�;x~l�U�'|fѕ� (?�v\R!$ěh,�D����U�
�q>*�(�b�7&�S�aKH��Wȇ�R:(��J�hG{����%�QL������ӆ/��	�_&lP����b+^��h���!����^(��<sD\����6h��l*��s��D5z��AӶ͑���>-�#a���RR��n>�S"�Z�<q�g�V�X���W;]�XHkСtz�[U�U,a�v��5Hŵ�O����dMjzH���G!V" a O-�O� ��'i���8�XL "a���x���12 i�	E��p>����-hj���0�2U.�:Q�W�'ZВ�f�ϟ48s�ҮT�ӅJ�F9Ж��A7�I�gΎ�HvB�	���04
�uj�� ^5��{��A
�}E�d��<f��m�F�p�j� 7��
�y2 ?�0�����?e��!� �I��a�Sk
���>�p�d�`�W�NBt@��i�b�∇�q��l�����UaA�U��	g̎��>5ـk�a{r$R�>8$��'Ĥ}r�r��W��p=q��Y�HD�զא�M�VCD��	��s'F0��
f�<I -B��f��
f�Yx��N�2�"��2�F�Fr}����<"����J1sa���_r�!�$D=EY$�"���(�ҳ���V�+T��-G��'ft@F�,O$,��
.rb Iu�3'���#"O`���mZ�A���VlW�v��	�3�)޲U{�/�n�|��ɗG�|c�KY�,L8�XӅ[/l���dM5�\�v�$[7��U8-ƬXͦ�z�j��5wjB�	�[� ���ZNZ=�R��w�*�@9�@�@�Z E�W�O"T�si��{�������@��% �'�\�.4:��)�b��hP�5��j��^�xP�s�>a��>qB�}�H��CbO�x���E�m�<q�Ԁv�lD���7;�2�)C��x���.��}���)L�d�� �\�,�BL)���W�NC�IE7)�vk�i�*��㇨O~>C�ID��������T���i��G.(kC�)� ��JS�W)�PQK�Y�"O\yEC 2�<����@�[B"OZě�f��OT(NO�;��l(�"O�R����v�8�㵣��D�B��"O�x�@� M�B*����bD@��"O�� .�A	�!��{���!�*OlТ"�\<w��}Z���h�����'0�%�D�	G�D�04cBd! T2�'�DYp��
/F�d�+PȢ�)�'}p�;�o�6`#�|Cm�]���P�'������L�=i2�""�6�F9	�'�ɪ�"�YɄ�p,s�z��'|-X�
://�ѱ��Ĝ>cpez�'����I�5�����I��*S�4��'��1"A�,T
���1�G%]j�8�'X�)e�1����𭅇^_֝q�'hR�����<�`!��W�DM��'e����Cp�\�{�R�LU4��';t�j䫅�!�`�t�����'���9 e�K����ƛU8�'?�����شW�~p�UI!w�d;�'z8e��c��|��e��/;^t���'����e[�.H�e�SF�:ި	��'kJ��Q B�z��񭒄 ��,�'̒�4b�D�t����z��	�'K`m��Ϟ�V%��hG6"�<�'��q��� \�n���l�S����'�
��M&>��%���]�Ț
�'f#�ԧ&i8��"V�p����	�')<|+�#��b�@AL<$r"���7BB�*B��zO���F�9q[�X�ȓ,{��+��_�is��F�-m� ��bYJ���"Y7@Pj@ lG���ȓh��)	ʃo�ݓ��ttx}���̱�q�ͅE�IK�����ȓ]� �r��-~�d�w�Θ1V:���m�D�+Ui��.L���f�C�R��ȓk����eT�/ޖ�k� �4�:��ȓ!(ȂD��O�N�A�_#A�*���_���$�O�֬	�HR�(M��+:���'�0*���;eń����aN��B�7+7"���(L�?"n%�@J���ا�O��2�]7�v̛���c����'逼A�C�,-&ɧ��L���(u�)��
��r9�<)��>;����%�Pe9G'���X�((Ů���z\�S��-l�5 �R툜�O,܄ᓴxޢX#�"H#�0tzO�+\�DL���u��W�^��}rN|�K�)Hm&\�A)Y	t�j]T�A�	�t�hY	D�R��M0���M�K(�9[@��H�,;�f�.
�`�� ��@b F��6�tX���R
��W�G�R8ap��0�����p$xШ�œ6H�	 	{>�9�FM�^�����M�){��\���H#h� ���ݖ���M��<E�D�J��:U��
�$̞�)��
5�pq�좄B��OFT��Ӊ)3�HP��L6jR0�A�1j�Ƙ�"#τU��ʓ.Ū}�'G�ά�D���țg���7'ytΌZy2O�!~{ܘ S��4_?�1��@��%��y<0��#ƘO���OzdPG#&�)�SU(�i��m�r vă��Igw��o"����G'L'����T�:j�X)�^�!�d�<�PL�"A-�hKf�P��!���N�>����Z��0U'ݿ4l!�dޓu	VyfD+�4 pƟ�%h!��޺!����n C���P:R!���@���IaO�M0�����+8R!�D�653�M`�%�$~-p�`��~;!�$řu����o�� - p{�N+!�B�=C���n�|�������#"+!�� �`
)NM��M��H�%�Na�"Op9���U��}��[$`x��6"O.�3eAؗ>K�%Ju���zG�� "O��	؞����e�4n;�q"O$���Y
U��r�� ,��Yh�"O
�{��H���Q�M��V�"OH�r�/ '$��ɴi�6Y@�v"O�<锠� sPb=���o����"ON�c��$Sx�-�A"Q9���qa"O����Ċ�4��(Q O�y?���"Oz� %e�";��Ѳ�78 Q�"O�L�oa�̀i=�L#6b$\�!���0�6���H�(�y �]M�!�d��u��;$/A!F PD�<+�!�d��~�+��� 	����Dw@!�X�;Z墳��IPu��Ǚ�%!�D��Bܠ� �*�n��sl�A!�D Ft��kݐkB�A�&˂��!�d\�4\X2l�.`��3C�<s�!��+f��u��#�~�(��D�!�d^=Ƽ3f���B���#�^�/�!�dα��+���sâuq�I+�!�$��`z,����[�^��=Y!��)�!�����2+0�Ь��^�7S!�ďL͢iR����܁NI!�$�I��m,b���Ҩ�=	=!�Đ�k`P� �o�X�Ah�#M!�D�9(�����\�Xy��@X�M!��[�M "����\$4l�U�􅖒*1!�$G ��	��OȯBk��P�;$!�$ʷF\��*�K��#fqx��=!�d�Q�4c��.{Z�%afn�=$!��g�z�cq�E��|���͆�2!�D�4U�0yIUH=�H)�uc=r�!�d�0e�P���n�">�ҍ�hP;F�!��P�h�%F�G����eh\�Gq��$ʷW�茒����M�`O�6�y� N�?��$Ӈ�3D��!�ehO��yR��k<V4IRDǣ":�3u���y��B�,y+@�Ps
�P���!�g��VB�T���c�}!�d�1>�,���D�Y�� �Eˮ@!��Čt�I��	!�d���%�;!�䈐V���3IF�$|$��#Ε!�P�s�l��gY�*f9K ��7!�$�:���q�N�~��r�-�K�!�
K�MB�FR3q�N)�e,xd!��	cܸ�S`�2Z��(ru�οc!�DY.��x*c@�5!� �Y�,C0)K!��B<F%���"�ʙ�U���JE!�\�,��p��"9��4C���:y5!��ư�U��M_��D��a���Py 48"0hQ�LZ�~m`�T�yҨ�/u��I���OFx����yboD�?�F���H�&=�v�;PI��y"�E�I�l���"G:�LQ�����y2�H����Z5�?9���؅ �3�yb9
�8�)&DӬHL�a�C���y��ήW��M3� A�<��mM>�y�ўD�P�Ь45f<a1�]��y+0"���$�	�3mt9���8�y�'�n�!�9_+l耵�8�y$ڎ�xp:*
M� �ڤN��yb�PV?��kD� C�ڠ��	��y
� �q�&�8,T-qpl� R{����"O8q2�I�Z{�l��n��ɫ�"O`�hI��@�,�2艛w�"��"O��Rq��^
�t��D�Kk (`�"O�0�fd|(�)�I̢F���"On�Cщ�.���r�=fy�h�"O~H��h��b5$߄[e��i�"On�e ��I\�-��(	�,�F"O��r�%-RT�!��~D�q҄"O~�2�f_�?A����G҈Z�7"O.d�Ή'�\I�p�ϦN�A �"O�i����-��"�H��)LH��e"Ol-aw�P6_	�Yh�F *~Sr]��"O" �V�Z�p��T2 &9`�"On��삛t�����D�MuLMBq"O�`)𪅬]Q���/��L_�A "OT�X���Ze8�W�@�w�XX�"Oa!�gG�L�@9�� Y�(!�"O���*ʈr��C��L*�F��p"O�q������Ү����d"O�Y���n9jí�`Y�"O��J�C�*(��!�":ڎ��E"O`����R� ��p/ɐH�&��"O
��2��F¢�U��;�Ҕ�f"O�L*�
��g0��M�M���"O�����#c����c��b�5"O�� R	���&0����!����"O��:r�;p���1Q왉z�d�Q�"O���0�Ɠ.v��I�#��;U"O��3g�?�VA:"��.3����4"O\�UC��5-��cV�Z�ƨ�"O�S�✎U��P�مo�0��"OX)��'�86j0�"���9�d��"O���/])S���P�@��r$��"O�Hr�(�@����m�?KL�!"Ozq[6n���@Aw*��)и�!"OZV�Y�Z�� �B����"O:� ǋȡQR�Y ��X��"O��q��J�O0�@y�d���Y<�yR�v� �Td��{�Vy�5���y�F�3<��`ȎF������yB�u9���s��8�ir�g�0�y����?�M�͖4�ʩ 4G���y2"��YĒ�:�(O&)����T�ט�y�˥p��CB����~u�f`�9�y2��[��D��+ O��y��;�ybH��Ux&�S��n�x4���y�L���j�����0����(��yR'��Q�]ѣ�đ~yp1��gא�yb�Q"7��"鎤	�
Qx3����y���g��9�!"H .���Ac�y�"%>��q���1ɒpɡ�� �y2G�4;�%�dK݌(��k�:�y"@O=$<*ŋ%L�4�e,���yr�6	<��	���+0�8�#��;�yrMՈ,�u]/#��X-B9�y"%L�yv���Ch_�d٤͟�y��L7o8R`�!Cбe�z�4k���y,�N�|� ��>e�x�yC.�yr���c������g�I�C/\��yb�ǡN�rM�4'�R���5��(�y��N�����FFE��i�d���y�M@�
$	��d��Cv�E�T6�yR��(Xp��]*?h����+�y
� �˃*�&�e��(Q	Y��h "O�}�B��<{Ҫ�*�'	7�p�Z5"O"��o�1~���� HkʬC"O�]��ݝ\�"M{S�R�t]�� "Ot����j?xM�ʕ.3A|Q��"O��&j�"K��©[�K9�x��"O&EH��P?S��4H�B�&�^]�W"O,��m�5Pr"�
3AQ�\�F`!6"O�$�ƩsӠ��Ǡħ]f��	'"O|��T/3FƁ�C@�1&c���"O�a��ͧA	�ȶ&E����"Oj���H�(}�b��BRR�؂�"O����j6>z����Q.�v886"OĥE�9[����Z������"OB�!P�C�\�t̓����"�[g"O��
7�U�@⮨bP�L;l� +�"O9���ݳO����1�߄im,�u"O�����qڸr��
0l`�@�"O���`�ۚo^��J-ɛ �H���"O�|{��/����Vk��J���[V"O����僮�pA+�lh ��"O� ��菈GԸ��dʁ��F3�"O96�7RN�Z�	�E��|��"OFD�s�ιXݘ����H6�dP�"O�A�(��Jg|�JB��'늬{d"O5��	`����%���p`S�"O6ͺ�O73����l�}�B�X�"O$t��#�* �Q���!w���C"O&) �al@b G)u�P$z�"Ob��$,��N��Z�nS�\�D-t"Od�ć$!b��R�K4���"OL�����,M�"-
�h����"Op���Jߘ\7�k��ɴYZ@��"O@5Y�)�b�B [��*�j��"O��ʂ�ޞ[��pU�y�`:B"O�s�'�'��� �����@�"O<��t�\�0��\˕+L�
� �@�"Oj\*Wo��r��#@�?H�"O�5���`v>������`M���&"Oؘ��mǱS�$i�OD	Fn�v"O��ҮJ�2(5�.�)-"�Xe"O�ԑ��RA�JPx$��.��&"Ojar���q"C"��`0��b�"Ou�sF%���n�"5C��p"O��K���PzQ[Ƿ�N<x�
h�<y��.b�Z�y�,۶���S#�c�<R�O$R@DЀaM�ܰK���K�<��Ɔ�R��9:r�K�^�C�.�l�<��`��B>Y���M�6iTh�I�i�<䉖<@X�k�oPL�H�8��e�<�΅;_>&){筛�_x�`�K�d�<����E�ҐH�̈́89jUh6�
Y�<��S�&?�T@R.U����Cn�S�<	I��H��0! P�4�����e�<�-�0٣����ܳ���J�<�-�5>'0<���5xV���,m�<�B�]C���b-E�l�|ԓbC�<�D���ؚ�^V���HW�<1! �u$f����I&XB�#r��U�<���V$ @  ��     �  K  �  �+  �7  C  �N  6Y  �b  �l  �x  ��  ��  _�  ��  �  5�  w�  ʬ  9�  x�  ɿ  (�  k�  ��  ��  3�  ��  p�  �  ��  �
 w `  '/ c= +E jK �Q W  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�"Od�:f���r��K����\ �ďw���O��(D�L/`�4I��L�cxp(�'��%�%�OS��=��I�"Ԡ)��';�+2O˅C�~�3$�A�x�XP#�'x^-Ȃ-�-h?�<�����{,�Pݴ�PxR��JSnUC��P0T�0PY�MX�˰=!�,U_}b�'9r,���e}R�����=3��'w��ё�����ȴ�G�&i`���z�O5�}s2#̩<�&Y�v�^�F��|�
�'Q����PA����![�F�>4�)O�=E�$둦4X��'�S.R�:\�ïƯ�y��ճV�����i��OM��I�(�O���M@�n��@�O��k�k7���D�'u��="�a�tRf1���Q����Ɠg��h��"]�΁�&`n�%E�?Op�~W�����T 5�a�'OH�<9�D�;v�tY7��3L��0�AF?�7�)�'��24D�>[�&�t*��w�T��S��0�G�3;��A�-��N�4\��q���%�]�b�(�X0��<� ᱧ��W�p���!O�<��W,��D �L�x��J�#��e�ȓc��D�_(�ţ�1�����6a�6�v����P����Y��u{�iq�Y��ڐ�K�{؞���g�*8k$E
�1".H�R�d8�U��#�P8��eP��b���闄r\�i�ȓ��ұ�2�6��Ȍ? �d��ȓ?�tea�'U����$˷5�Ψ��t�ވ5gE>(j�xӧ�7>��q�ȓR�jV�;���"�2"�h ����ɀ��(B��l2t�F��-}(����_�i��,K��)b���d`V���\b0Ò�$�O���䑈~�0���^JI)t�$�a{��>��'	�a�p'�.Ѡ$:��	�,Z�`�'��� ��L�P�sSȋ�$?�e��{��'���(D�t�)���,�~hS�����y�&1JjUa�ώ,�1��	���y�#^�_&ɠ�/Ƙ=TTQ�H�)�y���w�t�0R�N!?p8�JRiԨLz��p>��H_�B�r(�3/�7�\����a��*�S�'�!���*d�Q㮄�j�1�ȓ`��t��	 C��Q�p%ڐU���>�J<���$T�Q	L�FF�5'�����
�!�$@l�(l�q�]D�DbA�zx��	u�jfx�xw�M�I(R� ��'MR�|�ȓx��=�2n�C(2n�,"B.�m�<��F�`�A�!�� ���!iX��Ey�#T�Dë�)e �S� �y���C�P\2(S�%n"���í�'5a{�E'L@8�"�kE�ƒ���l��yR�0O��t�Q]:�^�8A�#�yB�	 Y�Q��.	{~p	F"���yBϞ,Ā���H3zt4]��T��y�Н-A�t���y���,/Аx��rr���U�	�A�z�9@B�+RP�ȓ��S��DcX0 3m�vM,��-;I ���1V(� 0֯4�LU��0?��4�5�!����uQh/$��T��	��~��9O��I��Nv$l�5JϚ�p=��}�,����)q�VK3�yB�Q
2W������P����y2��7
�ip'�K#����M��)��� Ll8���2�X���ǷQ���
6"OV!;1�>]��Q(#-HT���(sT�L��ɛGB��UdH$IND�i*��9xB�I!%�2AyG!�"u0Ih���0B�	=9T�!iCLO��V� Sc�T+�C䉽_8��(7�)?����JO	2�`C�	;
�|����˾#�Xa��W�7��C�"s��)Jc� 7��`�/0��C�I69�@r/�?��ȫ7(Y.U,��=����N�D�rt��^ItIkb�3�Oi%��RGI5���R�W�/k@-�H/D�� �$��D���'B�<��9+n:�	�<����?�|�R({�t�ǉZ6 ��8���x�<�!�˴l�X���.N�����r�'6�yBJH<{��� a �\�d9��J��y���"�ctA�>����R"�y��]W�bܚć�=��
��1�yb �E^Ti����]7��y�GX�y2�]�[��NR�5�~�y N[�o(R�)�[���U����1B��
%z��
�'�SA��EJ;w~��&̥�Pk�fB��9/	��:oH�3z��`f�)��}~��5&�N���Ξ �J@�Q�؝�y�㓅]]X}��#�vA���8�y��'
h!) �{5�$�ǖ3/�>uX
Ǔ�M�ڴt����(*�Jր+�d8��ۇ\h���3D�T�AgڭnRb4��bO��0�Kѫ2�ItK���I�H�l�$�F� 4��>-x�f
O�b#�	�[\�Bb��z)�$b6"O�ɐ��Ȩ`y ܘ��ٔC�� �"O�P���12P`�	E@�P�"O@��'�#En���'O�0���"O|x�1!�!݊u�7����O#D�Ԫ�ÝR�P��%M�8F&h�`
#D�$��˨o:F0 ��߿L2P
ZA!�1Q	�k^�*�:�HĀQD!���*�@8�'	���$��"O|<U큫S0 ����I��;u"O��uJ�'Nb�	vm�~fh{"O��kd(K7mh�PS�]�Ih<�0"O*����γ,Bt���^�U���"O���*��}d�(B`m�T����t"O,x0�<B3f �s�_���E"Ov�z�c-z1д�&�U/Eu�y�"O0��$�%d�Pl�(c���"O�U1t�T�Aj���)��	h~���"O
�٧�=cP�`����/�.m�"O�����D��s��u��r�"Od�C�]HA-��%�rd��"O��b�FY��@��iJ�!���ɠ"OʼkgKK�X��M�30Q�s"O��a2⋆oH�����F�TZ"Ov ��=
�\!`A~�V8j`"Oz�h����z��]��Z%�a"Oax$�
�M8�
�.�\���r7"O�����F:mPm9P*e�&�b�"OR貇 �(�2���X-!&���"Ol��$�ͦi>d�*�K�3(F���"O4,���ӔG�<�C�J�A ���"O����39�	�eL��Ayp�"O�����r�:����,�=AC"O�@�2fȄZ�(�R,���@R�"O�Ag#�2_���U�ç>�X�S�"O kc
�k>�%�A��<Y/�@b�"O� �[4�ȷ3>�x@n˫=/Hh0E"Of�q��(�� ��ML�]%l�Ё"O��ppH�q�(�k�U���"O���oF "���
�e�s�(X�"O����kV�o}�P�"�؅f(�	��'���'A��'2�'��'w"�'��l+�JM�����E{�&L
���'�b�'�r�'��'���'P��Oj�����@�-hۀ9�@o2k��'%��'���'�2�'���'���WdzuCC���-J$x�HEaW��'?�'Er�'�R�'�r�'�G�="+\d!V�@�xJe��4kb�'Z�'���'��'���'sB�D�#u ���_]zQ��h�!�R�'"�'<�'n"�'���'o�L�1�"��!AK [��)zBk�+kr�'���'�R�'92�'R�';��܉?���C��7�x8"�(�aMr�'_r�'�r��4�?Q���?���fK~Չ�M=�
!Z���4_#|�����?����?���?1���?���?��>�)!�K���:�Cg� )���?����?Q��?���?����?�[u@��sfƾ8�	�X�}2����?a��?���?i���?����?��#b�͓$D�8+�@jeg	MK������?a��?����?A���?���?���1�fD:@�Gm7j��'W����?9���?Y��?���?	շin��'�*|���� D�TL#�M�S���<Y������0�4@\9#g YX0�� ׎J)A�P~�n����s���I#O�~��C����9�Fj�'w�4�	�L�q#�ۦ��'��Ʉ�?���(�6�Ҭ7h=����J|&-��$�O$˓�h���V���U<A1ƬJ�Zd�D[C���qR�"�	w�'Z���w�l`hj@�L@�u�&+�C!�'�1O$�Ş3�1�ݴ�y���d-#�#\&V�B4��)�yB?O�a�	�ў��@pt���(�u�c Մ`�L�$s���'�'�6�.$�1O�5��)�*��s��:~�y�=�I���O��$j�H�'�@mᡆ�u���d�!h����O�$S9/��5���)��?��'�O�А!bB|�>��eI�"�f��i�<�,Od��s�h���� BX`4�Q�v�СNu�,c�4?N�4�'��6M9�i>5qu��,'Av�� �O(yi`PEp����˟��I�f޹m�g~�;�R���)~�\�"ڒ}�pä�Y�d����|�T������	۟P�	�$�CN)t���sD�Pfd�"��my�`l�P�Y1+�<A�����?L�i_&ł�o�+Ez�A�D�o��	4�MS�i��O�I��P�IJ�9f�2�W�:�(ѳ�l�U!�`#&�.\Z�˓M���`�OLi�M>�+O@���F�g��@���K�n�E�F�O����O����~� �d�<i��i�xLq#�'i.-ٴoD�Z*\��G.L=}:� K��'���'��	ڟ��'��6M�զ���42��u1���a��X���5&���^��M{�'�B�F�AMX��0����ΐ����!��jӗ^Y�)B��_95 ���?a��?����?)����x`�0�e֭D*��R�mٴ �X�BƮO�?Y��?�i���b�'���'!X��yRgY�P_�8ؤ��AFJ����McZ�;ܴoěF�O�����iF�d�O�<�lԭ%	&y��n��O�*M�Z�H,J���֟ q'�'���by�O���'��&ڐv�D�@G غ<�>刂^�_��%�	��M�K;�2��?9���rK�(��M���[�*g��� ��<y��#���n��M3J~:�'M��!�m�)H衸���LqR%Β�;�\�@A�R~2�O^��	�%�'y����NE�]H�+�
J�8���'���'�����O��I�M�ׯ�KPi���V���ƌ�%%@�����?鳾i��O@A�'�B6�,J>�m�0IV�f�A�hYxH��n�:�M�6��Ms�'����H������F��Y� �@���D�(�AN�O�\�Iby2�'��'���'ArX>]���yic�cG,.��$&֔L}n(o��|!|��Iҟ��	D�ҟ�A���k A�$�x�it	�.���s`ꅯf�f�t�Q&����?���iL�UnZ�<A��ՖM�"��)�'E,��0�G�<��-�
 ����:�䓀�d�O���\��p�b��L�
ઈ�d�����OT�$�O�ʓ����W����'�����<�iJ��ϻx�y��.�ғ|b`�>�D�i�6m�O�I+U�*q�VZ�$py���/`j������UBx��D���
{y��O��	+��B܀r� )� [�n�)s�$�y��K6q�p��*��x�e 'ʍs�R(d�TTz��OF���ɦ9�?�;a�lk�� �\H��Oњz�@ΓԛƩ{��o��bd\�n�<��*�������lC�y^��e��E��-���?))O���O���O��D�O~���O�TO�IN�<�tꂔaOz�q���O���P
7X�P���X�����OL�����&&��⠊��T6�Dd�����8b�4e��Gd�����@�|Z�'��"O�O��S��N�y�+���.�2���aZf~��q�%�I�L��'u剣Vn�a�����L�� �i�95����dB劣��(���:FIM�k��1rm�	�
��+Vaݴ��'���c�֌o�voڿs���""�$m����HY
E�`�	P���ϓ�?��(H�k�0��!������q�? hH�5'�cܒ-���L�L)}�f7O���O���O �$�Oړ��{�(	h�L`���=�h�Z�Bt����O
����q@�N؟���ڟ��Igy��W�`=�"	���"�L�8nR6�Tl}Bf`��o��?�Cw�Ʀ1��?A��W+9�u��b$GL��XUEP�R���"��O�@zL>�*O�)�O���O�0bI]�zx��0�K'j\q�%�O���<qT�i�-�$�'��'��F8��IR��"[C��"��-KA��+���5�M�im�O�럐LZ�'�x�����+���`!Ϥq~<�k /�N̮ʓ��O�O1�H>9e�?G�"=ڔ�E1?�&d�N�?)��?!���?�'' ��������ۦ�� �ԊX������<�x4"tE83J��	���4�?�)OL�dB}R�n�ع@�ϻ��Y��?n��acb�ʦ�p�4s���4�y��'zܵ ���?	��ORŚ���� C��=f��-f1Ozʓ�?����?����?����򉛇k
�
PU*;��	� :t�lZ�>Lȩ�I��p��u���4�����DA���L��A�9M�\q��3|��w�h�'�b>X��㦵Γ%�\��P�ʹM���h�ʄ ������D���Op8H>�-O���O�UR��P��;���Q���Aa�O��D�O �D�<y3�i�L�p0�'F"�'8JL�l�5Q�&���h�\}���dJuy��'��a/�$��f���L�O��Y"i�;+�����&ޭzwHبH~��OV���4����R�F�c
txs$�� i�K��?1��?��h���$C$�ӶF��=0tl�(���c��O�	oZ?kˌ��	��S�4�?�O>�;�8s4�����K^�o<��!;O��o���M�%�i��8X��i���O�ɸ����P��\h��栉����R�U����O�˓��O�������d��|1$)�]�-��$1ڴ4=A����?)����O��$*��X;a-T�R�Nŭ-�`����>i��iLP6�B\�i>U�S�?�[��e��р�aɻxܵrV-�:v��Z��^yB�١-����ɭW5�'���bJ�@�1C�]	K9k�H���ߟ�����4�ɳa��T�'&p6�ЮA%Z���/5�����g�N¶y��@,8�D������vy�O���]Z�f�v�$�n�}��"d��0+T��ↆG�`ɡ�HɦΓ�?��hS���	y~r�O;�����m�'�	z�(q �bO�9��Ɵ��I͟��I��,�IC�wC0;��ɷ���T"]#�����,�`q�	ݴ~u`�	���?��i��_�H�kϚ$OΘؤ�Ѡq�p���N��MS�T��:�4f����O�r	1`�i����O6q9�'Ũ��(����
���G��?��j��6,�O��|R��?���p��8�@���^�@��V42H�!��?�?�)O|�l#E� P�	͟����?��:-Lm�2��&K갛��C����I�� �'�6M�צY�ڴ`L��T����O�t �VF
&����A�!i.9B� c6�i>�2��'�l�$��@Ǝ*{�QYAEC�9�|;�i��`�I���	����.U�p��Hy�IcӾ!!�01����N�)=L(�
��R�
�����Ox��O.��|R*O.�lZ����CB�A�����J-M��ٴ}�&�ƿg�V����#͔E�T�~���؂j,XjQ��A�H����<�.O���O����O�d�O �'EU��B��ǉ&@��tVQ�dQŴi J�1,ۗh�"�'����O���'�M�;2"Z\05a��-,�2/?,^� b�i�.6�J˦��O���(��K�5��7Mk��J1M2 .,�H$eڶLb�q�f's�����@B�G\G��Ayʟ�U���2������+)�4���'�6�V�"��$�O����;B�(2O����� ^s㟴P�O΅l�8�M�x�@�	J����Vi[(7�p
��ϟ�y��'ն�c��n��qT�p�;Mc��Mß� 1��",�$MA�9�Eg�ܟ��	ן��I�8D�t�'�Ą��f��C�bm#"cF�T��,�$�'L47m��qEb�$�O�dl�R�Ӽ[%)_<So�p���3C�̥�u��<1��i�V6���-�J��IΓ�?a�֪M�|��^�_�`�K���;k�A#P��"3�D�O>1(O���O����O��D�O�����	�%j�50�J��r��i��<!G�iR�,�#�'O��'������9���'7�	(�o� �D��7�}B m�>y��iT�7m��E�N|��'��@��+�֬"D��2���t�[dΜe�V�r~"逪+�y��d��'�剶=&-Ic�Nu�T�Ɋ.Vf������bB���HB�Кj���R瓒j�@\AS����r�4��'f��ӛv�m�"�o�1|���7�C�e��d��*^/>��ަ���?��kNw����_���$���寱�=3��
-2��k�Ã~�X�Γ�?���?I��?�����bd��0&�ǒƍ���-'@K�C.�h j\ݟ����Mk�����d�OV�O�|�E,Y�Z�(I r��pX���ϊצ!îO|@mZ	�M[��*�R�4�y��'P�3&J��M�I�Fel�	"g\y��i����!l�Q�(�i�1�'�?���?qB��<8�XA�M��]�ls�[�?���?YZ�rX�p)K������,�M3�'p��qQ4���@�n��P�A�X��Γ\l�H�Y��y��'��fKr�!+^w�S�?��/\��$�j)H�$����͟���`�=/��������OB)M>q�)�����a)]�6�0�� G�?���?����?ͧ|UR,�Ƃ)�����(�H�!����򃍽[H%s�N�;$�F��˟��I������d^�8a�4zTZAA�"ß<X��)�AC.K{�A�i�V6��"-.J7M{�P�2
��o�@��O���� �2���5 ��U�`%�G�Q��i>��'���'1��'���'��S�Nk�i8i(t��@�$R-6�!�4�|��l��?)��چ��?a���?�;TU���v&�����2F;DL�@�i��6���u�O�i���	�$1��7�j��lםBr��������e��)D@A#o �	_Y�	cy�O_�!�"%�ܙ��<}U���k�:]��'i�'��ɫ�M˵�׾��$�O|	�BZ����M� �6�J�� �����^���	ݴ4&�'8�x+$ϐ/Pߐ�%0F}���'���j�X��m�Qy��?��6٨T�=�*޸HH��:�OجK;I�O�;	!�=�E��I��=Zu`W�^Μ���ضTp�Az�����C4Q�n)�3�T5�zp�Q�wE�)6���1�4)kq*g�te���u۶�2"):���,� ai�7��6WE,�r���ؚ����/�J�Xc�</X��-�!^� QS.C�;�Ss@�+��LB�;�4�a�*[�tq(�;j�P����U�w�: £(�(<A��c��&�4�/!h����:V��9��r���Ue��@aB��H�Y���������-ޫ2�QQ�
e����'T��su-&�I͟'�֘#d�JXCP�W�3m,�e+T�Bd��%A��<���?i����
2'%�p�Y,V;&HP��V(وU"\I�	џT����8�'EB�'V���i2,�t,^^	zl������'!"�'o2S���F�%��T�K�Ga��Ae�?t�� �ë����O|�D�O\��?���C� �O��h���S5|���&"�r�@ш�O����O����<wh�H܉O[�d%yJbLZ��]!pݖ�7�n�,�$)�D�<��z�H�z�kƃ�]��Aʭ�l���IWyRH��{�������kl�#R/4�)SC0��Xҧ��q�VZ���ҟX2�9§�n�1�d�0�)�1���4勚�6�<�U
§D\���~���
�PP��� :	�0,L M��tu���$�O��S)�<�O��L<!w�~��b��<2�V���^ߦ-i! ���M���?����Rƚx�O ��c�(Rh��K�GWJ��PR�n�؁�Q*�<Y��?��g̓�?�0/�e8����Ř:-MƔꦍK/��V�'���'5n�j`k1�4�����O��%�ʪ<�g�n"@���T}��'��oQ���'�2�'�be�_��2��؂cK2���a{��d�N��%��ʟ��Ryb�ߎTӊ�ia���dpɕ�*��7M�O*�@���OV�$�OPʓ=���V/�4v>uك`F/�8�!k�;��'�"�')�'��Ɋ-�谍
/��� ��T��:Y�v`<����	ܟd�']���kz>��`�:��D���du\� R��>I���?�����O�i��`h����c�}kL�c�_/0w̵S2Z�H�������Ry�P~$���X
2C rlz�rB�d&��q���-��ϟD�'���'��s��TGm R乕�@2'��A�
ܖ�M+���?A.O�Q��\v�ڟ��s��GY.-�����	TD&`���p��ʓ�?)���RP�|:��n����)�N�	w�� �n�E?�7��<q��! ���~r��r6��py2+"�@��^;1��I4*u�d���O\|�6�<�'�?�g�I��ZD��'�4�ƌJ<7M��}����O����O����<ͧ�?��"�r�F�׋��L�R�U$�4͛��R�
��k�y��i�O��PHY�<T�q-�YG� &H�զy��ȟ��	�"�-�����'���O�ܺՂñ=�P�@��	p��7+R̓lv�R�����'��O ��Å�;mx1ׂ±�rE�ip��V�F�������㟄�=y0�$`ru9e�> z0xr��e}�bE�-p\��O����O���?���	�H�0sL˯?��-�  0���(O���O�d"�	����Ŕ���X��q�j<��^
I`�%�vb1?���?�(O���կP�P�ӈr�<��H��Hׄ� o�7�O��$�O�⟠���@��Mc��4�b?@g�ј���B��{�_�����h�'������џ`BqF�6e�da7�,�����^'�M�����'T�R�\�N�XI<Q!Ɲ!	��)�@.��v�LDQ�
ɦ���syr�'_� �^>A�	ȟ|��?C6�{�,VLovh;R�N�Qx<��}�'za�2 ����)Ү;d,]�&�}9���qgޫ-��	՟<�a�Fޟ���ߟp���?���u7G ,[[dɀ'�^/M�,X$d����d�O�� '��^�1O�����˄r�r�qu@U?f������i������'�R�'���O��i>y��_^�'�Xv.��L/�~���46FV��$z�S�ONR�_�Z������ޖ.���{5)�!ys�6m�OF���O�6O�<�'�?Q��~r�
`h���	Ƃ��A� �xPc��i����ħ�?����~R�4-d�x�#AˡV��1������%[,˓�?����?1�{���Sf$0���5�Tib�Q���D��#��P2������T�'x"�\0_����a�).�T ���;��5[���	ݟh��h���?��^
&�ܙx&KO9��h��N^�a�5!Bv~2�'��Y���Iƪq��k���b5o��͘Q𔊂2T�=m�֟l�I��?a-O�B��i#��r�M-V�`y #��`�����O6���O�˓�?ir�A�����O�u����A]8!�h�H����2O^ۦQ�	c�����=7�'�~��&�8L�p���O$ش�?q.O��$N�B>�˧�?������� �� K5QZDVm�/`�q�B�$�<	��J��u7�SU�N% �J�J�v�a�"���O�Y˧k�O|��O���D�Ӻ��@;$i���6$�;U� ��Ҁ�\}R�'ՈY��)����OL������n@���-�����ڴp^J�y���?��?	�'��4�F�X�U�xY#,�x:I÷���g�Am� ���0�)§�?� ��A��:�q6Myskݿl�v�'��'/���Q��ϟ8�	C?��Vv,A2�P,��P��K& a1O��{$�Y��Ꟍ�	e?��i�5D�sh��Q�����Ҧ��VD )�'!"�'����'WV��@M�#�^<؄1!C�I&@���b >?����?a,O���j���1��?Ś���)Y�yb���.�<!��?A����'����,lج�2��OE�����B8ڝ3w"U�����O�$�<!��d�4��O� ��]�l1�,?tvEᖠ{�����OB��,�	�Tjd��=s�7�	�mXd����7ep1ZekF5���ܟ��Igy��'Gf��6S>��I�6��Z�i�2o��	1�Y�FU��4�?ю��'�BE��+���e��&bލrТ�pP�VF��En͟Ȗ'��b�2	�Vy��O^q��hZ�r)�-���A?o%:}3��0�	ɟdr&��
4b��'QV�p���I�NU,Y��˟7'���'N��_���'Q��'��$Z�֝�=h���
_�2�b���+^����?)�ǵ0���<�~�Ď��C_��7���d��(�s AӦI��͋՟��	ڟ4���?�����'+��'.�;W��=�D��i��a�Lu�^��SM�	xf1O>����<�����
�Q�@�5 �"C2�z�4�?����?QV�"��4���d�OL���wa���$!�,�3��QogHă�y���Y���n�$�O��ɸd�x��&�U�R�i���Zu�7��O����c�<����?����'l��z�!W��8Y�FT�l�5Y�O��;�.O]���d��{y��'��z��̌`�&m���Ƙ%�q�A��2:�	ȟ4�Iџ��?!��vّ(��}V\%y��K�W�Z� w��bv���'���'����\AGy�/A�{�,[��,+
i+'c����	џ��Ie��?����:�=l�F��ȸ�k�^�| ��]M����O �$�O���?���C/����O*M��*��<�,,I�[����eRئ!��A���?y'�ŉ'ې�%�X31�^���ř3��^�0:��o�����<��S>x�-��˓��E�Ma_�z�	?z�<;WO�="}�O����jz�b��T?��ëK�h�,%[	[;o�@��̸>a��#h}{��?���?��'���V�p�d�hH�C�Ѻq���\�@��5L�q�1�7�)��)5����!)ݙ9�� �g�6�b7m!9����O����O��	�<�'�?Q��٦Rp�E$�Pc@���,�X7mܼL.��2s��S�|��MC
:[��#�Ҋ-u�U��Ǻ�M���?��j����/O�I�Oh�D��������P�mM�Bp(�4���'�r����2�I�O�����`�N�i�	��iގ$��@�q����L�M�˓�?q��?��{�]'\�(�����x�B&��DS�X���2����	��'��*�" 2�|�$ʯ^�����P/��H0R���	ҟ ��L���?iW��","��YF�V=Q���8i�:`:ՍU~b�'�_�4���i�M�'��֢B�)���@�9��8nZ��X�I��?��ii�Bg�ڦ1�d��6X��C) �M�"�>����?�+O��$��yA`�'�?	ֆY� V�=Qă�`����+N]��'��O����*?��{V�x"���́����|�%.μ�M����?)(Ot��H���'��OdF �W�I�:���:V瀠-&�����>9��?9�V�8�Gx�ҟ\�2�"���ɹ��6p"�ћ�i�剟Y���4�?y��?q�'m"�i�YC���2� D.�t�  �c�p�$�O��З?O�p��yr�鉿?W Q+�̍�$���(�o�q"�f�C�jF�7M�O�d�OL��s}RP��k�*��3!�TH�a
� ��7-χH+��O6ʓ��O��|�µ;��Ѷ6����T��?��7��O���O
]X�{}�_����W?I�H@�x���c��Hrw���.x�&<\�<����?9��I��:#��%g��I��U�Sk�	�úif�e�	"�r�����O�˓�?��dX �s�F+M/�㇅!W)����̓�?���?����?.O�)
O֗���9_��r"�	
�p�'��I؟d�'���'`��\,S��ʠ�±��=J�j	0rH�OF�D�O����O�ʓ-:�є0���s����$�2�֭B�,��ӱi����X�'��'rg�$��D]A�>m	e(
o_�����M���?A���?�+OV��Uw����5��G�h��	��H�k�hX`kJ��M������M����?qF���<�(O�E�e��T�l��'��3;2�1kRȦ���ğ�'Zд��*�~j���?Q��)Z45����<zSN�Ɂ�ɔ_�P�P���	Ο������I|�IJ2RO_7|��3v ޑH��L�\0�o�~y��1O� 6��O����OP���D}Zwm��K���
?zA���x����޴�?Y�n*`����O�REX�J�{G��	���?),r�4l�H]�D�iTB�'���Oh�T�'Bb�')V� XH�p���:����ꚴ,`�m(Ƴi�ތbD�'��U��]����8��U15"�+�%@;S�����W<�M���?a�sV��JP\��'���O�Xj&LM�-ڔj��B'$ζAjкi��	ԟ,!�*��'�?���?a&��4Hl�����5q�q�5D�j����'�h��!I�>�.OJ�$�<����]�.M>,J��� ��a(��i}m �y��'�"�'�b�'��	�d��P{�G�\�d� "��v�u�1l���<�������O����O�!�E#!o�zh���H�x|�t�6M3K�D�<��?A����d�@��1̧Ag���aך_%�a�����`m�Ry��'K��ҟ��I���v�0�a�ԉ�Ȱ	����1��������O&���OF�N����S?�����藬f�����XV�ra��ͦ��IEy��'���'=�j�'(�lrb�y3j�fu�=h�
3֎yl�埞:u��W�ɲW?�Iԟx�S(<8VP7CD�#"X��G���T2���O��ON��D��Zy�ӟEH� ԙ�p�x�F)���i��	*T(����4�?��?��'c��i�����&@!>��DI&����+i����O^���4Or%��yr�)��S�]9L�U8��S��d��&M#+�d6��OD���iB�$!�>Q-OFLAShT6{vB���ڤ-�f=��C˦Y10f�@�Ily���O
e�Th �d��
���@��r�i�ʦ���П��ɴ/�2-B�O���?��'L~�H��=_��LIQBN2e�Nm��O�˓2��x����'J��'=R�c�a@�!���Wi�D��Jb�0���\��@�'�����'�Zc���!	�"���Q ��*6�v�Y�4�?�fm��<��?���?�����%.��I	S/��Y�vDہˀ�J�K�AT}2S���Fy"�'R�'> �������2b;p0�Ba���y^�$��ݟ��	xy(J����SG"��0�+&1�0rG���}�6�<�������O��$�O �q�6O�D�#��kvҝ�.���:�[S �O}�'0��'��II֥C��B��ԅ��p�e�@�x��� 8��Hm��X�'��'�� �y�\>7�B��^XBT	������_�o���'��R�t���ӳ��	�O����nV�$P�N���:yj�>9���(�I🨹��"�'������\�M t�x`林Dț�S�HI��G��M���?����bV���5�A�3�^9g�Ya�鄵M,�7��O��DD�J�dp��'dq�@-�D$�i��U�#�_�"qB�p�iU���l���O^������'E�	)"1:���F�O�D��F�9r�h�4-,�͓�?1���?��t�'7ru)'�U�i���cd�U�G���@|Ӗ�d�O���	�6��'��	˟��6�%B�kԆpn`��BG*T��oZ��	����DDu���?���?!��&����� @ȆȘH����'}���"�	ǟ�'��(Vz.ɒâ��u���r�5*�B�z<(Aϓ����Op�$�O@�M����0h���]:se�.�(�yG�U	u��O�d?���O��M��k0�_YQ�)y钶�٧�'|B�'��_�d*�mڀ�����17S*1���(��`ك����OZ��*���OX�ZM�����G��)4�_�y��M����=~�d�'�B�'�bU�|xI���'l
�!��aY�t5Fra"�"H��!���i���|��'��Ş�yR�>��l�L�<Q�G"\z��9f��̦��	����'�h�`6i0�I�Ob�i 7<�0c�oA;6%x��,.M2i�'z��'I"�G/�y�|�ٟ�s$Cʱk�^���hC�v��X�d�ǵ�M`W?Y�I�?���Ox@iV�3�b�C/�s�A�նi�2�'I�{��$.�s>Lz�ؖb���;gj��fv6�Q�m�oZ⟜��؟T��ē�?����(��9�5Ae���A��N:h4�֫��4��O��?Y�ɓE������]"��q�.�#u�@!ڴ�?���?�@Q(A�O��$���3!� mdh�ї̉6sf��Bek�"�OtH�2O��D�	Cjg�NN\�U�^[]��01��զ����T�(=�J<	���?�H>��(}<}��+�$u������mC�\�'l	�')�	柈�I[�pX�c��M&_U���F�5k�0��ʏ��'��|��'��˜$S���;�������Xsˆw(M�v�'��I�$��󟤖'OY9��r>a�!��IP4Hy�R9@��.��O��O��$�OFH����D�"��f��)����_�!C���?����?*O�"���c�9R�H�H��ȘX%�]�㬛�+2��h޴�?�K>���?���F�<�N��U)^�s�8Su �<i+�$�xӞ���O�
	���#����'$�\c��(�BQ 6���S!N9"qlt��}B�'���'KRP��@��L�qAքj3b��m��	�h�oZԟ�������˟h���x�͟��i��)�hȡ�*�� ��%9&��1�}����O��
��I`ܧvm`�� 0�[�fN�-�tl��G�Q��ȟؕ'��dT�ȕ'�6���Q0l�)I1�ֺdΊ�31�a�<t��,E�Z�1O>}�I2F��H�5�-?D��"�H��,= �*ش�?���?��I 2�Im�$�'G"g�F�9���=1����D
5w�c��I�^�	Ο��I֟�6�Q7}f���&&[pQ�1BY���3L����O�ʓ�?�L>�� �ҴEgF`0�-+XI��W� 	�/�<^���?Q��?���?��
�'���fA�(�zQ�ұ������?a��?q��䓓?y��2�$�w*�M��	 �̑��`�g�X�L�''��''�R�l�[�(ΧJ�T�I�kJI�p��E�#�tnZ�H�����n�8�j`��'���6�%Zt�lB��C
`HJ�O<���Of�d�O���Aw2�'�?��-C�%}��;1�W(�0Y8�FHz��'7�'���'X�e#t�ș��D��q��b���a��l���'���q���'bb�'(�TN�nI)�ǣȒ;h�M�pn�6_b�O����O\ݺ�֞:1O�ӓx��2�Â*L��y���#p6��<����]��f�~�����(@����;G��9��->�(���d�����O$�"5�)��`�L�+f��9 ��j`�KO(6mъC�:=n�П���ҟ��S���?�d*GC�� ��0Y�#���/כ����O�?����!$bբ�5����/TTŸ�4�?����?a�Ǫd4�'���'��D�.��<
d Jy6Y����k'�O���B�d�O����O�<�b,�1f�[e&M�9XR��\¦!��$x���'��'�?AK>v,��D̖�S�i��}�^p�񋌦
��ItL�b��eK�I;28e卒d�7��j0��G�Lo�q��v��y�a"OƼ
P���MZJ����t����4��0 ���ET
;��"Gi)DA��0@�d�� 5�������	z|��mLFo¡����"Q;�F�H����� � Q�c��5� $�Ҁ_*�x�5H�1�T$�(�$P�@�
�H��9�3�G7����a�7b	�m�޴�pnݾ$a�m1gD�AH�h��G�Y�`u c��XR6Y��O`��OJ �6�/K3��c��qy*��M�5FO:d:�|�Ug˖+.�1��	.N��A*]W��~�У�:؞��# ���Ǐ�O�'�,���ٛ�d'�	�O9���+�`�[T�_ 61��'l�O��"~�r��A0�΍ck���s��\�$���!�ēy'>� ��Oǐ b"�Y1zD*����Y�t�iM��'��ӡ(�u����L�ɴ�L]y!l��58���EV�����J� �&!j`#J9d��S�t��'�N�Kν:J�\��f�	X� �N�n)>d�R�.	����O?��Dr��w� ��ů��0;�\8A��O��D4?%?Y&� �
�8���M��e��!h#D����mŖU��l����[���bdM"�%s���V����_ bղ�*�@Z-}������?y�G#`�J�R��?����?�������O̘�S��V���J�z� ��!AП�f(� v\���^�*��	�e�v�B�I��:<�)Ĥ�7$�d�a�,�ܝ� �Ԇql��J�i�?�=�-K1��,�rFK�9�B-��}?��g	ܟ�	S�'O剞R�T)HV镪c��L�@R"�C䉃h���x3��.6��A�ba,[<�HO��hy҈ h�6-�S���J�D�4*RX"��)���$�O����O(�(e�Or��g>Y[G��e�Y9i�^�*a��	(Y���'O�4,V�l��m�ox��jdhZ/vb�W�E?|�@�i�z�4Qpg�Q-mf�p�J4�Ġ�TJ��F�Q��q4��O�����{P�ɃC�>����aJ~�=���(%<�q�J��eĤ��3Oѝ"!��I�M����%]39ĊeH�n���C}�]��@,X�����O�ʧ�<<�QL� ̴�rw� *T���+ݣ�?���?!B`�x��:2J˲)�lQ���@ Q�.l�q��>%� q���J�@	Q�Tpׇ�;f������&���o'�
s}��I^45�y�2CC!i���eDh[Q���E�O��%��~Q�T� �B=/^հ	��dwp�e��d+�Ϗ6h<d��UV�m��%�O�M%�h��%߸z�j����/CM��2��g���q�� ����Oh�'H
�z��?���cx������tdm�3�]�Z�hE���E�_>�94G����S����'�2����ȹ&�������-���.ٓC�T$jӮ�I�ԧ��"!�X���:!(�Sp�f�ַ<̊�'�"�����O��0WCH56�@tX#у ܼuRG"O��;�!�T��) !M�$�S�I��HO���;!Xp�՝U%��l��wHP���̟�B_F>vM��ǟ��	��$[w�2�'��-X5ƕ�F��1�=M����'�D��7�'��-�A��[��u�a$^���X�'vY��'�4��bHN�zH�p�Ȅ 01#�'-�`�t�'�6�^���<!���Ȇ[��͙�c:ڠ�@ݭL3!�d�N
�����E,��c�8n��GzR[>A�'����1�aӚ@�0���y��u�� ƕ�H#� �O~���O@����i�I�O���,�J\��'�OH��f�?�B�3C@�"Ҙ�2�'�R̪�,���?�W��	+R�9;mյ7�z���D�v8����J�Ofl�8��ab7)�))8��T`�n��۴�?Y-O�$0�)� �(q����h�!����K�l8��"O*Pa�h��<��8�L�(P�ƍ��8O���'���6����4�?����.�t�z�������Ұ��?bh*E��O�$�O�u�Р����<�O`��j�c��H(q�4����
������D"����jD��B��_n�(�ɖQ�'�hY���?�K~��z��d�Hĺ4�H��3� ��Ԑ�������䒝p�
)+�僿X��tӀ�<92a|�I$�$0�jį� R-`�+�h3�$�Ȉl��H�	N��Ӕ���'t�%�4{�\`���V�i�9�/T�N��t́�1O�v�b�rd�ң�� `�Q���ן(�� f�ʝ����y���'\�)�7��;N�����O�:�\�
�ߢ}B�'�R�'Z?���i��1�ꗚU~�1�f��I��D�O8���B#3�DNC9Dk���7��&x���"���&w�*�$�Զ��!n�&(P����&>�����O�I��H�jP��Ov���O@ �;�?i��aG*P�w�5��d&��s󬈙0����=$�r�eoV:1U��QL	&j�Z��d�а=Smǀq�����B	S�V݁A���?�����?q�i��7ݟ��՟��'��Hr����(A�l@9QC
�'|.���'�[��bwh�?_8���1-���i�<���_:��V��/D��h�-��ZҺ4�rƚ���'�"�'7���p�'2?�<��qD��?�y�AӔ$i��j5I�V�Xx���#4~�MA�a4b��?yK )�(@4G͕q>t�#���{S(�����@��࠴��
!HɌ�d�g��r��A��ʒ5�acTg �y������U�	ay2�'��O��5M tIȋ^!&����8,jB��M��hĤ̑�\Q�R�[Tf�	/>d���vyҥ\����'�?���r#��
� �  QMR��A�M0oO����?��I���	8��xǆXV*R2�&�?�E��YA�#%��	P�-��5ʓ��M�F��h**���c�|�x�)Yd���@o�
A n)��̔b}Z<��a��4��d�O>��a�r���	�;�V@s��yV�� �ᅁ)!���](��GF<֘Q�aF�a|B)3�đ:khf�!�cٍw5XX[�EP�9����q-��l�˟���k���X� b�'��H�*M���拚>�)���˅�2t� ��t,6�T>��|��6���c�ɲI�`�g���w�9�s�����J>E��]`
e���F�Eƪۨ(X�%�P�?�G�i,\7��OT#~��cA(a�vb�5k����*.��	���ɕ hx�m'������t�#<Ye�R�4�_�qy��Ä�6~K��J�U���'�,�7B^+��'"�'C�꟰�I'"]"�V:�P��5��y0l��	��@��F�w؞Lx�'�26"��S�Շ�ѫ����������T��h��y�r1��H3H7�P˔�B�q�X��	�i���	�MK���,OH�d�<�f��|�Z�Sg�D)X���p�k�<�%�:
~���ƚ7��tC$#�0�����OV�	�V�bY�ڴY������)�(;tK9�d����?����?Qc^&�?!����T�ߖ �>��tͅ�)�Xi�Q=���'b�
%�� R�"D� ��y�M��Z�S@�I�t�!9B ��:��[��-��1D%ԉpT�'�"��O,���'n�6��H���(�Lx<y�c�U$�ʦI�?AV�s�,��hōV,��'��:m���˴(2D�A��5� dO�(|~�Cd�o��(�O��k���i���'�哤2(��1���7T�<Ң+��N[�(�͜ܟH����lpf��-�jmx�-�-5�ꡫ�y5�In�ѻ"�F� M��S�F�;kLQ�����~[ju��J)0M$=R� �&R-Bd�f�<!��
�O�9?d��hg��<D:A�@Dp��=D���OГ�0��/"���:�%<	P�л5���!3z��(�)��<���M97������
y����fL�H�4(H<����8Ҥ,@��� ;G"��'��Ox�����?=��x�'l�'���Y o2D�l��܃u-*]L��l��"2D�p�A�v��q�"^��� �/D�ȀE��-�.��-j�2P1��-D�zg��.�����@�h�*0I��)D�xI�Ѻ#o���J K��	[4�4D�x) �׭[��;�$�#&��!�(D��!c��-��d����l��Y	@�0D����C�bӀT�Vg�	�.D����i��S2�Dy��^�-�� ��1D�� ��鵋�o��h�AV`�R���"On����`�H0s��5�`��U"O^�h�i��j����e��X�"O���K�y�I��*��G��)�"O����BZ�pvLE�	�6,E�}PC"O��"ϓ�Tv�i!�
G(��i�"O�PQH�g��I)�g"�L�
�"O���K�	r��!2w�^�,�("OZ�*�"ĺg����S	��=+�"OX�cċ>q��
��ІJ�!�"OF���/H�8i��D)1<H3a"Oa���Y1p�>!�7���`��A"O�(p�hËc���3���X�&ؒ�"O2�pB�@�}:%iA/M�Z�C�"O9�BA4{cl��⍎S{�6"O��)uYk[��HβD�I�"ONݓϤ\mByx��J-�Ĝ�"Oz@zq0��R!cO�T��H�"O�hk�+~�Z�C�����y��"OJ�R`̓�'�A�j�����;c"Oʍ檂��� G�R��"OЀB���6(Xܪ"%�iz���W"OD��qE�7��-�an¨@�$��"O����^8.C�M��n%t�z�"O�:��ēF�.�i�EW�����'�����7t�\���8"x�)�'�K!k�B�S^�J=��[��΀����$�`�t��I`�r}
'N]��.�be�	=����\\��
	r��h��E�/!D���ť,,�!�oa��j�88p%����	�:r�>�y��]�;�P��u�߾b�5s'�*G�X�G ��>�z�x'�i��}S�,��M�O�4q!��yGޯM~�Ku�L��l KAȘ#�xOΏv���H��V i��"z��(��c��k�����l�O�)�#�����D�oN�O�huH�3J���8@@܄$l�,�0<��B�3��1S1-)"�f�+$e�Ia`̊vb�R���/X�U�H�А׎,��"�!��=) ��%;�HE:㊴��S`�~r*�5)���i �P�����O��r}���&��5�S�OV{eA�[��Kv�by���'������<����eȜ7?����Ff�8d�@���;��Y�*ƽO,���R>0��W�\.��	h*�0S���=(�6]҄��)KZC��)(�pqK3�H�@v��� Ƹ�������
vcޜTH�XB�J��*Q��Q� ����?�P-*Mq�	��<Q��H�g��`�h�WF�5D`��pK�[G�|�ģgT�`�ȉBz ��JF�8bI(BU��*���<�`�ߡcD� P�x*�r��BdÏ�
�� ���^u������	H[}jiХ�U>�M���B�9���W��}����ӿf^��HP���<��\�C�2A��i�H�D5x��g�>E��'�:��тo©Z�� �dG��t�K�P.�,�v*��!W@�`�m:
�V>}+�)ɡ!���'J��#�>�\�y���>M���x"~��%�տ�,���3e���� dSR�Ze:P �sPUӔ��+
�� g�]�c��Qz	D	a��&hK(2V���w@u���O�d�sI_�9�Ys��\������'z���Ŋ�$$Rq��	^�2ػ`#K7G�D��ӡ�x�>P�5&�%��u�O�d\�W�|D�b@��R�:5�!��A�#����Ԅќ\َY���ߦ���y9���k��-݀0�v�˅{�1�';�l��I�?�2`5i�n���ԊE�r� �CV@pѶ�G�TH�jT,����97ʄ�>yv.�97�A�����̊��\�'��pՂn|P�'O�d:�>��O��ᔁF0D��(�ˀ+ �����OhA�@@�&��,���2eA#\*i��Df! |�1�g�>�TR�ax��I�Y����������g�(Uv�=�@h��0<�s/�[�@���'S�apç2�`��*f��5���5T0�=I�O�,R����-���(�Oծ�r���5\w����l�^WT<B ��I~�I<��z�H�S=��1�'�Pa�E��Wâu@�iLc�2���c��<1�$K%`��3�%��?�A��"C�tB���D�T8�@�4qIR}H�])f�H�I�K�O����ڄ�O�Q���� ��g����%��O�xt~.N0��I{����_SL�gI��D�4DC�0}�ǂf���)�3�i���;N��!�$�l��J\�[�H��1�����1m�s��X Q0��9R�E�R�ƨ1��{̓Ʃϓz �B�U�d��S�N�Y$A�e��bEn�6�	V� �`��	2C��ugL�0�B��ICJ��4�@0��0�6ϔ`�)i��i�$�DC	���0&
b�'�s�P)S�Kz�� ,ѹ%�Y��:?Y�IH�3�&��+j��}afA�}�Ӻ� ��b@Α�<�Ze�s��+T����<O���D48O�@��I2�� �*�6��L�U�$*Ld#���( )�Pj�a<�)���[%WQ�֘�>tF\��'Q�#�~�n��Y&C�I?z�z����9W XV�H�jw H���X�*��OJ�	$)������-!\<r�P֕Z�cޙt�����לsi8�A�-�+<R���k�Ho`@�3�M�� %�?�4�'������8_���fo{�$Ƴ&��z�H�<k���Z��(��DQ�XO�����E	s�8��Kؚ��ɜSC��aBA֞G�T�R#��v����<f�d�{�C�ubh���S����&�B�V?A��jޱm��do8t\�T�����\�9�� �,&��?c���$MO:^��l�%(܇Ղ��d�<R�����q �K��^�sY�M��"�m1�I�	���O���VeJ$U� l��w�v �Wo�0�i���"R}PQ��'rv!����^?L0����..�T@J��ޝ�~b�	=vpà
B"v�m�dB��hO+I߹4���`uD�2Ĳ�i�e�l8��X���1MJ4�Ư�}3���s�C=B�,�����\ʴh��l��>��'��2{�����el.,��F�'6�R}S��J{axriɗtJ>�+�⋒N'�I�`x�0�G�τ"v�A�	��Br���]<"
�[-�}V��@Q�;���i�o�M1b-)4�ĺW"	�&��!�"��4cV�)�'y_��2Ǖ�;a� ��h�ؠDx�;Tr��qa*�W��0�*,+Q�Sy.�%��G�
���a8�v(`UL�� �剦]`@Q�%�$�3������*�t��A*D_�j �p�����o$*:��"*����@��I�8���ÅԖN���Љ�)\�Fdȗ��,~�Hl���-83�Y�R�
�X�I�h� q�Fـ7K>Obt F�m��32�p,�"���}���It�@ .ڐX��'��rU�Ր8�QS�-\�B�k͙E\Px ѡ3Y����O����@g���!�� �t�;��*O�d!8p.�O��J �-RN$u &� 7 Tr�	�*�s6_��h�� M�A�0��?i 5xCP,MJ����J�;N��LCmZ�<ѠL�=?/���`��`X�4zK@L�'�\��d��;<�M	�I�g`R�#��ݥy�v�C�ޖ$��A;.E�y�l��{��L�A
�����>�nu�4�	8��(邍�46��P��F�c�თ�'��k��\o�:�� #�u`T% ��yr��WB (r�BA%�~N���u����j�>�9Cb���y*b0�O>)�3�B�*|���ƃU֦<3�A&�V�۠J�Qx��O2�ډ{����?Yaf�.hFH�uh��jYnSdݹ#E*a2��,3rqGxbnS.]��r"��7Ϛu�`j��yR%�#�:X7nZ51j2�-]�z�w�L^�$��r�?'��[��J�1S��S�⊌�i^�C�i��~�DJ�d�?`.�ٙ2�=`&�Ie/Z�P����'�^�A�a��P��EH��&Ǝ;Kbu��-�:GSL��g႗m��Q�,F�hX��q0�D>�.y��	)f��I�d��ǎAz5��r�n�`�o�X���S�.�j�觟$Q6�gO1O��{b�֚Y&��R��&VP�ӫ�gj����Z�Fq�S��#��LIĸ�D�"���.��"'㇈.[�\�v8Fx�ON� #뗨n����GQ�$�S��U����ie�'�8���܍6*�hB#bމ�.@�'Q��*-���B���kQ�� p����'� :T�(�+�D��r�&b�ʓ;�A+�I�X٦i��[�Y}���'� ��4��m��O���ѯ_�<)�A�Y�h��K�<�;+����)ڬ�˔�������I_
x@���&�K���\B�A���Oi�%)�4h�Qe�ES��ȡ�����P��@�4]�����)�O$H��m�0���ʥ����ҝb�K�,G�̫cˋp�`�ab'�	f?���ě90_`�cf?�Ty�ס�g��5��
 )��!�G��?�
�r�O��vE�!�DY�W��c��5 ń:�	U��0@��:���!�*]�@a��.�j`��FP�>y3�KA�J��b�H��[�	5���U���`!y(2ɚ&eê��T���
Y
��<I�D�>*^�2Go�?dE�m���4��\���3t��AR�ˆ,���J��9�ج�V�	���BZ.�Z��f�͊-u�]��Z���S�,�X`��$��E��hc�n�R�� Ԓm��[�E�n�i�� E<�B,�1����?�2Su���%N7b����;9�,E!�@�����剡7�ZX�$J�PMA0]y�T{��v1�Mr�gX1AUё/^�<a+�w��Q�M@2Yq�t{��7��'>׎t�FŽ$)����T�����>1�`Qt9�]9�
5Tw���GG"��ӣh�m�c!�
38��t�=UK =��̤y�2M㴋R�7��S� �'��d\
���3`&z�ʩ���:qƤ���!x��a�C��
0�:���X?��B, L}bD�͔���p�8i E���\�m�%=I�����$��P��a����#b�q��)�#gP ��q����T�p����)�F͋�,��3��Ĕ:��t��z�4ct�S	c�JM�Ǔ^�P�Kք�����qP �ƙ�8� ���j��( <0m�!�~)�=3E-��9�od�ӣz��2	��	x��X�G�(=�b�� B��Dr�3��\�&�kRj�~�I׆D����$�;Hg&�	��h�tlJ��	�p��pn�p�\��b�ky�K�+�!�g��"�h���'D�T~�e�b 8��}cf�ǉo�BuH��D�OR�	<,�W*��Xe��Ƙ��P��4ɒ�<%�K��E�n팘��\��� �8�IR	4�@�&��d��#ءC$�����/����M?���\��MO��^�'I�)��*H.1R�H�C���I���2.�xB*.%�N9��,H�jBx�CU�F�n��Q �6i�44���~R��O�Hᣩٸh��`��O *��eO'7���c#���x��+r�s`��Ć+x���:���h�h�8O?�Zȓ�\�X��
�6�)��H�<��I<yW �q��E!I��&���S�T�E�N�q`��7j�"-�Ul��~�^��E=C^�]�2"Ŷ�>Q��?:�$A6rP�#cJ��f���(@.���e!�	�r&�ij�_�Bd�yR�*�|��dAF&_�N(a��S5.��׌�tE���02����fE�#�-w/���'�v�A����sK�I�ݒ\B�Y`�'�Rp3��T�9�q.l|�����`QrЫ�@�vd���'L$���N����!�xJ|����C.��S$��k2u`p��<iڎ|�>q2G��g���sG�.��"Љ�-����NK����ء�F�1 KK�L�Z��ɡ��0"���e8r ��ɤO�Q��
T�7��ʸ1Y��5H,@��UH�1�\R����1��?��O� �r=�h�^daQ��!x��� ��1��*��p<��՚h)���G�yϞ����M�]�X����M�?�~@���	hyJ|�	���DX \���k%o�0ʆ�J�h����	�FJ��H�`�]��ֵ~��(�'@ThHh�u!���ɿ@�P�#���<�q�>�����G��ዦ��z<^A��i�� �Hc�h�!
�0ՙ�'�6P���z!�F��,.���s?0�:�L�{��q���^�Z�k����D�0}�Ņ)F7� �ALi�R��R�D�n�\�`p+�Z�����$�jUN����'����=2�1�`I�jA�{3M�||�'��y7E�uX�T;�� �)��{��&�b@��K D��i¤��t~蒯D�ܖ�2�h!D��B Láj 9[
���d �q�<D�\*���^B�cf��D8��%:D�\B�@���x�R/���a�F/9D��F�]2t�l3%oD������(6D�t���.k<���I�%`l\���&D�Ȳb��[� ���O�t4d�#�O$D���g�
-������GK4,@b%D�D�� �w���m�<��a�B&D�4�W��5u��i��L�)=V�j.8D�(�e嗥NZ�u+�a�$Ah�jd�6D�����T��aZD�׹r#4	ɢ�3D��2ץ�"�x"(�'q�(U���3D� �TȄ Z�Neb4�1��1D���0�Lq$�9��/o����N$D��#�.�=J�ع�gO5x���`�4D�y���ei|�x�ʐT� LI"�2D��x5H�f}H2e��5,��)1D��S@-��62�L�rd�X���f(/D�Dh�o�!�@����m�\iUO.D�̡��6#Cj�)��Y8&�� D�D��f3U���D~� �
��>D�,81C�|�H�LU5qY�$�Cc>D����� n���UĔ3Q�x���9D��Bqo�{���
+�1D0i�E5D�\�v�Ȕ:��@��HĢ�2�238D�,��l��8����e8�a(�7D�d!	��g��̺'E�Bor����3D�� �%X�lA�)Z�	�u*F,;��%D�����	[fL�$$+J}4�p#D���B>F��!��F�1� ��� D�$����`����`�A�QN=D��csᎠ^��[6#D��QK��>D��z䯌�!�d�c#�1u���[v�7D��	�+n�4���Ǜ�\)٥�;D��c E���&����0�$}���:D�4����E�9�Y�B.D�h�qM��!�¯D��@,�a0D�,��ގMD&)p�J�2xs.pp�e,D�$8P��9y��p�6m_'M�t�4A(D����,��$H8�c�݌~��y���3D��C`K��pW�5�6)ۂt���#,&D�� @pXre�`�1"�-�l�Z�"O�e��$B.6<4�r�Մ�ऋ�"OL 1b�&qr�t˱n�s��`h`"O>l��̇E�Ԑy @& �8��w"O����a߃3]��Z���&�! "O�ݢ��X5o��}�t�)\�x�T"O�xS�	�@>%�P�*��"Oq��5H���V��)�Peӂ"O.���O�����8WFL@�^��"O|-��*��&x\�Q�ʘ�*�hK�"O�L��ˇU!̸*�iLwhv��"O��r��#@�]"(�E�����"OX5��ŕ[��c��
�5�j�"O�̹��P�kC\�����.�jtɱ"O����IU
"Z��#��$G�.�I#"O(ّ򭟆Nꊬ+�m�1�fe:�"Oٱ@T8s"�XˢM�:(!��v"O6dڗ�
b�l��-p8��"O~��!�Q�4�"B��XR�"OBEy�D�5!$d0CC/H2m��"OJAڱ暢q~�IP�gW�r���"O*}��KW�/�L��YH-r�ώ-a!�dB3ٲ9w��+<ରqºG!�+b��)���	?��aZJX>�!��!�44w�
4d��uh����w�!���$Kw֭��ɏG�F0���ix!�D�l��	��'%0`	� �!�$ړ$`28kU�Wu����C��:�!���:F�X4S%FW�O�t#SY"F!�#`h��+]!��TK��!�D�=`I|���E�8M)W)��1�!�$O�r����ڊGt��3�9h�!��ļa��H�qa[H�@̠���5`�!�䍪 (�t��9w�� p�ӳ#�!�J�f� ��"N�Di��t�^n�!�<mi
L��h<ZDM��Z6+�!���U'�V7M�;�bS�W�\Ѕȓ9�!��a�97��xEk�KG�@�ȓI��4Yr���K����TN!M�"q�ȓ+lD��aٲn��t �eD3-����D�zsƐ&K���3p��,O����ȓ&��$�T��\Wrt[��,_X����\h)da�.CSD� ��ʤ�ȓ���`��R'%%��em��t����Q(y��ӵB`� �`�xz��ȓc�Z�JS�:+2�3si3%Y��p@�i 	��h�|s�"������<a�,e�Y�p=õCK�3v�B�I!pN��T�W����d��Wu�B�II��!@�*ԴX)���FV�B�ɮk�����	�o���fCX*�|B䉱G��tk���3A��xrt�ò%�F��'�	�l.Uh��Q��@he��,�B�[#�0���1,���a�O<��Oޢ=�~:AD͔'�|��wÊ�&a ��@{�<93@T�B���S�bF`����Ə^�<Ad���Y� ɝ*ETK�,�D�<�D �s��R�jʴ���A���x��P�C��YbD���-�X��WN�8�y���*	�|�R�͂'x��n��y�hX8.�@���&Z���e��yR<���@�)"ހ�a�O�y2ͅ02�H �^8~��� ����y����r��Eb�D�`z*ܡ�m˯�y
� �M��!��9IDp��;c],��"OY����#
�Γ,:E��؀"O��a@.\'p��� D�:�d"OJ���֛;�Lm���ʋp��,)F"O@�jd��|0�<a�D,Z�dHQ�"O���vB֝1��z�"ӣ'�����"O>�agZ�k�4Ÿ��#�\ 1"O�ڳ��&��t�叓nK���~2�)ڧe�T� ���a��c#���T�ȓ0�VAHkֆ��!��-�2��\nZw?Y��6�O��z��V�Uv�a��P2Uv���2�'��'�D�0��`�(���G*e��	�'�@�B��;R����U��<��M 	�'g�m����5!D(�㥥�=~a\*�'FsnO;w�Z�3q/��p�O"�=E��eH�)� ȑ!�J9IRb����!�yҤKBܒ*6�R������y�	 2����(��4l�=⤬��y�KH8���[�S�,�\�2�N	�y�E�+j�`
��@�'��Ը2j��y��Q�E�x�[AL]	a����&�y�㚈7� ر��I�{|�⊇�y�d��K�J����2f�sR��y��(>���"�A/Az��+5`�.�yb�Yj	v,a7h�1�8����yRC�gv�@i�N�X=d(BF֐�y��Y9Uj��'cU�b�<���ر���0�h�\UKfD��Qю9���"��ݒS"O��Id○6m����REA�!��"O �pé��ab�y`�J�dQ�U"O��K#`�4k��b!�6c���"ObYAQ��"F����+ZpI�("O�5�dQ�������$T�A�"O��v!\�k�h��P�6&kD�`�"OB�[WA�	amb���_�"iн`"O�i�k��Eo�P�.�GR^� f"O�!�#�a@<����PO�L��"O\�@��N�z4��� �Ӵ	�$"O��a���k��e���t��s�"O@T���X�I�΀�gJ�x�t��&"O�͙0��@�hq'>ĸ���"O ���o�:"u��7h�q)�"O����(�,pF\���ˏU�rv"O�(O?T�8E��N"~�8���"O��pc�HC���w�61��e�"OJas�3i�1�3n�+��"O6(����o%f}��MZ�5	Ȥ��"OJD��BE�1�BɈ�FEO���d"On�Hr��/3�B��(�)5 �$�"O&0h���4�Px�Nf�i6"O���d0��}f�$p#��	j�O]�5��$��nZ� �U�Mz�Ex��)�$B�W��l"
�$j[ *G	���yb�8B�f9�2Ô'h0��a���y�dW<K��$��^�ty34��y�h�+X��m��� �`Aڤ���y��b��ٓ5�ʯmjD�Ri��y��.q�Љ�H��y�|$��"��yF�6{��`�BmVp����]��y���$�Ȥz�Ùjpv������y���ixAr�I&U(�)%��
�yc�oE�8v��#O=r�MV��y�K�8W�tPy�iJ�^�U�	��y�o�2[G�0R�Z�U6��ѕ���y
� x�bE��6���B��J�4,3�"O1��G���HA��*�0�"O�ę���H��1��k�r)N�"O�9��/��|QU�A@ tҒ��X��I�q0y��D?f<)�2���'l&B�ɈZ�P�[�F����Q�(^�o�B�	#����dU\������ZG��B�/ L��⓫*Kn�(ÆX���B��(l,.�[GHĆ�@e�5KY�GR�B�=B�qi�\+��b@�3	��B�D>�0�&c	(��F�us�B�	� ��)Ӯ=����1c/A��C�	�@K�A꒫X���i�A-��dxxB�If��<⡎܏y.���E�1Zm@b��D{��$��>�r�b&�Ug��4�Ӓ��<���$]PMr�Jǖg����4瓹x!����M�sLL����#[bn��T"O�d�q�>I�����8"��L	�"O�|jM�8@ƌxpAQ���)pO\i{i��2��=ɠ����`��9D��r��ԔM��5��Àe��}��7D����; � ��<L��w�3D�4���;XVi��E���VyD�0D�ɱ�OUd�pʷ��M�j��v�.D���$� ����@i[BCU�B�9D�{p���x��ݨR�:)x�"D��JqO��X�h��Ů�x���C&j5D�X����'[  �� �N�Ƹ�wO2D� �$.Y�Q�Fd1�⍫8l4¶.D����ߔ\3~dy5%O�z�2L���&D�6�V�/Jl��Wj�!.�LC��#D��)Ve��pU�����i%D��	5�X$gJ8�8dɅa>&D�=D�$��7	��"���x�� ��M:D��s��lI����,� ��W�+D� {W	�.5�Y�RJO�6�9��*4D���t�o��i[�b�*&P���3D����a@�Zx��tHT�e��(�&1D��F��:�$T����%M��� �/.D�0�c)��p��|��hת6ϖ$� �*D�8�G)���&л5�)$����!=D��X!V
I����;c�t�	%O?D���ġ���Ir�睸``����0D�$�6l�N�Zɰ���R��P"�0D�,��L��<��ԅe��1��.D�(b�'j��C�Ӌ��2��0D����(٤3�p0Ԯ���q���.D�PJPJȉH� �.�30�Ҍ�Tc!D�p�B���n�Ђ�Z~�d�� D�|끋�#����#o�=B�%PW�:D���t/�7	����eZ�
����f$D���Q��b~m9���_&ڙ�3�6D�P���J,,U
ÊV�H^�@�3D���1 !+���5e��%+Ntإf3D�,�Ɖ3"�<���A�!�<XyuD=D���r�=i��*�`O�s1����<D���7#?�$�c��|\�����:D�h�Mt���˙D���0F�6D���hn2�`����[w����'D���m�Y��A�$�Ҽ����qh3D��#�B����B�6���F1D�\e��9����~.�1p��0D��gԪh�ZS"b"��ˡg-D��2Q�wp>����1.,5!d6D�� 
��3IF���,�.jRPˠ"O� q *�=��(q#�L�9gv��"O.1Ĥ��s��H@*]�5QU8�"OQ�6nH�$�`E �	ڙ(��i�"O�t���ճ%)�b3:����"O��K�i�/�M��T<"P�x�"O��X&kI�zd���!X�.
`���"O`I�Ɉ��P�Ή!J��Q�w"Oܽyɉ DP��g-H'�@��@"O�I�Cn dժ��q4"��"Or�2Ώ��x0��o-<:D"O���/r�왂���=M.I �"Oj���H���4PD�B7h�t"T"O�Q�#��^��c�g��{�"O�t*�Z/wv&d���̀:�,�a"O�m)�'ֻk7���Ϭn�ި�e"O�@+��N�\�4�(�ڡOʮ!�"Od�:��]1d�1a�'��:-s"O�4�0�I�Fg����у[wƠ��"O�4�$�2U����@v�F�!"O�Bp�j�ƍ��*�Bw"O��[�G�Mx�Մ�9���F"O�`P���YE��1��e#�a�""OT��
�<�Z�X��
��A"O,�^�����,ˆ}�,ݳ`hX�<E
�(ز���#W�J��Kp�T�<i�HȽr/��V��1���[��O�<-mNR�0�U�ܬH�G	\#Q�HB�	�}��j�M�u`���V��
jB��:)s|�0A# q�hLB���B䉖1ЖHu ���6�Z�*�:5~�C��	mFx8VN��p)"�Q�K�MȖC�	)}�R�ڶ��"��Y�h�b�rC�%u0��F���{�$��R���XC�B�	T!:�kJ�A�V��j[�B䉍?�v�z!5��a)D�a�B�	�F/v��(*�5*���yb�C�IMo�����T�����}W�C䉵Uwjuڐ዗x�����]�.�C�ə&�$�pGJ��|�f�!TC��G��U��O$��0y���1�B䉊'�F5�#���<0��yU`�-q6hB�ɦpwh��Vh��)u�5 �Jϒ-��B�I�e�����ߊ9bpQ�",�o��B�	?i�A�L�%0hy�B��q��C� n<4Yɢ�Έf��AR�#�c¸C�ɫz��}3l�%<Y9I
{`�B䉛j
�Lk��^�(g��hN�<	��B�	�x���C���Lΰ��τ^��B�I1�]r$��*0ÊIm4�C�I�}��,� ݔP������9ky�B�ɨ^'^L"�K<B{�-��&��Z��B�I��YR�Ę/p���bF�*��C�I2c���h�R,yFi�EdP
!��C�I4&�d#�M�y ��B�K.�C䉵�@i`�ݴ\���zQ���Q�C�ɻ=^�ĳaB8R	��9Q�,C��C�	w�NM �i�.��锩8b�!�D�G��`�5�	�MW��	3�!򄊳Ϭ��ql��Mՠ�	ť�0
!���$��䕘m�-2e�30�!��X$#��4KV@�[��(h��@K�!�$�6���v��>�&�� (�� �!�ԊO�,1".қR���s�&��J�!�� *�Z��({�ܚ���3_��"O���w�<f��;���*�u��"O��ibݱ;�f���
09�2�Xu"OȠ�7�TY-���Z�D��dC7"O�|9��
,�eð��:fd��"O����Cܛd�h���c��pp"O�d���F;$D�S�ڜP���"O�͚�a
�/���2U��V�R�!"O�h����018�s0AD�`þyi"O��ag%��Ox���c�u�&"O���]�`~`Ij��K�ErԘ�e"O�L`���:`��e�B\{����"O��!��z������zp�$��"Of��`�� w��0���v���B"O(�c�E�x=&U���!N��� �"Of���+�zr����(����"O�IɥA�1L���H6y�LS "O���-��f~�I0g�+�����"O�u�g��hh���Gn9��"O�Y���c�������js6�ن"O� K#k\�p3��zu#b�m��"O<d�uCͶ2`}�s��*-�ix�"O.=�G] BW�d�@�A�u7����"O�K�6i6�aD ��lA��*�"Ol��T�B%'H���E T�#��-��"O��CH8l���B���qP��p"O(�V�Lr��M8!#�14l�hB�"O:�0��y��FaX�� "O����'�!�*�Y��˝*~1�"OJ��5J��hT	�	~0 �*w"OiҶG��&�P�H�1<��s"O�]����t� 1SsE�~&�ԡv"O��!�#R�����%FRN��"O�٩!"��
Ԝ`��N�`a��"O"4�hG78&9cU !=�P[�"ON$���:��I #��I�#"O��z��� �T�+�!T���b"O���J��2�q����|���`"O���N΂|��A�t������#"O���#��6Myp�bּ}� ���"OY"G��8�[�kQ�VW�Aq�"OPi��O���IJ&a^�T����"OTDR� =R��rt�ɖ^��Lcs"On�"�h6�ㅮ�F��w"Or!���3�Ԁ�p�K�Etnd�a"O�9���Y�ޠ���z��|��"O��� �[0Aj4Cv��$YH�L1�"O		�HZ���
cKܡ}bu�"O�-b�	I1W^ld���4'�fi�"O�����2>x X"��d�H�"O��� cǒl3���3	�����"O�z%D�;Z�(��
��4�lȻ�"OP)�'l�#���C��Y�?�|XE"O�p�caؚ@K\��QH�&y
��C"Oz<��AL=9�(z���{��|�r"O� 1%���W*�T�#HI�K}0]
@"OP�c�ME�^�����3(����"O���F����4b� u�L)AQ"O��V(B�D�q1��at�"O���wkV�Qo.U�B@S�Df.��"O�#fI��C�jPRiʃ@P&��"OD=Q���#\�0d�2gX�m�P�"O�5qb��m-�5��hӾrώ�A@"ORи�b�-�>�#ԧ��A���5"O� d$hHMcs�g����Mc�"O�Ib���5�X�ɴ���t��"OB����-v�$d�GAtv�Q�"OJ|
v�A=��\���h���"O��r�BΚ�<]ȴ�_cd�Գ�"O�y���iLHa���I=E Tz"O�x:���=Y��0�N9@���#�"O�`h��*��x��K�B�X	��"O��ҩj^���WŐ�M�=p!"O\P��T���U��%y��y"k�`��Z�܎b!�%�d田�y�U� ���`�d3*ǲ(C�
��y"`�.)��G�+$B��:�� ��y��Z��t0�&�+<UaN�y��Ki|)���ɪzǲ��g꟟�yb�S-fR�#�;=�v��V��ybiPgd:�2H֜HX��-�>�y"�ޛzp�H�բ��v��EI�j3�yBÛ�2�R�Js��%xhD��D �y�A8,��@O�r3j��(F��y�O ����bX+h��H�0�^��y���>e�Y���ҜX�xUc0��,�y��X���<�&�G1
�uB`��y�B�%G|� �����D���I�#�y2�C�f@J�� uC���l�<r��\�v�[��:T���3�CED�<��Ś	L���T�ڙ��}�<��G+%RhR�D�35�� L`�<��\� B��8u�/ �V����]�<!5?�@��-Ԥ[i�m��[�<����Ahx���Wi��He��[�<�2fY�Ov�hP�͏V��x���O�<	�lK_n����T(�% VK�U�<	��0/V੐vG�F���k���U�<�vk�51nn���ꐂ��LäTV�<���ެ�d"7�ʾx:�#m�U�<�Ѓd6V� eޔ^���F)D�@뷎��WFz���ߜ<��㑢(D����M�BA��fd k-А�%g:D�l:p�]�tk�I���ن�y5�:D��B�k��E�vU��F��[j�"��:D�sX�44 a��XV��T�S�&D��3���g��`B��9N�hx�V�:D��QeȾ/�I�U҆s�:H� :D��9��`�jIz���\���=D�xc/��mV���N�,�/D��3���u-����ʆmD<���/D�8�B5y��@�s� ����Fm;D�\)2@3T&���@�81�#f�#D��+b��t���D!��[p�� b!D�L�7$Z�;Dݪ$��k��hC�  D��QόR8PAf 	X_�P��`>D�H�%I�&zm��mK�D�h٤�;D��a�A�9�`@K�ꊇ:�T���.D�ܐ����	���w%\�V�T���g-D�T��m�!t�9�cސ|�<����)D�$���9�z=)��Χ|�89��B'D�����lڕ롆���Z8{bB#D�`�bGO�žܘ�`��C��*pl&D�{ �ߠQn,�K�gL�{?@��uF D����-Z�y�3�
������+D�D+b�P����iW`�zBA�צ%D��3ᄋ7��sdꖆ�v��'  D��cQ�W�)��=R�FǸw�B=J�K2D�� �4r��T/�1#�
G��8P"O|�eA������'ۦA����"O:�`�<�*��Õz,����"O~L��O�l���	���?t(L#"O�l��V�&��b�ͲHPH�	�"O�}6a�[��IP��!0Vb�i�"O`}�Cڊ]�AH���|Ip) "O:aa�#��N���%�G�=�����"O2��Ӈ��X���#��;@�"���"Ot!8�ޝ)�\*�
�����"OJ����)j+N̑3*W�]��|p"O�!�Gk��s� ����Ww����"O�H9�cգ ���1Ս�xZ�9w"OxX��y�.�(Э�	 SB�(�"OLY�`��^Ct,@1OC`�d"O��Ch�P��DyGK�~?n���"O&\�%�6_`�E�(G;j�۶"O�ͨ3/�����1���(,Ѫr"O��A��Z�YHt��gЇ8����"O�q���;�{af�N:|�[�"O�8&��VCAZ�eL�R/���"O���@c�+}&�y&D��mBD ;�"Ob|��MI�a�Y�e��}I��1"O44�5��p:���\6S6I��"O�,�舆=O԰7F\�ˊ�r�"O�0��_ŞH�v�гy�|ͳ�"ORUHQd��8��Y�r@Z�D�2�"Ox�{b��4Ɉ�� �йqv��3"O��R��0`>,����O7Ut�|��"O���D��^l� �*pLQ#"O��C�Џ�4	��Mȑt���g"OTc��	1��jqOӽPߤ��3"OL��@��C~���p �=#̩�s"O�b�X�!9V����Yy�*�"Otɫ�@��uVt�QH�&���p�"O�1Z���$�,����e�U��"Oh��Tnǣs���(�� ��l �"OB��#X�x~���ⓧ8&AAe*O�	t'W�?�Zsrʌ��x#�'׈0�u�$`�(aKRf� C�xj	�'`����0�|#S�]I�P���'�xl�P� )K2xԁ2O'SK����'�2�p�ĵ/��r J�;9�Y��'�y�e��(���9ʒ~4D��'=J��̜.c���+&τh�'���XƄK����*�0t���' lQCEu6�����*�D��'��Uz�ߧ1d�|klSr�\��'����K�;�^E�S��%�T�J>�����$4�L��k�97���'�_)�!򤔷~�bT�Ɗz�C@I�3Wa�8�'�f�+v�F2\�nehG��"#y�'��UЋ�qK�@S���:���'s��z�-T
 -�`�N�x��U��'�z��#��^L T�GI&�`�'k�B3��#�n�f#C�<^T͓J>a���II(f��PK�c�δir���ZQ!��H�@M8��GW/n���1fk��0G!�W�g��q�RM���q�6L!��ώ?Z�*��W�L���P�QT!��Z�,����@21�\Puo_�N�!��-Wt  uh.]��p�����6�!��^�:�N40d�ɿn}��� 6�'ў�G~��7k�Pp�v��,5Vx1*�dG2�y
� �����D�T@zP�G�
�����"O���`� �d Z���V�L�0"O��YuF2Ìa�����M�T��q"Oܴ���� �z�c���8j�nID"O�x
��;��ѳp��,Q��f"O�dF�ѮadѕG�8aĮ���|��)��tI�X���;;��̒S�W�DC��;������J�R�l@P'g��z8<C�I�g8$lj�·�eKP������C�I s�n�𲏜J�^�A�/�%DC䉯rU����o�rU❜o��B�	%;��BE�I�]
Db���o��B�~|#a�ɇ��e*J/U��O>�=�}��$q��p���!�¹����P�<����(^�
fD��\)EE
L�<�QM��y6qi�Nš9�X��C��E�<�l·$�x��c�X��h��D@�<Q��B�����Ĭߚ!W��R�IW|�<�@ �Zphg��+2��Q�6(�_�<��n��Gq�J2m*E�h ��K\�:z�H�?�}�sa��.��8�uvp
�D�W`�<qte̢∀��f_�b-�QP4��U�<Q�.����֜<; 8լ�x�<!��ƥJ�F�*eC�"9H��C[�<iE+خ+�T HSeK�$U.(�ׅB�<IC�2KL����>K�7G�U�<�	�n�+�S77>��*p-��o�'K���i0#����D�mJ9�%Fԓo3!�"h������ۈ�R$�]��!�D�?���ٓ%�
n�� �B�T-k!�d�>F��H%B+���C���
!��u���&L@�SrvP�GB�S!�$�E& ���%՟8���
���(!�$��,�����A����T4C�'0ў�>y��GzP��ّ�ہ ���g�,D�$�kل</��Qc+���*)�gc8D����(�"ש;��a�#7D��
��P?uj� �bS�aLހ(�4D��HA F���T:�gP�"4�hCe8D���S��&7�����B�wEv �­4D���늗2b���0�N���%-��(��|z�O���U�á	F���fA q�Pd"O��ȁ��$S��;�j�rԬ�C%"O��Af��<bi�����"O{@�%�x1i5�����6"OHS�DY?)ġ[�M��U̘p��"O8)1te��gq
��g@c�p
�"O���b���}�j���H&!�j))��|��'��Oq������3�4I��ڍ_�XiYu"O*��$2A����:tص"O�L"fiƢK>%�rą`�x��U"O^�����.�d%�0P�N��"OZ-zу��F��1oQ-u�*�#�"O��Ӷ�q$��0΅:==~�c"O��h�$��H�<�cc��u����"O�mbE�1T��s�炔-M�w"O�[r�@�kc�=����r�ƝXT"O"X�2d:i1���� yy��Y@"OZ��m%?QVa�u����"O(I��.ՂS��Mxt@-�޼jP"O�|z4.�Hb4ps$/( ��ܚ�"O���ci
z'(�pu��
����7"O�3`\�M��[�m�G�ę��"O�%� �8
BHݩ�2l���"O� ��R�(��;H ����^(d����A"O�`��
���nq�`	@�J���"O�9`�NM#�\� ���,Eǚ��@"O�<�A��y�L9��O�~��\��"O:�k�P����Ya���"OB]�#L�A�p��C�.(N��(�"OLԻ`�To���&��*�r�"Od
�IՇ��{6e�u�e�v"OP��iT�e-v��u�F7L�J�*O���@d�-�a�����X{�'&�(�˝�IP�����>�9��Y��@�Uċ��س㇘6�������p$#��[�m��>{��ȓ$e�W��bm�Xõl\;J�@"O�L�7�$��̫�@���"O���2;�v� c�-/+82#"O��Fm:r�^�Ԁ��"fx��"O��sbM�)�B��w/�q����"O0�e	|-���׮�(��a��"O�%�,���z��.��_�d��"O��Â�x"����ǡ^��"O�֨I����A挑�f%RW"O�}�!�e�$�G�6J���!"O����� 7�T<�� �{�:�0�"O�xHA'�9`���E�k�(��"O��&i�eJ��@��Z&&V� �"OX��f�A���cH�_��h�"O��s�H��_�� #,O�
�1ae"O2�@'��NM,u�תЂ:nh�"O�0�!�(5V�؅L�$�8��g"O���)���x��˄.r�$�1"O��p ��II�,�w��V7PX�t�<)#��h=�c��7L�bE�$�BQ�<�7�PIEC,v�p"B�
*���X��Eْ���pp�c-��]��Q��
?��x˱L����!��'���u6ݳ�`�g@(X�Y*Q�����1�4(PsM%M&dM�
8tM��T̀�b,a��ν4��Y�ȓzyb���Ȕ�V9v)i��='z���1_�a��HH�y�
Ք���ȓ!��3�%��'uP�qG�,2|�ȓi��c�,%EFѠ���,�\�ȓh��7�R�$R��(%����'�<�`f�8�8�B��7*�(�'u�h�C�[���chL�~��LY�'�TY��-�@����*�p��'}`!i@�f|��e	�1�B!r�'�<!�D �:?M2ݡď�&@���'R���Q��&p�*H��ǆ�*��(2�'�^<�V�^8`@2�<-�R
�'=�1K6�]�l�>�)���J���'/2��2�A�1�]���ޮ|;�'��8ՆWB���sr	�~r�J�'v�:p�Y�_!�1R1I�n��'��Q�ǫȰfԌ1��pl�Y�'=v������sY@p�@LM2o�d�
�'FjAs�F�4=RL�-O�/�8��'٠�J���(m��zBj�*0�r	�'�"\ �\�x��X�V�׺Qv�i�'�")#��]��hQ�j�*R3�#�'�^���(L����{ �W�KE�,��'���;d�=%* �3�\%
	�'�0����i{x�P��®I�	��� �=�Z�yײ�KT�֜
�0$"O�5�2�
�g����`��Y�"��4"O���蛥#���x��D45��!�"O���2%A9a�1Ǝ����|��"OT��f��h��q'�F>n<lb�"O�E1HF�*d�A��aGQP�|�W"O����nƼ-Q���E�j��d"Oh8�U�4���a�7j܍*�"O�Q@��F�@�T $/
8fXN�{�"O�{�hƢ.�@���D�[��,�a"O���CmS��Q�T�5��T�"O����I�s�a��P��A�"O<���#�3k��E��ޢ���"O|=�ulR=��P�u��"�"O�!2d(ًF`�`f͓�
$Qa�"O��87j��l0F��3�Y' T�"O(�Qݔc��u{rm�S�@m� "OP�P���
.�`�b&��ud�9"OK_9)����'�LA:�L@=�y��!A���W僔<v���O�y"�S~�|�`uE�T� Ӄ�:�y�h�l�����$Ο�`�c$ƒ�䓼hO� ?YB��:| �H��J�p*Z��DΘj�<���Ơ%vB�ʀ��IwL�3 �c�<9a�ʲ-q���Ӥш8i�E"$��_�<�'�R��hiv���p����E�b�<�0�[����*s��f	��PnRW�<rH�I��=�V�D-(�`�"L�<a'�V8bd��b�ED3��l�s�<����:ZT8a���M�̢7�q�<�@jߕ.��	a��N=K~Ax�ĕk�<���!����EčyʤTpe)Yl�<)����(�ެ�U���`y6�#S��e�<ٰn�<LZ��u�9h0@u�Kl�<�2K�<5�b��0�F?y��Y��@k�<qW�Ut��AP�ܲsg0���+�e�<9��,R�ʦ�+V��Mi0e�X�<I�.��T�A�ɥ.��ؠ��z�<	��Ź���H�K_D�鶁s�<a䨐90Ԛk�f��?������]F�<A�X�qv<̳��#[*@�u
�]�<���7i%�<�鋩=��ՙH�S�<AF��Lmn9
Ba> !�4�CřR�<���N�i��Ц���&OLm˔d�P�<�NF g�!��ƷBS�l�E �K�<��ď�Vs��bS6d�J3d��C�<����1B��)'�'>0��F �C�<� �����#���#�h��$"i�<q!ٹJ��#6"�"J?��!C�{�<���@98ʘ|�􀔞%��j��z�I���?�}��,Zb��a�T��6�4Srʟ\�<��쉯7��`��A\u(u����Y�<�1���.���	��;���fHY�<�G��3�qc0+N�bh���k�<i��ޮ)�z�RW� ,ppYT�\�<	6@J,6���5B޶;��I�	Hs�<!�E��iYS#�ip�h�lGo�<Ae��
�if��9���("�G@�<����	d��C���vX@����~�<Q�
W��%�DL²�M#V��5�y��ֶy��Hh�A��a��}B� ���y,J�<��0dQ=0�85��y���?��ࡂ��"�� ^�y�b���P�F��~e����Kɕ�y
� � Re��+2�(!�e��4�F$��*O�(�B)��v��`��rVH��'��i��Y<������p��r�'����bg+<h8b�Pe�-�'�`��-(Ğ���LH/
t���'��hZn��x�M�`Ą$k�B�:	�'29d��p��%����:,���'��ZqoQQ�f��H�)[�
ti�'��]	��ڐ8�̘ҦHҬ]/:��'(z
���=��&E]	����'����UٔB�l�+�aU�[�X�'%Ԁ P��X{��:�hUL\�́�'e��@�vc�hKǃ8�~��'`���M���|sf��zy|P�L>i���i�i�p��@IE�y�潲��]�!�Ks5숀�b[�@�F�1��q�!�Ě� `(�O�:�Jp����tm!�:���i�� ��<K4�8"k!�DR����PC�3C�0�IbB�O0!�dКV��Y�҉c~&�IQ���?'!��P�,I:�n�,)�B	�a�X�(�O�˓�����i��Ֆ6@Z�g��E=�B��'�!��
!>�tа��L4u2�h#�L�!��H	�+֥R���R��W�A!�dT�7�\�f�Đ-�4 �W��2,[!��Y/�Hr`��%j+N��L$>!�D�O��@�͚$^ ����f�!��W� 3��E�O��x��	!�䙓�zYG�Gm��ӣC,{!�T\�νh2'��>�F �#	�)1p!�$ͼ5�~�����
G"))�̼m!�|ÎD�7��O�Mq��!�d�@u�L�8"�i���Rx�Ć�`���p�ǥ�0˷��X9��_��Y8gC�3UN5��S� �b��Ddma��D�HT��ŗ�	�݇�	F�(u�ߏ(�δKHҁ���ȓ(8�P�g��iW �ېeǶg�B���-�~�aOF�.1���%O3i�J<��d�>�Y�
K� F�����_԰�ȓr� Pb�H�"���s�R��.0�ȓ�	)a�I�N�����g��$��C�����Qf��ă���JU�ȓ]��X�ь�^;tI�C坻9�\]��6�����x���3#�+~Ψ��T�d]��NQ�j���j̐����ȓJ�p5��u0�-C�]�]�ȓP��p�4�[�|<h�h��v������P�9g��?0�iX���2]� ��vQ��J���0y�  � !�H$�TF{r�'���Ӗ_���{��O�}=�-a'-@6.�BC�I�
�Jt#�U2ʄ%�@%�:�C��?�:�,��D��.QxjBB>D����K�-%<����
M!����<D�X�t�M|�ޱ�CZ�B��Ò�:D��a"×f��e % �)]�5��9D����JYs�$x�d�&S��,�b8�:�r���]�ORޔ�!�*$������B:@�ܱ
�'�	Z"!��,m��@�c�>���'A��00Y*n�R���26�|i�'���qL֪0�Д���z��
�'��s%�֜Ｔz�F�ӆXz	�'����%��	�1��	?f�Q	�'ˀ%*B�L>wb�����V�y�T���� � �� r�j��d�Z83b�x�"O�E[�*�xI	��[����Z"O4��R�C+Ɉl"h�2r��+�"O��/���e3� �?&j��(7"O(d�M�5�\s`�EMN���"OJ=(Â�7k�T���aN�=7Fe8d"OĹ�� #��Ւ@�6G���p"Oz�j�'\�0�b���/�[ʠ���"O� ��+�(UG�	�D�C���`�"OhਐG�(=ƑbūA0"��"O�B�D�p���SM� a�.�Y�"O�����33�v�Č�h�V$��"O��iЊ�	t.q��T2X�T��`"O�UH��^o&����X���RQ"O�hb�
�}��q�؊0�``2�"O�=0n�<�2f.iܶeK�"O�l	W'_�-$��)�'T *ؠ�sv"O�ⶢ�&���
�:�8�,�!���8lĜe�eo#7���$셢1�!���r�@=hF&Q�_/d��d�k!��u!D@�"�! �$�3�X5!�d�W�B�JcJ;+r��lMQ�!�ā�H�l��օ�,h:4(��y�!�K�7���7���24� �� {!�D��$�:)X�AΥm������Ũ`!�䊰LtHyy� �N�<�� ;Z!�d^�*?p�U����
�a�-K��!�d��ZC��AHK8F�ȹX�C�!�d
�J���ڳ��<���P1�� �!�H)��h���"N��qkX�F�!�D42�z\�2ŗtx!z�˱=~!�;a >mʳ�� �x��)״r{!�D��D(
v��r�����f!�)>�X�T��1�,��ӄA�n�!�D�+ ��[Q�]� °� �CC�z�!�$��J�I��@֑F���YPb	�1�!�d߃4��yP��~�P�HV`_�4�!�Ċ.�Ȱ��K̆O���w�ܶJ�!�D	�m��p69oƴ@x 邪:�!�>3�na��e]�\�����i�9!�!�X<(��<Q6�+2P�@�t�L��!�$1<�]ru��g;l���� )�!��=��D Ы�%���q�EV��!��&fR�ӆ&б"R 5h�dʊk�!�d�'��1#b,U��ԉG+Y�!��<V�Hw��?J�4Ԗ �!�$�=^�t��b��{I8�(�O�F�!�J(o�J�y҂^�*R �(P��&�!��z�lҗ�E�%DNuP"O4���2m�V�sVa�*E���p"O���� �����!ޙ-3F9B�"O���V ʭU2T	����&@d=i�"Od+���9(NrHb5ꀀ���"O�*Aj���8�DiY� ��$J3"O�$�"��T���x��Ք%yu�d"O`���J��V��0�� '<(}��"Ob�+���E"���U��$Nq�4"O�T!���% l�}�7�� ���"O�R�a�88�<�sh�:#�f� �"OΨbR��)��!#�&J�B'�Y6"O$�G"ѵ#30�ҥ�Цxn�x�"O��XD��op���3d��6"O\i�B�B<c{����(�t� 2"OD#�L�}�Q�1�H-|�La "O� �E0�a��qK8q��>�ȩ)�"O��8i�7c��آ��1U3�M��"O~Xb��i�TL
6�Ҳv����"O"�2"	�!��!�fJ�gq��"O�(�a�Ҭpr�p"��NT���R"O��	 �G"h�X�q��0=�X�"OD���C,��!�AD�}!�Ps�"O���i�&7��@E� tf�Z�"OL����ȫ$<�\s!Ǜ���+"O8���X+�i��XH��܉t"O��r#�� k��]��CU���;�"O �� �IV�!�ˇ5^��c"Oh���#&�x[K֘q2D�t"OB�Zg��N�,
T��.�`{�"O�E�CY�����ڥI�> �"Od9bÃ�#.D�f��!g�`��b"O~� R��8"1�$з;�<�W"OR(U@у;��t��W
o|"��Q"O�Q�P�2�y�m�m��e"Ovݠ���{`�拆o��0��"OBؙ�i_4~�&9����;=�z]ۂ"O츫��T�dp�O܉7���BG"O2}���C4zq��`$�����"O��;d!]��.�Ӵ
�Lndi2�"O��8�؀$ԑ�	^	p_���"ONx�eM0�؋ 	��l_T8z5"O��ڵ��]��8C�F Z|@�V"O�p(�kZ�H�8=p1fLO&��"O<��4� S��c �{Mv@ C"O:�P�(W�%�H�6aP-�%�0"OBU��MZ�xs�m�#͘x�V"O���PU��A����5Iw"OhT#҇�Ca�B�
�?�rM��"O���@�D�m��`�l��`�J�"O��
�ۊ��*ϵ	�N�	�"O��2Q� ����x�I������"O0mI�,��Q#BP����u"O��I�j	a�q.AT��DPW"OV�'�c�@��'��N$�pD"O�B-=xG��)Ū��	�"OP��_x1H]�3*۲JҔ��"O���"V�_^zԡ��ˀ ��1c"Od5�/X�Ak0���� �4��"O�e�f�*TT�*����^���"O5��L�+����J�)Ndjlk�"O��r��ۅ!w����ʦp]$9�"O`8x�m�x��%�x��40�"O@(K�)��H2B���JАtba��"O�E� )[�12��w ��]��"OL�6���laa���i�\�js"OD]�4$�kE����R�@�c�"O ��@!P�B�H��n��p��"O�5�s���\dR�n}Dl;�"O<ɪv�54U�:�#�(ۨ�D"O�9��J'��k��A�V��U�	�'�"���L՞~��8{�!��_d^�'��𔎓��T�8�F�]� ���'�h8pP��
ٶ���e͔�F�'`�'태q�4(a�)�����'ot4���1)���a*����'A.�� ����4�1�\�~et���'1H��GM6P��(!�8{�F���''t�YG��#3	8�#"��~aVj�'e�0������N�R���(��@���� ֜���G8����-0`j��E"O��pE/�&8n2ؑ��U2f0ҁ�"O�z5�8B��1��<3Vq�"O�=0E���Ey��(Aa�|6�M;"O�����;�x`���$�u�!"O�4� Hɸ)�F��pNBV��;�"Oܙ2��ӂ%�xY���K`r�!��"O���"[3�єMАr�f�G"O��G`V ;�.��FQ������"Oȹe�<F.���"�y���B�"O.D��A�>\��٩6aG�F�ڃa'D��z�ȃ$U��zQ�\�e4�����%D����@.^t��D��~ 8J��&D��K���M���(Uu�I�J#D�,��M�XWV�!ը@,fix�{ƅ D�����6/<@"#k�8�����>D��Qt�D0�X�R�[f6�yb�j7D����Ξf�
$Q�)
TA��(5D���n���)k�;,.�pj1D��ٳ�V�o�6��5�X;sؤ�.D�@ �6=TT��!ɼG�Ơ��:D�L	u��!6��� #�9¾ ��E8D��[!��,�K7�@� V��*U,5D�0���}׾y�Dm)	��pPO/D�T�� �SE��PYk!|���,D�|b��E�>�z�餩˧oPJ��3�(D�ȡ0�ݐR��#�E=d�FTh�L(D�$0F̊BC�q��k"K�� &D��w���=Tx�ā52�HC("D��0MC�����4;D�$qP��g�0�w-�.��Q��9D��9S`�,aagn�L����j$D���2��~J��D7�0`�Q�=D��s����3�T9�ĩ�@�8`  ;D���M_��,��c�=% T�!�%D�|��&v�.Q���N�*�J	�p�.D�$B�ƚ8h����k@���g,D�4K1-̧G���R���'2YT$�1D,D���T�G�nM��qs�S�8l���'D�DsЏ��-|��h!��H���'D��B�,�1�f�{F
�}ID��'!D���C၀GN�L�v��[]r � D� �U�*D�ΐ�μ��{�*O���œ�r�b�1U��6=���˰"O�y#j��cS\q!F�#q �"O�%�p�M8I�jhI���� �"O��e L�:�I
��쁥"O��� �
�6�v��2ω0y�F��"O�1"���b/���ˉ�����@"O����Oڗ7�,����2�byP�"O�!�`̥%ٶ��f�ƾp���!�"O�8ِ#��\z�C�ПZ����"O��g@�!e���W
ͬS�V-"E"OJt�S�ڼ"jB���Z�R�t ��"O��#+�mo^��H@e����5"O&�U����0�i��/�ʭcC"O.S�ٝq|t��GgW"��hR"OJe!�B�C�y;6��I� �д"O�m*�`�8Z�\t"�M�K�	�"O�S���]�4��G/#�l��"O`�* �S���XV�Έ`�H@�E"O �[�A
5!�s���ɒak�"O�,�Q�G*i�0���ʤ!�
�U"O��c��^�C�j�ذG���%��"O� �U�͇}�p�&�p����E"OT���JU�10 �h��%0Id"OP<W��!PL���O8Te�`�"O���  {a��%*ѱ|N4؀"OF4�T/^0e�*iShR�
zZ���"O���GY�,�u1�ӧAu|��"O�(�P.F aK��S��[R_
���"O�!�3e��	P��H�.���"O(��C�]c�(� �JǼ�˰"Oft��R�
|	�i����"O�QeZ 5���P�h���4���"O4`�f���~vF��$�L'	����"O|i����kѼ0����b�3�"ObQ��	9L0DA��+c*y�b"O�uS�l�1p�ҍ�S&M�&W�Y�"OX��RnB�2 P�0�2CH�+a"O.Hp6�ѳ3ީ��f
S9:�� "O� +�-�"�Ι[�l�;s�p�f"Of�)%MI�@��T���Ql�t��"O�]�Q,+��d�2���`���Q"ONE�W�ʻG���Q��B�8!8"O���	�5S5�ՉVdš/����"OD��$�3�~��A�L��N��P"O.�:G� H�H1��g����q"O�i�_�uʸ52f��$]�B=�"O4��p� -#�BE�qo2�Vak�"O����#��~3eA��X)i�$U�"O��х`�.�`��%h^�T ��u"O8�`f�1\��I
L`I��"O��E�YTb|p  Ι0B�<0�'}�`���� b�q�v��c{�!�
�'<ѓ�)Q,n����B�T�*�	�'!j��Rl4Z��@Wd�D��(�'	H|���D=������80`��'��P���*��a�>,,@��'_rP�-V#@�s��(�(��'y4��Sg�Yö�ȅʔ.v1+�'�p`��!˖e>�@��0I�JP��'(D#��.��7�����'7n��#�1RN��W�	&�hc�'�$H���]i�hK�,K&,��h
�'S�=)��Yi����ڛ̀U
�'b^I(��8��|#mOh۴ݚ	�'�f��gI�(<��誃�s�L���'C�LBV$+�PhkS�"s�RD��'��IF�Z0]n�<@�(�"��|!�'� �Àl�0�aÔR�4���X�<��D�=��I�,
�/N(���IY�<���M0A��r`׽-f��ҋU�<!�KX7*�J(`�D; ��x�6��y�<1v�'PH�(���A�v�@	p��s�<a�� )d��r�ʲP�8$A�Oq�<�ց��X�B��)v�b�c&�i�<qĐ���҆�B#-!2���K�g�<�'���:P��
�-Ǻ�(��Rc�<��m�9O5���E��&�`�F\I�<I	�/FA����A�)r�D`bnJn�<y7�˾��8x�cN	Q�Pڶ�GS�<q�iJ�7��h����1k���yQ͉R�<i ��0�JI3Bj�&>�r���Fx�<�hYU��u)��N"����j�y�<�ˈ�>�zF@.�9�A��{�<���p��m�"�ϖ<��`��l�t�<!�D�T���#F��p�AăUx�<� �-���K�8�yBi�^Ut!Rc"O6���j��ja���I�E��!��"O��#֦
"�,�ʳgW�g)�UR`"O�4�T`�1yʝ��EїI�u��"O�`�`�F=z��ṅ�"a���#"O�S6#��n�v`Z6&]�Y]PLJ�"O��qA�"*`�kw�P�)g��i�"O�Eb%�ŁH���r矅3e| )0"O0���eE>/851��L4V��a"O�d�a'(v sGE	�1��=�e"Ob��@%D�#eb��儹R�J5y "O(0��%�"e�rx�C�ΏMz�@�"On�Q�ED�>�0E�7�L�P�i��"ORx���G-m��I;v*9��A"O�4��#�<q�B�z�K�@b��U"O�st�z��)��%��/�y��)\"�[��2W�4i;Ҩ���yB%�9Z��0�̖3T�H�D��y�H�Dh(�dY0H]�����D��y"I���AÖB;F-���jس�yb@�=6����D%?�<�"#fL��y2,߱~β�����>�09藯��yR��X��0��IU,>�̡'����y��YR�t���/M(X3��<�yRK,�`9hѥ�8ZP�a�<�y2\'7䖔���	�*ũg霱�y��9i ��iAl��p7H� �y�HŔ/�l�)6B
�yj�P0V��y��̰L.���� v�*�p�
��y�����J �C�����"Ǥ�y�
B&I �K�:)d4,�ѩ�yb� dfԺ��A5'�.�s��y2�J�� �A�lA�oa�a���y�nܙ����d�^ m��8ZcL_?�y��8֮�[�i��a�D�CC�M��yB���[�J�rHZ�\~�J����yRJ9L�,lp �L,G�y��NR��y�lV�E�l�ZW��Aϐ���h?�y��ٴ0��b3�9L:l��`4�y�B�\|�8���$~�^A���Y��y�ν%�9���Au>J�BM�7�y�)�?~���ɗa�ޢ1�Ԧ�y�mE$���ɣM��?�A���y��]J1��`d1~�\�"&O]��y2!ޯ!e&	��f�m�H�ۢ� �yb��}��$�g��ը"O����^(�|��dƳYK���r"O�DSEC3����p/��K@vA:W"O�����\�AFR(�h,=&H�)GOL�H�$٬rw��{�k�4IRp�W�C+9!��Z�Qrn4�G�K80�H	���Z�!��Ybo�@��վ0��`EI�k�!��զ>�������$���i�!��ϫx��e�X�[�d��`2#�!�$�-pP�rsE�c�4�YCo\�(i!�$����V:���䃭Rc!�ΑyT�4����2$��LR䢟3e!�$зy�0�Jq�I,J��8��O�N^!��I�Tw��§)ު��	@�/U�V!��'vRt��/����L餯�>v�1O��Dƞ?�2Q��M�*ŀE:�� �;�!�O�P���g����-�3"�x��O ��Kkx��B隺~�~��po�J]ax2�I��.]��
�,��-��/�����D2�)� HۓG@�@���J��J	w��2"O&�Ԃޮ9cJt �J��V�tDpA"O�`�:���EI��gv��;��'�ў"~���
KЬ��W-�De�d������'U�{B��,(@�9���6;�������y�A�<I���kE�67��H�8�y҃T Z�l�)d�1G-*��s�^.�M��'붡Fybh;��kVy�a�H�(�I7`�;fe����<iփQ3C\��"���f~�k7�CP?�F2�S�O�JD��7A|-`A��|K�5*��D"�R�⤆	7u�8X��ѿ2���"O␚,�!�iXP��<֒����'�ў"~
΋<,p���ψ.~Q�ܩ�G�+�Px��
Ⱦ�I7�#/���C�
O�}�tYmZh~�9O"�i>q�n�I�jU[���:������ֹ���Y �Od�B�vT|���l UbE��"ON��qk	�~Q
!�e��kUTu�w�>��>�S�'h&�h�4� M���z6��D$�͓���@���!���PK�Ę�S�Hk�-!�I'eAazB�9��]�I_���1�8��x��0/D�EsA�X�=�j�3Ai>���=Aד}�=K ��:��=+!͌vs�ik�H��+%�<��b/2:d���J�N�Y�G�6@dI����Q%�?!��qyr˟���K��I'X$t�0P���'��z�'�`@=R�I��I�n�p�0�HO��/U��Y��œ�J�$�J��A=�C䉽�����b�!.
�v�ӱ/�4O���h�%Uq��y`�hM �R1ꁧ��m����V"O����L�%V����d�v@W"O�yp`���0�(i	���9g�nt�"O\s��S�tkXe�w�4v|iI�"O�p��$��+J�Zw��M�<m+�"O"Tئ�ٍ0svQ����3	w����"O�"��Gl��9�żk�ј�"O��*'f]"U��l��+ھe/�+d"O|`�b�OJNl���"-|�A�"O8�4l��6g�}葌�	<���"O>�Wl� f�"��=AvB��'�!���#A��t1�Ũe����a�!H!��*�t�$DFۜ �ů�ya}�߯?�B�@�r�K�-��y��o�;'���p?ɤ�ۘ-��9��
�b���1�f|�<�`G*A�(�[E��4��%نL�!��'?ô�S��\%W����Ԫц,la{���-ge�I2����Ffju��J�Od�U��<ˑo�"%��Gg�S�2��*D�4�!�W@���e�Ȑ���@$D�L���
�Q�C�D�A 𴨂�#D��*��ԒZ5z4��>z}�p�A
"���➔��I�(E��Ì�rX��$V�*�M��Z�4��5.�'6˨ ��ᅎ�����8���@e��nƂ� ���kr)���?1g�9�4LC���q�L01��R�<�I_1\���`�DC�o��Ƞ�	�f�<����1h��G/kaT����]d~rV��F{ʟЀ`�NU�P��ib��gp2���"O~�RJ[.<GH�{mj���"O�q���} 1��' ��\�C���u}R�S<|�r��4�6��ō�A�'C��F8�T��*�s�tJ��؏)C��StH0ʓ�hO�S?�R��q�F�T�	q�gŮ4�>B�I�Z����&�Z0�5k�N8Syb�O����G���IÁ	�h�����\ar��ߟ� |��n�?�5RqӓV�4��?O.���LW���``�V�p0�9�6�P;<�!�$�o�T=��Q�&����MS��D:�O�7�r�$��̜֠O?0�ӡ�'����q��0b�G��`����\�!�Ûh������i���xҀܟP ��&���jA�@A�����瑙�,]�ȓ=~��J�I��x���t�r4�(�'a"=E���Y��"�۔ 
P�
�JBF +�0<A�<�O��p���h�<����!j������=D��Gkƒ"@��K� [0(Ĉ0@�7�OL�IqB�(�B`%����H�fC�I"+��#�X��)��0m\c�̳�)�\�;*����'=X��rf���[I!��] #tRH���f��:q�D�`|��U�	%yHax¯�'=�n��碁D�T��e�Ԯ�yRa��C,�W�A�A ���X��HO����٘.�8�9��[P���{� �!�Ď6%��R�M��-2�c�)>�!��Ķl�0�z6EY�J��<��d@�[���0F���Z�W8�iUȓ�l,�];�$�2�y��G�ה�@'G+z�.�	����y2mF�m��AЃ��wE()��.\���>����~��Ŧp�D r���-pa|]yg����y(�4C�޸!ag�Q���j�`��y���I������M9bѣ��#�y�@�&-�LɉG��E�P[� QeYў���i��4GE�n���Y��ЍV�ZX[B�"��ȟ�i���/�|PH�DU�#"���"O�$�Խ$A���/uh�s�Of��&�� ]�T����*٘DpTO[}r�';�x,L�g?@Db��,�Ҭ�
�':I���h��Q���ƴ 	ۓ��'��Rw��e�)���_����ۍy��)�S_Dt �Q��?c�ƈK4�A=	*B�I�w��u�+�!EH�|�CG�."x*B�I��F���ߊ$�:��F�r!��hO>�rf�Ҏ�����#9"@�Tg"�$�>�˓;�c�f�s����`@�5�Nl��>�p��F��!SbP����1�JA��1jB䐔��.C�eZ�c��+̪��O�'�L q��U�:p�pe�d��ǡ/LO"�  FG�*M)X�qF�)K��-D����O�#vh]���H­Qj,D�;�Ե}t�`�F&J^�p�&D�l�#���H�q�Ȥ	�8����2D�p+�#=;�l�ŋ�T�ʴ���$D�0�u�ކwJ��5�EkE��e�#D�LX��M	`s&�_<5���"D��ʥ�._D��QE�B5?A03cH D�0(��E�v�����TJ0���3D��Z1ᗺz���G��]H��6D�ʓK"rD6q��\��!u�0D� #�Y�(��m���Y,&�`t�3D��
eOW&E��X�
$*��D���0D�X8��ǂr��EK�<C��d�2�1D��˷nY�ߺ��`�W3O�p)���=D�8y78B�J�b �3�|)U�<D� W�] �B�{�%��U����;D�tˀq洑���Sr"��#l9D�@r�Ā-H{�h���I82��V�5D���aG�~j�|��\J�B&D�!���<"��X�%�c�<$��$D��l�Q��@���b�h豔	"D�� $e��,�
h���J9z, H*�"O&0%I��.���`��$^�ð"O��	�J�q��88�C�8�!;e"O�e�P��i�L�rg�T/$�k%"O�)���{9�}9��-DK@cs"O�����Ի>�����b�����d"O U1u@�/;�$�q�9	�4�C"Ol�a��� ,���yt`�~��y*#"O�m�AƉ=9���k��Uk�P���"O��P�Z�1�H1IR�֨J�`��u"O�LxG��
ˌ��r.C��pLp#"O� 1��A�5ȖH�0�Gq_�=�b"OD���/D�L���s �%~��	��"OPա���:]��9�UNݏ���B�"O\<RT,;=MtxڀK�45���s�"Ox��#A��"��5*¤�Hk�1�U"O�M��I�$u譣�W�&`���e"Of=���$C��hPrH�5sF��K�?O�uJ4jI�"��aK���>�x�e��?�"P�v��1?������gE�C�%HVm����� I�D�87�B�I�$�&�eH���������^C�I�#!�xk�E�|G�( Bᜭ!��C�I�l�P�Θl(�ăw	��+z�C�ɢ)�P	a�%�*7�P�Å'�2
�C�I$?2�t���Q�]�Fm��Á0 2C�/lZ����1EVu:AAPx�|B䉅|���i#�G�O��]*૏*(�B�ɋΈ4�%�_9*O���' Eq�C�	�^P��Z��×W����&�)�B�ɔJ �	��"�4^����'$�h�B�ɪE��e;� �!=z�|1w��9h|�B�	#]1.�J�'���xs�GH�lB��DXb�K0L�ܑ�C�I�B�I�\� ��ީ+9�����%�(B䉟r��p�GM�_�Xp1��כM	TB�	OUA�Rw�}��W�uv�B�	(ݬxs�Ɋ� ڥ�0I�/��B�	!�&��7,ýb��ձ�)B��fB䉋0U���� &n��,bWlߩ�l��;,�\�'��Dd�����װ(2e�V���shC≦)4�t-.I�"�1q�uF�=�逊L� Q���5��O�8�y�`U���E���@�"�x�R�'֘$A¨�7=����A�;���4$Je���9QWx(��B��"~nZ�T��AE)�*?�HH�ą��B�	&u�z����/͐� ��V<iZ��:���ز쉏��8A5��?�=q���IKFpq�&Ԅt"0
��`��HXbáS&�,2!��	�� q�U��*���_+ZA6�����V�a�䀺��3�
=K.������'���t�A%��W�Qh�xR�<��N�."9
t:�)	Hp�"Q(@��y�j�$9�a$��LM~�`�X��Y�� P�C��I�T����ٙM?��I-�1��':�"fl���@c��'��'���@+c/0��p ٭m� �(���%�C>���H�	$Wre�A�_ M-6�G}�;E��H�C �+���������HOz�,�#Ag��9 dUcz|�cƁ�1����, � �D�!�M
'�%����"j�� 2$�y!t� �%�	g�r����Ⱦ �*���F r� y�H�*���3r|�f`Gl�b�h��b/	�%�$��7]?���A*�A6��l�cb��9�剘Jx ���p��S�O�� c�#N����i�R�&�Ss�9�@D
	��)������$YP\�4o�(]��ɳ��8��#A�أ���'L�1�AZ� 	0��Hg�$�O|n��>;*��^��֐a2����d��Z��Q��י%4�e�� �L-D��P!�t�IR�dȺ\gkLߨu�2��6?��֨ bT�bw���B2��@��bU��?U�py�G�X��r�,@(W�>���
��G�ra�T��;6�j$���W�[���a���H7~�k�[��*�GѯXP6���N�/K���h%'�-��=�@�E*Fe&���jV3UyX츢�ہ#N�:��î	�~=CU��/��5訟�n��k�J�@���&�n�*��05��f��Ab���W�cO�~r�S�S�D�r7$���`�TR�#�,DTJX���]�t 8y���"?���E�m��i
�O RjPcʯB[Pl�&��'r9� ��b����0��mP6!�~к`�gmL/e=���gB康-ʄ���z�á<�K�,�I3c��[�& ���v>�`/Ĵ,���k0���Re	��b`LK�]�&<�vC� �A��i�uiv���e�T��MW�kC�M]ފ`�F��+��9�TU�p3V`$�,r&dR��0:s$V5g
J�)�A�2&�ؠS��5IĽ�rÔ4�X c���&>@Dݩ/1D�P�υ�&�ր�@�%3E�7MF)����D�l��� }K�8H�E��8q�pXtkV^���g��P_�Ry�X�뗝Y	��ɗ���wILx���R�I��
t-:	 ,Q��R�
�
T��݆|
��Y��w$��`��D�E��@�ڼ��	�[��-qEАu�A�����,���E�`]-Y�[�l*��'[��51�}�}�6"@�)��3t� �K*F���Z6�	B�t���Ġ)�B�1%�8f*�`䯁���G�
斉�w�=TYj �t	L�q���F5ڗ�դf�p�� �AJy��#~Je��׍qx�aDT��P�7��& ��Iu��j8�Bd�	o0� ��YP@D���#?&��2;��Ȗ���ZA�\��F�b��$�3��/Z��v�9>�:��[s��,���iKZ��:H�R$��2>��XٷD����ꄐ����w'z�#����>y���k�2�t�G�3^��q��)�h ��M N#r�;��L��ϿK oG S0�}���]yÈ�B�C��d,@�Cޅ���g��2(}.x�'R3�a�0��Β8����<�.W�)���A$χ+>���qJ�N�tY��ˋ�D�v����^�����O]�,��4)8����*KI�je1��$���.���G�36!��N��� �R�@�y�,����S�ql1O.���Ó#po�0��[�2�N�2��~�,p@F�#�?!S΄����e�K�=*�N�A�b��3���0_}
̓R�C#L�����πQ�@�i$Oж@V(�D���'�"Y(&�[W�OqLX�[�������_�uA4!G�$K6�8���s�u3�D yBx�ģ���������?1�wF�E	�b�*�X��p�H�9q
�'�TY�]�s� �j@e�5�ѸF�ԧ/|ԝQ'L.U��
��[m�VQ�B��p�.�*�_.3����V���S��5e�4�3+K�B0���Ɇ1	�Њ��Ek.p���+	a:�C`L�)�n5(0Ǖ4no����F�8�������xHm���K)l� �?Ѯ��M��k4���9�ɶj0������L����#J��]����N�-J����	�|�$�ސE�1�w��:eJ��� ���N��	��	$D6�b�GN�0��p��e�{�ja
�c��Cu��H��W�\�WM&G>�:4'��M��#����λ6���E�� �F|!4e�#�V1��^,�� F����@T.���U�I�l�X�-�		�Z���j�^.��@�&P ���0씍-�����ib��h���6t$�2 BI�ly��Q	�;J@$5;���P�dǂ)t�M]$���e���+$�"��V�F��a��X�d]؂� � `!rD�I�mȎ�\�� b�8g[Nc�(R��:bPTa�6�3R��� �J�&+¨K6��kŔ�B���hMXY�M��g�$%��*^of�)1FJ6�q�l��RD�	x�����WZ��b��eǪi�2� �)�`a��D_(X|c�웕+�$��WH��բĵcͺu��@�*�r59��<T�(�A���:b����	�(۸'��ٴT-w�"t�Ϊg���T,�MZB��'Y �:��&6٦k�
��`L����.T iz�
�C�p	9 ��X �E�$3Ӵ,S�V�jx�%�iK�((։A0T7pjG	;n���{���`�k%�G u���f��8N�$8ƹ�R��q(��&�-��A;��{������AfJU"#KG6��3����V��8ժ��T[A��9P��lDy��Ĩ)b�X�	�<f�!Il�cF�Ұ"D��	�3��v�2Fĩ)f�@�	ܢ;k�9�L�?U(/]�T8�Mi�Fӎ_ �CDʘ�7n (笤J���*5�z�B�, 3GLڸ��n�G:q��E��}8X1(a	A-u �����}T�h��#��:��Q�@	>}�w�m�� ����E($��MHIP`G&]���s��B�G0��a�x�MV�plK���+&Ș����pUHǶu%Ɓ*�  *O�j��PfU�a@A�e�I�w��I<
dXUrp�T�]�rG�ګL�dٓ�%bDI�E�I+u�����<�ᧀ9<}���v]F���Ar�0�R{�d\ �%D�
�9�G�; ,]��뇇tTV�� JJq�q�]%Y�S�@�>����D�6����	1F�dã�0YIBe���d���5�qhĸwԘɱ@� !$��J���L���̘� ��-������;~İ��iCH���t{>d"T�K�O�2)�r뙩rQ|�I�#�CG� E{"��?OB���
��}���Hї{>��qF��"���a�@0�d�Waҫi.�zbj	�/�1	t��{:�ڱ��&��҂AZ�E<�L�ס�G ���5��0h9t8��B��OvZ�H@�� �`�aa�� d�b�(p+ĵ	��K�p�4��d�	v&�PC�1մm��i�nYX!�$�?!6Z�i� ]8e��%�Dr�y����� ���N3�j���,�WC|�A��KE����G).�h�h5���� �4D��	�~��⌇ӿ�am>E����o�3vh����|լ��8=��3'��а<�H�M���S�N��C��˦�N,��l�3������G��dҁm�O�����ٙH��o�L8�� �I�."��P�PN�C��e��a\v���A��E�fa�p
��B".��/�\@�� ©Qf�%��?Cā�b�E0�"Fݳ���C�\()�Bx� �O�13 ͐�:Oҩ��-E.!��#H�^���T�ϩJ��O���EO(M��rh��=�
D�5�Z�NR�����_�#��˥n�@Ξ-���[�S�[�bH9�M;(X3e2x�	"x�\i7\�F��){f��w�T���g[&Jvt���C	2	V��h�^�q�U¤ָM:�0��ϏV��3���'N~d����	3V��̻&}JE��L7@<�h���L�A�ix�'ԕ�$PCD��>M���$��y��;���}_��	��O����GL�;p����'ŝ���q�ALx����=yQ��m����d�<�P����]H�t���.U��{�$�'>���j%�?�`\�򁋤Vʀ�&̝73���F�-�L*P�Lo�ʱ8sc0�nL���K$V̌�F�\�24��(cL��.����ƪsGi�f����R��7鉾H���iQ�ո"��|��ّ�b�<b�����
�7_@`�3�#���{�JN�+�(	z�eĶ8�4j��=f��誒� 6]�$�
c}r�U.
+�M�v�U'&�!�E���?��b[�m�X}�I�����7
�@���Ų@�F�A1ǂ+\�5`r˗�Z�&!��`���$�v�����sv�I����m��%H��� �� (�&L2�B&P)9<�����'��Tx�D�f���s��)
ֺ�*�'O:�rV�(:9����-�-�J��풠Z��\Ȁ�'�Ai�I�	2�&�u�'�>0×)ʏh��Q�q�2��ЍU�ɋde4IĤР�(�������}�bc&gYn�J$� 
�t�19_���ٳ9��H�	h����A�%��R2�b�`ŌY�2v���T�st�a F�TĈ�у��c\��1�V�v�5,X�:x���T<td����'����.Œ1a9E^(������.
����A.Đ5MQ���&�� hΟ\X8˕��7�|��U
�$:z���eD�Xt�!0��9]��e�`��TJ�U�'X�%{�O
k8P}RD�{��|��ᛳC����&C��qJ����%\�5c��
n3JI:���M��µ:@J	%TS � �d�x�����E�T�*Q�P�ֽ�w��#�%ӣ)�5]�|�Su�y��а�bX1?��A�l=T�΍����'�!�c	�7Y�n��;E��]����* ��V�4D��ȅ�	4cҮjf��!Gմ����>I�TX����hr���L�+N�dE4����`���ج҂��O�Nt�poYm|��!�M�P���)o����Ҁ�
N\P���6�K=����ǒUӶɻw��1���D�^����S蔢*rX��,�*d����"��:�P	Rb�'Ǫ�"�i�,7!�<�èU��hO>0���,�%�*�$QH|I�$��c����H�aR%�֗JO(X�L�+��T�ѧTBli���e� �+c,K�I/���v�X/n>���A�<6μ���8�O� ��Z25�hq��̫76�	�F�"
�;�)��PuƸz#��h� �02�haU�(0"�I!6��)���c��@C�EX��'�2�.�z���'A75N����Y'0�`!b�uzDa�'�p�qg�u���@��V�
r�Fp�V�)��$�0d����M>~%�؋"��o�Q�(�v�4l���p�?}"��ˢ��k�r!0#�Y)Hk&-�Qi�:"��#o�'x������R�s�b�;4�i���+ͨO쭸C�I�A�(}�v��?wFY��ƞ�:��0(dn�k����T_f�����H B�&]����}Pm�5�_�?�>�%GӬ7��}c&J�!	of�PpECQp0�F}�HY7g��&�3Q�>�~)��	q�8�I2G���S��$f�ܡ�G�iȔ4[��P�;�t�fI�t� �hޥF�ݡߚ�s��*gx�x�$
)}� E�U���	TR��"�2�Z�*�ur�ѕ��	E� �K�g�|�R��]�`�h�H1�&��K�+b��5��@�4� I���NdlH��� (n4蓯H� *�Y�d�<���O?  ��h7��Q8dz�G��c�`��p(��$H Ȕ�� �'����ᕜN�Tx�L؝ۦ�-*`����jg�'r< �ʅ|�X��ůƽH�9�JͼlϢ@�I�Y�j���D1k����VLK�y�B��Uχ?M�%��*�?j´h��鑎]��a��#Ph��R���!Q���J���OZ%�PIG�ؘ-�%%���)�y��@�D[���:��ˊ&�|4�׎
RD����+��H��G#~�� ������J� ��nV�p����5E�P�`��-Z��ɗ-�5*j�3�x�:��H��nZ�j��tGR��fU�@E.)��O�	�
p)��^�vcP�9T$R�(�@M�����u��1JGFH8�B��Dq�#�?I�L�"a#\A�
Kse����%��D0:�U�(��F
�[V��ͧa VYڂjJ�wh�����[��J:5j�}�JP���G��0�2F�V�Np���E�[�(d $�ъQafU�_�㞠(��Պ*��	bGl�(.��9�wc*/��b)��p�B���"~3���"�'��ZG��)+���C��#��`�i�!tR��5l�1 ��v��	\ӄ�Y��#"�<扞X��,s�a"o���x`!@�L\��UGؖS��e*cƁ(\2.���j�oz�U)%�ܤ6l
����ӎ�����Y�T��Ir�F@*Y;:ՠ���kr�u��!5�A���,��Feד*Q��_�l��ɷ,��|ɂ��,���m�O��X��۟�ܐ�[3�Ȝ{�HX=֜Q9剙4��������#-�S�rO۲�ƄS��9߈yiu�X�6��7-B9.p
8%曥.nP��H�=B6��b��Qg�y�r�Ę ���#��?��MR4(�4 �/�	'�Q��b��].	�)Q�8�\���k�;/.���A��o����?����B��_ c���"۩[7�A��敼i|81��C"2��,"bC�`Nճ&�ǒ �. b#H��'<�y�q��hp<`M¢2��0R��d��Ba�U�XPE�"t����G�)�%NI��'�"פ8,��	�C�7*8�e�P�V�x�:a��[�ip�T��$��Rp�؇�Rf�!�V�I+L��a5�{�>Y���Z0lz�t��D�Rt�З.C"!
t$�g)���°���^��ɥqFl;���=r�ڠ�HC�m2�g�4+�H�+�0��A�p����kͯ\��
"���B�
�Y��Y���؂a�/#�4ɕO�v�B�KǗ7�� λa��O��"�b!���d_2 2FAA�~j�M�dj�#�%����b|�c��!a�Ck7T ���-ǇFF�I� 2�N�y�o�b\(�ў`A� Sk���Oh� ���yY�y�JO!SƎU����m�����7A�� ���O�����J�xZ�I(fͶlR mM�PH��+;NZN�K�J$����^�Q��˙�L^H�C��]:W�$aܴnw�E�P�8j&��6��2����7"����Ƣ�<hft��)O�\��c[
t����1g�5@��Q��?���$���&�͠z��`��6��V�rBj޺d��:��8�Pɏ�nT-��͍�'��]�bd�ć
�6��y�Ʀ����/&�� �)ƋJ���,�*3i��r����Pb�XeVX�yS�W�U=a��)?s����	J� ��P!ά��	MR�q��sb�Ќ��V*Q_<��E��#x�@-c���`h�-O�U�,�&��1$>c��Y�X4��2ost�AbÃ���RN�F���UGր3?�(�a���L(����`�_w`	��I2~�Bg����0�N��)�>��Dܩ/f(؋yB ؍%�2�k�Aҙ3rV�;��O��y�M�
U´+��/��[3 (�y�č	پL2��@%KC��B��y�i^����,'(��%=�y
� �}��Ǵcقq��ᒗ~ҁ�b"O��x�\:P\6x�7`@6a����"O�1�C�)eؤY�/BXdM+�"O� ���)C�`1��4�p"O����A&Gm��v*ƤFP�3�"OzD�%��-�,�"�+��b�@�Sv"O��W��$��;ŬS{���cT"OL԰PG�6���ⵄ�0��1�"O��Ca�N�s?z�)�霕:*�}#�"O&9�S-��^�8��J;Dz���f"O��4�.?�0�bH��2;�"O�p�	�_004b�i�!� ��"O�lK0JA�*/,�a����{6��`"O>���ť�(��%�U.Q@��%"O��kү�9<l��̒?F&xw"O�9Х�L�6���
ӫXG���"OTT:��;$_�EЗ�S�NK.u"�"O �q�A�Spe�p'�nv!�S"O��'��:9lܼ!��%�X+�"OP][ ��[�t�7έd�6�""O|p(�A�_�@��ȹb�P��5"O�	i��U�8�R��܅�8�B�"O�|�#�$DȀ��f�P�~�2"Ormˑ��> 8Q���&��%"O�����),� ����2F5$�5"O����H��qk7H�ht� ��"O��*�Nk�ݰe)܀}cNE�"O,�˓J�j���B��EY޵P"OZppPDJ{����;(g� JP"Ora�di��G���B�n1!!"O�4��nȣ1;vx2"�&Z0q�"O`H;Q�S�4RrREX7�pj"O��� ��'{�Ѣ�B�b	TI8P"Oh�p��|�X�k� ���uR�"O�k#��~������EJʭk"O���&)�\������|;T�R"O��Ӏ�۽D���`l'��	#�"O&ء��;)f�*�� ���"O�ҳ-��12Y�dD�M�xI��"Oʥ�u��/gyD�b�-̈]Ȯ}�"OX� eF�({�Hsn�6M|��W"O��Y@�P;1�X�0��w�PA�"O���ҧʮv+��M+y���V�'����˟_;�ݢ(�&i�~�S0�Ȁ/�b%�O�-
ėX��PA%D�^��Ѓ�I�h���UgּF2PT�|��+��s5�e!����Sb��h�n�<!��G�v}{�/�;�e��fצ�XB� m���1'ݵ���s�̡I��	/od	���%{W��6"OhYu�e/.Ea��[);7�ӷ��埤A�b%.����:h�퉇Y���PT��A���{�Pc������3BK��ScaצcN��b_�>�*�ǫs<t��e���<*�����	���� aW�P0�	Y��Q��0� �6=:I�'A��F�j���~��*�z�Ҧ� '?�s�O�e�<W�[�a$4 ����hV B�pv�MY��8�mpq(K�b"���fT�@�Q����'�� ��׬��I�aMbJ�M�
�bH�A�r�ϒ)� i�#D�=�t�R�c��'�z�@RNR�f=D���c2��Ɗ'�"E}�Ǎd
�薞@F��qK�3�HO��`�C3	 �e@TkO "�����h�`0pCr��G��R����|2�)�"�ʑY$i-ғIj!��/�I;���iZJ�T�4cN2F���+0�ِc��9��DJ4O1�,{�+[9��)yɛB�@o�~�* $�5��
#�N\����Hn˓(�L"A�«*-nҧ(��� �@	�u����UǦ;��ȍp��G�J�H(Z�`��"��I�[�uq�� `��+����dJ�H��" 6����<)始��&L�G���4.4`����#z!�آ���m�dA�+��Q'�H�K��`�����p@I��4־��Q(&�ɵ.on �q#yƮ1��mS� Tr�:�X$�,Ш7lڳ|��	1M�y���7b�M�C�
�B��0@�y��o9� ���#U9ub���$2k�9[7n]0>8T�[f�. MXL�'���`N��t�� Ya�LZ����8%d��QUM�7M�
�"�Րm~X�k�fؙS�Q�dM� `\��GU�&c��i5�ѶL���3P ()��y��B�e��s��U�<��h��8"`T6�2u�P�8��>�Q���|Ƅ���
d>Q
�h �S�rA�S�Gz`!�犉� �4�@ѫ�(�3TW |���R�"�.�>Awp��JI$"�(�r΀+��1N6�.��m�!(!��	�v�D���OѴ=�BB�@y2�B�MD(i�&h�<3R�`�W�;2��p&�i���a����f6@�y mU�<�~��E`\.%qlt#���Ц��G��l�w]�_��Mc7�J'��ƅ�,�[��˓U�Ҥ�R�;=�t)˶�����*�\�����)C������.�@��"+�َ���
k��@�"�ğ/�@髀-(G�ൈV+�Ħ���5���؈��P��Ab+<�x�e�΅��J	�% `H��dY`8�)��<�T��M�L�d� ���2��KV���!N�H�L(���و��M�X�䌁���z`A_ͼ�Si*q�H���+b���
�Ř��?-�.m�*�B�
J�4]�ՐK>I��ʪ0T������(rH��U�	�}I�������<53 �:]������ (^�5JA�1wX��-OzQ���N��1(Nͣ2��I��S�8L$� '��p��(
C�>�dEr�� R�,�.�&ɳ��cxF@X�� 4�L���!ȰX���h�c�Vc�iY����/����:?��j��W:8q��_�Nxb>e��@�\5>HH7mW,t`�ԙ�e�+�0��CBr�l��N�-R�T�B�	�Y=.��m�n��7���C3;\�9�K�p�"1�r�A�Kh<0��e�"L�11G��+v���O�s��
�D8��2�lD;%M����ɳ3!�p �c�N�R��\B��F?��j��#@��54O~l"b �mN���+��5F��b�V�lc�%V�Z�޹�V{ܓz��I��\���(�M�"��S�	�f��f��>L�"�{���;	��
fon����"�Io����mB;:�nU�Cf���a�%�A�Y���� զ�	��S�7>��%���?�| "��[R�0����6x���a�P-{2��A�-���n}�����Z���I��iY!�8��A|��yW� 	W�9�M�d��x1GʛqhB5��e�%� �y&��{��i��	U��ɬK�<��&O�fc$a�E^�xN!�$�J�1�P�Id5 ��Y1=x���,U0�J�d���5�c F�B�Aa�(Aph
���~��2j�%X�
�S����bQ��p=��k dap�Ԫ^8ð�z��~L*Ф�0:Bh8��.3#�=���N��!���t��*�?���p%�0`��ЛA���BR@��<�a@�*AZR͋p�K,^�%S��O>	j�jT�T<	����h3oĸ3p��6z���ƿX�(��K���>�B˩j�3�L�j����i�=J"���v�P;�t@��*��x��B��o�c1�i�B�#ϓ��yG@�-Mʄ�v古lc��Z�E��y2��,_�d*%a�8g54U�*�۞���&Q�Kf��:�l0�0���/W�HB��O:b=:I�s*F�ъ6�ע[�l���sPDr��O?�azb��� 6��"��~��:em��p�6e�1A�q� >״(
 A��e[8}@Ӥ�;`-��M
#f"=	�
�ʠ�ThL�P�n�X1IVV̓Q�d��)F��� ѬM��0aՊ��tMQ���(��L[+Rn��͘b`�������
� �,�����)4j��.��h�TDZ�e�P��Mɧq��(0#�@5LM��1���ݞ`Z7M�4�d�4D[`�h�A�Ȥt��< 3I�4HD��ID�F9g����ڋ��k&{�t�9Ѧ��;6�5{g�t�Zh�P�3l��S�Y��@SSA�;ذ���}�r�╩̷2��c @O����)֪Y��\�9
Ę�M�x�h���4]�@�c�V�&�(�x��3,3���%�� >�b�@,B
%i(�B�O�_�F�[w$���"i�e,J�8�x�+ȁ���y�O��>ƅ�!j��\�!��%��c]�`p�q�����UDybI� z���jr�ނ\$��uJ-*���W�X,'S�5�ɐY��в��!{���rR��[)�(Ʌj�?�[C�Dv��	����еi��5+$� �'��*�2�<��C�����5i��1#4�@4&W {�z��cFN!}]�i����+!nt	�w����K�(��d�ͮ��[w}�˂��=/�TY��@�(�V�O/�f��4�؁h�l�$��"G������%U�&u�����-w��5k�m\�U@�RMB�2�`�c/�cSNe �'�.D��j�:���f%�by@�j$��$1�j��SOMbQLmƇ�G�ҡ�;yБ;�ܽT��m;f�Z�G,(�Sg:f���u���f�jt��8|؉��ݿP��q!��5v�Y�壀#[�9^�9f��x3D���E�?0�E�#�b�pe�g��}\�#=��H��LHs1 �+~�"5�3�ђ}������D�	0���j��?�%�'�.�Z|���)z�$%nZ#$�@�5Z�{
9��j��~{NI �Ƈ%|V�@���Z�ў�B JߜV����i�S2
�YイR��C1�P��R�s���O7(HJ�M�?�O���xp�d�¤S��<#ѣр�^�;`�	�zt���j�uXЉ�*��D."o8�'R<z�ɝ�B�j���̀0 =�7D�R��	d��?����_5rȼ�B���3sXH�J���M�VNY�VF���	�
X	�IT<o�eS5�
m�0�&�IW�W�_4�\S≏?��R��Ýr�`��7 ��`�C!Y+5�6�a'�֡Y9�h3B��?���� ҆xȐc�J�*�0��/XL>Xr���	5�1ɴ��2�z��I
zt@��iEH�z&�^%�LAt�F�i�R�)�!��g��i"�ԧG{xT�F)�V�j&�~Ө��(�
�������o���Q�țB4p�v�'���!�əF<@��'��]fv ��8a��@g��;?<X	 �&�w+֭ۑFwㄵ���Հ3op%xW]�h".:;5L%`3f� s-D\Xw`Q����5Ǖ��v1�|"�U��z	��rիቊ?XvP��A�A]LH`��E#�t��Z�`��I�f(^�7h^8n�n��D� ��Oͫ��͉C40�&)��c��9a�^"@,��͎�&*�4��#�b$@�W��I��M;���Q"B"�PU͏%,�<�3�o�A{�ςl�(,!2�L3Y}�`H���4V��0���&��$���'�Vر�G�3�Jl�3
Z&6Ү���(ŝK|� #�E�?��Yj��z�Pԡ�'�0�ZH�Ê{ӢM�'Gn9[��Ld$h2��^��\z�&���+$t@`!s���C��M��'Vאd�� H~�4`�߄;|`7��L���-���@Ǐ,)�)���	��u�r� �y#���I^:��2_�,��< a�I	"̶�뷣�%.1�����N�g�LH� �1\0Ѣ��$�ǆHF
�pS�Ձ-�D)���{o�lp��·�:��>1�aЈq�u��,Q�|,��bٟ�7�ܗ���O6
�4qX<�F���8a�ƦuzRμ\V������I�jM�$����5%ɾ(:���@���xZ�I�'����M�+�l4��Oѓ�\���B�R	F!~����T�$���	�-ď)�b(�����ZEQ�JX2dMR�)]� ����e�&&9{!fХ������9ʡ�t�,7�I	�K�!7v�£��On��a�6�T:�,8ƽ�ԡ�5�M9�K�:�n�0o �$)�:>,�i]�|"�Τw|@`V,ۉ6ot��s�_�(H�(Ѡ�ް{�旿:�J���
�d�9jQH92elٓ��
[�"D���!�̘+��Eg�0�!�ÂN��`�BЧո�Gyr�ۺF`�ɡ�J��e"Q�Ҵ�CD��ڒtr�B>*�-s��Kb��,cP�H'<>���3C���A�m�0ӆXx���^�}��H��I	$N͒���a������,�&��h�t�*n�mh�_~��D�I��K����faƦ���$�|ybQFL�04�YC�ԫ_�:u�a���`�<��	^ U��*ъb%P�C���!�>��Ţ��,��x���84�8��[,a�2J�`#@�Ӄ�%�*�![��GJȌW�, �	�-G:��$�!L�Eaa�+n��Z�o0O�&p{����
���.�(D�����7 Z!;q@�.嬹T]�I�0X;� T1��J`��O�n�X�
��ؗ(�}���	6.{��ū�N� ��^2)^�Y�bGۢ]���;%�PT�ᄧ�=�9���>T��X�aDKt�����v��s���@�'�P5�⊹{��y؁�̻f:��{�nM(����N��ܜ;��<q�D�T��8x��U�Q(�c2��+�K?"�Z$�R"lؕ�p��3ªZ�M� �o�Fx��Q�f"j���3A�'j��g�N�0`���)��9�m��A�~�Cf] h����X�m�8���o��+b��=~��L��9BGh�C,�O�BfDh�=aw(�4��p�3H�+�"�J��ŋ<Q*Y����@���p�`�v�^y�3�҅]t�(!�k��sP�GNtB��ݐ=�|���=ʓ 9֙KІCFTz�ݒ9�l�X ��c�y"��C*m/��1զ�� �"=��X�G�*��V���Va�A@�꒲b�Yjt��%9��L-z�lc���Z�V���Ҝw`���SK�%ٰU�e��^�<�9�F�	?�L+B��&^�@ٸŊ�rd�A�,�<ig��R5n����*�u�v�G}b&ۑ@�"Q'��A�M|�< iń�v�,��`�@i�<�W�BPA>�q'lӒ��)�Ly�6Q�Ût�&�q`m��
��ɸ��YI�� '�PX�'}�B� M"���!?��XH"�G-A�����H�}Vp��C��$ݪ�;1���G����'嗫;��	rM�:�A4�ɼx_d��-!����<��f���X@���<4P�NN���$�gN4(؀��;8(�1&��!,Je F��
F��s X�M�!sW
�Y�܉y�mI�g��)�4��3s�D��E�ܚ3؜�i�*9�V˒e���1F��<���X`H}@V�HR,�[4l̢{H��ȇ��b���qu��3C���7���}eF]�I	�T'�,ct(���x�w��l��pHF��9T�����w�' �%�V��5x�p�����G���1�Ef�X� ��i� i�,ъ�l�\ԾD���2z�l�&N�,Yɐ��UmK�Z����Gm�4��;U3>-AfΏ6��!K�G�^]�!�'p�ye�;8�Ԫ������v�inP�KΟP���$���l`��VfA���;.���0�X�ĸ�嗦J'B����vT�/\pu���9*������"�l��ꆛ0F��j�"�2���@BX�j�c�\/S$HKc9��`����5N��z�b��0���"�"�.%�����	�JQ��[��ͺH�T�2��5=�������!1ʌ�į,!���l���x2YR�E+.|f|�aG@./'D�+w���cTБڂGF6rԊ��źt&Mj��\*+rtT�g��)+Z�[׀�$g
=r��Zi&�!�@��q�I�Q�cҠA�FB?��!b׮a�����~P#'�pֆ�e���1c�1 �5rb&��q���UJ��I���1 �\Y+k��@�d�4j�%P-�7vj6��1c:t�,��%G P�|�G���$->�B�@=�4��e;w\]�#��B 8l�'-��)���G�	>dD�"B��Y!�J֢�d�PC��7'$1D�_՟4���
8nT)�"S G��}a��#�M��L�?Y�2��� <���34�\�O�t�%��I�0$��[�E����O~\bD�z��=��.W�`��YH��]�
J�[r�;"�x�	e�s�] �8#�"�sb�W yp�!��'
$iX�!��j
%� ��*T�������5�6�IP�Q�	g�Z�̍4���Rd� �A*W�����#H�6�>�1B1��H�/��"����W��I�-���q�2�k8�	8x�ɵ�E�^WX�Pr�A$uj��g�����$���J ��PQ�"~��Eb���(m�D���Z�oߦ�� ��5N��HQ��"��A�&i�k�����Mכ~	F�GFy�7_jB�)$�X�E2D��(z}�H�U�E�CF�˧��3�Z�X����W�ہ)"u���^#<����)_=~�5`��҆�S�x��Y�F�ĊI�n¸;��E�Q��)���C�I�T�,���
���8�*�.P;��,He."���>�0`ENB�:�rI{�AL�'\d��Ŝ)�V�1��W�u��H��A$� *�F�q ״w�"<��C(XF�%�z|hڕ�P� �j��e�+aRm���$Y�R����)[@��'9 ź�hPF��X�bjOvk�� ���Y
��ӡL�XY�f��q��#=Q��N,^6��
I�xw�L�RP�-��/�p�Z�mޜ11جc��>���yq��H�.Ua
��k�\�l�E��������<^
�`�ݱm\��Ҏ�D��xO��% ��u���Ο��h"$ָV:H aV,�?fƞ�Q'�ɍ'@d�s��g�$�{V�ɝu�Q?����G�� �rL�C���a�B�B��$�jdp
�L�IT�ç�>�V��$}Q�K7וa��]ҩO&훢�:q��5��N�'��(���L2)ƚH�Џվ"��q���By2�?T���Z�!/��D�zf��h��]RZ�X�'�4;�� J�{e��"Ə�+.�D�d�ę*E�Ԑ����!`�̆�ɮH�x�˰Lȁb5���eMD&L�����2 �Ѡ�y
� �9�FN�+��ݰi��J#�=�"O��
�.�	�bl2��ëE�Z	�"O�� E�Q�]��B� M���"O�=J��è-z�d{�i�e,<١"O)�P �,�`�8f��8�z9!"O��s5n\� ��E����;8s��"Ov��E@�$�0$��ol�B�"O���@�f�b�C��ڗ��Aq'"OzaS� D�N�̉Ҷ�D����s�"O�h8 C]�p�ϖ%��Ay�"Of���B�A������EpD�JB"Ov���yAt0�4I�6ih�P"O���eڠnX��z��#]"%Ѓ"O^A$K�0xr��5�pӞ�b"O�q�-Juݦi0���y�>%�'"Oa�!c�����Ԫ�]��� �"On)�"+�M�԰p��9�(�"O>���3�h�0�e�K> ��a"O4�2biٻ)�@��<xr�Ȗ"O��(�NW�+��̓7�֏*	F]��"O���,�W�Xy27� *-`l��"O�	p�Go��=�@�>m�j�"O�q9Q�D����#���9�"O��p�j����) C��.|����"O�$�����*L@@h	��0����"O���bI#��
��Ȝ`-����1O��I�+*7���q&�[������I);*&J��:ڠ�+� �
�����BR d�bT��-J;B�
d�0�?��U�ρ�&yiG��@0�p�5��a� �6p��ٴf���i��F�l-X�*�$�:�)q��~R�a��u��MZش3$Q�o*��8�g!X�M�f$ ��Ɉ0^2)@��k�`є�i�=�����2�<�[F��:)Rތ� 3F�T)۴�ا���$Ι���:a\0d��T(-���'�H��1O���7��0|*�iU��z�2e��r�^!�L�E�D��[侹J��iD&OK@�K0i�;>d*@�ib�DI2��Q ԠS �I#��4�0����#6�2s��B�Hk@/S!)z�}8r���3VL�O�O���ưi���X i`�D���(�4
�y �C,�
y�e���<E�$Ĝ�]�>�t���I�@Y�@C@�Cέ�u������ 8 a�t��t��"5-/�I��*ϐ�I�Z_�-���!a��K��/E{�n�'Q ̛$����;i�Z@� O��<�ٴ��>�3ĬE�J2Xh��E�Wg��1��OXТT�fXZ0�>E��KӞ\8j����Z ����?�p��#_�OQ?=z2�B^>������/|����#'�*0̓j/����'Q�g~�-�� �� 7�����׽3R���M P{�'f��)��@�6�k��E����pQh�>1$�OrU`O�t�j��Q^�I�4X,y�Ttr���<镮��̋L<E�$��)X) P�P��=��p�!��0l�n�nZ�J1Oa�D̂�0���v��@�Di��l�.� �y��O�?�A2!ʡCx�m�U��8|�� .�I(�?�� �<����=�"��L;���BB�N��<O����.%�)ҧ{�-���Ȫ!��]!E���nz~� &���Kn��
��)B�BJ3cV��#��\6���m�I12O؂T���'�T,.(�ȓT?r��թ�!Oٶ��gT�d%�9��a��i�dN¢2�2(H���UBNх�PY<z aV!2�DTrS#��&���$5�Eb��T�+vN�bcJ���%�ȓl�4ʕD���k����Vm�(��9<0�h�
`��h#��5PB���giƊŭ~8 [�\`��H��oD�h�d�=,�"�
�xD�ȓ/P�����=���aEQ����ȓ�P:M�y�L|�f�1B��݆ȓ��#�D6z�tI٢F$���ȓ�@i��D+N.Q�cCI�&�Y��S�? �����:_o���j��+���:�"O@L��e�(sՔ�C +j����"O8`�Q�L��H��oF�/N�k�"OD��"�8�L*S��;N=�-�"O@�17j��w�.t:�- 9H��S�"OҔ"qjH[B�t��l�&uEa�'"O����Cт`e(�8�ꘈ#AL�[1"O�yǋZ�h$ѳ�� 
,����'�
�B3_	}�L�EW�b�
#	�'�����x�(	q�憈`����'�*(����n���I%b�c:h��'RX� ����H�r$�3���<���'�>L�P�j��P���uB�	,�-���L� ���_�h��C�ɀw�I�go�7�$*1�\1K�B�	�(��X�SE	c���� ۂ�B�	�0@�0�vnҔl��#%K�B��= O| 2�Z%k��E圳M&C�I>k�)�pb�g���̐�5�B�I�l� �[S��.8O�hz5ț�Q��C��#�P��T���a � C�nC�ɤ+�ԋ�[)qֲ�f�֝FLDC�IsG�h��O	l`L����QC�I��$!�(���Fl�b�D�&C��R�)A�"Dʩ�4@P8t��C�	~�"@D�*D���"�:��C䉶K�FՓ%-��v Ѣ,�I|C䉭%���`�ĞP�t�1��^g�C�	^3��Q�KG�*�ɚf4xC�#B��9S���`i����?JS.B�	�V��� �&
�9�Nu��n�	),<C�I�<�ЇĎ��0�o��s|B�I.;<ı��+�.Q�u�R�4�bB�I&Pl8u;�L�>w�2]j0�Ζm,0B�IX����v菿	=Rc.X79B�	�wC^lq��@�l�����f�VB�I �����N�����F:B��\F��t�E�Y�(��� ��T��B�ɿ �hj4��;79>Ԣ��4p}�B�*̭q֏�v(�P��ԀwbB��!�R��+I�#��x�KS�*8B�I� ����oU���������5q�B䉌'�
�-y��țS����B�I�g�8�CC/u� 8Ee�I��B�I	h¡Q�)� ���'	c(C�ɒ��h�kEd0��U�}e����']��� �o�d�8��� P|���'�Z�Q¡_uT��cZ1*K
9��'J$(Bb�G�����N�U���8�'��fn��,Ϧ%��j���p��'���	1��M:	�W�-q�x�'Y	�j�D��q���S� 8��'���p��`��� �`��Mж�H�'�.��v�KQ����X�Ibd��
�'������I~�� �틌E��Y�'��A���� [.����I��P�R��ȓ'�&�$�J�K����q^@�-�ȓ���2+H�,{n���!A�rd�ȓ)n|�1Wĝ��P󋁰@��M��{}�:��΄��!��)(>,��g;�yС�2Y8"��VP��.0LI�3LD�#T��+���,�ȓ4�@EU�U�� ��$>�ĭ��5d��@�X��ܒ#��
,����S�? �I��nE�_�t��	U2S���5"O��+V�җT�4�!�{ת�!"O�<�枙{¦���]�QՒ���"O���h
OQ������}�"O����ɟVK�$z B�0d@a��"O���5��:ᰔ�� GrF�)�"O��C�@];��#��H�J�jC"O�@��a��@��E8|��,�$"O��jC�Ŝ]pp�q枫d��-�"O�śB�.��0b+��b�d8!""O갡�A����@�;��сE"O��y�㆟L���s�2����f�<����&q"��[���7vT�)kVm�<���pr�w�xJ�q�l�h�<��Bƛh:���@�2W}���DVd�<�ǌ�/J*��T-Kl�t�z�<ID� jQxVe$Ð)P�j�s�<1֯�r��Тu���1m��S�gl�<y B�	7,��Zf�	�g���@w��s�<��ģ�JX
��G�N(�Hfg�n�<�u�Xx-���� �8��H���`�<�6�I9�
Hh�iA	U���棙Q�<�ca�)q$Z, ��T'�$�$�M�<0i��<vʬʑ�� �ĉ+��M�<J��g�b�_�@S� QA�<�#e�'
ޘm��Y+�ݑ���y2��>�h��	�W_���Ca��yr/�1H��d���MhC�oY��y�cLZU�`���	��܋�B[��yB#V�na��2C�r|�9B����Py�d�; R�� c�.*�8y8�VS�<!��_�~h��I^,\y�E��ȖW�<�@���(�)�`�s�:�SV�HU�<ф$&~����@�'�H�;UOj�<��nPzH!�I��xVд�`j�A�<"
O��LФ�̢�A�M�{�<1��E�0��qWϟ�/���i �Tl�<YceʽU ���ʮo�
�	�i�i�<a�(TP�~��M�\a��q���k�<��.B�A�Ry�S勦%� }�QLNk�<�c��Y����N&�p��J�[�<���ǗZ�2�+R��#SX|r6��X�<q�F�<�A@�`b�NZ�<�P��P	J�j
EO�$�T-Y�<Q�e� 2�¼{a�W�.>ȍ�ģ[O�<� �̚Q*��Ԃ5�Qqt�S�<`a3EȠ̘B�B0ʹ�AP�<���j�.%�$�2�n0��FO�<ِ"F;�0���O>k� Q�c��K�<q��R�~Μ8�!��dq0h�mXI�<�4��>�@�Ҁ%ӏ/ ���EC�<1Tj�"���G�h��Q$~�<��O�'4��M�WgDt�0-/Q��B�I�İ���r����.-a�B�	�5jr8���Y$^�!�g�.c��B�	�>P��;�Ǔ9]���ӍK:`hFB�	��`��0�Y	b�6B�?H��C�I9<r��և�/0p�U�G/�,��C�	, ��t���c4��$�ʘ�XB�	�&Ʀ% �H[N�T�#�%\PB�ɂCʪE�Tg4\��cďI�pVB�ɽ$�ܥ tÛ!0��a��m:X��C�	!n�ų��& �f�	�'�2R��C䉊+�Q`4��ZO ��I�zVC�)� `H���!T�� M�9���"O� �5㈆of�E��kʭG-��{�"O<Z���$~�9�W�9$)е��"Of�2�F_ �Ba�C�X�<¶"O��r�Z�a��5�=�x�{R"O��f��4[{ڀ�p�
a6��e"O ���&�c �ے> 8��"O�����#2f�!D&S0u��"O����@�1��  	�19e"Oz�8��]�����Ř)�(4�U"O������V� St��9�"O�t)�Ƙ�Lt9�&�P�J�:�ѡ"Ox�rgD8q\hܩ&��y:x%0g"OV�XbL�rN��ҵ�St����q"O�ԫu-�P$R���F]�R��$"O�a� ̚oKX�JĮ�>d���pg"O��z$l���F�`�N��ZZE"O �R(C�x���(M���I�"OX��V�&/h����>!"���"O����y{rD���
 ��Z"O�ȲFoĪn$��@U��>F�0,��"O^@�i��~2p֋qgB	��"O�5�bcáGbB
�,��j0@)8�"On�rD+Zt�(�4i^`}�%�"O�@JԄ�2��k��1m�T��"O<HSI�@@ě��d��5"O2lB%`>qP���A�abȳ�"O��Ѩ���T�Q�٦�4Y1W"O>æ��k�ꭡ1o���<��"O�AK�̎�t�4�NH�F�#�"O�@��R�0Vl��cC�$��	�"O�LR���*{zbr��sf�iZ"O��H��TEq��U�_fx��R"O�)"$��}����Iߚf�r�"O����kpa�Rƀ�(p�p�B"O���6��BBj��ń#
Ii�"O�e@-$z���2 &�Lm��"O��[�?̈Q���72�($��"OzA���̽�bݲð���"O��b�˥]�e�3'۷�"���"O.�[�FȠA'6�x0&;L�"Kp"O��V��'$e�1K[)K��	��"Ot�
�o�V��U�0�V�9�j�YC"OFy�DG9wS�t� cU������"O<[�JX=i�h�f�w�P+ *O9�c��+O�HXacHT9DG���'�bY!S��	�b��h��`q��'��M� qsE7n��Y�'�p����Z��5����(r��Z�'s̑PD#աZ��$f�����'I�)3d
�&s�t*F��\���2�'���k�J�& KNU�Ek�Y1���'F��x�B�3�n�e�!eV��'�a�5LM�%�F�juϙ�i�Lu�'��&�.�D=��� ;
���0	�'�Q   ��P   �
  �  9  �!  �(  �1  -8  o>  �D  �J  HR  Y  __  �e  �k  +r  ux  �~  �   `� u�	����Zv)C�'ll\�0"Ez+�'M�Dl�Dpw:O�1"�'"d�?Y|��̛'"����E�;Bc�T�`��>DK���(R�9O %r�%e�i��#�?U2���?���%�f�:0������R�#���(:�\٥�HC��h#B$9ؘ��ǖ��u���!����'�M��	q����rj�7y`�1ud�$L�jq����O��h�ϐ�,���9�@I���
���(����<�����k��P�Q�C�Wp�i��"Y��@����h���fyB�'z�q��O���'S�Pi&�ؗ~�0)��I�#���@��'���'-bY�L�I$C����h�����|@j9K� or�){��!��)��	�<ywIɏ({�upd�˶w��y�rJCA}"?O��O|�	�.�>�u�?���+�2��@0AJ�"�j\� ��O����O���OR���O��$�|�wG����I6z��XWAG� ����1Gb)bt�'��i[T�iR&wݙYÏ��u�#Gs?�6����q0�m´b媵�`M5����iU�
��>��1�@��is5H
1G�b<8�-�!r����kۋS���8�+Oæe+ܴ[o���O1�	"n���c܊{���`�-H%Ct+W oI�7-ҏ�j�Q�O�"a��]R�-T3�r������t,n�)�MK��i�n���#�#ɞ�Ps��������R2���527m	㦝q�4.u1��ĚkDJؘEמQvĠC�_KؐsFBH>TI�u0C�=�����9w���q�i��7m���h���!U�񱴌�##<��+��i�܀�Э˞���9B`��I�OF8b�gc�ܪdR�`���O���HC�-cV9;�Gh�n�������?���?�rO��؛F�?����:ؾ@��� �J��q��OB��?a�����C�������������U�i����@d��abJi�i><��;��'P����p�y�G��u�¯ڬ-�8��2�B�K9N��!+X;�0<1�	���8�I,��DO^輁cv�����j�a�	s��'����io�ē'TG��mBh�[F$K.�O�o�6��pH%dA�8�z9�c�8��lY�4��$a��ulZ)Jo��	X��MR�3W�$�ʸв��w���.x} �-�9L�'�|-���'��	�\���kH��ن�D�Uy��jbÔ�$?���.\h��K1G ��B(ħ�h��u��%�!�%#�
�Y�R����RF��O��n����O��4?�̔�tH��|砽*cl��nb��#�'���'%�I��~E�傃{�@�� Y;80F�=�� .�	Wy�?��b2`H�t�iy&��67!.=t�'�x����D��Q��I���N�h��8�$�#1�.D��'K&^�'�@f��;��(D��1�"�--��I{1*-RO����l(D��#!H��fY�,َ<t�k��9D���c��z[(ـ���4Ր9y�k6D�p�����k�#eĬ#E�<Y�CF\8�QB�DU�l{Vb��)T�0��7D� [扉:5ø�5��{NVT`�)D� ��dJd��J�n�x�|"q�%D�LY���$f�*��'��F���)D��*��&�p��)��UKL�)(<O<[!�����I�����k-t��,c��&g4�Y����۟��ɦK�@]��Ɵ8�I-R���Y���ң/ח0�7��,#P"�H�x�����	�0<���	%���sU�إi�N�P��Ɇ�|��sJ_�!��2%�;@�����S�V�$�OL nϟ��a�kJક�қ9��+�Sy��'L�OQ>���#@>i��g��i8�}aF#&��T}B��2�M���[���!JY��@5
��(�6�|k�7Q��;����X5�V�Rb�ks�ڦxˆH�q�"D�@i�*H6���1��)�"���L<D�,X�HS=?<��p��I˦����6D�$��hD��>Ո3"]9sL�B�3D�Db���Q��1q��ߴ(k��k�/D��0''�[<��p��t��)�4 ɦ&���A���?�vӈ��O�˓@Vh��`�-}�,J�G]H��hp�z�Vis��5����IZʧ}��O�q�⠉�m�Dx���+�ԁ�2d*k�0�%�ʿX?��R1�]%%1��t[B	�~�A�yhB̀u��/�z��2Ő�H�H�<��D����|�I����I452�Qc�p�R����͙|���&��'Kf��G�K}�F�0�ˑ�#��)O
�nZ*�M#J>ͧ��+O�t;��A[4H!�6��=X�,2w�@� ��({B#�O�$�O*�� ٺ+��?	�OVDDR�~�F!ѷ蔺y�Mʕͅ'�(@�dk�O���'���wƗ���go�7�b�(�* 9��xBώ�B����'��p����2�R��ь�:k��aF%�?���?��2��KNԺ"$�&@3�X�C�=�]�5@�:ivtB���hA
�O��m�H�'d���l�~��Q	<���v^�]��	�4y�q���?!B��5�?�����/[��sʍ
��u�_��� �ؑI�-W֦�s��:1h�%�ALP�'��i�ū<���h@���P�B<���Յ7�-J�ǟ%[}�5s"c�2C��#?��l�8��M~���!)F�;�K��W�tcblG����0>i�b[�^(TUڗ,*;�H�r�\M��(����!:�.��s�����>4�Ivy��I�6�8�I�|
��D|��A	��x&�[�N!���Q���?	��L�6:����jӂeb����������O$7�����΀�Z! ��6��,�tڎ���K*9�#~�cE�$L���+�8�V���N�e~��W��?��]���&?ΓB���!Ors�1Cwf -UlT��ٟx�I������-�2Y 5��6��!�i�Ui�?1��S!wx.k|�5{�mV#R~^,���L妩��͟����K�]"��ڟ�����8��ʿ��.�Q�q
%/&
pC/�V̓I����ɒxw^���N�?<}�E���_�d���٠F4��	n�rIh6-*�3�	qZ����#�E�����.T- {8�%�ܹ���Ohb>c��H�T�y���W���aYR��Q$&D�@R��)
�,c�g̅4@.�F�O|�$M���$�|"
��9��xY��'r������!��کE��'�"�'���]�0���|*�B�)4�L���Y�u��L�w�X+0&v�#��ЪO�OQ��p=���/���Glƺ&�e���_'k��+�O���TE0\Oh�
�����
ѓs�ё	6��i���;gB�p�J9n�L��Y���Ȫ#o�Сj��))�Ѻf"OfȘ5��"kk��ϝ�Ub	���|��>�)O>�aG'Ħy��Οxz��)�vu��H�Wn��2��K �I�|�t��꟤ͧ
��	G�[�$�y�� �6.TtX��"$,��	�JjX#<a�B�p��=��� �Q��A
a���7/�O8I$��`�W�H��լag���f2D��Tf��$i24�0hӲe���Kql1�O�8�I0:���HRhֆf"qi���p���O���YǦ��	��H�O�$Y�u�'�؋�OZ�|}���R��D���@�'��fT[�l�I[�L��br��r���j`�ʊ82N �!'?�'E�/���d��L������ [��9�q�D�M���@��#sV�	�,���٦����D�OO�)Ι?�&]��EF�pI��� �8Y�y�'�b��8RmA{{���VaP5\P���8��?�gX��'��I���e0d���Sb�QQ�k@�7��O&���ON�� i�\6����O���O�(tK|��^1:��|��1C7`�6~�>�nfz-p3D�]��8�	�G��v��6��UkW,��g�x\0r�Y&V�Z���k��v��p�+�%E�0�^ˈ��fk����5�=��}�ɡ�M���Z��a�������$�O�Ȃ���Ij���2��o�,Xr$��hOT���f׆D�Vإ�$@_"���$�O���'��	Z���'�剰(.����R�P��;v���: \0�B�0�,��	���	���
^wn�'��,	�u�8�ZccR�>���C$	�(���
�'N�EY���1%����$F�/'Z�@�5~��y`@�mڤh�l�}p���(��7�:?3�4�`R�x�'��<~��Sˌ�V\�\��s���' 6�O���?���`��`^��Q@O��qpV�n�B�	՟�Ig̓3��8����C�Qy�ᕰ��'k�
jӆ�d�<q�4UQ���'~�$%>11��)���L��
�:�R�4�	� �	i�r�{�g�:"�z4�A��<q�ֆc�P�"3NNO�T
�i[�P����a6(8 �^�y�扺vCм��L�Yu�4��,R�[�����
r�i� ���O�dpW����[�]8h@��XF!�Op���O����OΒ��c�D9�.8_��P��k[/P*�{��&�O�����&��`�����Ԥ��2���<a5�Jz���'I�]>uB��Qş���
,�\�1΅�+`��u�PßD�IE��d�dV����O�ʧ��	Zd�8y�Ϫ;g6���Ʌ!`R�u�bvkW�v�|�i��S=YYB`Ifa"��o�D#��!�&-x�	�@���C+Bu��=�M#��i{��S; �`�+�4D�̴e��=V�ГO����Oܣ=��=_��_2mUP�f G>:�*D�~��xo�A�ɇ9x��0� �.|jTfK�%<D��s\���?A�g�'�
2`/k#�}�DȊ�{P���'��'���z�$�'���'��sю�<f<�3��vș�'M�P�DЭ2w�y#��7���a�'p%6D��"����#	<k��B�'�� �W)4�^1�ߐDC��9sP�\�e.�O-����;{L���C)�@��"O� ��Ʀݏ0�b��J�a�"O��C���+*u	«D�51�"Op�P���%�ʍ0 �.V��i�"O��A��-H.�|!�Q8X�]�5�'�*�'�D�"�I�K�$�q6�=g�N�	�'��@��S � ���BUg0`�	�'��E�v@ ��c��c����	�'�0����2	��xeΞN?l48	�'�H�gh_�D���@jC�ȡ
�'I|�Ӥm�j>�1:
-��P����� Q?e�f&�=X�-Q��\�q[&��3�.D�����7[��[�j]��p D��1��A�tuB�X�ҍ���+D�THf��?��e��`T�]h �+D�LRG�>�H8j��W�[n�	 C�'D��"�iӕo,"}`Dm�oX9�D`�OȠ1�)�MRT���S6j �h��AG�H�DE��'�E��Gр
X��*�c��6�D ��'���@��`�"i��� ",,��'��a�B:.jj�U�7�\��'��x� �[����m��s�Z�Z�'�좐�M�
V)�篛+}�8	�(Oԥ�R�'��l1�ᎫN3��.�G����'���Wa�ed��'�J#Pc|�`�'�����o�.'n(�V�� GT&��
�'��@
�d�q��2ê"H 
�'�l�qb�F58gt53�&��ڑ�	�q$l��:��H0РUSQ���1K~�NM�ȓ~y̴ u�۷P+T���y����ȓC�^1B!�D�9HȔ�ی@}� �ȓ
L!92Hp�L�卓�g�8 �ȓD�ԄxDK�Hk�(�T�X0Z��x�ȓ��*4�uLE�ҡO�~P�)G{R�
������`K�(�ؘ� o(G��TS�"Ol�5�P5OY��q4�֞XvjMJ�"O赡�Q�q��ȣ���*D��m D�8��W�w��)Hd"׳U�,�:6 D��؅b�v�
icv�-��X�k#D��Q&��qcP�'H�[��4��n�O� ���)�'_�)�nʵ4Xb +&�26Қ��'���
��R9xn	C�N�3�|T��'�p���d�R����'�!�`T��'fB�r�%�rGNm@BͧO}����'�,��ɡfT��;�Õ�Y�:�'�­��
 o��}[V%�V��/OB��'� ��b�pf���PD��|S�s�'沄����>)MZ �׼r�̑x�'�h�/S&������r�z�b�'	49"S�^� <yu���c� h1�'�*A3�
�;cx���-Q\�؉C�#a&t��1�DSg��8x`"i{���+x��5�ȓ\�����\�s��Gߤl��_x1�%��&n�q��$ǖ^�޸��#��k0��F�N�4�i��ѣ�'KD�� �ѭeC�4zLeɱ��u�<�fY�/Cr]� ��_����u�')~T�����5w������n��(#�m��u�!򄖻6���A�$ �3A��+A�}�!�$�z�(� .֩U0YB����!�M�P��� G+OPUjPː�E�!��Ր�T� G"�܅k�i��|t!�B1��UC-?�� !đZ�$�:�O?��@0BRn����0Cq� ��@�<1�OΞ�2 �T)|#��Д$�x�<� "�V���0���h�3�*M��"OJ��㇋3n݀]I�,W`~xxj0"Oɘ!h��o��� ��L*IvZX��"Onp�wI��:0�U(�bN�d�@B�V�<k�N'�O
�S�t���p"I
�F��"Oc�:dhXQ'�)RKz "O�"Ѭ��H����LC�e1E"O�*�^<k��98�}�Ƨ��/�!�D� 0�@��%��Z5�̑��Өln�}Bh�~+�f�阖�Zr,���S��y��پ5�aX�jZ	0D�Ój���yˍ�6@�e�a�݌+]����ĳ�yn�1 �nt�1�+Yג�z�X��yrG��nhr�[d
��P�.\�E���y�	�{y�)�u��=pĈ�G�ذ�hO�������d踪�h\�L�04Z���{�.B�I�f-L9���Y�w���q(	+N�!򤘾@�����i߭)R͡&'	kd!�D�"�j(���C�r)z��Ńz!�$J�����^y���J��$!�ާh�P=*���]lN!���L%|���
�O?�Bi���a����Q'ؘ� C�b�<����`��iƧƕ+������h�<�M��l�p�ȍ4/�1`\`�<�� ڟ�	裌O�l%��L@]�<Q�l
.	 ahtD( < ,�A�<I���Y����3�N6C�9HTBAy2���p>�kψ3�Z�`.־*�.<����F�<��a{J�˴n_�-	�a��M}�<a��;���%��#��Lq���S�<!�Q��`�a-Ȥ;7�0��h�<����X*�QӠ'�*eP���dx���H��X�TE1 ����0
�6ΰ�/D��xT��;+�%��g@(�����-D��R@O�=�v �3���M5@Հ�8D�����["9(l���[]�""+D�0[�A�9/(�d����u#(�')'D�T�`��'�J��1��%q��v�$ړl�ʥF���:�YxB#��w�E{"C��y�ד
+4<��nS�c���q�ԙ�y��(In��QL�n��BBꖜ�y2��i�$��FC��T$at����y��qK �:N�(u�S욑�y"��<J�nq�΅�L�豚sJZ��?Ys�x����(i[��$:��m@�[��u�'D�tKwgӺ���`P�hy����M2D����V�#������^�wS��Y��;D��b�%E	7�1�s��>~ٲ�"�4D�,鰡ޙ/���-��LM�=��0D���q@�9��G� ��6�WM�<q���~8�D�uIߧf��p���$ S�J,D� �W-2m.}YP �	<���=T�l�VM�D���V�3g� c�"O~ٛtNV�q\�Ԫb'�3?~N� 0"O<͸тI�l� �[QL	.Le�X`�'�h���'��ı�,�d�8��3#�JD 
�'M�2�aP3�N5�6H�jLtt�	�'��(�+H��<���S�a�^p�	�'��8�-�B��X���ދk�\=��''E�e��^Blu8sņ�3`���'��	��1|�05����;2I�`�����F�Q?e�F� �^���u�J1	qx�R��/D����H4��ۥbT�0�,=sT",D��v�ha�
=��)zP�ƩY=�B�)� >Z�5/*�x�l�*LNܣ�"O�h� �3o_:�(���"�Hk�"O6��
�?<�$QG��0 ��'R��
���S�c �).��%��t���G2c�:d�ȓph �$� !��-B#j� פ��'���#D�*��<Z�܎-C����I�����I6"ȕb�� !B[Լ�ȓR=29+�c(�~�҄G+�͇ȓDܬjaMمN�4��Uk
=P0�0�'���(�~en<�4�¶z,����D<4���dWJqB��41|Dx���?�H��ϴI32�K�| �ӂ�(�`��l6�9�ۇ[u|�s�K!%f�%��E�s��
If$�C�#�X�T���	�'w��I>Z�BIz�"�,I��!WfߚV(B��b>\Q�K"�|d�tB\���B�	�ﰐ#!��=;��9Ұ�Y8ߘB䉠e#��h"L%>nfI!��9<�@B��h�c�+
(��@
��ԇ�nB�	1k�������!����;�L�=ɶ#ET�O������MP����g�����'[��DfI �R�	r��]�*)��'�*�G��>�8y�!�X4�!�'�:�8�&Q�`��p�`B�;�B�)�'�8�b�,N:^��<��ߟ5�l���')�Kd�	!�!�AIS�vz����;)bFx��)�n����)��_�T�KbN�&רB�
?J��3���I� `�G�/NxB�	�WJ���E�3���O��#{xB�d�䍈K}�|0��J�jB䉎4�j �i�ZH�p���UwRB�Ile\�2��@Jޠ���;nY�\��^��8F�I�����r����Pɦ	�g"x�W��*Ѭu��D[\�0����Jh8��I����,1�|�g�W51� ��&B߉n���� � ��)��`�\����g�(~T��\�(O�A
7�B�a	�I�`I�*'jP��M^$z>ڥ3P�ĥ}�"�1S�?C`����!�(OBC�'�&6��\�<�:��տA�T����,�˓�0?��,�-���w�i�}C�b�mx���(O�Yz#h%}��i���@l��Z���!�^㟨���#w���ƌ���ϝ�NXPa�J5D����V2)����\�D� g#5D��Z��Q�d�J)�2ͅI���v�/D��;fK�H��VAB+g��pt�/D�f'�Y�d��@J��ˀ .D�@�e�E�`��c��B�)ѰB��K��tE��'�	3� $H`�6��8(m�}�	�'D����"!;Hބ���:.����	�'˾�YD�>`��T
oD���'�P\�t�02 �~s>%�'y8u�V���M�x�gf_w����'?@�'P�O� �'��>g%�eQ� ��؄�	�C�Pc3FR����b"�HC�s����ݣg؊=Jd!�z:C䉟p�*����
�^ۺ$�o$�B�	�R�LCW�;���ڊm��B�I��V�( ��	rE��dVo�,����5��*���ҥ�H<=��<
�AJ%!X�i�ȓ$�D������u�X���{&o-D��i%cI��i�k(����ro*D��k�JlHVt�2�@�P�����+D���Ǡ�2�p���5<Ϯ���'D� ���%E���))�5�Ƽ#rc'�	'��#<���X��_�y�Ŭ�Tj�:�"Oj9b+߰Zel��ϭm�.ug"O�ՠ`�.] РXR.9�`�B�"O� ��h�JF�~r*$ �*�o{u8u"O"��dX���9���=�� Au"ON=�dN�$B:�rBA���(2��OX�}��6:!�0�����w��-U���ȓ��t�g�ɪ>���6ɘ+*
!�ȓA,,���nӘN��g-�$l�ȓth�%���"\�����$U�1��}��-r��9	�*�jd�LJ����A�h	(ԥV�$b@��Q��I?=����D�29����Wh�1Rh�sE�9,�!�dƙ	��90b��x$�%rE*^3!�H/�Π�tc͛
B}:q�Ю[!��H���h1	��0������7!���'B���c@�I�'ezA��	џ0˶�M�M3��?�O���iG�"Ӏ�R�^���^�.�����?i��v�]����M{d��",7�}>�9vZr���NL`�s"<�� �S!���b�q��Ct��S*eH0�rc*k�l��'Do��#>�Q��П��ɥ�M����dCϨ%��j�E_�%QV�A����?Y�������X��D�
I��Q�W`��X���(�;?��O�c��'�F`j�)�ԃ��8(�/��b�
 �<��@"���䧚?��O�ܺ�ͩ�䔋���h� @c4�	<�h���RH�>��S���
�^�0��Ջ!�'�V��Ij���ɇ{k4�i� �9� D&0��$l?YT�O�T>�*mO��Ӷ�"N����K��s�8�q��]~%}�'�>��	9��'O�5�i�@�.��' h ~=A� }r��E��'ByIu�  ��kl� Dc��􉉒�I-H���'ox�'u'��(v��E� =b�C���,)��a��'&�]R����E(Bp�TO�k��!�탚#���H
�1��/-�ݥO
�m_�^����˹q:���`�5H\�*���O��G�4�ХS������[�B!�����{��ӧ�9Oh
���j���6-�v�2G�J�X���S�0�e�'V0){�'g���i�O�|PA�]�2Z��S���r��K�UU�	aPE��D�s�x�C��@�B��3"�Xu/�{hx��2+�O@���``�#%F��-x4 ���L���ȓ9ٶ����)zRU;�*Ѿ}4moZ��L�Ioy��'�rU�<��5�e;7�.\s�-Νa����C.M"�Ms������O@y�O�2V>��	<7.��0,�9:�ڹs���F��d�I<y���$�I�<1a@����b�>�x�7ȏ32!�J+f���Q��*{���&$!�X�ao0-F�İ����\�k�!�$S	N��� ҒN�*�f#˯~�!�d5��RW)C�D�rYbבG!�D�%�`�(�м���G��"F!���:��� DȮo���� ��8C4!���Eȸɨd��<�n�����t!�1�t�@a��1+�
q"Ýp!�d
L��U)↟�6��ŀq�S1e��ۋ��?͙H��R�&Y��/�'-�uX�n+D�<`wc� 9�(�˚�/�����(�	,�"1	�`�Y��b@�U�cȘd��.�0u���IBK��q�������u����a��#
�\���i� ���$�P��M��M�NXa@��A�X8��cA'Ew4���,?�d�B��^N$�4Ɓ ��1H�
#��a6�J�ufȱ��F�kr� �c�6���f���N��'��Y�,�:cb�=�IHj@�� W�t(�M>�O���	-���� 7zHP����o��O�D����k�*Q��!$܉U��=�Ԑ�ƪ�$�j�i� Wc���\7�`���S�I8nb�����4�?Ɏ��,�U
ihE��3�uA'�����'�"�'���P��߃A�أ'�ݓV�Tш
� �Q�p�s��=׊���EޖjBy���_�6�0�����?���p�����?1���?���2�0M� !�K���GZ�o���ADE��<w���'H���Ű��� T�M���Di3?�p�J+i⒱���L��n�k��5:�f|�6�T#I�Ү�9�|ՂJİ[�t�'0���;V;��G$�'�L��S;N�P,�䪚7�M;F�iVB��:���,OH7�L)t���6��B�c�'v��\��?F0��	3T4�a"4�ŤOV�Ez�W>��'|1'�X�)$a�֋p�ޥы��<�'4���f��힭��a�7V�dE���hO�>� ��k�'N$t@�P3�����R�"O�ea�ـq��M�V�j��+"O��æ�'M"�RI-mD�컧"O`|���D�9tr$y6�ʀ3�PU��"O�H
�`$'%i��������"OBq�A�5%�� �M�7���"O��RSg7~�r�J�FT�y� �"O ic@,o,A(���\�	�"O��w(�����*�;��m��"OB�Ձ��T�	�(@�P�����"O|�#A�	,����!'�X�
�� "O�"���ܕUM�
�j\j�KRi�<y��Bt����V�z{�aQ�eOo�<��⛉3Fj�{e�*X��Ey��Rj�<I��H�{BJ]�S�.w��(rHDd�<Dc��6+�(� 5 ��ؘH�E�<I⓴;�&i�둆B�WGCA�<�cL�;��88ڼq���Jn���ȓ8�p=��b<)V����m׃@X���P��	��/��i@��Y<<���ȓ�J ba��=�X�bN�@���S"*Uڧ+X�2�x�d�^�6\�ȓ  �!j��8!@q×L�Kܠl�ȓU�
0 ��3�|:��Բja$���F��k�?k��DOҮUʊ��ȓgdd.L�bbAD"7�ɒ�BHT�<i�� �+� U��[�%�$Da�JO�<�� ]�<�:��=1޼��tF[p�<���*>�0�7Ms����'�m�<Q`�T8T���i)'�h)Y��D�<i15~Ƭ���]&c��Q�צ�w�<�����
�*YS��;кC�IXU�\9��ń\V�iW�G #�zC�	<r���(Bw�<�R�B��NC䉸B����O �/�"M"  �	`C�<-��-
c�M,�ȫ���<��C�	�H�������x���AQ=�C��pvŸ��­��ѳ#]�[nC�	.�$mH"�G"��at��+&cZC��<3oz"���[�aAf<>��C�	�P��hh���a�dea�҄��C�I� {P�����D�`�t�&Z4�C��g~�c���_b Q5��F�vC�I���ղbׯ�LX8���!�C�IrT�����#QLx��J<hC��&$�X���NʞtPp��͔+unbC䉬/�6Z��_8}2����ӵzs�B�	�7�1H�K�r��ȗ�ѝbi�C��$	��E�r��2�8�i�'�@C�I4J�4\�`oU�N`�lȖf�A��C�&?�`I�4��J�dt
&�y�B䉞)zdb��!f�:h��'�cC:B䉴0�Tc$�	b��7�Y'3�vB�IY �Pi�� ��7bٓo�C�I�v2�ᗈ��z��}�p�� ��B�ɨ{����'��MG�qpg��B�	�K�u;GG�5I[`�s����B�ɯR����3)J<�!\�B�ɱF�B��D��+D�a�@ 	 
��B�I�C�n) �H�*��yJ�oȎN�xB�ɳ�� :w�##����U�4e�RB��!O����*	�В=)��%�BB�	�]h|asȦR�<ѳ�"	�l�4B�ɐ&�ei!�]� �J��)&J��C�)� �8 �U�5�R݈������c7"O>��w��c��\S�����H�"O��f�L,)\���D��_���"O����=p,A�UW���P"O�TI��]/xwI������F#�ye��c0�SP��<��34K��y�
�bx�A�_�0��x�r��y��#�~��B`ՙ!�L)Ab��y"�E�O��ecD���d}��.��y�e��z��5�@JMs�1�Nţ�y�͵�<-�D�Q�R��M��y�J�05xtq��H*��eP�y2��B�,w��3��Q�~�&i"�';�3bj]3p��GFQ�J�fU�	�'A�`R�����8ه�A�3Y
��	�'�DH�FU�x(��΂*يm�	�'�:<��KR�H�@p�A�8�L)�	�'��Xw�e�JL����8W���'^��x7��)'q.pQC��iִ{�'>���j�#'��	2 ����;�'E@u�`��$~o�%ʗb��~h�L�'�8u4P�L�`�'�#u�u��'.:�HuBѽ\�p�q�	ؼ!綍��' ]ʥc�'2��ݪ��� %��'�x��
�	T�ua5��A�'dܣ�c���i�lM�|"���'�� J�fH���x0c�J�#><݊�'����Qi�|�|���KMp���'j���*3'�uh�.CK��A�'0(مd��>R	�5=e�q��'
��1�a�/ߴ����B;���[
�'�4X�L�Y�����04P��
�'�l�B�ݼXr&���L�7;P	�'�${���������a�8�p	�'�l�ǖr�9��$N'X9�'�d�i����.T���بJ�#�'��Xr�
%[�`�l\�F�$)�'�IQ��'�0���00�(M�'q�QK''),J��.�>��Q�
�'f�q�^�2��̹"i�Z���'~�jV��+2� $��a2�@x
�'LVA�RN^&7�|�S'�`d��
�'r���c"/~�8�r��#Q�FX�	�'[�Dc&��ZR�x�!Z<A}���'�����M `f�pcҗ5l��[�'��iʕ$��.jhZ��=@��ph
�'���zs�L`Y� A�?���	�'ZH���¡
?�3WKC�8N���'~��h���N�D�CL�5�|Qz�'U�73\��H"���;[�d5�"O�
2#Ԯ+�� ����\։��"O$U"Ѡ�K�<@d�Nd�9"Ol���xq��a@�䅋
 A!���:?.�m�a�Ēn��e�$�ѐ�!����ט)�&Ɉe!��B� �#!�$��Y������7>�D���Ȃf�!���fVXYc7暴'��y��l�!��P Ě�bAA	�@��(>+|!���h��:�D���h�C�B�!�$��Z\ʧ�$Bs�y)GOS�D1!��g�ބ�$FL���Yj�(/x!�dY3v4�s�F������rHI7t!�t�r,��o<�T	����e�!���(���7 ��C����t�Q�b!�� $�򤘱5Ֆ�)%%D�QH���"O4m!�͒,.�T�xFꎚ6���g"OJ��|��:G/Z�F	���'k
��m��X�K���QV�M`�'`j�ʦ�
J�H����4F�x��	�'!A�S�턭�BB¥'�b��'�<\ W�I�Z�d� ��-6�*
�'՞�ۃH\ )�F�(P��5C*���
�'?�AbB�(EU�T���8ݨaH�'Q���B��&t����WaI3j
�K�'�ȭ���̲SzH=B�nD�'�3�'%Ҝ��g�0^9z�nB�b8� �'�����Q@�$BW(ײ/��8�'�t���(D��Fd��5��p�'ި��Gc^�eQ�La�(������'�y(���Z3��
Ʀ4yXh(�
�'K�i���:gE�<1T� ?^}	�'��{s�[x���s
ݭ:4u[�'�z�"�'̱������)��'l
�	�N�W��֪�s@Us�'�F銲HB�D�v��թ��h��]��'AbQ����3LP��k��e�")��'�>��R((2�is��A�F�Tm��'��hJf�%$~c�L J�.<Z�'�	�	Q8O]N(90�ѸC�:��'�N<����8� �5;�jE��'�|�Qqc����BD�M@�2� �'� ��diC�9�P�k�o΅9P�h�
�'%$E�vK� ߂���3ۤ�R
�'���rƂ9��	;Q"@�(�^�Y	�'U�Lx�J+_h�Рs���*r�+�'q�XjBa	1�����/��0fQ��'��8�aH?U�(�����"C�Lz�'
�@s�n�(pP��w�Ó4�|��
�'�n�[��!N�>m��U�Y����
�'Q4
b�ܛ ]
'ɚ5T�j
�'�n��s�[���Zf��7(�c	�'���h#.�~�#cF�$(�ܚ�'���S,ͺn�ҰZbL�$�$\��'o��#Q��~�����.Hy�'���c��[�2�HPK�/S��P�	�'��,k!-�g� ��*K��ĵi	�'�ب� �86������E@���'/�j��.L�R��4KT��Mi�'(�
�nj����۝� ��'�������l�zlK��Z {�D%z�'*N5ag!��f1��� }VB�'OL���X;�L�g��ӏI�<��dB3!GČ*R'�0(<��φl�<р�����@S<H-ఓc�Uj�<�
�>Fᐶ��-@Ș�C�ψf�<�E��h�хc��T��!��|�<q��J�M4�,)��5��s���{�<��m�/P��(a�� �+B�E�עu�<ْC��xǈ�@��|&<01�j�r�<Aq��L&>@z���P�jQl�J�<!�d�N��t� �;h��Ԇ_�<Iތv�Z�9�lϏw�8l�qA��<��Aq���T��3t��آC��<y����~��\���/3��$y�lR�<�����~(P��U����h�ŀr�<9bGT�� p�Ä�F4R�x�'�p�<�FE�>NC@��s��+�!�U��k�<�D��?l	p�eK�:H8�+2	�c�<� \A��\2mqHI�G%A�"�> ��"O� �'/GA�8�5�@$DՎ�j�"OX���!�p�hW.A���A"Or��V�TzʈD#�(&-�"f"Oz$d�ɛ9��'F�%O>
P�/4�<��H[�w�<�D�̓xR΍���+D�h���>�0��;}��ˤ,*D�D���E�\�:%�	:u,����+D�����U� q@�	j.
�H7C'D�d�D#�% ��Բ�-��X{ 4rCo%D��R*ɾ�̊eg��i������#D�\��I�b�^�͌[�8
sn=D�̰`��
<Y2h
��*�:�o9D��
�@!zR����$U�4:$D����� ��-Rub��IH꤉v!D�LaTa�,��pr"�Z��P���$D�<�B/ �M-~�ˑ�ڽz�TcP�=D��(��O�'Ǭ<�sa�u���:D���4����蕡1���n�Ƅ17$:D���JR�w��,�P�������#'D���E��4u��hÞ1��+�) D���S��ߒ
�Ó&Hs����/D���$׃<�|@[��R�gؔ۔F9D�p �T5(�'Ւ
��T��'D�ʢ쐧@�lUP��66���C �$D��;�&j�������?i �D7D��+�(Ӻ/�A�[)_����
6D��q�� xf$ ��>vx`���5D�4 `k�)�ͺș�eBt؂��/D��@�L�Z���ʵoʏS'l��2D�<ҷ�M!@QJ���1�@��i1D��J���
ZU���� o�"�Q��)D�XZ#�JE�d��wH�;�H�7D�x�N	���IK�Ʊ��j�H5D��r�Ţ�b�`�J��:oѨ�!9D�#�h�"'
����*Ùc�����8D����,��n,x��U�W���2G&D�|C�]��� ���D�&�BD"D��yq�ӱLx�d�"��򽐦�;D�|1�KS:��!�6-��{|��*8D�(2Չ�"��լD:=N��B+*D�(��(ۘI�����B�.!�O6D�r�Q�
<�s�U3{+��DA5D��id��?,0��k�H&x��sP�'D��)0N�]4L��@nH�O-���'l%D��;��	[[�m�I��ي��/%D�����<U�M1taљ|�b͸��(D��[�H�4�ИA�_�a42�;D�DӀM
,-,A;�/x �Wd,D��P��<�h�����vn�	 ec+D��r5���+Kd�9�B(7��}��&D���I��&U�P�aK��E��}@g�8D��K6����
L�8][`J�S0C䉫(��L ��E��
M�Q
:(C��,�&���+ Q��m���	9W��C䉂ae�E�ڱ7�P���嗇�C�	
/�:��r��xZj�r��A0�`B�I)9�f1��"���� ��� D(NB�	`ԑ#i϶?3,uxd�ΰQ�B�Ɏ9� ���E*?�F	�(H@�<a�h�8�Vi�$!�F�ik��f�<1M
�Z�`�1�O [L-��Uf�<yad_�q6�1`�_�n�$B��e�<I��'f �����L�c�~�pm�V�<� �7(�6;��Ð��ƼX2s"O �"@'�?�Y�B*A��PջE"ON�g��D�Z=)b���vQ�("O���TIT�"�La9&�@�LG2�z�"O� 
�	��<�l��rbա\�jt��"O`�j�]�-�ꀡ`hX�f��0��"OD�C�D�p<N���G*��"gA|�<9�_�HR�I2S�S"T�z
U�Yu�<�!�U�~�Xw˻MT�c�/�z�<Y!%�M��]q#��"R�c!�x�<)���/�$�0I��u?ʽ˄hz�<��C�,\R��a��8Z̔k�)@�<�W�ߔ0�j���G%`�X���	e�<!���	������7�4%;��W}�<a��G7.�1�7H�(����Œx�<)��	?�P�;�参=T%��'L�<��
 !JP��S��S L���+D�<��F�|��<��%�5��5#��_�<!v�Q[+�u��� }�rX�'+\r�<ywAL�������#�e�<���u*L!3$v�]K�j�<��`��l:p@�
[�r}<��	�{�<�G���J�`�ҁ��.x=�����_�<�f2C-j�ȥ]�u�:=Y5�BY�<����D��p�� O�^\~�j0�q�<Pg���Z�J		WL�P�_s�<���	�@3Ȥ����Kn�+�fSv�<yU���5�1�� *��=�T�Xs�<!�H� A�����l���Q��q�<9r��Lh�i��"��rc�J�<a��ӃxBh0�倒	A���O�D�<��H��q� S3�܇	��i(�C�<��˰�☻�N�B+z��e΋@�<Q��E'���g�}����G�`�<��'A6{��$A	�Yi���p�a�<�bJX�����N�
tz�Aԅ�a�<Y�GN6%��H7B�}�Jh	�n�`�<����fx`����a~\1� �C�<y`K!FC�Y��CƓ%`"=�� �H�<�d�8F�t}�EȒR������Y�<�t͉KFL�+S�K4�y�D�X�<!sFM����iJ�{�����X�<Q4O*e����դ-�8=��hSZ�'�R(���>�' �l�̄�Xpb��L�2��(X���훁U�t�����jmԨ�;]�Z�C(I߉���Te��.��ԝC�A3;~�%�f"O�[bM��g��<P�A�	���+�[�<���"O�N!�&L9�0<����@M��9��R�E�$�z���@X�H��(	�AՒp s�A�G��)	e�O�/����5E;��{�'e�a;an�0���b,] f�P�����
P�Y�r�̂!��8��HZ����ɶ�Q�9�dH�H؆N�xB�I�e�N|��)�>:(�H�_2Z4Y���{R��ש�O�����t��yҢ�
0+j���ٯgR4��N���y�+T�(h�l��EΌB1��_=B�H�J��NK�)[��� T���g�'o\4�!�G2lx=Q��H-Tպ�	����@Q��Y�\5�u�[/4�ܹaꇜQ�v�ps�U�"'��F+�}��|zAeF�l�@YSbߣu�°�v-,�I�p,�\	���YE� aE�)<�6�?ѐ��g\
����H:�Ƽ�.*D���VcR*6���ˠ!A9��0X�-��/�&�`��L����!��MG��%h��0H�u�$H���ͬl�2�0A�(D�X�O�s��6��B�$���E��M�w�0B��R@��⸮�X�����U�`tu�0 �w/^����4lO�"����>����|����W"�4Q~~�j���/(�%�S�N=?�bI���FJ"��T	ˆwϐq��1!mRc��AgDX��(��fBl��<A����3� ^}suo�.d���"���J�z'"O���D��-h��%��LQ��^=ZDND�܀�L�XO���ŃEd�>-�X0��6�R�TB���=l�rՄ�L��M�+�=G��ʑ���p��UÐ�	1��q�Aш\��
�&M�?�>Q!�V�e*�x�&���%���I���K�'�L��U#X!�$ő���QLa1�6S(��EB<ٰ?qW��^���+��V�^���@�'%~��a!���*�i!���)��2��q���9zhpQ��#�y��A.�^Y��]�%�H��t��~��ʟ@m�-B������S�m��ࠁ��$`qΙ�PJ\�U�C�	�;�Ҽj�G��r�:�^�?� �-�0�jqF��2 ��	)	fظ�U'U�Jf6��V䍶y����dN=$$�cG�� �遠%ߘy��M���-pDlp�	5F��Z9*n� ��U2�ȰD|2�֨ �])C�)K�a�T��$@\H"R�X"lQ6&E!�Đ%U�BCV�C�(��M
����	�b��E�?E��kQ����'hH`��y�R�y�O�IԴP2nԒ,| 4��Ɓ#�yr�M�3*�uq�����.�0�Ć�X��2P+�bt��ȓ�J䱆ȓF$D��b�^:Y��آ"31���ȓ1rP�@�D7o�8�2�Y����q��!��9�:���џ7�2�ȓg�]�2���)\F躖̓y�*y�ȓ���R��~����Eɓm�愇�iK�0+��.t�6]Jm�/T�Є�P;�EAQf��-�"U�5#S�A0�p��Y���E�gt�)B�W�b�v�ȓ;�с�G]�M� Ő��>� D��D~�C�BΩX�ʼP�,̣&h]��.r�L��n����3Żt�܇ȓd\��ԋÍ�\2��cX���h���d$Ĩzi��+1�	���*�x[�.Y�(�ǉ8���ȓN�h]:�χf�Ic�Д)u���ȓt�j�ў&Ǯ�!&%�4c,ԅȓ=V`$�b�ֱ`���;f��fz��ȓ#(e��?a�j\���̑R�(��ȓi�ȅr��If�cg��eE�P�ȓl�n��H�'FtԨ�1��h�%�ȓ3���蜗`�N\P�v0rY��>��C�IR�aE
�+qr䘆ȓ,�bD���ڱ �ȩ	E�ťW�Q�ȓe��� ��Q�~Ѓ�I���fa��J96)�"��3��{�eD�,�E�ȓb��-�D������/b>���tr`�RpgN;r�\)+rZ�pWPȄȓG�X���-�>)�������bzF�ȓ�r���-5�>)��([�&іE�ȓ3b�
��ӄ<~t`�3��<��D�tw���p1+�!Ѱ����-D�ر��ˠe�<�(�D��j�8�t)D���3�V���*�)̦F�8��v6D��p�K	�|����8lYaS@3D��bė	#L��Q�!�@��s�3D��K�-�0kF\ÄF/��c�>D���u���A`�=h}蕁d�!D��s�+�'�&x���%C��)vl.D�Pi���7��x�&�X�*�u��*D��
�]����%EpH�}*�(D�챁�̽i�<��4�=��-� 5D�h	��
$}"���K?�i��� D�� �#�FX���6��d� D�쒇�ҾK�bU)4O���M��)D�� ��h�Z	�����"���Xc"O�PI��@u��zVd�17� ��"Oh<���R��KFJ8��$"O��z6Ę$!�x5:E�~�V5!A"OFt
��\C)�д
�.s�4�2a"O`�P�U��8U2����*�"O�|�DY�$�~�St��8+���D"O�����)V�jZFOVg�f��"O�9" mN���)�DܐMRP1h44� K������M١;R$�!):D���!��1$�Y��רJ �Z5�9D��*�*�R͖��V�k��%!�e=D�H!Ǎ�3Mu�A��
�:�>��An9D�t0�c��UqrH���BH5D�4��Tb�RC#�5nn ����2D��Bv�5n'�A$B�2B%��1@;D����S��e2+�)�q"��9D������,!�8���BI�����j4D�tPD�5��b!�+��4S�%D�䊁�5�,���nϔ�	��%D�Pk�,�}5V��̆�UE��q	%D�0��K�r�� (���_�,�r�#D�8Ñ�9k�)�d�ߟT(<�p�%D�4��j�=��	�@�%~�����E'D�蓑�.EX�e:ag�5R��ǁ%D�����W�� <CP)ٵ#㎬PD�#D��q��H��M�vf��79Z8�s�Bh�<��(ϐ<�.`�@S�f�<��1��a�<�G��JCr�
����D0ke�]�<���3$�,}"q��vlt���C�<AVHQڼ���c�8/�8sC��t�<��.�W�0 k�;�؇�Z�<	�%ӝUal!�B\;;��X���n�<�rD5-��c�M��f�� t,�_�<)
J7TT�Y�PY�1BA�T$^D�<	�M�0F�t�C�2C)����Y�<abBߎ}���e���edtk�+�a�<y�'P�p�P4%�4�%s�,O`�<I"M�	4A1�Р0a�jA����c�<����Q�f������.�xU���e�<6�M�/��P���K��x)"*�u�<1�苰7�:D�ڲ>���� J�f�<q��Ϟ#�y��G�PC�� ,�I�<���<I�p,���1�d�
�,�|�<�Vf��e����!e��F~�!��	�z�<�E�N�3y��@e��u�-pqņ\�<�,N/ x�ThV�`<������f!�dڰ�h�gŦI�J��I)KS!��
���N�%[���1���1T!��-6�����Q�#�\�gn�Gd!�:hV���ǫ4f�dD���Y6.�!��t�!�eDى ۚ���ƩcO!�$۫�,%��a�8�p�&A�'B!�_y��AY7x6�s�E-+2!�B8p<�l����$z��1!%�B!�d�H�l��,}�ՒE�^4j!��Ȟ,�b�b[�פ��"��h!�H��.mRB��V�(Ļ�ߵ�!��2ra�Xb�@�!p��k� = I!�Ѳ'�l��&-ȧ?����R���1 !�D�
�l񷍗-v�Ҩ��[!��?c�fd�`�ְ5|����H�b'!��-
n����A c�f�J�M&!��A��ݺ�n@5���d)�%!�� d��Tb���鈲�}l��"O���� P�P��jTź�"O�L8��%:��A2���r6v�K"Or\�5 E9��-��*�UDJ���"O��r�ʔLAV]@%K�~���"O��e�%����Q�^�c1�[t"O�1pÎwh �6*7,�
5"Oސ��&J�1�D���K>�)qt"O�b�o;������..����`"O��3&WQ��Ī���'�	�"O0	ZR�� jx�����l��x�C"O�q�lֱ��q���ּF��(HF"O�
b�� }�9+t��C��/�yB��,<޸ӕ���bq�%�4a��yb�πZA�𲦯��Դ�r��!�y"�����iF�����E��E^��y�K���P��c��T����f�I��y��I���ߩu�<�cAI��y*�1�rc �'_�`��Ή�y�X�;q�j h<n�9��&�y2�1X���5nU�X|0���G��yR0�q��0L��B���y�,V�?���S��A�����!���y�G6-�����W�<��p�0F��y�As����ҞG~`��t퐃�yR�R|3�5���./�"d�5�y�(�+9{�a0��L*�4)�0�Ց�y�'�e�=j���;�1�0�A��y&Uh$|��#�S�8N��y"/��"r��;�]�Eoٹ�y�bϾ
��P�1��n,�ԅ��yǅ�N@l��׉����GB7�yr�ŁϞap��:|h�0�&̇�yBŒ�=���
GHPy���tD
��y�C�=�};�$�8@S�a$��yR��dVFdАb��>=,��mϠ�yB�/���q���F�)`�n��yBL�3��R3��s! ���%\��y�"��0�.���B�q?��[2LT��B~\Q{�GUQ&%�b��*��ȓ?�na�pb����z��!�l݄ȓv��0�$J��bZ�]�d�9T ]��g�lEjRI�8%�tO�y���ȓ	��8� �0(�ũ� �\�bŅ�?V�%D��0���g�
�pȆ�,Kt���I�sc����)?_|`8���R��@E"g`D��
�fe���R�^��D��
��d0���j_:ņȓY]�IA7���vwޘ+�+�L��X��V��[�h�kw�}�W�=H�z��ȓ4�m����|<S��Q;L6ч�{@�%K')�:Z���޲�&Շȓ`xp�`7o�<(Z}�#"p�p��ȓF~�Y#��.����V�bnل�}�V���Z�3bāS�+A2Bƨh��?��Has�˧6�@!B��f8p��O���偌�g�����.Tq�`��ȓA�`Y�#�3{�.)1!�Ia� ��ȓO�`l����D�9��L���-�ȓ!����P��ިKb��i��ȓ[��Qg�.G�L�c`���q���T���]��[���>nݴ=��;��ͨ��&-,E�E.�9蠆�!D�SA���B�"�)��*j�Ԅ��S�? �딮E>&�MIT�ڶ��Q�c"O(�`aG�@H� PF�M�NxT�FO*��ºX�N���$VL�p
��ѣ^!�dtV8��-��-̨0�kC)�!�D��I� I�#U�"="0yGk�0�!��ƹZ�T	�$ �[@� �F*�3F�!򄚻�&h:`HΚ3'LT�	�<�!�d��U�łGBZ�lj�E��Aí�Py� �U�����iIx_he�%���yr�̿a�VX9eH��<8v-�yr4S�0���!؆	<���j�y"��U� 2ƀ���,�U�_��y"_.@�����!���b��)�	�'�h� �G/#��C�ŋ+B.,b	�'/p=�F雃7�, �Fǌۢ���'V<����R"�X2KH2$�;�'�Ld�C4%3���v�U�#�� i�'� L��	��z(R�k�-)��L��'�H�b�Ε��m�� F?�~)��'��0�B��Z�u��+�~�l���'�n  ���&B;<��%Kԅ{ntp�	�'j6��pA�*����B�"�T�	�'�AӷFûa J��E�!N�q��'M<4C�A&�}RT�ٛ1|���'Y
��:�r<q�FQ6�`���'q��B[�k�Ęq�-ƥnt3�'���n.K���k�o�0rKص*�'X��FH�=xH,Ȣ�(7�L���'�ٺtfց&tθjgG.'-,�'��9A �Ys�c4���g�=��'n��3���(rh���b!Z����'{F�Q-�'Pc "(H�J���'s:E��Mx0&� OZ��"�'3,�`&�� ��؇"r��#�'�����%Q`��)d$U���P�'� [v�l�H�L�"LF��'KH�ZC�6T�D����9q�B��
�'<��F�ܯ\$`�2�Vx��y
�'�(Uॄ�M}2�X�% �H?:�`�'Mb�Scl��GY�a�U�Ў:�ȥ�
�'X�h�	��=u��+Ԯ�4D
�'ފ!��"�^pH3V.8i�e1	�'�h����؇&��LK�(�*���C�'�X�30��~�)��(��DR�'h���A�>2$���0�ċ Xp���'}"1p���j�T��0O��fO�yr�'#��{����d�A�N�e�8щ�'0�偕��
?p�5�мK,DZ�'IZ<��C��r���!ߌy�88�'���#P�[-4��wM�Hޒ��'��!&���2�60XgdC=����'��"�#ޏ Ŧ�v+�)Đ`��'��$&G2W�dsvH�(�ⴚ�'���i�����Q��H�8W*y��'	n	!�5g�:$����8F���	�'0Lx���.pn���M�Q��M�'��q�U��F���&�L��D��'�\)�	J�Z��u"�%z9��'ۺ��R�<E!�#��M���Y�'m�ԡc@4n6dXD?}b$��'%@��F3wSl�R4/LIɾ�3�'l*�������L�� >��ݚ�'�x��t< {s��'K2��
�'8H�P�ęh��|*�
�.؁
��� Ҡ:O�P$q)��	�3J��A"O���!,�c����˅?�4���"ON)���7=��X9sD2��d"OXm)V	��*6<� aΚJ��i�"O2T�� _3�)@/�g��]�!"Oj8�i6r���·��$ :%"O�Qa'ÈJ|��� KkZ�Փ�"O�P�ȇ)zY��EB���Q"O��8Ҫԟld�UA�-�]*uc�"O.� Da��*��(�1�N�N�i��"O�9���8�1�E����� "On��rm�8��
���<x�Hd��"O��ׂ,��]�r"̠[���9"O��D띂M9��S)2�����"O|(���1XtH���
�  ����"OZܰ�!H:"6�����Z�%�4
�"O>�C��"G^�)��6;w� S�"Of�P�	��±Z O5R\�'"O�I��T����:[�@��"OF�-����C�L<\v��"O�(� ���.^�,X���"OX$�j�>���J@-��e<�)�R"OB�@G�&�,�`��0:���"OZ)���+Z��d`Q�
n)�"Ob���F��,�Rܐ��X$�*�b"OF��G����j�j\-���[%"O�	��!��	�\z�j	�0�e�"O��c@��n��!jд��X�"O
�Ҡ	�pX$؃�h]:(��}�2"O�<����0m|Qc�l�LB�q3�"O6`餭��GF�E�IӗP7��i�"O`%s$�R�qz�����?�@� "O�U٥�Ю���0�E�Xm�x�"O|E2�#@$9.��-��]y�sE"O��)qE��f��I��F0��4�"O���v苋f��8�e�pbN�"O���tB�_pt��td]>k�=��"Of�*U&�V� GdG6\����2"O ��GI�p��1����T��"O,@��g]�<�>X�E!-"���a"O�	`��� R"��1�o\*9uPQ0"O�a�C�U,�u���Z��}`"OTA
g�&_e�QAX�@�r�X�"O��k"ˇM�Q�ԗe����"O��['ءm�$���	Vd~��"O��tR;z̚�Z���	U����T"O�@9�X/I�xC �6Ir���"O�QSC�Z��֍�2=�(9�"O��!��t6�%���E�w�D�3R"O\Ypb� �A!Ǆ�A�: "O��B�=mXijkݷ9Ŷ�B"O�E3�E�g7:����5I��Du"O,�te�3E̸��&^=��	"O��@MQf�4I�M9!�\CD"OIj��1��P�&�m�j,�"O�1�v*�+�Hŏ�U����"O�)�`��*Xv}�s�ʂ\�p�2�"O��"�dQ% �6�Hj�(��r�"O�L"eEM�H�F��V�9�HT�b"O��N� #��(���R�\�N���"O ȓ�C�9�R8z�(-j��"Oh|�q����)J!k��Q��q�"O�$�$I?���%�NP���b�"O�������J��8�$�/rt\���"O� �X �c�/CK�˒�3RH��"O�Q��7΂�0%�� :6q:�"OJ��aOS�Ul�X0Č�'w�.�`C"OdPU�¿Y
�i��c>�b"O�@�f	E.d��(�&��\}|8�E"OF����W{"�IӅP1�$�"O�T��(��%Q�x�rN�/x���"O��Q��C\��P�1p~:��"O������gI ��kU����"O��4mM�~}�IP���B� ��"O~����ѭ~��i��+Q�.!�9Be"O(����@2� �G?6���"O�y���\���u�ň�;��� 4"O$�pr(Gz�,|��!C���"O�A+�	����33��ye�1D�\!Bo�\Z�x��� {�(��.D�|P���/(�tt�p�U�k����B�-D�\�c��
3>�d���2R�h���6D�X�JԨo���p��w�����b6D�\���^���Z$kDRy �.!D��T�!Y"&,����cQZ�	5.4D����k_,*���nʇ��̚T@2D�X��J{��<�R�	�<��R0/D���Ӗw��҃�63���@Ə(D��c���p��ЇX8K��cU@<D���C�+6��]�$�9dF��A$9D��Ch��I���z���*`��͢��$D���U�O�JY�Ŧ�,R��!�d/D�0#dQ�G$j��^4U��� l(D��A�Ì2+MPH9w㜏+E�		��1D�pbЇ	z���Pl�]�n�s@*D�dJc`>�놆C+LdQ�@�'D��Ywb�=�ܩg�Ժ;�$c1�$D��"R��;fD�c*��?׼�� �$D� �3�++:�����A�����<D����h�,!Ɲԫߩ6��� O0D��{�e���X� T�\�I�Ԓi8D����h�aAb�
�8*�IRH*D�����
IV���Ǐ+��O58!�$�>=R­․+Y4��s/�:�!��u�쭩#�0g1`����&B�!���.�4e
��Ϸh�0k��J��!�d� 0��Xjb�ֈ^�Y�'�b!��5P���NŲV��d�[!��۸e�fX�e�ύ8.�4i^�!�DM0����0���r��M�E!��
0t6FE�էwP%re+B!򤞴c�,Ay6e�&a�-S����]!�$ثS-H���ӑV��)�ˁ�D!�D��#v5�'HD�lv]�䄑c!�''�ƴ�!է�,,�L1�!�d�_�|���[�px�5 eb�<�!�dV5|<,X%K;ɨ("vA>���l��(��}��?5���ԋ^�Q
�� "OXP�i�r zB��U�8��#"O�����m�2`�#�v�F)"O,�D���&�|,)��T	W�VmR0"O���� pʁh�;!�H��`"Ol�cT.��FP�������x�"O���S*�6�u��&?�ƀ��"Ol۔��^��E�?��<O!���8\�d��>uT��f�YW�!�䗎����j[.9�I	ah�?��z��dGK$|·֣+�}��"f�!�� ��r�S3_� ��!K�aĶU�1"O�P%���|�9�t�B���Iҵ"OV<sD/�h��XQ���b���BS"O�kBbH?3���!�φ+_����"O�
�B�/�}��B����:"O�H�­ԟ|"����o�zY�&"O,YJ����,۲��F2Zw&�1"OVLP�n�����H1)��ZL��"O�����	�����N5Y:���E"O�J�cɹR.�T��!a/¢�y�	E��I4f
�W��� F���yR���τ9a��R xD(���yB!_�2���`�Q��YJIȤ�y¦STf@�T�/*u��!�y�E��MH�BmLQ��'�y�%P)@�!Ѣ �3���Ҩ��y�ꂇ3�.������w�n0��%�0�y��UJ8=���]�?�p��-�y�K�e�9��M"�=�2�	��y���*�`5��M�9�^a�G����y��H�6yR�ʀ��8�Ջ���y�N+lbn�c"m�tٰHq�i��y�C�C�Jp���l�D���R�y�.Y '�$hpg��l��=Cé];�y�(!��C��9T&.���Gߕ�y�̊?��M�wM�w�4�!΀ �yR�߸Y��#�cHp�f���a�*�yrȗ�6M���ǻeXf�2%���yb
��~XM��L mL�=B�à�y��׶��4A�
^��;DC���yr"U;���i�$�òq�����y�'�^�p��7)R��,9g���y��6q%��"�Á>�JI��%�ycW�!`}PV��)s�+V��y��R�[�L�����0W��`��
�'r�Ѩ�Ԑ!�*B  ݼ�@p��'r	zA���]� �����,6L��'�J� �C&b�V�SK�<k�f(D�<�W�Ι`B��s��;) �X��%D��F�6� 9�e�+/C��2�.?D�,�
� f�|[P�%D���H�:D��X�&Ku(��A� 鳁8D��PA��K^�;�#�z%����N7D�dV���LdcW@ 'v���*D��e�u���sЪ�o�<���-D�@�Q��2LՂ	�Ǯ[�`�kCD,D��c���V��<eI0\,�s�I6D���D�(t�ܩzJ�?u��}���5D�0�D�̰C�h�W#�+i1�E#Cg5D��P.F#tt�K�ő1B���$')D��*T�ƚq~ T�m��1O@�!�&D�h������ i�ɄM�1E6D�$���ȃc:9�D��Y.��` �6D���"AR�%y&HWe�(��2�/D��HV��b͸W�̋�̄j�" D�@Q�j�1?h�X��k'4�تF�8D���F�1$Æ���Ζw�(i�*6D�Iw D��&-z��
:X���9�' ty8pN�= o�l��'l��19�'��T�z.��ER�}���a/�A�<��&F��ػJ�*�"���v�<�� ��P���'5"���!5cCp�<	V�6#`��ů&>��enj�<�k��a�M�䅊(<�Y����^�<� ���,	� !۷"M�~~�Ļ�"OP��P81�$�V�:`t Y��"O01�E9$�z2�S\d��V"O�c �I�Y�.���jT�	Bjs"Or��蛍;w0��El�V��p�B"Ol<���N�E�X��wk��$wL���"Oj谢kO!t���p��E;a��T��"O�ql�n:ƕ��N(.�6��.D�L`Pa[1_�\��ՀZe�X�&A.D��3�TK5(t���¢,��p�Wc,D�pj���8a�P��(K���3%�5D�$� F�1 W�y�eF�0do���O(D�D	󡐂('p�2��M�F~.ʔ3D���G)�)Y�j �"��� &�1D����cE�4�5#��F�d��0D��b�K	Q4���G!�}0�)0D�P�fL�0pO�}BB E����a�m���$S�1���iayK�7��uӥΆ�D��5�'�L5�L8pPn�<V�l���iP�Pk蟔q�����@Y$/Y! :���5��V��0��t�G�M�jt��~R���nGF�{��~b�X�X�JMTb1�P��X���D		u���dN��1�[?˓)͛�^� r���؈ЛaFҠd `ҡ�2D�$h2��1h$��e��q$�]��-\YD��eӤ�O����^�^Ǯ�1��͉1kԤ#�-ѐh����UL��wkR�@���?I��?�T��	�?���?�e�Υy1v)r�A'�����|���@���2/�F0�1.��|��ݸT�i��+��$"d1��e���b킵{u�Ջ��
� �vEA<[�`9�Fd�d�HુM!S#�p��l��\4��mr��D�gȘ�@Dc�O�(	 ��̡4  ����K�Iڟh��u�S�t`P(��l�c�K�o�Ւ�I��y�.�8�f<�!�g�.�����~��eӒ��<�V� `$���'��P?���H�]Юhwj�S�&���j٫O~E����?1�5�H�c��p���J��=ꐬ��(&�-�S����1�UO�}��c��TI�'L�y��59�Z��Vm�I��J��Z�	`,�[޳D�MQ�I���� �v �%D<�Br�|R" ��?��n����'��S|uT�����p��JF�0���V�����u���O� �ߠ:�@���чx�11�e�g��TX�4[Λֹi��P���RU�xy:��Y2j�.㰩���dW*K��%��ԟ����?�aD�X�I�A��]�s"����_�y*�e � ��K������z�'ϲyc���H�IK�}�)�B�	h�m���'���l	�S"Ġ @~�D�H��#A�j�hr(*w���ug��7G��S��Ԓ&����[�R:{����A�I� �G�H6-:{�R�a��lZџD�O���M�	5O�J�Њ5mҶ�
��_L?!��°>���O:Y1����%^�j2��E�'�6���]$���ƺs�aW�m]�(IS��:�0��7��W�R�'}��E��b�'=�'� ��lnZ�z�N$2�ðw�5�v�@�;�����D?���W,��U����A+��+G�L1'�Y4'ѝ!d0�Ch�� �v<�uE��M�ˇJj��5���O7�T�P.�# ��<�v�O���NRW��*�&�&���ߟ 0e�Yɟ�y�4F~��gy�'��ɔ7XX�R���(R��1��q��L��'S�9�������@�I�p�|Qcݴ�M3[Xu�J>!.����@�gD��*x�b�'[B +%
՚8����?����?iv����?Q���?!ձ^茝ч�4m�^�$h��4SĲg���5}�D�����I�3��	F�	P�2P 1NҳG�9`cA46�^Xj5j��n:"1��c�6y�����5a�f͒E%R�j\ �%�ĚE��O��a��ك�4l	��Ȼ,ϒ�!ҋ�(29��lZƟ�'9"�'/��	-iQ�0�DY�W�
��7FRO!��[�cj
8b-���	�d�,4�d/��-l}�	>�u��'y�'|q�� ��GF2o�.���Kϫ����%�%/p�5I������u*�=_�M�rǜ�7^��iq�'�&��fGN�.Т�`�#�'<�z	��n~�h�ҍK#0<m�Sl�N�(���GO6-֪�@�Ó%9�b=�$쒝l��D�R��t2���*�>y�'E�P:���G�Rup���!i�|�3�U� n�p��fr	�놓8�F�IbF
G�Ta8��n�d,�CJ��!l� `��ϣ]�������V8!AY8�Hã��=
rDa�نi�Sh�k `Y��tk���ׁ��oGV����n��87���x��dĹh&lqp��
q`��O�@H])��mPe�-h�y-8�ɶN���\2*A.�!l�9W4,M�Є�Z��-�R���qC�<�
=K�+G���V)�3�^�S��0Bdl�J$!X}x���W`6�b�����Wp��0��ȭ{	@�)�k��^�n�(ՇY	&��̲��Ğ0�v��EVSy��«Ȭ} P�0Qa��m�HH��JΗ4�ȸ2ǅO���(���|�y�'��i��sd�D?gX��я�$|R�B�f��D�H�sF�T�r�)"�Įa���n�=bV���o�59��p3�V�Lg����*B�z���[�B��MZ��O"L9�vK�S`�XQ�dZ��th�$�?V�"Q[U�i�h�b��*��H�gJ]&o�r�"`�5*�ɘ�)�D�	��JE�jR�T?j�CV�� �Y�t�P'�_�}tXq��+�Xy�5ꆌs��]�w�A�0��d��v�=�ׂ�	2�<5+ ��DB��:��Y�z'*�#J�3��<	�c�l�VՓ"䀂zzX�
��V6N5�6n?,I�'�-���Ku�Ԃk�N�Ӣ� ~~B�
����j|�pu˗*yJ�)���T/L��j~�@ M܇T�*H3��|<�˕�����IXu�B5Q{���'���p�]�l���e��}��,��@ۺ
ˢ��w�W�N���� ,s��-�Ǔ^� �҃������$߰lw�yt�U,Q����éj%��`�@�D�2!%��%b��GD;��B�G�r��R���'VA���>s� �˷C��!a]�J�0���'D��d�++5����N�w�dH*`��"O[&�ʂcЊ1�6U�Ӭ��x���p5#6XL�p�7;��e��oM�'2ph��$�ɦ	�r��6bT=���=,�@4�M¡.���S�F�!%�x��.�7�"���2j@zB�>)�J,(��b�q:4b�:_t
��aժ,P"�b/ʓ.�|"H:^v�?	�$m�S������)kF��Cq�ޘI� \����ܐ�dZ?���4M�R����QɌ+nL���+�L�@��ŕ\�P��!i��!%�,��|_Zy�E���@`*O�I"01Q���"J�ԳB
�8"�䘑��f� �����=Y��b-ϛ%�S6��r(�˵�ɻ$����q{��W����&$�/0������(���ɯoA��2c�m�V�M��S��ɒ��X�6��5�&*���� R�/Z�Q���hC�p�R��H��;��4BU�3��\"GJ�9��#<��P� q)JRV ���L��^���R�q���sG@E�i�ؔ�H�3�>%A�i۾r@ ��(L��D4�0�Sr���['@��j�v9�b�m}B�
 D��t��ӎ}�k���E�EH�+RC���i#�&
���\+$��2�ڽgiP��c��Hd�"�"��G,����Ů>@�y��W.w#��
tb��bbJ���DۓBp�qZ�@y��B�(|<�����*v '�B�:��B�9:�,e��bW�pY�Hq����yiB�����D����*��5��32��.BD�\1a-j�mS`�='�\�B�D����R!�]7��O6��ŉ�N���s׍>ut����]X���T��8q�>�7G^�K81�u%�N���[��¿w~�%۴�S�\UJx��m\�m�\ ��/͗`w4y[�}�ԕ�v��"/��`!6�w�.��|a���42�@x�M		�!���ESSb�C�H:	��d��@�2o�Bh@e�>1f��󐩊�-�vhDV]~�S�I���L���B.hr q�F/c�:R�Ū�(��<A���>���g�%j��)�jC E@�
�I�ip������޴퀂iT�9N��:��	�-�Dc�m[/�^��c^*%ؒ��"��O��򉔯:K��2=�.1Y�CX�O�L���(�b2��pM��a4��T�E�|�u vc�:V��M�N�S1wx@�&)��q�`E� E�<h#��#(m���A�S��$ r��6�4��)(r�X��$M�$Hs3��D*?Ϭus�N߰DH%�c�?#^��c�۴1��=3DQ Z4^-�C��*>΢mS.��CG�5#�?&D��s�X�0�1�`�^�ZF�sa/r,��`�m��	����Մѿ#
��=y�h��h�#al�m�E���O�"..Ej���"$��c�5i�lS�&cB0z"II�2�]�v �� )"Yb�@eI�4䉚Ĥ]ہˊ�?*x�Jt�۩rt���� �qO|pQƐ_QZ�y���"B�@��sDF2i��5%իf��=�V)�$h$iz�(@3 �r�k�l��]��AӤb�ˡBѩc����^���)��A�g |ت8�f,U3J�n�g�vG����i�Z9�Ԏ�xn�l���"yФ,�F���w��Q��I��o�ܙ�B�CL��uڤ,�@�i���I(����ą���	�n�܉��|��DE�t|Ґg9|#�p���$�^\ƥr܉�b��(��yq�O;:aЃ��>���ɻ9c���"�Ra�)mQHtJ�K�0��$y��� .
��&�g�'':-��Hئ=��ETl��jшX�89`J��0�V� UF��U���k�Sy�C�c�\�2-J���LläL9{��(�@��1�N{ ��p=9���#P�� �#��0���#�L�;��iR�HH?i��ǃ3}�j5}�̣1��':`���W�8ʧr�n�SlC(����-�Ky�i�=���$>躈���c�"|���#� |8��Bs��A��
=�:�!BK���$ڮ�T�?ӧ� �U�m(b�~|[U@DnZ�ʦaY�#�ܔ
&�G7��F����ŋad��4�� B�8�e�=|!�D�d@;�IʷAu�Bd�QmR@�0��p31�g؞��	5v����H�
'Fdӷ-�O(�����y2�@�z�N�R&P�N�((�����y��A�j�<if�;
(��`��yrBč@�,�x@(�+.��Ћ�y2)�p�����X!�4�PNU7�y"oT�J�"�s�͉=:L�B�	�y�#W<y�@���	�gb:�y򥎆a4�����䈁�JN��y�ǃ$���y�U4\�@���y���2�ju[�hB.}��PՋ���y2��O��C�~��Db6o'�yb&�
��qK�v��A��^��y�'��|\��a�߂SEl���-^'�y"�L+~�:$x@nI�Xb:����P��yRl��r�R"��M����3���y�L�1��4r֡��FH�r����y�"�8~��0�Uc̟�X<� �؈�yb�5W�$���Oɧy�V���J�yBn��y��H.�c7��wL���y�A[#-�L�`��(Pr8��i۴�yrn�4G6�LT�R�Z9˷��yR*�0N9^(�t �J8��+��	�ybDH=�tF!F�x�rg���yBj���܀{�̃@V�%��#͗�y��ۂ`h�|B �
�k�8:a�P��y"��+��kt�G���dP$T��yb�N�.3n�����49��@�N��'6��8E��7v��x��G*9��9�yb��*���8A��)��k�EJ�=g(���̦� E�w��L��O���s�c��M�bIɐ(,h��!v�_���y�I�)a�%M?1�a��A�<|Ɱ�� ����К`v��0ყ��c0/��*��	N~�S����1F������R&z���>�k�YN?�"	p�N���'g�á@֕"~���Ç�'"ќ�{6����ӽi}�x*��?�˱`��?ŋ�t��ܜ+
�b�Axh���3F��ɱ� ��Fa2��� �<9k��OȾ�,X��p0AA�AxJ̹�̛��k@� P����0|R�B�S�x;��<��4PA����� �z�^Գ�`E�Ք��c��-��?=�PbW���Ah@O݂r���!���$t�Q�X��) w�Q���	��:�8��W
"�V<:gb�w���IL�P��Zļkç��� �.�O.4�
�W��]��u8�|z���0P��/O�>�`O^�p��u.�L�iha�4�I
�HOP�Ov��I��O�D��b��ږ���"OzLR�m�I!,P�π�tX���"Ot�I�`C�w�2��!�M�yF��+�"Ob�Rŕ�@�0M���	��h	S"ObqHx�N�A��5���H�"Op��a�%g����� S��"O�5p�ѐ��:�&��JP�"O:L�$\��P�^��`C[��!򤚞=�&�9)YOe�i��K�!��ֿ
���p����u�p�qG���=�!�J�c��9���C�, �3ˋ�l�!��@�"Lib�\(�%̈�O��Pj	�'l���V=e��A�匃g|��'b���͙�8~T!Gf���Z(��'�4�J��A�fB��hcN��
�'��H9 
��2��m3^aF�
�'�=J�
��̼�2CB%@�8Ȇȓ?�$�i�ٖ-���H\k��P����i��WB2�/�V�<��ȓo��\����G#�d�[=Q�<�ȓ%�l��a��D�ȼ{PF�6H����Be���I9�f`��I�2Y��h��S�? (��@�ыF?�XI�k�1L��X@"OYcvdD�B�>3�埏@���"O�%��hN2n��!B%�ئBfhz�"O��E%eA~@zuM��zM�}KV"OP��BU.e�8��m]�3HH��s"O�H�.F/�"
_�vA�iQ"Ol��]�����Q��3G�<�c�"O���G,�F}��fʔ!�N�H!"O�z�I�8O���Wϛ�&����C"O,A{��0@�X��[�I���C�"O�ٙ 9K�|�:�LM(��U�"O��q� �
��8��(`h�\0a"O�$*eaH�l´c�-Y?No�x�"O5#v�O)Z��	3fZ����R"O��X�+]I�T:��P�sC��Q�"O�9ɰ�ȃ. �d1� �c+^x��"O�-�G�S5��[��\�X��"O�5��+�.��@��� ;8{Fq�A"O����A��22 �1��0�"O��D�ΣV>�LѺ�R�'�R�<I�g��g�R@pVl�j�F��bTM�<Y��݇ctts���uv:j���I�<	��5s����Ҕ)a䑱`UC�<aR�Ɛ;�P)GI�~Hhq1�Y�<ђI��KX�4R-D���D,IY�<�v����q�W*��)b���R�<y��3g��	�fՆL�M��C�u�<yg��-��и�">b���hf.�x�<��-T/s�������+s�] cKr�<6�����4J4�F�9t웡�g�<	�k��e�zh{qm��y��Y;��{�<y���?PXd)�.�IS�#_m�<�^�(M�]0����VPyj�+Dk�<�@'�P��V���q&�d�<	��ɯT�`(2�Ǌ1e��m��Tw�<A���kA������T�n��׭_[�<)��M�J�;@`,c��Y��P�<���@6e��j�M(*Ȝj1�\Q�<ٲ-�4�H���U���̚I�<逥K!�a�g	�0r�kĂA~�<6φ�$W^ݒ'�D�؜�W��v�<�g`ڕ?c�	J�L�Q�<� bL�<٥@ֶ�t����[Sӂ��F@K�<A櫒����s/D$z��p��PF�<�&h�����q	�>vź,H$C�<�,�� �ۡ��71+��	�|�<Q1,�?�P�"��+AΦ�Z� �{�<ѐ�"<	j�,]@񣔥�;|��C�I�Z����E�?��Ǝ٤[�FB�I�2�`-cקI>�6���/Y�%��C�I�3:�3��1��yib, i�C�I HHYQ��AT��J�)�
jFjC�I�p�� t�g�Z��^�txVC�	uqj�	��'^
�Q)a0~txB�8p�����$^À�
&d!^�B�I0@��Y�a�2�V�q�Ɓ�j#�B�I�etx��f�[j��%%�B� y�hy� ��%.N��F�Y:�hB�I_x.A��k�8�I���&T��B�	�n����"<.�,X:�/Z�H��B�YJ�P�\;o
� ��#�dB�IU>N�r��"��1�-��C�ɾ�"xQfB�+8����F>�C�	.PW��1���~8��U�E)�nC�)� �b�CHS�����˓�3��<RB"OVպ�:�μ!`M R�L�"Oi��a�%��٤���&��5�p"OrQ�`ǆ"Obв&\',�J4�w"O���k���,���	D"O�����Ş;���� �(G�"���"On�{�]��M#a��Me����"O �jN��hVx��Ed��f@$1�"O��
�G!��L�|2�aE"O$	��C��h����(�h3"ON��u�0qx\0+�#B��<J"Oj�Ck�J�ġ�#�b����D"O����g��,��M�k���s"OVtCԂY4�	�4�N<h�@ "O�L��"�-Gȭ8��R��]j�"O�x���̉8	��`���k�h%�"O�չ2�V�hT�|� ��9C�<�B�"O6 W�ȏ?��"��:F�,��"O cG&��rs�ak�`\�i'�}��"O@���a��>�KrAȚ^7L���"O��8�(�$+��q��]�K0@m�"OR���P>��BP��j/h��"O�u0����"	��f/КX/B�
�"O�Ĳ�J]�8�ʱ��$�!z���"OX��c�+r�*2�Y��a��"OZ���/�p?��bJ�N��mS"O���Sn�nͻv��'SlJa"O���䘐P:�E��m��|��4"ÒP䃚6����ԘfI��"O���$E�9ª���c�uX��Q"Ov�����pD�`1$!�U�xb�"OP�"$F�]݊�Ò�NXp�-�b"O�x9b�@�P�-*�*Ғ%pp��"OP1jO��&�0H�Q�U
^`)d"OJ!��IH�^ ��i�I�&���8�"O<Ԋ�ȀEBq9��zبp�"Oj9�taײVC�T C�8o����"O& �爇��YT�W�Ak�4��"O������I�J a� m�ePA"O��U�͒o��)2� G�����"O�Y �-�"=�m#.S���y�"O��O��):�!B�Ǡ
�R�J�"O���L�8H�� "��6l��ҵ"O����ҤK7n�*�"uL6��a"OV��E�T��Es2AHxd��"OH�B���3321�$̴A<��"O؍	!	R_-b�fŋ#lΞ1H�"O�Q��		7#Rȹ��P>d��G"O2��t��uPd1j!��_��B"O\��K<p\Lu�p��-m�^��"O��(7	�W"$L� PF�D�X�"O.1��%�r>h!q���P�����"Ot�a��� #`*��R�ċr��QB&"O�D��d�&^94��4��x|��E"O�="�E޾qD>E�2
�c��	��"OA�&I>�<��	�6���Y`"O�4Sq	.L�:���� 6P�z�"OT9����9�b��rm48��T��"O&�륁��948�;1�-Rp�� �"O�U�v��eȡ����M<ДS�"O��e�+ �-��46c"O\���W�a��LQ��߰�6=k�"O��������Q���1��`�"O��r��_e���bд:u��xc"O� 1�B��@@���H�)[�\�1"O��3�����Af(8��(q"O����N0=�Xǀٮ3z�)"O\e���ƅ!+��k�A)#j\�	�'L�b!��.!����#��0�(aA	�'t�����L�:?���r�\4-3�4��'����*I��⌘�9\_�r�'sR4��	ߚ+'$�SA��b���'��Pz�C�%&���h˦, @��'�j���g��K�4T���,�:`�'h��Ły0��S��E?���J�'H�rm� Hvh���#�3�$�
�'d i��E6�,T�d�.pƙb�'���ϯ+j<�9t P��B�H�'�rd��n�9A�Uz4dG����3�'G@1I"��zFu�` E��0�*�'���&���@_ =�GF^�v@��'=D��%���T�IbLs�J��
�'p"�"��,z�Йf��ewz�`
�'V$DJ7m�"!�2�����kT�PR�'�<�� \�@ie��:^�\��'d:H�4�âs����(��3j���'��y����7\�f�UjÄm��D[�'E���Ӊ�1�V�0�S�g��'l��x$��/�U���� lm6��
�'����v�[9j��ǅ3P�:
�'F�°	�e��X�O�>tƉ�	�'|N]k%,x�!/��t4�"�K�<a��8��]C�m�����YD�<�Q	�b��P��;M�D#�@�Y�<�j�����5 �^���r��]R�<	$BJ1;J	 !�	.����WP�<�7kC�Zt��ʒ!ц|8)��q�<Y�ƙ�T݂�m\�TWd��*	o�<�G�Ի��2�Q37V9S�,�s�<�tكB��m�%�~E�ԢB�F�<�@�P��h�b��I�Ҭb'mD�<qG��\��-��k��� �d�<�p�8Y���h�M �)��ENw�<!v�QP|@HCPϸ}Ćؙ�bPq�<��JT�a�����H,H(���D�E�<9w���B���p��(	�����DB�<�&�W�N�^��呢R�N���u�<���F]�&��#� !dX�S��x�<YS���(��1*j�܁Q!C�c�!��{G>	2c$0Seq�a`T��!�$	*\� �.�)>Pi���۴�!�T�_����g8Ezp:Q��2�!���8��X9\ֽ`@�CAo!��(C����/Y`�8�2�!�,8!�$��\����D�m�*D��� N�!򤞢[P���
�&o�����/C-_�!���<,*�J⩔:���GгD~!�D�h���׳C��$�Є@2
!���dE:4
�L�=\��L�d�ټP!��T/l�"��UA��~������!����d���)���;cq�"�*_�I�!��тh���I�{Q&x�0*���!��[�l@2CZ�+����'O��7�!�d�J� �  �P   g
  F  �  ]   �&  X/  �5  �;  5B  vH  �O  pV  �\  c  Qi  �o  �u  |  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�6x{3;O�1"�'"dE�>2��EN�%�D�j4Ý_�ց�Ф@�n���#!��a�w����CG�?�JS��?e3�f�x��x���4~�ABA#��j��5��Ėj��]�s�??����ƞ��u��|@�t�'oT�ɡA�T���,w�Ɲ{� �y^VxBt��O�4��a�|Lc���I�P��П`�	ݟ@�I֟0i&ˈ�	�$UyYD����㐼m����O,L��E���	�'bkۊQ1��'�r�]d��ÃN�
V��!BP����'���' ����r�R��?љ'���n�u
����j�8�^�s�@Fu�r7O.%��U5���z��GO���	�S�Dx�O`�����>����,j��8�p�F���,k�P=O%r�'��'���'���'���ɼ��h�Hy���!�$������\��4���'jӒnZ某��4J�UD�i����T�'*��i�Ę�.Af,�q�ކkT(d��+ғ?Y�0{r�7g���	c�34R�pʃ&� �С8���#4�0�3�X8i�hl�McҸi\���O�.9X�2eĈĊvF\2!������3�0��w�h�xz6$B�]t2�s�-}�����D3aBRh�U'^���ݴKl����N�vXY�	^2
p� �T9vв��4d�l�`�v�̨n��M[�%�
X��U�fov������#��#�k	s�>���,�):��:R��<"=�0�ҟ���`���n�n�Jxq��ϑ	lLq��M԰b�v�^�F�����;�|�;0����?QQ!�	c��c"�ոS��HF���?1���.�x��!�^�p��S
ݖA�����O�DS����m�h�d�U�[���s��T���D���?1-Or�d�O����$,�� �5���أbUئ��1,�v7�1�C��,_�V	bbm����]Y$�m��M~ݎ%�I���hh���Yj� �K(�X���ûo��'�VʓpS��xb����FX�U%��<H��ȟ4��`�S�'�y�H22�0Q#-��=���91d����?�s�i$��Q��}0Zh�q�G8?�iX��z�f�R�`�����@`D�c��$F��J�G6�y��TR\q�Q�IzQf���yҤ�,[4%���C $QdM�a'�?�y��CtЅ��E�%Ja!y����yRBI�0,j��#=p������yBՏ:�8��gJ�/NR=ˠ���?Q�g�f�����h��所&Bδ�%��D2��{s	6D���i�dL�*�H�MS����2D����!b*QX� �+W����	;D�Ĉ��*S�ؘ�R��hG��з�:D�� �ȓ}� -kW�)���T�=D�����.�\�!�*@KVa`�<��i�U8���6
��/7 z�EߗR�6�{a�<D�x����Vq�1�⋐�2��Ѕ.<D��y�	H0COT�Z�!)���,9D�`�c_�n�\���ُC|�=���$D��3T�� {y��B�jB#]�v��F#"<O�t��LC���I՟h�s���C?B|���4�lx���ڟX�ɣPx0���ş(�ɁeP����Ԧ�.ϻ2W�Q?|q��%� ��H��7�0<�Qn�5OFա���%߸�4N��ȴA���2����N�Otʘ��*0����OF\n������ ��&V�ř$K�_�h�{t�:?������(����QBE��qR�!��ec(`����>Ɋ������U��>|�dʧ�F�>��)� ��M�K>	SJB^E�!��2�O�8Ͱd�@XH��:��f,���U"O�#�<@�f�����8N*"��f"O�LHӃL�["pʂ �
���"O�A�`�ў��}���A(���"O���$N"��x�㈪[�`�2�"ODɸ��/�F�k2d�7 F)�bKu�ГO��C%����d�OF��<q�	σ~���-��!�a�]�J���$�i7�6- Ei��K���|ʂ���P~�� ���/�p#��,��J�]� �`�7���"�	��$X��'zNA+ O����4r�) E�qʵ�iv��N+ l�Ie��\�	ퟘ ���.���sE���`Ѻu�fNgx��P����-:QJ�≁�l.r4�#�O���W��@�4���|��'��������1	I��ir1�Qzĉ0���O����O��d�<�|''E�d��Ȇ%]�xb��y��J�2�衰��G[>���4�B�`��y�J�o���WBA�=����λ���یKCT��`F*(��t�7�G9]txEy2�W�[](�To08s
Z���E�$U����?	��D(����ڜ/4�Eѐ/�V���ȓH%5�&��(����GB�mx��$�ش�?!)O��@��@�S�)�jAZ!	F�HSCh�/4�����<���?��Z����D���0;⍀�=
� �I��@��Cm�9��ߦ_��I;��'Z��#�	�0�v�;�ɗX�FMj�\�{e��+!�ZD���Ƈ�0<)�"����Ik~��@��Qx�iQ
� !���Ӂ�䓟0>4��a~*�[��m��|J!g�[��@���&���^�����*��0�	oy��S	��6�)�I�|���Rl�@�S:B�T�S횴Q��h���?��ؽ
�r��s�L�裭]��?E��#�2C�f=�W�_�9��59�L�����x$Mj���Z����n0ڧ-��qB�0>�6��p�a���'{m ��?���)u��H�����F��	`tp�rW�7D�s�%ѱU�lI��A�B�D8!��4�;8�>}��G�p��xE�&!)�T"�b�צ���Dy"<��d�'��'0��
� %f�!o��hD�U"���!�@�g���o�R�`&��`�g̓@�>�� ؠ&J�p��7v,%M�!?{\��"�H0�J[�g�y��J�ÉY��8jP�5�V���4�?a�EhP�����,OZ���O�ē7]_,���D��/��h3�K�w�B�It������Z�Լ��>t��˓	�����ڴ�?�/O0��ۆ
�؅�uǈ"Z������QX�w��O��d�ON���ƺ3��?Y�Op��%'ȁT��T��bU3�V�$-��xR�Śf����I�.m6@@�R ����
�'����W!��y�6���0����?�q�'��}H�g����1�`�=C��
	�'',�Z���}��4�УZ�9���K>q'�ir�'���qn�~
�"���	��ޥi�@Q���֫]�~Q����?�#��?�����ԣR9fSj����9l���)E	DE葧�@�O�2�Kv��6{Ge�J�'���w�7S��7�S�ZB�L��@ؙNּ��	Q	a2zM�tG��SaџD�6��O4�l����*�lՓ�W�dX���s'��;��'M��'��H��瞑p�r�p���,;0��Ff�'Q&���`�K�<�@�^D������S|�p!l�؟���f�T�F5zo�\!C���qT���3���)+C2�'����S�ռB�.�O�n���Ɔy�I�JÆ;�`���鐽��d�=R�0F*:H7��SI�H�����d��3�O*�!� ���%>��r@�J5Qf�h��O~��e�'��6-�ʦ]��P�O��IB{Î��0@q��l@L>���0=�G_�Aڸ0�O�_��)S�ɀw�'r�"=�T��N��\�� ֹ-�I;��>��A�����d�%�����O�d�O��NuA t��k�f��� ��w��1��rf����'Z��1I\��Ϙ'�D���^W㐉JT���
tL��)EN�6A F�'��I�Y(��Ϙ'S6�`�-�Kb�[��_�!q��i������jc��'ў0��h�/YHDDV��d�J\�<���&t��A�^�D��ex�Oy�o9�S�P�����4V�����Rz捓�Bˎ	�5��ڟ���������O:��1Eʅ3"�B�◦�_X�pA-�!9-��"3�ȦXf���g9<O"<���L�r}k��IlN�!o-Z$.u���?@�D q  8<O y�e�КN�ހZ�5.������+�'�ўFx̂�r�;��4X���=�y҈W'~�	�h� ���3e��&��A�IB��,y4��'HfRA�ŏ5nW�U�2	_�3t*Ň�y�*���2ΐ�Z͞���I�ȓ}�d���*����� ��d�BنȓdjN���A^'^�L����*?����'��<���k[4��_Byƀ�ȓt�=*�KD�=ޭYZ��\{��	Y�~���	��!��J�^A��b�N�<Y��O;�~�զ�@+~�@�RL�<�Wi^�Dʂ�C��]���� '[`�<��FʦS0��E)�d�z���]�<q�L�z��,�u��44��b�c�<���&@��dʤ%^�BL� �័���5�S�O�T%	��(�& �CeY�Lt�+�"O����%|T��$dR�R<l\	�"O���-N�$��LYe��2K6�t"OF�Ӳ�[�(�e��A���R$"O>-�����LO4�I lK�,��c�"O��J*%A.�L��i����U_�D[�,�O�8���,!$(��\9a�:]�&"O� h����0A��{��L�d$�"O0,�TnuN�m#����$/#�"O��[1�C�F��t&���).y�A"OfV�yL��:¡�v���е*�]x�l+BŨ���+lX�):��26�s�+D�0��,i� ���M�>[��5�%D��S���$:�V�H�CĹj׸�K�#D�����&(e����Ő?p��A� 5D� BVgş���Y�)=2�����(D���kB�w�"�T�̱&n���'�%ړh� 8E�4D��X��@��,�!(j��RU��yr,/y�����`Տ6��p�Ui��y��^�p)�MFA��e;8��h_��y��Y�8_��{�j�c��Q@B �yR�ԃ\ܽI��0^7����iG��y�;wn@�i��HZ�r�����?��Kd�����i�4 P�ꎉ�q��ng�	�bo0D��ɤ$� �8x�̯d��`�0D�L0W�w�Ƭ�0�H�4��S,-D�(�'�98݈��t�Z�U	��3`)D�L{Cώ4Lp-q#D�2!��3<D��+ѣ� 1�<�q Z!U��8�E�<	s(�8�0�+^;bo����#mT�ܑ��4D�$ǆͫ�,����t�~��@�2D���$�P䩛��ʮaI���C>D�q�:H��R��9��4�'F7D��V�I+�p���D>w�<�#�?�O����O�Ԃ4�#��!������H�"O2}jU����)
#A��6`��F"Op� %΄�D$��s�<	�p "O���EV��؈RC0c�$1�"O<2�!�-:����gC��h�z5"Oਙ��V�"V.�
�Q1�H�퉇G���~���ʬGU��`��vw��8�i�{�<���&2�n���K:	����Fy�<�WjA�X�8� c�RjpL�pc�y�<9"��!�������z�D���`�u�<���I�O���h$m��Vg@Ջ1��I�<��d�nT	!E��(
��[V��Пl��*�S�Od��ZSo�������X�f�LYbD"O,����x<�MH��P�
3�"OhZ��HM�t��-���B0��"O��A�O�+QpQ��+O�C�1qf"O�0��*	hI�������A"O&�0�\���P�Ч!�rq�\��0D�<�O
(a���]�p8�-��ra�4�"O@����՛.�z�0�KSX
)�"O-sP�67�,���D�7:D]�"Ob� �.�:B2 �C -_�j �̫"OH��B"c岑�e����0�'�8!�'2D�1��,F��Rg�U a����'鸘"s�Z	�v��f�\4�]:
�'�B�����')
�� r�SC��	�'2h�2 E0�!A���(4�޴��'�FYZ�͎!� ��sٕ0�j��'�DY��E4��|RÙ�/`�������.�Q?�
ġ8� ��qΓ�@@�J��9D���@;b���s�&V"+����7D�<
��܋'\�`za�KC�|��J7D�@)5���DTT�*N�F��g&4D���(L8_,ѫb�N�_6"�hI5D��ʦ���M9��u�N�+�@��O�� c�)�jBQa��$� pS⟆y05B�'E�l'!K֖�Q���
c��D���� ��p`�F�%�N��%�����B0"O���FH��vUD,�`�£R�Z���"O����)t{���U�R�{���3�"OP�Cl�$[�X�X�͌}�C[���*�O���[ �����G$}�y�"OnMJ��Hx���A��V3Iwr�#"On���#)@0�aX�pmd��"O<-Ӵ?�<��ٸ+V.�Pv"O*����%
�ҝ�"Z��}��'�2���'c�=Idg�x��ٙ��$}��j	�'�.|r*� ���@��@�~9��3
�'vd(�FO6�����(!�����']=2V`�&_wx jd�6��z�'_^D�2�1ܖL�f!�eD�
�'L�!"�%6�\��g�QNY����l�Q?ىC��T�ۂ���6�l��� D�,�/�*|Q�k�Kl���� D����.�<��`.� I��()D��"��X?|'z]�(�,��xWi'D����ß�'��,���6~�ƭH#� D�T�!�C6M٘ ����Ё��6m��I��"~� ��k.� Q"M�=��ah��>�y�iM�V���X�KK&P��=�yBi�)�J]�ƃ�DNp z����y�(��/Dų�G�$Ce~}�R��!D���d.E�(�t����&,��DH;D�D{I�=J��h��g�=9�PeCĩ�<�U��`8�з*͜b��z��+O�^,;v=D���0L5W2~�a�A�<�Ȁp�/D�$ ��N�Ri�t�޺����4.D���G��}�$������"%���"�-D�� ӣز�ؖΈ�u��07�*�OZ����O
�2�hݤ6�0q0�֯CFܨs"O��v![�;
`���-�v%��;�"O�ujp�G8��U�2�7X�m"O�y�"������/]�T�"���"O�5@��nגx���_����"O�L�(�)F��YB'k̯A�N0X5�	7A�Σ~J5G̎I~��AB*Z����@UA�<�r�2f��(��B�l(�A���@�<y�Y (��!�,0s��]�#|�<�A�'QI�t�`l��!1Z�g�_�<1�Qb��L�7m�%=��P�p_�<ـ�����0m �N�P�A�������0�S�O�Y�@Hn~R1{F�>VOB�	"Od��.}gX�م$dK(T�	�'<pqU�%3&\ŸԈF���
�'U܋4'�P�����g������'�:]`�O�;-̮��D�I۬)�'*4�Q�j��L���@�Ď
)�t,O�e�'�ЭaFlƟR����'���<�A�'�$Q�AC�f ��v��3[N8���'$���	J.tRD��F��&�`��'�/v��E°�V�L^,�@�[6�ybϕN"İ�)��9�|��p����>a�aFh?�*�XIV��RMQMC��!�Kk�<y2b��[7�����s��t9���h�<a���&:μCc��:��41�AJ�<�#��$��x&�3MH��Ip�<a����1a���O�.zO��@VFAm�<��`�:y&x��a�)J�⬸��i�'X�̣��i^=m�*�8�?������4�!�DϗCZ1�w�^85Kcc]f�!򄄸teN���ߵ&0��VIT$/!�� ����ʝY\d�
GC�#PMA�*O�y7"ژ5��(b��!^�&8#�'E��B6���W�<���!24R��,�aFx��	�Iw4���U��޸)1��\>�B�	�+�b �a5t���A&0=C��<(���A�*U03Mظ{թ�d� C��1@��(į����`$��B�	o¥��b��R��� roG+߄C��!c��K�j�;C���(�j�F�
��	W�$աcd�~3�d��8DC�I?!U`�Uƍ
2��XB&O;#?PB�ɺ[��HSm�M��]��6~�B�I%9l��yr�*��\��b��e�>C�I�W�͐2�+MGE1k�:Ya����C�&����-eK�,�%i�� ��V�Qr!�d;g������6N����@�f!�$6,֜�`���a����@���!����3@%H� ���g�Q��!�$E>ܼ��@�0
��ȣ��<0!�$�"��QjuI�>A ��p-Z"ўtsSo7�'yrм�AM��@:�;E��v�ẍ́ȓz�м����\�h�+�y����T����w�"u�0�R.O !�"��ȓjZ,���+0 #4�D3~�=��+� ���Z9��x��Oi��ą�k\Lpc����i�2Ixta����ɈIT"<E��m�Ԥ#�!=4������6jB!��> 
B��k��z�Yr��>�!�ĔO
� ��g!Θ���D��j}!�D�6P�օx���G�fɐb�8+�!��31d{�+�����j��
���v�h�)�C ��t�D&υi����)}"f�^}�	`}H���	ɒ���q�8;}���L$��B�	Ou���G�v�� hdʆd�C䉾o]@���b-* ��@ư+��C�ɰ �8�����;t�$�1�lC�^��C�	�Yy���"�&�p�W
qP�C�ɺ:<�{ֈǹ=,�)F�n
0⟴8 �>�S�I
	�r CT�]�y2��p�l�*�!�^�i�h�Y����1Q�X��[� �!��I<Z�ƌC���L�r�bN��y�!�D�>���'�L�,���	�!�I�a2�a���/XڤajA�B�!Z!�$1������i�V���Ԉt�L�x��*�g?�ǚ;�m)��O0q	P<�c�i�<��u�<ٳ���)XAP���LWd�<)Į:��BŠʌ>Q�DxD��`�<�F�"_ʮ���F+�ȳ�Z�<yS/U1V.)p����%b0���m�<YVl[s4�kק�3cp�+����p�,�O����u���a���v8��r"O�a ��[��]K6#J�_Z��P�"OV��7A��D��b�*D6B���"O�]@"�\�B	���1P'"O�`Aׯb�`Y���S�e�
51��'��x�I�4I���dh���^Hq� ö�=D��"1ME�7iF<��\]����f>D��{��Y�I?2���ܵ��]�@�/D�<k�@�=T2
b�&2hA`��0D�2Ck�.��!��#V�(aX"k3D��t��B�(�&X�$� A��/�ɟ~�"<����*,�5E��|Y�ˑsulDaU"ODa��-�'E~E�iʋIR  5"O�В�j�
Y�֭cBA�K�@�7"O� �H��ȍ[�QC���2@^���"Ot��V |D� v �4��"O���P�ނ�lA:�I���`�E��O�}�Pi���7k�]�l5*Po����ȓH?vhCѦݶ"B����b�;\sv���T�����.FDtƃD:e��Ȅ��@����4��I��J��ȓs�6�� ��%+�VQ���
���ȓm�ȰcH�*uFxH�W`˴>T�I�Dy���D�=]0���I�ysF�#k	�C�,b�h9XV��g`\�g؉,�C䉀&�	ȗ�F 7�5J�׏(�nC�	�E�D��,�6!؎��E�w�JC�ɧF�P�F��w�mztGS�e�F�?	�KO�[y�f�'�B;�n����F�}񊑂����S`�'�
iۧ�'r��'��0�U�'�1O�I?3 ��!�.I�pi��4iѝ�ԛ��(�$8���g�Ȑ�ר4ú�E|��?7��J� ^px��6L�1g��g�!�$ȯ@N0l�Մ��D%�aۤ @}�}R�<!V�	Hz��w�B}����NCy��'Ҟ|�Oҟ��� �}:61C%��6��w�?��y�>�b���,J �P J\2K�H��+��I2>O��������K��� �ᅿN�)	2k�����~�K�����|ΓPon�)�˅�BA؀���S-{U�5�W����C��S.��<�OLdă��3Nݲ�HȀ�i]�\�D�C���U?���9O�5+���5Fbjm��nZIl���2t����u�Ot��O�P�*5�H�)�8Hҥȼ�Fq���PT��O(��&�S)-C$��7L���e�L�J���I�MA~�'���'�"AL�Lyݴ6�}J�)�&Q����sAQ�x��@�'�P=�M�\p��	�=�Vpy�����DJ���%U&	�AOʘ�O�s��S	!?I&(ʄ[jL��E�ߡ`>^���hې��L�-O��p��O��$֙�H�4�x�ʟ'�˅$�B��#�
^?qr��g~ʟ�d� F���3^���.T6��l�~e�*�k؟���էj����$�+4�$�9��%D�(��$�]�2��@<`��]N~Ӛ���O�ʓ�?1����|���@�`���I�(���2bԽo����'X��~����i�OJ��"�( �@���@ZqFT��lM{������?�'��	�v���+FmG+��E����h��C�*Ja��X`/F�$��-�ĈR�p�C�I?X����#M[���p� -��B�I=g�N�
6-�~�p���lҜe
C��ʤ�r�.��|�h��A���C�	$��,�s��>OH���m	�F`�C�ɩO��� �a��3,l����oqxC��/���ǁ
:w�p �A��1c�C�	�2��+��'I���׺7��C�ɣ����J�$�����@��w-�#<�&�)� �;���ٷ#2-GX�:��	D�<$�r�a�e	/?#�er�G�B�F�����P1KqL<��Gԕ-��� �5b&h�&��ڄE��CC�R�ɰg"W�0�h@���Z�P$4��	qJ��i`	�"�T��EN�f��)q�%X�����b���������i�����ʐ���`�	4�pp{�
��THa���2�H��+��G�| �l��xJ۴~<5�@-S1O���E ܸ{����'�R!ǐk`
���� �T>e�O�PE�' @�戚�g3B�M<��#ΤDɂ�"Y�"|�7O�f`�⬋�ޖ�I�F}|=k�튀��	Dk[�)��'4�9��(R�F�qӘ�D!�Ӹ=����a�/CXP��	W�B����CX�h�G�ޑDkV S�*W2�`�pT
3O�PFyr�	������iK
��8����@Ǯp���OZ���+�.A��B��O� 9�&� Y!�յV�~X
'e8��Ô���S!�=�9k�l3�ʷ��!�d�<[t���LB;���2a]$:�!�dN%�ZE���մZ�BȒ���!�8P�(Z��Џ ��tۣ��x�!�$�3%2�DH�
 '�X�jD�ȱH{!�� ��80�tL�!Q�\�V��u��"O��M�IΩ�_� nV�k"O�r�
����A�Y�U�(��"Of�jk�?d��A��R�T��"Or�zWŕ�Y��X�#_Tr�{!"O�����dVB�B�ߓ*&��4"Oti�%/��$Wb�(��L�6���"O���4ER�)����<STdɦ"O�-z�"�6m��X��FZ�dC"O�Tȅ�͇~�4�k"hK��( �"O�� aLB�u4S!n�*�<��"OR�C!�/{{�SO>�U��"O��a��U�������ҁ�"O���4̕�I.��S�Bԋ_����"O�����!�6�C��$%Y�@�1"O>�C��D����0�;"倈�"O��!p�̻X� �cV�1S�� ��"O&��C�\�4��լ�7U���0�"O�l{�jݚgE�J���6T4"O>�`"e��v֖R�l̺ٖ0��"ONmrǈ	)a��d��[�0y��"O(����31�i:�k>tC� �#"O*��6b�6x�l���jV�t�`u"O��r�I��p-8�󲉘P��Yc"O�e�0�,fP�R��i� i��"Oޝ�/l���d�t�p�@�"O|0�B��q�NL�qB�@���"OpL�v���\�\�*���"/zMaC"OxQڐ�%i��00�!�3>�*l��"O"K&bX�~�uc�Ќ/��c�"OX��0�0[�����J`�r �f"O�8h��߱(�`�d	��83]��"O��ڲ7�Fr �G2�H#f"O��zЕbY���Nۋ�w'*D�+3��p��Q ��H�wH�1�)D��3@�C�I_�h�l�J.����'D��pC��qfT1+G���87��sbm&D�D�䍄mv�#ѯD�rL��pf�"D��z��*N�y�pj��6�x[��!D����AP-F�V$ha�?m��0h >D�dY[�p�jV��&c�j\!��.D���Љ�4#�,�K1��W0|��-D�(�A�J�`	�p��%L��*D� d��)
�t�I�UBH@H�"�4D� �T��l���S��0C�$�N&D���pL��o����#������0D���s��j��c�/ѓ�e3�L*D��v@�9[�p���!�[f�)��&D�,'D�9�,5q�.O�23|��&D��JB��8y�P�p���\�N	��9D���#��	$z Ђ�G�
����Ro6D�����_�Ři��#��CT�4�l!D��Kэ\�a.���E�w���h�)D��4�8Uq�L9��Êm!�M��#<D����CT������B���%&D�8�A��Z�xR��*f,81�g.D�D����#Vb("Շ�
t,��bC/D����	�QMQ�ወ,� �c��?D������X�Zĳ� �:(Ԭ��(D��)$���\���aK��q���j'D�0��A��n}F�@��0���&D�|�C�d: �(���4-�&�Y��"D�|ڡ&^�x�&�؂���0��05	 D�������Ra� 4�]z��?D�� ��R`�nl=�#�7V�N���"O����]�s����d@�Eþ4�`"O�y)$�^��1��N�� U8�"O^	I�`�55,�c���4{���f"O4P�Ō�f�~�3�$�.
u�S�"OXe�bJ���Z����@�;�����"O�	��.+Y����G��eQ�"O� �M�M�P���
�6�j]��"O���7�E�I�5	�%3�N��0"O<�)���	8������K)�xɁ"Ob��⏒0<��B�����E"O<UH�섉lVDm��e�9h�"ࢧ"O�XZ��.8ؽ ���&@:��"Oj�3��K��c�I�TQ;"O�ij�G�9r'�{ C�1Cm&-�t"O�]C�*%S:<1ɰ�V�$S�ɂ�"O��@f��nF��bA�eJD� "OV��ρ?}ڎ��D�߽!A��f"O�Չr"��!ӦH�D.�A��"O�E"�ɘ|y@H�`M7�(���"O.��3G�?C�J��g�ߔ(�L=c�"O,m{�Q;<lty�#K��u"Ox(k֊2u�� ���V��[4"O��"�]*?�n�X�k}�TB�"O:xBd!��8U���TQ���"%"O@�6�ԹH��Kj��U!4W"OL�k"O�g� 퉵*߻`s|��t"O��X��	BD	S�@�5)��eQ5"O�݊'�q&e�qϝ�sT%A�'0��W@��V:P�`֊�%��k�'�p��c!�;` �����
.`P�'a8<*3g�4������?f��ec�'�|�˖�R�U#v�y�%]�b�̐
�'�"P�G߇4.0����=`�n-�
�'f�hB3��v��EScΜ D�!��'��9��Sy�@���#kz��'�(�A��2�@H`��- @���'�(z�"�<B �%�B-ܝ-���p�'����0�\2Y8n%ౄ۸YxD��
�'"F���0Q8ݓ�� ���'��d��d��J�� Æ��ְ��'h&@i�
�/�@i�@�^�����'>)��ױBF�A�ާ%�ظq�'��P4d�ZZ�M RN?#��ty�'	�;ǡ�&}@��f�1 ^~�c�'�;��9N� cf�+�l\��'��uy���Kh<����|$���'H�9��C	J5.��ݬn���:�"Op�;$��[���)C�R����"O@�QNO)1��iA%Ɉ����C�"O8� GYn>D�5��zO��"O��x�� jؐy����2B2�bC"O��d��:;u8�3 �n-�pf"Od�+b�W%X����Bc1W���"O��#	�;������Y��A��"O��0����DYBH �̝3w�X�"O ��G��\42Px�ˮdZ�\Hr"O�S��42BT9��$�e;�@��"O��ꔌ+��U�b0� ��1"ON@xF
��X�p�;G��ja"O����'U�7Lb�&T�<����"O@�8��
�[ ��`k�,V��!�"Ob�5ɟ�{"9 �#�
0���E"OĈ����$f�P�ɀA�� a��"O� ���G�"
~v��!H��"��d"O���F9���G-;��(A"O.<���=>�8M(!ëk$�	�1"O0�W�D�T�"�	�.m����"O|�G쌽,%蠫��]�(s���"O�L���Q{!���@C�e@��"O����W��Qp)��@Q́R"OD��T$��r��E��(]Xq�"O@u
�h�6s�]{�B�2G8�"O��I���+v��}���jU���"O���b��KH�9ڐN�S%�x�T"O���
�S 4���,�&�1r�"O�X�A�ޖsT��2D቞���R"O�p����F� � τ`�p��"O9�&�V܈��	]�g8�2�"OdJ�Үw��8�Ɗ'��"O��#D�~O�}*dݷ\�8�B"Ox����+��52u�ě��]#"OvLfƅi��a@� a�BP"O�$0��<5T�|ðE��3���Q"O�B�(�%;��;��]���2"O`1�`��q+�	�f,����"OF���晉�dhX��66�bH�v"O��٤�0�Z4��$ڿP�XQ�"O�M��*$���V��0M	0yRQ"O��e�!�zM����	���"O>�u(ȹU���၇̾fE�0"O\\�bƙ�t0AAG�c�r��"O ]�1	ѕ@���b�X�p3Rh��"O�}3`����a��REC�"O�bT�6u�\�����B���"Ot�"��VGM���`��$���u"O��`dBY@$�P���9�9��"O����K�~W
�QR,(ע�0"O$�k�MF�I�P��%�ӿb��)�"O,��/@�!YA�f�y��AQB"O��k���^Ͱ(j��![�H�C"O4�1$��Y<-1��3L�܍#�"O>���ƙ�^�أ��Dp���R"O.�H+I�D�m�$\�J�1"O.�i���#K�z���Xm����"O�a(Q̍6���.ZW��C"Ol !���=�BS�T�N:�s�"O^@���?jf�X�%ݪ(�u�7"O�UB!��E��R�e(D��"O�	�@�v@}�#eQ�T�Ă�"O�%����z�ة�7�]9c&$%�P"Ot�VZ1~y�Si݋��zQ"O,�`�I�>�=Hg'�GHE9 "O�4�C�L-D��bئ.���@"OJa�%N��E��� �E�U��d��"O,�Ʉ� �V�,�A�J�3� u�"O 09��CE_�]����!O��c�"Olx˅?	#��o,!�"O��
�
g#�X��bi����"OH��f�5����W�[OY��e"Oި[���3�4��֏UV9�	��"O\��6�M�G�jƎ]�8��a�"O��P���c(:E�l %O ��!�"O��&L���y�e����$��R"OలC�?n���c�*G5? *��"O(���aS	#�6�30H���ebv"O����$���.����0#�\���U����m1�2p�=<OUs� (V�"(���\#�Ѩ�"O� �5�#�<W^��E�Y�0�Z�Z�"Oڅ	f�;.��Ic�����(��"O��FNX�#�6{#,���M�B"O��#P&ߝT�p���c�*}��"O>��i=w�I��L�EHB�!�"O�P�3ǏP��ȟzSDش"OB�U�L�e\~�Y�oȡK<R"Op��J!%Ţ- �՚܎��"O�����nIRE-J����F"OTD I�#	] ���M�2%ĄH�"O���dͶSȆ�;F�H�K�l���"O�p+W�)+�yz��9O��x��"O�8�Z���b�@�iy
�'C���2�2Y¬mJR, �?��2�'��pԫ�;��a���Ǎ �ʝ�'�fd�􄂓s
�%���Y�\��̠
�'9L�C	\Q���I�6Na$-��'��UB���1,a"q�P�.��'5P1C��1InJ�0@�9y�j���'��)�OG*[���%�b�'��s�Q7\�jF�ЖL�:d��'�$��J'�M��~\�y�Ks|����B�a+��gș7�y�C�3P����:0~n,p%:�y�,B1z}Ҕ���J/"��kӠ4�y�0�ێ8�,�Ҥ&VX�\���'KZ�GK\9!��(��i]��,��'F,Y��U�&j�l�w���Y��%p�'VXHy���B�+�$S����'g�0��¶ʮ0BNA��N}��'s�t0�(�ر�tD���Q��'l�Q�p�W;{���g�5{H~`H�'�D�i4	^������w�օ��'�6���5Y��`�f#V#;�0}C�'�Jk��Sg�MY&�;_�`�
�'�d��䌌16&	�`
�8����'i�@Qc�u�QB�'��*�"�i�'�,� Q!j�d��Ktp�H��'"d���S�h��A,ܧh��E��'f �d�XY�H�۰.�("����'�nV �2Wu$Ըe%T�,4z�'��]sV�+��}P�K;:� �',��W�BBF��4gK�U���'�.%�-�#�uH�	���K�'��	ն� �z��	6Nej���'�f���%�
�P���G�^��'I^X&1F�����gпH�r�'��x�p�ʥR��l����-,�0��')(���f�eI���p��".��'�F�Z�WE�2I"�(��n:XŸ�'tY;@��@T������n�8%R�'��x�D�1�.IK,x�"�.�d�<Y�h�3rr�1�d��|�"��H�<�7+��-p��YGcކ+e�zb�M]�<I��jK��u��<4{���0F�\�<i�C�!ZM:Ģ�ޝ7%Fx�!��`�<� ���}��}SX(��ox�<���:ʼ��Q"�l���-�N�<pA�4�\�ze�G�F\"�iLq�<��"^(A��;f�������S�<�%�%� �WO 2��miU��m�<Yu�e�`����A�N)��Ol�<�W�`k�aiĄ�W��©�e�<As��!��U薦�O��B��<� f� c$\0y���Gw�"��"O�b$�Z�&&p�3�?6��\!�"O����׏"�� �U*��4��r�"O�����/wqfQ`�&�4R����"OX��,WT[n��� �"�䭘�"O�!�1��6&�*%*����r���+$"O�V��!iI�I*B�Ӊh �4"Of��a�zX �ۣr�V5�"Ol�#��6�e��M <�$�r�"O�܃�f��}�88,���ah�"O���� �[���[B�N;dE���"O.�R�ơ/(԰�`O�~�z9�"O��b	��&���C������"O^Eh�+S�MX����4�z}��"OE�6�T;_B�6˲��p�"O�hA�mB4GY����c�)���w"Oll8�7{>�SţE�r���"Ol�rǍ�{蒽�$��uш�y�"Oj]���%�N���/M�R�̒�"O��
���Rj��T9_&�bw"O��P.W�Ѡ�ҞFޅjW"O�@���
f�2�˒�B���h3�"O����)��Nb(Y��O��:��'"O�Ռ�>|[����C�5�ݚf"O��Y%��15�����j��%B-k�"O�B�����<:ǪY'g2��r"Opt��ɏ�$t�7��A!���"O������N�9�㰴�"O�����O�~1�b��;�0�u"O�9��أ0,�%�ł�U�Ċ�"O.�"�,ޠ~*
�J��Y;|Q�x(�"O�UkD��>e�+D"�9A��&`G!�#9��%��J`�dD0���!�d�7{� I�+T�`7��I�T� �!�D�_ִ�Y����<̮�I��	}�!�D�@�]�7YO,���u"�!�&R8f�{�@̧- ��;��^��!�[�.��� �4\%��)2z!�dI�f�Jh �,�
8|౒�ٶW��4�R���|� ���|x�R��m��o�[�<�q�_���i햝_2�!H�<����vQn��I>E��oN�;��Sv���0�����y��
`�@��2~�> �A����R td���	 .B6���X�j�,ۅf��ӧ�Y�a}�_2Jɕ)��3��� rB�j EP	:�
O*��!�Y�+�1� )K�,�~�S3��/<��T�K�4�$`�IBv�Si��kP! �/4��Iqcܴ&�C�ɳ�v� &��$ �������F<i�`."��L �B���Z�)��<Q���<  �Q�d�3f�B�J�A�<��.�j�@S��9t�����ɠ�:�@%��.tUZ�A�Z)>9��3�@~�z�c(�V�"�%�$j�|��I
ْLP�n�7 ��\u���SjR�t�*�s�i*���Q|%a��1�lA�CeJJ9�e���'Bh�§�Y.��ѱ��i�(�:$�~"rlP�(�N!>��"t�m�<���9%���礕�j<ܰ���
p�j��U�˟?�ZH���[q��F�T�Ozİ�`�n bB�ٻgЄP@b"O�$��eъl3@)֎Q))"����[�i���2��!m��&�{X�n*�Et�ٚFG�3G�|e���EY��i�퉏l���%Em
�U�ѯ�.bE�5�L#<jn�q�I$%}� �V(Fd��P��.ű2Xx���бz�LX�7�IS���AM��TG�a��K 7G�D��Fd�NZ�b�A����
��v"O$������W���l��f��!��I�K��zA���H�8j��K�>���=ݤ�2�T/W��0����P�>B�I�K������L��}{�'Y�`{t%�pͮ>Y��˛}I�٧�ϨO� �(�h��	h'˒6uZ�Y��'kt�U�A�mX|Yjp��i��
D���u4��ق͇E���Q��Az�*i��)ȑ+4x-:1�8�uE�3���y�'?y �%I E|J5b�<�H��)D��A�@���i�S�]�T�e�Tè���PF��jmB�I<E���O�d��2�M��oK��S��;�y"�Ō!�l,1��[�%ZH�C3�����ɗ˴���nN�p<����g:� ��	(=�d�o]��Љ����|�1���Cr�1� N1�2DG(\ah<�G�Ѩ��uB��D�`��}��r�'F��C��n�t�5D��
0ܳsj!f�C�I3j�䕒��է9(���$��C�Ʌ$�\�ґ�Λ/������_`(B�	�?*�`�%�?�. �F =
B�	
Hj\����/��Z�2ep�B�5$By*�����N|�a
�Z�C��?B`��ͼf{F �5V�dB�I�[Pj���g�B\��� ՜$P�C�I:S�B��́�`@~�!�.�%��C�	�F�X��A_2V��q�*�B�	�2�m���ď|�x�"�=7�B�bz.�۶�9b�!�5!E�CT�B�	)4Ƥu�֦Z?ji8���-nC�	*~Q�9#p�@�/0@Y�iJ�.C�ɼT�������ੀ�b��$C�I��^�b�eB���L��#S�B�$s������&�R�Aˈ�'ˌB�IS��c�zs� V!ˢ4�PC�	2J��k����9nU����O2C�	
fx��"f���2u�r�]-$C�I�_IY��T�9��H��պI��C�I3waX���@A#w�(��P)R�tV�C��@�Ɛ�`+��&�h�t�E.bB�	hJ���BK�"r<�|��j���rB�	�r�Zx�Wc�#�,�R�O�QDB�	MU�zĦ��~2ZyC"�OAvB䉚O��	�%��(]
��4�@�C�	,�P��,'{����o�w��C�	}/>��v�Z�-��\�E�!}+B�IE$�A�)���C�l[�n��B��w��9G�R�]?z}{W�bw&B䉀v:��F�M7vD�'/;;�B�ɏ#��|	�*�=�����B{vC�		e��I��U�J"���� )L� C�I�f���� a�8g8�y��@��T�B䉠q�`kI�C%���D�$�B���TÆ���=�xTT�F!;�B��;|t��Q���=�p��;"��C䉃:����d������?C��C䉿 ���0��O"�3��s%�S	�'�0�s3���O6.��fbE�znٸ	�'����E.9��;wl=l����'�rA����R���C�h�4d��M!�'h±�e��h�1���Oߨ��'���a���g�^���A0H�'�-)���(ۼ�RV�@3)J�Q��'Aj�%mTZ|���p���՘E��'/�U��N�1K�DI!^8�����'��h�0X	Sz�%�톕{����ȓo;���`h�0%Ҿ�9v���Z}�ȓ ��5�TA�jCx�RE���*��ȓ$"�c�:3����g83�2��ȓl�  WD�
(��K�m��1�ȓL2%CR�:K�:�Z�b��o�R��S�? �	j@� 3%�8�����xR�d�W"O$\R�"[���j����-�@"O��! S�O٪x�A$̈́xӐ%3$	�=B�������>RL�5	1<O`XuȐWP^ �G�@��8�qD"O��A�i���m�d� C"O\�p��)���g�R�3���2�"O�A)�<�5�խ���˥"O��J��R�]z������&���;�"O4��wDҩ9�J�в��%(fr	�"O��0)K�
�x��� �{��)xW"Oj@q��C����U�0�L��Q"O���G�
��7%��IP�"O�,�0�)����Ey�X�Zc"O����$�x��,����<{�=��"O���-�X�Ti_,�W"O����*s���U����"OH8����"�$�!.�e0ph�"OFd[��I��$�̃`H
89�"O�|3wI]�l��1�1,[EH���"O`������8��t�ҥL16IR@"On���H�9ON�"e�����"O�S(�}!� �Q�^F�>��v"Oh�5ɉ�E!rl�C���@��e"O��	�i�;��S̘�X�d�B�"O��f��-aP� &���3��5j�"O@�14䅖zp\��r�O�O�>%�S"O4�+3MJ�}K!(R(P���`�"Oй0ҤM �D���Ѓ`�J��"O�YY��I�N ��ˆL���L�9R"OȜ�q��{">�K⪌�����F"O�+5l��y�"�1!��0b"O��ҡB�4�QC�Ƀp���`F"Odk(W�9����F;c���)�"O�IY#C�!s���æ[�V�����"OT�EB�����'w���"O�,3�k��a�D|ɑg��_�$ب�"O:06�M����iAb���""O栉e"^�f��L�L=OFqZ"O"5��lE.�U� L\�a��	�'"O~Q������ 
 �6�P��@"OЈ*��E+%(v�{�o'~�R�R"Otxy�C�%X|H�Fo�M����"O~<Qg�I-i��������|(�"OzeSv���y�h{B�:Xh��p�"O�URB���b|��m�\�ĢA"O���.K"A��t����V���"OzͰ�d�x'�0�GV�GG�I��"O~�eA�Y �x1�+e��"O�%c�N�H��� ���.0�X9B"O,��1MΜ{�QI�@X��E"O��P�旆�X,RW�L�h.�� �"O��Pw�1!ܔ!
��4_�Ĳ�"O@)葢_3�(	(���}|���"O��bs���OC��{BP�h��}HE"O�ӷ�AM:� v��8Y��xXS"O^��Ù�#xzS#�3V����"Oԡjg%J�;�Ɣ�Cn��hNb��#"O�<1� ��[)z�[�#�[=����"O|�j��x�S󢊾9�J�+�"O�(����%�^�� 6>�}0s"O�	b*���n�藢G.��h��"Of�g�rBp�!c��s#"Ovl�u��H�|��r�V�PZ�"Ob�����G*��Rr��1���0`"O� ��	��*8�8:��A��̺�"Oܘar(H��,)��I $��)Bf"OT )`!Q.�50��QOi��a"O4�)'�7>Rֱ{A�܉zxp�"O��  �&@�"LU\���7"O���D)
������nA��Ѣ"O�����Չ9��m�M�)9,|(�u"O���oIk�\%sː�.m�A�"O(���	�|��l���
P��:"OF�"��5��pG�V��t��"On5��9O"�J�!�>@d�"O&��� �H0���14��A�"O���ʜ�`�pE"pM+(+n,�"O��a"mޙ#n<,����(!�"Oly��(��D�$Ҡ���.����S"O.t�pi����A���Ix�8��"O��;�F^ m� ��ӣ{��l�t"O]�q�]�?����A�t����"O[��YT��0���%��>�!�d	�S^ZTb�dA�e)�AcA��3D�!��
�^I[�Kر ��H�L�#Q!� !DY�Y0��?!�>��e�],d!�êJ�d�eOܛ~�8<zAf�N!�^#8�"53��1=i��h�=!򤐁BH�0B��a�\�-�	_:!��26|�%��3R�x �U�
�5"!���BcșҴ�ԵKnQ��)X�M!���|7F��A�t1d��h���!�$sƠ8���L�d��P�ح�!��]����������t&��C�!�^Q[$1P�ϕ�9�`a�E�%�!���
A�]�O�FԂ�1�ùn�!�� IJ8���kY�}�D;0 1n�!�d��Smt�@� \�����.,�!�D����Xɵ�."S�Ar"�,*�!�$ߨXTb=��AJGn�a@C�s�!�D�����T�
���z`n��!�$ʥ3���'�Z�|��8��ѿo�!�dH[�b	p��
Hpr�a��gx!�M�N<� h��o6�\�a
J�p`!�$�8_
<Ț�씺C6
B���ca!�ē�A}�{�Q!ФZ�M���!�D��*p�93�[�b6KҰL�!��)�����U�^�8�t{\!��:P_&�b�8M�ܰaOX�U<!�ޠq|����>O���e0"!�$��ip�P�M������{!��1q~�"��YN,��
v!�$Y�[g(���*f���h��N7U!�L0|>�X!�l-hf� "0�Ȉh�!��50��y *t�� �&HQ!x!��rr$|B#c���	��(Or!�Z��8��#oۨv���ㅁB	m!���+;NuQ��K�Yb��f���M�!��:)�`�s�Ú�\K��s`G%�!�䑃PM$u1��.!�e�o�	t!�DP7\d����f���AD�'qc!�$j?z�㰍�1ٖ�f�<eT!����$�W��1(����
F��]����̒�.��v+���#�?(����"OH�aï�"��r�
�h���"O@89dk.K��\ �8i��	�"O�QW"�O8:D���yI�p��"OؼSE�ME��]��&�V�:M��"O� �8C ����T(rl�%�ؽQ�"ODr 	�r��` LٟA�2qp�"Ob��U�G���2�k�t�n`�"O<YA��?Z�a#$ŋ�t
9�"O5"��X}2]x���[WF0��"O���	w��\!���4��x�"O�D�B��:�FūW+F:Z#\<��"O^d�se��!��$i��/�d"O�TI��Ԏ6o^=��'����W"O&���/IKQ�q#E&�V�>�)�"O��Ac��*!|�L2�"+nDH�S�"O>���Z�Y���d�M]���"O��a��_ :ʴ�%�8W�I(w"O L3��!3����M^��M��"OL�V��m���'D�P�Č��"Ol	*�0R�(�L�'xٌQC�"O��ɚ�;��5�� ��,��[e"ON�zWɆ��rS��7Ny#"O41+�Ј� ���a�0O���""O��� �U�*R̐�@�Ӕ���'�R0��F�tД�⇭
y�,<S�'�@����׺E�������h`k�'N��	�"3��$X�X&z �p	�'�r4I2❆!	�)�WI` QK�'C��2�n?j��M�v�������'Q��r�	��0�B�!L%�`a��'��ti���	~�J$� [�9[�': !i"�ю\ɣ�֒]Ǫ9�'�H�;�P	�&\!C-�`�<1�'d6 #3h�K��-��\?SL� ��'�̨S���|��i�. �Gf���	�'���	��G�I��`S��S�&�	�'^�I��l�9�DL�a�V�4`�'��)�F�a��i�D�;Hi� Z�'���H�"\>K��������'�H����=�ڐq���
A*y��'zd��$��;0����F��@ĲlQ�'�Z�	�g7~�p9AL�2:b$�
�'GҀ����N���� K�7�ҭ9
�'[����&	ʡ�F,B7���
�'6� u��(q�(�ɑK�)�F�	�'��$K�5A�E��f;,��"�'�.]�QÍ[�|��. x�'�<ӡ�E�Q*��aJ�
?r	��'o�h��B�<v"`�F)	S:B ��';DpI�iV�v���R����'��}����:/��	���21d�J
�'�䅉�FJ,�  A�+��AV6E�
�'�	����n)�,Y����Q�q�	�'�НЮ̙9�ʀCRjL��!�	�'�&a��Q�Iښ�B�?̮(��'Sj�J�Խu��4��oٙ4@!�'
�ݳ#ֈN[��z���3���'".%`$�$@�|8RgM�?~2vI��'���3D]�W$�F�ּH�'L6`��$4`�A��,ݡG��8�'f�8��A�V�0�?9�fy�'d�=��ǎ;�Ԍ�VhA).ƈ�0�'�u�!��\q��A6��&2�2\�
�'W��'�ֵl�``��-0���	�' FD�Si��x1
��Z"%��=��'�t��*|�@���9`�X��'�D��P
 ]G�X��,�z��'�=ae�Sqz�hao�<|�N4C���  �hRaچ_Hڴ�4a�S��-�$"O�P(�H��*�4h�Z�D�ك"O� Ɯ�tT�l P�~]J�Q�"O�L�ӌ�9�HP`���9\L��1"O��x��ۆ�z9�&,�f��-��"Od��3�*��U�#l�T���d"Of]��$$6�T����q�S�"O��y��ωT� ���F�@�"O^�`��7�%k��9M��mqb"Od]���3 ��
 �Q��r"O�!����'>���K��S<�����"O�p�ǅ_�8���R�ބ^sR(8C*O"��0`f��R%���H�T��'Z�
�I
�}/�h1ր�,s�]*�'�(QJag�FV�$�D�??�Ȋ�'��I��T�t���4k'���i�'v:���.�ҭCR��Q�T�K�'.�M��ѭ	�5Z�#1xs�T�'9���l��w������B&-�(��'H��#�iÆ�r!A�U�����'$X��B����Z�S�iHK.4-��'C�)�I�@wBU��I��~h��'�|qXW�0�=�V@�3�@�
�'�>��5�	_M.)Z�f�'xĮ H�'�̜K�N��pBf���ޒh�T��'�ڡ��J3�ڦd�,{&A��'��Tb�W[ѼTi� T�p����'�rMpT��!c��qbU���e�.�R�'g(�y�d
�h"h����J$� 3�'P�yG���t�08T�S�@d �k�'��`�K��X눜c���;�h��'�@};��Od(J�`�ߢǔ��'=�l��n�2����Ń�4���(�'qn4 �N�enXlKL�0N�œ
�':8���(5D����X.(�Ub
�'����1��(YZn����(hA�
�'�x$xwo�;X9�)����&�4 [�'/�t��M�/2+P�����/cT�Q�'N*��7 ٯ�`a!aٴu��EZ�'�~ਕ�ڵM�>M
A	�g�P�9�'G��ڃ$�-L����w!�eB�1�'��p�	B� A���H
H�A��'D�DVS�8\�S�
�98"L�	�'���b�^�/:D�O];7��	�'1N��L��Pb��Î>.�.�
�'h��V���1�f�)�љ�'���åM̈ft��E1!1����'�x#2��+UO�9a�HND|�X�'��I��"͒�R�i��?;w�4�
�'�0|23�m��SDf�7�$y
�'4�X�$�R>TDʱX�)��e�'�=J�(�$c:�YZ�"�%j�\r�'R8H#6HU0<�x�vً-i`���'7����)d�>�@�[��J���'�&�{wg�l���*� �>I��'���ґC��C ��ʥ ߷$�U��'O�Jt�W�#��e����E�T���'��M��$�$F�1�㔱<cJP�	�'�n�k�`Z>I3�ʕ-Y��
�'�|)Aw�ژ}�H%�e\�,�e��'	��������~�R�N<;ڸC�'�t�!H�R7�ɁC��7#��8�'��kc&ʇ�\zs %9��)�'��Q��%Z�� I`H�\.��	��� )�Un��o<��)7g����("OzM�E�Y�jF��!�|��J!"O�����H�&��Y0���?�~M9'"O����;+�@��QW����X�'��qA��JY�����O$v��	�'��!%ѥZ ��[G`	P�k	�'����(Ɩ���1M[�7���'l��kw�F�uv�ԭ�*��A��'��֋�	G{j�z�*۷9?�-�'���3Ѐ�� s�ޜ{vZؠ�'2��¢!G���狒n��}H�':�`�ЇQ���Sg'�/kcl]B
�'Ty
'�A+�r@צA�:���
�'�䠢 ��rɋ6��I}�	�	�'��I��L?B�Ԁ��ŗI��<	�'�xHV�Y0� ���ڐr�'��5���A*�;0�=0枼r�'�b�3шA2�^)�A�*��8B�'�
��toH�h4 �w�'H��'¬�v�ƴLx$৏M�$:ؐ�'Vft��fɳI&�+"�(P�N�+
�']<𠃂[����ËI����'�P�ӧ){��a��l��F�v���'�.Tɐ \}˚⭉-߆���'� �[b�CZ�q�$��'1h�@�'ۢ-)�i����{x�y�b;D�<�A��hل)U̬��|�s*&D���#Ȕ�GѮ�d�N��h��L%D��Q���*,&�c�Č Ai&��D�!D��q�E�`^L��<e[1Ç�!D�����CVXH��8a������ D��K�\����H
U�����>D���Qiګl�2Z��D X��E0D��a�1�d9�_��
�3� D��Qj�<O^�آm�8�6-� �=D����m�5,��E ��.0�.���
!D��a��L�&vzub%S+h�"��D!D��r!��;c��iۥ���Z��@8t"3D�,��,_�xa�xR�V�=<�,�&H/D�X����;~`ؕhn�Rj�H,D�$@���4���@gm_�!(����-D�(�],N�"ɦ��:�B�bcn-D�`����?��@�rKI&���� D���\$L�1���Y <��2�E9D�T��N� `i�$�r�RZ��i�8D�$�'
[?FH��"`���f����:D�ܹ�؀l���R��W�yx�qg6�㈟R���B
Z<0�ڢ�;#[*��"O\�xЈ�1g8>D�Pd�0!zՉ`"OT�"C���V���Q#R�;r4�G"O$`�R���H���G���5�"O.q� �p�f����?y8 Q�"O6�(B+C�6��]��g��kr~�h�"O` �@R�d&piŽ�ÚYQ"O�1J�䍎"F�rlK�\��8�"O��V�̏B�p���	��=ʡ"O��ª�<{�%Yu���⚨��"O~�
���,�𬈂Ղ1܊!��"Of4�B�zr<Y$�{��y� "O4t!�g\E8����7P����"O�dH��	�Y	�<Ц�ϼ7�$��7"O��I��
y"�|�f�Y�P���"O���R���>HR H�`�<=��8Cs"O���C˾�(�P�������"O� ���_�!��Z�.�Y��"O���uj�c0��� �)p�XS"O8HCp�
V��W@�1~â<	"O��觢����������"O�H��o�.��űvM�*� 	*"O��9D�?�Ѩ�쐐3�H���"O�{�� �� ٲ�N�J,�)5"OH42R�P���8uȟ�FH�3�"O<�)�0E�8�ZR�פ'||�	�'����D�ԑjNF9*2�X	-��TH�'\r��"*J���b*�p�Y�'��i�t�X.fg�HJ"!O<w�.�{�'��ReB�W�BT �=Q<��'4�L���ql�x���x�N� 
�'���N�
GqtM8���qzr2�'Ϯ���,Y���4��h6��J�'��8p��i�v���&\0\4,��'��p��(|�: ���'$��'<,�����K,��%�(M�:͙�'�ށ�Vb��s�(�!T?�p�9�'��y�[�A�t8��=U���'m��`l��9Ǌ$B��D��-s�'��q�k"�P�a��B5����'�����ȓ��ء0a��7���2�'d���:h���#Bh��'e�A��'b>]����> [x�� �U�!�x1��'7��A��E:MȮ��A�1F���'["�ʴD݊?�9Pfb""��j�'a��@R/��(�"W'�XXq�'���I�)	�8
��@
G���"�'JP�s�$��	�i�@� �*c
�'@$��f�]�}8��Y���4�hY�	�'夕����"Ѐj3%Q�L��'�`�r��>k��S�c�1k���'52�(��ǿ����i�����'�n�7�O$::XK�ҨI�~h�'��-[������	4*!�'������M�ܐI���#Y�	��'6^Y �A�98��ű�R�Bˏ�y�O`�̍�����^���.�F�<�$�I2<%L "�鈏x	��Q�.��<�����4,�K�
E�k<��+gÕy�<I���'�B9h�Xp��5_���ȓE�,�rP��}m��Q���9�h)��^Xm�rGNX}��e��5���$D��#$���Ǐ+o=@��C��a%!���`�5�×���Kdq!�$I�'p�Lq1E	�t��u��/GV!�d8_a�ѭ�6�2,c�� x0!�RЕ���#H�ظ�mX�V!�ć�$�J���-��-�^�	M]	f�!��)��5�h��1�:|ٴ@804!���/2���r`
�;𪉃'��6M!��4Y�慰�'��H�qr(ǥ\!������z���7�X� i�0'!�d̞�^��G��:w�^��HY�5!�DԔpx�����+N�@C��Y=w�!��W&m�lYR��C:Bw )��FS�y�!�dE*�tQ���.��9#g虴u!���;��Q�V�U� ̑���:/�!򄈻%H�r���z˪�	��<F!��W7#)�e�`�D:dR��Eis!� b�a�	�uI��Kg�˭ �!�d��!_F�kv��+�؉
t儮�!�� n��g&,v�k5�Q1"O$�3���:"5��z҃O�T l�J�"O�C�տ[%@��dE]2F�P"O@\�R>%�8e:wA0T(1�"O��C���W\����ȕHpc"O�c � 	�g�Y1�P3�"O�V�}`a��G>� �)!򄄛1��8����y�ʄٷ�׋d!�(]�s5��w���j��S&S!�ֹ7���+"�͡��I��[)!���i/�л��ˍX}��r�=/o��䋭�2���4���s�􈤷%me��!�f��i
  'KKH6i�U�����U��@�v$�WA1�S�?�NM���ђ�.\f�E��[�#�����>R���I�(zw���r� B)1"�o��GR>ט'nq��
Aj��p���e
Q'75W�KqӲnϟX�O���M�Ц�%\?��p2d�������
y?�����>�4ɐ�\RA	S�gWдw��r�'8�7���E%�dkG��Ԫɔa��Ȋ&��4nta�$@��	�0�h��4ݰ<��J�to�	�����_��q�(�:�v��t� ;������,���On6�Ex�c�5�d����]�7�����BfAP(��r���Pm(N��誟^]r�(�^����i��$��Ä�|�d��!�>V��dC��T�?�glF!�?���i������OP�drӾ��1"؃<�$�Qi�(KƬys"O�k�͍,�~ �A�Y z&pj�X0�M��iL�'��d�O��g��%+�9:�̨ ��Y���ՅVLfΑ���ȟ�
�ZzFLq��M2T�V�##�j� � �#�gy��֪[�Szٵ�	2-(��ʒ웮VDf�1��$p �\x%��Jт�������
4Ɓ�nc|Ƞ��&+(&�$������O
7�Je�h��%Zv����"��iK�D`�4�?�)O�$�OޒO�Ӯ,��Ѹ�D���`����CզB䉚��"�AF8]�c�ar�ɟ�M+U�i������4�?9����iH�_�|��?x�>}���b~��	dJ��������<B��@��� B� N�~��>PD@�C�B���!�*/�r�(�� U��<9���R�����"��0�U�g�.�b7.��<���D7~`���#�n���n�"��#�nm��П`��4�?9���9��E�"�b�AǍF/:x�lc�I��Mk��@*��<E�N�{�|-��a[�z��H�2�O�o��M�40���7i�Pd<�Qf��>q��h�ޠ���if�W���?�%�����ŀ<2�,�'���N�BS�������E�(Gg��1���0��!�J(�S�?���AU��=�B,�kбe̛��R�"�&� 2!\�Tܚ7m]�Qɸp�a Z�:V�#�˹|�1�.�h�DγN�6��˝+C��oZ%M���Ʀ�`�4�?�Οv����oԳ3?���v���ԙ&lĕ���O���dF�i��n�/a�R�paݟMjQ� bݴ8?���|��O<��hY��	b)q�hzC敡r6�h�	Пĩ����^=��ȟd�I؟X:[w���i�d�ItLF=5N�#�N��b]�	a�/L�q��p[�V���(*�!��f�iF�`�!3s�|"��B4�S���o��Myp�U�o�: ���1�i��� �p�a��j���f��\�H�@�����c,_-����� .%r�P���?�"�?�?1U��3[L�gyR�OD��9��\�`�֮fn�1�J8Bp��G{J~j���la��	�!-A�'��6'6\⦍�I��M3�>�e����䧏56�
�] |  �    C  '  W  �  �!  *(  �)   Ĵ���	����Zv)�ll\�0R�P��
O�z�V ]�n�1���2�����ӊ�y��D_�~!�$���dJ��c@�1q^���)�!E�n�u �,4|�Sf�����ש�:�h䈋3�$��E�f�h���ҙAiص�c�F^6��5��s+�-xW _�6��a�$��R�2Qv�ُm1���	�RvFL@��A=AԄ8[�L�/�� KY�W�P��Nǭ(��h��3;���{��'�r�'�Rk�~�F+<p<�n�����a$�R�
��ɫ#ך("'��H��Dkd�	���!�(�~�)vB�(&'��h��
�<�b쎝iʧk"��C F�F�XX��d�����A"d��bMo���0�����LJߴT��<����~�]�-|ȑ�'!>%�Ip�HZ��y�A��A�*�@��:�:�CVS��M���ɤA�*���]y�m�ʆ�i�dE=�%XlH(/��d":D��1�ߥP@�+ՊX �$��bh'D���U�X����
�A�P��Q�P-#D��J�Gӟ[r�Ѡa��0@R��M D�pR�X�a��q��nS�|�*Ds�9D��Kdj��n�Z`�ʑ�ct�P;��4D��[6)Y =�
h� �k��{"%D�C�(�/-� D
D왂W�F�C� D�����<R�֌�A!�;o��8�%-D���A�T9�l��Ƅ1(-Ƅq�,D��P���v� ����bT�b�'D��C��� =\����1z��(!�#D�����;^y�eC����|3n���� D�DxS`�E?HI�v��w�hP��L3D�l���Q�H�rP��߹ DD[`G,D��
6��*���b�K_�Kv����4D���U��kcX!�Ƥ"����4%=D���nI�.�faڄ6�^ɹ®8D���fר`Qv���B�K!�Tٓ�$D�|��&��\�nՊ"�/\0��%�%D��{�儯	�v��u�Ǔ!o>���K"D�H2�dѲU����e邥%!�@�!D�t�W�Y=j� ���:h�%b�,-D��p��U����j��Z�H�JQ! !D����E�U��!��O1H�0����.D���ۼE�\���Ŵ<���$�,D�PaV!ԭ_��� �k2p�h�6)D��J��/Q'j�q�	]�Z��Cg6D�Xh�dZ�"-�9r��&t��X���4D�t��Kčl��p٥�[8���"4D�|�d��W^Z5�v͔�/�Δp��<D����kǱ	
�`��1cg��cn>D�����2@]�)i�a��^��`�?D��;�'�+c�.���hS�<�`��ԏ<D�|`w/�)%6�aQG��g"���G=D��Ò���L����v�Ś+ D���S-�+�Vp�}r��YW��yr�� 1��j���x�Lj�K[��yr�W<@$i���r��䪧��yRjV����wm��V��牅
�y�J ,2�
�KʏQR��`�&@��yRCz�X2k��S�(@���y��TNh����b=:�#�y��7.�n\H����J2��
�yb���� �T���`)7��8�y�M v��`��8o�Y���(�y�Wod�trGP3	&�`�Ĉ��y ��"�������=0��!�D �y�G�4����Qj�� �TK�9�yB"��U@�R2	��?�v���2�yBI�4��h�!5�<�K�J���y�L8_��2��N��{!���y҉�4	���r)�	^T�Ê�y/fk�Y*G%�WaP�h����y
� v���G69.��	/�N��"O�8;�/Ƙ
*���ġл� ѩ�"O�G�D��zhڶa^2`Xq�"O6j�Ӣ��U0��ү B��"O������ZE���J97W��'"O���$a��Zi�Q��mO��S"OL��ʇ$H������:Rd�� 6"O^a�W�׃eF�Ԣc狨b�|�&"O:�xr �1p*�"��C
OJ��2"O@�9I;Jά(!�>�L�"O,Y¢	^6h��5��K��4�:di"O���E�]�b4��)�Z���B"Ox���9;֊���`�難"O�)�V*����p��pQ\�i "O���F� �,&�Ii�$�"<j� "O�"V)P1r���%B��kxE"O��p��k�%���r�lM��"Oɚ�ˆ-JŐ��� u�R�!"O��`��(
LP�+�]�}��0CQ"OX$S Bgle��囷p�v��"OdX��H�r�U���27Z���"Oht
faR�[�̌>'�A"O:��r�(=n&�x�`QmF$Ч"O��;��W�/�^�9�J�:Q�h�"O:�Jæ S�J�
��H����3�"OJPcv�L�tSs�-�� �"O��w�Ӥ6Yθ'd�al�]c"O\�J'��0764���f)�d"OH r�m��|�a��jı4��l��"O�@�p�BȤt
��Qf$ �6"O.�BS�0�z�B�-dIB,�"O(Y�f;M�$�����5�Nt�"Ozt�R�ыe�B9P�^1-��4c�"O�i��h��c��^�`c$"On�Rpj��a�x���اo�iIq"O<�� `�-��0�u�U;m�I"�"O��Xp͚U.|��@��/�\p�"Oz�t��O��h�b]�	��"O�u8wi�.>)�����w��"O���#�= ��J�瓊
� Lk�*Oޭ�Te|V=��o�6��� 	�'�DͲ�B�o�*�֫���m��'��)H�7>XC�F�y����'��Tl�!r��I���;k�0�'Z��T*\��@30,�,��X�'�D�;V(��r#�rR�_R�c�'��y�ү�;�<�5�TPgށ �'μa����R��
�gW�9&��:
�'�0a�ȃY�D/��l���j��m5 �X	�'y�i�̎#+�m{��O!���\flI�jU�먁�5.E���aΆ$n!�'���E�,O�`�5b����l4c����'O��b�U�~� i8�I�$���*�g	9`�\�������$J\���C]�;?2���!��I��yBM�{�2��)��	�ɶ*~-
�)_�9*h��A�8�!�đ$a�����fG��l��RNU�S��4����ӭ��8'
8� D�H�������|��(g왂$�&X)""O�.��5��y����4Y���/�iR�Yg�ǟL�@�.1yq��'�,�3/B?:4V܀q`��5%��
�'M,�1��ėL �m�U�OMC~�ʓj+oL}� ��&���0�WJ��,S���}��9��Ϫ ��z��%O��y"�ؙ.�V�h�4�����!8V� d��Dlh&�y0�
1�!�������g.?���XE�D�1�剙���jR!����Pw5�E�T�ãK���t�Ўx�`� 6�ԧ�y
� Nq#a��I.�Yڑ�^"��{v�R��!��*��]�.�!�ʟ'��O91O��"t�F�3q ���*j�f�k��'k�� p�������,P��0��]!Xvʼ�4� Q(� qB� �azBG�=1`"  ��7��4��ɿ��Oā��"\@-X�D�'fn�S`G\��V�t��(6� '�^P�<C䉦r�x1���O��pA��,�ʓ�H����#�l������n����V�"����J�7R�eqJĶtp!�$ETK�q�A�R5������RC�L
7\�,T���ڸzl@0�Օ����1�z9�U�ekb�z3��}A!��[}��;�-���3vDB2f�RK��^�iY�i�#�$�ד[J�r��V��A�
�Q��ɰ�~�J'E�X��B�F�Rb�$3Ӣ� >DQ@��#9�Z�"O�9�u�Y�:�0a�A�x���� /�vEq�ん�H��]� ���ffĐpM�iux�+�"O��G'����
���Lk���㆑�>�-�4�N~��=�g}rG�	�UJ􋇹tl� �[��y)�kf�E[��8z{ �/�3�M#q�ܘ(k�p C�'�BŅU�3���1Ə�{<L���w����t��)]��C�!�e9#�5-��)qN˻k�!�$ςCS���]�8�*I����}VqO���R��k�#� C>���2�I y0�M�W��l�<q2W3qP ;��͖\y�g�p4�?����O��1�˸GET}��M4mЊu�"O��`�6��}1� n�4X�w"O� �B"��t!8�[�nF�4[t5pB"Oؽ
�)ǘ�*M[�MPx�\Yw"O.����ʋU�V4��G��ddX��"ObH�MFO��!S#gʁ}��0S"OPeIc�	� v0Y#�`�>=}Ȍ"OB��2���H��4m�c����P"O8�3�P�z�Dj��^�ZPs�"O�H뇡8��k���HҜ\��"O���DfM�-A�Q;d-�^�JA�"O$3w�H2;��;Sf��^���ۅ"O�V��; �d��ʗa7*;�"O�Ak���Q����� $"��0"O6X@B'G��M�P
ɼT!�]P"O~e�h�i��]��J?P���"Or�B����
ږUJD��:)|h�"O*��,�2t&a�q�ψpB��W"O��c��P2/u���J�XxК"O���k¤&$tT8 CZ�3P:��7"O�%xc/Y�0X�;���kG^�I�"O�,a+P�H��Wa��a�r �s"O��C� ���80�Z�i�4,y�"O�Rt@�Acr�QԉH�F\sg"O����� <n��Ba	52��-��"O�$��m���
K�v�`��0"O��z�BWᐩ��o�	�Z�"O�)�F�0'�bX�w.�f����C"Ov\P�˛�<s<q�爵b�d9Q�"O��b�l�$��d��9o7���"Ot�딣[=!+F*B.�9y*� �"Ob��B��%$��j�,TuZ��"O�����x��)Ж�M�5Oe)w"O���[#M%b�)2���"�DH��"OT�a�ȏ.rJX�&D��p�J�ò"OH�ib�]!H������X !"O���AVR�$*�հ�	�b"O����˄G��a#��{�r�T"OB1��>���7��0}R"O��!���gŎ|i�A^#X�J!W"O�D�aKR�8"�T���8Z�6���'L��҅нD�z<"��I5��Q��� �bdd��S�șQvb!i!�Q��"O^�2��QjAI��n��C��р"O@���Y�H�qt��K�f�v"O�D�!��խ�iײY�v"O�QZV*B�_�ГSC�3?���0"O�H�2h�R���ǣ��-�)�"OXX�m�)FJ$$r!�]����"O,0u �=��G�*"&��1"O<Q�ɗ<��Bƅ\_&��"O��:C�"j�����B�����"Oh`��F�"3�Lbb�$Ԏ�p"O�yТ	>;�
t1Tj�@��p�""O&�c��C��h��@���V��!�$�8X�h�G/y����b<�a��T�00��㕔tmر°L�p/d,@�'4D�P�4K�s%Ic+�:4�|�62D��l��$x���*��+fV0��lJh�<��-�:���
7f��xq1M {�<�v�X��X��>w��ز&�v�<���4�8)9�,/'���׍^I�<��
��0�$)N�t{&&n�<7b��6e["���i?�hq�N�m�<)1��,�&��9���E�D�<i *�#2\-�WfE��u1eCQF�<� ��E��L�aIS�:�ar��|�<aT�W�f'����O*Yl��+�B^�<	�� ���ٱH˥6
4L�W�@F�<�唄>��H	�%ΣJ�����NC�<���֊y��)�G�� r�!4�X~�<�f�q�a#\@-90	NT�<S�\Y,h� ����N2�h�2��Q�<�'�ֺgK�d��+0&4�LyS��g�<�G�/t�8X9��K�
�D�f�<�%bG�8��͏ k�� �
Z�<��kAvQ�'-�t R1�	VK�<�W
P���K�B��[�K�<�wgԀzGt�S�MZ8ܰ#fb_D�<� @�I���)޿s�����E�<Y���XT��Ш�q��"ƙ!�D$M���z�A�:��UJwaX�F�!�$N.��0�Pށ��K2�!�Dǡ Chu� %� ;!l*���z!�DOl�!Pd�߷�|0"�B��!�$òS|i"b��  �N(�k��5,4��z���2�\ ��e�V,���1D�Pi��L�d[�;��QR<00e�<D���7gƏͪЫ��ϗW&��W%D��)�ݥpm&\9g�L4 6@��#D��UI�qXx�S�.���*t��($D��ȗ��/yTX�I��:\"�	!D���Q������g@�#XN��db D���1]�E�z�aLA�� 选;D���@ ��	�ԁ�`�1 ��7D�,sv�ЛX��iqd��c�ޜC5k4D��1�
�7d�)���Q�Q[%S)=D�(����%Q��Hf��*i��f�5D�� �Ζ�3��A5N�r���pb6D�<*7C?@�!��LhX�� 'D��C�HE��"�JO��XQ+0D�H##��5�8G���%������,D�(pwN]�s���0�H �;t�+D�| !\:�"6�>p�ܽ�7G%D���6R#��8GC�wĊ�aR"9D� ��(��TX���+V�e[p�8D�� P<2FDIc���m
�X�ƈ �"O�@���;�NP��+�)h��"O$�pW�@�!"��wiS=d
H:r"O$���� _Ƃ ��#]E��6"O�4�pg��(��C���):�.�yb�^�t�E]6�%�f��y�L��9�D۠B�9=�TXрM�;�y�
�1[���`"��>1���@�yBn�y[��P狇�}l����ձ�y�
2Q��DHB��J�~�2���y�j+?b��P@	¥6D<Q*����y�)�<�����e��+��Ys�_��y��J�R!�Q	0��*=��Z��y�e�%g*Qb���+�4|�@�y��ڵ=-J��ӫ�B��>EȊ���'��1kr-ҹXW�UH�l�96��`�'�N���~�Xjs��3'�Ԁ�
�'�����B �B���G�V���a
�'u��&�
za �K�.7��e	�'�ڱ�g쁡�"�r���aB��
�'�%��h� p���n
�W��'l�,;��9��bu Z�Y�"hP�'_�y�!�UL��{DiɊ=�F�{�'�M;4�c,T��C�ʋ!��#�',��'P2P��G�޹Q^��'����C��n(�[�x%��2�'->x��K�!����ܝ8���'l������;��ܱ`$e\�H��'������<?�"��@e /1Ld@�'�8 fR�r�j�2@�P��|A�'��X��Ԕ��a�Ʉ�)�T*�' r-h�]x������S��`��'Y�4×	�U}訸�%�.?���	�'�MWNʎ<�f�(�`V>P%��'K�dC��ΜX3�B /�%�'(ҤPgl9Fe>9Ї"ְj��'�^eZħ�ah��ڗ6��3�'�J<)���%r��V�C�<ܢ
�'�4uk���l���/�	:��A
�'�y1vNR
;��	�98�Hi9�'^�i��n�X`�G�0V�|1�'�B��"�Y���xhp���@�a"�'����K�+L��DQ*g�0��'�C4��7 Bе��kZi3ji�'᬴�FB,b;^�h�+��`2�'n0���k�T�&��	/D�"�'�������Rn�����+�0�3
�'����� ^<534���@X+	��,��'R m�7���C����m�R�ڴK	�'��C�+�(���C"Dk����'X��k��� BZXqp4�C�T���'|F��
�m�h���<��	�'k�����!^��Ȉ�d��:B�I'=?Ҝi���(M�$(�%�?t 2B��T��4FV f��e��N�K��D{��9OT)
�m��IU�<�f���=� �9"O�P���D�=��ؠ�Lu�����"OT��`b��CJn0��ˈ<���"OT@y�V+}�C�e��I$�"Oa{AH؝^���Vʆ�I:R� �"O�q"����f���wH��4�p�bD"OHcS+�2G,U����0^w<e0"Of�[H�� �z(z3[12k �R7"O��I���R�8Ȓ�`-�Jx�A"O� *k�ѳd�n���v�f�*�"O���c�ETk�耆�ݘK2�e1�"O�Q2�I�#?ҙ���T)S'�Mc�"O��P��[�zP�=��KN�P<��"O����Àm�ր�fAJ7`S>�Y�"O虱�g��Suv0�%q�6ء"Oj���x�^��D��d���a�"O�(8� c9 �k��A*�'"O�0��KM�y�n9kT�+��k�"Oa��οg�� �p�A� <��"O�-x�j�9-	E�ue��)(�P"O���W}z0z"�TV�� k�"O���@g�(T�DHa��Q�2��aPw"O�9�gCX;)����QŪU�"O��r� �n�p��R��'�"�ۄ"O\�H%�c�&%��j��<��4�Q"O,ɣ��R�X,H1V��8�2��"OT��1�^���9&��$=�0��D"OL5SbΖ���`Ò�P�?�Z��""Ov8�������(�`��W�X��b"O,����M�и���ϱ{�>�{"O��q�*Y��|���תu�~]��"On���%D��\Ҧ rgPX�"O�I2m��K$0�B�Оrhrɉ1"O�yS��ށh�I�.�=[f%"O�=��'K-\��R�صA'�T� "O�h���/*��@P���J.�K�"O�S�RA7�`��+h��g"O"��"�P.w��eQ���3Z�8`"O�����'t�Yb2M9Z�ݱ1"Ox̩��!K��M(U
_!h�����"O��c�h�`��IB5	�t�F��"OPd�`)ʒO��Թ5H5�f���"OZ�%O;:ي�#�J% �4��""O��+�̜�l����heP�"OPT�&�?!��1�ή����"O�8��.��;F�� ����"O�M�!9�L����,�u"O���reF�HR� ��σa���%"O�l;�����
iE��yS֌�"Obͫ��؋/��,���Z�rPp���"Ol�XSA�a-�!��"a7��b�"O}�Vh�>y��w��"����"O�y�0 ݓh�FM�Ék����"O�`C�5@�J
��߁!��["O��S	�
+���Z������b"O�A�5�H�$��=�tC�6�Ƒs�"O�-KbBۧS�` ��k�<(�p"O���>O�T�"F�H��5��"O���fƅ!/\�E"���G�`�!�"OL�S6��&<���� S�]pv"O�8�vKھr܄��@
.�|ٰ"Ol�����$B���\�ܼ�	�"O���O�=��A�@R,%�pt"O��xAW춴��O��48H��"O��*���9~h́�M)&��Q @"O$yCg
C�1�Jy�LKt���"O�tj�e�%@6ܡ@��(o���g"Oz��$瓶_6!p��2bX|�"O�����J	o�a�C��<�H� "O�QKg�'BlD����`/��0"Oؽ�$��q�t��3���9���@�"OFd��#G$jJ����+q��§"O������I9W*\�ff8 "O� ڐ:*��|ɲ��`��C�"O�Q�+W)i���O��Q~%�"O�H
e��/{�ћ�-^/�h�*�"O�pQb�'J=x���(�	"O��A���"5��seN���D�6"O����*O$
ܹ9��΋\��(��"Op���@�9|5���B�UN�0f"O`�cr�O>Q�j�B5�Yt0T%H�"O�|˰&�R���2%���'�Y"OR�Z:J��pE�F�G��Х"O�T�aە������V�H����r"O�M��W'<�)g�<� �sp"O�eP�ʅ�E���Q7�J�Ibf"Oz��ˍ>�J�i�������y�"Of�q�W��hQIDK�"x
q�p"O.�;�A8e�lz���#fH*�"O��g� 
NSp,��CפUဳ"Oz1$�۽X)�u��C��lX���"O��ȓ�  �P   k
  .  �  E!  H(  �0  7  X=  �C  �I  wQ  X  W^  �d  �j  %q  iw  �}  E�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�
�;�>O�1"�'"d�D�B��3�91���b���IWov���W��;���nd�%R���?ڑ���?M�A��iκ�)���XP ����bu��;uɐ�_�V8�Fl)#�(�:w�[��u��S�����'�t(�!�J��d���Ae���i�EW%
��TfB�O�٪a�$i���Y��զ2�J����ß0����r���=ͬ0����ِ���۟p�I��}�4���O�@р���d�O8��jEQ������1�´0��O���O��d�O��SV��OH@C!�'�����4���%��u��)�$���5�O\�	_]�g�̿d�m�2�G	K���y��|b�ON�ٴ�����)�9|Y�4�����%
�������'-��'[��'p��'�������Q��tC���*UX�1��ڟ0�ݴ6���w��X�'-h7� .�@�nZk ���� �z��X�vrre(dcÏ2�F�h����r�9Џ�	¸
s4�����%N�l�{p,�{�ȩ���]H8�x�d�;��7M���c�4���3V�ؓ���%H��9'�DPj@�JO"R�(|җ�i�������� �I��ۇO�hss�E�.p�(�$p�hyo�>�M[���

f�"�)� N��M��
�����*D�&f��io|6����ёC�Ԛ}��jSn�5qE��k�oe�8���0v4�i �ʃ%}��!O�C �ac�C���6����)��4@��q�[�$(�DD�J6mU:V��Ð-��*2
	�ϴ~��H�⊇$"C����:72�děQ��3��G�	l"�`�� 9���>�Iԟ\���B��Xj�4��Iǒ�H��ڳ	  �p�F$�Q�d��͟�'9P��8Ⱦ\�#����Mc`�_������1�.Qx�����0<	$����`�E�&���� G�����4,��t�Gn�܆�	9&��$�O,�'^2T 穇" bX�X�mڡf891��?�������ON�IRx0�# O�,!��z=�"�j�p0�"�**��d���&<�xH��Ҧ�?R�T���'��T�V�>��7#�(+F��(ccD=�!�ªb9�BB)M#o�@�sa8�!�DO�5T:d�W�B�ȹ"�m�R*!�  �b��󃍬pl���˿D(!���z�H�JG�5(^De���צa�!�䄈*��o�^W��`k�:�R���O?����@-����>38��afOp�<1�nG>ck̔{�C��l��= o\C�<��kJ�N",���Y�A���� �~�<�1��9o�$$a��]�B���9Vōc�<ib�"`�2��*�
������v�<A�CҖU�P�*�\����9���kybEץ�p>�"D
;v�t�
ĥg�y�O�h�<9cB��\���3&�:RbR	95�e�<R�S77q;��E�i��I3�
Za�<���3Q��e.�Lq�e1�@E�<��ޕY�Vmj�j>���P�%Tfx��RCI�M����?3�Y(u�4aХ�
a>0��E��?��.�Dl���?���u���a�M��Ɗ�h��T�S��y��.*U�塣ǚ�|�axR+�dN�)*#	B�	�B���� 0Ku,��ąدQ4󲮈� <8��/�~�	�Cش�?�i#]��zC�=���� e؞���O�⟢|:G��3@�W�\��\��ǟ�Y�b�X�'�>���4	�z1*��10AR1 ���u��ч�i��'�`Q8C���9&�O���%V
�Bc�Ͱh씣P3�C�Iu[41��a�'|�|��h��C�	�Z�+��V#9<������C�@}��o� �%�Ǧ�?�0C�I�(�MZ�:�Z,���ǵ&�C��8-N�;&���T8QuǕ�^��oZH�U\��͟p��ҟ\�''X�.�?�:u�D�G3&LHw$	6�66�����P�ݑ=v6��O�:�8�i�7}��P�-��O:^�xf
��J��3�U�5�B|;d�G��b>�kwH�w����<uJ�ų&4���c+Ⱥdpj6-�y"-\��?�����?���4t��a���V��A�z�a
ϓx��O��B`d3D��U����'3r��4R�DI�4CJ��|�Oh��T���I͘n0 �:v�A7԰�A	Q�66Bl�������������u��'��8�|T�B�B�wP5yC�#�:a[CGƀ��x��Y����N?<OT�uA]�	��"s,��f���qP@M�U��]%��#e.'<OY��n�8rRt�����p��@��U��'WB�D(�'B&҄��̄�^��Q3�dȿ2�t���
3���R;�v])tnE2> Y'����4�?	,ON�W+�ަ}�O8f]�k�x/�hk噦nƌ������O��d�Oz�{�R�#���9����W�H�)� X �3���<�u�T�2��@�'�����K�Hب1UOK��y��j��D�c��6+j��1u#!�0<	'&
ǟ�[۴�?��hH�:�dRQڦ�N��B��U���?����?9����'��'�)�%�;�$�F`�<�p��O_��B`|y{��H�k�&��c�(�?q-O6�˶*��q��ß�O�.� ��'6Vٳw�ל�r�
ąT<����g�'R�_�v8��T>�'��Y�����Y�k��X��@�Ox���)§dT�5�a�36�lY��˳U+�4�'k�����ɧ����#x{�pԒÊ y�*@�"O܌1��Լo�����IÜ�����	�h�2E�v'�Lj��D	N=�`�s���D�O��d8���c��O����OF��x�yz�eTI,�8@c���� �'����@�A��0�nAc>A��T�&/� =�~�����vHЙ�d�Gv��P3CoZ�������	@�t�U�	W�p��\`�'�q��*��L��T M�R����in^�k��	�?����'t�2@dMC��BQpH|��'�>|@6��uWڽH�kA�<�+O*�Fz�OH]��v�A�W���)뇆|z�}@$��/v���p�ܟ��Iڟ��	"�u��'(�0�V�A����e+b��TF�"yfH��i�g�!�D@�SO*�0+�	1c6���o^�5i���O$�0p��3BbD������͘��ڪw���'�O� �K�+M�n��l�3)i��A�"O^1;PA��SD���9Md�Qe�|2�e�ʒO`�7k�K�T�'"h���˔\��a�f�K�}qh�3��'8�H�o���'	�i�e�R4�GlG�Y�=zuf�O�%��\�"���S�I�/&l^L8r�'���Ȗ���{L<H�䏋L��B���f��4A�:u0���)�0<���`��Q~�2�R@`�At��H�F�����?���:�Cg!D�(	�!�,���I��?9k�7��{V풵Π��BE�l�'�����`�>������l*B�$�4xmj1
ڮ�6������O����˕�]�0) r�M�:]d�kq!����_>q�Ϟ?v�L8Ѷb����`�KGW~���^o2��㡙u:���'���a%'W?J�}qQ�Oh%BH�_��Mr3�H��
8��O�����'�7Mܦ���l�Ol�p� �@)k����읳l[�`�K>Y��?������O��?7�1�(�-%���6	G���dD2�c�.m`��9=D�2�N<x4��3��eh8��4�?����?�qb�?L�����?���?1�;H;�)aׯ[2��P4��,�Ȣ�Ð�D�b�r���q������E�RO+���L)�D'�<m�Q�S�� 4�Hq��Z(vtT-Җꐖ3x�BE�<���z;(��a��8��:e ҹTOYDP*��Ϧ���4�?�cV��?я�,O��$ԛ$�JQ+�[�p	9�J�<>����O4ʓ�?���L�z��N��d�3�"�ҽ ���<�$�i7�=��|�,O6p�ֈ�B��)չ�N��g�����&�O>�D�O����׺����?��OG���Dc��J;2����S����K�gϗ`2�A��%�c�數���*������'�)�$LΦ~媰*��Ԓ��� �3`��T�4��:X䐭�C��{{��Պ�n�'�>욥F�/�6X��/�� �����L�?9��it�#=9��D�4Y#R�#�*�+v�,�3��,}�!�����e�e-
$hҞ�9��'-`7-�O�=Z�4+[?��ɤ����+��3_HE)�אvސ��	��h �ПL�I�|�5��1��F��@��}2�L��i�TY:�	�(���g��	$@!��h�8W�|�<�I��#e�l)��ȁ?H i�����ۣ�_���D�'��>0n��"M�&	E �<�`�$��43�I-���6膀m�R4�"��69Ŕ�Ot��$zy8��'YP`�Ц������O�I��/[-hw�Ѹ���ԥP��'��O�Uhg�ϼ�DU����iG%7�>Q[F�@�<�Wh�*qZ�)`��Y�-2l�D~�<aD��E}�@s���n�"$^�<�WK�&�]kת� &�\��b�V�<)cD��O*��� gN�MG���R��H�<1�[������n묬��ȎП�K1�S�O�|ش�]�O��Ex7n�^=\=�@"O0]2�)�(^$F��`��:�`:G"O@�S늉�����+I�h���"O�\z�*N�;ZĂ������[�"O����n�RM�g	��{�x�!q"O6����}�ƭ�u.^���1�[���@�)�O�8�n��VC�8PP��	��R"O� �0��3+/D§ϔ�s�:�"A"O��큼92�Q�nL@�M��"O�-ѳ�C�L���+� q�"O�)hL�:��ܙ�c�/�Nu��'����'¼i��T��p�Y�m-��
�'��tȭ?"�m�`�G�R��S�'NB�Q�A�$?n��Wm��kB5��'Q����@�W��h`��7�`�'榽�cŎ�)#ؘ�v��1� ��'80�)�I��ce����
L�!��@���±s�Q?(&�֕R�<��&V�2t*!�'D�б�@�# q|h��NT�;Q"����%D�,����c� yP��V�3�7D�0"���d@nx��$M-%�F�A�3D��6,���a�wFL�H�V��@B6D�Ĩ��đ-��qw��D������O��"�)�'2��;�Ȏ�l��ab�B�T���'s�<�� ��0�����>O*��'�\aXե�8k�ʁ�"��!�h��'��#��I�b��lX!-��|��'��ՃW�jB�[#AW)&.�I��'�0M�͞>EԮM��d=!���-O�@��'ea�
J@,)s��K&HT�pB�'�� zc�ǭ](�A(B@\�KJi��'7��2�L&bL1�a�pH�,��'[�$�@�\4M�\ٓ1���n��Q2�'Qg@EO�Ā A�B�7�0�H���%b(X�l?)���F�Ę�~	�ȓ���#獂�(B�(0�*�>W�p�ȓc�Eأ���;b0ś7�7��`�ȓ3x,<�B,	d�f"0�+_*х�]m��ْ�)�����mZ��ȓ9<@`3���W�b5s���E�
�E{��Ѱ﨟��Q��}���*ԬE�k�T��"O��p�f_�`������׏M�%�"O�3F���t������
�
Pw"O����h���M ��Y`t�)pV"O�#g�SA��:⦍�rc����"OV�sb�#eD%�RdP,;:�
��'������Ӊ F�T�L�`�� d)��thć�=�@E(�̖	<��-�)�J��ȓ)�Da
���b!Z$	rF�NW���.R�`�P����ɠ�C^3XU��M����tk�o@����N�tFɇ�EQ�����
�'�Z�����4�X$�'7`���%���*1�ױf�<8�����@�!�D�����d�>-��Q���&�!�$۫w���A��#�p)���+?�!�;�N�� &�c>�C���)�!�D�ZjZ$P�fW{ �q*Я�*��}"@� �~¦�M:ب*2��x��AP�Ŝ��y�&�'�pM��xӤ$���@�y�刵!�d�@�F��^��8�a�K��y�eJ�G�b���W<�i	a�ϓ�yR�@5�����Q��	�����y�ꞁ"��8�&A��奚��hOtEA��өS���q�U�|Ţ�c�cJ�C�;���b�@8������)�C�I6�jH�U��)3iT�� ۶q�dC�ɇS1&ap�
�euN�1��]�,C�	�	��0RC䟨 64��M'
C�	/}n��k��
Hb| t�J�0���)��"~B��]-r�xH��e��(���!��0�y�d�.���
�s]T�3a�A+�y
� ���chOUh�C���!I *e�"O2U+�!��'�P$���$m�(�"Oư�v%L%�z-�%�A4�}�Q"O��r���l/��SW�@_�uP�Y�@�D�"�O�<�Ab��I�$��J
�lT�	R�"Oș�
�Cv%��ߺ1��XU"O*�+�C\'�()%i�'%�;D"O����Z!jx�5.E���J`�:�y��eX��0枝2ޔ=B 
��>����g?AW+*n{� o�utpAY��x�<����J1섑|��%9��u�<i"bg�t�v]��s���y�<��	PG����cF�MH�}su�<ygD'�> uM�NV���S[l�<�!B�<�z�"�+v�k�Cd�'n�u+��Ɏ�-�	��Cبi�� �˜i!��	E��e�C����iк[!�ε3>��a�M_�M̌<*�GٻP!��~��0��ӃG��#VNM!��MN�1�G�/s�����f�8q>!�d#�>��uat,��B�Z:23��4�O?]�O҄30~��͖4���c �K�<��I�q4�8���7@٪�AK�<����lh�s�,J����d�I�<��U�D5�!��4*"���/CG�<�(*/|�KT�Xdm8Ј�F�<�d^�1Ө�b�.Ԅ;30��dh\FyRdJ�p>�%D�����ҍ��H�n�!��L�<q@"P�3ݎAzSɅ=!O d)�l�r�<�6�V�����S:P��M	�m	p�<a��̤���
�DT�f	K?I6�C�I/cBzI�k l��13�ج:~���DE���>�Zx:aE҄[;626�!R!� ��@��)d$���J��`�!�B>L�M��:��8�(�_G!��ٚR_������!L�(YQ���L�!�Dނ��I��w=�������!�d��?�YYD��0Q%��$��<p�ў0a0�'� �!#�B:E���1P��ȓR*��Pz�W� /|����o&�L���)t���;b���Z<��!rkҒn�k�	���Ѕ�e���YRG�N���׏��ߢ8��^����OLTV&����Ӆ'ǀ��ɶt:#<E�D��&X��,"7�Ã8��Ia`#N�\�!��'#"���$�'6=��9"�ܣd�!���pK��{��9���q����-�!�D1KTX d�~@���k!��6���{&�ϱg���o��r�!��ۏv� ̈b@R�P`���Ȇo��I�6^���C#o�*��1JF$M��a�'R?hQ!��V�(�ƀCˀ�a8������bP!��F�2�
"��;bm؄��n!�$ц���1 #���A�FVb!��O��T#���7�� �E\:^�}2����~¥O�C��wI�8n�
l:�J��y��HCȥ�'`ǯ_�d�������y�G֋<���QL��^l|�ȧ ���yZrvq)5bx��\�f�$E@A�ȓ3LI��f
G0���D�"t�P���\ޑ�0��/�D2�Mܴd�)F{R��>����II���Ha�"h*�F���"O�Y��-�EbXD�@�M2
��,�d"OP���.}��	�嚌m;��"O� <��sl�G%��Zq#�x�����"O�Qh�Nq��=�s'G�{h��"O��0�u��yPp���m^ Q��'Lp,����Ӭ�b(�p`ӥh.uyWLޖ	�M�ȓ=��pC&��4�r)��d��I�E���	U�V�<���6����d�R<&�������D�ȓ?0�i��ж-���4F�_���xN�!�Ԡ� U�ԡ��B�<x�葖'��P��S2�@�!����m���B76~����)��u�AD�3(@R����p�j̆ȓYI��W R@z�z��	*@�TT���R��O(N�y���;n�2�3wh1D�P2�
C�j����1qU"���b0�O�\cU�O�r+aՉ�FF�F^ddA3"�A�<��#ɵ8�P5�J�/d��D1��D�<	��L,!���aA�(_{�p�ERj�<�V����#'h��s��Ճ#��d�<4c��Q��Q�r��2u
(��.Jk�<� �3&ẕ��!�M+
,"�(�^�'��=���� �+h(3!64��\2GQ��!�dE#QV�@v��Gj�]&�9�!�
N���
���we���F�X'U�!�DM�_�5)N]�RWڈ�T%ޔ�!�C�Ft.!+T̉?'���B�ў+!򤉞~�����m������1e��F'�O?��(��:W&i�h�YK]U�<�Q�� �6)��ݘ.�1�z�<i��F k�� [wHٔoT�`�Ǆ�t�<��CV/F�fi��aM��U��`q�<y"���2�@�N'!km3�ph<a��۬\�Rx�1�H�B!��&�A��?)J�,�)O`�l��M��1�?q��#��<bv%5a��XL�S���
�2=������?9��X�F�k E �
�q���J�^;vO�;!Z�:���n���	t"�g&�Q��D�q�'Z�rdnΓY�긠���NC� ׂũI��QX����m13aܪb!��el�^�'� �Q�1��#"�I,�0�k$��[��)��@��Ix���G�Qd��b�k,y%�)�5#�O|ԕ'T���u��= W�^���"d  3�Oz��O2��ƒ	qw��Ӄ톷O��u"O��!���mpӋ�P�^E86"O�ib�_	m��J�ʁ�6��LX!"O�|�oŠK`��&��r��U��"O�H�u�Z��$�,1q<41'"O�,b%%�z:�@���4rjB4��K��O��}��W|,Ā�
Ř��)�1�_j�V �ȓڐ s��L��Hi�V�^=V��ȓ"Ȓ�#�
�Jp(�4��"a�ń�P[�iA��+-��̳EL	 hؼ]��'~��e��#�$PYY���}�<�G�`}0Af&�,<��yeɓ���!�<�OT�pfיA�r�JO9�P�P"O:�`C�Q�f��x��b%�|p4"O|@pv@�\��q��m/���3"O�t�AD�6fX�������"O ��pBÏFvB(rF���l��\���'벴2I�0����mB��V�K�%D��:B�S7/�|�c� �+H$�
 �/D���A$Z^C��2��N���� ,D���5�Ɏ��1J�j���;�l+D�0r����"�D������-D���B[�Y:�)g��X��p1�ɦ}��"<���-�%��B��q����D��@"O^(	R舓Ӝ=!��_ ,%��"OTf@��m�i��/q�	�b"O� J��AE�d`��N�vY^) �"OhmX��K5S>pP`��T]��U�U"Ot}��	�T*
�����-�6B���O��}��e_0Qz�f�5�x0C�[��Y�ȓ6�ʑHq��xS�a���Ԕ9
\C����D'62xA$�n�D��&j/D�L���"%��H���3W �*D�`;�
�:lj�I���@��u(4D'D���t��;)t��0��''ʎpi !�OAh��'&�D��H�3�Kgbי"iv	�	�'��h�A&��i$���������i�	�'�z�.% ����](!��afCN�<!rg�%�,<8��Ϣ!ET9Q	K�<����z��(�ڔ��t��h�F�'�@H����>�������-����%��
|]�"���?��O�?A��?��d���`1F��N1�)�R��0|�U�ƅ,NA�Y��U/nh||�d��1�pGyR��z.:��ѾT��36��
`^�B'�M�l0a�#�1M�ɣ ��/�F�Ey����?��ib���2�;1%؆'MZa�kKҐ��d �O@�Cm)8�ZU3��E�@�
b�'�˓1:��؂(�I@r�ǀ,��u�'mB�'��t�'��|���Ib�M�T;��yG���-9ʢ?	��S�>��ݫ�m���4q���&��⟈C��*����?1ϟ���@�d@Q��F�w�Lr����'� H�O���<�%���V�ìT�{vx��P��eT��0�O谤O\�Z%�>�����j��N��:p�� �>� ���Z��5�O�9���h��D"wZ\���ηvEZ�Tp^d%)��>�$�>y!X���w���_�P8����G�&�J����?��E|�$��v��?�P�L/j�y�4ń���0�����&}��1}�)Ҕ���0�M+������;ՆP�3�Y�q��sy������#�ȟ�$�D�
c|�����+���)7�i?����p�T>�	�u�^�"� D��<P��
Q���:�A���f(6���O.18���δ1� ��D˪'�.Y�� ��2��x?A����?�M~��t�3y��	�+"���RL�= `)�Iw�aRbZ� ��)v���&���;�y��Y(���
��Py<Qj��צ�M{���?�+O<���Of���ƺ�S��4P׈�$U24���iRP����&����O�˧�?�ڣf�h���w���1��?�؍%�L�	_��|�K�����(d7f���ϰM�$Ӈ!)D�����H�Z�����M��/��l�t�<i#������k�g�Y�i�\�<�*�=�����N=E�<��s�J`�<aP� ����q��G'��1��X�<�b����J�v�*��!�^`�<��W�D���w,ܯ&z�!��_�<)��)+B*��2�^F���0��q�<���G[� �M^�R��a��i�<i��+�d	�"D�<0��M�R!�e�',�"=�O�M7�@�^~.	�EF0v���'��� a�H�"�*}`AO�*t�x8��}r-�J��+��;&Ő@��������[ae��<.r@c�l���#�
����4@v�?Lؠaf,^:,�8,[�.ARS!�X�
ubΩ#�:ԁ��%$$X@�A7PO��Y᪚>�� s͘R�8$�5�M���	 ���n!��-ͯD+,|�c���T���	�M���9�U�!�U���	AS�Y��	��ݟ�A7O "Ķ�N>�O��	X��P�"R�E��5����O��r�!z�	݁�����>$�F�'�!�GÃDeTt8��Q�^�D�(�a�o�	#:�h���̦���4�?��aS�_�F��dV�\�jH�`@O��':B�'ՖriՋw`�d(��T�Y�]9�*�Q��Cr��"�D�P�O]>�.��e�K�(�9)���>q��W%�0� �6]�q;5f�V�<IҭW$	ε3*KX�!�,�y�<�U�K�q  ��Z�N&Q�cn�J�<�AAQ�;�p�׫�*��qB��AE�<1��J+7z�� �%4��ꠦ�U�<9�$����:Ê �W�� 95��U�<��LI,N���FּC���P`@_P�<� L��)V� p���" ��C"OV�`�J�9�a�6�>,txy�A"O�$�Gh�:/��`��G�FTX�v"O�-!tdD3�p$�4!��LF�{�"O��J��$���n���3"O>=�����D=��J�̌�I�tEkB"O���s)�qA{A�0 �*"Ov!�(�4}Li`P�ʒ_�d�["O�I9��6R?��i�-lI���b"O��4�?���3�JlB%��"O4���="$���!ՏU&i�@"O����F�5�|lb�`�h�Nd �"O���GH��� 3$��(�n��"O�l��7�#���n���"O^�"��ْ�Ҹ)�K��.�|���"O@�������Jِ+�jju"O�X�k8u�����C�8['��#!"ON�`RAV� $<!�^>4�8X�"O~<taƯq@) ᑒ%�E��"O�Y�b�K�_(� 2U�*i+�"O�D���^{Ү��R�D`2"O"Ai�G%t����
D>�!�P"O�͊tdO�xQ���S#� �"O�}@�V���r�f�7U�1"Oź�%c�"�1�c��	��T"OF�Z�DJ�j���:D�.`6i��"ODUb�սC�h�H�#��N:�A�0"O�,0���p�n5��ȹ
}��"O��%Eۣ��t��"͊mHE1"O�A�g־p<ȅ�Gk�b��g"OΩ	 d['/,�(�E�R���-��"OH ʲ�Ol���R��<���Pq"O\eC�
6Bς�3����2�򘈐"O�!aC�d$�!�@�>m�|"�"O�܊��Qh���m�T�l��"OT!��@3_P<PP�T�X:���E"OR�x�@�Z���m~&p�9D�����o��!��ֵ+���Xs&7D�Ȳ2�7k϶��'V�0����qb7D��y��ٳ?��KGaY�w+ �sJ7D� �E�*((m
��Y��AI@�6D��b��T�A�@�p1'�h;���, D����q����A���u���!D�0���A1�4��ӑ2����J>D����+ƥiR!�Q(�~M�%>D�H� "�?:C"!����d8�#n0D�(ȡ�(9��"p�&4�f��C,D���m�����1M��5>�0�F.D���`IE�2�Z<r���J[<(#�*D���ȟ�&ǂ���`{��B�=D��[`�%hd�0E+�*$�3��>D����c^<������Y3g�ִ*�.D�,`d��u��u����:eE\�*�!D�p�`M�V�|�*�œ��Y�En;D��A�)��dl0�L�
���r�5D�(Z��O�T���%�
�gǸ�.&D��y��X�fq[��ʸnĠ�:��%D�����O�
蒼��Ɓ"%�\s�&T��¦GW 88�� ��ޛf�HU "O@����X0b8LU�D��Q�ιH'"O��QS�B�e�*�K�D��o��%bP"O�`�g�:eܨ��;0[����"O�x��bO��c�/U��`""Ora+�^/d�NL��h�2fQL���"O� \XVJZ�J�~�;�B�")6�q�"O6X;�..0��\6�c"OD�@`�	�[�����a�1m�l��"Ox��c�(*Bdq�n����V"O<1a��>15��b�޳��1��"O�PS���X٨�̓�[� ��p�<��)�X��o[����]n�<1qH٪o�F ��l�u?
a�CF�n�<A9R��"��Ŋ$`�\�Pɇb�<�1��	�.����Ӑ.�F�1��]�<1���I=(�X2A�V �D� �Z�<��N�AVbe�eJL�8�`h�C��R�<)��/f���DI^p���gPV�<���X�l�" G�'+�P��Lz�<IEa8+ZI/%�haT�*xhB�,��0e��;cH�{�,B�	"�=�͚���12�C��+�R(e�.}�~%`�h�b�~C�	!�:eQω���x35�޽q�^C䉿!H�0xt�7��4����&.��C�ɣ7:��*օ�-o��#Q��VPC�I|B�3EB^B�S���VC�	�t@�p���E�� �.��hB�B�	)\AxȲK� @�̛ĥ�B��/���*���D� (�ž��B�ɔV�@P�fY�h�^` ��^8$JjB�I:yT$8A.\��o����/�d5��Q����� ހz�H<�ȓQR�J�j�G�l�D	�J�ȓJS���
� V����[�[Җ��ȓ�����PB�p+\�#�&��ȓ[SH)���V�N�ٻ��C�0�6D�ȓ �|ekբ�%g`b��E �:[o�y�ȓ6��ؠ.�4���"�
ceф�7�fX�'N1ւh��ˀ�*�N �ȓT��Xqw�<R���̗�?��L��h�Ȱ�t�5%�
X��	�xh-���I`e��(0�! �D�	��]�ȓhQ��A"G�<,��MY��Hu�ȓviڈ�wS�GΚ��G�D6(贅�eQ|��c��*"�4I�Y0u������	+9Z(��W�y�4�ȓ(�,@b���)�-��!�.̈́ȓd���Ф��'N|���-�|�T��ȓ�(����.ot�;2�7���ȓ	����"�F�ӢVM���m��x"���|�e��"!���|N�i@aD -�!��n���'Y��I�F�o�~�HRB�p���c�']�
@��_'f�sk�cj�"�'��x���m��L�r&��d<�\��'���QB�M��|(�J*�P�	�'��Tf�;p��`��� M��'��� )N�A�����mK��L��'��!����`-�4X�lʖi����'�0�k��� ��(�$�	�'����)�4x�d��lG�O0��'B����1<P��I}t����'�4z�̍`W%��C��G�`�2�'�4�H%�9��=�b�H@,v$Y�'�x�7�N	6yF��KF�?�. y�'L�8Eo� 8��}�F4�Ty��'�v�ђFO`�L��h�+/�QQ�'�D�BG�1�l�'�	*tFD��� ����
�O��AY����FN�)��"O��֥Q�)��\�,�S�p��"O$=pg�	��i�e�2ǂ�i7�#D��#Ŝ����i�$� ͊�� D���1kM�,E�Lhf��-?<*�x4(!D���ぁ�A������C�%�U�,D�07�C��`�ri�H�B-��+D��;��mb,Ds��}�)p�%D�$+"@��8��ڶ./���h��C�	=W`г�h�R�	���͝� C�	Q�X�S�MD�����6J�#%��B�I�Zb���-_��d#�#Wa{rB�:p�`��v�;��@X@K�-�XB�|�y��@�=Нr� '�B�	�LE��Y��'R�§M�jҰC��kǆ�1���%/7��I&)ܻz�lC�ɮv��{�C�|�`u1`��&�tC�I ڠ��(�bG8���X%$BC�I�r9�IؕO�-b�
 AX4_`C�I���hɁN�0�L���l��
��C�ɬ-;0@��fO�F��X���B.��B�I�h-�l����({��� ��7,٨B䉣'��cs(�Z�:D{��]!H���EN����τ�y41��3!�$�'Xp=�7*X�V�G, 9!�$�2g��b@�|u�6T+!��4KѼ�G���6t�	���K)�!��W#r���< U6����!�dG�	>�}�BԻJ:��A��$(!��ä �¥��̲{&bp��} !��@�B��܊u�Vo�.W�.��X�ȓY�č	PH�2�胑	+��-�ȓڔH�D�p�����ʬ6�N���I��d+���;�� +H��ȓ.R���B�LO�#��GWFb5�ȓ4���G�ޑ+��c�ٰTk|0�ȓn�`����<Q�t�kuF�[A���ȓ1F�hՇJ�Gz�S�m�:݄ȓ@�93��
_e�)�,�#g)t�ȓD�rI�G��Jl�}Ђ݈@B����4��q�-�<5���ɍ!t��ȓ)�PT�G�B�[�6�ȆBëeK�m�ȓ&/FUrc��CWXMH��Ok��ȓy[�� ��<Nh��#ΎP@=�ȓwX:����és�H�s�C\q ���Y젙PR�\�	A$���p��,�ȓ}y\���H\$-��`�=q⩄ȓ��1�nŶv.8�� PJ�͇ȓ�N�|	3���G_F%�ȓ#L�Ak�nо)�N��q��7rf���ȓg��i�7�/\�(��3�*�E��aԩ�� %b���Bۋz�\�ȓ4��ɣ�g�I^�yҀ��C�����X��0j^$ 8ڌ�B��D����PJ�L�9>���
�~�ȅ�n��� ��,}��b�Ԁ)S�}��`�9�F^n�a9���!���ȓ3�x`y���
�� �	�=Qz��ȓ�L�!�_�U�h��C/� ��ȓnwP8��	ۮ�ro^L0 )�ȓ3��x�U�˪I�=#��	�,?l$�ȓ�r9s`:fղ�:��"�h��/����F��*����eJ#]�� -� (�(� �<1&4�
ϓ|/��p�'B�T���A�:B.Ň�S�? ����	+�miR�)h](\x�"O\�bA�"�h@��:Z��"OH��&Ǐz�(�q�A�Dv���"Oz�x��:����)2[4��$"Ov�*�k͌�C2�KO��K7"OXHp�T�	l4IHP��z�� ��"Oe0����c�^mj�(W'���4"O0�s�ё g\��#�8d�<��"O"�j��ߍm:���B̊�`6e��"OՊĀ^�9
|�x5��0X�U�s"On�4��-p#��rC�nSVm@"O��1���53�q�D��x�`!"O�9ڐ�ܤv �@"�ۆd�Y
"O6���%W�T�#a꘷Kd(�R"OnM�F	
�.Ŷ|Q��qo�D"O���׋D�f�H������
8"O�=P`G�,j&��9D��|��"OZ���)Qe��i�N��bĴ�A"O ��R��H��Y GF�wR���"O
4+���<wb}��C�"$ M�"O�Ҵf�1���Ã(I�F�i�"OT��A\� 
�@�"�+�P��"O�pC����|����`�&�	q"Od`�kA�W�!7M"P�5�"OV�s6���:�S�C�U��0k�"Oh��҆��n]�ӤH*WI�#"OH��ՇJ xd��DM�J�h�y�<�+�T֕�v�B��1RcE�t�<�"ʋ+@Vm� ��r3�N�<	��RU��!hq'B��|�D��<��N�)~4c��U:W=��yeυ|�<���XӐY��G�1%���`�Ct�<	�fF��}`,Ԭa�j���ls�<����4�$��7׳r��1A��CM�<1�����<YcTs]V���MT�<��"���feL40�<�aƯE�<�ȓ�r���Pp��WC����D�<�#.�:H��+�!O/B�$�b�C�<��	�ISaQt��k4f��u^�<yT"a3�	c"��3���`�j�b�<)��Sz���fߟ/�lfLXb�<a�"��0>��`��ѐ����iE�<�G�H"G�F	��΁1��a�EM�[�<q��^�IV� ƍ	��jQ��lFB�<A������ҕ��720!C���y�<Q���6�r�S�&3��� ��}�<q2ᎋ�P����1u�{W�Lq�<qs
"7��:�j<�Y8dK�x�<1�̚9ZXC��;�F��w��m�<�&�y���AJ u�`@F��g�<Id >P�8���G���k[g�<9�g���H�'�6y���	#��x�<�%�J����S��0{���I�<yͶ,Z�=�K
�X0��B�<ɱF�X���[���|�b�+�KRD�<�1*�(i��K�d�:#ܮd��j�^�<1'�4�$�q���n��jfl�W�<�v�U��00%�����S�<�1MB�]oR�8v	��� ���Q�<��T�A�%"aC�x��Xu��P�<ie�Yڎ���E��� �w�<�!F�_8|�[�c�T��a�	J�<�!���h����f
:�h9����F�<9��W�6�`����=i���A�<� x��.�'3V��R�	?ef�y�"OT��eˑ����2�:D"�"ON��2�E�@j$����y���*O�uj�	�	a6F܃�ϲ$F� 3�'V�pj�!T�i��s�ا^FR�r�'���[�\�ԅ�R"��$����'��883�\�P�]`Rɛ���b�' j���i>Wޞ�{�a�'?ےm��'�2t�P�KbW�����P�ma"PY�'� =Ig�"����CH�`.��
�'�>4��)݂rd���
+3f�#
�'G,Q荄U���p�YB�A��'������Z!ې��5Dy���'��h�V�y	�\����i>I(�'�(U����M"h�8��K�&؋�'{^�!��*Gz0���Nq�ԆȓH�8����03>��@�ηo��t��J��B�.؆2;��I�0g�q��;0��RF#Җk�XfJ��쥄ȓ1��k3�^�9}����O��  �ȓ���RL���(!�C�BZ�)�ʓ2��3�+�©ȃCP"�B�I���P��� �:�N2ū�(�B�	�@�i�1�2�(]k1��c��B�I7��P��D��,Qデ�C'�B�,2Xٰ^>62H;t�:��B��R�L��0+S0I�hH���5.�~C�I5|�,��E4�u�� �$�ȓE���g�	Z�>e�`�N(d:Bx��`h�Y��,L4Z�w,��=23dMk�<"BY� �V��J�@��cIh�<�A��2�H�ݨ�&�6M�`�<9�h��C�xXg��hO�u��`�<!wjS6:E���T�I���0��~�<y�C6d� �D�0�Ji!'@�<A���{|N8�&J��4��Ȳg�^]�<��(�0g��Q����O�$���G�C؟�pD�A�a���� e(��W�P'^2^� �'yp%a�ŖC, �P�
 b��0��$�d̰��e@0�S�T�^�9D��'|���CNZw,B�Ik����r�[)B4����G([��7��ny�$M�����S��Ms�aTq��"6� {^��hvb�l�<��LF�B���s��=/���b�e}Ը[%�`zLX$W�xro�O�@UYӅR�)?8�)��4�0>��A\4�(�3 �nB|H#6�ُJ-�]S�I8�6Q�"̗��?Cb�*��X
�-ۛi�0ܲ�gWg�'V���0�� �V`��K�wS�Ox����ؗ#y<�Yc&մP���p�'dP��bV37�,�b��I��dH�}�f4q�)�"l�jј�.�h��ދT��d)��C${O�I���8!!�D�5t|,��d@˔�|���g�DXA�����M�D����Ar��ϨODD�� A�
DV�g�R��E�Q�'u��D"B��ꉊ4�Qΰ3�f��m=^� �-�	ƺ4���C��~�.���0&Aa�^�ɢi�6��'��i���X�L��h�$m���yq�~p)~�6Q��̖�u���
�'�P�<i�lǄ\�ܴ;���,��4q�L��fIvM�q�]�s>@��\3WO��F���O����Tp��\�aL�J�"O�!r�K�qC3R�c�D��Q�Y0"���0�t� T9�ED�]��8�S�X��MC=s���A�Nl���	w����ׁ�b'� �rʒ�!��R;[L����S',Ȫj�n��l��K�<���VI���@�5��+�P�A���1�~�HȊ�$̤�X��g�1H
heS���P�M�A"O�TR�ȇy*(Mے)P5Vt�U� bXE|9���mTaA�J��>��4PN:Q���_�PeT/$��
�k%D���ĳ6���A�hՁ\�R`�U�ߡ^J=��+倓
�j}���� � Z@�n��6�܅툱�V�'U��)SM���}Z��K,m��d�b2"-�8:5��G<��$U�Vp<���\�za��?��RTh��@��$?i0E�F?�)Q��ϥ88�����<D�ؐ�r��E�פʆ0[��z(����%��f�6��N<E�-�=K�ݹ�nT.z,�&�2�y��Kl�ͫ�ܘ-P��(�<��I�q�8�h�A�p<q�-�/���t���?�$�&]X�� �&�3.1|�C��4BG�T#s,C�YH��6	nh<��,�'.��xa!��"��z�I�'9<pkP哋/�\s#24;�h��!�1�fB��R8P��B��Y�#�7/�B�	�� �v��B)v���FS�s!�C䉆g
r=C�D	RQ
La��2�B�H<Ix��U�b6�X�D�Z4C�I�8������9;�DW.>/lC�	�?Dzm����h���٠�C�`�>B�I�Zm p���䴅��"�33�LC�	�EX��ՉG���9�ǋABFC�ɔ%��P�ǥ�Jw�-��B��8C�I'"1xp�DL�kP�ע>S��B䉣8�P��mB� d49%ě��B�	=md����%&aH����0�B�Ƀ`�xQ4��������J;W��B�I2�I�R��A2���
CB>B��,P/ڍ#��P�Qӊ�J��]/h�B�	�K���9p�̳;Tv�Q�7�
C�ɥ
�$�p�/�_�F�b��L��C�ɌU�<(rϋ:`'.L(5
��R�jB�	3]����d��'Mi(��4�  1�B�I�^���Q'e�<_6(Z�-?w�B䉝[TDIb5
\���,�u'LC�I*;�4;v��S�@Ԣ��(<C�C4�ؕ�_23�Uq���$e6�C�	�M�d�a�T���!��Bs�<Xw"O (bj�>3j�I�I�yd4��"O�ik`珵*{�Y�@�еEa��R"OVmZ㍓�x�Ux$�
Nޅp�"OȔP��-i� l���,D�	9�"O܍�p�	�W$�d2r)���`̳0"O��$,�*��95�S-��ر"O�Q���2�@p���Ȩc�� �"O~@A�,�/܄�b��;��%�w"O�  �%ю}ʐ���pX.ͩp"O���I���m�wlؠ1�rr�"O�{EƄ%6c��PN��-x�"O��J��֥4��us+A�M��Ya�"O~�Csl��w�"�:K����"O��2C,ȽW1�����tn2�"O � ��B�iK�o<A�  K�"O�dqo��3T�y+2V�9�����"OlF��O�����L��hY"O̱�sIV	 ���K�E5rA�T"O��1gn
�D�MXu�?,��<Z�"O(A	�n�+]%"�
Ӄ7�Lt�U"O�U�vmO#�(��R�\Q&Ь1�"OT��B�9s.�Bc�Y�Uz!3"OT��GF�G�T̑t�8d���a"On����$Ze�$�e�$`�1BE"OT����Y�����oJ|)��"Oδh��h6�j��T�����"Oh	X�
5`�>L��O�U�^"O��8�+ιB�Q3'�B	fY�"O�x�Hϳ&� ��9y���"O� ��*�-%p��5�@9r��A��"O]�we��
��p��޷���[%"Otdp��G�PzEr7��.|��!�NO���z�_4W���e�2<Oh� E
�u���P��`����"O��A�#�2��a�P��X<Z�"O��(C�/��$���fu"O��Q�H��lY�������p5"O���Ĩ�����a�;N����F"OP=#&'�{��Aҳ�Y�A70��"OR`���VzDh�,�R0���"O�Q�pƔ	o��@5��.n�Y�A"O�tAʞ�h�`}�di�+\Z�3a"O@4��$̚m&��dK�&p@��"O�(è�N&�l�S2 2H���"O@Qkr
�oe|�2��5~�I�"O���\�4��A'��L�8���"O̘�'��0F���%W!È!�"O> �gDY�A4�0�e �M�.ٻP"O�X�ì�pjL��'�0c�"O�-���΀Ӗ��U�Lt��"O�{�K\���]�#�^�f�K�"O�A'���0{"��R!T�w��l��"O����Gh}8� �1 v]�"O�q�T�N�+������[gq<�k�"O6t�3jU(d]�l��-�-\�Q)�"O2�b���ڄ��*x�"O��#��\zD�NO����"Oԝ�LK8�xS���.u���� "O��T	s�����Я2����p"O�,�c�P�{m4�F�T�W�6�t*O$@h%�U��l5c�����IC	�'�jl
f�ѻz�^�A��\�S��uC�'g�8�e1!1^�����5~o���'��y��+~-��2W��~�lq	�'�D���<Qj���LK�G�|��
�'�><; �G5�(�aQ�.S� �k
�'��|8p�
u�Ƶ�`��O���	�'�jY"��P�z?"4P�B�@�`I	�'c�L2�bC9d9,h{B�%;���q�']�YX��Q�AJ䵙��֙/�� �'*`�QQ��=+$��c�;,�IK�'���gE�{$�e� �&f�x)�'�^��'K[�T��L�J>T���'ư!4A�nYrGÆ9l AK�'�t<�� 8�J�����8�@u��'w���UD6:�X�S�G�C� ��'%΅`U��2H��`�.10c�d��'��U��q`t(#�
�.��e�'߾�K��)mC,Rt�S�7J�(��'�	�&*-l
dMM�  X��'dу4�"�ɐc!ݠ:�iS
�'hx�aʡT)�w�R�t4���	�'X ��bk�s�:)�����Hա�'à�ңoTpG��p�@!O}��'��F/Q�CF�-qO��Kk��'^� �ef�����C.+�U(�'�n��O Jez9�"M� H��'Z:�h�י���L�	B�
�'�Xe#�ӻ��y�&�0l���'�l{�)W I�|�[�*ֵ_�2I��']NV�ZUA�<��FI�D�;�'��ܩ�&ŋ,��	�B�D�m�H-
�'Ȍ���cP�7�����H�3�UY�'.�e*�b�'�ܙa�dǸ�|�A��� tq�F�]�y���7��c*���"O�'
�	s���B�l�>H���"O��؁C�DK�اɂ�c�TP"OLuH4ǎ\J<�aj� /�l�J�"O<��*�7r��8��$��<R!"O��s��B>�^Uc!(��qܺ04"O�-�W%)T��\!W�(��a��"O��R��� z�e��+�����"O��Eؤ��E͏-kР�u"Ozq`@��)����>�<	�"OXs�/�k��IoZ/J��()v"O|L��i,j2j���GM3k��
"Onm!�"��J� ��e�����A'"O��j����<$�dӤ唳hz�`Z "O@Ai�ߍ�>YHd�*��	"O�СWj�.&��QK��0)�
xb�"O�M��M�i(�pU�[>E�֤��"Op!��,	n��W�:S�@� 1"O��P�P�nLn�K"HP�+��t`$"OX�pșm]�y�RE�#c��iT"Oj�b�@ID���s���M�|�1�"O<$��jY�Ŋ��/S� ��V"Ox)QS���F��	���-^<L�{"O��A ��qf��i�ݫo%\�c�"O���'!p)*����|��Q2�"OpL;�@���AZ� #�J��F�!��M��-H������u*tÄ]�!���,����'5|��!B
�!��		M�����X�|�=y#��!��];!}J��Ҡʭ���"�K��oz!�ϑ/�ܵ#�ڇM�.�����	8�!�Dʲ�.y�A���Bٱ�ɻ$�!�[�^�i��8�|�*g���!�]TB�*QꎅY��q�"H��!�D�D�4z%��P�F4K4- 'e{!�\�cH��%��`��ʒm16h!�d«B��죦⒚�`��ɛ1?U!�C������m[.{�ִ�F��=
8!�2x�5K�f�2-�"�H�iH�I+!�d�	ޖ@h�lV��qsH_.!�r���`J�f��S0��!�DK� � M�4U��}cd����!�d44���s⪙;6���T�!�!��|�Zժ ͜�+�h�IP��S�!� B����"U�E\*��� E�!�$ʗ1�Z�� �fX�9 �K3�!�	k�朸S�B#�ԥ*�W�!�	���"�#HE�d"��U�!�_�a�x� 6h 20��;WƇ��PyB�7LG䬸%���6f���y2���|���A�,��y�����y��B(1���@Ţ�#-�J'��yҮ�mi�� ��Y� a��& ��yb/O�Hfy�����0+҅���y��JH��9�Gְu>z��%�D��y��==Cr��4<{|x��n�.�yA( D1�p��};׊�#�0<)��C�V�=a%���ڬ�g[:@�!�D˲wKD��(�0��52��Z8!��ѹZbT��� D��6e��H!�	�J��s�2����3�!�$M.0��e	7~��)s�_�!��/!;�E9f�֭ ��E���!�d��8�X4 g�,� 6��ms!�� ��Tȕ)%@8i`�F�  �"O0 	ç��n+n%A�)�`���G"O��H4旘_�-:"ȍ�0Hz8W"O�p�ԇƩw0���T�Й9\�eR&"OHI�B�ի5|z�;萢Y���"O:`i�oy`����+.,�5"O~t9V�G!*Zy�F甌c�`�$"O�p�U�8{;�e�bK�L��i�"O�]8eD�0-��)I���¥�"O���ɑ��"	�b&�y��i"O�t�J�!  p��PL�$�r"O@���葕F�$8�π89��cB"OΨj�[h�b��w�³D�D��"OD��5�����.��+7"O2T����JʢI�GǄ�<���G"O�K�D�V�4ұ�K
N�8�"Oh@30޽�t��8�fd1�"Ol�ҲiОi� e"4iV[�θ� "O<�� �4jV�+�ȕ��z��"O�uKd�q��8��fF"P�¤�d"O�1��g�T@آ�� f��%�"O(M�A�F�\z��4��;m�x�E"Oڠzb���^zΕ��j!�-��"Op�"��ֆ~���z����F��4"Or��G�V !J�d9�
���(��"O0Ih�ƒ<"z���PIߚf)�#"O�$0"�?JpK�V�+�Z��d"ODpA�'��AY!-݆�z���"OJ ���Z,p�S�숾�n9ZU"O<� EёR:fc'-ց~~x��"O��A�,�ZP����:g�p���"O"l�,]�@5lr�\#gxl��"O�Q	TA�Dv�	�jSm*�"Ofeb/H�p�X���G&9S�\��"O��kPf_n��pp���$I�B"OR4�u]�S ���cE�M��|@�"O��	V�D�?i��@�ۂk�Je�5"Oai�k�9,3&Ɉ���:`f��zE"O�0 ���t�
�;� `�"O�qs��F6���<�z�r�"O&��7'�5ܘ���_�T�*���"O�j��[�f�:��Ô�0DC�"ON�"�[[����`�=0�ZP�"O ����
�5v��cm��� (q"OH��!� io����n��^��	2T"Ó3�n���tT!���&�~�9r"O$��6��J�(���Y�~��EQ0"O�����Rg�Qb��'��)r"OF�c�JJ!����o��j��A��"Ol�8@��A�!\,��H:�"O�! �'�(B�(��7{h�T0�"Of���
O�m�|y���c�����"OJ�qd$ � �H���� �"O��䈄3-?Z��4B_'#0���6"OĴ����'6A.����6|쀲�"O��`���t�f1�����d� �r!"OJ����z��Q �.�:'�BE±"O��C'�߿gp`!�U/A:E�|��"O<���Dl�"��0�Ā �K�"OiR����/W�!*r��(PMp���"O�EX��G)B�*�0�&Ͽq8heC!"O Pː)M�P1ҙ�be�!$�%�A"Oj�`Ʉf���Bd�F�ډ0"O�i3W��,d�&i�"��&y��"O� t�[fE��X S�h6��A7"OZ��>&\��3�~�xQT"O�t��19F5!E'ܹM|.8`�"O���K�,Z����D��y���E�r��EM��>�z����
��y�hH��y�EL�Ƕ���#V��y�G|��ئ��{� �R�M���yBg@>kp��rɛ�ulLh𴫆�y�l�:?,,	3���s��8�'����yr包呂�S�ؽ~��� �)�y��%)�)ۇ(�_���Ye��1�yb(��z��r$�P�r<zq"��y"NU�~���S�Y�O=�p�$ٹ�y���H�U��c�/zJr�0��'�y�L8
X���.�'lP��8._;�yRA�m�lHR6��#f�" �e�U��y�j�C)��yC�g[,T�%%ݡ�y�)���nh�֭M�W)%�4F��yBg�y먉���3PY�01c ��y��^���h"�P�A2���1Y,�y�`5�d��!8�	�#N�y2n �=f<��@�b# ����yҬΎa�$ 1�6^qvlB�N�1�y���D���b5KZ��uG_��y� Z{��5Ι�/���HC�yB�[�}�P{�`�:h8��$�ֹ�y��
>a��A�ɖ����4ķ�y�JF��7�݀�t���)�yL�"L�����6���)G4�y��&BJ�m�g
�Im�=KBg� �yR��),q�`�\9zeP��3�y�J�.@�0��q(��<�5��	���yB�\"uln��
86@Q��a���y�/�v��d�ӑ3*f�����y�bF�y�<I7��}���b:�y���2Ge�qr&.4}�<<{���+�y�fõ��t��O�q�dad����y��<Yx�L*FeAc�q3�O	��yb+O�L���X�%B �T����_9�y�CW=���F'*xmε�	Z<�y�nL~���Xy�|�;�$���y@�h�&�0��P�nJHJ��W0�y��;Vnm���\}F�i	0���y���Q��F��/���梑?�yB��
,�f)s�j�%N6��`ē!�y2�X�ߜ��Rz/�0åJ�y�/NF	�����˲m��X�4k̓�y@V�:�0T�����` 8�ac�W��y¡�xf�l �GPb��b��'�yBi�<P��Tp�����l��yb�I�<��4yЂ�'=����yBb"$�.��4�C�S��sׇ�y"�ų.�2��&�J1A�^�����yR�Y�p̤b�N��9������y���G=��3�"�T�YЊ�y�Οxi�3�g�(|a�"����y�������sLX���Q�Qa��y���/2�P��ۥ?h�J���y�Z�0*�Q��m��$��5pℊ�y�F&�:1�J�2�4�kV��)�yR��2٘�F�&�J[�hY��yRMXj�8�fO��8��A0�yR➬o5�9���۞����y��3��1A�^r���9�	��y
� D��1/ʶj�Թ�6O�.dY��C�"O��G�8���yîȮ5bj8�"O�Y�gO��t�T��Cn�:D�v"O`���SC�*��T,@"|��"OKGT�v �N��V|�$qf��yB.�
@]�h��!�<B�`�2�:�yR�U�8� �K���8h��9P&�y�D�q�D��M�]=��贃�"�yr�u��+'���h`�`��y��������1nN܉-Z��y��κai�i��i[()^�{�O��yb']�4���5)x�Q����y"��#H���A���l ��Ɩ��y�C��)��|RX:{D�ʡN��y [D�u�Ru\��",�/�y2%_&	���c_r^0M��æ�yҋ^.���〈dР�Z1M$�y2���?�"�V啒Q��=���Z��y"cǸ-�Lѣ�
NH��q�T*�y��T��`�����;�J T	�y�JV�,K��J��K�Tpm���R�yҏ�7�A�RLT"[^���5#�'�y�Q�H#F\{$�)O��e�4��"�y��v�Dī��B�pd�p����y�P�sdH�jr�`\�����y���7���0�U�NQS$�y�dY�@�>츱ܵE��|!��/�y����LAЧ�6%l��Ɠ�yR�7|�0x�t��)�:h�����y2�t�� f`�&^1�V�]*�yR�	����̖�9�Y9F�ۘ�y2�K�m���2fCн
��݈bF���y�l^+o�a�S	�$���K�"�y"��=�}A.�>��a�׃�y��G�5��u{Q]�9����u���y�%'0�r �Q��|����U.��y��%���R�J�|�F����yR���<�!�Ň����O��y�`�;ko��D�(~~�4�W
B��yB83_h+Q)�a��]�'�9�Py�ˢ e4�bB�O�fʉc7�J�<	���P�Ȃ��*@���@bE�<!�	�yB�pz���J��T�h�<Ia�D���,��*/!��  L�\�<�p��hS<I��ޤv| q�s#�L�<A��� zFx�'C
�
�؉JA�@�<I��GX��-��q��1�>�����(q��ڐ,ҀYq�-w��@a�"OP)Ja�c�6��9#j�lʅ"O0I�l�&�s���7Q����"Or�K���^�`��w�%Cc�e["O��'�E�W6�I@��-?}�ubR"OT�wQ�o��	PЄ\�ku\`{�"O������l�ٻ�(h&�Kr"O������H��ƣ9
X�"O��g�!����ϗ�G����"Of��F�U�/��Yp�۳q�T�"O���კ�%?8�#��9��PRQ"OtP9���>c�!���?n�f��@"O�8�L]�&vرР��g'4$ �"O2�!�8�,r���)�H�"O���O�?SkJ�*�����!��"O赡��{��i��� ߦm�"OF�I���r����tL�w��8�"O� }�s�	�^8\�{G,P��rI�"O��s��۩3ʩ�Ə'O�b��"O�}�� S�Qq��A�¤@"O��F�N�8�p�����u6"O<���%�5�͛��	rC�h��"O�͓�Nn���b$�_;PY C"O�"M 
2Eh⼲hy�ESy�<C�Ľ:#����\�12��#�K�<I��\�r1�Ij��
0s�N9��Ä~�<�W���2�xْ��E�C��lh2�	~�<yP%ͼ,A�@��Zx���3d�I{�<y_X��#!fāA�CߍrsB@�ȓ)&�x���B�~h�P�&IIOr6نȓ]j��/��Kn�$�rn-#`��ȓw@ �h3阳�r!w��Ҹ�ȓ�l��ԫ@�_n�@�7&Dфȓ!6�00g�̭M����q�q���w�pM��Iʂy��Άm90|��wlH"7
��	��yZ#�"ybP��ȓ� P���7`�zdz�m�k�q�ȓ��a"Bm/wF�i���=5d��ȓ&"�A&�S߈����R��rŇȓ����]������%�`�ȓ}�������-�;���j��݇�A���t�W(nq����ȎQŚ��ȓ=��q@�V�N`����Y
�����u�h�j�Z�WR�*u�
}N�X��[�!���� h�l6��P����A���X1A*ġr������"O�]���ڥm`x�Q�+�"W�["O�9���
i��Y��&|3"O�db卋D�P��t��t8�uc"O��bF�L(+9�䒰狗
T�"O��%ϻ{
��RG�{ߦ��f"OP�s��X�m���*s ����"O0�RiY�.2e��nY��j�S"O�PS��>�hّ��&n2�5�p"OP�2�	Y�����x<���"O�-C�A� :�)B\_�b�r�˟N�<A�ܑ��� �H�6Z�h��,H�<��F];�B��"����q��S\�<��  ���` S"=����̚T�<����Z��cb��)ҖT5$PP�<��i��&�^����w4�I#���c�<��J��G,<J�֓}�0�#@D_�<9��$nv�1�o#���B5G�<�#!�.�@5j�U�����^�<�T�*`f%qB�
 .	���]X�<��ͨhh��㣣��,�S��X�<ٶ��"-��q���Q?��c�!KQ�<a�M\�J��@f՚6)��كC�e�<�v
���֐�� Փ�@=iD/^�<�P�qQ�x�5�*o2� �"�\�<��u�I�Q�Y(>V\��%�WW�<6�J�N4zh!�W�x٫��h�<y���8L M�wf�rX8�����m�<9PKڗg�j����9\Gt!a���j�<�D��_�$�J��ùy��L�T��g�<���#nTe�wF�y�ڱ1!o
b�<��D4Y�t�J%���&����m�[�<��G@p� � Ȩ�+Bi�Z�<9�KF���<�͇�M�����X�<��ݸp�,�@��O�K6�sba�U�<��	v��p���wv�T�B�U�<� ��RǭJ1I�13"%S�D�v�D"O�Y²΅�"�`��G���V���"OP�4d�+YȞx[�S@ڴ�@"O��"��U�@n��:�g��-Z��q"O��A.͒Z�b�X�ɠPR�|*g"OL�i��	�pcDM�H��¶"O�l��_��y{B�R-V=:���"OT%����d��`��@�Rȴ1�6"OD�j��>x�
mN�a��lZV"O�Y��?Nq@)����G�p�1"O��q�E	����m@�.�B(Z�J�ON�{`���M�O?�ɥ\�긻��מ6͈y�e�˶	 ]¥ã=:騀��k���#&�8h�6�>I���H��/��LL&�+��V�nJ1�g�i8����A�Rm��0f�n��b������4i��s��#����S ��3�I�u�i��y0��'�2�f�p��/���{�)�@�,��@��="���檟d����̅�==�xs-=C6uy�0T/V�<Q�i\&6�,��޺��B�?xP[�@F�
�]�c=+>�'���# �`2r�'b�'�םΟ4lZlbX�h�e� 豉��f���Xt��mpXX�`��/ �Õ�W��bUA�=241%��'��2�d߈Cs�O�,� Y��R�9��8����&�}�8C�ȩfL9��'̑9wn[�59�$J���#�%����O�QQ�c�Op8lKt��<��'����І�9��RW���	T��w!�dE�t�z���J=t��zD䊺@V���4Qd�v�|R�O��tW��BrK��p��e��`G�Iz�q��,�tCv��a�Fx�t�ɛT;�ģR#כ)@|c,�|AJ��L�:�X�R�C�
ƮE MY>����(�LQ/B��EB�!� q���ut�*X�.av4��44�QɒiN�^2��
4� ��_3�����?P -)d.M�i厞nĝY$P��M���������?9�ڟ.�aPH)C�@�@r���`3���q"O*(�
����[�f��	6P� ��O�lZ/�M/O�xBc��̦��	�8�O{*��〵#�x��B�	6�l���ݤk>�$�O&���0ݓ�E�&�����E�+[4���L�pa���Q,�)�c�DhU���]�'Hm����b� �� %���Ƒ?�He{��ش�"0p��H�l@K��*7[d����SQj�~�V�	2�M3w�&��i���K'Mߪm�h@��Is^�	$+�O@�"~���*{�T�3��4]�2��5�f_��$Ħ��զ]:�lӚB�:�(O1u� ��b�����Cۏ�MC���?�,���T,�O���x�\����P ք�F�t���s��E�Y֩ !� �jAh9!TL̯s�x�t�\�4
����?�����U(k�$��H]����:�G���#v��t��u
d[�j�$�i�7i����%���g\���5v�^2�@A���Ns �r$h��M{Sf�������M����f�s�ā9e�4:U�C���<ٱ��O���>ړ��'���D�ҴIa�����O�Q�ȑ��ĝצqz�4�?A�i{ҏ̐dg�0Rl�"f#��I.>�a��"e������s���mJ��IП�����!_w�´iC�M�� ͺ~0d0! �[֒�P�"=*z ��D�%��լ"A����4�}���D|�ml^�!ȕ�(���SGރ< H��4yU|�2���|;��S��JP�혹'M>\���҃$�dP=%�py��H(ஈq$o��B?���_O������M�b�~�'�BV��#���-Jp���W�L,��b���>ؐx�C�uC��z�NZ*�*���I�M��4 ��V�|\>I�>IѮV0 >  �   W   Ĵ���	��Z��wI�/ʜ�cd�<��k٥���qe�H�4��6_2<<�3�ʄmn���s:�j�����Q�e_�c�7-⦅3ٴJ~�*�	_y䟛nSt���|F��Gb��*pH�A�IP���=Y�D3n�d7M�0e�R�3C���*���)�דc���(�Q�d-�.6��ɓ	�����ƌ
=���&?�,PtA���wL̴_��e�6�^�A�����X}��
W��P7�x�ϓ���{�OY���q�v*]*�ʐY��\;0�I��y��& W�����t
�C���Q��Փ���$�f�jd��$Nt�;�ͷ���ec��7�F%a��<� ��0�x$�<�Q�d�Z�,p��"D�kt`��c��컑�I�}D�i�J�Q�Ra�e�\��m��O5�O��Q�O����$��������YK��>� �3�\��RUk�%Z��1���@�
�nӔH���O�T�ůC��~<��^q��ȉ�&�/*W�Oܬq������(o��Za��vl�b�":39�I"#�PK����'���B�
�XZ(�\�EI�O֨9��˚�?���'p	���=e��7o c�Be|"<YEH3�$0k\�0�n��
D�(�a��/��dƾ�O\� H<Q�OlA�[e�`��bC	�F������'�Dʓ$����=R���O��Ē��6�O�-uj�:�O'��� ��L��'�`|Fx�#�s��&��T�pÔ�M��z�	��@��I�Y��H��I!E>qq��s�<�3k�7#stB�I�e�l�  �5;vZ4��"O0��7��o_>��Ǝ]82���d"Op�Zg�U$�����Zf��:6"O���U�_�<yR1��$}���"O�@���]�0�B��jx��"O��4��9/����]3"O��r@"O��bFւSvh!A��L(yL�Ě "OX��"ၹP���DN�$��09�"Ol��4L7�qJ�ʚ�n��K�"On$  �
k��d�'H�P��u"O:���,,KZ�Jr׻"�|ّ�"O�m�FÒ "��������P"O��0C�؍���c�E/Q]P���"O�噇����(�M���
M�'"O(�U!��|�'�͜w5�3�"OZmyv��nmH����>{,$�x�"O,8��;]H�ۖ�ސPXш�"O��r�� ,~�Q���^����"O�T�BP   h
  )  �  @!  C(  �0  7  V=  �C  �I  ~Q  	X  _^  �d  �j  +q  pw  �}  J�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�
�;�>O�1"�'"d:t&�����.}�ȕ��4��DK���8pp�hICAP
;��i��fݕ(e"��?���?j��~��e#�HծW���d�9gCL� �+_�Z�SfF\Pbf�b��+�u�͓�(���'�b��F%��%����)Hk�xÕ��-4"r�+K�Op�J1OS�#�r!��������"L�����������{'!�9�a���9i������D����ɖ_�$��޴���O�݊����t���O���!��/T��}��#�
�#�"�'���'��C��&r���?)�'���D�{�H`��5��Dc�ꔃ,��2<O�m���3Ւy��Q1�"��U������~BeǷ~Z��O8Ȉơ�l�ft�r�s�p����?���?����?����?�+�`�65`� ���6[������+��$��u1޴=����>u�id��
%w�2I�B�O�������j.�J�O`��g�~�'.����iL�Odrx�%��=�]c�զ}��$ 	Ɨ$��� �̛�f�Ni�Źix$7- ��S�?m�0%?�$gFF'	5��)@�S 	H��Uƃ��M��fIy$|J�cH�e��x�Ǭ��n=|�Q�⃧=�6�s�<(oZ�i��� o�"-����5� �#S-ܴU����^��Mo~Ӯ�mچ;�����^3 9��Z���2v*R�5Jb�!�%I ?�3�+� �"�k$�AW�d ڴ7��*hӲ4�Û%H�����-X�$��4>ZF���n�z#�$K���>i�}�	�b��8%�K-]�ʸz��~-,��'C�O>��S�w�L��2�V�p�*�R�I�O����	��H7투�M�̟@4�q�\�^�����Yw���'F�I���	�|�%b�aH��!�߅1��L:�4+Xp��DM7,��Da�c@=3Q��9ÓZ�f#�5,p���I%�?Q"HI	�e� �A�Svz1����{���pm�O���XMy"H�
+��1�B�o{������?���?Q���d>O8�ȅ�&`� �a j�AX�92p�'(
7��>;��r׀��f�(��F
�b��l�Y�������OV���T�ѻy�����[�`��r�"O0��e+������;\�9��"O>I�e�<2��|��[6��k�"O��"�D�+�&�z&	H�����`"O�={G�Ӯr%P���i�s��Jt"O�4J"dV:0��s��A;T�e�5�'��X����(J!�D�=����9-���ȓ|��q��<RۆMC'�5��ȓ�X��wg�3@3ԥ�H�&;4$���{�*Qi�鑻9v,�:���!ժ]�ȓr;nqy�IP��>D��S�,�͆ȓ?1F�S�A���"�l)��O�<���Qb8�x� S�TǺu����RD^���$D� ��NH%n���@�,`�uk�C.D��#F�W��<��Th�'W���)D�DPQ%X����sJ$C��4D�0HDd�-���6�Ⱦr
�ye*2<O�H3������I�����21Y@k�����b��4���'���9�'[��'�\� s�F�FA�6i����j�J��t,��9J{3 U�?���D�<X1BUPC�7�v��a�.H%�i�6�Y���E{�o��-3t`3��'�X���?�'�iYR
���*SG��'��z���0q#�՟�?E�dL��'3r�`q�� m[�Az�b���'Z�	H�O��7m�?Av����F 8KЎ��2C�|�oZv�Id�)�'QU�����Z�L�KpD�uh�r ]�yL77:+�B�O�X��
5�y�M^W���ʃB	�t���1p���yX3�L�p��
<V��D�ˑ��y�W1Lv��F'�UC�1��V*�yb��7W@=a-V˞i��C1,>���|R��e_���' ��'T�+a|nԑp��n�����O�6����@��M���i�8pZv�@$U�S���'��`��cEO "m%-��«<8"�i��M"�`������O����ƛE?Y1,։lZ�Z3�6G�X�ʔ��M��R�4����Ohb>�d�O.��@�2Z|���EH��L�7� wB��DPG�o� Y���D���%�P"z���'�F6X�)&���?ɖ'�Z��V���J�^������vM����H������'���'	Үݙ�I��t�'S}�	�Pe��2�z��7�O%����?9F�P��J�.���Z�Y���"ANSU`ȥo=Sǃ Ww�捨eiT��ϓTt��E9|�Q�QK<MX��E��X��̟��?1��)��v�	�m�4۰e�&[k�!��H�'!��`+M&��p��c��'i7��O�~]rA��i��S�8��
s��D�Դ�e��.u��$�<9��?���<�*��"ա ���&�Ɔ�y
� ���S�?��$�્<�<@�E�'��y �#UlM�t�''��yB��a��+g��P�V��@�/�0<Y���ݴ�?���c��R�dL�s�y���?�@I����?����?����'Ø'�
4�d�"���ZS��./Wq���s<�M�N���!00,�u��[��?y(OXh(@!�ߦU��럠�O����F�'���{ծĶ&d��[�]�E��c�'�B�P�cB�T>�'Tp�r��t�كo�n<B���O�T���)§k�	h���6���ѳ��/'zB��'j�1��#Bɧ��qC"g qݔaӃ�ѾM�jQ��"O`|kǇP�x�-CC�$:p�r�ɠ�h��TQ�F�>^&�l���&^�B0��i����O��
�E�*~b�'���'��݉1�|�eA]�\������ҩh�(�HZADb�,߉#�"��4�S��%��'���UhK�7T�A�'��d0L��J��a�n����oL ��f�ĸƘO)�9�Ic?!��1B�ź���$4�4ARee]�M�dS��٦)�O���:&������*Z�#k��TG�\�a�S�<�Ed�2R����K�H�v�Vy 1��|j�����P��N��iM�R�@\!CO�-";��y��ڂw����O(���O\쮻�?�����!%WD���Oڇe��!�"�#x�iS�'��%�K�2kҍq�N�L�ĩ�C��xRcK�1�B���F��:'
���Ģ�Ҝb��tc����Sk�m��ɇ.�%�e�_��y�-(�����H>[x�������$��&�|R�
�YA�'�?ف��<K6����%RU�PU@�?1����XB���?1�Oer�R#L�-c3\�F�FD_B�la��T�q�ne��7G���e��0:��3e.�c���?�DA
DP��#�rII���]�L� ��Oz�,?�TH�fņ0��%�%�I�x�ܒO��)LO�=���F+FA��F#d�P�A��'���5��c�É"(͌T�2MV;;J�\��Z�ʶ����OʧU�4�1��K���c")C����C�3Q;�|h��? bQz�2���$�,P�[%�V��O��S�0������E��1jS�R
9T��'��u��',��� �Y���ݤw��{���3�TJުby���K��c���� �'"��3�t���wӈ�D §o���c�P�mJ~���j����&���Iʟ���{y��'*��,N]�p��oF�N��`!�9hT�?�u�i��6�.��2)�b,�!$Cs\��P7�f,o̟`�	̟̃�(�z����I���������yJd���Ȇ4q���<�4�BV�.�^�C��I�(���	H�S7~�'���m&҆�H��f�5���^s���k"��d�
��f ߲<��Q��Z>M�W�ן|�>�C.0T����eJE��j�85^�Ul���M���T"�������D�Oxxp#ύ4��#�W�Lr��O���<������I�-b�YSm�&B'��!�H,74�Z��v"fӀ�O��'���I���tQm�('E`U�G�1@�{�J��+�f���O~�D�O�p�;�?������ж��$��͗�r^��#�P�Lm���!�<уTgȀ7�Y�6	��+� �Gyr�O�Ks�B���,�iQ�S�|R	ہ ܫPK� qNߗ?`�A9��ب'aGyb�Q0@�vP9#���)�P�_�|������%:��O�q����^�h�:t�
��� �B"O����R
X�f��� �[�T���|�t���d�<a�K� |���ş@�Ǜ�&��IŦ��h5P�;������I�a������Χ�b b��Z�[�hZ`Ć�fVQ*ffT�|u�rd�x�R�P���:ʓ�Hѐ�b�/��̊��	�bbnm�R�M5�e&S$X��h�1�@�2��X� ԑN�Q� ���O`l�����4:ҖmIaP,<�!/σw�'Ca| Q�Nf���)��p2�_���?�4�'Zb�yfMĲ4�����n�аr����'�J9���i�%��@��<o4l�HQ��`�k-D�DH�kU\��b.�d���p��&D�X�qF�(#ؑ����0�0y�E&D��0!Si7��p�!wˈ`4�#D�<B�,�}��{ua�S$J8[�� D��I�ܽ7~��e��&���O0 ��)�sU���N?�y��|Qp!�'�r=S0暇C<d��&ʓ�o�z���'��HCV �hP ���e�`}I�'�p8&�%<*E�W�a��`��'��p�CFڷ:ڨ��g,6_P,M	�'���j�lD2F��0i��^�$R�U@,O��4�'rq���G�P�Ȧf�;�8ę��� ܹң��T���Sb8��9��"O2�;e��5�Q����_��Y�"Oޭ�&�*.���`̥>���c"OV�93��+#+�A('	N ���'���X�'�|*�6h�@1�6�N�"TL8�
�'o@�@t��S�L)a��������'=��%�j�@U��7%�X��'SX��A �={_�y�� N�*դ���'�8В��j���Z%+űMٮl!�'J��5�����U�D
L8��8- Q?]�D�;g���ဧם�b�j7D����N��B�X���9u���sPL8D��2p��:<+�X�0w��-�P$+D�`���(e(�dxǌS-i�P�f�(D�@ U ̋X�n Z@㎬��i֩*D�p�d���2N�Dz�-G/Zߔe����O&���)�'6����s��L�p�����1V��:�'�� ���9�41�%���.x��'L�św���<��9	aM�+���0
�'i�%����$<�J��`�κ$pU�	�'Q^Lj'����d��B�"�h���'e\ۆ)�!3��$RG	�	�Y�.O2q�d�'�)��ޭ~��k���4|��Y��'���+�D�;���P#�!oDd��
�'�`��5'��܀�B;q���'���xS#�%\�^�X�m��ֱ��'t���s�v�J���G��H��8:"����X�QË,\����P�"�*�ȓ�I� &?�ʀI��C3��m�ȓ\h����Z�
�!�EOl�Z��Pva!,[<&��X"L����%�ȓ[~e��`֧d�^�c�lkZ^���CL����Ⱥ.� ��1�͜-W��F{�$�쨟>̫ ��%d�[��"]r �g"OVmZ ��v ���T�.mP�H�"O�	#Ub�'�Z	[Q�S=v8�-	1"Ot� )�*�"X�#�
�G�!��"O�E�sϏ�*��i�BMY7!Q��"O �I�F���m@C	��B����'垙 ���08Ĺ��N�!!4I"a�U����ȓ_A,Y��R�d�t���6�"U;T"Ov�[�8�ҹ�(�*	-�=2S"O
	kpA�$I2�#s�I ��a"Oܹ8fnC������&'d���"OU;R!�?֨Ax�j�i�^�Q�\��X�"�O��k��?�,�������"OĐ� �[�P_N,ix:<�a"O���@ܑB�dɡ恇z�>��U"O�=�@["}��W�đ���a�"OޜI�h��p��+��u���c�'RI�'Ψ䙠�����q�@H
�'����U3Q.���c�:ix	�'�̤)3�̓~(Hܰ� �8`*�3	�'c�����`rT ֯�5y�����'鼕������*��p���>D��@�k_7Hyz�ѮY��˰�"�tٮE��NT�R����
N�$�y2�ҋ�yB��L�L�D�?9�T���O4�PyN�V�,�7$X�;L����C�s�<�G#9���A�]�3�0!7�i�<qB PB�z�T�Ʊwp`��AO�e�<�£�`Җ��N�(�� Q�F��т6�S�Ox����Y�ak�u�㠒$wK�y@R"O�=��ܦD���#Ƀ3%,\`��"O� p<����6Dct�C����U�8i��"O�T�5HL|�~����W�D��|�"O �8�N�u�B�R�G�+/�ZL��"O:��fƍ �\-)'@~��+�V�؈BK;�O\�y&��"2�� ��՗%�.,0g"O�$c�
+ZfX�ZqF�6��y�a"O
	�w��-o�� �M|g���p"O���v��:�����X@I�r "O����YpdB�9V���@�'�z)*�'9V���\��^���(�ܡ�'��5x��\� ���a�R,�j�J�'�2!��DH�_j���M�x޼
�'@�`�DT�s�}���ZX�6Hb	�'�t���'@!d敐�g̛Y�\q��'�8ؘ0�Z�6����ˎ$Y�b��dޘq�Q?�t�MCE��ÉH$V�\�K4	%D�@g,�;KWZ��B̴WV�a�#D���K��9Q�9@�H�7Jm���%'T��aEL>,t���B@�����"O�0j�I�d��T���h���"O>(@�
�I#i�F�C�%��Y���'.V}a���S4{��G�T|\j0��.�%+#)�ȓ9T��1 �h��D"T!�ȓhFZ� �1Ӏ���}�4D��+�R��#�ӧ�$,@��}i�цȓY���"��7�:�S���5H`&ņ�}���p�b��\��|C&k�3 ��Ė')�x��p9�9��ےDg��b�fر�x���T���h��\�bp^��G�	9�Z��ȓ�|DM�3s�fL��8���s�($c�oM^�@��фm�P��xo�� u�౲#I�!�����^i��	1B�����ćr�B����| �C�	�L��2 \'hC6��@�8��C�|	|u��Ɍ[B��b�%��C�	���䣵�ȅb�(���ªh�xC�	(|��[a�,�8�p�#���
B�IT�M�r���U�:@b"&A�H��=���|�O�$-P�
Һ-u:(�eж$�Z%��'�^$���Yz���mɞ����'� �!� ������W�~`�y9�'l�`胎;W�8IG�	(r��X�'�)����>k�xWU�k�T��'p����!a���"�5$9`�� ���Ex����_f�b+N�r|p����˅<khB�	�l���M*~<qy�T�D�C�I�f����&݄Q2vm�oч2� C�	. ��#�L�(��KL?�B�������ޝ@����!�f�
C�	�E�Y��Is�iB�R�p��ʓ&�2\��ɬ^�z��t��C���;%m��<RB��,
^0p�Qz�����1�JB� x�H0�5{��� E��M�$B�I�g?Ԕ0�̽x���O��Y6�C�	�iTU@N��F��['j)fS����̖����"-����%�9^��h#D�!�]�(~(���+-��Y@e�	=_�!�$�Wd&���
m�yӦeI�%�!�$N�C\^���� oXpX��ÀZ?!�W<<�DQ�I�&B�Z7�Q�!�d��t�nq(u�&Z��UpWh�5V&ўd#��"�'v��bE<6	Z̰��Y�"
Pń�)���%/Ja� ��C�I-O;�Ą�to��u�{f!����,��S�? @qHS��%J���b��F�Q�Fp0�"O��D��^��)����v}X���"OV��T�4[��T�P�C��*�1��'�нH���S�D�Xq�A�[f�t�����a� ���'�)��J�D���H���6��1��E���H��}sPٱF&j�0�ȓl�ĸ��.�� �B�̤��@��(�}z��ų�*�A�#!X����������GMȬ��`�"����'������j�RLL0dm��1,� KM�I��A����� �� 0;6&��d��nw���gP��T�'��H�ȓ(byצZ5Dƶ@"���� "D؆��<��섵0�������a�:����5>��	�}9��CvIׄ	��D��D�UN�B�	�"�d�ҧ��$���A&w�vB�I�d� p3,
�@�TJѢI7�!��W9k�ʸz0�Z�a�@���J!��{��
�BR�W�b�c�
]!�DCJ@�Ȅ�Z	R��h�587xў*�;�G4Ld�e�"S�lbsh��!���A��C",5�5�¤�5Bǐ@��Bm�$�cG	���IrI���$u��wHȲ"�=#�ةy��J�3�,��#�L��̶nTH%���?޺�ȓ8���?o`�30���A���	�O� #<E�4��4+'h�#L�1T��,t�!� �9��,b�v1�����!�,Z����ʜ34�!��\�xo!��'p�y�� !�r��A�WY!򤞲w��h�2#B�##�(ܡ��:/��H�H	�0t
�@�v��#}RH�<i&�^�IB6M��=����<T:%��=*u���<Df�¢�O8�9d��O�d�OZCf���t6�퉇-�
dS�e�d���s�J�~�P��'eT����`�Q�0sekؕI�����<+E�QH�L�W��i""A�4`���[��^�X1(Q��%ۼ|Q��C�g�O�o���&jVT�����!~t lKC
�D�'�a~�啦ciX��r�\;���ê�.��>�4U�țTK�93D�lQ�AQD���J��+�� /V&0�?��g?��IصsN.��DĆ >�^A)���j�<Y���5pRP�Տ�4� D�O�<1 �N��{R`��8:q�gSP�<�ǀ�wW(4å�ڃ1����X�<�G%�A����'&�@dHy�<�@*L�G�x�2)�_��l��I��u[<#<����O0Y �gշ$+F����o9"�c"Ok��*U���I�@I2J\���"O�5�#���"-V<�P3C߈���"O�����Q7Q�r�8r��2"O���.@6��ź��m���	u"O �7n@�\��h��$xٶ�p�'�I1
�0D��(�CO���p鈵jPp����t�c�U#TYBM:��ȗG�����N�:<)C@�*e��y�E�e�n��|`*<��慷_��`�ģ�vP*P��2�A�b�ME�y'N�?�<���I'j�'IaKg��I4t��g5e^A�'4�*�L�)�%xW�V�*��3
�'R@A�ft#&�;��F*�	q	�'���!"�"���q��4
�]!�'��-��׳���`���;��)�'��R���(�*�q����������Ί�O�;$�[�E�	P���55��ȓ]؄���E7���yd
��@��D��n���
�K�C'Ly��(�,�����S�? �t5Y�ZM2�C	 Q��xҴ"O�T����_#bm���I.�T=ʴ"O>-�gM�-\d�3�(�-���c�
-�O��}�0-4̘�<P\��.̐t��	�'<(x�$+�'�)�� �"]�F1�	�'@Lx���+L �"OQhҜ��'8���� ��c��rC� D
�'8����X!eݦ��H���T �'��QbG�W<)D�M��a��@]���	�8��I�y��u�f�ϼHS�ճ)��7i,C�	�O�du�#鐭��9�Cj>#�B�	�
 !�&��KhL3�*;U��B�ɀ��1�V�G�O�V�2�Mɱf��B䉧{�>��!��4v�\��OHp\�?�E+ڻ��	ٟ��'h�d�(Ï�@���`@n�=�(������	ʟ �I@Ɍ��Ks�@u�h����l��(|q�tk�<(�����?K� ���:�4H՚�m'�h<yרG�y��q�" �M�
 㰬�R��Q7�ظC���RkQ��3���O`�n���'R��C�j�l�燢BH�)5^�d��I
@���p�k��9���\�%�b��$�Wy� 
`l TgH7���I#Ǿ��$�O��O^���-?�a�1�,�k�'X<L�J��Q�'�*�}���O�P����B�:P�l��Ib�O�6�%�\b��'����N�0��w��|;�E`�!T?l��zy��lK�S��'�pr��)3��L�ո���W��q�ɫ��I�=�2�'d �j�r���	bcP�Ӂ/�~؈#,����I��~��s��9dn��Oq~�����9\5jcEM�.A���'�X�',2�J��Z���u���j}�0�q�Й���SQ�'H��PI�P��4�'&�lb��N��z��rc�Iǘ�@��5��O���Op8�1�>Y��i�4�(���0-������S:#,O�@���>)%�S�t�"Xxf \?�1��^
���:�'�l��H���<$SP~,6�i�W��O�L�H �Ǣp�8x�BS��Z�CAڟ��	�{��>�1 埖g�0QҊT @c8 sA��O�Q�'�
#�'���y��ً�~Be�*,�%��d��u f�z�Ɍ#�?�2�;�O����-�8���폙l�nU�"O`P�d�9>x�:�j��Iʜ���i���'����h�I_yRY>�XhZY�7�ܿxi����h��6M�O�˓�?��V?-�	Y���'aZ����-w���P ^[�Hy`A�*��O6��Sg��J�p����.��Q0'e�!��Oؘ�z'�� �xt�'���!�$��VǨdxd��iS(LK�DN� �!��-Q90]
v��'��c�cعq!��(�,Ta�D�jE���;X�!�D1!H�3ǃB/>�x�'G�m!�YPr���%�Q�Y��G�5jM!�$،f�����C�C7� ��E�X:!�dE�3 �(�S���T��1!򄝯F��q2I�6�,�	wDUA�P����?��TnP2 @�9�o6(ON4��<D�P�4)�	\�(s��x�(���<���
��8'A�&xA2@�C,�3B�i ���~="�D�X��P��)�Zd9��4va (%A��Ҡ9"+G�% ���TA�ln<�ӫ�ު��B�.B	̀i�[��RQ�N�9�EpT�J�l���˒.	�OE~�X��A��A�[%�ɜ�LY�g�!�6ypܴb;<q;aI F�V��5�T�+�X�)f�'�2)mׄU�P�;�T>�O}�5%�˵l�v�a�-E,,*@+J<�"WjX����b�<W�F�����?`	��\,���>C�Œ e;�z�ģ�i=�'����3ӛ6�p�d��<�SL�\��Ǣ��Q�CK�F���NX��04K� �h)��[]rZ� "0O|�Ey���	H�Q����Tߺ���m�"�nqj���O��Þ{W��
����}�"aK8B!�D �CF~�K6.^>E���WV-�!� �<�r��Q��{����eD!��T�`��=�7K�2�𣃍�J��5�r�e�E50�΁��hކT�v���L��@c툉;K���qBT4��h�ȓe�F=�6��(:���� !nm��S�? �Uc��@,h�~\�U��09��!�"O��J J&z���O�(�Z5�S"OR��k2�X����w�P��"Ov5��a�0�p�x�L,y,2)� "ONP���
vj�8�]0�i�S"OPC��l�:����Ě?��E"Opi�M�|�8���\e#F"Of�8�e9��!Plj�"O�|Y�!�4ji��)`�-"O����u�$08���+V찤[�"OX5j�dN�'/�a袧asf]��"O�$xp��R�Z@X�`�V�~�G"OZ=��+ pq�J?6�tre"O�E���	p>�P�m �M��av"O��)�U�h�0v"H�p�12"O���菣v6��#Vb� 褻T"O`I
� ]#O���z���,T����"O����\�J�b�.T�5*�"O��"�$ (]����uK�4p�bR!�$K6"ǀ�
��Ve��MGŒ$R�!��&ƠE��HþN'�i!�.Ob�!��"ߨQC����@4 2o5!�$�	b�p�*T��G��
4��@`!��ʱ؁`��;F]2��@��!�$�V��aj��˭E�u����!�DE7|��r��Xl�)���!��y�0j,U�>O�ai #Ϸ'!�$I�My�<h�Ò`A��K��!�D��S����o)M#Hp±�6-�!�� pĚ<K�JV�)P��˙!�$�/7vn�r�
�U��H�b���F�!�d��Bp�dZ���;�P�;�-UN!�dU�p̘��Ǘp�<�O�l1!�ہ�T��t��xv���*̨B !�� {�La4C�;Xo��ժ(8�!�D� ���cR�,E�(U�C)�
G!� �(e���U�ma�Ѓ�2!�ѷ
�ީDB�rΕ�ֆ��!�d\$���bƍHk*\sGƎx�!�$�\�L���9P.,0��d�%/!�d/�f����P(�C�$�%}!�3@ٲi:Ҍ��8��+�A�3�!�D�x"�!�IͦA/`�2�� !!�N?o{�]�p/	Yv��րB0F�!��?C�J4��[6g��rB�ТS!�dV=^�����鏪#yj�)�O�1�PylF�]�T�;�,�a7�a����y"��2P��(�"a��Z�L������y"T2�ܕ�����j}R���y���3��Jp�@{)���"�y�(K�eGn�� 埨y;�u�����y,@�d�R�An�j-"b��=�yr,�*)<z�b��Eb���ɡ���y���8O
��ҧG�
]C��E��1�y"%04��)���N��0��&�y�L	5S�8��OR=Nčhtş�y����W=2����Y9@��
5%ڷ�y�+]�25�c��@�rUS����y��Վ@� e���"
����/�y�D�?H��b����	A�k��y�i�N��!�2LLi,��`�틞�yB`�)��<S���<Z�5�b*��yrM��m ��4�>S |[ₔ!�y�*ϙC� QQ��Z)Q.Z���ā��y
� hX�r�L��N"%�O.y�mCW"O%;�� a�Ae�7v���"O��)F�JYRf�RD������"O2�/F�5���CX�N	����'^�b��dVnUP� ҷU4��	�'�����٫.��l�E�XK,�i		�'�������^+Z�x��� C����'��6/�0H��GC�4vI��8�'��5���R�m�N8���aid��'����չ^~5�,��Rߌ!�'HV�XBR���9QVy��'�^��V�T�s��3e�E0]�(u��'r4y	!�x�r(�*e�v�
�'s��A�o��G�Z�{W-_�'2���	�'J��F�Y�d�@}��ѱt8�4�	�'S�r�Bq3`ͪ�gAh���@�'+��
q)�_pe�N�$a����' R�ygc��J��%��,J �}��'l��SEI!�@��0�X�:��\{�'l�y� I(:�)�G��9�ڬ��'������=0�p`���,@��'�Y��e^+#! p�S�T5�����'�F�$�.����U�E�)��u��'���(�͓3i��)@Dߋ �FI2�'䬂Pk�KA���[�����'�����D��7&BU����'�Xm7��Nxz��G��*~2T��'F����Iܤ
���7�EzJ���'UP�b�F҈R���(t��z�d���'�d��Ǎ�>v��0bD�>wY���
�'���C�s$$��2ɉ�y�Έ�'ֈ�SbԶ!���zb��DZ<��'��0��Љ9G�x,<JT���'upc�%\�Y�^"Sm�Q �
�'��y+ߦI�Hu�r�øs
 ��'���xc��K}��ّ�Öj��Q�
�'˰����!�np`4/X5~U��'��Ź`L��/2�5��7Vhĳ�'Ϭe�f��}�6 �����|x��'���xB�\�a�Q�ËX�"ف�'͖4�� K�D �B�፲~�R�'݂�P�f"C>�+F�J'�<J�'�9����1C�.0���ӽA^H��'�lH&%�Q��K1�W/���'��I�(
i���g�Vv6��'��5ʃQ�!G!֪NK��S�'8e�%ND�L�S�AɰD�@��
�'N`��ȭ]�����g��q��'&�ىQ*Z,S �ჁQ�7NrQ��'�`�	�6 �1�C�I�>H�D��'�6�I0(jn$�� �� �����'��!�u�Z$@��b�%	�	�$
�'�r�'H��8He5LB�y��'�άҗ��^D�kT��K
�ن�ls���R�Y)^;����m�/�i�ȓl��u�%��}1�x�Fn�%%�(����iAe�Y�L ��LΫ>��ȓt��c�C�/n(��)F�0ϊ��ȓU���L�\.�e !#�B׎8�ȓk��u˓��w�����ؘG�A��D���[���;��(dS`���ȓs֤�w�	0#�d�EO�f� �ȓ>��9CKȽst�$cW���9��]���t'N%M? �K��҈(�n���S�? ����(�1W�>�y�O��
!�iZ�"O����#�*V�^t���x��#�"O����A��@t[�,ʝA�Z��"OxIr�F'~*��:ˀ jA0"O<�� 	ͩcv�3A��"�<�Rr"O�E�fJ[�o�jAT���fή�S�"O4a������9$Ҋz� հ&"O��qΚC��X��Jt�
y�"O`a��_)3��!+"P"O�\���O?V!��DϜ3*���"O�p��	˨��3-��`�.��"O��jdo�4�e;׬���� C"O�I�M#b���Q�5�ॹs"O�����	H�� ��*$o���G"O�5
wa�

<y�\�����"O��:���8!D��Z%�h1��"O�@�W]Mb\9z���A����"O��{䥎����kdH����"O	�A"�2J�VXK0G��|i2�"�"OFI����ÄD�����e�"O���%�΢P��Y�E����a"O&ŸEO-?etUB��Z$8&�e�"O�����$l��|�B��	L�6"O݊�园{h�su �a���*4"O�D���LK�*Щ��	���I{�"O8	I2�
_(A�cD��x�Y�7"Or�R��"qL��Bc�9If<��"O~��b�>��l3���8A+�xjS"O�ᢖ-H9i�^�ñ��2p ,�34"O��jAU�9��� ���q�"OvkY%r=  ���S�>Q C"O� zr����iC�>gO�x�w"O���L@�u��Hyf��8�@h�"Ob=ɤm�)\�8����P#n�(�P�"O$�:P�]"5x��A�ꗤE�21G"O>-���r� Ҋ��\9"O�C���gZ<�� �<4k�"O�L����.X�gԌ4p!��"O@���Q�9A�k2�Sv"O���ȎG�jIz�Ee}�XQ�"OJ��2C�@\���Ƥ({��"O{��$,�f�M״N�0p5"Oplc�'Cw�tY���Jp���Q"O����L�=�F�+д@��̓F"OL(i�.��Z�Ec�Dӽ��]��"O@��fVkz����ď�E�0� D"OIX�a�[ߺ)���/�@�"O!@�T�0V�(4��q���w"O�"��f�j9����Yt��"O.��2Řg^ư����&4��"O����f��M:$˷��$[8,�Q"Oj����E���8�VA��m����p"Of]��6顐��7���)7"Oи8r�ݟYDT�h���O�X!��"O>��S�d�(իsm׉
[�D�%"O�Y��j�?�&���+pY>m��"O���C�,Od���R%��2"O�H�֏ͲgI:Ÿ�ؗ]�Jx��"O���0�=n�v�Z1႖(�Y�"O��s ��7<z���/A+��x"O�M` ���q_�4��/�3"9:��"O�H�K�/h���H��M�u&4��$"O"�HP.��x4�"�C|�pZ�"ڛ$�b��O�	"���%e'<O�0P��6p��I� �ҽ	a�U�%"O� ~��B��q��H�*D�7Z($��"O��J@"*Ta��h�k���2$"O���@�2��I��Y��5�b"O���C��x��ZHI#r��	�"O���2JH�y��a�L���KG"O����#ٱNؘC��=`�x��"O��k>j��H{���]jt|x�"O���HΪP��Y3���7b���"O�����, �n�ʁ�F�oB�Ĉ"O�r�+��^�n��
ݶ="f�� "O�h����(�
Ae�C�Y̌�#"O��;t�#�^�9SM��Q�ze�P"O� ����k�Lr��S�s7@t��"O8uY`�ʽ i��!@���i(,�ʣ"O�p���E�1ب�����!��{d"O�a
��N�4����
��`����"O��R�E%?�X
T�@&�(Z$"O���iT)1���fi� ] |,��"O�d�6k�Ґ��h�#���"O��x�D�m`���I�]`I��"O�ThQE�!6�i����.`��i�"O�����*&�sR@W�8].��u"Om+��ݞm�<	��Ǚ0Tx>���"O%`u��!q�{p�QV�Ri�r"O(x�0*���i���O�2�0�"O�ɇa75�@!�c��̐��"O�lx�.�"a� �lg�5�"O��%4il��R#I&_�5C#"O�0�7�[���`��7G>�L�%"O���� *�+]	XR];g"O��1p�0Bu�U�i��k�"O�y+bEK��ip�NN�m��"O��P���_���6Cɉ*в�"O���q�� �8�ա�h���"O��Cށ �\P��O,~��2�"O�}YFo����0�0�HQ�"O~1��4h ������,���i�<i�+V�da"t��B*� ��Vd�<Q��� ��Y����t���H�<Ag�T=o���K�+�&�C��G�<!���,?�ʢ�ީ|�$)�J�_�<aĊ�1���r�)F+:��b�P[�<a�f͢h*�Y�
U�^�����S�<	b�I6u~ �+§%�F���d�S�<fG�*H4(����<>ҝ��G�m�<I�j̐ow8���L�)��XE�^�<���;:ީ3�(��
�J����S�<1D�N7N��V,�2"b ��]s�<1B+]8Pp�/�ub��i��w�<�bC��AK��!���j�E���Sz�<�r�SN��8��ɝ�htd��A�y�<��	*Ks�Y���� 
���\K�<�QM�\/.���&n� �_J�<�r�D�}XbM�3��WX�ԑ��AP�<�6d�(\+dp	������ N�`�<��)�.w��0A����Q�M��< ��bŲ��W0m��I�cw�<��d�8���Cg�&@
]��̇p�<��$�;�L�� !� x�F�U�<���7f�6����� 9����f�YS�<iE	��"`�ӳ,����
�H�<�phG�W�VB� �1N��s�@�B�<o�=[ݸO=Ԙ�b���Y�<#�FE|����M�<2Utu@��Y�<� B���"J-r��fGQ/7�qR"O� !�J<��� ����[�j8""O �%��+���e�W"x��`�T"O�����	z�Tۦ��U�����"O4��dH�/c�4��"Ӹ1�BH�5"O��C�'Ů\��cb�\]Ψ�t"O���q���i/F�K��Ϻ~aN�X�"O6��u+�5Qz�8�a��HAR��"OD%pa�0t����b��ZD�I�"O�pb��;OV��"H�"֬�"O<APu��&dQ�}^��A"OT:ŎIv�I4�Q8iَ���"O�@X��ޔ�^����A��=��"O(ٚ�.J��^E��G�6|V�!V"O�����:?S.����^D��D1�"O$mS�jK �y�H2yR�("O�Da�E�s�N!��� G���T"O���7&�tAjg�6M�j"�"OV�;&f��,�z�C��VP �"O��#S����'F a�ա6"O�=3g��W���ƒ�FJʍc�"O�5�3�"+����0�R9�*�Pb"O@��'��8.B����*L�I�"O ���(�&
Б�.�U��]`�"O&i!��l�r5�k8m=FѻU"O^P��֕`�Phw*�"ԂAC"O<�Ygl�'J"� �P�=7�))�"O��G-�Z_���D�W7G!,�y'"OVI5�ܷS�t!��H#h����"O�A(��\?�
����(�tZ"O�X�f�!vk.�##�� Mx���"OD�Th�YQ ���(�9?~�}��"O&@��ȇW�M�b�� �j� b"O`;艵-u dђ�Cf��@�"O�x���.x��`�LG���E�""O�p�G�J�!�%@ᖚĆ٩6"O&� ��)-_!��@��-�҅�B�'ѨM "I��>�3҃�)'�� #�盳�jC�	�:�= ��'�p$��N�H#>�UKדG�x=����.N�Y�#%䕥/�8���+�y"bA6=�Y���X�y�tl��Mˢ�p+ґQÀ���s�$٨%G�n����9&��ku"Op���D��<��F1x���p�R� �3��\������c8��	"b	3LEFE��V=(�x	w�#�O�@C��[�+���̖+5@��׬�z
�y I$^l�P�	4�O��a�$<�	��g�q�Y�p��+�n��ǄY\�6	D	�@��<��M�R��������7&C�	�Y�n9�\�E�tdS&��7�$ ��䆓Q��tY�GW%r�|A�N2�g?�V�щJL<�!�섔)ڨ���U�<1�k�aF��sCN�Gi����%NC>6pb�Iw���{�N��	���3�"0�ea�kAd�Dd� \�l��,b���[�-�`�ɖL�C,*��]�b5�剈IT=3���B��l���7h�����A�_�ty�4('�	^$ȵ�ƣN\������/DI~����p(0�0 ��L�'��E�Q	7"O\4�  ɼe���#d�<{hnqQ�U�L���iUn}�6ͱ��1�>��3���D�F�(��IH�	�SJ4m�ȓO�ҙ��F.g��룭�{�&��P&��oh`�p����~Z�`�aRݺK��6=�R���R��"%� -�3Xa{R�J�D����d,�l`dg�R����_؀I�A��V�j�'8�p���*]��e�&�F�J�}��Y�Q4R���ENh��u
�)c��'<T�y fZ >i��?_��8��4D�����K�W	nj�Aނ$�P���>=߸%{��ƀv��,J&Şq뀣}��Y�T�R��Ⱦk�Q�׌�&`�Y�ȓg���� �jP�x��}xC �~hG�
��ɓ��Q�� ,�'������dB"J�ܕ���'�X2�G�4)��,	�-%�|R����LH����r����CM"le00h�)o��C�>�{��%�bI@&C&�$?��g�'yJ���ҁ$��("�$1D��c7�Ϝj���S��3m���5Ű�T��HT�R��h�L<E��/Gh�'%���F8Se�J�y�JK�$I��8�O
�}�l��gNV���4\{��Raǌ��p<E�@�q#գB��
��f��q��1��"�b��E�B?z�H�3�c��{G�XOh<�#��;VD&��p
��7���y�'�ް 6�Ӳsɘ�ȕlu����#�C�I�����S�_��9ծ�=_��C�I'6Ԓ��d�F�D����u#�C䉽wJ�]�G޸��&n�*t<B�	�J驢�C�yN�eh�c�B�ɠm�i2�ϗ�Y�*�3��$C�I*ZV�� "۪�.�`�N�a{`B�.V����Y�A aK���2�RB�I�=�@��܆/k��a�LV(RB��v�a�dǋSwjЪ�	��B�I�E~��ZkDa���q��R� (�B䉧���[0���3�̸�D�^$P�|C�I"B1�m8��0��-��.��~C|C�	6��(%��tP�F��7m�B�Ɋ�fĂ�/�:������q�`B�ɕ��S/�_�P��良(|C䉼<�d��#�5$���aċ�>�hC�	� �J��É�=(���	�.�{��C�
1��B�$L�\�@�ևOA�B���J�zQ��j�\��f�.��B���N�{��.	Ud�RB��ZC�)_D9S H�?Y2�
�-ϼQr�C�ɒ��,Cg!�#'5�w�Y
-!�B�'x�x�cŊk���!�R!+�NB�ɂ?�D�X�`Kz�`Ժ��_aC�I�e\�2*�3ZW4�q����0��C�	8ɼ����(:L�y�ē�0��C�I$dTe��a�C~q��V9idB�I5[���c�7��(�}A�C�I(0�@u���%)������O�6��C�I�)ʶ�)��ݙA�]�w���7`�C䉚f�tY�B%�'lے��č�70�B�24_����,��/�TS��A5W�B�I�=gr��� �!j�<��Όz�B䉖E�h��ȁ/�JPD��rC�I���y{��A�KW�ׁ	�>C�4S��@k����Q�T���K{
C䉝mX��C��>!\�c���h�C�	zS�L�d�K$�(y5o��
D8C�I�[�����+N*��X� ��+�C�I(x`�L[!��
L�y�iJ���C�I�#���٦J� �lU!'"�-M�fB��O�L�G�%2V���'�'b�DB��%@r�(r� ��M2Q��
-�B�I�tܤ����6H�3	
�.M@B�I6 BH��M��YڑS��֏'TC�ɁO�lm�֭Sfj�I�%��e��B��
w��D�`�:|1��B�WR�B��9x��`$�\��& ��"JdC�ɍ9�إ3�*Cp ��D#G[�(C��v�nYy�EIZ�� ��o�,B�	12�@�ƪ�yv����(�bP�C�I�l����9���ڔҼG��C�I?=i�p��j/�L+D��*'��C�)� ��1�ݫ6g�%� ��̖��"O���VMB�A�H�{F�_=Z�*��"O>a��Ā[�3��áS��Z�X<��w��!C9�;�M3<Oz(�q��0�(�biF�<p�"O8ĺ��G�V�P���,�,DȢ"O�͒��D5h�بKRe�xi�R"O�L�R��[�P2��S	�y��
�ju�6�*G;�xB���y2��Iᖕ:�"9�#��yre�<;D����z��]�!-@9�y�N�u����b��m�!␱�yrG�*7ӎ8P�E��a�(8�S2�y!�2��bV%+ �H��,�yBg
�`���Y�(T*�>��/���y���Q��A�I�#*f�ff��yMC;t���0��D���YH���y�-E�
ՠ�]�u�l�%��yB,(ܮpꄎ��r�N]
���y�%�w�DeR��s*�����y��!u	�Ճ�kjPYF�@�y���'���r�ݬ}�~!	��y�l@�=���9@��v��}b����yb���\5�u���:���8Rb��y"���X<�# Ժ5Ꞁ���yR���#,�xp
Ԃ�Y{p=�y���.^*0�*T"R8�v'V��y��ز�d���Á�'���*墄��y�ŁEڌ��C��0�}(�+���y�	X�~lr�m	��9�qՆЖ�y��^~Tv4��+@@o�,iŬ4�y"��Z�Ř���$���t�.�y⩇� �����g+���D&�	�y"GҬ=��E��X;K��Y1��)�yB�8t���ڃz�H�� ձ�y�.��7:N��f��X~�j�OI��y�e�(rD�}[@bG((Ԏ5hBl��yң�p�c&O�
Twj�uCL��yB#.5Q�Q�޴S��D%^9�y��K�e�P�eA��".8dᔦ���y2�XA�����	@P�ħ���y��Z�}�������r
� �yrk4s_F���(��n�t��G��y�g�4��1U���*��t,V��y®]�D;�C� 0�Y���۝�yҤ_�m���@F!s��Hs�Y��y�N+6j|qT�����*c�À�yBe�v=���0��a$��)b���y�VP���ؑ��3]�t Ґ�W
�yeK(;L�Y��KN�,<���ޕ�yB��N���EJ�ur`)`OT��ybi@��x�����hF\��WGA(�yB��/����Ma7fE��yBiSd��9��	�>FD�f
��y�j�Јk�Ă�/l.�I�c�(�y�瀇 nl��FF�.��x�0��>�yr���{ݚ�ӆ
�rADa!�ʂ��y��C�f��4��lS�!���
GCP��y���&'��T�a��9���&AA/�y����Z@	��D@O���$%Y��y� t|T1A�錴4��pc`F��y�������B�,1�xZf̀��y�O	�M�(˃FV!&�`�����y�k&;VFlX�� +$x(�C��y�(G�lp��I�$7���reZ��y
� �HDㅵD)@��gEKya����"O,)�JP�t�*Y���HM6 �J�"Oҵ �ŀ�yI����&�j<t��"O�y�P$#z��8cHΊ�e~�<i�kܗ6	Hhz�˗�~�\� խ�u�<�eo� I�(�Tٹ~D.���n�<�F��$]�Es�\�A�Q�v�<�!�*w` ��ɲT�n(aѣu�<��F0?y�x���)&X  ��i�<	uh�G�Ԥ*���.<J��rm�f�<qP�ӸS�* f��->���0��{�<�.�?o�����;o���P�a�<�̏%up�<qS�Z1��a!�^_�<�S��J�(+%#N�Ȝ1��!^�<y�Dʤ��U��?e%(T��N�E�<YP��9&��s��##�[F�<BeH�[<N̛� �&ـ��1��m�<�r��~ �(��+�!`M0Lh��_u�<y5HI�hz<�f��N�tE�3EMp�<Ѣ��$|M�eB0k
4�$�COAB�<QR^?j��pJ@�Er��i[sO{�<i��Si:��c�B
?��|���u�<	7b�8|�p�FR-fC����gIm�<!c�I�U�Fȸ�*�+�t�8ALO�<��	4^|E�m�3�Ȕ�E�<� Ȇ�l^�[�Gt_^�`�-�k�<IG�"<^ܸ�C�^��Y�N�N�<B̵5nL�[T���ZAf�k�� G�<�w���#�b��A`�6�����'�@�<�c]-^D$0�N�BX�A� /�d�<��̂l72�ie@C�(¦(-Yq�B�	��Hs��ٴw�P��/�B�	b(40G�ƞA)d(K �:8)�C�I�W�
��C:�A���u�%D��	0�!Q:, ��l !�A�-D�
rG���,�����,�&��1#0D��	���v��SR�87O�84d/D��0v.��9r� p��.���c-D� �&9b�E�&D��]b $,D������%{!D ���[�8I�%�$D���w�>X1j��!#S@Q�m$D��"p`^���(;l��4�g$D�D{0\	�y�'�6-2�"&I#D�4���W&f��3�dy[���ed D�@k���*`�}Zv&Գ2����`!D��c�i�Q�'�"vLƐr�K>D��A��1�Fa�ЉaĦh$�:D�L���L"
lW�i�����7D�����D`9�k��
Uk�`J�7D���P�jt���j���ڇ*D�������;�лR�	 {$j�� �#D����Q�m8����Y=��b�%D�sRM>sT��q��$S��X�ӭ!D�xpb.��	��x1b7,�D)AP>D�X0f��#���"�E<)8���a"D��K#�Z�U.Z�hF�7.��̀��,D�0�a�)P&d���B� �ĵj��*D��PG�EB�`ٰ��$U��-�V�=D��Ӕ-A�x��"�����p�??����ӠD�09BV��"kȱ���"C,$C䉮:����p(E
b��P��(:x��C�	�*��r��Sά�a��T�
�fB�7v�����x@�(��	�TB�I�5�,1^�t��D�J��U�2B�)� �X�j�[���%�%]��Q"O�"�H�<E����ߠ3�*E9�"O��z���}W�`:G�3_�V���"O���.؏F]8}�1c��	�`y�"OZ�X�HW=b(��5��i��"O�)��
�x�p ���06�tS�"O:���+��0j ��+h*b�c "OƔ��昒PqDac�.?)V�0�"O�+ ��	bir(p$�
/|��س"O>�9v�L;&f|��2���h3�"O"��� �ce��顭�H1�� 7"O� gf�(�\	���> �b"O>aA��Ez�X��(eM� "O��2�B$))�H����;N�ʵ�"O��B2-ӴM�F��MY,�}3�"O���I�S�䘀CƏ ��H#"O�M�TgL�_�BqrWO5w�v-q�"O�M�5F�)b<	aHK�N�.��"O��� >9�lh3��w����"OZ�a!O$-�hH'�1#�� �r"Or�c6��0�l%xU��h���"O�Uhe��+$2�!dh��Êq��"O�����2I"p���L&gH�yE"O��2��@:D�|=[`W�Z>6�k�"O8�+�*W �����%,N�i�"OB̊��j��J4
_:pl� ��"Oh�� �N/Z�~�2�ȼp;����"O$-� ���^�rň]."�� ""O��Ps͓�w]�i�`�S�"�(Xs"O���"nQ���D�(_�2��c"O|2E�D3zd���4"ɸUkG"O,��b&�6[�%[��WAP* ��"OX1���E���Մ�4�P�G"O���a-$�n���՟xe��"O�M���..��m���R�E�`���"O,(�BE�p@ ���ךP5l��"O|e� A������ ǜ4&*�{t"O�13�E� @������"OL��7��70. �ɡ�0S�A"O"��֒x(؀���H���6"O�h��ضnvL)Bf�2�g"O�H��bL2j�a#���$b��"O����S!*���㖗9p$�!2"OB9K6�I�4_4m���͗O
�i3�"OlmcQ��!ZB���Q�9�8X��"O(����NV�5�O�tb,`0"O���JV#s6��P=�t�F"O��c�����Iq�,LM3P��s"O�1�j�=��aa�KLG�R�"O��S��*?"|i��j6~Q3%"Oڀ�q�=U�L��E����"O�pР� >��4�)�f��"O�@z���=%�8��G�)c`�9r"OР�׬�$|��q�(E�����"OƜ�a�,C�2Ykd��$J�"OC�ê{Ԟ$��5 Ξ(��"O���_>N@������ +�pq"ONi3	�#Q��� e�%�,��"O�A��r(J�gD0��e��"O�����ڢ!�����G�f�N��%"O8�jw�:&,�C�;9��4;a"OJ�@�
�>NE��2B;t" p"O�E��bȇP~�= \(+�([f"O�����S[-��;��" �1e"O� @�adjC Fr�]�h�(Ȳ�g"O��bj�t�V����ȔRa����"O ]*ч�9
���	q�&e2��s"O��ے(����˴�)har�s"O@M����Z�z��t_�{2��e"O����F�2x�p����0f��.�yBEZ([��$;6�Af������y�fӄM�aX#Ŏ2��b�>�y£��ZE��0-�,�Qc�=�y�ͽ �Y W#���EmB�yRIW"��IKpHY=f��Hce���y⥓<z�����)�v��ŀ�H��y���O�>��5bD*_�`���b̚�y�EY#2�b�+�V��a�F�yB��:h1� �%��Z:< ��+�y���*aj�OGb��b�.���y�	��9.� Foٸk���#O���yr�D3+�D�#�:k/��&�0�y��L�nM�mQ�c�7Zd� �B��y2��+-�^L��D9
[�!p�]��yrG�B}�f!�����7 �y�� Y>�Y��v��R�a���y$y6Ċ�'N?;qZ������yb�]sx g`&��)i���y��X�FfH���ab�83�B,�y�CB&1�܀n��A���A"���y⍟�$$�t���� J6h��9�y򫐍l��K�NUoI�M��[�y��55V�p҇_g�L��B�6�y���_�x\��_�>E�A��y�b�VI.�b'�9$}�T�@MR��y�'�qL] ��)�4T i��y��pEn�Z����Z����N/�y�ԇ>�����I��J�;��!�y�Y�BN����%��=�����yrh˄P����U�.O�<hV���y˅J1��*��-Lbzxc �F �y�.}�L媄�?B�6�z���y�-� /Ո�*U�):\���aOO��y�F���MBԅ�,cl�a���y���"�x�D�μyff��0K*�y��O��"ū�C�);���6�yrbжaR�c@͞#�����X*�y""ۚhFmz4�Q�<`��^��y�tA��
ab�PQ��@Ӷ�y�o�!��4c�Ȗ@��)рM+�y��
{!68��),1�VA`NJ��y���<���K�M�.@(!����yr�S�=�EC�N�5;x�q��ߊ�y�$O�\�tp 2��33�x��2/�,�yb�_�;.�����f��C�̙�yb�^y����#�9ք�
daR��y.J$n������R���D,�y���<"�`N��ypT���Ґ�y¨�7������vF~@�"��y���)��{aC��strEARlť�y�܉3'41"���{�t�*�!�,�y�Ɛ�-�$���EՉ~��q�·�y@I2���k@��8=Z��U=�y��&&�(0P")�'Q����7� �y�7ƪQ�#��8��*w��yb΀56g@��f,��<��/���y"�
�C�q��%�&�j%L���y�% �5�BD��@�!�����G�y
� `�hT�E	��t�٧@l�0�0"Ox�L�s�2�˶F�
R���"O�Q��ƺ-X�8(c�I��.�j"O���
'NYvl�gd�� �~��P"OXer�E��lZ�1T3S�t]��"O�1
�OP5zT\(�"X�Lj��(b"O�h�\
*�0�i�Y�k�<,�7"OxT��j
�(�10�c�Y��	�"O�US� ���N4�"��& yW"O��HFVsnJ�Z���U��hӇ"O�2�iSRӴ�:����*�"O���"9��X6�>шL��"O�]�'��Dz5P���1lȾ)�@"O�,�Tʖ  �Q���R��l�"O�ԡ�J�y�q�&��bD޸hC"O�aV)�Q�d�byC�d�d"Orи�HcJ�م�<K��4"O�	 �ܕs{ވn��M��$@vL3D��R�A�(q��2����Q]XY��3D�Ȩ�NՅ,���:���@�`�)�6D�X󢈖'4�����!Ǥx:Ra��"D��$*��Ǥ���D?(
�� ��3D���A��~)�2� ��\��4D���eNǂ�Xƪ�,B�|)�0�4D�� !��QP,��Q�_��Fm+2b2D�$�L��Q���1�ʒT�����2D�X��:6�N�kP)���v1D�X��L�&K�L	��<1b©
�H-D�|;���z(2����)F�r���i.D�l�$�H&��(�B!��m{:e 1�0D���^/T��)Y�	�g�f�Kf@/D�`i1�Bn5໔d��^7T�K&+D�@����$�(��EiT�viHըQ�)D�d��%S�@��*�@�7~���.+D���@�/j��,�a��6c��Y2�,)D���%dS�II��%��''��ba�9D�؃2g�
S>��K��N�\4��L;D����3�"��N�=Pj�+��5D�� �
K���2b�H�o�4���/D��C!s���!�[�RD.m�'o-D�p�#� R}�y	҅T�E�2M�G7D���2'�\�nA�����Uk$%�5D�p�BB�|�Hi�R#V�%w�!@g�1D��9Ӥ^�;�J�p��R����;�	#D� �Մ(�\�������j�	Ũ3D��
 b PŎ=�g� g�hɊ��1D�`���Ș$�s⟚���
b�*��䈟��JЁU��HbS�؟*7
��1"On��s�A�[�X��M�
 O>(�"Ofy� ���%����l�48�\�b"O(�����0� ��?=V��"O��Q&K�4h�ci�#��r"Oxa��
j��0����/��Q"O i�$���Mz�t�`т"ODՀl}L�i0DCS$�Љ�"O�lJ�-��kw������jjp�C�"O^Bug<�}J���H~�A�'�г`��b����(�J�!�'\�;f'$&��H b�U�~Ux
�'��pd���q�ds�� Y���
�'�f�9���V\���V\(����'�|���Z�W�d�9��=��t:�'-~�{�M�7����`��9��	�'C�٧k �8�hHSnA"������ >%���kЈ� ��&QF��C"Oy"WᗥH�(�I���ODl�"OP�(�m����'S3��ZW"Op�� N�+^5�m�zy&%�"O��T��LB����b�xa��"O�8��$����`�ukM  �±ɦ"O�����J�(J�S����G���Kg"O�����Z����)W/L��F"O�ceNK�F��Uy�Ĝ4�xA�"O.�S��H01�H�;p��0�����"O��r!���\�ǏV>b�V=�3"O�њ�G?z"@��ߞP;b\�w"O0Q#��7K���q�P,�\�R"Oz9���$jVLI�%@ N��pq�"O�����X3�]9f��3����"O
d+"�A)��t+���M�p��"O�'c�3Gȳ ��39�n�J "O�����'_��WaH(F� ;�"O�܈�䅫�Ĝ�Ŝ%1�*�:�"O���i�R��%�,x�@�`�"O*X�7�5!q����R�4��<""OPIkF�`�����J�*arT�"O�)�cK [5�A*��8P`R��"O$	���B`�~H�3I�.j�51a"O��sꎉ2��=�egƕ" ��5"O���cl�%1sԘ#D�k�9�#D���aר-ִS�A8_���m!D�Ԉf��Q�R�9���.T��B�3D���b���v����΢"Tn��3�$D��+�H����3O�qu@u��6D�XZ�$� A�}9�b=i�Դ"5j3D�$��퓊�j��DM�]�Ę��@1D����$F�S9�H�o�\Ia�#D�D)bi�>�t�Q�Xkڸ��#D�\Cu��9��L
D��u�d�� 4D��Pr�.Kl��'�m�h�"g�?D�8����,��`��C1�"Q�� >D�����ʥ�xѳ ��`�60���9D���H
8�Z-[F'��mV4k
6D��xv!Ή@u�R ��K(2�kօ7D���R��@��T�$,�h#����3D���cHF�Y"��ğ�*�|�`��$D�(�(�S'ک�*қl�z9@��.D��6DD�t���F�.�${7D����۟]��L�#;e<L���5D�h97*���|3����6*��VH�d�<0TQ�f�آǒ�MMҨZ�H�{�<��χ� �8�1��6������P�<Q�!�%m��� MI Fu�- 6ɀa�<�b�)^��:v�\>j 2(�1)�H�<���ٹ6V��1�i6u�A�@)LY�<��)�#�v�����!j�]��%AO�<��� @�ԓ�͔<��{A+Kp�<�Sb� �"-�K�~��l�<��H:y:�Y+�3_�l���l�<ѳ��b ZQ �������Юq�<�׆��:bR Q4�͠lR��n�<���� }@���H#^ �U�Ѕs�<�ѭ�~M�1C��d:D�<5��n���*eͤ0�~ 3�K�B�<�� ��h+�IS�Ō IH]�.�}�<�G5 �,Т�ɂu,aS1a��<A\5 �E�R>q����/r�<ad>5rIP#�ϐ�G��qʣ"O� f8RL�� ��/B�v����"O�}��l]�Q�Xa����s�AV"O��r�#j��)��cM* �
�9�"O2u�0Ȅ;��B�BH	i5"O���cE�/*� Z���ne�"OD��T�ϗ)�6��� \�/��X��"O8a��Q�qT�t��H}|T�c�"O�E�n�z�*�DO/=G�B�"O\]�D�N�#r�����9\�1a"Ob�s�хt��iPƃ�/��۳"O�г�(��UF�X�Ϟ]�MJ�j�Ot�Ce퓉�M˫O?�	!�	HVʬjB�UF�6���EԘR���k�'D>f��R���bB�>����d�w�S��d�� �U.(Mʣ�i�dd��Џ�t��J�IYv��3�D� �@]��*��s�A+��N�ȑW�'~�]�ig�����'d�u�2��-��)�`��N��5Pՠ��HT;c�����쟘�퉖�J�C$���V��s�\_f�<ᕹi7�1��ɺvk^�c�rAH!TY�ģ^a�2�'m@Z���L2�'���'+DםΟ,o�+͚H[9��i�u� %�V�$� �v<��Zi>�Q���}��	�o�Hi�v�|ri
�a4^�k%' P��S�G�|3E#K4QpDba%٘�s��h1���<#�Q��k��$��.��@�F�J���!�(\��?��o��?��i ,����� �
9.��
+tNX����8e2z<��F�0��%gSL̼�N�9���a��u�|�o�S���?���sy2�U�B� �p2J�r��u�BS��v��H�'��y�'��=����^]�!��Аs��`��F�]~<���@�T�E~� �hR`�P/3 PĚ��Mc$$j`�<�>�#�k��y��tn~�ڤFS�NOz�ڤ�'��p)���]���m��_oa�����>6��O�� ����DB@Ϗ�!���e�H]��E~�<	uY�x�Xt0d� �3�|}���w?���i�66͵<�4튠7���'�"R?]�� Ť'.� �!y���� �%U6�M
��?��� aX�s&e�=k� ��=Y�Fx��}�%�2�<��K;(�d9��դwQ�H�F�"c`���l�"��������O6p8�^�j�CD��ϒ&���&\Z�cFiP�@�����
K}�j��?Iиi<����67M�8%"4�� [%ZMa`l�\w���	J�S��?A$Ȯw� ���<�"��΋W8�,��4�?ڴ7C&L��G�Ag ��}j8���~����i-R�'z�� 78��	ן�lZ�� �C�R]��ߌ�X4p�+���̌�#�U4�(MpC��,�ФC�l����'�zYc�����.�""(Q�s�0�P�Q�4ZmZC̾1U���gY^i���!17�P�Aʭ��Ƽ �U�V�4J�1εI�p�r��i�h�z��?	ոi�b�~:L|n�[���s���2s Dt2�C���I�G{"���K��×�Bjyz�d�@�Q� ��4��f�'7M�O� �g�|ݡ�W�H7U��L!�ݼ\  �T���?��КIR�� �?���?�	T�N�O�6�N���NC~��U�V ������%61>��� �m���b�L�?���C�|c��OJ��a�U]5PpӀ�F�ZZ�R��[զecHo*큒k �T�v�t\������fmZhS�' *ܨ�ϗ��`�:׍^�9�*�I��OT���O8nZ�-���<q������z�$$`�
��1�����%ò����iA`u!�	T-a�4RT�EYf��m�Ӧ99ݴ�䓹�	)�	�nOҖ  �   X   Ĵ���	��Z��wIJ(ʜ�cd�<��k٥���qe�H�4��6_2<<�3�ʄmn�.(��f̅3V��(�87�ݦ�+�4>��$<��uyB ��<�Ty���Ѥ������G�9S0��4|�0�=���%�1D7�Q\�:I�Ň��<�c�p��	��v]XT�ʂ��I>�.P�łN�:(���&a��֢s�LYʵ���^!�c�J��-��(Pl}2.�#<$Tz1>����%�ε:@cA�	�j�F�.Ar$� �w��I�yr�C�0A@喧�$�Z�"�PsW�I�}��7|
H���"8<Sþ�P�`eaea�
�˓9� ��nQ�}��Tkp��������9���y�d#<Q!)W*��)E0a���AO �d@YP�I3(���h�Z��Y7j<C���Ci8,|�)h�E&}r{�'.��=1UI�jR�IJ�!v�V�"2��ʦ݊�ቮ[N�dхĉ� �����I4]q��P��8
$b�TS�I�j��I�5�A� ��܅0�cL�*��� |�#<�`0�	�O�TaAFS���bK�#���t�Ɉ`�X��'�bh	w�N�[�:}X�G��>(ybHJW�'��&�t1�f՗,�<�1�� <dXm�������	(S'�'�����h��OB l,����b���xy��Z@?!�l]?��	��� \w��H�A�
h��'i w�)����;�O���H��b#��KF���Q�6�tD͢>�� �4�"<���5D�ThF�H�_2���A�<)@�� 2  ����C���q�.D�l�#�8d�l���R�{�LC�i,D�� N�{L�;@�°�Y�XAs"OT�j��R,������.�I٢"O�l�A�D-
5��2�NΒ"6��Y�"O��+�ƙ|�@=�t͋�
��?�yb�����x�,48� ̛����y�D�v��s���g�J�;��4�yB�Ƚ#8�a� L�`�ĕ���L!�$�"G"~D�ԩ��S4���«_�!��m�e;��S5��4�ӭܮd#!�deB�гP�ߋ	����U��6&�!��]��,=:�f��[�~]��mT�t!�dC=2݋�N�'�e"rbׇ|�!�����s�*07�d��Xu�!��_6:\��3Ҫ�7".�t	CDܐ5^!�DZaj�BVU#�4h�U�X�4m!�D�(>}.|[Ӡ��id�#�N?    �  *  �  �  ?"  �(  �*   Ĵ���	����Zv)Cll\�0R�P��
O�z��1Qv�i%��/��Qlр�yb��Z���Jc��?��J��ߪs������I�<7|�������ݚ�-͛J��j2@Q66�X
�ڠo��	�����N�9 J:��� �:OC��j3iZ�5���c��&h�St��� �����O.:���3�0S{����ځ8����$��A{�A�/� _�D�H�&�&3�@U�u�<�Iߟ��IڟT����$XM�@
i1��		sf-c��gy�AM�$����'
R�bt��^H���S$FlY�I7|��tŎ"d�$I"�擽���	�p���Հ���1!��K��Ξ��@	�\�M���'!��ٓ�'yB7me�,O������b�&�vY&�#1�ˆ@P��r�3D������H�֡Y�!�spAP�fl��!Dz2�H��V���bF� {��ɅcL	�b��)MdU��!�П���؟��	�u��'i"0�阁�'Hre�����'��l�.&{_r���$�O�����OD`���xl �,��dw�Kax�x;w(�O�����D��Re@\q�j\��QR�<�c�,�[r�5��%kg�x�<a7I�,&�6����"9F��f��J}B�{Ӳ�O��c ��'L	0(�a@աNvH�a5�i�j�Z���-q���F/v�:�r
�'܀@�s�іt���P����'�� ����2'�
0K H$����
�'3�tۇcM�=ņ�Jc-�!D9$�
�'��c��ƚEۘ���� p��'X<�g�+vc|�"�NNt�����'5n#�GMb�zh�c;-v���'�$�[�Ki�� `���a댼��'��Qu�	�6��	K�⁑;���'��y���0��£LD��)�	�'H���v.ɿl�XH�ɕ��P��	�'�L����I�c3���ՉA�1R�]B	�'��A11�%���A�#�h�'��$�ǚI��kL�X�Td��'��PA�	�p�a��Tj.�3�'WX`	eM3sV��� �9OQ��	�'����A�$C��$	c \�@\���'kn�
�ޠ0�ȉ��㝞���y�Ϗ�d`�W��[k.�����y�b�;!��`�&��i)��s 	*�y©H���ƯP��eQ�fZ��yrm�qNĜ1u���9�]0X��y�m��^�rP+���6"<�b���y��M�3n��7/Bz1t]��J��y2���xy�w�5l�^����O��y"m�%pQ2=둡�r�գ�f��yr�<	D�[�J�9e���5g\��y�O�� ��!���@
�	x�L��y��X�����N^�
�����;�y�Ȝ�U�5�g!��s�&$!�˔�y�R>H���c��{J��)��yR�!gh�a�d��yCO��y��N�K�
�q�gKЀ����yҏ�B"�4Ip��F Jȗ$�y��C48`����� >?�-h!ŀ�y���l�Vm�voT,4dx�C&���y��ME
5@�bO<@pܙQ�
�8�y�� Ű�����M�|�r��=�yB.ʑ\�P�j%nߩ��Y�_�y��V9� (Q��Wy週�VM��y���5B�lj����t	�q%!��y�kӎBQ�"a�!Znv�;�b���y��A�^� ��`���)�%"c̙�y�/"צ!��[����O#�y���4"<�U2�#��PϺx��e�=�y�$�(̥1�&�8V
��D��y¨�,(m)�H� R��T�Z��yr�1�v�xp��$O���G���y
� �(��d�$�%1���2Z�&��"O�e��O�?$�1�X�&0��"O�L! �/+���c���9,>��ٵ"Oܹc�#_0�\`���?!$l��"O(%�ԋY]L�p8�㗍+�2�1�"O�h��wKD�{#��4�c"O$u�R�$�@��R<�ƕi�"O�d��͞2���I��tv���"OF���E�t(<I5��\a"4[�"Oh�YR�]!t�5f��^��Њ�"O�S�նuF�B����Vh�"O�)Cn�:L��9R���
��h�"O�d٢��.�����_��
�"O�h�5�}�&�M�c
����ݍ_+!��!F�&};�����hh�G�!�!��_�p��7�(���[O�!����l��X�v��(��$լx�!�䃀]�� �9?Sx��U%�-{�!�.,m�����G�iך�J��0�!�D�D�ް���
>�(�EĐH�!�DA+�2l��Ϛ�*����SY!��:dzE�DFEl^X�5�	&0!�d\��^�'�A�i�0�)B!�$�<yhD=;�՞n^f@��&��e!��[�
#b�wBX ;�E��D~!��оn� [R΃2F�Ɲ�p��{o!�$�!��a��9D�ire��Ux!�$׼u�T��f޷;��91��2q!�dįEn�hD�H�|��9�2f�*:�!��B~�͓�Aί�0EP��!��]�\�W�̲2}x(UJ�b�!�Ĉ w7ލ���Q��TY!!�$J0�= D��{,����Xq!��� Ak�jg��[F*�"�$�n!�$�:}��cm�*`�L��b�6Q!�$ľ#|����,��<���-�!�R�F'z�¢�@"-�TA��!�61�!��L<���c��	�*N�G��7!�dt*�i��ʂ�~��� �_)!���K�2�[5��@l��&��QF!���b�2	��c�?�T]@���F�!��3����79�:�Δ$�!�d�(*.�S��i�(��+I�F�!���TXh�#5�L�du�i�W�[�/�!�ږ	�f5ȑ̕?k��ȗ)�7'�!�$�2 X��̗ׄv/�����
!���(��:!�<4+��7��gq!�ϫ.��,@�C�<y|�Q�#H�/N!��ʝ7G�)a^pd��� $BK!�ėl��nBP4)dD�P�b�;t"O�tٖl̛zВyq$+�� o����"O�����v�P�	HS����Q"O<�V��u���鍉q��qʃ"O�Z�k�~5�w�#s�x�xs"O�9��Ss�]Ru�R�/ؤ�[#"ϱS��OD�}�o����	���2�:v"O3&N��TV��.q�E�."|u�v��Tֆ�0�%��a}�ݼ)�1r�Θ�E����4����<q�ƈ�'���0���yrPF��#Q��Cn�P���y�����ӏ��.�
�5).�R�'��1!R$R��\��D��˘(>#>�1��V�J���r5b���y�Q�dņ8�K�%F���u��&��HRd�.0���@�G�h��L>�w$�+g�茢�ɔ"�HSgO(<9���dC��
qS:�)rl�U < K2���PG0t�թ��=� �<2����d!��\�<�!��'� ��t-�w�v��	�E�I��N�]���0AN.��!\W��B䉕^l�r2�5I��p@�+�!
:z�*\�dG��t��փ݂Φ�|��C]��y�+C�'w��� �F�<��!2D�rG�D$V�4����.h�,&K
7JEb�Ah��i'?E�<ِ� �Dt١��
�4����u��Xٔ�!r���fWIVL���*2��%OH�z�v$�`�ԝ�p���	�-j�� Vc� +��J�`ˢ�?!f
H�}���!�"Ѣm^YZ�k�:bZ ��fX������a�1(tn���'=�d�g��_����% M�1�Tr(O~�懇�t�6�ZV�Q�w����'§.q��ر�w#&L��E_N�D��.�5j2�O6v�a���>q��y�&�K�f��ch6?��g�g�y�G�N�à"ɯ��<��XxnԄ�I-gN�Ѷ��1Gb�g"E��Ycv�-��q �� 1�R��`�U���C�-*4�J�;Nv^�{�8O�i�T�Y��p��"�3WE�芥��	C�N���O�0`��䀧�[\<!�D� 2&�F*>$� %#rA�?1�I�~rQ��	 WiR��(�X����D��I �d��"OP��v��)pQ��	Z�Z��ۅ	E;,�X���
e�#�g?�ǄH	Ȟ�)��O?v)h\�Q��{�<с�� L��@���4A�X)��Φ=D�Y�[(�ԑ"�+lO�8#M��u�L���E C���u�'r\��h��1:�	�v�S�{�XB0#��`��C�V_�P��	_�xH�3-�*Rvb�L	����]�X|��I�>k�T�Gd�L�B'��4 �!�$Y�~V�	(Y0/J���A�����c��P�I�F.Q>˓�RMbՆ�;$_8:��ٹPW:��ȓ�r 
��2N�zI��K�����	�p@N,����S��Zӂ[ 0�H��F֢k�B�	9���PAÒ-8x�T��k,RC��( aP����
l��Pp�$�7>*C�	�C���τ�I.�1��F��7��C䉸b�&�s�o�:w��!맣Нox
B�I�9f�1�5H�l`�`�a�ЋS-B�I�ao�|�S�T�G'�xyfi̲|L�B�ɐ����5�Z�����"MTB�	���i�G�"�2��gB�8kRB�	 -�N��W�öQ2.Ma��,Z
!��Z�t��d2s� <���Ӧ��3!!�S�l��0SF�3lQR#AK�9	+!�$}���a�v���hSlٹ!�d&S��M	�Ծ�$ 0#��#*g!�W�`��)� ۶1he�f��-W!�$p�t`�L|��,+�F�!�$�'�!����70舠��N\�`�!�R�:KD��� &0x.x����!�dV�>�:�ˣ��yk��`>!��Ք(�Z=�P%�L6�<1PCF*!��
��� D�.BX��@�D4!��P�ٓ"��6u����5+!�$��[`�l�`�so4DJ]�D!�26t�t�� ��,rZA��鍜=/!�d�9|r�ȖF�#ZP�$J�m!���� {��ҽwq���B�	e}!�Y��0��@e�!S2Y���M{!��A�p�P�
5/\X� e$1r!�$[�~B��	����T��2b� f�!�d�!r�0:�Ħ)�b��-M(!�D��k�x�r���1��ɤ�i'!�DY�0: PQ�� R�|����}!�d�W��j�%�1P����,�y!��U�E����`��;�bY!�d��$���	�iø<��/0�!��u�*<B)�����уR�!�� �i�l��&	��S�L���AE"O�8q!�8LTLڄ�Bu�c�"O�]M_�73��ِg_j`Q�"Oj��G�ly��q6Ɓ�7B� �g"O�ԋ�ɞ@`1�3D�)X�` �"O�h �$�P}�86+�8�F³"O2�� �+RT0z��E�>��"OZ�q�lV0eϊ���қ&u��"O��h��	 �r�bA��.��c"O"�S'�.C�J=�&	�f�4� "O��C�\#g���3��,F�%*�"O��xP��<=�*%Yx����"O��Z��)9����o�O�,�"O*�X�KE�=�|���9�F�t*O28�K4_^��D]<w8��K�'�젊ա�#Y�P��@�ךhfܰ@�'��!��U'+~-J�+K�TȔh[�'\&���#F��`k�D]�S^�@Q	�'�H���-t��Qo��Ay ���'9J��V�]HbX)�T�������M���@��B���5���׼<e���A�ten��2�)� ɫfo���yb�\7`n5���67
�bGl@
�yr��#�J�Qo� �4 �e+���y�j q�j�(Q,} !����yrk��r�2��p��=/�M�+�(�yBn�< �A��{0lS���y�cɪw��,S6O^l0�x` �y"�Ǡ4i0,�vN�6\�ب�F"�+�y"��{?^���DO,R�D���`[��y2��+Mg4R	O1Y2r ��y"�+�]{V����Y���Ȏ�yR�C?X��ע�>�<�QB͍�y"�\��%��C,`��1�s�Z��yb��*f��5r�(Q�^{�X+C#��y�W+C�����BR+]N���s$� �y��!f%��a��Z�~�H�+�yBC�D�t,�G�֤U�"�2#P �y��:Iq>���)��G���k�/��y�,ژwx]���_�o�E�TL̂�y2�+>��q�l�}mB��� �y�J�� (
Y�WGW�Q����9�y2�ƹj/�j�Ò^8��D\�y!	�wEZB��uO��CG���yR���I�xY�"'oǨy��l[��y�RR����K3jB��2��)�y��R�r �BK�v�
d+�j^�yC��� @�o@�22��*'T��`�'S���!� G�|$�d�(]bY��'�>��g�0�DhJ�Ĕ|<1"�'�J���l�#�21Q�	{T- �'Q0%�S�A�Tz�8@��˂�\���'#N=����	�fչ�關8�h�'�Z���@}t	zgL��r;�@�
�'c�m�`�\'qP���;>�H��'&8)���G>Fqΰ�R+Ą3�����'�<,�f�$츒�A;|�⤲�'�*C��E�6Wl�{� ,zCp���'��0���D��u*��n؀(�'\*�8rˇ��j��c�Y]z<a
�'I^���U".Kp�b��	g��-�'K�Z�C�k.@)�A/.��
�'�r<���B�t��	+��O,5ܑ��'��9[c���b�a��L�0)�i!�'�L����FM!�).Z��:��� ��	��XVqY��Z�h���3�"O*|h�C�$e� ���z,�f"OT�;,E�mߤ4��-��%)��R�"ON�襅[�xe���t�I7>��"O��1��}FD�9���x�"P"O��	�;\����T eR���"O*�8��]�&M�{" ��|��52�"OF�haN�n�0Z�.�2��h�$"O:�+w�[�@`���&���Q@"O(q���ɾ}�$�Y��X���"O�8q������^1P��yb"O���kW�I�Hp����|Z*Y��"Olp"$mL5VLH��jҔ�F,��"O�i4�C��m���_!R�0t�C"Od�;嚃Jd���glS�?r����"O���Rc����D��9�!��"OD���,���!���4S��]��"O��j�$�[���!�"�*t�<"O�5k�f�#9� �Q���v[@"O����c��P9�������"O��ksi�<��J!�)�\ X�"O��X���~6>�@��
z^�Dr�"O����Y�"<+�oG>3��pq"O �ThB�7C�aQս-h���U"O,d���
�28��2GS���"Ot$��Q�܀�BG�B7���W"O��HЉ*9�0�:��=(5v"On|� �)EUR��A@Ȁ3���%"OH�3B�ˉS�
L�D�u?�c"OJ��)ح`Ă�`�mU2p��I�"O��Yg�X�Ȃ|����=w�j��4"O(�VE9��l���1�9"O�9��ȍ\^mk1��6Df��"O��;��
o����E/j)�XBa"O�!�e��+e��x���ՍO��(�A"O����T�iED�(��T$B6
e�"Oʤ0N%ubR�x�!�= 1" �R"O�V��-9H�J�`Y�a0֌H"O����Gf"��� Y
8 "O�����l���D�j*P"O0P���4MKl5�7��6�� "O`I�e� =&�j�� �K]�#u"O�( ���6�Ȃ�ŎC��"O�4BVM0n��h�1�P�6m[�"Of��F��x�$��u��(��!��"O`(�(�1IS4��c�A���	�"O�|C���{ڶu�+�(���a"O�������BH� ���=d����&D���K�C|��C	��`����f&D�Ȩ"��40q�j#�>������#D��µ���UUH �1�I;JrRB䉅;�4P�c�1ZzPI�*�8�HB�	�n�l�"o� i���1Gi�~�@B�	�N�2�Ae�O�)Jt���(5HB��,>�$��N�t }X��S0E.B�	8�`��%@"c"��9���[�8B��wo�,����-�x���T�(B䉲f�X��l�*6�-�1gzq�C�*� ۣ�0�)`g���C䉞$��T�W'�j���&Uw�C����{�n®C{���W�ޭ�>�{��x��aH�2�l���d��a��3D����d]�y�6	r/D�������4D��1U�2i��"�"Woz�q�2D�� ���S�V��
"+�?˴���"O@�*�@��ุ�
�4A��\K"O�0��^Y8p����l>U�R"O�d���3��ibec� 48��R "O�mr7Cu�*Ca¤g8D#�"O��B��T0}>�{�G1.-��+"O�S���}#n=j#.&_
R1�"O򕂴o��B�s&�1���f"O��R�����	����6����"OX�w��$kG`�
��@�E�X@�1"O��jE����*� u4�1&"O�rG���g)�9��D�'syZMH���I#�l��"B��J��B�N���C�	���u!p!B�_��)��L�[�B�	
��l��9e�Qb�L�,w�B��i8
0���+I&���V�H#B���6ě@�A�P��3�#��coPB�	� 6��@7�E��z���L�d�C�I7.�6$�vft
�����2#C䉼+�i���&_��|J�Fև9��C��!oj�t��3`�UXg�3#��B�	�	�nō(�0�p�n>��B�I�tǞ5��'۠�.�iG�w0C�/[����3&3D�����;�B�I_�tP���l�0�;�dD�|��B��{+����E]�����sD����B�I�k�h	5�N���mj��=ԔB���8 &�
k�͡��W8%vB�I>#R!@vC�B(�dp�(�:%.C�2f4Aq'͒nL����Ä�(��B�I)p�b�@"k>b�P�n�t!�ط+q��F
�t#�i����)m!�3Q"m��ϊ:v`5 ����	�!��X=�}'�A�t���R0 �!��K�f�a���J{��C+��!�D �_�9��2��y�G�
-K!��#Q�EZ LK#G�0限A\�_-!�]I�(�(dE���PSt��7;!�$�*���t�,VN �_�`!�9njH	�EJϗJD�xهOůO!��΋}G�����9,@XrU(˦V]!���3pMtȨ���~%�%� �̑UV!��N�N�ك뚇B	�,r�Ε�5�!��7-^��pg^Sc� K����!򄄣��aɴNR�SQ�-(��9�!���g�`!!�%V����4�!�T�\��i��惵"2hQ�OQ�!�(IN��&A�"$���A-O/`~!�d��6ukU�G�
��'�6pq!��J2:��Kf�s��=x׬W�0�!��9Kb 1g���fLvlP&��hC!�D�r&xk�kO�FCZXzPl�^1!�^�,ai�i661J��ӼD!��`dh���5��m�
N�	!���}0��]$.r��R/�!����6,(f���I2�P�C�9Y!�d�=�.���%d�p��l��
W!��!`�^�z��ƄR�C�� /I!�K�r�tY�È#T���HΩI)!�Ćt���9�Kǎ~�Ӥ&��?�!�D�/��I��,9�������I�!�$���&ȓ%����(�HE�$�!�L���|p���(o�|}*�h4'!�D���\�mȍq�2��3e�1&1xB�)� ���Nh�$��&  ?L|�t"O"5��D�K�p�9��S?\x�f"O�i��eǄ
���P�:"O^����K}���bg�x⢥�"O�A��d����StZ=�ч�b�<Q�m�o6�U)!XO�y��ŕ[�<�` ��|��Ca��=����Ą�M�<q�-D&&8:v`9�vHs��@S�<I7��M )�o#,�3
R�<1���������C�<�MJM�<a�(��m��9'�[:� %�`�S�<�0#�"$�h0�KϫvP��K�h�<	�C�	�(�"�⎐rc"ٛ�"L�<A�M7�*){�gK�TW|X�1��c�<�����G��ԹG'D?+�X�ʇZ�<1�(K~	��xm�9R�.�qmTQ�<��i�13�h3$-'����͊H�<��#�1N�`�@#E�Lw)�1
�^�<���+{�j�葬
�G�!�D)�Z�<�p-�:� ��ݟ!d�[�*@�<R�������.�$m��*�y�<)�D��� ;F���`��p�<��L�������Ȋ(@��P�u�<��!0s� h#Ŏ��;|	3���Z�<��# *  �   V   Ĵ���	��Z�wI
)ʜ�cd�<��k٥���qe�H�4��6_2<<y��ʄo���+�􀷅�5��l��#D�#7�6٦���4Fs�*�I\y��7f_��k�D����ة�L�G�ԁ�%�vJ�9�=9��9g��7��,#�U�ϐQ�8"�'�Ir�dT�smÄ3m�"A��y����
0���p�2�NS"bzpw� E��0�B�w}�%�6f�^}����
��zל���G�a >�(%\���b�c^4)E&\I ��_?��?OT� KU�� �82�S	:��	�4{D",�@�p��+��I2���S����9_�PL�'� ���*���'�"pR�Ƀ�,H!����6���'��GxR��m�'cj0����y�6���"{t0Bed6�>�r#<9��>�c-�%X"��V$�(�f+*�-�O�J�{�)OJ�͜W�L�*WCW6�MS'#>�C�#<c�B�p��x��Ĵ41
4XU'��L�>���;�E���.<��{���m�us�f�,?x�'���Dx�VI��x:K%��@�雕�ا;Q��s��/��#<ia �O�8�h�5LF�$�ӎؾ;�j�*��d�>�O$� H<�O�-���Cb'��3Y&D�ѭ�x?��� �RxHOFL��b¸	�&c��1���w�R4�I4���f�DGn<N�'�~"Cg��w�t��3MX�Z�Te��W|�|�$�6ቹ!�$��B�g�TV6�k%B�
&����'�(XEx"��z�'NV<p�K*-�<a��%%ڍ�'�vݳ@ ���W��o�<�Go�� J��Խ!��P:��Q�<�'d�rI��B�j#��U���UM�<�B�#��PK݉iή�X&��K�<���\P���ɤ���B��؂��H�<�R
4-h�8�'b��QiKN�<Y�NG��Ǫ��fJ���bEFG�<��L&�.t�Ql�Q��pP��E�<��#ܮZ&���g';7V����<��'E�k{�d�0/��I�4XZ��}�<��d �E�� �L�Rj� �a�<�B�E�`MVM9�lF�N��F��a�<�� ePP%@f�ϞV���xR`�W�<�4*Z��Ɣ���\�5���"��l�<�"��2]���'	��2ސ�+�H�C�<y�6Q�\��q�z6�����W�<yF�ʎq�jDʓ�> ��W�<��	�&-�2�{��t@n9Q��j�<�HC;Ģ�    �  :  �  	  M"  �(  �*   Ĵ���	����Zv)Cll\�0R�P��
O�z��1Qv�i%��/��Qlр�yb��Z���Jc��?��J��ߪs������I�<7|�������ݚ�-͛J��j2@Q66�X
�ڠo��	�����N�9 J:��� �:OC��j3iZ�5���c��&h�St��� �����O.:���3�0S{����ځ8����$��A{�A�/� _�D�H�&�&3�@U�u�<�Iߟ��IڟT����$XM�@
i1��		sf-c��gy�AM�$����'
R�bt��^H���S$FlY�I7|��tŎ"d�$I"�擽���	�p���Հ���1!��K��Ξ��@	�\�M���'!��ٓ�'yB7me�,O������b�&�vY&�#1�ˆ@P��r�3D������H�֡Y�!�spAP�fl��!Dz2�H��V�d��� {n�����f�r��N֖����������u�'��?���:��'����[�l�"Y���n�[�@(�O�1:�Fȃ;�V�j���a!ǊͶޖ()ʲ1Hn�(�f0<O�8p�'Rt�� �qU
�
�O�Mꄸb�%D��ئ."0�`����cq���?,Oz�<�$��H�رN��Rl8zUŗE}��x��O����i��=�dJ#���w�Y�&�ir�3�؄X]ʴy'�N�LZ6\(�'���bPM����K��U�)�'��)�A����M2WL�H�p%"O�@�OL�H2Ld+&H�ii�h��"O�9c2�ȝ7�@�l�'1~qQ#n:D���� ø.��X��)w��A�A8D��r�+ԀA���%c�	0� ��T�%D� Q�A�'�Dո�˃R��C��8D�4��'��?\X��2 .Ӫu�ի1D�p;�Y�tY8��@7n�8c�A#D�а�!�Vr�+EcC�^��
t� D���JK���i �M��{We2D�T�R�^�P�l��	�418��!�%D���B�8��X�!��(]�@B#D�ر����x��S���b�� D�蒇�T4�<j�� /j�XHPF	*D�(* ��C�l* ��><���*D��D�o���P`M�2o� ��C(D�lAbn��FFX�!G��A�����9D�а�B���*��Q�Ug꼁 J'D���6 �t:)Ҧ�Pe�8��7D��!�-c�^�8�	�2H�Q��&4D��ic�OZ&�g�{K���"�3D��2�g�*�~|���'�Xyw�.D�|Hb�	;_��dy3c��W�@��4,D���n�����[	T�9`���ybO�5V�y L�1&��;T+�(�y�B�2�`�F�_�.H� �#�y� C7)��q'�\�(ke���y�l´uB�5I����X�H�HMJ�y�MZ�E%R�RþP���¦R��J�'������=�\I"�iĞ���Y�'�|�T�K&��I�Q�� ���Z
�'�N�E� �� [�@�H��)	�'��C��W�l,��瑄\�����'U�5A���o�C�F]�i�8py
�'j"��`��%:p(Yǋކw��$��'H:)��ω?��j6���i�4��'ðĠ��M�F�Q�Ի�6���'d��zV��<~�p�3T*���,��'�L��`Ԥx�"T0���?	���
�'a���A�$kj�킲e�,�8X��'YX0�C�r��8Ů��%%6�Z�'�,�ap"�D��ybm�M����'��D*wl�<a��%��_61�ب��'���0
T��n�YT���+ll=��'��t�$��R��|Z���Y�x�h�'�D��gcL�C:�x�QC%Tt6���� ��:@�prE����)�H�*b"Op$�@��5*$���I(4��I0�"O��Đ��h��E���V��}�f"O �:W.�4��S�sz$̢"O���cH��k�$�+��[��*q"O\�Q�f/8ⲕz�k��7�0�X�"O`B���(C�X�{�	L!���"O�!�f�6��9š�;��Q�"OȈ�\j�@;��Y?���r"O)�A/��imN��n x�x��4"OD� �Kޯo��6ƍ�q�BAs"O�ء�n��Zc�䈲%�:j3�	�"O�X�e4R�I��g|bxcC"O�q��I�Z��̃�'ֆN� �"O��X@����mh���R��D0�"Or00PG��0�V	��mB�+}H�x�"O�"�,Q
D7��``���i��Y�"O�Q�Q�N�N��"g���!-
I[�"O�����-�ҭ��׹2��g"O�pQ.������D�*F� �"O)&h]�f���2+��,�@��E"O��K�	�2&if��	E�S+��a�"O~A#�H�
ގ� �ʃA7<�`�"O��C���1{��e�G8+$L)�"O�<C��!�l�3�\�:��]��"Ov��fc �X����U��q���s"Oz�[Vůd�ޘ j�*N�R�J�"O���q R�"E>Xs�->���:�"Od�+x��٣s���_X*�"OL�r�dҿ;�.�ȑ��7#}PpY�"OR�I6�ݪRj��0��+Aa���"O��0��7yԚ��SD�,_Դ""O��B� ڭF"�eX�H�_D��8�"O��Ą�&4n`{��B U[�`[�"O�DBҩ�7t�>�lRX��c"O��χ7Oyj�+��>C4tI:F"Ot��B�!3e�=Z���\�$�"O2��!41=@�ccU�~�5"O� zqd�1#�d�CC%Y*=2$��p"O2�)�H&�V�!�k�*`b��2"O)�7F��,�nm���ԝi[�4�t"O��K�f�8>�V�xk�KsL5I�"O\`���\���&G�2Ig$ )�"O` �V�F~��v��<c1��S"O @s�G	�+}�Ǔ%6��c�"OF�X����Z/2h3R ,U�4"O,%�*N$t�h(re\�E��P*B"O8����Y$<�!�ǭ[���5"O��!�+^�%��[�-Ɖy8&=�"O��Y��"#�Ey��#7(��ل"OL ��z܉BЂ���"OL���G�Q�.|J��^6q��d�f"O������;�5(eH�=/pԀ�*OR����B8O�ܱ�D��c��M��'�F�q#[.�o� ��Q��d�<��'}�>�I�C�6�%޲�,�����}�C䉜�"���o�ZgFă&F�����$-n~�I�	�Y �}H��\6(|�x�_�1v$��I,v�|�z�O�q�v%ϓrݎL�#dA3�Z��W�@�ՆȓU�I�2-
8����#��&���\Z�Xa��T�O��%�57~�в�ʻ}IJ�'����C�+Q�� B�7~"��3Ə�}䀸���O�s�/�*����H%9����K,\���ޡ)�f�R�AY�-�by8�Y�き��`p��UZ��(���%����S�? �|HSn��l�ИB�o?몐��'��dY��*=���ZS��E�>�+gk�3s#�M!p'^sU�ar��yrIL�A�ॹ��^�UR��N���$�v+��:&+��y�.��6�	��(��e+5$��F��ق��T{�TD:u"O� �6��c�k�BLvn8axkG�M&�&0+��T� g�O=1O4AR �&U2�s���J�P��'h4@P$DZId����
?8��Xrs��H٤��@�K1��g �w'azrՐAZ�#�	��Cq��@����OHj%�H��#f
�ctf�A1l@�oJq�@n�N9��Q�̐G�DC䉕^�A����blZ��tnm�˓K���kA
Դ�x`��$?��u����Ԩ�8EI��~tލ�щZS�!����X�B�/2��dÔ��xm�h�%A����� �,_��щӞ���ܰh�.ʲ�ߒI�kF�Q��Ԇ�I0C��I��4u7`�A���P!�F�Z�$��@Qs�=t=�˄	R��4��/_�.(a�d�xh��&g/O�uC% [?`�`ŉD�Uy�PГo�;?#L�1Ś�yD�AjW�J!Xc!�čqc����;1���[�K0"Q��)�~�	[��81�����	
�J��� %ʁ�6\
U��u�!��M<dB�ӭ8��\-(�ɒ���e@��M��;�g?�G��;^Thq�E�6����p�v�<9 ���h��D��Q�ء�����1A�
�SH�V+:lO���ti[� �`���,�]H� �'���e�)U����3N�v������&N1�v�Η_�C�	�挣u�X�Pjru6�M$�Nb��z��S�!�����T�j,�+��l�1ѱ�I0.!�	�P&̊��	62�� {��D�q
a
�L�<�Q>�':����f�gV���W�SuDćȓ���	G,YW0���ʆ],	�I,pń���[�T8עX�W(��gH.g�C�ɂ#�R��AG�]x�䛓-@� ��C�@r�x�k�"x�( �E
N x��C�	~kv8�d+�Q��Yk�C��!_8�(�E��A�<<�`�YVB�	�"o�#�dK�%&�W�\�"ZB䉤Y�v��oӣE��(1#�}1(B�ɪd�*\j�����$ę'?%�C�	����S�/<j�����lZ�A��B��	}/<���O��}p�9��j%E��'�(u@�0�,�*�+���*�'��x���B#_E�@  ��d�l��'2HAxǆH?�1�-�O�"i�
�'��zT��in~��Ɠ�B����'P�54�՟B6���'��	�'���B�Z�?��<�Ѐ�5��œ	�'��y�a�� 0 �5���A�a����'#�����uA:Y��g�jJr ��'(�y˱��2`�ja�e
��p�N%��'rz`�
ØH��@I�[��VY�'N�J�o͉J`����A�\��eX�'����%' �z�kRa�&d��'���k���9lrQˡJP����	�'���9��Qk�}8�O���65h�'�(h:���t  x�P��^B0R�'�b�*Ӫ�=Gצ|s�)F�����'1Dhd��'����d�(>�r�h�'���P�+��?aM�b�'G����A�SRMP���n����'�d8
�R8<6� `�Ə*}��`�'̤j@ǃN�H�FȆ�u�p=��'u��z@�?�,�8��ߩ_ox���'���2�&M�)|��$�F�Vt�
�'�s���i\ԝ����0�� #
�'Xmp�-�n�Ѩ1oך\��'��$�2S&G�4I���q8����� �`��\�1k���QAP�Q�Pq��"O��r�j�3n��"p�D�.�JU��"O����ؚ1)�$ �`D�g<H�s�"O��{�jY�*����l2A<ٖ"O�I�e
ǣO�j<y�Q/l����"O��G�F�}t�뇣�j|���"Oʼ3WU�9$`��z��4"O������v��!�#�Nm��"OhE��i ��0 �Q��Ԁf"O��[��L->�҈��ܾ?�d��"ObS#�Y2������PH�~<yA"O��	��I�G[�D�5�ܽX�j�j&"O��z��N�[v�Q(�Fԛ{/^	`D"O�\��m��o��!�A+z���� "O�؀�i�Z*m�d	!72ay2"O(`�eCҦ����Ƌ��u2=��"O 5'32�N����S�c"O��bg���~�^1ҧS�cG�)��"Of(�1�ƆY`���F�?Y*��"O����-U��0veN�>V^4B��O��xY�쌡3J��� :��7-U�L�(c��?��e�q�V!�� W�H�&	�Ԁ�A�M
I>!�E�� �C"T�V���g�ƺd4!�$:v�-�F@��V�)t��Q!��r� ����˟6���cĩ9?!�dV�q���e�#3�~SD��<�!�	
K�[�b_�ך����0G�!�$�(��%��S˶ۇ���!�O�s�0@�5�U�I�ĤK���7�!�$œR�j�fd��S����t"O�H�!����I�!���UK�"O�4;A�V21��		�O6y�p��"Oy�+8��)C@��?)�ݙq"O�D�&�b�<0��jV�k:,�@"O6�Z��Ί]�<(2�Oؙl��I�"O�#g��]�.���=W�9�"O|؇��9Y[�!�"āYIz�v"O��rF?O��x5aU�䦙�"Ol�`�N2� �4�X�"O��@��� `T�2S�T�SC"O����
B�>)��iv�̆��d"O��i��'xҲ�  ɝV��1�"O� .]��X�Pǉ7\���"OV�c�[ u��pb&�2(\8��"O�A�E��=<=�����L��C"O:X$	�8�(mQ1�S�{��"O��[���0i0�A(E�2�x"O	`�kӉ$b�
��s�.$�c"O�`j"��
Z~D���?r����"O��Ch܆~Wn�I5K�:��YP"O�E���,d�� 7*B��6�"OZ�	�DI�}$I�A�-��"Od��sn����&���U�b�J$"O.����x�v�9bh��$�0"Op���0�L`i��+�Ƒa�"O�pX�hS0l��)-�� ѐp��"O*�� E�.���(І.����"O@��o��o3b�R�ˊv��Qk"O�y��/QxI�BO�F�@�ۅ"ON)�'C
iS�M��!B�7L6���"O�����P����_>k/:�P�"O����M\�Z���#�(� �"O&ՠ2���w����DM�y�xy�"O
�#�<(`��uaY5�4rE"O� 0Is��Ѥ'`C�$ـ�r"O(��ĺ'?�$���ĀYÒ1d"O�Esh"bh���(��m�L���"O�ÇH�Qg��h�F&��A�"O����>k��Xk�`=fB�"OPmؤ��;h�C�D�}P�u�w"O��� m� ��|���!t5<��"O\s�.	 +��a��-3�� �"OLə!�ZL�k+J�F��]i�"O�������4�Q��3��9Rw"O���,�e� ���[3�"�)7"Ou
&��q���������H "O�<�#
	?L���h�`��P"O\�%e�+�f�Y� �"OZ��'��)70Y���ΨEֺ��d"O��s�
�?y����^��!�T"O��%�pH�5�ug�3L�ĭ�7"O�ؚ��0,I�E�2ZJ�!r"O��
w���?a��p���'Ut�3"O�L��➀9{�$s�Ʋ+���"O��B�d͐K�����	!=��D��"O��b1�^�1E�M8"�-f���C"O��QS Ա!���;��T�I��"O*(7��/t�
�Ҏ\�-9F"O��*�Ç�-���@���D"OR`���f��q�P"@ 	�"Ou0s�
�"�(d
� [�lfX��s"O�mӶ��=9��i��.�-V� �� "O
y!b�Z�:��S��16�T�*�"O�)�lWU��$�Μ�&H��#"OD�����WH��Z0��/5<Ĉ�5"O�@Z��@ �\��%�8IV��Z�"OV��`gE2�<J@�B7��)G"O�aB`�� Z��ɃPA2l$t�;$"O2Vޔf�Ze⊻H=����A�<���̟3�Dʃ.���,乐	�e�<�p�^�SN�����L"+��MӖ�T^�<qg����x�B�I�M|D�rĞQ�<�Qi�=� �5/��lE��d	R�<�����0�D��tm��7��Y��k�Y�<!E��+X��ݳ`�]�5�ά��ISZ�<!�NW"�4����ي���ˑmKQ�<�����=��S0HBݣçK�<14�ʉ2�Ш�NRy�\�� �	]�<i"�AG�4��$���*?�U�<A�jT0ю���g�bi����b�f�<��&X�.�9pv�H$H��t'Wa�<!�m�V���Z�����p�IB�<9�ɂ���j@`Q\c�h:�LY{�<!W�F!t��;�#�tWJd W}�<��m��Π(�lЍN��f�Lx�<I��������i�Wn�u�<Q�,K+hS\�Akؘk@U�RSL�<id��}��'�y��Q"}�<YƉP�>�L��BL�-�X�	w��x�<��ɍ^7~����
8�
4��*Rt�<ɀÞx6�����>��a�G�<)˔ .����ܱ#�m��f�C�<a��Wb<�
L1.=�]BѪ[�<1�f���1�,:�BF P�<�2�����R�ϗ(R6����<1��d+��s����Y���$4�dq�ȓL�D�I��-�^\qI�.�T4��Im,1�0cW�)�x0a�כXpх�S�? Б�'CЫG��� �%6�q��"O�����dp��N�
�2"OFÐ�QK��qfS46f��B0"O�I�&A��&A�;Ċ�-u6je�"O�؊0@ԥ/bdɳ�ɀ)�U0�"O� XAJ?yL޸0��Ɋ3���"Oq[TW&S�J�ХP�;�]Q�"O�q���U%���C��S!6 �['"O���ѨB��d!���Q@'|\qD"Ob�`��K)nH�|�ӬM:!��"OD�x��L)*N
�S���+@(,�u"O�c4j��{�� �!��v�(h��"O�����M0:�cB!I�X�.�[f"O�退kݶZr��o�,$�N(��	V����
 �L) D�_�#�ʸ���G�!��Wd��C�ɀ/�JXVH��|�!�̩l����V�ɌGS�}���R��!�Č�C�̉�E��& ;�LA��!��W.����#hڴ.�s�K*	!��J*;-Z��& �*$���)7
+x�!�D�M����I�����"6+H�!�م3��pfl�$;I����Ӯ{�!��U�`�����Y�R3p�مD'�!��\�5KDC_28���-X'R/!���o~~�;��P�uc��5N��!�A�%���C� �&YD�H�P'׻�!��\�<G���G���A�$0!��5�8ત���W<��26&�}#!��	b�^���M7N� ��e?�!�D�2)��ÃҔ4���Q a�!�D*[�<��l^>AU���T(ԛ/�!�䃳<RJ�Z�h]�cTT��&b_�tu!���8���ŧ#ޘ��@T�It!�$�df$�K�h[%5x ��O�Vn!��W�hA�q�.��pU�?8�!�DZgC��X���<�s��L�n!�"3�E8�iY�2�漲���(f!�d�;j�0`ș�n��"石n!�ğ�܅�] Y�G�.���	6"OJu�1HV~V���A���N��f"O�!pe`�%t���bB.@�B���"O�A��3�h{p�����"Ob��$W�=��4Z�!W�v�bt��"O4	1�B�{�R|k� L'd̨a!�"O6� s���v�*���O		�t�`"O��a�/�a��a�5�^�,�vẓ"OpUQR#�%2��=[�@�t��Ui�"O ̂��4�h8���?#as�"OXT����W�N`�w ̨����#"O��q�ٹ)�A[� �'����#"O�@FL4�q�S $�0u[�"Oʐ��O��d({G #��1��"O�1��r�X ����"n���xV"O���*
�R�dUHP��w�.��"O�a8� ur�8hجw�:�j�"O��#�.��Wr�s�fĲ?��+�"O�A�T�o �87� f�	y"O葢�LS(d�dq�#9}��	�"O~����ґ4*
3���23�*X��"Of	�֣�0l��Q�s��&�X�"O2Xa$ M(�<�O݄Va�(��"O�9(DC�:k��ɣfܬB��i��"OL��6��?sN�eزbF�(�0q�V"O�!`�D��6ܰ�OZ��E"O� �8"&/�#fD��	��{\��"Oji��這ts�ܺ�-�2N��"O�#Ř{�XʷM�NKZ5ˑ"O����R,|�x��'A(�b�"OZ���-_�&8ꑮF�F�h@5"O��27.ws>��ūX��M�"O�i�Ս�18G��mJ��a�"O�4 ��	�7�`e2��M& ��J�"ObqӬިk�YQ+�,P],��3"O�y�5��?���9�L�.Z����"O
,����>O0���Zm5�x��"Ou�#,R4M�4���3D1��Y"O��zE�
�P\���x���"O$Q)&8GzZ���Y^���"O���&c� �&�[�L�!X�|A�"Ox���R+Y�h����>Y"��bE"O&q�Rg\�,1�A!;�V,(�"O�0¡G�'4D0���Ru�8�"O��Xq�S2��˒�G�=Y���$"Op�HAȏ�I�6`��IC�>@�)�"OV��C��2uB�� c���6"O���B�ͺ
(Y�e��]����$"O�Erv�W'pRl�BBZ}���R�"O���✉T�P)�b�VF�(��"OLm�b�
  �   b   Ĵ���	��Z;t�J�(ʜ�cd�<��k٥���qe�H�4��6]22<���ʄj�ևݪ(�䱑Tu��@��M��7����Zݴ1t�+��]yRfO6d�>	��X#�J�2CĂ |��p�#p,���=1�f.&.7M�1�biy��C!V)����ΐ<����l낊]�[�!l�XL,��<3-O���I�Z\R��Q��(�h���H���u�' ��1PB���$GX|���,8k�M�B��4�T��b%J<��&�x��F|�ΧmH�$�'-e^�X۴O��0i��@+
<���A�Ř/���e��y2���moN���������'/�ȓe���/�$e#�O���t/@0GB0fH
&x���կ^*��p`@���'�~�Gx���-*(��IFf�.	p�`���B�#<AGH?�]���@���"���~HB�ĦNHI�O��h��\�',�uS��4|���j��K8:tr�4�"<� �.i��	t$�@�L<A��ȖH��Tr�Z��"<�A�-?�"O��Uz)�/? i���ey���[�'�@�?Q��(:�6=���QD^��Ф
�N"<aSa(�<l��D�OWH�n&���+l-1O~���$�/����#��2��ʁ"����G?��)m�O�p��4��i�e�] a�2�K�^Uo(���!���ɿw�����F�O������432�9��۸x#D���ƣ��'�JDx­�V��= �q�F�5�8so��E�I���l����t^HCŦ�#SJ�Q��" �.��C�I�*}z�  �ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��t    �  o  �  F  �"  �(  5+   Ĵ���	����Zv)Úll\�0R�P��
O�z�����@��?�64�r�"�y���}���c�Έ��Q�0ē�1�읻���:N��t��n _��CKܼm��C�L*6�^�Ɩ�-��}{f
�|�xI�mL���d	2
D-��,a���R�XЈO�.�x�rXs_@]!` �1n�'�"�D�c2��t�u�`��#hl�	X0E@�/�nX���	1ƴ�s�H�7.zX���'��'be�~`j�]��i�Pb!2��#^�1�ə�4]i Ã@��dSud��$Z��% ���@�jϪe!�5 &��z\��x�o�?�0ʧw�:��#�iV�**�26��4n��5�G0>E9l��4���֟� ޴I�<A���~b�S'���t	�Z.Y�S��y���|��*�$��š��� �MK&�ɋ�|�Iyy"��X>��FoG  �,� 9\R�K���m���'I��'�f�]����I�|�wiײ}�lu��O�6TC�'��@�­I�eO�Vs����gîyڼqw��7	�� ��0�R�Ї	��$��}ZB��,O��`�hG�M�̕I�ꓺ5�(�TJ�	�H%�,�Tj�O @A��d�����B�O#T	{��˦�s�4�?�(Od��;��~z�g�i\�T����k������J�<	�N@�"�f"U�8Ld򃥐A}�>,O�$�"ǿJfҥ���H6�	պi��T�!�5vZ}j֨3jr`p�'K؍���*�>Lk�EƑ`�B�'�6�Q��	+��aI��� ���'��D��T,U�\
��ȵ(�}��'q ����V�s&��p̕`
�'����t��7%Z�� /͚$�v�H	�''��Jvm�4L�"���Y�
��	�'�h���ն^�,�2�:V	�q�'7���d�QBd�;�&�OEQI�'"X �E�J(S�h̲3�ā�'���)�b�g�r��T��Z�����'X21�Ѝ��Jㆸ+�'��W�H�'��t���/Pv�]J�瞟L�p6"OhACoȪi}��s��
��<��"Oؒ �ڒʖ,��A�k���Sf"O�l閁�-QZ�2s ��$:�9b"Ot9��O��kr6�[�ɐ�eN�R5"O�����X7� cFH��)M0�F"OP��E���؂�O0C2�;P"OL@إ����h$z��)͔]�P"OD�A�C��5��S[iF��S"O\X��D_#jۘ�C7���l��"O���0-X7	Z`�K���lAb"O2��7��b�z՚B��p2��w"Oz����;N�x*Vaǹ{%�"O�y���PN���9t��$T92�"O8�;���z�����@"Ot�r(�6+:�T@��.��p��"Ov�[$������!w��t"O�0H�Ȍ����ך,o���"OB�C @ h��0V��/E �B�'>�����$-�m��޸W�!�
�'!v�%j�f�P���ÿ`���`�'ܒ�#)�;^6}1�����N��y"�-��L��D
}u�QySҞ�y�O��Yx�Kɉtr�0E��y��D(Oh`9�%D�i!,9��M�y���weԽ؂#T],�Zb����y��8+�t0�g���T�E�=�y�K0w�bs�k߀R 8���=�y�ZP	��*DhI�����R˂��y���uȖL�� ��rF��yBk(�f@tfN�K���^>�yB��Cl���>H�i�AB&�y��@��\�t��{��9ۥ�,�y2��.@�4Ó��w��H��I.�y����?�0xw�U%\�2	��JN��yRC�&quf��1��=P�p���D��y
� ��ڴASc����W�K�hƚ��"Ox�IĪ! l�2��G�X�<�ap"O�|d�ۍE�x�)5%�8�;�"O�X��mϸN~h1�R�� �Pq"O��JG�
7�R��g^0S�hȈ�"O��H��߶T5Z��4h
�g1�m �"O��BV#̧^�F	��3yM��x�"O�Q�A-^2^	�5'�!����"O�8�� W	�9)����<�"Oڭ���M�
�z�9vʔ ��x�"O���Į��d+ꌨ>6�1��"O $�EN�(<MvЩ��T�Ijd+e"O�a3ף#c���ƅ��4p"O0�p�T6Kv@a����n�F�z�"O��z%�C���F��&��"Od���
S�.L*+�jP x��-��"Od���&��@}K3jT0	�)ٵ"OX9
Q��q�FT�h�	YQ6"OU���ؓ)��̃�,�5�!��"OF�ӲhT�|�X�R��'֒�r"Oh�27"����W�B�6l2"O����%�`���V-1�I�%"O�r��C3�S�f� ƐQ�g"O�]��FB��|� ���F5,�a"O�E	s�_�8;&��"ƥ;��C�"O��
�� 7n�6Je4N�(c"O�3��šLJ�p�B*3U%V�""O9��Y,	�0P�
�'"f��'"Oе �;/ ���qG��F`)�"O6���
V	�qI�e�)���"O|�B�2[�`���]n��0�"O��8���Pq&�Z��-A/�A�"O�4�'��*/��{uA&�{�"O���A� JI�,C���2-�i2�"O���� G��Q*�W�؊�"OtИuԫ`� ��H�C�EA""OF����D�B��:clK^���ɓ"O<�c����@�����̐"O�HB+F*_�j!����S�h� p"O��BV%B�1�u�c�btr�&"OV=�����0lt\ˑ��@T&)#"O�{N�?�FP��-J�aP@xQ�"O�l�������9Y�Y�"Ox�P�L�?ܘT2�`L�M}�Ms�"O>8�2cT/��A٧I��XZN��w"O�����T�vmҠ��]�ވJ�"OM�ej=L(*���FJ�|��0"O���c�Û2����&�,Q~���"O�8��d�
�Bp�u�P�l|�)"O�PF���X��
Q����[6"O؜[�� #5���2dk�J��!"O��)�b�N{��`�k�[���rr"O�X�a��>��(��L��4-xW"O�K�-�wF����^�.�@�*ODx̛&�ѡ@hB
��%Q�W@�O��}��J
⠁�c�'
�@��_�@��� �|��i@8aq�X5�Ƙi�*� �ѷ:��*�Of��e@�&+�1sN�9U��)��'�� 3w^�yվ�+�h�O�U�#�(-���v�C"�H��"O��S�Vu�tx�e������P�|b���NA��Tm�xun�}�6��_z�{��ѥw|B��@m�J�<�p��D䘲�
�� *V��X*KzIpI�	;.�6M�*W�BI��L>)�f��.6
1tDD����E(<I���5r�Qf�M1(xY�A$���X'O�<�V�������z
� ������9�q%3��I��'�@�b��Q�ka��]
&`�l�҆"M�$:��N�{��������yB�3hv�!s�o����0�����*_Rp3�i�C�y`�$�>EQ-`�D��ț�Iq(9�!?D��QPїo�6�sVcԫwa�岅�9E�|�2`'���&��60<&?�xI>���eC0�"��3�~D{� J�������v��-RB!I�QJH�D��;� jCB�e�������T˴��\>���łvi\-Sl@�#��G�G�;T�ڤs�l\�A��!����h~:�y7I�f��xH��=IvD�34��:Ө]����N6[e$���͢<iBb�zYl���K8�5h�����?š��uZP���-�2Iw��Z!g4D�H�����kV��+Bpx�7���!8� �柞&E�vM.oyfU&?QaH>�Ү$�F��7�[�q�P�b�jI����֦�!��@�_>H���, � ��Y L4�tr�+��!8Ʉ�(>�f�xC��s��I$gDI����;2��)��^y��I�rH�3�	�/V�k��6%�5���2�"O`P���w���L�4Vy�%*����d?�!"	#4�(Q��b�O�i��`�B��A���	�"ܬ8��'N�3�E���؃f�_� 2l{R�D�ys^�8�C�]y��9�g}��Qܴ!�`�A�Q�1;�`ȯ�y��S0.��y`��X�M!���M��5p�����\؞���"�W����"P�[+����H+\O��
P�ƪ(+z5�&�'��8��!��3�����+Z�i*�' ���wΕ!�n͊�L�B-H�}��������/�[G���An���SH� D��<��p(��S�(Q�+\��N&b갠��u�'j��E�,O.�ô-��q�:�X�N�6nP�"Oy��_0:WZ Tp���]ßp�G�l������#�p��^0{�vI��m=D��&aQ/.��Вc_�+���z�d(D��B�]�,�j�Y�B=�)�-:D�ܩ���N���HK�i���q4�<D�`��	;��}s� r��P2�;D�P�5�_#c�컇 σ>�����;D�`8�<^ ̩���RC�T�e�8D���u���aD<Jdʖv���YE'D� A�N�h.�F�._aZ�S�f$D�� Q�ׯŨt�R+'�Q>D�0�¬�h����!��r	'D�����I�,���Ǐ�L�4� D�<�T�E>9:0(q��P�0�ԝ��.D�ɥo:X�u:�c6T_�R&,D����n�3.F���A6Y����G)D�xk�K�>�V @V�4}����*D�@�G�G����R5<5b��<D��B(ױD��)s6��1[Z^%J� D�\�d��,� y��-�Q�q��O#D�k�b�=&����'��g�RL�D?D�����J?}�:؁�B�=ju�I'D��-�S��]Xf�0"�A%D�p��a�k)���͛-%��%�)7D�hc��ȐG��A���&'�3�3D��SlI 7��J'�	�� !b��0D�\��2�u��\�k��q��'��4� k�6�<�F��l[����'$��S0�FRlqq6AO.7	:0	�'�`m�㍎�
����Z�4jm�	�']�)�!F�;������2��Dc
�'����#�S�7�h���+[�	�'��!�E��$�H�" e����U��'I�a!w�	3�8,�*�T��A�'Az��5�ˈ/� ��t�>&<�
�'���!���aMz%����"��+
�'r�"�N
�-)�ԩ��Ñk��:��� �EkU�3A��e���L�;���a"O^h�Gf�5.ڜ����"�A"O�X5,����e�b�D�l�Ω��"O���G�cfj0�L؞(��\�2"O��"g��g�`Ӂ��r�<�)�"O"%� ���S/f�s�IBy��ᢢ"Oz�C��l�N�p��l�P���"Or$��D�-ZԥS�-� ��<2�"O�4i!�<�ty�0�Q�/����"O�QyF�؟}�r!�%k�7KR�r"O�\�����@A
��|0�#"O���T�_G�X۰�֕Q���r"ODE�&Ŝ=�`��B�1E�lu��"OX�pQ�|z^�Џ@�s�,���"OA+D��+)$%Jg��>�����"O�ݱ`�
,�\��6���tq��"Oz���}�T���l�S���4"O��ƌ^�:���@<�@���"Oz=+q)�vMX�5�@(�D *&"O|��3��z��bJ�Ӻ�� �	�9@���!�0�ԩ~�6�O�,[�t���GL����Z�O�!�$X�(���G��:J
��	ݽ#�!��ƩD�Zdxa���tfT����@9!��-C>AX��� l�PHaՃ�^-!򤘠'�h�WM��|�e��cװ*5!򄞺%��A�D	'z(�z4�%*'!��s�,㧫�2!ǊL��o1!�DF<E���O*y�"\h�-Y�,�!���:CӾt����`�L��7�D��!�$h异�*e�V�R��$��=�ȓH]�aBB� )t��Yj��'�5��}㔅*A�&7���!F�R N[^���ii��AΈ��ޅс���w��X�ȓcC��ꀋ\�V�!)Ё��s��M��	S0H�&1���r%�������4�2+ۭ)ڀ4a���o<�(�ȓbYDA:C	X�#��(��b��U��9��G�ȳ`V�~��M��S�t�y�ȓ.�1&�^�4i�g��q=1�ȓo��MPG�	@�
h��]�쑄�ʒ�Ѓ:W�]ДE	 /H�ȓe6$%��D�*1s����#d�ɇ��J�V�$ ��JF�8b{�n�9p���2ʎ�J�k��'Ț���jI���#�b6%'B�ȓj!����'V�J����U�Hs��ȓ$��e���[�h|��B�>\�(��7��Ec�g@�aƔ���J
"��a��]@����d����pW�Ý�����c�x�[��U���*k�>4�\��Sq����LI�f(��ʑ�C9c2`��VM$]Ar�K�A�tZ2�+F���b�\�@$���"��& 
gݦ�ȓV<v�x��]p��Qb���ȓ	�-����K�Р��I�)��8���bO�l߶<�u$��md�ȓAhΘ����4s���Ň�Q'�!�ȓ(t\�8e�ڑ>o@��+2<L�l��[x�A��D�L�mӣ��豆ȓ��� t,��zf������̅�C�9�FfK	�����|0%��u	a��m/|%�q�0P�̅���$���J�`Ĥ}`&l'��T�ȓ/R��1!'I�Ah]X��>���S�? �	��ڊ��a���*I�T+�"Od8�M�����`��H�]�F"Of��0��n��U9�7���(�"O��1�ύ H��{��խ(�`aR`"OH�{�E�N�{�l`��"O����������ͅ/+�(q��"O��g%���j�eW"J�^��r"O��rC�h�dP���`�8�6"O��r���:�RH	-����pq�"O|Yh�BFK"|��"�ӄg��t��"O>��D�tx~Yٴ��R{�	�"O.��CE��,�u�a̓�qg� 
�"O�c�ϑ�@��]JDL�qKn� "O����!9[�eb`
H�7�� q"O�LRd'BT8QZ��	n��V"O��zWJ�|V��*�.-^����"O��7�ñGq�����Y�H�Q"O�� D�<' ���o�)|��t��"OM(T\ xL�1!t���,�vmQ"O��S�&��4jb� 5}���3�"OX]"�坺AO���gܐB���:�"O0q#��ɂ_����� _�����"O$���B���|���h�|H�"O�A��`͸;=�2�ł�<Y�iC�"O�� �,N�,���d� )J��5"O��C!ȳLw���d��g���#"O(�9֮Th���@��:|i�"Of����z_�)s�*��̱�"O���P�h肩�A�ʾ$�H��"Ob�Y��M�Q���2�H�?�6U��"O��z��ei�p�,�*}¼�ȡ"O��"���3��
�Y]҄Yp"O��)��E��(��L���\6"O@A���� y(А1�ŹG�z9""Ot���%�/��+�h��p�Z,6"O��8Ҍ�rN�(�
�>s���"On��'˅
���`5�P�����"O�;R	�2�1#�A�F�^8!A"O�B "��P��Ћ~H��@"OXus�J�}�<K3�	[񈰻�"O�d9���u�B�`�+#!���k$"OМ�@�(���K��
�܅3#"O��S"� a愒UKՆN����"O��c�k�f
�]�pJֱ,���b�"O^A�`�J��=Fd�(�<k""O�aD����@�^�@|p��"OBq5 ّnt���Kߥtq�iy�"O�2io�� ͒=�mbâ]!�y2�ɍa} Ф33`��j��>�yBɇ.M>x2��H7�P9`�eӼ�yB%H�Lc�`�����3��� ��y��A��Pq�%���4L�;ǈ���y2�Lx�I`�ceʰ2����y�
%,	�I37�×o=�A��&�yr`�"~�*1'Q�b�(��JK��y�.�Z>
����T�D�r9�S��yB�9�<��^�7���tΆ�y�$�1D{,�	/�43�)*&�'�y��	#.��5d�A��;n?�yR-�!���AuHZH'�`�B�
�yB�k$i�0�V�DD@3"˖�y"�'���kT��Nkڀ��4!�$X2	�'j.M��]��������'�����U
�(�h�LO��X����� ����V겡ᲁ�jnt"O^����S���IB��x"OT( ��d[��@Bf�&$��"ObA��ل��b%*T`���"O��l�NdR �2FM<*xr���"OvY���5c8���T�q�,y��"OL$%�|"u�!߳���s6S�F{����.G<r�8��B+m���%`α4!������I6 X�a�Ԯ�0k!!�N�>{e�PMؾz	,�Vn��~.!�G�>jƩ
�j�9���:p!�$�tԜu��c�2Mr2��4MQ�o`!�D��-D���KXI���m҃TU!���3#Y$z	ٴ�R�"6�_�=!�^)V��ɲV��#=�	sk�b!�"�@�Rc!�TFȠ�1ʚ�!�>%��" ��1�Hl�2�'��A;�IM�j���Pc�̖8��A@	�'�T��fٰ	n��>18J�3�'I�4C%Q(}�>�k��-W����']�Xը6W�d��W�M�	�'�Ƒ�J��)y���.�����'��!cO�A��$PE \8 ����{�� ZXI�P(��B��y���(~a��1�
S�L&���@���yr��8;f�#�Q�Dh.q� �^��yR��t���[ ʣi����4R�'�P����Q,2v=
�՗i�����'������X���BǩБqS���'�H�5��*V��p`�[lĪ�'�p4I4��.$%��K���V��T�<��	:�(0	�C�02��i �m�<���A�/����ņ��f;(-����E�<���_ �
�iaiY(#�UJ�
B�<�p��<W�(��`O�!���y�B�@�<�0]S�4���ؚ4�n䩒D�H�<Qs��,8Մ!�@�G ����Y�<A�f�FM�w-�:ך��"S�<IU�ӦZ�T$�Ō��L3����M�<��A��v��Ek!��&�5q3(E�<��ׁ0��	���e�4����C�<q5Ϙx_��w���3��hf�<����:*����`Ez2q�&A�E�<�2N�/p���t�F�Jp��[�@�<��եb�Xd᳧��H��;�)`�<��M�����U BSȊ�r�k�v�<��HK1����� s�"�� Z�<I�ρ�i�h����8c����gT�<b�J F�>�� 	�LX�At�<Ƀ�хpR)B�"F�J�)	�cLr�<I��4�-@b�	��yр�Bv�<��n�����F,B.d��Gv�<�Cnٔ7~�`j�`�%_�<�!0�p�<�ҍ^:r��V�$=�:����n�<i֋E YT¡��J	 �2ك�jf�<��<t�8:�+N���1�%�^�<a��w�`�I��,te��Lq�<�BK�򬽒s+ͤs�N��o�<Q����t�g��2h�]����l�<�rГ7=āZN��.AF�Q�h�<aF�X��$@R��F�D�i�n�h�<A�eS9%Ld���:VH�"��Y�<)�(= �t�"#�p���g�W�<��DCI0aH�!ͺ(��Z�o�Q�<� ��T��$j�hs�+ܒ1�"� �"Oq��*
6S@��R+�!"��6"Oh\x�U3����O�e�4��"Od1�#.Oe!P�ȋ"kX$��"Od"�J�J���!��~�a"OX�S`��1��DJSE��p���"O*p8��P�#-����ۢ6���0"O�� Fj�;���y�-E�x�����"O�]BP��1N�ƌ�	~���"OV񻐄�P4X���@a"� 	�'rȡ�J��ls��4�B�"�̊�'9R��;Pv�ySbS��N�`�'p D�D����y*#ʇ�P<��'u.:��L&},f(���@1"ۊ�
�'�xd��KJ(.��1�0G\��	�'�2�9�Iʙ=�.!���%J˂�a
�'��� k�k#~pg,��v�`
�'Sr�UfE�k.�CFK�tx t�
�'�fdhc>du8�0��ǖW):���'
�aHV)HIA�;SHH�����'>�#�%�-B��`�ץ<S��ʓAzThz!JC�$> %1`LϞ�ȓZ�����%�`���ź%���D;8��ꐝ.��)W�?]�r9�ȓy�t� � @�?   j   Ĵ���	��Z�tI
)ʜ�cd�<��k٥���qe�H�4��6]22<i�ʄI}�F�>A�,]��#��r��A�7-�M+3'��y"���<!�BA=&鸜:W�&��P�3H۔e��[�A�)r�������Z�FÆ z���r��*�4܁%�7��$\
46v�# EJ>��Չ'�� $ߓ��
�7T>�z�e�#`&��[��ׄ
-�#����/�'g�8�5�ZXP���U-ѯy�H���ގ` ���=��A-O�!�ɒy���H&ƾ��A�'�`%���~EJSh$$1�OX%N*��`�%�~�+��YM���RG���D�	k��b��
�}d�+�ՠǙfR6� �1K(\=
��B���(x�e&G��h���D���d.7cN�K�cM�O�����Ċ1��Ć�#,� ��!`{��"*4{�<�#<I��'�	�/���f ��9�#F(Q�X��7-^�O@ų��d(�Xh��F�.\@�)� ś�v0X�Ĝ�O��K�O�) �ϔ/c�l���K��8�r�W�p*C�	(N��Oj�aj�2-�����Rr��I��Cٞ�O�)#���ɰ�?�I��L(��$x"TB`t�[x�#<�c�0�$�
�����,F�r��K�)łl���ʵ�O^PAI<�G"G⟰�GN�1X���T%<#)����O�t:O��kRO�ܟL����M��SQ?�2��ec�G�v�p�P �G�]g�2�I
�ċ��>IRa�m�L�@C، �v��D^}"oBx�'E�Gx�e�i�-�W`ԕ�}#Ei"�y"�Um d  �y"�ݬ:&MS�b�87�D�CI���y"J��q �4
I�M�R�-�y���_^�H�/Z�'"q�g��'�y�o�"f�´HU�Ң.�537�P�yr�;���H�G$	�Å��y2 ҋB�8�����&f�����ybX?y�v��呄�8����y�O6eL�!�"�~BP:�Kέ�y��z������ds�͈�y���Bt,��a��`���@��R��y�k̢Kh��C��3X��#�+��yBlE�_q�X�+�
K\I")� �y��N�[�^@��G�1DFMB�o�2�y2HD'`��<{�dҷ,�B��2�T�y2W�]u6�с$�#�]�0� �y�WD>HɣG�ϴ����yNE;Nv��C�
�
�RC�V��yBF�� �LzdF�W��B��yB-��[� ����|�D9jҋ�y�O+p3�42C^� q*q�R!�yr��j���a�2X��p �4�y"O+��@b!�0��(�����y���<Ѥq �F_9i�&$��e���y"k j��l)f�Fc��MC�K�-�y��&P򩺴gH%[��YA�j�y2EǚInQzᩝgB^t�6Ɣ�y�gJ�F��ьv�f`��]��yre��F�H�"ŤM'$�NYҵ�@��y�B�8I�<����Fi�5�G#�y�i׹I8,%#qC���d:%	�y��F9K� -j%$�fd�!ʺ�y
� �x�k��E^&{p@�=F(�X'"O>�#�h�JC����)
zh�|��"O�,+o[�D��Ѹ�.Q;ZSZ�[p"O�|�O�1A�� �홨L?���%"O^�!�-�y]� Aި%���+1"O8�8t���su�Հ"�Q�j�pV"O�(�p�݋�sd�X@�$%8�"O$	;E�()4̤	��@8��P�"O��*�1��Q����Tn�X*G"O"�[��ԛz��y`N!J�%��"OFt[B֊~ܸ�A!�#���"On���]4s�ASB	W�\�18c"O�iV'�
^�ܸ���O�t��"Or�ɴn����51D.��AFu��"Of	9Ń]�2l�X�Ы�!W@$��"O��z�nU�YKl��o�kT�:G"O0�u�ƛd�Va�4��?d���"Oҙ��G¤_U���nPQ��s�"O,�9�B\;~i���.ŎW5���"O&�IW��:����L�0F.��:f"O0�"�(�'|�E���P�0�g"O�!�3*Y T+*�  ��7n��Tb�"O͡p�9%�\9�>(P�3�\|�<���J�"���kW�ԅ)�te��ds�<�uc[# *  �   M   Ĵ���	��Z cwIJ(ʜ�cd�<��k٥���qe�H�4��6_?><y�ʄd�V�k�,h"�l�A���օ�0267���հش=�D8�IBy2 ��E�@F�4mBԁ@�ϻU�,u���:$c �=�G�"�o�6�"eZ�p��7O�|�	3��
;2���<&f�J$a؏U�Ɂk*���Ȏ;q�I U Bd����:~�(��(�,{� .��O|p$)
�=��'�D��*ʟ?#�PȓNUoO���$DlPN�o�Z��ΓC���͡<q�O�e�P˩('ąm��6$>ax��L���p,O��*��J�)7�jC�䙲��Y�y!_3"���Ƈ,5PVN��yb"�w�'�L8Fx"c�J����f�q����w����#<�)T���%sp�����T2����&�W��O�)ێ��J���'�L��I�=f࢙R3#���:ͩ�461�"<���9�@�&9;��Ȕft��CV<�����O�H�� "<A!?A�͝] ��pON6$��s2�Ly�B�'����?9���JU�tȃ\��~t����2ܒ"<��a$�L4���H1*
�i��G�9kp��l\= �1O��	����1�ē:,�"vɉd
�yY� �%G, ��4NJ#<ف&6�[?Q�L��v<�k��o�z��%���\��P�l��O*Րg)"��'H*ם�f��`eύ$�R��Ʈp8��=	W�(�S��'�$�ޟ�B�kB���<���O �Ȋ�� �O����
��~�z0j�	Z�iR"O0�p�  �x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��     �  d  �  �+  �6  pB  �M  �W  	`  l  �v  �|  ,�  ��  ��  �  H�  ��  Ψ  �  Z�  ��  ��  A�  ��  ��  �  ��  ��  �  ��  � � 
! �/ �9 8@ zF �L N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'*7͑�X�-	�&z����g�8�Y8W�����4�����'�B�z�ZESt
^��D9��0$��'2�q+w�i��I�|��OP�q����t��$/襂Ц�/7:��<����3�';��hc3�_���4�Z`�-���i�		�yr�I�Ц�])	�ْ��F�%X�tC3��hv������`����ӻ_5�6�x�
f�p�H�	4ܕMZ�(�yB;O ����9ў�Sោ�H�?y��y�e�^m:���Ǉ~���'l�'��7��(�1O��P��j�������_������+�	�����Oj�Dk���'��8�vjM�r���R�J�Rd��O���Y��� 0�X��?)0��O~�
�'�	 r�i��β8�Q��ɧ<�)O��s���VF$hA��R�Ǘ�$�H�Mt�h;�4grX��' �6m;�i>�IG��!��M��䑲B��ZV�p�<��ğ|�I
V5ֱmX~2=���S�&�&��`��n�؅�!��Cy���Þ|�Q���ɟ���Ο�	��9���,#0胏I�[�@�(
RybDi��J��O����O���;�2@G�R4Fܪ�h\$,V<=�'�6m�증�L<ͧ���'	
���;(��2�l *g�ˇe�I�)Oj8�H؄�?�$�.�ĸ<ikט"�jЮ�I�v̹t	[�`ܴ�ĵI����AĘ���pw
��m`�qa��(͛��dQ}�*t�6�m��M��NI�p#B� �.��,�ڴ��lM�4�ua�4�y��'���2�?�z�Z� �S��5�C\4PNx�PCR7a�.ͱ*��y�'v��'���'"����'W�RGh�JJz��u �7&�B	�R�'���'ON7�\0CR��d�OR�nZS�I�Pzl� s��(O��r�I�H�4e����M���i����Ru{��:OR��R(�Nd;�j����x�N�N��]�V�A��R苐��O�ʓ�?����4�'���'�pr7G�	~�Z\2�b(% | z��'2�'֘}�E��I�0{�'���'��7-���9�h��@aȘ���d����1O����Y��D�O�6���kq��0ʧ�b���C�QIV��D��!���)���(�.��T���D9���?����'�r\$�L�q*�4�2x�%��r�y'�F̟��	ϟ�����b>��'Y6��tW*mr�bb�p��B�|$X��e�<�Q�i�O�p�'�6���#�}�΋p��IQb��o�Hl6�M�i���M۟'���w}�䟨X�)O荘 
�7_��ݻ�\v���!�1Or��?���?����?1����8�RLu�Q�L�3W��lz{�H�	����A�s��1���;k �z�8��@ڄ9���:��c��V#x�,�&���?��_j5oZ�<Y$I_��8��7S�:���D�<1��H�rN�d�����D�OX��S�-���惋�7D����Q6Z�N�D�O����O`�X�f��r�'��΋;��8��'���:qgF�g���|�A�>�ѵi�6�\Y�	�S.��F���0?���a�&�$�Iܟ�s���n�x !�WLyr�O��1�	�_q�&�&mb�qe�ԤM���y ����y���5����� p�%�aO�H��m�d%J��O$�Ӧa�?ͻ]r�,��N��}`{¾
�^�)o���l��G�PAo��<���2���/���,�͈PӼ�Y��.&��������$�O����O���Of��S-:��z`%�B����	Ȥ��˓M��6-۟O��`���'��]>�����SV&��£��6�\4��ayr�o�6�l���M3�����OM��NG�`κ]���\�g�UP�j5\v���["����Q�ɟ\�ǘ|BW�("��Z̈e ��6(.*X� #�O �m�"28�	�{�`��7��U��tI!+�V{��	6�M�"��>�ղipR7�������C�2�e/H;m`򵻂��3�f�m�<Y�ZWh�;d���lez*Ox�I��� ��x�a ?����.�x0�q=O����o��b�
� �(�(�ʓ�?��i Hɟ|$o�r��?w5$��d��"<'<�3'p���kO<�ig�7���j`��|�f�	ԟ�sw92��qB؋*Y��#�Q�zS��'.��%��'c��'<��'J��6`�+^�Ł CZ-)�xsf�')�Q�A�4�J|[���?����9��a��N����.�E �	���$�֦�4~���t�O�I�v���&qХSqoĚW�"�# ���h8�\�@ݽ��	�?eX��'��'�t�в2��P��UX��� .��0��ٟH�	ܟ�'sUbA�*O��nZ�+8����xdYq�V�y�I�C����՟d'��SRyR�i�p���E�"�Ԍ��a��&��l����ݦ�Aݴg�H4!�4�y�a?+P�@7D��?M�'�BR�ڙr�ց�`gU\AJ����qC^�d�	�(�I�P�	Ο��O4��C���4)�� &"7Uv$M���n�ĵ�f�OL�D�Od����Ʀ�] �^88bT�N^N�{�f�2���47㛖�3��S�0�7�v��F.`��5�EgŞc;�%s�u�� F��\{R[b�[y��'�"�U�(酪٦�U�B��eq� F$���'���'I�I��MKF��?A���?4�F[�T��t?hbB ���'&�6_���x���$��8���p��'�9$H�{B�O�$�=z�+�	�I�ʓ��2N�OH$���G��+h<f�u�>@bԈ0D�럠���`�	ş�F���'G�XcM��NI�����ޔZ���ڶ�'�*6�2:�ʓ���')ɧy�k�@̂���9�$)�!�yr�d�ČoZ�M�ĂV-�M��',2O�S��,��	�F9;�$��$����ؤC���5�|�V��G��F'7��P:�KݯXh�	'n�'���^��i�\xy"�'���8��Hוp�� �*]�-�$UzF�a}"�gӒmZ$���|��'��дx��,�(�Qp�M$Xkv��錩���6T�&]x��ܸ�T��F��{w��*�߀��0c�
(�s�70,��e��|��SW.��0cf(���XZr�F%dn0y��ER�Ol! b����⦇��FA��R�����Q*�^��4J����?���1(ڣ/�il�F+> ��gR!p;ue� ����c�%eEL�\���cQ��!���(�7j�,�ie��;		PP�\�
�
�I�h�i"�ǟ3Y5�/�-^��!�-��^`Tl��&���
8�6OV�]�Z<IE��ws����*��]��5Q���n������65���ǩ�Ӧy�An�:<��`��|
 �"������?qM>i���?	�AW}�Q���qP�T5yp��-P-P�O����O��D�<	��ҩ�O8�p Z{{d��E)�l�*oӌ�$�Oj��?9�fPm�|*M[�P�b�-cٴl��A��f�'nr\�TJ�,4��'�?)���'�	��P�T!g+������%�'8��'���Ҋ���'E��4hш! ���hܠ�dQ�=Z�nZqy�JN�$5$7-�a���'^��-2?y�W�/�D��5j�
,��S�������Q�cy�O�����36��Ж�6Ir��`T�*N��n�=�0���4�?��?A��l؉�����<�5�q��H��	ܴ	b�n�`��x�'��'���y��'�m���ɹ:�b��1e�16n�`�3�s���D�O���S�tvt&��������&��t)(�6LQ�q�'��B��Y�O����Op5����O����O�cBN�@z��ԏe�\Yѫ�צ��I����J<�'�?�����dN� �\�1���@�Z�(����	m���!�a1�	�L��ğ�'J�B$Ȋw>��/5U\|ʵAƾ�-O��D�O��Į<����?��$������6t�F�PhA(-�$�<I��?����d0-����'J^��,ւC�����BZR��'���'�Z������ᓃ�~����,]jTq�*I�j�f��BLn}��'w��'c�	!�Z�2H|R ,d[(����1���Yc�5
���'��'k�	?:��c?a'��:)7��4�ʱx�t(�E�~�D���O˓'� �������'��\c��-&���&0�B�%�jL���4���O���D�|�1���d�����r�Ru�A�<L�p���3�M�/O�tK�E��y2��<��M�'�Y��JL���@�HM>b���ܴ�?��Th��/O�S�?O��u(�5[�R�gS�z��e³�i(�!�f!|�h���O������'��S�C: �x�M�!{�|�s-ʇu<e��4y|88`(O<�d�Or��D�O:<@�&O�(��D�� ~nfQc�ʦ��I֟p�ɐH=� [I<�'�?Q��ݐ�CV�0�F�ڵ��
H�K�Q���I���Ӄ8�	�d�Ig?��C67� ��.�oӀ��'���	>g��A�'2�'��d�����It�|>��Б����	�S	v�8?���?�(O�dU��$,��e�G���O�q5�r#n�<9��?I����'(mM�� �p��V&Z���7c�dc�8��������O��$�<���=HV �O�L�YW�ԫvJPiҧ�'Yl�*�4�?1���?q�B�'Ԍ�DD���Mc��\&]#8[�)
L�R���SY}B�'ER[�����*t4A�O�.��3K��`l �s�f �B>w�6M�O�㟬�	�j��`v4�$߅~���ۄ]�y����Qf�z0�V�'��	ϟib����'4��O�б��(�&Ҽ˥�X8���#�/$�	��:�?� b��'E�.)�F���x�c�[*P�'�bkD��r�'�R�'N��Y��=� Z�12�"M�L�WC�
T�(y1P�l�ɧ$��\�`�6�)�Ө8Q����%B�S`,ړ�(7-��˜���O�˓��*O�i�O�]ka�^v}N��E�D 6G�t�1������T�D�b�"|��YZ	;e]20D�0b��h�����i���'C���n�i>�I���7�0r� �+7[��W�R(;X��(��D��mUx'>]���`����0���=-�h�)C� O˓
l
�+)O���O���&��=?Ɩ��c�)6E.xAo��P���L��TЅt~��'��Y����#(9�}XCI]Y�p�H���\���c&�Cy��'B�'�O���� %P�bd� ��t�J����R����J�9���ğ��I\y��'tZС�ҟ��s�NZ ۔��Ej,~�zu���i�R�'���$�O.4#��-K�V�O ��qF܋a�ECOI)����O��d�<a��8@p�s)�X��Xfz�O�c�������8����i\����O��*f�V�p��'D��+��H+ EE�ڴ���4�?),O�����-��ʧ�?�����2@4Ȩ@�kX'B� (��K	CC�O�ʓc7V�ExZw�t�8��D<+��a��زSș�Op�D�%����Oz���,O�U)?��]H%Zedr�c�n�\0�	zy2���O�O=
L����YP���a���e��qٴC-�<���?���?�����4����_ E�Z���5U7`Y��޲6�D��'�PTA����OfS��m[��q�dȋf	P�������ɞ__�u���$�'��O�{�D¿Q�@��qBG�]g�u�7(�O̓7L]Z�����'O��OH� ځ�|]`��[?�Q1�i�mQ8����p�	�=ٷ��=?�D��pH�!s��0���y}B��Z=�d��O����O��?��(��)�&HD�Ȩ-e��v��D�M*O���曖�'R�O��d�~P��2p%
�J��]�feX� Kd5�Ð|��	����IJy�'[xyP�ПB����S�I���#F�N�P��i(��'c��D�O0�����%o�&�րC:�5���l�xT����	��D�O �$�<��Z�Xy)�^���!L�H�HB�͞�Ёʓ�QT�lZџ �?!��S��̃���U≲ 8(D�GMJ�yFX�Sa�#>zd7M�O���?��J r�'���PP�u-˔f}�5"�,�o�BT쓇?�d�-S�d�<�O��p��!P�<�3���-�.���O���%����Oz���Oz�)�<��Ӹ]q�H�����{&��]�'���D0vE��y��$� �F��Ap��m��@2�IC#�M�3d��?i���?I����)O��O�5��Klx�3�3S�6�@1���y�bA�p��c�"|R�;jHH�g���D���5�l9�i�"�'�"dD�'1�i>y��ȟ���+ �@�����&t(�6E�O&܄A��ON""y&>Q�IɟT��r������ :5�����2��lڟ��S��\y��'`��'cqO9���R�QHQ�S���78���R��C ��!���?������OB���ʌ�d����s��[��(ah���ʓ�?���?9�2�'�1*�B8q��!���ܮP��%�&��$�*|��O����O"��?1��µ���?22�Q#m�:Eq��X�M����?	���'�b	D2Y�n�ܴe>�Y'l[�zCG[<�i��R���	ן��'2���$c�ߟp�� ��Yx]���ӧ,����h�?�M;����'�r��|`L�!H<u(�!�J�Y����H�KæU�I[y2�'$.�3�Q>9���0�S/��@i�K�DX��Alܾݾ�#�}��'����J֌Ә��i�+S�̬� �K!ռ5yB�2�	Ɵ$B�	������h�I�?5��u�T�<�@�	ׂ`*`9�	�$���O��!$��1�1O��v-C��E�Z\8C�B~�ܛ��i?J���')r�'�r�O��i>���)lJ�	j2��#0	HI��%ܳ+��ܴa6"l����V�S�O	�ɭW�n��5�<G#������w�^7-�O���O*4��<�'�?���~�g,�|S�n�%i�:���
� 8�8c��
��T���'�?)���~2�ʇ*I��X��)o�\� �i��M���k6�9�-O����Ol��4�I$9�K�XjX�P5�����7Z��k�HAn���������$�O�L�@+P<c�P��#�u.�Qa�(R&&� ��?Y��?��'O����K�`r�Tb���(ʂ�R`�җK�F���O����O(˓�?��߂���	KI|uq�f��TN�E�CW/�M����?�����'V2�BB.��ݴ@|�U��F���i0mK�S �M�'���'�Iȟ�+7��V���'"�\0䑨hj| �tgzT��lr�@�D/�Iȟ��FE��G�.Oб�ck2�\3�(G
+L]"V�i#X�\�	�,���O/�'�����)zV����;tiqPeR+,�b�P�I.m�����0�~�Lޑy(���%K^�8&!�#dAQ}��'gF�9��'R��'���O��i���cU�9��A�t���i�&�sDF�>9����{�N@\�S�
��(�u����.T���+p�Pxl�2C�\Kݴ�?����?����	|y2DA�<�-�!�fujQ&��,R�6���/�����d�(2#K=[13�n������i�"�'bB�������O��)� ����G��9�|��QaO"Mآ�ƹi�"W�(�C,l��?	��?��'��|I�bK������HA%9����'aH]@p �>�+O ���<�����O��Yc�	=	�*X��F[}��E�y"�'4r�'���'剽P.!� ��ݠ5�u�I�Z�F9���,����<y�����O����O&ȱ''R!��ȳKO� �>��\%1OL�D�On�d�<��BBB�)үR5 �)��ęD9�䑴(�VR��Z���I`y��'���'���0�'�j(��@2b\��uLQ�#`��&.j����O����O��jd�z�X?��I���ً����3�H�Z�d�$DP<�ش�?�(O&���O,�D�7P@�	c?�f);�)�ʾs������ɦ����D�'�V�`��~����?���i�8(" e�z����WoնyL�y0T���i��'�*a��O�����h�ol��yp-5Fgjɺ�.��M++O� XAK���I۟��I�?)��O�nW�Q��m ��]��]�gl#`V�&�'a�+�y�\����Aܧs� �O\ )=9�Sƞ,5�0m;&��ܴ�?����?!�'j���}yR�5 �֩�ZY(�����D8 ��$�ܴw��̓����O��h�^; �c!*�����)�C	!�M���?��H��,�X���'���OX���'=�R#��F��8�i��'�xI����OL���O���¬x��uZR��tp�l�v�ĦU�I����4�?���?!��>���{?����A۸��T���}����A}Bˉ��yr�'T��'���'V�	"�Z��LE ����%��<(БD�է��d�<����D�O���b�$��"�: aT!֢ϬBB��q f�eB�D�<��?�����d=!c��'_X͊���22\(qZB�7�b�liyR�'��I�8�	���1u{������O�9���R*tu�\���O��M���?����?a/O|��e)�z�t��5&�R�)q��ٍ~X������>�M������O����OT);O~�'<ѣ�%|��m���
dk�4�?i���N�*�8��O2�'��D�X�9�JˢD�z��p��V��?Y��?ygP�<qM>i�O�
ݘ�H�
�� ���M(w��Q��4��$ƌqn´oϟ��I�d�S&������ч�y�J=󒫐%7��)hb�i=2�'v\I"�'O�']q�laCF
ŅL��%��:A��B�iyP��`�c��D�OR�$�\y�'��	<R�R\�ԫ�b!�$.�:��[�4[��?�+O(�?��,JX�a���2J�v(��9�x�;�4�?���?A�OSd�	ry��'�d�A ��%�ŌaR��� H��IJ��'��I	y���)���?��A0�hs��l�ȹ�A�R�
�cA�ilcP�9/:���$�Oxʓ�?��_�ܕ���@��4iP�3��,�'1fQȚ'���'�B�'RX�x�&�$Kn J���]N6y	楞�q�2Q�O`ʓ�?�*Ob���O��ߟow�xI ,�%Z�f�/F8�2┟$�����	؟D�';d #@�u>u&��vT\ p���qGne÷�sӴ˓�?�*O����O��	u��ƌ��C�#Rp��EZ��E:!�i|2�'�"�'&�~��Ѫ�\��ƞpIW��o�y��n$K��-�i��\�\�	؟$�I�+&0��d�ć7x�(��ե�{��=�TBh��'�r_���$������O4�$�����,� B�0���m�-b�29�_8��'�"�'����y�|�՟p��J�k`��EH�w��!rd�iP�ɂn �h�4�?����?�'g��i�c�FM�B7v��E�C9�� �x�����OR�I�2O���yr�)��qd��p� Ұ-���zF*1����!M6M�OH�d�Or��VC}�R�`#3�O'$����"��k���P�� �MKg��<yJ>����'Ԑ0:�L6�$�5G�4C�bqRq�`���O���Kh+��'��Iϟ��k��,�6.ɊBf�q�C&^�L�oԟ �'�> ����i�O����O�,�4����|)Z�nM
*�H�W���u����MR�Oz˓�?,Ox���\����	�	�&/�.S�$���i�r�>�y��'���'~��'��	�~:��ue��C�L���C�w�T��fG���d�<�����D�Op��O|	ڔǓ�~��Ivό1P�0(!�Mښ;r��O����O��O���JtӁ6�RD"Pbх��� �뇐Oܩ�&�x�'�'&�'�쐋�'J���]�*a���R�Pi2�>1��?q���d��,�Д&>}��?C�H�d/Y<D�@1\ʚ6��OȒO����O�m����P��]y����1ӀNW�%��o��\�	xyBɝH��|���`U����>K���U�2{��H7�t��͟���C��]�	~�{ZB èd;��K�.��}7����K]�a�'D��a�wӨ�Oa��O�~�3d�jc��R�|	��ǫq��n�̟���*N4�}��Bܧy2q�dA�hq�E!Ql�>yn�?�.�*�4�?���?��' f�'�҉��LtW���X�	$�Rߴ3����䓦�	�<1���ҌKp̉1|�"�QP�΍�P)�²i7��'�F�E�^b�@��o?�rlYJ6ZC��
�oX!J��_�J{`�<����?1�eE��k7iܶ~��EN.9{�c'�i�ҧ�(#��O����O�Ok�8d�`|�0�T�VBN�3w �T�ɾZ��&�8�	�����yy��H$�=0R�.T�| X'�QR�;�0�	ܟ�$���Iܟ�)� r� � ��m1�	�IPx��!j��<I(O����O����d�2�Z�|�%-�,�RPہ�\�,t><���c}��'��|��'�Bi��yl��}Æ͔ �,�h��h�B��?Q���?i.O0��@Beⓟpj�Ha	A$M����.�	<\��ٴ�?L>���?�0���?)K�tHT���X["���_`0{�Bf�6�d�Of�f�� jf����'L�T�Ԟ��x�c�]6{��Cvn�<U
TO����O��:�9��BbE�8N���ء`ϗr�F�;�eʦ�'d�+e/�h��OE��O���6m�U�>�iAР�6sr�El�柴�� Y��z�Sܧ[BVrD-+.�*̢��߰0�oZ��m{ݴ�?����?��������a�8�ث�Ѓ^6���G��6�u�b���O`�S�O�b�	K��;P��!M�����У[��6��O\�$�Oh�
g�<!)��������f6�Ap�	N�V���b�*�		T9b�D�Iݟ�ɛ� 1�e��6Z�쀳"�M��	�4�?�6�I��?��CC����$�4���������aI�	�kt�J���25\�����H��؟���py�m,%��	A�$JԎ@d&)�Z�ǽ>��?����?����=6װ��E���Q�n4�2����\2��|��'���'��'�$���۟T��k�kS��t�Kd�*���i["�'���|2�'��*��|U�ݴ5�hA�-V�yd��3^���'��'�2�'Xr'��?H�ٟh�B�"pg��p���.��k��&�MS����?Y�� ҴT�"�@�	6cU����	?\��Va׌Oep6��O.���<I��ݱ^~��՟P�I�?��ca��2%�@�d�XV��U&.�M���W�}��Ov���*X��� �8e!��)�N4J�i��'���U�'�b�'C��Og��5���~6H ���Sj	Yp+ͮ�MK���?���^��X�<�~"tJ�"rˁ&c��2TG�>��6-&s����O����O���<�O �ln�[��� DN�(̥аf����`{6b�"|�������!PhtM^�s��x2�i�"�'�rJ_9�`c���i?ї�N�N��wo��j��(�b�X@�o�d�<q��?9��RP*��0{(pŁ+S�HbF�i��Q�V>O ��O��Ok�ܸE��IC�-*�tpu͛$'���+��b���	��t��ky2& �K�����nF+0ER�ʇ�����ĳT�(��Oj��,���Oh��L�NLv�y�g�/�P�1mI��8����Oz�D�O�$�O�Q����Ot�q5��&�0Y��NG)�yZ�,Ʀ����,�I��(�I�w��E�2����<h���!L�~��\�'��b���34�r"��k&XARO3�'r�R��E[�x�
�#�I�:K�\���Y;t��6�+�(=��ѐ=3��}�Ty)IQ�����I���-;��O�I��d���	m�D����&3�`�+�(2���U^g�����ʡ���4K�(�.7�y��Rx�x0 �a]�N�jX�⛊k�m��j 14�t��ǿ2�t|�0��#a���"6���Vٜ$�i�	5�v��%�[:4h����O����O�����f	�,{����c�Y�&�Ҳ�U W�N�����1��O�l�f��&If�x-��Lʖ�i�C�Z�pͻG�ȑn�,A�����J߬2!^��#�1s0TJ�ΪI���*c�'^�6mEFy�'���"��H�eVg�H����"�y��'|�}Rj�6!=��%��9�kU��O�PEz�O�2�G�U�,+��ُ;��B揓=V�r�'!��)�od���'��'����� ���#�,�vH\2_#�@�&���T�T��C�,��քͯX2�86L�?�=���#PY�p�6A�y�p���L&� :Z|���D
��
d�g�'d�� @����ЈE_�v��"�'N����?q���<��D�s&Ȱ���s!:B�+�I�<�Qf��U�ġbU��E��Y�H�b������2vg~�oڒkQ�!�Љ�f�P���Hz��l��ß<�	џt�W��ҟ|���|do�Oڐ�GU7a`(صdЎl�zSש� iؔ�Z� ��<�%/Ś^��\k�"B}� p����Q(6d	"�&1x�����<d	���ɋ|瀄K�'�es�h�vB��+o�xD{���'QP"�随 �����L��V��B�	�u>�{6oF�E�*���jJ(w�����Į<r�Ϣ���ʟX�OJ�`%��:��={�%A8�xG+�4V���']��Mݜ�b�l��>�27��O��-+c��{q�(yh�ӗg٬Hh�<	v����`Jr
��I&��G�����@{�X�{�¼w4,�L�["��<�"	ҟ(�Ip��L!R2O�[&:���cC<��͓��?���c&���܌V�
P+�+�s�H9I<�wD
�d"��s��a�	�DO�<���D�:w���<�O����3�'���'���K��� A֥k��'F?h���K��n斉�Q�j35�\��?�O@1��J�ehH� @�\NND�D	���`�f������H�;/Z`�_j>�NB�' c0��L��<�V��R$xa2`�O4�D(?%?�%�8��ɿs>���:Q(z�X�,D�� �\���('�
��K+`��U��3�HO�S�vRZT�HZh�r��(O�N��	�	��!!�,��Iß��Iԟ|�^w���'����ȱں��*\)�����'P��%�ؿg�
��� #O��!*��i��qbU-$H�!��O��AJ�Ħ�HSLCY8�0���6b4T�˔ed��s�������O���8����F�uT}Тzd�Ȱ��-i�!�DZ9�Ͳ�Y�LsE�44ZhDzʟ�˓���F�i>�:������ɗ��7b�qAp�'
��'�"k�*;r�'��i1��6M�O<8��%�8"CTja�5���'kphZ�tۀ��4���2���g�N����<�O��;1�')46�ܚh�>���ń�w�� B�8h�&�mZǟ��'5r��?��^�G�ū�`�/�(�%�<D�H��J�>_�}���]4m�0a��x�l�O��b�Yj �i^r�'n�S�:�a�ᣚ�pl�UA�D^U���YR@՟��I͟�I�ojp��<�OzЀ�)f1�&��/q�8Q�򄀈e
<	��{V&����(Q`$T�Ƥ@P�<�U�����40��F�'��+I]�)��A$J��'	 #����k�S��y2�Y���g���d5ʱ(Q�0>�єxR�J}��|#�珘�Q��y��P�6�O���|
�DS��?����?1ӥޝ{����1h	l�|��C;2a���i91O�3�R��JS�\�@$@��Ԛ%C�D��H1��O?���=Mv-�5��8ʆ����BP�����O��d=?�So��?�f�3P  ��&�A�VD�DYB���<1����>��H�)�t�k��,W��@����b�'��"=�OJ�� �%֑i��9�#(F�Wx��B4�'w�-��!�V)ze�'��'��f����ܟD��dYvz�xcp�
5�.iP�������#�Z;F��Ď�|��d �zNyQU��'XN���=4&vة �'
F�9�Y�x�͐/ҭN
Jܸ��'��a���'���,O4�d�<Qg���iMv��ŷJ,���G�<A@�ߋ2�&1�G�6\I<U�����{+��D�&�ٟ�'�+�z���G�!����
�
�hR�"ߟ\�Ißh���-ے���Ɵ��'+`l��Q�M�L
����@
I$]���ã �G8�PC�)�� ^t�nچz=� j#n�lI&9�ѥ	�#����&�2�~Ӯ����7T%�e���y@d�`�����	fy��'�O�S9Ua��S	��k9�=�a��y�C�ɮL���W`
�^��y�Vj��`��)��ģ<�a� N���'�2[>�sc�#]��'䀗 �)X5"W�u�F�	����tL�e 4K��o���:$�*S0�)���Ԣ�%�����G�D��
%�A�2)�Fh;c���R9�W	
1.�ԝ�O�lH�W�Q&Ij峖�þc��Z���5;��q�dn��$�O����X�69�I[֯�`F0�+��'�O?牮^�,�p�%�C����U�hd��_w��7���'%�93\X��T�x���	B���S���ş\�	Ɵ��*�\t��ȟ<�IR���I��%&l`�B'ܺ�H��E��{q V�b3IA
n��,��O�1�C�"�Bݠ����U�f���-��60.�I�cذZ�M�3[�<9s0�-�����aO*g̀���Q���
2����˕�W���ن��	^p�Ex���'���x!Ǆ�1�ra��7_���'���Z� �:G�.����Y��iJ��E���$�'b$͊�b�$����#a@�P,� �'2�U5z�=��'f��'��A`���ڟ�h���?*�h�x�l��:&i��G��`hf䋪vJ�A�퉽(�hC�B�P��L �+ϊ4�	�?g��cMh؞�2+а�X=F�#5J�Q;pOP�Lk�U�A�4�����O$�'�<i D�t�H��Ł����ȓql`yXR��.<�b�9c �Db���0�I�tP�L�B)Ժ�Mcnܢ.��Q3��.��PS�O��?���?q�u�5��?y�O�d�ZDK#��ֈ��C�(��q��Z�l�v�@��p>y��%0� ��4x4<Tj�iIDyz�D�F����%.��ͦ�B���1�8��&S�O^PǨ��M#����$�O���''U���a�l�KL�DFl	& 4D����o��qo�m�a+��#$~�B�mp��O��$Ű(��Q���I{��B�18���C�Ж7	�8¥i�$3� C�'��'��1�Eˉ*9� �T f�T>�GR�py3Eh��>65p��)��B����vڨ�2d���8>��ᐬE�?%� �γ8>�yEI��XRf���(=���}��	�M����@jJp��Z7ys@i�E���O���䄀���0��	1t��)�-�N�a|R+2�� 2���_t�"l�禖
^�.� ?O�%j�.�Ӧ��I�4�O�: p��'���'@vX�S&��k��ء2h,_�p��;	�8!�.���E�u��W9������Ͽ��H��V�R�r㩊��B	X@ ұߞm
�-�>�`�H���2c"����&g�RC�n�/������t	J�_�^a��@�x������L�r���O���?UE���@	y ���"<j|���M�0��̓�?�
�_����U&F��$E>4��Dxr�?ғ��� %��1��`��h�Z��#�b��O�!�g���Z:`�D�O���OH��;�?���LAb� �MR;1�8x�*�<��K�>1�%'�|]�,��	�!�V�	Q�,+����.=D��	U��)b�D9d���ɻ��u�@H�1����	�T����l ��������t�'C�T�0:E�
;j�S��1:T��Is�"D��E�Վ,g�����X�d��A���HOBʧ��Ӽ�C�*K�Zԁ6aV+^�t��.�w�<᧋�#�xY��_?Y��
�[�<	,�7+�t�k�`ڔ�<���m�<9 ��.)��ӑr��49��b�<)�B�h�.�@�j[���8�a�<�G�Lȡ0���h�=Ků�[�<1��V�	d@���җku��
�@U�<����)�0��U�@�B�/H�<��iN�U���DB�Y�N<B�C�h�<�B��V�jkB� iܞA���X�<�`Mp�)��/�O�2d�Q�T�<�pd��
�dh��`v�.RG�<qf'ش9'��ȴ͓�������<Y�h��X��=�Ua&�6E�Q}�<!tK�>��
�~��}�w��x�<P��>P5Ĭ[�@C0�و-�u�<Ƀ��#;��\�E�K�h���,	��C�I�	�ٰ�C؝"�H�f��	~�*B� OxvM�ah�nU�����Y�6C��/y	6t�"��&G�^�AEL�2$C�	n�9����LI$e��B䉬2��b�(u�J��5��3��B�ɎDv݀w�B�)?�ea��
�9*$C�I;K��0:C���y)��ŉ`��B�	Nk<4x�п.,��@T�X%�B�I6/�p�t��'G��c�'�E`�B��q��d�΅�x�,����u�PB��&"qT��r�6!�h��=z�TB��9em���0�C�/��0
P4�C䉵X��DI0��>(�RhS�iN:b�LC��B�V�Bȗz0j�%F}flB�	�9~�,�,ة=�^��0.D"<��C䉿b&~l�Œ�JU����,rC�O�t�f
�M<u頥X'*vB�	54�������)6&˗V�+�XB�5[������E�`�QB���W�>Y�ď�;\e�%	V}�)����%)/�|�;��IS��ȸ0�푆r�%��R;�HyU���9Г�t7��]�$�Ihn) ��
z/�4@�ȋG��OԐqAHڊr�dm1��!0�,	���'RV�� c��u��CcA�4�ȹ.buAp�̵	��L8��(t:�!v)F7D�]�T�ܤ0�{"��M�&�&GJ�yR�S�!ʉ��D��0s�J#�R�WG�<㵡ĄB��P�0J:E;�D(�hB��Ebp-�8}��E��"O!��Q�]N������W�(1��� "l� 4��ʫ86�p;E:O ���|�G�D��;6�|a)���fF��gà+\��v|`���]qh<X�cI	d�D�{R �<��ǁ!����Aśc�� ����x��ρ,�v�"�I,=�ظ�+ˈ�0<���0�r�#��:�V%�cH);�0WāF�<�#ɓ�Y+<��5k14��c��C��=9��T0�>�@���H�9���Y~�LJ�T����w�ı"	�%[�d��''��:w�O^pI��ڽK�^%�焆�{���'~�d�!�Q*g��Q�l׀�l-��O\6Yb�p21�f-H��נ�~*���ꆍ��	x�¸RJ�hV��B��gO�ąҜ�B���P�l"?�B
��FUX�B��%<�,L��-ٽ.��(ԅ�k?9biڔ+A�TCr U�j�L Kb���L��_d�P�=� ��(���!M�Oh�xZʜ�ҨO^AB���>2Qt���N��% ��h�BS���+	w9� ��f�05sA�#81�r�	�Oj8cB CW�<���~ʟ"@S����`RHJ-1�i	���à*���b��@$(Jx� d�<�h��+���iJ5-����D�߂�)A��X�r�Uі!
���,���2�~��9O*���
�~W��q��'Lqt$�F�B
8,���s͝�]�qO哭����Y��"��p�p&��]���͓Uhp�i���O�B��a�,�Q-���։�$5�������7Z:�s1�	p���u(�j&�i>��EY��M�v�\�R���u�يf�:�zt��)wȢ>)a㐪��jb�C�g��]X�VT!�&�>2�a��BS�le04Fx��'�ʍ����`��O�05��fU�l㰑X��C�gd`�����*e��'O�����;(��B�eR��qJ�{�'��p�,��M��9(��D�hA����h�$�O�E�	''�t9j�O�YYg�>a�*��lĖ����9c����ç:F*�X�Bd��[�ȑ�>�{�'a�\� �!I������-{h���'���� ��t�^ݰ���}�'a�]�t��()���zď[�e\X!�#�/��	��HO�ӌ|���k�48�U��DKL�zaQGh�lwD��7 !�ʹ��`�6�Ճ/�OW�@�MV�`c@G�b��:��!�{ܓ��I�";��X�'E����� o
5��l��K#�Ek��<M+"9XR�Ҭ,U�ɱ9VEp��T�٪����(-��ȹ0J̜Ye���ME'w��(a�ڌkS�)�DT�;V"nތr�\؁����J��O�hՊ��xSD�	%`^��l��_�-�DĻ��O���3�	�i�`%��Z�@fְ�̙!3�$WB%p7�܄ N�	�Ǔ,�pL1f*��
US�*Y2<���ʦ�4#&"\���@Uy���NuHEYw�hY'�)An����L������u���N̡IZ@ҷn�?
�q1��:3�LO-��j��<y4"H	L���O֘�`�`ik���VG`�x��]"u�sta˅�0<9��;o���m��K�.M����(�V��%2�BmA'mB�x�h�_*0S�xʪ6DA@"*M�mh�L�Oi���B1m��P!��!$	 F�>�FH^�BID�-�8X*��Iz�E��`0p7��p�Kٞm�Cw�{��Z(w�����)O��Xq�ªt�N�2a��Vպ��5�i�n]Z�&�)�LpŢJ0��q-O��y�e�.4� 8�iG�k��[���-d�v���I�h' wMP��$O���1��8H��OJl�	�g	���s�`����kA$dʧ�10���D�#��(�s�
�1'���o��$aJ�H�>�IlZ~�I�d� E�ɸS�xxó��.H0�K"�>�
¶K������bc~d�&I]f�'v���e�2*Fb1c��ȸ_�HP�aOh[��C�L��;���*���}r�*@�]dJi��'����C)�NX�|��\�R����	�5D��
�3?��a+�����	�O�\��W�l?�F]��E�w^��iY4P]Ȕ!���yRƦDy�-aF�N/Hmeh#IFHU`mH���2&Th���>O䔀V��@�vd���w	<����J�Ut��R��bhX��'�@�ؒ˟9?�d�b�ΰ6��Zc̽My�-[Zm�f`=�3�I.Pn|(�)�r��(�E?WT��֧Br�#�	�R�t�u�0�j� �;R
�8��l)ƌ�d��yө�C%�fdӦ��>�`�� ��)�F�Ѻ<\65�B��Nf\�a�"/d���mC�n�d	�' �V)�ĊШ�5�(OeZE�ڱK�l�S8�h���'� �Ng2� A,�=k�$ 	iɖI5�)��$	>L�H
4Húe�ș ���u��ň��$K$����9�?	��Q�A�d	P<=�)���@�'�x���	P"<�"��v�zaQ�O&5Z2��Q8ݸac :7d���b[�SLa*�˽{���wO�9+�&4X6�$�.��M p
O����i%*4����$F����P�{fp��I��<!t*]���aJܴ����4Ĕ ��֟M��YE�b�P��@�/���
�p�$�D�ڣ3����h{���AB�<y�	9o fp�5�ݯX��F�ҳ���d'xs��̻B@Dm���#7T.٪��<�̈́�I-0����oG$��%�ᆋ$B`�P��%F/�z8�O \�I"b�H�$� �ߑ�z���Q��-V2o@z:�_ f�8*��-�H�6oS/I�<T�">*P�1����ΰp$mߤ�x�e�=ˆ��>IX\Kԯ��T0 �eǯLh�I�V��� �]?��r��_2VW��K�O>ld����� $�;��Ş$\��Q@F�>Wl,C�b@�C�^�IA�d�����0`�����X0h*Y&��i��.�� 2���E֡��i��af��d_�@�$�#F�o��}	�MI����2Or4���ܕ	̄ф�O���'�$��߭+1kC��� ��"B(����>�OF!]4*~ƴ�1�"6Y�@w��<��t�O@-/b~	"�O~�+��O<��O�����=�jx�C �hv�a)�.=p%߂�����d��`S�a��,Cz�J|8��Z�E���,�2ܓ�D��3և;R��8H���	��鎤eZ!��`��~�s�(RnA>v�ޔBa�]�RD�"��be�!g�\P��$i�@ i�l�I6Nޕ@e�M�����Z԰�f�.��q߿M����U-+�f��$O�P����p�ފM�Z�?� ��(1YRK0:8�KPc�O@�l�a8� �C��@�f���X,"<9�<c�&D�J�&G|T�gT�S[ �1
��T�R�U�S0�� H���H�)rYB��{�<����$��`��	�9<�!)�!�?���ѓaX�uf�\�6�F�^�81�y�M	D���!�`Ơ'��MH2�O�"yr���E�X��AE�w. ���#�6;�h�(�F�T�{c
�+|�bL�煖�"�j�#��)�<�����6��,ֿ|��l0`�.�*�c��qMb���"�@�F�ӈ�9�$����>m¼���'�>R�lex�C�,=,��"��j���a��F��$�?A2ū2��M��)��B#��I��] d�P�(��ɔ�x+0�	���Χ�?�O�f�K l�^>���#ڸr�Nu󐡝va �9�����y���/6� �;�wݎ��Ņ�{7U*ӪF�]���I��X���s�'-j��C̾t՞��E��7T(ג�d*L�~)��Iɖ.B� h����O����D0z�P2냲m݄�C�$�|��˛Q�"]�  +F�"��ǵY���[ ÷z���h�~]E�DX��+�/E��v�ӓT�|=b���"~RU�	!g><K���fm\�}r�'��@��ƪ!K��!�L������Q+$�n�69Uzޅ�%�
;.џ�Je��pH,e
�U�	p��D�������B� �^���*
t�֝A?�O"8�F"�#d�A+l
5Z(��A#?=��a��a �A�xB�,|�!��k�%��J�0v�0U'��*�
Y�8����OT��DH����%��d��D%���^I  C��/N�(��D�3ݱO�%B�\�x$�A�G<8x:��:�T�6�2��Ai :��� ��X�P�j�%�X����-b@n����	�<ӪO(9����$�G�+��a��p-����'N�bz5��6N�~�F���O U�c:
��Y�|��ժ��ĳ��=Edl���ǑN	\���	)5l��VB��^�^�������<�P�&�!�DH�!�>m���4�sݱ�S��0`�\K��?u[�l�GD��:s�,bЮ��ǓMv�i��o�9E��`�
Q i�*|&�T(��a�P���G� $��yb��z��<h X���ˆQ��@
Srrp9�O�"aD�r ��T/FE�>a�.ū\�E�u���a���`�L���۾FU ��T���w��`�H�d~2��7on���(μ�iP��?��'��`iD�MP�w'��=�HX b�"�dQIU�4�r��'���O��������<P�Пrֲ�qgh-)|�X&�#%�
�+c%876ѐÓ
Z$%aS"��}�QR��n9��MR2v�b��U@��[�0�
��O��'8
	�v��!��|�0X�#��3R� � ���G�<���@� u� ��K%����e��aj��!n�5"t՚�l�c��H�1����Ɣ'��ѱ��b>I�.#�*� N�.RzX�9��R4��O�P\� (���B)3H�c�0�4�;��8  oq�<o\�a�f��g�>�����1�O`�:1/��'V�`S(��<���Q�fޘP�i��L~ T�v��!!t�e�	��O)���D��mHC��M`�̝�lm��J��R�]��3P@�$N�H�Ү�T	ay��J��hc!�@�y!})�đ#9˪�x�!�R��ړ���VA�韤�PѠž�?	fP�Dk��:�7K��B�t��l[�v0�y2C��t��d��h���Y`b��P$�(Cq@���f�<�ՊR�<"�1�'�Fӧ�s�<!r�
�6�n�I���H�����v�,��x��Q�k,�Q��/Q�l"`�J?Y�C �nu8I[�bW� �tcP ����J��¨P�|nZ=R���Q$�M���O� !
A+�� ��1s	őGd���P4��7P{D�Y���0`� �\��h�C����	q$	�>��W�]��$B
Ǔ�h���g	�����g2� �H��F��1K4�O�� ���Y�pB�O:\�%������$c��27%à���0=��JB�[�`��;)_���#޴5䄩�Q)�m��O��##DMl��XyJ~nZ=Oh�2'O�1"�Iu��:%[t���Yq �8r�V�=	
�W�6T��U�ȓn\L���n!SlC�@
�\��(�F�<�5��h�Fd˔�4y�=�e�,D�|+�n�'�P]�-�-,��)t+D��B�ڥh�q�9~����n'D�\p^
li�T{� �z���A0���X�B�I3�0�܀��[��yB%UD��U���~!4���$�"�y�	_�4��8��G�nY(�v�ޜ�yRo�h���M5�P1����.�y�D_~T�fb�?�
��ͅ�yҦǛA�����#�<�{�냬�yn+X6
1��%ӟr�Z��F�-�y��C�7˞��dA:u���iӜ�y�W.��Dz֩Ĭ[8t)"C�0�y¨�9�f�Yn@Z"��)�gG��y�J��,e�d�"6i�7�T�y�d)�l���D����1�v"O\4�rh�;Z�hEk�aU�`�P�"O����<e28��^�T�z B�"O� �lJgM��b�&��fmˍJ��"O���!����v�a�L0(�2���"O��#�E@�1��T��ʔ��l�3"O�x8���Z���8���G��%"O>U+@���sǘ���"O��B&�8�2L�#�,����p"O��Z��)Xt���'DRT��d"O��c��Z�����
z��X%"O&�HB���RL�UK�.�/$���B�"O���cˎ�s����G *��W"Oι:�R�o�n�UN�o�
DR"O�d#�Y�Hղ��%;$"O�(R#��-�P@2M�Z2@��"O.��skOp��������t�+�"Ol�D���n���@)@5Zp�Lcg"O�9�n_�i�>�B0��OHlxad"O�cP'Q����Y^��P'"ONy退J�K�lh�1G�B�i�"OrE�s
E�U��=�����"O�b�F*k�Ȼ���1&�p�k�"Oj1��ӛ��l#�J���0�B"O�A��i�4{)�yn��FR��"O�eAG�׆�n�S4�Mn@p"O��l�M� �pJ�>d$���c"O[0!�
Hh� �� �a"On9k�F��4h��]F��"O����ƿO�-y�&H g�xmz�"O$���/Eh:y��Kߑ��@P�"O���w��z%����i�v �"O\�AȒZǠ��/��E�,U!�"O)���L�	�S�ߴOYr�P"Ovdذ�MX�N@�'�_%'K��;5"Oj��t���P/�ᡥ��U�ؒ�"O<�A�֐=����qO��E�&i�"O>�ʕ�C�UxPhGN��}��ܠU"Ol��W��'��QF!a��A`r"O�$��ODR�����|^0QT"O�	�g�<]���bfC�,c��"O+J�;��r�����D�5�!�\L�e�ĩB: ��+�,���!�D"T]��G˩� (qƁ�!��T�<&D8���6a�� zb���!�䓐!�=�`I~�΄�I�!򄎅*�h�&NJ4�3b��J�!򄚧�%��J�b��Jҹ�!�d�NB�	e��Z���Vb�>!��ܕ)h ��C�C#$y�`ѐ�!��B!r�,�)�@]�	"p@PB�C�!�H9�-�B*�*#V�[G/A�j�!�d̮>��հ�GЀF�"�-.@p!�X���v��zZ<+q�!�!��/��������9���y�!򄐃Z�trQz���Y��!��Wi8d8y��1W�v�#��H�!�$X��j���aД-�nM*�i��N�!�s���i�d9.�U���v�!�Q�o��p���
✤��DT#�!�10\&�ʳ�"l��%����!�d�<@X�qt(	�6�Lr��ؿb�!�$��-��s���m�VX�7h]!�dé$+�Tc���=bg4uIW�ʗCC!�T�9�D�P���&f6���Y�!򄄢#\m�W%V�$d�K�BY��!�$�YX|�E��d�Y��Y�!�� DQ�k>��� v�{�nD��"OB�s�·y�5�Uo��2|�i�"O�Q�PC��I�yX�2 ?l�:�"O�](��f%���"�'\( d��"O���Ae;V�Iq�M�%M�20�!"O��x0�Z�XX��^�����"O`R�(-����U���
�d��S"OVm�0��'�p�V-È�4��u"O�4"��Q,D�H`Ȱ
��U��"O|�z�JL7V-B ���..`��"OlXad����y!p������T�x�MGG�8$�g�U����'$��ҡ!e]���#ԉLH��ѥjTd�<�#C@^���"�%%6`�����L�<) gҽS B�ّl��A"���G�<V��9���8����L���̝\̓�hO1�̘����Tr����!��!%nib�"O�٨"��F���k�^&D+*|!�"O�4�A��@t�MB��ͿZ%��(�"O����M�0N>�H��Є0b͘!"O��t�N;$�9�,��X��C�"OB<0(W�n &%��k� ��Y���'�S�<1���g`1n���
vʞ�A��C�I���a�3�
9WL��"I�8-jC�	�x��]�b@	��X�W-��RyBC䉋%���Q3ĺj����ۊ�C�I)Pt$dk7M�"������rH�B�	>L��%���P϶��E[6DC�ɃQ���Ҁ.�'I]����oد"��B��m&�F�N)iS���⭔
����>�т7Dh^1��#��Z7r�[��S�<�t�V�*W��@�Q�*����H��~2�Ts�O�t%���"���+ah�Ru�t��'��
�aϠ�>ٛ���K�iIS�)��<� �R�$�5-�¬��mA@q�ȓ5d��/
$/�$��D���Ԁ�ȓ1j<K�,]c�6|�U�ٸj��4���@?1�"#_v@Z7�:{B�`⣕z�<)Cc�cR�3qAI�R��=�GW~�<�SK4TW���#�MɌ-���p�<��fE�V����lG��b*�W�<��`D�t4K���Z�h2gΟT�<���NX��7B�#0qJ���E�<��N�6����KLy\f��d���<QP�K ���C���N��LZ��X|�<Q҄Q�I<-c�@��I�� ���B�<91ȹ\wvq���V�d�D	�B�@�<Y�nH_��*�˅�3P��hf�u�<��o�57P��3��Ҏ2��`P�V����;Cx�D��(t���M	�t'�D�<ߓS�,p�숬#�D�a�A]�h݄�d1���L�q�2\�@'Fx6��ȓ&��)�%¿k�vH(��Y�X�!��j�6�� L߈U�Z� �޵\�هȓ%�H���S:�3$���_���ȓ|kh$J �ϓ>;���V��a踍��!l��ʲ��[3p"l��@Rs�<aF���:&x���eU:*���ffq�<	�f[�.�DɋtD^�1��I6̙t�<��C�&�JE�1�J���ek�n�o�<��H e*�a��	��Q��i�<)��	+i"P �A�$՚�B�N�<q%�5[���ڄ玶1�r�`EM�<��oH%x�n�����/]���kOH�<� j9�@"�|����L��M#
%"O��+���\�F%IwJ��q�"O%H�$��^�"�3��XN&.�X"Ox��D;�I�)P���K�"O�I����CqF��R��@�"O�#c�
�p����r�z06"Ofai1HE�gH�e����y��x�"O0��7�N]���s¨�b�X��Q"O��[�Ǎ{�d@c��7uG�@�"O^8 ���q(�t���/wU��f�����ɱ$�aRꈐLT����6e��d,�X�b O�d!�e��7��	��$D�x0dG�;�0q��[�Zr&}�t�7D�`+E�*?WrL�&��h�V89w�6D�h(��!��d;v�X�!�8���'D��	�fj`�Z�bհj��k��&D��zA$X2&�JS�)�1۞��u�?D���ĢM��A�b�ϛ �H��& D���2(��&����+��!v��h3D����#3t�ր;b͵=d�P��3D�x�ЅV,Nxh0�I�x��A�<D��`CY�`̒x�tl	�'�@y��K>D�p�ԀL��6�B�`�z�!��:D��x祅��4��0��E��A+D��ڶ��5:��2dG�.��H�7o(D���$�[�Sh�C(F%E�J��,1��蟚�Ӱ�Q�$"Q��g�����@�"OHMۓ�@�cele���ҸC*����"OP}���M-r]l���k�&i��K�'���"q�N/@_���AS�.1�=�'�t{p�%!0�r�5��p��'6�dr�!�)ZH��B
	�d��D��'�b�ғ���*"�س�ֶq�L���'��YB�E;VX5pn��j�1��'�
�R��PW=�(AJ@��'�8Ԙ&N�'��ق*L�%����'���P󣖛�bR��7.C:|(5O��OM/U*��
$AA1YZ�$(\On����ȦY-�xR��ށbU��&"O��zU�D���%E�9����"O�pZaˆh2���A�����:6"O���A&R�g�����[=i��h�Н|B�)�S/5u�R���I� ف@��J��B��	h�0�23�(}i�t�Ħ\�N�C�E/��g`ȺS6Ь+�B��=�&B�I,0�a�lK�h�����+=WB�ɂD(�eBc���L��9�B�	,{BA��dE�h@���3�Ƞ��B䉚�B���Z�s��٣���y0�B䉊�t%�`� 6� �" 
�onlB�	�B�t�Q��N�U�B�Ksi�%i�2B䉄߾t��Ur:Ԡ�P?\�B�	�׾,B1MIlX�!Q҃ə&B���@���7Q�9�"F+k�(C�ɶG�@��%mG!)�VzcI	�j�B��#R� �!����,��dH,�B䉧9[U��S�@���G#M�B�I7p�闂��?�.�����*�>B�ɄYXB7C1k:����'�0B�.���B��ոwqܐJ��[�B�IA=֔q*��EĶlʥ�^?&��C䉿8�n�W�J,�D���_�[�C��Qw��Ul\�et�네@6Zw�C�	&O�N�1��B�,A��@ +VC�)� t�kR�ɪ=����.�]|��"O��zCg5Xc2qitMK�G�y�T"Od�p�M+aj8yc��:rq��"O>�YZE߮X�j�d�x��e�WZ�<�R��4�Б`�] \�:�su�]�<��\#�
����I=U49�DC�B�<���l��4�b�I<>�2��J�h�<I㋓�:�� 1Ť�>1�h  aƍf�<��O�b���d�"z�dQ�DZ�<9A�Ӭ{�p`��P�a��5��c]K�<Y�LR�:\�p��9�r`+7��F�<��Ԍg� �c��̋P�����̈B�<�b���M������_�!���D�X�<�G����]���\�+v�X�D��T�<)�.�;g"[�
�%;�Z(���S�<A�bq��� J:����S-�O�<�d�8*�bXc�G�
� �0�ZQ�<�W�0%�dx�l³��'�̋T;!򄚕tR���$�W�|�q�̷m�!򤌩$��yѪ�͌�+g̮8�!�� =�`��iL/1��U�B&͙#v!�D;Y�̽)����LI�$�ȟ$ �!�ĕ~Pd�e��>i�M��,P"]�!��%i`�*��U�`j�0� L�=!��<ɘ�r��O�@Z���`Y�:!���|m�͒�j��L�F�ϻ` !���Jx��!ϙz����T�E�H!�޷*�B	�co��i��B#@�!�I�~H%��F�-}Ƥ�{	ٶw�!�$��g2�-�����H�@��燇Z�!�$��l-�C�˥��Q��f�7j�!�P	=a���E[�8��Ht�7E}!����un�up��N��p(��*Sq!�փ�F�㰊� $||r"l�'!!򤆅y|��b�G	CI��kƋI�q!�$_�9V.��Q&�|V��JkC�b�!��.C Di�%c��kO(8��B�G�!�D)��Ӷ� R5� sR�Q�Py2������X�N���RC�	�yb� ?d��]Z��K�g�X��W��y�g[�*���6�ʲ\!ҝB����yB�]�al��Z�R�&��ׇ�y��W�d�"��iW� 	��(#�
.�yrHR�0;�m@����p��Ym���y�枷��e�%ժnX����^��y§�$�`��D����ia*�9�y�拉'��0�O�9�@�k`� �yR�U�ة���:%lִ��U��yB��fC�\���\3à�X'���y�̿DmޡX��!��i��� �yb$��1��(���P�h_�yrh�	'P:��֩�:3R�0E%��yr�Rf�t��/N7s�@e�E��yBoۢzgJ1qR�̥:�X�"�(�'�PyR�f�ʄ�U$3�`HR!��V�<a�JQ�`�D���bXa���S�<)nT�).X]ѣ�Դz���`��Y�<��鋣��(��lA&&L�(bp�T�<���]����&УO	x2��T�<��DΎq��ǭ���5�QNT�<i� L�V$3�,�5���h lUj�<q�뗳R(�c�9�V��DB�f�<) b�%Z~���gK5~���I2Cf�<�e�Q�a�d؉��. Ԏ\�v�PI�<� E�4��?�,�@�lP=5���"O������Z� �?�j'"O��S� R��x��#F��	��u³"O���-T�c���� wƄ�xd"O`�f#�q@�P��_H֕�"O>d�'j��E>�$P"�T�<d����"O���7F�I��+բ�!��h�"Ot�aF$�=X�J����_�2���CQ"O�uX@.�M\<cg G@�$aA�"O�eiЭ],gn��4��6`���"O�u��\�t�H�y��q��x;�"O�JRl� ?���m�/2$	�U"O���~������Z�4-l�#"Ola�sl�$n
!�%N7�E"O������9-~�1Q)�4Y�p�"O*x���?c����Ӝ>�x�"OB\�B�0�"�S$��,)�6Uك"O�YG(@;B~����AAs���f"O�ݑ�M�|,�P Ӓ�ɘ��y"�.D}d��b�w.0��&oݻ�y�dF�,
t2��N�]pΑ��(�y���Z��%D]�I��!zF���y"�Z�-�4�{��HP������V��yR�0lLa�%޶|fzm��	J7�y�.�2y�le@�	�r�r�[>�y"��`� ���}ZZ0+��yb�J&@4�s�f��#rv-Q0,���yҩ���tq�q�'��U`+�	�y��wNZ 0�
Q������_5�yba�	{�|�$j�.3ҀA�n��yr�B�E���"�E�(gߔA��1�yr�Y�a �A�"�Q�5��y�2�y2千dp�<k��^�.	�3A'�.�yRM�4N�u����d������yB#܊	_Z�&�L�~T-(qN���yr���uA�������6u�`c��yrb\�)�bIh�mR�H��ٲ�o�y�+)�B�ǈR9���Ղ�y��H�L/���˂,8����kR;�y���'>�� ��I�)^J5zdCЁ�y�(��
�0��E�2yż�B�o�y&U~*�͊�)�6g�$�#��0�yҎJ�Cҭ�B���t����R���y�e=}����Ď�t6r��7����y�/"K���2�?`���ڂ�!�y���4�L%�h
�X�����ջ�y2�V_N��P�T'P�4,���S��y��\'R���f۸{�l��g��yBno��X��V�\�T��W��y�M��84�xA��Za��*�W��y҈��*����$/��J/��y%��yҫ�$�j�!m�;�0�s�\*�yr�����b�7�|�"� �ybE^�!Q^1{q�0O�U�A��.�y�aұ%C��B�U�.EB	�g[��y��ȍ|��b��|I
x��R �y�*�!Fm�!I2z��!����yRaM�N��#�%���Pgަ�y2��!w��& �̞�ȡ�ʭ�y"��-gL*�8ᯔ�M*�����y�¿O	��1���=�6X�5� �yDI#[�%��#��	��+υ�y���{ ��	�
 �ȁ$�M�yb�E�e6֔)A�I�^F5{�ş��y
� �m� ֳ�	�J�=�R�k�"O�,�7��k�L4��X�o���"Oތ��,��~x�D��"O��ض"O�u��C�,�ٚ�K�"����"O
�F�E3t�B�k�m�E�J!b�"O����_�'z�LC��,�6U{�"O��panԽ	2���B+�i�W"O4X����,55R5W��Z�B1H�"O�8�un��J�A�S�F6���R�"Or����<n��b��AFn<�"Oj���\ ��,P��A��S�"O������p�H}ie���?��@G"O:�`�ɂ�xy�#!@4����"O�݁��B�G.�E�5�՘�lPS"O��!�%
�m��#U'bx��"Oȥ#$cK<M�Q�C�քlb����"O�`H7�,� �I�En�Q�"O
�ȗ���]��A�w��Fȴ"O���gW�H!�ų��#	0��ا"O `�4�P={?�����"'LPI�"O��P�)M(^:�,��cъG�@�3"O�=�V,�&V_�4g$͢ Sdс"O^�+��Da;b�k��!?�T�q"O6��e�C 2l���APԹ"Ov��5�Λ9"L�BK��H[�"On��©	 `����B�Vh!0"O&�:a�E�0�0r-�e����"OΝ��g�d�� ���Ā5��$kS"O�r��MT��,u�`�Gn ��y2��+m�ȵ >F��ږ�̰�y�kUo4;��R *�.�f����yr�ûbݞY�#D R��a��7�yB�"3��p���њP$݋Я�$�y"fR0��0@�[�F[ �2a��1�y↚�*���O�72��S���yrhN*3>�����{�tY��I���y��L=�l�cP�:�b�K�)�yb�ϊhncS+S$b�Vyq�ɒ/�y�jPM!�(*fiՎYȲQ�tg���y�
e�%��G���|4퀩�y��8���1�����ɰ/��y��oD�1@F�1
6@s��y"B�d�
�ӕ��u�0`�gA��y2�[�[��d��h��o4(A����y�+�H�#U��m�6ܛCJ\�y���L\t($m�TK��#M��yR�Q)Ob ���$�(]�P	���yR�+@�d��Tc�T�s��y�#��k�̨�֩��,���B�')D�,�e*�=J>��M�@��A '4D���4��i���3&U�Gvx`V�1D�$��Z.u%`�cd� �8q+D���n���ڳN�<��$�g�-D�x*Vk؇�]�$��ARta��&D�4h��N*!���ؗ�C�j�W$D�TH$��+�n{ �7��,[�4D����h��X�f��d!r�6D��`t��~r�y��Ζ#Y��*��6D��!��'y�U��ē�2�nz@�4D� g&��<)r�N�lf^ �A�2D����fـnD����
/8�8�n3D��`N�
�y��ݯlR\�Rv+%D���+ިWM9����J�<�a�"D���@h["B۰#T<p��,D�� l)r�韷z}x;���C��0Xu"O���fA<{q�a)�͋�l�����"O^�
�N\&J��A�͍� �\�G"O�� Ѩ]�qMv���/p�x�9�"O<�6n�{��0i*��%����F"O`�����b� d3f�.{���"O
ʆ�\78�2���I�V�;�"O\�V�[�^�qC�T�����"Oҹzq��4.���E�Q���Y�2"O3����/,81��Σ0���S�"O�|A�B��T�v���ܪ���"O֝"@���*\����0Ҽ�*�"O�%�� D�|(qdۣ^҂Ę�"O:��t��=��(�d��Y�"OTXg��6�X���,Y����B"OF9�A�� 1� �A)SG��8�"O�!���|w�P���ӎR�<Q��"O(#S��*A�̡Ӧ�Ts�j�"O�D)bU���f^I葯R�f:!��B�ʔ	P��2e̫���@Z!��O�(�=ôj׾7/B)Y�iǦj?!��>p�����!�>�� bC	�7m!�Døh���r���:Mʌp��
#!���w�$��@�4eK��%��f!�$_5�P��G�o�6��'�\�r�!�d�9p��	��͖�`�1%W1TW!�^!'lZ$墂�v�I�T�T�!�dQ>C�X)�aHU	7t�h1�/=!��G�%�6�T�,d@@�J�#�Py�GW�CW����Z)uY�����M�y"��!G����dF�m��h"��N��yB�J�$�0����dAPu)d&J��yb��U�k���X��m��g��y��/M`��T��7J��$�̎�y�×���i�<�� ��_"�y�WJaB��4�Ӊ5Y"�6%F��y�.^�<��Pn�8,�d���Z��y��W1��KN�=��<`C���y��%J�܉�e�р
��Hs�d�!�yr'�t��ehQ	�J`����#*�y�����h$�)D� ����"�y�Z�� [w��e<�8��C�y"�-(�P�[��ێs~bPuI��y�ѣhҦM�w*O����K�#� �y�S+���茙��-S"�[
�y2�q�Qc��b��@�eV��y��u
Y3�!�%�i��iȺ�y�$^.)r�y��%EP��,��oъ�yr�0(������	b��B��y�
�R
h����%>�2o��y2Ԇwn,1c�ŵ��2+ܖ�y�(�	it��噚N�%�t�H�y2!'��3�o�I�Z��ì�#�y�$�+϶J�D�:�Iʂ�T��yb�48�頌�;C��PZ�d�1�y��B��&\8�B�A�8�H��-�y���fa���GU�4cW����yrW�p4t�����U``��y��C�t�%��H�	�v�c���yBo��F�Lh�wK�6.�J�����y�!/s��s��7-D�\iń��y�c}��h�HY�~���y��&��ť���r���J�y�!	Gm�`@f��!r��!2����y
� �����3#Z�!��0�y��"O�ɀ1A��=��t!�+C.(-�!"ON4S
�hΉy�KŹX�,���"OBl3"�̥M8��A�؅e�����"O�q��!ެ�M�1)�s�|H"�"O�����Z����	U�]5█��C�Ʉ%.���;Z����)�B�ɑ,�R��k�+O�IkpI�RGB䉇��u�ƌY���1g�M�օ<D���S`��/����+̃s�����7D������!��]��r���L7D��X����Z6&�O��H%p
4D�����G/`)�:T E
� �0D����AޠSWD�b�T�\��+D���4L7�!��
�K>�C�$D���@�Շ9�n�ن�Q�Z(t��-D�ؐ��F*�T!KAǛ:b&@ې�*D��p��A�9dqI"mGgk��Kr�%D� a��8g��|���B5^l�����>D�X@�f�1��Ct��̕`'D��a�.��J��b�=<��T{�%D�I���s��l�3�]!�,ɥ�/D�tkc�ݧK���S&�Z+?�Ě`�0D�,��[EN���%\y�iM9D�(��B�77���Aś$���t�;D�\�"�� 2���xfL֡Y �U��;D��q�Sr��|Y�dɡ+����r7D� 1�jЩF&D\��!d��QZ��"D�\�U���d�aBK�(c�k� -D��@RH�&z����(_��3cd*D����(3�����ޓ:-V��)*D���vk�&ULL����.�H18�*D�4�բ3Gv�@�˪%�����N5D��y�B 8�� x�l�74�A��i?D���` <iH��Hf˱�̍�T=D�`�sχ"[�t�kt'�/QQ��q�-D�8؂k��5�ؔ�"I�z▁ra&D�Hې+ȶ:�����C�d�N�h��#D�(�d͒�1}�YQ��@V�i.!D�$5�6<����(#�MH��<D�H�3!�`�&�qH���A�'�7D���͑�/v� � ǆ�B>�i��7D���q�^�y��y��>(�r����4D���u���A"<б�?���S�1D��)3=0h��`�.
����/D��C��:6��'B�l�|��vC"D����τY�m��B�'$FR0 �>D��i—J/�u�A*��ZN��5�;D�8Jfc�b=�q��"���&��td;D���hJ�\$8�%�ܞ3�:�iE9D�D�S^j�l�D���6d�r�$7D�����4� �c�mX�B_i ��6D�@P��T�1�z��Ui�,���я9D��s��Jt��=��@���)�&6D�@)ɞ�rs��Nǟ��Ibb3D�<i�g�u�U��+=�!ɔ1D������>���o�jB"噐�.D�ؓ��݅��9��/L�`") D��A�a%}'D�Hc�-GZ԰�>D��x��[�!p��� �(\�0,d(/D�ܹ�4#�b�C'�"W�θ�P�(D��R�V�X�,��!�E�D����(D�(8�gN:�HE"�{T^�G�3D���Ɖ��^�!�	�`���`�5D�� H1j��y����`��<�<	�"OFlC�Ƙ?�f=�Cc�+����"O�ن�ۄ-��a��!N��@�"O�,Q
�v`2�+��'$�(y��"OVy[��!�q��Hz�pI�r"O~�3� ��j�W��,���{�"OD��gK'��Ź㊈+W���""O�@ң� <n]k�� �#k��+c"O��.U�_�V��h�8���0"Of�Xd�� �D`�G� ;.�Ѓ"On�y�h&R"�Y8�)ׁ:��a�"O\�t���3똝c7)Ӄro�MQ�"OF(�`ʓ��\�:�F�Qf\��"ODt0M��p|�g�ޱdz���"OPy��4�r��C@R1nn���"O�=ГiS�7�n�2u�ϗDt xT"O"�aF�:|�x��V��!�9["O�q ��n�ӆ� 3[XR�"OT�qf[���4`���E�q�"O�i���T,N5�c�U��b-rC"O����@/�)�.E�N�`��$"O�<BQN�a�b[7�M�ڰ��6"O:���KȕV(
U"�*���6"OJ�"��T#tbܛ�_dΊ�"#"O�eMW�L�$��[0o�R�i�"O,p���.w�x�[n��E��Ѱ"O��PЪ� �ڭq������"Od�7M���9ـM��_�\"Ot�KF�Tdp!��K��t�""O2ԑ�ޯB��hE��h"Ox�"j�;�J4�*~Ol=�"O���d)Nc����/HGM����"O^�(��F�Ӣ�� D�|�"Ot)1��{��k�X�JA"$��"O� ���\�v��e�W��0hUyC"O�D��D 2��ȃ�	Q�U�����"O��jL��\�DJ�ΐ��J�j�"Ovlb���E�X��6ϛ�y�R"On�{0��*�%���3%e���R"O��Q&�.Hj<P���j�<�P"O^}+w�J/l��T�2��\ˁ"O�@����@�䵪�f� w��d˦"OEz O[2B�l��5��6�"x�"OPa�gꐾB!\!�Z�o��h@"O�*���%�B�+ � y�"O���1���$5�R�M�I�|��"O�����*r�L�� �@?���""O.qq�؄3�\t)Ђ*&`L��"O���@�U�h��س�hL�m3�E� "O4�
ׄ�9��(�ؠ%:Prp"O���T-H � �)r���"Op��.a���RO�5*~�hv!ɨ�yҧZ 2T�D��zO��&���y"隅g8]Q�'K3g�f-��.ڮ�yR���1�pN�.ڠ!!,�y���)(hs�I��ϊ��wKQ3�y�	�,?��Ui�
�����7�*�y�oH�e7z[��ʱ�����O�`�<�3��0�R�pU�@��j����d�<��@+�p�%J�}صy��u�<Y1��� FR�8�!�_���Z��n�<1��Ng��iJ���=]*t��h�<��(�����a$�2bh�qMPy�<��̟�*��=0�A��Bcd�9U"�~�<� �9p���9[$&Y���]�&"O(�a!.
�j�֝����Kļ䃒"O�h���\�~�$�S0�ه�z|"T"O��9�k��:+�iV�ֱ7�ޙJe"O��5�{������J;`~'"OT W�н<ry�"Lr4��q"OZ�(���>m����bAK ~�8���"O�8J����mS��H�.m䈲"O���i�h�����e��
�"O<-���@�r�R�M ��Lp�!�$A�~�T y�A��@ @Q4� J!�d�<�FI2� �c��b!��!�G�3h�x��M@�m�b�Ѧ^�Rs!��_�����=m�����i�!��T�r���݀+���CQ�L��!�_�����Δ�}��!�LܥG-!�T�` ��1���L�DYCa�@!J!�D�M{�i��A1�0%�sA�?!�=y��!�����Y�E!�@��!��X����q�é/�t��)�6!��hZ��Vᓃb_&��!0!��ӛW�@cUΗ<2���c�J�`'!�Y��i����	u9�eѠ+��!�$����;$W7m�R` �Q;b!�d�oHkëڨ[%2��Î �!��ĉI7�M��/ەY�e(thƒ'?!���>T����.��S�z�:��*U+!�$�
�2��BJG2O�v�Acٍ$!�dZ(_\���S��}����l�!�$�����L�o#�,{��"1l!�����G�؀Z��Q�E33!�d�D��q-S�l1�3$�1!�D�+"p������{z�+���nC!��ʅ�a@(9~��éXz�XL��|rt�"bȍ��9��F}x��ȓ	�RIm��d����� rb��)%x�� #N��X��"�Z�n��0��[� c���m�0�a��1d�l���/]6�k1nK��F$ʧ�X?�M��'�d��3*��Б M��-BZU�ȓ/U(2��I�r9�%H
$jl�5��n.�I頃��zɞ����1�NU�ȓG>�CQk�2&Rz�� X0�V��ȓ*��-s�N�&/�ְ3奂��B��Ɠ^�P(�@�� (H9)tϓE7�����hO?*��#X_����#̳h�vq"Ԉ�I�<Q��%N��]��.W(��b�{�<��_ʒ��+)!�  o�y�<	����}��@�"|�[UǛ]�<d�>	�f@��N�q�X �G$�]�<�T�H�h��E�u웗" ��`�Z�<���_-e�.5`��G�
$��X�<9�,�9Oژ��Ӷ=��[E��K�<YB"�6xNT���T�I�N��̈}�<	��,GR8J"��lx&����{�<Y"�
R�����	=n<�UydI�O�<�+���h�h���?E�a��YH�<��9�& #�L�[Z4Q�(��y���g���d��O�����K�7�y��<:�Ȁ�2B�F�
�y ���y�."1�����ˮ?aDEYN�yB�LX���	���+0���y���y�m��m�dH1�D�-�Ҩ��䞘�y����
���	���\�H�L���y
� nd���I�M���vDܮBkj8��"O�YX7ϊRjX��Wb�	, :u�"O�ѠW�;��#�� �0ٲ�"OH�
$�
�Q���n�2E"O�hm�.��c��@��Ts�"Ol� �f]�W��U���ڸpk�"O�Ր����.u�!��1��)��"O)�aM�U���	�8��KuO�H��	��k@vQ9�nA/@l� !��OXC�I<��IyFB�.C�T���h�(�C�ɑ<` ����ݺcȔiuM\-J2�C�	A��U�e+�g;n���E�C�I�s����D���u�x�Ǧ�VKrC�?T��	�_L��Պq�л��B�Iz�Y�!Ԓj{H,���0~��B�	'�\�����>p��qU�E??�C��e,��K% E]Ȳ������VB䉽`?4�I�G�8E��PaC6XjB�9d���J�N��yb�P{$(�*V�C䉇>����%1�f�cW+�<+�xC�I�jD)���L]2���̊16dC��:08�$
�3LpN�9�ߘ�C�ɯk��hcʚ/� ��\�B��C䉻+����L0L����O� L��C�	Jd�P��m�
fn�9r��)�^C䉊[܀I�jE&\�H|YJ�,�VC�I�r,¸9e�� �j�"S�X4i�TC�	,�||��JY��R�[�DDS�C䉤
&"uh .�B(|���Bǝ~g\C��0ɢ��
��: \X`���9(&C�	�_�ٻ��|$�X�d+��C��	o�`�dK�~��I>_C�C�	<W,ԫ#��-�R�7�ِto|C��_�m�r)͍	�>������_�rC�I� �,!Ѭ�9ֵI��B'Q,XC��n�z%�Z��ջ��L�D�>C㉏0���)��:Y���r���k��A��3�Nq�fM�a�~)%�b,ԡ��0�aH�1~� �p&EP	����ȓ��:� I�*�V
���d�ȓ\�ʠC�_�P	!VL��K��ȓ �PA�������84��>:l�ȓ:��8S���o��"q�ޭp���E�`;d�Q����tX<�,��IWy2�'�ў�OЀ9b'݉@�t0��J�H5J�'��aHAJ��Wy�T��h�%��'�1ZV��8Q�}�cP58��թ
�'Q��`fX=^�±��i�$:���h	�'t"X�@.�4������Ȩ3��AZ	�'�`�cf�@�	_������/*��	�'��1�Rǃ7l`dq �ȗ8a,���'�V�!�ӕRS&�:�A�-/�TA"�'l�}���� RfֱI��R� ��'��UZ��(2�h6!]<O�9*�'
��p�=^�h��A�>�P��'�v�"��J�D�S&:����0D�hb�R5����nO�m�´�� *D�`�ҫ��`~.uJ �o�� �M&D����!ғ5�
A8�t���d"D���RG�� �tKf��v4ف.D�ds�,�6m�IH�Hw?z��!�9D��%-�	u��M�ҥT�M\��6D�xY$*M�5#<$(2�U�_0�=c�h7D��e��9���Ţ�RӦ� ��4D��  I�pE
>1>u$I�Ϭ�"O��ⵊޠN�!	N-M�h�0d"O� !�֓AD�` ��Ր?���1"Ox�X��)�h�33 �)�2\x�"OԤӴ��&8���
�,Q�|��%"O��C� ��5�Jyq���<Ur�"O�<J��<\2$��M�±��"O$!�f�X�v�<I�@΅�'�AK&"O�B1#3J>Չ.m�^�#�O$@�iП~K��"���.�]QĊ�OB�$8�O�X���ER�XagG%5f���"O���JQ�HJ�h�B��"O��*C ��9�<���@�*!X�"O�)"/��By���5�6,��|�1"O0x���۝u2� �J�D�ީ"%"O*8�V�G?mL�-蠈��.�ͫ�"O`ҧ�x����$Ж�r���ޙ*��'��(�e�D[�\�!!G�$��hK�'.���$�"^�� ����40!�	b�']�ظ�Λ���2�gŋ&QB�(�'bP9A�&��m�C������
�'%�Pdl�y�L��Gה�ȹ�	�'j��[rΟ��@���M�	����'
n��tC܂C��Aрi�V&��	�'��pE�=Ӯ<�F@�P��x��'�4�A$`���hR�@`���'�QI���^4�]�!�]�"��}�
�'�>(���,(z �H�H�8�
�'l���@/3FLV<0�/��
�'�Y����&a,̑���G�V<��':�� �V�z����L�9aFLQ�'L���f�ډS�~�X�%��o�<1��J�7�$y[V ժ��|y���m�<!0��KF�Iy�1"5h���U�<a�nȮ ʔ�8T�.WPp,S��S�<���G�lI0�"@�,�Z{�Ef�<���޹ �jy0��̠;�d���L�<i��i?$��2�uMb �7F�K�<��і{� )��X�w����f�n�<A�DP29E��;�D8y.
p�\b�<Y��Q�<,(��b�;f�1%G�s�<9Ԇ$u��A�P�Z6Y!��I�<�%��UFqx�*y ��`eg�B�<�3��4QU[� N q_��Q�V|�<�2�U�I�(M���Y�H�8�0�
m�<�1HhSlx�M�UlAЁ�j�<��Zb��h��D�:+�:Xy�cD�<��9]=�lX���@W��pcc�<1G
�17H�a�b��fH$a�%�x�<y��wyL�LDO1t̀ң�[�<I��N/[/:<����&���趥�O�<��B��q@f|�c�Ӱb�͊���d�<�`6���5��,r� �c�<Y����U�&O0r�q�u˒v�<y十�a�"4��c��:�d��-�p�<q'��E�i��P5�2��k�<��ߊo�\��QE�-n��Icϙg�<�LEHZN%STe�e`PP��`�<D�	�&�f��'D�ꨈ�g�V�<�wI8y.0mB) x��3�,�^�<����#f�Y2�%� uFdy���P�<�dg�4&D0ء�f�� s�8;D��I�<ɢ�Gy���ũźcǀAfJB�<a��3a�0�x�J�ck�r�'�G�<� �!�GaP�9&��L�~i%S�"O�]�w�$,�jr)	"78Hbv"O�d���n��9�3l����"O�(j��wj�8�p	اn��ʢ"OhM�,�5Ҏ� e6�	K&"O@X3Q��3i��A���,-�5�"O��QU�\�d(�c��[+R�[1"OJ���^r�er�E�*bP�@"O�	 (@P�|�RD��i�U�S"O�M�&4h>��"����j�c�"O�Q�g�>E�T$0Q�$,ƞt[�"O|dD��I�Lqa��	
�d@�"O�$pe ��z��cȲ�ec�"Oj�	S@�!oE�d����S�"�"O$0ӕ_�Q�,���A�:���#"O�$��bӥA��t:�C��M\P-�"O&09A	�.,�*x�s,X�NWt5"Op��S(��0��4ۖ�ơ.1ʘ�"O��򦍊!0 �P�*#��"Op
 `C�����ݼ�U�3"O���E�8+��r�L(CTl�Q"O�mjRE��|h��k�2+�,�G"O�Q���R$Y����JػL���"O4�!��)bK0X���ȒG��Вg"O �+�3}�,�ABU�s�822"O�IS�a��A�����&[y��!"O�Q�w'7gS��C
�0r��"O��JD�E)r��-[�� �0�8Z�"OH�fG��e�� G�_?]HP:f"OY�p���wO�	x�<P����"O��O�b��x9�c3C��bd"O�a	�JE�b�RH���f^N�I�"O����@W
s8ы�+M�U��pF"O�y�(���Qr�	ܳ�����"OD����hi�m��۽�:E�w"OzѨ�蘹}<�bc��R;dQ�"O����G�@�p����9&��K�"O �q1N @i�4�F7.����4"O�]�A�
^�rdI��;�"O:1��5;_*�Z�#�E��8�"O6��C�8��xa��Q��*��"O���4���R%��`]�?�T(�1"ONȳ��U�K�НwO�00���A�"O�]�v�RSd��g�!�n�"O@���?^>D��+�	[�N8ч"OH��çY�<�0��I��HXq"O 0� �T�>�1�PT�R�h�"O
�P HW� �9�1"��a`���7"O6����ù#�6-G�bH��4"O(=�����$�8�S�ϐ�L0$dY!"O`P[��K�rPQ�E�V�@ ���"O��K2�T�0FH*������f"O\${ i1�:�"o\$y�"O\Is�,�y]Tqp��_��a��"O"u1M+iJ�P��T7�4<��"O|`���L��m�&=�HtЄ"O23�)S$S�U�Pl�w��]X"OT��t͋?��H�?�6$�"OP��V`]�
�|�2���"7�$�3"O��Kg@P(m�ѳԉ�H��%��"O��ꡪL�p��"3F�0<���u"O2�3q*��� +ۍS��!g"O<Y�$?:���BJ�GP!7"O�Qd�EeZ�|r)�Q9=�B"O� r=���җfb��g��5�3�"O��e��#y�&M)4�]-Z
�iw"O�\�ek�<T&L�DG�oL��W"Ou�!M��6��RG�<SSp�K�"O�0s�V#Y�u1�b�O�Z��p"O�� s�0W($����d�rqp�"O��!c�2�tD�'C�"�l�B�"O�����;w����U��~q��"Of5$��=R��S�^�Hz,!�B"O�9U.��l�$C&�Phpf+!�!��U�*�B����v=����4t!��@_in�'��^��y�`N,iT!��7~�s�ID6O��Y�"��!�$�	��)GI�L��P�$6n�!�[oP�Uу=&��H�c�9u�!�$ہ(�HQH���nyS��)�!�Ę<F��bL�S�5 g�ЮVr!��M�w~Y*Ѫ\�.j���ּvJ!�dL�s.~Ye��5d��hz�L�!�$�M��x�å�'�(#��Z�* !�$T�WV�(��Z1^}v��d �BI!򤌌h��"0��.���OB!�DA7�qi���SRq�A�ӱ Y!��e�� 3P�"<	8-av�ȴ9!�D�_D1
�#��M�0X��B&8�!�䎓�~��cb�?_��{�FP�v�!��2F�.�z�GTB萡#S�+6c!򤄺G����O�%Um
�c$@�	U!����Ǫ6�<�tC�9)F�� �"O���iVW&��K�k�	f=����"O�0)�S�B��C��p�.���#6D�����)_*e��+ -�d���j4D��2�M�~��٪��=izC=D�̒d�I�.� ��E.z�9��:D����K/-*L�9�j�&}9�w�9D���ߚH�
%-�4> 	9�9D����W�I����O� 9Ɛx�1D���a��;��ѣ�ΚZ���c�.D�h���[n%fK�G�~-+Є.D�8G��m^J��%(q4m��I2D�ء�j�*V���d�E67"eप+D��{fӛK,U0W�޹9�2��#6D��7H;9VH�s7G�]�"��5�8D�T���Ԥ!i�=2����@���Q�)D��&
Ԭ+߂ݰ`�15�Ĝ�-)D�3��*s����K1�� �ƃ&D��a�iB�m�u�r�� X:�8�%D�{P�
�T����� ����1i7D�̂rJL�ETΩ���&/�4lk��4D� *���芰�Y�"�p��K4D�8����(������LD��:v&?D����~�h-Yb�2g��(�M"D�ܣU���2�$��@J1��E�-D����B
h��-������k��+D�A�P�HЉ�^6^#���p�6D�p�Q��	ި�Za��$.:����%5D�H�wk]�
����O2��1�4D��@G��ɰP�#*��Z�d��6D�8�q.�l�nH��Յ\,����9D�(��� y�����R�j�J�`!4D�DbRc��%�V<��І�ju��L6D�4`v'ą�1��~(��� �?D�H�g[�!m(��ǡb�X�$ ?D�8�Cf��q r���

04��:�>D�� L�ie("#e6 �CqV\3�"O���!�"��"���FD�S"Oؼ
�_62�$t��aQ5I���q�"O޸�%�-u����/@8<�Bah""O��K3�Ԩ5��$��*<ԡ�@"OZqQ�B���jы�d�	'<8���"O\�Rr)�Yj��e�8@�b�"O�]a��_�QK�X�B,lA$"Oj��)H�H�-��◂�ޘ2e"O����L�.����T�X�@�p"O$e*�N�9J�.�Pd�: #Z�JT"O�ȆV9*�dz��H)h�"O����d��h��kF�)���!"O���̉b�5jRa��#ɂ2!"OPԑU�,���Χ(�`��"O��b��+�-�=l>\(�"O�3��e/$�+Ϙ�*m(�"O�(2���5<\|���U,)��1'"OV��3F��K���P
�y�Hq��"Ox�*���,���c7*�
h��4��"O"��` ��O.����G&Ɔ��"O�1��S�G�LQ[ n��
�X�1"O.�I� Ê y����5�N��r"O�I�S���OGBU�R�
#�(�R"O�a���{�4@�C
����"O*E�W�@@���n�(��@r�"O`���#1@�7k��s�p��"Oj�#�_�v��go��<m�|�C"O�}@"c�2Q�@y�Eў/�	�"OZQ�%��f����#�<Mu���"O.�{G(�j�#P�6X��[%"Ox�����%(r~]�5OB*@����'"O��E�Ζ3��8�N%�8\8�"OV�{`l�1���Ɣ*nn�x�"O�d���!91�p���@Y��V"O$EAKWJ:1�#)ƴb���w"O���#'
�c9&u�wH�`��"OV�"fQu+2dG 7b�U�"Or�sdUn�T}��E�;[���"O<|�d�X�3�P�Iu��XkB�;r"O�ФM�Kv�$*�9[,�G"Of�r׬
�;h��S��)Gg@H�"O�i�O�c�j����+�F@Ju"O��d�.���`���y��"O�e�U��P1f1J��� o��a�"O���p�/�R���*��Ps�"O%Q��5P�@yEƚ+J�$m�"O� �wǓ�x� Q1�ĝ�ؼ��"O�=1�l�b�����I�6���"Of��?�����,+B�9!c�<�Eb�yhN�*$�T)a�C�<��
�|�F,J�D�T�b�P�!XD�<A$�_-J�ӐH�_t
ipw�N}�<IEDU[�Y����xg�Ux�Ax�<�Ł��҈�� G��+`8l�PIO�<� L7#@%:�^�{�ia@�G�<9��U"N�B���r_r�8BjS~�<a�ePaF|�J'9�1AdD�r�<��!�?/�Ȫ�X-]���91�n�<1��^�H����N3T9S�h�<Q&?Z�0�B�pʌ8j�a�b�<���M�%���DE��{r,}��&^�<9�cW|��ԧ)	(j����Z�<�Q�ʽRJV%��
*�ڴp���\�<� ��)�����HUA��J�8�"O|�ᑊ	Y����r)^5}����"OB;�j�*5|�E.?��"O�Dk�*�t9i��ړ����@"O�@��i�I`) "؂u޺`�"O �0Qm�% ��c%�C�z���"Od�(��ȥUbB-�怄�z�\��"Ox�T'�H �C�?��5�"O�#K=It4=c�KȫT�l�Q"OD�%,�>:���*ՠt� � "O�}h��.@5ڐ�#�V�%� ��"O��`hכ S�=�VBS�pL�5"O�0bK�x�0��A�
$7Z���"O�4�'���9�X�b jԐH0�Y��"O�����l2�S6j�d"O���.ѣv6t *G��zT�"O\�1u�	M�����.AH�1D"Od-[��tiְh�iR<\ �{E"O�u!�?qS��%���|�F�#"O&]��:ގu���Rv���1"Oj���1T�$�u�ژ5hxہ"OH`��NI4�xq e�!J��w"OR���I�b����Q-,;���"O�@��]V�PY0�0(���� "O���#��+>��x��
N���"O��°nM�y4��B�5:�xq"O|�Q�A	�w�R�:G�Ī<���"O.Pa��K�03~S���r�x�"O���%$��F&X]���Y)H�i�"O�5��ϛ�Yo 9ѢgG�H�j<Pq"O2a� �HQ�L� �f�%T���"O�aVF��a��AKq�:h���"O,E�F�Û0h�40�E;-J1*g"O�(RD?&|�	�n�=K"J�9"O��¤��������tz4�"O�p	��X9O�\�ST ��NDd`�"O���'�X*h�ح�t.�I���RD"O��bh����P�BvƔ*�"OVC
�����1�'�`��r"O|�Q�"fh=�ǃ#���x�"OJ�S .�Nb(K��$�ɉ�"Ob���m�O���;��D�Z��e[�"O}	�� 2g��H�W���0�89��"OzP��	G�%4�aV�J�A&F]��"O�XF'^�E�L�� �2)�	{�"O�mk��"A���`�aL:xm��"O�MR��F64�L'"���2"O*�H�DՏ-�����@G�oKX�b�"O�t8e&�!��ّU�.*0�
�"OPd%&Jq�~�/�l�I�2"O��2��$>��v�<,��
T"O��O�4�������96�*���"O�̸!
č?FM��h��`��"O2l���8�I�I�O�>�[�"O$�s&�!tʉk%� Bt"On�P�P )�����S�WA�M1�"O����ׅW����V�=64!�"O|�A���9=W�ɢlQO:`�A�"OpE���ӟ=�͂�+�<�2<��"O����\=`D0��K�8�fԺ�"O<l��Ý0K�l|pk�4-�j��d"O\)[��1R��b��I]�� "O��U�ťFqƉ(�NkpEys"O�� .�1�Ȥ���̟��k�"O� ��3˗�J'4}(�E�q⺵��"O��hgjg.
�I�Ȋ��,�d"O\�@�L�^���K�A�
d|J`�"Od'D�L�l�(�J �hn��p�"O�u�a!��A�.�J��Zp{�"O��񑂝�b����E�'8��"O� �Ə��%34�!�ϛ�]B�Q��"O&ḱ��97�iXa�ωL%�8a���Ҡ�)�'�D2p�5L���9c
�3؈�ȓHo=���#1d��b��Q�f	�ȓi��aԅ ~L`$��i�~!��#if	8�&ҿ&N0��c�k6���r�����GקnP�AC��@����8�0Փ�n�ڦ%��-̗Z����ȓ������
#E��AIL�0�@��ȓd�B�;�n��U�Ⱥ��
�d�ȓE�� q"�JF��M�$'	mά�ȓ,����צ
@��e3��Mkrԇ�	b�'�P-Kf`��m`t֧�"��	�'�L1��he��h�� dT����O<;QF��/{�p v
�+�n�X1"O�	�˅�rm�1k��V1�����$;|O4�q���,���x�H�&\�����{x��" � W�H����е�0|��O(D�d����$_����B��6vL�i5f)�O�w��;��f���W�n����}�'N∪��J�Ss�x(  �'Y�:�%L,w��%sk�v��k�'���9"Jӊ>�<l�S��/l� �
�}\�8E�Dk�#�p\��R+NTacB�D3*:���'�Lx��%��� Y��àk(%��'nў�>�B1?O6�k��*e����)12֭�2"O�$�PN"�M9�J�|Θ��%_����	 �����%3�5Cp�W$Q'r���0?����?2:�Z!�<
� ���H�<��F0\�B�_�>Nr��Y^���n���t���r��*�PP�O�27��P4C�<�I����ɵ	�Ȱp�4~#n���&����r�/<O�tr�	��Cش!���ȁAB��R�
OH��6���8[cd^ J����;�OD�'�Q>��ӵ�E94��>������x��j�'>, Ѣ�֕0�L8d��IUT��'6pap�-q-!d��I�L٠L<��k-��r�Oж���\9o���zS��s{��'+���!	X�^��xz4�p6xb�'[�KA�d��gE��QqhP��'U�i����!Rɪ���v����I_ў֝`�'���Q �B�/]����*�&��A�ۓq1Otli����)*�����mPA�"O8t1�)W�1����۪tll�H2�Io�Oӈ��׈2D�N)ZU(��,E����'�1O(���L�FN� �Ǡ_���A�m�_�!�֊��i�V�4��:D!�d�l+��#��\
yH��FcJ?!��D 8c�&-F��B�&�!�D5JR�|�X2S3����+<!�Di]��۲r%fPx�C>M!��#D���M��t�鐏�`!�D�6{IВ�o�(؀D��/!�� %�£���ڸC���r!򄎴1%j8 &H]����S�JG��O��=���l@���=��i�c��?��rg"O�\�$��I�.i0�n_���s�"Or�:�'�	K��u@S,ݔyA!�i$��2q�'���ȟ�� ���bꔗ9��ᔏǯ'�LP��"O���A���Z��`Q�W�~�ıZ�"OȖ'ʡ�"��GUu�d���"Ouғ�0�1#���h�@dB��-�hO��&=�����F$�Q*�=�!�$��)�V�2��$R8a���ۈ*�!�X����cU$:��8��םcG!��S�|	�PcC���("��H!�]�9�Xu[��P��33�ѽ|_��ڟ��V�d-�c��I�)]*Z�S M63`����@�xar#d8X���co�Gx��)b����0�V����:&�މh1h�f�<�!
�130t����ġ4S��h�i�e�<!���
9Nؐ�DHH/��`2�_�'��?I�Q"2R��>!ꩡ�(o����	 *�
�p7��<!��h�,��J�&C�I'��L����<h, h7��##�<C�jg 9�D��I��a֏��e"���}}�x�T��%�֝Q0PL����
�Q����2SC�I�.��8��f'^*�(ׂZt=��	^؟�zpBW4���p֬P�&��	!	7������J4�6��Um@�7"O(}��C���1�T��O[H�fY��8�[�P�O�>����ύ$w�9�ˎ*y����We0D�T��a�As����k��F$0��hO�Ӕ�v�פ�{@�3 ��m�C�I�Z����A��K�0ϝ~��˓�hOQ>U��	E�S���� ���ݔ��7D��ۦLF�eu�ū��ƏU=�;��w��&����	�c��)��Oa�jP�R‎������<���>a�����ׇ/��[B��j�<�@#�u� R��7��;P�D��Olt�-O�Ϙ'/<A@��sQ�X$�(*�'��8�"��D�t1�g�_�u����+O �=E����R��B�	''�@�� �yr�Ȗi���*� �vi�ы�MK36�O����M��G���#0[x����n�IY1��m���:q� UYG"J;K�`)W"O�,�$�Qh�н2A"̧V4����'
qO,�(vl̃�4�Va\�L2=��"O��1S��4��� �H?Z�T"Or���AV:-����"�WC��l*'"O��r�K�
Z|�c/3y�*$�x��'��@��ȹ\�<ԡ7DԮ5��ɪ�'9���G͹].:`�f�*FN�Q�'�v�T-�.�b|{�&�<z�X��4�?A����i��(	SO��(�uᔹ.�^�K�'��Y$E�
l�,�e��waZ��'�������h�D�TW1n�T�����5 ���"b���/(w���'�0M���&.��KC@�'A�������_�b�'�a}�4E���\n��kc$���y2�H2=2Qs� M�d�1���ē��D+���B7Z��R��3cv(d�^�%!���-H�d�	�%��gX���	\/a7!�D�!�)	ă�#A��g��8��ȅ�	uј$����N,�R#�T��Ɠv���ɒ_2�Ƀu�C�}��Vy(�-M3$��O66@����� �|��R��5	ң�!Cy������4��"?ٯO�c?!�PM�p0�"bU
��X{�M,D�0���,KfDF�:<8��3�*D���r����(8�(�P�(@B)�	o�'��I��R��sF�U�Xb��G�FC�)� 
]92�МA�J���d#����cx��XWǛ���1��D1.php�-D�Dr�K׋le�봯��w��!b�+D�|Y�B��� �.�(
.���@�(D�@hƠP�b�����=�P�*��'D�C��A6>)Z����C&�Iڲ&:D�ذ�o*A�|�9�[��#�L6D�l9�"����$3¡Q�xaj�s��?D�T# !�	�<�K�k�th��!�?D�\r��\� �6�!Rn'���"�n:D�0"�J��	����ҡ��\!P���8D���i"E��HE�Z51n��  �3D��ж E5:�R�����-��c0N3D�x3�@A<]�U�3��p-'D�t��B:�b ࡬X\ �� �/D���[�K�04Fc�D��QX�;D��z��;v}�5��2�*��N=D�� �C� d����d&�p����& D������4������I��*�=D��:o��@��Ȁ?��t���/D�(Uh\�d��p2 "}LT��wn,D��@6cG�T�8�`B&WB����)D�����P;j�	�j��wo�y�@)D��8��=����w�
,Ԩy��g%D��s��#��d�s��3}���Y��"D�`��D\�9�� �,U(YR����%D��2��V�Ĩ�"
��E*U�.D��[�$B�z2 \�ԉ\�u�,|��"'D�(#� ϊ�ꐇXO�N��b�%D��PI�):� ���8�r�c%D�\�r��3~�0��M+! if'D��B5oI�Ch��U�M���:��:D� aq�MIԔi��OM	3�t|I�d7D�H�dï���eK!Ib����1D�tzҤ\˘0:`	l���Y�'"D��ja��E�vE#�Ar�N��pj+D��2�0�`�&F\�"�����'D�La�T{��7�lt�����9D�L�j�)���A" �"� 6D�hDEC�D�Ǥ�>C��䈣�4�Ol����Z�-X��'m��c۬ �e�6}���"O��B�c��*�4��.Y�P@�"O(� +�
1��9Z�_8G�,|YE"O���N�4<�b�#�c���f"O����˿#�-;�Ǻ��Ś�"Oj��E�Ay�p���*#_4U"O4H�s��FA��ر�A�G= �S�"OP-�`Ů��L)��ŋ*�L��"Oj� �bZ�~D�P"��;)L��"O>P�""[/y@
�� 
[	�d;"O�3���j¤���Ap���;�"O��[e��K�XpF���fB�E�"Ol�����ި�R�C�2�z�"O�����u/�IPs�U� X!��"O�mB�F�BB���e䑵I�>���"O�ؙ���v�`����Xz"O2�3͘�j|���R��*B��ab"O�T %MȚD_ڜ9#!�e���B"O��G!�Rn��a��0�)�"O*8�s�*`��	2AT�T:1"O��S��D&'ШYr"ϙ/��1�R"OR�a�E�+����b��:�� �O\Ű��_ B��O�>�����8<@d���>i�V�Y2�$D���l[�0Q<�pr���V.>36m�<���	�%\��4�X4�0<�  h��o��*�у�[=8z���'q� uU�O�)0��0 �z�	��4��0Al�i�����Gg������)|���׮ف�Ԣ<р*�"Ea����I\�x���O|�ӅI�pV	�7ƌ�{�����J�<i�B!����G���ʓI��f�,�!!�nw$�Xq�+=����'<�PQ�U��!��@
�@��Z�'?��1�B��L;h�s���<�,���#S.	�ă9a�ԑ��>����$Ġ�89���J�a�n�SA�Ls�Q�r!��,����r�@`G����W�ֲb�(�g�/������A3~�f!#�At��04� 9*���֠�>'����
B����bL8h���ē;���3��S�t?@�!w��i��b�������Z�l�@�Sg���`K!�$C�-H(�C��!B5r��"�@�!68��C�7�8r�F/�  "R?�1W`P <�X�ܞI?�+�$#���9��Mq��b�a�8�\D��0���U��d��K����5!�3?q�তN�
2S�i�"�R�'�ю���a�Ea`�����r>rɉ6h�ٴ����|& �$Mi��5�I>���͝j�����[�dM�7�B�\A����Hz�M	�a�.ae�uH"F���� ��gۖ���?�R �_��<��$���S�^�ƙ6����^�&@�z�F����\�dhQi���l@��7Δ�Z�ұX��֕�T�6П�.χ6�:�������" I6/���ݟV1d@� �L�q�çI|�`C!$S+Q�<(6dZ=o[����F(���Ӂ`O������|J��*U�(=H^��q9T$�7����w���m|�D.9C㪸p�/~u��K$p��9Z�ńk�p�矔��]�իE�ϳ��M@#D�K��E��Jٜ��/X�4@� �t+�"�ňԍY1��IP3D�H���	�Iِ�qoY�x�}��#A��Z�L�P>F�g��3t9�'FD� �(��mW��1d(e��-Cs��S��M�ր�<E[D����B�Z�0�b���S��Ԯny$�%�S*��`_=GRVњ��^�<����u�#A�|ء0�N#D�V5�� IU��1
�.��� *�.TJ�|lZ1F����s�G�̩��yWl5��93'XRW`�+��M�t7톞9c�8ઋtȮȪ��|�c��bFA�1NؗZ�0�]6[�Z<�쁦Y����`U�U�m�I|�@���kB�c��p>5�W��\�����ԹU�E�e��#��M*�Q	%�q�S�C�7M�;I�4:�D6)M��h�!^@���,OܨpD� H�b5�f�R�;}ěӪ�BR��pW&�2M�<ّ�' �A2O�2��Cg��<��!t��va8����<s�X�G�RL�z�
.��6�x�,=���<AGH[8R���D �Ա�N~Z��ҟhLN�9B�\�Թhf�?E|&��V�E�%��|�uH
d3z�c�'^}"�S,D�Z0�s�ez0��5�hb󥝄#6�5;�(�7B����	$3V�U"��"~�	�qP�²3���VbŸ~��� Nq�>+C�κn"^���́�B���7�����;{���;_���q��!=�N<�EI�3z"�=��b��1���.N��3�!�I�O��c�@,N�<�tH�~��xA�n� d�H�1*A1�	�z��H!��#a�X`���H/}2����Ub���Õ�}�|�T/�s����waL�;2X��<�G���?8N�'���L��`aWHN}ިۃ�T�i�  %��7B	�'FO?q����V�B R��'��ɗ-��(|ǣhܧPF��.�%�2���� :lw�	�1�
Z�Fp�Ю¨Id����\^���'�"����?�]!�P�;7�S�nJ}KӠ̹��$žr >Yq��T7��)�'���� �B�O�~�y�dM�5A���R�J��<��$O�DI��
��ޯ�� �B(M�n�)$,3L����E����m��Llɕ	�m�~�OB�ȲkS.�اu���-�:ݠh�#.u�G�o�����<�lx��4xwn��Z�],T��1��D6EG}���s��ICS�T���1�ěŸ'|�82"�] ���`9�����F�%!�����:~PL�c����>P��cq�H	$����Ņ�8���
�e�3�EwxVp��+S�j��J�M3gaBL(G��-�,�Ѧ�k�بq�L�����V�W�7� ��!g��B1 �) ���3�'�j0�C�I�*����6�B/P3�8#�&�'*�вiۉk�(�#ɳBg�M
�AS�+�������-U:�kf��"0����n|��v#9]T��P�F��=�>���\�(On�:�Bw�T��_�g�$L�w!	UXVX0��D6L��i
��}�%DEZ@���b�<�=!YhYT/�)1�X��l��(���<���L�,��$J�@�E�,�����Ԙ��Ώ�xl�v!DSհ�ۤ� ���Z�LE�nVq%���L�a}(_�3��7G�4L�J5�ق=��5��C�/u{�X�A�(Q-����_�?��j��6E��b%��ywb�)�5Y�Ǧa<�𱧅Ɨ�y�0��tz��Y�Z�P�wLW?�hb�ȏ't��m�� �z� �1#O$3��X'K��_�D��њQ2�6퇳Fk�В���<6:S�T'Yr|0{��-H_��@��3DJ}���s����q��.=7�!biH�GdI�3��g��¤�Bc���9���9�� �&.Jw2�P�)IA~#=	b�R,<Z����>1�8�K4IY !$,�³�>���3i�F��%Z҂�.>\�����=6�(�d��"$->�҂J�a0��9y�H��f�H�+�N-x�ƌ�b(��SQ�=N��e��P����I�AZXT��.ZO[���� ���qtŅ5{�����UiӬ���\������GT-�D�p����,R�a�$��I�-Q�u����cYNH�pgP�z�h��RE�7L���Eĥ3ƍxA�$�9q �`��s� 
�I�����s�A:3��X��'�A�K3c��#C�iJ����]�Tjd�v�R�^��}y&$�4�U
աG�k? ���X`B���㝧V`p�&c0]��qa�D+��U؄���V���zC�S�9�R���]HRXYP��5�2��3..T��u��	�H�q �%}b�I2��5=5P=ô _�th�ǦI#�`m����I�)��&{n�(!��';L5��� ��HQ.�QÜ�Yc�1!BR����X��
D %�	�Qǐ����$ND��$�Y�� ��J�@B2)Ih|#�f�$ 5.�ӈکS6 �D�4Un�}r��OP�"�!��#;��b���f�)�T(|<��2�*rM��3	�$X+K<�$�b"}؆&΄qS��*"��M[�T�!ob�lHgE	:eVѐ$��9�M��f~���o�]�@ &g_!k�@s/�q(ވ�Q�Hbp��v�$1����[�ճ&%Ұe�z�)�戎[V`��U��l_:9#�.V�a���V_���e�c�n�y��^Yt��*Ռ'�����iC�J|���EJ'bD� ү��9� �D'��-X�|�0f4�#�F�*UA��h.t��h+5�C��-P�D���Å-��I��Ri83����$Z��i�R�����}A_��4�O�8g�TqP�D2�<�5�\�lxژ�R ]�bﮭ�2�*r_"	P�IBdz2�)0a�Lֆ�"œQ�>�Qv�y�DMX+s^81(	`|8�i�᜔K۞�bgeΞ�p�ВU{�4�B!@Yˉ'��A�������X��$�jN�#\< �Q˙�7�u�c�V�0af��E*�C��3����M�f/r�F�X���tm����g�.}k��7M���a9'��ͺ)؀��N�"YR�+�v���욀	ߤe���S&��qG˿Ƣ���M�&Q*�k�8�~��T��d[�H+���+�/HX����C����牯b)y�ߔ~�4����B�PV`�g��]��N�l8�5�����dϞ~�2��� N�Xf��u(Р��IO=���S�ڈ[�"݆�IU����W�D�H�v�#!�U0a1 q��S�6�14M�GŌ0F�&]6>9r�O]�D�L�r�g5$��M���7FP��5sB̘J5!Z@'C�d�xg��9�\$��{��U�t-�E�HP ?�`�#E�b�^�I�b���9�p�ֱ59h�2d�Ǹf���y��^�
H��Fg��8���=:Ɔ�;��,`mx��U��Oܓ!���!�J	^�B��sK�5!�"E0bJ�%��؅鄮:��]�j�$ ���*!ri:�,jӌ��4� �+k&�;���=r�b���|�1��nC�W�������+d���ׇ��~�ax�CX�ĝ��I�����A���Ĝ4/OnD�D�X J/`��rgn5,JfH�T��^^k�i�@�9���F���S����Zy� m�r�x��ĭW\ H农	Qh��!ҁŪF�� �I�Jr�@�� \�J1䟎q�\�a�F	Pi���!��B�� ����Cf��:PS�@��s&:���� =!h���I <"n�i�jC�z�}�DCƇ} ���L�+K�P���ЕO<pL�7���y�x��d�E~� M��cǅ~Š�,ǪI�^��  �F%��ݐ:��U�Q`��(^�#=�N��B�nɟB�0�p�C��-�	�t��� ᢠ�V�	�ZX*��0.�\�,`5��lE� �!��N������%�D%(����ˊ+�J��_/^�LD�ᢚ�?���
��8���u��%,���S�.�Z��ӡ��Z�^�@)Qt.p��ȉm8`ZЅC�)��v*t���	"x�V �)M�(Z�	�9*���w)T�7���O� ����� {�X5[�+K�**1i�;/���q�
x��V��
����C�@����Ĝ�|%���:j
��������N�dK&.P�<�pmZ�MR2��j��9�#G� * �}a ᝧ#(:<�&��` ��2J�!puA=>��r�:�pX�L���c��	p�61bPX'�ϴ������N�l�2�`��T�ސ���Ye�l���B(���!UjL:6��(�%&�hOz�⃌�m,b}b1%��f��0%�G�<������^t��FݎUl���,@�o+rU:��l��P� �;��������85�1mO,$U�0Hu�]���0�3�O��#�� \2��c��OE��2��ۼ��,�%CI�b���X0��)R\��CQ�i�|)����Ha�j�#��X;dIXU�F��qhF���7�O��kCB�$u���*��� E�����BmH%���#��mP��<|�h)f�7'4�I�ꛕO�g�FjB)2��&���Y�v��!Y�%R"x�l%&4�����C06�&r��&@(�\��*ͨl245��S	V��	٠	��4����mE�>Z�U
]�Ty	3h�E�B��@US��#>q�$H��ܛ��V)Q��2���O���@��x]ْ�Y��j�;QĈ���� ��/\���!Ndq�.Y�J��  �g92��	�/��t�e�4�.�O�@���������8��@ARL���	��<Y�}��"���� �n��X�Q��h�'��3)θ��Y>(�@�Zf%8��|"+Y�f�XH��l�����b�ƏC��BeFܙ=�h����)Lz�1ĝ/Rḿ�i|�����I��
妜>��I�a2|�F,@�*�`��e��a��{��]0t��@[�`I)�K,P�)� `�2�U{f��N������<E4���6���c~>�$k��)�&�4��l�Q�L+�GB�t�|�4)ɘD��R� P)|"P'���O���i�*��a��bGÂs�\�T鉙G��f`�/q40G�ߗN��0g��f�+-�2O�h���3�0�	�%٦q4�!�,O�!�R/:1�N ��i2T�ֈ W��0*�J�k�nŒ��1[��LqG���oT85�D��	ܲV�ƬP�4��!���y�2-�SN@���HAR��ۄ82����	!~�>	� 9�L��2iЍz��`B���AyW� �@\+#��L�`�;�x���Ͱo	ʡ*B�O�g�dND���2��(�` 0Qẹg�|�ďz?Q7�)kK�O�Q�@-��s<����2a�@z�O�=#6I��Ɇ�j��p���U� �B��h�vD�HЌ4Ɋpo�?��'Xճ�I��0���'R�$]b1@A�4tν���N8"(e
�lҤ|1�]����"%V�4yZa���Eo�aҭpB�##p�e�A��
Q�ݒ$S��rb�ظ'��	1ˁ�^ 4Ę� �F�,�B��+D��QkG튦r����oݔ;��Ĉ�7rܺXBg� 	��y�c!�)@��q+�틤v�����]?��Zd��?��i�W����/�L�a��U��:%a�:Q�VH�%/a� ��e�Pb�
 Cf*��Y<#O4�r�*OFUi2�H�~�t� "�R�����%Q�s����'!F&�"a
N�ERAjw�I>{�d�r�iL�� E��6�J4���i���� ��S1�e�@�éF!�6G\���8��B�o����`��Uz�5z�$3a7�<�$�,`]VT��G� vL,[փːJ���Rf儗zp�J��"�	{u�5�k�,�(�!k�r9�[u����1�"��Q�2����9RH2�zPk�.�(�I�:r:�.�	��"V��C�ε�ào���sTh\.�9Y��99@�y��8:R4��mN�C�%إbX�A����+���0�H�5>�����H�J���J!x��x�3�Z�Y�t���U:� ���7:����EV�J�B� �3�nh�ȡ�"D��k���6[�D���%{�u����7[G��z7&�6~��}Y���4q��%<*D�I�9���#K?jbҡ�F:Լ�D,�V���$��!%:2t�H�	�l"H:bJ��i��PS�m�1��!��H�^�Ö��4�p���^�b]�$��i���!��pi_	pԈ�����/Gx����@�gF�I��Y�b�Z��Z(Z�� �@�\����F{���=a�#W"?ˌT��T�.�dh��؆@� E*V��%x\J���-�Hx�]`įS�g̀@��Ŕ�.�ft��'B�.]*F,�&}DPY�GsDy��>�<��D'Z��Pg4�I�B&�1�i�0\�x���T�r53Ӥ��Q�(J7��7'���1�H �5F~� ��@�u��x{�-����'7�n�@��������ɗT��ʆiR ��yx� ҐR�B,����� ��
C�1X�&}���S>�@�O4l$@���Պ�1e��(/�541!/�i�ڀ
���l�p����kމ�����X"�Դ61rXa,���43#&4�1d��lgp�(��lӱ�p��4�r�a)E���1���'aѺ>2~���S����<��cC�S�2�3�c���ɏm;Ԭ���" �f�� �a?ɑ�M�!��C.��''NZ�G�b
�ڒ�[M�-sahU� �-"	�,ʸ��T.8lO"	a�噶6P�
���'2W2��va�#Gj�ek��/M�p*K>a�U/L�t"Se8i�O9 h�,��	��`1�B޴:�n9���d�&a��Xx奋���O`���U'�% �ݘ��5�B|��'Hp��GD-(��SF�m�չ-O��҇
��}|�)O��|b��B!n�a�î(^���
�F�<�T�̮J��	�m@�[]��!oTE�.�̀'�"O�����ť6� 
�)��@QH�ۣ"O~8V�M`t��ұ���3�	(�"O4|�ՃR�LM��Yf�}�����"O.��v�G�,�yB��l�(	r"O���5B�l�h	�ǆ]}(X��"O��Ǣ���x5���0U椁G"O&Љ�4`�4�J���;46��"Oh �u�0KAt�H'$)T�z�"O��ß�8_P��Y <"����"O@�YU�V&^�ɕ���=��F"O��r��R�{�h�+3J��"O�� F�:@ՈE�m�0U)^,�"O���	\�V�qB2�ئK.1%"Oh\I�̅Efq���D�4"O!��Ǎe���@��k{�-"O@�"�oΈp�$���8YL�K"O���4j8����dݳ1�X�"O��plL�nB�Dyq���Wh��e"O$��pGB7d��P����_�["O����AF�&%F�h  ��:�j"OT�ɂɋ�=�0ȁu���w�ru��"O���`!�0�`#U`՝D�y!"O�����{���+f���଀�"O�x'��JД鄈�$<ۂ�u"OD�2KU�E���a,N'%m<��"O�ݡ�Ȋ+H�*�;g��	T�ha"OL��レ3��*cɃw�Z�"O���(���R!r���rg!�d��-�h|�m�O)���g:el!�$�1j��s�K�.��JG��PP!�Z<l��j!"G=�8�B��*AX!�$&+(,H`��7��K&��TA!�I�
�
�Q�*��ݒӫ�TH!�D�3P�:q��>Q �4�QK�/t!�$�9.�zj2e�Ig��*R��&b�!���JU�-�b�,lD�����GZ!�D\�K��(��3�{F�OGN!�F� ����B�7C�8Ν61!��S�-Kf��g	�a;8��m6!�dķ"�V@�b͆-��8p"ݦ !�dո����dE!$���@�]�!��A�-�*��G@Χ(
��vi!�?d.��ƁU'o_��a�D+N�!�d-%@0�� H�1$��� ĎmD!�D],��$��j��:��2ӏ��J!�� x�C���4�֌B�i��[�̫�"O����S)D$����I6, *��O�L12`ID�Z�O�>m�5 2	�N������6�~���:D��V^�ef�B�
]5���p`ô<�JU�u�2T�����0<A�b�@�>���ǿ��}���iX���� QmRxsp�ڈuL$��傺j�ᢒK�B2���A�'g~M���՟�"رFǋ�a��k��$Z;wctUҰ�(ȩf�+�)ߚn����MT�k����)m�!�d�8���A`̗-4u)E�ۨa+��˱� �l���P�S ���)��X���ܕV-B8Ѧ���g��3�#"D����劲~�tp��X�A
�cͪ{Z�,;��3�|8��[�D?��3�}%��"\ም��W39_	E}B�@�q[:$�]�r-�cQ�{. (�E@�XZ!Dex�&�ҕ��'RLR��%�O�0��� B��53�j��r-�'�';:\��i��`�v!�WK��l78J��1'���ɟt4�'!�+D�r�E��L0��8D��q2$R�t�d�Zg��+F�c���&F,�'�-q�(�ɲdN��(�'g�v���AΔ!t�9X�'�j��E���`2P`��Ǻ �-��{�CݐxӔ��~B��5fv&�"1k�/��ڒ��<> �h�MR�		6�߀P^< �'gF'��e����^&�<(��_�B��B�P?[�#��Ƕ;�p��J�),��'�`ӵJ�+(����%Y�B�pt�C��5X�\�j�iB%_�JEzs��(�<C�d��c�6L��4���H�t�.�$d95��G�	[/i]ʜ*�l߀ �|��	�g����E�+F��%@ +)^��X6�[�mW޴zTL��t����yw�<�Q��.^�ʡ1� ��~2�Bw��� &�͠��|��SB��hŶf�š!j��";�@p��b�JlcF@Y��t��o>���4b����J�7!?�Lp�`�$U#�!�Lh�4����N�og�Tz���H#�A��a~�]{f�j��Pь�׍O�P�+��0#f��b�)~L��4N]�G�D#� F
,���'��L�ܭy�/�#	d��`��<�DN�E�V%#`$�.�*A���A�`�e�QLP���.���dV�EV!��¸NX�0Sw 2Zd�XDeA�V�, "�!řpU���e�te{�f#CV�!�ۊ[#��Swf�O$<���u^�����?vf��y���]�!��(P���[УJ�`A����݌ޔh%��>8��oZ_�ة�!�z�$j_��w�	��\ 0��pz�ȳ'>�b2�x�^�3DF�He)&B�M�'s��hs�	͢#Ȑ`А�iޅ�Aڪ79������� S���ȟ�j�C��y��ah�(	�V�j�S*6<���/_��SE�G
����M�:?H�XU��;(ώ�JB�bӸUP�ǁ�� �1�e��^D0t�%���\cMj9� ��i��a�D��Jz`����'�8:��I�>��ú
��rD�Opr�:�R��2���a�!@\d�q�!X��f&N�!��9n5�p
��<ٷG���d��h� s���K~z�Uy�p��p"�'D80���9�R]��MV�,��+@�1ږ�Cao�E}�-�'��sޥ��%F^d	r�# �����o44L"�Ĕ%� *@m ؟"~�t�l��pȚ�.l!( -�i�X{'F=��-�ǂ��z���˴��@hZ�{$z@����l	�Dϻ;]8��EQ�}~R�K �H�x��Y�.�"���^ 4N����:�ɀ5K��Se,(v\Pc�����!'�R���ꐯjH�dD��QB�(2h�[�ْ�����@)�U��	���@&-^%X~�feA�Y����l�e�1O���l_�`��a�5�d\,��+��I��� �YC�������$5(t�$���E�hY;o�'
�@(�3t���4��F�jY6�bgE�p�=����)h؀�eR.3zNh��'^1l@��p G�lU.��'�v�1���yW�	e8LF�07���9�?Y&��a��c#l!}��I��c����p�f(
d�H/G�ΝP�!@�{_`P#���"@���2�H����WEǷt�r R�h	�B��䉋,	IR�@nY�C�j��<#0�
��'�i��*�F�X�#�")�p.�*&T ���6VJq�>����A�$� H03��!%Q�tQ�/��Z	�ez�m�y@X���.��<!/��:6GK;Q��"@�	i�^�[bb�d~���GeV<K��P�ڦF�P�@`X�SRp��d��p?�7¶ai*@ ��)e�䉕|$0L[���ة
��3fO�`��4i��dؠ �;P�96L�y���[� �)�&�e��4@	$�y�B)R��af��E��h�ၠn�6�Zňg�:�IDH˂0(���B�P��1��R�A��08s�@"h��(�r�( s+�Ea��蓦���0=����4NT�)ナ�C1(�6M�4dE��X rA��n�Xm3��6x(�������`٦6�hOl��JS
i�])��W' �Da�󄗔%�l92e�<T�$�����6bh7�+D����
�R��庵灭X��J�]LmzՉ^,X~Ђ�P���ǟ/A�1i3@�\/�TJ�m_�n}��R�N��2
`-�u"ɦT�����'�,G�!��W\-�H�;]�t��棍8]�� ��c@9 �>��d�h����E��"%CP
H�=lNE8fJ�,.AZH��钳�����fU�d�b�b��4 ���9fXqP��i��d���ӓV~�EEC�h��)@�϶*85y���[U6D��j����'<z��2a��QҔ4h���gjj����;^��P�噳<�BHj�Ɨ�lO���ՉM�$S�	�3���c`r���鉠+q�����2��D��T�G�1): �����D��A".z���C���|h��� -�G�/I@=�u��C�x�f�R2��*@dU�[&�I��D� @6M5	A�i�n�JKr%z�Kפ�N]j��˝�ײHy��?rO\�۔��9��]��ʔp&�VN�(p���:G`��}�r.D�S8Č��*�:b�*T���D�@�O`�28G�N� ��L)(����c��*A2�cti�S:���'I m��,��Q����h6�
s��vi��iMcph�aO���GI�o��0�vGQ6���(�Ā�M� 0�a��	h$�5�DfV�x��jR�ܰ��\�Ilvy�ч��1^ �Q����i �!��V'��r#eӟ�R�1��\7\MBIe�co`�c��5!�U��䔐fU\� v�:4^�q#�=ʓ7 @�jV��W����i�_@��/`'JE�j8f�H�	!�"~:N�J��S���sf��O\$��ㄬg+��ÈA�� JVI�Z_�02@�;3�tI0	.�����`�@��E�!O��S�O�Bw��jP�Ec\X���<[1��X��PM��t�D;b�		Ex ���QC`@x���>_9�h�g����ᐄ^Lĭ�'A�-;�'���c�C�&Vl��R�?>�<sB�H:3�>�R2��+���^����q�XbΩ�7A1�M�&��<0���p�@95�.�`��?j+z�+�~>�C#Ϣ��Z�\�N���3��h�����*#��9	�9�P��V ">i��
2��F������l��s����%ч�Y�*��h�EM��*u#��֒^�q���ꦉ���psK)�.�D���̆�`�XCJ�Z�B���\�l��� 	7��I`l��� &��i ~��̭b��,�k�`H ���6w��)
˓>z�#f��A�dQ�#��[�D���$��̏�~jT�����E@���`N0_��@�����(B�K��8��lO�z`L���$�AG:qS�D���e���5[�`��x�Kڎl�����%k��ؓ�ֹH���&�h�^`�&� �Pq�(�T�x��i� *j�1�4!/Yk�J����E�?M�xB7����<1�C%'�2�U�[�:rX��.�'�,t"��B�W)��SGM��qbC�%�"�H�"��?{H两���QZW-W�n�j��A�
��X�5�]t�~%�a�G.s$��H�Ex� A�錕&=p۷�λ"zm�b.f��Pi�c�zR����(��!q�I̔%:~	�7�9!�&E]=%�>��2c2Gk~�s��A�/[	 B4	�/�I��I-���qGX�/�L��u�n78���K+�*��h��\�@��6�S�1^��ʙ'�D��H����E��^�hqT�D��\c����P�idbS��<�0"�I��]"4�D*�	�<�H�*����M��a�N����#9v'$i���C?��s��[��a;O<	��Q&mz��.݈H�6�@�$�� 
��c�.�;=��mc
D�L ��0�ٺU۳�1�FD�\w,x�.�;g���Z�e)�yWğ�-��<�f�X88���$:E���b��2m�*�����-L��k	Ó%M�9�d����@t҂$]�un>=�'���d�S%�>�3s	Y�$��$[��m����tm:5K�^ �Zp���ܡ}�􀂰�שWg�t2ʅ7=�zb�U.���b�M_�4�Q�S���(�$�-���S�CAw>nZf��L�ueT�{l8�qΦB)�eQF��%XRN��p�r؂ѯ�+]v	[w�ǥ.� ���G�/�&M�?��K0��Wqj�+�q�vŘ0�� �txc%'ֿ:V�!7��
5���-��Ttl�#���s�x�ɦW�e@��4*���!MP#=a�
ӪG��� �m�h!�c�$�2�J��́ p��D��j����E��0D7�P��MO�vݸ��ˌY�x-�$x�P""h��0F�t��	�}!�2#f�"���!��Y��1�ׂX�5nBpr�1B�h�UI��x(�s��$&����dQ.�HM��h[�A ��Q �.IO ��͔tx�$�P�Y�M\�%X���
x�`KB��>�����F��Ǡ7$��� CYHU�8���
�D�Jz�u�'�L�"D� �HE�Gb��Č;�O�Ũ�T�څ~�d)wnS�t�2A��N�<�P��JW�p�4USߴ)����s��*�Nђ®�n�zM�랜<z�U�I�-�?qrń�p|I��
c��u��IWh�'p6�:e��&�*���T9�6M��'��SK����(�d�W��3-@u��ތ�:����t�N�ZBU�'���PNë�ў�p�%s]�4�T��-@ �(��݋v[<�`g��H�P}��D�d� g�C�rX���U+K�xfn\rU( ��M���	�$��-�Z bC&V!�0�P Px�H�5��!F~�S'�� �ftr� ��\l�$j���q���F�7i��FnӒ̈�����D���K҂͏Pr`!H\L΀��pl�f�hjVlćf ,Fƻ,���4JOfD�tj�D���NN����t�EE�81��N�)�����JnJ�$��A�����jЖ���o0Uw:�e%��q[:#<���&ܴ!ׇ4e��P8�J�>X�l���~�1�kP�)&$���G��m�[p�
��T����B\}Di�&�E�f�E|rBIjX�����ٚ��[&�4����+
�|ԁ�J]�]&��@�B��i^���������O:9Hh� Mn��Z����ˑ�4=4%xE�Ѷ!La~r��%�<e�1������/�"���!�(I���E����C��!=�� "��� X�P��8��1ʘwb�T��an�~���B>��B��6(��U�*Rn
�Y4i�JX�oE�`^�U�A(�"wрu�v�L�Q����"�M��j�Z|��/�dY�I��On�����t�hљ��X����V~ܓnxM�C���AN�&kζ
��&��<��-`�/��x7�>z�(��F<���r狏r�*�˗�0\�fLȋ��L*P�K��YP���hc��+�\�%��	-���\�,8é	�&�lʥ���/��Ụ��3�����I�6�v�CoI�^gp{�	�h�
�B�.7�0��$�%�@6����.O�E��@�wލ(��2M� ���|�� ga
bz1ˤ�2=��i� N�sԅ0��ֲO�9��;��Eԉ9O�x�E�Ze�	R\�8�ӭ[Ntf��v�հea�>-��?Dc���u%�8OȜ�u@ɰ>yN�+��_Q,ݹ��M�\� ��G�=Ah����e�>BҰ�� ��:~���x_j<�,o��`4C�)��U���FC?i��"r�m!�O7�j�G�0�zr��ܕW������Y�9:n�Х��%V��@�D(M����F
X��a
�.6rKΕ�T�X���'�:�f�ώ��\�f�}��@I�N�)����Q(��;f�@�N!����Km>UӳfOy��TyN��.������%E<d2�cM6+<�Y��ݤZ<�@z 'a8�+�ɐ��� #�nVDIg�V�4�m�|�>rT#Q$%�����LY�
c,�����#C?
q*ҌM�-ˎI�;{�.=2�#P&!��Ի��h4�����4 �見�c̸h���V
Q�ɷ\�(83v嚗b��p��,C�t`����0d_�I��fĸӅU(j���f�H�,&�a�r�ǔ:PD��v��g9�x���+:f@�C��*o���3��5)+�U���8U�V�J�x 1��
�`igM��]ٸt��(�w�1�`�q���O:���M �T��� ɯo]��� 5+s�\34�Na1���)�ʈ�b$�5$�)��Upܸ:1ˍ,L k"�r�-O
+�"O=)j�w'M>7q���� ��"���R��xp��{cgH�l�[��N?,oѧ��<5p�֝iˀ\�#�
�_"�����]&l�`pҎ,R|��B	;J��q���dɻH��U�V �"�	�B���Z'���N_�H�Ht*�h�RG��9x��e��&���+ �
D�`]>s��i��bRA�&�z���=	��[7��c.<A���<������q���h��$��M�.�#���0�q��H�����~����a��%h�ş4w�^9�9�z�R6+�1P�q��w=�l��G.`��)x����u�P% w�78�t6-ԋfr$�P�%Z�
 � � �TR�Xf'���y��lA��"�a4�T�#�5�%�)����B����T��,t�eY�I�<*�)��D�L�
������r�Q��'	�}��-lyՓ�d�M5�Ԛ6g�	`�����g<OR��$�̯o~��`���n|ͫ�D��N0���f�c��wduH�� p:iHE��M���ׅ1(�m#@��F�n����UJB<)v�XДQ��`U΄����Aj��(thۄ(�xI&E�:�̱�&�C��Q8��պ+��O:v&�)��|�]rf�C (��� ȀA�$�6Q1��C������"koCh��T:��C�Q>�[��Y:D��*�*_�V�R���>_��{�.ȱr�n��E��)'��G��0� �"��-̕�B�-P&ɸ�)���� E��B@╪@�q����@�:����nn8y�d,�5cq�	B�J�P�8����N��HF��"� #�9�����tY��{����6$�;�`�0S^4�IUq�aA@ݳ ���<Y��@:f�e�}:�5��$�.)����K.2ܳ^Oa{b���C�~�{K�ݔiQ�z]�HS@X>$V�0���V�	�$T�8��-�T|dD�O~�Do�;u��8�6�$,�h��_y�'Jڥ�dI6{Z�,q�~:R��Pɦ=HeK�
~ov�!�v�<ivGЯ�Ne�v���0���B�e�sy�%[�y��bSKV��9A6h@�V�J���8�o�RC�	~v&q`ŋL5L����H�:�`���$@�axRF��U�Ω��B='���(�.� �y�� WN00c�Y0O������y��KA0�y�#��=�b����ޚB�I�~�:0;�䑤 �� 4*��&�B�	�.먉zT�E/Z��H6�G�jHB䉢������5QN�|��Ks\B�I�u�J@�� 
$x��H�#n,B䉀^bT����sv!X;?�XB�ə&�8)a�J�"\�qdZ�t�<B�ɨt�"x[�-]"T��� BX8SJB�ɵY�$�B���O�R�Ң���K� B�	Y1�p�T!��V*��A����C�I�c��a��B���{ुq7�C�	1���hn;��3)ݭV�C�	\���0���x���v˖�w��C��0RȀ���	u��%"�':��B䉬Q���R�L50&��G'V>C�	�5�n ��LC�6� }�e��"��B�II��㖫rT|�f�M�/6B�	6Z�E�F��?u�R�1Ww��C�	�z�LL�#�5
�"����. �C�I�InR�����{T��#�рB��C�	��I1ň���Y��H	�tC�I��n��aaL���%�3I�xC��F����مqp�87�R�F����*��\x�ʜ�=��UR�*��v��� ə�R�qO@H��l )S�N�it��W���} ��,lhi��]�¼�B���^��Ҧv�t�C�A]J��ç���I��;��e(�]�{y��A�}��=hw�R6d���`O�0|�l�e�Zp�DܩW�Zp��Laʤ�QƋE����:�0|��"��cf`˥�t|�d�ҟ;�(�19}¹i~�����T��m���WH�A��`�c�x���F���O놩���F4���BnK#t�8�O�1���铸&;�+E��o�8*`!��@c�6M��(O�?]2g �
�2�P�!�g��8%���s7Ġ0K�dS>����>>�lH8�*�6:���j	�����s���yr`�
 ����i�
r)�h@�5�!�%��(��Y�<)dS��b?��t�<G��m��k
,>Z��JD�H���{O��4��蟂d퐄pW���Ǧ���!be� �M g�:?I��"���S6>x,"Ri�(ꆌ��m�R�`���<��4qs�I*A�@Z�Y��O��(�A�O��lyӁiS�=��]J��DO�����i̭8� �@G�/2"��f@�LH�'3 ��F`�؊#)A�π ��r�FΤN�8��$!�J����O$q�'��O��i�S�U��I�t�ĢxH�h`g�W$uS��O�KJ<E�Te�ey��B판!����� ��y��^��A��a����8kT%J���'�x��͈)�rO���ڴ#�Nb�b>E�RH�=Gh G���W���;��<?!P�d�\�#�y��Iϣ[P�h�d�B�uQ�!Q$,��)��֟ Q��n���I�����k�zA t)�m����y
ç��M�dj�*-�%S�D�8pڄ��t?�y�����?q:�c�֟�r2��?���H������$��`BCe!��mm�U�a�ֽ0���jw�\�cV!����=J�� ��4e��ö�U�<��+K0�D���D҆<��SS��K�<a��K/%v�2�,��|Bn��D�<�E��N#޹�ݺ�|J2�u�<�d΂�!4X�#��4��R��Im�<Q`��J}��H.}f�.��<�� z�����K?*:��O�x�<�6� �6�̡E�З-�`4�sOO}�<���\d��\�B��ncn4JW�b�<��.�4وr��<wò	�Ba�<i�n��|�~1H B4U��U�woBG�<q��_(!�ƍR��+�荊E#�@�<Y��f{�aq"��`�Y�V�~�<Y�ì�~�ƨ�6�8P�Uy�<����(�\�m�{��q�f�q�<a�$�8B5ʬ���|xI@�Nm�<�2(B>&��چɏ�Z�S�j�<���:ߒy�ţG�,�h3���b�<�Ҁ�<#���$/�)(��
x�<��(QZU�r�Z,R@��l�<1�<qx�m:���wm�z�@�s�<&f�%j ����H2�Z�x'i�q�<�6nLZ�:���Y*{��9T-�b�<�&#6�pTn® Ң [�J�^�<1��;W�>�/�}��	��A�<IE��E�8��WѸ��!�@�<	���ZQ2� �j�6�:�2���~�<�V ���s	9�Dp*�L�{�<�T%Ӹ����q��WϬ�y�ɍ\�<�U��N9T	�d�#V����r���<�r�J�:�����εc�䄡�ɇa�<Y��(l�Ƚ�����H���H�<)#o��� �3%T�A��P|�<ٱN\$+ \��,==z�{c�a�<!�H�0{b�RbAC>$�`�*�d�V�<y�h��� p&��nDF�R�O�<��OG	$A<)���d����VC�<�[9l줐��h�f�dy�AA�<�Fm���`C∉�$4�Ak;T�@{���m� �B��Jະ�9D�L3�D��bܡ�r�A+8�@�"��7D��y F�.(��e�[2���f*D�D��,)H�`Y'�޿�ּ��H*D�\��"�&%� �j���#?pX͘",D�$P�&	&h�8\�� *��
�>D��ȕ�\�a��V �*|LܐP2�<D���Am�@"JY��CS�l_|�b��4D���Ù�d���s����x5�e4D����� 3�D��6��E��"��4D��y�H@x���2;B�|��n1D��b"�A�t!�s�I�8�p|�@�<D��G%&���:6Lχl-�q�5�;D��*&�ںL�
}Un'�	�Ҧ%D�\�7*�fd�Œ3L =4��C�	>D�� �����ߓA�R��T'�����"O���I�x.��!�a�L��e�ȓ@��p�jAj��ٹ���>�����E�n����>{�|��Md�ȓmM������8"���6@�#L�ȓ
AJ 8��c2𥸦K"S���ȓ."��3C%����!C����8x1G���u 	��֙%�J��ȓ@T �M�K6^��$�`��`�ȓ�&��׌ЩU���ՎcU��ȓA�dI�䀅k8�%��Q	3ćȓ��lz�Fͪ=:���a�*����xzJ|8s+�t�z	ɔ�Ӛy;��ȓ9����l�uҚA�c��"d����1����@��Y餤]
�X��ȓ�����G+f�#�`�@i�M�ȓT�`�X�
�Z}�pC�$N��i��WN�9D	�e��%"��,�b���s��`��q�p
��Y�aA�B�I�O���!�g�DT�Q��"4ߌB���+�E�(+p�KE˜� e`B�	�dո9	�&-o���@�a2
C�1s~y&���a�����H�'�C�I ��eK2l@�=�j�rSH�|�C�Ʌu��-Ӈ�B>dt�t ��M�?�C�	�t�H=;p%����o���C�	�ֲ�S�o��X7(y� �]?�4B�I�S�&Lx4(@�S����"��*nV,B�	�Mf���0�SFM[].C��-R*m󂝛� �D�BC�[���o��[�\�#�J�U
C�	yv�8��EA	�\$+�.M�K|�C�ɤY��`jC�;_��Y@��"4]fC�ɾ-��E7m�^��qG =�:C�ɍC�����^�=�����D?&�C�ɺfB�@�Z1�Mj��C�C�ɍ���2�gS6:宸����L'�C�	/l
�R�߭_׼<
'��[�C�	#%�la� 
O�@���!���Jn�C�I��n���ЀJ���&����C�	�J��80�AJ{:-�>A�VC�	�5~��r�ʘ�M�A��C�>xC�I8��e*��4�!cIHa�VC�� �r5p��Ŝq�X�0c�Q7*`4C�	���YV��&"zXI���f��C�I)0&x ���9:]�R�РAB�I�DOx��coϢ"�kP�^��B�	�4�4�P�g���Pӫʃ5�C�	������(d�a�GH�91�C��d"	�`ʛM�I
��E%s��C�ɗE��I(/`QA��W9��B��0(a�Ȑ\Q���d����B��FA�(��킃P�������7��B䉻F�4ukq(�6t�x�$��)�.C��-*���!qJ
:��<���	:v#�B�	=U�V@ҒV�VTĈ��	;K �B�Ʉ�΀@$Ö�]Θ�0�Y��C�ɴ@I��� �	Xb����8?��C�	&�"�h�i� ��B4�qhJC䉋$,��A�k@?^������@�o�~B�	DS>p���� z7�%���%�hB�I��~��w��!FIpųr�.6�bB�I���"�E|��E�2�Y4/u(B�	:h ��Jx�J%Z���,��C�)� �e�!!̦��9�ƫMv���"O�"�$I�E�l�QH�',�TT��"OP8s���J�N�Jh(@����"O	�(CL�%��]�4U���"O���E[�	\N\�A�I�I��[�"O�8�1�1L*�I��_9|Q�@1e"O�i��'�7Uw
���C�xj|u�`"OH�hv�-a����ĸ[�(p�"O�I�%�%w�<Jv�o���BF"ONᠣtVB��p���J����"O8��iQd�TJ7C�5P�$�Q�"Ox�H�CGy�([d��{r����"O����Ã~tAZ#�>��"�"O��2f�@�`���M׃b�0���"OT\i!Hґ\�P!s�+�pl��"O�U�O�(jɢ�
5�rD��"OviS��)j�:D�v	�
st��"O�� �zJ�8!q�D-!`��q�"O84;C�
�#�0��uR�h�"OV���!Ӹ&(�N@�C�]�"O�Q�UAA�zP�+�"�˰EKg"O ��@E�s��P7��|�N@�"O�����W*D)HD v�z1b?D�LJ$��0�Jp���[��>�(<D�d��-�/:���PBD��7�0��ad;D�Q��H�i�X��!�/m�.�!���)�����\�>�t@eh�>C�!򄎽G��]�V���
��JS�a!��!���B�"#�:�0AJ�U!���n~���) �% d|є	S�+-!�H���]�!���p{Gɟ�B9!���9l@y�������h_�!�AY>�9"Ə�=���{�ӸV�!�݃�<��D�4��A����!�$M�k
��1�R�u�|�����!��ɮH����	��2x꼙A�\�h�!�>6>h5�� Uf���g"9*�!�dD��I�u�� W�.urcL�0d�!�DL�|�u�OA<�����+!�$B�lJ�����N~��ٕ���8�!�Y�p�Z�
)hVɁ&�o!���CT��`��49\!�A��V�!�v�t(�qC .V ���c�*�!�$ь1Jb��E��i�LW�N�!�_� �n����>�
��JU�\�!��R}�Q�����T��)X�y�!�$*#��O�)��p�A�7�6D��r�)
7�l���L�X��;a3D�̋G�[�`b0�-8��q!�>D�Pd���P���B�<�کc��2D�P��A��K���ւe����D�1D��;�@�n:("5�5>6�y ��0D����!*&D}�����������-D� ���	<t���q�n����a��-D�P��u�L��#L5�A ��8D��!w/��P{��q"&Ύ"
!�5�6D�H  B�(>y�tϋ�e��$0�.D�@�'ΆI2��" �'q�'#8D��h��ۅ}^9P��!���"�l5D�t[��Z���PQ7�4LT(ץ2D� ���H�A8�M�$//8�A#�5D��ӪTv�īE �On>a�#.D�Xɶ���}Ȫ1�I?0�Xt�$�*D�4�S&ΘC�Иi��
�i�+6D�� |К���T�8�zT�ҡMĨ�@U"Oz���Ƙ4Ϧ�c2�X?�8�"OB)��e�1��%+W�A�c�Q0"OB� bL[�n�1�%G�U��]�"OL��MܗA�Hdj�/C�~T@�"Ob����nߤU�F`��o���p"OF|�ī�E�t퉡OFK�dT�"O,$9U����e� ���%�
�e"Oz���i/��5{j�"\�&,�'"O�u�Q��,/�`x@Q���I�*]9�"O̰J�꟠RVxEA�'G��d��"OƑ�*��j�9Ra�Nz�R@�""O�呓�"�U��+ڎ!w>�y�"O��   ��     b  �    +  �6  �B  �N  [  )f  �q  �|  ��  ΍  Ô  �  Q�  ��  ׭  �  x�  ��  <�  ��  ��  Y�  ��  L�  ��  ��  !�  �  � � � !- �4 �C qR �Y )` lf �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;���ē]�.�X%���tM��aF��m���d"O>P(DǄ�.���w�G�AB�"O��UjGOV.mI%�]8Z�y�"O$X�Q��L�"c��=�� �"Oe	���0%�^���a  )�6E�c"O������r�ꑺ��O����e"O�%+�CdeM��1O.̩G&�eh<�E�ߒu��P�L��SF��h�]���	@X� 4d�N�F<�bi��E�Uzo+,OpR�O��dW�e(�EGߎxB��ݢqĊ��ȓE����E&6zn��8$$$��A�<�<O&�s��E�π �Y�P���.i���x�ЪF"O�)��B,]�X�S�b	|9I�O�=E���7` 
`Ʉ�F/e@^��G� /�y����`1�G�A?]���A7"���y"'�XPq�'T �W"���>!�O6�zee�82q��[�2f(-�3"O�a�b_b����E�Ie6|��"O(Q���r�F�A�E:<�|�
�'T�9A5f�cG.���ZS�bU�'�^�Ӕ����v!�'O��Y��'�����$r�LI`f/ˬB�ڡ��'���vOSNxX��d� 7�(���'�S#�$]墭�t��>#��e�'Z4݁R!$(\���gA	l��K�']b�qH{�t��gӣi⸋�'J� ��-�J�Jw.��H6Ű
�'F��	&E�J�K�e��y,�9
�'5 ��uoV��P�
# RA�:��'��-;C�P ��hY���3zR���������9��3� H�8�Gh/D��aO@�k���4������Ĩ,D�`T+��QB�"[Jh�����+D�X*t��(^�R���F),�%a��Ot�=E��C�#���IU���] �E�.G!�d��q�ɂ�!�'�~��Лg0�f����G�U����9����$D���S��&��d&��ɕh#D�,)��Q�4�(�1.�BG6̪�@ �SK�#"G�_�F�zY�#��+L:���IC�<9���@Z�(� bU�x��!�K�w�<fET[n��#��B8�����r�<�p�B A_����Lԃ4J�e�w�<i��gM�L���;?��P!���o�<!2�L�.a�3���EQ�P)�ğo�<���S i���X-/l�����h�<ѡeˌP}�K�o�(Ejt�����Y�<2mX7#�B�G���&�h%s�'XS�<QB"�v�J���"E�RV�L�A�VN�<i��J�J��� �M�:y�)X�Ǆs�<9���"h9��̀$(���s��p�<)į	�� i`g,���N!��_l�<U��Xۮyp�(?1���%$F`�<��d��*�����!��b�~�K'A`�<a�D�E������8���k�PZ�<ɴ׬L谜0B�ƴj6|��O�<�dEU#G�[�Ɔ:3p��l�a�<igF�I�� �c��U*F��V�B�<��T�H�۴$;!q���4�e�<y���{��Eh��.pTb$s@�XG�<��^�1�����"��(��$H�<�5��sLt�Q�� 5rUP��O�<��w��<su�S�)���(W��d�<Q�n]�B/���fؔ���C��w�<�֭��4]�4SG%#7�4�m�<)���QtHܻQ�
j���Z��i�<Ae�Ջ|�(=Sd�w;Z�rA��e�<�u�ԌbV4
6���'7����l�<AsJҼq�aSD�5 ehD�s�<��L������HQ8Ny�48�� j�<����Nr|��V^�{ �#���q�<�o�9W#��#H�N�Y�w�Lk�<Yp��Nj��&�q 1�m�l�<i��0�hq�g��l�,�t��T�<��i��	��H1�K2�nAgZT�<� R�s���'�ja�ԀJ:;�8hs"O����&�bљ7�O�I�x邀"O��G�/J�AW�K�aQT"O��Q��"��(1VkKN���"OȤ��Ĥ�L��E+�8<�h,`�"O05srcJ2+|5�	�S�I�"O�0�&��2A^Qko�6z�z�"O2��D�%<I���B� ��ȡ1�"Ofܪ6G�%Б���S�*~]ڒ"O�Q�7���DRn�`͘��,2�"O�9R	[:^Vpx/���L`�"O$�������(�5�$j�ePr"O�MX��P�[�X����YEn�T"O�����n֜CA�7cA�EÔ"O�$8V�\Z��%h�oԚ�d"O8b�ϊ	L��г'M%r�81��"O��*ӢA�/�����O�%��h�"O4ٷ.V%f�2-��Q@��ˆ"OH��C.��g���I�AH��P���ȓlj8sQ+Q��q� 왋F�|��'E�` �Mh��ţ7nݢF�h`�'�^,)I$j �sꅇA:T@��'92ᰧ��-D̄ S�>4�P3�'K0��*8��8;����,��'���sc���O��]�"'ָga0�';н���!Vr8�0g�ݩg�Z,s
�'F�|�Q�B�dy�C��3;��Q�'�ha������x�
�;9�0��'nM{ E��~M����ə!bo�$	�'�0��#��<���a�`ިN;����'���E�Sd4���-Q���1�'+�=�Fd����p��	Q+8� �'�����	#:%�4�\4?.��	�'J)3OJ"X�T	䏊
�`%;�'��%���5EΈ"�`�T�����'��Q�a��0.2� �ԅK��d��'K�K����4K��`$��2-r@���'�p�#�6�t`q�V�hJ�
�'#zD
���
��j��5�ĵ�'W4�hC�pA�E��H�0�����'(t���R?�V�:�g#1 q�	�'���P�J�J ��A�(���	�'�Pݪ��FA�iB3-�	��|�
�'��]3��ӭ9�����Ʃb�J�X
�'�J��#НÖF�]��t{�'ִ�J�)ncH�(���V�~�Y�'Ǡ�3��LY&��p�Q�TѾ�S�'�v=�D��$<����)M�8��'�x�� (f����񨀫q��}2�'<�17E�-B,�0��Y>�}��'g Xt�ǿFB����ם����'�%!�+F�P���p@B�	�L��'�t}#˞l/�؉7�
V6����'�*��e�l馤P�FB��'��%㖆�$]ad��6�O&0H�"�'��(T"�.7����e����4�	�'\
�y!�B���#�-�
p*0�'�F�R��Q?lӤ�"EP�~�Dq��'�~��$Ƨ
�:u�T�oQ����'���b��M/YTf���#�=_�Dp	�'�R��`i��w^�䳀�GPWb��	�'�L�k%�
�!�EA�n��4�rM!
�'}����X�IRR(��'@q��'������t+%HH�4bHAs��� x��'̔3�����؝fb*`h"Ox�S���8���P�?_��� "Oܙ��	8��$^*5�6��"O��@�0�!RH�:~[eCF"O��D�	?͊!�`�̡X����'���'���'j2�'�r�'5��'�",�BO8n70�2a�IPN���'?��'|R�'+��'U�'Zb�'1Н��%]>D��s��h�Y�'*��'(��'B�'r��'H�'o���Dě�A;�pp�]�T����'[b�'���'��'-�'\�'Ul�@���(=�d0���ux��I��'1��'T��'IB�'���'rB�'t�ADD.8�$Z���;ܜ�ZB�'i�'���'C��'���'���'gnj'�.##�Аr�"�tXc�'���'��'R�'Y��'���'�J}PT��%+d��X��-vx����'d��'���'7�'G��'p"�'5vp@ta\#fM��A�̕z ��p��'�b�'MR�'z��'��'
r�'¢YK�W��3�Nʐ`�NDa��'���'��'��'���'�"�'�Vq35A��&݂j����y��',b�'�b�'K��'�r�'�b�'"$�f�ZX��`�K±i�`���')��'���'���'�b�'�r�''���
��e�D|J�
�+H0@���'�r�'�R�'�B�'d!~���$�O&	���F�����gB�f���Qy��'�)�3?邵i�ΝiSH�2�8��J�&^k�ŀ"�G���J䦩�?��<������@.�>Mp�*sL
�D�<y���?� *�M�O
擓��J?q���'�"��C�\#^�X��,��ß��'��>4f�F���9tC����lzĂH��M�@�_s���Ob(7=�h�(vO�.S�<S�i��LmZ�{��Op�l� է�O��ڱ�i��D�� ��cF�,�J��o��J7�`�����8�4�=ͧ�?��k��>�¤E({�$�3����<Q(O�O n6A�Bc��h���7u��IA�M�����L!.5�O���'���'��>Y�Ej�]�`�S�{$5�$@i~��'�zdx�k	 ��O�x`�I ,�RL�=b®tc��%fd�8�.+���My������$WA�4�jC�6�v�xB��I��$��q��3?b�i��O�I
�Hlx��+(���KW�n���O��$�O�$sRKo�j���d���t Q S�z�XT�� u v�T�@�����4�6���O����O:���
DjR+�띔#o���,�(˓zK��΁�`�2�'�b�O��䟠�q��*)��C��x�ԍB$��d�O6k��D���K4^��j�
7Lh��Y�F��3�� &��$���Ia�XPV�O�˓���b�^7<]�`zQC�3a~00����?���?i��|�(O�lZ9\���ɍǼPy�fۤ%;@�E)ҹ����I(�MÌ��<���M����a�����(6H�eF6E,�\x�
�'�M{�'�� ��S+�����P���<b��f��8r�Ö1?���͓�?���?���?�����O!�8���,v���`&\rt�a2�'���'t6m�6M��O�oğh�'�$�hQ�5w$����գU��8�1:OH�D���o���Q�-�|7Mu�<�I+	�X(��ꂱ�����EJp�)BY�
��*Yn�	^y�O���'B���^�B9���T�3� �A��Z���'��Ɂ�M�1�K��?1���?������ ��S����ܚic�9�t k~Rl�>�%�i�6-t�@&>����8H�];D�\	%h� mk�����B���'M�����J<*��+\�O(�#��
-;�\j�C^6$�u�#�O2���O��O1���G曆
́FaP�ĩ�1�|Ҡ*��na4�'�B�c�F�?���A}�ef����㫍�a��M
�b����˦�̓"?"l�<���1���Fi�؅�'p-�*MPj�h𠁈6R�:�'��ß��I֟L��ɟ���G���_�$�� yb-�"z$6	H�n@�j%�7M�N����O��$���&`lz�aJ�N�Q氭��%�'E�NA� �M{�im�$�>�'���5Ξq"�4�y� �4	� e+���'�j�
� ُ�y�RB��T�	�@�'��i>5���
]�q�� �.pk��p��|�b��I����Iߟ��'�7킯w��$�O\�$C7�"-!��6rY �8�̕�s�>�2��Jq}�i�jpo��<1�OD���"Y�-k��HUI'$mĤ˰4O���U�2D��{e^�����?��W�'l��	�]��Ac �='ɘ�v�ۻo�&�����8��̟�6�+�'�?�D SKͪA��?�h3�J��?!D�i�����'���c��"�4�f���Q�4�*�&㒿Vnu�e8OZ�mZ-�M��cy�\#ݴ��$��0o~i��'^�r��G�^w�H��l �ue 8a$'�D�<�'�?Q��?i���?"յ$��P�lܙcuҡ	��������=Q�*�П<�Iџ���q���'�r���
��3S��+���0�G�<����MÜ'��O����'�R�e��c�T�I�	|4,(��Yj���Ox8FD�?�6�d�<!A .wJ�I�Ӕd����Fh��?���?A��?�'��D�a��,�韄!eb�'غ�CgGD�(E���؟���4��'�X�2T�Ib���dL:�j�iѣ-�<�`�JJ��| �Nr���Iϟ����Q=~�T�3?�'1~k� p��v����r��5/��6r��J'6O�$�O��D�O����O��?%Re�N�`Jc%->��a"��h�	埈*�4I@� ͧ�?	#�i��'����-J�W4$��f)� )�^4��9O��kU�6ie�N��C9Y�V7-e����l�fy6��+g|��r�L�|9Gc�B�h�	[y�Ot��',"c��S�`��f��s�X�2A�@5f��'V則�M3E͎��?���?q(���2�Y��L`*�/V��xh ��|�O*ul�;�MS�'��O_�TD��4�0���o��sq�Hg�ǿ'p�(B��:[�H��O�����?ѥ.��=ga4���ٺ��AAg�)�����O����O�e��҂��S������u���?4�#%˒z��m�s��|x�OZ�o�D�j��	6�M�M�-Am��P9)���Ű0ٛEh�V̀��l���.B�hy���B�,O�P�ݹK�,Sv�L�
�6I:�;O���?1��?����?�����I[�XЌ
�%Q�a�΁W��7�!o)2���O�������<)1��y�\���9�H�br$���i�P�7m���	
����4�\�I��^�%u��牨!`�t�����{�ZMW,B:<5.�	�j��ݙg�'�"$'�Е'���'Z�4��҈~J�� ��.��'m��'<bY��iܴV-�	��I�!'0[1�0U���.�:+���?�Q�0I�4!��f�O �cX{��^�Y2d%Ԋ�c���ܳd�ʓ7�
�.p��'?�Y��'����-	J,��$�c{`0�A�Вp�^,��ğ���Ɵ��Ih�O�B߱ =�a��h	��䝣)B�|�Z�L�dߴ���y'���l����SoP>'��*feԆ�y��j�*nځ�M;�%��M#�'U�YbdL-�S�l-Ԝ3�P>Z��p�G�j��d�А|B]�0������������͟4R�,�3��I$��� ��\�d[�X�ɫ7�$x3��O6���Oz�m:Γcp�k���/��8V�9s���V�x�ܴC��.�O���)���U�6+�M���%�לB� ܲn��R@ @��<ip���j�d��䓀�Ğ�cO��I&��`�~IH"��Tj�D�O����Oj�4�H�s�֪n���O]�X��
GO���S�ͯou�$���U3�v�D
J}�#f�>�m�&�M�GLVH�%���w5�2��G�lon���4�y�'�~Yx�-X�?]K�_�4����Xg@O�#����N� z:=��#a���	�����ҟp�	��(������hAlh1įD�/�^<�q���?���?y��i���4�'�7�(�D3�=h�O5O�4� W>C�l<'��2�4����Ok���b�iJ��Ot0#a ξ����կ��p�AfU�"ޠ��XؓO�ʓ�?���?�����������(�2�1��� ��?!(O��n/U����I��h�	X�ԇ���5���&�ڲ����$u}�CeӺao�$���|���>?i�0JJ�����D�YF����c��7��HWV~�r���0���>��]p%
�*���0U�ˊi�P���?���?��S�'��$Tڦ9�S�K�cy�y�
���h@
En�0���'C�y�L㟌��O�m�<:Jd�@��
i��0�H@`"۴��(0��?O$��źq"�0�'I��n�t�6-$$�U)��R>!|x}͓���O���O.��O@�D�|��dN6�콋uo_6M؆X�"N�`V�&J�+w���'�r��̦�L����ۨ~�X��E�7J
�I�ܴAC�v�?�4�����D!�H|���:��kVJ�!&!|T��mRAI�P�r�(W�O�m�N>�,O��D�O����θL4��χ���{��O~�$�O����<)��ia�H�7�'}��'M�9��Φ ��7*��f4��A����U}�"nӀ�o��McvU�l�cd�A�|-�ׅ��
���Gia�����x����@��p��i�'���ZJ�Ξ֟x#��Y�DJ}��#|�L������	ٟ��IƟ��I��"����M���t��!,�H82��"WFH՟p
ڴs�xP�'�����'��	���I�m|0����]2Q���j��V8���MKѲiv�7�G��7�<?�#LC��I)YPH�� �*����c��J���H>�+O&���O���O����Ol�`��x��[�j�؈arǪ<�p�i4(ES�'PR�'��yBKՉ��3pA�9-�ti�1KMb�+��Ep��O1�bu2���؄a���u����iR�n:���PB�<VH']���lZ���'��ɅY�=2��g���H�Â`�P�	ȟ@�	؟��i>!�'z 7�')p*���Hȼ�*�A^9wB�Z��d��)�?�Z�X�4B�&�'0N�bf��;J$�x���R��˵	��p"����haw� ��$�)��u�@	S�9��� 9�a(a��<9��?����?����?ي�D����XU\�k�P�����=P�b�'iB*v�쭑:��������&��I�A��=��yw��uM�h��U�<��Ov�o�	�M���4�����4�y��'k�\�3�ŧ-c�@)��8�4a#%؛M@TT�	�2)�'A�i>���ߟ�	�(@8�e*f��|�f�_MA������'S7���#!ʓ�?A*��zd-Ѳ>5�R�f	�`������l¬Oo��M{�'��O#�d�F0� ��O�?HKb��t�۶|�n��.ɧ��\k�O��i[��?��F)��y�șag��C������'X��D�O~�D�O
��i�<��i@V����/&vq4�'F)����o�	�r�'f�6M$�ɧ���ͦє��'b�V�`�oN	,%�P8�Q,�M�v�i � {�i��Đ�c6&Ô
A���a�j��� ���$ �Y������4Jɋ2�i���'%B�'���'B�'��${��4Y"��<êXsg�^)��(zߴ>+�\����?i����'�?����yw�S�dL�j�Î-wr��r傅-�0�Dt�,�ny���:��rjʉ��4�yBH��C�\�B#&�����%���y��E�r(�	)_�'s�i>���T�J-x.�,���sȳA���	͟\��Ο�'.�6�LKap���O����N����$��oB~��#�\WQ��p0(Ov��|�r�IA}BaO�.$8�'���V}��J�/�y"�'�z���5R%�\��O
�	(�?�u��O�]"��]���1�"TP�؝rS-�O���O���O �}�;l7ްs4��.d�B�h4CŞ8c氫�K���[���$˦Q�	R�iޱ�D�]:r-�X�PESq��U�p���4
���'/�`Kt�i���O@��a炩|��N��eu�Y�E��x.T����1L�&RJ>�+O����Ot�d�O����OV�p!�B�NѤ�����R��M�D'�<A��iu@���_�d���?��O�F� ֘�	7%԰l�Р�"���7��Y����mӨ�`�S�?���.p�0���?�x�JF7.�`��g-+R��j\��規�O� �O>�.O�iYf�v���At��6ft�	ip��O��$�O2���O�<$�i��$0�'sޔ�F�iRV���j�3t*M�'��7+�	���	��Q��4�?��� 8\�ȉg�x��%��NR/e�H�ٴ��d�:n�T�����ȉK~���Fg.̑�%×vB��+SbP�q%��rٴ�?����?����?�����Օv��aA��7tv� �KN�y�'��Ad�8�i����a۴��_�LX2cJõde��%�]c�L`M>�R�i&�7=�ra�Jp�~�Z��T�K/)Ȭ#�"̬_t�X�D=VD��n��u��'��	��	ܟ��ɜGO֝�2͌���Ⴞ~�8��'�R_��*�4>��0��?�����IR�}�a���2¼iՎ� 1��	������ ۴���|���U?�$��Y-1���!E�pjF������k8rр҆��D�*�9p�i�6�'�̨!�>Po�İ����Dߚ����˟�I˟���Пb>�')X6퍾X{�q;�G\�Bu�h˹Fީ����T1ܴ��'�:˓�M[��$Y�����A�#�t]�wi�jO���'���᧰i��d�OT�˵��K��ԅ��C*�t(ӌ��B�8���̬>�d�<����?9��?���?�*��y;&B��+Ք���FӒK��U�b����4�z�d�����'?�
�MϻI�1����S2"i��1uu�T�'盖��O��d�'� !ײi�����>Kn�P"�>Ҕ��l ��
�����i���&� �'��'<޸1������(���	p��RE�'_��'w�S�!޴v�h���?���ix��h��_�8xa3�	�K�y���F�>i�i��7�/�Ԝmܒܘ� �f>|1�J�f��O�-�#X�%����<1��v!��oZ3|���c����퐼���Xg
0rb�'�"�'�"��˟�36�I���1���\��e���Y��$3ߴP�e�'�7��O@�O�.O"+i�b-ȱB�B,sf�K9-��$K��޴�?yr�ǵ�M��'��c�Jt�YA]wH�<j��5oDR�jW'�,�"]�UϞC�Ify��'���'�"�'J���*&g�Y
�d�IF2]�`�Ήm��I�M��o�?����?AJ~����L\�pO��sMN�)����6N։2 \�Hڴ_��6O������O��9���#F��[��Y��Ô0
��{���:��G%crd�|�	ey2�M�h( ��&�E�*včrQ����'�"�'��On�	��M���?��lJ:�|�rb�;@�*� �O��?	$�iQ�O�$�'��7��u�	�O5@���r�����`)���!�P���̓�?� ��2?�~�)Qw~�OM8��,1 ������!1�"_�p�Iß��Iݟ$��ğ8�	l�'R�s�45D�Y�F*`�c�B�-�?!���?�4�id渰�O���e�.�O�x�$�g��@bW!W�X�Īh�P�'8 7�B�]���n��<a��%��ٱ��0:�S`B����a0M�)?������䓄�4����Oj��D�?�8����!�P@FF<����O����Fގy��	�ԔOx~5��@3izL�w?-��]��O ��'s�7�Γ�ħ�*EZc�$}pQ!�e�by�� ʸYP<P(e��Y�H�'��DI�ϟ����|�b����l�P@ߙ9���!�ϐ[��'<r�'*���R�̐�4
����U��&X�6`BO�8�`�"�"1}Ag��⟤�O�lZ�|�$��!㚭mB��X�S�����421���
Л�3O*��Gy�����f���"�.���A4r����WC��������O:�d�OZ�d�O��$�|B�.���F�h0n���IXҡ���?����?i�'����Oz8lz�ɘCQ^S�P2���.���pg�$�M˖�i#�6mW}�O\���O�>����i��~W&I�4mG!h����D��~7����&$"�@����<�(O����O���r�J2z�2i��� '��3Wm�O����O��ۆͻ<��i.��W�O�2�'��9!��өVh�H�w`K#"��C�|b�'k�����n�dm�Z�DH��a��xx�@�q�&!�a�ͥ�y��'W�\�(	��$�P\�p�Ө"@r�C�D��F
f	�)Q��A ��W`ʟ�IߟX�Iuyʟ���g?�*���.v,����˫R�q�� <r����ɦycCm^������0��wyr�y� F�u] `�ڧ@�I�U폮�~b�i�7�S㦵2bNզY��?֨N�|r\���z�? <� 1C�(� H뵦{�\���;��<����?����?���?y��G�7�R��R�K�fRze��L�5��d��5����R���ߟ\��?��IΟl�`��+�$� ˍ��`��VNC��$�Ǧ��ش\ޛf �' �2�b�V �ȸ�&3���4�޾o+Z�`/O�@ w�ד�?�Ղ5�d�<	���4E~��r�;W�h�!�Ƶ�?Y��?��a���AN͑���Q��	�D���?�"�M�\8�ͅ�B�dP±������@�i>5�'j 7�NϦ%��4�L�DB�Un�r�Ŝ�����ٚ�MK�'l�Y$��!J����?��Xctx)�TÓ/��TBUOؕ#m��'4b�'���'M2�'��HH�u�^�Vyk"��t0(��>Od���O $l9P���)śf�|���5^�v|�QJ	�m�0�P�և;��'M�6m��e�	�w4�o��<��IW2��Bl�)#�$�S���Tp޼ �%�8�N�n���'t�����I����	�_m8E��R��Pd9�×�?�~����X�'4�6-��4���O�������C�#K4˷�DE!Hr��1H9��7������ܴ���|��'"��%���R{�;g�< �h�����"uGT���gZ���d1Ŷi�r�'�(p��ʌS#�Y����F��Hcvi�ʟ��Iٟ�����b>��'n6M�=mQ�("�KN{�eچ�M$ĝ����ܴ��'�2�1�����Q���ڰˑ�#Q0���"=vy&7��Oְ�a� ��ӟ�G�$Ef���>�剼DL�ԓ�G�
�|t�q�>3f�	|y��'��'�b�'RT>I��N�"s(YU"	�+u�l���2�M���D�O���;�i�OD�lz���1d��>��!�~ƌ|�"��M[��i�v6�L}����ԝA��4O�|����	�la�acժD��!�:O.p�%M��?��-(�d�<��?�i�~�5򕥗.)gµ(�E(�?���?�����T���3�oDy��'a����U+�� 1�Ů�0�;��'�'=��?I۴�yX�dH�P4w�("���u�42׎|�x��3"�%�p'�s�2���1��O�e��k����Y`.��0��2#�I����?1���?���h�����#ipͻ�/��\䬢cC5:"��d������>i@�i��O�N�)���@F��y=;נ�&�d�Φ�+۴Dě�M������"v���f]��Q�����W�yT��C�>VK$��{y��'�B�'���'��'�2�vꞘ�I[oP�pk�#W%" V�ntx�
���I܌��g�'
��d� }!9O��*5��>6�f,��g���3v�8P��t��O�m���M{�ዹG���|����F�D�P򬰫�b�2�&U���L
=��A�6Ɋ<4m�I%3��4�G�'�д$�8�'��s�ӭZj����bĘ �Jۑ�'���'h�����_�����r��O&i�WM�$/I\h*�̵y��T@�1O�%n�J����	�Mb�i��6mP>\����-GvƔQS�̵\��H��m�&�5��E����{K~���A�ե �F�a�BK8s�F�"�9O���M����?���?a�V2���e��|ju*�&+�۰��Xr�)�V���<I��?��i�ͤO�An�j����6!A���BA+,#~�P�����ʦ�8�4�� ���MS�'p�#�5��8ScȚT�*7�^V%HE*�)�Ο iђ|�Y���	��8�	��,�h���H+r�X�;�d\:#�ȟD�Iy��o����'��'��ӏJ���K1���9@�R���"5(�{h����M�e�i�T�$-�)�98���:��y�'&.�TB���s�:X�W.�K����b!��Oj5�K>�Ԯʎ�������7i� �C���?���?����?�|�,O�o1XDة��ӻx��Ȃ	)8
а��>1&�i|�O~d�'T�6��11�p� !ݙl��{����e��o��M#s�B:�M�O|�6a���b��<�k�hU�t�D�]��Y�Ҡ��L�'<��'}b�'���'w�Ӱ?|5!k�,K���	GDd3۴ ���ޟ��	p�s�TZ�����Ƅ�I�\L��H ʜ!���؃Ik�ir�d�<%?����Kݦ��Y��*�	��=x6D�d�&��T� � �O�IO>�(O���O�D����d�Z\��Ad�O���O����<A��iؾt�O��d�?kh�T�!� NT�kgE�r"��H��Ob]n��M��'3�ɖ��@�Ԥ8���0���%��x���Sy
A�T��^�Qib��֟,�F�&Mvl@�C���,�r���<�I�����pF���'Z�H�s��hִp�� 4|�d�'�6�:����OFymZC�Ӽ'�U�k�,R$�>OD�@��<���ijb7�Ӧ������'�(ʱ���?��5,T�Q��MȕA�~�d�"ic&��'���'[2�'�2�'x�+���}�B���ѯ/�"ɂS����4]N���Ο ���?-��y"ʑ�4h����䎣a��x[b�P X[*�7s�&�j���	e�O��ܐ��
.:����,��\���x�H8>��lJ�\�����  ��+Q{��@ybN׋@�<�j���e�H��k f�B�'��'��O��ɰ�M3G̴�xt��]������"�Z,�1x��
ݴ�?L>Q�[��	̦=`�4M�
�Ғ�(5�SaB.k<�B�O�%�M�'ya�7]��U��/P�	�?e_c�����ٕC�d4�K�<(Y�-(�'���'�b�'�2�'���)q\D`�A��/GE�4P`2O���O�nZ2e��|�v�|B��<�@$���DdX�3����$�>!�io�6���8hCB`���	ܟ�+p-/� .�K5��<)BH29�~�������?A��%���<y��?����?A�l̻]�����gV�q���U��?��������y��Oh���O��'R��R��u%~��6l�2cvb��'|�3t�F�z��=��O���?�"�(Mv�� s̉#R�t�xe�S;rL�@�U�	0�f��'��BVٟ���|&^
3|� �S6�X]��j��UNr�'��'���T]��Aߴ���꣍�Qk�!���$���7}BFo���t
�O�qm�:�p�цK H����d1�bY��4 ��)Y��6O���V]fT�'4���I3 �ū�?/� �3n�8w�`h�����Ol���O��D�O^�D�|�s��;x��|TV(%Z�C
�5���%V�y��'e���'�t7=�"����B�>���ܱ����e-J��p�4��Ş��x+ݴ�y2�M�CM�����9.:��)��=�ybd[�~c�+�49E��O�ʓ�?����49��f[+^F(�s�WC��T����?����?!.O.�m�@j��?��b�0�@�s�űe�FY8p �?�I>��Q�|��4k%��O:�/���Ս�7/�ܭ �(v�8�Γ�?��Ʌ�:���t����$㟌��@��d ����2Dӥ�TH9�L�$���D�O����O���5�'�?!�fô/T�t@��$��,��S0�?!Ҵi��9��'|ҧnӊ��]=oy
�@�B�K�����V�ɀ�M#��i��ɚ4o���?O���֧^�\�(��(&زEf/q�!V낽:����5J"�Ģ<ͧ�?A��?Y���?	���
(�/�`�7gպ.	L4�'ɺ6�������O0��;�ӓ\(rE��c�3�<x��Nvc8��O��l�	�M{�'��ON��'��h�`7%�h�'C�l�ؐ��*�vѻ�O���7G��?�v� �d�<9���'��m�΋t9N��b��?��"NA3a��?ͧ�?)�'f �nŝ[����e/F�b$��$)|!���p��Ċ즁�?y�Z����4ٛ�'	F����Ʃ5�v�K���׺		V(�X�f9Ob�]7G�v�0��Gk�	�?! Yc��<��0Տۙv���ا���y��'���'�R�'��	&
�T��6	����.ڀ3�t���O���H���3�r>�ɩ�M{J>��-
�T�j[`|Ӏ B�!ڝ'��	æ��ش�?�����M�'�R�[�,2��A�CY�TQ授4 -�B �㟔�u�|P�������ϟ�᷂I�r��Xqت:���XL�Οl�	؟lQ4E��6>����I柈��՟���|
���,6�x ��N7cW�paFU~��>4�ia^7�k��'>-��'���'�2j@1�*]r���b!m�/>>P�P9?I�'Dxh�����:������޺Q-:iZw	V�u�9��?����?��Ş������Y#c�aQr$�*8|.<ݫ�d��:"��
���~}�n�����eY2c��r"V
da�0Kf�ΦE�I�SK^o�<���i�܀@�Ϻ�F�<!QY����r�mI�pA�^�<))O����O��D�O����O>ʧs�J9��6GW:�[hU�h�w�iP�T���'O��'��ON�.c�󮈼i.h9��cN�����9Y���o��M��x�O��D�Od�Ҭ�M{�'���Cq+Ѣzb4[WT;rN�ax�'��Z�����#�|�U�<���x�o�&a3b�%�d|;��D��ğ��	cy��`��08#'�O���O�9B6L�Ĥ��R�<��ȕ�>�	���D\Ȧ�cٴ�y�S��pQh��P"8X!s�M?L#��i�Gk�<�	2+�$�$Q�fUN����E�O��*��v\���G߆��Z�r�R ����?����?���h����T�]����R��\J���j�T�$Cצ���ԟT���Mۈ�w��i�?4��u�g	�t�JѠ�'q6-�������'�dn�<��L@Ƞ3&���4�'�P+g�����M�<$H��5-��䓤�4�����O����O�����Ud	Q�"N�*��/^�f�ʓ5��*ӄx�r�'�2�O��՟��"��8�8�e&(�-��ϗ������ٴ�yB����O0r"�]r����ƜclrL��(?���������Pd'���yEؓOʓln��m��HI�3DńV�L8i��?��?���|(Oam�[b�l�I�RBA�T��8-�	�F��]PT��I)�MC����.���8�M�i��)X8iHĉ֚j:�p���>QYh�H��it��O�T�1j��������&�5�e*pm�I����as��\��y��'���'���'Y���J�B�z�kEӹh�cJ?l�����O(�d����ũ5
ÿi�'fy
p.I�t�A��ۙF4x��0O4�ۛ�g�v���.p�n7�f�����YR h�$�:R,@$�bcW�gI %�%jH�KXB R�	jy�O��'�bF��an�����0Q����]62�'��	-�M���?)��?9���Ҳ#	�[���c�(t� ��R��<����������4]����'� 9b�I\X�����9$9�<�q*Q�%�6e�eI�@y�O1���	"AC�'���u��z�
��c��B�1��'b��'Z��'�3ʟ��O��;<�D��$.����G9 }x��Ό,�?9�7d�v���_}�|Ӗ|Z`�"1��1 @�<Ŕ�P6/�榉��w�Um�<Y��.�\ڶ��<�'�D1��l=���3C�N��'��	쟠�I�\�	ڟ �I�`�I�E7dc2*ț����g�c��j��I�	瀴�'r�n������޴�?��A�|Ќ��R��s��bC�9
B�i\�<���?��	�[L�o��<� ұ{gd^ ��e傻W�֨ �<O�(�e�?9$L-�D�<�'�?��k�)���I0���M"b)',B0�?I���'�?a���?����pC\���O\�D�0�Q��G�a1RU��i�~����(O���^�	G}��&6*I2u�҄&������y��'�,}c#�1AN����O���@��?�BO�O���
G,]s6\c� �%UJ܊�m�O$���O\�D�O��}���3:�eC@�OA#$�f��i�����	m�& �8 �"�'�B6M"�i�)�Ơ(2���Ht���{u'y���4F���@}�<P�La� ���dQw#6Qc�$��\ ��ξ/���(� g"�'�̔'��'���')��'��$�i�M�H��K$m Z1�^����4Q��m(O�d6�	�O�0@I� ��;�AN�K� %��F}��}�doڧ�M#���$�O���a�dd�EX��іa������$\� ��R��{�剁7vY���'��Ify2]�<i�NK/!/@a	�EB�kȐe�E��L��ܟ���ܟ<�w�y��y������`���[��P;g� 4"��05O>8m�A�I̟0��O�To���M�1�i�0��vJT;M	w�� �6]�!�D%�v6O��d�&X5�U���y����B����I�r�^�pW(1����8Ra<O����O����O����O�?��a
N/V���1L�����ϟ������ٴ���Χ�?q�i��'2t�P���-r`�Z�hW5e �E3O��W���r���Ѳn=�7�r���N&�K�,��<ѠL)tl���扶���P��vy�O�2�'��	W�o�TШ i0e+��puDE�B�'��I��Mkp��7�?i���?i*��ӓ㖐4��}��=1������O�,m�M��'��O�����/�ՉC�ӳ#�|�#����&��9��()p:���O����?y��=�DĔ#
 ��LH�-��՚�ձU�����O�$�Od��I�<���i�0���[�Fq ���j>6�����sR�'}�6-'�	���$Uߦ�XP@�&" [���-9�Ճ֋��Mk��1
���ٴ�y��'L��$���?�`�O.��֌Q!��
�ӎd�Ё��;O˓�?���?����?����I�JE�mc�	*�<�Fł<|��m��B�<��ǟh�	w��w雞w�����柭;K���7�ݷ%���a���O�7�i������'�?1���M��'$�)���ʵA�x��EKs��j�'"�l��@�$�|�X��SϟT��
�#L�<I�ə��1Y�)�şX�I��|�ICy�(p�R0��<O�d�OrI�V(I4{�Y���-Cy�0�AD7�ɭ���O&6�?�䖳}�P�TLû'[��*��ގ}���O���eB��(7�<���uP lھ!�2&�=0�Сbw�Ő+>ZP7�ۑ+x�'���'��ٟ��q�بG<@,��͓:��j!E��ܴOt��'\H6-7���m	&@Qq�9���2k���>OT`l��Ms��L��=[ٴ�yr�'L�IAsǜ��u�M�/z�����<�|1!�&Dfr�$� �'?2�'�B�'G2�'�0I ��1K�A 6fq�IIrU��r�4�5��?i�����<	dn@�'���J'_0r	(��T��<��I
�M#�i�ɧ�4�O����K`!Ч�3p�X�UFڳ%����V��J�i����3�y�XN>)-O^���eDRp�@˳,�J�r!m�O����O��$�O�I�<y"�iMh���'R��	�G�Q
̅��*�=+�9i�'�R6 �	����a޴�?I�E?e'vH����F\����ýf���ڴ�y��'��M�⋵�uWB�myB�O	J�4$�7
1��D�
^�Lu���;_�CP☫m���NR
W}rL�&�=	�	Z�G�B�Ր���1k
l���D���K�
B4�IC͊)Y=I����4��m����?B��<ҤAսX�x��ڀ�^�qd��Fk�>�<�w	^�	�p����Ŏf�N���.b���za�ЖY4\�h�"�x���[�� �xS�Θb >��am�)��]{��9{~5��a9�^��Oڸmd�9zrdP�v(n!�n�5��;���-S�Ud����ɡ�2Q����A�F?�}m�������2�����?����~Ҫ;D��2UꮖP��l�ԟ���ڟ<� � ��'�?I��?	bǆ"���P�'k\y��&�A�f�'��xj� �4����'���=$ab� OuX,Y�%O����'Μ�ɋy��'�"�'�剢K��1����
Iz!T�$|M�����ē�?���?Q*O �d�O6�AEG#mZ$��&֝v9H8�#�Y/t�1O���O(���<�@�(��Iռ`��̰��̆TlX�r�K7@��埤��V�ey��P��Ȱ���*��ɗ#Lj=
���P*������ӟ��'�ȥ���)�B/������2*�D�!�d�4�Jn�Οt%���')]������Bp]�wE �%!�!FE�1�M���?I/O�[u��a�ޟ��s�	r�1g�i�F�N�8�p��`Ӭʓ�?���9E����M�p	�?W�,��A]�C�%�a��%�'�<��Ea�4��O�O��x�6�wݱ�\��a�>I&j�o�fy§N��yB�?�|�'��RN�"`��Q��Lr6��ߴOV�-�2�i]��'r�O��O��Pm04�,�`xB�z��4^`o��u�����$#�9ON��� ]���x���3(��� ��
@|,�n���x�	�!q��?���|*���~�/B�PЀ�WR96Q��#UB������<� y��?i��?�*������7�ל	TԌ�u���
"���'�8h���*�4���?�D�@���j�I5�E�����L�` �'NH�y�'b�'��<؀ d�5�ۮ#��Y��Ń�#ňi�B�)0�'E��'P�'D�	-`�6a��% h�Cަ[}�0��>�I쟰��󟴖'�piCp>�pƫL�f�X(�Jʈw�J��0Ȩ>����?�N>�-O��SP�X�Ȟ�nJ����G�OZ.M��H�>)��?a����Ď�g���$>�'�Z���4g(2�ȶ���DЩoZ��l%���'�@q[��d��ms�[��^>$�<;�D"�M�����O~���ħ|�/O��酶l�a��¦}����l��{���>Q��-�,t�p
T\�S�$�֯R��1�KFbn�Z��+����OT�b��Op���O�D�8�Ӻ���3q���ir�ӷ����Eh}b�'���X�
�1����O r *G�.A��<qJ�'���4o�lp���?�-O���<�'�?yU.��Y>0�7���z�r{��
�5�&/G0;���y��i�O�d��@�
#Qع�We���UP�-Ʀa�I�����2+��������'��O�8qj��8k�{ebS�M�R� ��'l���?�	�Ol����4�'��"	lF���W(a�,��pf{�����2��?���?I�{B�A�	H�T;%�Z�X?<�tm��Gl��9��\�i�lxy��'I�U�c�� ζ�9PL�Rk� i�#V:��	ǟ���֟��?��L�J����Cڪ�����72B�l�7SF��'@2�'��	��{�O�p�b[�J�c�F�s�@�u��E��ҟL�	L��?�Re�QV�l��D������!n6*��5f߮�l��?������O`(���|��x��24B�o�	�r �Vܨ=; �i�����O
B� ���'����P�����e�:�P�4�?�/OR�$o�y/��˓��'
̺9�,q��'�	o�<}����/{��O��$��f�qI3�T?=0�L�k�����=R��i��J�>	��=�P�����?1���?������ބ��4i�L�*{Äx��S�(��:��%��+4�)�� k����D�1cj9RAUAxb6-� p�d�O����O�I�<ͧ�?A���n��Q�������kD�ߦ -���8=�.�	�y����O�aʢ�ڌ"�&u�$b�>��q{C�ܦ�������P0J�����'{B�O��� *�!p�H��R�ǅ^�>D��d�E�#����d�'t2�O�ՓM���v]2@-
�h��i�R/9KS�	��L�	��=iU�53
� �O�t�B��G,m}b���p�X��O"�D�Of��?11iϿvV9�'� �u$��$, �H��/O����O���=��X?Q�Ӳg��z1�_7��Is��Z⦍��+?a���?�*O��dϫm��!C�$%�@!�$<Bw�U6~c�6��O.���O��p�'�"���4U�9�T.?dv]p�
��Dd1�'�"�'��Iޟ �G��n���'z�K��6��i��J�>!�jǍv�|��1��oy"�_���h���Ѕ�7Z�U��&
��n�蟠�'��ۣ_�������I�?͋�L��0V8hL=e$ pDO֎��'�-$�<��y����W@�T�����
�tR��	�Ll,L�Iݟ����P��PyZw�<Q�_+*�K�>����OX��X8[��3��Ic"���F�n����* ���8Y"�'���'���T��՟��^d� ��1d̷J�,蛆*���M���ߤl�xq�<E�T�'��b%B�! g��u��5O���[��z�4���O^���U
���|2���?��'�N��䩄�smB�c`�N�;��(�! +�I���3N|����?i�'�xC�"јfs0�(��ġ54.�ˬO搘��<����?�����'x ��
�<^���TF� Hz,!�O�PS�/�%����4��hy��'�t4��ŵNd�=�GC�;o@)��U�A��Iϟ�I��t�?��6��zeH�5z��*�ʋ����
�]5(y��'?R�'j�	ɟ�� f@*U�E<_xu����Z�rTr�������	���IJ��?᢮�<<�(nu���S�F�-VD� F��w���?�����O�d��|��p�܌*�D&�vP���!~���Rv�i�����O0Q�'.�!{�'�<�k#�JU�p�c$�e�����4�?/O���W�z��˧�����5�P�!E`�XYBiO@FP%s���n��?�$B�y�|�<�O�"$(���5� ���X����O*�DƊ����O ���O����<��C���jT��2t|����+C���'�2�� 	?z��y���%?j�b�I��ՙ�XQ���0�M[�J�?	���?Y����)O�I�O�Q���5�>-{r	��|��0�F�������b�"|*�iH������!��%�2aْT�5/�M���?���})d1�*O�I�O4�D��$�H	 7 �@�A]�2\I�f�ޘ'�}�Q�%��O~�d���y�	�{��@��_-�b��v��>��������O8���O\➠Q�B7G�<, 4Ɓ$�����>�&�Z9N�R��'b��'���럸�� Ɨ&���r�O��vl�򔀌�db8�'��'��D�O���CL�p�8�a�����2��~�je���|�	��'Z�R1���b�(�PE�	1Z��d�!'%c8���'�R�''�O���ن�r˰�i��yD(��r_򤲃���^/ȍۨO��d�O˓�?1����I�O�<� �(���̈́�n�iWG�^��:�iP��$�O�<+�B��:?�'���z��/%��I�DҀ^69�ߴ�?y/O�$�zT˧�?!�������I����/D�V����1�U�8��Oz����XȌ�ҵ�T?��Ώo�d����(ag �{$�>���f������?9��?���������&�R�t �	&Lj���V�����<An�-7�1O�����S�ל
Ĕ��F��*��"�i�����'���']b�O�i>}�ɕ:���AC�  ��q���2,�$AjڴPi�Ȣ��K�S�O�bM�甼��N��![d�	)(7m�O��D�O����<�'�?9��~��%7.8U�s�Y�ɮ(�fL<Trc����Ĵ�ħ�?Q���~�Ɨ����U+X=lvP�E�)�M��Qj#/O^�d�O���>�ɓ2�Q�jU�C���DL����?�ʴ����Y~r�'HR^����dJq�&i��r!&��C�4k�0؂C�Tsy��'�r�'��O���"�1�d�@�#ҜUQ1�ݚM��aV�Ϭ5��I��D��˟�'�摙�m>����\�!X����֍^�ޥ��m�N˓�?	/OL�$�O@���"��KTi��Ȅ$M@���W�l�Qm�|��ܟ��	}y��	&���'�?�1 ��"U�M!76��S ڶZ�xioǟ��'���'�fU�y��'�"nI����bʏ��rdj�6H)��'�BQ��Q������ON���Ձ�cM7ur���X<@D�̺���z}��'�B�'�B]`�'�b�'�� ��՟L�;�'�5 �q���FR4���i&�	%9�@*ڴ�?q��?a�'4F�i�ͫF�_N�N�X,J��G�wӊ���O�uln�\����=��&H댜  n�^qԑ�HĻx66Mɛ$��lȟ��ş��S�����<�f�O�EP�EK�I&H̬���V(�F��:�y2�'�	b���?9eK
~\k��7f�ҔY��	k�v�'%��'s ���b�>i)O$�������9a&`�U�R�Y� ���~�d��O4���� ��?q�֟���w0� a�yƺɰtiߌ8���޴�?a�7e���Cy��'���ß�X�$A���ϫW������˜f�n� H���?���?���?�-O�U�AŊ�0d
��]���r��&*U\��'p�	����'q��'��i�LY�0c�R�C�`xC��7w�h��<,O2���O��d�<�A!ֻ��@�2�����@��	}���B^,���V����{y��'82�'�,`�'j��G��6Lz�e�+0\�X:�g�>i��?���򄉌~�`��OrR5 �`5�C���K��r���8WtV7�.�vR���Iݟ<���c&��Io��4j"�,���	�x� �ُXAnZt��Py��
�ꧤ?q���� ˑ��|�6O <u��Hbb@��	����	ҟ�{T-�'���i6��.	 6ib ÷�^	m�vP�4�%��M����?����^��
��C�9vlD8Æ�=-�6��O@�$�+�DEU��'oq�h��hv��0�o 8x�/��#U�N67��O0�d�O���f}Q���b[ *��R%��r��T�a΂;�M3�[�<Y��?�0k	��O��������Тޚd��ە@�%[S�6m�OJ���O���wkUU}�R�@�	n?!�eѻo��5ۗ"
;ef 䭈Ӧ5��yB�X�yʟ����O��D�;�R@	�&B�0]k�U��Ɣmʟ� �g���<	����$�Ok�V���3�K��f�� ���I��MD�M��Ș'��'�d�'*RQ�����I�z!�P/�m�~�j�.?O�����O�ʓ�?�)O��$�O8�$��4Ouy�E=G�����ܠRcrMr5OP�d�O��$�O��$�<�j��(��I
>%? M���7N� @D)�'��&T�<��fy2���Ms��z�^dϓ"?,��+��>*�tc�΅>|�ڗ�i@r�'t��'��IY��s����$ȮD�"�{�b���٨�J�x�o��`�'���'�ro�;�y2X>9H��[�
U���e#|���)�������'K\P3��6���O��銭b��M(G��@�B���/�#�x�'���	��tCUI��'���'l����P�ۻ@4�R���W2$xopyr'�g_f7��w���'��t
6?1K/?$���r����$���	ß�+mP��&�<�O��$с/�~����8ň��ԯ+�&���|.�6��OD�d�Ot��W�՟l!��M��0Pa,U�"X1㦌V�M#�F��?�I>a��D�'SD�@'Ǚ 1U褙�L	2V�
}�#j�T���O���H/gאI%�(��ɟd�<�t�k��̋r�����X�KЀmN�R�J|����?Y���4H�E�'��$�1a�)�x�p��i�rL� b����w�i�9P�W�M�A��F�l��%�$A�>ɢ��2�?,Oh��O��d�<�bhI�&fA�G	H�ո [���jl4��Ցx��'�B�|��'��`��mE���-�8x��HW�ڢ��G�'���㟔��ܟd�'1�4�!Cj>��v��hK^�B&�
	w<�)d'�d�O���?Q��ybf��?��ȉ��e��g��uMTh��/	���Ɵl������'�@��4�)�iǡ(�ba�s$���lpkp��Ev9l���&���I��`ڦ��͟��O�rq��*5�`��L��X2���w�i"�'��	mBj�J|����q�̽	�� �k�'Yݸ1(���'��'����'��'�i�I��؀�B���Dҷ��'"�&Y�8���M;�^?����?��O� �i�s�ԶZ�I3��L�v��]��iuB�'����'A�'�q��P:�L����`�kE8y��!�i�(8zrOxӒ�$�Op�$�'���	�d�M"��H�naj�;�ⅵ4Nt���4$@�����S�OvR��An.�"��ɀQ��p�@��]m�6�O����OpUᤫRR�	��d�	a?��	)dE��@��ˡ"M̠�U#Ϧ%%�pIw��>��'�?��?aBJړ~Wd��f$��p��㔸v?���'H��٢m3�4��<Y��#E�F��P�ҞK\���Tʦ��I�J��	џ��	��(�����'f�D���rp�ʒ�W)a|���#M�7I�O��d2��?A��Z�\lU��W�6���{�n�0.�������D�O���Oh˓o��5:��|`���#�x�X����\QS[���R�'KBiþVb�K#<��!SKh��Z5g. n��?a���?	)OJt���\�h:��I�CE�n!Q㥝���0��4�hOb��I��0�� }�-��P ����c�&��K!�֫�M+��?����?�5��?���������:)ҵ57��"F�^/Md����Cv����l�		�t�AA	9�~���E�Ḁ ѭ�Db� ��O�'	ֹ�ly���D�O��$� ק5�n�
Ty�r�[#��i�H
�ē1�X0!����ēT�D��4`�8P��wiP2�nڎ� ��۟��'K���'n�[���Q`�
6���恧r���m�Mӈ�'�&��<E���'6�̐s�+�@�Z�=�v���qӬ���O��dԉT^���I�O~��#s�d��WN�!���*L��Ɉyb�ÐU� �0�d�Ol�䓌+�h1G"�.T,L���$� *R�mП���;���X���'���>yP�3��=%��6R#P��BDW}RƔ�_�'���'��'��
O)y�@��(D���.l�z����'��'O��'{�'N��'�XC+X���ѫ��%z@�	1'��>3K|�B�O��D�O ��O�ʴ���D��E^��3������5B�2'Ѣ\l��p�I�(%�t�	�<�e�+t�t7-��T��Aj���7�&Xs�ʘ�(v�Iԟ��I�@�'݄��n�~:��R��t��*gԒ�X��n�;&�i6��'
�O^��&G �	�V�[3�ڢ?��\�sk�Sg�6m�O����Ol�ď�%)�˧�?���
�*O(ٺ-J�I��OXF9����W�'��'SH�c�ʄ�����SͲ�O��uP�Cq�
�]�65K>��m`��yB���H��Py�f9�	�	)�'Z��QC�7?L|0���@^���!�:�8c�eJ����a�?S
0�`��>,kޤp@�
�T,.HSd"�鬌�p �,k!f|�Sd�:IH�kWIĥ7s
|����"0Q��sQ��|���%�:Gy6���f�0a8��Jë+�nФ�۴Y.6II#��$����p	F�j�� ����'��'B�c݁��矠��*M0=D���	B$|��@ ��\�:�*R�A�j�`��t�G%@�����(O�<�ጇ��4��CY]�l2�e��̐p��&]w��S獡#^��cg���Pj
����1�q��9v�0�w%@? 5j��Ho�T�	��E{"W�$�Ca�S�@�J��Ls6�Î;D�����t�*X�! �!i��Ѣ�k[��HO��sy����t��7m�eN�� ��u��D⠮̿r�����OH���O���@J�O��x>�㉂;�x���̏��0�/U�%�5h�8�T �f����.R���憗@���8Q荸r ^k5N;cp(�yT�������;cWr�'�f@Y�+����)��3�.p���o�'��� 2�PFO�t#�.ò'8 ��'nxc@H/JޞWٿWЌ�`u�l���O��W<D��S����A��F�2f�#a�3���!�]%-� #��'���'x�sA*�)"t�4c3��4�T>eDh_�1~6|Q2-�4kHhR��)��t�a�n��^��X����'z�6l�4�1ntR,@@b��~��tEy�)H�?i���O��l���Q8Gb�@���]�U��'���	
T�����X|����0>�3�x� D&K�8�w#���Q�c�R7�y�,�A?6��Or���|��/���?����?aq�UV����u�@��əB��۞�Y捝+f��3܆�*�hc>��R"�~-h�+@�f�N@��F��q�*K���6��pk6MH<H4��޹5�~�q���w:� '��=�8R�+6�.���O2pL"�aӮ,oZ���D����d��E�`��[5��S���ϓ�?A��٣��� G8Le� �י(8�Fx�*<ғ��)*9�X�A�Ϟ`U��3j���D�Od(Ƞ�W:*�8���O��D�O�d���?q��F` sƄʛ!��eaǙ��;L	�ɀq��D�D�X|!�*�d�=u��P����r�NZ�������f�B6�Q=1�V��S%�mO�D�Y���'������՜cp0öE���	�'�.��qfU�VE˅��YQ-�S��yb���(c3�Q����c�Æ�ybOS�����@O�B��ؒ�#�y
� ����B�,S?�ɸ�g�"$IdĹb"OZX$��d�A�riL�#Hf��"O\%�tj�,d~���gڛI3� �"O�	��@V�����تR�l!��"Oj�;2� 'v��D�jΜv�aB"O�Q(0lv�)ʕ�H K�%�$"O��a� <�H�(T�]P��*B"O��2E
�:�f�{"|$�$"OH0(%��j�؈؁jsL��"O�7mA�@���x����
o�e:�"O��H�Ɋ2@б���K�YUv��Q"O��al^�e�`}�Q�N�O>��2�"O�([s���|�|AI��֖�:�bs"O��(��L�צ���n
�z�<��w"O��D�1�����l���q"O�T�kȞ�� '�J�B�A�"O��@��qހ�cRIF%�\� "O�xR$昐�$\#Qh˭��q)�"O�`�a�.)P�I�@��m~8��D"Oh(	r��g�i�d�>_m�u�"O��G�nz~�qӥƑSWJXh�"OR9�Ue�.��X7�Z&bL���"O.��#n��?����n^�Kq&ͩ�"Or�hrʕ;��r5-�nd2p{C"O�5Ad"`PT@2%��	J
��C"O�l�� �Z��HfA�R���
�"O(�k�_�s�@s���F�L�"OT���XwU��f�K"6�����"OZ�Iv�,��)�덻DLr��`"O�Ei��[KU��h�JQ<l��Y"O e(3��#y}��P�o�6m��"OⰢ'��!7Yh�)h�n�i[$"O����
� NucAQ19�,��#"On�`ˁ�z����wL�aR��V�ov�I�a�O��`$�"����0�	@���8�Z��@S3Wc2��P��q��P�@\{��ك+v8�R���9|w�q� ܅'�<����B��1=�©#�,Zt���	" \��F�$��С�$����,8� (	W�@�H9�Ad/D���&�U�bd��L�eej�ʆ�-?�	�k��)���������5!$�����V�x��{jZ\!�_�1�t�@�g�Q����e^�31hdEF�>D���;{�vx��i�"�Hp.�HkXahAG"����*��|� !��M�"d��R!l��8��	�ϠX���U�TC
�z�C�!| �� ��?�\�ɱ��ӀF��<������ t�aȁ�O�.G<L)1�U��0<��[>�RUz�mR�Al�,P���F1�4eL�5(��So..Hl�*B����֢'Xw��!�O?7T���� �	�)�]��B��M��	#6������<C[~�)��Yf�O�b�T��'n�A�$D�|~�P�'�,�0'%��ųs�#OR<*�+׊o�Tѡ#�I�5�Eɶ,ݓ�� E�O%ZՇH�1��6��L�8���x�\��Q��Q��K�G�>�:���4�O��`��+Xj�$;�+�>�!1$�78����P�y2��揽���A�Q�<��4{��O��=�E"�X�0"����p,K	�r� �Y�M�D�ȼS�oA��?��B� B͌�j�������/(� �Ę�v]�A��4f���C#G*%Đ��5���-.H�4� ��gR51�ܑ��`�:�?I��:=�U��	�: � �u�Jȡ���eŊiyb�K�<�$�K��(;¤ͤN�}bF�-�p,�b矒�?�`�ه�`�� �2���ēO�,�j�w��QC��$`��I��]�0x�0��'�~A���O�T�84�(�0�s��� ��H�NE�s2C�����$/j�O�4h�tɰ-�E��0-F�D���'5h2.�?�� @K&�����O�2q6}[b�I9y4T cv��P��)�'ހɳDl�(e|v�cS�	!"����$�0� �c�ȔJ��îR3���O�蔱6���Q��l1S�ă$�a`�'`�ZB�q������ƯI���r��etP���,<Hj��	�?�~���w����T(NX�@�&�H���	�'�p$Q�j�jE�UQ�����W2�~���:]��9����|J1N����� t�y��#�n�P3�KU"p\y��'ߒ����#5:� �A��݀�o�i
���а)pf�-{�����'sl\�PӬJ�y�L;J����ċ?�ٺ����0�L�6��O�N ��A�}o0�AԢ֐?a"��'z:`A�֔!�v�x�	��3!�p ��P�nL�`��g�H:�'r�����i��)Քc�T�uN��Q��"O���&fؓ3��BXP�S$JS�\����"nȳs��r�D��O���W�!~�J�yR	]��SF"Oڌ�c�iwĒ!�E�����ݘyVj�r�PY�����F�s�h�BG$�� �D�+�Cl�az�_ 	�Д�)�+��_/ 1Kڶ����D�e�<����m&x����'��U�W�{�$��������96R�|`��I\!�ν1Q�6{v ���'���Py���Nt���s�֭2�D�z&�]1-Xj��@_��q㉈7E�c>c�\�RF3(Ӟ!s gJ(g�0Т,�\�VN�mJ2�� ��=�4Pr�N��%�0ڢ,��Rن�	�$� `v�K�Ddtr3�&\����$�[ܺ$ Ǩ��y�6�"�`��@\2�(�m���T��'��D���ӵ-�-��n��"��qI�!J��Z�'�2�@S�Z������ӎ0�\�!� 7���PGI�lc����GHQx�p�ޣq�v���AO�E�4pPg���<c�OR,x3���zc1��	�U0�!	Q̘�}�@4���>	��Q��P�� U����=�剏0�� Տ[�Q(:�t@͓!ߞ�
���Ȓk�l��"�
��R��r��H!1S�sJ0O�����/�
��6o���>��並k�5-<L�cr�̩5r�ɆoRh��?E��cY�x�dljw�ҵ+spE`��ߎ����+����D���Y1j����N�O�t��E�^� ��pbb,.���H�'��<���_�u��{�ϑ
n�(PJD��1m2�$��Gh��8P�'1�1O�5�0�@2�l9"-G� A���O�4�4�0;Dh�V�$��
-�m���P)�A�#^� ���I��2y���_A*m�bE���ě�}r)��i�
è�f�DĦ�X�E��x�Jï�"�E `�/D�y$���tV����	�O��ɗ"-?�#��3V�[/D'�TQ��<���P���)@dY$,�RC�	_�r\!�/�=	I����
N&���)�����45���B���f�g��L����+&�1s(V�/�����GQL�KU/=�X���
��9Bf�՜}2�#`�T5���1��'Q���դ+[�q��TB7�x:
Óf�X�04홙r��0���ғ,U��mߎ-	l܃�ˀ�A�x�{B�?�ybǘ�)d�*��
3nDR�L���D�!U�̩r >t��8�q!�n�O��̳'bE�� *�eے6���'G�L)�jɭajrHB��b�rMX��ɖV���Z&&f��G�H�Mc1�1O�4Jd�\&"P���<|=b��O�5H`d� ��y��MΑ;-d�x��V<�(��(����<�SB�I؞Hpphǵ;<2���g]�Q�$��`�-,OxeJa�θ��ix!���V�V(XW�ݣ/�j��)��O�&�y"��<�l�6�U#8�Ȩ�$�߁8�(���Ot������M|�q�A޼�Β�;!�9X��֕j
���ΕY�<Yak����:�E''f�9��M~�&�>y'����m!�I�i��O*�3�]��Y�DcϽV)�����'�<x�1�_�����(x4��D�[Ȥ��7���!��\A��#�(et4�ĠY�I1Od�D�X�	Aa�t�\�5	��(�&��%�:I��OY��y����X�IR$ �ƾ��7"A.&qJ�k�y�"@,���	�ZGf��Amԛ{�N���#�3�2B�	����G�	��6�g��}�@Qj�m��|���DL�2�P����Y2z%k��;�azb, ����Op�١%�(�I��@	�#�x��"O�Hz�l��@�	Z��X��T0���Y��DKe�Oe$��r P)l;V��FPm����'�u ���Q1���F@�j�8��'��{�ۑJ;[�C��fӐ�(�'9���!���$���+`���J�'���3�����Z�q��+������ ��R��5�~�@��.4�2�h�-1fP�':x0j�b0�3�D?f8q�5@T�R5b :�C�`t!�X'���M�,=�$�����P�0m1�
�		��c�'��sc�r���O��>�V��
�!�>�kr!��u���'<|]q$�
!D�ƨ � �8�A�'�����$0 ���I��
@�J<q��$�5�t�[@�OhP�A�A̖ʂ��$ݾ]̮��ȓ<���aP� u�	�!�p�@���	G��r��L<��U==��0��N21�dP���rH<9�o 8�zE� f���a��O�x�F�@ CP�S<� ��Ie����/����49��y#T��ɽ2>�R䉔c�V�UX�M"H�"L������1M!��ȓX�֨	�[b
��e�qO�m%��Y��W%,�,��K<�'�D�ȡ�4O@p���T��<�ȓ/2P��M˞**|9�qh�f:J����U��ɤ%�d�j��L<�!B�~� �1Y�f���W�MYH<QNЦ~Ӕ8�pX 
����}dM��M��E�ࠄ�	�]�H�si@�l���c�"�����ӂR�^ei���M��"d체��F��l���TV�B�ɓ]&&��Q��6%[H���oՖ@�O��sGި)�:<92�o�&���	�>�2TZЋ�{�B䉘 ��&-D5FU���7ڪB�B�	s��P�''�S��ݙd��8>h�C��1�HA�/ˈM�6)�c��=y�rC�ɟ]���0�"
�ۆ��MC��p�D��IR,��S�|��C�I�l�J	���1��n�5��C�	�5"��T�R�=�e��-�ɢB�I�$m����Õ/��Iʄi�;Gm$C��:;~�q%�%H��X�Ԩ�N9�B�ɂj$\a܍r�pDAT�M��B�ɒ;�\��G�(���J��P	��B䉱V��HPO//EH����W`C�ɘ1 rH�cBA�e���5j�TC��{8��1�H��t����e� ,�$C䉺}�F �a��2J���m�C�ɔyP4M�B
F2�T�Qw��.��C䉲k�С��$��b� �5i!GdC�I�5Xi�d�&b�;$�ƶG].C�	0)�,P�v��$@� �uA#r\�B�ɞ[�����JW�J��TʔOG!xP�B��<*Y\��eOM�$c`$��O/5m�B�I4���l	,$�0���m�.5��B��0x=&lMz"�Ԉ�L�39�~B�	�X.�QIu,G�Y�̼q�
ܡT�TB�ɂ=G�e����+Ϧ�����JB��5Ohec� F
 a.)�b�d�8B��!9�`���FB%d�M�R�
�)}tC�	���Y��!@�RABG�*�@C�	*H����'O�l�	3��*��B�I9p_��B2	Z�+]2�!�Q��B�	�P-T�Z�ؿJ+�����)��B�	�`�Y�W��Z��p�Un1�B�	�v����Q���ԫD�޻d��B�I�H����b��&&u����/^7N�hB�	�-��pk�U?G8f����� X�C�I�@�8��A�`D��ר�",fC䉳ZG��	P��%�my��+||C�	�^D��eJ�5T��B򬏩X�RC�I�1�r� �!H�Y|�ٺJV?|B�	ު��gU�dv��G�6q*e�	�'��CW��5�f�h��O�YDx��'7��aə��$�`J	�php�'t����ʝ*g�m�s�ߤu�l���� ��9��˳E',����ߞ��K�"O�EQC�=���BF68��4� "O`��NDu�	�� ,q�JE"Ob����+�0��Wh���k�"O4�J�!W4iN,ɒ��[:�Tp�7"O�A2�o�/tP�hM�;дJc"O��B-����b�U�2뮄s6"Ox��cȞ�FiY��IG0���"O	�1�ݓ o�%rE��Y_���"OH�HQD[)A.��Tn� Bf���"OvM�P��.�䌸�*8(\p�"O��
A�ɥk��1��K)�xx�"O\�&J��|�(�W iR��"O�LP��

^�R�z$�(�Ҳ"O�-�'K&q���h��R0��Y�"OH �KNH&d=0�9Бx"OB35�Ϡf�0�;�d��L�Q#T"O�	�Fa���t�K�c�',C�`�E"Ov���&P-6ت�(Ѓ��K!�mڧ"O������2��'��̨R�"O���0�ʧl��\�ċ���\	�"O�(סL�5~T1�Ð�e�@���"O��h��Շn�l��� ��vhVp��"O����\Q^d��ު:��MI�"ObE@�OFU�ldj��� Uz"Onuitoٓf*f���cW�@��#"O�\�w���H��#�"?6��S"O�H�e�
�#��0W�  ��'"O�A�Dk��E���$/V" ����v"Od5q���E�~Ȣ%�6I ��w"O��SE�׺[u*t[�`I')Dt��"O���ˁ�g�� �� ��R�"O��헌?���RD+ۻ�I�'"OL�C� I-I����L@qo�Z"O8 ��\����c]�``�!1""O�i�@�G�g�̐��X�A�BD�p"OlmBІ�8*���c�8@�X���"Of��"�oު��" S'j��Q� "O��B6d��p���Ha�Q�g�"O��B����HhkD�ܹ1[��"O0�W,C�2K4ta!	ϴ-[jm��"OĽR��'C�V��TH��II��`P"Op4Ӳ�Ο{�.��'צ3� ia�"O|���ЬH����(� ����"OZD-97�p�� �53�E��\7�y�OD(\O��Q͸;�J)��*T4�y��}0p{2�N�F2H@�6"�y2#Z�FgR�2�Mݙ5,�E(�?�y�C2;`ht�*�&2�]�H��yB�׻M$a�r�.-k���^��y�Aj0��`%�0�z��ա_�y�-?g�!a6��,Rw��*�O	�y�f'2�Թb�D9[�]���>�yĀ={�x1$ْs�P
Co�;�y�D	 B�JBF�&��Yz�"ԅ�y�R������&�p�#�MѶ�y�h��q���Q��6t5�@31펍�yR
�#e$2�	C��2��t� ����'fDP8p�^�&�Z��F�M�PU��'�����Vw e��"�'C����'%6,���׆#}�aa���G��H���d-Ob�˕�O�?
a:��*]x�[�"Oa����{jʌ�uWDf�Yu"O$��V	����B 
�N$&,�"O� V��5��e�~9��!	>ht��"O����#!Hx1��Ɓ����"O��Q�b
�m���ȣL�F�8$;�"O2����!h
4��Fc��� ���:LO4��ӫ]kD��AK�b<�{e"O`Q��ȉ�h�~I �g��$UX5"O�H��/hF0�9�g��T5�E"O�� ��E�R�P� ��;F)ؽq"O�lA�e�&�����!&j�#"O���%�:Y����đ�59����"O(3�Z(P0u����}�a*�"O
P�VhϢr�fu�&�:*��#5"Oe���:Wh؁j��dY�"O\��6�Хt�N��������q0U"OX�	Tcɔ&������F�N�Bt��"O"��wh�>�=����t����2"OS�J]thC �a�tLYV"O,��A���6$�8Q7i�-�ؙ��"O���Јuђ�в��nV���"O����M\ʌ�c�� � tـ"OfT�Wf!LRZx9�.�yv�1"O��0�`�	a$	Gh�n�~E�c"O�cӋ�!�"@�cEO�y���A!"O"�b��!U	̈�q��.CDRR"O�q+������D���V���"OI�SBOq�
8���"�ލ��"O�T���B� =��@�_�d��g"O�%c�/ 4P�(��%Y�
�N�;P"OVL[�jZ�3�p¥��/|��9�"OD8��?z�e:��"$��=I4"O ���f"dR��t@R �¸S6"O�ë*m����M�b"Ot����	�&����_�t�V"O�h�_20se���^��#�8ШO�#J�+IxJR�-e���w��|�4C�I=v؞AiQ���%G*����#5drC�	�J��!yal\�bL�1�C��<��d/?a���Q�tᰠͭV��0��NNf�<��e��;�XMÆ�F�4��YR���K�<��f�L������L	0�����LG�<y��˳Ay��#$
1uT����^�<�Ɩ0��%ѩ }�D���^S�<a� .T���r��"�,�#��RO�<��"L��f�2���+'���s�K	H�<��J� ��W�����`��Y�?.!�BCvHq�ceĖ��uSm�!�$�.#^�!E �dZ �)C�ѻ�!�${��IXc{LAp�]� +jɇ�	]�%�ɛ
7����@�L���ȓ";&����e\L��T����n˨����>4P%�F�J�CG�B䉓6�"BoЍ.D�%�H�B�I�^H�+����4�!RzLC䉨{�~�`���3���Pa�@�?7�C�	�ٛPE%>�1�����-'"B䉝%�t����M�h�ژ��C��R�C��)i@f�8�&JA��m��@ �C�	{�����-��T $I@=lB�I�����5i������'��B�	*��@�1]]�к4��%w6B�	�k����e
 =^��7-Lu� B䉀�*!�U�n�ӣ�/E�C�I����5F�*[f!�	�PC�	�|^:�p�̉#6n��&�3J�nB�)� �4�C�V/J@�esԎݹ(q��X�"O�]��g����D-���.}�"O����X�@����M,{�h@�u"Ox�����<�xU�
)Ì]�"O���c�ɢ&,N�w'RP�Ԙ�E"O^��Dɢ(��X�Faq�^�ʅ�IL�O�s���)�]�P-�I�T��'���Օw�`"E+L�ZT`�'���5K.P\�SR�@�=H�X�'�������Z��0BN���~a+�'�<�+�@Z�z��t!ӈ ��5��'�L䈇�Q�8��y�JA�ͼI�'��2g�C�l��tS�N�:P��!�'�p�ԃK�&h.�R�KM�&`��'4�Q�Ĥ�8Ƹ`��_�x	t���''�܈�hJ*۾����-x�.��	�'��,	G-��&NB 6	R�i�be�	�'�v!�rM��L#q��
F&IO�|�ȓ�����g�EbU����}�2$��Hh�Q��M!�ƨ��A !�C�	�S�����ѐ9}�iZ��ۻ*��C�$=p$�¢�Sk�I���1Td�C�I2T��8V��Vsv]�Gk��Xa�C��?u<��Q��V�$ء)�) �`C�	6)c�� ��8
�D�p �:zrB�ɱh;�Ђ���=k���G��fx\B�I:LR��:���2L������?|C��6KV��h���W��h�@i��^�HC��$B)�Lѱ�
�~
�P�*�7R�|C䉅v6�q�+\3�x9T@��+f�B�	)LxY��ǞP��4����<q�vB�	(2���(�R�l0��Iӓ8,HB�I:nȡ��"�;�R��� +RC��/E="p�j�J�� �ː9p�B�I(Dc8y
C�~A,�s�aUNB�ɑW�F�����lo�ej�i��97�B�If�� �v��+&���j��̚yN<B�I#U�~!�+�FX��ѕΜ��(B�I�$8�4�c�(xJ����WQ�*C�IoJ����n.>�j�+W�1�C�I�>fԁ�)'e�6L��'A�r-�C�	�I�ƙY�	�*[1b��Eqp�C�ɛ�"��^	��6GY�g����'�Ԭ��l8B�#�A
.6��E��'�.�[� S�X㤄��5�m�ʓpY�U�c��W=�m�3L�j�%�ȓo ��3!P3
HZS�v�,�ȓV.��@�,<Hʅ����%.F���e$�
����7�8��X�D���ȓ�<8jDJ�8rZ.�`�+کXCJ؇ȓ��i��"'D�C͏�9�T�ȓ�z}Bs�>[6`���4v����`� �Œ'PN�a��8v�P��J�z�	\��
��$"��e�~9��j���fhO���Q1�č-D�D�ȓ]/�3Eϋ�7���q���0i�ɇ��p$�0l�1Z�=E�Շ�'/���C���O� �9wY�8�Lx��<l-4 ��m�Xi9!L�j�x�ȓ/֚���D�5x��A�i �MD��ȓ��ș��+�v@!�CL�v�bl��|2��C�G�e1]R�	X����ȓyB5cG�]%{ ��FK�=>��,����!�R�\�M�ܡf�Ҟ��d��S�? ƅ�RG�%KƵ� �oor@��"OD�)��5��{�J K�<A�"Ob��С5�v�x�){�DiP"ON��%�٧+�쵁�b�2R�Rh��"Op��@e��0�t����[�$�b)�%"Ob�+%�O�Q��l�r�8@cvTx'"O�\1)۽\%�����6CaZ'"O0!��@3~Z���o��W4
Б�'�z%���MY�z�h�%ȅ�V�Y	�'�>�B�W�o��7��KP�0	�'�:�;3e�6�01!�ET*K�,�+	�'���J,&�0$��!y�1��'�����=r��\x�[����z�'�x��q 	68h�(�����Y�'�*(��K�/����@�A�~��
�'xYX2�:1��k���D���{
�'��+�ۦ%���PW"�%� h	�'�
mз��
/$��ړ�H$h�h��'��=I�D��`���4#<���'��Q���;Dў�jQ��$��	�'Nz������9𐭏�G��A�'�,�
�m��P�p�T�BZ`B�'4�����<7E�)"��o1�u��'n�����:7���V�͕6����'�lA�h�,u,$�UJ�)`bR�Q�'n��Q*O<0iZ�Z��NEL}#�'����@&Y��9�#�pr�D��'�( �Gm,�����-S�'�ƅ�$-��R} ��T��ڸ��'X�a`�S bXAuo�>�
���'��UC7�M�;�p���y"�k�'AƱs��ٚ5��([4�o�Q �'j�����1RV&��c�\4a��m��'"Qȱ�	�{��YV�M�PJ�%��'��H�bT4`�;v�٧@r�$(�'�dh���Z5����$Q��'µ���.]>�yE�"+�Y��'L��j*�VƙA�5VYp�'K� ��S@,@�%� �����'��x�:Qz�w�CψU
�'b܉a�)Y��yIP-8�
�'.���U��^0@i�V|UF0��'�= �Lپk�����$!+P��'o�ew��<4��@VjV��!��'e('���)��졥��2$��b�'}�y���"�r]¤�OAXţ�'O��;�(\3rgt�ʦ�ʂljYY�'8>��ƥYa��r�
�XƵ`�'v�+UlO�����̋�"���'�L�a�4Fx�� �#wGz�2�'�����3mM&H�"�&h�����'�z`2L� �갨GeӠm���X�'8�(8!$_�!���[�(mn`Y
�'�  �����	w��8exrؘ�'�����Ő�.��3�ȕ��j0�
�'�0�3f^�YV]����%�ș��'��hy�(��& �srd�/���'l�O�D�JMj2���W���'�(0��C�s�t�F�7JO*I��'��p��ʢ|
��yפZ8E�P1��'�8�KBY̸�	�*;��yB��9��h���4'y�\��	§�y"h� RB2D��NL�O�3�e�y�؊R*ܪW��;�*T�CdB�y
� �T�W���|9c'�" QhkS"OdM� "��L��&F�Z�pKs"O8�f�İTa hh�gB.Y���a"ODe����\)��������JL!�"Od�����{^��Kaŉ�0��MQ�"Or4�%ҨS)�l���>�tyR�"OZ��6 �*Vf|Y&T�f���7"OV��7���>���bX"�Ԡ�5"O����!G�v� ���O,]�Z�j"Ou;�o�/}��x%���e�f��"O�dKb�fw,��L�,�䷆"O���@"F��q�I�n��I�"Oz����M�;�ڈJ�ϓMi���"O���pNH�a=�sLG�(c=�d"O�����Νg�r$�̾`l��{s"OJ���R5C*�)�/��5j�Q0�"O~���Lq�NT�� �$}��ȗ"O6���C�1`��y�T �I��a�"Of�ňΡP��]���A�
*���"O�x1���* �>հv��U�Z<]!��?0��\+A�Σg6��kʾ2K!�D���6	b�R�&<�{U-�^[!�pƱ"�����Kt�G/rJ!�$+#t��a@�;Z��A6C�!�䂸%�zT�a�Y�z����_�=�!�ٰJF��K� ߖ��F���!�)L�@��� Wݴ$90�K�!�$	Μ�@El!s]�qcq&��N�!�d�1T-]*�.L�
R��"V��;T�!�t�f�j�H��7��Xg��^�!��J�
@L�x�L]�s��$�y�!�DH����.J�e�*���ȁ'i�!��/2D�HGH	6��E��I�?k!��j�t�Г�߫eގ0ۦ%ء%M!�$�	� I3T�,�L1g�^�wK!�dG2����uf�%�f� ���m1!���$e�v	9�@�5WԵ�P�͆I�!�,z/@Ȱ��k^.(��'��n�!�$)fl^4�u��"CUB� Fŧvm!�DR�2�Y �O�I;,�	1��ea!�<�bi�+  {��.�����/D�`b��L0C�)��`јG�$I6*O��9�%�N��sb'�c�ȁ"O`)x�k�9:��ʢ&@18� �"O�|Zè��S ~�c] D%�5V"O�����Z7\�vtc��B�j��"OV�;��R�W�!j6B	+v��"O�aR�؁*�����!�"d ���P"ORe��`���� 0a�i�0ڰ"OF�B���(v$A� \�uYH ��"On(��'<�lhb��ԅ~EPaB "O0�'
��m.j@�@�I�_34��"O��#6���A_�i�l�*.���"O4d��K�;�J	�T!�+j���"O��O�(aZm�K)^Ø�˵"O���M6'yl�+t*ָ���x@"Ofh{�'˹a�����(�%>�"�A�"O��J�g��������3
9br"O�0��$E�v�����D�Yc�A�$"O�� �
te4�0$�����A&"O��4N�#-V�E��D%qM�Y0T"O�$ٱ��c�<���fڂ7Ӡ��`"O� ���N"!�Ę�℀ ɔ	�B"O0�� ���^!3�#K_�(%� "O� �uX�,�2�['��BG"O<�@e�XN�ǯ)q~Y�S"O���2!�;�`�:!44|���"OV��&�	����e�#>�}ۓ"O2MC� x�Hj�A;:����$"Ov�xp#�_SJ��$��s|�0h�"O$d'�b�(m(�Hң"_��%"O�)��cϏyP�chG�X?�e!�"Ox):q��>�� :aG�(2��p�"O��X��٢9ڝ�R'�p#x�z""O(a:gJ�_������W��łG"O:�0b
*[�6�`�H��ا"O6�a�HFWI11dĞ��u"O�����TP��&��W����"O�MH��K70xD�SC�<(��б�"OFA"aP�@�ɘ�"� �N��"O>��ӣL�E,"�
`

�y�"O,X!����g>�b�#\�q�6�!"O� �E�1A�,0Cց�J�>E�P"O ;4��'�i� ́1�H`X"O�,��+�G;�1�`�F�Q�\Dc4"O �)��$�R9a�4R}R"O"D�n^>Cv�L	wh8@J�-
$"OZ �)T�mi8���6 :��"O�D� $��1�B��+��D"O@#�Q�`�!���k縹£"O�k�6R5L�c��Y�)��!�"O&�h���;�5��L�,A����"O(��dF��w���bfGS@hL�"O(/)pt�0�H��\Y� ɵ�䓘?yӓ3�B934x��ϖ	z�Џ
�y�*G` lذ�E�d��1���y�&��B�l�e9k�D1��y2@� :����4��Y�P��y���/����ޥ�)P�ŧ�yBb�3*�=Ӹ|)R2�̒�hO`��O"|2���3Fh�Xe�� Jp���\y�'�<�x�O�9B�-SԏZ5����'3��cS쑱P����#���@b���
�'���_�ֈ^��Ҙi�F��J�!��ɏ4N^��%�A(Ec��@�K�j+!�-7EЈ����;J�5�'��b	!�Y!,��Q�7G�m*t�1R��^џ���͟��|
&HV���H6�\�!B�f��B�<�b(��fT	�%��1UR� @}�	n���O��P��a�;9M Y��M�|���x�'E0���mM<~xrU#F&ױ`��q�'B�)�i]�h$b�[�bMkR���'�⌚��R��ۃ,^D�9�'���SAA�p���@��P�$��'�	�ff�<��$����8xI�Q��'�t��ShށQr,Q��Kɗк�r�'z��p�͇^�J!�U� J-<E�
�'a.�K��M�Q�(�A'�6���K�<�fÕ�q���-��#*�K���K�<�0By@"�����k���p� �I�<�af��l&�9u�ٜbvBa�B�Z�<i�*��E�j�@���EW,� LVy��'�d-�� �[�:��D&W�tJ�d����)O�g	�#3�$@��&�-2�l���"Opt�$�$�ժ'&=�`(R�"O�Hu뀛�XL	��@�2_.5��"O~q���6����[�i�"Oz�1dAU,g�~�q�N�=PK68��"O� ��S`��X�҉�m�`6�1"O(��%�<]�p���R3r<��"O� ����~�f�bd�]�.�>-�$"Oh�p�R�
Y>L	p�G=k����"OlYb7G��_S�Ȣ�#%+��x�"O�@���6([Q�8c��r�"O����:jC���Vc�u�X��Q"O0��c+�tu�x�>Ж(S�'���!ؖ��@�E�]ux��mC�4V�B�ɞ����S wbf�36�8Pf�C�!���-�qTB�3U��3�zC�I�3`��xץ�O n��I^�/�JC䉤[�< P����F��E�\��8C�I1:<LH���`!e@қ|��	��4D���Eٕp~��P@̩谁U��OP�O*�S�Oȴ��! �<�P�A�](O@���"O`�We��e�v5�DM�f+���"O�P�ٺ	X,1&H�}F8��"OLE��8|E1E��xcHpv"O�Ԙ��M�o����DF�=2M:�J�"O�@:�'JC� M (�c7����'U�	�(C*�o�!u�@�M���=��څ��@�X�'͎<����B 3D��ȄϘ5q��aI���e�0D��:�g�@�Z([f���L�Z�{T�-D�l2��ͺU�\$���$K.l���+D�0��/رo&�$��(Т+U��	.D�Ly�F"�A��
����g,D�x�pG��D�����ѣ]��5:�$D�0x`
�W��(�!�=��$�=D� KP/�"*<�I�JۅW�L�(8D���ѯ��/��/�.k(Dp��!D�lä�R�0�2m{v%Lwr ��'+D��K���.-���#�kK�aP<k�.;D�� s�K�=j� 3Ź<@��D7D��zV�Q�3<�1�A���J��4�@� D�Ē��B�`�,�rn�Q��>D��z��]�y���lZ�/�b �'K0D��Ty.q�m�*n�:���,D�l���_&g�ز��*�$��V�8D�����@"������(��1#��*D�@+"��?N
|b�d��.D��TC*�m`�نᓥ��!�K�.Z\�ç.LC�I�{څXw�W�q*JU�0��wC䉉;��L�5@T�p�r��0:C�ɽ2e����ϮI����UL�Lg@C䉧|o����M%n`�I�o��B��'7T�T9�匀H�H���Go<C�	�c��E:���u�N��c�Z�H�=!ç2����pfE|^v���3d��u�ȓ
����� ̰*Ĕy3��ƬM��=�ȓO�Z4�V��;܄�My�Ʉ�_ՠ��Ԃ�c��I��� 9A�����r )�2��j��d�رK+�P��d���S6$^)o����MIfu$���H�v\cB��LZʑz$�n���ȓl���y�j؅,72�s����m���w��W�թ@A^�M��:� Ňȓ=�.L��舂M������@	:�m��t�v4����Wjp,p�(�~<�U����X�텁lm*���(A~`h��d����
�\U����)J>�u#"O̈֌ƌ���b�B5�2=*t"O����Q�}J���.̞h�<Q�"O� lZr!L�rȢ� ��p���"Op�k�g�<S� ��x�^E�W"O����Vqv���J&0%B�p#"OF�(pM�	p�N�s���X�4K�"Od���0H�L�c�E�p��Y"Oؔ
1c�}��D9w�+7"OU𑃞��n�i"j�6	p�"Ob}#�$S�~y�9�(�&8�젇"O���DB_� ����mؗ����"O (�JN�(e�	
�
�m�q"O,H�3�M� zZ����7:��jw"O�T�%!<Q�Ɋ�`�o�}��"O�ي�� 'qĤ(!�B=�RU"O�1�o6KKf�
a���8Qh�$"O¬�E�Ǜ ��x��L���R"O�m(��z����e-آWK�dʴ"O��Z�ꌀQ%�USC�̨&5��c"OؙÀŚ�kJ.\�4L]0j*���R"ON僇+]��9�jܓ;��If"O8�I�N���a���?{���"OD���H�O` 1Brj�9U~t�p�"O8`�ć��6�F�1��ɔhzn�.8!�dW�f:�
���zǒL{D�@I�!�D;sK<�j.,j����M9H�!�䀕j�r���Y�g� ��Ӌ;�!�K,B�F�R���l���Co���!�� �0���� �H E�T���d@�N�!�$�(pc�(Sa�T��9��ތ9�!�y����cJ�0�&�r�cO�!�D��xUH���Oo��($H'\+!�DО#�h���"Yb��Y�d:!�d�4e��\�"ȃ;_
L�wf+S�!�D�K�ԠAV�%�ڽ��3s�!����+�̭��G�'�m1@�J�!�̈o <-�r,87Xͨ� �8��'-a|�����LB�|��̂'�̻�y��	���{�/K�%��e�G&C�I�J�.D1f"̢�r�C	^�V��B�	2=���1/)dOR����� |8PB��;/a��q��DW:�[sG\�=U�B�I�A��b@ϸ`e�"o�9V�BB�Is��YQDP�b@��E�Z"�x�O6��9LO����Y�0v����ă��4{�"O���4�®�Ʊp1*��P��Q"O�s�eR�D�`�Ё)T7nƪ� �"O��c��Hj�ЍS/
Q&=�"O<����0��x����VDʄf"O����@�-�F�c�Jn&�ɳ�"O61�fo͊)�Q H^���hr�'���'��'��\S�c5s��+ �sE k��5D�l@׍���1e���	;@�3D��1 ��n�@�����nF����>D�L{�E�l�ޘz�m��e�Q.!D��K_�}�v5�"��,gF�T��� D���4�
'G
�X
�

�Wk���+D��h�n	(pa���ƪ��z�@ gg�<)��?I>���d��j�.E�3���Z1 }zT��.I!�d^�a��i3�_�`�5�DOD�wC!�dٔ	��yÆ
˵O� X�"�¥<!�d�6��dS` ��F��I`�C�'!��7bC�+�£n�6=���._�!�ƻb%q�l'GN�)$.�'2���]��pl�6���W�F����?Q��?y��0=)���	���MkL�-�7�Z�<�  t(f!�!d��dA�#F��s�"O��eO�St\��fi
E����"O�����4xF�KZI5"Oʩ2�ː�dO���3,�	��@J "O�a�7D\&$x\��[KL��a�"O$�b�NP�i�<AH��6.�9h7�|��'��!@��7SB�+���>�����'�� �jP��`�D��3k��[�' ��9�ˑ�bdh� ���07_v���'+�6aJ�5�`���x��'K.T�g�hp�s�N��с�'%v�!ъ��5E^ms�ɈK�^�<)�&%<�z�3U*�!wHH�F]�<�S��<ȉR�ϝiiN [t�F[�<�� �{z�9��L�q0xaE�[\�<����'$U ���@_;
D�R��q�<�׈�2�\L�vg�_��|�N�n�<�n�$V���@%m�/����n�<��"ȋM$�!+�jM�S
eK0ǁm�<����7d�R�����3WE���NUe�<I��ԫ4�ek��/Ԭ�8��d�<a��Ϩ�Eq��K���	\0�ȓp�4T���4��d2�@o; ���qޕ�K���i��B $��D�Ri�t��O�z���ȅ|��$�ȓf�����(��${��8+�.D�ȓ?�e��+�)]̰uCь}����f%��p"�,l�T�ъ;�VЅȓy*�Q�`�Y�^���	79�=�ȓ"��������!���<p��X�ȓ�sR�?r1.eA��T�+�H�ȓ3p�(�!��l¨����^~�ņȓKF��w�сAZ���ڱ+4N����f��BN ��Ӧa�.D��p�ȓ`�� �L�#�����'m�i�ȓ]��y��� ����B�!+-pY�ȓwԢ���c�}}�Ec6n�'t�j���HiƥY��E����N&+ì���a~f��c�.3!���uE�+Xּ�ȓ\{�!�v�Шk��uZ�)^!v�8�ȓY`�b�К,� ���D4 ]��-��i(�!�+`��b����t�J5�ȓU��썍>����ҡib@�ȓR Pf���O�p��)ŚxBP��ȓgt����A ��y�Fj�2Ozֈ�ȓ]Cn|�dmRA`У���<M��H�u
�钻?T�g�9ЄȓV䔰���U�Ÿƕrg���ȓ"��UnF�R�B��5�
&uq4y��=��\Pw��t�ĥ�f��8V<�ȓA���H��9�U�m�m?D��~������K�!�l�8���*nF�ȓU�,Q�DB=8I�� E�iO����
�d�z��ar� �tkG�{����?�H�J�b	~�(h �U5κ��ȓ5�,����zL�gC�5^Y���X�ؔEW�7��D�Y����ȓS5�Az��=!ʥPX�Їȓ5 *uba��3rv�a
�>K?Ь�ȓ=6	��N�����g>�*��ȓR`�5�>.�A��O;q�n\�ȓ{�V���OX�d6�h7'Q>#U\	��"���GQ�A������Z=�Y��r
T�U�B�����f���,�����S�? ҅�ĆA�h ��@�2��az"O:�چ���M�}��O|�X�"Oj=��E/
��|(b%֭[]�u�P"OF�cs���TpRg�[�HJ��"Oj�fD�D�8�9�툍lP���`"Ol���� }NI2�ҡOn�ё"O��f@!bŀ�.�64����"O �+Ƣ:u����M5(||�p"O:8.
a�α��+�'&J<�(e"O(]�A�֪���B�aI�_&Խcq"OR�/��`KDD]�s*B�!A�	~&�'r�'a�Dl�D`A𪙈��ڥB���y��Uq`�xaN���ABG��y�W( sf�yq/ֵ�`h��D�yb��!A;��A`H�	Q�Q�q���yB+��y*�4�#|<0�5b���yR Z�zVT�B���( >�˒!մ�y��Kx,Ac�D>z��Y"2�H%���?����T�H�.R�E8Rm5s8��q�÷�y���|�)!@�<Y����ћ�y�@�"�9&hX-<�d���?�y�Љh�IӰ�#;�lq��Z��y�%�3Wp��#P��20��`S���<�*O��<���"U��?�r	�`Ě�v�U��x��9���U2iR��q/��u��'�0D{���S�td�@��D<X�8���?����d��,�#�ܜ{P�)�����v�ȓ9sְ���Ĉ;H�	$D#s ��ȓ(��2 H9~�X�2 ��k���ȓ��(�$�߉���lQ6� G{"�'c�IX̧��d`a�Y�drb�x�G
[�LI��V�H�9��^7�h�x$΋ ���vu@h &�қK4)��"r-��ȓ7����De��b.����'��M�ȓ*mLaJ��;.W���_"]2���ȓP�p��D��X��A&�նG���["o�Z�:�h�������8<O
"<u�6rM�`Zq�:h
�a[ ��R�<YAe-0�A��ߋ7��poL�<�燺E.�j�&\"~���E�LP�<9I��vD���׳,C�!�F�d�<Q�ț:|[��m��n�~��jMy�<��ӤL�6��ެbN`9�V��Z�<��޿-=(q��ǆ+�n�2��OU�<q���P�R��6$���+ѠCP�<ib��n�zA�BᙍT0P�HK�<6c�;`;��b�o�IΚ�Q�I�k�<)f�)8s^�0uh�`�*Ë�b�<)u�:y�6(��"�*t�X��IOe�<��	.,�z�M2_t�	�aKG�<AC��;2����C��vRdi���z�<A�K�@꠱��C2*��I)�$x�<a6�3,�t�#V�V�����-�s�<�)E#ag�aՆ{��P5��d�<�"-D*ż�sW��z~�A�%��H�<��E�,��y���пY2��C�B�<p������`��=l�9�WNx�<�B�9�r���&\�aC�� �v�<�r�"	� o��M�.doΟ�y��N�8Xԑ�P
�\��1V��y��ـ<��xpUD�Er����$��yԎ\�t��ΩR���iѯP�y��F�[�nDCd �&{����1�y"���6aN�3#����)��_��y
� t̳��P�C��h�b:���#D"OtU��(C&h%;��K9n���E"O�ug�
�J�I&�[����Q"OBq�AOD��+ɓ� ���ɀ�x�<�D�\ɀ�h�,�Tբ��i�<�q	� 7�L��Q�\�a�0��u@PP�<��A�)%Ԩ�+΃8�ZKV�L�<IwA@�d�D+�h�=b$�eC�dn�<A�Lڧ|sDdB)���e�U�Jm�<�v��U�r�8D��j �Bu�<ac�M�7,�<82NC(�ґ*��Zn�<y4-�i, ��&#�!Z錨�B�n�<E�<�������\̓$�j�<!��G���s#I<^[����D}�<�E��7qg"E^(����5)Zy�ȓ;kF�	�O�P*�	Z���
K��L���:XcD�П=�8��/={=�T��=�6)���u ��cB<����ȓ#�2��2�.�^�*�N�8 XX��Z�q�͍�
 �ϟۘ�i��6D��PdH��(��JḲy`�i�5D��`P�S,9����PC��Kb�)S�L.D�(�E+C���Pr�D��!t�%�!?4�pYu���__�|�1�*ui�����$D{��IH�	G��8'�P3v�J@��TʪC�$:]J82�MNu(<+0��<X|C�ɠh�� B'ΆF�\1����jU�B��	r�|�bR@�t�4�"��\�lB䉶�R�.9D���R�>%ࡪd�|"_�H�	S�O�R "�)�*;t!�S��X˲9�ߓ�?���yB��
~����SaH	g�yXV"D�y�%M9��r�j�8���J��y�8 ��B�N��y�B��C��=�y2(���p5�#`2k T��'i���y�oEa������Hd��7�_"�y��?<�$���A]�p���$���O�"~�6�~0��E��^�B�zu�V���<)g�̵0Ѻ1��l@�<Hz���V�<Q�B\�=gK�A�\�ulR�<ɑƉ�4�N=�Ά!<�� ��g�<1���'Q����	Uw���
e�<�q��t$��W��!_��W�<Q�H?87���d���
�J��AS�'�?IRэ�0VM(��GQ�Q�.���ԧTD��ğ�o��8r k	�e���J�g�.T�!�\�'t�s�*��ɸ�	��گp�!�DA������Ia����R]�!�$0`ݺ�*!��T�8L��fG�r=!�d-3��):u��1"��������!�$Z�4G�����7P��q&�#Ya!�[,S}ƨb�m5�L�ZS��)[!��/c��P���Bh�+�O�VB!�$��}�аB��� bS0��W17]!�ĕ�'�\T�u��l="���R�JU!��[i�6�4�R16ݙgoL;!�u���PP��
Tw�m�wd��!�!�$�<�v�RQ/݂x�032�*=�!�B+)G>}���]���wE]�i'!��S�4�`��H�-B���`$�,!�$�+x����f>P>�(ʣ���!�Ē�j�:�	٠c=�Ess����!���
e�	���ܥkB���% ��!�䒿FP0�R�dڣN(4���/G��!򄐚WN�F*͞4|���B�ǝ��{B�� b�y���>iǴ@bD�
2*����"O0ԑ.�[�D<%�ۏs���� �<�S��_^z�� �ɓ�3L��'�!�$�X}2�TeVY(+U�S)�!�$�8&���í�$?>���	Z�w�!�d�2g�!�ƈ�y�޽�a(��;�!�AZ�0�"Pm�P	�!�$M�sH���&�V^}U��h�m�!�D��"�{�	�*x��w�Щk!��W���"�i֧�+�Ġ�F{��'�� RC��+	�ԫ�.ɿ6����'02�HD��(z�t��)�E^����'�l0X�c��̃�.^
?�D�	�''T=�"M./b�q �EL����'����D]!0l�p�a�4��ر�')0��_��h��G�)���'{@@A�͜X�D$�g�Q)�<9�'az�v�'5~H0dH�$`2���'wh�	��������K.H{�9 
�'q�I個�k�^�a�ћ;$��8	�'����J7��m�r�M/1�, �'�樹T�&L�:9R%ˊ�4�^��'� ��%��1B���Ԯ�1�l� ����<�� R >JT1���J�wvp�wd^��y�5_���2�*��$r�Я�y�+���P�Q���@HV�,�y��T;'��4:��L�yz$@����y�e�'$�vY����(]�`$�L��yR�M��I@��M	!�����I��y�I�<^\� 3�K� 7B���)F�?����S��H;���z�����BFF0�#&_c�<yD
±Eb�0Q�{g�`�b��x�<�.�9�1�2hۓnH�(E��o�<9Q��>�^�" /�N�D�H�j�<q6���_���#�' �1J��Qe�<A�)�(��t#B����:A���P^�<�aM&q�Zek��p/���ICXyb[�H&��F���Z"OU@�C��+WIz���y���X�RD���Tw���ˢ@�
�y�k��E���X�o.�[�l��y���6�$�r�`�9k�X�&!ț�y�H�mt<@���d�>�X����y2H�
*�! �C�k� ң�۞�y�F�`����� k5,T)6���'�ў�On��ف��%z����5C�����'��k����UGD�U;?��}C�'�����X\Ȳ\Pe�hq����'��q�G�!0���x7nR�`�x��'��A	� {���S�ə]P�;�'�8u;�@��u�� D�܌\�p�
�'N�a����J�
\rc�Q�[���j*Ọ=	��Y� ���dihU�Um�KJ!��C���1P�Wx/���f��/D!�_ C�����Er-����� Z!򄃔W8��#�!S*@; �K�|a!�E"D"J��fk�qf�����`�!�UPdDdځ:B��rG��7�!�䛷=��:ꖀ+6��<��yb�|R?O�mpu��$\Ф h���}`�]B�"O>�2� �*N�z�V�Z�=_��ڤ"O&8Q�l5�X�!�<M��"O^�����'M�*��$��L%4A�"O2�Zq�˱j��de�7k��sO��`���+q�}��-G�$�84���%D�� ��Qcހw+�k�()j�H ���d>�I}�_�U�K�=˴���i��,`�-DB�Sx��Ӗ�� ��䐧�P(9��C�ɺ^t�c7m.AYx���j�j��C�I� ���+���1,��tY#���j�C�I;{퀘 ��*Cht�f��#��C�I�*,��woB�*�Z�;�U:y�C�	�\���H�K�+?V �3o��p��O����6~H���A�i]�x���!�䐅SVR8�GB�5� 蓥d��E�!�D�{��xq/�?�� �Q��!���(yP���`U6��x�gE�:(9!�Y�k����+���j�#C?	�!�$>V�t���g�5��x�6�ʗ�!�䀤��a��	{�����L�u�'�RZ�|F{���-�H��P /�b�xA��-�!�DC�!w�Q�ׁc喤w�՘+U!�$Ԑ4<�BC��]�"D�1a��A!�D�� �&�T�W �l����B2#5!�A�6XD����H:l��I	�.F!�D�7)��Y��*�dɃv&�!�č"O�zH@��*�P���I� ���_y��|ʟ��~���o����ۃ�[1���HE.D�,*��H\�����|���@�<a���S(c��� �̂y|h��I�U�B��R�64����	SFD�94&�:t�B�	�o��d� ��~%��:�
��p�tB䉥rDi����@F�iS�O�(hB�	�ub�B'Ej��s��͕Rm2���O���'�?i�O��3�)!��`�a.ݒZZ У�"O|�q�[�Բ�A��\%lINq�"O���`����С�6n1� �6"O𹫓+�)Cy�UG
k#���"ON��6�E�v
�t�����`�:�"OT�'ƍ\�v��D�eFb��"OZA @hJ�V�,h�n	::��@�"ON%���4ONa
fGܱ�R�ɒ"O�TA��V�<Ǧ��Ĥ��*F"O�]Z�EVL��|�W(x��AÁ"O�� ׭߉R��Ex�ӺWs:Y%"O0܈ AD�J�t��O_�2\�&�'���;n�n�����~q@��C��7e�C�I�3w�{�� �z=9woјVB��2C��cA�xƕj�@�+�чȓ^P�(��%��E�Bj9�ȓHWx���O"f���b����j܄�5��d��T�D챷IRt�Ȅ�?SN�s�	3���)�V1u Ą�or�H����'L�e���%�f	��r�L)�6�׃:��iBTM�<h��9��N���v��5�����mR�Pؘp��Lɶ�����%yD���&k��ȓ7~�u:���$	��A�������ȓ}vDS⦛1N�������.��-��Qtd)qG$@�<�.e ��I�-KLE�ȓ(��:X��#���<�
b��[�<1�F_;q0�!å)�"}��=
��KV�<)s%�n I@�bP�x@�s�_mx�<Dxb�
�2:�(
�B��;S���?i���*�T���A�
$a*�.py$��<�.���C	tM�Q�B��N3�m�ȓ1��m{C��pp�p�ħw�`����,|q� V�����U�BV-�ȓ0µ���֝] ���A�]��9��S�? z�C��6CUD�P �]�JJl��"O48s��6[l�� T#{��xq"O�8zWĖ�G�RT��oe���Ä"O�\S�i� ��T��KN�х"O��3P�T &���x���?���"O޹H���x2.���˅��x�+a"Ox�h���۪(R��w��z�"O�aꓭ	�Nj~у��I�ʬ�q"O�8k�/8���u��7:���f"O��[^�E�cb_�Vܓ��E��yR��*� qxP��;G�`u�D�?�yg_D$X�s"h��u�S�X��yҨ��-Ibe;�㌯c��Jn��y¡B�S=��[��ڊ�
���.҂�yBD2���`�E�7��D� ���y�N�"H��� 舫x�>��4���y�fE0\�@"� z�h���$	��y��b¨�[2��%�p�{t��y2bʮw�69s�ߎ'Pr����y���A���K��Ҋ�a��%�y"�kp͘�%�/\����C��y��"jkXiA���$�S���y��(# *��c͉I��#S͆��yBʞ<�B�
��ؖ:�ڜXrƬ�y�"
�s�\(s��.�*� ��;�y�㌊E���f'�!2�hy��9�y2�	;n�xi欚��ӯ���yB��_�<�s�#ۛ5m 0A��y�b^�=��(e��Z��ii͘�yҏ�#��त��c��0ϛ��ybm�~�9RE��'-H�����>�y�B6Ld�m��f'(��(k`͜��y��x��)�`e����H�&�yb-P��1bK����c����yB�[�3|@y.�8�3�$[�yrE�/����F��)K����S��yr��2c���5N�,�b�9'��y�ԧx�N�JM:r^|A���R��y����o^�[Q�5a�t���Ϛ�y
K�A����-9e���Ĉ���y�F�e�H�ە	ēU��Tf��y"��Sd�FD�N�(���E��y��M�`�0���&��!i�2�y���"���q�A�Y"p��y�	�!1V�јa����~�y�
��y�钯\"!3o�E,�6N
�y��#"���p�Ѽ��C�G�	�yRB�:��iك�M���Eu�B��y�$Ffgĸ���W���q��cؿ�yB��/Z������P�T -?�<�ȓ����Q"�.ZF���k�v��?�
dR4.�8L���ہ�ò~�"A�ȓP2�xCc��`>�a;���+\=%�ȓZ~D����h��S"h�V�B}��ΖԳ6�ޚ6E��Cѧ.��ȓ �Z˔ �`3J5�GX"��ȓH��X#ϗ���	�
x��!��Z��5`v�_�$'���b]�~�a�ȓUB��OՁC�H����.J�`��%
)sT	������̫o���ȓp������49 �C��C�xȘŇȓ7Tl���@��cJU�#"�+=�n��ȓl�Y��k\�5�Q�i�(7m�X��/�xj����jba���K�����S�? �ix��U5¼�XR��e �X"O2�9CƹQ�����G�\1U"O���	D�-���:��s�NmiE"Ov�CDg�tz�xrw@F�Ԥ  "OV�0p��O#f5� S�W�Xm9�*O�%��K�C �e0Wf��`��C�':N!	�ɇ5|� p镡�+��
	�']p3gA8%�Z��!��Y�-2�'hRf)��j���MŲ���'��I���Yz��$3'��&0b4�H�'�&�k�M�&�`Mi�/¨W&9�'��ܛ�J�LN��{��#���'�� a�O�&]P�#R��/g�H��'���+�E�*tj��A��Z�΀�	�' �uJ�n�+������S�}`	�'�`�1 �35
,T��E�L��QA	�'�TB�̈́�-��u�EAS2F�����'/�yȁlȂ�t� Ƭu�L�8�'���r0m��J���z&�:n���R�'�R����aR*,�%/er>�I	�'4Р���3m�؁3�	�|���'��[�)ˈ?t�У�C��|�9	�'4&�3�͎j����Un&�m
�'��h9#ퟵw�v$�U�W�|+�']�0�V�4!/��D�H�~=�'�xy��A��HGIjt�{�'�Fᑔ��;
h��Ʒ5b�4+�'��!�D�ƶjg½�`�+X��]�'ot�K4���kfd�ȶ��HYlx�'�r](h��M�"h��ϙE�H��' Z�h��(p�0�;#��k��8��'s�
�.�<QPI�BJG2Ոq��'��|C%�E3E[d�h�E�R؄��'�y�f��V ,���a����'����̀�
{�.G/O�v5�'�Ax�$�'/�hh��K5R��'���",Ӽ`P��r,��H��x(�'�T�@P)A�d�C��SI��ق�'�x9��:�֐�
�=7]�5��'�n9E*�������G��\Xa�'�b*@.��Ur�lw.N�{ݪ���'��u��-{� �v�v���'R�{���tA2M���pv�u��'J�:��DJʹ���Wvb�`�'���R��ۧ/�L��E��Q�r���'#D���!N=#��۱�H'����'lF$K��A>?�=���	o����'H$��ҁY�A.�i��l�_ �y	�'����@�T20�e*�Yʎu�	�'޴[��Y?8$��;�J��`�f�(�'��]�l��qh&�Ӈ�\;Nyb�'،l�5$ۗ%�|� �=U�P���'G�8{�$Z i�e3L)nx	�'h"�!Dl�WD��@�II�C�ji��'�8,F,hj<KǤT8����'���x�N�F=xx��#|�>�	�' )i�l�N��uQ �u���!�'^����9VH���R&z<�̀�'�:؂#"����}A�� r]J��'��P��\|��-�`����D{�'q)�aHйC-L�g&u��'�pY���ρc�����'%v=���'��+㧙�<�@�8jIpEy�'T�QA3�+��؇T��h[��� ���֛s�<���_�J5�1X�"O6�12i)yj�8b���(��"OLe $��0� "֊?1f���"O^��D/�{$l	�ֈC�B�ȩ["O���iΆK����ĂD�h�
l�P"O�y �eC��`[T"X'
J(�%"O��x� ,9B��0$�ݺ7x��"OJM�ܬ'G�q����l��I2D���D'�tv `р۷	����.D���6���^�:=�D#2��␈?D���%'��QC5�ĳ\;����:D�c��ܺ\ERm4r�\�j��#D�l�Ƌ��N֙@���Ym��dI D���W�B2l��vV�O[`�Sh>D���4L��K�������q�8�k(D�4���2IA�#^��X4�$D��PJT6���E%�mi��"D�@hD�f�ȱ�d�4uJq�;D��QCE�k�`��$�7�
���$D��Zv��+n���0�/Z�}�,�
$D��E�Z�d0 �e �H����	0D�`���"4A|��� �1��0�6�.D�ȳ��.p܀E�|hfa��o"D�ar),?�H3!�%�&eS F4D�؀��$�����A�E*H��Fd&D���.3���!���\�`9; �7D���'�+*��erP�V}ӆN7D���@��
 �	��E�)2�y�F7D�H�r%Hh��s��Ɛ.V^�(�6D�ʁ!@�u� .U��{�k�r�!�91,��шLd�<�h���	�!���^�N���]$�����?}!�[�r�D��횰�J	��F��u!��P���K���6z�,Yc�]:[�!���	�(xh���(l��P�^�^�!�D\�f����1ʏ]d:R�\ !�S��dA�A�C3�� ���#�!�W�"-P"m0� ç�Pz�!��3è`tk��hJ��yB`��d0!���%!y��]��`I�C!�A�@��m�&BC�o����![��!�D��#|p<�G�d����i�)'R!�d�!�<���ǃ"�|��phͤdF!��D�lKpCs�£|���S�
	�!��1L,~P�i��>q�ܠEG؆]�!�&d���P(3b&I�i^�!�D�~�x�2'�:N6 ��O� �!�䎩��؂ ��	E�}sc�G�!�D��,��$3EG�8+p	@�B��f�!��D�Fx�Ƌ(Y���d(!��3H媤�����LUڷ�͔&!�d�?|�d����^4$�qdW!���B����i�	]&y�����!�ē�GZ��*�[��;#��_�!�Fg�%h��F+uN�+C�j�!�$��t���,Q5��i�wF
�_�!򤑻D:n�z!��(`2�CcK'c�!��+x�b�hQ#4Y��}���2��=�|*L>�ȹq"�E��#��\�<y��M����7 �U����OX�<� ��'��u�3C�>���P�V��D{�n(0^����>'�`��Wװ<���$�6RA��s��D,����P��	!���
�8�e�Q?u�ٺT` 4W�!�� Œ笂�:�Tb%̦`Ҩp9@"O���u��D��! �ț] �<�q"O��Be�.B�L�r�� h��=���I�+��?�`a���L����j�b� ��4D�pa!J���r��=rbU��J1\Oc�l� Kˬy��X�`��H�r ��(,D��� A��6�`���U�,�d��&*D�lwIW-E��zR�eRr�s%)D���*:�V��anj���$D���E��G�>����T<>�Id%D��Y�
��ne�����6$ ��e�0D�X����$�H"a�)d;�(S�h|�$���'�ɸ�ħ��'�X�8dd��n��)��B�4(��P�'E�`���jC.p���A���iL>)Of�}�<.٠e+#*XQp��߀�<)N�<G�D,��T8`(���G�MZm�C��M#
�'���� +��-T���KH3�����'�ў�}"��|sZ���_r���3oWH<9^��z�/N�,'V�QT�C�u���� �����	�v���9M�4P������>��O`�	���	 ~�6}@n_�m�hu��Bk!�܂|L
��"�t_j���
��1O��=�|��R�j 9��l���LIy�<y ��4\��֌ϊ�zM@�Y�<1���>��KF8�����Є#�� q�<I�"��9���I�
����w�i�<y`�Ô^�@�+�BՍ�B�(է�N�<��"Hx-�`�G�E�^$)�K�<��'M9L��q��+5BX�h��$�H�<�'��kZ��Gřm_`�e��D�<I'�N��UAũ|�6)+d�C�<	����ء �Ŗ}<Dz$RC�<���5t������)k�dաs��E�<�qD�9<"C�?n�ع��c�A�<Y���:YZQBCQ�7��t�JC�<�,D+(;V�P���2�h%H�\F�<Q��AG��K�$Z�h�>� �C~B�'���WL�/�j�@�JʼC��4��'��1X�f�4���ƅY46�8��'R���Eq9&j�,(�H<�����Ц�4���ۮ��պ�Ɨ�!��A<l�X�{�`��~����睽F�!�dD1p�DK�� �S-Vy�4'���	����I8�1F��"�ў1�E<W�����M��(O<��D 61����7�C2��e[�#�<"�!�䚖DMp����"T:��" �!�dʃ$���he�D�C�,�=T�!�d�2lk��O����.�!�$��ff�s�B�|M����i�$N!���GtE˧EB32�}��>=�}b��>��L˘N�0:�C�+:�Bt�A)F��y�EH��=y��M� vv8! ��yrd׈)֨2�KY$�ʴ��旭�y�iّC��T1R�##O������?��}"�'�g}	�3,2]��%��)݆���G��yb�Ã;�D��N7sXƇ��y�L͢u_��RE��l.I��ڍ�HO��'
�$<}��F�p<�DD�0�xhf���y�`�>%,Tl����w�:���Ē��y���4Td$�a�[,BO���8�0<Q�R�'��U�t@S�?��bsc�L��	P����O>���" �8Q��Q�ƌ!:AQ�ȓ'S�X0�Î\��	S�a�$����ȓ$��R��[�z̸��]"��$��	c�S�? ¡PU-�%?	�x��@V���iA"O	�"�L-���lZ -4�"O����a��z=2p�V0���O��E�!���)cI�'  M
�-L(x!�D i��aȽ*fvU� ��= J!�	k�$�òĞl3�y�k� `B!�d�&��d��cY+G2��b��/�!�d�ub�����V8(��:�
ѷi!�6�����W��k_�dk�Dڐ�p?�2��,E�>[w@�qv�B��H�'>�YsfR5��5{�`Η�Ip�'�2�Z�ze1��gʐ)g\�g�;D�L�p)\�ߢD���M]��1�&D�H��b�q/n��O(౰
$��hO���i""ѢL4.ղ��Ħ@�e�RC�ə?�����.�~���P�
�+�2C�ɡ[Xq�&�(p\ְ��f&�B�I�H���`�E$h����#ڇ_��	_?�-O�	ɟ��R�&P�58I,������V�<y��Q�T CUF�Y:.]x�G�B�'Kaxb� &�DQ���ip�ȸ��O��Ұ) (Y���-BF��U/���C��\��
#p�X�'ۍiV8��퉾��'U1����{���K3��+0� ��O`Hi�,R���J���7IVMQQ�'�O��&.���;�6oL�1I�"O|\s�%[U���`��C�<��cü�PxĜ
H���j�wV���)�#�yb��oƈ��"�̜D �xdC�7�y-˘<22m���[�\|�T�ь�y��	���{b�ı��䉘��0?Y.O>勶l��:~$��5/�p��+��x�'��@ ��a�<#W��/yq�(+�'m�YE���7�h�`�9w�� 0�yR�'�dP���%
'.����u�L�RA�R��z*�>��2}�um\%���:#E�sl�1�'��+\O��J���9$��q��Y?&fxP+��'P�dU�W;�)�D��y��)�3��)c�.C�	<�Ѓ��J7x%I�Ĕ7q�?1�'���)P��߰t���K���,B��C�"OL����.B�T �i�6"2<��_� ��)�'YPL� ��W`L*��F�|e��Gx��O΢=�;i�&<�fƠL$L@�WO�i�䡅�T� Ū�cJ��AaoD Cs !��4��()��^7Y����a�V#�$���Ly��rV�Qz���4G�$��j�HK��x�IA��y��6��Y�DA`.m���y�N�O�����Ư[��9����$�yR猎*�Bd��?e8z�	�`]���>��O���ԣ-M�\�e�T�BCh�#"O�Rw̎�
�)�Ŗ%��2T�xB�)���'%���%�X�^�~��fb�/%C�)c��ak4�D�%�|X�4	_�Z�LB��8���Sի��l^4=�0���?�*B��2G��{�hQ�	ap@�qn�4B�	�"^t���낭+4��:�"	Q�B�ɧf��4��A�	����gƗV C�I��Dv#���P؂���V�B�lb̉�b��6�H�҂ڊ�'A<�+��С�5�]?w6����'�a�5�*@�t�0����nUb���'��[��F��Ъ@���=��q�'�� ��ݐ��� L���|�3�'��("'�=����(۾`��H���� (x��B&�t��O�	Zڡ��"O�}0�m���Q��\�+Cٔ"O�iX�!ě
�J#.ˍ>�Pj1"O����84:�6lF���%3"O��
`fа~F���j��g���"Ob]A��	���)Tk�v=J���"O��xH�����E����"O�H�����,1	�o�b{��A"OxXI��̙s���;P�}; �%"OR���-ߴd���H0ɩ�"OZ����G�`Nq���R�/3x��7"O|L�1.݋X_~��$��'E��"O|�h�A޼a���;�|(��+"O,̣����j8Ja�_�`B
la"O<Y����(�\�[��S.b����T"O��@�W9IQ:QAOgnP�R�"O� IR���!��p�@k�+C� ak#"Oh�k���c�DL��J ?/����"O��Rp���z6<8!QӲ&����"OY9�L�?�mZ��͛�.��"O<�H��J,j�=�TX�L�0`"Oj�Q�ݾH���`���@vj!��"O��Q	N�@�j�6#�>�0�v"O$<� j[)
�(�͒+�B���"O:����ǈ&˖�Y���b֒��7"O4\R�≵Bɀa*�/.ڌ��#�'I`�iP��7�Չ���2@�
#�ˑe�޹��'`���� �7M	�E����Y�`y�'�|Y;צ� <��W%I�_ypH��'���چ��	��J��L� ����', ���O\\z�Q��x�
�'�ڔx�f��Al�4��IF!Vxi*�'��	+�hْC(`,߬L�u��'pVD�Ui�/R��!�	W3j��R�'���Y��[XȺ Yg'[�Y�dc�'�*=!���~/�|�FAј_� ��5���[6̜ jy� Ceݫ u�ćȓv�ZpR���C>�К��$B�pɇ�Pi�(8�ߊwp�:��-.�r����𨠪!^T"4b�kܭi-�A�ȓ_��!�1C��S(pC�k3:���s���h5�@@�|�ԃM)����T�݊#�z�132��'`�|��ȓT��UK����E��q�3�t��H�ȓ~-|��ꂖ�ީR��@�}5n�ȓ8�60��
����#��4��I�ȓ~������ A,҉瀏d�TɆ�&���	�"v����Qj�(�\$qB��q�q/��O����qJ�T~�T#,c8�)b �<o�B@3��ț��x���2,u8u�2eX&�@���*K'l�,$�b瓗)Q�aR�ML��x�&�r��	ԩ,�.�
W �)T�� ᪇�lNQ���Ҫ�(ptY�eH��|P��O�����&^�$�dP1C�L�S���
B�K�<m桖'tJG�(�3���2����S0Y�]��j�=4�oC�:
<���h���#
�Q>��/��h\����B�IX�ےkO +�m�����:4"���'�@ys,�%I���"DіUtn�i3n4�JU��� -Gyy%���4��SkIyr�
*:�Ɯ͓C��%�4	�7f�-�� \����	5�
d1�P1v�>!"$�($C��zWb�gnr9��Fؔ�
��I�w"*i9Ffgg>J�m�O��ZwB2��Lh���R�g;�5�3�zCQ��w$�lȈ!�"��b0���E�x@��I=~���%��x?���WUA<�����[�b��JyS@@4Q?͚'�<W�'���۱F�As�֫S?�!��I?�p���d 2#~�R%�� {���Ñ�iӾ~<~�Pg�I�v&�m�� �i::��$p��@2�♷(�����3nS�%?Ѣ�k=x{�i�CG_W�@��T`Ȯ|�����g;~�%)E.eu%p�O���>r�A�n��M����2�x �Ô�tP�mi�.:�9��A�<)��Q�	��PN~*_w`l�B�رy�xA��Q�ϲ���W7@L\|(v��Q"�Alʋ"r]Std�d��|)u␘�Mka䃯��d�S'
� ��s1�}8<���o��\Yqa��UZiȧ�<aUeE�z�J`u��Jcx�{�/FSPV���'R�L�P�J�-����?,� AE��"�]ˡ�Y�:ʶ��S��Һ�%o�h 1H�o)��i��� !�2o#4���kN�<��q� A�<���K��X�Ӏ�2 ��@A�r��g��9m, c�&�`TA1�߶"�H:��	�X��[b/���US�.Ȥ�P�uK��$���^�'�h
�Iw�TR���+@a��)�8�0�G�96m�P,0 �U�ҫ�Vt%�_@P�p̱�q�r�ÎPy�'������h��)9���1Jj����Y	4�R�d�|,@9��It���OZ�R��L�r=Ka����4�{�cy�\��Hǵj�����;a2�6-�����m]�4�Ej̆�����Qk��!�X��BL��:{D9�W⌕.�Ar�ME�Ux���/O�h�g)E4�FɱF.�W��xK�z�Tp{��F�]� -x'��Mߪhj��F�k5t�5
Q q�9�D
'e�|��C�,]� w@]�Oݴlz��O`��e� �P��� 皔;����D\V���K�w�m��k�(N�^`�E o}���X
Pa��b��/~����&<�(
��BI����V)
TdA����#	,��\Z��3��?��Iт �lz��=g�����X��͈6�
=/QX�V��&e��Ʌ)��iE�ܛ�A�m�YJ��Q�^������˾+_`�v.Ц���Ʉ3d�Z�
��Z�SYPU7�Ű+�T{�����"��U�t9H<�roD���Y��0���<˜՚�#åE�F=(3��7�pX� "L�^46\J�*�5�b|�G�
"�����D�X9(CmG%4�bp�BM��uGIS�?V� �s4���ƊF� }�sa�8DN�%�x�C��9 C^ı�GB�I`�X���?��
�)�G�(��ߜkd��Y�*�S��XC��@�HP����f^���J�O7@�<�\$�lk�OVI*�
�;R`W�V3��P'�Ӄ\��I�4ܤ�цF�z��J��=s��J��̩ch��WI -P.F�#���4�t%�!'����:��Zs*�!3ր|p0q�.s�� ��O��ë xPz��@m�?�9�F*m���c&�F�&z3�h���v.��c�t��@���ؖ��$���	PG�R�Y�4��� X�;��"�w&25�� �X�!�')ڕ�l�*;h9 Ο���Z�)��i��4?�|�#�M� ���jt�
m��X c��>�� *�D���F�24�d�s�������i���h�2�a���؞`�@��,L���iC��HOH��u+�mL�U$�d9����p����<�V��C�׆(��()gK���cA�D;�pqȒ��v����dh�=�B��3�x2$���(嫈��Ԕ��
�/���֐��*�I����lAT���z@�M�	�n��P�ߝ��A@�CQ/G<PJ����� ��ޅ'=�J�!�$;�Xi �8,O0�৕�6�\eK���^d�׾i�Jaf)i%8	�!\�n��u�Ua*nܭ��"A6Ʃ�]'^�,٦��B�
�=A�������ah<�� �x6� aBB�Q�����C�8�W�"-�Ku�[9e��y���y4�81�8U��KHZ缛��R� �yzwJUJXā�xX���sçs�q��G��F����.<q\y�4��twx��l�+H����O��Xg�W	�B����1���#��I�`L
3�bRj�~[��=�Vi�:/|�) �!�@���F0��Ɇ"!B h��F���"O�}�� HzԅB�6��,�2;O�����&ʐxc	M-��u�"� Ixց�~B'���[��[N�.X�1����'.�r�)�3�ޥ]U�%c�ʐ"~e�eb�۟O#�Q�e%���
!�G��v����~Z��L1M�&�I�J���iRJ�wbLq��_�_=
�P�k�'֦�k7�'
�0�ve��2Y���V�%8^-YRM��I��,Å��h�:�s�C�'��(�$�nӺ��Uݟ\5a]�pY���DB�m�Yw��fg�L�џ�Y��'I�X���Z�>1>�b`
 #J@p�u�ӿP����l!+�Q��'[V<��,O�m���8�➥�~��ɂ,=�@)1�R
hXz��0��Wx�IK-�}�чoGL��B XZ����w:���U��4� ae�!'P)R�`���_�_(���S?!Xtv���&�(���'L��!0��/4 ��)q�.�T$�J�h�Q�2�p�zW��JO��1��4,2��
�(u�88���	�1x�w��������"Eh��p��ֻt�M
p�<LOb����ZH����H�P�rA�C*ܹXRha�ud�M��(x��>�ҽ˥���_B����P�|E�sj]:�y2��~�X@�r��V8����Z�f�)E~�bBHŘ����a�X���H�o!:��P��*���u
K�W��8Aq�	�ƥ���,X���"5+�U|6�}Ӡ�vW�.�R��ą�k 6��/h�d\�T��05:n���
N�?Z��Kvpc�(,��Q Ĭo�zh؄'21=b��r*ϐ:V�¶m-����膷#��p�i�&x#�7�Z<ԛ�M�	~2�H2W�ߋa�vL�g��W�hJ��V@$;�ޭ�a �Gs\��`U�l�}�sJ	:��gU�\X��� �>�̅�a`�BxB�e���o���%�l�
8� @�?n���h�W21�� �D�U6=��O�����ƀX[�����<�F@�$���(�&��X��ɓi��Ha8t�`�ln����ߝ;�@T�4FC�
� ����P�ёsDG9[:쐊�A}��
�hG!�?����)I!�W�\/3�|jQ��Z>���x��Z#(�#M`���!W�Bi��fۓ�e�BI͊~�52uL�[c�1Q@��B�� {�9"ulUYf��*�(��|ӎ<3e��l�~YCA I=Ӟy�a�	2PU�(�v,׵�����O���2��e���PpD�l�6���d�*/���zS Յ (FL3�#��`�^���(2 ZQشhev\j�L�	0��!uF ?��H�!f6�#2��=�f��J�2J�q0!ϓ;JG^��ȗ,�`mBS��,�˴�>�f�BJW�5F�q q/�IAT���זD�<�K3#Tg``�CP`��HTqq�ø60F�'�� Ғ��uep�RR��.uT�g�!*��}H��S7`b
,����E�"���ϙq &MK�F��I3@iC�J�(K��y� S�cd�ӴC�2���ڟ`;�k�,��2g�2d�N�ұL[3���� .yDM����cK��)��b��e�H�ʁ웚7� �X���Z�~�:��01�"�!�ʏ�!G���%�-S�!K��V���22���<i%�25�6�qUʮ�dRu�97�t@��&Q� �����	K%P���#��5l%a2+�>k��lJ%�ig�Ÿ�AM�%C|���M�O���Ɇ@����iXã#bHXPYv,/h ��	0J�<iQ%Y����O�-A!%�3��5�'�TXԸ����S@X�vd�Z!镭Z��5:�z���46����J��њ�SA��?}��
_u$��fZ�@�:e$1Z��8��-\���`��&�f���J	!H�� ��2��9v[j\�d�n�(%�iB�ሠ���`kD��r�W�V��GZ�?�"���:*�x��O���4��.I��Q(P�4��q�$�JD��ʴ�_��`#�	Hu����d��L��M `�韰y�t'�LI����e�T�S�� 7�6�	TZ2y��\q�.��TSjs�Ag��?�̪�ԉPD��f��9cY'̴�q��'Cd �fN7.ܩ�%b�+�αP��i��i��ݚ]!Ĥj5�1o���@V�Wy��	�擸W������+rL����.n̆�#��˯;�@��-^	�n x����am����cO7y������t܈牮<�`�Gmߋ�`4X�=O���HTb�@@4쌅$_x|3��I�R���@HUf�TpDL� Wh\s��
��Y�ū�1�@�"��xPj�)ԋ$X�.�`,�(���G%�A��M��O�D��>zU`��럤X���Bcn,F)�2lS._F�p��-5�n�"��T+�>�����rE��
��-	N%���^D�p�D�5�$̩�B!K�̰Sf�� ����'�"�T���eW�Q+h."���N�?�CF�F�#��'g�a�ׄʷit�����%�~���f�|A�P� W�-*�]�𭗹=d�e���u��W-/)�I��M�=b�u�g�� ��(r���KP\	��?(�RE!P�ʣe"��TeU�2nT̓}��Nh�C������������95�daH�KI8�(ɸ"I`�S�����Đ��Q�:�OhbE �,�y���b�&X��@��ɖӕ� ^|ܓ���Xo�S&�4� #^�N�.��0
 5	t�8�^n��Q��iڅYM�h �Q���y��}�U$�C���'�$��]>��դ^�a酆] eD��t �q�� gT���`�2W�Le��mP]`�-v`՘N��'�^�@�ͫ�Zq@�G�V�Z��T�P���jQn��e�|���������Չw�([u�) @�;7��	M�3�0�a��ٮ:�	������
C�Ý2���za#�82����1�%�F< }v���Υi������W�E5���θQ�t�6K��<snI;�	����p����hO��f��gv��@�l[p���1H�fe����`���)�(���yV���eq��H��Zt���'1���Zw��!�%H4�xX�O�2��!i��I�%ڼ� &�B�3g-��ŏG35�f�zU�<*�����˃\�lss얫R۠��n8on��'`�\��F�ޔq��E����x�Zщڌ"��50�8'G���G�$"��ٛuL�*��Q��@�q}�i�l]�[�^��Bl?q���0��k��T�g٦nʆ�Sj�
4�����	ϴ-y�Y�6�Y�s���(�n�n��`�'ؤk��7��.Dldq�vE�]�Δ��%߲I�*�j��V�mSr�����mR�	�t�S�<���^����߳L�8�"t�@�o8�a�a��80Db\*d�H@c@�F����n�S��G���Y���k1�M�?�Rm�4�ݪd�	&x�E��d	�7B�h� O�K�d�ag؇xF��5��Ҥ!��y�q��@�h�3;����Adٸ���haC^�	�C(�+A���>���G�f��b㣄](haBd ��%)���� �*��L�b	�@)�wE`�5&�eȢ?�x��U�\�h�!Q ^/G&��o��>�S��̾&:�x�
��d��2���PQ�.���l�%���O������yÔ�`7��5�Т��g�$iQ)�rhJ|8S�A�hSl)��M��$��F�0�ز��W�`�8Y�B�qo��/McO`h�wω
t�T�!o
)��i6d��e�EƦY���)��iV$4z�����g������a��8#�F5=
X{ �߆a8n "_~����)0rOB�;���$��;11O������r�Nȃ-
�+)v���a��k��H����8֮p��W�	X����Av�^�˃-��,&d�Ҁ��)�u��O��I��_�+rʈX�
 W���	񢀙S�ٓb��H�P�����#1�,��%�1EA�7f�h�fg	?3��L�e4yCfJ'h}��{���wĀr� ៮l�F�I�6�aP'�(f iS�������`�%d�bb&_(i���0k�%�
�LYC�շz���e��Y �p�6�rOߏ_Ůaq���B�ԄJ��:.T��LZ�~:�������8���0ʧf��ć9GxJ��&I:;�(B��GAh�3�g�m�����j�m�@4��EyH��FI�8=�65λ:o(!���߈F�#����������RRy�΄T�H�����'%�}Y#�L'!��M��ǌ� (Ieg�	f����bjX�)~��!�BRuX�pf���,��y�rg�<(	��H?E�5t���!
?V�H�K.p2x��a#ל+������Z���&ӧ]�f��A+���,
�/��w�ī�`�5:\���a��I8�}��a3f�i2z<�'���U M[�	$�z%aґ�����K�.�ɲS.=�an��''��$�S �p5A%rݽ���	�4�t@8]��zQ��Q7�ͻc�NS<�{����r��=NoDH��̋'P"��AŐ�Z��t��j˾h��e��:@��E�HcPh���'
Z4 �3�ē�y��]�R\�z���&d��`/D�0?�'�)9�䠂�e����$ֽr8T�3�(2��I�fJŹ;ÜI[��´<�؉2��_l�B����q&<P�g}R�7>�dLJ���(ت�Ω�O�Qۦ�ҎL�z�P���Y���!U���t4f�0��
b�[��$���ǃae����ѪV+R ᅈJ��N8��(��Z�2��(�!�4���BۦA���ak����Op丄� o�bQx���|��$(��!�>�;T"Ƈn�Q�G���~�C��C&��.�� � ȁQjڨ�a J�a��	A�4@ef��
�4j�FT�A ��8�`ɃUbʴ�;I��%����s`f��ǈ��Mx��I�XY�u�	�2K��;b��� d�'mE]�	��
�!|����G�~ڈ�I�e�1M��#B�&��O�`�§�6(���(��=.䁃��?&��iQ�L�BR@Ѥ��@��k�pT�q�#'�'j�~�SF�Τy�D�E߆<xDI�&��:aS��	2H��7�uJ����;,�V˓5�%S��i�ҧ��i꼄%��v؊22-��%�¸����`*��q$��" ��}��	�f��݈�o��v���C����x���Th !��ǎ{���4���?I�6�4��S��7=F�u�Z�m,I��"O� �ׅ@�c�޽{��\� ]ab�'_&�ܹCE��hPU?E��ń.B��Ud[8N{�h��$|�!򤘨����&o�1]��ѳ��E����y�����N.�$�0*�Q�� �,C�j�0�ܔa�/�K)�l�B�'h�d���YT!(5�� GD��(����8�@�*�rm�*i�DՀ�B����	�@��ȨO4���*��-�Q����=Bx��b��!�责����y"ʘ��\U���]8�Hx�T
�:��䛗v�4�+�{��	ӏ.��:�k�KV$��E�v�!�2 .��VKHNL�B�@�=�!�d_�a��5J4 �F8����
!���g8��#��3I< �B!���y�x!�&	->�P�Fn��t�!���e�r�Y�k�2���C�LΦO�!�$�E{��
'�L7w��5P����!�_'At�z�AY�'u h�k98�!��>2K�����	�uyt����E�3�!�$ȶB�"���G�%^qpq���ؾ�!��C�+Rm���վe��U�؋2�!��:F9��D'�����RE�!�dZ�e3z�IS�2̠�kX��!���s�>�A��� }N�G�̑\�!�R>ql`��$c��PC�w!��.�l�OJmD|ِ�R0Qm!�	*���1����y�a�
e�!��m�ִ�DAv<��#��ES�!�D�,[$�C�hքI0�d
�.�*9�!��	Z��B%(80-�&���!� Rz��a�ƴp �]a��	
�!�#��{�(
)s�<����K�!򄐄�ʍ`��'t�.��/	6�!�x�����Y�_z��M� �!�dU�`P4,PbƟ%%`�A�mQ3i�!�d�?�Y�D�ҠBFp@�@���!��ï<�&-BmÌT�������!��:5�F ��	H�~_�a��	A�~;!���`�%B�&�`k|���"j!�D��A�@��IS0Y���J!�dʴ����CI�_� ��BT!��%	�`O�tǢ��rm�
U!�DG�N�P�k7�X$L����1���H!�ď.5��:"��E�ұp��P
9n!�DP^�Ɓ9Al�F���ib��]!�Dש?��@?cL:�!�!�D��jH��g˶'�����8[�!�d;L�9P�ƺl%v�Ȣ�Wli!�$�$)��\8�n�P=���D�+{b!�DϥISCt����%"�WT!�DڛR������F>,p�ꐁ��m!� �X�i�{Zd���G
`j!�D�n� Ke+X�@b�-E��� C!���2"��-E�F��r`.�6NI!�
�V>�",փ|4�	����.'!�dS�o��e���D�(7o�.1-!��+y�,�����n�`8qE�����7�$
��S n�d0a��9uCM�(�0@Z��� ���3��04���2�`�A���^:r��if��"+�������3�!�g\$��>�}���ѿ�v�q��/��ic��W_�'M���M�����!M��'K|�Ӻ"�,b���(����7��޸�K�!�� WSd�R��L<�S.Y�r�8;�βO���!�K
�`8W�A3R� ��雞q����cnF�O�i��
'r������[��I#O� n��l�Q�b�����I�,��7� /̊�d/�|���2�� x��ВM����w�?�׾]�!a i��?����T�\���h���h�7}��G�����GͫH���Y��ܙ��c�vH�u*�}���g�]�Q�X�֎�[�&D��k�s�ر��;a�rL%?�B�&L#V A�ǗaܨQ
��#ʓ![0�z&M!R(<	���dֺq:��C�?���(^� �e�T��0̦�Qd_��
Q`������#O�� �u:A�,��/6׬ijP��e��|�SBF�!���B#-�$�h	/zk*�A��~mv��F��̯4�� B��E�Ɔ�R\���V�k}�'Z�vX�0	�$O�h��vP'��IH��&?]̙�P%FI�S�B�z!��Ẅm*U��8��`ytjK���S�%i�8<W���J�&<��ˇ�9V����/��"���I*ӧ[�z�+O�j��	)N�d����]�%�,E�UkF�<����k�^�TlQ��� N���)J�������'�����BU�l�����q���ķ?����
�T P��;/�l[rF[��1hV��F����Y��r�@Y�JΊ�р����׬u	��;X��t+*�y᠁�W�h��u)O5��Q � �0�w�}��m�)`M lcpD�0����)t�I�Q}J�rRҖ�~}��\�C@��@��"_0M��Vn��=3T�)���/�&�CfH��$��Ӂ@v��Ϟ�D
<U��ع �	�ܒv���q�@��?�! �s�9��>°�%R�QǠ��,r�|k�#�L�
�u�-����5"K6a��bH$�M��N��`]�і�%+\����
M-�� �Q g��U��Ҹ"&N���"�O	Z��'J;6�{�?��=L�xL
W�D	��Q��Ӫ!k�᧩Y7hh��*���*:��f�}��a��F,%� �P�S� m���ٷik��*�h$P�#kD�((�^�pH�e�c,@�8�R���Oy������
�ʋ
:&�G��i[�Љ�B�֥Ђ뗥|8:r��E�uB�O\�*�jm�wC�#&��<T�P%@�ڡ�BkV'~?*��@�B�]�9��+g�E`�p�ْ	�:�љ3j�p�Vx9ȗ�/�&찃I����'�.��i�=�ݣ���E�T��%��8x��e��n N�Do��=\�(� $T�M�&�'�@��Ce0l��E�?�����+I�nx��`�n����W�h뾹��/�)��vJR�h��f�Z�M�x\��Zh��)Ie�V;m�M*�H�V��Ͱ�T����I�b�'w�$h��ks@�)�'rY2�X?�xfN��U�\"~���ĞF�D�2e��o#v�,j]��-��J��U*End��Ǭ8W���b΢S"L�
�@�0h��[wwF����1���`)-/�`R)��|��l8�+�N��9|��d0�[���ÉեP��%҃G[*	n��Ƌ�F\jٱ�̕&=y���� ��g�`"T�-�B]�3G�(p��Q&�%CPr���'�@�8�R�O��#P�:e�􀠴0��J��ӉP%t��%�B\3hpVd��HE<�.����bn���dU�5��P(6�C�7�Hx&��?CN#3��bq:���1f�)jؘBH.���"�S�A W���x�*��p�<n$p/� @D���Hu���NC+uB����(jK�{�Z�(S9d^�Q�3.ǐP@�bF�x��I6�iyRAA�|4��W�����Ɯc�Z���bUW}�)�#��:W~�F�T*'Ny��]�?EK֝+=�43GjO�(��s�P�'y���b#N�w��=�#�p�|� %��]�Iu�2fU��	X�����
�P�]5\$8���fŎyLx��.����m�Eb)xg\��G���Y���+�4_.,��W�%�d�2?�v�	��-B�
���N�X����je��X��0*1�W�xv�IǍͭT�����A77"a���ĩ!�q�����@_hKC����F�"���8�:��ã�h1�t{5rj4�V 0h�bV,E��U)���,E���*4�E$j�Bi���`�:��Z,Be�`X$B�<-�yX�,�;�`e0".�{��ɅƓ�В�G#zxf�:g�U.[�j��0���H�5��ǖ�v�J��)�:�
܊�'�#x}h�r��Ԭ_�d�ϻ3w*ћ"nA�a&�P�f�%s�Pه���r�\�{��wP�Ԯ4�~x�MK*��% �Ϝ2���)���F߶�����!��])���p� �I!�\�	�&[�c�$a����=��"ȰUw��vIX�H��|ͺS�B�#��1������m��"O�ݪ��V�iҏ�3�:�c4O"�x% �$�1 ��:C�պ�FBW��~�'��?0���adG�T� ��+���'�|��5";�3��ȘhY���ɚy0�5��@_������ڏ0V��HRjH�����x2�9��0O������i�����b�j�L�W�Co�e��ϩ�0>1�h�4~R6�A֥��$^�����;5��Qf�ÙfX�`���-X���dW��Lˢ���B����<}�D#U�T��
#%�P�B4�*�N�5C�2���#)ϋR���R�I�x6��"�
�&'z�#*�S���GC[+3���XBǮ2�J}�'�O�>ɂb�P5x/F��2K������ʦ<	��K�Jw�9�K(���{�߉�Բćߡ+&���1+
�B����E�>���qì�$Q��E���=|S��Nd#(���/�G���g�Y���΃�#o���%F'eeؕ!߸
�(�kR�NXO`@:&�X����C:"l���u�F�a]�Ea8B�F��	2:h��n٦2�p�-�ifJ��7�'},��ΘH�@�)5�l���R.����7	�Y!s�w0��r�_�
G�p��	Q�6�n��W��<�@D�.$��q�4)	�`jD�g�={u�#?&/��MC1;��ĻE����S�V�f�&���T�+Q�0B�D;���afSM:D��2EJ%�Z��P:g���i`�X�R H(�(z�L3�vDžC�f��Ġ��x�M+yFV�	�I	��ێq����=E�|������0G��{@D�{4�>Y�
M�f�W,c
ra�� o1����M�%kX�XR�u��Hڎc�h�3�b�-|4Е��0���Rf�<}р���*p��h��,b;Ȥ��Gьx=Ĺ�A��5���RV�͛9r ���#\�M���j���/ X2�$Iq�m��O�S���!�|�o��R����q���aM���G�I����Fs4��tf� 5��<qb��+@3ft�1��Ofxj�!
��B�C�Ԓ��'0<��$&��N!ґ�
sv� �5����S�I�����ZPz����K2����Q��ru�0�E�V�u��I���xa�g� �H� E�Օ.�����LG�z&T(p�U�L}��ʮ^�|�ɗ��%�\�P�M�(��ĺ5�,D4X�4RS6� ��+���E%R��n�`E���q�<@��K:[Y>	��-�L�Pe�	T��ڲ�ٚ��K!]��?)B U��9^�� GQ/���R�i��e7�
��8<ڢ��}~.D6,�m@ĥK� �� S��Ύ��
�B�ˋ�f@���p'�	�NP�@�B��9�X}f ����z�k�gB�!*��1V�>�b�F }�d�J��#HTC�C_~�*�D��J��;Yt�X0/�V�d 9� H+>��Q ���u��3�8��㕝R�4�����_�J0{P��:=F�y5+��0�,���C�O"8+�A�u�(9⺦�XSD�G
Qώyk�i?@�����̶C�n���f�L
��A!��BS-�=,J{� 1�V1��+ٯn�z�ʾ*� 1[�ԁ.��њQ��2�����P��L�I�g��2��K<.��� ��W��d��Yb��am&�H��P�yr*�9Ư%F�(�bF�Cbd���4=�����h�[��\8�,L�u���:���q\�,a���hx�\�2�ɪ7X�a�U��)R�J�&��'I���� ��L�#؎j	��3t�Z�n�2lJ1�8��� �z�D�4%>z,��� 5t�Pa�@���H#6mk�C矐��H�HXh#M��M9�	�F�L Q� �L����h��<"�ő6����W�:�L���[9QJ ����d���r���+0�uC��5�
�@�/���Rc�v��lHs]�А�kBW5�X9���6���8u����(t!�C�%bt�;�o��W���P��Q>�x�f�?�(5)��2<�f�H�jbN@-hq@��tdFqi��/'� ����ևu��E��̣^�B�0!P��4 ����1B��$څl�5���_V<=c���\�J��0У�*$�U���F��4��ׅU�Հ�ꝡ���k��4xY��	�>���a�[FX�B�za��xF�r�tD�d�D-�9�W�Ka�R�I�톄ML�xg��8�ʅw�dX�$�d�$@'�&tE���h�&l �(%�C�Z<x�'�(l2%gG8k�6L`$(D @xl�U��(]SF0a�'�;f�H�;3�O�Y����%eDgz2�K6�>0���u;�@8q�G;d�B�c-��X��Yh���{�0�u��q�@ ���&H���G�2]!��)�N��{��p8B��/}� �E��p�D����'~H���K�7L�d!H� �������B�O6}�4.ւU��d_�?+������B�`K ���O�`����C��2�ER�R���R�	J⤬cd
)3Z(a(���+M�h�\w��N (1_.q �M͡(M�t贎��[��8zte��
�������OD��5��"ER��0�
8�BL2�$�	ژ'�FD*�DT�[�vq!͆z4�pA�k��� 2#W1�P���H�q�F�`�I#5x��~>�P97�����x�AԾ��1��PB����v�i������'��<Z�@K+C䴢��L�O�@���KO"AaHLѡI�5y���#B�?��#d�E���Y�Q�ʼ�倁E�1�O�¯��	�ӖHVNm� M� a=�r&BO'��`'��RFB�%��T㴅U׮(VÐ.b(�T
�΍6��oM'E��Ӈ�ߕG�Ȩ�d+�)l��\D,�;z��Ua���K�T���Ox����!Qn@A���u�]!� *[�B�;
�X�2�#�җf��
���m�5mR<�2}�@Oj�	�&|�e��l�s�=���a����dA�?�� ׯZ1EP@��)G�AC�	v��ۈ�DO�����E�<D-�v �������/(S���d��o �R1�������e<F��@�~Z�	*8��9K�LH#"�z���mȺ~�����2%�� qĝ6٢-�/R<S}�\���+-�\���c#bǨm8�n�d��Křk3Zr�LU��'^)�P��B�0c�2�b���k��H�0(>��X��_퀌��{G�tEJac%�څC���ť^}��*w�7TG�]���/O��<Q�BJ�8{���&莤m�>ي4KJA'�X���.n��p��N�.M��0y�B�=v�Ȣ��&h�V�8_������w�zp,�
I�4���͍=�$JGA��� ��\���F	���`T�a�Bdzׄ�_���K�k<E�� S��W30h��H8 ����0s'���c$Zɂ�b��sM\� 3r�ıd.��kWH��A�T�E	D4C0'ɟL��E�JP[t��|��ٴ�'Y�I"Wc�����%z&��	��\�f@-,tԠq�$K�1b��5�X.6��� �zh�jޗ.���@AB�%bhk
ߔ���G��d��O_�! ��P�O-ZRt$n�D]��%n�r��6�']dX�3�<���D�z�Y!�I6}��и4)�0��UQ��i$�1Ѧϓ�����b��g�6H����@J����&�a��C�C��Z�!����<�"Ze�2Dف�,CF����JӦE�'Ǹ0�F���G�@ g�O&Epd�SOE�C|6�Ղ���لȎ�th�H�HB,	X1Ƞ�OJ����W�4����Fo�
h��1�拚VGz�x���h�\�����Xm��!�dW6�1O����W
	�60x)Y�~x��g��9��X�p+'��Š���8p؍ȣI͕�&0�)��lXȓ��
�u�O2�T�H%M}�iV���<��ed����'�S�$@1O=XB��!K�y@U�N0Hr1��уa<`����h�L��TE�
ZRt�8��B���&i�/K^䰐u��
�+��j�BՂ�Ŏ�XUz��CF;{�2�@�AJ�C�N5�r$��6"��PD	���%D恙�	žE�Z��pET!]��`��ٟ�c	'!�p��)E�P�ް1��� vdz@�����R�Ҭ	��ց"u`��(���Fn�>��ٚo�&:�d�;Q�_�k�~츳J��t��jG8��=��.G�:��ݒd�'>�|�C�?�P�2�m����F�0d�ӭ��,"�I#Ø�rp�v�<(6��.RR���S8Xfh�U�Wd_�0�$D�;X{0��fV [�d�y��KMCp����^kr!��햝f[�d�-?�n�2"h�3���B�&Y�p�e�F�"��0�{R��C��!��ٗ_�R ���P2bD	�!��R4aՌ_T�H�l�M�DO<Y�2��A��D��[���AT�Z_�'�"�2@۔UP�C�J�,�ްR�'6�YaEAD�BúH����)@�2� c[�u�oѲ+Q��ꐽM�(�2�ԩR���3�[&7�P+P.�.�L���I7�6<x3�`�+�G[�}:���	�T��ظZ	h�% ۦ#yƜ�0�̆������F�]�Mj�w��/M�e��� ��o��Q���4Ȱ�;=�,�6b�N�f��Ǒ�I�r ���!h)B9���G+yy�dhǂ;�:4�F�հM�n��7��	�sd�BG�0�$�MӨ��#>�@.�_�DrV`��@P�}2�#���R0��:h� h�j��o`5J� �������	΍:ե��@���R��.�>��:gM����nRP��1Ʈ�<y��H��4�P%)�b�����_z�$��N�-3wΙ:��!.�@Ő����� M��`����e�N�D�'/n�C�
8���`�-1��#)f�S��O��@c�/4�XHRp�W>QZ����I�73��Rc	��yg�B6���,�����3��+�p?qѪ��;2<X��C?&��/G�s�(����w�`�T<&�hjwg�9k�!`׫/B=$����һ���psg���(�	�f��Gؑ���T$�9��u`�锃D�̡!h��&�z�s� ��D5XD蜚���)r˖�1W(k�?��԰�aι�h\��jX�*�Z!Ppm�<�QA�*`��t{�`!}���psՀ�7m?zA��10�*A��J�� ��͂-|��0c�`k����e�5!"IB�] +�$t3��<��[��cD��>+3��X�II�!�
T���F��� t�RB��I���uC��S�"O�aqE�ԑC!BիS��:)�]8��'�H	d"U�>}���[E?E�D/�w��\����T(]ф���!���f�4�:�$Y T�����m��e��$ˤ��.VuAJ}#-�Q�Ę�*Ǉx<�h�ɜD�¤�(5�OPyIԊ�=V<��I��ZD�cU���n�VLFI>�&����Qt2xB�CH�Q�����l�[�Q�deGC�E=�L��C��A�a�w��X
�^�!�$�5�`Bf���SsPePp)6t���	~ J�I����Q�5�� F9?��Ի�cN�x�C䉛}��h�t!ڟ�n!Qk�+z�lC�	<Pۆ�H�	B�hr\�脏��C�	?
��=RP�C�E��8�A��&#U�C�Ʌ �ʄ��O��Bc�l0U��R��C�	.��P��KV ^�<����dS2B�	�?1j�b�U�\@N��f���B䉜	?�;ug�,~ Ar���noB�	:]�>��!J˫�� ��Y/4��C� {q^���J$F��)
���R��C�>o����E��e�,ʢ&��f� C�	�>	�0�o�M�&�!I*�B�	4+����_��hm�S͜+0��B�	-�`��+V	u},��cC_�l�B䉐1�x� ��_�Q���O��?��C�	6��պ�i�>o����힩�C�	540X���Q�td��A��� B�ɐ?E
���gG06Vv�g+J�����Qp���W�A��J�e�J�!���z�2��#��>4El��2�l�!�W�oIp����͏=;4�I��ף,�!��z/�5a�L3�� �1~�!�߮�2�@f��2@�9Y``_��!��4���[��_|0lZ�aĽM�!��P�v�t�[�g��S�6���5a~2�<�����&�dD�G�clN��-[���'&v�ㆍ��xD4�~BńGj�%�h�=�l��}�䑰2z�1�#�W�)���.�Q`L6L 9����P���b�e�Y���S�O�Je�u��)v<��sl0��h�r�]��ɘr��_�)�)�1m��³ݟ��D�'����6F�5�½�4�]�J�:4x"�O�nb�Y��4W����I�or%�s�بy�m��N�+6=����8ƈ���O\��	�'q4L������ Y�k�ft� g�;+��ɰY�$�#���Z��MC�{2f·!ߔ��D��/��D�1r<�̇��0|�F*Ug�� \+H��}��Jr�dP8V����!�U�)��PIpx1�(��\�n(��Mٚ+���ɩE ��zec�u�)�'�^<6ȅ�8����B�T�g�4q�ͅa�^��Þ|��)McL��i5�Z�R�F�t�ۈ>�`8��
_�?a�4��|f�I3���@��1w�L5A�1O��9g�,�)����t]X�>PrIQ�ن��}��$���)ۈ:��[�J2L0��F�C���.QQ�"}�ׅ��(w�ܺ��t�\܂#$�t�<!�EvW�|C�GE�h���p�<����$}�-��E��"��pC�B�<�c�Ӱ!� ����g�1���
d�<�c��bi�x3g�^�M$RYPQnUa�<a&�P�y+r�Q@N�l�Tp�G�[�<�Fŧ_C&(�Zt��(hማs�<9��� �(�3�lG�E2$��u�<qfo�&'�f!Ѣ�f"ޝ{p	�p�<��gԸ]�A�GIp�����́n�<�$Ͱ��Җ��.r���cOo�<�qI� ]�}Z��*p������m�<!����+�,�#��ӠT̎a{7_A�<1uÚ!b�Ҕ��,Ƞ%\�t��<1`��1_�tT��w�6�zEh�C�<� �0�T%B&V�>@�E�!Y�  ��"O�9@��[a9�eI#�vx����"Oz�0@f��PI�t@F�VZ��(�"O�r2�02�M1��[�9K��U"ON���)Ԓ`g�K��[���"T"O��X1��m�P�Å 3s�)V"O8����X=}G/�A2B�#�"OP��3�L3Ik� ��G�#n�Q�"O�dK�$XLz2� 4�Вn��4��"O���G��h4w�Q8%:`�R�"Ov���cՊ,9�M�g$P$�.x��"O����B�a���Bڶq�"m�c"O�*2GۂW�LZB灁�����"O��e��-Z�:1�%�!v�|11S"Opq�0nO� xy�&#A���50B"O@T��O��wa�� (�%ht��a�"O�,"�5S��M�q��I�0yu"O2���HB�(��s���7G���"OI�Dרi>ҍ����>/�M��"Oh��qúQ>u�(��4!���"ON��@䊯ㄸ�"(�F�[�"O�5����l���Qǋ�O�(�"O�Ց#��I�.ȡ�
��4�B�"O�!+"���p�9�C"��F��a�"OFIK2��0~j��C�/wj����"O�)�L��:�S�4�8�"O���b�^���q��ߢh�d��"O�B�XM
�m��bņ>�X�0v"OJ�q��K�X��b��T�����"O��J�ƕ�$�i����r=
�"OZ Y��R�!b��dA�(�؄�S"OdM�S��\�l�:��I�tr� �"O�1H�ϞF�x�z5

�#�(��D"O^D���I�1a�u	�,�D]�A"O�e�_$q���2�́cO0�"O:��Y�58�C/Y��s�"O��Yr��4J�,)J�J�~>��c�"O֠s��U�X��=�焕1 1VEK�"O`�1Pc�	К��`�Q X�A"OM��5ZȆT�!�G�~R�`"O�dh�/Q�<�J���J�)��(��"Oٸ���'f/� �kW3Z�ċa"Om;au��y-i����5��(�y2�I(uޘ��̟7����*�y��O��`�ᖭ��-ǚ��g�$�y�F�?S�u�G��1%�
�ɖA�;�yb!��WD�)N�������y�Ŏ4\�<2!g��b��yR�&k��X��a���xK���yr�'%�*��P��t�>ْ���y"�5
�H`"'a��i�NXq��M#�y�!J�7G ���&�#p/>I�1�
�y���n��1&�=h��43`����y�-A��$�͎sN:���O��y�I�H	��f�R�9��A�� V��yB���(�<<�G�.9��������yR��)/�*8�|�v���g=�y� �l��t!���l��m��+�'op�C��đ:�p�@�*fl��'��DaS:)�N�`G�xɚ��'�4	�֍͏ �Ԕhv
�\��Xp
�'�P�sPlE�0ph`RB�E��@j	�'��H�v�AbP=�F�³4�H��'���JRn�
4!-�(h���� 4�����hP3��D90#0"O��㗎�:i["��)�]
hx�s"O2h����X����Џ��9�|��a"ObAc ��E�(J �ݽ�10"Oҙ�B�,�ͻ���"����E"O&�rL �+�(���A8
��8�d"O����j�L���� �
�H�"O�Y� L��-x��jClj�*E"ONI�-@~��(�j��\�,!�"O�Y0wM�E���J��d�N���"O( 1�n�*�`+�)_!Ғ��"O���"X-~A��[��4�C"OR� ����&�
爌�o�����"Op�p`(.P ��ƍ�x�� e"O� ��Eh�6]�K�Êm;�"O�h��,7���a�+�41��"O�5ZR��zg�u���8��,�`"O<�s��\�P����ש^ i�"O�I+�B1�.�I%�ԏ&�vYQ�"O��CR��Y���csh
r�����"O:xj�bڃy���S�]8�����"O�����LM@�%��󨤰�"O*�ʄ��Rs����$��I�\�&"O��y�j�lq�@���A���qc�"O $a- ���"�D�f"OJ]���K�R�d�0�- �&y�q"O�0����)/�`��b�[�� 3�"O6�PʛqhfaQ&�B6?��պ�"O���!��<~�a��H��pQ�"OF�r@���`Kj�8�*S�]7�<@"O"y�a,��g�"L�I��
$x�B�"O�� ����:u�i��\�?�ˠ"OҸ��dԑ Aʠb�#�<{����"O���W
�	�4:�!�*K��QU"O����.!jD5ϐ�n��b�"O4����<�ir���&�2�"O�9�"�S�*� %�a��# ��"OL�(��_/BH����&��2�"O���S����Z���L��a���"O �Sf �N�`PC�)��"O����ܫ�z59��Rl��j"O�h��F�1��Ѡ���p��x"O��[A��\��L�U�D��"O�1�a�BG^�(1�-b<�ШP"ON!��ꅾg}v@�F�+T8*�"O��+҈�L�<���Q�}��8�"OP��C�	�rKvyYBe�^���b "OHc�$زi.����DC���Ȅ"O@)�r%G3��$�c�h��6"O ���Iˀu��8Ձ��k�$�@"O�p�V�d�� �`!���'"OL����F0r��=[�%x3&��"O�͢5*/<Ԣ�@��Ëv1����"O�M��@�^��,U��=r�1��"O@4zW�L���Y���x�8�P"O�lJFƗD�<���H=Am���"Ol(�3��q� � A�X����!*O���F���"�:o.��2�'����`�(�B�HO>a��5P�'�b� �b�d$i�/�5)b0���'��	j��Y�j�r�����!�T�)��U P?b�J�d���Pz�(�,!D�tB)ܯt���zq�*%���?D��Ɉ�,����$e�F��TK=D�� `4`�f2��+�ǖ�)�z�P�"OREA�+@1AFv���F�;��*q"OtYx�L�+d|�� c�yf�SD"O��D�@+P�q
��5O$�R"OT��p��9o|�`Q���GG�`��"O^��jD�O�^����W q���"O��H��g]D�A�4��dp"O�`����>,�΍�-@4C���[�"O]��݇&��b��U�~�@�"O����ýF�Dt ���6,�#"O��RW�۴��y&�e߰#�"O���
�6p�eyS$�U���"O�b�ML"x� �����Y#�"ON�8R*î�Hl��ӓa���)A"Oܰ�ԅ�
k�	���J:�A*"O��p��xN�9�¶_ &�H!"O���'�����!@��	�"Ob	��U�m/J��w��9P�-�Q"O �ؑ
@*U"jER��4�"��"Of,��ã {�ARAʂ���l��"O�����R�����"j,A�"O�İ�/�
6�.%�s�ʬ(���CW"O`�-�K#�������W_�I�'�N�����&lACI�RF��s
�'�2@v�Ʋc��4�4GݯQK�T�	�'I�YI���CS�@�s�
8r՘�
�'3F(�Ӆ�-9 (����d����'�TQT.D�;��W��B	ԭu�<�`,V�Ac��2�!N�b�ݚA�[�<��O�OrJI��KQ5T,0� �W�<���!b��� A&�qfKQ�<y��ѤO�����G�7�|U��+�P�<Y1���`ݚu��'��(a�N�E�<�eGɽm+~PҀ�Q���JE�<Yp�ĵL�Xx���!���s�˂A�<�SMB�^T�y�S�O\��-� �z�<��H�ň-�c��5!�D�bp$�u�<Y���0�IF��5H�*q��q�<��
T:<j�E�/%y��p�ko�<�1���V�tx��@��dLFk�v�<1w�� 8R�"v	V*Mo%a�+�z�<�5���d�`\q�_%J�b�x���b�<�3�x��JblŶK�Nͻ��D�<�e�ƛ8��P�,54�Р�-�v�<�3'F�hʈ�}p�I��JW�<IUA�?m/ �s��߆��0�ɆM�<��*�d���t/J�B��0f��K�<��E��H�dW��� ��,E�<1��S̰<��\������K�<Q�-Л;a�p�0WsH���N�<i�o��Ǟ��A�[VG̀�w�U�<����~��&O	���k���w�<�ԣX��b�@F���Vc�̣�F{�<�~�LB1 �^�T-���Xv�<�*@&�JQZ3I�
Ѡ={�c^�<��R�p5,Y��f��`�~��J[�<q�bO>&�`pҲ��6s�2�S �U�<��Ή��:��m\�S]����LN�<!�HN���Ł%0a��:���U�<�E��/;����"do�l��cU�<���!$65ɑ�M��z�p��M�<��j�"#����-�G�,��5��K�<Yaf�u�态D�`�(��S.E�<yD _; 8  ��     �  d  �  �+  �6  oB  �M  �W  !`  �k  ]v  �|  �  [�  ��  ݕ   �  c�  ��  �  2�  ��  ��  �  ]�  ��  ��  ��  ��  ��  ��  � �  ! �/ �9 L@ �F �L #N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7����l�ƀ�M�hX6�	W�~����qܴ�����'���#qd@c��U'K��D!l�r�'hjeyV�i��I�|j��OP�'jE���JU%n�(ڕnկc\��<����7ڧ}��僐�S*	(����+��K F8ږ�i��M@�y������.v ڰ��ě+��x��Ɠ�Q���	��������C� �V6mm����B�#F�����n�=|k�o�ΓM���q�����'��Rd��dR��k��<+�e��'@�	R�	�M�S̓��a(��PQ�tj��_���`��ͬ>)��?��'d�I�U�0D���Ћ)X��	I"�b�?�0*�D���|� 
�O��`��,&D��R�7y����b��;�t�*O���?E��'�tS3��f���IqXR�l��'��6-H�x(�Ƀ�M���O�`#cK�!T′���0J�:I��'���'Mb@��<9�v���'O���L+\��9��L�6g��YTF%>��&�ؕ���'�r�'���'Ǧi�1'�&�ᛱ��$<?0pQ�_�0ߴI�������?�����<9�b��{�U2A�V�GA�#�{���)�M{p�i�vO����F�iOqn�4�$�K�i��͙a��T"��7�_3DA<ʓC8�x7��O,�J>Y/O�,9� ̩S�
' B�'��`��'0H7m�6+���R�'nĨ��7L��C왈7'�D��?�S���ߴG$�F�sӨ�q𡇇Z������!]�h��FD-CGv7mg�(�ɻ���A�O�pŖ'��d�m����\,f����6��?�PCz����Ɵ|�������៨%?��Ɂ��p����r��a�9d���	֟��	2�?)F�}>i�I�'�$�D)�*4���=�Z�A����M��S���435���O֚�Q��i��d�O `7�H�:XJc��u�Ls��/E%�9 ��;��O���|����?���ޠ����V7�.��K�%?�� ��af���+O��o?i�����ܟ �I�?�]8c@p=yЏ	DF���FS�&�ӟ �'�"�iA6-�@��?�V�M�����CD1%�@4
蔎nXx��D�9#B���+�Oz�"N>��"� ��H���F��N��N"�?���?���?�|�(O,�l�"�~豱��'�8��`dC�tg�H�^y$rӐ��ҨOd�o�%e��PpCLZ�k6�4-֖�q޴m�%H�hj�&9On�Cv�4�韚E()Oh��a�Bo W�B�,$rPK25O�ʓ�?���?����?�����z˼2U��$j�y�0O$eN��m��,�I�I����	[�s�H����0(ً[�ƀHB���f�87�Y�`��vtӚ\&���?����@TNm��<�3�]�CJ8!!��^�[��] "m��<y���SH��������O���@�?�̙Be5c4��;t���v"|�$�OR���O�˓(j�B�����'2rȆ'������ڰ��2�$��|�>	"�i��7��A�I�r�Z��6�I!`���ENt��	�� ��@)'3���FEy��O����	9T�H_��x;�n{��������y�lU�l�ʈ)��qE���(�"�o�p|(3.�<��i��O���
�����Y-��z%"�AU�DVЦ�ڴB��&��1?��2O���ۮy �Ai�������'�;�Ä��*@%���I��䓫��O��D�O���O��W-,y 
��z��oޏ"���vI��/���:��'���O��90�'����x�h0go�5�����)�	,��-�Mkǵi��7m[\��?q��-@��h���JK���ԸƸA�"NԔhW��u#`y�E�O�\CH>�+O��[�������#hS>��,���'��6m�9���D�"&��H�D��["�i���<5b�d��=�?��R����4Z���fb��ĺ��#! p���B��)he��}��6Mt�D�	%� ���OB0�'��Tv�� 8lRb�	�x��&̒"g��*�3O��$��B[H��	�1�(!��e�%��d�O���WĦM��M#�u�i��'���Ǘs�x;�d�|aV�� =�EȦ�H�4��s��.�M#�'b@�_�4��sd}�6]��BY�E� ��'	C���ן|2Y���	���I��2kх*&,S�J�H~�(bp��ޟ��	`y��b��u���O�$�O �'Q��M�V���d�ꀠNO����'����&,tӢ�$��S�?�Y�"� �%����9+_(<C����5�Փ��ۉ[�,��'J�D�^o%�����8�'��U�#(�<}���j�Jo��,Q�'���'���o4�$�'���'����9STb�.)dM fTB�����G��&����O��4�d��O\�C�O�%mZ)k\<��vf�9$8М�P�ӓD� Ȑ޴<؛&D�(o��1O
X��)���A����T�OpM/o.��:��֒D�ԵIb���mKdR� �	ڟ8�����I�,�O���,�-q�
�qA+U�z'
 Kw*r�@��7.�O`�d�O�������p[�!I� 9&R�Z^-+;��!ߴ
��v .��IX?�>6�i�L�'�_s����̟�?G�pCcv�n��L���'Y�%�H�'ar�'��S�D�e�go�17#���'i��'�V�$�40Pj����?1�k����k�D�� /[�;b!��r�>һii6�@|�I7*� u����`��50D�q�N�ןD���	�����gy��O�,��	=��(B6�z�X�+��u5�1��5�R�'���'�b�����`�j��Iv�|Xc�c+%�x������Oys�\��8�4�J�	a퓺dU(y��'�Li00O��o�.�MSW�i��X�iU��OX�1S�Ї��a� P��X��>}�����(*�ΓO���O��[��B�-��M,-�^L�T�����4U��ac��?�����Oov ��&�!SbT � "F;�p���	�>��i�f6M�N�i>m���?�0�ԛa �%�J�(��uX@�0e����f�RyBa���f�ԢHC0�#�##5�Sf�D�f}j��9,�\�t��@�*�j"n4rh,KEv�'
�nE���,,U�p��Y�_l�#nXi��bD4-�U�v��=JX4�cB�Ns�8�ᚽ{v.�ST�@>+=��lZ��&L�/·p��(��E�7��������w��,��ȵQ�HPZ���5�*=�@</-��E�K�T��+ЈOm,R��ïe���w��	���X�G &E��g@H�B�8��"$^�X���@Ӊʿl*ܤ��9 ^��(ժ��<B��Dr��p�A�RlӤd+ o�u�e��~!���� �-x�����?�H>9���?�a C}"(."R&�# 	�0��5�q�J���D�O����O�˓dG�eZ���ċ�ta~9�"ܓ^�"�F�l��7�O��Ģ<����?)6Ņ� �WGH_k꜡G̧R,��:��i���'��Iun�\�K|2����1N[hЦ�8o��rӧ�48�Dn�@y�'������O���MہR�YA�7-�2QJLU�E�Z��M�,O��qj��-ɨ���$����'� �Q3���`B�� %H�ތ�ٴ�?���5rF̫,O�)�Op��x҂���Q�V�i�xI���8�M�#�>%ߛ��'_�'�$�;�4���8�?�|1�ClH4a�P��Ќ�%���oy��'���Ϙ'��~�˗�n���krH��x6��O��OΥ�a�O�i>���֟p�!��>�V��qɛ�Uۦ�0�B��'*r�'@<���y��'r�'�D����e����΅/��q@�f`�6���'��$���͟��gy�ΈT?p���BćtE��h4E֦6��O��;���O��d�O�ʓ{(Y��a֕^���	�K�,b� ����]�'Zr�'��[�l������s�1u�Q�JN7W�N����,��c�4�	˟X��[yr��f����!M�X��֊�.�y��, �)����?q���?A,O^���O|�"SV?IS� J�}���2���� �̽:vb�>Q��?����$�dD=&>5�r�Jrd�a�_�4�����M��������0v���j�X�C�g��JuB�c��*c�i;��'�剛r�n�I|����:A. J@�vh`��䅆d�H�n�Ey�'.J��O,b��M�peԧiDljĚ�?�Ġ�ЇGަ��'�T�Flu����O!��O,P�M`̨�a�kVp萩��Uo�ٟ��	.~Q���)埉'��(��Ê�P��YpE�?0(P�4`�\1#�i��'	�O�BO�)�!2� �]*�F�i�b]��n� ��'J"�'���y��'�����Խ@��8�i�Q�bP:v�r�8���O8�D��Q&�����4�I�S%�r��t���K�2(E{�O��d�O�YP���O������0�-�&|ZZ�c fݦ*ں��!L{Ӳ�D���ʓ�?����?	�{ �0&�b4��A�B�쌻� ����и�ե�Hb~��'��_����Q�PD��b 1`̜�P�HU<��q� py2�'���'��O��d�1�T푷�8���-��6���ū
����џd��Sy��'q�a��ܟ�-�FA��P���ǚ����S�i���'�����O#Ӆ����f��-+,|Ӳ4h@h℃���$�O����<���cU�y�/�v�d�-o�\����&cے��U��$e��nʟP�?I��M�Ų��F�I�4���"�.Q�x$堑�
F,7��Oʓ�?	�GS��I�O�$�nakG��C��E��L��ȄA�Cn`��?!gdW�D���<�O����@�8!R^ȊhԲ?�&�ЬO�����&8��ğ��������gyZ�� �,stJ�	G*%�HTG_8��1X�L�I�{�$�5�)�)��A����o�8�����(dr7m^�t��O��d�O6�i�<ͧ�?�gQ�h�[�[�={���Y-^j�F/R�P���y��	�O�t0���0�ES�䎿A�DC�B�Ҧ���������i�^앧�d�'���O��Hfl��*wz���Ѹ>m����Et�^�%�c��ΟX��[?12'��1_ ٱ b�2�
|� ͦA�	�<1B(�'��'����#5����$��L��|�dLȠT���$Mʘ� 	4?!���?*OP�D� JO�H�&Ŕ�I(���n�_�\���<q���?����'2�Ɖ2���1T!�[06�Õa�Ŕ�X�������O�į<��� �Bt �O��#c�&�~��mD� q���ڴ�?���?)�R�'���$���McV���Dh��+G�ά�����V}��'y�W�t���z�z�O����%����Ak]2M6Ja0�'��~6�OH㟄��	3���\n��2 i���+	���nm�p6��O,˓�?�w�] ��i�<Q��<�j���j-�RRɓ�<ld����<! Jr��u7�ܸ&怳�@��I}�ѡJӪ��$�O�q�"@�O�D�O����V�Ӻ;1E��l=�x�&�,G�P8�C!�L}U�\�3h=�S�S����G�SD�b 01n�6�7
8��D�O����(O�)�OR��f�]���Տ@v�L�R�(C_}Q�O1�l��ۃ���Y&,P�>d�IPɄ$㦕mZ۟ �'N��'\��������t?y���!�`l���L<��u�'8�1O�{�;�)�OZ�����R���!N���b�=?���KĤh�T��\#lpʓ�?A���?A�{I߹w�&�ڄ�6y DdC��[��$ՉI�N4�֝� ���L�'� �yyHْb'V�B�`ө��_^�}��V���	���	^��?�F�ӵd�0�Ĉ�$O�2͘�]+#��Q���\~~��'`"P�|��Z��N_�Ũ徲�j�	��B��$���i���'R���O"tꗅY1���j�5?�ܵ0�E��[�byjkK��D�O��D�<����H�+������K'd����Іw6�X`�+r��o�ԟ\�?��X��$!����I~�VD���.-x�|)�GX�r@�7��O˓�?9�����)�O����,�8���&؂����|=Zab���m��?yPd��<�OѼ��͓>S�� �1�� �O������D�O����O���<�;|� �!�F�Ao�e����v<�'7�:x&m��y��-�G���:�#4�L����5�Mk$�[�?����?�����,O���Oh<��	*�b�*��[
�(ׄ����s�)�3.c�"|R�'�k2�b�����)[�"!p��i	��'��傭?�i>���ϟ���M�|౏��NVR��Ԛ6�\&�dls��CK|���?��'M8�IW��a|���c⑻a��Y�4�?Q�l�����O��d�Ov���6NUg�f�0B'"�l݉$��>!��T�E~���'��'���؟�+�ӖH�����\,/����O	�8)�'�b�',����O2�aǅ2Dr����晏1�� "`���ոӘ����֟\�'����>+m�ɇ�V&:�Hdfc�ZF�ǣb�F�'�r�'��OL�$X�Z�tdְi .8���6}����a)�O^�$�O�˓�?A���&��i��c�� ~�n5��m3D�Ԙk#�c���5��x�%si�q�xBo�7Mv�iPB�yP���M�������O��̻|���?���g���:�,S��agl�nt����O|DKV��{�1O�ӐmRĘ�Q�L���]�j
y���?� �?y����D����Ӻ{��
$,B�9f����Ό�f�]}��'�4�K��������O��	���K?-����_%'���j���8���O�}�8���O��<ͧ�?a���#&�z}�DE��6߶�e#�`��@�;dlV���y����O���&�;[T�m(���4M���H0����I�����.D䔧�T�'W��O�:��Y/ܘ�����,0o2� g��V̓21�-ؐ����'7��O�,cf��s-���h#J쥘4�i��H��t���4������=!�DY,��
4C��n����ʑA}�	(�"���O���On˓�?����,tʚ�m`�뵬[�1�)O����O��%��џ��T�7� q���u�: ���](n������>?1���?�-OB��&D�@�S,-4�S.��8i��(�-ˣ	n�7��O���O��$�I��XD�t�Ԉe�V`h�MhF,�:`u`X �^�����X�'����;	��S��ಇ#�/QVpX3�]I1@�RJ���M����'��A��~��8�J<��_w�y�CR�S� pSE�٦���ky�'��,��_>m�I��P���*+�-������8cQ
h�8��}��'P��
F+������	�?[����a�_+�%sj�eF��ϟ����ҟL�������?i��u�.ź'�NiXA��\)�5b�Ӎ��d�O��X$MΜ"g1O��t8�%��tLXH�h]3U$� Q5�i�|��a��D�OV�����1�'��	!i�0Hb �A
���m�)YI<�4D���Ex����OJ$�a$^$@W�0���)%��\�%J�Ǧi��؟���� �F��O�ʓ�?�燎 ��+�35��p a"����Q�i��V�Ĳ���?���?!�ޮX�Rp��	 &`��4"�(Aۛ�'6�]ȁ��>Q,O��d�<Y��C�aM�NX��Ӈ�F	�8�!�j�s}bN���y��'�"�'��'��ɀU$\T!c)��(9|lT�Q�$�����E���d�<A���D�O��$�O4�b�r&nH��W$
:���G���p�1O��D�OP�Ħ<U�U2��o�z�hr ��h�,��s��r �v]���	Xyb�'L�'mt�!�'�P�*el��w���V�_&�Q{�$~ӈ��O�d�O�ʓ8ltk�_?�I�}/"���  m2�@�ڪ\Eb(��4�?)OT�d�O��N.}�Ib?�I�O^��H#HѾZ;P0�$�ަ5�	�,�'�Z�$�~���?A�']���a$��Ę���=# jx��V���Iϟ�	]Z����D�?�S�ʈ<�^���t &l�BEj�t�08l��iq"�'���O8&�Ӻ�r�����ڀT�Z�ca혆^����'���8�yR[�,��jܧJ�e��h�/:m�c�
E�m.�m�GU��4�?��?!��V��	JyR,�0��]A����U�1
",7m�9>��7��2�Sş�
7�V�m��r7%�o^<�:'�;�M����?Y��_�P`��V��'�B�OΤ�	�%N����m�e���jS�i~�'���*���I�O��$�O�l�u�ݘ+�8�`S�B45��P�g		ߦ��	�~5��޴�?����?�����SP?	�i=2����'Ar1;B�q}���y��'���'���'��Iw����%�30n3AK��R��}pu�_��d�<����D�O���o�PX���f����.ߙ�(8ҋZ���D�<����?y����$�5�xH�'����(��t)����\�V�lRy�'��Iҟ��	��HF�k�4IanM�[)�a�<zmB�	�A��M����?	���?�*Oz�i#A�}�T��5�&5\�R�H7O�x�"d[��H��M������O����O��k�6O��'�l�Bf�U�
Щ+H:���{ܴ�?y����U�]�U�O}��'����ʜ;J��r��X#S9����Ѧ'��?����?!����<YO>1�Ovf5�U���K�:�bO�qܘe8�4���Z�;z
�oZ̟��ӟx�S�����fD�D�u�`�h ��fҴY+��i���'%jઘ'��'q�D��b��Xea��"KcH�X5�is����l�,���OT�d���'�剆��%)��̾abB��7!����4~J�T��?�.O��?��	�B�nl��ȤW��Ik�*�`��	I޴�?����?�b�5]���dy��'��DM�[F(��k޿r�4�"Y��K޴�?�/O8�
?O��������X؂�+l�x�	�V>kh{3�ǋ�Mk�=��
P]���'"Q���i�Y�"�T��2� 4�V�8��I���>�a��<���?���?����DW�H9��1Ǟ�?� �b��1P���y}�W�$��Oy��'���'��	7�MH9�2勝����'׶��$�Od���O��D�<�G6I����頄�P
>Pj��aL >���P�t�	Hy��'���'���8��5� ��X�֜�Q��l(9
�Б�M���?���?1*O���r�^M����5�D��N���ٗ�#���O���M{���$�O����O���66Oz�'���s�ˇ�|�ʅ
�5C ���޴�?�����z��O�b�'��t���℈��  �(�/T	��Ó[�D�	ϟ��ɟl����E��^��Xz\���C�]�~�S0�C��'NF�e&~�z���O^���<�קu�
3[�b17�[5`x�QA"�Y��Mk���?�%��<��Z?�uܧwf�ݨ���Q��En����nZ�W��t{�4�?��?������RyB�Ɗ�,dhB�;=\��̍�f87�b� �$<�S���� 	W&v �0凍e�& t��)�MC���?��V|��2X���'k��O� �#���@�nܣ�̜]�����iqX�<Y!a��?)���?�#��!5k��Lʍu�uX���-b���'�>,�1!�>�*O:��<���#�,߫���A�A۵;�"Ƞa��զ��I2u���IƟT�	� ���`�'��`B�L���0])g@L�>0��"S�D1r����ODʓ�?����?�uCYМ�j�$Q.lS���!���̓�?a���?���?!.O�SaU�|�k5$�fԡ��%�ެq'-B�I��%���	蟜�B.}�t�ሁja�h�Oװ&�P��Y����O���O(ʓ`Rn�Z��t�Z Q0�����K��p �N�T[�7-�O��O���O�ћu�$�+$w����"Q�Ai�h�6�v�'(RR� �B�(�ħ�?A�',w�X���I�*���b$�"4��l!��x��'i��:r�|Rޟ�%�UețV�0��f���1Enq�ӿi��ɌL)��2�4"���������HS���c��d������/Λv�'m���y��|��ɒ�;���4��� ��ӱ�]����t/ 7m�Ov�D�O����d������1�C�^*�@��n�:xQ�%��M��)��<�K>�,��ʓ�?Q��Ӷ�`�bI 23��� ՏL�uk�6�'^r�',�� 3-�Iӟ�%�Ȍ�Ć%B*v@�5�7P�T4�>a�"a̓�?9��?)3��%t� �`�d��k��6���'�Z���=�$�O�$���8@�e��>dhmSb�P�6�^�zeR��w�R������՟��'�T(x�n%vbb�S�@�$Dh�d� Wpc���A�������� ��A%�%R@�ڤ�ױx�t�J�O��<)-Oh�D�OҒ�R�"�+�|*�O��Q�.�KT��i�܀�FGy}R�'��|B�'�R�@:�y2J�`<��q5�\?��qPfM '����?)���?�/O�)5�O�S?D4P�Qm��P�$��0A�zMpߴ�?9H>���?���Y��?1J�X;�7x�D�!��u�&��@|Ӟ�d�O6�(��А���'h�΁&#.���0�<��M�q'�&u��O����O�m1��%��h�6���et�P+G.�&ITh�����'v^�@��`��(�Oj��O
�#"jl��P���]P6hF��Uo͟�ɹ���Iw�Sܧck"t���~�V�V�j�nڅf���ٴ�?����?9��j>���d��qz|݁!�B�h�������o,�6mW�5v��d�O|�S�Oc���&������u@dd�I@�7��O��$�O,E!1I�<�+���$���:ҥ�+>*:�9�ۍQ*d�Q�9�	� )�b���I�	�&s<0��O)aw���)0��Jٴ�?i���?��^)����%�4���ڿH�x�P���u|�*a�@��dֆG{�U(���I����Ioy�Y"v?p�
����k3ܩ���ιzY�uhwo�>)��?���?ٍ"K�;WxJ�K�.Y���"��f�92��|b�'���'���'7&�iFޟ��ڐ�(�\�NA�9���f�i"�'�2�|2�'�rA	)R�h�4�Έ��6x���i�::�u�'���'��'f�jǯB���⟔�l���q�ón��ES��M����?��!$�!BL�	�	R Q$͓�úa��Ki��7��O��D�<񦊍r*�����?�H!/L�!
�po��V�!B�å�MC��$Q�4�O(���$����-�l`6�@�jM����i���'��!�1�'��Y���S���i��Is�ۤZCR�3p�'F�f@�!k���D�O��ɗ���1O��m8��J�Gz"��%�	�lCB�s�i�ji���'�"�'qB�O��)*� ՠ
�0Xp�Z'8Ҁ����Ϛ!������p��y����O�����]L��1����	��Y즩�I��t�I�e(`Ր�}�'%�$�?v�Zx*#��.V�dH3,A�S��O�����OD���Oڙc��Ǉb��[��«yv�1"�i���I�*�|�cM<���?�O>�1Q��}9�cXj��Ґ�V ,FP�'~9
�y��'V��'��I�q���32F�d`l�q���5�&�;�LK����?A��䓿?I�
���PV��"�:CЎt^�X�b��U��?����?���?�BC���?YV ρ&�H���I�)Ҹd��d�g��v�';"�'��':2�'xp8�Op���Gs��x�������ڧT�PB��	�L�q�*�"H��(TD#�����h���	�nV��a;0"O��0�LO�?���Ή�rc~����O��	��6vI|�KC#]8b���&��z��WE�> �E�2���uPf��K�!{
jQ����?�%���T9Z����d&a�a��S&8�%�FL�?Gr�����obE C�_/v�����87�@p���#���5
Z���I�� ?8����L��l�Xq��%#7�n`�3�'���'D���%E�G�uY�&�Ep"F���n&5�b���S�d��'Dl���'lO�l0�dW� �zEDO�]��S�fG�#��S��?A"@�It���+҉�P�"@F)$"Ġ����A�<�f��y7-�.�P�����z͜�K�K��<�����>A�cr0����"���!�y�'��#=ͧ�?�F��&��y��I?v�T����?I��k����l^��?���?9��tW��O���ON�R<�&�$�:�k����$x��P0�I��&'���$۟ўhb�G�s���$,
�Bڀ���?�mx��*�9�ؑ��ɵ?�=I��@�JIY���fIT��F�M^?iBH
˟��	z�'��I��1��H+H�:��"KG1:�B��*Ֆ�(�c,	�:t{����Rc�J~���)�<!�=W�����P�-�!/]W�F����E�]�r�'�"�';R���'R:��0#��M���s�ŷe���t��4GZ�h�G/V[���E�0<O�a���K�TLR��G?#��uc��?12 �Ai���Dz��0<O<,�A�'���I�/d��3���!�:q���ף�ў�F2(@�I�u@����p~ )q�M��y� ]�6��eC6c8�h0%ؿ�y2��>)O*a�1�Y}��'d�S�	Y�M3lL�ry�m�A�]&
n<���J�П�����$"@<�ı(0n0B^U��S���j�Ha��'��X���(Oh\:bB�	z���!P�̋�ҁA�&+O��%�k�p��V>)�rB�0�(O�� �'���	Ԑ:�0Q��-J\��jヵ,�d3�O	���
c��-µ�0v���'~OV�8�IͨPj\���2rԁ 02O�}�fE@}�'�哣Bc�1����,�I~�� 6-)c�q����O.a�-O�U��)�2�Tj�<թ�S�T��'+&<Z�)_	p(t�Q�I"n|ܡ8�b�?�,-vdM�:�X��%!�JN���c���� P���{����F<mŸ9�7���:���O�S�SM�I!)��buEϓG ��h��61{�B�)� X\ 4�+At9R`(�����5�I��HO��{t@Y�)��$	��P"c���ߟ ��#�{5
e�	����	֟0	[w��'�lt�T�0�ؔ��=/��x�'�^�q5`I�R��q2�)O���ID�(���)p�ďQZLy�A�Ob��D	��J��pNU8�����H�H�E�V*:�� ê���FJ�O,�� ړ����.8�^\��I� j"���㡂�nJ!�D�m���h^^�Y:4a��B�Dw���I�<a$$��i#��D[�p=�i�WF�� ��D@��'���'�J��'>�j�JeӚ�2#�Y��)[$H�HD� fH'	�|r�O ��I%�����A���jU�N�$�.����;�&c�*����p4(�g$>b��7+��I�	fyb�'��O��+.����^63�t9d�h�zC�	!�n :T�ļf0|�i3M��H�*�I���<qA�І;y�&�'AB_>�"w��Y��9��*�B��u,P6m@��	ܟ���������B�S��o�@l]B��G�E.�A�#�� �(O:��0�
4%�>UP&&�.
*V@��0�Ĝ{�A7�tQ�I��M;��i9�^>c1KU�0�x�"���6v����GU�D�?E��'�bz��
fn�yg��'I�M2�$ډ'�@	8�.�2]��hA`�мB�]˙'%^aȗ�m� ��OX�'_D!X���?	��J����BG97��!f�0��(/������T>#<	��?�B ��IW<5Ų�Kk���h������O�l�f��`�Ι�U�@�%D�P��A6m�v���O^��?�D�� i~݃'��JǠt*�N�&Z����?1�>�ԥ	6dP<!nܹ��U=t�j�Gxr!'�S�dJ�[�U�Ʈ+2�1`�a."�B�'\�L���>v2�'���';��ǟ��	�Ȅh1��t),���Z�v�>�I>(V$[�G |O&嚑�_�@�&@�Bߴ�;�O�q.
�6}�{�J�$_D `5mX-y�F����9�D V�B�'F����O���4|j�-T2U��`�0gDD��N��5K$���!�z�����I!i隡��fy��	����1d��X��H��@�٤��9g����Iܟ �Iݟ�1��ȟ��	�|ʆ!��-c*h1�4$ɚT��y�t�y���ri*u��I&K
5��	�E{$V=h��<��aI�L�����6�O6Y�s�'97��]l|qH��cJ�UpD��:�,o�ϟ��'����?%yc�ޏ
�.���h�A�x�T'(D�`����F-p�� F��D��1#z�4��OʓH���3�i�"�'l�S&��rGPȞ�٧7iŹvC��Iǟ8��JT \D&e[DM��k�\����K(���*��eP$��7#hp`a�ү+cQ����ݕ��q�A�7B����$_t��@̂B�^����2/�1ڍ�dZ�]���e��mZğ��O<:��.  �ze*�;@&���'��O?�Ʉn<�$EI:Map�YgML����$E�	����!#�3R�!�ˉ�h���'���9�!�ٟ���ğ��S�,�R��	֟�ɘ8vl�`lȠ@ \H�
E����q!�0�"���ŝi�*��I0����i��\�X����FCS����C�5����(҄]4�ј��_2�K�k�X�0�%�I���M�1��h�-;�(l �!Ͷ.��I�d@�O?���u����[;?x���fk$:!���f���ȵg��B�/^�"<2�i>��	<5|���B�,E�8����;lP�I���X�fAE+���	������[w���'�ȭ�"֛;)�-��(���)��'�p2i�z|a{BHEXZQ�%�T�]8���Ũ�~�V�J��b�'pL�S�W�|!�fF+���hd�'�X�q��'d6m�����<A�����>�hq��Ë��51��
�!�d^�# �}��SQ��AeeN�zHEz�^>��'�4X)��u�,�ㆉ'4��lX ](:�H�U'�O�$�O���� *u*���Or��8�J��C���m�bd�'r���V,E� Ў���,�O��B��ϫ�r6m#O�<U��2��$l̟a��|�n�0�?��i�� �����b���P#��J���l�n�d�<q�����i��[�DR��
�0�F�yd0f!��@�U�b�c�)���>-��c!}b��A}�Q����������O:˧P�@��+V�X� �j�y����%K��?����?���i�nlr%�[�b��UQ���'H��P''S\�����?!Q���ă��)�r{���ED�/B����)@ʌbT�V���<�� �Q���o�O�n��O�8d#&�	�8�� 
��N	A�'���'szm2tJ�F�
������E��h�:���� ��R����i��33~�(T<O�豒��������H�O_hy 1�'�b�'ʸYw��]+�8@g�ٽ0�zա�� E릡@'D�BY
�M[`i �'��Ͽc2	�T��6&�6}��r�B&& ���NQ+[
(��$j]`*�{a@M�8�T]�u�ӯD����ʭzҤ@/oȒ����Ϸ=+�i�����&M��d�OH��?D���V� `�����6������Ut���?��,�8��&BT�N��1X���Z�X�Gx�� ���IIu���Gm�8,pyăN(a�����OL�ha��,<<����O0���O>t���?Q���"U�w��!_v�����'B���U��A���Y������3,��]ɂN�� (R4	��bQ��	�C�LY�vFU�s����dL�H���sd��
8�Fy����F��$�G������-*�t�'�2Z� z�fB;�T��l�]L�I@PB%D�Ѐ2l�V�iXq:������^#=q)�ޓO�.@�ȣ��7s��pZA�̑),!�פ
�*�Rv��*h���p`�Q�!�Dú!�APРO�	�<M[��5u:!�$��p�b�5�+r �xc��,!�$/X#��C��.xuX��BC��D!�D�KW���a 8^��2��T&B(!�U�fL2�G�RB	J�Fھ	!�Ԧm�a��]Rᒜ���$!��g���&.�C�8;�ƨu�!�ŝ!>6EK�>>V� �U�M8�!�Ȭ]-��Dl���|� ,�<�!���1O����#�g�#�)��!�d��G�ޑ�cjߞRT*Ԩ�'%�!�$@$�`���	�FVJ4�(H� �!��	`E>�5Ǌ�^U@,ф�5@�!�$��U�fn7:�8�c;.�!�$_QL��'�̄# h�r��3�!�ءzdHH7C����I!�3A!�$܉�N�1�U)?��hUe� 7!�� 1�D0�ӷے�BE�81!�d�6?xH��,��9�y�L !�U%emP���j�
5�d�Si�-�!�d�$l�LE�@šw�<Tx��
�!�$�->�P#��:�lb�M�?L�!�D¦Y���0��ѪR��u��, �{�!�$ ��m�1�.Z�V�;�БE!�D_!D7J��'.�҈,�!m�9!��[<�r�r޲�������"O��ڂ�Ӱb7:T(�f\/!ּ��"O$�TnM�x�4�"�:MШaȢ"O �K��		#�,��v�	 dώ)#�"O�uj�d��P�B�խ`D�8"O�4���׉lX�xЇ��6Ga�=!�"Ov�#���-]й��  pX,#"O��[���*1�CFA�f^]�"OT�OZ)C ���
@�U֖<kJM@{��0@J	;-��d��v�Tl:��e��EOڄ�;y(�E)����n]���E��kr�]��9��D2���!G�٘�L�h��\K�č-s9�s6�y����	����a&��#Nf8�5�$ϙA�F���
D7#B�&�H(ax2�_,7�:�� �
1(�r�c�e�L��G.?
�D�y cZs��xSR�d� ��"�{b�K�+M<I`�#��[���q��ޑ���W:M7�8�e���GW<\ju��I��d��~���9����)��SX��d�D�^�{Dj�b`"O�`�u�z�!��X W���*�?�`�!-�8�eA�i����p�S�D$�kژY9�w�P�CtI
��ԙ�D���_����''P�A�#B�8p)��'r��fИ�?!ֈ�&4Йsd(�T��Kf+%&�QjF���v��!T�J|���	x]ax�����5��*,���D�T%-Q�H�0R��ei�텡
	� U� ��)aq�M�6^�{Zڎ��pJ��T�v�85�}�Y�')<��fj2���b؃w�^(��\/V���b�4G�0RH��b�n��-[.�yRږ�����wK�!��_J� l�M���}33$�fgl5�Vʶ[��Ӳ����Q�j�"�䙆z�b"J?n�X���E����� �P��6�E+��OJ^sT~Iu�M�O&8p��X>i6s��&pg\TY�h�3���ѲhR#��H s�U��?1�Y<m&43F�d�? 왋a%C�5��%�%.'y| ���بO2%Z��A"9"� r�� -�|���Md*��c��y�n�bb�7.�eb�Ù{�n�����O�s�L`:�����~ʟ��2��T�t�k���e���s����
�8^8q�떃=&�Q�⌌4�`��1�w��9�Ӯ{9�\���Td������(s(�츓�ڕz�N�B�Ț�H���s��:w Q�8��5��d��ltjE0��S�ǒ��'E3h�6�t�j�9���|�>}�JA\���#b-J��F�:-��y"�b^�E{�fU�cP��F}�BQ&����aH�"�J��B�F�3޴w�� W`V9a�P)B��a��|�� �3���k)F`< ��(���	��	Ӎ9f�D}� mB�*Ee��\��+��� ���%8�@a��ӟn(�]#�F6�?�
�1BC����|"�N2��Aw�P`@�Y�S�r��an%?���I�Ne0�;�,�:T(.1�H�I�U��4V�RƘ�t���\�\eP�/:�y��L����2�?��M	#L�D8QE\".2�'�r�y�	c	29r&'�d)��!ǹg0�3�(��اu����~�p%LO�V�����L,�p��(B�5(���HO��Ѝ��W��$��*�5Z�͖a��9E�>i��|z�3n���g'�b��D$׫tH�pq��;*���G}2'���r��D��/Wg�;gA�hA�U�"ﴩ��o�L�*�{�E�<I��A	n��d�ߟ�ɖ�H�c�Z-2�A�^?0`:��7s��Q��	"?�p(_=.f�̡T���?a��f��D��`C[�0������~��@��s��K�Ș��~2�O�d��%N8Nlu���P��-��(����� D��G��	��jp��U�Z{�	"#<�C'�Z|��BD�A%�N )���<��O
 ��V��8���S�E���� A'�T��%Bݷt�0�[�.O��Pr6R�XD�$�Z8O����$lB���F�=I�`�u�p����G��4�8�g^��fГCj��ē��̢#?O�Rv��T�+�ۧBȣIf���+G�U�{& M�Yq8�ቤ�������A�͈ǁG�d�܈#�AH�A:>�)Gl*;�`���ky�4Z$����1�6	+0@�te��Ba�/}��]�"4!s�e�T�~�r�g�!���$)��P�L����)Q��$.���h�؟rb�����#j	���k��+%/V��s4�����xrɔ�O펑�@�%�F��n��m�� �H3KĽ��`� L��?c�T"t&�4-����V�� @�p����S��J�H�H�D��� �T�锯�j�e��`�tyr�C^�$�҅T)�y�A8h�i���	98�"
���>	�+T4"}4I#*���|U{�jV!#|���E�@t��Oh�I$e�|���fŌ��C!�>Ati�����#�ݥO����� �]�'�\��V�&1�	bs�c��0�'^��"����Xj'�;Sʜ���-~� dI��6�z�1��9,Oz=Y� TS�Pf�Tz�	����!��؉Dt �'^�g� �b:}*�蔨��(}P�����q�����"O"��A��5s~��:�L܏yR�8� ��_�hY1��N�cH��Ş_��u�q���1�O��� )҂d!ꑪ�/0D�t{1�$	������T$�����\�W�nI�'VR���?��Ϙ'RA�/� ̭��g	 T��lZ
��8&��5��-$��R�?m�ӑ[�P(��JENԈ�@��dB �A�"\-Te������@��ƍ<����REl��yU	�$�h�ʇ��;o�TP��!�����,ON�Cb,�.�`ȧ��"Q�m#D�'��H�`:'� 3b�cyiwHY4Z��Q�K��P�<�Ѥ�yҹ��9�$:mh�*V��� �����* "�����X̣�y�&�3�MH�tPH��T�>U S��9��0�'�N�0�Q�u����iK�h�0):@=OdZ#�O�	�5�b��G\N�4� T-ʉ�@)��OZ�ӂ! ]	@Ѫ�:Mr	u��i�r �ia���D!��T�Z�ц)&?���	�}��r���	pB ��&��XD�q�ӂ�	��>��[�1�N00穌)l[2̑��B�Q����wڹ�2-�>�>%�'�<�3�5O�|H�wﾘ b̔�lO4}A�![ ����MY�YB��T�3W\0A�o/Xa��"�[4>�i!(�`rv�D|#ܺX��y����m��QD�Zz�h�s�H�]0.�X���d�d�����,T䡑6牳n3p|�1&�nI�D8-��1 ��\�*�Q���D�6��%�>�����I Ft�)�H�X�)��Ѱ�q%ٸ�	B�6<q��	X<I��]Rӊ��/0k���<Ѵ�'1�غ�RS?������!�
gH��7IU�5枼3�g��]r�r���_��Pz�B͸��4��(S�� &(����I�="%�!d���I.�qOg�]?l�"XH2�QϲMR��Z�0>y�e��Y���G�Z��kҠ�NȀY��KE|X~�� Ŏz?A�RM����CU3<�~��$͞�3J�����K/<�"po�0f'0�Gx��7�衁���l�h�A�ή�yrN�<�ɢU�8G�!�ЋU6V��P��{�"��?	$G�Z��;f٧��9O
)�ҫȱ/��u�v��4Z	85��n=�=�'H)/�l��C�O�ؑoy�t�r�����w	l�2塎����P�)Ϩ6�ѐ����y�e(u�hG�-y	џ����

��a��5� ���$���@��T~�}�!�[@�I%E~���k��>� @�aɬa=	� �!I=扆�ɌT�KE �M5�� � 3�FS
z���j�*�ظ�w��$�0,�	; ��I
���?���'��k�� s3��W,���0냿9zz�Y�(#���aL��#�H��a�{{����Z�t&̲pc�DVDĿ<O��KwB���-	�nZ&%�T݉����4' ����<���9*���Ӡj�/N}��PZ�p��fo��b����TJ1�h�����̱
5�C*h��捗2Q�QyT�����s ���,Vx�"�*�y.b`�CO΂Dm\�`e�6�����*:t�-J���@֦lѴ��|��S�$a�|zL� BG0]1|4i�!H:ay�)bd�z�t��'��( fl��y��\�[M� �g�R�c�
u�!Ps9�T���9��@�]� 42�]�_E� �g�B�#z�ODlL��aէw��h�f��^�	����[Q�ٚ0mӊoP���c�.q��˧<���ՆxF��bR�
?+�ɗʱ:qNL��,f�p��
�q�O��	+I2	�E䌏C�F�B�jВ[��� K�0���: g�	*,�!�!ڧ�y	A��hĻ�ƕG&*�=z���ŅV�;~}�lC�6n�ѡ�	e���:L���1����Rb��= ��@#
>s��(:U�m��S�$�Er��8`�Ӫ#�u�p&
)�)�ózA8�8��'�p�*����q���]r����A�V2V����#o��"���([��$״@G{��;[�V����Y�r���e��L�D
�	4Ak�[F�_���'�P�⊙L{����@�3b&i/��A	���T951&T��-e
he���vP��kS�1��P��Fv�OJ�ɹ�"�h0��y���i�Z�h�T#­F���ٔ/���1�q�6ҧ�~r L�S�"93g�Ӝb�>5hd'���91&�38�+��C��� xu�ɿ-ǩ�0�5O;6���&я.��ٶ��N��]�kSj��� `ݭ�S�'3�v�F-�-%,ሔ�Eh{�$/�v�B�'�"�b�	�<A�-��b�#�d��@A�mR@Я[�r�jqx�'z���>]�Q��<!��Q*���y��Z�f��g�>M"�Z� /�q��$�++茐�bX�eF�l����:(E�O��*�M1Rԙ@*R/���0	K�2]�I�����ٟDA'M�)A$��W���`��N��̸t���&��m�:	���Pڮ�QygR1�6�>�Ӻ�I�sP܌��	ҫ'�$��H4�t�:��8 �x�D¾ C7A'OZQ�AZ6B�)@��E�C�{��-�!�D� �	�<�,5�Ӻ��(W 0���������L���(w �q >��3F�-���D�+���V)n� P�'�0��@�?�
��	�!y�D�!w����S�����	秘O����(;i~5+���6b��й�Z�o���;#��dd��Q��[���N?��_�ģ F��j��܁�}E���CE=}{��ϧ8��iQRe�������2��L�<�0��	U�{�la*dc�g4ޥ�&JP��[1�8}��?��a��3Wθ�e�G��@:\�־!9w휛a���r�A�c0���d-I�`y��
'T��K��z!�А$��m%�P ���PH*���?m)��wRɿ>�f&x��l�r�@c�\A�B\�*�"��P.#2\@�F L��q3&½!��ђ�J��~��u-�ty2N[�j�2��5o�O��O��A.Uo,(Q�5z�zw� >(�>A'@��AJ����L�;lT@u�e����'(h��d�)*?B����P�X��ɸ��IY d���ٺb�گP����O�=�Um�/q|n��6g��'V��r�ȃU���8-�YJtj�9.�1��?�@%�ɪؖa���'n΁QA.��e8�rw̨�p<�PoI�2EA���r$�+�#ȿOu��)W�a����Wf����T?˓���g��m;��<f�Qc��J�68s"�'c�0� Q���d/=�R}ٷ��%F�0�s��[��ɞm$.0 J���/O��M�@�k�^�����+E���!�V+�y�,��'�j!�bnW�(�B��Q�r�y�Ϗ9�	��'��l
�� O� �y��N�o��(��i�m[�	�����y�Hϸ���8��Q1����y�c�,A9��Ń�**T:���y�-V����9�-K�j 0a�D#�y"�:
@@M9���&�.5 �N�
�y����p��k4L�,��$@�yR��0����	I9X�}��%Э�yr��?6�AZ���z��e��4�y*Ɣ9������Uz�xPgI���y�ŀ'R���W: ��������y��]� �{�d
G[�3�jI��y�J�=!Ԫ��R�,?�D�Dn��ya��*Pz�7��l���ئ�y�NJSy^\�vCJ6�l���O��y�(_l�.(�Dl�+A�T$y���y�KT2c8�@���Ó!���t(P�y��@&@V�����f؉�%Â"�y�`�3�j�CEd��^erphW8�y
� *�u@J�a����F��)�E��"O��#��	���hw�7 ��"Or���ǲf��ɫF�s�,�g"OTZ�
I�P��H�rnH�:J\�	�"O&E0���,����g���"Oƕ�$���0�fъ�K�,0𥀲"O�ŹgB�{Q�����<sd\��"O Y��e�
%�:L����^j�Q�@"O: ��UJ�� [b ڜ,g09��"O����΄?ȱ2q�0,_� t"O���Ԏ����+Ο<r���"O��zEe�!N�+��Ы^g�
�"OV��a�9�
|�UIT�x����"O����%״Q�.q��'�5'��jf"O ���'� Aqt�8�k�@|"O��rv��  L��A����2��(��"O����]Hc=
��W����yra��Eʔi�&��7��Y���7�yr�W Y4���Ζ1�Npjqb�yBO�E�"�����.�DT�^#�yr�Y�B��DU#q����M �y�*�
��8SaKE�=�LKT���y"�ǧ<���y��4~�i���yn�g���[SJި!#���i�y򁚤J$|9�*]hw~�*���y����)2C�Xd��|���y��2V�(�0�^�\?r\ۧ���y�J�'��lRDT�R�0���O&�y��V �]2���{Ũ�ӕ���yB�
��Ez�l� {�.xZ�o��y҅��s�PR�F��E��Ĩ��y"��)b���-DAjX�Ĕ�ya�$|�u�,��X�F�"�ybh
�$ m#0hĕ]��yK����y��P�7����ch�2*{P,�4e �y���A~L��׬ӈ1��ɓ��(�y�,C�00��Z�yzt@��.P��y�g�&��\:h�y+�m��B�;�yBQ�\+�,���Īw��5PE��yB�^�6�cDp�^���G���y�aW�p�L������$�9���y�-��nH��@`�K�� DFL,�ycҀz��8�7E��KP !��h�9�y""P&^3A ���A�N�K�J�#�y�jab��3hM�2<.���k�y��-��49Q�F)�Ε S���y2�	j�ޕ	��%�����c�yb��>h)��+�.�xPA!��y�� ���`d� ����e�-�y2�L#�-#�B�.c���C���y&�$�!���&T��ݡA���yRƆM�Z�YS�ֻ�~A	e_+�y��D��4
ÍK"?b�at��yr�P�O�� �+��B)F��S+P?�y�kȽ`��lƚ=� `a���2�y
Ii�`� &Y�k����E� �y���V��A�Y�DMh􄅾�y�יM�� 

�F\[����y�ʾ{�`��i�7<�1k�+B>�y�b�h|�b2c���d����y��1Cx�zԯ�,^����ɥ�y��K%�lZ�!�7R�$�:ta8�yr��1v�1[p�����	%G��y"kgT��35݁�\�ht��y
� ���R�ս}� �,[�z��"O����f�D��8��MѤ���0a"O��3���&hQ#Fţ&��-P1"ON�p�fZ�
U$�1���o0Y�Q"O@��߲�,�(�n�
L�M��"O��$CQ���Xa#퍦.T"�D"O���cAVc�8�ʴ�\�T<*��"O�Y[��53�6����Q-e(Ԅ�"O�0 ��c)v��6M���IE"O����
{p�ib���G[b�aC"O�c�5jzN9����N����g�ID����/R:mj�D��dE�V/;$��]I9�љd�!/�.�J%�ueZB��M` EyDKZ{�x�JR�u�HB�I�O+�Dj�i��+�`K��B  @B�	�3�`��W�L�f��rA�t�Tb�@F{��TH�L�U������2�I'�G��ybI��6�@�9/�8�����#_	�yr���Sc&5���ً,�tH爞�yҀV�A�b< v#U")��2��݈�y�&���IC��]�!	z:P��y"�G�z��j�@߶��͙Rk���'�ў���뤨54F�e��A$9)�XQq"Ox҆�؃aP�4��ƀ�ly`7"O�� A�:Bb����2�*Qr"O:�`��R�b�8���jߜ1�f��"ONd��m��y�ԑ��ʊuAؓ"O��Ň�(?�ry�#H�mXP{f"O�AYSfH�t��+�@A&����"O5x��l�4�B�؎)�r-���'��	2�"�2dϧ[0�� i�v�2C�	�	�i�pӣ[ �d	�mF/NLdc���<+�~�F�;Evl�&��]��hA���<��d��^�gV�S�
\a��Ŀ�hO?�	P����"n'_ߊTx�B�z��C����LR~� $,��9�C�+Sfr �1��%{Ͳ�pǃ�=tZX��Ĥ��#��W*-�.%��HI�v��H	f�$D��x5ϕ26�����2S�����>D��ħ�?E�y��ٿu�X��<D�dp�gօ5�쫑���U�̻@ 5D���$�K�<=�#,@=.���pf4D���X�v:����/qĝ�2+&D�L��b�V �s�%�Z�0��"D�`R����NV�U���;�@-Ȧ� D� *%f�&ܹ�	"]��t8�� D�t����gu�̐@؋2U�8�D/ D��7� 7iD=#�ė�\�r�#��2D�hS���d4�J��
��@����"�O�扖�~�Z�X*�İ �'2Ib�D��1=������2i��A��9B�	3wj��Y#*�z �D��e΅ �C䉲CKTLae�\
C���"�N�^�C�I�e;�:���3uR�`҃ͣ��B�ɦ�������)�T��%A��|�B�|ʬ���
.-V[�a�;u$�C�I������	�^�<��B�ؼB�5I�m��jЙՄ�3�ģ�TC䉲X�p�r�eE$dT�|C�@��}�4C�	�	\|t�R�Ն8ڒ���c�A-�B�	>kAd���#Ï1(V�E����	�',.B�[z�p����)-���'J�|�U� �PX� p��><��ũ�'J�t��BD*D)p'Z�-`�Q
��� �x���JK��`p��@�56��r�"O�Q3%�X	la����%N�}+��ku"O�yC�G�!YN���$��J�@,j"O<��c��
݈#J�
�E��"O�XQ!ՑD��h�O����@"OH��B�]��Ed�R��k�"O~�v��
J+�u@�()��Y�6"O����j��r���s�ɕ�Q�^��3"Oi�ٚb���Υu�\��@"O���s�ʉ�ȥLAqf�隰�����#l��<@���?6�q�
r��$"�pB�@H�q�-��͗�Z�lz2-%D�l3T��1-l�5J�1n���y58D�\�O�21Ӿ����;U&��r�+D��؀aV)w�ݩ�B�p�VŸ�	7D��/�Rz�i
;C`t�2�Q{�!�Y�7�B% p�E�Q���BJ!򤛘xǌ���/ L�D�8G!�d�g����G�����	A�cƧ4�!��U�||����:!�Z�y7�"I�!���.����uU܀�Ӆ��p�!�d��}�H��q�'I�Y8�X�l%!�D׬|Bѷ!�`)V� �JE!�$�>�f���ԍ�\���V!�d�>y<�}pD�ɂfP;���a�!���/�4��d��Dq�v.K���E��B���r�jRCJ�=�(�f\=�yraV l_<�%�8�c6f$�yb'Z�L��(�A�й{����um���y" ��u�p�1�/W8v��:��1�y�a.\U���[[&��t�K8�yB�ٵB�w�J�K��Ъ����ybD��z׀�&ȊsB�`��F��y"hXx�A=o�Xh�á��y����qnz$)�,T����0�9�y�ꊮ6��JQ%$J���ѫ�yr�h��m�5K�E~�j1�R�^����)��@�@��p��M���tձO$��� 1lGT� GV0Q�~�2AVm�!�D�Ț�"MG;R������ˬ-�!�ď"Y�@b	�)��!H�&�,
+!�ٱd��H7$ɳÈ�,-g�	q�|"�)�S�k���p��]%��mL�6D8B�	�o�h-#E���m�9�P�H��B�ɩQ���2�r�5rw�InHB�	'^�
A���K
<x~ݘd�&)ªB�ɍxJHH�@O�M�l����E	3~B�	���@b�OD�'��QB���C�I/+L^��m��,{!����-_&PC䉙BT�� �:l���W.mlQ"�'r�h�r��:�ά1�b�#9i�A	�'�,Da�lǮ&7Ly��FA
,��U@	�'�' �U\��b����
�'4L�ղU ^]�2.щ�
�'6�9�
ߢ%�ִ�A(Q1r�=�	�'�ZX) Z�q�`�cg��q�䉈	�''|p�s�&/?i���n�t٫�'�r(*�B�?d�J���+d�����'$
4��HQ�2U�ibV.ަ[��p��'n�q�pAX�FS�hY&&V9�����'�>����ʖJa��㥧�ze��@�'�X�Q��L����!y�4i��'��\a�&M86ђ��A���x�'sn�:!d�f�$��d��'�u����  t��P���g�M�+�f��F"O\�hbʖ&cM" ����40��"O>L����Q��q��6� QA�"O����T�ekTm����2-��` "O�АO\��T��R*W34p01Z�"OrDە�ɛr�h��;+�8y R"OT�@��<I u��N��4k� ��"O�5'lڨ'F�3��QX|��"O�<Y�a��6��e�D�8�vm�"Oΐ㧂�6ni�!��&Ú$"*OV�9�F_�RL"�I �G#_o8��'��P���U O���Hp��4���	�'|�u��B�@r�(8s D�TȜ��	�'��X2B&ڠ^��Kʟ7T��	�'GjA�&�ϔJ5I�"�H�-@J< �'@IHs�IҚ��G�R6Kr�KQ"O8hx�/��(J�i��)j�t���"O���dʊ�Y�%�w�	�|&Xps�"O2�cw�"SJ<��j�6 ��"OH� �M.�J��giY�Q�B-�"O�Z g�Izu�K���-b�"O �*cD�-��<�V��]�"O���� �=$�F�Ȳ�ߐSz��3#"OL�j�
�Y{<I9&�8r���"O^ـ�aR D�V�YT�;�慸�"O"�Ag.ƿfs��ЂR#N�av"O����A��{l��ʅ�������"O{���qo�!M䠛�&�Q��`�ȓ�\My�$����5#��T>{��P��_e=�"��(x��
�nR;�,p�����w�G�9�6�"�D=!K~݆�v�zu���=��-+�&� e��Y��x�z���a /\@���U�R�<���'���嘋�rH:��),��\��}��A�%W�Tmj�)�
"�
)�� �q!�ƍ�sc6c�ٝ*,���x�m9��>����G�r�����K���a�� ��)�!߼X]���ȓe�:�B��J x����#��`xx�ȓJ�8i���!I���CT�g����ȓ����R��m�� �7�[�� C�	PWFL)p2�(3�O�rƠ��W,1���D�L�ڣb̿h!�d�ȓ����s�W){��`���&e�F<�ȓkq�b�	 2�đ""�� #�t���N����8��DH�Ԋ]�FQ��p�L�� *Ҥ!�b��O�����,dPa(����RlJ���4hލ��3LD���T�P�4���F��]=�B�I;Q6��'�G!�Ҫ�+&�C�	5޲]���*��x)���=m��B�I���/@��+��;3�=!��X�<��M)A�ND ՠ(C���P�TP�<�DO�LRR�S�DHti�� "�Pe�<d��o�ฃ�#B2㒰@�oUU�<�Ԏ�!'�ڸ��aV�J�PMF[�<Y2��QFN}�!e��1{�����P�<Q���>Vta��e�6mzHa3r�J�<��MӅ~�Z���4!;)3�@�<y�D$B2�&�1�|-` f�c�<IҥF�'yȥ�a�1,G��s�
y�<�"nF�*���rC�w�� yqBw�<Ah٬f�6����<t0���g��Y�<���y��a7b#i���ȠC�Z�<� �0I��J�E��Tl�4[�"O�� O�=_d�4��hOWc�%"OU�V�C/>�6�i؍y�tp�"O��]�wt�}m!�T��"OBLj��1eP�8��d~�� �"O�@5.ۼt�=p`
�
x��
�"O~p�.S���8����Wl��"O��8��Uo��AEh���(��"O�)fʊ�y6t+T�7#�8���"Od]"����hր&~�ѰE"Oz�c�ϐsy@l#�l�Nz`1Iu"O\�i#���	�W-� "x��!�"O&���j�/R���zE�w�p�0"OƀZ�@�XdF]d�L;.�fy�"O䁋�B���@�+��j��)�"O"I�fb��9����gΚ4�x�Q0"O�5�g`ͳA�ڜ����jv���C"O2Ԫ��D�!hz�"�Ƀ�]���"O�Sc N�@:�܂����3���f"O4)�E�فg�dD����B��	�6"O�k����d���p7F c�,(P�"OX4�S��Nn�!HC���-�����"O�� b�92�VW��!.RH��"O���!+)f$�!�u�SJGZ}y�"Op�r�HV�ZN�#c际/dz�rd"O�;�#Y>P�����
�(Y��G"O:5�ӯ�/������E�y���*�"O��{p�L@�b�eW�:���e"O��R1�64ٰ�*Bc�I�(�
�"O~�cЅرw�*�s�a�"��Hh�"O�X0WEW�I�T!��M�!1yb5��"Op�P���6>\�MB��#g║$"O$�w/S�9B1�B�C6
Z*�Bd"O���ǡ�kƺ �ƢP�	�ԐX"O�[Ǯ��us�0���)'��H�D"OzP��!�F����0 ��yQ"O���p�+{P�l	�O��Hn�t��"O*-ɰ�2���U��F��y6"O 82�荳W���ŉ~M$[r"O��Y��U^Za�0C/�c�"O(
��r��<q�ڊO�x�a�"Op��(N�[a$��Q��3�J��"O"M1&T�<��쓔#: `5�g"O��ĂL�À%"��4"OuR�ƀ'Gt1��!��2��"O��B��^�%j�I�4�X<a "O29��(ɣPl���TW�Ӏ"OQsրO�M:Ru �^(U�
�iR"O�=�$�H�M.�2�OC�X,p�"O|qC�_.<�L�F�	)���"O\�7� MIv0 �K�P�9�"O~�Bc	��14�Ճaeٍg����"On��#A�1��H�Ζ%[�´�7"OH�Z!,	D��X�Q�[U��c"O�T{���
Pv`�`�M>DMcp"O8���
�#2�-��j�)Q�\�#"O$DQV��p�LP�郃"����"OB�h7�SZ<�)x����^���P�"O T���d�vy�6�ٜ� �#`"O�`z��^#[�����N�i�f"O���@Aȳ!�U�pȞ�c~���"O:|�ӧ�ju:%ǜ�6Z��1�"Oh1����}��tyӦ�)S�%j�"O� ��I������)>�0�U"O� Ll�$��3MӬ��V�=8�x��"OF��p��.5��x2$ȡN{0�"O,H�DGq[�A��F�]��r�"OiH���[9�Ei�EADD��b"O
��B�V9~G&yQ�dT814���"O�H%b]�lDƄ�U�F�x�Ĕ�P"O�-aS��4T�z�Y��t�H�"O��
P���I��q����<G��!�D"O@��`D;P�N@�ǭW�+�E�"O�|;r��l"d�)v�
$�dB!"OL��f�2��� ����X�F"O�,� W�~�T�ȔcK6uM�"O�� ��B�6�)�b2qHH�BF"O:�����36��Q2ab	�O�D]�'"O$`�!�@~n�X`!D��~$D��"O��9��!�R�S�
2g!����"O�l��K^r�s���슰"OL�e��8T/"���t�,ps�"O�i�Z� |lv�]�[���H�"O�!���0	��[0��@�n� �"Oz1 BќE���,Ĳ w�u҃"OތsF�����̴/ZP�)�"O�heʅ��f��%�O�:Td��1"O܁[�]>���A��ZS̩3"O� ��R�%� �"�L�)Uq����"OR����m|  ek�<�p��"O��Qm�/T��s	�!�h��"O*��Jœ����D�W� ��"O؄xNO�S(tJP!W��X��"O��*��M�H�h��Z�?�άQ&"O�����K:b�`@�ޙ.����"OT��C.C�>��Z�H3HQ�S�"O��p,ܴS���`�8w�dӆ"O��2NJ(}v]˲��5Y��B�"O>t�%�ӿP8d(��$`c2l��"O��c#��9,qu	���z$�IP"O�%;��Ԥ/��)
&M#^���"O\�J/_�0:Y)6�%��Q�"Oj����#!�ꭊ���Ut4K�"O(4S�B�G�T����ZrH�5"O�5!�|4L�+m�Ky@�C�"O�1���,2�eE�Zs\��"OX�X�0`m�i����*��e�"O�5	�\�8���p�
�U��Yp�"O4�P�8-5ฺ�ſ~� 5iT"O,M�2�.R ����F��tzG"O�P�9"�|����	άD�c"Op�,4�#N��<OU�6^<z;!򄌋mR�l�rDՒs?�lQ�oTH!�Zr����i���\���k�%�!�X't��X�G-\\w`DJ�G#�!�Ě�IY�x��A{qS��`�!�d��9�
,	EGK���(O2O)!�� �l��A�G��Hd����!��*�V�`���4P�H��[�1q!�� w��4	�d�M'@���U)n�!�Ąw������H�<����!��̞q����f�jI�#��!�d�%@�z���-^�z  v�j�!��вI� 9�)��8m���F7Q�!�]�*�Ԥ{�iF������#ș�!�6}�@���Ж$�t��A�R�!���' %�C����!��Y�y!�Ch�T��\�Ru���͗7!�� N���[<+7̔��i8I۶�(u"O���F&W��;�*�=>&xy:v"OP���(K%`>�`�ti�-�z�"O���Ɔo�������i�Q�2"O@�c�����z�m^�u�ZA�!"OL�s�Ά\m���smZ�wVl`c"Oe��D1o��QҐ,�
w��	a"O�,VC�w�:��ג�h� S"O�P��#J����!�٤C�P�R"O�̢W$�8h���@bC��8h2"O�[�"P��p�C�'$�J�"O��7N��t��L� "R	.BVr"Oy��Q�l ގ	���2�"O����07۾�!��A��P:�"Of(�ajثU�d�����F�FX�w"Oސ����Ԁ���0M�ؐA�"O\;5'��T��Ч%��,�"M�w"O����e�2@.�R6J$�4"O����Z�_��T͐J,6��"O�<��F�]����C��n)��a�"Od�r2��7���A�)|M�C"O��:S�X�
#>�1��ݤW���t"OZ��G�ėE�Ɋ��7Q�%!"O <����;"�09HƮM�o\2��"Ox4pF�Ei*pe�U��U=.m�'"O�����
W��4���C��ي�"Of�2A��~��x�ԵnB�P�"O���pHۃ�.�y5gŁV2�mke"On�ҳ,؛/� M�GVu�8�"O|����-%����/�X�v"O��"��.e_x�j�f��z8>EzU"O@��fmI�*}����F*Y�d"O:��!��L�f��E��T��`"O�\q��ш3����T�fVnY�"O�9��*PGj:X�.Z,vH���"O4�wfG*/E��`�"�WD��s*O>@�)Bz��k�c���:X��'u�8Ӄ-I:i� U���N����@�'�>���[3�<9e"��~��y�
�'�Ē�f��Kg�H�o�zq�'��Ѣəqq`��E��)aZ�lS�'Ҹs�
ŷ`$�RuJֹ�� 
�'�6�I'NV2
,���d��qxFP�	�'�BE�UFH=,r��u��5^r	�'�0�!&�* C2E�(�XL��'�l��C��|�x��f��T}h���'����A�8{QC��W�w���8
�'`���D���(l��@!n�,��	�'*բ�"�%@��ȓ������'��ɓ����� 	 ��`���'�VyÖ��Y/�	��g'w�6x��'=��g$ܺha8��Tm��i�����'���`n�!���6a8V���'ޥ�`�K�x�8B$����@�'2")w�6P�l��d�%�@	�' H A�+Qy*�����'�X�0�4�%gE�H�d�{�i�<�Q�=D���6"^,�U!6"�]�<I�H��&�Ѳf��.�0]r�'t�<Qu蔕⾥��&�|r%�r�<�Ї�6�R�Y�ͼ
>v�Y�%q�<�d.RXИ�"�\?2��I���x�<�ժ ,]Ϯ<Xq�Ʉ��z ��t�<)Ӭ�%U��xz��W�S-�p"�B�X�<� ��ؠk �V�V��̓d� pD"O���Ѕ�
?!�hC�	�~ ��E"O��ČƢ܀E���ÓSLh8��"O�Bd� 6i�j��G2Kp�"O��Au�SgܾLX����F5�%�D"O���AIF�QB�k�h
�|��w"Oj4�4�_�]�  VM]P�
��g"O��v*U�^s�J4�V�=��H�"Op�b�`,x�8{���I��L��"O��ARJ�%V�DB�늵,�!�""O��y0��$\p0(�����=Ƭx#"OL\��+� $�Tx�@�pV��ɡ"OęC�p7���eʒ�����"On��c�|�(��d 
�0=�t"O6����� 6n��dީ��4�B"O�����][��1B�̈́¢���"O�(��d\��Fu�tf0UGDY�"O��f�V?	�x��R(V*G^Z��"O<0˃��a�Dp�E�+� ��"O�=�Q,�55�0�IFㆸ����"O��9d@Y�<�Dس��4�Z9�7"ORx�&ɉ	Z@���a�	m���"O8�	�'!U:�هMҘ\L�4"O,���(�9VИ#�Y��S"O"ę��T �J)�%+ZB�1�"OD0d�C)b\e�D0~-� 7"O�Y����I���*Ѐ�"O9�oW�^f��UB:�"OnhRh�7n�l�8�e"O�U�6�S0C���{%d�� FX�s"O%H�F�"4Bb1�5�B���Q�"Or�I'լ2��xC�N��^�����"O��&āG����v����@"OFD���Q���+�l�'��� "OB!*G�͑1Z<;׊��0�Ђ"OĬ�E�f����'1#h�(���p�<�'&�N��"����o`zi ���q�<)"�G1F����گH���ړ�j�<���<3�l��`�4?�( 2�`IO�<���7,G�� �
~�f$k��]v�<y�F��01�C�̆l4±��u�<Ya��0���j��7��q�s�<!��^i��9�R��h��Ug�-D��S�CO�A��	:�W�Shi�C ?D����ה3���������
�8D�p+U��a�ؓF�;;�JqG5D����)ԄgHn�KR�K<���R8D��Qwʎ�q |xq��;-$���D!D��Y�LS� �@�
�x\�,�PO2D���$l��!An b ����남1D���s����ScMur����4D�d�HϊL鐆��wf��A�$D�ܳS�����CI���F'%D�,��+-9��r��E��is�&D�\�{��k�D�.F7�ɨa#D�ԑWK ������M2F�^�!n4D�`b �ý? b�ӇBσL�,�*E%4D������U�~�Ѳ&��gnR1�b�0D��S&��u�*��J
(X	3D���ƿL��5͓�"8��1D�<r�e�%�-���(�=X#l/D�@jt�Że��h�7��9��,�P�+D�h�2�#�"'����(h�*)D�@�Ơh᜙�0,4X?p��E�$D�� �l!�,F}`	ڣ/`+$��""O\|��E�sȖ�څ��D���7"O��R���?y��;ҍ��e�l	��"Ovyj�TXu:,X�C��Z��"O�,���7EМH�fO {�z���"O���'��24y֐Ӆ@J���{"O���"�Z:}q�dŮ1�!R"O,�2Ċ�u����k��Ej�"O����@����TB
J��Ux�"O>� �9R~=(g�{���"O��A���;�"��E���Dv"O�ŋ���!="]˳�
>�H��"O�8 ��.c�Ļ�+A�wż�J "O�*�`ԧ:�ؘ��#R@V��Y�"O6��fI�GQ��ł߬38P�i�"O"����*f",8�B�^J>�r"OfL`䓇!:%BRaDe���"O�sdf�&mEJ i�`X�=����"Oh5I�J�~�$�A��H7fwJ0q�"O>�å(l��G����"O��P�e�'7�:Pc��(����A"OH�ȑ�#j���S2�2(�Q"O�5�u*7Q��#��@��B�z�"O�x7�T!2l:�%ʚ*D�u("O m�"ݪhK�!Kge�Rb��9�"O���tNĕFwfx��	�~RB]��"O�ͺçF#W3��2B�Ȑ""Ob-w���hj�A�4c ]0L���"Opt�s��<@�����#js.�"O@0���z�P��v�� J�dJP"O�:1&�-�@ �CX/)V̥�q"O���Iȑ-3�ҕ��3)j��"O�\���X(e�����\��xP��"O�}�2eG�r������K"�""O<|��ɊX����ͤ4�j�Q"O>9�$<`�K�>�| W,���yBd�"B�mi$��>�qC���yB�\b�"dY� W��}��JU�y�CJ�[f�����Dr�A���)�y�ʅ�D��pcх?�h�1���y§_�
_�k��X�>�b�!�׀�ybb�s�X�2�L=8�j���DD�y$�`Sf�2�ɘ�=״�b6��4�y��:U����.�1=N��ĥ�-�yR� i�n�pc:`P{,��y�.�0u����'B�")���y�H����퉶4�=P�o�yB�A���M����]7��ؓ�E��y"����ʹS�
'Q�R��g@���y�矓��y� �]�y��hj�,C��y��J�,U�󔮉 ܊�ӷ��5�y��5A�A �
�!rX9�Fg��y��̩!�("#��$.4��(+��yr"!P_�;� F���y��	D١��
n���K\��y2�Χ�,�(�%ߊ��
��y��nI���� 6�*�1I��y�\�q��	k5a��[��u�����y�Lv�r'��@�
� ��yb��!/r�%H�2����Ň*�y�gZa� }�Ǭ�&?eJ��*�y�KΩ8�~��c�G�
� ���!�y��F�2����`���7�(��hV�yV{�E��jka��xzJ�K��� �$�v���4a0D��i�j��6"O2ш�Gn&z!B��"f�f�a�"O���C���C���QR�Ջ?���"O�E�0nB�Oi�8�j�6i) �� "O�+�o�9e'��Gi�#F2�P"O𵹃�S!_N�9d�H�T#L<X2"OP���n��=1��$1�db"O��#��L�������e�,hC"OFT�b3`M0t��L�:F��T{e"O�X��G�fV�uYp�ݯW�Z!:g"OJ����	%�@e�r+�:~2��"O��c2%�m���
�IG�QS�"O�O3� dB�hՅH7��"OhP��E�6���[�H� 0����"O��0`�_	<!Q(�6��u"OBL  �A�BRѲ�`�~�|eس"O���������A#&�?[�
��"O�� �
+-D9��%���l8�"O6���;r��m�#�
�I�T�+r"O��2��+�ɀ'N�\	��3"O�8;�E��x)��ؚ�_�����"O�<���,a�^��􊆼N�t�0"O�\:��+k�çJN8�``f"O�����`�\�A�IG)����3"O����lB�Z-R�֦	�LX�"O>0��F�Z�QU�i��\��"O�Es�ǒ]�鈶f\,�.�"OH���\����Xa��Q�����"Ojp�-��v����܇Y��=��"O�s�l�>�� 1�ƃ)X��i�"O��r�GN.%(��*2%�8T�� bv"Oȁ�4&�9�2-rPJQ�St�= 3"Oƅ��'��-u��y��V���r"O�@Ò�	PΕ�H�%_x��w"Oؕ"�jǤ�G�7nF\Lɳ"O�� 䩛��bI*r�71Fa�"Oܵ ��C���R���� p"O���q�w�tdH����`+�"O��)�H\.>�`�w��8�	��]�<	v��f�X$UmU�o����<����a�P����|A��B��&����SAI1R p��;��C�	��:�A�0$�Iq'"�8,��C�����@�W(Mֈ��uߠ+>B�ɉQ���R���*�!�R "I7�\�Is����t�@1��"�-�S�_���J!D������+�!DE4�1q��>D��R�?\&Fx�u -CT�բ�o>D��:ŏ�	/���0hSrA��J�e<D�� �˜�[&�(��I��
0�$D��%�}\��'Cƨl�lDB� D� ;�ٻ~z�l��@�p��SP�1D���5f� �5��ŋU�&�)i1D����g�k���jVM?��`��:D�����Kd����6mל��F�#D��ˀN0T�r��ē0a���($D������^[R�a��|i��=D�ВBb* ۞%�5n��Bݐ�:D�����L�Z�>]*�a�<+�h��l<D��� �c��EV��"d��u<D�HK�oZ�4�j��7�ӏT� �ӏ:D��˱EB�e 
)�G�O�.+�x���;D���k��t_�0�!����v(� 6D��Ôa�r���1u}���i?D�� Z�o ,"�`���<@���D"O�yH���30�M�d]%Z1V̘�"O��CeK�� q����s$���"O�����L��P#&��/�@�"O���@��&��,TxF"O�Iq$.ɔ;B���$��-S�"O�p��N�W�ڈ��I��np�5"O01f�ȥ9�ܒSFF9Vj�:�O�]+a��<�8�pV�܇��0�)�O�B�I<�.� �ƨc9N0I׃D�LC�iUD!�� |Z��i7���KOt�	�'�L9��[�n-��"w� ?C�2 �'���x�k3B�J��:�0#�'@�T෨��LpP�{�%��:� ���'"T�j�=�J�����-2j�UH�'b�A9E�ǃI���T�_�Y��'Mj�q�Ƨ����CgSE8<y
�'��y�F��L ���֮w�<�C
�'B�ӷ�D1:-��	R�R n��d
�'�򩟡A}DP �ϙ�V8h	�'U< Fn9�J��O?��	�')���"�(*�<`���~��E�	�'>,;G�;`n�9a��$h�����'��{�*R�r^80�@)S6a��'G�p��]8��X@�H�'�:�!�'�Z12s�Bqðh��I*T'8���'oxMjA���~�����6���'�D�r��۲�qSskưj����'v��F/F3f}RE "�W]��k�'7Xl#�,  A����X?Jh��	�'��i�)D�hx�`۫Y�Ľ��'�D<bhˁ ���ǚz{��9�'�Bi�Wo��b��S��"`�0h�'̀zԢN�
4�{���
n�J� �'D����@C�f�Jx�G � g��r
�'��eXc�A�fHH�F�X�H�k�'�jI�$Q�q�XP��d��9�"OP�#�/F\Nd��%��Q��"Ol���h���aE�����"O�1�
�2b娄D/�(,�p0"O�)pUGK�x�6�:� �����@"Ov���I)g3�I�F��Mź8�"O��j6�/a�����X�8Y"O�ԓp��5I�H��gU.��7�'��	��HG{J?�v�Y((�<�W@Y?N���{qL!D����(�@ȲF�(�<����>D�d80��l��:�.3D6��p�9D�,�ҧ/N2��C�(� Q"C�*D��)3��?��XIADP�/w���& >D��s�B�DIcY�H�����!D�`�L��*��y�e̓%G��D*�F D��(�b����@��I�/N��г`�?D�ě�)TJ!��̀�Vn��0�>D��	� He�>��5"��]f�p%�:D��[uq8Bf�Vw�qY���,�yjԓ|ּ��0O�[�T�)AKH��y�eƖ^~��@Z"�E�5����yRI%lC����
������y��L�(u�u���� `�wO�=�yC�<J|LK�O~Zp�k�&͗�yB㕡'�0<2E�Z�W���G���yr
�D�E�5/�$ɖ`ь�yr���4�)�l\o"~	:�%��y`�*p)`E��g\*o���2� W��y
� �
���}�l�d�W 8�B5�w"O踱uN�"wJ 2pfV�I���Xf"O����˖0X�ָ�ϗ�{`�J�"O*� R�� ��y�c������"On�XRm���e���C�!��Ww�"�����;S��q3��[>�!�\CmJ�2�Tvp��e��:DK!�D@fN�C�#4d��Mڀ`K!��%j�q�c�W/"e4�*S�ړ��'d�٥�'d�Q>�<�X�s���h�(�( e��a!D]�<�j�{
���/A�oEi�o�s�<�7�M�$�ƍǎ: �� Ri�V�<!�a��>H��ș�O:����G�W�<�q�_����<������o�<��/�c��q�Y��($�D j�<!`%�	af$m����(V���φQ�<�d��
�0XbE�ͶJ0�Ū2+Q�<i�	�-��T#D-:�V�R��_L�<����I�(Qӵa�!kw��BK�<�0����i�b�$݄yʤ��<�%B$�$R"�R�q'�����u�<��iU	N{�tç]�PB�)�
g�<a��M Tr��:s�Aj�p�y���e�<�ы[�s���FcX>��ܹP�c�<������PC��2�p�F,J�<��Bv;�$�g�<4 k�UH�<)�`��!I��In��]n��P�Ak�<!��(n���b��"\j K0@�j�<Yj��k#ڡZD�R+0gvղ�Sh�<Ѳဴ.ޔ�`�̤r�<�z��e�<�P4@�N�Xэ^%��@J3J�<1LX�`4LIs
V���Q��EJ�<��9$k�(�AԆl	��B�<!SK�)�3U����E���G�T���xЮuPE��TR�1�@�N0Z��|cH���#]g�� 6F�.�x�ȓ۬���Bߪi�΍��(ąȓsZ�Qp����
<�ah�%�\��ȓH+8�3�+Q����,&9H5�ȓD���0��S�B� �A���ф�V�1�3(�� P�A�.Ά\,�M��w�0z� ߋ�\��v��)s�هȓ-�m*F-��Uʚ(��ŔF�25�ȓ��!��m6@A��� ����ȓ1�sFI&dz���G��K~��8U�T�ф�Y�$�+>��|�ȓn\�\8�g��Yg\Q�@��?_�~%�ȓ��Xp��8Dz���oL1] �Q���ƙJ7�NO�S�ײ�,�ȓ9���� ����i�.j#�\��h!lq�U��"���@-�u��q�ȓ-DLy��kW�4�BI��ɒ�B�`����aP��R8ZԼI�C3'q���ȓ$v���'�~+��1�j̚s��5�ȓ1��aQ�G�\99!��g�V)��hȞt�'H�{c>8����Z��ȓt�1����/��0�d\f�Ʌȓu���`�D�v�	�sI���d��8�ǎ��d,ة��H����&�ꓧ�T��(w/��}��U�ȓt� a"�!z~�mx3��6]� ��k(�r�U�������`�X�ȓeM���M�<�r��P12s�q�ȓmİP�2�߆@x��Ƙ!6q��S�? V����	�?���_"/z:{�"O�uᇨA�	���2�EP�]&C"OB�)6B �9��u�Ӫ�'{j��[�"O�@)��yt��GO,^�{"ORĹ�$�, ��(y�K-p�<�*O�P:�ʖ�_�.QHɕ_���
�'�#�g	�D���Cw�V��t4B�'��PI2	�
 r��Z����k��2�'���y�M	 _�e�u%Z��
�'-�q��ߵ[Av1b�>�xɡ�'tP�� �6�&Sp�U�O�8�	�'p�Q��N08�Th����G���	�'W���0cҺn@��!��7B�2�	�'�̭;傓:(��l���A�
���'/�1���#3z�(B�"ҟ}�~��' A�����1���GXȂq��'DtT�פ͇	�z����ӣ>x��'*b!��B��I8��	�68��'E�A�v&V�;�Ε�"F/�|��'�R�bk�<��|�n�%���Z�'�8,P�J�}�Ÿ4"Յ@�D�*�'ɖ�;G���"��W�����+:D���n]�h7 pD��5�6D���6D��
1N�:��(�k���6��2D���C��/ȊL�b��E5��s�-2D�$��8]��5�9T^�x��<D��2-�^�D�6�͉6G��V�'D��h��}���/� }9ԉp�F%D�t�fJU�
a�����ڡ�Ԝ�Ab6D��bA�����@�!k�Ab�5D�4�K��(��ZE!�.��C�?D��2�L18�rE��/��qe#D�����_�s��!�Ǒ� L8�s�"D�X�g��={cB�1�]*���( D��2�l��g�9���	�4�2�>D���m��n8|�Ao�f�ޔjsO/D����e��[~�J ��P��Dp� 8D������t
�MB��p���5D�|�v(ڳ	G�$�5ᒐ1��K��4D�(�V�АhV1зe�g-|�dh.D��XC� 2	�)�UM�M�8%�W�8D���Q�Y6$�x�C!I'ei��8D��b�!���D�lf=�w�5D�4a�k����x�J���2�[t�1D���և��Fh0�R�&�VAZ��3D��xw�ҁ�<�P��R8�~�(g#$D��i!6I|F��'��9X^8 k D�S�ݱ�L�yB
U5�tmj��?D�<��f�^��8����;%�:�B(D���u�Z��~ah�c)��Z�c'D��X葡 �R4G$-k�9z�!D���x��3�B����C�$D�,i�	Z�Bl��%�, ,��j>D�t�р��H����^�����0D����I7k������)�b� /D���b�	&gjؘ��+ 4<J��d�+D��1R��%zu����"�#���b3A6D����"_�(Z3��:U��RD�2D��I��%?���ŋ[��D�I
.D�d�f�Z�M� `�fN(?�ش�V�8D��Q��]�-pjɛ@C�'�0pVC7D�4	&#�5=f���i�_��tydb4D����L) T�!�W%[�<CT���0D��U�̦&�0x3��h�4Q)'o.D�� ��f)$gx`Ă�%��>���Z�"O�����}d`��*�jx��!f"O��F��.a���
e	r���B "O��(��=�0����Nu��"O�k�O�1`.�Lʕ��d
`� �"OP�@�&,�xH�E�	�v�Z"O�Ir4l׺j(L�A��NAъW"O�<YѦ��M�  �˝�q-hp�"Ot��R��%�tX`������A1"O�Dc&��c�᠑�ŕ/\,�A"O�����ÑP��h���� �4!��"O0h����g��0�WH�V���"O��R�'s츘�g��,�8��"O����[XZ�f�
3�.��E"O��y�)��̈R��2�\9�5"O�ţuS�"9�x�+��I�R�@"Ob0A��΃F.���a��5�Ĩ�A"O��TC��X(u�F�@� 	C"OF���/0���[ `��{-�v"Oj��� q��X^�*�h@�"Oܨ�`G:-��m��k�萈Q�"O��G*�����plݖ�,�C"O�$A1'�	x�e��jƱ\�v���"O����i�@}�I�l����d"O��H_�S�ʙ;ǭ�3�<���"OZ��I��-���@ME-� ���"O�Ӡ��7k�L��㐈r~���0"O�E� �]�+��R3L�-2C`M"OpyU�V���3�k A���"Ox�s��̩RGV��iH@��y`�"O��M��O�\Q�J�(��P�"O&�PP�'5�H VƄ�fQ��`f"O�=:A���U�=X�o\'WܕKc"Oՠ�j�~7R�(W��y���0"O��2roG�X,~���F���|�Ye"Ob}1�/[.b����\�dq�Șd"O<#����/kڌa5EL�q�p��"O,u�0��~�)��.��=c�"O�`0��O).U �Ɯ���hC5"O��9A�ɾ30ePO��b����"O����۹1*p�P�@%t&�k�"O�0(![=��1c�/<̳%"O1""b	�9���A͇1�r�c0"Ob�٥�N>��e�̙R�օ1`"O�arVNH�*�l�C���.5��"O|���4�lq{ �[y��v"O�2ӆ�-��-�Gj�??sr��G"O"�ñK�@e��g˗�J�ĉS�<�d!\�3D|��sN��m|R xV�K�<���u��Y�I#s��M�d�]�<9�+1jH����x�G�Y�<�$�� 2@���p�ɞ�f���o�<i�B͕4Ś5�G����[�,Fa�<A&�m{>r�o�;g�`���@X_�<A!.�!O@��bǘ�k���BJG\�<iv�ѲN3 	As��
>Kr��CJRa�<	dF?_�-ɴڅ0H��b���^�<�"�yAL���r���B���\�<!t&Y�4�(*T�a,�JS��V�<�7!ˉY]6���.E���e�A�z�<�u�ɴ2Z�b��{7����l�<�'� 9�n�����LU���-	A�<�Uޟ?�Zjd�1#i�$[�(Qz�<a��U;W���J��k�L�0&�M�<� HH����0���˰�X
L�P�;"O���QE��^ȐA�!V>'� \Z�"Ol-rWᛞx &�K��"�<�u"O�	�W#j�ƠZ��%8�l%9�"O�Y�������J6/X��lkU"O2`J�gǜk��� �ΉX{\h:"Ol�s���z�l�GlY�o,���"O�]6T!`�q���zŒ�p"O�`�A�F�@!$,3��F\Zh�"O�|�7�R ;�g�KA� ��"O�Q�g)�'��U����/:2y	�"O�}�C�';�f�PvB��7�E�"OJ�cbA�>ሄ�����B�zaz'"OʸY�M�q���㣭�;No��R"O�Q�X�|�����.o[��c$"Oq�hE4���Q�L�h�`X��"O$`W	B֢�X��K��9f"O$�Pq��5R�B�Ↄ�dD��CP"O�Q`!��<^�.-�� �'b���$"OʅP��E)9�����NŌ`�l%��"O�u1��G(9�&�A�M ]r�99V"O�����&+P0��Q�ܡ2bl��""Ot�CiM2�x�aJ��}���R"O� ���U�Y��iT�r�xU{D"OVAs!�3Ҝl�pC���H\X "Of�0��.\�fň�(ҵQ:���"Of\FF�4H.�Q�Z�\���z�"O H���;Fp�9�F�"z$P%+"O������7�(��פԟ6A�B"O�AQ%�/JPx��[�PF`��4"O�M�%iE�N?x��E�( ��7"O�ta��j�8�3�+%	ʤ0�"O�I�����H|�8��[�s���*�"O���F�ٲ�:JG$q� m�U"O�t8�,[O�P��Hԭ|��Y��"OHh	��@�0�5y�'U�<)z0��"O�8�@�(m�T@R���X#�,1"Op�C�D��)� ��a��
�ֈQ�"OP,�`�F%�ݘF�ۚ�(�"O2�աM|���Zqĝ7[����"O��YU�v��xX`�զ#w�4��"O�l�d/^'ew11vh@�!����"Oh�ȅg���xu�ߝh ��"O�� ���b�,q��h�h	#"O:�R�ѵ�� ǌ%��iæ"O���o�	��'+E'P��@�7"O�iea�^nV���̙s�t��"O^�:R��%:vab�
�(`�~)��"O�)(ō�I��� e�iA�L8A"O$��4oV�5jp��Z�Z,h��"O����iՌ-*�(p��L3|!��"OHPZ���C2� ��
Ai�x�"ON ��X����(�
r8b"O~��6�T@"��R�<K	�uq4"On�`�" 
x`ũ%gy��Ar "O�p���2n���c��+����"OD�#��6.����9�<���"O��r�I�j���]_�Э�d"O�	���pvr��`/�+�.�P�"OL�0v�T��(Į�?dب2"O��o�n�l����|�f�Q2"O�$�-�:nr�(��)w�H�zs"O���� �~�P��P1� M��"Or��P��i"�a٦Ǉ\|*�k�"O� !����p�k'�G%\oR���"O؍q�)�>��(�1"gtP��"O��lZr�t��@�W�d^N��"O�Ȥ�ơFE� �썫z�0U�`"O� j�L	��ˀ)T�rhXR"OL���9B�Z�0kҩ����"O�X��Qr
��UD�7�-�"O�#mQ�0Pdl	U�_���"O �B��Y�4�QĂ	?B����"O��!n��K2^����lAD"O"p�T��0AU(�1�JW���9&"Ox0y��"�ِVKG!q� ��"O�(8u�QC>R$Xvj;Kc���`"O���0FݯV���"w��Q69{�"O- .\�`(��8pgH=C�m!c"OVD�@a���ťi+NyZ�"O�	"��Թy@� �DmP��:h91"O�-�V˛w�.���b̼V��Y��"O��+E�]{O<PAӀ`�z#q"O���Ս�*}x�-��LIA"O�A�g�q)J��r�ͽ��	��"O����<�ҽ��W�V��`"O2����"�,��0�߶m1��w"O�E�#&;�p�pGc�:���"O�P�C۫`�fL�b��3)���*�"Ob�9�b��*�$J[��srIW!��ȏw.��e�i;\��͒9H!�d#nU ��ܽQ�rQB�<A!� 6c�X��L�=F�P�H�u�!�DZ1�,\z��Q�.���rL0P�!�ȂTnyC�E1n��Xi��0�!��Z+6�b]
��M&�B1 �G�<#�!��_7�	�VH�$!Ras��J�?�!��ڧe�|li3��c�$Mx�KMRg!�J&y~P�R�S/Tر��	�/�!��ءr9�c����2DpI���!�Č�'�$a��Kìn����U	�@�!�;�"\"�	$&�:`����$-�!�Ƈl��A��H>�����w�!�$��Pr����g�%/�	����!�D��x2�t8��S�x4�i��呬Zo!��΄i%����8��sE��)n!�dU>*e��*���f�B � ÷@\!�؛t}�	��	2^���d��9(!�$V����⅟�.�T|i�I+>!�%`�}�(�C�n����]�o�!�D��D�n� ��6.�t�B�����!�dS�C�p=j�(�V�(ݚ%��n�!�d%V�ћ��
-�TEC���.$t!�D0E��x�����z�� !J�^U!�D	�+6䄛��~�� �����'*ʡ��+
)_j	cE�{W�(!�'<u�._�bd4�q��"y�X��'����!X�f9��Fl�4���'J�)���X8�J���|�8	�'1aQ�OOC����Co��`��'CѓW!S�:���3�.5BJ���'9~����.^������? &YC�'���;�F��z��z#��(5���
�'�DmТ�P>x��9�⍍8Z�V��
�'�`�p|x\J��OO���x
�'\|�[TLҺ?��H	e��J5�E�
�'�HXJ�G�R��!��6F��l�	�'p6�#��֩k�>]�劚*?����	��� �Y��*��z�A��"T�<�"O��!��._�X�2HC�X ���"OlX�E�/k�*�	 �U�e?\|"O������O����$�,�M�"O�41$bT"K �	�*op`hq"O��@�?l�-���^2L��bD"O����Č�a�s�2H�r"OLa���ԃ2_*�����K�8+f���{#�)§Q5Z�+7̋�@d�(�aǝ��d�ȓH���xu'�) pd���K3����)&�LQf�ʱ!��|��Z�1F��ȓ*>���vc�.D3�p���[X�4)�ȓ�8�3�lP#1`��Dk�p���ȓ\!�l!���
r0���k�Fe���ȓU�&����J�ad.C��1�=��(����bţb~���V*�N�ȓh�����L3Tc&$�64��,v왨��[�Z��re�lD��Ii�'ώ(��P	A9ưy��|p ���'O�T[a���[Ϩ���-Y�
z� �
��Od��ׄ�Ჵ��O8NĘ*�"O�$�vO�as��X4�	U]28���d(|O�щ�N����a0(�`����H�'Y�y2�ҥX�����Ŗd����KU��yBl��je	�\��a�@Iܙ��>��O��H1	�%_@�����K&&D��' ўX#�^kw��8��;���:D��z`��]���Vc̮-K��5D������Z�#I:��\rկ?�	a}��S�,��5C0Y�>���(��5N�(�ǉ<D�P{��U�mL�J�� ���U�y��E{�����<y3D2C�����уTr��2a�l�<�&C��f�Ƶ��$�!I� ��Oy��'B�x	�K�M�ܐ�wI*%�9R	����7Pਉ+��U�| �s���B?!�D���T��{��qP���_��c����M~R)i!���O1ܴ����C!`��1}��'�dXӑ'K�/x�:�Ҿtx\9�{2m1�牾q�2����مDR4%�R�dC�BቶS��5e)Ǎ1�:���	�� �1��H��#�'k�`�%^�T�4-��O|]䩄�əxT������W,�g��+3� #D�K���;7����m@�J���e>����'hQ>�;Fc)�zU�Aa_(��\�=D�����I�R@��ҤD��_�P��;D��gdؖd�Z���T �9��!6D�9�T,8& �0��<g���p �O�YG{Zw^Q���s�C�l{iS��W����m'lOx�<���JWO.x֢1.m�����<1��\�&�n5��K�a<��jg�~�'�Q?��Ȉ��Y�'&н77:1a�$|�\�<A˓U{��
j��!�@%���^HŅȓ~�(Re�th�A��I	&x���b�8E�1�L,���Фm��$�ȓt�8���Q%�l�Pt�C�M4��H�<��@Ŭ&�d�@����مȓ~fh�!�ܼy�y�)�2H��ԅ�3�t�tȒZ|-Q���	� t�ȓ7�Q��C�gc��7��.y�.���=�bu3�HHl��i��Ϯ_H�ȓ~��0��Ed^9�%�29�ν�?	���~�H�Us:����f��7	�V�<�I�H�:���4��D���P�<�p"�2`���� �l̴���l�:e��m��fyb�&��� ��`r/A�R�^9+$ʅ't(��@"OKw
Յf�ȍkEN�#�Y@2"O�����1.�h�:&䃮$��l�"O����*��c�D�����o���[Q�I�hO�ɚ.X\���I�e�Qdl�47[!�$���4��OEV�E2�[�B!�*J"��J���7��X�H�+:!�Tc)�l�q��[$k甇!��D�.b��q�HҒ�?��	П�ˀ�$(�q�D�{���}� �q��=	 �ȓ'�B�f����Y�7n��<1���?]����f��X���˒!=ހ��&>D�(c���;9�����N�� �<D��X阓�T}���5R�|RF);Ⓝ�(�REB�
��;�V5u���<O���D#��,�ծփ!�Z� a[�)�!��@-*~,� (9m��0c��?n�!�D�>o���#GC� 5�F�U�Uu�D�>�I<�*O&�O�nّD����o�4	$��֯�8\!�ĝ��T���\�iPT-��d)�OΡ ք <A���H�O(ѸE�q��\�O�,���@�$Cf�P�E�gO@m!�'�#q�A�F�J���,J)�T��O�5K-OnӧH�̽K� �
o��Ѐу�=�Ib�"OD����=\HԐV�&n.������`����X!:��@���!Iĩ���#V�!�ę�8�p����ķ%���cG�*K��Im��(��|��ηM[�\ $��yqv�"O@$��n�2�d�u�+|Q$��<O��O��󤟯y�8Iq�?B�	 %�1}FaNk��W��/r34M[�"߀�Z�c�L'D�<0!,� o����a�X7$� ��`x�*�'��Ж��g̓\���!땯UU,�j0OFLm�ȓ��@S���(�O�
����'Aў�|� �;�j=��<����cZ�<�@)�1I��X�h	&]����'�⛶
VM���h +ޱf����3D�9t�L(8�n2���$p�b>�(c��b��v#��%o&�0��,D�py�ɩ��u�Ġ6�N=�`�)lOv�p��+�(Ӿ�b�k�4�h	e�3D���#K��-���Q)9Z<���$D���֢M3>/�vb�h``b�>D���G�?e���`�K�E�$Q7�'�D!�O��"BA�b�|RV�F=_���"�"O�x�Ŏ�:|	�2B�&���[�"O��i��4���.�3��U�#�i���s�ܕ�@��6M6�	��6K�<�C�"O@��@/����ȁ�tz��w"O��)�++2��% 'Ez��&�'R�'�F	pA�P%:-(ұ�9����O� ��c��C����>+�U��9�:ܤOf��Ę�#�2I`�HO?x�����)n!�V��R����I�*	y�쒱	�'s�Y�)�S(��p�w��@숱��v��C�I�G���h����+F��1�ZC�	�u�>�&+1ͬ�SC(�:X�#=���ҍ��-:�p	ԹF����'+>p�ΔH�t4�sF$x�4�b�'L�KϞA��1�+r�I�'qiS�)���E��x�豓��� ��O���O_��z�)�e��(�C(���'��ͳ�.�8g$L!�C�v�) �'���d��&X_H��t� �_���r�Id~","��q`��ȨG��y+@��y
� X��"f�dDhe)I>dX���Ixx�k����J�Y��Ϥ�2�B -D�Ps�Ќr����*��k�t#��,D��: +�R`~�9��J,j�xY�N+D�\b�HϾ
+���c�2j�<bD�+D�0(�$<(N���.��&�:
*D��#G��*+�0X�&�;h���"4D��R�gX6)*Y,���Q`.�(�!�d�)-��<�F�4��X��3.U!�$R R��i Ek�U��e�	�V!�J"k�.W
'���P��$/%�P��G����JR<	��r�c˜�ؠ���v�{�i� Y� @�Y�4���#E4H�� 3�Nɑ���\�J�ȓ9�i�E�G�� A��cZ:Gĭ��\B��
��S�Y�v�ZR�K,8@i�ȓB���aV4�6A*4���ɅȓI��8b�Ωe���Hw�	b L؅�:aJ�x2!O6u�X5�sT7z���8 �5�ؚo�d����f ��<a>�+��M�i�,��X~� /#D� q�İ?�
=�T4xވл"*O�<B��

4�6��Ƭ�0.�2f"O��S�Z�k%I0��3��3�"OB���b&*��R��W�=��rf"O�3�(ʗn�J�)���?@yܕ�t"O�<[��&p��т"#C�k�j�"O�*�Z�:rb��%_D�z�"O��D��9��*Q!ֆWzh��"O����>j,�DB!`�/\@�m��"O�M�rL��xM��� $a,\͛�"O"��c��_��؋���yl��W"OT��gC�)b:	;R���L
P"OlT#LO,R�(��G-��D� (��"O�`s1n۰,�`�&�-��	�"O"�#��Щ���5XVf� �F�!�$��WG �h��47�R��^�^L!�dD8gWZhrN�/wOj�`����!�$F�PJ������3\0f��@@�9!�dQW�)���B�
�\�@��W�*a~K���$�b$_&�kl�4T����+�yrO&U䠸�A\@ t4������y��܅W6VQ ��ʘt�>Yc���y�@�'�X�ig����gmE��y�h"�H!�TM
�d�@$n�y�F�f��ٸ�EU
	e���;�y��	p�Rq�0����HW�Ѻ�y"A$���2�Ћt�"�(�ܔ�y��U��a��l	k �����O��y��"Q����g�S(n:���@��y��3�d��6�^��U(�-��y�l��~�r�`LӼQ9�>�yb�US=.��㝕>�0�s��]��y�fWT�!�ħ`�$�҇���y�홤7��!�!3�vd�.��y�!	8�����گON�K��ţ�y�E�<|@P6���F[,y!Nb��'�`�be�GY/0��*V�yw�a��'��h��=G"9[S��A���"�'X�H��G� ��'J:��'�±��EJ�=�A؄z0*�'�܅��b�("	�Ib����(�'bFY��O�ɧh��	�OC�H�����Zt"O$��q�ޙ"x)w]C$T��tT�x��h�uF
�H%��Q�� �`ay��HF.O��a��'��=ѓ�ǿ2X��΄l�j8�P�����b�дI��H��I�x�DL)�g��qK�Ȣ��&���<i2�K&z�JP��3sO��J|�p�@
)�����%�Ai��S�<�C暲c�r�^�@ءЭ�<f�9�"3��� �τ��z�D��'�|%��f5(����n�>0�����'M���`&�;YvD�+0BB�?N� {��e䨻G�)0\�s��3M��E}2�Țw�6Я;��6b�,u�ޣ>!�����ܠ� �k&��g��#'gȱ D*��s~D+t��:b�8��D��F���#��'���ᥩ�S#j0�����6�=���^�n�"�ƃ>)N�HCmQ�_����u	W.U(~���I��+M& �QefD��r�iB�@7|!�D�W�0j�� c��ł��C�v�E1��! v�,`F��~�04X�^?1�C���l�h����Az?�t��S@
իDD�zK�E� �p�%�&l�e8��:�|!6	@�;J�@y�w�6(AT�$N���ʕtΐ�!�.B�B��}�4AI�lN�TEx��I+�L�+��B�e�VH�UeF�@�@�B�D?M* %�H�f�>E: ֫�_Rv`[tNȖ.oR�S`�x�����*Z�YCe�7|������'��㣃ÈQ����~B7�H�>�h�B�"�^�)BR�P�t�� �ӨG,A$�}�u��� �� ��ɡ;�|�
d\��s���'a�i�*�d� w4��*rl��L���'T��1斑ba�䈐�L�|���Tv>�i*�_�5���1$��>�N�x��%DJ���OM�h�s�Պs2�Ab�Dߝ0���!OQ�m��X:�2J�سe�;�Y��'���q �Ĝ)#����X>��At��8�ǟ!o���3�o״>��U��g��_�)�bL� �ba�#+�rH	ѳ*��� O�69��e�17O5��_;��X���U�8�R��\�r���,���pu��<�/S�0V8hj�CT�J���񵪖�[� C傤�]����g��ڑ�U�$ט�B ��%~�xX��,�^mC���M�1�a� ��-��<��G��h�5� 4J@%I���@x㓩LZ���Y�E�Q�d�iP,�;��XЕ+�#1BP5�?��3K�j]���g�y��΀%<k�4�ܴJ�) ,Q!*v�-��Gm��I@���	B�e�� �����w*�T�n�/m�BA�G잺"���4B��e���&n���Q�_�|��Y.i�Zu��"���$H�Z�`)&$T���UF7L`�qmڃ/Ā����  ��8�v�>+��)�b\��b��ڧ3����ʀZ�ذ�C<6d�j9>?�,@1aE�	R,�#񃁧�~��c	B�Ȁ��<8h�qj��=:���D1'��*�%^
$��	A�S�_�H R�.Y䭔'hx�L�:�L�7�	�qD��֪Ό�s�^= �ܣ�I�1uh�˒ᇗqd��3�@�?B�dC�G�/tl)'����䛚>2�i���2�k�}��i �
�4{丐�F� 2����k����(3��
;m>�]~��y0�*�9�@8�b`�v'���][���v�D"(����Y�F>�����)h"B�)�
t �������[V���2�N�����w�y������Y�a���rt+a���\�@A�$�	�9�2�Hp��	J����M�B!<��0�	�|�v @��܄H�һ
{���7���� ��L
w-(��H���q`ט�TLR'�/`�����IQ��X�o�
 �(��� +߲��$�
%�b�(����d�
9�"M�+OX��B�G	�0�B6�T�yM��a�&�-��Y���!\e����wn�'C����	;���Ո�*���c�+�uw��-zШ��2	ψiaX ��"��`�,̒���,����Ƅ"j!��Z�,�.|ܾ���)Ίjd^��;R��5VY��i�c�mQB)4�Z�Xs�ew< ���'r�A2B��u�O�������d�dK�+5RʈP0j��,�
k��
�V��U�	7���A�a�D%k۷Tǒ|S�'ɰ��S��;}�vx٥����L������O�nߖ &�k�h2u�Q��*c�@�p� _�<!��2�&�R� ��4X �Jf�1��$ݖ(R��1�B[ G����cC��HqOl�a��%�X�R�̂���N�*Zd: �
�/jT򡏉ns���J8�"e#��G���`��I�&肱������Y@�F�$\�]S.9|���(p�Ya�z�02EY��!3�������_�K� ϻL��r��A�-ۋ|j��ȓ?��E� e�G�=������K�'_��b�a\�4H(��	�?��Q��E��B��g��������B3d
�غ��&	X��>݆鉂mXFXۤ�L�n�|)� ��;=  C(ͼyaH�p��[W<�K1���5��쫗� �����Œ�7D{�%Q�j]���

�l5a�*̘'�j3�!�JW��6 l���� �׳Th���.l�v(���]2ƌi���)U�L��( �3Ď����~��˴- "hs`�B�V �����_�J�<�V#,/r�yP�ɲz��5�d��myr4��֟��.�!MNPa�=bf(��A@cV!�JG� �T��K�4qi� �4>��ѤdHMr����듕B��+c�[�H@���'IN�$mA� ����v�i���R�OT�*��4��N@�L�̑���^.t�@ݺRj�#8�D���)���RJ��`��~�\m(�W�Y��M�nگU�2]�+Vr�:M���ڶ��+�'t�zEH7҇]��yc1�	�k̼�#ǋ�b��ۖN������[�:s�$0�ˏ1m�L1�I�nǨ�CGK f��(�n`}TP��k�*�)���C���r�*��w�
p� �-ғ o �!"�{F�չ��`�	d4J�C�� 3Y��i�� D�
�J�(�U�5�  �ui4mP �@l�ɦ��gf�b�,��V́�@��!�p[~T�R�	;D�z�r�JE3��D�|�Z����NU��2��+���k�OG��^$�%��q}b��+��Wtn0!�C��̱�C��
�2�iU�7�x)�;|f萋Ts`(	�#�ܕ��Gvӆ���P՘�r2@ڷr��s�g٢	��1э�*#�a��Y2`q�꠫Нђ�Zb��6p��k�X ���;C����<�`^���)t�N�5OɈ�K�����(]�FO��{�1�7N����*;��d�v��=��J'CH�ړ��F٠w�j'��9��(?� �x�-�O��B˘ O�Y:f��A�^��5l_�X�̸�W�^$`@� �%ʓ@�V���,��^�Ԕ�租&fK� ����IXC�R5P!��3>�q�O؊n���X�n�֐=��~���F�YG�L8�2<�QX5O�m��̒��K�;Q�!sbjM60�f�PC�x¤�oh���q&_?�U��K3aFX��֦b��UÚ�&N<�����:h�HA.�3N�V\sڴwԦ�Rg�ډ �ƍ{�i�oG�P(�m��wҪ��f����	v	|y��&�*Ey�g�[D�g`V$����<���#�.%T��kӤ3�B��ph��;�n���w���s�ޤnLH�R-�M����q_=D#�e�v�6*��l��+�-�>Qb�5>�:t���V�$q�)Y0��p�ï�����H5Q���#�N<Pb��r�T5O����vy�ݙW	m�(�D��;p��4F���<YP)��s�!P��M$g�>� m�<!	ؔ����AA�F� +�
��A��J2��;�/��Cn����=  1��'��]d�Ѓ,��SL(bo�(���&�������lY�'M�)3ue�Ҧ�Y�@Ӯ���߱TZb0��KS���87'��B��P�iZ^
���υ��Mc� �5l2E�	0������p�x{�F�t�F�P�B�� Z�8�{�!Ĭnr�!K 7-(@<�˂�Nز�G�B�@�"��_� �+1!ŭmu��]�4&�"��M)*	�8�a�(#��AR3�L�rȤ�2���#���	�M%TuG�03�x�����1��"Շp�vC#�y��3�㎋N$^a87�17�l����iz�a�I�G�*�� �d���ܷ��I�ӓC0��ZN�}�<�Z��(P�XMc#�4:���B ��}	��jE/�45�X��!],���'�PEkC᭟h`&м h^����Z9mlA��Μ�`�lp��'�����M���9�KKs��G㋞I��0� hL�4��t�sFIe�"�ra"R�D"ڑ�h�Y�x��-*E���ųW�`��=�F�
�*գsĎ�l�6 g��Lb-�L��9@��VhS�p�X���*�/�8��T�\%@��=G�y%�܂:�>�1u�W!�
�c��U��9�s�ӟSez���'����Pb���b���5Dx�|��O$(��LP+}�	��G�|i���MS�o�Dz�t��H��3p����8zt�x䬉.;x���c�!Y���~;��ȥOȡT�6�+�Dk��ЪT�F�<�4�h�<PMpD�޴Z�����B�e��ɏ
�B��U	�o+j��;G'�]�Gc\,-9�岗�6#	>ć�I6"8�kD�_�y�!��.Ų�:âQ9$�^��q'F���aL[�0*�CRk�p�$A�J,ø�2��9&�R�ϓj$ţ�mY�o�T�+v��#�nxGzb�?7��E����5o!�!S�Iݓ@2��C�޹Ķ��f��e"@�ndn���,�h����aڷ#
�a��V8|̦#>q��ɩ�p8Rb±,�8���/w+�����G�#"( �pA�tE��2�b	��x,9�BC�	>� �D��t"��B,I�kfXЛ7�),�da`�C��$΀��6�=��>��N�S�]ZF�Ω������Dqa��%g𤊱݀�xP���X�a
�Ꭹ��-P@�F��·��ѩ��֥Y� 5h�a�ȂG��4I��⧂�)<�`��S�M!D5���A,]����҃��Ms���*B3��u�Q�RZlء�%r�L�J�#M�\�9��|>]��Z+$OР�i�b�J�GxB�t�n����6SB��eIҩ{���@ǯG#�0ԑ�#R#^���B�P*@b��:��~48��kH�'��j�F��v�$��g�IU��튕N�BKF(�-˜�nmI%�߬]���@d�E�Nئ�1�O�P������N�G@\Ӵmʞ �pUŭޗy5aZ# Ϡ�r@�K
�pI��$6���	!i����C�#@���2!�{~�!��@�1�J�Θ.,�Y���#l�6m��E��%�u%ÿ-��<�;� ��a�Q>�� +Ae��
���ɉ+��u�P։EDL"��N5�5K<A`���A��\�$��U�z���䗚0 dr@���H8���V�~Dn�QAC �`å	Ϋ&�2��Q�W�>F>����>�~��ăҞQF�I�5�[�Uv�P���J�n�>݉�g<q�~���*F�!i��.��Orh�kWl�{�rX���L���d�V�'�k'���,� ��V��axrѻVA�1t���2M�;m�l,Xg��n�SG�Hy���]7L3$��#����Q$�-��ٓN�P��B���C�x��<�O��8/ܡ`P<���B��`���*��'��5R��k�.��0�F�I���X�oݣd^>�F��?�p���:�����C]Y�t�!�Ed�d��'h��[�탥s���0p�)��<jU�w��Sa��n����W�tdWȘ�?\�  ����"�K�7s��k�S�Xş�@D\Pi��f}z��� �'�<5c��3*�>
�B�28̰�����0�˂�\�H88M��"��=�D��!�>�����/"�<���U�L�!���ɡM2���.������ �9d潠0�Ȏ�Pѱ�l�Zn��!_�y��`.��̤���8`�����I����5 �Lt�{S��-p���K�ިO򐹁�<5�I�"g�<�t�S�M����0n԰ݾ����үO�*��4�^�T%����.���o��H����0޴�� ��#% ��O�v�QQ��1]C�P�E�Wy��1`�x�G�k]LD�d*@�X�|�!�H��ɪ[!���AӁ.�f��H�Q�����*	 �B�֝d��<yա�)]*��@A@?�!��C���ǆ	�G��%�6O��$ ��O�1z�΁�}���S rh�3d� a�P��J����޾5*akQ/]uְ��t��y[�����5�ȅ ��˭O�:���>�ɰ��y���	G�qeKN;it�0��m��Y��КU�椫Ƨ�*�H1��OE�1�K�jq��r���
y���_�b���)�`��(ř�A�y_�i6ȝqO��g��t�@�)O�����/0s�
��󌈡>�Bp`E��Z�:�K'�A>8Ƙ0���E�PM������w��s���:�RPP�K�_�.�+�� <sQZ4b$n�gYb����+r9�'�n(�#� kbt�+�8)/=2g.�2.4��pp֟�MI�hаpA9��ޤ����R��)�9�`��q�Q��/!~���͐2	diq!j�������-�-o,y� �+W��.%�a��J��n����7�9s���B�&�
���ʺ?���͖�*�`u ��S�t�;��P�n'Z-�-ܿ!�`����(q��Fb#T���{rN��՞`в��j!P5�<��ѹn+�򲉀�t!A���f�F����#(�@	g���Dy�t֍��]�5��ɀ�u,8a��n�AŊG�y��tj'C�scE�O�����i�p?�j�AQ�wS1O�B�A�rXlm�t��9�~�8w�P-x�Լ@��U��p=��g��R����VN\a!A�H|�5�ǋ{�بDԔ�j�4��XЧo�I�? p����W.2h%#@�/N6=_��b��C)�U!"��z�hi�)C�"�ڑ���&����Ee�����+2>V� W$�
��c�^L梍js�ČuO�0@�;Ee�͙���+3=^�0'�@��Kt�i��E�D�&u��!��ݻ�pLڦjݕHG�t�g�EʉS��'h��4=�4�C��L�N������E��eF�qm�<t*A���yRqI��<Pr�yg&�D��q+�%�]�=�5��K:�(
bޢ�N�s�?S8.Y�D#�B%�=���3�j�[uC��K<�<"D���L� �	ֽQ> A�T�O�G�|¤�w茺���%���Z$-A�H���P�.�ɬ"q��cJ�9��$�S����8=�&�k��t�?n[H`%��oY�&��0@�X���T��)��p�"�L�3S��}9QP>����ޗ-~塱�̞P�����2}R#Q<�z����%1�pĻ"�Π:?��sj���I��-wpT�G�;SG��~��e�"Ǉ4y�<�$� ;�0 �'h=�'�y'�B�3�����d2G&ȓD�*6�V�^�Б��H��I�t�se�4Y�w>"�k�� F��2�K�O 쒣C�8FZ�BD,Щ������������d�r"�����-�e���!Wq*�3�O�a���j���K?�ɷ��=*U��s!|<���ʳLI��k���7*�ի���__�4��z���H��vm�Ū7�u���X7
�3.炅Y��[-{��O��I���{��Ah�H�0z2���ӏ�iIL�X�@G�n/�"?�M�|irXc"*F��ӣ�6=��		m������_6JB��?b�2��w�]���A��u�-Oڭ%c��K# �:O��|Za)�}kN|:�A>1����$IBe�<y�o��%L�(fC�`�t�!ä^`�i;֘qB0O�Թ�<Y�Rys�f\h%��"OP���e�,`&Ta�'L�)\���g"O޼�0�U��$�4�C�IH(���"O�ؐTĞ^��2^O�41�"O�9�`��~�(B@��?6 �1��"O�Š� ��三��$Т#H�{d"O�!�!j������ƀQ�Р�"O�Y2��� ][1A��r���Ȳ"O�;�េuD��ӀP�Z��T)w"O�`(�c��1v�₏�|y
���"O��`Dɒ��=�/��Xi �h�"O���U�E�J��d�ԨpX���"O|��k��g������&7����"O$S��R����:�B�E��Yg"O����֯O����S-Kp �"O�-*g˕2=J�p�#e�w~氰�"Om;7+�?8.�8��3!�ĀPS"OF �gI�h��ɛd#![�셻�"OV	k��>/�ֱ�3�E�2dj��"O||�a�V-0��v��~F����"O��x��%؊J�M�VO89�"O��آ��Ĝd�fLĿ;4���d"OpEYM�'M�y:�����( B"O�j�gP s�P�����:"�$�B�"O����-��p�@�4�ӚIDFPc�"O�KdĖ4%-2} �h�<XL����"O�u��� �o�6�"�Ve2���"O���E:xX���׿g��AXU"OxԂ P&5sP��!@����"Op�"�չGN�0+�$���f�"O@\�s�!!¹����C�$�s1"O|Q�O�/�eb�$íX,��"O�td�H�����C,	+��S�"O��3vK
��J�B9*~�5K�"O��S�h�<��[eH��Od��b"OZ� F�]e',!0�h�K>�dSA"Oz������iRH�v���"O��d��jF@�xAԝX,d��"O����D7��Q�b��"�"O:�)V�[�W��i��GM�h���"O$m�A���z�2=!�'��B�\4�"O0��c����b%�e����1"O�����#�$3s�9W��R�"O�`�f/Y	Q��M ��1��]"O��1�k�ik�� �"�\{���"O� j�Ғޥb����"���K9z�Bp"OYC��^"�pU��F
�Z4���O�(��Ҕ6S��O�>�R/ɚZ"I���J/S�f���� D�dA�ɝ	���x1�F�t��Ղ�<�c���ԙ��֋�0<��H�J���sV!�5G�)BJxX�|C Hr��%��*
؍�Jݕ\0�Q�o�P���'��� U���6���� j����
[���8%LR��<���4���e�%Bf�-0�)kP�ˎ$!��-j[ ���[X�u���>: �Ѻ�� �j�����L����)�矸a��M	R���[ߟE48���f:D��k#eƨZ+؍��˞�Ic��X�7Sf���"�=���a@��62��3�w�
p�@��]�0����@�A�F}����	�8U�=��Y���+q�\�u*�t�C� �Q���!���'^�29�p�1�O
y$%�V�f� �F�%5\6���'S6�p��ql�YnZ�y��5�������ȁ.�?Jh��!�֙����P�
t�2�ʊ�4�ȓ=@!�Q*N9f�B��GE�|�x��Գ���flU+9~N8���G��ܳe�@���"?R���3Y�49��J��x�N�8`N�qOB IB���O�Q�pÝ�d�<�xsń"<�VXz���$Yp h�MZ̦�@��O��t�J�g�U���*�j6�X!��XВ��3j�5ȶ��C�msl��%9�D��oub�ХX;�ՕM2l9���pڟ<rySh��m��ƨ=�h�Bv!�1�z�!���8 ��-Q�=x6�O�U�$̔�iP�PX� ?T��l�2.P4K�\}Ȧ%J�Q��S��ɗ.�q˄��lY�Lp�`Y�;r.A��Hb�Z�!D�	+X��4��oF� ��̠AHR��E�)������:=��|�G��$���`��K�;�主l�'|W�|���I�d��N�?��X��E&	���@��K!;��a���%
*ik6��`�h���X�8����#��%kƣ������$��L�{�44��G�-zqzq��Mn
ܒq,�^Y��j�K_uä@���0���I�w�����!��Mi̢�'^��Z�k_Z���ZC�VZ0�lX�'�L��&N��1#b���U�4*Uf�:p�ܰ�U�ÔO� ,�	#Qe��{��L�J�L��ĵa9<4��C�+.��ďA$r�BH3�c�=8���I!I�hJ7��6d3.��#z��]?��x��,���K�� k���vIYv�����$���i�.-��O�;[�ū��?睢6/��$k�M0�j�6W6 b۴2�j}2Pi�^G�I�ƪb���,L>A�K�5l�VA��wv]
	>��r N�ur��IA�'�4 ��@�� � �G���4iC�=���r|K�?�>%p@��(�*�A@���de��Ŧ�+��:���/jxf��``�?CR�ɋ^�����j�G�9�d��W"�[aˇ�5Zla�C�rI 1$�d�FC v@4(��س�v8A�EV�8a08p'��|@[w�>_&�Sj��jk u@pG�3v���'����T!@��Ρ�"ρ��Ot��b�Z�l����p��6E�$�S�H(e%���6j�
}�Hc$�Ү2s��Z�OjX�#�["�λT��-����(H�p�S1���|���A��z�Τ�d(��& ���S��y2̲l�b���D�v� y"f\�qT�4����[�L|Q�a%n�2'�O�d��΅p��&]!�y��̰<��Hi��Kv�R��qM���~�&J�$Z����h~"|�<�$*ԏlt:H���3�}���#6���S�{��Dcs�XO`�⒘i*����55�]�O\�Oלhm�	�rj�0�	�@N�-M�Ё���)��Ȩ�y��������6����r�J�"�:�,�oJ��!��ݒQ2��S���
Jl�10��pY�%M<qC �4两cb*�1�O���Ph�s������*��K�k����ibǩت(�J�� MP���=��'v�����j�;%0Ȑ�y\����8�,�I��J͈��Ȩ?�S�O^ �ԣ���xQ��I�+l��}�MDK6�H�V�:�����/ݕ5������vq�s	K�j��QI�'�h5Ư%�MH��pz�l�N���(��#�O�N�!��ؙC�K���&��8�X�x���]�¼T�5cc�I�d$P���-am�%#�s�'f�L��J�5* ��R�8 # Њ�{�Gܐd�	C��S�~�9��r�)Yq�מ6~<t�A�݂#l��!�X�H}�	�W/^�1ҁ&�O�ztfD�N+��A�2sg�%�f��CoV��4b��h( S�&�	o�7�M
�@�ɣB��d��[�l޽�s`Y���Bu��H�nЫ��?D�D��W�hn���&D�(&��ۥ�]w�`��F�=lcF����Z��E�H��lg����&E=,,���kğ���I%Dͪ��EC)
�Ĝ�2/!LO�|�¡UaiVA���Kb���# �>�)��OږS�-b�L<8
� �#	��A���� ��ܣ��+�;(b�(ãN���ۀ�@����<ɰI�����SB�6;�sH������NY�>%x�����!(z��d�Э664�0�$�9Ie�Y��8I7a}lD?�}��/�JG6�91�҃w�R�+��4.�Ě�DR�:��D=�A�R�ʯON&�!��y�-U�(c�E��@Q�=;PD���y�NP���m����=i'lh'J�i���1I����&���p�p�Іn8��A�p]?l/xP�
V�o�7��kdT�S	B!���7"�5��8�fE;�"�⌜�|"�H�Hs�A�e��C��A]N�I��xc��"��;c&:���"_$Q�>��&�/���{���{#�qr��~l�#=e(]�]iF�� �)V�$tXd@�#P��1ۅFD��.�ru�G�J�Hܱ_oJܘ���*Q�4P 4�
!U����hW�yv ���ɛgS@T��jȥ�l�����
���l����2+% qIeD�>A���x�N���;*�r:���%f�|0+ć��H�&�����v�R|*f	F�Es�)�'r\��zn��J�>�XֈNo^�)۱ŠA��,�\�J�O�:�x��I��l	P*��[0��YȰ́7^�L��Ơ��t�
�
��y��Ṓ$��c�j���*V�0�����/G�BnW��r�"��\!z���҄ �g�~���t�? lDX1d��Pa^�Rѥbi�Đe�G�K�(K���$� A�FM^�|Xhq0QeT�)��$`n���U��G��BQ蒡k��ɠd�d f�[.�:9����HB�ؓ�e�����3ʓ���["����[�D֐t_��9N<#0���ql��BFz9!'�"��{�c^���1;D��O��)���$<�I�'�"$�����
I@y���g{�<Ja�1�%��c�
BlW�ap81)U�Ɔd��Q���E
~L����̓�UX|H �)Y'/�T����z�4Q�%Ǆ`��aҒ��|J�١P�R�V\2  ��Z�0���G�+I�E�P�x��ϥT�"�����jMY���$Z��d���-$p(0�3:`�j�X �<��HR3v�")�4Z�B�ABfAj�Ζ%l`��U,E� �Ӥg�n�I�3��Z��;4��{6)�6��%���(3 �г�˹b��8�\�;��js��>8��3���4���nY,�$��I�:fg~9�E���o��=���j�֝�[tݫêۿlNQ��c�k��^<�i+ @��P��t��{��]���ڷ
`�0-O������n�0�E�T��M��^�2��2OP�'�hY�w�N&?���!�xX�Ԫr/Htd)b#ɶtR�9�I�#��сU489$���Ek�2`I�jʓrBe���y�\��v�#��8��;<*���O��m�&@qR-�:=���E�&(j CΖ���5NX�8/pϾ�'�F�{	��cC$�e���j�9q""%��E�4!(��	�yۜ��
��ё��|�&�$[R�Fi"	J�lJD�-2扯TH�L��lZ�3E
Ay���-o�<�
$J�Mľ�Z�����(�-WN�X�L�-6Ii1qL]�l�2�K1i~��샅�+=Ujѱq��0MƮ�)�[^�h��3֝��<!&V�▋v��YZ�U�3F�+Ys�,/��V'\�!@;ba¤�e���7�+�M���bgĠ�S@Z�Wʰ!Q"�Z#c0&�p�'�z��,�B-Ѱj�S�ܝ���IGl�!�8�����9�~�Kv�u�1)�.ê~����͇�<),�"��d̝j8�{�O�c�E�GD�4l�`���ڌ_�U ��DF/�,�P�h�?'��ACE��v�`�j0삈V�$���.T�� ��o��Ȁ�F)��6��U�I��e;�D����0��R�9u��%h̅M 
ew�v�6�s\�S��@�tb�p���h)��9t� 0<��<+7�E�0ᇋ�BnPU����Y+N9@e�Y�`�	��4	?,h����T�axBD�LB	��؊��i0�� ��dȝ�Z� F�,|����9ش��u80� mFЀ�D-V�7f��z�j����7A�T�d�kC�+\O��QpjU5X�؈���#)�����H�L9j0ze!�	��-��M8�M��	GG�4\
���GV��!7��N�x�Xt���CG��Ű�Ä��9+���X��Y]x��H����u�ੱ�d�c���˘,u����ℙl@�z�P�y���bgjϠ8-F��v$��e�9��kX�u����"D�<BE�+b�}� ��v`q��7mϑ�lkʽU�>���A��]6���c�7f@��S��V8�X�p�5Zp\�z3n�^�n9�3�Ԋ$��U�e'E�3��=ٕhV��Ol��P��nR���t
�yF�-�3�ƚ	��V��9L�0�񷄛�;I|��`�o!s�Y:K�4��焚#?Fb���a�A���(ΐS����$�	<RhR
�����ĕk�|4Hu!�9 "D�s \�PFF]��V�k�B �:�1 %��h�l,E��	!����Z�w��@�dJ0�x����
��^_�D�w���gt�-؂�()�興�NG���p"*��/���R�i���s�XN^=�%� T^z�A�m\�>���a��mRb!��4f��O.J��L�O��AC�$b� �Y��)a%����)Cl��#n2@:֯����aǀK����+C'g�TJ���<Jh$ش���"hZO*ړ2ϼ�Ku��=��!��gӪ�ְ:�l�PMZ���Y+t&�R�L(7Ŭ�cEdē9���2R��ΌJS���F\�e��A2$���E�&� ��ؤK���Dndxc���=��yD�ۈu6�� 4��4��|��+�Dв�Xw#@d|Ho�	~fY�蛵�x̉�w�^�Y�jG.��q��D&B�x�'%�4p����g"Ęi�.�$�}��?1�M��FK�e��M�Pa6<^"u����c��9.^��I�cӕ=2�Q�`&
�?�3�[�8v\,qFn4s�H� ]a�'��G�5S}�� B�ݒl(�Ɇ� �AwNeS��"�<����g�TIq��1j���Go|�\�9ƁJ���<�v����O�h৉�Q� C���
M0���|�6�X��2��� 3-��H��IÌS��( L��H�	$w�T�"&��9~(�c�僯j[�-y��� �O
4��jؖHB� �N��t����A�O��E�A��U��X����)V�D*JD�H5. p���5ﺥ���U#\��!�,S!>���'�|��SΘm.&0˗� +G��!�"v�r$I� �z��d)^# _�W����ǾH%��В*O א&.
�]������;E��ٵ%�J�B0ӕ�$%Y"���Ĉ����9�MϬ)y`x���X�H�N���A�X�M����$KJ�yr�W�{t=�Uڇ!�}�0D�&%|�>�gW�W��2�ĺ�vCBe';��b�`�.c�D�C�0 ])!"�Y�P��rv�D;�x{�%В!6��2u�ɱe�i��KӤ8�.U���ՁZ��q��&�<Y�sO�X�'�t�j�e[	x8�$�@$��t�R)V�#V��HQ��MH H�a.·(�b�2EZ|4�� %��\��w:l�%MCN�TST*�.\�*O:1Ja��([_<�Xu
��H�p<��+�P�Fyx�nV�ie`��揕$3��U���t�f���Ɨj�N�qb#Z�U�\M wohv�F����~rF�q�����@���<s�Noj�8ǫ���8�&Y@x��̧^L��C���Da�Q4�K�69X�+�G,�D�x�G-�b�P0c��n��H��ARn�/W�6L�xq��J�S'V��1�Ӛb�͛�eV�Q#~$��-` ,�y���>zZjQ8E↠J���R�0����w�WU$t<����.f:�9�͌uft�+˻J4=��)��`�F!��➴0�XR�e�!�Ȧ4鮌@��ƻp�
�Վ"��� ��߼- �26+;J�xnN�����b��,b`�B��Ԍ&��@�+�</2�j�a��G��gA#2��Q���H�+�"�O�1Ս��jK�i! �(!p�`$QS�"��F�?y���>xU|�b��G9A��t��e�HR�뷅�/vXz�k$��k^>D��@��|\h�2'冸B��X�F�BM	\���4Z�
̰䬆�kl���Ԩ�f,��թ�I�n��F�I�V� �a�{bfC@�5tjtTJ����� '� �QX��֜bx�;��Y�yh��q]�BJf�i'�!�121痪��u�V]̓��iXT�R#I�@��vA�R�X�v�Q�gG0��nE,j��(���.m� iVDS!L�D���P�^�]5F�5���ҹ[b����^�W����m�>������;��a��ϻ ��1E���&ã���^gꘫ��TO���hf M�1}�u��IM4P��4j�b�T[��ږ��͘�C�J�����L�4u�i��[�O1Z���A��C��k�v@k%��J}��d��|�C)U^d���Y�0&l��X>���Oh����%F�PY��i���8j�Ehg
K-=Pr�{e�[�AB���&Nw�����E�9Q[��I��i�QHW��즅
!�*A@*V�ع!��}�"�I*���J@� �gޔ�Sr/ܗ+�OĨ3W��:+R�	!E�\y_�x�������V��XM�7e���� �ެz�~- Q�T�{[�t)��K=,A��1�i�D(n8�$׊)��p�JS�yiĂ-E|��2���������G/n<�r��	.��)�
�T�
�`���#dk���n��TyN��M3*z�F@��'���1���:O#Z�)5"�v0�(�dȀ&G�$�)�ϊ0���cD@�k�D"T�S�� ��L?G��6h@&�u�ƕ=/�l(���E��dN	|��v��`���f����IY'�X+��M(����@��-q�6���ʹ��ʧp���Q��G�pD捷f����|�LA���Dc�`C�J!�H��݁26��`�B�xzP3�$9 ۴ΊA�O�o�� �3�gӱ�����cq�A�t��+�d+`�H�P����aM�L%���B�0 ��@)��X����3�,���q.���:�j�B.3eZM�R��p?)���b�iS�*��'8�j���-��	�B���`%��C�hDnx��a�/+�~``�)6lO0�%EV� |`�f��]S}��!�;S��̹sb@�4i`��M>�c"��5hb��%P�Z�O���h�pC�=Z���8�X�q���\�D/V�3�Nѓy�&�O��� tl �7����	m߼Q0�'�.����&Y��6 7줙+Of &��aPԸK��|��ޯ	tq�͉G!8(���@�<yv��(.���(A��t�����~��[B�?O��h���,�cd!V>b����"O|�YŤ>
$�R�Шp$p���"O,̸���	���s��W3��2"O��+g)�?22	�ƣ�.���"O���c�ņ\r��a�w�6q�"ORaj��R���z�!ɋ ��p�""O��Ђ]�F0aٴ�=#$�p"O�kr
ܕJ��eà�T+ D"O�tr"��f�\�Qh�E>����"O<Q�j'.Ŷph�I?&�5"O���1�F�3)�#-Y�:��s"Of����T�#�X���.=��ժ�"Oj��;S���@C��m5J|�"O��i�J��P$zx��I�j�����"OMH'_�&\,ʳGЇa�^�SC"O�Ez��2/�>�0dGE�t�쬸"O��q�bR�@\<��c�-"NmYf"OZm��"��a�v��D/�!�"OA�n�<P���۹-�Н��"O��Z�kAeH�,�U�ȁ0"Oz8Ss,R�7H:��␧U`&���"O��EfΠ$zz[�C��
g��3�"OZ�XKٻ��Tsc!�8Aa���7"O¸���,�>yxWꇴN@�D��"O�0� GH�h��]Zw*C�>+��r�'��=�e��?|��4
Ǆ��4R� V�����{b'P�|���賌$��bj��>MA��B����vA�6Gpvxٕf��J.��0�i�,��Gqt|хF/�.�eJ%LԔi�v��1g)�X�3�i�2U[���!6uJ�0��X>�±lF�-/hq�F��N�t���K��d �⢆Q���W>p��X�>ĚbEčh\ӧAˁ����O�6m?�S�Ӭ��$Ho�(b:@��@$'j�Ov(������3w��4ڄ�M�yF�A��
w���$mQ�"}*4�]Y#����������鈴�2�)�S��]�u�G�T�JY��7vx�2�n�^fz�@M��0ç�0���f�u�|��9B�@��.�+
i��P�>O
�+t Nd>Y!��X4�Z��P�����1ULЕB��aH�'�~�x`O]�S�e����/[1/*\�C�6DX� ��K�����Ł���Ӓ0Pͻ���1n��s�CŵD�)�#�<K��'�6�G��tjïÑr��H9e;E�p�b�"�>6�8!�'P����\�h��g}J?��w�7��t8p��f5k�ϝo�Y̘�{çes�xBR�ݔjK:��ߩfp��'�貶�)�y"Gϧ$$�>�  u[��)�9A@Lɽ3�0�u�OJ}�'��O��R� %�d}��ʯ$��(qF�/G��ļ���P�x��	�� ~� �E�<	x�R����M���I71�$��)]�:.�v��'�Z`2���B#��'����i���<�|�#a�(Q�G^9�а�RF~�,���(S��ӻjj.q�r$H�U舛5!?I�Z�I7�?Q��.�)�'Os�3�UI`.}Q�!����$�'�Z��'+��O��qB�W"_�\�	��	._d��3M���~��<�2�����/�?��$WH��5�L(��[?,����1l��B䉉{1zݒ�'��X�\�c�MA�΅8D�|j�J�	I��0�&Ɍk�p��6D�yUbpB��
D�w��qi�,(D� �A�4���k�M�$g��X� �!D��dΈ.J���a�Y�>@�";D�+�)OL��%��<+JD��c8D���@I��M��X_iV�K[�B�.Hr���cF� V̓���q�B�I�T�z�J�9E��1�#7#6C��+D�ACrΟ17�z5;��T.PKXB�ɳ���20B�X��80�E�96W�B䉵@w�T��Ϸ�K@��*,�B��C�E�V)�!V�^��!+@1�B�I� D� �%��ژEZ"��0q�B�I
U()S��ޤ4�b�:��U5JdB��7h]���f,Y��Y5M�790�C�ɍ{�DPa3lI�={C�E'�FC�5`l���hB2h
J�2U�Ǉ+�~C�	���)IW�J�;;8��F�Èx�rC�I<%��8�O�
�����/ �YE C�ru��n�. �\I`�^|��B䉠O։�It�D�����=V�B�ɢ#jL�x�c'~HB)� �P1'��B�	
]� )b%�~N�-{p�n	�E"OB=���?��� ��{XfE�`"O
��C�(Iz�%�%VU<ِ "O�\���E:���m�9���ߚM%!�dV6����פكw�@��� !��S�9R
 RƈB8j�>���B9#!�d(d�!IfAP>n�t�8�[ |�!���
������& �!�ĺ\�!�DU�+4�yR�M�F�Х�A��!�$#P���kU� �4�ǹr�!�ę;�>L!/]�B%�HZt��-`'!�3N�F���L2wpx�	���=!�d�7 Zr�¤@�X�q�DC+|�!�ƧQ6X�� ȉ5s����� �"e�!�ŲB����V��^s2DQp�I�{�!�$�=,Ph��o�
Cv���O��Py���/?2*M�5��j-��V �y�L�_�:Xk�"Ƞg�,��)J��y��ޠ!h�D��G6d��9f�2�y�΃���i4�X��b��S�yb��C�Q�ϑ�&Np��tn��y�	���)��%�:�z�e��y�o
	��-c���"^���6���yb�^�nN�H$��9ژ pF��3�y��\�E`z�K ��9�E��yRˁ�D�-A2$X2��MK,�y��Xy����]��"e��CK��y�S� &���Cd�-{�$E9�����yReJ5���g^,���.�yR�X�D5�0ꕧ_=_|�-�f#Ď�y2�E�'����"�]��M�`���y��x{���jI*!� �@�(_8�y
� v�s�lY$r��h�ۍ+R�}3�"O��A)�&J
T�� .l�Z��"O��A�	� ��@S�@θw`<�C"O,`Qp�#t���� \ju!�"OD��6�� F���ÅW��(J"O�@Z �u�T��\�,|�(�w'�@�<���
!�:1�UAҡ.Dx�8�BTy�<a^vj�]1��Þ4'�Ȁ��s�<�d�U>_=$ͫ�&�	�`�S�� s�<q ���_>�u['Hˠ|*U��J�<��d� �x���HY�s��p���F�<��ˀuۀ���7@@�ӄ��\�<s�D�_L�IѦ<}���s F]V�<I�.ϔ8`>Dk�DVn���oP�<a���� 1��D=\�D*H�<!Q"z��l��N�/����LGC�<a���0�.Q�ҬL5��<��%B�<����������ArݫƁS|�<�b�֞)����v$�"w�<�O	=z؄��J>)���M�<��ǁ8^��[�:F�$D�əc�<!qd��?��e��)�+_{D}q�)�\�<���[�gl���F�ƥf(��щ@B�<� ����v������[� ԇ�!����v�F3f�����싖=
�ȓ`	>����	�!�$�P>q����ȓD��E����a�ܝu�ǷMAع��%I��Ѓ���|���(�S~d��	�*M�
�#�t��'��&B��L��Dޔ�"O�~�ĕ���L��t��ȓM��к�,E��,�R`�1�V���YvnH�«��+��y���K����\�pqruN1��1&�	;4�b��ȓ^!��O�2Ԥ� ���8 ������� �@�zt�# �*���ȓ'Ah�i�%ٮ� ��3R���ȓydl�B�� >�%�7�U�rp9�ȓ b����н8��L�B��o?�%��<�V���'�'U0�顉
v��Նȓ �v��Ë2�P�GR	v�<t��D��Ɩ/َ�)P̕��68��r�t͉��rB�� ��[q(��^�~=���^'i���V��2V�L����h9��g0-�H|*C�P�L�(���\tp����<�����0F ����L�Ѷ(��)��`�0�W�7���ȓu� ��Q/ެc�`�:5��@J���}e�A�?L���fR�-\tՄ� �x��7-�/d�V,R�N)G��e�ȓS T��nJ?m��!*p��(��Y��v�V�i��Ƿ	�3F>Aw@=��8"��$���hQ��)�:�v��ȓr8�t1�i�/�����h�<~m����T�Zy�����Z��1��N�8�Fm�ʓt ��z�.ǝ{F�S�R�B�	_N��[afJ�S�n�!���=~"�C�ɴ%���Ň<B",ɱ���hB����*��̲X�m��bZ5M�C�	+>�lhR��
<� ��ֽsQ(B��-c=�U( ��D\�s�%V�{�$B䉩Iid��1z4P��կ2~�C�	�}^��GhM@�\�`�b���C�	�:X&H`�@;
>��g�+r�RC�*>��2g�*�rh�P 
�o�C�)� R�i"�U�qf&��G�ZFB�T"O�M����"M>�]��.ЧU\24�T"O
m(7F@�Vf��ٴ�JK^�p;a"O��1���*�hV��?hځ3"O#�%�p̮(Ha8P>���"OD�t���
��1���S�&7L�2�"OP�K��U���RĮH���"O����>��Ӏ��(T(v��"O 	�`��e��7"D4�b(�"O�uʠ�D?�HR�K�<l��2"Ox�BE*Ǆ
Мa��e>�Mas"OJ,�2$�Т=����-K�L���"O^�x�"D����5�\(s��q�"Oj��
����D�;FӆD@U"O��ҕN�,�b�ʟ �,1�"Oh��Y36���!ULJ6\$����"Oؠ��1FE�T��5K����"O����I]p?���L���"Oj��)��M��+ʘ0�*p��"O��*��a݄ѭ�9����ƔL�<�wKP�Tn���V�Ɠp��r��I�<ɴ�3b��A�tg�BV0��C�<Yc���Fj�������B}�<9c�'��iz�3oh	qÕP�<���:q�l`yP���?'�T���V�<���`���8���<��zd�ZP�<�&�w3aER	>��V�a�<�c��r���f��o݀d3c)�^�<�D��U}8��n�@��\���`�<�a��y�X5����Y͠�V.�a�<��K�+ �6u	�N��e��jJa�<�$f�k�Zq�A�E�$H� �Q�<	�=: �FCP�30ɳ��S�<��H�2T�23"\|K�)(�^B�I[����@&@�
�I�F�M�h9�C�I� �W�ճX�h
�Y��C�I�Έ9��Ҁ]�a]�V�bC䉴)h�51��#e�Z�y3ꛨ:�\C�4dX� ���&<mVa�!H�S�zB�	�sѾK�a[T���*EdB�I�A"5#r���`�D� R��&>JB�I�ob��F�W�|8��ٯZ4B�	�h?p4*�M-��ɗj�XB�ɑ+f�$ң�$��0f�f�*B䉍G8@UKӄA��V�J�A��;��C�I�/k&1�&��1S�>|�BhZ&��C�	�s�j����O*��u�5���6B�I9���!	1Q.�%�5� >H�.B�	+LXЍ��h�^.֥I��ы�VC�Ig�Lb0�_���Aq&�s4"C�I��a��M]<2��h0�H >y�B��!3DY ��T.���tlמK"�B�ɚ%��s�	�#�d�A�K!,��B�!KҊ-"�A�+� ��A��e��B�W-*��H3Y�Θ1�d��E��B�	�+��xr��-u9k�F&a� B�	�	�` J�j��+!��"RĄ=��C��Y0�L3��?:E��� $Ā<�\C�I5[ވ�Vo�K�!�T+���<C�I�;lLI��&<����� ?a�C�I.�J�2Hé<�p�ǀjb�C䉦J�RB�$3�Rmѓ�]?-&�B�ɾyÚɉ�掃L�4��G^�aW�B�I%I���ڑ��	SK8U2�e��B�)� P �G�-W�ҝ �Uj�Y�"O}Q�Ɋ!4� �J���
JC0Q"O G��&��8Q$o�\$�Ya"O���Fm:<!�U����bi�M��"O��:���YnQ�R�X%3"O�`;4� -���R0lD�3h��"O��W�ּ.���5@B�E0��q�"O���T�X�02�@�0���i�"OR��p�P.�!sJ��4�"O�ĒA��? ����� DF�^�2"O$���̹m�=��J��r	��"O�p�q ��a�
.YN\EQ"O�9#+��k��@d(�XZ�%�"Oj�(C   �Sf�
�FY+Na��I./�$Ȃ�0O��
�J�X��QfL1_����6��6ܸ�'T+f�4�5�٪m��s�
�u^��ц�^����jOi��3�� �s��"܀CÌ�:|n&�QF�A'Xr��x�b�t��c�dA�rk����a+���S�ƌrc��a H�U�.`00BD:>�t�H�� ���I��<	KV��~��� �7	����Y1&�~����mxI�P�?>��=K�+	�h��F`W5��ś��0#�l����nLD�!����÷ A���?�cU�(��ca��
<�4 �h�1����A	:�������i@�(��3�I�5�pP�ܾ4��ʒ��;U��i{R��03"dBWnPe �ቓ{@T�فa��w���� Ȩg�9(�@��o0���mK�2
t(l��i�F�,{Ӯ�ѐ��E��h��j>٪�*�Ʌ<�:)s7K\U�� 
.�M+�'��qd$]%�F����&a�v�+"�@F�}Q2)�rPQJ!�$a�����v�d������P���(M��A�.\O|y0����)C�X2"� 0ʍ�a,W�p�H�B$� &+� ���rYxG�@7-I�%0�Bⅵ24���Xc�����P�$�Ɛ����28u��dX�zAd�3��I��`�4*�(�69�������3��B��B s��X��*n��-�.N�c�:���7:����F�1��V��!9��4����r��ٕ?�6H"��.H`���!k�T?��Yv\5S�L
C0��A�2$���Z�"� 7>��t�+>L�2"X�v(�=3�;M:R�:A�U�!���<� �����*��BB*��p�����9O��ra�&�ج�/��>��ͫ"o^�.���
u�����	�+�txؓ���Du���E�"&����F�;(4���Z�8"=��aq��i�c ��@�-Y2
P��Yd��bn��Z`� �W׆	��匞@-�d@Vf� ��h��Y0[��1��ak��B`� Tx�Jq��!h��6AL�^V����J0!�(А�E�@6��~�Y8��9��E�N/p130��<Ј���,ܣYR����b�2 BV���f�x [��V;�$��e��Q��N�x<�P�'��,����
�;x�\��GË{���*��M{�4T.���O�v�J���F�B�ab��x��Cђ2Ъ�d"?$v���

0CM�)D-�T��"�z��L�P�1��'�H���ޝ@�4)�6U�Bժ�ĻiF��Q�@7�j@c�(T,9�Z�ۖ_�@�$!cǷP�P�cI�l��ـS��p��yBG�E��E
[����t��YH2�$D�qO((�3��T�8�yN�3�p�!0��\�Ru��΅�=�$P3�� �����T�m�N0���C�4�d� ��Z�LM�6�ă8�0tQc�>@�B��'ʥ葃ɶ{N�uQ���	6yI�]1 �Ų/�n\Q����<�p���<D+��I���1*q�ۜ;t�Ux&���7Ƅh9Y%�L�&�Νe����M�"[Hh��D�k{��9&!�j���	^V��4��1n2@YI���*5���@ԸKN�4�V�T5��YZ��ԟ��I�䕛�@@�§H�V���S����&��hs�@�Ј�p�BKj�	���B�S͒� ��O&����F�|`��*��-/���k`��.xvt�����6�n���_9� �◧�-zm��zc�G-/��{p��xv�u9��˗_���`(��=� !$��T�u�m�h�,8�(�<���í0� A��'�Xq�)�#,��z�g�d"�k��H�E����NK.Ct�uBF�=�@y� -��B�%c*
�1�IF���J�oڎ:|��c'�RP-0 @���hܓ�c�MU0{�x��3�]�*�ƬQ���p�J1��k��'Ò.N����m��eȆ%��ԏr1*�r$
>�"D&�١(�P�HGcR.O�ȋ�Mödˎ1��J]Rđ��DN0`p����<������ŝ*=@�Dc��nzV�C�
�	LQF���A�S���Ձ�u3*�b`�BQz��vc�\���C�� � �@�+k=�D����2t0,�z@��S�'��q��՜P.��h�+Эy��C��I�qCD�y5bȋ�
ъׯ�������R+��H�됭y��k a�t�i�R���d�H���}q	�*��*]�*�@�P�V �7�
!�� 
�e� HT<�0/K<[�h$�N7m��a���S�!����	���l�f��>�7e.J>�4��Ǜ6h�Ip�)�z��!�wl�lV]��C����鉄N��3&�iRMm��h.p�a�;f������ڶe�x��G!��]�A�<�юBq�;6���c�"���-�d�O��#p�ё^"X�p�B;bS��{R��*�F�[�nـ���D����!H,��	�CN����0�mQ=;<����]8� lZ�ľ!�W��|�+�hk� �kߟs�4�p���6�8��������1�'o
�E��O���t���������]�T����Le|lb`
��.z����	�?�Ʃ��в-��y֡õ�7MX�tǺr��0:�8���äVM���[�SŬ\���{B�J5p��$ ���)D�� p�����8�MZ�(6D����J��p:���c_���b�:�,G����j1�EQ �ʓ��)c7ҵ��&���T��@��li�NiC4=����oM��1���sD�A8�I%��5$P��/tzm�r�[��Iv�B:DT�ȓY��Qa˂ *�HY,U ��=�ȓ���������V!���G�6cq�ȓi��k�(T� �Dgm؝� ��?��1���ܺ#+@M��/Z|�Ұ�ȓ	V�ٺ����8��F�]>)�ȓGT������5)��1	�ͺ-^���ȓr��C���r6=�P��l�ҝ��Ov�hPaF=�̩ �씬rr0��[8�P�bc�2@�	����~p@م�E��H�q�P�A	lq�cސ
�)��G�*�"e�E1 ��/Ύ�R܄ȓ|hH@� s�R��t��81:a�ȓ�f	���� $���Ȉ��l�ȓv׆ђEIV5b��q`��vdx��� ��a��^ߒċ�e+κ��&��{��W2Xb�{��%y���ȓ 4�jX7v��xc��X�V00m��a�x�f�<o~��s)4����ȓj��|3� 	�{v�I�al�O$��ȓR��@�A3Ze���3���p&D�ȓl��W�X6��1A�͗%�0A�ȓE;^��f-D)���n�!W�\����V���x�d<���G�=��0�ȓB�t��!�ψN:�!;�%^w/�����"t�/�8zqJi�Ǆ_�DR�8��z��5Z%ʲ�ļ��Թ4Xʥ��S�? p�3�V�I؞0y$���t٠]��"O8��p���B8��C�'p����C"O� �	Z]�p-Bc��;���KP"O��� D� ��ig�/X\|)�"O� ��U�	�R���lQ+�� ��"O����	����4� KX7�v���"O&ݙ6�)�*`�@+�$J�H�Xa"Oz���J�M��P'���Y�8�zp"O����Q+�����\�r�t�@c"O`��cD�"gD��JQq�y��"O��`�*��[��5R�Hո}|���V"O�4JѠ�#59S�MS�V<�P"O��w�ִPw~( �F��=}�mR�"O�\���Ö2��!6��9h\l)��"O��a��N�N�\���'���jv"O�� '�Z]p%p��Z%,>\h["Ohe��K��d)�"%��6��:��'�@���M�k���4l�����",n����\�6��C�ɫS�r���͏;�b��'��h`��O`���]�ic��*�
'�':>�x�iN$P�N0a��#.��lHu���
Uz���ˌ6if*��!6<u��x�'g�E�6�3��I:X�0KD�	� �*ucJ�wr����i
<Y�@�O�w\�ԩ�@����`$c��B���H����Q:b���t!׮X��D
eb�OX�x�Oӄ_�r��)��m<0qa��ipج��(=����G��9��A�	�'(6���Xr�\�A�������O�ęcV�-ʑ�E#�ߪՉ���G�5F*�s���N;@���	�
�!�ĝ	c�b��R)�5����$�������.!")�b��Y/|9��݃	a��r2�1Oz(sQON=^�L���Dx��'�H�	!��E|�oڏd+�=�׉D/?.$��D7���2h�|�R 4�c�A�6��z2gݥ\L�	��y���QGO�+�ēY�6�s�.ޙU"ळ�K� �"����<2��1��J!vT�@i�B�Rap��l�)���ɢ�r\�P�:�Tp�L<U�d� ��أ��f/��sf^*}5^�3���KxJ��"{��S���T7��afo�>7����բA�&����'Θg���k+�H�$/��ם<`�8x1�%�1UO�98�J�'P��0R�CXbK���NdB���!c�(Xq%G0VK�㞴K�+]�;F�T�D_m�`�x��5gH�b���#}2+�::�GA�A�
U�n.woʀ�qň>B��9Q�AڜGG.%��M*]��s4X�G���>	���jt��7�~@#�h�a~ԠAA�Se����<?�q#.�����;l�AK�σ38���Rwr��f��lP�h��$?�-r'�.8Z�G��5��<�'���Y��?�$�@IO���?�y�o�&2րc���!g24��ʊy���0��M�W=`�3-����ϙ�'0��2�u!ť���5��.x$i �)ē\> ��NK�b����GSR�N0���j�`�l�y"e�i�����3�t�0���:	�!�I=0#�`%�"��LᱏR�1��b�S�d=�����,�Ac	<2$�`"Ui�O��#�#�<[�"u3� �rw$P@�C�P:R��嬓5V �Gg�<Y�/W�J�N1��C����ߴWZ�+���/Yt�Bp�N�?��m�W��<cH4�%/c��H7xST�+�D`Ӱ����qr��֯*{��A&�
�S Ҕ`�7LT��c�<Yc"F�(e	�Ύq@�E��O$Z40�M��G �+HV@� �9f�����D������x�sf���)���"AۨNZT6��.��e4S�8\�;*��A@'{�p�g�Z2imTԊp� sH��}��9�v&n�g~��0�u����K��$��u��\�L�>�K$,�y���x�
^�",�ي�R=Bϴ��')ʊ���H������!�%ѱ��Q�D��f�Ni�]`�"ړ�e�|�Bٌ�����W��A�5�5q�a�=찝�k�6b��1-Їb��وnZ��|;&P��c'�ιmd ��c�Y��`H�';`J0���,(�ԥ4Oټd%8�XS&���1�PD����eW�ȥ��Q���7�sȜ豁?F����3���p����M ��$�m���I��:>|���)��xf�|8�f,e��7V6Wkl���L�Gb&@��L�zXheS�&��|a�l �6���G�4Qf�VGf��t�̀f��l��ֶ\Xfy@4��N&�D�8.������,OliX&�"j�dQ��ߍp{�<;�C%�j-���V�d���P'J1g4��1"-W�o�~epV�^tq�'�n1:�M'�p�Q�B0RXs3Hߣk��Yr��$,qO� ��KNi��� ��D��3&H�~ ���
�>c$��&��yƚ���A;�$4�S��'� <�c�R�m ��'B��B�`)m8�z�G#*���.OB��pJ������ٓo����J���̹(K�`���6�W�ZPB�$���v�^=gVh�@�p��+�a��o���؃��ž ��53W��A���ñK��NRD�Kr��t/(1T/?������!��!7"��yg'�'�Dc��\�/��'�W �p?�5��^ʐhA�A�Z�B��E_f�w��!>��nU�orJ yA%W�xO�ty�A�_�X1���J��>UI�BZ�[�8e�5� �Q�á(�� !�5�%��\���`���`�8G�_|���m�Y�,I�׌w��I`q�ʿ:�le����� �A��e8��x���S4^[D���>OT��Q.�5�,m�5Eňy�i�W�T���d�0��6[QV����{Zƨ�a.ڥ*�k`�jY	�t)�6��x���]0X[D,�<N��`���\��1�u 7@���$��H�J���}�x���{�T	����+��nԷaJA�� Q&�<ȉRHߵMa~�� %���`�,���H�a#@�["��!ˁo�"Q�.U1mDʅA<�<��S�	�F�YS�^6O�\��?;���:,��6{���4�I*0�����6[K������}�p]��CޒJ���l[�@���c���yQ�`�$N�Z�yf�A�W��yG��WX���Ӭ��z���P
j,@���}����Oϣt4��vBջ;�݉c�|��<"wC��l!Z��1c\�9�`���c�6Y��1 �J@^i�p���O�hC�eZ$Թ$�Ֆ	7����#�0.����M��tJQ�Q�P��0��ڨ�>�i�H@�7%��7#��ʡ��T��PU�� [c�p�jtg�6�Ȥ�F�E(�]Y�'jl0��I��,5�!Z�
l:N=���Fl�F`Χ��8��ա\綤�4�Q�z�L�����;J��u�*M���=G*�Mp���n�j'%�%[��3���-�@�Y [H�3�Ӓp@���¨D���A�;c�01)W$ȏ-�F�iP�"_^�+�vL�԰"HE��4��GX&Q�R�� jM4l�Á���Mv�MJ�ND���0Y#�I�4d���hJ����	V���TE��C�A0y���c��b!b�YUdA�?����K����i�bW��$��?JP��$&N,23�]�U�K��p��s��*����05�}�3�T�O��P��בp��j���#8�j���B�gjt�Bl��|�����V)r2��'/�T)Чo��?�r�:�G�b``���~����-��3�t�ޞC�r�b�!�!;D7��b�N�����[*�т$�{o �@�I�>9�����`�*Ex��'fR�4: ��s���M�,!�Q����H����>�B��Dn�U�B�M�59��c�T�O� 	#I>��)���6�aԍ�,t�>�ZC/\�%x J��A���BwhC)1�F��U)���8�Q���.q�$�"�T��?���#6K�$����$J�L8a���	(�)B���y�DY�d��S�'&��qC�������w9�a@�n×KkX�	'xzt�C��U�(@�t&�y.Ё��ƾ�M˰ꝅ(�Ȉ��BO:��ȸ�A�N�nԣ"@����$��x�'�I� �G$a8�my��׉pZ8�V!�6r�b3oNVc�c��ˉY$2�E�*3��y�&ϻܲ���� `^��"��NUk�;p�J](*�5���e	�D_��	M:@N, �Ajk��-)��J'/$�!�hȆ9RYYA˟�5���q���v��p�'OP@bPÝ�=L��AOϖZ �k!D��7򣔜��@��A�JZLrP�"Ô��`o�G�ԍ ��ܭ ʀ`x�,��B</ Ѝ0�C��&΂xH����^ S�m\��ד`C0 qVL��dl{P�Hf�t���Nq0��7�ayR��5*��� �#c���*w�B�^qs��MLJ�ZJ�,q"��A������Ě�d���"ߴ1�� �ٟP+�]�f컵��Y�&0�P^6��E{r'W��~��u��$p��V��e-Վy}`��f��q�	�>���S���o��i��c��CQKK��?������APv)�<����'�x:��0p��DKBoI�"MN�`�#ɺ+�ȉ5'���K"dՉ5�r�,˱s��TSω�&DZ�03�� !P�1��������;&��A������?�w���ڔ3�l�zT�1����R���i����m���MG>i�Dy�K�W.�K���L�f��V�t٨u�*~�1H3��&m2�i#��'gd��*�6H�)�� �u�VY�FG),��d�퉊!���奇0��L��#FpOp���=YOn�qs���[=f�9�ǺY3�ك儆�4��|o���ēxԈB�g
7-r�  r��!9�`�f�Wq�'ݶ���@�0�ꈳqb؝_�R��W8.0,��)�4},�M
�!܋d�r�oZP:!��υ�H�:�k���.q?^dH �k�V��t�C9�n�,�$Ӻ\��pcԞ��&�x"��)?
�qRļ< ɱLs��,�P�lH�Sb�-Cx����,Q�B�9%�F�;&��*��ǙiR�
�l��R�h�IN-��'KRA������¹}ʎr�d����Is��v(�P�+��A79����شe��rªN�p����m/�z�R�it��t��&D�I F�"���ڜ%D����]]�r�H�쌰!ج�q"��U�ـU(F���-��&C���E�\�z�x�L�1#ޢ�IR���[~<9��!�
roR�6�].�!��� �9a�J@����+�0Y������=�4a�n�@�@�R���!q�^�NV��fo)�:U��Йh!�h1p��<�HE�e�N�l�Ї㉁ ��e�V8���{��7P�}�n����� S�x.�Tɲ�v��@JN8$��g�.��aɡ.��	�ꐃa`2�$�e(HK��.+l�U��AOK��]UЌ��炜8���@�D�e����9+s2ȁÉ\��B  � ��u��t�V��gl�e̝��^8A��� שŚ}��y����.&��`X�t��9�ǄV`L��AC�\���N@�C�f| %�D<(< �5`y��(��\��Ĭ��%$&PD3�K�Xː�1�Y����Dߤ$V��!5) �h���*6m�.(���xr��U�
􈆈)`Ӳ�B�Ȋ%L��%� l���b�-J,.���8d�W��}j8 `5
��gw�,3��')���됒f
ӳ'��Pڤ=c���@NX)�Ȓ�wT��J��
�[dD�z�61�+{�`!0A�=CK^=���S2q�'3^aʀ
�3������oqJ� �O�����%2������G)HH�V�9��uj�-++~���Yj�|�2v�Σj9�����)	.�m��O�,f\���JK�l��D��nR|-kpvdZ��ŧ*
 ksn�/5�����%�LHjp���3��Y�2��jxfL
Q��$ (
C�n\6(�L�RH
7(f�[FN�7�XTa �'�J��aH'���a��|��5[��ٙ}�H@�
�3�L�7�_2$����A�' �����Ηx���؛~�\:�
Ywp�<x�$
�Grr%h�l���0<��e�*&Y"�3k�9`�:�%l��4]�-���N�7je��ϓ!Sh���#�P����:�:A"BEF)�<�<)J��	w����|�&mCWE�z���3��m����q�N�˰�#�qPO^�n�`�l��&i��� :���RPm߯b�,�0 1��"9���r`-�o��db�i�5~��@����=S�M:V❧%��D���%];�Ā�ś'e$�y"R)H7{��l�C�8Y�I
Bݦ�5� :t�0D2xh iϱ�@�x��	#$���S� �L�؇���3�6	�TN�EyP�
�h�|KN�R��0K���x�'U�6�B����+1�8)��N
AsF�RH�y����E)���ĖvJ�(I�GJ�>#��I�"����~Z�"Q�lNjII��ː!s����Z%�H�)a��p�j��Å˚Ϧq ­E �8�I�8W��AA,�#�\�EyB��D�ް�4�3z�N\�s����y��ͫO6D%��HD<������A�̔���1~�Rp��i!�t��܄�$-� km��z� ̶|�>ظam�Mׄ�[�'�܈���n��i�A�]�Jd���.7�J���P�I��m`�D�.]3��*cʕWC��D�On��EcL�1�\�Y�d�H��i@��ʍ�N��	��n<\��#ͻp��O��Yw��ʽ:a����O��8P���7)�`m@t��a�����ϋ�p��I�b�ׇG4~@)vh��>�,x��6*�t](�C�d���қw��`�0MC�m�p��nE�Y[�ؠ��η� ����+�R�lڦ���#B��)cx��?�&\� ȧ�6�I���=b�1�V%�LAR�s3b��Wc���zy��@	%�,�c�[��3
�6}Fo�/ɨ���k�?Y_�4� oS�b�P��R�	Z�:铵eɱ�&Yjfo�.ͪ�ȕҽ]V�(��/R8j񖅚
z�m��F�*�B�a���kQ���'Mk¥�=�,S�1�D�X��
7� �#ݖ~���Aڒu�q
q:�]� ['� SM�:�p�㝖�%h̓3Eӆ]��#_�q;z!���ɉs:9�
Y0n! ��A�WR�o"*���o?炴x�S�o���f�>�v)���+9F��S'O�]���3#�FWX�!#�8w� ۥ�\;?�,cD��3T��C�ϱY��9�C㎰B^�@�/�Љ.)Kxu[AGϊE�h	+U@ȕg�^Y# �V5q�xTj2W�\������'�S���: $��J�؇�]d-��2 ����xґՎ���Y� %�$�@�Τ�D��'�ܟ`%��p�x�g�V}�7�P�j Qaۮ2x�!�@�����H�������UI��(�
V�hP��[.2z�!��^��jY��!�D
�!�OD�-��p�f%NgF�a��eH�@�`ј�J���F�?,θ8�	]�A5Nբ��ln>�R��1'�H�Ԭi����f��*��<3��]
@9P���Lޓif0��H
d^��Í�	B<���!��n�qO�����I5AZ  ��O�o�@0��O�	�Tkte�cE��RgVK���+/��K/wrP4Y%$��et�l�RBI�eN��w��VJ � ��M*,���ݫw�9*wn֬VR�P2M��F�v�B1g"q�h�B!E��$�ʨ;d�({�'Vl�μk�2g��Z��ƥ5�d�1E�r'�;�M�# �`Dj�V�W�N�h���f��B��F�7މ'(&aa��96t���!8��Y"Ӕ � @�#!� C0Х
�cK��Ĩ�;<"4Cݪ!;��q�⒗�@H��F�6_΄M�C�Ɲi� �as��\f�q�eL�=S`́��I�8�RMR�
L�BI1dM�aSTd�3�G�_0��H�T�E� J�ń�<jj�5ø>!fQ�. *�i3�Я�B8�R���#;6H+#���g@,R��(���@�HO��� �̨�M3#�Q�T11t�A���q���u��ՙTZ�I'�;�CD���Dҙi�,�PBLDK�������G�{��4�C}hA$� ����=1�őU��݈�D�d"|b�'��4	wl��t���#�׵ $^�iH��qŔ6-V�Qyb����L>1"�,"��Ւ���-�hR&�2!'V��K,M�,��ڒ�|�'�
�y�-O!`
@�i�H��>H؆�ЛV��
�@T��6���-'EJ���υ�8jX�qŨΩ���䈉7S��8@�͋;��zb
O;(��ib�W#J>���c���=9���<>`��G*oӎu8D+6���XF$�(=rn��F"O6�1h�xϦa
S�J�Y��Y���E�2�9�S�?ΐ��E�̥8�P1 �F�l��C�3~`jXcwf�1
���æ��
��C䉾8�f�+Ռn�Ԥ�GĀ8��C�I�&�$p���ܸ�����"�>V�^C��s���8P�μa�t�FG߽Xh�B�	'L,P�{ �6bPSvCɾ`FdB�ɰ,���e�N�q2#K���"O�su���(]"�g�mM@!p"O����k�  ��Х�� ?��3�"O�	��Y��i�pDDg�Xu��"O���.S&GS$i*A����
�r"O�x���<d�t�ը6���P�"O��㶧,� �c�΄%@b�#"O��)BNŴԖyHt�»,D,R7"OXsF�UAH�Ёɕ�/��h�e"O�� PI��J�� ���5��x�"O��`��կx%`��7F�
W$�97"OP��[,e� I����̠�"O>�`t,�%X*�Y�O3xҤ��"O�0�)�6�vtQ'lA�>���"OBй�a��p
t�	<g;�H "O6a`�ϧA�*L
��B�T�0�"OB����>}>H�bG� S��#�"O0yb��I1H)��:��F*'(��"O~����{{6��qi�!\La�3"O~�{�A��xk�x�Q�f$,(�:p
��G&�p )���ROb�'� 2��F�N;N�*���l޹��
G�l�딍���M3�!PC�����t�BUp���q������M��4I���M;#���"�:�)7��lY���<*���9s,ȍj����wJ��M�W�Q�=f��A�Oq��Iz��)n� e�E�ǜt���h��yB5�)6[u~6�W4�)�&� �ĉrW���]yJ�:(	�Kbܨwd�˓y� Xش���'�1�� T�AT��	����� q��I��Hp����(a�DBL3
8��5(�	q�\���N�$�0���\�Bꕺ}���S�C�T	8��0,?�)���J�
 �`3�m� #�X	�⃺�P��i1�)��Hp����>�b)B�A�)xs����.;~�'���O=�ă����+��U�V��a���ɠeM�Z�0QeOE�gx�I[Ԁ����'*�a��U�̩�4�����'!
��tnM'q���O�>Q3�V=~�r qc%V�8�-�q�1�h���
G�7W`�������e�J�JUZ�H({q�j�d�N]4����t��n��B�"|�*�*8 �
(��q`�	�OF��҄`-�6mU�4�<	���vU���	�3���Xt(-@w9 ��[�5�26��2��Ȏ���|㤆<�V����F�f-� ��[af}�Bձ�?i�H�"C�L�Fv�V�2F%���'^���WB`�`�_�f�lx��#H�ri�`Dvy�IR |VL�ç\7ꔎ˕K����CY! Zte�-O,A�Vb�e�lم��"|�d��O�J�q�VqLX�w ��<���>Fna���U~���_�\����N� �Qh���eo��õ�O<�U����[�f>�Zg�٣N�|� �ƣ)�a`���/u��	GR��H?gJ���c��x)�D E�o#��{����Z��@
t�D�𩍯�
m��(ѹ	�� b�O�;l�	"s�	�l߈w�&���^84�p�WO{z̑�O	!�d��ߔ�)��.ad>�S��[M�!�$�M����N��_(�l�bꞦ}�!�D�<��\8��U�d�PC�O��*�!�$B�)��CBC�5�����$R�3�!�$�vE~���˛"f�l)�2�DDt!�DU8NҀ����w��%�-�>Mf!�$2Fx���bbʽs�th`.ܤp!�$��O1���F!��o�,ph�Ƚ]l!�d�=w;�Aw�[�-���&lW�<M!���~AڄI�Vk��aA��[L!�D�-7&�1���7!YЈ{��G�_1!���?�p��w M:Gp�nٻ` !��4l�����i��%^В�n^�(!�D�'|Pt�!g+�Z�2�nF�T!�d��"�F� �Q>z.�W �904!�ߟt+�	;2E�.�Hl�E�J~!��ؙ8����`o��/��Hq�h�=a�!�Ē0U3���4�{u�*��� �!�ݖjS��[�9hN�ʕ�%<!��&[��$�C聚YV~��M��k�!�DAl�����jNN�j�
S�!�d�1X]���j��
��Y�)���!�0b��z��ܼDژ��S��r�!�D	�#�^p��!F+�F��vQ�P,!�)/�x)� ��%l�҇�H�!򄟢ZK�qӂ��6(z�Ȑ�^!���r��e�JC��)�&�1�!�2K��tQ� t���&q�!�D��H��X��g�b� ɓ�n]�!���ba����%�� �̽+!�d�h�^ir�A�)e���čU:N-!�d�[��#'�QR��`��7,!��+ܩ`��.���[���6!򤘭-Q���G�8�(=�(E E�!�$ĞfN�����rY��Ns\C�I�P�``�2��19B]����DC�� )�� �bEppV�M	GkC�I�s <�y���-1�n�ô!L`�B�Iv���ˤ%�:�w(ǛSv�B�1��-C��H��J�8�C�)� �	R�E�\BͺW�],!� ��"O�QaGD��� l ��S��zA@"O8xi�^z���ɏ��ĕ��"O,���@�'����&ʃlf�[�"Ol�[(�Q$8�֠M=^�	��"O ��+J�Z԰�
V�~U�|��"OH��Ɓj6����Z1�	�"O$�KR�-+޴B'o� ua$"O��u��=g@P�MG�8�L��"O ��� yD���3̃�Fl�h�"OT�" �):~��
�Y�Qd��b"O�$���81��a2NO�_�ȱu"O�8�E<w��ԛ���UD^)�2"O�9;s�ݸ"�6aJ�M�~Z6�Q�"O��ϰmz�T��M�:��jq"O@x��)R�t	 �̼e,i��"O��P�]08<hy�l
a0�x�"O�ejg���M��D2��ܭN�H�R"Ov-"SΆ�b��̘2?c"��B"O��S�˅���R+؇?z�h��"Oh�2��Ѡ.8�8�]�:B�0�"O�ժ��
�HH�iRh�,F��"O*����ʭ<�~@3��B�VT��3�"Of����,5dX�%&�6E:�"O\y��ǖ�1��%��d�2#3���"Oش���3dU�����X+Jm��"O��KH�,>�BA��[I�m"�"O�i��a)\*���#a����a"O<�K�k�u�5�sO�1^�8�"O�("	�?jZts��O"���"ON�c�d�/Wz�Huo͹t
|� "O����팲��$�ٯ��$	"OTT�`�H�R�D�ʁ��)��,�g"O�Aɔ ]7莐B�oRf���qp"O0�oS.s؄P���t6���"O�Q�E��9����ICYz�3v"O~��0��}thQ��J��0Z8�@�"OV��υ0wX<���G!h:j��"Orؒ`�	m*7�D*A���Q"Oƀq�׊:&���gd�]��P"O����ɀ�9(��e�Ĝ���z�"ON!j�D�[�0u��J9)�2�k�"O�Q@�ʔ"�=c�.�?X�np��"O�<XפA�8�����BC>F<��"O>�Kqڝ{z	�!N?���V"O2@;e���`^Ld�&��#y���7"O��9p��<,l*�O!YӞ�*"OF����9����W��0���"O�+cF�4VBb��-�b�l);"O�%�G(G�L�q�b��p"O�����$=�dm���
�`vD�0"O`����1.p�0�R'8����"Ot
t撀-DY��G#-��a#"O�h+ǬJ�Gy^��t��^ԂD"O���tO��� �+Yt�x�ٵ"O��C��X�^8a��]'xHp0�"O���jx�Q�IÄ
�r��"O�P'�Z�4�f��u�U���T��"O���J�O=�,��I *����S"OH�`�Ӳ( �!�� ,v�x�"O|�sd�H�XUѥ��'gj��@"O�I���ۧ�P�&�ʔq�X�"O�R�M\2�Rx����D:0Y��"Oz�8̔�b)J5����$��"O� p����9<��mCfM��|��D��"O�t��!a�- ҍ/m�d x�"O�A�`�2wv�Ѳg�]�#z�M{"O�Р�ƛ�S஝��Z�g^���"O����/Z�H��qOF9 iա�"Opa'용f�P#�Λ(X�^���"O�=x�o�4R�1�3K<z6M80"O4��3��
0��h�;Oc�M�G"O6��R@�h� R�܂+O��;�"On�2�ެc�6TӢe�K|U��"Oz�BӅy���D�HH��2"OpLz�)S�f���&��
���Y1"O�<i�H	���Aǉ�(|���r"O�Qg"ŋz�6�)���(Oh�P[�"O<\���#t�r-�ƧtY���"O�S�@݈&�|�����+S��`"OD�#\�m��@��^\4��Q-
!�ׂMh ����X�Q�F�^�!���h~ ���M�:k�y��G��!�� �l�F�P򮗀S�d��i��VI!�$A�9R���U��(>�ɻ`	Ŗ=!��\>Ɋ`��A�34
a���4g.!�]������-�i�x��m?;!�d��" ]�G��()����mC!�$Is%�{G�\�|������!�YM��(��� ���j�$^4�!��R.��Z7�ݬ�d#��ϕ\l!��Į4����̓Y�\]r��fo!򄕺�)C^�~��@ !��7s!�J��4�"�5.(y#�lU!�d�=0�X,��l��u�r"�F!�$E�]eb�	gծDJ���@ɶY�!���M6�ip�n�
2҄�@�"C�!�C�r@�����s���QHL�Y�!�8L4�9Y2L[�0y� ��G��3�!��D5��a�E�EwR���懊%!��A�b%��c���?R>�뇄�!��R]��u��!mC�M�e锱�!�'%0z�J"oJZ���r��U3�!��j�D�'?�v�p$_� �!�$�\@:�#���$���/,�!��>$I����4B��`���*�!�$�c�n�X��	W"*�#%�9{p!�d��y��2A��4^��z��N�To!�� Qs؝���)M�`u���,d�!�Dևu҄���>����@=E!�Ď)��
O��v��吰�R�3�!�؁S.�%���<����'�53�!��K>.����0`�$��� 3�!�<zb��"ڙ0{�(6�^�!���ŵ�{ �W`Ք�(UK��i!��I�|L�QB�%�(�2��d!�䋢8��\A���4�f̂��O�
O!�&^F���,qo��i�=Pg!�đ�b_�,�S�G:4Z��6���t�!��d�({PC]�$,��{r%K�
�!�D�1m*���H�f+��c�M�1w�!�D�:��@��aQ ��J �_�!�M	�R܁� �:���2�E��S|!��M�rm~5�EM��s��tŚ@o!�O�}yp	��vA�5��aF�zk!���,��s�&#`5@@U�Ŋ,O!���Y>�����vø���捽S9!��j��J�o�/�8p�1�7nC!�� By�b/ݍQ�֑)Њ��n�z�"O�Q��K�K���U�q����"O:�����b߮�J���5Fi~���"O�uȂ�ՁH�@)gD�	M����"O��m�ȩ�FY�/0>���"OzAP���E�l)���X�y�&q�C"O48���ͅ(?�xb��0"\�R"OQp oMV0
x���7Z|���"O`A��˄)d��@!�ˉ!���7"O|�z��M89�P�C�!n׸�ʠ"OP�sb��>ޢA�#��<Ȧ�
�"OJ-1��M����s��C��^��""O ��E!V�C����!S7jK:(��"O8����]�XuX��b��b�f�� "O�aq7�K oWJYJW��j�Lt��"Oиs���C*���bO �b_�9s�"O��7��Z��DaA�F=)���e"O�ۇ�EUքx"�̘�7/�D�!"O��0�)2J�1�k	�R�K�"O���J��0�4����S�Z�JP"O��*�l�a��&�4}zZe�6"O~Q���n�~�XgؿX Q��"O�9�'W�|D:�`P?Mrd�B"O@�[�j��E�!OZG6�Y�"O"9���9$�\�`�-�uĴ�S6"O@�p��|l�ږI]c�ԁx"O\xq���z�����0�$�I�"O�����V�
���i樁���۴"O쌹�g� 8�D���J	�^t0A)"O���   ��     �    �  �+  8  D  ;O  �Z  f  p  �x  e�  �  -�  ��  ��  $�  g�  ��  �  d�  ��  ��  c�  ��  .�  n�  ��  ��  ��  ��  5 � �# $+ 9 �G UQ �W �] Ad �d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�)� ~�ȠB�-Mx$5�2�	�-��a��"O5c�CO!	b�l� �, �6�q��L���Ovl9�֥��d)0䢧�L>"���'m�M��U!:��fG�+�V\
�'�0yVLʱe %[s	D�|�Je�
�'�|+��D�n��k��K�i]��Ėw�6�R��È4WP�W�n�a{�@���d�ONL  +N�Wu8�Sģk�L���"OH9SC��F���
cY �b�I��h�P!���2>ƹ�'K3c
��B"OFS%��-I�2L2��O�7�`�ARR��E{��ɚ�)�\��&�0f�p��f��7Y!�D�Y�`}*��P�Z��qlk��$��Iìb�Ĉ7N�6 ��2t�C�I-�̕K��>4��7�vf�1��'ǎ虂M��h�p��wȝ�"{*(Î��~�TЊ�$b�!U��9��	OnOf�( R�'�v�Y�	����Dоm<4��'f�#=E�D��A؄U+��τ$�6\��a �yRJ�;��"��ڝ�p���
S*�y��B�.b�SCB�3���݆�y�a"\�l@�S7d���'g�
�y��ص�i��	U3�M�t��%�y2d��ch��@����G7��F��y�-�%�<	��J�D�~|IƆ��yrA�
�0ճ���vL��5�y2I�{��$����q`����&�y�O�M���b�C�|�a�'͛�y2
  ;"d��`d�s̤�kFй�yr�ñ0�dXT"����@��yb�[�@�\M�D���m�@�%c�y��Z�U��ȁ꟬lҔB�
��eNh��<�O�dZ�.ڃy�:p��a�O�����'�>|�H�؋tHY.�N��7���6��M�aK����'Q2�'tN\��cĕ^���w�\%�x�
ۓT��	A?!S+�81h0�SC�ŕ`�v�aƯ�K�<��O;VTJ�hT*O
̙�6i�Dܓװ=�������h@�K�%K���X��C�<)A�ːa-H!� ���Ƭ#��C�<y�d�'Dx0����*Ms��x!@�<A��+eHR����<fW��%�;T#��C8�p�F�π;���[7G�=�M{7m<}��)�S�#���D#]��9:���Q�C�I�px���ē+g�5I�M���c�d%��Gz ��b��x�D
^;��x��:�xҠ�2q���PA�5$�)�b�5ApC�ɔm��Ȃg�T<.�x���Ȓ��C�	$'�I�%�	�36��%뉌q:�B�%o���e"Ү0��e@����sSn��4ʓ��J����H��I�fb����ȓR�`1��/=b�Yu��JJ�=ۓih�c��4#^)�@AL�/ؔ��0yN!q��EX� ��ƾ�0���y]�b8`�r� ��C:y�Ѕȓ�
�@�[�:鱓�Sd����8�fl�7�Ĭ[�DA�%��*<t��ȓT���*bdA�-�"��ҊZ*e/� �ȓ[���w�@S�&|����JM48��_N�Ц�T�;��I��V<RVT��Mە���<Dht��/͛�\�҆��@�<�4�ˍK�����o�!_����D�z����>���3e��tJB�5&Q��,`�<�rlU�!6�2WͥB����gZV�<�V0�u��
8;|*mѦ��z�<� ��4�Wp����#oT�%��"O�9��K��c�6}��ˆ� Q*� �"O����FT�VN���c+�8~N �p"O��X�j�6��l�g�49|��"O
���dY�9h�.¼

�R�"O��A�����@�T$�u^F$�P"O��Cc�V�x,�¾�f�B�"OX �D㈅:���D�M�4�.�@"O�IC���}�D��#^$��"O��+S�_�u�~i��C�ZX��4"OF:��,d^���c�Ⱥ|꘲�"OH�bq�^>l���m��p)�"O=��	�i8ȱ���N���G"On��FɊYʸ8��çU�H1��"O�ݩg��Twu�Dƌ����0B"O\0��΄<����7�Tz�"Oh��F�,`�]sp��3x_^���"O҄����J<:��D4A��1�"O��r!!� K�` )��I.q/V�p"O���Ы@��P��:�~�+�"O���DaG R� 	��@̹ R��"OH��؆U���!`�5	TM�Պ~����B�B�,�4`�C�>#�M a�y"�˰!�5	���p��R��˾�y�'��=��
<y��w�^�[;41��Mk�4��6���)5�h�I#aғy�0	#B0D�0��虈$5�����(-��a�-��P!��	X."w6�c�ΓK�J<��ӑP!򄖿IBb�1�Ε>��`q��MB�!��ҏG�aS�!��y�a	,N�!� ^?��P�`
	���b7�V�&#!��! "%�2D�N�`$s`�Rl!�Ĝ�C8���U�-��t�PY�!�ѡ=$Ɇ�V��<0��+��M!�������&U�(��vJ�~+!�d��Q.�@��CU�֔!�k��f!�$~"F���-�,m�Y��P�y�!�̋ X�5���6Tb�U��"��)�!��t��y��Q�w���u Q�!�MS݌�9�(de��a �m!��0-��=��'q��;�^8Uf!�d��n&YY� Iꦙ�P��!��'9Ȁk��E��sQo��'�!�DO�=��<���'Jr%�g.Ĺ�!�D�/]��=�&�F�E��8��l�:<�!�D�'0r��NJ%}��CrKK�[�!�D	j�HPP�g��z�H���
���!�0�ɰ�g�]��i`7��0 !�DH��:` �L/Q،4v(�8s�!��� �n	X�g�R��$�7���i	!��W�e ��5�"�2�Rg �[!���I$�A�n��r\F� !�߬S��Xy���1p�|�8Ѯ��p�!�
~�0����dKA+n!�$"aKf ��NĒD�Z��c�U+f[!��)z6���S�Y9����E &6D!�dO8F�(����D�
ܐ���D֗%!�!�fA+c��#�P�ѐ��!�!�$(���k"����\s�cл?�!�DH�X�:���%�^�� ��h�!�&G�չgLB�1��ɧ�M�i�!�LǆRN-�P�����o!�D�NPDt�w�h�E�pt!�?;��Q�n<"@pЋ�e
N}!�� ����Õ�:�:Qȑc��?V�L�"Of��w��. `�ơZ-.)z5�"OU��H��2��M�D1��r"O,����$m�!���n�=��"OD����&j�2�(B&R��R��'���'���'c2�'nB�'b�'���/�� �~�qJ���j�'&B�'<��'���'��'���'���bS퉸U\�{g$Q0�T��'�'���'��'[��'	2�'���'s�T�òa�����܎?5^%�S�'���'���'5B�'���'�B�'��5�A��4�� O�O�Hq҆�'��'���'��'���'��'}��+�5T��#V�&��zF�''"�'���',��'m��'"�'�^�h�b��~�`=PL<D�I�$�'���'g��'�r�'&��'�"�'�v����/�zD�$ ��r� �� �'���'+��'8��'�b�'��'��%&钭)���{� G��"���'���'~�'WR�'�R�'���'ߢy���

i�)�C>�X;��'���'c��'�"�'���'+�'	��Ye��*L�|p�3�W�_Є�'�"�'XB�'O��'�R�'"�'�����
�d�ˇ����pV�'�B�'C2�'��'���'��'�XL;B펚q]�x��U}��u���'��'���'}��'�2$u���d�O�x඄�=Vr�; K�9�Μ����GyR�'�)�3?�Q�i�y���G�&���NXW�M��g$���S��?��<��l�|�GD;u�Jъ�ӥM��p���?��*L��M��O���,��L?��F6N�2&F�.E`l(1��3��,�'��>��e)>+��c����A�������M�D��@̓��O�X7=�Ɂ�#I�H��IgRY{6�I��O�$}�<է�OДyñi�Y+>!�;�䁬� ��vGx!r6O���,�?�vg8��|J��b$Jݫ��B��$<��	�Fpع����#��������9�	�8,�joL9@@��7�A��5�?W���I�@͓��d�-2�ʰ���S0[�*��W���5������p@9Ej�c>��`�'k�I�I
�2���N��hvV42�/9�f��'o�Iş"~Γ2r��!���=b�\�s$O��Γ2b��
�
��dB˦��?�'ZU�l���8yb~���RBM��?���?Y�&��M��O�����3�8�b�\#d�!� O�K��Ol��|���?��?���V�R��5�(�^LH]#nИ`!G�<�üi	`D��(۴F���'[�����H���'/<� ��V����֠�j"��i3˱>���i�p7�����zL|��'�0��(~-��z�`+X&�!�H�6_GL8!w�ݶ�?�AG��|�T���u��9}"ǛeyrAA�Z�x<(�h\5?V��Q,F2�'���'�r��7%���M�B����)��T�i�%N�;��p8B�<�`�i�rW���I���������ٴ~���c�Z���Hp�?B�R"�㒤[�� ��ia��O�\"W��*�������5�_�HZ@~�yia&]8�Iş��	ߟ$��؟��P��]��A���0;� Ǉ:hlu�Cϗ"�?��i�V��9.{�ɾ�M����T1@P��#,ʪ\�dM��Z�h�^oZ���D���� �4��V���M3�'v���=��cHԘh�@=QK�f�B��U���􉦝|rS�������ٟ|�@��N-{��ֲ
t>�����u�Rd��zy�Eq�h�sm�O��d�O������`dƐ�W���*�n��q;O��VPy��'ݛ�hj�l%>��m+�E�D�нt޼�@m�!D1,P��e��[
l������n���\�Ojt�4l��C��5J�;<x��%�O*���O��D�O1�Pʓ
ě�Iȉ
�"`ˇؓ^2LlP���_��H��Y�4��4��';L�NF���Ru��L�/O�d苇_�V�$7�ѦuXbd��eΓ�?!D$��i���^<��L6hl�b;�l�vHɓD���<����?9���?���?I+�"�:��%G�\s��O$$)j�(F�5��l_ß����@�y��'�7=�|S�bO3ywp}�����y��������@�4�yV�b>Uj�&Oͦ�͓Ht9�S�E�50�H���Hlh�=U�q��A�Ojx�L>�*O���O�|y2�C�cZP�qd,ۿy��r��O����O���<IÿiF��;��'���'hΠ�Fa� y`�t��ȃ1?����'�'ID�z@�Ho�&%�L#p�����}����l��ej����=o8M���m_v|�'_�D'���@�!�'s�2R�� w��p��W9N<����'#��'m��'5�>�]��)R�-_�Th�ѻu�h��	�MC����?9�CP���|���y7�M�m�cj�ub�尀�
��y��a�̙l��M���M+�O�+C���Ԡ�?����cAx5=���P� �O˓�?A���?����?��E�H�gM �y�JH�ԋ�5K�h�3(O��o�bR��I������?E2����3K�L�G"�@p����+լ=��OL�l��-̲�4g��O����O������e�~i���O����3P  �[�
)�O%	D E�?�0j1���<i������E&	
�͐��?Y��?1��?ͧ����Ħ���jXڟԃ�F<d@���倭4w|����U��l�ܴ���?�\��h۴q��Foj� �R@��ұC�� �,xRD	N2f=B7�~����O�,���O->��'F�$�p�� `��@���J�N�c��_��H��2Oz���O(��O����Oړ��xk��ʈ$���G��'X_�L�0��'!�lq����O��d�⦕�7�myBbsӼ���<	c��,E��Aٕ �8!�p��%7G����<�ش��c��Y`f}���ğ�1*�;k�4Mbd�C�z<�@%��0a����'�8p$������'���'�Z�Kl͗V�ry�+�4J�:�	'�'�2\�"�4uvj�@��?������֭��Й�\�4�HB蜠	q��,@�O\�mzm�=���|���x0���g��Y��#�b�>��� �M�>�<I�a�\������$���}���$�<1��F[�&��Ҁ�# �D��e^��?9��?����?�';�5�%oE����T��ɒG��'hf ��'J�ac�ވOlt�'F 7��OD��?YQY�����7b��7z�"� �%Fн2��M�%�i,t��c�i��	-A~Z"�OX�D�@�fAǭj�@5��)��A�X�����O����O �d�O����|�%�3*T=s�P.Pq���'L�fK�7gR�'����D�'��6=� �y���
5� �kn,�Y�	Pئp�4C�����O���dT�[�?O(4q��Y�yU� 8 �%Wd8�ۑ2O�eu�� �?	E&:���<����?���C>Af�hk ��k�H�LQ�?	���?����$�ߦuɷ�ߟ���џpU+R�0F	p�o
�+�|���YG�Y@�I�Mնi��O,e��>�t��D��81�D12:O.�d�	[�¡�E,ˮ˓����O�,���u�T�{@(�)yU��R��C"��R���?���?9���h�����8W��T�%΃������ρv�r��
�!�&f�\y2�wӾ�$!�4�%�q���j�hС�j�'^t%d9O�<n��Mq�i���z��i��O�\;�%�*qA�"c�~�@�S�Uƶ��w��Iod�O�˓��O��3��Ѵe�r !��N5��``��d��4(��ј.O
�d'��3na�52Ӄʹv&� Ҳ�C=8����O�o
�M�7�x�O����O
j೔!D*  ���2����e�gzB�BT��dC�<m�
C�_y�� Y�萱���$�f�G��1c	"�'��'��+߷&��I>�M���1�b�H*o��q;�H%Ho�3����?���iwY��3��$�ڦ�a۴q�fAY�-e�E+� O��<P�� vX�p�i���O�P��ǰ�:����S��56�>|���Hv��L8���UIU�r�'t��'�B�'��'R��oB���"0ir��f0uu��&~�����'r$�O���O���m(�dҵJ[�5��%��W¦5RǆV@�8Qoڱ�D��ɼ�M3ֳiܪ7��p�7Mu�P���j㲬�ӹ��[F�p&8�@�	�,p��4�	�u`�'��i>����H��!0�t�H!	F�k�N��4�L^�����,km�5�'1J7]B;����O��D�B�I��;BD�D�Mn�����@����O�|�'��6M�Ц��ش"����톢7E�B����O01ȵM�u�*��@E(Ke�i>����
޺+��'���-z��B���N}de0C��.R�֔�	�8�	ڟ|�i>�6,ϟ(�'��7M�b<*�
�ͮS2�0�'B����':2�4���$�O��n�X�N�Zd�W)YX$P���9x���4P���\(p�f���R��-I�$�~ڣMȹg)tp�e&ʢ-���/Y�@�Isy��'��'�"�'b\>)4��3(����"�6ӱ�:�M; ����?q��?�''�j��OT6=�8���ֲw�X����(���䢎ҦUz�4<W��ϧ>�'����q�z�4�y���:y;ȹY'j��(Y��*vA�3�y"��t���	�b�'��)����&~���`�a�:*��1�I�pc�4n�>��)O���
6r�9�@�3#� ��ɘ�K�����O��m���M���x�dڸ�V)���A2U$��Pu���y��'�lB��Q�{�J�pP���ӊF���Qӟ� K�%N� a���-c��	���ٟL��ğ���˟�E��w&&�Dq�6��I�������')x6-�V6���O�0mH���]�W�Y��
�J�T@x��_�F扭�M�i@�6��=B&6-r� ��6p$�ڥ�OI�%�e�Ɉk�$�Bf�<&,���� a�	}yR�'w�'���'�2&�-7���8vaI�r���փ˰/'���M�����?!��?�H~b����=~��<�fݱ-Dh��ST�p��4�����O��>�i�ּC��H%Z|P�E+E~ú4)wK�s�URE��<��$W�cB���������++
X�S��LX��p%�Ϟp�����OB���Ot�4��˓4���P%q��B�i�2HI�O<:Lx�S0�J!R�h�,�O�I^F}�w�&HmZ��M�Ԏ/"�hQ��F�|�sᄐ>'�X�rݴ�y��'u�X��]�?y�V�����e2��,A10(���O>J�����e|����ϟ��IğD���%?e���G�Z��'�ޮs��d�QCڻI�A�3BJ͟�����M��oH7�?����?�I>�gW�5]´�Tk���c�I�F{����>���i�47����&Kw�\�	�,��l]d�v�1W�A�JZ�abT!"g~��Fos�0�Ify���u�ڟ^���O��Ă"}���6��0��M�H�=Z"���O���%Dy"T* ��d�O0����E�Shf�@�B�aĩ��H�M���Ɍk��Q걮C�<���M㑲�*����	�c�cB4m�p�0 d�K�
����]<92�3���
*�I�?͐gO�ǺS��'�剈T+�٘�X�\���D�\�Iܟ�I��
�`4+�b��	ğt���?	�]w�)a�
[/,'� e�'#��`�m?����?1I>9#��?<�Z��� ���DZVR��'�L%!'<Mh2���=D6��� B����&fЂ�J�Eo
���?)�3� ����@�V���A��V;J�1��i4�x�'3r�'���'l�'��S�Ь(���*0�$c�;"�h��شw�q��Y(�?���R����?i��?ͻ���%�Pr��4-Z�78@�b�i��6��ܦE��O�������߈DQ�6�$�#d��hH� ͥv�b�m�DAF�����U�Od��|j��0��<��n��14܉���3����?���?))O��ow_�\�	ɟ���;b��,i�&1#M�k�n/��0���>Y��i$�6�{�ɘ+x)q��ĪYh��"�����Ih��V�k���y ����&��O��!�b��G�cȊi�p��q	�(���?1��?���h���0i��H*Bk�?e/���8K�R�������Cyb�sӀ��9T\�)��� �B�3'��va��	��5�4gu�F�ѥU��8Op��Q��½C��)�$�*��_���k2���|ؖ�c�;�Ġ<����?9���?I���?aq���Xj��@�:L��A{��?��DFۦ!�3+Z��I�x$?牦g�R���4������i�/;��D��)Zش0Ή��O�,�����Tc�mخB�6HbR6!�3y�˓W��!�"�O8�1L>	*O�D@��By֍��̈́���n�O�d�O�D���<��i��Zw�'��H���Ώg樻s&8I�r�Ҧ�'�"�|�O���9�M���i��6��fRX:�$_�lcԈ)���|)�F�o�F�Iן@b�Ě�4���o)?���uak�ʍ0���9�"�
r��q�H?y���OT�$�O(�d�O^��6�5F(��Ӯ�!f�	��țB66��	؟<�I�MUh���^Ҧ5%������5{H�É�=U�f�������.x�h��8�M��'�b�ߖ��P���1=����
Pɚ�,�ϟ��|�\����������|�ꔼz��� D;��J ,Sퟔ��Zy�	bӂ��f��O���Ov�'n��}����(_uLT���Ҕ#P���'�T�3T��/tӪu$���?UЦ�G�T���S�z� �$Nmh���e
˥��<!��)���DU=�?)(Ol�p��;(����gԱw��Y���O(���O����O��M�p�8<zȽ<��ihV�"@�q@�ٺc�@�^-
��X��'N|6�O���|��S�`޴?�9��ƚU(�� Gۈh�ľi��7�^��7�c�|�I>|F�
�O���L��RH�x�^9�1@��v�ϓ����O*�d�O����O,�D�|b�� �V����^�UN@�!��6f��V�yz��'0����'J�6=���� U"q�&	S�\f!�a,���}#شD�����O��DA�/3��:O�<s1.B;���b��t$�I��0O2�s�Ȭ�?�G�0���<)��?Y�N�tv�|��JhV$��@b���?Y���?�����d�ۦM2T 	����I���5aؕYԸ��l�"u���`�(�N�$s�ɥ�Msǹi��O�x���"!�j���:�=�P8O���tҤ�aC����V���g�O:�[��BQ�w���JP�e���Rx����?A��?q���>� ����?��O�*)�^��U� l�%��Ɋ3�?��i���3�'3�������<��Ӽ3QnB4o���N� Fq`�.˴�y�z�~�m��M`];�M˝'~@�Ġ�S�hd��Pg�3!�*�q�(f �SU�|2R����p��ݟ��	̟�:�-�a���C�ǐ�N� ��H~y�-~���[�@�O���Oⓟ���]�$O��D�OG/v�̌�'�6�B�����ħ�B��VOm����[��с�Y�g�i#r�L"�0��'Ǿ�Vg@۟�2Ó|bW���aL�y	����!֖��X�#���(��̟<�I��gy�Be�JH���O��c�;Dΰ���9�ИI>O��n�Y��Y����MC&�i�"��Na��$kH"%�HZ9��h�'�i��d�O��7,�ꢙ���S<�56d�P�1kc-�č�����y�'���'T�'R�)^�{�>d�҈�
*�`���$���d�O ��O����� P|y��n���OƁ�҈+m�5�2�)k�^��զ|���' D7������2[�(o��<y��u�81�$��^���D��7�)q�PF�D۫����4�����O��$R�n��r��-S��� #�ޅsK�����O�˓j�6��R���'�"�O�w��
�p��b�	t��a.��yr�'`� ��vl�p�l����'��oB\��X��$/y����h�>m�����-ضcJQ�'��$Z��D�6�|r��$f,,��2��+5�Xu�$�J4��'��'��d[���46�L�e��}T�M�W������@h��?���K
���|��'��^���B������Jߙ٤i3��@�d��7�����)F(�Ҧ9ϓ�?)gďC���������^\��@��A�'3ȐbU+�#S��d�<)��?Q��?���?�*�4����J�"`���Y2���4LWۦ�����ğ$��ҟp��U��'1l6=�z���-�A)0�&*[(�TK@�ʦ!�4#�����OU�th��3��7O�xriW: �� �ُF��a{�'�ҡ��GǟLzW�|�R������#���52��k�?�Ţrf��H���x�	zy"KnӌP!V��<���ix������@K�@�r�OTَ"�>�i �6�
Q�I=��U��)�He�
�n�\�	�h��#�!b�T��My"�O��e��9#t���9h�Ĕ���� ?X���)-I��'���'���۟� U�Ҳr^� 0�b�b,���ϟ��ߴ�,�q+O��o�z�Ӽ�%Ł4OKfãG�[���ۦnD�<���q��n�,>Xj�l��<���]������� H� 6@�Eϗ[Ӽ={c$�/_�,�R�d+���<ъ�Č4*�x �@�*-6L��-��b\����M[a���?!��?���t��+�^����a<�C1�ۘ��^��sӂu��v��?A���pZ�'�0SXpU�޵9�P*��5g�'��0a��ӟ�I�|�[� {�� i���@��[�AQ���*[�@��ߟP��Ο�STyBOsӔ���M�O�e��*� h~ A���:s��:V<Ov�lZO��&j�	 �M;�i�6�AM��z%䁠x�=���3]��9�-y�T�	�.v_^ ���XB�ʓ�J�;`Z�;�]0E��H�AIE*�,���?A��?��?!���O'l���H�v���2E H��@�'�b�'`R6	)��O��n�X�	$t�f܊��E0v�P�ZF�D-�NMZO<i�i��7��}���Ӏ�I��dB�(F�-Lب��&1-[|q��A��+����R�'e�$�Iwy�^� �I��D����<�(]�_� 9���շJ<�2P��$~,b�Oqy��c� l/=���'���O�'LC <RLJV ��L��Qn�4�y2�'e�I�M�i\6�l�'D���2�N̺--���,�W2���A,"Cp(��"�D~�Oo����;	3�'��B��(J,<��t�n�r�l_�\�	ڟ��	�b>]�'��6����H8�l�=}2��v�͜|�ʥ;�ͤ<C�id�O*��'%�7�ܡj�ʑ�
���7�*g�$nZ䟘*�� Ӧ���?�V�/@�)�D~��߄S�%c�B1x�8�(pB���yrU�t��I,\C<�E�G�W�j�@�쀾�D
ݴ!�����?����O��6=�dJ��խи#������
�V�5��45��V����?���w7��lZ�<�@ȃ1d;���2aZ�r���K����<����;���=�䓹�<97� [��Q�p�X��Zp�CE�X*ܴ1�Ai���?Q�TS4Tr�(P�~��T��r��(�B��>q��i�7�����'܍����NȒ���H'Y��'A)��P�t�)S"D�I�?��Q�'�8$�Ij�@E:6P�[��x��I�CV���I��l��П<�IJ��yGa�J��|���0g�t�[�A�D��mӖt[���O�d轢'�4�iޡʁ��*�x1�աםy�H�!��|����4��V~��U!Ƭd��>�ܙ���L����@�wx�H�LQ�>�Fy"fMG3�䓿�$�O|��O\���O��1&�Lx��Ȇ
D<��*C>In˓3�f��=/�<�U�'6B�O�&���_��s���f�f��Z4`L�䄔��d�Ezٴ[��6$,�������Sj�̃� "pЄ���$8�	�2��<7���9I(�St�'pP$���'���!��/�,�a�擶z��QA��'�"�':����X�h0ܴ<�B�X��R2 �x"�3�p� ǻg�\������Hy�'��f*f�&���^� t)S�)>�c��Р+�7�:?ѳ΋?���i�/�䧈���	}���㐎��f� hT!�<���?���?����?���D� �i�����[< �Mk��X�eV�`��'}"{�𥢧��O���O@�O\8Q�#D?�p���@��,���&�Ӧ��O��l���Ms��m��u�۴�yR�''����� �@���S|�XJ A�&9+:��	
N_�')�i>���ПP��-2���.\�q��/��z�	@KىM.�ٶ�Ry""z��$@������O$������uL�&(Ѩ�.O)@���SC6O�d!?����M#��i
��z���M�ڸY0���b��\���ܻ_��xagl���G˶����&�ua^�6�1��R'g�T���jF�a�r�zD���O;5٣΅)��g���]𰈚nY�7�d���nC�u��Ɖ��c�n�� Ȉ35���;�U(s�y�p��G�$�P�+�83Z(�ɳ�Ӹs��Q�{����#dpӚ�s�Z`� :�/�{p�H���I7fDR��/�&0P��#J� �@����d��b�W�[(���`�F=rl� *�0D�5XF%G�4��dB�L�q�Y��	�1<���5�8ѤF������AA�":�� [�1���dB� W�����R�{H�i�!G=L�|H�J�i�� �` �}�$�7�����%�$�����+�%HDD�a4԰�a�l��"c��	ߟ��	Qy�KR2�擠kJ�x5�95X��B'��<-ꓻ?���?a)O���O�	�U?q���Y$Zw���p�#:S��h�&�>����?����T�{^�%>�r��H&]���u"�%-X@�)V�5�M��������3y�����䗳.�a�A[;��X�Ƿi���'M�I A�^$yJ|������Co.	R�"ϡ'��5X��9�P,%��'���b��i�?�h�-�<�z؉�^ J�\Y�FiӺ�}	U�ҺiE��'�?Q��Y��	>|�|]{@V�P���'n�>�6m�OJ���&u���S�$���V[�l����(�qa`*�/{30 m�R�z��4�?A��?��'*����e�5�r�����7���FT�|�7�!��˓�?	���<Y�p9�����͸[H�KS"4M�8QS�i$b�'k��Ϧj��O�I�O���8��D �m�(w<	`!��.�����A\1O��d�O@�Tw�H����ľm�Ȅ5*ן0v����Ol�挑h�i>������'%S	@%�c#��<A����L�2f�v�'+�<�y��'g��'�剝{�`�w��Q�8�!��]'Bhy�	,�ē�?�������dC~�b7��+7�pH�]�e�4ё�d�On�$�Oh�O�!�4��UQ�
L���i� A��&�{�\���	ğ $���'�䈬O�y���^+}��(e�O��� :�\���I�����yybh�M
�b<� ���V/A	z� �*���k����%�i�r�|�[�L0+;�ӥB�U�f�.F A��I5�6m�Op��<y�
���O���5�oH�G��JA!/�p���Bԭ�ē��D6z]>���d�Ny�X�T��
�J^ ͎�l�iyBh�WR7mM��'��+0?	�a�#ٸ�qM��i���Sɦ�'ҖU��O�SF�sӐC�Gs<�p�kĘ/����i��� ��g����O`�dោ�$��B��Yi�If�C$	Cԥ�ش|��!+Oz�d�O�����O�{�h5�`����[�ha�'�����INy���>H�i>E�I�`��
�Р��Dϻz�h��#+ 3��8P��7��'>m��˟|�f���cB��1ZM��F�/a��':p��[� �IПl�	k�Y@	��1��` �Y y����'\���A�ؼ����O��ķ<	�S�d��e��)�>�򠊒�gPQQ&����Of�d�O(�(��g��c�!wy҈��$�>]*i���M�I���?q����d�O��@i�?m�fIϵO��� G'�+&z<��g�>��O*�D-�	şBƷ0FBeӲd���E%`.���W�]:Sn��E]������'1�St�����H���<? ���&�Ƞ�LU�E��۟L��K��?�r�
>ְd%�|�N�3]8!r7�V%G�N��G{�j���<���Gh��+�����O~�)�&,�Y�6란'��Q	��>���>I��۾l9�"S�S�D��$f���2��+E
M�f�����O�X�@��O.�D�O���
�ӺK�$pZ�X7�]���Ajl�H}��'&�2�⍴����O�e��bX ��=��DAt�|ŉٴn0�;���?a*O*�ɪ<�'�?�ӭ6�ruX��~̬;�O�9"���4�	X�y���O@��"E�3Z��:��[\���xe\¦9�I֟l�	���ȗ����'y"�O�5�׌G�TZ ���o�2>�R��'�L̓I5�)Е���'��O�p!�g	�F��A���]+k3����ibReӤ �����	͟��=Q�ݾEjX��f��[:�<۱&^}bcV��� )�O��D�Ot��?��n?'���^)^��pd-8�2����<1���?�����'yB+��)H�� 6.��4���f���q�ж���O����<Y��7|�4K�O7�X��i��!�aƢh�����O���?��۟�Q�)�4]��7퀳��X��D�5�J���	�"y<�I����|y��'��A�V>��� /=Ѓd�$��5#Ǎ0����4�?��V�`��8�QF���T�R�$���Ɲ�4���'���֟�*! �h���']��O��h�R�E�/<>���*��l�&�	py�A��O�nC�uQ���S�{��⥅�"+����̱QG�����������?՗�u'b�����)O*�ڀ`2���$�<�6��K���'(�́ҩ�zR�2���%���n��`
8��Iǟ��	ޟ���Ly�Oq�mN�Ht$���C�E#.�b.�q��6T(���U���P�PH�]ӆi�3�B���!�:�M�����I"����|Z���?Y�'O,1 t(�"q�m��A�$�(�+-�ɍz�t�+K|����?	�'b��AC��d�t0���Gմ@�ڴ�?��G��$�O����O8���'@�KI��	��\352�Bqj�>G��dT�'Qb�'0�韸����Q'�!��M��(�&ގo��u�'��'Z��d�O�݃�ȓ�	N� �G��9f�C&e��`��4`�� �I�T�'�򣎤)�����.Z�ѳ��S�o����������F�'���'��O~��� l��Q��i��İA�>I�a;�㛽_"iЬO�D�O���?��lB���i�OlؐQKC2MC. 3gb� {��*��	����A��?�g/�R��'�8:L�[Q9q Ԕ4t�슑km���<�����.��$�O��	��K.9b�%�J=.�1��!\����>i�EP @g�h�S� ��8�F3��%#�T���KO����OD%���O(�d�O��D���Ӻ����)!--� �U�{��a��Z}��'P����<Ș��O��1�� �?Ve����ӽ ���S�4mĢ����?���?����4���dL5:��H9��	�a�0N�XNZ�n�E��8�n&�)§�?y!��e=��7�
)ST� �\$W����'�"�'{����[����h��k?��նfv�P���D��A+���F/1O!�n�d��П��IO?Y�V-(f�kr��.`E�զ��� '�8�'MB�'���� *l��ᰃ�8���i���(O�ɷU��<�k1?����?I.O�����a����Y�"��h�E�,#�<�4�<���?q����'RA_:T�L:#�ɏ�@4���	}v��*����O����<��,��\��O�(��!�R�o���Yg(��0r�MSش�?���?��'�ڽ�Ţ^��M�2/��6�����̓�A��4��b�}}b�'�rQ� �	8(�}�O��$ȧ|����3�L�e����U�Ce��'j�O2�$�<s	h	�x2ɰ4z�!S�T�Q�� P���M������O&4J�D�|���?��iin�PW�2e�L��թǷD����$�	��z2�Exnb��j{VL���/אI�h��$�i�'$r�E��'"r�'���]��=� 0\�NS3��賈:[�*@*EQ���	x�~%���-�)�S>K�SҺ�0!�֥�t~t(lZ�I��@�	����ϟ�S`y�O;BFгN@����e�(B����'J� 8["7�H��D����ݟHXf"��d���ԍY�N}�WȎ��M������owf��|���?�'��puC��WV0��#[�g�E�c3��8�J��I|ڞ�?��'2��Zd���)f��d�M)RfP��4�?��h�,���Ov�D�O@�0��H��~%�� �ܖQ;�H���>Q�G�WHq�'��'��Iß��D(}��`�f�5U�����ۨD�H��'���'��d�O$�U������W�8&~��&�
_J�}QƓ�D�	��Ԗ'�r �!W��E�8�>(�7�?C�	U�C:\����'�2�'��O����!&��(��iA�-���.��ͫ�m�jw��!�O��D�O`��?QK9��I�O�� �L�����tlۉ%��n�馭�Ip��?�TCA>�h�%������/�Y򰏏l�R;C�m��Į<q��0a��P)�����O2�i�	mN�I��\�V`	���]�SȬt�>y�0�(%�f�NI�S���I�P�J-��I�0 ��bc^�M�-OڡkSe�˦��	�(�I�?-b�O���(ݸxaR�T�4K�tzh	͛�'M�n���O��>%JG@�H��p�NGg����s��,�Kצ�����I�?��Of�$��pQi+m���#�;gF�ɱ�i�t��'abW��������0��:8by�FAɱ:�fh�иi2��'��#�������O��	����6��C��4z�W�Z7-�O�ʓF m�S���'��'ԍ��,B5�,�ThʵW�NDC��tӘ���>#��@�'��	ǟ��'�ZcF��o��bj&Y��	���Y�Ob����$�O.��O��t�N��!i�xơ*�)$.�9��B*c��I{y��'��	��t���`�&��9�nu��!
^�F����&.���(�Iǟ���؟l�'���d>�!#`&m�*Hk���	ǴY�tEn�ʓ�?�.O���O���И���4V3����x��}Aƃ.
�6-�O��$�O4��<�� <����R
91�R4��O�%o8� �M+�����O����O~ �s���sӖ���腖!?���#�t̙��iwb�'��i���r�����O���I#(7�$�X�y�P��`�3K���'���'�Y�y�\�X��r�e+C�(�"	�fƃ1�����&�Цa�'!��GCe����O �$ퟘ�ԧu�K�|_8Ms�2H��C��C�M���?at���<�K>Y���S�<��x1sB<pt2тN�M#/יIe��'�B�'l��Ƭ>�,O��F�v���w� 4����a���bJu�$���*�i� JP8j�p��DH8|�̲a�i?��'����Y��7��OT�$�O����O�O0o�l�Z$�q��@1��m���'�割}KR�)���?���o���#��H�C{�rf�1��R־i%�L޲1�������OV˓�?�1!ށC�		�f�&�[A��o��,���y��'���'RRX�K3�N����+w�u��o,���OL˓�?�/ON���OX��Ɓ-��EyAk�Asν�&
�-���=O����O���O|�ļ<A�b�8V��II0�0�6놜V�eJIo�S���Iiy�'���'VDQқ'7�� &ٱ>����@�2��k�>���?����Ĵ4@��O62;(�HyC�^:y�J�!��\e�7m�O�˓�?!��?�����<!O����*#�@�2@� � }S��}�L�d�Oʓe`�1cY?)�	�L���J��X#���;Պ��D%T:�H!�On��O���
E��&�d�?�K	)Tti�"Q$�<��Gy�`� �$页iV��'~�OŲ�ӺKF(0���7��(+����æE�����cc�s�x��tyb��"#�R݂��1Y��(��Q��v�9[^�7M�O*�d�O>��T{}�Y����χ�mF�|
S��oZB����6�M듪P�<����(������f���5�D�.Nr4�V�H��4I��4�?���?))�&u��InyB�'���
���!�@Ӯ� �	'9��&�'q�I�Fh��)���?��
�"�agD��G�-bw�p�i0�NʿSn����Oʓ�?�1-�P� *bܸ��	�`0���'<:u��O��$�O&���O�� �L!jc�DO�RѪ�jy弉#�f]�J5�IGyR�'��	ǟ��	ɟ�05�ڛx��t9��D�P�Y��#�%���	՟P�I��,�IӟT�'�ā�i>���.,5:��`拐�x�����Nh��˓�?	-O��d�O���� |�\�F�"E�;,^착Q�.���'#b�'a�X��0Sዧ����OD+���h�`ŀt )M )���Ҧ9��hy�'���'����'�J�`!HQ�T8�S%N�I�x�m�֟��IGy�jܕ%��꧊?����҃�U�R=�4��N�7]��b�BL:i9�	ԟ��I˟�ڒ�l�L��yݟH�QCׇ���FJ[/w�yP�i?�I"z5y�4�?���?)��Z�iݥ�0�H�3��VőN���I��d�d�D�OB �3;OV�O��>y��b Y?b �f#BiP�Tc�rHk2��̦��I��I�?���O�[�Ĳ�ʓ$1D]���
;�s�i�ze��'QrW������_��� �dY����de܃/�B`:�i(2�'�r�L?�듕���OX�)� 4M3�L	�X����D���sk"�"�i��'�2�,�yʟV�D�O��в c�Y!���s�Lɠ:���n���\�D�����<�������Ok�ڄ_X ����QHQ�և��op�^�Mkg��<����?����?1�����ΰ]�P���g���0�aj�z�"�ѕJh��?	J>���?��i�2i�hm��Q	u��zDd �ef�ϓ��D�O���O�˓#�dQ6���VCR.K�6�;����T���%���A����	�w���h1zKS`��s��5�aF.0N���'�2�'k�]��(f��ħ�,�9�(�1GC� ���C�q�؊P�if�|�'g��B7��>���?
�(�l
�#פ�:�!צ}���H�'��Q�E'�i�O����й����p�Yߐw<I<���?	%��<�K>	�Oa��3ggU�	
l1B�T���4��$ж
l���)�OR�I�@~�o��iQ�y��a����k�a��M{���?��`�<1J>�/���	|t��6ǀ/��s�)��?��7-W�1ӒlZ�t�	��D�S��'p��1�H}��AR��ۇH�.c"�7M�-����"��4Ed!'�P(H��\ �h�vj#hΛf�'���'��ek��9��O��$��4�q�N ��E��2s�DQ�8���@�ZI&��Iß0���:#��3f�
<M��҃�l���4�?��m�jV�O���8��ƜɃɓ)j�\�YŌ)=�$0aTS�trC�c��'�b�'3�O��cΐm���@EB]�T0��[DGQ�1��Od���O��Of���O�P)peJ65*I	��4./���#H�vd�<����?yK~�GB�Tn��ND�p3I��8���jR� �bȉ'|��'������	1!8�����3^��9wL�g�r��?���?q/OXp)�+�]�|���5јT=p$�FE��u!ڴ�?�K>���?�#X��'��I��"�3I��I�U �6�*1ش�?������W;j�t�$>}���?	�qi�)!� ��%��V|$�q��5�ē�?��k%ϓ��$���h���MKb����M+*Of�ch�������d����'���2���6��x�%�$k���O��$' _��d�O~�S�[�@�С�S�u��A�_�Qmڹ������I�<�jy�P>�I�N�Z��Q/��A��t"5�] �M�s�v�'���
�U�1r����6$
!�W�@ao�򟤖'.� �'��Z�<��h?�F"R,���ZVDďG�,q����1O&4:��{�ǟ���@j#�_5h�R���A*�܉���M��1v8vU��H��T�D�O��'�0�{C�O�3��h��j]:=�T9�Ox����*�D�O����O����O��1��iZ$�pd�)Mj���d�6�˓�?���?�L>����?Igc��w|X�����4d�ъ�_	?T,���/XJ~��'\��'P��'�+|�I�?�z0�G���7��!2q�Y�nP��W�8��M���<�ɇ=��xU�sӤ}H��>T���(G�3HQ�M�!Y�P������	Ny�����'�?A��ڳ4�`�b��Pke���7�P�*����'or�Ė�NA��80���#hL��e��,�`�#�p�4�d�O��d�O�-�r��O&���O��d�\ �f��2H��R� e�B�9C�O6���OXd�5F\�M�1O��%hB��)��Q [eN|��a[�:��?q'@�?	���?����*O�n�~��݀�ٿc���ҮO=����'q� ��$R�y��t΁� l�����s��(+�E��M3����!��f�'�R�'F��k3�ɉ P�P9��ǞX�E�vF��� h�4feV�Ex���O�Ձ���p�ΚT�f���"�����ٟ��ɜ.P^dH<���?Q�'�7��(g�\I��IC[�(5*�}�J��'o��'�bL\�+��pѷ�C�q4QI���& �6M�O���#Qf�����f�i�u�Tg� T��y�Si�@eB&�>a ��d��?i���?����?���
"��Ek���&%��I�uF��~����?���?������?���f�.�B�@F!X8$�7A�Sp8w\{�'-�����R�~y���F�ƸO��9����21������0q$�T��'D��Js�͘˰,�G��Z�J���{2L�-g!|x���Nc�$ �D��K�̈��C��/�T�i6)��t\��u�2��`� ,�p�	�ď:^�@q�ai�?�:1��/��@4xB��,(��[�*�D�ʩ����2�ک�uA,QF��0�#,+�n�#+��V�JbG�GU�3�͙�1�g��d*4�q&��?c�H�=y4��p� 4c+^�@1�+�?��[�Ē5D���l@[�ʧ��̿b�����OV�Q#F�3ճ>�OzrEѰ'�ѳ��1�k��B�L#O�n��ANRS�x`�O��1�'�X7�Z��O�!k*�z�ˎ�=�JM+�&{9:��$�OR��$H� ���Qn��^��5PAMT$rax�2����в�(�Ţ\�n+FtQa��M����?��8��@$�:�?	���?9�Ӽ�!��7 O��@� Ή;/� p��-$�H
"�3i�g�#SL����L>I�Ά'��)����Zr���3�,L�#���<+"b�z�\	�}&�Ȫӧ_}n����Z̈́|#������'��	���|ʌ�Dϑ/I���ě9YgF��@��)d!�� �乂a\�.:�RGع�, e�������?��'d� 	�l�]�>�JSŌ� Cn�!�D޸Qh��U�'B�'_�lq�Q����P�'Q����eˎ�:��I㬇�o���n�5mج䘀�	�����E�D ��҄(�8��ǘ"���qZ�	Vl�A��Q�4��
UlE��G/
x��'��+���1�fWܟL��[�'l�Oܔ��]�%�Y ���(a��}s@"OD�#e!M%3����*�/nB��xd��P}�[����g�
����O�4�A��YVNh`�H$b@j)8���O�䐇�v���O��(n"�ũ⪚=r��Yt/��Aը�	V�� 5M����Z��3O�1ڐ�Y/Q� * L�{/�5�5�!�ы��¨7�ɰ�A�2T�v�8��%�(O�Q���'��R�KPoZ�~bFʮ6$�f�7�	n���z����]u�첲*��sS�=˧"*�t��46X� ǀ�k�dq�G�5;0�d����ױ:����'�r^>Y��+ߟ,��D�s�� �2�ļ^�M*���֟P�	���h�fg_�a:���Ab��?�O��v�:��4�ЙS)r̛���{�*�'��4��Gֵg�"u�=�&���I���'|��j��)-hIă�;@�9�OT�(��'������Că��7��(�RF���@3',D��Jg�F=Y<$�{�ɜa�A�&e+O4Ez�ܬM�R=�d+�?�b���a*���?y��z`慻a�ɦ�?����?)�Ӽ6�� L9�h�Z�ٸ���Q,<��F�I�+��[�
0�c8�3�D��'�A��;V��	1�6P�ycd͇��䆓s�n9ˉ�L>9f-[�Gw�IV�P3�څsF���?��OX�������ə�Sd@O�?Ό��B���Z�HB�	�S�
�A��Ƭ,����al�
�&�����O:,�}���<xY@��5FF1#���#,``����O��D�O�y���?A���4�C�K�$ڗ�Ѩ35Q���~F���r�'aJ����V��i
��:�h�Y2�_���V&F��{Q�%}���U�L�����m���o�`�D�<a���'���KE�IQ�҈��� ��H��'�M���9W�x!��(�b�\�9�y�ƽ>�,Ol)0W#���Y�	ΟKR��2sr����m�tiyW�B�h�I�.�����՟�ϧRi���A�V�I�^w����
^<B#֜�6*^+8��d��H��1� �|���4��;$�&&���Yu��p<9P�T��T�۴*ݛ��'@ �J��:���1��Pq��T����u�S�O-�g��x��t韃2�"=��'��6M:kR�i��%]<�U$��2O��d�<��"JC˛F�'�B\>��g��˟$�G�^>O�ix�E�=͊{fi�d��f3���4☧�P����\Z����.:�z�� �:}2�Q*m�O�A)G���rǰ��j��v0��>��+�ş���i�Sa�('2�Bc�ߞI�4�!��.��c����@x�����c��~P��̄>!?L����p�'���y�ڔZu�!��0	�B���h~�z���O�����l�O��$�Op�4���B�_���k@�R���r�&�	e�J=
�`(��{@t�B3�W�Bs�񁣃Y�%�Vm�ybg�;����}&��b�D�jS�F;���9Č�r�r���Oh���C����Y�H��R�)��-ک~�VM(A��>)�Ɠ76X�u-͗KF���F:X�'h�#=q���?�,Or��g�Љ&�`��!�D`�H���
ZE�]�u��O��d�O���ɺ���?��Ov������"5v|�҅ �	���ui��(�0�'�X���>&1�,zT%]�I��Ԋ��A�'����[��Ԙ����z"�u���?�R�iې6��OX˓�?I��LM:Fҡ����6PS�Mޛ�y�c��H͐�o�W2�
q�"�'�������^%@�m����	1�t���H�&H
��E23��%�Iß���D��I�|�fNE�}���#��ͪ�D}��M�,�h9�%/T�G�2ȫvfE�Ti
(���$^'f��Y�c֑4&��!���nR��b*˥��y����� � �(��-�"4�	��M+�iq���jz2�ӑI�^٨ᓭ���I���?E�$�Rf`����̎�S�<uA�/�x�cmӼ�9�돗%�h�d�̨^(�y0q��O�˓��q����|b���?1�'`�ݣ��Vhv��0�5{����R%/"��R��?17�W�6��$�g	�E�@玨G�`��E��:n���$��&j���Ӆ�L0��	}������U���2T+�${�b IW���ӼAx����#�D�g�T�#h�<\�\�:�C�`����y���?��7b�4����!Q�M��.D���']�t��[��O?���#!F.O�XDz
� S��X��F�4�<�$����㟌���'z����؟�������i��S��@|�Jd��P�n���zu@^���H�TSvbV}�g����#-ݪ.xa�i�7�x�IK>q�/T����>�OER�c��ڹ8�e;j��	�0n��b۴�?�䮚,�?�}�'��F/o����k�7v�f�� ��pC��������#�M|����G�s�����HO�˧��4vLe�"dI9gL��"ƅ�fU!�䉨^ྍ8a �"5����%ϟzS!��	]ұ��E����w�KM!�đ|J�9G_�y"H��ʕ�^�!�V� �D�d&��s	x|��� D!�DM?X�h��Cƚ�$]1�Q/?<!�D�
k	���.YYf����dQ�~�<�䂆2Zg%J�	�*i����7mM�<q��_�p���S���khv�ҁk�c�<��d͗2~$�V�(���f�C�<Y�b�K�"�c$l���4���i�<�`��l��I������Y/�\�<�I3�^-x"H^n�Q�Y�<y�D��Sn�T�Q��>�ڠ��DR�<��.�%7v�,�v'��W�z2nv�<��hնpu ur�����i1iX�<����B�I��� ?�F��!ES�<yt�Z�	������s����Ӯ�Y�<	�햮8�Y�4N�&}X8 ��U�<IejÑ[�p�`t`_	IA�-���O�<��狱uԪ�9�,�J"���"p�<iP/��O<�B,�'v�TCefOn�<i�圹�~����$1J1���R�<��C��
��	��#d�@�H�,[P�<9c�u��Yq� {0�qGb�<���a��e٣j�[9����`�<i�_iz����{�9BC�O\�<Q������yN�iV��W�R^�<Q!�#jX�h5'�oS�T�c�Z�<I��?g���0$NV4;���`p�U�<�Bەq&(��5�-'����p��R�<Y�!L�=*}��MH.#qj�ا��O�<�j4��}�c��-n\��S+�H�<q�c�"p�~Ő��Wl� �$�`�<q�7/B�f%� \46h81�ST�<�n��J������ۡY��m��f��*r����ˁK�l*�1�?�P �?ZܛN?��ǃ0����(:oZ�����D�!�ه�<�sM�fu��/%t0|���ȃ8�4�iTcɁ�M��~>z�|j-;�OJyRH��?".��'^9>�K�b�0>��)Nw+��("��?/I䄣��#>��喼�>T�LV
 �;$�S��n�i��S5��OF1p0��)E�̃Ǩ.b^����ቔ_���!fl�3B�Uہ�I	<D���F���r�.�fe"	�a��-#vⅬ�gh�`��I1zc�ࡇ"��l��xG�|َ�3�<>���Ȱ���0Y��I>��7T(9Y��(����Bp��SL�:i��t�F4,�!�dU0s,���#��
'�`���+� YF$qC���;Z���]�C�9����'��(cQ��'�<91�K��^X���/�`	��kf�|#G��;���d�I(7[��h�d�%Ex�{��r��35	�b¦�֌��#�ށ#�QZ�'����Ir>t����It��؁��7[�T$kG��2n,���ue�t`�P�IM�VT�ba�N,��qz�.��������V������H ̙�e�M�A�1a��1>��,� ̄�?F\���#v]�0�7�� �ܸ���]�����ô�)>��#��:u5 �
E�k�OjA�����)=�aY`K�
s�*Y(lQ2x㢁�Tk���q����r��%�5"�|ZdC�:�X+`I�?��k�~&^A�$AɷnD��1+µ1���c�$����׌HW���1���wP����`�=c]����"E꺈V���).([��I�;c��
�ũ(�����u��U�7�_��\��'~1�SO�K2c 5E�l�:��ĉ-���a���zW�1�..�����b�,�P
Z�~��JƠ�2̊���l�2H%��D�$��(QĤ(��*Jnj�)��L�J`�X�@�k�l���F�B�Ne�*�5n� ��RǦ>Yw.Kp�,���uC��?�CFhl�5�C�s$J���xbc��joX�x���y
� ��� �H���HU[ߠC��Q�i!�	�d���) ����	S0��PJ�&���O��T�mD�9��Y���\��kE�L7�V��O�m8� ӂ����48���b~ȁ�gː,~R���bD��
��,a�"4V�R�'������3�$[�<>a&��mS�1)�I�}��h"��B��x}�2@$s�maVB#?	�.F�����"D�E�X�F!�Phb5Y,O� 1gG�I7aZ�,���~�6���h�a��f32p�UI�(s�R�I��)k2+�1�>�{yb�Ն�i�.L5T4Ta�m��x�LM$���j�I�c>c�D���Q�
���zW��D��2&%P�ON���O��xS��	��O�^�Uj��J�n�x���N�ʳ�T_�F��d�_.,"�oӉF>>�tY��T��È�!�``p�
g�	v�����Й��I,{ȁ&��y�)(1e��
��'lh�F+�-��iK��C��M��H���'1h�h4)6 T�H����'Y8���V��`�'d:i3�"�2I��U�N?���ɤ2I���֡f�L]ꃯ�*I�M(Gi��Yn�Ʌ~x�&�hRǤ<ybĒ3/���F̄O�P�!M�!N<O��4K�DK1�1OL�9@AC>r��S��	U��l�sĄ�C�4�!#�Ou��S1ݦy��)ʧ���h���E%�8j�����(؈b'a"��V��J���|���w���M2��h�}�n#�F`�&�p�9�W�(��+�Y��mh0 ́t���y@� �O�	�O�#2������h1%�����s �_�Q	"�F1"���C��D��<�~�C#2��8��'�>�ƳX�T�$M�S�������r�'�\,�֓~T� E�,~���*O�� Vn�+ ( ��CP�_-0�FS��� e~��p�
-&�����0ʓ4'\)�����E!B'f�V�%��ăR�LB���etb  ��<�s�p�1#;p���jt��<�$�[�″J/Q(�|"."�X�O��;�"���4bR�C�)��u~4x���<�3�	��y��  ��������$	�EV��x"/�-� Cf#�>!�`�+G�-+���	[�O!��a*`�)C�k�)�f&Q�O[�<2T�A'4J\��У��g���Qt�\��ԫ��'$U����8@��{6n�08Y���B�̻
� �ɓ1���V/�7:��T�`� U��=	�ʹ'�fm���%@�
2��@�'���
е3����ң�
 r�Oĕ�A��d�)X�"�}t��O,4�t�$I[�:��p4#�Y��DyFE@���`��⍓�[�'�u秘Ͽ�6�_�'��u��\�I�4�ga�<�U"RZP��p�F(K�Jt��h���"D�-�.�4��(O?�	5Rx,��f*gE>͘PFؽ���'N�}�5���;��h�B���-F�tƚ� �1JC�ɖa,y0q�،�yr)�t��m;΂'S��y�CZ�7�ݪ@�ߩ����a�+c���{׈ˍJ���%`��O�V�0��i�(S�d�)�r:&)�4��A���g�r��$�=2�"ٲ�k�I�Rl�F�=r˺���I&_n�͓-_ȕ�CfIޠE�a�G]�@O�$�֨鰯��BE���� 8�&ʳN]�=%�(6%�K��E飉Hb��p�m�0@ꡢ�=O��`�ny��
:^�D링X."e��r�e&��/1�Hp �X8n@rͪgH̙+0�	�0\����ǁ�w�p���)���I�u�;w���;VFL���J�E��YY�B��#��@���T�o"TPY�b�ux��A6�K�UP��ڲ�B�0#����U`K�4�%��mk,��cL�C2�[�Ђ�!�ָ��[��Uh��D��]���nA����:�V#S r`�'�Xq�
#ƛ�7�xp�*49��Fx"O� b�"6N�=�P�*�I��E�69	�h>}��I�d(H��0<���Y��ɻAD�GI�� H�b}@WI�$@�Ƞ��� ��q)�'4�H  ��X����H�(��O��+0�]*�4a�N\LK��ෘ�$kƢ��(��-!Eg �?v `�Cu��Ɇa�V| �Sh�Q1$� �E�5w�����H	g��KRl�� �-ɢft�mK�%W>Ob-����P�(��̖$�r�� \aN
�%ق&�����C1�w2���3������*S!%�q1�O��1���ib
����+-DpȄi�i}^�Ң��H����R�O�I��j�6uFA�p���B�8e�0U�<��
�9~�lc���j����1O(���m
�[�>q�`�A5D�K��K���$}ᨴ(��ǥ1 ���P��; �2��Z�2�~].���5#�M��<���S�3�Rx�'�lx8���� ﰄ��釵"��H@�'R8xHpJ*o�nxi�ʽf�zi{6M_***U��K?��i��'�p�p��D�K&�c�c�m����F(\��d��y����U&p�r��T��~��M��;*<!;�d ��c� ��S���]�< I��4�1�b�,3�\�� �͂�@h��E���ә'� �[*(��Ip�O�0��OD��¥��e� ��N������'�.�1�&ʾX�U�7��53��a�s��fu+�얊y�����!G��'�͡���#Ø��O��0�H�f������Q'I�P�i�Ob�i��Q�~�׀�YF�k�$&�t�>x���ՉN�dJ�J�0�` g�"��8�"|�'������	�aZ��C�ظ`W�H���$ �e��q2`��+��Oɧ� �XGo��{.�8�m�7��$B���u�,���'޼��SJ^��p��E�YLV���'�%$1�!�޴���l�o��'֤��Al���D@:~� 9�"H�m56�lݽ  ax�8W�m��!- k�$(�JJ�f� V�&�"�C��W�z�*7�|2C��S�j�j�y��dk@�?Z�h�ϏAx�ؐtB���d ��{fK�)Ҥ���6~�"|Jg�G�b�t��q"^�{��Ś��F�pNnt�<�w�G{���D�T�@�&)I��9�0�O�b����D�@*4�R���⌃K��+2��$�������b�Zi24uB�Mțe9���p띞(~a{�$W3^�nXW��	K=��(��S�v�RS�5�J���3N�;���%Y��3��q� [ro^�
`#��rM&-��0�DY*�y��F [���i6aQ�L�9B��μ,��`�"͐x"����K�-!1O����J�))a�t(�Z�8��MB���r����dF,��Eb$���.:J�4f�|�ѡV� k68��-
x8���A�<���߅lZ`��U�Q�tڨ��V�I�O��\ʢF�H���
,5��'>1�=r'V2@���x!�Խl�^Y���t؟���^� 
n9�`��14���`���nl'�1H�L=�IY
~�6Ɇ�	�P�	���hc�Q�4��"H�d"?��@�k5�eY����e-`("P�pU�q��}��`bL�n�|"OZ�#Љ�!�+D� �*�� �����Zd��℉D3#��I*e�P^H�|�r�3`�����RֈYr�i�<y�aO'��8qa��r7�E�����3��UPT��3WVNq*sI�-��h&>��=Qp挶`����h8Qo�1`�H؟ ���;)�쉩�1p4�s'Ǌ9��)� Ə�^S�PR�O7򬙅뉀A���-�Jy��Yd��	#�T#?�Ύ�,��q�wm� /�\9{�B� Oj�܈LK�7�U��KC��4�"O�5�w.C�f��Y�m�(a0|z�T�4yA��)�pdK�©bt��9��WS�O�f��t*��=�����WU�,�	���Ҙk�����.���. B�DV�S\���b���bIi�� p�t���X��ӽ 0�T��$Y1jqxC*�ObI�����"b�"^���`vGG�*�D���	b�!���-&�t��d��lml��j�l嚵"�gN�����$K;[��T�b#g�K�g~�Ib K�O�� �	]�H���bq�0[�ܑ���*Ʌ �-pO��#I*o��'	n�y�?	*Px9$�"��@���){��͖	U��B0fҕq��B�6u�qs�-�s%�� �ܠo�fiQC(G\r2SB_*`���B`&�4�ɜ�*M[��Y���9�G��;+U����ɼ?*pb!���͢tJUT��5lN����v��
'TdCq�'�|$X�HN�X�@j�5�s�'	�(!�@ٲpy("�_7.{���
�'(�����Q����ڬn/���	�'=x���┒e�
t�*�Y�:�3	�',���%�'Z�|�0O�'N|<#�'S6�%#��gmD�c�LT�?P��'�Xh�n���䞏]�d�z�'���
'�z���1�ZJw����'��\S �Z�g�2])��ԙ.`�Ԙ�'s����!j�t��À�aֈ��'p�0@(֍���'�-"H���'5�H�v�,�>�'���n����'�2%�Y�T�)v�Љq�'�$JR�¨;/Fd��iP%7%Bya�' ,���M�i��� jޅ+��'��Z�&<���t%X�Ф��'���+qH�*����g^�N�b\�
�'� �����%[S��!XkJ���'�l, Ci��>��܀W���R>�R�'�I�ぐ�1��*�C��E�}��'0JxwnD3"E 5H�5?T��9�'�d��Ί�l[��Ke'L2z��2	�'�L��� � 9Q􈞨4���	�'�&���$­&�Z�k���+��Yh�'Ә�V�ű�BP�BI�5)�tP1�'N�|Ij�j�tZw(�/,���B�'���D��[�f�{c�],P��\i��� ����[!djf	�g��<q"O�xj��b�h�#��}���au"Ob�� n?�B@�#ļ\��M �"O����cb��iDĀo�0�"O`���\�-�J���	@/'�p��U"O�U1R�ώAӪ�8�kX"?�t�D"OF��'i�6ƶ]cvJ�i|ؔ��"OjE@�ǔ� |�L��鞍x����"O
ur&��7)�<� �
Wf��1"O�91�6�@�c��@"FPL]ɠ"O�yd�T�gu6����0�;�"Op5�bG+#�� gM
D̴�4"O���FQ�B�P�G�;��*3"O�\
�.[�&Ȣ���I;/�*�R�"O��A@��(���;��|z�"O�EA� �6 � a�֪0a��S�"OFؑƦ*��$�2c$W��DA�"Of��NC�*���EO@�1�ԍ��"O �C�Cڍ`�v4H4��a�Z��T"O�jc���?� �1@��Y���"O���U��9��e� b�Kg
��0"O���F�*̌�ub�>+�z���"O̓�hK$G�<t�V�V�x�T�8"OV\�uޛ����e�[���(I�"Ov$*Ȝ@��¢L�*
� ��"O�d�&/�*����"9&����!"O�pxA��y�H}��!(t	�,jw"OD� �cR-[��H%`�	s����"O*�6��CD	�fDיa�H�s0"O�� -)F��M���
�g�09�f"ON���%��\�n��� D-S�d�aC"O�	H����$��i���M -�V�X�"O� "��!?ӜUA���!(�`-˳"Ol�G�L=-��:��0&F���"O*�J�k'�2�z3/D.4.bLy�"OF�0V�- �t)3Y-�>�;�"O������j��ƃ�*~�&���"O�U�2B�)$<�����y�S�"O�����Z��z�j2���Z����""OhQ8��K�|5N��O�RE��"O����(3~0�%
]�Z$.T!�"OJa�sሞӒ肖I�"�	�"O�8�Y����9�%�-���"O �ҶD�,�P8�E[�+, 1�"O�)���\�f��QC���E�1"O��2c�K�%<Q�2��#|�};�"O�ers	�& F�B�"؍G�. �"O∰�e�0cL�ɀ��(�"�8�"Or��W�St芰�1��\��%"O��9��C���qQDn�+[�J��f"O�A"C-C�o0�䓄mW&i�P�I�"O�|��̨~��Yz��a|llr�"O~�8Ra��K�&�;Ui]�`�đ"OڬY��<�֙�g��Wd�� "Ox����Wp|ℋ�!���S"O�l�AÔ�./��;Є��`�L�:g"O��{�I�-<S^�+e�ׁƬT��"On�a���u�P��(��J^���"OP����+m��X��4	���$"OF(�a�o������Y�	���"O4𡆏l��4hfJE�#���Z�"O���� ~�5+r�Ѓ'�@�X�"O��beH��Z�� ��/EK��bv"O23�NZv`���nQ8�)�"O� ��Q$)3~�ޭ:��O<k�Ē1"O�Pi�*ƻi!0�Pk.0ͳ"O<H�W�8�ĉZ[gɔPj"O�L���L|.�2e,X)��(�"O�+�.�V��\p�[!��Qj\�4G{��)6還��J=�,�S�i<H�!��K;S���j�&�4��BcA�k���x�����oޚ K~!�5�
�`bf�16�6D���a�<#�<4SnEi�0�귄5D�d�O�6����sI�y�,�YQ�4ⓐ���
 H�<q�x��G��Tٚ�"O��p�A0��3���M�n�a�"O�� �M:��)'����5H "O8}�$SI��}K���-�6�K""O�#��S�h��i���#tP�A7"OΑZ��ĥ&�����6k&��"O����H`<�s���fOv(��"O�\C1F�9m��i�שO�+^�E� "O���`
-�F%)E���(���"OT��c�̀4�h:�#� ��@�"O�aa  m( �*x�<eX "O:� �&��m���"hǫ	�V�6"O�x��瑯=��IVf��Y�%�"O�-��ER���w%[4i	�"O�u�A�8g5��d��}�S
JH<��u/�ȋBA��.��B\�'y����O�VL@��'~�H�@x�6+�'I�� u%Q<;�!S�M΅����O��=E��	X'FbUٓ��!�:��V��2�y2n%Z�8�	H�F"|Rf�[+�y�-��BM�>C�}31�/q��`H	�'�6��Pi��x�� �$b&hش�Px2�K�ri
ç��u��<�.���y�N7I���pU��>ۖ�*rM��yB�ͧg�셙�D�2!ȚY!ReU-�y��1eCԩχ2�ܡ��-ʟ�y� v�0�A�I��r,y�)�y�LU�he�X�shB�>��N߄�y"́7v����#Ѽז�gꄰ�yB�L�3T ��EGp��%�7�y↜�}�H��&f��a��޲�y�d��y:��ѡt����;T��X�ȓ+ƨpB�#@�:
r�hMR�b�^d�ȓO~N,�WlV�����n�^h6�ߴ�O>�?Y�K@9S�,�t
	T9�r
�A�<)a�˛<��*gJݚu�]�ƈJz�<i�ˍH�J����.>��A��t�<iD�ܱ0/^��H��%�r���kWr�<	w!�1��p�bڧM�\Q�" s�<����R\|à��/E�\X8V�q�<
\:L�b��egk%����#N�!��)q\%p���>}��!��7o�!����~H8cKХ��xb�ɍ<-!�d�/\xZ�4*��9��xA$�y!��*S�ޙy"�l�R2���!�բ'�L�+�t�v�R���h�!���s�zd�G�M�L[E�ֳ-�!�+6����T�J��:���f�!�Ćg�<�
��]@YJi�@H�3�!��[�ib���.ՑQ>��@�o�!��N�?��dQ�'۱dY ��>nm!򄄌Q䄡[��@���l���Yr!�Ժ���v��-��l����V�!�$ΕI�B��Wf�k����j��}�!�� ��CE�(v{j�z�h�'l����"O��)2CD�p�ˡ��wh~l�e"O~�1�B�~^�X�� /a�-A�"O*9�1��A���b,��0M�����jx�����%����$5��`�T3D�p�3�E!:����唬24���5D���j�RWb<�g��� ��i5D��Y��
z"D�!��,J}��@qO>D���晍 '�)�5!� JE�� ��?D�|�� ,+����#� pjmp�( D��:4ѣeJ
�!��+0�h��n8D�h���D5)t�tX��mMb-��:D����@�*{�&1+��ܵ5��tK��6D�����-p�����>-]����6D���@H2G>*���P��*��i�`C䉠Y���`'
 ̐y��M�u��B�IY6��z�Iq�j�rץ�W|B�	��f��c����5qN� }>B�I�>�+�x����"b B䉢$����
4� uJ��1��C�	�(}�)B�ӎO�>�7�ցh9�C�	*8N�u: mB>�.y�vO�/�C�	��D]ʢĚ2KgnP�R�ˡh��B�ɀE�Xo�4$ʓ��?IBbC�I�S,v��)+-�4#d+�	-!vB�ɇ>��y�����4����PB�� �@�X��	$� )▌N�C:B�ɟXFV0۠M]e?�5�PF�@C�	�}fD$SЀ�t���IL�Q�6C��-PZ�k5�۹v>�@�.̬A/�B�ɸlSb��RF/Kv�	�:N��B�	7��a��l�:U�AȜiM`7�-�S��M3�����>��I��N�Vc�lC�<��Y�3�d��Ɵb_X�����<Y��]3+ X41P�߰��t�ab��<��E=m��D�Q�z����t��q�'�a��LA�s�����NƷ~�"�@AZ��y2�V$s�v��#�y�~p@p&D��y⠟�"��u˔h\�H�����k��y��[�V��1��@BȲ	*���y�O�G<T�b ɖ:�20��B���yRN$U�4ZgH�?/IB:�'�y��EA� �,crY"����y�K��}�+ۀ,'J�R�y"��J5�Hi-E�x �1�Z8�yR�ƠO��9��fRDE��J�yb�����4��#tHO���ybLH�$47f̸�13���B�!�UF����6ۀi��͇�J�!�-)%��P�Cm���,D �!�D�3��]0 ���N��"'+�!���T��ģuCZ<	|�u�!C|!��/���逭ͽJ�ȲsK[,k!�<T�ACdF
i�@9��䀽T!�䟕��+sE�k���J����R!��F�3Y�L3��N�����%!�ē�=�<җ�څ{G��+W#��!�;'J��`0̂.M*�	�'c�u�!�d��tx�h7lڎZ'��j�!ߺM?!��۾v�P�$Y *o�����!�rf��A��S��(ׯM0c�!�������GH�ֈ0��ثFa!�d &V�"�c�늦V��	;C>�!�D �E��m����.��Q@WH��>t!�� �;�&�P�
0@i��p����"OZhR�힒){.iC ���`�*#�"Oj�B��� O��k4�Ɉ4
Tly�"O�P)�3ׂ(+��T%�ҬQ�"O@�t�U�@5bb�#���"Oq���Ίq�r��5�
��&"O�(r�B%a)���B�?O���{5"O6E�Wo����ʥ`�\��d#"O��FD�Ūb�H�@H�6"O8�[U�hD�Jb ����w"Oް O� ��!�eחH����"O(DY�gJ>9�-���I��Z$""Ohhi�����Bf#%t��"O�iZ�Şz����</a2�H�"OD�� �!oNȓ/P�$CT�A�"O�}B�җ|?j!�E�\3~�r"O�Q�#ԙ�h��A>|��$"ODq�J79�-���NR����"O�$�1���i�l]M��bE"O����)Q�d0i�l���\$�"OL��e�C�0�ʀf"m�Db"O��j2�/!di��a�aP��"O��@�Ɖ�T��8�Z�HZ,�1"O�ā��E[�x�ҕ�/ ���`�"O$�P��S�F�(t�Y
FxΙ��"OR�:R$׭=^�m���\D�جI&"O@���֌|Qh�c̊Ѽ���"O�dCG�,;���H���O���(�"O(1��.6���1C�*� ��p"O|����Q��SA�rM�$b"O���,^N,�� ǎnB��c"O��!q��
�(4PV�J��0\03"O�t��
"�C�% �n)4|��"Om���0��)X"�2��4"O]��	�.� �	�/��1CQ"O�X�.B�M��T�3b�0PZ"m@�"O��	�2��Ȃ��L�mZ���"O$X�S"A�w�H�F!Y�]A�	Z�"O��kѢ��}���y1|-�F"O89[��`���pF(�Z/��13"Oz�Z3���m�y+�G�k �)"O�����>�r�R\�=����"O|�	V�Ǘ�\��T���/���"O�੄�r:�=�u̒(�"�"O��J��'��u�E,���t�"Ot%���Ƅ09ހ��KB$)�
m�"O�`(AO�0G��Ԡ��U#�=��"O6a��#���A��k�8�P��#D��AAo�Y|��
���C���#��"D�H����rǰe�c�4	nr0@%D��"�ˀ`s�+Q���@�#!D��Rc�^�O�}S$Q����&J>D�8z#�1+Y�ljDh��}��O'D��(u��(I���bTlV�i�DP{�+D�PR��?=�@�C��	�K���vJ(D����$�}�n��Co�H��#D��zU��0֔�&�W-���3�#D��AL�	��Uԧ��%Ԉ����%D�P2SD���n��R;6�,�t#%D���%�\�'��4�R!�6TV	a�l#D���5k*RRH�S.���TL D�`��,�
��IRA�&��#�>D�@J���-X�Gʝ�"���+�C<D�$�sJ�3ఘ�m�](@�;D�� �h��.��p�I�W��"O>�c�j�I��k!K�ua
�y"OF��ā�~��d����Td-C�"O�Q $�N�Q�.�
CH�'"O"m�7�;	��y�M8'b�	�"O���X=w��y�r�����(�"O���]r�	�J,��"O����Ú+{R�a��nQ����"O��oD�]Drᱦc�"KX�Bv"OZ4 �a�D'�BC�B��y�"O��"���e�t;t��B����"O4�)���Mc��W���8�����"O��a��e6��!P'�B�A"O���W�Hጨ����9\ۮlZv"Ob�8#%s���Cb��f/�I�#"O��f�._]$���@C#6�x�"O�9k�kD2D�%k����c"O�a�O٫PI�АF@^<^�k#"O>!���\�f����������7"O�u1U �/Z�b�p�(I�)�>���"O��µ�H1d�	V��<քdq�"O���v�A�M*�k��.s����P"Op�R�F�2b��'��u�"�"O@<���R�e��ř�Ċ ,�e"ORH�ڃV��p+�M�;�q��"O*��� ��,k�,F�j���Y�"O���P��O���هa��]H"OF�J4h�k�8<�4��fj�\��"Oj�k3��rx�˱I,7$��'"O�aG���>l� c��"@4ލ��"O�����N7d(>��U��>!��d"O��ТA��rFR%9�	
 rb�Hf"OX$��cV�?��10�e�j���ʐ"O�����˭6A�a*A��e���U"OЂ�(
bȨ9���:���à"OB	����o�t�bܣV��I/�!���d"�1
5u��h�ĻS�!�./�X�aԯ���S� b	!��U&4��,�#ϖ1%T4B�_�O"!�d�5n�#6���z���nG'f!��&ER4}��!Ѐ��J �A�!�$�
*��x���.n�<��L��$�!򄈴 ��|r%DS�qef�z�iߑ%�!��2�z��b\�k��<ip!�$H*.���X�`P�a����2bA!�䂪6���A�@'^�����T!��(S���@�s�(sf�=:!�D��O=���I�sך��6�753!�_#��yA�mϝ|�(�k���w�!��C;S� ��2eXn���$
1m!��&'��ub�P5@R�|�T�H�ak!��24��㏽sO4��FAN�`!�EZ�Ԭy�'΀<?6��O�#U^!��H.S�3�.D�@������7[!�%4��"����ݱ��E�tx!�D1STĵ[�lܝl؞i�aL0R!�Cd���Y�-���H q@M	N!��3!3��I3�V�p��;¯B,S�!�D� �� ��Γ�I�¸�q.[>1�!�$�x�P�IM�97�[Qs�!�D��qj�u"�G�@���)rY!�$U S����ތ
G�X���2U!�D�?#�����5U60����(Qp!�U�&�[ve�~5x)dO�Iq!�� ���1qf6��C�#t5�"O��g��8X�A���ud~� a"O��`�n�1��I!$h��J�T}�$"OB�r�HFl<�P�1T�,��E"O:�C�n�p�8"��S刨�"OXQ���[�M�X�����^�|X� "OX���d� 4�$q�����4�jW"OH�+���"��h�e�"y�����"O
�AO�;��)��!W�(�P"O�(��GA0-��А��	F��xr"O���&b�8ش+0�֔w�X$"O�e��P":�]B�-$iȢlx�"O����T�w�<eb�l�{����S"O�	��jT�Ae�����/p?��D"OV�����*r���F�Q'
y��"O搱��,R����;B�L�0�"O�D����-|V�ȧ�P�d��i�"O��	���I�j%��&���"�hG"Ou�WbD�=���D�� ��!�"O�(�p��~�:]8�^\�|H"Ot|��d k��A����XJ�"O�``��ն[&>������q"O�P���M4\�	J�M#݄��"O0|[����~.���!δT���B "O�䘦��G�i �.ӄ�Ȗ$�y�IY�xF�,�'��rs��{���-�ykI��H 5쌏nQ����n[��yj��|��ͫsH��%T�X��G��y2�^�o�:C�فY�l����y��ؙrX���U"��kn@��yB�M�Zɬm0�3)|h�o���y�+��M?rE�h���� F�y�2<�Ti��0�l���^�yb�]$x2�#��јx�=	�z�<)3 ǲC�Y��D9D�z�4
�d�<���L7B}�7�I7j��T���^�<9�f��[����?=J�M[gHZ�<)�%)Xc 0��ʽA@XD��]�<і�ռBC̨���=.��\��$�V�<��Z�ipP���[��D�ɆEJ�<���~K���1�@|��(VQ�<I���� ����	l�0a@�M�<)V�R�����NH��Qʗ�t�<�p��$��ْ�G���Ge�<!��?�$E�!��
������\�<Y�D $dGm�SHA<Ū�H�R�<��
��fA������̰'�N�<a����%*�SPam˖�z��r�<ap�*t4@ʕJM�K4���oIq�<��	�J�.��D�I���u�v-p�<�VÂ�\rČ�p
B�IR���.w�<y��N��/�.%qxQ� ��s�<)�������8KX+`����{�<��M#+佁���&d�zكF�r�<au���"c�Q��ѦcpХ����n�<٧�@�m�������`,b�S�k�T�<S�ٰ�$=	�mY=�@�KO�<Aw'���`1� Ꮪ3�@�´�FK�<IdA_|��9w�LI
y*��WQ�<���Wz��6�Ĺ�5nV��*B�ɇ+���⎍�p�P�a2�θ<��C�	W��%��H� *.l�F�A*x�&B�	#�|�S"��`�h� b�/gFB�ɫ_j�(S)P' ���v��1^�B�)� ��$w���$/kW�<�"O$�D
ǐa��P��y8�Ѣ"O�0�f���3����	
��P�"O��R�'6�����n`�"On����O�Tp��+	�=�g"O���䝋���v�©U�H}��"O� ���W��г��1t��<�V"OX12pO@#k��I;��D&��l˕"O���b%����q�Ca�e��:�"O����wK�w�$4�:AY'"Or���ٹ@\Ⴁ䏬4���"O��	���	X]��B�CG�
��#"O�@B��X�t���R0�юa�(b"O����	g 8u�υcl8�"O.��!�%B����	28.U�"O���2d��lR��3�&c�H""O��{�X�$��T9�v��9��"O��!�I�:1bU F�O���"O08��(dHYP����2�ڴ� "O�e���}����U���.�L]z "O�-�R�ۤURu!���.j����"O*(��,�r���J��Ӷ�-�yrρ L�ⴺ����`��0RF$���yr���<�\�4'�-Gf:������y��a�������?;z ��\��y���	�,���E.0������Ȉ�yb��?j���4���
`4JT��y��=�00b��J3<p8 �Z"�yR�P�eä����;�.�1�&J��y�`�5o�H��f�ق�$�T�y�_'E�Q@W��K^�H	�ŏ'�y��'P(�R(C#�Qaj���y
�2skP$X��7ST�ퟬ�y2*��V'�:�D؇C������±�ybL)�2s
��m�"���DĮ�y���#\��;��ڻ_I�������y���#�0ɉ��b�Z����A��yr��&.>���N�Y�\@�o؃�y2I�6>��e��R<VQ�)��n�!�y�j�sI����#D|CL�yR&�:V���"E�T��qA���y� �(Q��!���ؘ�	P��yR�ŕ��p��@�����B�W�y����:v�;�Ң{�Ą��K	��y�B49_���d'ל⶘F��y��֠�E+�Ҡ�uJȪ�y���;u.�1��	~�*���>�y"ELwE����٨qA~�{B���y��V1LV��+�B>x����k��yr���P�q�Bǖ ��<����yҀ�jR�(�ƌ��x 'џ�y"J+KEz�)\?J%L�g���y�"�#C��H�a�E�����Ҳ�y��HQ�Pɉ�O�'��񃷁�:�yrIGIj���Y�T���A�T��yb#�:cW>�RA�"PrNM�q��y�� zPU�EaA�w���W�$�yb�NI%��!I=n�ְ:'�è�yB�*,�: Rˆ<����Y��yr��}�L:��^𸚦���yb��$�d@@"�!'�1a��/�y���@�R}����#�FS�c��y�E>Abd�{�(�;O؝0����y�^�
Qh�(�'��E��Y��y
� �Xp1�K�"����Ǡ*e�y�G"Ox��@OW2�z�Y�*�C���a�Q�`��I�5����C�# �a�#��U�B��St\�H�H�z ��ۨ<��C䉈P�0��ˀ���Zq�>@��B�I�u�R�̖@| ��f��y��B䉅|��Y�҇�;7PՓ���)�B䉷]��X�2����C*�㟌��I&�����CaҔ8�0���~ʓ[�z�0��EI���	5��)����<m �Ԅ�*�AKÇ�;+���F˵%1�|��+m�q�G�ߑv>�{c�0o8T|���pA�*�z�XsddC,fV<��ȓ� �������:S�f� ,�Э��d�i��NB�A�2�������ȓ~s��Y����c�84v���X�'�r�I^̓7 �+��=߲��t��.Ac(t��V�������	gt�[G)ǧ�m�ȓ~n������1l�T��aL&]�fȅ��`)�T�_�&��s��-C�u��O%>$
�J�SN���@\g�مȓ4�0��nӠ.S�AkDGҔ�$����b��(U�Q�î�7�h�'�a~�F߶M����b���6�	p!��y�OҀ2��	Q"՘J�3D�#�yB`D	4X,��DoPt�(��%���y�	R#P����퇇QB�x� �yB���"X�ҡ�A��	����yb%ا�j�9%f�	+ެ�c����hO����ؘ��-�� �~��KTFQ�W��	/�Ȅ�z3�H0l�x~"��	�4C�ɫ_���d���"�Z��v� %�C�
öl%X$hdX�Z�@C�I,t�(@��16��E6C�	�>���CN��hŸ�8T��U18C�j<`X���u�tZ��)"C�
�P����%|�d�p@��˓�?9	�D,bP	C��E�( (s��5N{�i��e�4T2���!W
T5
8~���,�ڍ3��C+d��Z1n�>X���0�~�#5hڏ��u�e��I0.l�ȓ#El��'� -���Wh�J��%�ȓT��y'l�&h,J�-́]����ȓt0&�AA1����ƓN�Dܖ'�a~Ҡ�@������J���Q�J�y"��2_��!���"r�YC��I9�y�CG�1T�t�%�P"k�X}{ࡑ8�yb��J3h��>gx��k�/���y���2|`�W熁cfd��!F��y�*jx,mԪ+i:X��f���yf�:@ab��%��_��æ1��9�OӃ	F�0�.ēKׇ8֡� "O�X�+ĕ<��h�� 7T�%"O4�`������(�l�ް�r"O4��w���������i�`"O � e��3���:��OR��T��"O>��1F,g����m�%�D-C�"O������'�,ݩ���Cِ�0Z����|���O̮4G�?�r��taǻk�B���'Q��P���5[y:��t�=�P���'�aS��߯K��TlH,B����'MV͹f(O�/��3q�M@����'�<ErrK��_`��ٹF�j-Z�'U�����]�U��	�_b^D��nT�<� ��@�"�:Ex���E9 ��qT�܄�I�*�p�z2�Kw8nu��U�I^B�;x PBUM`�@"�I��<C"B�ɧ"(���̛�lL|�Q '[�"HB�	(���[�%ޡ�F1{'`�4�B�	&~*F�s!#¢m� �h��G 1ԬB���VM!G@H8!ܛ�Oćx�B�&|Q2����(7����DXB�I�b�P��� ��uYg�n�|B�	�S&�8"U�
a	~X�($B�I%�@@��	�sX$R����4�C�	�["���aN��TЙ�"�6NR~B䉀[ ���V�c鮍Xנ �LΘC��61q0���O��q˄��>OjC�F��2��W$7Z��b]>,B�IK�����"�2:�H����El��C䉣�XAK�KQ�_���U큶Dn�B�	�,���1�M�T�Б�⟭j��B�	�W\�8(c�H1,��	�(J�>��B�
�ɇh�q�@��;L�`B�u��m��mڻ:WZ��v� 7�B��#T0�th�=1>�VB	<��B�I �0� n�֜r���"bC䉁�&	 �싪(���آ`I�pm"C�Ʉ_��uK4J�>_�ٓ�m��2��C�j�ȩ�"Y�Ua~0A
0ϸC�	�#R��V)B�`�j �L�C�C�I�or��0�����`�@�>C�	�+�a�)�|;.)�hE�]��C�I0Y�� 墆YE��x��R� C�6HN!���E=g��1�0 L �C�ɞ3s�9
��Đ�bi���QVB�I+7�(��L�f[.��R,��|B�	�4�v�"��{���
/DB�ɆI:��R�L4=���g�@
��C䉮.���P�n5}���p�_	m�B�:bլ|Jeա;���G��+IUB�?��e�o�D]�(�(`�B䉲#`Ҩ���r2��J7j"B�_~2�z��ں7[4+���@@C�	.M�=�"��t,�Azri�1��B�IIy�(��k�(@/����f
�J��'�E�OR�SH@
i�%}J�
�'2�d�A��]&�s�O��W�)��'�4�C��ɝ:3pQ���?w�X��'^�e�u��P��{"�յp7RLb�'\4�X��T�u����Fo��)@�'|���d�X�?/��ڷ�I^�d��'�<�����Hx�gAZ�\|N�H	�'��xi�LqN��ǩ	�,`��	�'���#�<l.���@�4@I)�'Z��Α.m���(��ֈ&����'8DH@��[���O�<0�F�)
�'�"�J@�t~��Gd{6\Y�'��0�#��kG��+�
 q�`��'}\ ��B�:*FƩY����pzĘ��'�*)�"U�(o�A�"Ă�fP�A�'�2R�-Z^�cB��:�+�'�	0f�''����'[�Ҝ��'M���f."(��J����6	�']��;%��E�^�ٖH�������'0��jGʘ\"|l�*	:[׎�	�'�n�C�A�n��TY�f����e��'M�T����0|���6�0������ $�y! �'>��q�l�t�\X#"OziR!D<Z�2��Vf�I����"Ofċw-�6����|+}�"O���ANB�B���m�	r��q"O��!��I� ��x�k��
�.��"O(�طE�R�X����M�7"O�y3��D4n��9��+�QJ�"Of��S�K�0B%
3`Y�iG|{�"Ol�2V;s�`�gM�8[�`�u"O"L��Mӊ9`Y�S�ܡ~~VtBD"O��{�ĭW��!1�ZB��s�"Oh���B�O��e���	"1��(D��%�L�c���ԏ |�@��!&%D�8��i�`3tU;TlQ�!�xKU�=D����E-M��P��*[U�|�! D��ȷ�гf��r�@��-t<U3��2D�$��o���S�D��a�q8�1D�\��cU%N�u�W�8,*�2D��<u�l����7�����p!�3�̰��A��i(� � Z�5!�M �������I �X��n*!��
B� J�O�s;��k�-Ļ7u!�D�\��y'�� !2 �v��*b!�ě!,ߎ�� &��[��1r�(.~!�D	�z8 ��ɉ(��jԫ�U^!򄆅~���J�*�V�����K:|!�d� \b��#u��:p-�`���� r!�d�AJ^�{3(���Ej��˒(!��̣{��"ˣ8����@`\V!���!Ne���/��ph��,���!�.�1�u�ݕ~}�P�a�@�!��9��ׇ�!V�(���(`!��R,8��q�P��?��"Iƻe�!��W T�|E��*�
\��UHBa�!�$J�m7dq&)�t��*S.��B!�̈Mz��j�d��G
"Y$�+5i!�P		Ŝͫu�B<��*���/Q!�DH�0L�ÀD�F�����T�/�!�Q�	WX\�c��}k
(�H��L��	ܟpD{��Į8Q�_�30.�C���y��S�V)�-x�9����y��eb�`�D�,�!�ș
�y�H�xR�iC�9D}*׀��y2��G��[���f@`s�y�A�����c�J�P�i"���yR�6[�b1ɣˌ/I`�@�Ь�yrô*�hɲ6�IC��W,��y"�A:mP1S�
b��E)�װ�hON��)RH����ż�~�ak݂M�!�䏈V��嘧�=4G�Hz�@L�@�!��]LȢG��_@>1��.T2s�!�DʗwML���'���A��և�!�dYnRmx�E@�y[ˆ�!X!��/)����jѣ*h>x�!�'z:!�D�;�^8���Phas3/({#!�29��ŉ��|ּ�ˍ�4!��T�2�yF)ҧhD"��ר�!�$�����@AD 48�N<O�!�=�f9
C,�� O2)j��*F�!�D
s�V8[��D<H�3�9X�!���M�XA#�LBF�+WO�x�!�� ��x�GΉV2*a�1O~�!�ĝ!cZ0��@�.͂�)G��9K!�D�]��Q�D�ZT�=KHUh!�� ��p��J�L��x��܅P�h��"O`�&��q�Q�7b���V"O��9U M�yg0d�de �N� ��R�p��J���5!
8b.y�#H�#�U� 7D��2!A�3���9&�/~��)cVI4D�"���>󦹉�&�+�T-c&�1D�`��f�0�Ġ ��(P�2�Q�0D���"g׿GϮq�5lԨ?j�D�o-D��Ҭ�
�p��6R�N����k-D���ݴՂ�#�/�Z����&D�����	[���D��aj8�c�$D��Kd�W$?;T=I�M˥y��Y��>D�(�f��8DD�� �> i���D�9D�H��q�8�1�Lx-#<D���gAX�����@ΕM��e<D�����Q �T(��螠w����	&D�4Bf��9�(qΛ�6�Ha�bD#D���C.�'P�������=p�4u:ea#D�8��-i�.���&ish,`ч"D�tK@L
 N�`�a�'s]d$�Qk!D��E�ƵY.��sj�.�>��!� D��C��ԋSG�-�d聘Pk($�+*D�Ȉ�)��v�+E#ަP�3!(D����A�
���j@/�7f��+�� D��2i�Mqv0�`'�ꂡ��H D������;�Ɯ3��Q�N="�*O⭳���-=M�H�c�]�"��͸^����{|:Y�)��Q�h���K�K��B�I�q��āG.�8.��D��8B�	�G�P�&�J�A1�r) B䉜6�P���gR'v\���ϡ}B���0?yʧc��Ђ�/\�C���#@�l�<�g흦1ඝ@Q��R��E�j�<�fd�]�*�c� ҭ!ò�� �d�<���}��i*�K�4+/�����x�<�7��KA�M�H�&t�b���Ox�<a�!E�w1�T�ag�J(P�Qt�<٥)C3iv�ŀfa
?K씁�*�k�I^y��'Jў4��\�02��Ce_(��(�J�<�G���W�*��ԯ��$��md�E�<�`�S;%1XeSr&D�R�]
iW�'Yax�`ѶE�r�G�&Y��镗�yR�ԈnE�2�c�3*H;���yBi�n �L�ǣ
�%�İ E$@��Py�&Q	q�ջ�" �OG��e�YM�<!ALu�]����Tb�hI!�s�<�Dm\�uxE ��O<~4�E%�l�<Q���Y���tᝊ`?j����AG�蟼��e�dB3mYO��9�Pa�Y��2D�\{��^���Zf���	�1D�H�^&wƮ�4���;�d���-D�`K�f^� �&�Y@�hl�d�я?D�[�4'D�I2��Ј����/<D��q�>fuT�iQGM�g��|jVN;D�<Qt$��LfA�g޾3�{7+ړ�0<Y��_<sTzH��-�]�3TU�<1� ���%<0���H'D�P�<��/\#
�2�� `B��m�c�<i e��l �k�_7S�j%�Vc�^�<�#��7h1�P&O���R�+AX�<q�d�U�rhF�-9Īìp�<�@bE|%�4C��Tsj���Ct�I�(��W�k1�[� �,i��)>OLE�F�<D��jG�і'�������=)�0y"C�/D�� TH`��}�>t�)�2�����"O<X���_&n�8|�QWI Ũ�"Oip�@J�vp�g�	,MP=hA�'��Z��'���
<i+��}���!���6��1�7d�-G����X^ơ	�Ƅ��z�R�H�U��'��)H7��l�P4���B�4�ȓ)~��v��K�"�N��T@���p`�$R"+�Qg��IR�A4��4����Ā��grv���>�Ψ���H7 (ր��Ñ�tm<L�	F����k�+)1�H�S.ޡ�
��ס3D�<��K͟ *��u�߱��y{eF=D��j�E�5&xY{��d)��;D�@� )_`cE֤M��7B4D���FU����	�H_
U��dy��,D��;-��Y���#�랞}����W�?D���ܲU����ħ�,e-��q�;D����]�_�tm
g@_�1�*�Bԩ4D� �,T<5��E���-`�T8Ea4D������\�qpv�	'�����0D�|r�F(r�DH���0F챸�-D�T8�NY-(`�F�.��Q�g.D�L�1,K
Y,���-�?@��H{�
:D�P���Ӷ&��L��F�e�
H�WE-D�x�vh?qP�4 �i�53���&&��0|B$n�� ��̑P���n �B�T�<��K`�q�cb�5�<ɛ�eOP�<����@��q�tɐ�1��� L�E�<a���g�uR�I=Q"��� D[�<1�o\&<,����8��L���b�<i�����r�噂 �Xh���f�<��FGk`�1�E�&N����k]z�<aƈ9�\P��G�I3!ٰ@Pz�<i��ȭ4�`U� ��%2U���i�~�<�	Qv���D*S(.�\m��
y�<�������h�AZ#~���3�t�<��/E0K�T�àIS��a`�Ct�<�0��B�`]1"�ŝ �������E�<	v��\�P׍E�Sw�� &#E�<�����C{���g�:R�b�@0�Cf�<Yg@B^\-��L�5ޞ�è@b�<�F��"}tB�Y�F^ '�$�cNNE�<����fE���W?0�����@A�<� �Y�m�����EX;<�9���^r�<�6�fLQ20�\�@��`�6�Ew�<i��A��ˆ�$�~\xCq�<�U�5D�R`�G�J�g�v<��p��0=�F�>O{ؘ���B�,��$�F@l�<����Bb�q�H\�`O�88a�g�<IfeMt�,h
�cXTD�`ENTI�<��D&�0U�u�Kyd�X0a�I�<�Rɍl�0@�A����@�A�<)s�ܹI�ʄ-Sv䤤���B�<)Ro@.\��h��Æ�+P6��Bӟ��	g�IA��~��'�|���]'?�6�:uH��yRFԖ}C���1�U�lz�%��D��y	ˮ
���tB��Z�6�!t' �y��.���a�蒿J�L4K��P,�y�g�X�U�!�M*-��������>����yrA����SC�L��m�1�y2�W:Pu~�Q�nT&��̺�N_��y���v%8L!5�#9D���j�6�y�1e妸�&K֍-T�E@e�I��yre��(w��e?�,�	��ƾ�y
� `���B\�^��d��#=m8]��"O�p�T��bª_�>��Be�'~r7O��q�e�3]�ԑҤc+ ը0c�"O��K��M�
}�'��N�j�"Ox�J�I
9P�D �
�I�xP�"OF��ed�6_%�%�����"O���h�X��l
W�Гw�>�bG"O�u�� �P����N
_��iq"O�
���#�$�rVɞ�3�h�P�"O�e�A�RJ�s��W:6�ִbO��B�W�]�2)��{�����-D�|
�&���F0�*���)D���H7X�(��3�#w�ŀQ�)D��Qqd�%��xi��E ��0��2D�0��%1��T(�Ar��s�,D��r��'@�ؕ�ͅ���)�M D���3g�c&�C���)p����?T��b$�  �33��F�I~�L3�G�@�	Hp�G�S�f�`C�;D���4(	<Π���!DG�ByHa:D���Tu?ĭ��. �8�ⱑ5�8D�BS�ݛ%�e)�õB$v��%�7D���Ϸ!��}iC)0��hA/ D���Ū��1��bW�L�0s�=D�����6X��T�ל,�R,p��O���G��'���#VK&'Wn�X��	�RP8�'���$I�&nєe��ɘ(;�q�'�,�
6�\ 
��@���~.�%�'i���n��W1��f�ۇpՖJ�':�����Ԯu�-	�E	%j�UQ�'��ţ����Ũ�6R�xp-O���P�㚈���٘��0ꁯ�+U�!��7ZȩbZ�F���U��!���* ���������)s�H	�!�1�hݲ�C��)ɴ�� ��!��F9��ĥ��Y��p� Ȱ�!��Y�,�D0#��ۊUi��E��.3?!�d��1", C�Ǐ��t�p���m-!�de��[� �)�P�#%{r!�ʰ}���j��Y�y�N�1�ڊMc!�Ȕ��b�&ȣ	�l�P��M (!�ĝ>6ŘriY�i�V���	ܞv!�@�f�(I�nV�G��J�g�"=!�d�B�R"�B��I�w�:�!�d�V�Q�@F4�Z	�uIѣw�!�d�(�X0��$\�8��+����"�!�Ę$��H��fæLP��C6Q�!���k0���Q�� 輵��e[��!��R'�,]p'JC�a��d��_�!�]1N��oL)+沔�p,K.�!�;h� �s` =k �K��;>n!�dA�V/Z�6)O6h@hJª�&�!��E��Rڧd�q`��̜;j!���T1���r��K�0�!�KK�.H� �C��H��*	"p!�$Z�a��X�aA��~�"iU\!�D�s��}3pd�j�|i�g�L!�D�D�|q��.�.��U�� `�!�$_��>d��*�lĨ���]��'��'�f�	��!x�,��$�=w�%0�'Ĩ�ᕇ	�%G�x�ndK�mFs�<�OXm��pySL_�{Lp���E�<ybN� ^� ����W�
t�D
�@�<��Y�Dg�]��O�/5 ة$'e�<� 8��� ��,��E������JR"O��m< ��bB�F�V�� �|R�'n�a�h�X�$�s����h���'�$�D� �pq��*�� ��ic�'���Yr�˃Z��R��w`!0
�'ֶ��4a^Ͼ`�ˊn����'��k�#R����Y"`�nК�'�N���¨�a������'�>��Q�K�*Q��{�/3�zUi�'T�i�!�Lp���kL����;�'@�.57�3�,@d�5BNl�<Y1�$���㳃A�X xӊS�<�qY�H,H���[^��VI�O�<�o�Ur��h�I=0{�!J�<���+�@�ҪQ�
p�S4ƞj�<q�C�*�-c�^�������c�<QfT�2��a����$�n��!�U]�<��j�x`�d��G#m
8�{֩�N�<1U��-6^�pQ)1�`��ŕJ�<A�B�;+.�A�K��0�B$�JC�<����,*nh	�R���;K��EJD�<� ��$9h���ҟ�ڨ)��z�<�d��\����jÀ Qa�M�<�4�ʾ���ڿ�n��2A�,B!�1rn�k@	K�B�&�D�!�
���A�J�$(�C���0!�]]�4�P�i�U�L�TIV
w�!�D�6T¢H��l�697�`�\ �!�Ď�{�����D�1Lq:���*!��U6̄k�{�.D�U#�$>!� 8{F�P�a�I��5��@�!	!�$Y�7pçjZ*'��I��<!���x�",�����)���z�!�Df������	�F�WG��d�!��m�,�����3fM��D�~�!�#CM�7�W�d��eb�"G�U.!�7�aB��[O�F�1��*!���2T���ݭ���4��"O� ��L�v�
e;�Na�Ƶs�"OX�1�����b9�¤�2k8���"O6���/H�8Ԋ�C#L?��(t"O����ݟlR�q�'���U���@"Opy�a�_P
$������*ON��L+N~zI�э�#��k�'���(6����h�*с^���H��'�x<�B/�nv@��7��%� ��'��m��X�Yܾ�yw�H�����'�Н�6��!5���S�����D%`�t�J�C[R�rWE[�~G�Ԇ�d��lF�]��HAhF5;���������0���X�d��
5)h�B�I) �{�KX�0٢@,� C�I$�I�%���!�\)���S9��B䉕��%�8�X��,� �B�I� �ʉPw�M�b��ʅeY��C��Kj����\������eV��B䉃#��h�����t;��%��B�IZM�b����r|6K8df�B�׶؀@b�
D>TjԤ��X3NB�	��fM٧C+� ��l �"�B䉥y�4\��GY&�ı��	�m�$B�ɰ,$`Z^X���e�=c.h���?D������M��Y���ƋD#Z�br,>D���v���0�Z�/��p�Z���7D�� �x�gAZkKN��4���bD8H�"O<AU�6J/Ƽ+Afˈ]vTc�"O(z���!Ph��2�D��6�x1��"O��X�F�9���a���=��t� "OҠ�`��QpY���X�<T��"O4����r�L(���ً�|ma"OJ�H`�M��b|Z�&P����A"O~�:���+p�`u�W2**��Q�"O��J	�q �g�@��p��"O�e�oE�>3���� Vcv�`�"O^Lq�G�o81H5 ˹USD\KW"O04#"�<C�Ԓ����^RȤ��"O��&�j,�� oL<-O�]��"Oh�p��c��$: �W=65�AҖ"OLq0��1L	��W�\�1Bv|Bp"O��i��M�m؂I\
Be "O�9;0D.���*�g �h$�d"O���@G��o���wƙ"��Z�"Oya�+S$qb���44-��"O��f�==�X�{b��.p�-I&"O~�jЃ��S|A���$(�NHp"O��3�./R�F��c�#%e����"Ov�)�.����h�"FL%�"O������	Y_���#���'IJG"O5#i��zݚ́�`@t9�"O`����Q
\�q)�B��;`"O�"`�13���:êY�28�" "Ozar`��{R P#���#{Ĉ!�"Oʝ�f�3NӀ�:7J�d(��"O`\!��@� �z���ɂ=:�P0�"O��[�+ۖt(�iҷ�9̬�˃"Ophf�ɏ]l�@�)d!<;"Ot�����W���;�c:�pt�"O�M �%M��� 2@>��c"OX�󈁒(�j�d%�(O$>ة'"O��� @'.<cץ۬Kr���A"Oz�ґ��(4���A��0y1"O����/�&:<	���Rz����"O��DJ����s�� Dx�H �"O�Ik��M^,$jWǁ4�(�"Ojqw�5'���*�E�'j �C"Ov��`�ZCN�x�	�x�R�"OԄ�)��v$Z5�A*[
mpX�"Od=kc�٨c�49B�KA�j1͊�"O�����B���up��'$�8�"O@9[v���Rd�ŋO�x2�"O�����l,�p8v�˛5 ��S"ON�b�ٕ)d�9��˟�#&�)`"O����'�e��Ia փ}�F!��"O��y��Ͻ8�,hс��8�D��"O��$֖:�� @qB��vIt"O4��Fʗ\���с�: ƹ:%"O����t�FEA��]\)"O`�z���#�n]8e�N���G"OV	��T)?���w���i��{�"O�} q�Q9y�.��4�^�gW��!�"O2�#&䟋�YA"�?w^��""O�!��M<�Ȅ�Ǣ��Yx�S�"O,��f� #��=RbB+J���"O���BZ�b��5�C��J�H��"Ot�y�/^�G�<PaG4��c6"O���C� |�|��A��3$�X$��"OZt�g.�a�)X�d����"O�#]i`�
{hh	�%"O� y;h��B�p-�↕~���"O |��� )�SFA!Aeza��"Ot!B�L$7��W�P��Bm1�"OFK��/D��+���8x��@�"O%˧%]u�OW%Z�漻#"O�a"��Ɏ'�L��mI���"O$��m\�tz��b�-�>�2�"O��`,H��L��+\�D�,��"O%:�%\�'L�Y�D*�zD@"O������&I�$C�{�N�A�"OZ�QhI�x|]�6܎��UЄ"O��rA�O	=�vY@Ѓ��"'�G"O 8 ���)	�i:逰Q�����"O��t��B3mȯ�q�"O�8�#�E�.�����T���`�"O8�{�Aܘ8]�!`H��a��i�"O�(`ɆS3�$覆I(/��r�"O�|+7h��2���e��[#4�#""OlE*T�o��Xg��C��R)�P�<)��� Ȥъs�N�y9^��2�I�<�dO�.��MhF�	;�f��%�M�<� m��(�zQXp���z�6NKL�<ѕ�L�`�� QD�[%Wcd��EP�<9pdöGx������x!` �#�M�<)�L���+U�#����`��t�< ��y��0��ǂ�`��eEq�<����X��M��,W�r>���( l�<	qK�Xx!%g�_�I�"�r�<�C 364���K}A�\Ӷe\m�<Q�OE��@��,d�
a�h�<�'��q��	2��,C��f�g�<�'��I>���JC%@���&�g�<�l�'@:��䓤')���Q�_Z�<�’��T���m� �)W�<I����c�ܘR��]@�U|�<i�A)\	+$�
H}��i�~�<�C*�7G�$���M9\�Ud�<�DJЏf����cn��̒�*O`�<�J�Vi
��' X�.��rv�WZ�<9��F�����Ӑi��Dr�m�<9`�	�f�fu��?� ���a�e�<�v��	JCp�:s'�.9SxD���Wb�<QS���u�[��@�{f���[]�<����o�ة�ǡ�kU@uA'��A�<i�.=6F�9q�M4>Q7\D�<Y�Ɉ]�|m����1K�����_h�<��� d���[�*��EZ@� T��[�<��I� 
�%z�蝩Qؠ�5+�X�<��R�a��:���%k��`�|�<����e@�HH���mhu�z�<��K�U�j(�3��23B���K�t�<�4��78o�z�*�y�Q`$��V�<���0ΤD�@*�7Z��7/�M�<��Ҧ$A���Y�4������d�<��+Q�d��y���B�z��x�GEI�<���F��dU�Æ��R����OB�<��

�c}�hp��	�/p�ƀ�A�<�R��$������H�Yף}�<A��m��Y�6G��n���C*�N�<�d�vH�����?}��� ��OK�<I�'�!Y���)Ԩ�9�RA5�|�<9"��'Ra҈Ɇ�O�|5�X{'@�m�<)D�(�z=Y�%ڳ.��8+u�`�<Y C�\۠U����0l��R�@�Z�<� ��*�*�4/��3M�"���v"O6�kR醩uP�e�ǅy���*V�	�S�Q��'k�*Hc�����>F�YB"OT��r��X%� �`�o|�`q"O��p�0?j�r�.����"O��Kb,�3A��Eb7m�4)d8�
#"O���X�]_��^�p��� N�y��x2�a��#�!]�r��rǕ��y2��1��ѲQIY?XĤ��Ш�y"i���,���:�NQ� ���y­  i� }ك Y�J���{ǀR,�yR�e�Xt���ĂL���e�
�0>YK>Yt�[�Aj��I lo�i9t�G|�<!D�ʳ;�YFhq��騐f�ux�d�'���B� �~���#���2Z40�'6�4�c*�*)�Bd��̀���)��<��	�fE��SDI	:i8%�����<���Ӓn~Э�R	�&9VL�
�c�.c7B�	L�"��� ����s��.D�C�	eLҕ�-!G����6�(0��1��{�I,D���L(I�J���i״�fC�I�_V������Դq'T�_�C�	�w��D(0�5|�	��	�.
B"?1�O�b?�dEC�y�N�h��J&N�s��b���'�'*����"$�� j��Q��YC�yb�)�S6)��ܫ2-�$L(�BC��-�d�3,(�@3��˧@��Q��=0䰸V�(�IQ����FI&vdXJ�E\�}D4�@�!#4����g@�u|0�C��T����fHE�<)��`��g�<6P�����ID�'�"=�'[
N���Ğr�UQD��(?��X�r�i��n�X�O��>����Jp���`	�_~E�DF�+�|������OL)�ѺG����TT�l�!�"O��r�I#~�Z��.Z: ��8{��Oj��D;}ғ>Y3�)x����4Nǽ-���B�. p8�l�S��|�A�;`o�y[R�3h�8�/7D�����Ίe%�|�G% �&xt8D�4ғ7���h������M;r� &/ͫM�z ��"O���DB8
jX]q���+=|*]&"O�i1�l8!��� Xu���d"O�A��נS�RB�	2Y��e��|�%%�Ӻ�N�lۃ�
pi�D�ѣ�K��]���%�O$��/$$� �J%,x� ��ب(��ąȓ��q�����@��T+.��1��IO�q3X��sd�t����Q��?猱�����+��Q�'��-���H U��i�*8��y��'
b�	6�څB�Р�dP4'@j�X
�'�e��TFle�1�� 
�,�
�'�<������)�'�  J|�'�@����'V�����  HT��'�P!���#��! �/�2�0��'�Ρ� �u1��a�ʟ���Ԋ�'��u ��K�J� ��%/�.�&�0�'E�X���ft��ٴ���|���'m^t ʖ�Gd������ �P���%�'B���Iw���{Q"�4	����Xh��BE#B7�2ͻS#.dw,ąȓS�P���΂�*|n��h֨YR2�&�P�7�����'IQ>ᙄ�Tu;����HH"N�2-PC�*D��BDjG�S.�E
�I�Nb�ikfe*D�0��f��(��2��"JԪk�E$D���@j��݅]6"ڄ"#��h��ꓣhO2�Gx�핞;��A�0K�%b����!�y�K�Q��*�D d1� ͦ�y
� R@�l�%
2q���]6zhN	�C"O|țq�T��¨2�S�d|$0"OjP
�
bԣ�h�4I)����%��� ���Y�p���ǀZ4�5dx�LA��&D��Q�k �r�@��xi�Y�b2OT�=�HN(H�P�3�H9�L�sk�v�<QvCz8Y�ǯ\�NT��%u�<�d+�:�ڸ��.�c����Gy����?�� N�y���o	 Ǻ�bCJ̓��=q�(E��!�6��(�J,z�KF�<A',��r
a�.�HaH���F�E�<96LÝEʖ��1���X�CLFt̓���?�<��'&~�Qԍ�?�Ԡ�dX�@����'�|�[��C�hP��C�\~�pi�{"�'#�i�����Y|����s��}����<��h���;Ră�d�[ǓY�<�k_
N�6�𶩞�`��I�Q�k ���h�rX@OT<7\�%R�CD"�(�B"O�ك#��,k������0�p	� �'�ў��g	8�$µ"�/{M���s�&D���1�J(�pdۂ��6l���f�7��w��� ��򔮟�":db`��?ĤC�	�K�ܭ�SE��AO�T��i�'+��Ily�|ʟ1O��Ss�U�j���g�+`���"O�\*��9Z��Љ"C�U{lm��i�8C��\5FU�e�T
)T�#t����|��V�p�O?�ɘx��i�W�V�t��-�WK�:�TC�	2z�Ri:F ~( ���= �^㟘G{J?E�f��<ypB9%F�)W�	PL4D�lۇ�6'����̮n�=(p+-�ߙ��=���K�w̐��|�P�Bv��JX��'���1O�IA��� J�D���ǳS�n� "O����@�Ex8��F���v1���'���ūoR)6mݼ���[B�ό,
!�O;O����""�!	�r.X�!��
o�9��݉D����CB%f�!�d���d�@�'U�E���[�g�����	V��'���F%�(v��B�	!]���Y�M�"AE�M�3��W;�C�ɉB��H�$䜷R�0,�@Ι�9�\O��6�)�uYx�2�N�,a�D�%��@�FB��8���C��` �P�t��H3bC�ɫ����g����@6�%�DC�	���@$�
?)`�8��n���s��7�B����dͫ ޕiDę�%���8�L��'�Q����I��H�X�O`-&%���ܯd��B�I ��3C��� ��7j'}��"=�,O��|��A#S�~@��(Ğ ��@����Y�<�)&u�(�q�@� \W�<!Ư	�AÌd[r�J�n/�M��X}b�)�'m�fd
&��!��T�*w�$�'7�}��M��r��H�F����y2h�%%PőQf_�x�mz��#�yҀ�&v������N���"Ѣ��y�'��H}�żdߚ��v�@m�%Ɋ�y��F�v7��'���9��#BS$�ybL�8���i$�ϣ5N�8��@���O��=�BJ#]�4��-QD}�e����y��R&9�lQ#��J�+8�}[u���y"�)�YqI��d	� [5)��&s�V-��f�|��U�� �B�p�9:�|��!O�ꄅI�ZS�M�@ ȝw�����%��4(��C'Q�x����.��Z�D�2>��̂4y���S�? �ЋV�ځEa(�[7 M�"��h2"O�E�q�S�����ÏȬ8����"O@� ��2��0���v,��"O����IP�|J���Z*E`X�"O�"�A�S@���:d><���"O&����˄A�jQ��!2�	id"O�T1�"X;؄Hb!%�/b-:m�C"OPd�W��	u� ��õB(��0�"O๚c��Q!^y�œ�N
���g"O��7
�'P���	.9c:}H�"O��X����{(�:s (j(Z���"O>,0���e��b�Pq��"Oq�R�_�$I&�2L]T�L �"O0��k.e*-�:�%"O�I4I��s�Z��e��  �\��"O.L�d��z�,	Y �1z���e"O�IC�B�9$2Ga[s����"O��P�ԗ@�nI�s� a����e"O���!�8����Q
p����y�(�_�d��k�=g@�h���U=�y�؞dlh�Z�vEZ-���,�y�G����2Qc@U:)ĈZ
�y�"U�*W�P��jP/�V����#�y�ˋ"~rrԐ�,�?�>쓦�Z)�y"n��$m��lS�~�4E`&�(�y��1t�nh�Is�nP�i]��y�Ϩ6�H)��B��j[Ps�ȥ�y�o�3�艗��)j���!k_�y�)ثr{�����Z��X�!S��y2�"7^F��1���A�����ڜ�y�%�x^����k�7B��d�u�Ƽ�yRˉ�Whz�r�E�1��)u�©�y�#�'�LT@d+�<�b�fgB�yrDR�P��-�l�=T�my���y҆=j�=h�Ä�)p�(��M��yL>�<8�m�!�ΡK5���y2AX���C)��˔��y"f9h���#��x~��i4"��y���0Q�H�E��1J Zܑ�֜�yZr��xC�ħW쎐��d�xA,Շ�Ts�l7�Ư5���#t%HWX �ȓYu��bU�#"U:�3�dD D�E��~{`�iE���x_^@�'�C,W����3Ʋ����N<�����)c�4��y�>}5nӥ>Rl:���,2d!�ȓju�՘��U��� J� �>�^чȓ:�:�y��P4�fX{� ��q�ȓ+�eze�E:C���*�K��E�ȓ?�6����M�|h�E��Q�<���KU�E�� �h,��M&Ԟh��_`�Xy�É5=�����%��ȓ\A� �P��z��	rg�<1-�Y��(����I'U���g`W7G t��=,$��R�@�|%.�it��,K�F}��
s� CBN�=A����%�-u���ȓS����Ҧ �.	3��ê9V��=��!Շ�~�2��	��(����^&�((����T�!��S� %�!�ʯ��˵83�8QpaҲ#�����Ol�xX�+q��@J��Zj�#tO����#R^���9�!xĀ�x@ W�,9(��hO1�و�@|M��	�s��UH�D7u��u��I'M�Ʊ+'�U���!��M����{���U;ܼaB��̖��`@6D�\k�ȥ80	�Ȁ�|F��R��<��"�eXE�K�"�ԡ Bi.ҧd���B�A�5�e����#��Ą�S�? ���FΈ="Kf5[Vϝ�b=Nu�@���o���䖳e����T%	.�'f�qO�x	v�/]��A�6��y�h��'Ѯœ�N^�(�@ ��X���H��ĉ:�3eLF=��e�A�BT�����Q�f��$�%V?����2�W�L0$�'�6�g���&�PB���+s��h�я��z�,0�%W?*@��R�V���ʂ%J|	F"O�\���;3g�"��4�6�	���z'F̸A��SG���I�p�ۨwd�u&�k�w���h�C�X	n%wJN$bbЍȶn��g�4Ѐ�{�����1�H-��'ױ~���T��--�S��U xsn�G�M}���rl��3�D1ڗ痰z��8yOm��g��@���;RD|I��5+k� ���pN>��?n�(b��عQBvQ bĘ>0�J��`
��$18E�$3�����:t��#�h�P�E�?)0J�!
Ll|iG�u�R	�E�
%�b�cs� ::�py䑟���FHD}`X�bȂ�cf�l�Z/g��Q�F*�6�fK�|^Z�y��_<Gr@��%�9g���"���0W��Â���>1�,�e� %���_&W��:��P�jV�0?��YU�@*3�f�q�ԭ��	S�TF���;��<i� X-������0���M�݀B��-}]�D@�bi��`0��Y�f�矬i�bj��U�n�jT	�&�%�L��6(��$����@4dnd�Q�o��a`@�hB-Ys��&�X�ə��!{P�;�H�!!c n�R�yP�ܳ,��k��՚6t�'����ıPdX�XPe[�ldSg�O�`�13��O:N+u����4SF�۲1�����~�I����3d�M�;L"]Kp�[�
� Kf��-u�*���1����2wU��3���x����ݗ<���(ոT�l��_+:����Cd��C�B�!��Q���gU�p	4�
�20.��42�T�C�+��h�w&f��iыr@�M9�w��&
�9]N�`3Gu�F1��n��������3zT�!�Ε��������\* 4>��1�J�V��,�C��
lG\��$,�,U��KJ�#96���+y������ s�X���ކ��'RʁZE��1"�"�^�%�&59��ϢpK��I��(g��Ahrn���J��[�=<�Zv�_�#�"99��O!vH��I�Z�m�t9K�I�P���Jve���FF%��녪82�I�H�d��@/��耂&�j<�IYU�C�3R0Q�HP�d_��iJ��Q�4cE�4��V�c��@QU���3S$a���>Q5GJ)|f�Y�捝	<��m��n�:sE�<���6.:����͗n��Q���Ne�b#��򩎾a���2C�S�~5hDT�uB��sV�L?$4�A��!L@mHW�<e���#c��z9@bD�pO��֭S�0%��@��>��Uag�� i�|�z��S3̼�*�uW|���6�ӕwRt�ƍ-Q��A�eDUj��H�4?)�-�p�$XC�ui��D�dm�3b؁˲iµ�[�Rg�YD�>٤��E����N_�����O�""RU� 䝝2
�镋��Kl��bB�	C��1�N�[������%/@q���'9̬� 	*B[�� m
AZQ#����bą�lRO6a�(K�ܮ��M!I)l�9�K�?5�nIB���*�vMѶ�R�R�C��i�L��%Y,,���;��{d���D�6jY���M�6�x��g��*�"�c���(��r�\6���,��B��61�H���vhN�i��4
Hw<  n�	�T��`��=�� Y�� ���l��HDy�	��JI� r4�'	�P���`ڃ�y'^V��h3�]i�@��&T�0�Ah�{
�F�O��.=
�|��%lA"!��U	�,͘1����Z�,	�b��]�.��q�ز p�إ,@�$.�$ʍ{�P(-l�(A���;ꄝ�f`����O��b����.��i0�0�l�*�l��`	�*����#���]�f-��*V�K���"*��<P��ɓ*|d�h$Gb=��K�@�]��ɣ<��Q�^j�Ū���8�d r!#o���m�2Y�)��g$�5;�h�GmF���V�"C�	�~P�r��t�6X��E9;@��@G�,B��P8��B'�Z��3�Q�y\�R��u�<DHR��;>I睾)����!��0|�cT\������.R��i�ć֟7���?Ƞ ��	���d�I�/�Ѧ]���3,A��c.:e�{�"�t�q%�Ԙ���>̺E��<Hm6)P�2��*z��՝cи|Rt
�%5�����G����8��P�N1D((	<g�D '��Gр�#U�'���[�� tX���ƆD,D ��X lOIY
�*#�h��ZT@�� ��H�T�Q*1���f�E�A
�`�,N�OV�J��ɮijB�z����mM�$kM�!R	�g�J.ǐxRiE� �@��$(���+6胥�X�	���0
��p.Y��	+�L&д�g��bu.]��2G:��;P/����Ù�^Z��. (*��'�xpy%�����c(�d*z�`���W�� �A�L��J� >H�`�_�t�"�����f�!��E��y��ӫ]�"��6D��^r�8O�Qk��G�G������0�j1���5'Y||h�/\!?�Z� s��/��YK�EGC��1�#(��3�|��k^6#P�lS��֐�����."#��{�	�&�|%��	I�I�,�b�|�'n�*�$[��j˥*�L�K��Z<t�|�g�Q�M��D�¯T�b����q�O�~
͋��
�,�H�S޴~1�ع����u�DБK�x�3��]9F,��[�w�'��}���H�v��*��E+��{���6mM�i[EB��;�\��&��<-.�!�3��U"��s��o�L���"�9��U+�8�^��)�=.)�=�c߷W'�����&�H��RhR�A���A�'=�yY�9*�6�Zt�[��+����"�X���/@�����8S:H!%`�7* �Ԭ�=�L���"P��)c"1H�������X�B5:e N�6.	�T�<��'N� �(���=Jl�񯂯`�XX�.�5f��Ė�6�zViĦM�� �#��?@z��aoC�f�D��=p.\��ֿz7��S�Ô(�й�C��)�f��ؼ�8�<A�/C�,�ĕ-2g�bh�m���r�K۪w��:�*`��yɦ
O�!���*��qh�
�8O��
bKڨp���"�F+c�Xpq�$HŚ�+v`��\�2���P�U+��"�Nd��!c�c�+I1)"�(+R��/ 2�B%r֩���D�.X��oۃ2ś֌�@;���eK���7m��t���C>��' 
F��h��W���g� ^$�P޴P�0P
�:8��X�D���8���� �0����OH�d���U�d[dv��q�K6yÐ-˷D� x�ሯ�I�$�ѾhS�O��J�W�p��ܫ�h�{n(T#�j�ZW�H��H��ᧇ�u�L�$�"J�f���)"�H`�� BD��&J�$���C"(O�S\�������,b��Q��'��\�˒�(UҴ�Gj�0�68�3d�� �T*��9y�451ӯ9C��H���'f����
Ӓ3�>$�D΋��P�z� �!f�Z6q�0Xi���|t�n:�p���:J�1eC[4(L0���3�X�:P�5D� ,s�'>��!�T/ �"Q;t+@�9��C�]=����h�~-06d� K ,h��3���h� F�)8F��c @��z���-�Of����:{�)�*N��P��F�-0V��� ��h��Mn�	4��2w3�a��U��."p�ΞCQ��ݖr�J!	Al�#���$�;�k��h ��ړ/FJ��T�qԐY�hNS��-�"��zcFEk��o��@Heڒ,G@��g�Դu܄u�F�ipr�p�dͯ>� �yc-��m9*h���tI����2��S+�;H`|Q�b Q82/�a���ɶ$��4账֗+�KÂ�˒xc"�
Loly��'#�i�l��hb#K�Nj!Ka.}2��sգ����>����2�>����J:R5f	�w`�Ml�I�Y &`�J]�vm��0��ؕ ��M�x �J��jw$�_خ<�4��!�ao�*^�6��ɦS��H�'�z1����$�@!�rI͡x�j�K��ף~��!�I��+������580j�G��q¾�����G��T�C@�!vT�
l�;=�
�X�I59��DA"{*���B�T���Ŀ��y����<��M�
�*ӎ�#s:ٻ��ޔU����_Vl�%P ύM�Te�L?8d��[����� �%Q�����&�p=���.�(�Ʌ
�
�.dJ��4.}��J@ʓY�� �OB�5*B@ےGޯ�&��J�
�&pb��.y��b���tq�@r6 �q�1@m�$��x�ˋ%~���m�lܜI�!	ධP��I߸��&͈�0��@��
'p���m�iׄ4����㴴@"�O�|>X�:�)U>�J4 `\;8�aybL��6yP�@P���s{���'�e,�9�ۏD�R(���1�Q��$5��P�m� �$�1/�f)�1	҃[G�Bb�Zf⌞Ql�8eE�)����0}b`
�$^��w�� F�T���j/ ��X1��>|�f=r�śE6,�q��R"DG�H�備8e��Ab4c��D�>�D��^+��[ϓ)�����>}b�;T\;`��!�B`ϓx��ػ�AW�G ʵ+6���-�0�w��<yl�{�"}yۥ.�v��3���3D�[D쟠B#���	T~���#�M�+TP�1P��d�"��m�n邥T��P1Y|~H�q�	6|��L��*�]}��8���L�'���.�VD�N��g�l}���a��r��'�)��˂�"�8�GљX!��!���RBX-3w	˽G?��{5�Oy��q�D��u���$�̼R>АT'��QG^9�I�>A0�'�@{�(��]�|=�N�ci0M�O��R�'�i��T��F_lE zeK�c���,�$n�Y�V�J�:�`�s���'Dh�%����/i��3�׺r2�H$晣9[L���iK(�լ\D=�t��#|0du�f��\�ҁ��1KW0���V�l@�E��	�FiKG�hԲ`�03 �m2v!J*��q�D�B%��I�2%���W�Vm���v&9qجSffN�+TlR��ʪlt�m�cg�:dg���%ףRd����Gڤ?|�=*Qb��v$΁wM�a�AϜ�9<��Ѡ�-O�C����၁��e�@[��	L��usTO֊Q2t��gIj��OX�A���8�MY&EmHa;��H��e[$O��1O2�$#�A�(�z1+ņ_� laƓ�T���	�|i�b��%�t ʀhS�\(h��k�(�bPp"	G�( R�,A:t}\��7�#�&�ڢb�3{��{�g�
{�,����r#4��@�ٱq� ؃��}��k�Bҝ3�=[��-�p��G���w(,����w�4�۲���{��#7B�U��IЩ%x\���Nb��D�M$�Sv�YD�i�u��h����=d�M)�a]�_�>��f��O(�{&a��G�q�J¬l���¼f�L���dϧc� {�	L���(��mN�t*�- ��<�F���Dt��FG#H��M�@	�*4ǋ�9D���4�	���Ғ A0Ct���äثH.�$���٠/
 Gxr#��[`� �N͸w�zh�d��1�~҇��ui��s�c�:�ՁeZ/5w�G�]�C5 P��!�^��b�����J�KZ�{� yR��Ǟs�
ma	�(&���>��m��gp���P���X���K4����HϠ~�:!���o�3�ۈM?������x�(	�� ����#J)������¼ ���&�,ժ�- 4$⧯Nu�D��Łf��4K�I�u�;���f@(J���5}e2�M�[8��;�AE a

h�w�'SZޔ����>gF(B� �7xQZuE�;]5���_T��e
/8G�@A\��x��E�+P�кd�~2���`���h��) X˳oH�Lh� �r��0��uN��>���dF��.�te���	\�t�/��Jc�$��������X	�4K��(�m�0T!3@C)e�l�s�'7,�=Aab>�:&iW4:�E��>d��L��e� �^��N�hD9�m^�MM�̸B�ΑI)�!�&�$��X�Cˢk��MZ�eвHT01�rmG���X3�9s]=��eR�*�V(�K�0�ԥ[E��KS8��mՁC�����;w[9�4Kі/�>q#a�E�� O�p����{�G	9\���:dE
�J�Faq��58|��ӕȜ,DZ�����2Q�1����z9>�Y0$I;6��S� ��	�Ԫ���C��[#˘�S �%�@H �0.�a�dh�=@�fP�4Q��g���VȊ����e�#�|�ƴa��-J�b x��P?5S��S�_/hY��� �2��t9���9C��uIF�)(��k��ؘB�\ r��C Yȅ��e�+��)rw�J�3@O���1
�$!�zA�!K+L�p��K_��q�V]���D�7���qJ�$&�da�qEK*A�\��+ݩ���A0J=�DR�!�?&mbE�$ 0�t���0��⑧W�1O�<���ХR��l� �2/�~ݳ�bH�PΤ�W(�T�q�RM<I"�p%aM�}��ܩ���)�z٣BH�S°���[�A�ҍ׽���`��AO �A�#T2F��P��#V7HŹ�+����l1Ĥ�"�#���(� W4k��"��9��x�2�
~Y�fʀ*�ȸ�@kH$-j��I��6n�
��"��
��p�����#q�-p��[�O	T�t�"B\��ł�'�a���XE� /(�yI��/w��KΟF��b���[b�h��K����sa�I�7E� �@W�Q��l�@��?`��1���$f�H����k1F)��8- �yu�Ɯ8��3#\*+�����Sxv̙�A�9Q2Ʃ��O�Y%gF:���(���F�X�^�(Vi�s(�S+�V�~��E�D�f��`g��<��U�>�dO-c�P����i�?  �#sČZ�-A?t�ĭJ!���~�a��+��k)\�P(�@�%yΘBѽ��eB7*���:Ի�N�69��k#.��]� ���ί�O��eO]�lq9�&j���a�[����F�k�<A�ʘ�gؐc BՌ#	b��'����F܂�japKT���sEl?��.����Z �͢�U6f4��'v� �%`�즹ڦ`L'g�Ĳ���g����t��9Rtq��FU�^BP8��Ċ0-2�3p�W�mj\��5$�boD� ���'M���eEW4d�4�IEg@�~�d��jO�\QxU[�OV���9O>a*�.��ʼ;�@�w�:��S�O�G�Td�P�L;r2�i'��j�����-ͶG.Y����v��
�D
?O��|S� RN�v�A'-�$O�r�QM�AL������%�Rǔ �L��LF����$�h��=
�H�*���`��CM��`��|4
��qFSq�<����f��\�Ћ�_(�l�$�Qs�m��9r6g�A�Z#}�����[������NF�ح���n�<���%
�0��ƍ8:S�
�_!�U�� �@�S��?Y�e�6r\zM�#!I��e���c�<��$(G���b�C�1�����T�<����
>PX�돹C`����z�<ɀcM 8�P�0vQ�5���Y��i�<�������d�5W�h���m�<Y�[�8�t!��ϓ�j��XAJ]�<q� ��uu��[1끰 ˞�2 �q�<��B�0>��aQl�/4��c��l�<A/́>�DБċȧ������n�<�������VA�
YĮ`p�L�f�<��������CdH�	ؒ�z�<�0�
Wp���#X�� ���C�<�mD����x����x�7J�z�<1���P4	�s���I�T�s��L�<a�LO9`�Q�ጇt��9��J�b�<!�Ӗ~r
�C�`��r��(BG%�b�<9$&\	Q^��p�kظ38R�@3��^�<y�i֢HZ�#�H��	�&ѳe	�w�<��(G+~| ��C�1qIz���Fo�<�F�^�V򀓴�����f�<A��H8�덿<JX�����J�<	j�R���r'�Hx(�qE��@�<�p�	i�"�Ѐ��a�\�j�b
B�<y�)L���)Cщ\�O��e�SK�~�<�GnٖV�N����}M�,
��a�<y���s�B��Hj�"����C_�<a���4#��}��U&0�$Q�6�V�<1��&h��t	��ԉS��x����[�<a�˜=�qF�ބ+�Nqb�Ci�<��H
���m���QE����B�<�C����"!9�K;Q�.��W�Yy�<��N�0g dq���� @t�<�ub�T� 5 ���)�9C"�p�<�5�!i>���u�K'R�
A{�$�p�<�V��� ���E)	��*怇o�<	�OKe`�F�B7
�x���a�<��-ʳ ܞ�r��;t봈r��3T���@��%W60�q���!�"y�f!#D�TX��<vV��vcM,l�Rq� D�l �j(��0��FF]6q�U�>D�l�4�_�(l�Db�N�M���A1�>D�1C�����*p�!j�e��a=D��R+ǦH��+�f�247Lɛ�L,D�d�C'DI���P��"Gw~��!D�ܲ��ŏS?uA��P@n� @�>D��uǞ�W�n�S�;II�h(D���O
R �J��R�f�\�׬-3}*�{��m�OX����]X���Qa�6*�
���>��	0���0�Y󣗫[��+���Q��'�jm[���>�NK�zp�d��Q��r�j�uH<���HUdLŨa�>�u����\���yf�"���C9|O� �#A�S26�I��(?nF � �'�$԰w��"O��1���}��BL�b/������4\�0�a���y�C�F`R,`HQ�Ka�%��3����OPd���h�J�OtZ(Tϝ\��0p�g����

�'yvY[uc����4�c�*![��y2'�P>�E`�+�=G�:�eʘ��Ϙ'��@��W�S=��C��&���{�3���;ҡi�|�Si�'7��D���Z���b��+P�Y:�H',l:9��펬7^�z�� �������G;�� ����G9��kY�4|�7��1Td8y!� ~r	�fO;�X�"��()��͂ ֥"V"O��
��Q4.�L!2�*��<(�@��E�+�M��Ԣ�±�s�L6mR��J�O�4��	oq�V�k�e� 5c�RE���z��`�1$I�	�4Y#�5�)�'p�n� �W�����<(�8�۔�����	����W��z�Ḧ��Ֆ9�����DJ�ت�k4�O5�~�7*Ĵe��
>G���I�h�i���'L�Z�ԑ:qY�)�t|k��"{ �LK$��:Z���S�j��bB�ҷ��Aۊ����+�	w�a���qƀT�d��Y���S�E�v$�!A�D	�����FX"H�t��X�~L��p�5!��9�kI ����m6w2"h*�-f!W�i�qOz����	�TQZI�va���ʐ�O�"�Vic%Y
b�L��)ͫT���O�W���H�̄�ڌ*U��|��LE0`.��؜w�h� ����up�D�'vh��J�u@>����~�#?U5l�CrIՍ���OP٘QC#Z;Z4�� [� ���+$��V�. ��D�M �m"P�ʼC@�Z�¡_6@V��i�س���Q�R��
�4�4CF/_�\��M�1k� �@�SK;vܢE�D(��+O(������X �O(�.��4�F5w+�h ��$��)�#Ϙ�qlD[��ȇ�b�[R�3;����AgF5t,��ֺ'��˓OY�x|\s��X�D���2��<�D`PiȽ2Ռ�v�z0@�� &'��|sf����M�.�c$<��������d	 ��DI޺k<�!���].$�q��ЎL��7�ǳG�X����1����|b���x1z�ݏ;7
1�E�̜lH&5�#iD�г�\!����`u�����ħ'��\3�M«uhj$���Vt���\H�T���A���!��צM�Kɞk�P�ص��:7���RǑ_��I"b��vJ=�!4!��Ale^k�Nu��/���	AO>�P��4�> ��/(*��+S�ըBo����E��	��$!���Q��u�&Y�*VrM����6���
-O�T�U��)#H���#*���D�/����pj8�ʬ���(����%u\��E��S]����Ö�rBqzr�>�L]��� ��[AC*ȸ�$�GMF.S�	Ӑ��a�H*EUtQ)FmHw�O�j5 ����q�Ab 	��g �Z�	�T�Y '��%�B��@P)V�~`�a��p�$i�d �2�wnr�	V��n���dKg�*�!e&c�XU+�'Y�(�%	k�gy�FWc�6TвN�y��Q��ciʬ�4nC�/�n��ghߧ3��fL[M�"d�B����q�H�@�@%D� /Ʊ�B�I�{	����� T�JP9��ܚ+�ث���)���W�̒UX%
��"jܫ�H%U4Pr3�F����&�|�Ly��e�4�`��!�xҡLl��Xq��<{���	�8bD�5Cף�ȉ��ƛ{��.F$��[�C2=�q�'�m�r��"�>�0����Cp�LV�ԋ]%��k��קW��8��1��W�V�� ��Q��ȟ���#
��h2ř!/JG�L�A�.8���Q�� �҄�����S�Y���4K�/HB�l@Q1�bEI��>c"�)�?f���`��qO��a��in�ɪ�7p�3��ʤP*�%����p��  �9 ڼlrEB�	�01G�^�?`�S"-��V&qOD���`���NB�%�Be�V�	I.���N��s�0H3∕$m^��T�U�G�R�qjT&bވ��ć��L�9�IĘQ�PMb�-�p=�@�2|h����BW�g"���#�h?Q��G���SqDX%(`�ؽ2�b�l�b)����胩�(���ڂ��� ��J��!��g�<����'��	��S%W���GN;-q>U"`��Q$i
�~���GR�����%�T�̨�.O�����4.�!E�G!K9�� ���z�����3�ΈK`�įp��;�m��&��1Cj��J�2�4{���@g$Հ6`X)s'���[/��
����-xW�τ�UP@�:Z�t��r�I�Q��{w��w�`7�U/P:PUl��k�>�������ʰ��0Vz %�֫:��O�yp_JZ��$�A�r`*�mء>�����·�!y�d�&`ږ5����I�l�2�'C�D�jLzFm�:����$N�-$s0`)�I�6���2�-k����2No"l��K��ᰤ�;k�LXCAڧ=_$��T�	
A�ˆŶ0�a�󅒿M��0D��k�FDK�!�$;R2��;m{��(A�m����.�=2x�'�!cp��I���eh�h4H�pa`�r�TF@.A��h��V����O�I��W�͏�l]�j�#���qQ�٭=������6��	"p��F�O����)ŤN��؊�"T��X����\=m�TD�I
-(/Bq�A�Ũ{-�����&J����B�Ԧ�N��"�>i�򐈃�2P�@�D���jf8q *�;@�S��ջF~钦S�'1�40E�Ĝ"{v�����t�|i�,�J�^ H���:Id� B�G�`�����ꅁVvn�ÔFO�r�xq�4V�@�@ꎍv��0���R�1�|�0���jo
��$�JS�'s�8ɳ-�-2�r��b�9ih��tG�=�P,��3\]�� �e����FE�l�zh���~ �HA��
�VfH�VM��0^U����f���*�ƅ�n�4h�g
`�n��%U-%���'~ �06��Y�@���ʣ(8$t"�gd�~��enխ$��Rョcy�}�˟G�m�D�'��S��7~��)�:J@�9���;7,�i�׫�F�q��D$���+d#����c�mG|b@�V�S���K2<�Vė� �pK��g$���oMj-"���U���J�y� y	e��7L=�v"6;���7l�rV8��cԲk%P�<�f��7?��Ӈl7Ya��r�R0`%�MB�OS�G�4L��&�9+d*=s�b��� �3$�ô]l�	�g*�m�R8A�6P��ڦ.	�݂�Q=tx�k��K���T�4�S��t� WΝ<7ȁ�0BߧJ�,A!� ���d�?DN� �����xҨ��nOx�ñ��˦�P��L9j�	�|<��2�fL,-�Y��4��XP� ����ʆ	����-iRh��Z#��8E�.5	 �^�#@44� b�,18@�S4ґ	��b$�#�����#;�J�D%�UZPD	���y��<��D�KQ>�eD�n����l>���C�#=P���4�q�&ƙ0>��E_;d_8�Ac�rfv�a)O�E��$ǏhK���E��M{w�O#R�s H��WP!��,qL����pX��Zb�0]��qt�s�<ac� jZy����� 8��6%� �V��O��<P�!Ɂr�2eCrk��jWE��� hW嘍H���a�Jh�v&K�HOx`�",ƌ �jI����>tsE�$.�xĀ�iW�U)��3f �!1f�M�V醄,�x�k�]�c �F�L<.�&ـ�z�\���lA9Ei�죢�R�|�ǨS�	��L��+�8���� ݼ�?� �K%k�2�ʳ�]���CH�:
��l�˂�:��5�A@�?;�(��@&�>�����bް5�yɡ��.Xg���h,�#�P�!\��F�>��O��Qe�6!���@���?�,QKIP��|3R�_�UR8q𰃋0����(��"���hUES9�S�	٦��$۶'2��7�
'i�]��lI�y[b3LO���7&�X���V�Kq0R"�W[��S��;TbE��g�#%��Y允�<�HܩS�w� 9r��~b�N�),����U~�c�	�t��ی�MJ`e��>\� �g��L/�ؔ��"VQ$�1"+�a@kq�>8z� j%eB�#��6��h�ɔf��rR�X�R�R�y��O�ġ�LՎBX�	���Y(���$T�h�f/QEj�82�ӑ6p�9[���Vh��X,���T�y�N	�,̦/M܁a��@�~0�h�$�p��d���]w���G���JF �ܟ�OJ�Jqa9����B�r�hD�����'�������(Z!>`'!�?SZ,��̦�3K)�r棍~�"y�E�ِU�D�2j�`<����J'Ye�zR�Q�-��v���)!T�3f���@Ł6�8��ccQ�'��\j޴G;�( ���q~|��$�IȐ�{ԃ�:�`�0�.��W�.ՉD�t�����l�� �0��qj�'T3Oh��J��=p
��	C
�avR�D�دFf�3� _�3��Y2&GձK`��R�V�ql��� ߣ)ĸ�#���B���)�GQ�a��Q��r=S�,L�p�쳖#�n�x$��b�d��+��m2�V��5�@�av@�}��c�o�t8Hc���g�d�4�(E�
��N {��Q���E�XC���7�@*�r!"��ڡ\V��I�,p� i��Q��z��e��;��y�D�K��V�Zoʤ�a
Yx�@
�G/\��E�Y�/��K3��9 � Db��Y���тn��6~�aB�c��B%N��5iY*��+��46�q�aF(U�X���nW!A08��[���a��F�> h�E��bJ p�!��~�	����Z�0
����MK�ON�xD��k��È P�®!��`3P'�n "��\�y(d8xw�*M��e��I�������8vSFAj�l��_;��3����u뢢�(0�kE?<���@�]7(#�p@B�c\����Aȟ
��U�b�I��Ml� �,đ��U���D�z�"*��k��ø!����	 ����`2��8@� �32�,/��2	��/�}a�M�t/��"�H�.�x���4;�<�bY+��<��дnEq�AJ[�[�Tb�� y��D�5��!��)A� ��|B@��hNU���Z�-Ȅ��HV�f���x4H�
%�	7�Ρ灇�p��R��{H�T�B�ȴT�� B&n2��Q��)��TK��"!g(�6cHJ�\�∉6S�� B�S�h9�0����*��q�I�^�ލ�C�	n12��	�H����g.U�iT\�	DH� ��Vǎ�2�h����ÿ!#�����h{��CS/�
l� �c�"O�^Ԁ����=0�b��m�|̓>z`Ea���l�b�3��&2UĘ�'��Ո
LIn��aGGέ,�n��M��y������K�up���2�Q�~U�h� U���Hq��bx��#��$�HhňK�����b�n�a�"&-ֹ��#��Qh��=r�"Rb�l�)AҌ^�g�v�C�!  &�6m�%��y �M	�ڑ�S�F��$�Ҍٰ`���$��C���� Ȇ`\�y��eh(Pq�<a�T`\4JQR����'���+��cZ�a��l!DYH�N�c�����(�f��4mR�=��������.���`p��1��}�����`�@S&L$L�� ��,��D�V"�7dq�6�^܁ �S�m�P� �M3B�h;��$ƿ)��)�jK�8��@�-V����	TX��q���a�n��g�a�5e�qa0�9�+�*}6�maPi�D��k�jS6in�"�'�r��)Tn�:e�0mG}r�F)P��I�C �д�I�����]f���4k�!u&��4��(E4v`����H��8'���OΒ�B$c�7Xl���d+��yW��Mі05�N<U��(t�!��'�*�tb\�u��9A*�]�'(TR)��6���xwN5	}�X��e0-\�3�؈t�L���*WT%��ž2����.��p�l̻M�H%W��~,��� ^���H��t�!�q!�3or�D$�ӷ9y�P0�%B��Uitɝ�F��������< q��F��D�	�R�iQ�Ȁ�P|1��1C���� 5�	*IҔ-H"Y|��"��U�4��ܴ�L���N�_,���VP����|�����tuhUi��n�b����Q�:�����-��`���G�&�<!�Oy,*�ъ{�a����
�&Ӹ����P�]��豤����1�Gh!%�E�M�ORDP2su�Ƃ0Y�����%��qGl)1�iO�X�JЫ�i�&k�P��E����h��B׽zr�����_NV2Q�0Z'*+p�ۧg,{'؁UǯMkp����!4z-��zcV�4�fp�P���pk1�O.=|ir��
��(���I��;%J]��X�sĄ�f�P=a���7Q��=Z�o<AF�MA�LD��mU���B�j�"Lߨ�R%NБ:��*��yT��hp�.x-�C!�,1}r�ş�"�J��V�9��rcgF�}\��XH<��d
&s�>�)6k�#Jdq����oK�LZ7�Cd�:<cDצ/>"t��
'r�"�Q�+C�"J`E�r���uIY���zT�������2s1����K�B.���Hٹ"< �<���Y�&(S�cY�
�"��&��-��7�}�p�N�d|+���
~x�3�Z'	n�D���!jj�hq��5�Eʰ�td)F�o�=�oT�d;e� &��fb�`�@�֥
�r<����z�@A{6C�lti���n�PM��'�[g� R���v�͈�zy8ɠ�Y�$�$�b�g[�O�Jy�W��2���{Z��%ۿ� z 0�/_�1P��'��#R�!�� ��Z�%��,]R�_�76`4hr/�)3S��'5er�p��8@�Z@�j	�,A~�0�,}"�[o� ��`�B$� ����A�8A�Rh��I�.Bx�H<⧗/hu����j�==!Z\���M%tb���H�-�2��C"MY�h��/iv����ʃ�?'T\ɴ��٣�q���
���U,Aw��$&���@7.��4q:�	��S�w2`@j�}¤]�� ʇ��5���[Ԣ�2x�ɋ6/L�jm9�?F%�뗁Y�m���D�V����sdb�1}�ś^w�&��5�-}��З�/�.]3A�*� 镌SM�'��y��O�	\�Y�V"J?@h!bkX����I�/���m3�d[2��E���R#��D	%ߘi�5�J���犉ɲ������\^�CSa�% �M�'ٟ��E�U�4��D�?+S��q�%!Z��n:�/R�>�2�������F� \�X��i��1����]l����+EM�g̓wh�t0�'�%�b8����
'�
�H�FNGr�jrOS?�e�%��<I�烷PGZ����[�r�����^�VtE�E� �8��eJG�.��zbcS\�&5@��7:q��X�(��e64����Ңàd�S�J��¤l�C�
�e� Rv�'����AM�gt�18���eӖ�IE؞4(��n��)�࠘�.� Q�a�˺2� ��!�Z����'0U�d�_�g���'��b���To8=�d��H��҂ J �l�;�� 5"Oι�Am�l5�0�揊-,��c��+��y�F���O
��bO	5|��f�	��`��"OT��F���q O
��%V"O�dk��Am��!i@ Ѝ\S
�yP"O��d�ԓv�p�/Ȼd�t�rC"O@Q�ɍ�
�6�y�G>s[���R"O�J��"6�Y��.MF����"OV��v�Na�e�5g�k�F��!"O��$���6�ҩ�E��;O��4`e"O`I3�
F5����m)Y��I�3"O6 )���J��B�l�rL�٠"O���䅀#���J%O��Yj0"Ol�5/�̨��0Ǒ"tŪ�"O��b�hд'��ۗG1Nf,U�u"O�򷢝*J��� V�E'DLb���"O1��쁺?�>}qn%a���"O&\���ۮe��Ŋ$��#
j�i�`"O^%âN�,F�B1e�ݦ	�%c!"O��J��B�ad%+@�C�|��"O��#�'F�)����%�H� #��@c"Oa��lQ�N]zb�ʄ[�\dK "O���� ��@&��Q�剫`�r�;�"O�1a$���1��35Ò�~�,�Y6"OB�P`��"X)����[�E��zq"O��c@�; ܖ�����l���"O���K
�cV^-��f�&+(�"O�E��g0v�Ve�f
V�&t���	�.�k�O�i�b��A���ҳ4ܳ@Ø���ЙQ"9#�a�� 6���Ȧ2#�O��ӂ��C"�	�$�/&	���:,834b�Цar�%��"@a��E<uK~�Ya���U6���.]V�[�ėڦU�G���^V��S�O�ij�l9>S]�ڞ�)�w���i*�G�#k��S>�@H�"=?��TkCf)���&I\ʦmY��G��y��0�&�G��e �TkL4���:a^��7KJ�E��C��d������z����OU����,�$H:���_3��9G5O��ʠj�$#m"����4��{���|���C�u�ʵX�#@=7<��.��?1�Y��|�����&���3����f�Φ}����}W�=�p��?�.�)�x%��g�}P|�;`U}x�@2~�|��<'�N�=�O�HH۶dY����v�(1R�TJ6��Q��B�Qc�0�ǧ	�f,���X�NDإ�wNUk��)���0q*��<s��\�h�B�: *R�K>��P0Rf i�.� Q���C�N��I�<��I��uG�7<�%�qZ))���򁍑o���y��v�6%�7^?�5:��O�������FiK�h�&"���z��oݛ&B��m���T��_��'Q�J|���L�"IB�UMT5n���ó�M�@	 ���B���x#���w�@����-F�J狄�Ni����J$m�J��rD�<�7bl>��!�*Y�x��$-
	Z��HD�1(���0<y��"��`3G֨UҸ��`bS�jVZ$�`��tss�&dԮ�@D�6�nx�֌���)��CR�k>�H�?O���w*ڂ(=&q����"~"4A��$���ɚU;ĩ���ȾB��X�j�j��]�0|� ^��#�߱G��e�Hò�r���8s�sԑ�`���!�pk�F+3�x�J3&B���!A7fX�IfM�4bW�#�3�	�����/�i�l��PH�<�`C�	�\p��$��<5SlLbE�2�"C�	^&6�:��O"i�:,�E�B�F�
C�I�2A��@�.5m?֜C�\�3ϠC�	w�%� H�+|���x�A�4M�(C�I�r^=��J��<�|�#� ��DC�	X��R>H|����Ռo�C�	�8�q;4�'I�ts��3Z��C��&.0�0U��;[f��SK��s��B��^��`ӁJ�T�*���P!M��B�	�f-�����],�����"��OƜB䉍g����AN��)�V�����L�pB�I���� �T;2�h����3�hB�I"8	������Y#N}!2K�%@B�	9�ء0w-և.�����
~�B��E���r�f��xm��&�� ��B�IqX�2V�� �4���q��C䉈T� �������f�`�՛��C�	�K�rԱ���7�Vu����7VC��4<!�I����X��5f%�%,�TC�*,����N�� ]�$a�.�bN>C�#�h��9`��<B!bE��C�]�����A�s)���%��I��B��?:^y*"@�!5bT ��^\��B��
f]�H���9Q~���Q�SC�	${n��%�L)Jѡ�a��l�C�I����SU�<i�*YZ�MΝ9s�B�	C�p��� ��pk��(~P�C�Im�n���"�i�0��p C�ɔ��l�D��HI� G�Jn��B�I�L�I�� Q��)@��*H�B�	[W\e��-��D@��Cc).�B�	�?�HX��P�'���aaJ�k��B�I�¦�j�-_���@];n�B�	� �d�4�U��B(�0�ضtbB�� o:��SG*L�.���iWG�^B��),�}h�C<ye���'C>B�I4�����CÀE��q��l�>D�B�="�:9�u-ڥQ��q�d�]'eD�C�zɂ�ۣ�ۣ-���U,�*-BXB䉜&ł S�&I:y��kwHPc�pB�	;`��l0*��H�\@D,<}�6B�	4+U��0c�? �Ȑ��*?5B�ɊQrV� ���(����/[6��B�	�P�8�:�7RzCKi�rC�ɨ?��D�H6/2�ܺ"�U�D��C��'.��!�j�'��B,$|��C��CM@0XꟖS���QvMN�V!hB�I� ���N�gu���v��Y�rB�b��ZtG��=]�yS�Զ+h�C�I�*��Uk &A9	�<�#å����C�	��Y��,��^��c��N7�C�ɭ
�Y� M�t�`�KK?=�B�*Y��A�Ø�Jx&I���ʑ��B��$"𤱩֎��y/�C@T=w��B��6tx�n�i�(qӕ�S88QlC�	�y�^@����Y$=�U/�z�.C�"��h��e���P�~�C�I�+�8���O<i�XI���/\�B�Ɏw`�ī K�(��,X��<�vB�	�+�tE[�N1������jB��&\���W�#h�@$+�$ݘoB�)� ؝�2�ɹ/e�*e!���|�a�"O�|���rf�DAt���j'"O�Y�խ�A��r��*�截"O���gL�6�
$af�1�M""O�Y�F>,&��׊A+E�G"O�8;��ڬ`�*$�`)m�"O����m��<�@N1�fL!g"O�l�G�L6[ǦHʥ,�5��-��"O�,�`�9�v�!�U?W��ع"O�DRRkL.J|Э�"�i<2�"O*)y�lׯ_�"m��]t0#B"O�C�ꊋ,�.�#�R�x���"O�Swf٦_;���"Ǟ ,A*�*�"O���AF�����u�(~Ύ���"O���V-8��-��V���2"O���
�N�����*׈^�B=+6"Ob�!O�$Ѯm� C_�i�7"OuC��:E���"YK�9�"O�@P�͐�)��ዠ#�N��XP"O��҈����h�+C��08�"O���B@�B�R�� EG�#/��h�"O�����?�0ю�� @�j�"O��2Uo�ĺ|@�׬  zG"O)p�U�]`��G��m��=��"O�i;PcŎ/s8�iWfX�E8D"O��:�j�P�x���EJ�+1�a�1"OƩ�t�_Hx�����d�d8�"O.`"a$Z<;�RXP�H� 0�)�"O�ثr�Ł''�A3s�X�/��E"O@��gX8�,]%ԕ��"O�I7���4�:!�V��}�p$��"O�@t��#f�6�b�A�%�*���"O�uy�k�'%$��ɖ�
�`�vS�"O���F�F"I�&yⴊ	 J �r�"O�]�E�ź-���r��PB�(y�"Op}�eě� J��"C�?1@T�r"O�������ا"_�M��肕"O��/�RZ�+�l�0ep�q�"OF2�bN�w�I�*�+)g<�"O�!v"�k���{�NE45@���"Op92���E�,¢�˴HI��"O���Fv��X��;G�p0"Ox�FHC�nL褨�"\����b"O&)��"�-L'hG�4z>u�1"O<b !S�{D� �Q
�1�mJ�"O����I��<��4h�II5p��s"O����+d��iŹ2 Z|Cb"Oxm 3N�3�����!*G�-�q"O&��&���/#�dRt�E1�Q��"O{qф*ix  tM�"vb�"O`�B n@&r/����S!S>���a"On0B0MF:�<�B�ҟbM�1"O��!�C�?��5�%���HE"O�:���R2�z�MћTNY�"O�]Y����,w
!�pL�i���r"OIB��?��1t��>����#"ORP�E�ŋ5��S�*Қ�%�!"O\M���6�=r����]��"O�L17(�G��$1'	��XM�p"O���IA�#�!��|�X��C"Od��bΎus�P3��E`�Rф"O"�y�Hw��ao�(�&p�2"O`�0��dȪd����l�Z))V"O�-i�A�����_�B#�"O� �l����;�8!w�:��A�"O\jf��D'z%qC�Hy�~�B"O0�p��HA�ތ�#�ƉL���"OdȢ�"w�����6J'4���"O��yR��}u��Y�-ΰ8<�"Oҡ20��
�4홒c� 8�B"O��f��Tw0�Y6cO�`�P��"O��a䄙+B��%1f$\�P�h�"O�5k�Π�Hz���9�z���"O�
FĿj�z����	t��ܰ�"O���D�{C0��1��	��� "O�� �@H.iWjMy�h�Bs"O�I�$/��8��Yҕ�l	xƎG��yr���	�p�P��_�Z�#�(؟�yR�!vhTz�CēQՐ\;���y�n�* p���L�R�KA��yb�.7,�b#g
@K��8���yb���	J�it+��p��'n��y2h�"#��kW�U/|l�+�솆�y�Lt:e�5�z#��;E�1�y��ɴ8�������k԰i$�"�y
����ũWK��c�%Q���y2%K&t����膶-�T)� a��y��գlq�%j� .����b;�y�
�f���p��
�����ǎ��y���h8��E�H�&.�gh#�y��p;�h#�N�$��11���y�O�#������	o�N�1Ό��yr� �߄�P��M�9�P���%ܮ�y��i��ѣ�2~�z���,��y"�9*Y��paj.�I�`���y�A**��a��ؕ��s�D��y�C�0u��;�e� #�}��Q��y#߃o�lH+$�!|�V�{t�΀�y�LL����C�J#af�bdeO4�y2j@�dbL�%��YFF`����3�y� �5*y�ӭK*TMX��qG.�yR�׷u7�ȳA��9�2]�`�M��y"hO:^�d�k�O8ľ��P
?�y��63�l9$!O74#X�YЩ�6�y�n��~�(0;�K���P!	��y�d��<�T�����#�a6�y2�	&�@�� �{.�˦�ט�y����D���J�|Q~�9'�P��y2�>a�I�Ћ�? �(�%�^#�yB��l�k�ɋҡ�G���y��֕vӾY�0��"����'$&�yR��2d a���S6; `G*���y���~e���O�X������yR)�5)sԃ��@�"��#N�4�yr$_�t�"��v��>E��t��yr̓rԼtb�h�n&�|�SO���y�m+*Bݘ�)c��u�c.J��y��{-�a+`�\��x�-��yBLO�X��Dy���b�)8����yl� tbE- q��	�����y⣆($��8w!Urmʝ�'Bʀ�y2c)T�~  ��)t���R����y��ى�@]���L5r������y"��Q��=��+�'�����K��yR���r
�T"���%PT�c��Ǌ�y�={����Bg£;`�R".]��y�O��Ri�A�V芐C �Q�T/�yB�y�P9 f� ��)SA�ζ�y
� �|��cY �& �N�:G:�I"O�]yp�E�EV�(g��[�,��"OHp��K>0�n�SEM��b�>�k�"O�U��*@���52��тc�<�S�"O
L
� H��N��l�
<?:e
A"O���a�
?W�6�R3ˌ�3�6��"O�xkؘE+��SFϑY���s�)D�@�g�    �P   �
  �  K  �!  �(  )1  l7  �=  D  GJ  �Q  ZX  �^  �d  9k  |q  �w  ~  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl���2<O�1"�'"d�p&$�#f�<b�FX �~���$P�0�ȡS5�ʸ?8V�媜.�u� G�~�dM�r�Th o,�DS�F�"`���d�%�]pv���ZFZ-���[!k��ם�y����џ��.��:e����@������h�^!I�
R�?���kư�{��-K��6mB.D4B�'e2�'��c�c��Sw
B�y�=z`/Z#,��'���c�Dx��	��*G@^�?����0҅�Y�R{�1�0�C#H�Z�Ƈ�����ן0�	ݟ�)r F����N�OX�I�?����6j䬃��-������Tu��\ϓ5��@�`F���^yɤ�Țn���'��+�$���{� ]*��?3��  ���;QfZ�� k�N����O����O����O����Oʧ�y���h1��0��V M�6d��?��i� 7���ᩪO �l�+���xش�$1��� ��!`�	��#׀�Aa��q��R�����������Q���<;�� �$�>2)�`3���Q��]��#�THb�o�-�M�e�i����O��I�J�D>H]I��'1T���������t��-��#�5p��H"V�(�(�J>�j��ɦ%��4]��V�X�~�n���fι�Qs�Ow��3�ߌG/~|XV;�MC�i��6m�?�X��D�h��at��(S��|�B����pATN65�����b@.�*�� H�6A�D�oZ�Mۅ�i5$O�'r��qբS���Am�l�h�R�#�]�p������G�(�P��!�F�m��6d�r�9�IZ+������L?@�*�/&N�y�	_��?��InѪղi����\,r�P��P���RK�#.���<����?��O{BU��)�?}ɲ�±}����y+�<e�L����a�Ti�S�'�x)Ң�)s�܂�L{�� �,���鑧ľ`�b��#���0<�ħ�ٟ`��=��Dj���ɰa�k�,��eǜ�R���'R��)q�X�0��B4��d)�1=��u�.�O=lZ�m�4x� ��Q �j�ΆO*�5�޴��$�	_�tn�ʭ��H��DB�t����²M�R�;��T�[�	 ���Xr"�'H�1Ɇ�'Y����(���	�f�B��DA�%!�0��3��j-D�K�@%Z����	ѳ�h����@�"�\)���Dx|�q���J���OX�l�5��O��?���Z�
�|un��ņ"P�S��'>R�'i�I�.||Sa��h6|��k!  ��=��` ��Oy":��`#��)n�6���▤���g�'\�e��d��Q�`�`D$�ڠ��DZ�JU� �;D�d9����!�0č;.�baA��9D�L� ��c@F�'�,QXv�3D����6j�x���	3,���R�3D�,r� G��Pr1���O5�H�4D�tPD�D�%F=��j�QJ�<���o8�S���JI���&-V&u��`U�$D�<��L�:}�4ų�J�#�8����"D��sC�\�p�f��$�|hI��>D� @�76�q$OɒP���Į;D��PL�mE$��A�Gp6`S��:<Ohrt%�Ǧa���4XR���d�ѣH�S���B�h�I2Qʊ$�ID��<�R��H�Ϧ�B��
_,#�L��\z�e��q�	�'BP��0<	VܛUl遰�]'&�rh���+�����ȏ\P��B �-)�2<��ɜ?G����O�hm����Z�Uǚ�¡��9l�|�`H�FyR�'��OQ>�F��XV�\�fϙmԱx�I>��Z}r���MsקD|l�P�n�e ��g�_�x�v�|B�θ
iӵ������P�F�up)P S�9zf��X�y"K
;yGFQӔ���]{�bS��y�,��|e��������A��˽�yr�{���xc�]�wn��J#j��y" Ώz�樃�K�9p:�Ec��U��yH^�!����j��?�Rj ̠	��V�|R�N�F�4�'��'���NH�#�d92��Q0�B�N�� (�#�&�M[4�iU�S�޷ �S9��'��p�mB�#��'�X�0m�T=i��`��@�q�h�,����O����VM?�@)��C� \����)uFPI����M��X�@�3��Ob>�d�O^�$��N�H*�bA�{^����
/¨��dYt�m���K��L�����#B���'�7����1&���?і'\lU��`�n0i�V���b��{���t�����'+R�'�B@l�A��ɟ�̧ج�uK.��� �'?����+��k�4�ѱKضQ#�x@	�B�� Pw/�&V�
��FZ��Lh��e�C��S���1q v��ϓ@��{��
�7U�̡Tc^;9Jn��Ɂßh�	՟��?	���T*?p�H���!V��lr&��~ !���,�m���S�	9�5�'&�$_��'�R6m�Ob˓ �u8��ih�S�kc��a��G�h�NI���JmQd��<Q���?���7%����$�!f� ౑`֏�y
� ����nW;2�����2w�ʴ8��'�\��	[�v�-�H2�y�䊋i�&��O�-DH����Ə�0<&iN���8�4�?Y��k��\*�;_YR�����5Tn�H��?9��?Q��䧵�'�� b�ǝT�V\�1��5�D��#j�,ȧ#n�j&+ p40�Qd®�?�.O��aGզI�I؟`�O�|��%�'W0�#�N?-DI!�T��R1�'��C^8h��p��)6&��	K��(S� *����cV,k��-��܊ �S	9f�24�����52��EW~��R�o~<�O���ɒ$P�8����a\�=���O��;��'#�7�Un�O��)��N�.��� �e��6#��	�'�2A* ��Ԭ��/�J��TЏ�D_G�OB"zs��#
�Vϕ���m�2�in��'�R�A&z��	��'"�'�"5�v��!��	W�m꣡���p��۷=ǲ���aU=zTX�771�1OX\�# ��)������	�4s�E�-w���3e�\��@���(751�1O �4+^�$ʌ�*�R�0@�л��'%��%�~��'�ў�2���s���3ǉ=U��+�^�<)�>��E�׬7$(ɰ�!�Sy�� ��|����$I&x�Ո�区
��(x�L>?2��!C]��$�OJ�$�OѬ��?����$DC7p�&qi�	�<Af8ԡEƣ�����'���H0e��z���x� �0!#}�g*�MS�8���d+��bA�'T�8�t'�~"�a�!i�<.NZ6Ĉ;�?9��'6��PG��+6fB<�P�%Xr��ߓ��'|��)�G��$�f�A !ðUo�T�K>���i��'��-!��}�N���O�ĻCiҜS��p�0Eˑ�X�	�d�O�drS��$�O��$Rg���<Y�w戍ӣ�=j�.�b"��G�y�
ÓX4��T&�C�̡{뎌�?�GkJ4=����/�*�c�m[V��YdG�Otum7��d�y1 X��#˕V)�p�LO�{ �	ޟ��G��i�1i�d��㝖RԘ��͟0�'ў�S�?)a/l�6��� 7;�X�5)�蟨�'�658��>I��?��'�Ȥ{�X��������(���3(?��{��?���.1���c�8E�<����%���ST���c�8qэ��v���c5]D�ɝ%vf}�PG�(P�B���
͒W�Eq�G��s�������?i���5Ez:)ٳ�,��"��&?Y�g�8+�4.�F�'�>a��K��{u�x:GgۺXk���q�&���O����O�˓�?�Ο��r5`�i`�S��l�Py�V�	?�M��i��' �h1qA��[C�9s�š�X�#6�h�,�D�O>�dV�$Φ�ieB�Ov���OF�d��, s�
ɨ�Zg��]肥IJ�"�Z���u2�p˕S�j̺N<9�ϐ�UC`��-�q,�9/�Q�`�I�U}�1�XS�b��08ʧ*��ԪflLҼ�»�8��$�/ }L��!�T�M+��i�2+ S���Y�$��2m%V8P&��y��J�Ψ'ȑ�Iß��'�r��>�Ǔ �
Ms�DΨO>�u2��sy¢n�@nf�	|��^���'�!�J���H�2G�ԥr���/E������ߟ��	矸�ɣ�u��'��?���Cd�̼g��x��V�y>�}�1�L�.f��$4�����fW�'���!AA��(O��۴�	�#�LA�	<�封�>ob��H �B�8���֔!NpY�eA���(OJt9�ל`�\�u��!��Ƀ�K`�X�Gz��5B�l�C.�ڝ(4	]*.B��i�-�4��ɏنXR�|�/pӰ�D�<i��^�x����\�iS=�0�[��@&*ܛs�����	�0�����|�'�؅p���s�H���X#Y��]0#��
b+��1U��h��i�
�||iE�'ʓ~+�<H��[�P�f�$3⤀$h�)}eT�dK���\�-��z�DI���8�J	�u�	��M�*�P;��!��$B���R�ۮ-��&�@��	�y�Ց��̺N�2��B������Y��8a\���!��sئ���Ol⟈ID�$§�y%�4df�qi���R-ĭ!�d5�y"ꗷּYpd��9J���0�F��y��!�H��r.��5q&��\��ȓ9r�(��$(	p�+"��wQ̤�ȓ0B��b�R�+%ȸ"���2v�l4��4F�@2Sc^1=���R$�,4�B��ɛL�"<E��灦HQX����ɬaDp:wk�}�<y�I�-�T�@��>�*<U�}�<'���M72���+�����.�n�<	��(���y��&i�&��#��<f"K"Α3b-SY�D��![|�<A�=L�\�����~�ʌ1�-DOyi�'�p>I�`Ba��%���ҌȀ���]r�<� nX��Z�#Ǻ�H���9��$A4"OڥKR%S�t4�A W�ڍe�<�q"OR4z$Iv:���ٝy��U�"O�B��݄HbXQү;T�ـE�'j�${�'�8�A1!�-R2�q �.a,8��'TX���^!lg>y!�c�.��di�'@�@a`�8(��Q�3NT1:�$A2�'�6�A�ڳpX��`F�X*:���
�'  ��k{��A֯�q�TA9
�'|
�[v���:
�!�N�;l�:� ���� =	Q?��5�V7X��`0�lظe��� `k!D����U3'�s��ќ{����P*>D����@	U�,����pl�ȃ@"D�ܙ��Z�IFT�S0�L�b3(t�"D��U%�w�4�A���Y.�# �"D�L��(�:��aId�#!RQ��L�O�mS��)�`b ����:�H���G��K}����'�*�8t�:��Ӷ��>7��h�'{���Ϗ�#�\��vC��*s�\��'�$�Y7�8v�>ђF���<k�'���� 	�,q�����(8F�@�'����/��%՘����˥?�+.Oh��A�'R V*ÙqN���"���(�
�'��=s��*R|��$��r=LE�	�'%�i�� @�ڙ���9t���	�'&u��CD(-�
hz3LU�e���	�'�0ݣ$��'xsZ�m#.��M���'8�@�'G�rr.�/���BkJ�aۖ|z�'%¡��bƛeh<0�(S�Kǜ0x�'���B��F({9h��`� wņX�'R"s�*�(�V}A�G�)9�註�'�.�`�H�#4�I"�3|T��'Lغ�b�D�����q���k��DF�lIQ?5�(�Rx��Ë�+X��c�4D����I&�zux�l�.*%r���E.D�8[fG%�, B�z���Q�,D�(Q���VT�4A�Q��mrA�8D���عt �S&)�q^�Y��2D�d
��5���"ͰI�<���O�Ă��)�'P:�a�����hV��gOS&/��@�'`���H�� H�E��'Lh��'E"<� ����x�FD���l<k�'#RX���ւ��XZ���r�^Es�'�8�4%O#En<t���f<��k�'�p�����cq�"��Ԇ	���K,Or8���'_�=+g�CJ��l{��Ȁ{�f8�'Z���S�J�1� B��r��p��'�P����3��A�&�N �ܐ
�'vY2�bN�"T�ͺ�jA}���
�'c~��a"";(t��!]��Y�"s�t�#�5�c�O�/�,@��Ш:�v��ȓji�T95��WK��p�*_�����<�u0�*Q.�����ND�-�>��ȓ`-,,B�JVU�Qx�b��K�⹄ȓxpz��7/�&.LL(��@7����2�`݂�B��v=���/��S�L�E{"hӘ������g�B3#�ꥑG�		lʀ�"O^{��W�#-:ղ�ȐF�b�Z%"O��S�,ݰ>^�ݨ��!Cx�ē�"O�$HB��d���RG�h`��"O��sV#,4����PL�z��Y6"O�q����j~��Ɇ��ifUC3�'S�\Q������)��L"0u 0�c^!`�D��ȓ#���L9f�ֈ{�"�'SH-��S�? .��.�>Ax�N/A�쪆"O�Z��ڏyH�fT?j �W"O��A��5]��X����,b��[#"O��X���=�<8����lha٧_��	O1�ON���o�.J]�����|�0��"O����#�!G��)&�F7#�B�P�"O�E�AV
A�	'�˸pF�PR"OZ�C�O9gZݭ ���A�^=�y��>%��$`�&D/�Љ@�ɞ��>q�ha?	d�s�J0!'ß~j Xs�Sb�<�1�S%?�Bi���
B4�5�e�]�<ٕ�l��DZte^7��`�"&QX�<������`�׫@�c�`�Kl�R�<�A�7YA��cD	�.V2�˵.�Q�<Y5`ƾ{�`��
9 6q6�O�'���c�����}�J���&�y��p�����!�$g�
��&#�b������3I�!���_� 	
4�V���*a�<�!��� fU^̙P�$,y�9bAU�!�HI��\�f��
[r4��u� t�!��5#-4A�-��Krb�)��!!�"�̫�O?��%]�R�X̀ǄK3L�t`�*�v�<iSi�V���F@^�
�H����]�<��NKH�)�q(�'.��q�l�c�<��ɔ4t
A��eL�Y�$��d�<��h�}��QI'�Ra`3b�\�<I*Au���:e�J�G
I�B�YyBK��p>�3�)'�F�B�r��%X7'�W�<	���T�:B�Y*d'n��1�R�<1��F����c�=��̂%n�P�<A��,(��BR�֕V�zLk���J�<�0���GށC5&ҝx���:���Ix�d�p`������C��V�TK
7 �Bŀ��5D�T��?lsbɹ�j�U$���4D�lac��D�^�c�OKЭ+T5D�� �I_�:EKv�
3����J.D�$锊Z*��脥Y�\4�9�0D�@s�cD\%��Oݰ~)>)hb�-ړI/�D�䧏�� ��!�vUl�G��y�[�3X�e��
i� ى��6�yb'I"���1�)]SX �1	���y�	�<'�8��l�m;*-Pq��y2(��a��,k��J%dy\1�-�,�y"��%�����&�1`S"��?�� a����:k�j�h�4`խ[[u���d=D��i'���8H�}�G��M��8@�<D�`����K�V�*V�siYW�=D��S0c���Ġ6���G���gc>D�٣�ͺp� �`1FQ:0�r	�A�9D�Xv�ţ�p�KkS���Љ���<92��S8����m�:��f��", bhJ�+T�l�d�4R:���B��H��U6"O����>7p���b��xy�p"OL����;(�H]Z�ؿi�C�"ON��f�/i\�`f���Tc�,� �'�P�H�'�Td��&�6#�� e�C*ɲ(`�'�䜀w����L�fE\�1by�ȓK=x%���\&Zkx�ë���݇ȓ",ZdA�f\V��be��F�ȓ<4�L^�0!D����t�ȓ�.(s�U1I~���"��E?R�F{�DY���f|�A�Rz��JN �Z�0�"O�;�J��3O�h)��օ��0"O��%b��K��9C�X8�
�ID"O� N��H��o�� �3�v��"O��	&U&z��/ˠ=͆�"7"O�}�b%�
<� �Ҡ�-Q��j��'�|U;���~��4�Dȥo�<���DLHN�ȓ�rEB�
��8H�H��2,f}�ȓ4�@͉QH��k�.| ���23��a�ȓ:��d��
�~�]X��9F]0���9S"4�`(*8��)HP��9]�
ć�-���K�_I�f�Q6�ŵdu�ٗ'���`�'�t1j��8���v��ҩ�ȓ
�pc7�� A�bi�&�M*1ZH��J�X@��ȤV����j�]��1�ȓ *j@�wlD �*���iW0OT�i��P�"�-��{��`}R�gPx���v����BցN�ՙ$"]�|a���o%D���P̗150dY H!q鮄��"D� �J�=Z���(�y�rx�.D��P��؎B����Y�z�z!:��0D�|JGI�3�� )]Z"H�H�N3D� �uȔ����˙�?]����.��e/�''�ԝ(6!��{|�ҠSw����UQ�L;D��r`���^t��ȓ�8Y�!��7�@B�
�F�N��ȓY��(��@Ah�"���Ů��'���*� ��P�P�&NT*	a����Q" <�!��2"��Y0c	C�J��=�	�gM�#<E��䇘)c�� �Q�6$x�3�`��B"Ol!�0b �{>�׀\G	�@�D"O
U����Rha���D�f�`��q"Od����5��`Cf�	1M����"O�m��(_|��!�R #d��TQWO��F싱;�r@���۝�����OF�'��	��'�r̋@)FԦ�@B��?��S�]ƴ����1{��Zc�P f�P�Ƀr#�4��ퟄ�I�u�\�Q��ʈ[;���V˒E�'(������H�L��h��G[4X���E|@��$q�/�w{(����KB`��3Z�l����-b� u�"�f�'��I����|�s!�<�r��DC�0U�pR&�hyr�'��Rĩ����z�ƺe�JTq�a剬+�dH�W�D?1�Nc�ȗQ[f� �օ�x�����Wbh�թP�e�v�׭~�<��Z��t�R˒7b�V ℊK�< ��6����Gh�m�QC&ZOrP��W(�uhY�,�v��L V� B�	M�A��K_�'�\%蒡
w��B�I�g�\1`�1j��dx��1f� ȁ��{��~"b	� E�u�ͣ@Х
P����y�A
%���+W��8�U�"ߊ�y�B**��x��J�';{�-�����y�o[�@H�@yA��J��P���y�J$0��C���,J��� s�R��y"��ce� Ӯ�k=��P���?��)�M���q�G&U�n��({x>A@@;D�y1�8p�b�W*�30��+��-D�����=yV$y��e83�DaSD�5D�C�H�b�8S�Ϳ*�>-�n5D�9�ǀE�4����<��5��.|O2�2��>AB���0u;�g0d�~D����d�<aD�8&2��5i�>b,hأ c�<	�ǓjY6p��(;D~�`����J�<�r��ih8���J71����R�SC�<)T�LiH�qڅ`˴g��D:bH@�<ɔc\&�M�$O7YȊ�#� ��'{�i���~��F�E+2��6N]�1� |i@�h�<�5AמN �0uabZD��	�d�<!���u�F0+�V�_%	�Ea�<� p9����1�0� EA�*[@��
�"O�������B'g~�	�'��}ztiĠc�4��H��o�&��ƤX�'"�>�	 �@8����=
$P�fBB�	�u��{U��[���vi��rrB�I���d� �NL�l-�$��c��C�6_��t��@�H�F-��\��C��k��q8�g�2;p	 d�)1�C�I�r?`�H��}��Dj�.�+���1k��~�ɥz	�т�g�e�� ���yB�ݠ_ֽ��j�i�f�PI�	�y�O�I�@�HP�*+�ԩ�G)�y2Q&sS��㎝%q�*� �-�yb�O��<���j�ع��c˘��O�L�֋�Φy�Iǟ��'00�JI��'��	k���4���yӐd2���O��D�OJ��B��Oxc�擫s����O=HG>��%��v.>">I�(�F�Ow6�3����,��1�'G!aЈXQ��n� �I���Ox��i�iO+-a�lp�[�RN Ly�'������5G�9����PJ���k��I7 ��oيA=�i���=EN���?�����|�����YZ@7�ǆ4��9MZdџ0p���<`����2S�2,��K�BF�Ot	��x������O7�0�4��RI�U�G�ڼO�����O��K��\�O�s�̨!d�&v/:� "�H���U��$T��'��'p޽K�\YI| f�=Y`����0 1��ab�'e���S��y���$�F�)S�ìMI�p#'H�\d�%�M�ԫI��*�F3}rD�~��-T*~�V�;���^��U���K���:}�k֗��RM��h�	i�H�dn�Rɺ ��Ox��F�>ѥ�>q��RF�DS��!Sq�V��(l����E���@�<��RQ�D�\�OJ���e�
-N��]��b��䴟D�u-}*���B�]�	,9��x1"57�XE@ࣃ;#A��C��Hy2�����'$DD��,�MM"yt��;M��zV��?�4D��p25dP��|'?�;}����I�lD��� ��iC\�c8��d����?��m�r��@ӷ.�N�X$��\�<1Aɜ
{b�X�p�݀0�<�Z�K�����Iџ�'/��'A�	f�\c����$��.9��,q�;c6���4�?�-O@��F�4�'F���$�\�Y+,�2������PQP&��ē�?q��OH�MJ�5Q�A�G_n���B���ȓ-�x<�B�W1�0�A�b
�}�(�ȓ6#���A�M��})BM>Gz���ȓ^��[!H�K��9%�V0v"�M��c�Ddq���6r���_+?3����SF D�e�K	�����H&>lpt�ȓh����B���J�VE��B-lf���X(����r�|\#�+ا-�1��L����h�n(�)ǝ�|�1�ȓ%Դ!�⎔/"��֍I�/�|Fx2"4�S���~E�4'�3rGpDp&+إ�y"�W{���d��m�����9��'�v5�2��]�)C@��]�=�7�U�'���:a�G�x�[��.o���a��&f�EŻ���/�%��!!�kȨL���4[��#���
�Z���/&<�)�@ޢ	�����o]9b��#Cќx�]z�K	<5���0A� F�`��R�'�l8�0�З2,QjشF�܌J�C�+k��}��`Hx9��hT�'_"��zmLT��E2�T>��O*8X�������xZ�\Qi��J<�v�!.�,8��	���c�Uxx�$J"� �<��i9QH]*@. ��KQ�F7X�'8`��b��ot�(��"�>�$��F�	�b�b)��{|T��IzX�����	^��;��.X��!,%OޅFy��4V�����R�!!L��|Ia��O��ą:$�Q&OZ�X	�x��#Q��G�j�0(�r��]6��(j���y��+g6.�Z��J_D��G�yB.�  ���9D$�
SV-1!惝�y�ȃ�z9�	T��:0ژk0�%�yb�D;)i��yAT�"��t0��	��y�K��>~x�(d������x�쁫�y
� �(iw��B�b���A.Gn�l`�"O�p�dS���U�U/ĵnsN�c�"O(0x��ׯc1�p"���p�Lx'"O�1Eγ!)��Q�L�.�j-��"Oz���O/ZR٤��+:��)�"O�}��EK�1�����A�W�bp�S"Or�)��1�9�/
	S��`�*O���G�	�徐��D�dnd�'1�Q!7��.W�Ь�11S�%��'��3�lŊs�J��b��(�h��'B��bdX%~� 'Ă�:�!�'`(��C�y�"튕&�8�Ł�'y��� ��l¼R����~�;
�'W��: JJ�4	���*4�tJ�'�0Tx�ڢaZ�� �dQ*�Hp��'���Q�T�{�2�3�j��'@���A�3LnX Y�뇉d����'y��Q�F:n����DL�o�B�'���ņ���-�c������'��X ao�ʵ�Á]�ft���'�$IC��ݗ[���§o�]�� 
�'cj��S�K`q2�\;(�B�'OX);R�̂U� )2���>QO���
�'�lu�}JM����S�1
�'|�yoś���q��Lk��	�'�����'��?�!cA�]�?��A�	�'\���"c[�̪І�4?v ܹ�'W��q�%N-
>�xs�5��a�'2y���:�P��h�0`ʰ��'�-*3h/;��i�s�7u�6��'�\��v/�!`���AU�5~�y�'�.0c�ĺT��rMG,�����'�&�'a���ڡ[��^�%��y�-U.o���E�)f���Ĕ�yb�Y�89��.�� I0d�ҽ�y�h�>y���ÃV^A� ү�y���n��`*BA��za�`	M�y�@T9eAjM!����x�ઋ1�yRO&"W��R��˭4PS��'�yb�߳ckа�V��,~<t��U���y���E���8� �q��ze&�!�y�mI.�ޡ{��h����I[�ye�\L�d`K����5�yrl�" ����*ՁQ�:0���V�y��B=9xd@�mE�G��-��A��yI0na2���F	*p�vB	�yB��2'M��!&�V1Q�ʩh�����y��LN����'ʙ+`ڍ�R'U9�yb�S�{�RP�3����z�ZB�M�y�B�2[��Ht�������aH��y���4O"�%��׋8��I8a��y��r*t��ǫ2�,��ԅ�y�aI�O�8H�.ɶ"��]��W!�yrF]"g��Ź�j��F�*@�آ�y�H֔s���3ɛ+1����O��y���O[��X�jI��@�qN��y���F����/�Z���H� �yr%��V�Bi1�]��lp�A��<�y¦A�^�z�pdi�/�D:����y��)Gzvʰj��[D�� �,�y����ԸAJ	[Q��������y��RPޥ��7S��L�`�L<�y뀖xܠ-��j�35�b)���\��y��`^�@���(}.婴aT��y
� ޝ �`��;������M�vES"O�!�Qƹ)�X�k���{
(P0�"O�h��hD:N���H���2gY\���"O؁���?\h|y'�)XL�%�*OJ�Z�I�q��J���i%�	�'VF�y2h� ȵCW��Y��'[�Ɉ�C#o!L1Ў-{m�8�'$�	�L�J�����vx�8�	�'�z�z D'�}u+V"͐Ĳ�'HB�EI�<q�%9Ta�,��2�'&����l��,i�`
�n��'q�eA��*�asej��T)hu��'�t$"#��6dj�B݌w����'G����54ۧ�@	{sh���'7^:�ƍ	��<	f훉L�pc�',���HJ�v��8�e�H}�̄b�'DD�Qd�(R��5c�+�,�#�'��IѰi�:|�Ɛ���3u�M��'
^t;�Z�5H��d�_;Z��{�'��̰#EĂq�Np�$D@*U�!!�'x��j��}G�3D��{��A�'	�,��E�d�`S���*E���'|X|�0Y<�+��>rƢ�i�'v�  �ljy4dU�p�b��'��xu�[2V���@�?oZ�'4d@2�c����P���'c`�
�'��1!��6�
�`�RI��Dq
�'uj-�5j� ;5��c h׵H�b h
�'�vx��m��c��|�wcO<^�Z
�'":��o��.q�u����;4��'v*��%�	I>�%���3��u��'����`ӟInj��L;W����'��p�!��t�<A��Ʈ8���'�1Q�%��T��C-e����'��ice�(^����/�7bn��	�'%� 9R"6D���@f�J� ���'P�P�3/ˬ
�2��R1>���'�8(ɤ�''��c��Y:4�����'uxX��<j�0�Aܓ2i�t*�'�J��S��2Xi��
�L�&A2ı�'��KW�Ʌ9��YF� ��i�',�}a�/+b�F�AQ��C�l̡�'�P;��E"&���AK�4+����'� �B���DE�1aa�H21Ne8�'���)b��' ��݋0���' N)��'68����"�B��
�%SĹ �'���OĴ~|��A�'L�:�'���w(P�t���j��G'(�z�'ԨKD$�֤1b ��0t��'AP�aң�=fX��W�7	�����'	�u�p�
�Hj�� ?$� �'��ҫ�kj�9�K>s�D�@
�'�x%Kq�15�� ��eZl2
�'����ea=�l���
�'݊�S��V!dPv�B�ִ}>u��+^�9��*�g��\�2�ѻ]�L��ȓ6�vP"'%ڙPs�Hю;D-��'yʽ('
 S�<pc4U}���ȓx|(h�5] ��wl2I<��ȓ  �c��v����O�B�2l�ȓE��,m�$@B�ª	JBm��8D�0B��Ӈ,�P�1�,�f�)v()D��"ǫA�!t�٨�MżKW���%D�@���)����+d���RJ#D�� �ؙ��E����塆&l��P�u"O�������$(�!��[n !�a"ODE�+2kf�� �V�m~�I�0"O ��n�T;�u��¾Co��s"OT�k�F y��� �F�J[J��"O�+P��
������i.h@�q"O��ac�:~JtP#�Is'2��"O��0jD�H�8�@�o�� #F9��"OH`�"�:"50s��.D(\�"O�)[b�:160k��U�-�� E"O�a��D��Yӕ(
����D"O����Ӥ�Ј���R�~T�5"O����$o��m�Q/ћl�&�jc"Ol9�î��H��C�#G��82�"O"h)�����*oU�O5(�T"O��E��4(B��@��C%֕��"O>8{���<tXP��Q-�`"O,MZ��1�lMB�L�T&��o�<��$S�
fr��W��y���8m�<I���/����#	,#������R�<ID���*�8���"̪2�>9��De�<�գH*L��i��w��m 0�x�<i�N�^�sk_4�`h0R��^�<�aA�� _�QQ�ɧT�<틡ǉu�<y�͚�l�DI�צ<5�}��_p�<��V��XZ$�g�~��F�LC�<a�)K�d+��_�9N���@!�e�<I6�8S�2Т�	T�S�6)p��Y�<iMN�&>j����,�@��fF�a�<��B�a^�EsP+H3tA��;,Qe�<���;Y���k �m��TC��[�<A��.��dHB(8{Ȅ��I�o�<A���WH�h�ɢ_�xi!���m�<q��
vTe��N~R�T��j�<��C�e�A7e��^F�@%�M�<�qn�V�zP�7�
�;�*s�B�I�<��@U���- c��``i��_�<�&�/͖m�FJ�ɺ�6]�<)��ݩmݮ��$�61D�\Y1ZV�<Q��S)f�X%&#۴7�F<��fDj�<��h��h����b��G�b49v�i�<a�U�:�(�ɅAW/`��ŉ�a�<�&I���d;�Q �0�"LI�<�ĕ9v�\P:�B�f�<�G�F�<q��Q!�Z ����j�0�q!NB�<�&Ct�����eO���	�|�<�ᕤWňq�X?�R�E�^y�<wm����sH˷%V5�vf�I�<a��Ps� ]���IK��w�
M�<a0c�C�P%����V9脀 J�<I���l�N�ao� Zs 5��N�<���R`=�1�t�_�f����r�M�<��	C�n�VE�.��7l���_B�<��kO&I���c  K[��S�d�<	��ڣЬ��2@R��,��V �^�<���@#�f� ��+���:�[�<!���'H���A���|�D("&#�T�<!��]�0R$0	����;"�Uz��Q�<鳧կN�>� ���:���&d�I�<9�H��L�������f�`D��'D�<��=K+ ���[��y�;T���ӤU(Wk�P����]S��?D��@�����k �`��Ah	d�x,�h���	���nx�|Z@�32|�Y�.V�VR4j֩5D�� � �AO��DT�SoF7łS"O~@�w
���	��W�p�Y�T"O�,�𯆛]F�}�f �^gX�Y"Ov�Su��dhց�-͵Z��R%"O�]*�A$��L�LQ(>�ΐ9 "O8\�4�-���hӂ��d&�rD"O>�s�)04�sA��4j�D"OF�iF��Nh20�E��#Iz%ʤ"O���!��4�|	ZC �˒�B�"OH��'�^dJ("�կU8Vr�"O�LI�� alF=�g�-;�p��"OH�A�c&-(ue�f����"O�в"^��p$��U!�"O����ˌ�E��e�T�?��Y%"O����قPD�0G�I6{��]��"O� bC��	CDH�+���p���"Ozi	�:8j�aq��0?4�c#"O���6�V�
ܢԤ+M*l��"O��0�˞. �����x�X��c"O��1da�&�f�sS`�� V�*�"Ol��5B�d�"Y��G#q
���"O�x�T'=`� �{�Q�
O�`hP"O� bF-rH�$Hٴ|K�=��"O�y��
��B �X�&���R"O�`�S������ؔ��	? �e�E"ONǇ͎pa�j��(o_|��"OR[�D�(�>�"�A�UD�X@"O��*'j\;]��E�<����"O�}�W�SXn2�+��J�~�t��"O�4�n�F�]2�+��(t\�"Odi�
 E���"�!Z��b�"O���P�_���B�ML(F$�:A"OX8���hԮ([F.T�^`&�RT"O|`�'�2R��BCֺNX���"O��D�ںX R}ӷC�yW�Y�c"O�Ⴐb�[3�q��/J��k"Op�7�*��XIb+֠�>�R"Oځ0��u�����k��%/�d� "O~�(��
l�1T�@�Ay���"O0a��Z'u:�	a�>Kw|�I6"Oz��BáwΝ��]�R4l�"O(��gڃ?!���7�< �P�Q$"O ���!u(PD��)�b"1"O���׈6�,a�H��J*	��"O�	�F6�Qɧo��\�H"Ot	"`��#����n̈́�`�3"O��rM�y�y��j���9F"OZ`��J6^H�#I�͈M��"Oh05��L�E��-޴?[@\z�"OzM�K,E�& �0o��k�6p�C"O�A�Qj��%��!Ju��=q��0YR"Oj%b��Q	� ��e�!O���"O�`-W���lR�|�f��C!��Y�	���#�OՓ���'�[ +u!��I.5[f|�`�S�������"bl!��My-��O��Z��QQ*C�>l!�N,
��a[���'l-;�]F8!�DCl��Y&(W�ʉ#��#Nd&��ȓb����&,]�)8dI����(\��1�$@�f	U��bӣ��>��Ѕ�4�� 	�c�M*���&42���S���y�L�b�j��N[,�lх�#A�5:��*��鈷�!*F4�ȓhRtM�5錫4屮����@_���S�? ��;��Y��}B#Ҥ"�ui5"O@R��J�s��D��I�/�b"O����`Y��  I.A v���"O�:�����Pb�'̳t���d"O�`E�/�� !G	`|���a"O*��P�F9�v�""F�-=c�P�%"O��Z��5!d�����~��"O��`��%��#1
�<t`��"O �۵�����G�� (0"O �B"�ٶ>߶Q��\�Vޘ��"O(�����*a!�J[{�m �"Oj��&&K r'Լ�s#Ǟ>	�W�f�<a�*~���p����¡�dO{�<)B���8��}ʘ�tB��0[B�<ɳ��Quh�qW$ل]p��Gn
[�<)�)�%${T�u'�:Y$Ѓ��T�<��(��FtA��L0{$V��$�HV�<)dD�*W0�����t�����(�T�<�0��L��:��2I~�]�W�	R�<cJ�pQ�b�GT�x�ʀom�<	�ٟ
��-(F��w��6��R�<q�K��,6��IF�hj�J�P�<��BQ�4� $Y����W�R��ōj�<��.B� �!8%@Z�R:�m���De�<Y1	ȧ*�h��
z�4��<I�! ";�(��e���p�`�x�<Y���N\��K�蘋nSݑS�C@�<�����1��$�A�W�/����$�F^�<�u�M4.�li��ǰ0�k�W�<�)v��f^�/�.y��_~��(��{�u�E��lT�{� L�v]��M0������=�8�r���E����f�<):2@���l-2��K;T�v�����M؋,�����
��=��"O�͂%X\�p��@�4$���"O�q��� ����'���`��"Od!��F�+B^�`%M�L
ٰ�'���@	M�9s��k6H)�8�p�șD��B�YZ͐���c �����0��">�%cR�Yr��a����k �=�W�(�4�;�.��yRb���؆b(l�d�%I:6�U�2�ȦZ�(m�\�"~n�-X:�I8V�M:Nu��h��� CtRC�Ɂ���M��]�Tz֢
P�B�(��V=P��	Ǔi.V��G�/Ll�1f���j��	�qd}2S��W�R<CC`˵'`�4#�-z'
t�bm�t��]���(�dOФGt^��s��	=<v"<9��׮m�2)0����	��I~��.��\��A�(J�N���NL�<I5$E�i�4lC�BI�6b���(���R��R@�$���8d+֘+�	G��'�r h�n�-~Ɉ���F��z\�	�'�r|�Pk�s:���fFWv�ѥ!׷I5��2�+ڪ(��cpm�:�F}�!�9+�]HtnL=Sb&8£��=��=�cB�$�4��#+S�3ִ�c#د��J��[AD(�G[�|������F=X�	�.��e�A,
��Y�>q�8�r�hd r�0*����6+�mq�a<��E�ҏ`"xC�^Ƹ����]� jj�s+P�	4>�a�:Z��d��F�y7�D�3�'�~RiX$gMVzv�	�D<�q/��y�HO/[�M���>-@)d��5	�U�ɴ+^.��
԰�(Y�]w�Q�Y�a��8@Rm� ��DcH�b#4lO����`	#�l���Ӫa㖏�	^��Tj�'�-[%��مh .yx��$..�&���N�(3�	8 �Y�}�Oi�cO�T8�A� ��Y#�� �0��K$_#@ۀ�_�"�1��A.�y(�����rQmɱ
�H��}Ҩd �WU�����d:`Ћ��O�d�Þ���p�E�L#b�$��Q"O���˂o)�}��d�5g����Y�> ���5e�8�L�F}
� �$pG �?.�a+���qo6�Q!�'�DK��D�����H����O�d� �#�DDI���Qj�6c:�|��"܇^�m�/�Y%�l1��
��|&?��$`��k9X�L� ���)D��0���G}�! �hS�UR�ṟ<��)@�@E�N<E�Su$�Z�p_�y���x�<)�R,-�R8� &ʔxq��A��X�D\�iq�Y��o8�pyԋЉd4+��ҍ��-�.�O�t��ۃ���_#/$9WɌ�M�b�� 4�$���'oF�՛ՋK(r>��r�9�8x1��	��d�v�ZN��!
َW-!��;���"��ҧS2�!sȈ�K�!�W���Ii��O�S{2d�g(I>%!�Ğ(��u��G�.urqc�܍m�!򤗹d����ھcj\iRa읚Q�!�ʓiu(D�7nU7~i�4:����!�$A$.#\��ǝ>[����^�!�D	�<�D�{��.@"�u(́h[!��(I����`�d��5Iկ�3!�DF�b�=���m�\��� �D!�$����<�b`�n���p
�9!�Ċi�*��JK	�ycqM�R�!�	�!�Tq���+�*��d��,!�ϟ�mDZC��~�:�����t�!���&ˆ!UA��Xl#t�	��!���������s���,	.!��K��╅�5OfB��a�F[!�$G!L�x�1U�Q{Sĝ0cɁ=�!�d��_A���V/�
��MB��88~!��8�x]������ �T�+{!�$
&<]T��>Mb��2�*ߋCb!�BFc`��^�aCz츐꛰}c!�D��4��q��EK�+�����*\)w�!��	�4�:Wm��T�"��6@�(�!�dע�t���M�_x�x���j�!�$E�n��,0�KYm�6	�ȑX�!�dm�ޭ��nU�l�t���+J�!� }�`ݨ��ߺ,3��@'��2u�!�D֎>@DX�hֳ3%^��,>m�!�]�&���Y��� ���,Ǔ{�!��=��@]4h�$8p�F)5�!��|n ��cE�����a�^��P�ȓ(�ΩPw�H�7�V��5��&#A���ȓC�(%BP���" "|T��J�-���V�s��+wgޗ:|�=��f<�#挎(GVI���K�\�q��2��X��8K��AD�&4g�Ȅ�:)\�Rs��fo|p����%/T�ȓx�@����84�p	$�/����l!p����Y�p�"�N�\����ȓ}�Jq��eN�YX�-�wI�4uC  �ȓQ�&!�u�Zx��UΔ�
KT5��K&�Qt.F/eS��B�M�9I�I��^mn�xw��<=4&A��4q�e�ȓW�X�B�;6)~��AH�2��0�ȓ\m�Uc���9�pr�̇p��i�ȓe?���T�Ҋy�6<�#��2C��Մ�r��H�\�)oXLR�U�LG������u����I�]��M��!/��ȓb�����Hs쒔"E�@�%D�dZ���0j�x����	`N���/$D� �mD�x�`����P�-�`���D D�B�'̽�����D$��if�!D���ݓ]�i�����g.<��.D�� ^E��"-"�j��$� �"O
p*�)>w��r��rP-�"O��Pc���:#�T+��%٦�F��٩1&@��pAX�i"<O.,��/��d�e��+ �氱�"O):���8\��q
��=D��53"O��z�+��D�	��,B�"O>�[N�����(ǒ����"OX�SfB;X���uE-mGL� E"O���"MK�L?r)00n:G�0�"O��p�ڃZLh�凙�ez���"OB\	C(I:b�X8�f�'bx�9@�"O�-Jv��2���뒃ؼV��1��"O���ŵ`�F(�bмhh] 4"O��k�h͘�؂�S xO�l��"OV����%^�(�Pm�M����"OX�"(Ԗ>���C��2$մ�	a*OX|
�AD%Y
S��Q�f&V��'�V���H�6��@���X��I�'$�����(M5�tR�G��$M4!h�'��Y�jɌa(i���?
�V��'�dXLB/��`� �ؽ���;�'&���@U9x����^M80k�'9���樔a	
vJ��x�n5�
�'�耢�&�;����UNZc$X�	�'{�D2�zyYO��+�`�	�'��l�h�!�D@(7ɲ� ���'�4Q��O�6�.�!N�˲ 8�',�ܣr�����3��J6A��R�'��DO��rIH��Mu��E��'�й��4�x�{Q�X#����'�|����_/z��ɲ��	�P��'z���b]<��i�ӒH�(��'3j�Z'��T��d��KR;#~QQ�'�TY���Q ��efM
/.����'V2D8�K��<��(�d/ݗ!�~L3�'�aC�)m��{�늀q�`���'ޤ`1�K�4���V�׸_t0�H�'�$�I�K	)Bb��V[�"1��c�' &Ya4WkuP����<��
�'nT��щ�YF2�q�H�9�p��
�'�]�uʛ+c����Γ��D\�
�'�&�23	��w[
a�@B�f�P��
�'����m���Q�+W�dȉ	�'lVe��F�80H�ɧM�x�")K
�'Ў���C�7�.!F�ЉB�J�S
�'��D��ߦ�Z��Y*4���
�'�B���D;�%p5��4����	�'�Q9��M�:e�5"%�]�`��x
�'¢	�c*�0Ox��c�i�p�X	�'-�����e�'M��	w<��'�H��"bܼpÚ�R� R�	����'���D��2s8Y��j�}F�80�'�b��)bબa�݂^���
�'w%�ph9*�T��K�XÀ}Y�'O��ET2)e�)�+@8&����'/j@��	HT�� �㋘t�����'�p�T�Ϸ3H���`�\7vdA	�'�\��ᜆmB���P�u|4$
�'���&N�>��!���U�ql�y��'�d����@�Q�	�d���'��P���=�>�״�3a���y���n�z��!b��j�T�����y�*�J�\�3CI^�s� HAՉ���y��V�q�|h�ƀ�q��H��hM��y
� �P#�f۩Yqֱ10�؄�d)�"OHL3p��K�Hk���zz�,�"O�ɓ��Kj�r}�v/�,n�<�D"O8����+o���W.D�MVT�`"OjE���R'j��:nM�
dD� c"OTҤ)�	�̅B�&�5cڥY"O`��&���:��rfМXj �H$"OH�pD�$Kv�gK'[ 8aF"OT8���DS9���_uE��q "Oh0�� �b��WDT�N%B�("Ot�蟛+/ܨBƃ��a��"O��B�l޴��D�w��1K��0�w"O�hG��M�pCg���1"O��;���To����I��Phv"OZdH�,^���Q��ɰ�Q"Oba�vF�Nz>,HG@�3�.�y�"OF5���Y�?��q!ϋS*�A"O~9��+�V\E�>#n��0"O.e���4�����e�+��س�"Ǫ�we;�NA1���.��(d"O��HCDTW���Ԏ	*��Q�"O��*fDǐI����҉D�MjA"Oh���i	�n�sQ����J"O�`$��<-:�hx�,�����V"O�!b�\/�,,Ac̍ ���"O6P�A�/4����$_R]�2"O6dr���x�`8�7�ĝn�:I�6"Oĉ#�ł)�1���F
aں�@�"O�)���H�L)QC���F8�"O<����4s�< �q�Ť���"O�$�G�.�Z(�ȋ/7x��"O�����B� Qp�j�0'�,�"OPU{��Ӷt@$��H�%\{�"O*e��ʯS��=l�9B�"OT��Q&�5>�	���E�om����"O��F�ڻh���@�ܨ	[V�#�"O�:�'�		����uG�q/N�a"O�(җ�Sl���� ;�M"ON�R�k��0�~�8����h��"O��S�J)�l�JWC'a�\�8"O��o�.>���*��H�%��xI�"OR墦�)7׆�0� ѥ3�$t�"O����´5�PQcuA�K�i�"O�ѕh[Qkb�ץv����"OJ�酦��Op5K$��.:h�bt"OJ�@�/�?p����6ʘ6$��[�"O�IX?L��<IDo�Y��{dO�Z�<�tC���B�͉j%�f)Z�<�Ư�@���+֕X�~E���GU�<��.q(�)'CG`�,I��U�<�����/7�Hv�(N��=�'��R�<a����P���ص���bPW��v�<��/Z9�*,�v�������1��x�<���>���PEy�F�y�<�f�Syd���9�z�y��t�<�㊜�}��ġ���ze��Q�m�<Q���\s��J0�B�H{�p1!JYl�<�E-ʞT�b�S�V/�& �	H}�<���#"�0�Bb흊�T��@d�<�lB�c�vH �A�(��X��'f�<@�V�#I����Ѕn�ZT���a���=iv�ë0��8�M��pI	�j�Z�<�"�	Q�j�ѥB�-B۰q8�	OS�<ف�͗B�ҡ���Ѩd�e��\I�<� ��򮜊��1�0����"Ov]q%C���`��ʉ|��� �"O~�$$�h����p`F����""O.���晳�l�����tQg"O�dڕ�A�+��̫�C��:�CA"O��I1/��G� �z�)�"x�6(��"OJl�r�E	On��$腃 ����5"O ��k8;�ub%GW08�F�:5"O^1�����Ўt���$颬�"O ��1�� g�R��eD�65��ɖ"O�)a�R����³dP� ���t"O���E,�Nl#�Z1 "O0�g���t��_i��9��p�<1����h|a��Y0�����n�<���F`�恙���;	��us���B�<yah� 	s�J#�/6��]�f�CE�<��&�{I�Q�U�K��Mk�"�V�<��T�r�Ԩe\A�����KP�<�c��k�nJ�`�ڌ �N�<�p�B�"�dt"քǝ`zeX5�SH�<i�vj�چ�CB�(�A���i�<a�A��*|�}(�
%�h�C��f�<Yw�֧0�r5"�,G~ �B�~�<ن��3����"�r�3m�y�<b�J��a�Qb]�KRh��.l�<����+M�"HR ޯ�,���	c�<�e��0���S���PD`�2ծ�\�<!�@ԍ�RlS���tX�Q�+n�<��C��bդ�
��������m�<�R?uX<A�Po��4�I����k�<ن/��]L�H�`�.\k�%��V_�<ɇd����� ,[�"��$�Z�<A���1\��B'.��t����A�n�<1�Kيo���0�cAY�B��Og�<��dN�kh�;jP�R���&.�{�<�Sg�zZr����B���w�Fv�<���4i�3�K��'�e���Q\�<q�J��y���hA��(�XR��[�<�0Ď9Gd�;�C]����S��|�<q��2"�`��i�Q j��ԩPO�<�E�G9 ��@c�Gi���¥�O�<����30ZD�GX���@b��OR�<�5��^���1'�P��F�Q�"��ȓz*��¨�&]b� bn_�{|�a�ȓG�Լ���8��� ����)���I�y��ۼN���)����x��u��29����m�+�2TYWk�)K$�ȓu��u�
Y�8T04m�06�ȓw�y�c_��i�¡��.X�!��tQB0�7��w�>x�	+l6�!��B����d+"�B)�@O%4�����L�ۖ��;t6�
U�ȓD����w�ы7�z`�%��4b�`�ȓXJ�r%*EW%�-���*�]��H+�L� ��&-CBY ��W(#ц��LăG�Oo���1ЇZ"Vu��ȓR��������4G�S���\��ȓ0'N�r��� �(ٔ' �H���.P��`1�N�n6�=#� M*J�n����q Bk�	�
��ЀR�l�L�ȓ4�݋�_"5q�T�B�H�FL�� ����C�n��90D�]��ȓS�N� ÿ�r-���"a�M{�"O�s%`Q/hLӐխY���"O� ��BS&�Q����#?@Q�5"Ob ���?b��G�@5[����"O�Ӥ(�S����O Q���&"O��u�@�rW�@��Dܷ~%@���"O�5�\�,�T�����1�]�F"O��jWc��$DH6C�*u��"OR��!Q�	&�	�N�"a+A"O��@��Z�C��!��N&N�9�"O�*��P�N� f�؜K~NAKP"O �D��\���PՕwl�]+E"O��K��	R.��`oR^&)��"O���!.R�O�E�Հ{�����"Od�A�h� E�`
!n�	4$���"Oʠ������"S��*a�`V"OvE���@�{;J9vV�"��X�"O�)H�H���X�K��H���;�"O8�q�E�Ur<��I�,d��k�"O^�@۶y�.A��o�3|�> �"O�YT��.2������9�����"O�e����X��(�à�S�D�C�"Ovpr���)�*
oP3�LE��"Oj��r�[Z���T.�G�j��s"O<E��^F���
G�M+gnV-��"Od�)�HWr� +�OI4f��j3"O�c.�q�4ib0��[��7�1D���c/��[(�Xi�Ι�CVB�c1D��z&I
�5���2�*Iu�UB�K-D�4�fz)A���
b ��M�5�!�DV�b�n�"�(?@�Ѕ��,�J�!��Z w��a�@��&��ezqJ'6!�Q����7 �p嘕ʑ�a�!�DV�S\9j݁n�\���If�!�$R�^S�TS�E�%htmY��ܽI)!�dǂ��@A���Q�B�:�F�+6�!��=ӰK�@� l�6%ɺ6�!�d�*�|(Q�$�����WY��!��ٙ@��p'(�9���P�匕n!��V!�]��ْ(�4	jd-V�!����!�*шx�E#$E<�!�dM�d�
�b3��rP��JҤq�!�	x��۰j*<E����Ȍ;p�!��4 �N�;�l׮e��q��� x�!��ٓ�T�(&㛆(*���	>!�A�aS��U����)�G^^Q!��h�D����JB��
5���^b!�d��#�R��$�H�7aP-	�R!A$!��^�n���4�Jf�1:���<'�!�$�=�v�Ic�'Vlt�*��~!��2+F�=���k�-�4��Wu!�$��)�=3rJ]t?d��L�-�!��4c��`B��q@*h��S5vX!��6_Y�������1��/uA!�Rhv%(�oC:o R��u!���f�&3�͓�s⚙8E$�x�!��ȃs��X;@�Y�/͘���_�	�!�䗏1ڌ	d/L
O���8�f��G�!�$I ښ5K�H��Z,��'L��!�ą �$��d�
~d�m�����!�$_%X�)C�B-Ny��ϔ�{�!�d��U�p�ݡL^�5�VNCl�!��A�&�,�dAJ	M1XYZW&X0�!�ВOXp�zEc�M L�IucM<Qb!�DB=c.�T��H Xn�Q񦡟;0e!�D>l��H d�>9b��4�E�1I!�� ̔۠�E+@^��@1i�R��Ht"O�%a�b�%[}�W��wv) "O q ��թ`�� �U�'T^d�h�"O�]if�W�N��4b�8vz��v"O�hH�� 
���'�K�m_�=Y�"O��vnӝgZO
y�5f��,!�䚀g>͓V�]�#=�y׎F�Z !�$1g��i�66x��h��!�$��s'�}	!�R�D� %"�9<!�D�<Q�\Y��M��^��c�D�i�!�$�9��8�2fƀgQ���`��!�9	`~ՉE�ҌmI��%�ǯx�!�D<x�$-����j-YP�ڂ�!�DƟ}wԉ�ƥ�� ��uJ��-�!�DPcGrq���R%#���W�O�!�䘃b)bĨr@�{�fH�$M;M�!�F5�Lآ��"C�F�qv��jL!��^1Db<�[0�ĺ@u��Q��HI!�d&M-��`A׳$�t���H�%�!�5 ;���̚��:�6'�K�!�Dڧ~���1��l)�֌��Is!��]�����M�p��f+�	 X!�D��0�R7�[�d��!�sD�7|;!�D��7��xC�m~6���� <�!�Ę�|S~	���y`ɩ�ʇ�!���Bąp�e��p�&J%�!�D�b� u #צua<�����+l!�� M���E�L�W��-�S� z
�'<�t��`Q/\������ E�HB�'�F�#��P�!��]��옰D��P�
�'7���V�G*V�)�䗱HP���'�� ��VbƍA7랏��	�	�'����ϛ�4�ъޣU]���'��˓`��B��"���E�^3�yR�K>2��*F[E���d��
�y�d��M2��C�%:�5q���y��|�*�3����ʙ�����y���:��E ��<Vt��H��y2�Uk�i7�D�ȬXFަ�y¨����F.��}x��w`ō�y��W�9�Uz�%2oˬDpVѮ�yB�5u�Y�ʘ�c-i���y�ֻK��t�fA�C1���d�R��y���$b��"9^��X4W��y�nB�G`��E,h����y"�5���F�ܝ$Ց�D��yBo �1ըܹ�)��+ !�5��O�"~Z0�E�!�4���mMH��1:D�E[�<	rH$T��0�sPfb��SET�<�F�>S#��P��j�֝�"*�S�<��(\�h3�]����=�̭`��Q�<icK�>̠�p����)�Rh(DJ�b�<�@D�3�@\�g?=bB��t�<�C޿r���E bx�ЫdQY�<�VF�� em�Qc��pf9���S�<���\0/�j���8C��xy��JN�<��I7�؉	���6:x�Q1�B�<�q-O�M�`A� &Wq��l!� i�<Y���.���BȄN��99�)b�<I/I  �Fm꓂·?���#QaQB�<1���Kg�a{2c�v.����@�<��.��4����Ĥp���%O�~�<13-^cjD��8O��lFS�<!C��&��8p�*��;7��I�<� p�¦	'O0��iBh1(J�C�"O�""üi ��`���`͘�RA"O� D��N����@�ŴX]����"O�q��<5�Q�&Ÿ'B��sB"O�=��Ț=e���I	 TL�{�"OE��Ϡ;���8d@A�qM0��"Ov��H6�`�Do\�I�6Չ`"O����L"S�z����Y�I��(� "O��J�i�'��d.B�6�nt�5"O���&���&��� �#�J��$3D�`0c���T�	�M˶2^n��� /D�a�*�E�M� ʰ8�&��
,D���F5+:���C���a<i��&D��pB^1J�x�q��/P��=���(D�$P�)S#��P�1N�:/��˰�#D����N�|��h�  	wE���E"D�{���-V|@/�Mx(���?D��adDҴ
�^c��S���T`=D�����	)I����]�j4�M�j-D�Ա���7bt���F��[�xcċ)D��b�,��0���UJ.@vԊ'3D��	!A��W��p��n̨F� �rfa0D��x@��x�ܴ�� &�����e)D��@Eȕ�9n^����ï� �p�<D��:%�6Q���7���lO���`?D�h�T��.>#�� L��*	�����)D��V*�	�2�۴S�"��0lZP�<�&�u��(������a& g
!�$U�N�`��k�6E���`��t�!���s����M�i���dԢ�!��X߾}��N+��8�ƅ�v�!�6c�l���D�%�v=i�eZ�S�!�DΊSU2��A�>pۚMk�EP��!��h<��X��q�V$��^&t!��'�ZP�X/'OB!E�];Ig!��
}p^�*Ɨ#	gx���ر?X!��[�F��0�A�^�EV��P��W0!�Ǵh���q��P�HQE^�yE!�	�4�Hr��eSP�qw� E@!�D�����c�Q%H9��Ή�H>!�D�#����j�9h�	�6	!��Ŗ+�@!��N�";U*8��iN!�dǹD�H0����:L*�K���!��Vt]ɴg��*P�5a��!�$��&��Q�nX� �L�ʂ�ѝf�!�D�Pv0��� V�R�.������w�!��G,���Y0JV�S`�x�T.�,Fk!�D-mHL<:�C��u<0�ڗOÞ8!�$K�t��-�� 	@*:�a��N"�!���8w@>�������y0�ԛ^K!�^��}���ܓbx���C�a�!�FY��ɘ���*)`�pGW�b!�D�0p��ʴWE�%�t�^�YO!�������Ǒ$D8� i$�E=IH!�$CW� �po�8ҝ���	*]\!��i1������HhŲ�pt"O���nO'#���`��B�F�c"O�l2$DP��/̥W�0	30"O�EYr�ҏ~mR�1r+��Mu�`��"O�*�M,p������-a����"O��;�(׎2�C��I�?����"O�(:��:R��i@�U�0����@"OPu�b,̬��@��*{.1��"O\�� �s*�S��
�8	"O� 4�!��ފ^�D(�%̜��h%h�"OJ��$���q��,�Մ� �B$r%"O$�j�)T#m�t�8'M�f�@Q"O���v��3=��9A�Z�x�D�"O]	�c��	�����o�*�Z�"ON� g�
�8 +�$�q��Q
"OViRAI@^,�p�4-�ya�"ONt ���> �|�V�[�)8�"O�]��@�"LP*0�aCW�I���Q�"O$A�����d��A�)�t�["O����a�_��}��+m�T�ᑆ�O��e�\��Mc�O?��<F��	"�1A��)�P�j���k���FL2�h�U)݋��¡r���>Q���@�(p�8���͖y~D�`�iM���e��l����$��H8�ʋPvpH8��R~�s��(���9\����L�%[ՒI�wӒ�;��'�"jz�V��-�禵r�.}!��z�"D,7��$��ȶ����͟d��	�9�ȥ�Ô�q��S�.µ05�<��iU�7M?��ܺc�K���W,[-���w��)v�', �ˡ��?	b�'���'���]���l�	1h��%E�c��(C���d.��[czz��v���J��%D�����a�Q�`�'�샖�M�"�=��9&�!1v�#h�t��,[�h���`"�JV�U�X\	�#�)�Z�+�'�9c2̒
gY�(P��/I���H$��O<�x���O~qn>���<��'���D�
5�mz� �	#l�j���!��Ģx�lu�A��@� ���8SmL�1޴(!�v�|��O�t^������|�^<S�Շr^�1��b٫Rw@4z��Esx�4��+r�4��H�Gv�;�n�!X�����$�b
	�.#h�ڍ����$x%��$� N3DY��J4�_�=�}(��!���H���B��=�ڴ���
C�$�HEy�n�'��%�H�	�WP��B�
 ������� U��=�񌁱�M{�����Ŧ��?ydџD@��/Ŕ�5 C�-/@�ٙv"O�a�bv6�ӧ��/M&~0)��O��oګ�M.O��aºޛ��'�BW?iP-A"*�x�r�F}A:���-���%���?��u�����hS�<��1�� �] �L"Ժ��D�K�L����ᮞ�|>�I9�.��Q�d)sHƀ\�n,��FMT�H�)]�3�vDѧ�դ,���{��A� 52P�T�-��kqnԧ`�
D��O�dAg�':7������1	у�9k�����(�5<��ـ���?a����'�(9j���t��-�T
څo�k
�4�v�'����|4�@�*^E'$�)f#� �~��΍`��6�O<��|�0`Ή�?9��Mkq��O 83�����g�6p���th��"l�1`,|h��B�Ó'����'��Yc�}
���"�^�Xp��-5��̐ߴg�P8ǣ�*+P-�����*�n�c'/	wo���RF����Ba����-i�"|���UY#׽iR:8���:m���M����~�s�<]b���xـ@���H�v9I�OH��"���'����ŗ!G�@ݐ���\Iv�K��$V���4�?��i�"��^I���Mqd%Pj�͠�)Կa^��I���d�aiB�������	˟��_w�r�i (�#"D�%܌u�o�9IBf���d_""6��2k4߶���Jo *�i���N��|�˄/������"=bqP�GA$Ap6m�):f�C��" ���A�p�ăʌH�nt�G�Q7���Q�~����a�1S\1�(�e��.0���		�MC� �~�'�[��[���/A޼����u_\a2Dc���x��#�Uң����<"�.G�M�4-���|�^>Y�>�i7 >  ��PDxªM�c�= �%G'($
U8�C�0>!U�ҹ,ײY!Ӫ@<p+���a�3;�MR�gT�U�Ќ�T��QN�y0�'x���	Π
�b0���7B�h���-�s�
�%�:�#�A�k��re	�GP�\ҥc4J���y"/XW�V�i�"O a��7���U�b���;� J�P��d �4���i�g��W�A�`�5	�1���>J|g��{0 �7�
|�!��V�@��9+�-GtE�fg�(z��HD�����tHN4�V��;��8)�	-I�1OT `�k�fg�@0��݉1�A�&�'nN�z3�M���A�:[� B�� ��!A�.��`6�
 P8�A� �0=�S�Ј|��I`る�>80��C{�'FZxj��Ƒq9��:���5w��]0ଔ�rr�=Z��ۻc X`��kّ���IcL���y��¹N��!�?���{sM�]h,��B%��{º��e��WtИ�ûJ�(����w~�K7★(���ŋɰ22�A�'�4Q��J�A#"�i�_�M�t�E�]$T�Y�.[�Rp��2@����B�㢥j�y2�&*�l� bT���3rA�0>��叱k��a�fO�aƎB�Z!<�CEb׉אi����8���B?P,f���ɏ>�tKS��:2����@"#<I���_�4�3����*N~�a�N��$�^�_0��#b%Iu̓[8��c���)_�=��vI�<H�`�ߏk��D�'��Wd���L<&1���s����O�5Qv�c���'t���Ƭ����'��+���2c��S$Q
TBۋy�����lWߟ|2�I� ������-/��F���,�8��J�:&����Oם:����!�*,OLQyae��{�d�ѣ>ti1 �3^Q�6M!eU���k1��<�he9��x��	~���l�̌� K��Oda+5�c���W�9YX`���@BEH^!����6���������>�|��ʑq��!����=�=�UkVA��� 	��n��/O?�I��!Cp)ɒp0���U�zGJ�k�}�ߓ���I�P�0DP��L�~�*�� ^S�I$:ʅ��?�
���!���N�e$(8K�㙒X~��Q���.��<q���e1�5{�OV���q$A�*x��oX >��� 4ثO<� t�:㌒+Lj����>s5�!1!�	2S�t�8焂K�O�8p��"��Ds������y򠑭��b�b>�Dˁ�,��G
�_;N����'D���'�Н]ͶPr��\�d<���-��'G��1�𙟸�������rE��6+N`j�4D��KE��`in�P�� �8'.P8�钽P\X<A���XW�Ҟf��t:�B��&t���I�{T*=(I<��J��M�5J�&C���IBY�<9�F�|�x�� �bI��a�X�<a��P�U��	��(, ����P�<��8i�$)���ѻfh�dB�	�	K��С��6�*��d�VB�	��&@2��=|�	�2��f^<B䉯��i��H
R���'ғ,���D��@�t�q*Gb�.q��f!�"O����R�&Ɠ�Es��3�"O�xx����oژi#��X9G~$� "Oz�E�#<��}·�r�]B$"O`x� �0/u�y �$Օ:@"�8�"O����:{����bQ,�*���"O�!����#@(�AŁ�Vg�YKg"O��f�Y/M���A.��hM`��"O��P�1+��=�D�Kۜ�(�"O���ȘV�1���o��	�"O ����ϙs�V�c'�ԕ"�*h�%���
GN�k��|�\�^K��ӄԨ���q��(�O����Od<�qK�?nh:��#o��"OLM����7�Z��U��{�N����9�!F���=~C�Ũ�S�f���ƕ��0=��^�^�#cJG�<Qw�ο@��肤�/���c��<��DK������,S��^�9�h�A�gߒZ�n�H�dސ^�~��K�01�?防W��"�x��@.�����)6?Qq,����=$���~���yu����R�q
�?E������__~r�����	 8���Ӳ$�y�b�@1݅=C�ɐQ��q���|I4! �#R�-Y�A�c���D"�O��H�[w<z����
!�`t�W�'�F��
��e8���'l���(�u�\�;�j�X����'�=l���S���Ӈ�3 �蒌y�1$��҄oہ���:�B�H�.L&��ROIe<x�0"O�Q� ]5,�N�?r3N�t����S������1�g~�"Fa�4��ˇ$r��P�@C��y	�O����#N�WS�H��x(˄˥s�nm��'�i�`
��O�@S2`�`�#x��:2�!LO d����;^F=�U0Oxy�6��,	�b�"�.�<U�\B"O�}�U�==��� �@�16D��A�5>T�B��ٕX]?�k���0Z�ۆ�"�"R��?D���S�P���\ 1��>tx�<��^8M��`n-?9�-����F��ڽ��f�;N��s���W�zdۑ�܉k`a~bjťy�tā�L��!��p�F|�GOF<äЁ��4�<�{��0c����}k3+�� k@l��?D�0FB�=3�!E� $��a��>�	  ��!u�?�"8 +�ZP��(�v��0"Oxl�#'�YQz���:��|��Ƥ>z1O�\[�3?�QkЦW�z���F g�=q���K�<� F�L�� ѵ@7&���Y��p��(
P��|3&_*p���KB�d=X�J�	"LO�C���$��-���acX)J�f��� �&B�I�R�V�)���w�>E�mF:���?�Bڎp���<�}���1@x9�g�J�� RN>D�K�Z&ad����3 ��4�����@��c��p�'�g~Rᙍ�H3f�# **8a��yRb�_�L�	c�4&�ᡇ�v-��5���0?1���t^B	���@�zۀ�k��~��H1� G�i�������fΛm�0����C60=���S�? n@s�B��k48���^�sX�*�"O��G��
�X�cT���5�
�q�"OP�j�?�V=����=r��"O��Pk\�2� �YD�[*_NU�B�q����'\��ꂅ1�3�R#>�@�W��i��"PǞ-�!��*FD�D
3P��M3��S���"��K�4�[P�'� �2!�/WŠ4��^�A	�Z��a)+>�>t�'��`�+ �i��iu#
J9<�I�'��0�$+דm"��d�^�2tЊL<9S�U�@m(���iU�O�0QB-ʅ������VL(h�'vr��3 ��u���B�-
',�L���'V>��JPĹ0���xS[��# �V�pJ� �.G��x��W0��0�'i��c~��`F@�Y��$���!}��z�2m�U�G��>{��u�P"��I�y�����$<
�"�*�5H\1n,rl#GF�m��ȓ��(+3f��y;��I�oѻn7��%�XS�ޠs�~<K�#2�$E�YPs_�b�jeف���`Ԓ��ȓ7:
`�CC�x������^��ą�0���Y�H��=�L8�Ǘ/�d��ȓF3�8
��g���J#ْX���ȓ���઀�f�@�Ā��W�Ƙ�ȓ?+�<Q2,ܡMv�M�5�� |>��ȓ=�&q 򨉺݀%㣋޻�4ɇȓbπ1���]ސ�҃�H�Pćȓ	� ��M�4w���k'�9B^��ȓ>��L�e��fB�6`dq�5�ȓ�(�:UAֲ.���2�<V��ȓi�Q����~�p����r� �ȓ5%��� �Q�4[& �2�J���>����Ci��VM���AO_���X�ȓQ}.D��G�c\�2#��Bx���ȓX/��/5C�$���UO�dh�ģ&D�����Ɔ6W�<�dB��$��2�)D��т�_)d��7�6)el{��&D�����)&��٢B)<,8"U�%D���"�X,)�((���-)���#�"D���#k���1;�@H�x�l1�f D�L)��.}��j�E
&l$UHԫ=D�Ce!#.Z�#���ɑ�I:D���GK�f� ��S�]�4l��	�,D�(��i��[e$a��o`��`�5,+D�TA�J_R���"�\�6����b)D��*V��i�d`I��Y���D�܆�yR]� ~�ӀK�Q�^D�F���y2����8���^�Q�ڕ�B��y�5'F4�(��=����D�
�yb��%(��Q*P�/�>�qCL��y2-�3�Z�����'�B��%�_��yrj�9Q��0G*ϼÄ�j�㏋�y��
f�Ҩbp�ջsHL򃏘��y�(�(y+րp�e-*�h�
� �y"E 8�Tb�ռo��m�
�
�yrAJ�+vX����a-
1�E��y��#�����d�Wd��ť�y��*(�8:6C
9E�h�$��y���\-���ԈX�'����@W��yR��� N�����\����z/ �yB��B��<��cJ'M@��q�
��y���Y�����>U��t��;�ybj��N��q���ĔG�"x(`& ��yb��0��pk�A8>H�y���&�y��-H� 9Q�n�C�q eC��y�=A�������j�X� ��ybD �mJd�H��Y�W���a@D*�y
� ���Ѥʀ
�q3E�	{�{�"O^��N�?vGt�Sa'4}D\�W"ObUyV�@�RKv��Vȑ�
$�)2"OLr�'�9��̋���z���0&"Od��O�jf�BO�+lJ�"O�Qbd�������.b�2%"OΨ�WNO>*'�,T�9v�����"O��3��D8� ��$.	q0�B�"Ol��ǀ43�e�4c0H �"O��B�^2d�U��\�f�~�X4"O8�
�G��Z���T�U�T`8q"O�`�Ѫ�V����e+B�{eйY�"O� ��d��)Ĝ��3醍W+�5�U"O�P� �[�xI�d�˧,*��ذ"O�1(�d�B T�x#�Q�R!�YF"OK���Wy ܣg�)336(Ҧ"Ou�bi��:�D�M.���"O\�t&�X{�� ��5+^��Q"O��	B, J���,g,8�'"O*�`�eG�J��}�d�,�d�C�"O��s�iR#,`X�ZF�Is����'"O�來�TOB��
I�Ѭ��g!�],v���������̍Q�!�@1>qM��I�[����FjO�q0!�M?;���{�O<q�T�	��!�M�X H��ԉ�0f�ƀ!6��*�!��ݚv�@�p���%�zAaԦ��<�!�dĄ�����Jw-�� ��éx!���2�:et��&H�ԡD��1�!��X2��o^)L�,hH��2!�J� �x�Z�5Ѐ)iG�1'!�DB�}�H�� Ƈ4�pU{͛
!�D�ch�k� Y�S��{0�/�!�Ā�	g$���g�.��-��Q#!�$)=R,aP�-̀P������!���1���r���l�HiQ���!�$��R��%y�ʍ,-���*Gk�>$�!�dA;�2�QS���l9У�M�z�!�d�	��Q�c�8݈�P'�Q��!򄐌6���'eT5'2t��혜^�!�$Z�/��9�G��ZsReӑm֑F0!�B��\���蚦)Z�d��ŕ&3!�d��%���)a !��U��Ŏ2J!�d�A�<YK��-�f�fG��T�!�	 ^�0#B[��9"5$�/|X!�䙊B�f1��j��]}%�fA�I!�F. �@0cT v�у�A�[/!��N�r�A b�i�8��l݆-!�d�(xu�׮Ov���-X�!�J�?��]*��\�r�gT!Ux!�$Բ|���`�=w�<,(�e�*�!���Tꆍ�TC��n��� e=\!򤘿G�ŋ��_�VK�x� o��O!�_6���ꄊ��U:���c.F�
�!򄏫"1�B!�/r�<=��,��4X!� H�P��Ah�pn���K�&nW!�D�@ 怪�wXhZFT]k!��	K��1Qwaȫp�� B�67N!���Msp�S6U�����*~�!�ĉ�H_��`c��%�N%�R��=4�!���Tl�y`�B�}�.a��}!��#�@�����x��lh���B`!��S:QWba�����McU�=hK!�"`��[��7X�HA�W��'>!�� ܭ1��Z#AV@@
�9C$��g"O.x��̓/;A�
�HA>y,,p�"O���� jI���ӜV]��"O�D��cS'8d4����ݻ53��D"O(!�O�7-�C�C'y+\�ْ"O*��
XM��M���X8p�#�"O�}�%�FLiv �w�;���"OV%�B��	QA+#���{&mP"Ov ��ִp p�M6'�会7"O��sff�jP�����1c��"O����P�>w����-��Jh�!�"OF���֦+߬��7��1 9ry8�"OZ���I�t�.Ua�,ʵs�4��0"O����䛍G0\����/@.F�#�"O�Ɋ��X.Tb�}��e�X�x� F"OX��Ċ�t|n�Q��%)ϮY7�'Oў ��h��eF�CQ�N;\Lv�h�J4D���K��<�H!B�R��DI[G	1D��*0 +{Ԇ�{�%Oi��y�@*D�<Qk;(�<��%�5����B/-��p<y iKv4M���K!y�80�&\W�<YF�=��pA�	�c>X@�V��H�<�q��j��C٣����+[`�<Y�������!֣O���G/u�<�U�R���+	�qC��¤�Rw�<A�Ί+
�$%��̄�8qZ��t�<��[�����zn>�+��u�<��F!%�Ҍ�w�M�D`����y�<97c�$�2�ja�;Ev��CI�|�<�b�G�rM �� b.�ⵘe��z�<Q��1^>V����Z�VC`�8�Ɣ]�<a�k�U��y�>=D�S��	B�'7ў�'Wʖ���%8��ˡ
�<o|���ȓC�>�S��X.4l񄅻T~Э��;���y�I�<��ā�.iŅ�Ic�%5�(�%G�-{��3�I�(3��E��R�1��޸�l��b�I�L>���ȓ0V��ړNH�e�����W0>	��-�0��ΎQjK�lZ�/	(��'������" Q�x{�͂��\��L����LQ� ��m���5:�X��ȓ�&m�nSQ:N���AB�i���ȓa@ب ���}�V�1�U5.��A��($0�C��ͤ_�Da���d$���j�r�82��|�4tp&ӣb����8"Ds���u�)�(������&��8A+�.q�b���͚N�lM�ȓi|�y��^���"`і:"��ȓ����KJ'_j��p����5���u�������'tЄ�M����$�ڸ	�^1-��5@�g�1����q�����M��W/�)o�q��z��"E�T.]��G�(�
�ȓq*�eH͏7xD�s�� ^Q��ȓ[�8Mi"�3){��SV�;C<���+�����8tr�	�clO˂#�[��hO1��Q��o4pur��ŤN��� �"OT�A���l6*���h�,��a"O6M3�kޢ]�*� 1G��X\�"O$�p�(k�"�¤�8���!p"OB�T�ح�క�+�P�	R"O�(�#n�1;�T��Jݛ>�6���"Ob�i"m�8��s�E�p"O��#S7\� �L!�6I)�"O� 8Y�6�Űh�֌r�%W)4�¶"O�e�"U&������^1;�$��"O�0"�,���x��M� b�P�S$"O&yBU'�/eP�8�˛�M}<5s�"Oti�̐	vs�\�d��/�x��"O�%s�Z?u�&�qedˁ5��Q�"O�b�^�MÏ�X���"Oz�t�LG�@e ��]�(+��2@"O*QK�h�_���;� Ӽ)&�q"OR���7 �]�ab�1dh\�"O@� N��.����M�,8�"On��B�37\���#�<{����"O��
Um]�j���!�����Br"O�h�l���6K�T;�!��"On�K��^ 9��� 4��/���0"OzW��5!3j�	���1#\�3"O&͚ �P=$�%i�mL�Hڭy�"O��0D��- ����	��ȁ"OFĹ���rK�LP@K��f�u "O��xPK�+X�F�T�C10�5�"O ԫ�>lԩA�̎Kv	
�"O��ȁٓ&�j0�b��
#; =��"O�}��%�)���)��O� x�@�"O��%�W�D����$��(�	���'o����� �Q�|8�A�!��U(�B�I$O�B	�B�z���HwFɢlJ�B�ɸd<i �f��C���jQM�1�B�	�D��m�,�p�{�%��?TlB�	�UT���Fe	%+��A��[&�6B�I�RSh�{ׁ�5P���S兜�6Q:B�	1V���gЕ2x"�!Y�j��B�	<)m��%I�6vp<�3d�+Z4�B�ɬ?�j�KC� �ib�15nC�	>Ұh�e#/5�t���>4~LC�	h�NňF�>���K��+�DC�	7L���f H�Kc�HȄ-�;pC�	�	�|�*�6E�|@�a�p�B�1]|h)w�B�*��!
�5BʰB�ɪYg� �7�pm����S����`��<����fur�E�?\ub��ȓ1z�}�Vl
=	# ��!L8h&�-�ȓ`��-�C��	%��L�t�M)5�Q�ȓd ����Y�b�j
02�Y�ȓf��Չ3n��fB����	��e�0��ȓz����)H.* ΍!S�W�i�����رj�#��>���Q5CT�ȓh1"	h�I�b' �&�ڳ%N�U�ȓfn�p!�H�r���(Wb �cL����D{��Œ!�]iD2/-�-����He	BN���Q'�ij���ȓXiN���T/z�ltS�φ�R�~��ȓE~x �K�B<x�� �W>n͸����|�Gׁ9M��j��C�`Lh�ȓO��ŲGL�*p�r�J�b Q�	������'�Ę>$��RB��G`P��� �"�@�%%@ܜ�p�H�~����ȓ58Ƹ��\�1�ƭr�&�Q���&�P�i�ibH�:��G/��I�ȓ���k�(��I�~ȡv��T���ȓB����P2�>����f_�͇ȓZ��J2#N3T4p���ͩ6�D�ȓ��h0�̛2]R*�c[�k�Є��d4�`-�0 {~i�� .1]��$cr����H=c)b��D.�m0܇�S�? *��.�Y�	��`'\�Z���"O���B�:h
,k���@D��"O*��`�\(#��j&o��@��"O&�:c��2qb5� @6�t�"OH�  L���D*GÞ/N$�5��"O
50��ʑt ���, �M��� "O�={��ZCb�Dr�,��H�̕P"O Ii��"a����Y�nDyW"OV<! ��R��樌	�&��"O��c�̀ �4T����0W����"O����`�5 � !lH�)�JQyG�8D� ��3iE���$��[:E9��5D���G��3u}��Pw��3>X.Ma5D�Hc��A�8/��q
֊Xg��4D��[�KM#I4\II�ԫ`#�e�EH0D�`���L:��0#���+G`	:�-D�l�1o޺6s����Ϙ�&�||���)D��A�&�9|�{��C&';DXpR�<D���$�"����R��<d&2T"9D��U�UđbǊ\V�U��$7D� ;s�>V���q��m�g�5D����Ҕs7�x���X+|-���3D��RE��AB�Dsa�	3H�,�W�=D�P�$���ty"���F(N��� D6D��B-�:%��P��ŽkrҴʧ7D�p郇�$@6P�5�4����+7D����j��ִ��ر^��9ӠH"D�``�"��-�r�y�$��H��-�-D�dB�/�3�6�kH*df���C>D�X���5B�p$�!F�~���=D����eɐH�]�B��Rv��<D�Գ�@�e**q bb����Q�b:D�$ ���@���+����y�Z�Z �"D�09"kԢFC�T�wg�'�\�꣮5D��a+�&x�4������[0���M4D�4ca�P�L��,c񁅚S�K2�6D���S-�'�N�����"o��\:Bn!D�$���[v��P6J%{UҰ�S�=D�
��X�E0�sD�]�`�ڶ&D��"e�J�ME�Z�-֏o�b�p��"D���f̌Z��Q�s���T�@��!D��/	?�0Q@s�\<UD�$?D��A	U<��ds�-�aVB���n*D�(��c���t�7��;]6�³c5D�����P ?��E 3��8�hI�K D���D�&R�<�f��?Y)B�[��>D�8�1i�-s�(Q�wǫyw���?D�L�"�շ~|e{���,�
�H��<D��h��0T�x�G A( ��t@�'9D�,���g�V(�f�C�W�>4iC�!D�$��/��hPR���Tn,�`I2D��*��G�-����kug:D�l3�G�O���Q�[�0Z�8�%4D�d0�b��w�9�*Ү��V#3D�l{Ԯ� E5�BC�L�4�S�I%D��1��L=��xRw�۱y�N-[��-D���$%,_�j��G{9TTr �6D���(^�;�Ƞ��ڨo�2�@�c6D��c�_�O��s)�3&���F,3D���dҭJ/PQj51Tu�
4�$D��+�̖M� !�A��'��8�.$D�X�i�<����"G^�:j�\��#0D�8x���^�h�ia*iܤ<��!D�"ҏדo&��! ܕ	�b��wf+D�� h�5�Вjqd���ζP"B*�"Ov,q��@�{�Q�d���>,y� "O��#R��Hl��FJ'$�A�"O�Y8�+Sprxhٳ��V�%V"O��{b�V^�
و�g�Ic8�"O����9Ii�A�FT�%xx���"O�|�̗�#�n}�҅M3)eD@" "Ob�Q�D�4W�0x���]^^���"Of9M2��A��/�n�V6n?D� ��GD�I��B�O$�u�� =D�Ш�W8S����̓'3`��':D�8#E`��d�k�'�W�AQ��+D�P���ߎa/P�S��;�@���6D�t[�̔��Y�F��"Uܱ0��8D������TZ���D�?3��u�q�:D��hC���D���F�K�;�Tc��>D��زDzB�#��G,rN�A��<D����(q�H[�BF�����ń:D���/C�}?��0�B�pD,E.4D�sQ�*V�x}p��߲<m�ab"4D��Z&��$Qmx���/V���%�3D�@)�M�8��=�B�%:�vX���6D�0��)��N$���.�3^�`��b4D����.}�d1@�%�"�k��1D�Tѥ`�:?0�Fj>X�V��3D�<�h\���\k�
A9vk`A��A/D�B!I�a������s	�.L!�dV��"�!'�\afH ;!��C$=f- ��۩ D�6g�}�!��9J�`s� �6R'\Ȣ0÷m�!��;f���`l�\PŪޔ"�!�$�	l*�q�,� "�H��e	J�K�!����� �)*-^�iI�!�Ĕ�5*$���zh�ѓJ��!�C�L(Ӭ-/J��r���H !���hb���w�
�p�����i�!�æI���+5h �2��s�����!�$�4Z�l�)�i�� <#!�T�l`ZB��g2΁��@�!�D]8G�3i�:M~��"��3q�!�+	b���C?eV9��OJ�!�䍑T�kA��a"�����E�!�$��(k�PY."���.9�!����ꕁVh:t�b�֣�8B�!�$A� �h���3#�ģ�%� Vl!�E&/�H�&̤0�<��$�V�RO!�d�7w8��$hJ�A��YB�զ2!򄟋(���!f�IY���p�O62�!�$4RG����G��j�xv�٧[M!���Z�nICF�S Xr�b�5:�!�Ĉ�7c�Jv-ܘ����R!��n�X���:�p�v͡o!��]�T�T�P&K�I��D�o!�$[y͂�����c�V�Kq��R�!���[?����,�~�v
�k�5&�!�d	=B���bƊz�n�#���H�!�DU�LmT��"iU1B�^�)��ͷ) !��$?�ޡӓJFh��G»V�!�DK��]8��э	n�Jc��7!�ձ[Mz}ڷC�(V�h�7�7D!�$πCZ����Q�>R�]Iv�##2!�dQU2 P0j	</A����
"!�9k=�e
A�]�-H�R�.��Y !�DN�,�`Ycmޠ|�M*�#�1T!�� v����?X��+ʘ-v�$"O��ڐ���U�.��#+��:����"O|�
����~���&)�1#�~`�4"Ov-��#��
�*��D��½#�"OҬ�E-
#K�� �T�-�~
�"Ol�ӧ�m@"Q�a$������"O�]@���$��J��T(�D�Z#"O@����T8:h���Н�.�a"OT��WF�6M|���b�$����"O|%���[��0����ݮB�:��q"OP񩖇'c&��G��5t�@9b"OD�!u���)e4��O�PIyw"O$�3��!w�z���*�V䩠"OR�0�Ɲ�tU�=Ф#�dA	5"O\��}Kd�BQ�	:�<��"O�4��D�O\�Õ��.���C"O��cIV�����`B�p�Ҭ� "OT�&��gnT�@̑?�b�"O��Z�@0�F��RV"�bT�<1���#d���n��]�yCǙg�<a�`�r��@�t��s3�M1���e�<����f=x�J'!��-Li#�M�<a��V�p�X�qC"�G�\DIb��E�<)�a��
�p� AL0�XW�<Q��C0 0 �A�u��QeE�S�<A��A�S���`@�ϋ�r��N�<1�M7-�>�y�&C�~gHaj�h�d�<Yl�0=D �W��8�L�@�΋a�<Q'B�i��=�2�+<�r%N�f�<�&��>@mR�#�&]��i� �h�<�a""���EE!<�u�"B�k�<� ��Z8qf�ğJ~,��!�b�<Q����b������@C&�[�<Y���s,.)�#�_�<`̥A��q�<U�I�O{|YR�C'g��U�n�<�%�7�\�B�!¤y�����)Gh�<��fO�W��!���)h
��7��e�<��
3=��s͉�F�ၧ��L�<��o�8
1h�p Ļs[�0S��P�<��d�?Y�|�P������L�<�fCQ��3��9)����f�D�<��kA%T+��c�lۏFr ���~�<�` ;|�iȀ+ր���R�|�<����e9����GQ�:(�pb��u�<��40 ���*X�Q��X�䭇u�<ѥ�� 0H�1�T�6��|a�o�<����n��Qц�UWr@	�˜m�<!���X��
��|0��HR�<� M{)��|	@��ao)#�~B�I�1:�@�N�5���e#A%&�bB�I�?��X@��@�_��C�ɧ|��I���onX�ZE�BE�C䉌2G2 �wNH�,T��N��&4`C�	,G�uk�"c04��BIP�6ÄB��/ R�փr��U�fL?j~\B�	���C։@�d$��Js�,	�"B�I��&4ۂe=Qx���AQ�T��C�	S�4p0V狔]j��)PNLM�C�Is�B|0�(Q,"3�̑Sk d���?��?����$$@F�ϬR�M�D(�
�y��.�j�'A�O3䨨n�6�yrm�U�②�d�/�B��v!��y�6 h�yj5%��R�+&����y2�N"X�f��E)�\��Z�0�y
� ԝ��&��@��f�˳i�8���"O`yaDE�^�p��7�^�j=�t�A�ILyR���X)��g��$�PbC�Ke!��O0o' Y8U�I� � �*g�ǀ~T!�dS	���Њ�<!�8Q��GC!��	�[ލ��ϖ�h�����,'!��#���¬N�\ϲp1'KX�!�dX+dA�xb��Q�y�d��jP�r!��Ӗ8.Xy�ri^�*�"���FAQџ$������|�B6�T�{P����D:pM�P�<i�C� ��I��M���Ź���J�<i# ��W��Dr���B���S3�G�<IP�I�4�:���ƃ�4����ĨJo�<	RF�2�6@+��D�0�;Ьu�<�SJ�6t�����c0�	��@�m�<B�+ .p���ܢI�2��b��l�<���R8���Is�US4jEs��'T��
Ս΍kf���1A8s#`٫U2D��+U�}R.ðj���8k�J0D�|�e��4�j��^�q��Q��/D�p���u�ƨ�p	��YC�]��/D����-j����4�וhx)�4�,D��q�[U4$:��Ŷh�4*D�6��B��k���V�X�b��NL�<a�DRCR�ڲ��9u�x�9 ��D�<�Rg�<�:x9��R�����VE��<94C�x��
'Hҽ+�D���V^��%k1D����h����G�#iI�=�D%D��yg�Q9\�.(@��ً��-)�A"D��� �@)�J ؿ
���*Q�!D� :���{X@��A%���A�	-D�h�j�q�����D��l�8�)D��rV���~����kK�hsׄ�<�+O����#��)�A��&��c$.��q�!�ĉ�FA��㳧��#�0��G�#�!�dѾ>�FaʳxhXl�#��wt!�ڿOzRd�!�(� TsD��
b!�D�>\4a�����A�f�ZsU!�D�o¼�K �C��!�~H!�r{F�!����h�d�ʸk!������rr�ʑԐЄ.l_!�d�[�I� �L�Ftb�ퟋ,�!��Dm@��! ,	�*"Ԡ����W�!��X�ıb�R"	���p/F�E�!�4c`�(�jӬ	��xQ�ěOg!�d��a&�!ye���^b���.�.D�!�D\���[�I�|��bpm�)|D!�䐿f�@�0��)��(�k�|�!�� S�z(���WkUd24EܒQ!���r���(+7�r��Tj�$C!���	A���ED�<��3t�)!�$ľA�\�A��R nJ5Q�Iў,��I,9lK�.�0u�0�TJ�3�B��e��p`0zībkK�,���'�S�OR�e���+phf�R�[�	>4�+#"O�2���*fm�I�G,lPJ�"Ov����{����P B�]`��"O�P�������J0"�&��"O�,��fX	Fl�h��"9�L4k�"O���ʓy��V��-����d�|�)�G�"Q1��"e���Af)@6���?�S�O���S�Ɔ�|���:�c�
)�F��1"O��pa����`���Eu����q"OB]�PC�*L�u��)\#��Q�"O� �!�(=��(S�^��<M9�"O"	��Ɏ�Vk�d�C�Y�)OL�X$�|��'���>����0HI$��d%��{ c�<	w���p��y��H0z��M�c
�4��|��|��D��
´;��+�H�b�m�<2�!��5��d�(�����pOF�s�!�ϱei�D�c�Aw{`4�$�"!�d��� gM�Ye��"��L
�!�$E�������� D��!���'�|����3WW"I�U,�8���Ȳ�4�vC�	*Q#*�˃̒����z��U:���d�C7�"~��bC�����'����k9�܄ȓET�ຄ�,^$��B��Tk�E�ȓw��C
ٿuo0e���%�Vd�ȓ1�0��e�U �Ar*̞W����ȓv�2��W`C�ΜMQ�l��l7:��?����~b�%[9(��j��
�`�`���YB���hO�'
8�9�DA�.q�HU��'o�6�[wl����<E��'�0i
�(��?��=[0B�\�b10�'�Xܳѥ|��GH4M�>���'�yxЯ��n�"�����?�4P��'sDt�Q�ݘ8���C�31�t��
�'�l�@��ؙ@e���@	��W��1���hO?!Cg��b���4`}��5�h�<	c˂�Mhek�ծ=((�BT!�⟐F{��ɚ;;���2
F�M!lUcD��)FB�I�'^fܒ�%E�c����C� t$B�	�?/���m��P;�]�Sn����C� S&��\ %K���C řS�^B��dM�$�Y��a�jX�˚���;?y&%�rh=33��K6t��ey�<y&I
<��qӁo��e���&�Q��`E{��)�h(i9u�P�n���jX�4�|C��-$)E�R�)���� .�.x�C�I=!��q��/͗ Z�M��C�7��x�a�<$��Y�GB���C�I�E���w'�*ފ�CIڔrӲ����O��ɮ;���y7*
����B���0�zC�Ɇp (��Yn8�@�V��.,�T��/�S�O��Ic#I�tډrCL����v"OL����Ӓa��u�4��+H�:�;�"O0�Pr�M2d�,�R�� 8DV*e"O���q��)F=�HDn�$��W�'���"G��$��J?T��w!�?qbHC��<	��z`n�T��`��-�#�nC�&�*���ؐk�h|�Q��1˞��Oj��{�'�v x�@�YI��Aqc�g+�'�f�؄��7Y�dq�	��� ��',5��D��4aES{.�L��'2�0�ԂXH�AP\�o� y�'���+�g#$�\ P�,P`��8��OP� f@D��Y'��r��"OL�:�e�]&V�Q��&x���#�')ў"~����)
0d��L4Z�đ��P��y��H�>��£OB-Pm��9t���y�)+G���c��	<I&��/I��y�A4�z���K�lp@���K֕�yBd�F�ڒ�!e�����%�y
��Nm,���X3gG&!q&B7�y�hC�<~�c��\��BA��y�A�|��ԤV�\� :���yBd@�Xc�|(�B�Lx� q�ė��y��?>X,�`K�G���U�Z(�y�h��
hIрǭG�"\p�I[��y
� h�c�"�.��)���c�J�{%�	\�'8�hCF��v��:��
�`�+V�'�ў"~"��W'7��k��O�y*ѳÜ��y��>.�	��_ o�
�R�H��y��=C��z��e��X���y��ٟV�^l����[ P�1
��y�cܐyҔ `���L4$��)_ �y"i�'.��(�"U�w�|!!M���O,��?a���T�UB�P�������$P����yR-�V}H%Q�ʊV�|�nS(�yb�
�7��iy�D��N�\17`�<�yBHݲ4��5��,G��5	4�Q�yRUd(P9RӤP�:;@�s&��y���?.T�i��o�<1�M��g �y���38�]��#4y��t0�����O���.§4�d����L�s:��d�א8%聇ȓ���� b��MU����&��v�z��*�.�D�Y,��f.��[�TD�ȓi�A@$å��8ۅ5"��1�ȓJ� i1�@@�~S�bƯ'^�����@�ۍ7j�D&^"�6��ȓK%��q��T(Rٺ�@,�,�F{2�'W?��/�3¨H���:@s֙x�N4D� �Ao�5!���4R�Sg��2f�,D���D,��A�������A�%D��j���8Ch��z�$0D�� 2'�h�TԢ�,R�1%���7�8D����δ;g��� #���8U.8D�,��	J�~�z��O��v� �<D�X��ȬTDZjpKLI�J4���:D�p:��Q�]0�PA�--$��ah9D� @�nÅu�bXɞ�3�ꝑ�<D�@��E]�IX�0��m��bd��b	:T�02fF��4��cQ*u��`�W"O0X Џ��"J�:C�
��-C�"OP|ۀ担q�N����J�n��Tc "O~-+�^��p RT�U�]u*�d"O���j��|j0��/8y���"O��À�M�E���FN���F�y�"O:5�W�g~�5���ϙZ��YA�"O��0��5�~��2Iމ;�%��"O�8�` ȡ^^��g�"���2"O��J�gV�oh�:UȂ|�@��"O�C����M�ȍ�1�S�K��l+�"ODi�D�0�"��䝩5�x���"O����>l��*��C�Dn��hF"O`���F"^�A���3GLL���"O&��j�V���[����d�0@"O���%&9^�F䡤oM�[�d��"O�<�hu*,m*g�A�4��"Ob����F1	}�H��Q�&���k"O^��C�����H)f��E�x��F"O��c��#�LxP�NRV����f"ON�@3ژ1�H�$�;z��r"O�%b��3D�M�#/�N�����"O~�)�+8(Ҩ#�.��'���6��Y�ȳ��i��}�����nPS�+�D�O^��� "Y]D��ކ4��3d"l'!�Ĝ�JT��|����#�
e!�	V�T�3�N {^X���aW�%�!�$�0?/hC���z8|� ��
4�!��лz�|�Q�똨%&��z�V�1W!�;c�nd �Fk�8�"\;�!�$%�Ԥ�v�4A��ҁNC������Iz��� ^�J��E#p5f��$��2ȂuYW"O� ���;��a���W,���	g"O0�+�5-�B����MB�X%�"O�z�
S6�hL`�Iʜ�Di"�"O���f26z��5N�%TD��"O
��F��5f��r�,_Op�"O�Y q��+X�5,���	H%	E�m��Q�H�S��I�{a~@� ܋K��� �ϝY@�C䉋A8���СZdJ`�4�K�1/�C�I A������3��١'ʕ�(C�ɹScT(����!p�!ܕX�FB�	��H	��ϙ/�ڹH! �6tB䉺b��2'd��<h�xP��;:$:B�	�L$re��G9�,l�c��	v��C�#Q_����L2Yn4؁@iԉ�jC�I�_�F̱�J�����w(Q"�dC�	�k�&H��FS�	[ȉ��,	��4C�I�Gz҉���Wy����"!(�C�� Ӗ��W�V.|�k��Z�Y1�B�I*����`D� f�6K�%c��B�&3�J��2�ۓ-��@�ǓNFB��o�ٛ!�	9L���d�+Q�C�	����G"A� ���ƍ�Da�C�I/���!"-ҋ[��*��L�Q��C�("*�����	��8à�
�uaxC�I!<Š�R���b�\��cE��pC�IVT�(���hGv��򤈡z�t��>��|���
�jw�u`��]lGƙ e��8�!�� y��y
Q�Z Q8��wc�8H!�dџW��Y���%wN��RGiM+!�Dч�Hy�$���K2.�)�I��!�U/0�3��_�z��Xy��R�!��ؠ|��Ĉ��;�l��%��<�!�dEP�!�E�$A��vH0�џ�IO�O�B4!��Q�N����A�D��'�Ĥd
�Q���Q�:	�
���{�J����`K�+��u�!�d�&<�&���d\>V��ѤjαXD!�J������\�EE~Ux@i�N!��ؘ�����M�f��E�ah
��!�D����f��%7i�Y�ӆ��'aa|�
9¶�ӄ��`B���y"��(̜� A"�����2�ۗ�y�Dޛ"�0�Kd��b�D�B�Y��yn�8�����j��T��\�y�����#�9ic�k�cF��yr��$e�-iv�(u&za,��y®��\��5!�2jʪ���g���'aў�Ov�
� �1-Ju*��ڤG����'�d]�
^��J��S2"A��	�'��ӷ'�
�a`�#t}��'n��Q�M4$H�����	�z���'��=PP��(p��3�k�#�<��'R�l��L?~씋&
ӡd�V��	�'e"ećX@���EW)Y�X�A���?����������K�� 0V
ŀ�K��һ B��m��$�*F�7i@�f�.�C�ɨ+�0l�sD���	H�Ş�k�C�IT� E����8Rj��OپC�3	Y����C��	�̀	dٮC�	{E�m1 "�̨�d�W�B�	�3�ni��� ~�t��A	����E{�O��d��TT�(A��f*��B^	_3�)�'*
&�
���-h�@��Y�\��LX	��� >h�4E�"6���ffI�II"Ox���bE�E����Dȴl��њ"O޴�ƣ�(4�zfe�(��=�"O�I9�Ja�b�"A.��.���"ODW�h|H���Xj�����P�I���OC�� ��aqD�%@_)K����,O �D1��p�'� �c=&�(e���ݴI�$��'�n䢥��WHTh�"l��Cs|L!�'	ɘ3��uVH��ʞ�?���3
�'�nѐ��C+|���e��>hZ� 
�'��ӧ��� -���5�K�2>�h��'(Y�h�jؠ& (�̂��D*�`�I��B;� ���R����'�ў"~r��Ϳ4�v����(Cff$x��yRH�j"��Y�`K:wz<P�Î�?���S5X�|��͓~}fe�Q�Y�^�B���a�8ѸrG�) zN(�D-�J��ȓ&z̅ I��S���(w�U<z1L���F0��Pq��F���S��R7Zj^��Io�IVy���G�(&�p��+[��E2�n�(��C�ɸ9��UK@�ΏU��Y�a��e�B�ɖ
W��dd���	aFA]�wp�B�g�(�rC�ɒA�H�h�ۏ ǸB��5JN��¤�V  m����^#�B�Iie�)*��Nh�TiiA�A4��B�I(#�����!M��y��ԏh�|ʓ��$��)w����MA38$e*a�"�R��A%D� ��S�(���1�dةF" D��kp�Z-_�T̛v#�"�h��ad?�Il����	 Pp��#i�2Eֆ��adV�LvB�I�fH<�g㍊)����a��#�dB�I�M�����K^d�Ԏ��38B�Iuʘ�zv�0*�L�/�:C�I3_zpuHs��wmn�ɉ23�B�ɝGw��rE-�fi���H
��B�	�K�IH3Ɛ��P=.")����?	����S�O ���rAX��Jq�RaNd��'��*@��#�R0/�=X�&�P�'zv@� �R���'E%A�*m �'��	GI��V��9�3���8���)�t�������'�59��x����䓺0>�5��	
��\)s��V��v�<�`G3F𱒇� {����b��y���hO�'��,!̟F@n\��VD�ȓb]�qG(F.8�az�J���LɆȓ��d�3*D�����e�)Br<�ȓ,�Z���)�*�
q����1:�2��?Y���?	��IL�c�
Ա���� �sp�,(V!��4	�!�e�߹&�j�al�  Q!��(W�[ԉ�(z&a`5���Iğ��IS�)ʧl[���%Z$&{p�Q� �N����c�� �S�NUjM���X5:D�ȓʖ)k2Ϙ�EP$iQI��y��1�ȓ8��"�G6�j����(�G{B�O��1��i;I���Ë�f�ՂM>y���?�t���?�b�ձ��Os��H��<J�Ju���Z�B�H
�'�0:4�
>z�mX���.>�^I�'Nv$2�I��ܽ��� "=e>�I�'����8\�Z8�J�9#&��'<�ɣW���kN��# ��>'�zY@�'�&���́	�dç�ėLR�9�'Q�aÐ�@�C����W+�t���S�<dExb�'���xp`ۀm���#Aٚ�y��G�}�(i�6,o��\�@���y
� �0+��L�s�� Q�^�~�|�c"O8Mj�'�i����C�09��i��"OR%��m��T�f�h�m�"V<:02"O�tу�'���C�TY��T�'�'�O^��!?�);���ᢘ?{@f�E��P�<1f��6N���J�	�:Zl3���h�<a�$ό�@�!L�cDݺ��{�<i��X�lRX��	��z�e�\�<Ѱ�{�0ZB�f���u
FX�<�QÕ�=��PL�|�9p��V�<a@�K0�ҴB��Jz�(]` �V���hO�R^&�a5�$�Q�cLn��x�ȓH.���J��U�F8�-�Zo���	_~B됪W�J�R3`ʴY�h(�t�^��yrf� h��[��Y�"��GE��y�'ՠjƔ�Q䜛W�� a�)�y�[�M��9��P\"�fٵ�y2�ΫN��@2��[M6�kl߅�yRn��3U�T�'S�E�ȹ@5%C5�y�N�5gs CI�P�h��DGۆ�yrd�2ڢ�(�ʜBt�X�êT�y�Hٍyr���@ϻ?�Q�")��yB�лz��Q��F�<�t	{�$���y2IK#M�A�#M!6��U�a�X5�yҬ�df�#�
)3��	X��y�Ƃ�v:���ֳ1�$�Q��*�yҢѨR����������B��.�yBL��z�2�A���a��oE��y��L�!>9Ġ�*>�Q����y��έ%��S�I9N�QF虑�y⢅)Gtz9��#�4�ڴ���yR�؀EX���%ɕ@r�����y�!ߓU�ܠ���t���aumM��y��)P��Cr��>���t�P��y��[w�D��46�&�s����䓒hOq�n5��0��)�F�i`���p"O�)��"��\q�n��r��"O��j�b��QrT�Ĉ�"O��1��E��Z踄J�?��p�"O��(��\8"�Ĕ�E�PN���B�"O���a�R�`  	f���_ƶ�QU"O$eB0�F�q��oS�f����&���O
��&�Q]~G�FS�D�F�Z��	 	9#��Q���5aC9A����K���Q*		N���b��o^9�Ɠg3�"Q��6om�c�oT�KҮ0�'���v�K����Β�<5J���'\�ppU# X(�Aē�/�ȹC(O�$/�O,��M�
�z�j�G&EL5�5"OZ�r&�O�����:5t�"O�(9��_5�
]k��?Q�=z�"O��� ܕ0���񁯄4D��iy�"OJ���h�
^$��R��U�:�(��'R�|��اdע �� �4��9sdF>D���&V� ��ȡ�G<<	����I!D��� �_�p�p��--�n�H��,D�l0�
3R�`�ǫ�s�`��4�,D�X!'��7;��A��=U���H�*D���'�ْ�ĵ2Q�Z�	,%��(D�p�!j�$�NE	ŮĴj�V�{u"�<�I>���O��k��i ����ƙ40�tB""O��Z���U��\r#��z���1"O@����L��
Ɓ�AR�3"O�`��C�&!n�� �;H����"O� D�`��W*ty�$��&]��ku"O�4iVhJ�*�z�#��̑VV6��"O�\``E��U8D�B:!Gd��a�'��|"�)q�ƿQY�]����6�x�B�5D�����i�z���D .e�f��$�1D����  �Uӳ�\��N�K��/��B�����c�n�SS���.�}+VD1�C��	f� �@/θ!wzy��Mr�tC�I�A���� �.ٞ���+L;H�~B��xON�x�n�[ll���G,:B�%BĺI���Ww7ZD��K��+А�	H<�'$�k�P�h�b���|k����<AQ����g����#��� �q�`��J֦㟔�	>!sU�'qd����~{�~-���5D����@�� �۔k�`���!D��
���Uy���]�\�2�C��;D� �����]�$X��nێ5޼ᨦ�8D�8:#�X����*""M~ VPS��O���8�O~Xg��O_�	#R��*o&����'!��$.�Р��˹C� ���aéL���r��`b1�+:AL�͏�_ɬԅȓ5�@��h�8���i��z���m��c�9�Lиb�\F��E�ȓf��Tҵkɐ����ǗU�Ṙ�Yq�\Q&���
A�,y�$`�'�a~�n��`M�H�NLي%HS4�y2A�M�89Q��w��52���
���hOq���x�6�
i��	8�����"O �0ǃ�����P̏ ^f��A�"O6��cË29��"�=6=5j!"O2	;���>d'�KP��o?�MZ�"O�<����\�HФ
� Cx�3"O��)�G	$M�V�P$�ۮ%�n�(�"O$� ᄆ-x����f��X���q"O����c�#��41�U�]P$"O�e�� (-��8cJ�1U��c"O�i!b���}�w� w�,�"O ��a�4��	�#(R!Mn��w"O@� �� �Bݨ@�ӌ9 �(�"OZ��d�8=��J�>a"0PB�"Ot�hN
`D x$�_$%��d��"On��r��!4���dH�e�1;�"O6� teπT� ��Ħ��D��"O�̙¢�:����H�'Ά�{�"O�:�@U�+Ɣ��N�&g��1	D"OX`���4+Cv�k0�_��΅�w"O�tk�N�>e�*�Fѽ��c�_� ��g�S�O.-��	�z��Ր@�+���'����:"�ڹP�ˠym2�C�'�,,ɲ&Q�����A3�,("OJ��Qn�6L�P-�ƯӚ$L�)��"O��� V-%v�Ń%�I�FMd��"ON-�S��R#Z�(wMĂC�(�;�"O�=���(���ap,�v��FV�xG{��酴^��H���G���B��~T!��A%-u�y .���0y@`�S!�d�?BZP�) B:z��$��[�!�N!p�؅�� ÄZR�W��1N�!��>mܪD�%N��$Y�)@W�!�݊J��E��)�;o�:�'+֕k�!���K��E�ʹ
�XسhY?c�!��HZ{�Y �p��uS�4u�!�$-/�u�aϙ8���IW���S!�D��*ފ8p ���ꨲri��%�!�� �c�Αg��t�Eg�8%
]0e"O��Y��7ZT3G��2��Z "O
!�*Әg���Ae�U� � �"O�,�"J�iX�	@ �N�B�b�ʰ"O��0d�#F��l�s���fc ��$"O�D�AE؀F�81#Q�\pd�0"O(��"�X��tR"��r��	�""O�5��E	=�ޡ�� ��y�6,"OhQK�%����G�*��A"O(<0���Д�T�I�N�p�{�"O��{�瓥%� Ba�F���"O�H2�ȊdP #�.�=)^�D	�"O�2b`
YL��! ؒW�"Or w�Фw��I�P�Z�l���"O����ѕ?�|�ޒ"�u��"O�a �"A+Qתm�UHT�
�P`yA"Ob{ǚ�-�f�RF M�.� V"O��@��4b�Rb��}�$��"O�0�Zi͆�r�A�=��G"O��4�l����L~q
�"O�qB��f@�:%�=#X*d��"O���pc��2B��Ʌ�V3#U���Q"O� 
�gO#� ��ᐚR8�U�"Ol�Itg�e���J��/l�U�"O�ei�Âg�<�5莝����"O��9׀�`�,��጖�pw�(��"O�,��l�6IY�I{Em��|�c�"O�X�h[�M����l_� ��A�"O�!��9R�\|�6ҹc�j�z&"O�Y;���CrE��
�"�B"O�$�f�5g� 9xK<jp�)p�"O��*&k��a��U@qj�o~�-�p"OĀB%O�.FP����!z�%x�"OP�XP
�O��QE�\֞�S4"O� Iw��:*}pXk�N�+a:H�@"O*)9���Y����`�Q�l��C�"OTM�R�
����v(U0n�x�h
�'������*�LLq�6Nq�
�'?�E��Q�l� `�*Cz8(!�'C�A�
�!	���0�W�@�fi2
�'o\�+GBU#R1 ���`�	�'*`��EʣLf���GF�t��'a.@�똚�R�B��T79��Uz�'���	�/�*%�%��$578`�'�R�
��9 � ��C1R1�' \y�G��0C���*�T�Y	�'�d���%�Cp��Z�F�+´l��'3<����D)W����V6X��qx�'Vt���b�$2|S�#ҞI.�h�'�pᠴ�ʌ���[whG�P�e��'clh��`	�I�q��?W�z���'�Ԭ�&怫t�@0�ը�?z����'�
�a�S&�5�HO�k�\���' ���7H��uޤ �,�h�(���'����.�Fȱ:�� *h�=��',xA;�ϥ}�j���SR&	�yIS,�HrQ@j�};�k
<�yr�Ċ�d�+h��f��HX��ȅ�y�a�6�2�j����h���tGܼ�yF�N�J��W��]�� ��NZ��y"e��A��툱c���i%�Ü�y29�ر��`^Wx�sSeٛ�y�N�h�f���AI&#����R�S?�yX�;�s��L
���
r�*�y
� �h)c�W�"
�y��Pn$�e�!"OpĢ�B�nc� Wcm ��&"O捩F$K�`��P�mO�0R,�Z�"O�!���V�V�:u��_��x�"O��	�&g8Hx�3.�	e|2� "O���c�<��1�l�-n�F"OVB�a 0&���1Vl�r���"O�/��[��s���df����!D�Ԁ�M.7W0�qbD��oj� �=D���G�.SXY�1A�O�����!=D�p���>_�(��u���w։���/D��K L��2)��-P�D,D��0u`_(#^a�a�KV���rr'D�ܻf�N�`R�QC@�ǒA��y�&D�r'ew֥[�ؑIp�sB�$D� �IYjoJi�����V�@�g>D�l����v�$dQ��B��
�7D���Ҏ��g��ٹ�L�*�@��ŋ D�(�@j�8�1��B)hTF���<D��H�d��d mJ���-#̥B�:D�D[�F,M�L��N^���	�:D��J�W?H.*���o�SY�6�4D� �t�	 mq1C\�)u�4D��c!ξa͆Dy�@ 0�A9Ѡ'D��c�o�x�2���
Q��$�g�:D��p��]l��j֫S"r �H�6D�p����F�X�	c��O[*��4�2D�,Pa���<`�g.�0��|��%D�(��tFΌ�꘬b�T��-D�h�%�ۺV�ɐ�B�Ls�|��	.D�H�n�-|��+%�Q�'f��2P')D��
pȀB���ۓK
 *�����%D�0� ��5yl���e	�8B�a�!D�Ț0+��XP��
v/�(a6~\s�N>D�$Y�O�*Z*��bt$1M�����<D�4�\�#*!⒩���z�"M D� S��t�:���/aO,���3D��u��<�{�,�5
�m�C1D�HY�'�, ���+�̍�.C,�.;D��	G�b�r�bŊ]�
�@�7D�Ġ���L��=�0`ɔ�YZ�!D�@�U��>A>%��-_� =��<D�P�f$P:Z&Jȹv��Z(�Pd�<D� �b�<4�I� �	����g�/D�|���d{HA9��0��0"�I1T��If��yn����ˇ�k7!�4"OhEBs�6F��㇊�-Mh���"O�0i�#�9+/İJ���	Y9*X��"O"��-~��ڢ�߳Z4��w"O�!8W�E!�zq����7�x�%"O�YG#�1wh�2S��1� �"O����
2"������"!Ҁ"O<< qKZ�JT"wV;E�Đc�"O0LhO*6H��2���;\d[�"O�� l�4T��b�CBSG���"O$=��d�YgX�cĉN����yb�>M����sfD��<Yچc� �y��k��}C�A�y�80ƧC��y�ܓg��sՌ�-��0�բ��yr+	���LS�rh�%���y�F�Kl~���膗k
$���ᚶ�yr+T�3��웄�NZ.�Ce!ߍ�y��1!`D0�� \�6��TrQh���y��7f(8�k�� �X��f�]!�y
� 4u��%D�^�$���IY7���"OhYrh�%M�&9��̎���"O"q)Îԁpl3Qf$��k6"Op����/b�0|���&"� 1"O�d`�f��o�*�H6Mܫ9� ""O�9�"b�-z�Ġ-Ʊopv09"Op��.�;a�<����54T�y��"On�s��
}�N�a�ٟG�e0�"O�T�D�،OV`BQ&Øb=����"O�H6�ѣ�M�7eL3}04"O�\9��62kg�Cev�[q"Ob�&#&:��!e�<Z{^��S"O��`�i� �6Ku��k��B#"OfD��E3!$��d!ւa�.t�S"O*K.��;L\`@�C߆�y"O��3caF�gqR<xP@�r����q"OMxT�5_,�M)`	о{�"1�g"O�5� �"N.d`�F�W昐;�"O4�@��~���s�%��9"O��HE�-`!���	k�>�3�'�Pl�p$��:���ч<u�l{�'$�жcR�\ AKW�dI�	�'u�İa���V�H�p�j�}f�*	�'��4KlXazu�ǅj٠|��'䲌`𥗥  �뤈��dq���
�'�ʰ�4��+	 r��dH�c�@@	�'d��sf�| ������_6����'�	��`ۆF�`@��Q%�z���'�Y��b�-,��@fE�4#Α��'ښ	��Ā$����G�&�y��'|��QjH Kz�ɷdB)S�e��'�>��V*HA�������0�=j�'Ҳ"���.(zK7@������'V6ra���豙����U
L��'tv+���}�HE���R�	q����'%�2E@ѧeW�tF�{[^aP	�'�u0���7�U��O�8s��t��'��a���g��avi7q���'�p����4@���z`*	�'�=W% �5��2ix(��!D�: b8p�i��!���a;D���Ƌ_����bI$���)9D�0�C�ߍ#�ڬIe G6d>��[e8D���R�.���G��D�5���5D���NxI�#�,!
�@aa@?D� s��R8T��@�RE(qi�i�C?D��8Q*A"#YhaI��";uxhɷ�)D��Y7���8b�Q3�m�\@>���&D�tKU�!")H�pB���4�g�"D��sv�M�1����5�@�`�٨��5D�ȓvĜ���b��K�l̾)C��2D��s�I�{
^ �,��Z=V�ra�/D��B M�j�zl!��@��hP�2D�������4�F�O��h��*2�O<}�O��S����K���gj��~��̋A�2D�|�5lF�K%���?g F�2D����G�d�8�'቙H� E��O>D�T��'�+u�aX��=@�(Z�#>D��	'kN�e�� �&E�j�d?D�l�Ƣ&\�
���G�Q�XX*��9D�p�̏�/�$Hjbf"k\��M7D�pҕM�.��@#b#���j�0��*D���Bg׷sfN`�p�P�te.��T�(D���Vh�1g���mK�a|ހ�si%D�� `��#Źd�� 	���rM$S�3O����]�Ԍ�ĂW�#�蹱#dS�n>!�$�2�ji����;$�ݳDҡ�v����X�r���efF��@�o,��hO���+���ڂe�m�a8���y�x">��I@�<SܙB@�%����n 1!�ǘRG��r��۽Q�����)!�dЎ
dȜ�whU:Ǻ)����F��O����5b�B���w�ΰ�f�2��7�O��#�)O1�*�R�����}�"O�X
cj��o4���eȯV��	��'��D�t�>Q�4��z����I�tn��*��DRn��yrI�o��q�+�@^�鲤)L	�0=y���W:5fHhAgKٶj�bĬԮ�(Oi�� ڹ�voW���p��hV�vn�%��E{��T!�
B�$z�߄���KU��y�`�!��Ѻ%��ީ9����'?az����T�؉�W!6�^���'J��p>i�>q1B�5��Pj\��i RƎßLΓ�~r�'b?��O�N4+�
�>��f%Yۦq;��ɧ#ĢZ�#��!U�	%��W��{��n�<��!CI�$�����&dS�ٕX!��Ey��)�OvXrf�ɞvW4���E��9��Q2U�@��	p�p1�W��;r���y���Ysh�	�a~2	�G�t1��p�a������>���<��d�Hx��Q.��YGXix��	D}��'�icfg�N�[�,�R�1�'A¸# ��6�p,Yf�J!H���'��M3�ǵ5�d���H�@-v�.ON�=Ys�Ę�.�@w�7��]�QmR73��	a���;��DC��	���/��q�%�7�r�L+5�O�`崽��)!����(6D��y��;=�HHS�+ {b���#�uӈ��m̓e�Q?!���ȍ"L|�ad̚Ίɑ`O>D�(2S&7� sSO?dXEԥ<D�ܸT皣J�fM��K�4%8�$:D�h��Ȇ�n�P�[��	n���o7D�pRb`�Tl��@#�C؅Af5D�,�pFۿ-Z���hHH̚%C5�1D���a�
�/�R �¢�(4d=��;D��pb�W�%���|rdX4�%D�h8��$��
��Q��H�T�#D� Y �"3,�i)�`�' �@g�5�O�II�F��T!r֪}	1��+?"�B��HM&E��Z�[,@�F��0��B��)�L�K"K�*�@� 蕭-E���$�/U���<ad*J!h,�"q(�{��}�؞D!�Q�`jqJ�G�e��I� ƀq'!�P�/R� ��i	*�d��c�!�D��7�VL����a�B��S�HD���D��,T#Ԧm`G�H�\�����!10!����B��E26.���P����9+!�#0�@ԲLG\8��C�ߗp!�$׳xsT��Ś� u\h��b��P!�$��x����C�)6���8���)�OpHP�{�����&�Qwo�1IGh�!BL�:ǒC�Ʉ2X�ar�B�&V<���g�mfC�Iڟ���G�F6er�AE�Z(��
��2D���1�]�/�
[d�C�X��;f`%D��ȡlB+'@�5b��η��d"��"D�4��ߋT%�T�G?V�N�6͟jy��)�'I?���!ʗ�8��T�����K�jчȓ'�
pH7�� ,��@���Z~��� D1A2�]�%<z`#���BD��'2��z�S�π ��[��a��䭟7M�R�"�i���o8�Djs�Ϧsf��Y�'6h1�2�(}�)�ӫU`P�A 2^p���һߖC�	%m.t�f�\��z�#�Q5#%���&������?8|���Av���(lO�Lyb�'oX�%K����!Y0����	�'4Xt	�B������2fp{�'L"�I�`l8��,B>UX�bO&�y2/�W�B�*��F�Ѭ��1c���=��y�X?x�`L��BK&I���!��N��y�L�{
C�	J�"�qAk܌���;��&�'a���0�ǉv���`��Q�;�L�ȓQ���!��6h�L؄�Ѽw��<Fz�g2O^���'�#[��8ũ̻b �%J�በD��Ix����Hȕ@g��P��A9E�p��"O P�G�B�enp`��^0X�QA��'f1O�PL��6�Xc��W$V�bհR"O���Q�D�a�����F����W��;��)�'M��2�C���([�"�M�rl�ēR�J�P���
� a��Y�"�8��>I�`+�OH�wj��p���C�ɋB0H��"Ov�eH���R�P��V����xb�'B�0rA�I�{g�"&48��x{�'�h$�7�
��>U�� �(��p)�'�LEӕ���8LXǈL�I"ы}��)񩇘N����kFƄ�ZAMA�2�!�d�;w��5`#"��`�0E���["=�!�$�O���Eɐ�̚Ē�K�ay��'[qO8��4��%W�A��툐A��ȥ"O��a�FгA�9�r�P-N^��"O��� �ϟ2�����q�.���"O�����,� ���3>B�0:���3�(O�c>�j�&�
�� ��%X8H�����$?�S�S�k�u�s�W@� ��b�tB�	n���bR0Ն�q�C�;�^��d�<a��+W4Aq�JE"(��+�W|!�E:6)r�҇a�'o�PH�-�/o!�c ��x���;��S�?$o��XF�d�K:SR�ܘm��4 P���D/�S�Of�!@֏�y��0�S	�2#�TT	�'�hI1*�7k��p�+p�h�'G`�A�#�3Z1�8��%?����B�)��<�hT9�, "t���Z��&F����'�a}�J4x�4ȗ(��~8
YzBJ�y�� &~�XƦ�eGɹt� :��?A�'����G�Q�m1&�_a��
��'�>E0�iq]��c'#�2;[�����5���2��3�޾4$p
	�T�(Їȓt�<Q�G%O��!1@� �d�dH�ȓ4O,|&��6q�z̐��&*M�)��x�.���.�� 2̤���l�D�������9��m�2J�ݚl��{���*'��L���bko�D�ȓA莌H�郭iR6H*w�g���ȓn��4[�L��,.�`Z���[R���ȓC��@[��ˣU�|˕�A
xt���'4���AC�h�8DB��d��B��a�r'�8lET�qҭ�i��Y��
L�)�B�Y=!A���[T���W���؁Ŏ�D�ũ�FA�u���ȓ]�*�䚔Jæ$z���c�V]�ȓ}c��G���Ň�7)���"O�U�G�(I��!�\x����ʡ�y���*$�����)�g,Ξ�y
� ^l���TPґ�jL�+L���@"O��� D�<:N�TKR��j,ne)�"Oz����5�̨��T�(�T��"O���`�Qܰ�Yu��n�ف&"O2ܺ�O���
V��?R+x3f"Oh�k5σ�:H�|���˖u�v�9G"O�-�f#��5������K��� �"O��ң�k��2�"�f��EJ�"O����G�\�&�BV�N��j�@�"O�a� % ���E�3m��3֔p�"O���Uj4sy�L�k��'��"OJ=� Z���ēd���3j`���"Olt��%�@�iႦʂ h��2""O�P����8 vdR��R�n3h !*O������p#�רc6x�"�':�!��Z%o�VT ��<
�:���'����&�&I��� 3��i��'����B	�{�y���ܒ^~���'۰a0VKD�j�
 ����L���q�'���ZTk7$5|4@Ņ�6TR0��'����$G]��9�U�^�'�>4�'X���cf�\�2Tݞ	����'oL��K]#�D��&C���)�&�2��	j��U<k=9�$�Ш@��=�d��h �92͆ȓUD��F(J1=��u�f��E?�؆�2��|pCV�J��0J�^�V�r��,���杸>ݪŉUD�8XNv��ȓ\���6�ǄBN ��m��r|��ȓe�TY��~Pec�*DZXx��tq� Y1�T�W��b�*�0���\�x�҄O�
z?��z�̉�X6� �ȓ<Xข1��0��7C!.�椆�k�(�I�BF(m	����5���ȓo�T`Icm C7�0��]�5�>d��2d�H���!��`a�JM�M�"���H1�̀���#��I��ވL�d�ȓZ�s(�U�Y���" �P���;%�� 2�U�|0�a����񢕄ȓo��% ֨M��� ��bZ�a���ȓJ[L ��(�$q�(Y3�^�*��m�ȓ0�x�J֣�a����t�>`����Z�>�;b��6�N�bd���p ��ȓYU>)��U�04;T�ҲQQ���9,����|B��.\v:W#\O��e ��\���
��T
�o �db�,�)T=��ȓ�Ni� )�,YP����?^�'�����׎>X��1��f�O�(͈B�v���A���z�0���'LԥA!�Io�t{Q@�1O�6А���v�с��O�q��!�u�g�	�?TU�I�Yf�l� z�B�������\�`7+J	v���`�/c�$��Et�����r�p5�T��:���F��U9b�?��h�9,��h+P�O5nX����|�)�g�2d�<�J��2?��pF�0D��� A�+(*�1����	����f��DYq�Q��&l�w��7z�l�pE���(��4J�h�Q ��ހ@Uzd�u"O&e:��I�&A!qL �%o �"���$u�� ��Q�4r�Q)W�&a2ׯ�&I9�{�C�3�����9(�(��'�0��<����)�$��G�1=�${��@'n,q�h!RhZ|��U�X�"Q�y�"0��Eg��Lj"왑A�3C�T��.�3�*<�@)Q=�I�7*U9HN�)�#�6dl�rE����9KN�=kA�k������J�z܊��Yy�'���&Ko�O8�ч���vu�CM��B���)�a�,��Pk;�MY�n^�g,����J���!r��ϻ"Z䘉��\�HM�F�I�;�%NYʽᐞ>!����u'f#]��V�,^���ŉ.�bB���1K!f=�ℍ
W�䰢��"U�9�t����'��\�� �*���ř0 N�d��4Z����5�0N�(8��.Gb D1�I? ,B��
�S�(�C�5�F�Aʓj�0X%�Q�g3`��<��Oƈ*E�ĨL]�=
� �ǀ ��ys̏5Xu��+5�[c������P)��5��Q`-^�2h����ϖu�PT�����)[wR&<�%K:®����E%K���[%BP�ʓ�$�f/���]�!�t�_��B�'�԰��N� .�T<ZF�V2')�0¨�o�5��jĠdp+�&���S/�����D�߹X1���d#��.,�@J��5��õ#�<L0��I�U�tM�'n9Y2���D�Yy��9~�����wN��X���-#, �Z�o�U��L1wDڎ!3\�Z"��/`�xE(MsE��0bc�/''��'�޴x�g�;x���R�$E<`\��4r���ǭ�%MtTJ�S�����?5� ��iP�Q��33����;D班UQ\�2Ǭ�^����Gr��J��q���еX����s�4X����]Opz�:�lI�}{�t;a�f�����-VԐ	�ƭ<y�f]�2��L�6g�h_�c�����Y,SҘ�O��<5#�i��k�GW�/O����΁T;\ ��a�'yv�D���Xݴ�>��JK��ͼ� �մ㨰����?��8Ѣ�I�	}He�A.��)�S�M�*ւ�� ���矙$R���A�*kǒPاE�Hh����M[��R���l�~]^`��FJ�Kٲ�K���
��t�EĔMa����]��ល7l8	��&ݕHD�ܙ�̂ �#�#(g�}�N:�<� ���3f.=�"��OK���Ӭ�"�3&R�>Y�`AM�
|Ҝ��b޹Rxc�#�����`̻*���'_:` ���5�~�����T�0 �RA��{�'�*GԌQ7 ��dE9Vx�����sj}�ǠA�RC��#gY	/MĨ�@֖{ t ���&�r&O�"�&)�6H�m��	�@�Q�m�	ݒ��C�%P���X��$�˧s��T{��T3���(�l�0b��@��1sZ�qc�މ��%6k�w��HK����|:��_1f�����aB�B�P8�����) �(��0i]�'.8�ß�"���:�H"�S�}�Fi4AFH��9"�ě#1֐0���уI�`%��B��bN�-B��H����1]#�zFdڠ7ۆ�7�x��t?D��Ò�p���I�z2��i���:=$U*���B����M+`�N�|Q�R+2�v�sF+p��RA��FD������!Q�P��GY.�(d;Ԅ�*Y�8b�`+��X�X�>��'}��W�;rEP�C$L�'161
m�	x����:E�,lj�C��uڬ�����tHF��� <,R�mJ�z�� �;4Lqa'�ǝO8���I�EܓI�����"��<z2��g�>C�@�<�&)F � !�@����s/�a�:B͇�J�l@!>�*i�0��Y���ہ%Ev 
��P��̩��'r���7ǎl@t�B�"͡5E�e�#��6GJ�)����/�4�D�>o�D3Ԥ0oGz�P��"3N���8�P�h��p�C��<y���F�2�B ]��
�;L,��G�]h�6�P��46�4��6g$N����>V��`[jR)i�h�t��K�������mv���DA�sV2L�2A��D�O�my�eB�(� � ��h{���A�p^ d��-@����FD"�U��J��tF�����Y�BB�	�vT ��ω3�|� �q$��G�+������9� ��M;�D4l��A5"�l�;XȬ�P�I��e��4!e��?�i���
qܺ��mG�;L�a勇Wo�����g��Z�#D [�D 5�/��AHo"0X(�K�Sf���J<i'+/"�Ic�H�}u�(�����'�b���d�o�Y""Ofd=�.׊Z� ���@ՙv̡Aaˌ�d�.��Ы*N��@���p`��2,O�3��u!��˦"�����Oa���U�GȬD��	W��8֭O��@�T�
�(��� E�g�����XT�(�܇R����R
�*�E}�e�c|�u8����^�(���Z�,i��_���+E"շ,$����4��=*1. 8V(RE��B��3�^#��%"��'<��XJk�����#4.��S`�"�t�|Cv��6�E|	꼻�˻".*��'D��~>��`˺'%:ĺ�&RVÆ�㡌��8�x�dm��j$�!��	>�(��!�%KѦ�� &��Tƈȳ,�.�ēp�ݻ'N�V��,��S6�!�-�<y�2�JU
��>�4	A���p�͋WN+R�� �㋓�0�%i'͑�$�����R�V�f��c�˓�KMZsf���鞩O����E�
�(O����/ǑYth0�2�
�3h�c���M+X{%P�/�����1&nԍۤ �4P1��H5f��'���h@�@T��s�FFQ@d�5��%6�ƐB��N�'�����GBYPD����'2�֌r���>�4�� ��y0p���6�8���'R�] 8\�w�Bk�m;a���Hp4��Š�z>d�K���2���G�+\����H»w:����LM�:��ӂ�i8YP�Nv��y��tP䰫��Іr�` q7��q�(���8|=A�T���S�9+��1��A�Ms(tHq@X�5�b���2*�L�dG� ��{co�x�I�"�꽋��X�=V�0K���G��q��_9��	�#��UZ��	d�M�&�����)ز?_�5��@�����.{����j�"vQ�U���r����Z�����\�J"=)g�΋T��a�So���t #��R���;���F���	ǳT�P*\�Ul(�@�Ę�r0oZ��F����A�DL�(SC��t ��Y��O �9"B5'`4#=��;Y��1$�
 ��(s�!4��{�U1 �x�rl	?+{,��F�X��B=C2L�( ����炩i
�}kphT3%�p�2�,�=-p8��& �6��$̏�.�Fm1·�3}�1q�3:y��%�)n*��x��� C81��NUС���]4o�8[bd�<)W��Pg��Ӵ)�3'ln8�N�_��x�L�!3b��E���OЈO��Zv�MK����k�����ʨc,� i�ߝ_3�A���>"���"�b̐O�����Xm���[��
)c(���gl�f�f�PF�W�L>8!���y�X�y��'�lX2���GLW�&6&x���*������PpjaybCB.v|��iʛg5�qg� 4&|m�yX<EIc��O���r���5�D��zŉ�ӅO�D0@��DQ�7�J����[..�D�3�F�
K�q���pc���+
�'�|�t �HT\ȡ�8��l��bL�O�$����dكkK�!�p�OI��zp���v	h��٬>�d3�'f����Wی����L5v��Z F��zH��-=�Lc�.�.b8�q��1?i�M��+݋|�Zl[Q�S�F*�&ܥm���ꄴ�0�y��ɗ���"����H�3�ӈ*��MI ɚ)�����$:54��,ߕ���B�
���\�c�
-��a����.��Y�I����� �'|/�i�@* ?�a{��Ż,@]�tC�I�&���dU�Y�0�� ��M>�}�4�ӹ[IX��eHS�p<���c�N��fK)�SdZ��� ���gD'37�Д�	�h:H�������X��}$b� h ��A����+�AA�,���c�F�5�|�2 �ő0wϺ�6HK�;2���7�C_{��k>�ئ� ����� �n��<��$�\@�R�Q� ���O�^�I�'��d�:.�
4v�X9�!3��Yq*D�a�ҭXS'L�cdm(��X��F,FN�?])��J�HeP=�� �	d��"��
6����D�>�c%f��L���Q�P邙#|�f�ŚIU�P
#Os=�IZ<xL�q���
���ć
�2��ѫ�
�zRn��Y���V(��	�l��t)!a�kJ	��E�� {�t�΍�Aˆ���R"+�'I�o��h��Ӧ(����N�<:�h�qNK���x�i
0�U��ޓe�ް �ߌKX8��I6p?�	!֭�����d�ýX˄H��^g�ʜh�I�NP6��5L�6r�"�
�*��f��*��1N�Q��Xpb�e�)K�	�� N��8r]%��ik��!\���!N�Bq��j�5 ? )�EGɲ*=�d(U��yC���#Yu�'�V���B�8K9�l
e�S�/����H�X�T
@�Wb5K'�]qx@�B�)ƔN�
t��%�uҁ���1ᤘh6�6B��Trs�A4C��"�.�c��Ms�
̤5D����&_�Lpf��%4��E@اG�t1RE�Bj�5�㏫^�QT�A�#R�x(�f�� ?�� ��F�@I�e3k�:U�Q���b�vɻD�3�E�'�M����P4�}�tƍC�lܫrnѫR�Dk��7Jb��0���=)����%6P0�Y����F�z���NЩ�E��*!� �3���!jĹ�bő�p�
̇�	�=1 � �n\�-�~��� _�Gԉ�A
� OnA�� YxT���Z�-rD�i��ٱ�F�O3����ꑡJ`a�v�^�	YiT�ʒbB 4�	jw���.��k (Stn[�P�eÀ+�UTLxh ���C���@E�7�ƌ:0A4^�Q�G�o3�Qwg��!!C�ܗ{��U�V�߅��<a@%\;s���Ϊd������ Y؁k� ͌_b�����	8H6�"�E�u���uFO�`�����R�Qʽt�C�*�(����[�Z�88�r�ϯ��?DÈ#w>���gMYB���)�-c�TIR�B}֬�e���:�"�M�#v:�0�\K��HQ�/f�DQz⧂7 &	K�LY�v�X�`mݨ/����	�g�8�{Tb�1m�RYIDl���Mx3��qutY	�*�ZDZM��z�$g�D�*����H4�i8C&�spzyY�"�9~"iA� S�&\���a�R�G��'O�Py�ߧF��sW�%) 
@jW�
�p1�Ej$�	9u)�`� ��I��� D�� ����/�1("U�t�Y�Bqb�2l=\O�{���+^D�	��!f�\��^;4M̉���#��="j"q��3D /TR�aB��#c�^2����c�Թ&^@!���R&.5�!��~�'���!U��W�O��yKc&�&���"vf�[��
�(�52k�1qB�	�eg]��,�!P�zas���$����f�_��,ReHW�6c��)��Q�-M����[K�@R�dIR�y��$j�ҧ��P$j����$�%Q@��yu��+n@ʈs�.[,`p�H@J
�N����V��s���`�W���\VHEk�&9�(O�5k���9O�: piJ�B^`m�:OΕ�D� �� 9�e&?��;Fb��K�($p�I�GTrq�S�ݲb&����08DH��x����X����V���G��L�q�7�C�����g�-R��U3p�� Wٺ�A�)ΟG�P��$�@�?J�
�"���)��KyܫáA�Uܴ�"��A�D��t��?>r��6fg��l"<Zne��( ��'T��Ki��83AX`�dg�����BFnI�t�j�$�al���P�պb�μ��.ǩuK��b&�����;`�ޔ�dΆ�sA��λ 6���FR=�¥!����c�e*0C�j0��g��Z6�o�����?�@�"߳:�,1�aG^N��ts�CS11���07�ܐVF�DJ4r2"-cCkȎp[�!�dK��XW�34���$����L��P��d$	�#���!��8|�T e`݃NJ�pRA��F��wL�V��$��!���d9~�@m24	�3���i�tXL�rf�N�Fφ�rY`��i�;.�|�P�� �W��mۣ��1"mz�s�Q8l�=W����0BUҠI���E������9ch03t���u
�mH�,N9]�%�&G�B&Q3��̘��8
�bY�4��UzCB0�� 5��u*��Ѷu�ܬa��
#1-�ps�$5 Y;��wm:A3Q��'= *�/7$z8�)w��6F�}ړa���\t[�grd.U;$�%9<����yw ��{/<EU��f�(�����(�H�Gb�VaR��=.t��� �$x)4I�O��a�F o8ɛܒ��P��B'){h���f�?N���IQ�ը�?��&�Hb<ͻ�n��D����P�yo�'�H�14MP�uO�9��nW�}V�4B&�ŜG�qS'䚱N�d��7�	�g�@�4-4sF���NW�z[�<Jh��G��%g$�_����
6v6X�uʝvJ����K	=0�|KW�!�		<4�`�� 'Y��H�fՔB��r�  �0�2�
F�_kPY��\.sdSC���g*��զ�@��z����2�*�J��ÌZa@E1t��7Nd�8ӵA޷g�N�����I��D@��A%��Qb��/�!;Պ�c�`b0oۧX�F5�ȲP^l��I%�p�����m�� Sq�$E2�|RM�8\�P��PB����"�O(,����9�R�\9O������'%P,t��k3+!��=}�uJR%B%��Ò�]�L��'>�ϻLr�q��Z_�^&>&�H�)�=�.� Ȓ/-�4}�"ދq�Fd�S���>����S��ēM���M�H�L �W�N�,9q��a��y ���ʄ�yq�lۢ���|���M-J�F0�7�N6-;e� ��61N�Y���1M�Xl�օ��b0^1(�ㅚ�T=����4o[�D;��D��i�f�z`fG�5�6Hj�C
Hl�X���|��q)gå2v��q d��gZ�(��Ä'3_�3qkO�PǶ�ǁR�L����3��4R�;�Z�h��pÌ��[�_����46Z���۹m��P��K�x�؁oD�����L ?��X*�<�W�71��b")�z���/k�O>��J*�h���I>M��y�{�D����{p)Q,XE�ԧ�1^�D�ڣj�ZN�[1g��j~.�%*�+<��eo��y)� �f��|b�սy����E�Z�93�)�Vţ���X�^h��'�AE��O�0�O�6+�b8ʵ�W-X�,�b�B�`h�B�]�|ц� 憊'I(��'F�k�:7�И��D�t�>������J
!'a^�`����]!��=�`IF?*��s�~�  c`�\̈��e�"u����T"O�  �X�dG%PѤ�@�oK�fq�PkD�I5F&�P���(:JU� �*m��� ��ˉl�.B�ɚ*v�0l��&�u��KU��tB䉈?ph�p����Y~N}����7'�`B��.524����+&��+�*�	!
�C�əI#n�"CE�$���P�L�C�	�,/� �,�2*�,r�l��:<FB�I.��Ũ�M��Q�����K�yBB�I�M$Ԥ�G��26�Q3�ˈx �B�	x ٣M� ���U��L'*B�,��h�l�
�0A��H>Y�B��%#ê�YG���Kn�K"S
�C�.l�ؓ�A�ђ<r׫�7[�C��2��)��!r@�[1��n �C�I��2 ��Kn쐒�'łB�	��y��LW�:�L�D�ȟ-7�C�	�Cr�!bw�l�$hb�H� mSbC�I5/����	g)�hH#�$�.B��8<�(�,��:Z��i���q�B䉌j�n�3�Z�n"�1��P\��C�?��ĹU�Q�g�h�� �Ca�C��X���ª��c�^I��L��C�	�ḫ�PN̂	uDBQ�Q�"�C�<
��y���*2��3/�B�	o*%��eͿv��xak�/qRC�	�d�PHy�M���#+��B�	�p�!�B�W��KeG�<��C䉽����!"�;Zz<��̂�i�tC䉻	Q�1�7M	((} �5A�2xۼC���ЗCP�n�:��r� 'b�B䉜"��a��*@Etbu��c�xB䉧!Fu���	*![��ѱ��>�DB�I�:���0"��a1��I®�!
.B�	"n(x��Y+��#D��zd�B�	8���r�ߢ�|�x$üe�C䉜`q�̀�a9�.��4%�2BC�I�7����"A"NJ�[7�
&(�B�	�iG4y�t�0,�^�Ҩ�,��B�I4V�=�Q�
�ewʀQjĥ_�TC�ɲ*��cT
��K��b�C�� �B�l7~+&@��xln�[֯ndB�I7qF�,ɳڌ
��"g��K�C�I�<j��d��<Hį-5l�C�ɺ`Z�K�G���5���	 '
�C䉣a���	�n���#�mNB�I�sA(�vΙ!;G��5@V*^��C�ɦV���XC�Ҕf�N5ӆ"�(ƸC�I dXz ,_ �\=���F&Jΰ��$C(Vͺx����>Aa�[̸豒 	$#j��1IUO�<YDH�(� �A�G�#��)���8�O)��/A�C| 2�a4��Е�bG�L�@���������ȓ 4.�A�L�!G�rm�R��r���#C��6�z�'�ܙ�4�>�3��H�X�c`�B(AN�]�vm�<���d�$z�,P0�cL&J�x ᨏ�[D����l��P>�x�DO��������?��H,�?z���jCnD�x�B	�7a�l���ǩ	&�yſi#̘Bģ�)@DWG%}�T$��'��\�W����ř�A��"�p�Or��cc��sO�%���h�ˏ�i�	O������� L48��c�K!�d�V�LE"r+>#b1����w%.) ɕ�&���0֣k�,i �bS V�HM*b;�1O����c��E�B]��ˆ�xxF�'�FU��F6zl�^tXs!P����Q� ÞDyFn��0Q��]^5�'�t1�%.�2C����e���RE�L<Y���j"f��)�&��Is�US�2��Bרl���r��P�!�@���e�	��RR�X]�Q�p�e��3!�?�
j�I��xs�ՆWd��aM�,S�|@�$
	�12TM ��]3�p�Z��GĦ�'Wf���f�� \�S)Ct4�[��r���k��Ŏ:�4Ygc�p�$#���]�7W"\iSk�8bx�5"�fU�m\X(���7�V�;��أBk\m���D�4P2|)�kT9a|��c1i� v��-�Jmqp��Ea�$��S3�JY��.}H'd	���GZXyv�QP̅%>/�D��ؘ{��<�&�&-�L��&m�����h�n��m�>�ț�s���ZP	.���0Q��U`��Uh�:^��u8�l0?9#P��ܺ�)���0��c�Ѱq�R�� �١$����e^L4��H&�@�:��C�w��K��Sy��:w�U;0oXId ����w��-ʂ\�z~���n��l��u����)P�������M���FJ_I��=Ң%�~ZힷQ��T��^= ��A8a��92fe1y��uCQ�U��3v�X��?�7@�_?�%Ɂ�`��=2.Oz�0���)"�Q��A��{�	!�� *{t�j�X�F���g���x���G+$��e�Q!D�{y��+ )||�D��v~�r�҈][� j��f7FB7��)R�2��%%�!T��˓Z�B��$B�*�F�26'��M`	�%C�^���L}�"�Z�mR���Q*䏕o������-f�(y�!�$C�Z7�C?�lm�eL�'	18u�d��@�b�������1�'R�p�Q"XE @L:���&��ϧ!�M��E���)��ݲ|ـe�G���cG��� ���KQ-
�\��y�Z<uw�(��ݾכ�aK�|����I��]B�xh�H�.[�@�c�0+���I ��R��I�o4-�B�;�3?�c��b$��0A��rr�T47�N=� ҟB6��N)$�NU[�K�j6�A����E��R*O4��D�C˾�9 �NW�Qb��҃7PL�al�����Y5I0�DJ��	���'0�>8ce�Dƴ��aŋ>]z��V�"�-��S����be+��`��k�>h��ɕx8��:���8�qc!���|���6���P��4X��UC�>?a�*m��m�VNH?
�.�x�F3ޙ��o���@h�s����V.�Jr ��"����;�O� 4�E5	.�߈�f�w��u}����Բhf}#��G~�WG߃O�R#0��7 +v0�t�2ovUC02�`���.I�h�T �ՅGmv�I�=�(��O,4r��̫����D�<���Â8b���UD/i��A�=?+��c�F��YN0��&��8'��"[�o�Ԉ��xRg��m�|��w%P�7�^�,K�@��7 �7H;DٓR�]�۸'��]d�L/R6�0���CЁ��>&�	�I�{˔l�D
�h.ȨP!�S�vÆ4�l�K���<�7,�H���Ƣ�>)����r}�1�V�B~2��G��hy�mF�X فt��U��\"f`�5Y�v�����J`��yE
̧f`Y��o۠^T�oY�1a����,\��4�ç1/2Q�3o�%AҰu��lٲ+�yI3��?�nmj��Z5̌��Ж7%"M�/���}��̙�(�Yͻ[�
�xf�̠Q���H���C4�����f]�c�� �<����[4��Rq�B�A8.�mp2i�	^�r���	�dp(f�^"�h�����)f���r�D�����өE-Q��z�i��*/Xj�ə�*�:bF*`�ܙ	�@�6H��It��**�bh���\�T`D�7�۝@�Ҥ�B�'��ћt�Dj�x��)b3�z�'�Ԁ�1�Ǎ2�Z�b��ڢr����̻Ld�8��E+g:�JG�޽H�NdB�1T�"D!@h�$�O��Òm�#��<pW��:r��=(�&�`�΁pJ�<���G	(C��oB�a�nH�$,�p�i�5��Q7,)p`YU�^=Fu��)�O>H�𤐂��ɀ�

�mtn��҂�,n�8�YÝ+�����G�(#䪖jә!;���"
�ns`أr�n�ɜ;D=���@_sf$ �R�|�#>���G�C��(�3�O� �J@J���?�b�J��֮ND��q��\�ց� ��P|Ŋ��	1A���U�]	
cay�Ϛ�!�a�|�Z9��Ƙ�y�!X�r�,��T�	�n�v�[��BG��y�@� ��f��ը!A
r��x#��Y�t��@)�)³_P�>)w�7#��=Z����S� <�A�
s�P�r ����A�vn͏^�nD�D�խ����]�j������ƕM�L����:��U��NL[�xl��+u�+M�?��`��RrZT!����� �V��˒j�놝���_ Zr�he9������X+l0�,��GX/b�|��h�$�����-�2K}��bv��<I���2�ɈKր�d��`�l�D��\�I�p �bt1:+]y3"���arP��,D$�	��B�7%<�#!��s(�Z���3? Qq3BS���E�'�3/�$!*$��kl�`{�D�Fs��b��FK<��vFO�s�F8`��D�Gw��MR��X�O@��(4��dmd`aO
�'��h �(ЌB�n$qֆF7���0"�IF��ȱ18���G�N˂j�=+�zӑm�W: ���K�'9���l�?/�j(�m�S2�#���:�|퐕!J�lm�K��F+��BV���[���f3R|��i�"K.e|��U�J8oj�c�ڙD.��j�Z� �q$J)n��
!Sْ�n_0�M�Q�
�m��Z�Lқ42��[��
�O������+�8�9�c?cg�4�A�@GТ"��a�%:��V=Ga�AD�ʠpu�@�Y�X����L?��M!dn�! ��'�l��ϓ��tJ�˻/�N �FK�~�*��@��$2\����LE m�L�wϒ8�ljJ9*�\�֡
�<�ЮY>��e�H��)8��ɑ��� `�[ӊ<�D�=�c� �P�	�s�����!�&	�0E
#M�䝈��~�u��J�$7�^��d/_�+���A��e�曫���s�#�?�,P��;3�ޘ���-�d�;�A$�!�h��n�`b��8$WP?�5���[�H�� C=t�:Y�S�߈a�h�$ ��6X�3���%8B���AT��`Å<p�.u��Ğ�e�b�	�O7��{��X�U�8�H�Cٸ��٘�i�|s3*�%js�׿��Cw�V32���F���-�-Otyc@��]��agEv"�aq.��4���v&x�����BaC@1�9�h��P!5�t��癷@x�� �N�c�=*��>@{�MCD�N
4�6�Q 5�`�S$g�5Gv��P�N��H��Ź��4� Ŝ���9@�a��zUZ����9H+	3@B y+%�ڭH���Ã�;�v�A��RC���I
70���m��GM;%�z�,MqFƖ9~Ҹ ��
6�����' �GD�q���,w�ўX�A�40`�Y ��n��1B�$<�,#�Gu¤�R`�XMP1�!�!f�|Pa�[���y�����I�wĴ��k�H˂H�m>U�v�@;s�v��[H!��(J<L[T��9q?t��e��i�����4a Ё3�Ǟ_N1��(>IQ@|{6 ]�"����A��[L(`GJ�S�.���O(���%�|��p�B�#��#>� �)A�yvJ��"BT�`�2ԓ�2m���''
*#D�8�B?\z1Æ)��zrN��b�
b�"�ӵ��O����f�u��G��3^i
��^kmN�Aۓ ���s#m��]��$���U*�5�H�Vڬ0�0�O*I�H�c�a��[!�(y��ʳ	T���ܴ|��'�"\�s,�n�HM���H!��	hfڡ��O��2M� �pkG �i��V�[4LjNx��Q_��3��#��A�ܴO]�!��T�#��"��I۴��'.���u�
� }�)Bz>�jaD�8�\fA�?G21�#8���{�pJT�ưҘO|�tRtG2V%ܜ`D%��P�e����$L�FI:!�B3DRRl�1���	,.A�d
T$1*<SE�?a���d�b.�[�O'�����g�M�ҥ16�>)����ݘf:��F&���m�"6�"�s̀-
���Y���0r1�l�p��Dj*ղ��ڜ'o�GC�zb(	����d�PH4ˑ)�8M�ŠpJ��ҵ�O* ���ФA�&A�dT@�g]&y��b�)�N�q��Ƅ_)D�BDɞ:~��}j�
M -�ēQ��ي��G5{Bޭ��ѣB<�+6��{lz\���]�=�j$�N0dH�����5xG΅�3� G6�Ę,zh(��W� ���I*��{��'�2H�X�A��,��p��)���ã�Ⱦb$�9��0x�IJ�H98R�ػ���v�~!Ч�%���Ӄe�?j6�iO>�f ��^=ll�d�L�T^2�"7
Q`��Z���Dh�n�D��� F�(���顪�Q�T	R䭁���2D�4����X9p��c�@�@�>i�l�v���'Yz%�p���l���.B�r|��3�֐�����+�6(��9Qn	��	^�|7�\�2���'�.&rp�1��=t6��フ[�hx 'e'�Ot|�Qg�2(*��w���TT��SX�K� �b�+{!��` �*9���
��3++�����P@���K�M�����1.@�Q�c��R��2
�')�ax"�ͫ�`�0@b�W�*i��k���*�pfd
q ��!Q�5I< s�bN:�x��/�
��p�>�H6R�r(�<�|�"_�+Dܐ�㨜%Œ�s��X:�����M�A7F�2s�N�+�ɘUw�����ph*=7C^��*��V����4��]A�`&l[�$E�:�LZhq�%�;<O4!��ꑫ^
%�F#�DQ����R�n���@��h9��!%]?H�$	�vJ�(T��#ۛB\���ĬSj��Be$��vU�80� ]%9O�*6�:�O�jdKF��{����V�T`�t@�6'cuɤ��w�LI�ŖN@Ts�fPJJ��g̀�R�@L�� �4#ee���(4X�q��ֱe��%r��y�axҪ�"��	#wo)2��k�-�w�]Cb74y��`UNH�Yk�A��' �|SSg�P�H�%F��~~�A{w�mX�И' "�c�_%l�~ɋ�JI't�	N��W�U;"�^Ȑ���ap\����-}�D�SB��8�hz�G�2��%�R	$���c���p����/�zU�񈉯�p=�7��uNd��SM�|%t0
�)�"{4$<j��*9B�t��BF!&��$�����pDv��y.` ����y2k��zݤ���B�,}x�����v�ўp+$�޷)�>������"�Ѕ/��)���D[�g���ӻI"n��,ʀ��-�Ve�ywv����?K¶<P�ߑh]�e�WG�|��5a�FK�:2AU�ޫm?pq��H��'i���3}�����C�P�⡚fC��y���Z1�ܶf�r�i \#oN8���G)�U#��t�)�f�R(�j�2�!�c�Q��e��/����V�1,����)��<	�eR��`p��J�[���(����VV29a�G�'"�����
t��C��H,v̳���?DE���M�=��TbF������	��Uء�NE��``�P�KC�U�QW	 \P��e� � u�d�^d�h�ĝZl�LYMHK�yȁ��%T^��U�� �e��%w|zD�D��?C����.���̉$�O����	ҿ?0��Ճ=�Tm�#	k�4�;A9�B	�s(Ն>7ޕ�ƨ�>:<��ӈT�;�JY��c�m���3�r�H�ӽiuڤ��(��(�1	��A�.��'͊�M�4;�jh�OoT�9�K��fy����G[�J:����f� ������4z���d�)d�-!�(4&d#ڞO1�ͩ&��'R��S��=�hP���5��{e��8��������j��>dZ����-M=�n 0(M# <��Kv�_�=��b��K�gH*q��/�@�V�#��ϫc���;��{�ޑ����}�X "g�^"btN��=ak,M+�F��;�>��4O�?�D�3vF7%c̸�̂;H���s�E<bj(yK2��>�,���X!;�F�+��vypB �0i�[���$�֜ˌy2��0'�¬��+�>"�����1G s���8M�*��)3L�u���:��`���]�ְjs���n�h���m5�j4�O�+6I�a�v�>��x��gޑ+�D_�Q9�:s�|��E81@�Q����&�.�+OǮi*F�k�ߒR�ӹx=rE#�b�'�h b�딚M;̬��(�U��8EgǡP�F�ᤣ�Oޕu��	Uy`4Z5��H1ތ����y��Zg�����?l.�l�h�یP����Z�ɳfB�l�z���-Xc��a%��k$�d��V�َX��A�P���R�F 8������0���E�=+�t0�)�j^t��yihYd�Iî
<X���d�/Y"�L��=-@��+c���!L��ʵ�:|ɨ��˘<1���3���,^ ���wl���C��	�%K��;�BC�~������D1C�pW��X�X>��k7BB7}������5^˒-�5#�:q.2�)#���l㖕2É/lU2Ȣ M�0�\��0�>Њ�eB��X�I��̶h圙2�ɂ/mT0̲0�����wD�I��*ע��ga@pCJ�y�`L&�6�j!͚�{�p�DE��%>	̻<U,�p���� d�; ��܃ÅS(N�e��Q)D�K�N�<T(�@��~��P�xAN0�����yi���"GP��ÀGIQ����i�& b4%J�|zuL ��Jĉ�.��FR���`�ș2���*k|	��C�$xp��h�/�_��i�2Ɩ�x:L@���d	I��x���߸��dyAȄ��d!vc�D���!���^�ypHΔf?
�X�Z��p���@u�(��G#T��ĸ���
WF����ДUEB|�HZ�M�%z����,qh�T)��G�m{"a[Ր&�Av�2`�u[� ���T)��<I��n�8�%Ėj��	Z�LXd�O��X�'�I��@�"aю0 p-h�{�G��Hg�>�nDF���7Lϖ ����ap�%��!Co��A�0�MKLN8%�4�>�O�d���4&q��äUk�Y��'l6\SB��<M��Z��(���G�? ���)�n��3$�(Uf��g%9q�0%yq�ֺ?B���$غx{�qBR�hOb�eR:D0�/9LM@!HSm��#��z�aD=<$����kJ�AXT���&�>��=���m���Ad�|-(q,B��yc��Q/y#~�1"O؍C�(״aA(-�Q�Ɓ`d�c�	�:t܅K��z��r-Ҍ8*�|#�B�=`�C�ɟQ��I��X&��凒<X��C�If���S��W*���uÑ7}�C䉩x��a�)͛;��x;�g	
�C�D��0a�]@zd�`�D8&��B�4!k��y�*�--��#A��U��B�ɊQ�TP7��+-���E.��wN�C�I<k;�����V8L�@A��	3�6B�V��;ei�.ņ��$���=�C�	U������J�d��|T���'|�B�I
���3�)S�}ٸ����(o�LB��5ZF��q�M#}�TP��"�<F��B��2�f�_'|��P'/ֲV��B�ɰM�n�#�/SK���O�1K�jB�	&[�Z��u�٥.o�h:�Jؐ
όB�I�8�e1�OO@I���򮝹j?�B�]o�2�d���5�T#A�~B䉆J8�1�\�H�p�Z��
C�I�F� �b��1�R��GB�^^XC�I
kT"����ór�b�K����C�I�.���b���-�xX�G§\��B�ɾz���cab��^�EJs�W`pRB�ɒ0�t��S0����#0�VB�ɢ]D��w�	K�!�HN�`B���ܤ����FiР+� FhB�I�}J�# j�ؼ���#.�^��W����Ha�gb�>���ŚzD� 'U�(Q@D*˧[MR�r���8�tZ-Ol1A1��0|�R�!�@DZFBJ�%B�! ��R(M��I�)��!��&K�Q?��K�Y]�jɄ�0��!��n�T���H'��q�,�l�)�'F��ak6��"s'4�)E �:�6ec�	]6fRh):gb3���:�~2��߈R~���THg]���˗�SY�'ϸH��s���h�e���h�K��y-�EO6�$��Nľ�b>��!N�X�$QJ��u\���7}�ȵH����y��^�JZ��s@%�!z�ȩ�Ҡ��<i���ȓ!Tf�j�VF	������d��g_���d��2�-"�M�e4�݇�J^�a"hL�bU�C�[^�(�ȓ=�8q�e��i��i�7/��;��U��`XP��cNƏ&}�-� �Z5(
�Ԇȓ設S ���.4a�-E����ȓ5�F��+�:��q&�Χ?�\�ȓD톄0�G�p�sF)F!q"����1��Ɉ�ɘ�Y�лi�8�x��E��ˢ-N;P/p)�e��=^6��ȓyN���D"�2:�dA���=x�h���g�L��ՅN'��5���*�1�ȓrXz� �A�J-@i`�*_�,`��_�");���Nئ\����:�8X�ȓI��:R�F�P<�䋑��#k��ąȓ^6%	M�?a�%��A��)��cd����ۃQ�@X���Y9�2��ȓn��K%���
����(*x�ȓY.\��$R�%y��ʀ���xPb��
ޝ
��}kj�
}�I��{�M��K�JL�R����Z���v�%��.�81B4��J̤oY�D�ȓg;z��� 7f&�J�I���Ї�s�����L�s�����W��݄�Ll`;E	�-�����Wb�U��S�? 6��f�5W�Z�{� Z+4(4ؙ "ODq����24�-t�W�K���H�"O�(��_�&��X0�´`����q"Op�K����P����a�����"O��(���k�8`�� h����@"O����2��q�f�ȝ)����"O2�K�G�D�9���έJs<P""O�|R#�ܬO�F-�.8e\m�3"O"���$��B��4���"O�� W�m�6 pn
�TЂ�"OP�2��>0�|�d _o}2Uɐ"O
zDХBi�� ő�4c��"O-#2�'e�Z8���	�yct��"O�q��AW�cU�� �o@PKV�С"OҠ3h��'�`���$]�d/܀��"O��J���&�h�s䂌x�X#3"O@�u�� [@I����>��U��"O�suoL���$�橗g��yU"O�s7aA�Z'R�A4K��3���p"O4]�.�/w�+I��7n�10�"OR�3F��1&IP�b��@�[WY�w"O��Q���0W�qpG�^"!���b�"OT�q�@ԙf�0�kkZ��"O,+P�ڝS 
��4-%&6]Q"O\�2�Q5H�P�Q"x0�"O�԰��G�R#.��fL�_ܪ��"O��B@-K�/���q��'3��9"O�A��J7O>.�Z��J=��u+V"O }0⥙2<cd<���Wm�diu"O%�fZ�K5P�t�̍b�����"O$�@�B0[R4�q��/h�>��"O��BU�дkY�@�E�ٙ8Ҹ$!�"O.���dՒIj��a
�D"O��vF��.�1�c%tq�$:0"ONĲ�	�L"���b�1J7�h�"O��ۑB)�ژr�a�( ,`�"O = ��D�!9p��d���8R͐R"O�y
 n�2&�{��X�f�qAS"Or(�$ѪY��`1A"��z!�M��"O��X�ț�M�\�$�
/lh"O4�s!I+	:��!�AH�0��{�"O�$(��_ >��݊�S'�X�r%"ONY�d�&c���k��oF�2�"O�8��)�1t�\x�5%H�M^�W"O�ք(��rǦT�`!0k%"Ov�S%�p�M���4#h��"O$���^�)���P�A��"O}{��m�z���ؾv�P5	7"O
���E9j���&�) n�p"O �s�Qd�f��P$D	�	!"O�]Sv�9�������-Ԑ�Y�"OD���VM V��q�C4�n�I4"O-0DIF�n�����=,���{�"O"����0	0v'<@�Hr"O4{e���t��=bW���@��j�"On0�PLθ!٤�X�'�/zr�+"OP�@�ؠ"f��TH�Z��"O�p8#�ٛ3�  ��o"�`I2B"O�9��vC&�{��E
#��ٚ "O�Lq����M��`���9|�[�"O�Z��?Jx���O�����`�h�{��N#G�����E��
�H��my����1z������$%�Ć�|�*�p�	��,t��f�]q" ��S�? ���<}&59���1�xHi�"Oz!��ܤK�v���m�?�B$�V"OXu��b���b�+R�U_�q1d"O��Xb)סr��pza��
vE\@��"O,� (T>u$t�A�bI��9"O(�� H�m�P=0�A�946d3�"O6y۳�G�}�@����v(�D��"O���@�d���Kb��#��"O�d�����<P�pvK�D��2"Oh�h��\:/���W�?�}��"Ot����:7t����B /ٸ��"O�ݪ!������*� k@͙@"OH�YR�:"_��5ώ�G
�4#"O:�#@�=�H��0�C)g�eXG"O�@��*m�]c��(��H�"O�d@��������dB������"O�����8�xH�'�E�JK���"O�!"�m�4LS�4�wl��"G�4Kb"O謁s&H�?]"���76J��T"O����Q)Y�Rhk���G2���F"OT�˧,ӴX�� #�X q0��K&"O\X�*�A%�X9��!l�y2"OZi�j�!&���kЄP�^�t&"O�I��N��d�S$Ӽk���"O���A�?_�2H#��ػ�*�2�"OD�3�I���Y���-_pr<��"O"и��éQv�E�E�Ik$a1"OphY�G_�w�J�+��� Xr��h�"O��k2�8��laS�""^�aI"O�㑈�""B��豊 YBRmS�"O�����	]`�E��,�"OR�X��b>~	;��C=Ny�ar"O��$�Na���� �  !T�]��"O4�1$M�޼x�a�-V:	�G"OH��u�Ue�^�8Fc^�L�ʦ"O0(����4(sD��8>;T��"O2��q"�'�����f��7�$�"O���6l.@��1�$�1/ -Qq"OyX�.ޓq��t�P�G�	zI��"OJ,�g�.%��QV
�%�"Oh;��ɳ]���F�Q�0�0�"O�(����s�8��� }�d9�"OPD��mX�c ���ƈ?�v���"Oz��j�%0���*�����%"OVSDؿrP<e:�Z%q�"O֐!4m�9Y��xb&bK"�.��"ON��go+T�4�6`����&"O��J̞n��`��!�06�~!�"O��AP&�ua3��,%�V"O"�p7�@���΃4q�p���"O6�j�GT1tĨ7�+D���p"Oht��M9T<n�XW�8{]d�"O���"��R��U�D0Z>�D"O6���g��]bZMr�"؅EG�i�"O~�VJ�����ͪJՄ��"O�� ����@�9Ҁūe���!"O�Zb�Y�~�8�CF�����v"OxA�5�ϦM�`�W[?~�
s"Ol]���=qJ�I���p��q�"OTU��сr��5�e�,|�8s"O~h�փ��s������N$�R"ONl{҃��}Q�N���1��"O���4+M0y� M�O�{ꄁ"On�H3bå_�@5�Fg�&�zI�s"O� ���a T>�(]F�F-Lg�DЂ"O�mucR�N3���dD�3ZL@"OR��.ӑ,���B��/�Nt��"O0���,@ ���k<��	V"OZ��T]�2(J1�°I��b�"Ot���N�I]̠�"��/��4P"O�Ya�䝡%�p+���
Ni�YQ"O��T�I#@�q2�6dd�)F"O]0%*̑A�9�aE�B��8(2"O.�{5�Z��T��fĠY�4�:g"O�|1�jv�[�&^�P��u+s"O&��E
��'"��`��&_���r"O��k&'BO�v�$���e"O*�h �R�E��q��!%��,U"O�5��Ϛ3�VL�� d�����"O�囒�Fv�@Sj����"O���4bٺ1��@_'��B"O�H��Ppy�`bC&2�ڠ-�y� �d��š��م!�s�n�r�'}�+ƎS����5�̠�(��'�ȸ)'%��Z�����M��i��,#�'��9� �&Sະ{�N4a��Q{�'�"yǥ	2����C�\����']]����V�����%� V���R�'�� ���ѲQ�� �C�:~���'۸x'��<�L�ccE�/Jn���'���!m�v���N�(��s�'��U�(��FpVE�R�Ѷv*N �
�'Qb�9��|t�"�ى���
�'��D3��Üxld�u┨d:Z�S�'t(8W��2ڴ$�3rN,��'զ�G��KgBd;/�!*�pA �'^�ؕOE[5���cܭ!�ؕ��'(DB��[c�hZfB�/M�<`��'�ʝ"�̋�E(j���P�����'�@$�!L�!&4���w��3	��2�':���$��?(zL������R�'AH
 ӤMS �9f$��|���'�zF��lt�0�Ą��t�����'Ɋ�C��1'Q�9�D��l]6e�'�4�s���=~J�C��$HZ�'~(�)s��%ErP[c���`��c�'x2�Q� �"�I�O�<[�����'p�Pd�5-�T��u#�(M��U!�'�$eكK�} ���᧐�p�u��'�"�J�)�WˎU��D��HX��'ְ���n�/2�.��"�W>/���'9l�S�@���)U�Ђ�L���'~�P�R��\uڥ�Ɖ��6�@�'���B�dI0s���;w䙽�(��'������B*D���E+O��q��'��0����<�����Aiz�"�'贡�H�j�����8&�$�	�'J21��]�.e� �s�W�.0��	�'>��J�A�Ug䀊 	Љ �>���'�{ע�z���;�O�nY��'jv`HSI������`�T���'iph���Ք5B68s׍��U��89�'f���Eߍ @0�Ɔ��9��Y�'�� ��Ǭ\��p���ҐG�:Y
�'��i�  ���   �  �  �  '  j*  �5  0A  �L  "X  hc  �m  6t  '  ��  ֍  2�  t�  ��  ��  t�  �  T�  ��  �  V�  ��  ��  )�  l�  ��  ��  =�  �  �	 F : ]! ^)  1 n7 �= �C �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'�~�����|���ZW��tZ �'�R�'�R�'���'���'���'�jp�5*��I�x!�b�7<��'���'��'��'���'=B�'�xt �j	Amtp��@ИS8���'���'[��'��'3��'|��'���Eb֖_�x�b��ڠ-�b-Y�'[r�'TR�'���'��'���'UZ��)���pi�f�0,���'���'��'���'���'��'�\���A�SJ
hbB��,l��U�#�']��'�"�'���'b�'�2�'(�����{�f��D�;��'��'I��'��'���' ��'1�����^�p�l-X���}�Ty��'�"�' R�'fB�'y��'���'����F��
�1RN͏@�"+3�'pr�'���'TR�'2�'���'~&Y������ֿ�K"d'�'�b�'��'��'���'-��Y2c@6����P�y��tkS;5��'�b�'�"�'Z��'���'?�<�\-qD�ѕoSb�"&M3<W"�'���'��'���'�`6M�O,�J+"�I�F�]��9��L�I�*��'��T�b>�z����5H2�9+0�˩g%���R���J����O|0oy��|Γ�?)�&�$�<!ⱉíURȕ��Җ�?���{j���4��$j>a������<�N�IV၆"r-Q��F�.]�b�(�	ry��	p���w$̳+OH�����(3�@`�4^�,��<)��4�k��Ƒ:�.����®���Pg�ҡQh����O��I}���!�0��V<O� Y���>�<�2�%��B�� �5O��I��?!T@:��|J�{%> ��G(ƅZ3ƐC������D-����z!4扨-yx���'�[�p�h@�H�x�̍�?q�_����ޟ����D�2�T��#�	+!gZ���a��O^���!H����O9�?��g�O��È�^�	�#(��@t�pç�<Y,Ov��s����I�.|RL�<N��tb"Er���ݴGc(��'�b7�.�i>]�w�3iy��$jݵ=�����~�8�����	$vv�]o�D~�<�"!���_ۤ0 ��ʍ%.�aXW� O��8���'�T!��'6�i>��ǟ�����\�	�<�B�IԿ	����&З;��A�'�~6�F����$�OR�d�|���?9�B�,��òm,-h��VD�7M-�	Ɵ���w�i>��	��\8vƛ(J,p8�g�.�@���9��oZe~b�W5,"�h���?!6*��<	)O��*��{_�i�I��O�����O���O����O��D�<���i�V���'��鱓*	�{�N��':���kq�'��6�<���OD%�'�r�'�2�����f�:�f��Cd�_؉�B�i��O��M���s����߹K�S>�y��ʷYA�q���t�t�I����ԟ��ğ����Ń6A�䄃�eH�P݈I�UF��?9���?��i� ���_�,�ڴ��56��b�*ԴZ�I���0
w��AK>���?ͧ�(�ߴ������g$W�o��i��#g�1X$挞sD|�	�����O����O���^�L-��3��-t���� �O�V�1#E�l5�ʓN��ƈ@:��T�'���O�'��E��0��H	�hqDq@1	J�y��'��ꓙ?���OUR�Q#'�i2B��B���2�0Z�L�pFS#]���?1	f�'�t��I�4�	YW�MkoP#J="yx��m���h�	ßL�i>����8�'<7-.����	O�lu�EZ�{=���H�<����?),O��d�<)�Z�@��V"R� (��jW�N�����?�ԩ���M��'�����M���d	zo`��%śg.(�䭆KD�Ķ<��?Q���?���?a)��="#CU���D����\�T�C��I3��ߟ4��ɟ'?�I��Mϻd��ԩC�7v��Yxc�3[U<�J���?!O>�|*6Γ<�M��'o$�j4	E���(�pFV�tb-ڝ'�P�Q.�ӟ��P�|^��Sܟd8�nȉ@K����,ִ�,ږ�ß���ݟ4�	fyҠu���+�O8���O:d1�׿��Qb���	]��y*Ç"�������O����@���x����FBњ#l;?�4 �f���7瘝��'d��D��?1fO\�$�^���B��\H�c���?����?!��?َ�Ix>1C�
��7��}0��4C)V�J@+�O�n�}S�����<�4���y7d 7|-R��6oL�S���E�ɺ�y��'��'H��豰iU�i���	�?YÇK���HS�Ř|<��&�C��'x�	����I��t�I˟T��;4.X���']�:� W�ʳ":�'�,7���BT��$�O����b���<�'hԔ3<�"����Gla@�-��	�|�?�'�?���$z�M�m��U:FP�2�[�)M�Q���Dڜ�/O�4�dL��?Y6O�ON� !?O��M�R��m�4ga�x�3Naj����?���?���9q�=K*O<o�-y�d�S��� /N<'��}�B�eQ����M�O>���3��ן��	ߟ�!C%�L�� ]<>��� �e�	�el��<	�� ��JS�*��' �t��� ���g�#<Q(L3���=z�s8O|�D�O �d�O���O`�?Q�䬉�{D^Qk�f�8�R�9�䟤�I��|C�4���'�?y&�i��']�H����=?T:�	p�N�HR�|r�'��OQ��c�i��i�!�GI�!,⍹$@q������I�K�'��d����l���P]��07.ZU��uq��@�	ȟD�'C�7uD���O"���|27Cz5�8������@&&�T~¯�>A��?�O>�O�b�I�ˈ06�LRr�G5�İr�)�D~��p�@���4��89��I�L�Oz=����>���C�J�?P8��@��Ol�$�O����O1��˓D��v��m��QҦ���Ti����"�F��y�F�'���y�T⟐	�O���\��FTۥ�X�q�U��(��n��$�O�5�4�q�F�Ӻ�%����(�<ᷥK�
ͫ��A�]� ��FM�<�)Ot���O����O����O��'V�t�d��"�=�p��M�"ೡ�i��X;f�'b�'�Enzީ�uMS%'��Tcϯz��ɀ"�ڟT�	b�)�Ӣv_~�m�<�'��+cW�� d� N�ջD%�<9ve�
A>��P=�䓉�4���$��.���H�zc aQ������D�O����O���E.Q6:��8�I����8R� ؗ���K*�����	"��=�?�T����ߟ�$��x�g^1K�*���Y�r,"'�>)3�&VǞY F�x̧RƖ�D�8�?�!�����q%d��r�KlϦy���� ������D�O9ǂ�U95�5�;���2���\}�`uӦ�Yq��Od�DMƦ5�?�;���qJ��B�ͱVϗ ����?)��?q��1�M{�O��S���1�*"fҋX���P���8�$��f��)�$�O,��|���?	��?!�6�� 2� I��ƈS��6�\�*O~(n�Fmj���֟4�	@��.A>�a�c�����"�@́��80�T�d�	i��|����?)4�X�{ծG��>W���SFC 1pz|0UM����O�����k���O�ʓN�^8D!�, >��H��1p��?����?����|�.O*�n��u�d�I�y��@TM�z��9��J�7d���ܟD��sy��',��ӟ��iޡ��)"��5ȱ@��E����Yf@�B�iM��O����������<��'��R'pdF�&��|0t9���<	���?)���?����?�����V�P�pta˴V#t	��%�T�2�'2�r�$���:����զ]$������0��U9���f��7�4�	����'ߜ�e�iY����z����t~D�s�g���կ&���V�oy����#�Fpr��_2�ܭ�-N�u����4\�$(:��?���i[�=J0z�C�@Ж$���:��� ���O6��$��?A9��
?p������+N�a���#����0a�3\6�����Jş�h��|rE��-B��`B�%H��4đ�)��'oR�'Y���[��1۴?�N����3;R�Â�W.O��!��N�?���'�����
n}r�'Q�is+��t��ܸV�ŧP�,��'�ҏ;Y`�Ɛ��ʣ'�12�T�~
eY�zl�S�Y� ������<�/Od���O�$�O��d�Ot˧��X)��N�&��E�W�L-wٲ�(`�i}6�ۂV���	�?��HK۟���)�M�;Bs8$��ۃH��X��͑!v`L ��?�L>�'�?I�i����4�yb�32�9��Ȝ�@�<X�b����y������������O����3"P4Q�hĶ����B>�T�d�O\��O ʓa��b�b��'!M�^ަ���V"H��5/&��O�y�'^��'@�'f�f� [�� z�`��D!��O�q��E�{	6M/��	j����O4)x��\�V�TX�A�3R �"OTa�爑SBQ�PK3�zM@ ��O��	�0Ժ���Ob]o�\�Ӽ@�S�S��d#ׇ0	��q[���<9��?���#�� �4��$�2]��)��O�����iV�=��%C�Q<tJB�'d��y\�����?]�	���	��;�b\�h,M�0�ڏ`�&q�5�nyrBg�~a�&)�<�����I�Op��Y	�.g#�;�x�x���crʓ�?������|B��?�,ǵk��m[��#T�]��P%1�h9q�4���W�U����'*�'m�	
I�JQ�E���o��\@CҊ/�����Ɵ���џ��i>	�'r�6E�gAX��M�$	ri�T*�8[�^19G�T^��$U����?��]���IYy2� (} Y�r`�
RT*i�-,U�!��i��I��$)P�OS�<%?�]K������nb��i�:7"4�	^��  �g�63NQ�w�2y�V�;A�M����	Ɵ����'�����|BhW�M:���Óed�Ԋ��/6��'����4(ş}��v����h�w?��s2�&+�|��AY��x��O�O��?���?i��L�>�ʣ͔:bZ�av ҃G��1��?�)Ov)n��@A�	͟ �	b��5\	ئ�.+�>A�t�5��$x}r�'��|ʟX���Q�b�N��gT(Y����u�E����:wi߸}��i>�%�'�6�&����{� ��Sa�-\"��,W�t�I͟���b>m�'հ6��o�
10w�X2=HI��a�V�\c���O��$SǦ��?$Q���ɧ�M��CK�Z��,#���//� ���şpV&���'���҉��?���� �=)��A�72��#�O�����G8Oʓ�?���?��?�����	I?$=&����	/�MS���)��DoڣPF�a�'U����'C�6=��g
+/ 0Q"��2ު!薇�O0�D ��IލU��6�z�x g�+m5H��C�zV�9c��i������O����a�Qyb�'��]������~������>HFr�'���%���0�M�������?!��
{���%�?�|����?�/O���Y}r�'�O����� .�����3fϲ�1s<O6����V�F�ԌQ�Z���S<Y bFM���!宊�x%���E�ڵ��;��^Οp��ɟ����E���'��[��/�.5�aیr�AR�'uF7��+|�4�Y����4�h� +{�!BK�q�x�1OR���O��$?O�6�#?���Z;��)�� 
LH(V�M�A���b�J�,!�H�H>y-O���O8���O��D�O�����e`n]�q�]:�H���'�<��i�f��t�'d��'��Oerb�Y���҅K��O�<h�o�2<X��?�����ŞF�h�r���+�� �R�>!�Z������MS�O����^��~r�|_��re�N<�.py������N�����ӟ�	��Hy2�d�`�Ѵ��O,��gbQ�_zxh�γ1}H�aŢ�O6�n�M�@��	���'e��PR�ڗbȴ�bP�8� ���A0=�Ƙ�@ ,ϛo ��%�J���-��CJ�pb�����L<Se9[X�	ş(������Iğ���y��6�x6#ǯ�j$�@�˙�N��(O,����M�g>9����M{I>iR!�&y�
J�d��!޵�䓫?��|�Q�,�M#�O�T��玺�
��0gK� #�L�Q��D���#�'Z�'x�i>M�	�L�I���0PC�K� ��3d�y�a�	ǟ �'B����-�	ڟЕO� ���h�R]�����Б:�O� �'���'�ɧ���(w�2���F�.?����𯑷5�^�r����!$B7�Bgy�OU����P@Ԁ��/*c�i���'{��y��?����?��|���?�)O(�m�K��3/&u>��*f,Ђ
8���gf�ٟD����MH>��Y��	����)O?__�T���L3�ʌˤ�ٟ,���S�@o�<Q��>�	�?��'^~ V�Y;����q#I��9�'��͟��Iџ��I�	���Z{�a	�;I��(��']�7m;)1$���Ol�-�9O@�oz���n�f0�@�����x��k�ޟp��d�)�)%n��l��<�P��fcЅ��/1�[6��<q6FV�ZK���@8����d�O^�$���|�����^a"Q��,
�R�$��OX���O��^��)K<0���'b5S��� z_���E莕;b�O>��'c��'W�'	t2�%�^H�7�p8�]������ !7�|�rc>�	r�O�D�5-_$�3bo�,�:�z1�F�z!��ڠ<��X��ݰ@���+ɾDb����ş��7��O������?ͻ#�X����'?�xU�äz,�Γ�?���?1�cC-�M��OB�2)���d�<C���>V���AK֚B/�'��K�'R�ɋՂ� $\e��`�a��O �I�� ��OB�D$�ӝ�^h���Z�<��*ۭɶ���O~���Oj�O1��m��e��G��J��V�(�ޠ�0Јs��7�ky�ŕi�D�������$Ī���F���t��t-��@�`���O�d�Ond�3�r|�ʓ��i^�^%��>j���/��p��[��[1^b�m���D�<���Lg����0�'Ed8���Z�9ve�9J��(�7È$��f;O��$����X��<$����)���IF�s.�x%O�Q�r`��?I��?a��?a���O����F5["99s�ʇd	$�B�'���'��D߼��)��$��ѩO�c���8�d�W�Xɣ%��@�	�H�i>1�0��ѦY�' lt���B����O�c����d��g*���䓲�d�O��D�O��$J��������y!�G�=F ����OZ�Sڛ�Tl���'�rY>�Յݾ�©��֤b��)X*?��W�(�IΟ�'��  �|9�ӽ{�(�����dǂ� �ė�.�����A~�O,I�	��b���yR��M�=ZjI=vA.]��Z
96��'��'�ʟ��R0��<�"�i�M�EJ t,�Z(O΀���]��"�M;N>��'y�	Ο�Ò��p:pq��̊ �L���������Iw�vm��<a��|�Xt��?��'�j\���o�����Ə`���'��I����P�I��$��P����$1̵��� �����!2�7�� |Q�#���O��D�����O2��J��wΔz6O֖#���$ˊy��	��'sқ|�O��'h�P�5�i�����\�p�荒+x���PN��x��E
�� ���֓O���?��.��#�퍻O�=��D� A��?Y���?�,O0�oڈC����'Djȝ2 �����!�BT[�M �"��O�5�'@��'��'�Ʊ{���A�����K�O"���!�7�Ta�S�	F���O��FL�84��,��2��굉�O.�D�O�d�O��}���^dT�t�5���j֧�8!Y셊�W���\�Z��'��6�4�iޥ ���傑J +2h����q� �I����;M>nZt~2Ȋ<�i�g�? ��cr���.�� Jti�/$A� ��2�D�<����?����?���?�Ef֮:޾8y��%>V\I��\	��d즱���J۟��	ޟ0'?��I�w�`��EV+$@�`��
�,�O����O��O1��$;`�0/F�9�'�>��b�/F�Q�̈Q#h�<���>�H�� �䓒�䛣4�VD:�Ԭit��l�p{���?����?�'��D�릭R�J���c��E2���ʞ{`qP�e��0 ܴ��'듍?���?ٰh_1�hJ�C�	#-����eJ�um Q�ش��dK�>i((�	����:o"��*��ݳ�zX2w5O��D�O��D�O���O��?)"!� lt9��t+��; 'Kџ ��՟p �4^x`ͧ�?1��i�'ČuI��5j�y�V��
((|R�'��O�����iu�I1cs�9�͵J=��r�N�auJ8�a�ɠAc��6�$�<ͧ�?���?qQ�ڸ0�x�r�)M�9�6���?����$����agH�ԟ���\�O�h��$H���j����a�����ӭOn�D�O�O���yNp�@�_(bj�Q��^�DA��䄞mTU#� 3?ͧ5
��� &��e��ث��� $m���T�
�Ii�<����?����?)�Ş��ğ��q��$��"��ӑɌ��y�D�8 -�'�$6)�������OX�!��
2?Rx[f�S�l} ��ъ�OT��ƌ$f6:?Y��ďߞ�ryB�\q����܇#��۔u��d�<q���?���?Q���?�)�xM*�"���*�H� 5`���g�����$�埀�	۟�&?��ɞ�M�;P���a���QN�A�@��8~:���?9M>�|�5IE��M�'��m`F�8gL���
E�q�'ƈ�r����hQd�|�P��Ꟁ��"�j�f���B	I�:�Б��۟�����jC\Xy2,��`�aA���D�O�̐V䈅���o�`Z�W*�O���?	c\�����%�d��MȊ��x�g^����@Je���ɓ'%�jE ލ
�E�'M�������:��'v�!(���	�#�n	 ;�4A��'4�'�R�'c�>��I�p�NI`�C �x_T�14hRሐ��
�McQA�*��D�����?�;���?j}rd�7WI��̓�?q��?1f&��M��O�7]K��� =A�@<[S�	n���Xpkx�n�XN>Q(O��D�O��d�O��d�O]��lԵq������#��6�<1��id�\���'���'��O�үB+s�Ir%\RI�v��|�4��?I����Ş5<Dej��� rRPh�ca���x��f�8z�(�`-O
�2���?��<�d�<�(�3K�เ�E�͌ ��Ş��?���?���?�'���F���Qh�����D���r��C��|�Ta34N�̟`cش��'���?���?i��(2�!��i	���2M�>��)��4���������Ol�O��Fܷcr��礂�9���ӳ#A�y2�'|��'	��'A���U�y���ea̸��Ē���w�T���O��$O��h�Iv>9�	�M�K>)tEϵ:):�P�H��%~M��ia̓�?�*O��Z�yӮ�BW�\c�T�LX�B��.���l
�4D@�$լ�����O����O��d�)2� �E�I��<�f���*�����O�ʓF�v������'lBR>�h>z����b([4˪}D<?�wU�|�I��'������S�A<S��@�#IE�n��Y�q�+@�B��F�H/��4�*=3��&��Ox4uh��G�\Mi�̗�P��e9W.�OH�d�O�d�O1�F����ڪW�DqT�Z(0�(�s�ɭnl�s��'�Ҩ`ӄ�XR�OB�$�K�|@gK�pFN@Q��V�R���O�`��GkӦ�Ӻ�e��7��Ͽ<�$A��Mè��w�܄��u����<�,Ot�d�OH�d�O����O�˧>b�J���6x��:V�\� �iyj�ˀ�'V�')�OUr�q���<i�z��P�U�,�(�T��u�j���O\�O1�Dٺ�}��扨'9� ���ߐ),����ꖵ�l�I��Y���O>�O���?Y�0g��(��Q+\�J�V�����?	��?)OplZ}{|��ɟ���C��r�/PJ �b�)��.�ȴ�?i#U���	ʟ�&���F�4U�āѷ��q¨��B<?�/�`}���"G���'j��œ�?�3D�n��18�@	�J��S����?a��?q���?aI~�B[�|���$Z���'B����#�a>2M��Vg���T�>��'tb�'��I���7�ְ�AeX F���QI^0Di�	㟸�	��\����ϓ���L^5En�mM-+^! M4��U#���y*2�'�P�'�b�'=��'w2�'�b��\>zZ�j��QXT�KR��1�4=ތ����?����'�?!q��;Vn �R�;!?�)�v�ˏh������t�)�[Ov�p��� g%��*�[&kL�q�gP+7�"(�'C��0чޟ,�0�|�W��c�a!RO��B枥�������	������hyrhg�.��f�O~�dĜ9P.�Um�&f�*9�&7O�o�g��v�����T��ퟐ�r�XJ0����6d���{VnL3+�^%nZM~�ٲ1+�PF��w^\=�#μ3�Ԙ����JkBlj������(�	���	ğ���덺q�|�
���5�	ӱh)�?1���?��i�a(�O���h� �O���A�3;Iƌ������<(���*���O��4��Q�7&y�j�+��P� ��v���aWhUb��N�A�lp�͊��~ҟ|RU���	П���؟�*�&]	:C���3Ö�p�� �g��H��Ly�z�8��.�<�����^m�hjW��m���rW&Ǟq�ɸ��$�O���/��?��%搟b������iu/J�ZL��v �	��FA?	M>g/ �(�QDY�R�D|C��
��?���?q��?�|j,O�io�(c������4D�����BJ<�┥ΟH�I8�M���o�>���a$6��	��D����6�
H��?����M��Ond�Ǉ¼��O>�Y3���aT� �˟�V�
�'�������ܟ�IƟ�����ӽS|��oD6�Z�P��2J��4$j� ��?	����i�Ol�D�O�n�7�6C��5|�L�*rM�[A��d�O
�O�i�O��d�"R��7�}���# �2 ���C���(u�j�
b-g�,����$���6��<�'�?A"aG���%���ͣ|���A���?��?������������T��ٟ�"f M.h��W���J̾��j�o�\�I��	J��I�I+r�$�:�O
�n�j�V�I
U#S�M�d��4�Fg?�����<ː�\�����p\�	r���?����?��?�O5b�9E�'�K�2*v���q+��,�����z��$��yچ�<��iB�'(�w&&��dd@�D�0	�&ڳ�@j�'�R�'Y���]���3Ox�M�}	���'r�"44�H�ʩA�CX%v(ͣ�"���<ͧ�?y���?���?��̸E;� ��Dʆ١b��z����M;�eH�����O�"|�$�*M�0I �D�c��L�����D�O��i�ɧ�O1�9�BO'}��y�%i~���� �2}�\��O��(���?�t%2���<�Ջ"-�	�%H�i��\�(A��?q��?q���?ͧ��DW�+�V�@8`��"PN@��P@�}+2.�ğtz�4��'�@��?����?�"���;֦PQmB'?F�`,�:!��}8޴�����M��؟Ғ�����]�5{�-6�����!s���O4}����OH���O����O1�p����	 b� *p�T�S��MY�(�O����O.Uo92^I��П��Id�I/i���r�ߐTd��F�F�v��&���	������+C5o��<��^�8I9T�ڂY�r��C8��\xs,R�F��d:�����9O8�X&���[D4��c-��?u�M��ɿ�?��kП`�I��4�O$6 �U�� 4Flc6�ʞ8��O^��'wB�'7ɧ��UV�r�в�T�_�)p�Z# N^�`)Ίc46�Wly�O`T���k�܀��U�EF��UeF���EX��?����?Y�Ş��d���� E�r��jT�P$����%f8!�D���J�4��'�L��?y��4�����u���a.��?��X�F�!ڴ��dưPC<��Ot�	9�<Lb��ʬ+6�T�⡒=bz�,��L>턼Z�BJ %
iCg��/0��#�Ϧ?̴2c��3~BČ�SN�{��fC�x����4�z�@sA��v�$�ė<�P1Ѣ�A#:�#>i�O�5�P�a�h�"| 8�%ɏ:.M�X���8�~xbW��(J��xC�狊!� P!j�,`9p��ʈ0:e���G���G��iC����`�£Lh���T���8;��� Jr�jťːS)�)¢���\��ũX@�\a�b&dS�M�!zF0����T�j%�Ħ��ɟ���?՛�OD��Vc�	M�Zy`��F�:z�@�i<2�(`�'��'�3?��	�TH���@��]H��A�@պi�R�'��`\���d�O��	�\H���Ǣh%eHDJ�� ��}b��',I�')��'w�'Z�z�3�1-WK--��y�i��*[�-��ꓣ��Ox�Ok��lV� dED�l]t�)�@��	��3`t�l'���I����	qy"J�} &���	��$������m��M؇�>(O��d9���O��$�#ٖ��U/OZ؀��T<R� �[���O����O��ǂ�'>�^��h��M�Bu��c��$��(1C�i��柨%�h��柠��A�Y?�0��b �p'��yTtc�BG}�'JR�'�	
�f�#��"��-����-G|}��@&�	g8��n�ßh$����ß��$�R�	��a �T�a�,x��i���n�Ɵ���Ey��p��꧉?���bS�g�D�^�n9^IG [W���3�x�'��`E3{���|bן��hrI��W䩳gOƀ("�([�iL�`Wh
ٴ�?A��?1�')"�i��f��|&e�[�t�&��@eӮ�D�O�l
0�OȒO&�>�V�*X�AP�#T���(a�d�:�k6�����	���I�?Ѡ�O
�R������.�8�Qb	�+R ��i�x`z6�D(���Hh��>����ͅ�; ���'hٌ�M���?Y��c��)��]��'F��O���e�9���Ӆ=��ar�d���P�O����Ol�Ė�X�rh o��D���� ��{���mΟl��N����<�������p@߅T�nH�T
�pt�U���G}hʠCT�'�R�'uR]�	GZ��3K�7p�=��g%|6`��O�ʓ�?�O>q��?)"g� ��`�+�<Y,Ih��>�B�H>����?�����x��u�'"XK�=)�P���l�61-�~����?�H>����?�B� B}�A�C@�ِT��-�"q�p�ø����O���O��G�`���R?��I�CJ��;^�(�H0*�%�
�U�۴�?�J>���?1N�ĸ�� qe�T�d��K70�6@jǷi��'��ɹȈ�K|�����N��>����NЮQS��%�,�'\��'}��yZw$dYb��ĒC�ܸ 0���d��|۴���D�>4�(o���I�O��ITr~R%Ï|~$�CbL\$i���(�M�)O����Oa%>m%?7��Lz���Ŝ7v��0�*3��F�ü��6m�ON���O���NV�i>�`2MC|��8�"��U� ��P=�M����?�����S��'�b�7f��ш5��@�H����DE�6��O����O,���_�i>Y��k?q4D'2<�s�ؙT펙��iSڦ-�	F�ɭ�������a?Y��D=���Z;�]��$�ڦ}���{�T]�'��꧉�'�0�b�%b�@�㇛�p�p]�m'�$Ј$1Op�$�<��S�hm�SbN�e����c+״@:½���ɶ��$�O
��+�	�p���Z#팅y��l���T02�@lZ�'�Zb�l��Cy"�'*a��֟б��ǐ�	�(��"Ϛ��!�b�iir�'�O,�d�<a�����q�s�0w�dx���%�<�"�D�O���?y�����i�OZؙ!o�=�5�Ŋ��hJ������Ħi�?�����dP��'�Nx���(,`L`�v�1epvt�ش�?�����䚒u&lt&>���?��:'��1�ߦq���`���J�rO�˓�?1����<��*�������TRd�c҆!U���'�r+ܚ�R�'���'G�4Z��	��EKS$��y�|�Qb�5bY*6��O��oDR�DxJ|�s̖2gR�P�l�˨�z�,������,��ӟ����?՗��閲~���q��:yt��k�HE�3�x�'�(4X���I�On��7���<�>	�ã�Y�,����������8��t\�CO<�'�?���2θչ�"�=p�Z�Br�ƼT%d�k��i��'I�I ��)�|����~� �A�>�,Li�R%��۴�?IP,�����X�������ЊJwYD}3��ȁc$x�'�t�� ?)���?����䑎?��ݓ��^�/�j�c��:x���
}�	����H�IqyZw&^�BO7tC�-c��Ԇlm@�4�?�/O2���O���<��hD���i�#�`����> ����H�Q���韄�	����'�V>5�ɚK����U���dvb�#g���XUF�j�O~���O���?y�Q�����O�����V��8y�oڸi�Z�Qǫ
Ȧe�?����U�'���z���3!ײ��a�Ι�8��4�?�����kĈ��O�b�'��땧PX��UM��X�t@I��Ĩv���?	���?aa��<�N>��OVBB�޷ ����a՗�>�ڴ��ţ=���lZ� ������Ӂ����i* ��G�̸��D'�0ꢽi��'�ڔQ�'^�'�q���q@H ,�r$zJ�-�����i�X�
��q�d�d�O����0�'[�B��M��ۧa���Ǩ~!F��M��(��<�����:��ߟhE�����v�!x�$�A!��M+��?)��x�����X�ȕ'���O�8�1*�> n�(+O�m�`���i?�W�<peeo��'�?!����4`D�� T�r$�VpD�`�g�3�M���6�<�Y�Z��'�Y�S�w��a隭CW�J )�:e\	�'*@�'���'8B�'��X�dS���D�R��/;n4�R�G�l�  �Oh��?�(Oj���O���
�%��P�b��*,��N��)=��xw>O���?q���?�+O�S��E�|jUÄ�l�@Jք�`�d�'G����'��V����ԟ��ɰ����
e��������7,�� �ҍ�ߴ�?����?����ެc�X��O*"�Ǵ)1��ZFXҵ��^�d$�7�O�ʓ�?)���?-�����ܴ?��(���-O�(�l�;�oןL��By�&��b�v꧁?���C3m����GÆ�C�@�[�IƟ<�I��PZ�)s�x�Icy�Пle�V÷v�)��Iϝ��r�i���5#��Z�4�?���?y��"�i�U��"E�Dv�P��_C\H �d�R���O�2f<O����yb����J�@�C�/�5z��{���,s�F�K>z��7��O��$�O��	~}�T�����.d� Cݒ5�\�a���3�M{pJ��<a�����-����`�� )9�,H0e��;1���R��6�M#��?y����Z�H�'e�O$ͫ�@�#��℃ Q���i}�I͟D�%�~��'�?9���?��OȺ}�� v���6X�HӒ�B�^��F�'|^�9Vi�>�-O:�İ<����"�5��4��ˊ��T!���U[}"䗃�y�Z���ݟ���kyB����Ba��j�0��C������>Y(OX�D�<Q��?i�����f^ry�pk��z���Ҥ��</O����O<�$�<i!S�]N��ƀ)��-aP��8v�n$��	�yI��U�4�	Dy��'��'x8�R�'Y<A*
�7M!�qPr�P(W���r�{�B��O����OL˓|_�,yUX?��i��r���n��Hb�ju�
�Ѧ`tӸ��<����?���4͓��i�dQ�0��2)����ߗ7� ���4�?�����$K�_��]�Og��'��D���kj>��V�X\��yW��Hc�>!���?���
C����9O����o� ���ɃLa��QЬDn7�<��'�2~��'���';�ĩ�>��;�T�[�H�5`�h1�CϛV2�m�����u�l�	矤�'rq�� �A;�@��
��gG�CfD�
1�ifLͨG�pӄ���O@������'���/�f�e��0K]^�c8&�a�ܴo�&�ϓ�?/O�?��	�XF\� �^���K�-H�C* 8��4�?����?��bNz�	Ny��'%��̗�:(�L]�R��Т�*ߍPX��'���'~$�������Ot���O0�k�'�(s�n��U�J��KЦA���6��mɨO�ʓ�?A*O�������*�*�h��@���h��R�0��B}���	ܟ�	���Nyb���@X
.�C�><���BB�qg�>�,O����<���?)��k]{M(s��`%.�3n'��"��<)/O���Ov���<!����U����&<�(��cA�h���a�*��FQ����lyR�'��'a  ��'x$�R��E�����92$���`Ӯ���O��D�O�k zu �Z?��5$��	�+q�
Q�m3**��4�?�-O���O����_��$�|n�?r 8�F3h>*�Zw#Ly��6�O���<��L�M��͟��	�?�� ��7f��xE["�D�pB��)����O�$�Or=8�<OT��<!�O�`�Q�\�<!f9�gZtW��X�4���U�7�ޭoZ����	�\������t�w�����P�� �'�L`���i�B�'�R=c�'>�_���}�Ul�f��Փ�/Y�{$�A�R̦�X���M����?����zV_�ȗ'�01a	\<��%;E,�U��*a�!#W5O��ĥ<���t�'����+82L,��T<M��mr���p�D�O��DBa/F��'2��ܟ���j���H�+y��E�O�:P mnZ� �	���㒨l��'�?I��?)��k!ܽ��0k�.�ApDPk��v�'�I ��>�.OR���<����l�we�ݣ$,��P����a}BcW��y��'���'c"�'���(E��� M:��c� ����&� ��ē�?9�����?1�Kd@5�.)&�S$�V�3}< ("Y@��?����?�*O^}Y����|�d�uR)ISP�c�����n}��'�2�|��'�B�1u�D\>��͈�hܖ`F8a���-��	������'YX�Ғ�(�	��
��@3tPg%��~���irӘ�D$�d�O���F�i���5}�j�6��q	��S#kϔhP"���MK���?a,OT��[�ǟ��6L���,ĥ_9Vy�U�lw�II<����?ylN�<�L>��Ocbp8g��	V�9k�.�9��ش��d��^Ȍ�m������OV���\~A�,JD����L�>��p�[�M���?1獄�?AH>A���Ɯl���rLlR��C���M󵯚�OP���'���'�tf*�ɝlR���)o��}�&]�N#|���4F�Șϓ����O��@=�h��Q��'[��%`@D�=��6m�OH���O�q:�gY�I���\?)vM�/�H�(e�(Ʀha�.[Ҧ�$��X��x��?���?�1�I!Za��
���_��͸U�#u3��'�Ęp�4��O���*���Fp���06V�@aL�6���k�Q�X���g���'s��'�O�̥��C�*��ƈ��)"$@_5N�D�H<y��?�H>q���?�V剁ri�A��ܦ745�w� -}P �����O*���OT�����7���b̑ (�0 ��Ɉc(���W�T���X'�P���h��w�� �']��]!�����6�Z=��L�'P��'��U�|+���ħ�V�)�˜�t.u!J�_@�a�i��|��'��J0v!қ>��(շ��5H_�s]Z�ٴL��M����?)O)��(w�Sٟ�s�� eI�=0��D�AB�c0]0d�3��Fy��'��O뮜#6bAᘳ]< �0�	
��v�')"k�6��'B��'��DR���{���ӗ)�jl~ِ��|<:7��O0�K��DxJ|�%d[KFT���u�hbƞ�=9T@	8�M���?����BQU�(�O�z0Q���-!���ɓ�K��H�Gq���d7��䓺?�BK�#Y���zd̆�K�rtK4�P!��v�'��I:JѸ@�'��	� �<��ak��I�+�m���U:�I�ħ�?����?9�-� Ҡ��ě!I�N%�1- �{K�V�'��):X��[��6�2�$&Ύ��so��05���䇜,/b�'���f&0?���?������B�)[��b��-C��a ��)H-j�ӣ�Wn��T�I��?���k ,|��d@�d���1��I���<�<9��?	��?A�O
6pH�O3��ϸ�	��ҧ6i�[۴�?	��?yL>�����%f���L�o&E�T�CW�(�R�Y	��$�Od���OH�>jM|��oN�B��Α,|��<
3jZ?U��F�'Q�'�R�'ɾ-��}Rܔ$\��ZR��,axn�Y1Z��MC���?��O"��K)��O��iH#��e0oׄ8��HR�	�&��Iӟ����>���FU	Qߐ���b�lޙ7N��M#�O"1pG%|�е�O6��O���O��Ӆ��� ��c���] ޔm�������G�\#<���'IJ�Ur�B˳J�X���?р�߉�M����?������x�' (�3����xq1�
A.*����+hӚt;q�)�'�?	�A�#wMX�bq�A3��E*3����F�'-R�'E���1���OH����x���h*�DAb�X�M���o$�I�|�c�X�����I΀ ��T*�9R��'��&�hp��i�2�[�~�c���IG�i���=����Qm��:�u���>!�aWP̓�?����?��O��h�n<�<�Cv�Y�3�h�K]6�c�`�IA��ğd�I4}�l�ڧ�?
�}ӵ�W���%xf�8�I^���b�˚#F^�E�to���Xs1�^�()��"(ͱ�y�`�>S�&%H � �@�k�����'���S��ێ[汪����wW&( Ek�>������.͎$H�	��'�(�8�
@9l��mJ��ȹ����	!�a�DX%:�^�	2����i�S|Q�%BkGkH���wq(����'dc0�gV�m�A�Wй=��25i��=�m(S���P�e�3E�_��Z��7H��Ct�
 K6��rWʉ- ������?1d��C�@XrÌ	?&z�k���wYJ�S@���ۘLl"L�ԥKۈ�*�����	<|�d��V��'���شr>`�V��^���`��uĆ�l���P%1�>q���'��iIs�'h2��џ,Q�7r���!�
ʐNN袃 5D�����"�D��c��)m7 "3.O��FzB�n3DAb!jôOB<܃3��?���'E��'yb$8B-N��"�'~���y7�M�&�cuʚIhDc�T 3-�X��IN�bYn���/|y��3"�|�o�y�*}��2�y�q*�3y��l��ޜ���dR�#������L>ņ�x֢Kb�	O>L�'b��?�Or� ���4퉖=J���;8�AR�_>�\B�ɼ#�J� L��4"��4GJ�%đ��'����0��j��M�,
�d�Ʈ.Ey<Q+��+H�����OF���O��;�?!����DH��(��t����)F���pfʹ]����1F?>�\�k'�'lOF}I�/D�YgM��`�,jf4d��꒔,������܌?m:I��I>������jZ����*�$��O|�d9ړ��'�N !�,2{��`<S�<��	�'/��fͯ7���f��0��y��>�)O��
��]}��'[�А�πRZ��Q& R�	��!��'j"�!e��'a�	�h+N�S��^#/����F �h2�쉯GA2(�2�ý+����I&�̹��.F%�l,j�'@�9��F�C� ��kZ�n����Ǔ2Q���t�'��1n�� w�LP�D�$6UZ�ҋy��'
$�˳�d�fxa�0�*��'��7�K�u1 ���OSS堬�"�>V�$�<I�M��A5���'��\>�R��
ԟ�*���13G�p��o��z�ퟜ�I�  �9��4������#��WՂ�s"�͏��)�N!}� ��(y ��A�-]��s�-�D �e�J~��&mY��P��2�Y��B��Իecb�'�7m�O&�?$k�+�c���/1����kd��'��V����C�p8��M�'��9*�����p����޴�?���i��k[4<�óC_�?���у ��듌?q�IR ���?����?�׿k����5tV����E�直Q��S�A�>�5��

��1�|&�|�l�nຐ"t�^�:����,"���X���#���W�q��'�$���c�VY�E�R��p�U�'"�ɭq�N�4�,�=їm� �T���N;b� ���m�<�F�E�?�i@W`[�$��\hQ �h~rA?�S�$V��3U&X�K��AX�G�	/����i0���j`��ǟ��I��@�	:�u'�'0�;���2���6KK��k	_�GT:�jC+��U� �FB5�O�L�5��^���m�?#$-Â*ƠKq����&'�O���7Q!e��T�͕+��q�Vt�"�'���'��I����?B����\���F鼹P!nO�<�"�_!]ߘ5�e��
x�X@���P̓��uy'G�:ꓥ?a��\�a�b�1�}H$ʴ�?A�Z�9����?��O^�|�&��*W�I���>A�mZ#4�G')$ l�S�#O�1q7���l�\�h�u?QѭʳTS�����s�[�N�I8�P9���Ob�$�<�c��bъ��'(�����p~̓��=��HS�}�v��a盺u�����	v<�i��`���48�H�����3YT��*�'��	,ƞY�O����|"�I��?IgH^��8�-ڈ@(���-�?��y�dE!� �.�S���*���'y��Ce�_)І�_�ft�@�O���S�\�^�$����I�#}�ꎗN�xs�m]3W�(1CQc��f��'��>U�	�h�
	��	�~�R�ԧ���0�Ɠ�% ��E`�Q!�T������HO� 1�����Y%W�V5�)�ĦU���<�I�kgbAUm��I����	��u��*
Lر*O�7t]Y�S1O��8��'��,*G, ZF�T�S 4��{�-����<���XO$��e-�C[�����<ܘ'\����S�g�'����AI� ���\��C�)� P���C�ܠP�l��������Z����n}P�&�N����8���x-�$8��?v�h�Iݟ�IƟ�^wV��'"�H�gG�x(Wܢ���R	C�̂#OD��4�Q�J�t��TC�u�� V�	�0!�тJ�:��hۑC,�40g� ���y:��'&�';��'*�O�a�.	-��q���s�B�"O�@+W.H ��Ӂ�Ra�P`D�d�x}��i>y;�ϩ!�B J���7�VqZd/:D����Y��5ؑ�ӑH~l {�6D��x�@V�S<d�K��̄1�^�(1g:D��Y�	+
�]k�I�*@ST,9D�4c�oV$ @���C�h�ay��8D��0`�_(v~<5pA�6lܙ�s 6D�Hڔ	Z�4��0aߑ
��A��6D����,`<��I] `��!��(D������>g	 I�)��t��IU 'D�ț���4����Y�d�($D�\���G����9��\�����"D�\"��1$Iu2uDC"lD��b�l%D��!��M��Xi�'p�Y@V� D� 0Eb�>s 51#�*�$Y�d�9D�@a����#�|���T�l�H-���)D�p`��>�`�; m�U���[��2D�X�U�C�Dp�Q��M�f��͐��2D��ᄅƷ|�>��D�K� ]��Zrh6D�4 ��N�}�2	�H2��H�3D� *��h�Xd{���1Ί9u*2D�� ���;Z�Y����~U���0D��1��L�g�@] �IŤgXI�4�"D��ꅨI�M QTK�.Dm�Պ�"4D�l�sdōjnBa���o|,��k0D�,BQ�
r*��(���-����,D�|��
�/o4����`��� e*D�HK�)�T ]sF�R��إ�)D��t�Q�v�ֈA��D6.��e��&D� ����r��P�G����Ub�2D���IN[Ґ)�sJ�\�8`/D�(�0��E��#'�F���,x�(D��iӭ�=��3s��i~�4�4D����C1`($aE)"l�|Xx�#3D�(�do��B/����^.��3p�$D����N�;py�-��a��h��ms!�!D���u��!n����O� z��)SQ	 D�`
��V��a�p�!m"��;1E>D�D���Ä.jRģVc�'`v�ӧ=D����bB�4S��q�EL.1n��$?D����Yp�x��y���i�e
$�y' 7�yp��Q:p�����`C��y"�ӊ1�x�9����U��D��S?�y7 Q4�� �O�n�QR`��yB���N�n��S%�Tx<%����yR��#㮉*3�ղҽ32�U��yR��6Gnޭ���v6^���C��y2`̝W2�p�U�@"Œ� 啱�ybl<,!�,B�ۊk� �˵n�"�yB�E	1cx�� ��c���2&"ʅ�yBgQ�4�(�`�&ۑ\�]ؕ'K;�yҠ�.FJ|Z�M�O�\U	_��y(M�?l�t"���@�ɹ�(G��y�(Y&��9be��Ѝ$+��yr�R5 :��FA�C���x��G�y�b�&T�{�DĮ?dP�Wϣ�yb��o��aI��	�I�&e�!��;�yN$F�3�U#F� �R��y
� ���3�O�g�<k��G12@��"O~E:d$FZ���K�O� ��H�"O��Iah�����w�@41�HD��"O�(H�A�D!"��e��O��tQ`"O�X�W/�./$=����k�t��t"O��)�P5>�$T�O�7���q"O�1Ru�W(��!�md|e�"O����#�!��,�TcvPA�"O��(�J�U[XQ��D�z@��[�>A"l�D��Ho9��i�?��rv�<#�L�|�T���ϊuj�����-����s�OM�L����|h�b�\��4AԌۄ	�N�"~nZ*�D4@C'�p� 5��3��>1�HE�<$@1��4Ě�S��B�jU��:��)����+yrߓI�dX�K0P��� ��Y��`��[���Z�+��S��$�a�G�-�Y·���L��l(]"��yǬ=D�xK����p����@����zRF;}�@�L=2]qu��/�v5�FP����~�����
T�<���8�H�h��ҵ*ߑCXa�s�ص$�ک��-���U�ֈ�}/�|	f��_��,O��z�-(�s����V�\PU*¬V�r������	�f�(��Sb=:����A�E�A�=�X��Bم+r�X��ÊŗPJ.]�D�S8�xkR�
e�t5��-�;��{�A��&��aSrGGc?�OԱ�?��t��k��4jj��C�J&C R!����frh�������O J�$�#+˘ȣ%>�Zu��Ò	��5��Z����\�~����H3A�V���Sސ�g�$-�}�%�
?p�2�i[`�� kPcO���'h�!iTk_�J������S�4�S�O�8c%��j<�qe��Ǝ��F��!r�Ȍ��g'���:��QCn~+8�1�`-#��D��=��y#'k ��1�#�_$��g22�Ce� ��9��FB�0V�lt`d_ 	��H1]w �	:!��F1�2'�W5��h�'����a3m�RHrQ��V��8���U 2 "F�Ƅ)'T����1l$���)Ψ���)B�Ȱ+ L�H���VD�>Do6�8�H�h@ "�Ȏ<!ń�A�n#ړM��!!J%PH)�;<x|�f�J�+�F@;���?&���O�Af.D���C�p��c
A�g?�5�>|�z�#☗rH1jQ�i�$0Q�3�ɦ)u$1 U���}��x�%��V�.�C�� �Fϖ}@���H�(r�f�I��<,tlؕL̴�#�OX�ڴ#�t��hCb�,��C�'m v+��8,͉�Eɕv�ny���! 7���Ǌ��xޔ]kK<Q��Y�<)���=�~r`��F��k�'r��4��c��~rHM!xY����A�^��	9�J@���4�:�7&��2��C�Oֶ�	�E2>�NO,m�
ЛD<Н��@:�{�p�d-4�p��3��6�teH��VBA�
֝9k��<�ƽy��iAG漫n�';}� Y�$!�9Yp(T�
��y�I>Yr,\H�OK��I�������&��a#\!a�.,:�yb+L!.-8` �*�`@�`�И'�v	�f��&�L!�� -Εp�4!���ێ}2C�gl��ja�-h��i�t���';�MH��IC��(à��}Y�P�rظT,�52�g�Lz ۓmU��p7G�7J�	Ӗ@��?�t�JrF��pp�@��@B��;��G�sR��'��hI����<k4٩��%qaj0ZT#E��yb��'jgX�B�A�&����rE�%,6�|�r�E	$���!�+��'��#�k�\��w&�y�Vhγp�L����а5X�q��7���c�
�B5(�V"oX9��a�~��c�8��i�'>��*P�B hd"��%扶o�acA�� ��L3w��"'`,�>�B�
Rl�B� �3�,p΂�/��T���	,�v�V�(���ӧO(:����a�^p`�V�,LO�"׭��F3D�1Ea���;�']�9+�K?�v�*ufK�sM� ӭ���D�3A��_7Uj ���)��X���@���-d!��C�8�A�)#z��ʣe���na2@��:T�P�r"�ά8R1OP�p&�ތx�&yx�4�):��[+����X� �P��'�D��"��,�@���X�\�:�٤'�X�x��<٠/�5Ux��tT�j͎t�q��̓>ER-2��>A�|�wfA5U⼄D|үY�A�vԙ#�̵/{�-��B��P���Xd	��TҒ1�࣋{y�i;!jݕt�XI!%	#I��鳓/���?I�������x��) ��9�>hI$��s}���b� Vxx��'瓶2�@9��O��C�|̓�޹j�mY�/@@�ɖ��G��q���fX�T�?E���D5�H���@Q�2rHIVC�A�NUAE��)��)��i>咖���e�杞dG<{���.O1���C-Q|���[;<�B���� H����c��d���T�'�hi
�*6�'44�p��Dh�j-K�$"<�AS>�DU�8�h��Cl(�zT�a�?�T����D�Q�C��8LЎ���-҈��i� X����hD�0�GefI!��!L$����9`����̧^�� �L�0�L��V�{H�}��?��?�����Q��=`�g�n̪��DdD��@ 6ҼD��@y���1��� Ԕ}KR�{�� �7_i���<@b@L��)� �,I�dC&w�v�a�A��,�5@D�ɴe��m����0鑗��F�M�����6�U���csÂ�ÈB䉲F��ɰ��Y#L�0X`D��z�d��-vL`@��R�(�)#KI�)rd�}Zt�R�t�0t�g��Y�$I�v��}�<9���|Zd ����r�lX��ώ�1ʣM����H��		���fhSp�n��D��J���T�C.J�"��-�.Ȉ���v�h�H�D�O�f��6ᒬH��9c��Fi��t�e�5S�rlZ�/_4f2�ʀ� �\����6犉#�6�ۓ':s�Td��:X��]cTe���	�)d~��"O�aL;8�:ɘs�ўD6F8�`�i���b۠��s�/��Q�(�Af�(�k�\�����	lD�x�"��N!�5B�DEI�mҶTO��K��Li�
X!pGD��lI�,��4Ε�BT?��2�d;����G��҈Z���(�z��קt"0���Yl�Z�,N�tP��̊Z��#�.C�u��P��L^'%�έ�ߓF�q�ś0�^��
L�8���<��\�?��ݹe�
�}pP�7�P��O����J�/P�9sU��]@8XS�'6�d��%c�\p�uc��S�si�6�X0R���ȈL�����)�<���ǡ�)\T9��l�<3��4�s"O��6GU8[;@��t�3 � )�PG�9m{D��1ݙW�8T�L���2OE��㟼���S���qT�J�3���C�*LO�9�u-ù�⍣D�M�g]\�)#ɦmm�����[#n�+�����M�R.�<:7���ɺr�Hag��j[^�#%�b��+\��X%�ݠT��)���,.�p�� ȸ�u���=\tw��6!D�124%�+�y��G��X�%� [L������P�r�M_�5�I�͔�n�,�B�C䒟<�Z�w[�`6F��
�x�)a� �1��'?�dB�/�+�Bt��˛�/��"pI7�9�!%���͘%���<���Ѝ\A���ԓWo9�$�@��$!��ͫg�N1�'���	��W%+@Z ��������'f2 ����K>:���#ɂ9z���y�/Ѳx����a*@�OU�(�̈́_J˖C,���A�'t4�&��}��7M	/ Z�� PM^1���O4���3?i��]�J9.$Ar,؏d�� 0��v�<ၤ9f������ʀ̊�Ѧ~��� �`A�i>.���I�j��g���)�KX(eF�ի�n>&�P,� C���Z/�!���:"�����6B�5H�`�!�ս!�^=B�Ɣ3 Kb�<A�ʍD��Y���0v�E�	�.m��C�0B�B�	�,'1I#��.Ű�cr�EI�8����	�Tr�fR�PG��OPK`gԷG8�����E�,)�5�Q"O,䊒F��
o���+R�\+T�[Q�Z�H�t٩��U�p>ѳ������V����#C�j���k'�0.�~��vS����l�3jv�d�>W�!�S"O,ݳv�D���<0U!M!2�av�$U6A�bp�����&��a�B9Otҥ2���?R	��"O6Ti����v��'�
�s�:<(�g[�&�h%�<+��<�R�Άv�X\ '�O(P_�1�TFe�<�hQ�T�� ��K�!SU�5���i�<qp搼�yq�@�
%��w(Bi�<)B&[OP��O��$^<B�J�I�<)�N�S� "Ąu
(3e�z�<aeI�4��q�E߂=�0��*�o�<�5�ώ	�VM3�CQ�6)PX�g�\i�<��(P����B�:a��jš P�<�6*J�t@<��%�H�0�atv�<ٖ@!�29����1T���c	o�<�$�Y�9���c�,1%�q���`�<��#cI�1)�D�'=�r���)XY�<��Γ$�n��ώ�4���K&�S`�<ar�P��vd�� [�
�� 4�B�<	�M� kO��(��H�
�svc�@�<ѣ�P($�b��"aғD ���{�<9E�̑
�px�-Г6`�	!�,T^�<9��s~�/Y�:!��̈́��B䉝V����Ч)>�l��H�a��B�)� ��#`���Q��9�� @/%輪W"OF�S!@�FnJ�f�Ɔl��"O����e-�K�'�]��"Ob�2A�Y�]6z�
h��S���t"O����G^�C�,�tǍ wXR��`"O�@zj
j���¤8C�T��"O��Ұٟ2�Ƚ��C�;=�"O��!C�Wm6aR3C[<= ����"OdQ��-�'���qL��7/b�b�"O��Ђ�]�6,���E��bs
�J�"O�H����hQ2(Sԅ�䖪)�f"O�zҌԉ'����+-v�6��D"OB�S�$@�nH4��+�Z[��;#"O�����;n\%jĈQ�uf���"O`�D� ��ɣ�0K~|��`"O�R��09zBe8�G�S�*xj�"O���O&}�%�FeX()R���"O�����>T? ք�,
�v\�t"O��A��6��a"%�$����"OR�c�Se�,I��T�V�ll��"Oxp�kQ?^��Pp]}ڼ�y�"Or ;��U�e�%�߬|�\tP�"O"D0��eP��2��YƠ�S"Oݳe����<��o���z���"O�QC����
�x���D$f{�!�t"O|�5&��\W�!p#d��;��Ua"O��[�#n�~����:��lCe"O�P�J�d��P�R�_�\ �"O*�xX���*R<y&~ �"O�����W�쩃�hD�m>
��"O4�p�P2>]��3�}��I�"OR�!�lY�$۬�6��:�� �"O��񅫎�6~�i�!�D�6>q@B"OF��ń]�J���ɤ�J�&�܅��"O�hA���r_*��@ Px�� F"ORD�G/�<P>��� hZɛ�"OXHy� дHaO�4F�h�"O<�p %�$%ʹȑ�d\F�-��"O 偅���D�95��-�Up�'�!9�Q�W��!V�e�\x�'��\+��V�\І�VY	0���'7�5��FZ`�_.Tj|@
�'Q����e=3�H{PN�\�C
�'1L��5��r~�H`FB�[�����'N]P$た\�
0Ii�P��b�'��Ñ�F2|1gН1<�|�+O6���J�!�:�`��<dKUꛐR�!�A_��Ԉ�.�.������6,�!�$]�ty88��N;|����ʧ�!�d�4wYhIaD[7?>����3�!���L�d��4�C( �H�ek�]�!�dB�M� �
S<�Ы�* !���I��	�J��)+�(p�I�F=!��<R��u� H�l�=(3h�J!����q�6+#m�� ؠ䙏x!�$F"*�D�b����N�\i���Y2�!��bI8�IeL��N�l�Z�� �!��9��@0C)F�:� o�!�$��:�@�P"�_~5" ���O�!򤑂J�b��&+	�q�nP��Щ�!��R���!e�c�88JdGQ!M!���G@^M������(�H�*g�!�DD�E"��	�nzLtP�(�Y'!�D�P��5��ŉ�bg�Ⱥ��L!�� 0�ui�"z !��Ε�{>EI�"O�P�0���;3&H3V��.xul���"O�Ds��M�4�Z٨�N��ogT|��"OȘ��.H��|���,Ua:���"OLy����k01�`���DU�q��"O,-��"F<c��܈�d�>'�J�R"O����
)�1�c-R�9� H�@"O�]�k��i�~�ƍ��W�����"O�XQ���������R����"O8����J8t��
X�xz��D"O`��bO	S�t@U'"rfV�R"O��S�aL� 2�E�.xF�e�"O0`�Ǐ�.q]�rC
SH`=B�"O�\#0 ��:�*����E�>4���L���X�ue��jp&#��H����!�!�䗱8ɪ�c�.\p���1 	9!�$
�B&9���N�R�� �0e)!��;N=}���8@n2%R��O5U!�$O@y���(Z-_�arUa�8^��φ �|��ߩ~S�K��1�B��>ctY�흊4��M��"ȩ'Y�B䉒_>�[��P5%���@s(�q	�B�	%Q���F��	H�-��%-/�B䉣P��LEa��Kל%sՊ�q+dB�3;V�S4&��*LA$��PaC�ɳ$R��? �н�V�R�	��B�&P,K`�ťM(�!kŔ�x�B�	�c%`b%�=`z��rER�Qk�B�I�D�b0�@�T�2tȲ�L�{��B�	�
��xQ�l��"�
��J���HB�I5h�n����2r�AZ��_,r�C�ɻ�B��w��>,K�qQA�&�B�	�#���q�Ħo!���v�T6	�fB�4i��}0e�N7/�NI2��p1C�IMF� t/�W@:��4��,�B䉒(���C@ͨj��0z�_5w<>C�	�j���0~�Ĩ���mp�C�i�j"�C�B���a����"Ї�O�&�3Ɗ;}�@���"�'}�ȓ�LBT�ڽ\��c�(��(fLB�ɏ<��U"�o��{���b!Ϗ�!-lB�I9GN̬8td]�h�	é41��B䉨�f���Y�+�1q@�B$GT�=�
Ó&�m��nПK̸t
�ʌ�vR0�ȓE_p��4�d	�*%�C�	�g� �r+��n��T��nl��8�I ep���ԽbW����#7��B�d��b�K�"m���P-7`.B䉲����w�ɝ>��"�� �Pa���E{J?�C�m�w��*4�]���%3��&D�8���G�mʠ�'�6y�)Q�M%D�,h���(��E@pJ׌:1~MV�&D�@�U* ������2!�09�+�>.O"�=%>�bc%���)I�酴J�8��Ĥ �O��|�,e��[�m���H��L l4��9oT5�W�1c��Z�U"u4݅�2���tI�q-�8(ק��( 9�ȓF���{��+���i_�h��чȓ�x-AAH��YK���.U�s�z-��U}֘)"��?@��Af��%y����H� 	 �,�-9}L�k&*��	F8��s������a��\s �./
���	I��!0�
={��58 !��X�C�ɺ$Ӣ�r�D�|Ҭ<��n��!�� �l��K!uG�T(�+эZ�l-��"O�j扂�qZ���L�_�2�K'"Oh�a�ʨpP�)�K��_Z1yf"O �p���%b`�,0*R��ku"O�@��ŕW�laz�!�0(ЈC"O֌��ѓ^퀍K�Fղ"� �"O��Xq�# w���ħ�Ȕh"O�)!�.��0��`PC#�� �"O�`��h�J@��
#-��w�L���"OV,�v���|1�L��&!a6"O�1`"���Mf�H P,��9���۰"O�0K�N�9`�v����!p�X�x�"O
�)�`�Ahi@lB>5��S"Oz�p&9��tJ%�YS���X"OL1���/ I�%Y��Y�B���"O�A�g�m0<���dt�|��"O��* MЂ�>�!@� 9쥢�"O�hXS�D1rO���S��a�x�b"O�
P؛��c#��T����"O��٠�"̬Y����R�F��'_^���`;&Uh�L �xҪ��
�'�����ϗ5��� ��2~�p��
�'�0��e@ MP-����tj��	�'��ɹ�A#�`���h9����':�%*�!�g.�:�@�6�q�O����T����j�	q����C��h!�3�TE#'LH4	���a�;ng!��_�/|���.ې<��]�&��:0!�Dӡp}[a��NHtay��L4K!�T=LMYԏ��<H�	kE�O�!�^�0�8e#K,N<�M2d���!�$�:�����k�H�0�07�B�K�!�d�<됉p0I4���R��ĸ��yR�]� ��r�C�}��%��ğl�<�v �	��ɐ��?.��a)�H�`�<)�C]M6�Z0'�$Jy�Q���N_�<��!l��V샫c���0Q)_Z�<��ș#T��q�b�}`b��]U�<!W�t�ZAAg��&e��|ȅ��V�<�%�\�m�"M�@�K�g^���'�U�<qs��#k��#(G�W�&5b��]�<�RK��"�^A�QB�n�V$jD�[�<�5��q�X��5���?�X��M�<F�J�!4 �G�H St0a�GEH�<Q� 7��@�wc��T��Q o�@�<�7�$���ǙQ����a@�hF�C䉸K�����W�>�v(R�S��y��+&���M(l��(�y���K3�(���J�XI��c�.�y���������$�=R�4��	=�y� �0#�
�as�ة����T��y�K[�YL�"�<L�谦)Y�y��b��ܪ����U0F���y�gZ&�=�惚�D���c/�y&�-j��z��z�L8!��В�yR�аh�Z�������^2�y"��LR��ǎ��<���c�V��y.�9Q�7K�:.�^�[F�ҹ�y2�������a���"�Ҹ��G��y"�Ľ&�H��$lC��zE2aHS�y�f��/H�`���M�ژ ġ.�y�I�/FZ �w�N$\ږ%Rd"�y�	�l��S��_f�֌C�y�L\��"���WZ*�+�$N/�y
� rPaա�=X���z�
?�Ҁ"�"Oҭ�4,ƞ8����C�l�.�"O(-��Z�l��+6��G+�XiC"O�h#��~�:V�S�<x�`�"O�Y�qmQ�,=B@�IY�fe|U�"O��!@+�2.�)�I�ad�{u"OP�(g�]!P1`u*C@&<8=Ȕ"OT� !��S�p� s"ȵNr�("Ob��+ۋ&٨E��+�$]騬��"O| ��BCw��@�N2	����"O��Qi�)�h;���y;>���"OΩX�P�;�8R�M0�U��"O�u�BQ7a�u�K"U�*b"O��B�[��}�R �-Z Z�"Ovu)�K��E�j@a�m!(l�у"O&��f"��L�LH�ČNx��"�"OL���,� Z]<�1�lG�E�5"O|1�ۆv��R�$����"O��&c�>%��s�_�p�(F"O`H8�ʖ]j1��D^�J�� "Oz-h���u�ISf�IR����"O���f�+[6�x��n���9C�"O�B��E8^��<x��r"OLH	�DN/R�&��ӂ�G��@�"OT1h��"�0) �݅�^�x"O�TRp��j�3�I��2iCs"O��+gh^8���f� k���s�"Ob	(��Ce�\I��\/ v �"OU�CN�W�^� ��/v��}�@"O��dhS�4?��h��F<�|��"O\���Zt`,rWв;�F��"O,�a�g��D�����p�dc�"OT��ǚ1&7��p �Ńtq��"O.�#��+�6��"�9{s��"ObH#`��!��x�!�ƢD�6 ��"OPb�
"9��p�������"O����i%��!��hԣ ���R"O|Ջj�0�aG˓~ �Z�"O�,��j	!Hx� �E�!{��\٧"O~��� ��0=�P��	)p���s"O.9�W��?�H��Ղбi U�$"O�db���+S��Yu�ȋa��Q�"O�L��GZ�O���R���MG�`��"OJ�v�U�!����#"K�U�j�"O���V��;1�[B"�2TLݚc"O ��$��8��|k4�$0J�y{�"O���Ԭ̋4v|P����uF�5P"O�Q�FM�5
h�m$!9���"OTY�:3r�#�
�k�D�0f"Oج�f��;��Q�Z	G�lq0"O*Q�rdW�dT*��@w���"O
��!�[���䆗*,j���"O���j�l��I5#�6U^\��"O�d�W�[�k��H1p���X|� Cg"O����g��B�0`ӏQOez���"O�h�$bJ8`��y ���-^�4b"O$���l&`��l]�Ma��{D"O���ŀi��tx6ldS`���"O���� UC	~j5��;4��R'"OZ�K!J	y_�dQ�I�T��I[v"OpĚɋ=^�j��%���~����"O@�"�Z��lr͜�c��%[�"O� 3��ޒ\`�E� l^]��9p�"OE� ��5X !�Qʒ�6�z�R@"O� T]�a�k�^-��&\�8���V"O�X�h�$S朒5�?�\��"OL�[ǀ7in��ac�Oh�k�"OtT��˝�|o|��U�U� ��"O:���Pr�&B�X�&��v"OZ�XΒ�?f�*�+s����"Ol�{eρ�)˺�sF�ϔS�2!��"O���Z�p�d�؁oWX�>x��"Opi�F#�|�\x�dP�F�T�s�"O|(JdaV+Y��0��)g||��"O�Y�R��JUp']�4ZZ|K�"O`:We@�b�ec�-d3r�u"O|�j�W�QR(]�R�f0YP�"O.���c�;Ld�9�d�O�]���"O�`�̿^I��hD-�p��Ȋ�"O� �W�5a�"}c�*ۭ�*$�v"O$b@�ڨb[��q���U����t"OP$�c&O</X1�'W�${�d#�"O\��t!W� ߄)i5,�4&מ��G"O �#J�we�����
�#$=z�"Ob�����3t�|Bi��@��D �"O�x��\0"e���+���"O�|J���$zҔћҡF<i<D"Od$�7 ʴE�rx�^pR2l"Oz��΄F�]zv/�@���� "O�D{0�87[>8CT���p�0��"O� ���ߢzN��P�W1P��"O�P3�Ο>oB)�E�ʺ@�@<P"O�0fh�5�JC��P��>�b"OTeK�Z���)����jt`�"O]��ݒ�fr�-ɪM�Y��"O���a��?�6�X�L�J�>��s"Ovmh�OC�SV��U�Z�A��%�y�լ9�±��hģN�X�Q�߬�y�\�+΅�C(N�|�n2e��'��i�r��%�<��O�#Y"j��
�'���9���+x�@D#�*@��Ѩ�'���ݓeS���Z?+Hԉ�'i�U�c�ܢZ���
�h�;\,���'���VE	�S���E`��8O� @�'�*h��� 6�����5*^ѐ�'f�M"��������w/M�XR��i�'3,���-�2~
LhDŐ]I���'���BQ�����H.QY���I�'0�e��I!y L�S�\�O��'H��V
ގ���@Ǟ�u�0���'ݠXC�$O;:5Ps!ȋ�8��e��' �����UʆdS4fЫY�|(9�'|���b�Ows�,��Y�M���q
�'�R�BE	�)�TJ!L��m�1S
�'0�Cc�%Q�ع@)V��M �'������G��ቀ/O�NYX���'$~y����k8�s��A��ih�'�d����r�hx��3>�}��'�FTCd�/ZV�jG�M(-n���'�<`J���i�>xA+�*z
�!�'<LQ���?{:�Ѩ����$wL��'����%�/�0�
�H!�hm��'�:h��L6\���ɡ�Q�?��� �'����ٶ71�b��<�T�
�'�B*�@aX���7� ��
�'o
p�E(��|�5OT8'���	�'K� #4NL $�l|���-�F]��'n� A�Ӊd��ݛ�%?_�l����� 𙡂�0��Da��R�r@q�"O��;�䇁��� �#���vDk6"O�t���g�@ �ԃ�!��a�e"O�`#E�$̙3���;���"OLa��Ie��� � �3k�4�ٴ"O.���^�MJKQ:j�XbE�4�yλ��#�� ]���)��� �y����m�G�D�N���%�؊�y��,O�t�bg	�L���,�2�y���g1�0	�ȑ�7���1CM�;�y§�=|���SJ�3{O��ӣOſ�y���T�d�U���W�i�ᐲ�y"��p�TX���%q-�)kfZ/�yQ%Vv8�1��N�dZ|a;����y"�%_ ��R��k����vfF��y�,�$��VJj.� V�Y�y���2bz�VgH\�)UFץ�y�� �q���`��hBDoŷ�y��_�u,F�@��G�Y/���
1�y�lU�2����0U$Ԁ�	��y"�;wq�����S8E�`�9�G�-�y�_
2�ր��댁l�D��!���hO\��3Q��@���8����F:џ�F���0R\Z����R��� �����hOq�ܘs�b��S#�d��[F �j�"Ola�W*|�=HE��)g�6I��"O.P&K�-�$��Ą˙s�j���"O�Ġ�m!�^��EiOYpTi�"Ot�@C�7U�:U[(�ak�y�U�'��Ⱥ����[nx��Ve	�ܬ��p�)D�x"@���6@+㣈�)u�б�-D��0�b�NdNi�Ҫ�'��xk�)ړ�0<!J���d�������!z�R�<1P �;*:���E L���qd�P�<��LȊV�����l8�9��P�<d��i����UM�I�fe�t�I�<�-8tC.0Q0Bԁ+����G�<1 �K�j��9A���;sL�+�j�p�'�ax��.OoD��Ƀ$o�8!:�#����<���G�>R��� ��6��0�ΚZ!����V0xbK�8� -�v����!��$:AD�� �h:�k�"�!m!�䗴v ��jSoB�s��!��X�Z��'�ў�>��1pw�x�H\9`��@�Q#9��7�SܧhL ��ԧ�l56ZF���g�H#��͟d��5Q�ϛ%��=E{��OȂy� �;e32�ڞ��y0M>�,c��`�Ӎ-��-�gO�V~Іȓ`X��'6��}���"?~!�ȓF�r��%�"jO� S��ڟj�
D��S��xĸP,��6��D2�k����C��$��y��;j�B�j����x��C�I#n���Y����|v̈1����?����) ?��+b[�KED���I�<����;��Y�4�{r�mS��K�<Y`O��X `�YЦ$SPnũQ�F�<�2��{KNA����0I  �m�~�<OխC�*���[�K׀�#3��}�<��UvF��$�^ AmH;C��A��0=A`� �JlB�9# _�O/���U�V{�<��q��x�l�9jv��P��z�����O0�$��N���
�nU�����'���S�%�g�p���<�(��' RYl��;<��B�Ԟ.k�%���� <��b׎ }(�(�Ý�F��q�S������|�&��CO��P+|��"A�-6�C�IN)&��P��6"��5�t�O��x����x�'�d�D��l�Q�S+�x ���x�
��z�u �R9 5r"F
�y��Ăr��9�M��*����'���y��]�wRIaf!�r�0DF2�y�i-�`jDjq�e�R��y�ƅ;Y�|������ 3��8��'Gaz� 	y��%���4 ��KAn��y�A�� :�&Ʈ) y��!9�y$�"���5���'Bz�#P썋�y2m@�B*J�C�3{x��4��yr-C T�Xӱ�Ψ�����y�g��)����e�_>o�0pbC���y�J:�0�3��LQ����T����0>1nR38���ѣݥ?N��R-]d�Ik�'����<aD��Isuj�!A8���[a�<�V��v������on`AkA�x�<�T�1|�
8�T�:K�R\�C��?J\�YB$��Q����E՟B]�C����b3C�:Dp�eC��Q� �C��/pu���!��*�q�^1Tn૎"�)��lN֎�"���#WX^B&�Y��y򏀰<�j�S�lQ#Kn<U���D0�y⏇=}�
����Ќ>� �����%�y�E��ZĴ�#me� ��װ�y���eH��t �"U}��hQ*���hOr���@+[���kakŭ(��TK�
��x~!�U,v���%	/+��hC�nF�)�!��I#�J����@����#��2O{!�DǕp	�£K�El�}�`�MI!��kH����٘Kh��Ӕ�Z!a�!�ċ'@�<}R$J3�,������!��_z��Tb�
|8�:3*���!��W�b����I�p|-Q�
��!��\C,�|yvN�U���cB�7��O����xg*Uh��:E���O�${!�đa[J�;��@�%#TJ���S!��@6��tI.��[p|:��"C�!�64�jL[��I�h�1ɖ�!���)�`Pg�_�"9H�'O�!��5I��x���v�8�c��r�'Vў�>��>Y�a��6UʚT�§8�$*�S�'�Ƒ��L��^A �Θ�o �t��	b~R�.���.��җ\ @�J��
�'��#G�� p��f0��	�'k��ImQ�=�aS��D�2<��x	�'E���/Xǂ,s��#�����'�`�0����У H#ZBQ�I>������1?v�k� K�vXF@Ƃ��+2!�G+x��z���
{AȘ�C A�,!�D�!z$�5�ƤKV���<L�!�J!�����%��DK���A�
|q!��U`�d��@j�?\B�P���!�Đ7v^T�WJ՘!Br�h�/G�!�I�Qi�焦j�lhq歁$.!����4@���V��)YWBƍ<!��L��1��Ց:{䍑�Ւh�!�C�0���t/X�Wu ��Y�!�DĚN���nmb�SO	�!�$	�gy���g��`�`���z!��Ta $��OE�p�N�BUI@��!�$Q�e�p1�g�����a�`)ȣXo!�� "�ʎM`h��lDj��@�"O��Y�LN90#Z(Ɂ,�)���Is"OZ����IUR�È�;?�d �b"O��Z�fQ�3�j�����k����B"O�
6���1����0�W8�T�p�"O\��3C/w�dʄ-·v�>�1�"O����.��P��A��'��'��6B׆��􆛜_��@�ȪB�!�Ĉ�G]�rdB�
����흄*�!��)g��I��D�������&�.�!�� �)f`�i�m�>w��mC�LO�!�G3� L�g��J����i�N�!�K2F���-�0�Rq�o��T�'�a|�E�'�<���'X92 �j�P��?�(OL���P� ��`i�iA�X
��6d�o!򄘔V3��hs���y
F��6B��3|!��D_�\J��Fz^�����Mx!�d��Y��u�vJJ�
����!��SPnm�En�0��-�6P:�!��j�$D����6�r R�횎b�џ�F��M��2��p-�<O��v�B:�y"��>��ip�+��E$4k%@՘�y'ԹBo���g��<�P�)�
ŷ�yB-Ln�R�C��A-k��TnK��y2#����!c(  ��<�'
��y"f�2-|����$�Pˆo���y�e���҉�1�Ѽ"�As����y�	ՇjR��#�#=�ƍ��ɨ��<���D4�\@���#�V�X��ǚ*F!�DV*L��0��RF�0S��,[+�y��	� JmX�&�WHf��*]*"B�I4�e�����iX(H���+'B�C��6q��qm�c����va~C��1R@��A�����p��OE��h�=��'���eZ�u|�[��Zܰ�ȓYa�S��>�h�c�FIa�Zȅȓt�>9su�B�m���5� �r�4���鶨��F�A]]��,��F��ȓ_ЮL��	\t0ؖ��'𮹆ȓc�l��3,����[@�A�Ky�!�ȓ7=��IE	j���EdF�%�0}�ȓ��-�rd�(�X��s��=�DX�ȓ���h�G����cs�<i�x����T�f�F�T�����6<N��d&^���#�����*s����ȓaP���2��9���7����qզt���c �#6NM�Q`v���$����m��镎�3����ȓT%��`�8r2s��W��%$��G{���M�v"8�;�\�>-��b�X�y���V���<x��T���y"F�T��z�㌮~�t	�$�E��y�&S�#( ���B���tɇ)�y�j]���
��;����AG(j�)��#%|LR#�϶5n��&K��j�|��ȓ!������Ի)�: ��q,XY�<�ǌ�0���@P��y�ҋ�T�<1��S�F ^�䁛�FsМ3b��w�<���߄mP��1�.F������p�I}���Oܚ���ɗ?��´�:�pQ
�'<z���Ƃ�Ϯ�Aw�^���$�
�'��5R��8.+���(� �ک�	�'|` ҖGр�,֯.�d�I>y�z^�I�V žDz��RfEI:l�p���S�? ���
 9�FPk��l3����"O�������#]t=�w�]"D!}��"O��&֞�(���Μ6n�ű�"O��Ђ���v��(����c\D�""O�Qc
$T^|X)w ��E�x���"O& Z�/߹')SRA�"6T�p�"OU��+L�oB�(���Q��"O�ɓ�%��(���!�0|����G�'����ʱ�iY�}����Y7T\B�ɵG�J�(���4����[	2B��7
�`��E�$O�q�%n�����0?��Iו6�z�pUbY1|�:�*����<a@KZ!�&���
.O�Z��v��~�<�Uo��B�(t�"��	��[cN�}�<"'V3{Ĕ�J�/=M�Лg�a�<�5�& ��l:�l͹}�l����`�<��Ŗ��!��H=�2��І�R�<9G[0)���ql�UmyfKAP�<�Ч��@r���	�B@��NZK�<!�@���䀐��	Yj�@D%�]�<!G�	y'���BgQ:�F!�*�n�<QBF,�.�el����C &�l�<AA*�,�j�`�/c�l�K2�l�<�aF#����G�"{�.���͈k�<a���@��"6���+�0����j�<��ܤ[P�J@����D��e�<�#L��M�����DЬ7�� ���`�<�BE!l���#Q�Lޒ����Y�<a���3h��c�G�-Z郔'�Y�<y��3M�!�c� OA����U�<���*��p���oV���N�<��˝9_C�ة�X�nI�y9%�M�<i�@�s�^�I�*��9$�MG�<�o[�r�,�@d�d�T@Q�Hn�<9�.��E���i0 Ô~V}	$�Rm�<��F]�S��H�sĜ;E ��*&̚k��hO�':�!J���;l��g�eI�ȓ�M`Ʀ�)�(@T��!�r	��K��|��k�h�I��Ɇ�D ؠ�ȓDI�E�J�ʅJ
��!��|�<�V�ι\�p���7�ؔYâv�<�w#�;Jz1��.4ROd�I�]r�<�+ۊ`"�=化�Rg�:3I�F�<I0b�8.�1!���N�����E�<���Ő՘��D���:p��DC�	�F��-b��ڢ,v�UkEOW�(L�B䉘?������i<����V;,e*C��	h�P�7��D~UkQđ�N@ C�'��哳���/*�T8���2:w���d$?��-^�	E�l��}��	���t�<�K�
vŎ�cal@���Pƨq�<�&��?>w�t�삁W��`�)o�<���M�w�l��Ũ(?�J֮]A�<��K�z���xg" 9JV� R�<a���v�He�!
9ȼi⧛K�<1؛x���᪛!X��a���k�<�m���(	 ���!�Fi�<) �¿�\���--�xi��Ky�<��0pkH	�*D���bNL@�<iEK�� 6<8��R#p��J�I�d�<�R�P�V�~�4�� 8_��R-a�<)ck�X}h(�6�0��X
VT�<��a20�mb��:�
�.�S�<90�3eD���U5t�����Ux�`Fx
� �)�W�ϓ{?D��`�݅)ٸHW"Oj���L6_&� WC��*�vtI"Obe���y�� ����q��jC"O�Y����Аj�D~�t���.�S�)�b�6{�Ԯ8���G[�{=!��-v'��i�� ���1%��5O!�dߟH�
�A����[fEL2!�$� �$0�ƃ�:�t��d�!��Ob�=���ukƢڨQ�>Ts"��4_\V<�"O,=k-�T��d!	A�W�!k3"O��C�B��E�g�;@�~���"O�����H����MJ�"�SC"O�)%���W��|�7FE#��RD"O��D��[��� ���k��@�F�z>)��`R�r�
P�r�_�i'����Ĺ<�+O ��7�&�J�bOC L@a��p�8��"O`1ƃJ�E��x°�U�<n�b"OJ���DD$���&�/Hk�,��"O����
��\�-����f��KG"OBI
�7v �M�񯙿
c�mb�"OTP%��
�����JK�h1"O� qwjİ&r�Vj_��
�����Oأ=�'X�x�0ԉʌb��Ԛ%H�6d�L��Pa~U��J�?��zχ2M���ȓ%��e��'��Y��P�߮3f8؆�?�\��bʄhGN'G�D�ȓ\~��$$:�y�Q�D>\`�ȓu�@P�"h	�{���3�J���l�ȓ�T�a�׏S�TY�んu. �ȓ��M+3 �-/��MC�ꀕ;���ȓ/�2��������sEm�i�✄ȓM�e�T朅1D,AS �%v����ȓ4�4�����0q�+��!=X�لȓՂW\�!��=�� �<O�x�P"OLa@ ������`ƅS? D��"O$�@�HZ�0+��-(��"O�qb�/$�vD�&����D8�"OX��U	��E�.���
�����"O&�KtC��u��(q���z>��E"O`�{�����ʅk��g�P�"O1��M�c�N����7-hL<�'"O)@r%LY��p2 'ϖM]���q"Ov���C��O�D�[��P+LS�dI2"O�|�!� ]s��y"*�%�>��"OJ�Y�S~�X�`@#G]��0��'��	�6�����Q+bp�$L�4C�	:�v�bi[�W������FdC�I4_��@����)hX��.O�DB�	1#_�ѩ����J� �B?H�8B��*.��eR�b�r����f��(�"B�	+Xk q���ڷo!�B�ɚ}o`ȊW��(�İ�$�\RivB�	A<z����	 '��d,��O�C�	O�8����՛D[�FF�`��C���%���{%�8�|��"O��O��a@FXaB�P��p= �"O:�r�Г:8�z�M�;��ʲ"OL���k���Z���S�;�HH t"O`�cb,U{JQ1��h~@QQ�"O�� 4ĝ[�q�L�k��c"O�mj�̕
N�ՠ�JH�,�J�Jd"O6��s�]�|�:��ށ�tt`�"O�@�TH�02�IuGK�N�z�"OT@hb!�4'��M*�-�Qj�H�"O�  �r@�P=�|��5Ɯ�S{��a�"OH��古P�,�4@]�A�da"O>�HD�c�u��Wx����"O�iX&@��	�غ%,C�Bd�'"O��(�Œ.�@����1+���Z�"O`P闇 ��/�/�TY�"O��X���E��̈:�.Q�"Oȵ�0C�7�6AF��l.��(C"O��!g(�M�6��!h��H�1"O8QѓҒy�L ���Һe�Җ0�y�ŝ�b�B82gb�	@hZ������y2�I�o��EI�ď.Mdc���y�%Od�}Ycˈ%��DQ0���y"E��5�0=hu#�O	�tSd$���y�۴>w�M�F�E�vh�S.״�y��?w'�4:�i��:��8��)^�yB�,{�`	�$̎�1��$��f��yRG�#��L��$�te�ä�����!�OL�H�%��T�Z�:�`G2pq^���"O����K:�$�QW�Ę`"%p1"OB���u��X:�-E�NL�$��"O~\h@�4F�t��FT� V5�"O"�@��%%T�Eo
�U��'|�cF�D�[ ��k�	�R����'5d``��uQ� ǂЌF��)�'v��JU����&Ը���'�R��
�' <��SF���(֫P�1B�
�'.��7�(O~T�ȥ��*+�L8)	�'���*pȉ�.��Aش`� p�h�	�'? [��,I�f��qX�� @	�'�l�эNL����AĠt���'�He��C@q�3Kքp�R���'�H�3�/�-,�}�[�lY�-y
�'�X�h� ø�����Nxr	p��y�@��<ҕ�C�=*���[aDI��?��'���F����,���Ƙ
L�0��'�Z����K�_~�XYQ���|Q0b�'S��)Y�?��e��,=�NA�'�p8�I14������*�T���'qx�Q�Um��H@�E��� u0�':���eV�Xࠨ�b	�(1��'(f�2��FĂ5zu��*R|f44"O�����;tV�z�HL�I��"OH��!IK0��	S�N0.<:�I�"O�(Y	ͭO\�3��G�rz���"O�|���ÆcZV<2�D%\�H���"O�y��@M?u�]�t�+}.�˂"O�2��R�"�X��vbI�s��Z�"O���5�������DBk��R���D6�O �;�Eu;B\�g��G��a�1"O��y�HW�dU�e�4%�����'�p�e*W*��B�D�V�9�'^~d���<�=�1FN�B�y�L�edPi�A�;�ވ:��P
�y�	T�M�
����N�:c���Q&�y��?��!�i��+��I"�4��'Jaz�(P�}� ��eω#�xs����y���Z�B�D�i��lZ�(G+�yr.�.p�v #W$װY�R�3c�O��y� Ҥ1��q�P�Ь(ب�r�c6�yB�S�efACǉ�P�l(����y���B��4Q�HH�H�ƭK��ݫ�yjkh�� ^u�x�0J�y�U;��%�2g��ӇF���y
� �U)��-wy���T����"O\
E�6*���I�*�>[e�U��"O�X!6LЁJ�&������{"Ov	�Fg~F����A;;�����"O"�[��?S����&I�]'��"O�hI�R����bfF�l� Bd"OP�C�\�&q�h�#U�z�Q"O�5z�/�0{f���fc�<-�ꍂ"Op�
�G% nd�#T85[��4"Or(��ʓ@� ,٠a@I����r"O����#�;Q��x�31-����S"O(��Aa�q��mT����o"O���#סK�^`�&cD9%�� $"O\�(wI�2J�xl���O�b�C"O��B"-u#J�
u�L�L���1W"OL�[�O9�lڒA�C��0��"O���.L1SنB ��y�D�Ä"O�E+���.n�T �a^��b@#"O���M��z$�����8q�D���"O�!�DL�}���R�-
�>���˦"O�@1VeE�7(j�����/;��"O>���l�Τ�����$<h7"OM�ӊ��25��:�U5��D��"OH	�rlF+g�x���?Qڌ��""O"p�Eꑍo�P%��aײX]d���"O�V���/�Ea��@X�B�"O��R㩋� � 8�).,-��5"O� �d��0r 1�Ph�$^$L�"O��p�I�&�v$�I��`��E��"O��*1�\�
���*y�z�cU"O��fF�i9�ybP���2����"O�����e�4�+�^����c�"O� 1�Ō
<�P��DUx��+"O��bV�DrB�1��)�9y҂ �"O�̪uk���I���&#f�dp"OL(��nS<j@+d'�4����"O2�93��o���p�����5;�"OnT �L�d���W#���W��_�<�HS�"�9<�E �-�S�<��=>҈4���܃DЮ9Xc'Q�<9�n�$w�$@�T�CV`3�^d�<YS�bj��1��.:��T��G_�<)��X+[�ro�)-����!�B�<���+�e{�ʋ#}�KUHOi�<�`�?30Kd�
�xt��(i�<yf�Q<`�ѧ�P(~7td��K�<g#�?b�H������ � �-�]x�8�'���"c��5�
1�`׳[�|��
�'ۮ��D�'L��r@M�6F1
��	�'s�p���Y75��h�į@�8z�z
�'M��D`�+c,�aHܧ4h
�'6R亳e0$����\t����';>�$S�Y��A��.<u�BP��'|<)�e'J5g�n�2�Q�j[b 

�'�*������֠��D���&��
�'��*�c����K���c%Д3
�'����g�,-�QfGA7' *
�'2�!pV<H��9���	v;	�'\�9k�A�6�.y{5�W&����'���A�?&�$49�ۚ���'�(��������;���'���	eU�f������-��"O��3F�V$dn�ȦCΫ\n�#q"OZx��'�z"�?\�@�"O� �x��S�Mt�R(��j��D2"O����Ι.w;Z	���(~V4�W"OB)r�gM}�FQY��S� VR�X�"Ob�xŇ��b�����D�Dd@*�O`�T��G�6A1U��,^�:�xT��OPB���&��PփRA��m^�C��4x2%RP_�'�����2�JC�IQO*xQ��:����d�~4ZB�I�k�(��o"$i�AӦ!��R�<B��&E�|pb��T�m�&a2A�+ �&B�ɋw����^� 
%�U�$-0B�I�~�RA�P��%Rl.��ՊJ��<�&�D{���+�����g�Z�1��,�C���yo�����j�"�p�3�Q)�y��?nb�hEc�#h���B�W��y�삽R�� &B�;a�~�9�bݘ�y���ff��W���*�x��T�1�y"!͔S� )�G6kE��Th���y�	 G�T0R��j^�i�5.��y�'�:m쨱�h�N�KD���y�J�Z��U��@����)3ɘ�y"Ϛ+B*,�bT���%�r,
��y"�X�q;������� ť�y��V�c~����Q1l�(BPKC��yU@�*y�1G�Z�x�����y���H�����d�e����5�y�l�(bX`9�'V4��('#�-�y��8B�0�K�R���B��y��3�0-����*\��	��y���gk�E����k��g<�y���2K��x�'ò�f� �AǼ�y���D?hqG�U\�,H��G2�yB�@�+9 �cd��a�تvBօ�y�WM�ޜɴ��_�xI!q���y��ŎI��˷h�?DCN�Y�j��y���S�t vd�$�b��+�y�����$-��~�#��^��y��͚��c�>	&�C"KW)�y��H� ���FQ�hR	0"�̉�y�j]�6J�x°�X6���y����y���1]�o�$�t� ��	#�y2��;^��}�Fď3<�6D����y��;�.9�e?.6huP0	�y�!	BnF6�0aEH����Yi�!��\h�=��l�[)�]�"�	b�!��>g�v�d/3.�Xa��&�'|!���e���x2���n�`�"�p!�Ǳņ��J�W���	v��Wb!���f��iЕ�N]S�b�a:wU!�D x��8jV� J�1c�`[�H!���7�F�;V�G=jE��)s��:�!�d�t���z����  n��F�W5�!�$A�\5�=�pƻN���m�js!򤁲0K�� !��c�#j�	=�!�����`��DM�N�Rw��	!��.�p�EY�z��8w*B�	�:E�9���"Df�� ��:L�B�	$@ P�I�<}�l)��1�C�I�b�0b#�+�8��A��F�C�>'Bi�a�@)%t|S�$'z!��D�F�BMCDS�	3�A�����&�!� s�\���(��1���®+�!�D�g��bV�!l �.��O:!��'6�J�hքS2*B�a��.H�!�� �d��.0w�\�{�Ù[$Hã"O��[�Nߝ2��`З�W�A$�'"Oe��.��K�"e��Ce� )�"O�p��ߔf~@$���֨K��}��"O�"�k�qRΥb���O����"O�!�1�X-N�ȡ�4k�(�"O�R�`ڪY��m�q�F%�"Oz�z_)n�KBb�H�r�+��t�<aPa�3r~j��1�3d}V��[�<	v�ɓ��e�%"�1�`I����<i3�����2fB�!��d��Jq�<�&@N�~sfQ�#� ~�J���/�C�<@�R�l�Sw땢U��9�uz�<�S\����ǝ���Ш_�<�"惲8D���h�p2\����Ea�<1sL\&J@�B`/D �!�/�s�<Q�֖dz$13'�'3����.Ll�<�+�4�4Pb�c҉cAE�#Ym�<iw-�2��͠3+[�`b�#2�~�<�d�;'D�D"܀W���Ox�<�� ���q��LQ| �"�MHt�<��@M�d"}� _y81�VCBo�<��G�{�N(AC� �D0���i�<���[��d]	n"tBE�l�<a��Zx�1!���w��l�eÆs�<Y� :R�ְbE�/c�Ƞ� �q�<I�C	��1 �%�?;�����DMo�<�A톽nh{T��#|���
�g�<	Q.�<b'�)�	�&TD�y��	d�<�UfL�A��	���C#��@U�<���Ӏ,3p0�A�ӥ#��հ4N�R�<97��f�:T�֋ӇG����f(�Q�<���|�<Qѡē�t}f�%�S�<IEɃ/9V�02b�0u:�z��R�<A�iD�НX��Q(K� �@CTE�<I�o�O���;�&P ㎜H#�w�<	d��@G:l���E�l�Cchv�<�#V�4&&�22�R"�"�"!��q�<!�(��%��\A��/m �)�b��l�<�t["6��њ �@)Z �]�4�\M�<I���Ӿ���K�	/�+C%�J�<�BMM:>�tA���"������]�<�W�#��j0�&^|r9Z`O�X�<9��Q"
�VD`Q��$G�F��o�L�<a���@��h�U���QP� F�<QVe�-���#�Q F:�P�A�<afk��,��:�AB�U�v鐵`�y�<)��ȍG߾�;Mɶ<U�]���q�<�� -	��R�F\��J`�U$Jq�<9\N���c����`ĂF��!�$�2c_Lx�$�����у*�!��Ro��	���+�-х���p�!�DG�F�(�dS�8	�}1�=�!���N�Mj��90��i ���!�D�sN^$yB�Z4Z~e#D�:�!��W�jp�"�(O���+��Z�>~!�$�;<�Bȥ.��"g豢T�N/A�!��?d��j C[�d�颴"�V�!��ϋ���r'�`F*t�c���!�=
.�1b98�ؘ����lu!�DO'p�� ��mߝF�E��Q�pg!�d��h%�Ԙ=a ���AO!��R�
������xARX)�/!��ث_:$9��a�;0X��ĕ�j!�� L5;�cW/|�C���>0�P"O0R���-aӦ)��e:�:"O��@T,��e�J	Xp&��d�RQڠ"O�����VÒ�S�n÷�"r$"O��� �����l��,�*�"O��ԥônL�A{�m�	f��H�"O��7�p �ݸ��_�Ph�:�"O�SF��bąH� ��[I��8�"O6�b$�:]� Y�͂�$2����"O85 ���%��h�`L_4_,���"O��	D��fHW�IjJ�)�*O.�I�k]���eO��)�'.�hǆ�7����
���B�'~��t"-?0��B�H$
2�Q�'2B�@1'��B�:���d$��
�'frY�v�G�$d�X$';Vg��A�'�68H��KK.���]�H���
�'��BǂӌP���Ίt�؅R
�'6(X�#��-T�a�#Ѵo���
�'��ՑtmOr��ˀ,Ѓ\��H
�'��tZ�h�R�Cp��"(
.<b	�'>0��d߅$Y�t;!�~t���'ͤ�Ӳ(����Yj#��͛�'�\<rEL�? Yk���@xd�'��azЎ^�d��,X"_�� �'Kp�A`�E�8��ɸĒ�
�'�0Y�d
G!������ݳo��k�'_ Ax�B��t� �&�Ǥ7/�m3�';H�����;W���o�_�9z�'|=���A�F�
�8�=�	�'�R-Jt�5�
ȹ��p@�:�'�^����6O���)�Z���'1��{���-�`�SR��!R!��'ᄄ
��Dmnv���dS�'h�8�'������% K�6d	2�0��'�!PA�Π;���,��r-~dY�'��y��&M�2!D�[ŧ�=v9����'h�x#7��(<�|h�΋#n2z�*	�'���rSN�'�������e ���'z��"���k���(��ʊd����'���Z�)܂V��<���6c�jA��'eB`��)�Z�|�r��֊�x�'䔽j�NR�M�z�3��/���y�'���hQ.Y@�Ӳ�͑,�8�'��@p�������+Y1V���i
�'��5�⬜S��5֍P:b	��'�P1�\l��[�,W�Eb��',��V�S�wM�LJ�bǝD��I��'�6��cZ�s"��NΥ<�q*�'����%a��psL%���G�=ޚAQ�'* ڇޣgz(p���B&3����'�݀�B]�:V\��4�@�0P�0�'�@`���6Y�&�"[f����'��$��K�c�Z�Y3��)T^�$C�'C�b��� >ڍ�bV?,����'�x��#��Q+��+b�&0�j���'լ��b�IS��x�Vi�#� $��'B�(\u�:@I��٪"�hi��'N8�R2��]X(���$F�`�'ȡ���.��w˓ HT:�'��1�Ǌn��!k��N:z��q��'
��gIL2%������@�"a$%��'9N\�RBV.q���g��p�'O�`h�S�M�hp�v� e��b��� 	�g)�&���N/��q�"O�5J�b�%#���E�D/m�J���"O8�� #EM�~�kT��8O�N�۷"Oh4�GrrcŪ�1�|C�"O��3��pbԩ 1�L�]�X�H�"O
`�C�&J��6�5�8���"O�ݨ`�s�T˷�ݥQW�Mr"O�Țp��;���3,`�@�"O�y� '?�h�щ��R&ى�"O-��� �8���@Q(_5�^��"Oĸ��a߿x){��]-H}�"O�PQ����;�
���Y =����"O:	i�j��x��!���RR�v�P&"O`hHܪM@��r��h�"OL$8�æ}L��2�@�_�m�#"O֝���I."(��E�A8sY.��"O�,{@/��ձE��
V��z�"O0u�R�-BC�aI�� 9Q�e"Oց;`#W.����%W��;B"O�����s�ԕX�H�B<d �"O֩���� )����M<*�p�G"O�Yɰ膩 �@���G�$Dыp"O��eGۂDĐ������>\���"O�if��f�z4���w�`�"Ojx�B	%(I���h�
 g"O˶&>d��[����E)I�y� Ͽ
���[5��Y,F�h����y�T,<]l�sg�7F�(Ŕ/�y"�	�)�	�	T� �g햩�y�m�#x::��(�`��c�O\��yA�_F��@����T�ʭb�Ɂ�y2c�	�N���!��\�CfFP&�y*�=�� ����?~��pɅAƼ�y�IUr�0C�m�Ic���܏�y⃂ �Bd���u�`$�`��y���!��d���q�ؘ0�.���Py�� �|p�D�X�~~R�;�EK\�<�E�T�H�p�cVs7�ȈY�<�F̛�3�,�#�J��2C!�\�<AK��V�H\@�H��o�RA�@��[�<��I��2���.K'\G��c'�Zl�<��C��(�ʌ��CO$Bye�q�<�ь�6I�!ie$,���y��B�<p�Q��R�D�I^֝��E͹!�!��>��"k�,u.���'�^$<�!�䍖?��Q�ɜs!"��"�P1!�� �̉`�B&�8���!�4c�!�dD�Y��1���̫����*�#>O!�d\#X�$(��v�X/�	0!�P�-��L	TC#V�M�!��P@!�$ޙiY܉i�7 Fv�bw)s!�$.?D��2Ŕ!4
x`����!��2.<�w�S�@��1��A<�!�$��hb�����N�lά��C'�!�$��5U7ʃ�s,ۂk:�!��J�o+���6!Ƨt�q�#ߢ�!�d��K��Uj�Ybl��@�8x!��,1YG��p'��'�N!�$�0B�dDq��3�ts@j��^�!�G	����&3r[�(T,!򤜀Y��#PHV�Jyn�8�s!��ݜab�4����m�^` ��S!��0%D����"$Up!�R��H!��>�(���C�+���b��>]!�� �	�G��R/���3jX�;(N�9e"O�\3�(�TlC�� ���(��i+ў"~n�	:"]
�g�=�Ȝ� K��?_F�OP����(b�lJp�[�$k�d2�,¯���^�� )0#C0�X@�I9uD�8��5�.�S�'T;�L��h�!�P�u� gBԅ�e�L5H䩞�6ǜQS�+t��Q�On���ˇK����93�\��"O�2��ec(c��ƨX0��`"O�q/�R�J�W��	?(֍k��'��	6 �"D���
-|����YqB�I�&>Lб�^�*�(+�O�g�BC䉔� |�DL�b%���'杗V��B�	�eP3 ��	���!�+?
�dB�I�)-^���)��drs�KR��G{J?%�2c�/�@%�ͼ+yH��g�j�=E�ܴ��@��S/(p�qw��X���D{��'3�ؓdO��QAn
?/�a+�O�����X"��mݹ`H=����	W+�	�<�J�ЦOq�j��"
�2 Ҩ9@�.��J��7�'i�!��؇dl<��{@�V$�D�MH�	Ex��)T�r�R���� ���P�DY�=�a}>iC�C�Q�p�ްf'��(Ɇs�g��rD�C[���iƲ����f���'h֐G�tcv��yu�P4���L��!�p�A�4D� *H#	�Z̲���-}$�P���T;�4��SF{@�;fIؑxR ۟<f�|*�c ��y��{��ѹ��U
j 
��3���y"�'=0A �O$PcPd2�I8*4p%q�'mڌ�R�*��k���*�����'m�(�P��=\�&��f�O�"�li��'>%���N+�!�ך.6�)P�'���a�/�<ƙ��O�z���L<�r�"|OU)� d`�L ����DH���Q�O�U"�c;S_�	�e�]-u�  	�'B���g� x�B�L5����O���D�4D)�6����	!#<!+A�C��y�"$�z��G�$l��D��yB"�3�����gdv��Ə��x��'�IZ�N�2-�&��Lʂޜ���'�a��ȩm�)���.춨���N��y2iLO�2h8@���<MA����yb��/�� c��	"��wI���y�nΥ#����FT�O;&�/W���'�az�n��`J�9�, BV+�N���<��k�*#��<C�Ӱ�*l�$��@
�B�ɣ.Ԥ,Z�hf�=5st�@!LO�X�>`�Wr���Z��Y�q�� 3',��<���&"˪EksLP`�jYZ4��y�<�U���(���a���Ф�V��t�<���2f�(����4H�9	ap�<��c[�C�,��W��0������k̓�MKS��>IO|J˟�m�!�����D#��?���q2������'cʽѥO��D)fx0��2Z9P�6&2�S��?�&j��c�! �N]D��"'ȅX�<�(ΕkT�E9��؃�|yz�	�?���'���`cT�Y�uNU�͟�L��� � 9��ۋR!����F�"���ȓyl��2�J0Q��Tj��ٰ�B����O�'�Z`3�K\����j1�$Xz�N��3��'����E
�i��\`U%I�O�K�t�Ik�����>�6�ϡU^VP)�'Q�:�ّ��o�<�!�4�0!*���<��ᱠ�7؈OH����(D��ɲ��ԕ5@`'%M1!�� p}z�C:*��p� ٦sH���%"O&i��U�I*(-c�\kB�����Oe���i�Of���@Cn� � ի߰w%ȥx��x�We�����̅Q��Ӑ�|��Z��-� �=���'o�S��?K&"U���Ucb��@h?+.�C�	���r�G5^��)�-�% �P�,�S<��}�pd
�M՘@��D��Z�xQ����Q�<9%��I[�x�HȦIx�����c�<YU��*k���AɞyM"I���J̓J̑��'�H� ��R�B���l�"ap�q�+"�Dܖ�0<a���MVB=��� eߑ��J�͙�<�L>!*O?%���1����BK�_-�x᳥=D�����.Z4���bLK��J��0?��O�Ósl$rG�M$r��"�ߑR��p�ȓ*����G!4Q�4C��H�<�;�4s��oDC����q�:�M��y��X�]��!�#&�8:�R����e��D�>��!1���fV������az��=	\\��?)V��d̮F�!��1�g��z/�9��$ma��"O��Чm��*�R��R0̔�"O���
®�@�{��V�t�5He"O�u��HGWwd�qw&^(g ��6"O,��[M<���� w�(��"O`�t�r�:Q�r��vO���0"O��b2�-e�pm�*]>�H�"O0(��H��L�&	���	~=0P�"O��r�;�8���E
�:-4�"O�Y��1FL�<I+E0E���"O���B�Ƹ4�b� H�`����"OFU�A�V���dȚ(���P�"Op,��. �q�$��1	�L�c�"O0�2
G�z(`��0�����"Ox����m�`4���  �^E�!"OD Ys�ԗF��5:�A,Z�ne�7"O���� J�;��4����*�z��'Nў"~ZЏ�y�ɢ��

k�O-�y�Y�">�b��S!_lTS��@�ybDPn>�+���eϚ���"���0>iM>�dn��-J��q6��/i��H��^�<1���?)d@`Ri�)`���@֨K��hO�1E{��Y*T�kbg��k�Z1��+����m6Uis��5!���W���{� ���$;�O:�PCg]DRڅc�,̏e�t�(�O���&_^����f�3e;d�"D���,�R��R$�t�S`�!D���W���!Y� �wj��/�ȱ2	�''�܁��� C��!���$�C��hO?���5v��S#��5@\� ��<��ضT�<�t�O�,�	��NV{�<y�UC��<1�BJ$��u��5T�X��ث٢a��-&�|���:D�`���{�������Tlf��i&D�����\(2�`

Z�t���8D��S� �@߼�I��l�BV�:D����A�;pZ��dȉ�C������7D���%�N����wd޹rD�4D���q�G�b#~���N߹}��1��M(D�`� nO�`�d��-�{�l�� '&D�̐�!<e.hb"V
U�h��4�6D��1�"�:b3�AT�y��\*g�(D�l`�`ӧ��|eb�m�R,S�*O�]I��0y����Ǒ�Ȣ@�"Ob��RL��NVi�էK�1�\@YP"O� Z�2޴bz������o�^鈲�'��/���9�G҅@Y8�$ �27N��ȓn������ ��5�C!��l�$�ȓfy���rJ#"��F�$|MB%�ȓM��`W�;4��kš�
��1\L)zr�\+J~�y��!E�cȶQ�ȓN9.Qq�Ƶ�d�W �#|(X�ȓx�蕸���3�2����$4t�t�ȓu�x|�'Ý n?�h`w$7�i��yGj<3���.vH��v	ʞ?+�ԇȓF�F�SݺV®u�� +�1���T��u@�(r�͕�[�]�ȓL���@��s�I˓��
j��ŇȓC�Z�J@a[*�J��� Uin4��l��Au�$<�-�@F�{�rU�ȓ	���@U4O���%G3�ȓ0��pQ��2y��U��l۾�m��F���(Q"��(��=��l+�h��p��|��)Eh��:�l[$��@��v�d�##���X0�D*��Ԣ3}Ω��V.8 NJ�������Q�i�ȓ9�.D�s�FZ�4�F!��jk`������ʦ�Ė{8�A�D/[�4U���Y���g�n�Vcؠd:\9�ȓY�Ju��cٓ-���B�����b�(0����!A�H�p��1�K�<D��9�F���K�/�$��C��J�<�T�>Vf��ad�*�<�k�A�`�<�&,8'����.	��ࠀ��^�<A���%*2�#r�� �)X�V�jąȓ������KL*�!���L1�`�ȓ%�ֽp���$Nvyat%�,{�*�ȓ:�D���d� �Q�mơ�ȓN,�KE�H�<�0�"*�|�ȓ�α&ߟh�t�p�@ԟ!8Ҡ�鉷M�~��
�fNH�n#�Z]�i?Pn8C6ဗj�FC�	�xT
��􏛑<�D�X �ŗ,kC���`6�V�I(�C����B�Id�Z�`�#d ��^���C�I	�!B)�6&&أ��<<2B�	1$�T�����\��̂�e��C䉕/��iuH_� $�1��>	�C�I9Pv�:�U�I(x����0DzC�I�=�"Vܪbep�K֣�a�B�I��T��X[��2fiԅ:��C�	��F��M�>E��:�cH�'��C�	��lX$H� �)$�ʬj�zB�ɐ z�hp���=Ghd���F
nDB��-�&"`F��l0�3��+ �ZB�0�$��H��p�����i�n|C�ɹ.w������0p>��Q��V�8[NC�I�h�Ѣ�=Y<��!AmT�UZZC�3=�5��F?�F���s�6C�	�!���[�g�8���[Q�Ԥ	�C�	�&u��*�E�H���x����b#�B��1�A�0�V9X��d�%e]=x�B�	�]V=J��ѕ�p �M،L��B�	!Pu�yP���f�ba`t��U�pB�I{��� +�M�z9�U�̞$;<B�"���g�P	�2AK1o7�C�	+.�3�nD�>Q*�@��8��C�	#txص��=%'��Xr��
]'�C�� ��YH%N�8,r��C��C�I�v�^I:���bU�]p�	y74B�)�  {�!J/)B|�!�XTR�0w"O�XTG͋#7d�HR�+]^�G"OhAP�.�7 uz�H!� ���%"O.��
Q��e�1) Y�f�z�"O&��7��0a�9xC��ɪ��c"Oij�D @��[�!�'I�8P�"O6�(�K�!?�ě��]-���5"O�����6%&�����i�P+�"O��oͮ2��q���K�GX0�F"O���<w����Ɓ	*p^b�QW"O"\Pw(ͦJ�Q�� �Qd�S�"OؽFk�4�恊��W�'F A��"O\�"�f�2��I���$$��"O�!a5��$k{�$��Z�O�Qz"O$����*"h��qԎW����I�"O@ XG�Ø�0���+����"O�P����ݶe*d�Ӧp��h�"Oz�C�.M��;Q��('0HI��"O�h�� Z�:bb�Q���X� �u"OJ��/��h�`��E����E�"O&-�4���0��4����.i�>�sQ"OBTx�c_�>8PZ��ګxd�Q�"OHd�u�ܗc�4��Ao�B�� �6"Op��Q�۸1O
���N�1��}ʔ"O�*�N���r�{��ʬ�Z��'"O �����]�H�cю�}�<ms"ONX����h͚��*L$�!��I�8|���%��TT-9��]�oq҇�X�[U�|���<��U��JȕD%ƥ0�6'�B䉦#W ��-~8:�f�+z�On�x��`�(4A��d�#f&����K�i�x	�G��<F�|2�_4{)��H�!5���`�;9�v�H�b�on� B�[�J���	��䨲�qD@@xP��).V�<A�������rM�pGFL``�
���i��]����F�ή�˵N� !�d#o��!I��K���@�왿�9�&��"f�X�t�f̖��	��o�Q>�����II�邬Y��Eʆ�E�Lf!�1(ƮI�ж�YzT�#LВHp,X�aӦx@�#L�A��T�Ʌ������'����b�.`���#3h�@�r=*
�i�5(�5z���+]k����$u���h�-�-C�ܩ�V�]�O�xͅ�	�E�z95,C�um~y�0�Z.?h�<�C�@�n)i���venY�Nڟ,;n�R\ws�D� -�_@ĩ�Mnf�M��'WNcB��� �zWʌ����wń2 �ӑ耮t������|PB(S8���$�!U�P @t��6J50)�"O�%�3N»>��<C�+f�-RT���9�4�Ӄ�"r4��R&�� @>��vd��=9掐�H�<2�A���"mx���6bۭa�Yc��P�]�<�DLW���*ƮY�B�ջU.I�I,� -Wz�z���qh��tnκ-�,� Ř���O���+��vx��A�,Ϊ	[B���K���@�:f�\���aR}t���Iu~d�s����Js��h���wI|y �j<bb`<�'���c�˂�Sg�-cÃا=ML `��{�'e@��V�։I�8PR��C�2��'�J\��f����zB�B*F�l C�W!O��1�faH� :6�:���1�r	�d�߲m�,rb�ª���P'r��y�����FLU�Y��z�ʊ�9��D(j���?y�ثk��8�q.�3�5Iv��>��Iq���%B��[�`�>�c�MP�!�8����}�'{��� �0H�O� ��Wj�g��(���ɇC�dj�H�=W8�ӕ�Q��Q���#j_���"�9%V��#��ĸ-�v%��)}�sB�<��Z�r*�Tx��.扯_�T	X6/�<KK��A���Qʓ]� �G�1MlR0��/S���e��dr����zם�t�,��Ã��z4H5{��ѽi���ɟj�ہ��W�az�ě1@������I Zj�Z#pD�9;4�J6�,�� ��2+�h!D�C����-�V�!�9#ن	�c�3���B*�������t��@;�#����]�q�Bpo;2c�P����]�uA��(��s����z8j ��L�q
�r�O����CA/b�N=��]�T�#2E	5�d���ɤtJFu:��	�'�f��E��	P�(P����$09������1m̥��Bo�mJ#�I*}Ҁ1�V��P�,RCF��&�(�"�p�ɓ(�R|)��3A{`ʓUKDQ�� �������r�4Z��Vl�	1Dsl8�Yw�51��lB(V�d�a��<��I�'�z}h����<� |!r�V'&n���F.AV؄mא#lqA�F�J�d�����K�r"���$	ƮG�S�<qt��0t�T�[���n?�� ��%F�~b)Q c�L�LU�0y6��s&B �۠nϞ��0�BPy2��U�V*�D��|[�lZ;]��a�?kT����M�Y�џ4,36�����ͫ�ħ_�l8���I�|�����
�'���%/�$�����M��?�`�f�cG�s���ə'^�����)����Q�*�<i�/�<���1}��)�'S�j�Þ�(�I�gD_*d��Эu0��A~A���剷J,�:��W|x���N�pq�L���2Ǧ+���&?���G�sKZ&
��q&���y:�0H��,�Չ�[��|��V|Nm�ǃC(x���bG�X;e�U'x�'F�H��%	r,���)_�Zv�+��J0�AsaE1v-џ�	�	�\�>q�p����;?�|���*��C�M%�M{��׎!0�Lh�^~���isf�1 �)Z�ؠ93b��0h�)Olq[#f�;X�H��|�2"��$;P�%iG-Wk.%�0�r~2�X��LZp�'s�1�1惭8>U�`�\��@Bc'=}�aܸ)�5�����O`j'���:0��Y#V�}*��X8�p�
�/�6!`�g��l���͉4��a9�cC�Hr����� �OV�Xd��`D�<���&Y,�t��ɭFm�邤�R��O�b�i0�V?��4�&��{$�	�'��ZA"G�G\�[���>����O�$��lY+O~�O>�+A%ȵa��Uc�ԁ,.F�g(D����u��(W��9l�ᓤ�&�I6b��A�Q�'�*�p�&�GL\�9�͞>	΀�	�'@Zt)!eѶO$����bD�� �'{�Ǭ�v�L0���?��M�'bP��,F9
.4���V�e��d�'a�1�0o_2�s�KW�X����'����
.H�@�d�78Ɗ��	�'-���E�P"D�.�af+1欀�	�'���h"��\��@�s�$ �"O�8��R*���`�,P��"O�m���6R��˄�ƥqֺ��"O���A�8VXT ���!<S|�Y�"O*�:u�Z)%L��T�Āy3"O���7��+D�\� `�-P���"OF=�)D��H��V�9�>H��"O��kP��MC��� c�8چ��#"OX ���,Bp�"�".�R1G"O�D��H04f6a��)qs��@�"ON):2#�3@n<���݌SP�d�"O�u�6��*a��5{�-ٯp^p�"O����oA�1'F��@^*D�P!P"O>�H��^�S,H=����>Ա�4"O~$����/~"��fƂ�E�< �"O��SaI�K,°ڄX�I��(ܾ�6��i��Y�\c�H�6�� �P�H���	4�-D�k�OַV�k�F.��5��ͱ7�bqsH�g��|��]�tʷ�GI����V��<	�/O;�d-1e��!����>s�r7�i����'�~�!��D�X��QٕzI�]Ys�Y/C��)��(��F 2\���('�ߵ�H���H��Q�0�z�Z�E)oj�<�"O��!���u6�e�I,gL��1�Q���{'����j��A9�q��'J*��%�@�
��%�"#@�+�d	p�'K.���R<=3��fE�����a"K��"ٓ�C�mA\��1+�h��|*�*��R7��Qǆ7H��`E�>O���-�>?�i"'��*)�6[� Ǆ'��[e�=�x"3PwE!򤖏I0�R.\�T'P)3 \��	�q^X�xńM�qwf]�e����G�$O�)8�� "qO�f����W��y��
�}�&��è��A0S����gOC9:�B@���[�"mI~��y"��c"���@�Ӗ�>��FG��?�^'`>$L��Q�o�,�p
 �6�`6��FAɀ��A	ӓ/0��7�E�Cs��A��3Wj�G§ށ���"��a�t��Ċ|j5Ȥ*Q'L�Q��Al(�Z�"O8��Sb҂
�fx��$���<��^�p���ړx�\��ʸ������g�π ��a
�>DΖ=q�$�h��Tx�"O����J��߬l�5��N�ĳ�
މ�0��m�'Y#��`>.��O"1OB�I1AWb�ۄ![v����'{F�aQ�Y-�����ȍ+y�Ȱ��C!dy����J�=�Ș�)̻i<az2i�&��}�r�7|˒D���-�0<Ivo�� ߬�V�˽#`�����g�,���I��2LD�һw�I���`��#͆�+�u#ӏ2P+H��'V��f�`�N�0A Uz��D��l��7�~�K!���ty��D��y҃U9f�P��!�){fV���?
5L����$+ �D�RK�ᓈ�L>)���j�����ʹ)f���H�F(<�ō��p�i��J��=����Pg�|�	��[��=�D�P`GL��w��?r��K�OCX��j��}��5r�(�����+��b eJ�ju2Y�*ݾ�y� u�"EA�=>���D� ��'<:���$��
DD�dD��r�	."\R�-_��y��V'[s�P�Cl������Dt�%���\ܓ:Α>�^�`��2���q�:�ӱ�\�|z ��\w����͇F����c,�:_�L��ȓN\���2 ԋ��5�ɘ}����m�T٪��؞cAq�h��������!I��эlǮܰgj�}5
���ڜ��w���]�6T �J�<�j��ȓM������M�=pL�&��݆�XH8!s�#�$-h�(��A$) ��\8��0�&L�}�)emU� ����IN�{!GG=#��Y�HI�3HB����bգ�!�%�����: ����)�9�� Ͼ82��7C�h��V^he�U��1	P�Q"r�W��Xd�ȓ!��	��G��!$'L%iż9�ȓ� ��Y�;��6�T�OV2\��'V�=�`)�54�j���i3C�J�X�'a<� ʎ���
 �
���'���3�X��u�
����!�'I�\�Ձ]�MC``4\+��[�'�c��Ho����	j��
	�'f\e�X����̎xe����'�,{s�U
K5	a��вogQ�	�'��!2ֿ1�~�c�lۨc�.���'��tjP ��X�.�!3�ޫ^��8@�'�v���M�*ffNt�CN�Snd��'�B��e�>Ev�sl����I�'Q|p��4$k`9���X�F5����'�ruq�`[
�h�Q�.��7j�y��'\��i�ρz�^8s#V))U*�'���s��]<,� j'�·$g�Ԣ�'�� �d��>����6��WC���'��q���Iv��LiX�'S�@Ys�!y!�U#]"D� 4
�'.V��,�氱�4l��Nk����'��҉��L���H�6�Th�'#���dזj�R�J���7��U��'�v�ʇ�Km`|S�iH�g�`�'� @F�1�d
�(�Mk �a�'�t���ֶwn��@�ν,��p�'�8���H�'D�@g��v�#
�'YlE{0��>. 0d��3
!�`
�'@p��
�H�T��4a�� �8��'�4Q�0%T�k�Аrԋ[.�Z9��'���DN�-F.�+VfU�J�'Ԛ� 	�Am΁��k9�	`�'��nJ;���C0�J�<��ݘ�'���Ǭ;�Pp[C��2����'�r<s��j��`�"��2�
��� �A�
�qIZ��G
��'AL���"O�����MR\5�P;
Nh��"O<�����/MƬոdF�J)d�h"O�t[bgʀ I"��`�-+�x�"OX-xP) � _�X�@dU�7@�w"O��	�2�yh��W;�@��"Oޘ��e�>&��c��F+*��`�F"O��)g�3�ne��%�Hc^�8�"O���E�*����'��9q"O�5 _iW��q����P��jP~�<a��˦cX�$�2��mqo�t�<� �	/%U���g����#�_q�<)�
�5/�;Ą�f��)P�/G�<�G�I�\y�́a�4�cA�<Y�Ɖ#2��I &䝴0:Q:��|�<iA"̫}�A���7��l�΀x�<�'�čn���z`/�@S��	e�|�<���RK�,:(��� �D�<����T�\[�H?�\� �B�<Y�*@�sI����ǻjr� p��U�<!B�ObA�֨_�F���h��L�<y�!	Р�hх��l�v�<7��0�,�J,ax�3�n�<I0��*�|lsnD_���{#Dr�<9c�"����+/hRT��L@n�<��O��?v8 �4d-ǀ[��So�<���\1F�Ll�k��x�ıå�HA�<��X�u�gd�*u�D ӑF�C�<�&W�V�87&mv�c�&�S�<!̉�pT�H��n��2�l���J�<y$�Ϧzr&�����N0�ݠ�Z|�<I'��`����C9�t)�� ����ppH��9J:�$�"~F�6鬉a����X����=�yr�y*��Z$�*?Z4��L����T�"�^MЁ"A���<�1' 	d�����l+#�U2�o�t8���	>^�`�9bC)H��ɱ�MȘdta��H�1�2��ēAd�YC2��*O}�9���"�b�Fy��En�q��+M��vd9s٫5s2�8��#x��C�"O�DMԌ ��`�7DZ���Jġ�c�P�h�O�zD�-����2�W&t��M�r�I"LvxvmI�y�a��z(8*�Ń�r����P�~ba��+��PP#�.�ayѦA���0�$�%fC���#_'�p>a��H�z��u ��*�]bUdL�T��ԯ4l~��	�'H}��ϛ]�pp1�A)1o>a���M@U�AΙ^�tb?ɐ!�ھ���C
��`b��3D�tiS]�E�- �\ �C��<M�u� R�T�
*O?�d������Д=�T�H�l	�Z !���N��d@���z���+~9�O�-��4�j���` *W�h�ɠ�`Ϳ:�@ܳd�'�DԣDM��K�4�H���(�L	X���z�<Ћ�"Oh�������{4n��mK�Qk �'�H����37�V����$x�T.�
ynD�I�;B�XX���5��k���`��U����,*��F|�&qYC�&�(��O���ia�	_�BըeL�Q�r�ON��D
,a����$�r��Ac`�T�h���H���]5�{��F�,��!�h��s��O��	��D覽��#�8�x`� ��c�G,��ڳ��"w�J�҆��E�\K�"���<J�JĪo�~�j�@�A"�x�񮊡p�Z���4���f�9Z��D/2Z\���?%B6i��Ǵƣ?aQ��H���p�E.� @xKv�	3CL�"������ �
�{6GQ�3;��pbI��y�Dp��8�C�j��c�ЂŔ�mMr��PE�>�{��<ف�Bt��pk4�ݾ. �HQ����$TGk�@���� kݑC�T��b���8��������Ҡ��c�d�Y��'7X:��Y0�#���8D��A�"�E��]q�#��`Z�3d-,;@,���?�ݠl�,`鱂P�($Z�8��Z�0� �5�[i��
*#N�T�.X?h37
�'�S�g Dn���×�s�P�(BAO9fzZ)84�K�^;`WZ�4�4Js�7� f�@��4�I)�!��$|@�W�	��d���*H��A��(Z?�m�2�o����<Ǌ�1
�(G���F�ќTE���W\�L��6T��B�>�%-��2f' I�`�w�ބ<˓`(I�ߟxZ6��D�x�3�l���E�O�%
`����6)�҉O�:�2<���*���6O� �c� mS.�b��!<O4��DE,�<JR�ݐM7E��%���"1�A�%V�����J_(��l��.���u�Ij��넭G�nk�-�S�E,/4p#�lF>�p?��o����MYw�O0h�|m���@k�$@Y�tG���X�d� $A�bU�!����#�ħBʲ�#s5D�@#�F M�u���U�'�V!�X>�&>*wi�pW]q�gA'z\��"�N�!p�Rc��Q0q`��O�	\�AU��Qȟ�d�>��y�AƝN�~��L�6.��uH(}�Մ�2��S�O7� �C�_�,�J}h����pX2�'��-���U���� H',O���.�Ew٩���7faR��k��C5h
���`/��4m֝�;AF�1�柄d+X�q�z|�Y�b/2j�����}����+T�D^xQh�&'���1�S�,�N�[L>��/�Z�dE���O��a5�
<�H�Cf{e��e�'�WƎ��c��2a���<1�e�O��p��g�#q'B��ig������u�Ds�O?7R�<�ʽ9�+�>i���Gg�?��I/n+�f�KH�S�O��!׾�E(��1�Z����g~B �.g`�p�'.NPPn�8i��ı�K%_<�1��$}BmǖO�`����O�Ģ�� ��S��"CPv	��Q�]dZ(�
��+�1���D$\rDȱd��.$T��[d�Q�'2\d�e$�O�9Y �V��A�!eT�1jB2��� Z`�EXw)ƕP�O�d�,0�P��U�V��tMi�'u��1��+<���*��:7pX�O����v&l�O>հ J)`�҉�J��gr�d�;D��p)F9S�&a��)Ȱ7  ��+7�Mȅ�'��y���Pw:)��� ��p�'�Vt���5��L $qZ�l��'dv���KT%?H0Bѣ�_�hQ(�'�J�;P)
c�|l��GD�~�P�'���� ���1|���Dƭ�%%�W�<��
�(X�}iSL#0��iS$��y�<A�^�>4c4,����a�I�x�<��섚\\��YS�Ԗj���Jh�<6"�H|��a!��in�E8���N�<���:�,�����<�D��`A�<)Qըh����`���.��D�B�<1��ܫ/|�9�!�5oSfx�q�x�<�F��LZ��E�D/�6��AL�{�<�WξA����Ɨy�f���"�}�<)���C ��K���E��{@�y�<!�C9E�xr��[u���f�r�<��($�:Y�_�EZ�j{�<��;,� ��;"4%J���X�<1�O�>������A�:4H1"�	Y�<I�� 
r����l�z`=Z�gNW�<�&F�rd��h��:y�b�Q,�S�<1�i	�F�Se��4}�����@O�<�t'J�:]x�ǰd�DuɄ�P�<At���fN�+��׭Dp�l�ƫ�k�<Ib��B�(���+31p����x�<�&bH���"ή:��MB&�B�<y��_3v`n�t��.iL��z�H[x�<f�#y"&�B!L9��|�<���ޭX�%3����l4z�y�<Q�%]�Ɣ v)R���\����v�<Q�]>ob��GG�x�.�ǃ
q�<A��J�z�3����N����7kXi�<��ٶ�����$2��(A��i�<Q� �[����Z�j� _r�<��'��ҹi��!#P1����m�<�F�3ڹ�6�հvA4XK��d�<0/44��`3�
p�z��A��f�<���4�b ��&�vD����J�<� ��
G��!ip Y�s8�'e���N�KX�h�b씎!���0�L��;�d��F�$lO���%�ԭp�*��#k�dḊR{�=��@V�$�NB�����sI�
8���	�#T���� �A�_�h��V�o[<� �L3�4x5��1J�C�-��D��-�39Fx� 瓝𚨀R�M6j�6�'�-E�,O�P��1H��U�䃁�wt��0"OȌj���j:Ȝ�g�ѭC���C�L(tx�|�f��}�a|"!��c��M��+>k�0��T�G��p=�/�6
�*=؁�x�9t#F&x�N�B@�Yu�Z�� a%D�T{��Z�5<~��х�X�ٱG-��ܸc��F�?�#2�U5Q��8!�u��� 4g.D�@��+�ʂ�����2�x���6
��y�l(}b�B���`:z� 0DX�v`x�B�Q	S�!��z!Y�P鱴��9���A�_b��U��JZa|�̜�K�l��L��Uʳ���=)�)�4H|޵�'Q���5hKz1dL��g�"�¥�	�'��a���-�%��-O�^�q���\+7, �G�d���'\���bƖ4�|3!��!�y�H�������* �M�y�*߅H�!��A�v��Bc�L�<ٰ
�4=������O��qI���}�<����+9�R���,G�S��а�]z�<�D��!"�\��L�[��0Ɔr�<a��>l�	j��ޥ5[��P�)�s�<ycOZ�[	�e����)?��p���g�<�TmG�~���CρAɮ|HN�k�<)��&v,�AV�@�G�j�c&�	{�<a�JR>lTU2i(Φ)��oPq�<�R�
�V=�bGDROĔ���g�<���`�j0Q' �#"R��t`�E�<i��D����J& �D]��NAA�<I�	�l��-y`��&�����d�x�<	"�X9*1A� :Z8�Q+Ʃ�o�<Q嬘�/LdY�alL5~yڭ��N�h�<IW�`op4����7���D�R�<A�&	~�
�`G-�0 ���T,�u�<y�s���;��Ev�s�<�A`_�v�B�i0�P:(��Ӧ&
`�<qď�5G�j�q4��8N6np�`.�G�<���O5�B�PA��ED�פA�<9ue�9�@d�ҫ�4��ax��U�<�u�$�j���*���"�Q��4!0��G�L�f�-T">I���6i�	�k�W�  ׄ'D�T�!��x\�uc@ꐳ9)���Dg)D��i�!:��	[���/�-"sH#D�أ��˷%�
��c�x]F���g4D��A�F�(g.���d�(iZBIS!.5D�B��=�V��5�V�Q�EY�5D���D���;�p��%o�`���>q@��W��H�<EcC�T�M��hBg��X�,��imJ���R��@(O���T��DI�W��7m�(h
���'%U�]�M����z6����oӦ�"�����ԧ���	-vm"u�AF���q��e{r瑦R�"~*2��I۴����R�@:6휖"B\�Ey��	ƻ"���AI�1�@��_�zTQ�P�W�O���3!$��B<���gQ�7^-X�{��[���'C�b�'���b�!��U.1�O��ڋ��i>a>V4��g�)|l�u2'�����5�hOq�����r$|��E��t�A��1U�b�>�O'dc>a0 ����)���=}O8A*��4?�CO#{��t�D�/}�𩈣s.Y`g�ϟ'���hL:5��f�������$P: ��)�p���8t�\&c<�y0��S�L�G�^C&�a:6�s��8u�{>U��O��~4�۱�̥mE�3Q�X�&��W3O�X�F������	[�@���mI-1^z)�o��s߲a��hJh���kY�������� |�bR���Q���]�Ƶ�3�'Čĉ�.�_�S�O]�\�ə|���1���,!(N�����5>���|���.u�`m�<Z��hC����(����{���Ipa�DL?,�ر`�`O'h|�z�̉���i~�r��)�)k�.��R'�L9@�)`D�9�PB�I\M�x�!GB X`�l��FCBB�ɫ8^�:)��pW�m��^�lB�	=�P�B~�������b)B�I�aqrk�G�>[N|��T/�)P��C�	!�F���l��0�'��_G�C�I�e�$�¨�<����É5JjB�	�C�Ҕc�g�>��t`�R�B�	}���'ŏ)��5�ņ��c`B�	�{ǘ�ٵ.J%B��1���\~*B�I:m���W��O�h���_,PC�I�%֨ɐ��D�<@(s#'�3/"C�	kB`��H;,�$��	cUC�	~<���r�E
?�P�aQA�|N�B�I%N�<\@C�O=p�zm���=e0xB�	:p� 5SgNӥ/��<�q�Z'{�0C�_��}Ad
iF��w�Y�?8*C�ɣ*H����*�J�8�&>@5�C�I�_TQ`Gȓ�Z���Rӂg��B�	T���e���,���,]�OtC�I9~���h��C����T0DC��zJԉWΑ�H���b�;J�@C�I>#D���H[��"Se��e�RC��T!<�5K�^����vՆB�?{�9�� �4r0��*U��B�	��0�"c�|��A'J�&VrB䉒F�I3K�I�j�jpe@0sddB�	���躅	3~�L�q���}S�B䉫wY�Hr*߉k�6d�m�1ѴB�I"g��K���"u��{b�Z:6<hC�I����n"��]�1�vfC��t{���W�ʎ$`�QqE��,4C䉯F�P�Q���pi�p��?�LC��&-�` �Mϊ1�4٘���y�.C䉟^-6�@�įq;u #��dIC�ɍY(��0�9O� J�ˋ��B䉪]_T�p�� Wm���q�(B�	�H�S!��[��a�4o�(B�	� �x	���	i�0 ��6q��C�	�0�<�+�J��7��� 1j0fB�0�t� ��5R{�ݫ��P.}MC�-"�B�)[�ta��b&.��B䉺4Q��Z>1�R���[�|N�B�	�@=�@+���1XH%����?wj�B�	3�ޑ��N�J����/��B�I�\�B0�<P����g��B�	%�l���ɾ �n<����1O��B�RE��A��T�mJh�4�̬w�bB䉘E��e���_�6�"tÅ@L�C��2\��Aq��>Zjf�o�|C�I�L
"�jq#8���)c̪	KFC��''BF,IǠͼ'�z!��\g-C�<G��9�$Q�v.��� \��B䉸*�����X5� P��M[�_q�C�	�H�T1�H�@�� xT���d��B�ɪJ����%e;aoL�rW. �y`B�I�ӡIW  ��P��X|�C�	�d�0��c� �g�`���ͣM{B��sHI;�J1�T�*���qi B�	2a�^���/�!7H* �u�yC�)� �yR0�/d�ܥÂ�m �!�V"O��R"_j�&���'Șz�%؂"O�P����S�"���f��.e)A"O����g41t�I�rE�h�nTAp"O T$JӦ9�2���#��X��"O���H>u2� N�T�T�[�"O:��d�^�!X:�Yf�ɀ9�P� �"O ١����%2�����r-R�r�"O�yB����N��#hԴ^����G"O��Sm&`:�b����H�"OXMW�E",�sg̉�U��@��"O6%�%e�(^,��`
K�H���%"OV�IPB��@�4lkd��1����"Ox���K(2�`�ڕ��JV�`�g"O���󈄫#r��gk],n��5"O��#�in<X˂���*���H�"O�I��_=<��aJ��G>@���"O�LYrI[�#޸�qe��71��98�"O�<��%�[�D��eЖ? z�"On�#r�F�hH�Y��^34<��"O(к�lZ]�Xq���Ĉ�6��s"OԬ`W��0 tH�BE�J�F"O�8����%<�z���12jļ�q"O@À�ƤiU�.�1,2� �"O����ѯ%m�BV5I�y��"O�	��c�/f_����8A��z�"O�H����*"+�9P�"���t �"O.�����E
�9bF"I� Y�V"O���*@�LƖ��!��zW(�{�"O��x��c~�����0c�l5�"O ����v����C�X,�1"O���Q�)I8�X��-5�4Ń@"O���5G�o�ųe�u�j�"ONXv�״_K��;��D�:h��Y�"OB8�6 ȷ)s��"�(�iN�j"OV�Y�S�I")e�̉o\mC�"O��� �0\���T���:8�/�!��B� vЁ#��(����!��a�tp��O�0�ά����8�!�T��:,˂L��	R�I�!�$���<���@%h�HDФ(װz�!��*��)��̐Z��cQ�ё@'!��Ê|��L*Ā�7b֌�Q����/!���)~�ˀ�Q�0k�>!!�x�����C�I�RA"P/F!�zKnl"�}$ъ6����!�$�14#��X�!'8b	ru�P/C!�$=
T�x;j�6Q0|��ߩB�!�߱��90��.}��|A�4�Py�E���x1�N��=z�z@Ԝ�y҃
9\����ǎ�1Ҧ}�m��yr� 3J���fލ&�%����*�y�+,� \�%�$�:q؅�
�yRQ��	�L1~Ezu ��yb+ػ�2��T@�p��4�I�y2�P1m�P*�G�r�YBT���y�I ,?����8Yu�@�C+�y"�@ �U�"�$XZE����Py"��,lF�#�E�Y�������S�<�d�N#!BH�EK�5��e��@�M�<9���]��β��X��K�<Ɇ���W�Fux�l@+6����O�~�<�DNY.`��ő�f	�K�z��I�y�<gH�B��9�,:j��YrH�L�<� �����((°b���#Z7�I6"O>=h��
Y�!3WjY 1>�x�"O���E��:�4�G�!Z'$e5"O���φa�&E���!�m	�*OF|�n�T��%)���K�\X�'A�ʧJ�%)8Ȱ�Ƒ&4~��'�����W�`|������Q�'��x;�@�l����g'�	
��d�	�'�l��ЃZ�V��4'�6���S�'bh�!�ț`x�I6+Q�0�����'�q�+Ee�� z]V(;�'����J'5���lo	���'�`%��X�ڔ��Ya�����'����`j������
T��� �'< yk���:	#DD"�K�0��
�'0�u��$�K�H��B�M(�o@M�<�wb�	Z�dd!��6]�*��T��H�<�4��B)��g�	;Zk5�Ec�|�<��B�T��P�s�C8�Z���Q�<��$KA:�Ȓ֊~�X\	���N�<����p�=*�Q���|� *VL�<�7ˉ�9`�S���Q�O�<a%)�'r�
�aٛa�r�E�<a�搐)x�1J^�%V�II7̀Z�<)�I�k4>`3%�Tp��� d��R�<A"�M��x'��R]B@iqiBY�<�p��9W��a#���|&�}�s�U�<�c�AD�%�b
�+�� �MT�<A"��*��#���#9�l�k �.T��K(k��X�ժЛ_G�Aڶ�(D��p������ӑ˜p�]I��%D��Z�`E�~ia;��=R����Q�#D��ZcfY���;�!�	v���s�"D��S�* <K����JM2�hj�#D�hy�g�u8xͰ��	+u��e�?D�����."�&��B$ǔ�y2�=D��!g@G�Eon!�׻2�PH&����yrG�0��D(f�ը~������yB��c����'
�R�)��X��y��˟��� ���L�}aa���y�`T�b�*$sR�Ĥ"yִ
1���y��4:��h+���I��I��J��ybnH�¥
�;E��ݪGƑ��y�#Q0�S

�{@p���0�yc0%ṑL8_����i��y��uE4*ޔ�s����y� �*`��d��-HLQ$%�.�yRk_wk��S2b�̄�ق���yB�:�xd���򈫂�y"#�i�`$��O9|����&R��ybܺ6�Ќ����,��X��喷�yRi��R�p��8n5L��r���yR�I�q,�$��Q3p�@��J��y��8x��dyV�ȝ<(��Ф��y��Ʉb �BRiH�58������y"i�����k��0�q�/A��y�G>�͐��[(�5���E�y�ㄧs�:I�v��Od���ʟ�y2��-�D��@��I���(�*��y��"^b����؁luĠ�	��yg�D���C�ǘa��!:�	T:�y�f&|�@A�F�Mz�ލ�y��+eR�m�.� $y"dT�y�%�|��Õ8Q؄�q�!�y
� ���/�F�b�2�ʃ�O�a"Oj�Bb�!M��$��k.pֱc�"O���,�%F�`1�� �Rk��"O��N6al��S'�Rbj����"Or���B+K%H��BFU:�j#"O\`QA�3k@q���!oҔ�"O�m"���p/�]iZ5V�!"OX�j"C����E7H�
���"O�b�	   �