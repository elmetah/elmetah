MPQ    $    h�  h                                                                                 �%@=S��cI�+?��::A�����WM'�O,������
�@��qM���Ś�����/CT(��7���)+YLJ<����6ʼ�!�cTͰ�W4�{<.s|U�A�?�4D�����1w��7x.��vWz�0�������c֌�K�c��+�*���n� �D���L_j�½ �(5�%|ן�z*�Ρf��Ґ_9W���*;ԗ~��&γA�Uk���W�����]���pF��l1U�%z۹zjԱv��.����rb�ɑ��/Y�m�#Na�Z�\��q�#	��e6�%����a�?Ow��j{���}�����(ӏ�e5Do�H�`�D�����wNv�wz��C~��x:�ڃi�7�����=�ʡ�ݡ4����Q���{�����u}����~j�1��JUփos:��-KY�\� &�\A�j@i|l�a�U��4�cV���T��A����ޑ�_']y�{��Ȉ��w��Y��M��T^B
�~o�v-&�+K�'(��qg��W���`����rc���A�\�9VG�[��.����,qD��-~co��Qq�:�Qo`��POOMJ�Ң%�V�+��jV,�%~��#�(*[����f�V�%/��6h;]T��a��3���)��͂��L���:�G��)�'м�,�8���'�	����2� �ʟڍ��R.�`�ݾ\�2F~37f����'�������?�����@5��޽���і�0Vg�^���S�s����
IV�s]��<��w�/@ʧ*��w�EQӕ��c�mP��Ea�|�h�(Xc��X�}~����|��@�rg~�T?J�9�6F��ϸ�l��R�u�׀!955�歀� OPY��A��ޒ7��2O� 5��.�Eѱ_X��*T)���B|�1��E�����ݎ��nJ@!FyR��?cπ��TL1D��/�7�"���gf���= '��z���o�e-�J�s61��^�Z�W0�O(,Hc)��:yA#q�=�}3tf��"!R�Q�+�/,)�����1$�v�Zye�t����] U��R�J�T�B=��[���^�0�ꢻ1	oR�s�,Q~wKI���kP�>Eݬ�	�?)�Ǯ��,P�av��)9�p��K_������A5|۴׼��*?��fA�53q3qE!k<M�̓����Pܝ_K V')�ś!��NC+}�{+������a�5�W���9S��a�lH���7�mV�(ʭ�h���0H�L#>6��������C"<��$l �����P9#2tH�����/���.���(�/P�w��/�����L���� ��]\my�q�K�ᇂ�ںC 3��\� ����}͝��d`ی�>�K���d�2Ѥ�������~g��N�K�O[�j��d�&|�q��5Ҽ�!<E�J����_q�ݲ�Sj�7竝���)bR��U~�rh0��dZo��mcܱ�|�n|��탞L��Z�`��o�'�bP����D�T9�QЀ���aS�3k;�;+�7h>V��D¸u����3��-7�]@�<��|��d�&�ȁ�a��@}v�f�2^>a�(����]�e5U�֍u,�Q��Ӧ}����w�m��gb0��YMT��kw�	�
����n� nB��6ua���Y���{�'N .
'�9�>��O�1�理q�Q���.o;o�]����EK]��m��:	'vvN�%&�C*�{R���@���a
�^�M[r�9^�1�xHS�:�&f���Gyd���g�#Ih'��X�X��G�fե��ߌ¿|ԍ�lN�/���+��PS-�൑Xsȯs���3E��"�	�̽+���[�p���N0/���?��!=��ȗ�0���I<�}q/�z�W������&�BՓ���C+K���jfƠ�<h�4�f��*�	����"E��I򍒡^C��;�_�Z����ie�@��o`��w�U���Vo�����������c(#�r�qH�eKx�T@t�B���h��q����Dl����'j�����7[�L�f����d��������c- 8c�ʕG����^�9_��;O��E�L۞�#=4�P�S�L*���:Y�+,��C��o��MhBbqJo�2������<Hy��lō��{+��$}~���r󖁮~��]�{ ���ݭ%D�(�� $�*2���\q�hwi{۞����^��Gdr9I��L�io��䖁�*�؏g���P�uK�Y�CU:��>O�J@5��c�5�ESR���P�� �f��?b�k�5Im�uA�hc݉�6q��!�6��M�w�f�Y����o�h�ڜW�4�tM-�M6�}�y"�^ Y;�+��cXG~����ު���)�Cxm�!�%S; q1�4�����픗�J�O^�1�����	@%�@/�PB���>�����@E!6}A��(H���;���'(Z�6t�u��P����R��kD��ڜ�nT/�	��o��e'0M_	�����_S�a�el?�ݝ�<G�j���!���f7����D�u8��.�τɺ�s��ыO�ɪ�뽛2�b[z�˵��OTG��g�	���tg���r�2ߗ�t=-���y��Wj���.V�N%���\�ށ��Y�MQ��`b��\��:���y�P�A�
"������RH���������W�� L.i�%����-��o�]{�/ɒk�����òm��?ÿ�R%r8�q�4�ȼ���:�� yr�r�{6Ln��*��Y�����'��FC�E�%$�~���};��B���E"eIX�0�Z���@b�E��c��`�-[���l��{AH�{)Y!Y�)�Q���s�F���B1I���l��FYir����BJx���g��ş��==�ߞ�2b�n�ˏ:Mn;��s��/��<��-ߥ��XS��Z1��B)Z
�KYSj5����	��+�'q._��6A����v6Pnc�?������e9�X�b�
��MFR���az0:r�K!2�#�������?p+uC]	�]��m�#����?xL�[���N�7��i��N��(A3-!zui�G�<����l���,�͑�r�d�V#�6k�E�K�ݨ����'���V,�a���V���P��v�L^�W}�2͜��(�4�.0� Yc�b��MZݭ�H�gי�oé��T٥���×R��4��]���pA̕l�wF��q���Yұ��W��OΦUmb��4�/�`G���m�u��\������Ǡ��%S��\B�?�9t��w��(��}	d��Ґ����5�IKH���Ds����~葒����*��t'�~�5:> �i�0���h��¡�x}4���,����SM�uxQ�A,�jK���Չ�UQͦs#
�h߈8x !��b�
�l�Ei�݃a)�9���V�E��%A��
�9+��qy')��!���Iw4Ph�\�M�����FB�+�~���-���K`���'.嘴l��P��X��c>{�A��h9Ѽ�[��.�a[���l�{����oDsQ�M���`�t^O��m��%���ǆ!�G[�VG�$�ئ#��[�s����� ���W��;����:X3]6��
��h�m�G���Gv�)�ڼ��8ڱ�'��ۅ�^������5Tu����.���X�}�¼3r]��r�����`�^�m����Ƅ�8�W����ǚ1��+��g>{��<�n~�U����M�W]�5��7D2w�v��b]X�,[��Х�p��0|Vm뭟�@tj|m������}E���/��!��d�r	��2�?� ��-��Yl-?Q��Gp׻O^5��{�*O�!���_�ޭ�5�0�ʫ۲���gEl�X�hT��c�ՠ��'g�������	q�,DgJ��Fy�	^��;z��om�DM$���ү1�.ۅ�G{'r�]z����e�t��N�x�ø��|z0�$�,��z��Ժy\�q����X]�fRo"�^HQ?9��꧍�~���u��5NM����9�]�S�@oERH`Ȏo��=(#"[�3�1����,?�G0s�IQ�/qIh|�k+�z>�c����i)ԍ�	��{La��U��?�p`W�_5Ln�z~�5w�+�B*��7f\p ��3L�kw� �ė��Pe���Kۗ�)�>�!Ht|C�����ҕL�讟��WI�9.���ܥ@H��L7��Ïە¯�����C>Q^��?1��C]�J���#���r�/H�#�V�+�
�/?���B���q�����*�w$�/����0�g" �mfY0m���F# ��7��u<:N�x���{�i�}K�h}hC��_�Y�n��n����uk���S�9h����űF�\O�A�%�F�|d�������Em�)���_̊��?��R�ŝw�a��$�@ �U��h+@�d�h��(����8m��N������6Z���j�'U�Lߞ��4�T�Z��[�_��h?�'��6{�7ÍފO��_T&u�Փ���>'�-Һ,@��<��R*�A ȁ���pPvݑ32��a� ����� �W����,�ը����J���6u�m�ud��lb��ܞtZsMϱ�kR�ãD�p����[i����?a���Y��{�X�N;z�
��9ʅ�ת꣏��[q�zHl�,�	K�o ��ͧ �EFo���P:ͅ%v�b�%��^C�{R���[�-�>��9�[�y�9#]�1/[JS�l&����&U�a8�g<��I�o��J&Xl��G�ޤ� b���P�צ���N���F�"�� ShJV�,C�Ȫ��� 
d3 W���	G��+�D���޺O��I9� �?�+o!XRδC�m0ב��0}�1��u����Y�ꨠ�&�ؒ����k�+�5�������뜏r^J��$"��f���x�ք�)�<�T����_�wxڑ�4�F����J?��Q1kU*[�F�o�8¢_$�w���b{�Mjq��e�ntx�T�t��t����7���h����ju�����7����!B��2d;~���h��'��-�z��+ZG4P��_�Tw��jo� m���j�=�q5P���L�kƻ��x�F/��q?�JU���gB�?qE�������T�n<�*�G�_�x9T$�}yqc�r�8Y��qw]��J{�*���2�(��7$,!�W�+q�,,i�"�}-�^��˘I�T��k��������ES"֐ҏ�뒨���DU5t����J������5~��S�ޒ�M)�I� ��C���k��I�DGA6/jc��)6�7�OZ!���R�wO�Y�T�����he��W�r|��y�-�^�ؑ�"��^;�qnD�+�}�c���ŹN���.�1-�C3ܛ!5�~.�;��J�ʨ^\��<͗Ay�O�1�	�ĊRw@ �X/ϯV�NU��X������x6�,��eȓ���;����8��)�НC�`���!��͸0F~���OƢ	q���Zo8�7'��f	
���2�D�D��� e��ݘ�n���%����z�e�۶F7�Puӂ�)�I�w�}�.�Ѧ;�%f���^���zr)ܩ�`FG7���Z��t����M�m�Ҡ=�f*�t��W�s^�W��i�7�m9��F��BM��`](�\&WB˸Dr�k�D�����J��S��R��%�>sFצ4O�;u�L�%s� �η����̍�X��/$o2��\U���m}Vߋ��S��c%��8�y54��ۣJ�:�8	y�:�Vsn�*\�Y���LA������`�$ZW���e��%w�a��eD���j�Z�Ĭ�[�<E�ֱc�Tv�hI{�5"^�q����{��[Y5cQ]0s��F��U�&
1D4�c?��e]i����!��x~��g��:Jn=8�q���(2�n���Qh;�3�s���f3��(���b�S�&1��)�Y`K4@��Ob�eg�	�\����*_|��A�Ji��gPIMT?:���4/y�p�
o�Fm)���_&|K\C7��Z��|���1��+0�	���U��#�X�z�/��E���k�7~:��5߬���(��hgu m�7ZG��L����
�`��W�?f�#⇛��/���4!��>�\Ụ��ܕ�1�R�X����Zt�G��W�	����Cn��� �D���M�+��C�gv8~�*P��x[�D���r�+�oq�])K�p<�	l�8ۛ���hX�l؟Ӽ��>�{b0=��y/A�s�ɐ��\�����B��&�%��W�?q���i�C{�}��)��(���P5zD�H��ZDΔ��]7E���u��i�Oj#~,�e:مi�I�N.]��Q=��3a4��\���!�1���us5O���j�v��/?U�6
s�ګ��lӳx 7d�=�'�i�nxa�����NV"��̾A�f}ߔ䳗��jyB�>y�户��wok��XM���:+�B��~�.�-�K;;�I��31���`����`c�uXA���9LRG[�G�. B��B�g�����o��Q�T'�x��`�d�O�.�(x%Â���!l'Vbts#�>][�i?��T���E̲7�;�6GԼ����38|�&���V�B=�:��G1�)���a8���'#ą!�����Ɵ�:�..'j��ӷ���]�3�tq�����%������H����R��T��3�~�̄U�&'�g���kK�=%����������]B
�2�wG��������;���K1k�Hm��؀;��|ȱ7�����sϗ�i�I�Mr����0? �D������l��;��:�����5ku�voPO
آ�S����o���R��P2�0��E�X���Tߺ�Ð��B���;��hR��g�Jv�y�_o��������?DȈ
���R�lk���'��qR'�UzY:��Fte#$�)T���2��>0{�,�k̛��>yw1�q�Ǔ3�8f��""W�lQ����̧HA����1�Ce������]KO��Y�R�Ҏ�y=���[��0�ԡ�� ��'��%]#s�
tQ�I�W�k _>�	�?d�)���dAF��Ha�g��fp;M�_p�ϽWY5r���r�
*�d5fw�+��3'g�k��1͹�����S&nK��)�נ!�0�C��5���0��jX��W�W�9I;$�W��Hn{�7��!�^����_�Q��oh>l�b����[C��
�ZU߸�	���_w#�YHF:���ܾ��.�l�)���%��wzf�/n�1�(ݤ�OW �e8�#*m�A��A�:�8��0U�i��R���D*���j}	>�Z2ԌɠQ���jٚ�Lњ����tqo�*�T�A1�O�� ��6|�����x�1*rEA����_'y������m�'����߉��{�U���h&�d�W���,��P���ˡk����Z3$߉e��'��H�Y���O��T/��6�L�ם�iɕ1�#7��̩O�z<u�ޡ��]g�yg�-m�@�X	<_�+���\���������sv��2D��a�-�VRY�����~�,�H���|���P�ђ�m�F��Kb�������MJ��k-=	�<k.xLֆ�����?$�a�W�Y���{��pNv�Z
]خ9��n�1֏e��q��%�F���Fo;,a�B_EA�V�#u�:�"v��%u[C��S{�6���F�;���0[y�09>|�1�]�S��]&ܜ��}[5�ů��	g�P�I���N�`XG�jG�v���AՒ��2��r�ON��?��<$��5S����M�ȥV�{'3���	�s�+��A�I�I���s�Dbч{V�?��!s����N0�� ��}<��p�/�I͟�cn&��5Չw��]�+������z������7��?�������jֿp��׫���/y_B�(3�|�Oa��6�q%>����U�(s��oh���]ߩ�2�ܭY�_�(���=e��ux�t
ta*P�V:���	)����o�=�Cj������7����j�4?d�n��h��b��-Vݕ���G�Ł�_���o�v�1�1����q-=j?UP�5�L������aRR�9�ֳ%�/���BQT4q@��z�ǎ14�!4<>���"��@�����}t+��ri����j�]��{ַ �Jr[A-(�u�$gM��q�Iiq���X��^Q��EpI�^��᧟Htށ�&��А���&�ݏ��U0����?J{�����5��GS��ɋ�\5�S�Z �̂����k|n)I���A�w8c��6�T����!�"���w
8�Y��e��h@�W�O�8��-�߁�3�7"���^V/��"�+�+�c����T߁��ҒԌP�C�jS!PtJ�W�;���f��CZ1���A��� O�T1[P��0@��@/
/?�黮����z�L��n�6�h9���K�/F;|F�]����Z�+B�h�"�I��H�!س�*����w��jRo�v)'���	%�`��J~I���e�n�ݓ�3�� ��<�/���ۑ//r{Oun���$L������v�����ɠQ��s1���h6z�����4G�mP�y��9U!t]!�(�8�b8=cOεo��W �Q愁������ú�ϏMM�5y`X�t\��	�s�.��0�� ���Φ����R~�N���D��a1ӹV	�L=����g�,�#�S�/k��L�����om��F�����5Q�%�#�8��/48���^�Ss�yh7��1��nLߝ*��PY�sS���K�Kb��{W~$�O��mߏ1)�����e?����Z��ܖv�qE�c����W������o�xf{��Y(`�Qؾ>s�E�Fnxg%1?_�Ͼ�,�=�i��3��ՃxY��gO@����!=3
��T�u2؏
n��S0v�;��s;�J_�#���SA{�1�)P�TK�g��0� �8	�;���&_7�@A�!��lf%P$W�?uDٝ�~�/�5��@e
*c�F��%�We��^K��p�:���wh��t_+�3	���+#�t#��g��@�#&At79�6·�D�V(�!��&u�-��2;
�JM���	A͇H��#�_�{�ؘ��Ɣc��������W�G�^�Γ(ۊ*^7�B,W3`�C���^t�$	� �P��sZM��2�>F�gѹB���n���E��\��M�����]�$ p7��lB�)�V�D�˗f���sӗ�j�yo�bˁc��ø/j�Z�T6�ɫ��\Kش���ϝ%�]�RhG?`��O�F�^�}������M�@KD5_GH�JD)���ȾQ��ë*ͻ~g{
:tQiW��ѿn�<� M4��ð�:�\wb��;un9��8j�z���UG��s�t[��gn B�y��w�i��as��ł{V]��%��A� L��U���Gy]3������w�bՒE,M�Q��/SB;+�~��J-�v�K�ރ������o���>��c���A�R!9��[h��.[B��ݰ
b�E�>-�o�.
Q±�����`�tjO �����%�HW�<����V}W��O+#i�[2�8�72������;����nwG�3��a-��W�=�<��lYG�X�)/"f��p�8���'^.`��������@o�Fg,.Bs��N����3�'��Ԗ��rF��p5n����.��ƻ��n=*�gi�!�og��&���ʔ���1���9]���-4�w�e���"?����S�&�V�om!Mʀ6��|#d��Y���0�x��'���ʶ�
�r8~2�Ng?[���g�l� 9vl#f�MV�15>0�qXrOa7�rg���x��&�櫑D�k: E�3�XҰ|T:�	�K�,�]3N���N�C����,tJ��yo����ϱ�C��3DCj��آ����7�˅���'(߶z�g���Xe��O�ػ9�+ (0v.,Y �E4�y�h7q��^��f�;�"��(Q��(�@jΧ։28kG��W��%^=�o�r]���c_R�� ���5=d�[���].���s"���vsG�-Q��tI^SOk�j�>������)6jǿ�:]3�a�Ji���gpcT_��Ž�O	5m�m��8�*p[�f�����3(�k��Tk`���BܮܕKQ{6)��!>�C�`�,�x���^�F9�W��
9d�����,HI��79�u����Oy���*��>�\��5�N�h�C��ޥ��2��Ag��F#c|�a�W�%�����i盪��� ��w���/)=�	�Q�XX �}Z�6�mJ���<�1��2��덚�n���G6�����}��w�U�J�$Y��|��ٵ�����lƯ�т���<�cOl�_�O����|Z�-�Ƽ��l^�E�א��%�_��$����ѝmM:�^�UO�h!Udk��Ӟ1�����7�|ڢ��2�Zε0�`x,'0E��%�j�PT��8��I��kt�,{.7y�w��$>ƕ��u��]"�˴�`-j�@��5<�U��3�wz�#I�w0�vSH�2�u�a�:��7g�����'&,�L�d�����l��m�7�x٪ba۞�`4M�~�kߣ���� ��B��c����a��cY�{z�N�r�
��9�s0�`�ȏ �q�,KbӅ��b7ov���ݪE<�@�~�:C��v��%}L�C���{��ݑ���X��o��[4��9Y��1%��S�0�&J�����ү�g�#kI�EI��GX"�G4/�V�o�E����d-&�N���<��vH�Sް=�bxmȠ����d3vL��V	=wi+�
��f(�AZ,�?���־�?L�m!���9#<0����g�}�i�k�ŗ�`��~�&e ���8ݽ+�ݳ�;I���y��Eύ��,�Z�N�\iY�@ ��_ݒr�����u_�����K�jB���X ]h��YU`j��oý��3�M����7���`"��e�x���t�i����痘������j�xΟj�����ލ7lf�z�O�Ed1��z��ϝ��-�_󥻷�G�ZJ��j֊������i�O��=-mP���L;�ٻk\��|�����z� !H��I!B�Aq;S\Cfp�I���<="<��>����{�q��5}oV!��r$�T�σ�]��{��糅S�o�(�wy$���ovq�i�ˋ3��^�j[5߿I�Π�!ND�l�1��I�W���Ca-��*�U+��O��J6h���5t�JS�X0���u��� �/~�PI;k7|�I��BA,��cn��6"ȏ��!�b��Iw�кY.����C6h��WOO����
-�ءώ�V"P��^q��d!�+��c	�|��ϖ-���C��!k�t��;�{��G��u>�~:��5�O�Nd13�gĀ[6@���/E����B���!��/��q3�6��Q�[gor��;W&����^��D���#�������^�Q��e�U�?
 ��Z�o�e;'a}�	@ի�(��YncCB�e=6ݎWI$��қ��3��[H5�l�g�F�u	�d��҄-9$�g���'�]B�N��?�z�D�~�G�݄�:�Z�TH3t�[q����HC�=�W��j�W{����E�_��c\
�o���
|M"�`S֟\�Ñ�.H����!�{��é"��ɀR��
i��5��N;�q�L�t�ȶ)1�Vi;�?2�N��/ڇ�����0oms;:�zU�p^�%C�58���4�>z����n�y�ΛMn���*��Y��C�>� 9����$Ph��q�)�lLA헅�e:��A�+ZI6q��"�E�}Xc���ޅg�k��ӣ�RAp{Zt]YC��QSm�swìFM;�X1:�V�溇�Ri���bx4ճg���p�=.I ߯�2�y�n�!��@;���sT�S՜�>����dNS���1 ��)�X�K����ڛ�F	����8n#_��A����@oP��N?���Q�*O��&��
���F��7�ҊːqK�ޭ�)�rm��>7+�$	eK_�#e�>����,�:�Y}_6�7�[35���U�(�0��S�u:{��-<ɏ�mj�>+�8�)��E���#X����C�ά���i�X�'�������������Ł2�=�gW����_�y���� �|��M+)��9�Xg,[纠ɧ�� ��:D��(w3���]_�p2�el�|�p�����b��ruѦ�,�bf�q����/���l���h\��Z؏���Q��%$-l�M+,?�@+�
ah�y�k}z]śc���{�5���H�ؑD�ĳ�+�����
�P�~�Y#:��i�� �ſ)9��
A4wV7�zH��`'�$�ui]{R�`j|�L�&��U�iUs�M��\P	�� �[s�ы��i��9a�g���yV��n�yBA��v�J�חK�yx�o紈m�Hw�M�-�xM�����S�B��~�\L-�K��惿��i�����[�i�co˖A���9B�p[C1.�b��x��]�D���lou�;Q�.4�n�`h�hO;:b�>-3%�.�Ǘ��x��V���j��#D�P[m����/��3q�h��;I�J
C.��03�g��n��9eq�8���goG���)J`�vr�8k��'�z��WyI�����Fg��Y�.]����0����X3#��Cl���äo;++�w�&���a&�Blީ�ɚ����pgO���������vP���g�]x��(ܼw��ʓ��*���1�������m��s�1m�|~6���K���i���[Yڶ���r�hC���?����")"�;��l�)�舀q�l��5���la�O�:�-����#������l�����E=�Ẍ́%T�A��}Z�x�3�1R�DK��ЈJ��y��%yl�l�5���nD����ï�	ґȅ�%'��3zϡy����e�)����t�(�!�0qc�,��o� �Sy��Oq���=f�"�D}Q��
�i��7�Mz��̔�ƌ%�`.��
��]�z�Q�LRya����=�4�[Zs��J8+�V��^��)s�KQ�SI�n�k��w>1�K�u��)����"���a�M���p�w_�O�Kh�5h�8�(��*+rf���!93��k(~��������	�}K)/j�!�	�C��g���f�cο��:CWz��9���MEH$��7t����p���"d�k�>�b��hJ#C�ƥ�����˴@�5#��|Nz��w�zG���_'���w0K�/�
�$����% _��
jHm�V��7����ڦ������H�u��϶�(�}9���P���1e�7j���\�ѐP��d����ǂ`���7O��V����4�|�ע����秲xE>���ti_ݵ�pz��Ý�h&��1}��]U�'�h.Id�f�Y��--N��,N�Wi��8�Zig��[],'f�A�Ϛ����T%�H��!W�Mh ���'+�7�;�B�Pư�_u�)>�8���Gh-���@�.<0۫�;&��Ww�����R��v���2zh�a����=շQ8��B�,}��?�9��"Y�.m�H'�	�bM����M@��k��D��^d�!�4l����wa�s�Y�M�{U��N�j
��9�.׻{��.q�������+o�z��x|�E7e��ٷ�:��yv�^�%�C�C�nK{���,������n[�P�9t�1�S`�*&RX�$R��{�r�}gmvIԏ��D��X�GoL��V�e��݁裒ND���͋Q0�S�����ț+i�131#��	��%+s�R��T{����:d�1Gp?��!�����50h��5a�}r3W�f�w����ٜ�&4[���C��F+7�Y�����xߜ���{j`�ue���m��e�5o��y�����_��,�����[�,�ۛ%� �U���
��o�-��>��h<�O������]De�tAx�Et�������:Ź�Ӧ۰�����/jF�&��	�7����Rc��jyd��x�Uȅ���#-�)����GEs��!�֥�'}z���Sۊ�=�:}P���L��#�&H~���Б/e*�۶��9��B�%gq6�0�q���ީW�8<4������,�%o�}j�StCr��x�꼋]c�{�o~�������(���$�.����q49�ig�\��m^���И�I��_�|�����6�L��ęj�c����8�ũ�U&<��lhJ�
K�7��5��SoEǋ�L�퉘� ��5��+�k�-IٓlA�h9cI)�6][�� ��!7�c��w��"YIe��[oh�%IW��R�nJ:-������"A�^��E�?�+Z��cD,�Ŋ`���z��B�jCd�!���
;������y���y�ޗR�EOJ�81N]����@�2�/������fߧ0�E�,�6�@���f�M�u;��m������0���8�O;�:�.�>8H����o��چ ��joIum'xV	['���Y4�s~"�e�=݉2/��V(6NV��("�G���1Iu��xᄈ��_x���/yɖ���)G��N5�zC �ySGHn9�����o[MtS����?߃DL=��^�e�hW�E ��	��]���G�J���E�M�<�`N�\7������������Ä�����R���;�OG��׊�����L�ȑpJ���}b���I//5ć��SU�/��m�ݹ�UGë��%ެm8�Q�4���{l���
y^���Qn�/d*-K�Y����]�p������a�$ˠ��L�Ï��$�20@e5���BZ�i����Ech�W�ԋ���lU�)�{h$Y^;Q�;�sRaYF��Z�H�15g�t�至�Bi�c���mx"g��J��1=)���
YP2N�0n18&;���s��\�7�u���s͵S��T1;�n)F�Kż<V^��6L�	��:�� _��ZA0*�b;EP���?�.B��%����^
��F����M����K��p���m�8�B)O+aZ	 R����#@���+%Ҳ��ᄯ��KP7��P^��:1�(�{���u���(]�� ����v�Sy�}�N���#�;���YƘɘf��0�0�O��M�N����	���`�e�8zW�l��c��ʄb� ����N�QM���4*Mg�l�[����R��K��n�� ��]�72p-@Nl�h�̐��V��o��MH��	 bk���
/ ����	��@�\fC�jI�ǌu%���H�?�����Δ�}�Eś>��Ӷ(5K��H���D�|߳�!������u8<���<~�W�:�v�i�T�_�:���ǡ6%=4�Զ�U����i���Oud�;�y)j7�-�A��U=3=s�Fm�TpP�&� �Ψ�X�i�a|�{�FV��[�A���ߥ�9�?�y����F��HG~w 9,��=M�{�K��B���~�#�-��K�����;�g���P�Ą�c*&lA�z9��[�{.Ѣ�� 7X+ ��A�o0ڱQ��f��S`C��Ov�z���T%�4+��v3^OV�G2�F`#��[���mM���è;�%��m��3�;��q����3��K�%GbF)e����8F5�'�洅�l���d����i�jt.x���D���y��3^z��q������ʬ*�Ne�Aט�$�|�*��!]�������g�,/�O�:���Q��9�l]H��#�xwX��Nh�E�z��F���ǄXmWlՀ, X|�(O��L�f����8��6:��0Orns,��?�&���;�V�3l��c��קH|5<	��g��O�u������O��2�G���OE�ԺX�x�T�0��[,��A��˫��잎�QJG[{y������'a��1�D9v�~`��ymH��� '�Q�z��o���Ye��o������a0aC�0l�S,�����y�6�q|i1��D�f>�"(�iQ������2�y��h��arȘ��͇�o奝�]�����yR4���� �=%�[5sӓ�3|��O|W�6]=s��QPIT�}k���>l��m�)�7�u£�jVa�p���� p��*_!�m�栱5c ׃��*�f����
V3�	�kc��͊�	����d�%K�޿)JcE!4&,Cr�*��R�ǟ�}��[�W55�9����ȃ�H��7�(��/��ǉ �bn��C�>�ڭ�+;NCL�CI.å+����̴�eE#�!��E�u UĨ��W���vX�_Lw��a/���?���ɾ :�E�Um���2���I���a_��n���N����T7�)}�ԐK],��)���my���0�/��?���%MR����2��O"�Mx���|PD�|N���&
Eٮؽ��(_8��+�t�<��cݪ�p5��,=�U��rhh�d!���[T�Hii����2h�s'@Z9<�Vb�'�X>ߊ�C���6T�����{t����:Z��"�7/���y����mu�h�*�->��@���<p*�>�]��T��D��-p�v�~a2{�a��|�gb��	J�]�,��t�-�6����m�y`.Z�bר���M�˷k��:�0 ��Ѱ��ǖ��px�a2�Y�K{0\?N'��
.s�9��g��폖��q"_nXL�u��o�Q��;�E2�)�4��:��v��%s[�Cqu�{>}����a��p�%k�[��89���1%�S;t�&���N�D�����hg()�I���ܿ@X�{G��륌����C0��A�N"���2��,8�ST�u��-�Ȗ�Č?Q3�9^#�	3��+NP��bB�w��5�'���?�:}!�>��/ ;0CI�pzD}t]�aOF�Z��ۛ&Oq�������+r��q�����S����64X�f��R�/i���p�ᒨ�����_S�~dm����݌��k����=ZU�M��ZPoyF�S����ʌU˹ѐ�b�eRax��LtrH��_�����z�ۋ���N�j�Ou��T7"��Yfх&�d' ��0(|�7�-'�6���IG������M�������ح��C�=;h�P�xL���S���{��K泶l)�t,B"��q1�!���ǿ���r�v<�0+��i���z�rY}e$��\�r��`�x]��_{g{��A�,-1(��+$xq��C�QqO}i�Z��H$^o�kr�I�Ț�׆}�y�h�g��?�	�>W6�G��`�8U!��D-J�ͪ�R��5jyUSJR��9���$Hk �U��.�k��I��^A"lc$�g6�9�R!�w����w;b�YdU4��
�hшWū��	�a-�*��D3"Ƥ�^�`�Z~+5�Fc�_�%Q���~�ԝz�C�R!�f7j�^;gͪ6����t���r�O"�1io�v�%@l��/�l񍺯�� ������6ݺ�Q��(��;���.�d���լ<�����U~񹢽�����d5�u#����o���'ג�	v�:��b��"es%*݄-�ډH��.i���Q)��"��#=Du?�E�>̄�#K����x���\�q��Kfz��&�t��G�n��Ll኎ot�h6��߾e4=4�J�`I�W1!!�CP��{[�Y���%�9뀴�MX��`I�\���ˤ������q�W�_zɖ?��RO�~� -?�x�ג緹��.L�C��l�S��ͳ�2��D��/� O�};�J�mi�ŋ0Y��ب%y�=8���4I-��6ߣ��q�y���¦�n��*Ȫ�Y�X��J�|�����$F���'E����[���ce0��MZ�'Ɩ�B�E���cC�-�TB$��8&�U�2{�{oYy��QI*7s-�F�/I�10���,��n �i��4�"�x�@g m6Ŧ��=$'�e��2	�inLq���I;^�sʈ:��M����V�Sr9�1V�)�׺K�{���S��-�	�����_h��A.g%��U�P�4�?&Ԕ��� ���~
[cPF��S��5���'KHDU�yw�h�;��3�+�r	;_RA��#Tf�f��b��%��N7j�XkV�,(��NT�upv��#�;�[)��n\���c��k#�&�LRa�Ĥ`�t`l�w��'����@�D]��(ѹ3Q�WD#�t���?$��>� c4��ɋMa���/̝g��к���
Iu�0s�ބ��[z�]�q�p(��lSu�ۇ(ӹ���X�8�(�Φ*b�W��/{5i�>�����\}#��E���Ǉ/%Z,��C*?q�咀�wίOb}pN���D��$5�n�H�T9D:
[�IZ��OV���Z���%~v�:E\�i���O/���S�Q`A4msB�0���m�Z��u_]�j���\U�Qs\_����?� 3D)�����i�a��ԃVn�VBG��&A��� 
|���7y�ǥe�3�#��w[���c�yM�@���HBl�=~�-v�K��&�5�=�ci���j��c�eA+i�98�J[��!.*ꮇaS�w�O��o��kQ�a�d�g`dUO���t�N%�Z_�M\���$V��`��#��[�ܽ�������";��^@I��ʨ3��;Q��o���.md���{G�-)�<e�l��8!�'sm������돟��w��.�N�ݿ)��T'3�C�y���Ҥ%>
�7�\+���!W�����8kt���g�KWc�y�|��,��t�$]��B���w��[�	;�`���'�cӷ�cW�m�+�'��|4;�늪�Ɂ���_�1���5��r	���g�?l���ڹ�q�nl��>F����5מ2�b��Or�T��b��4ڪ��)�"��fUEs�{XÌ�TKH4�|Z���Uw�'e��Ե��Sy�J�Ɣy�������f���D�ZQ�Y�s�Xh�ʅ�YH'9;�zE�I�7ve""����[,��10g-7,j��v�xy��q��l���fy�"�}�Q�>��QȔ�4,h��^��7��|V���.V�@��]���C�Rﬤ��m1=�5D[�T��N!����-4��sxM�Q ��I��krkQ>��S��Z�)��Ђ�6ca�C�@�p�dn_\ ����5^�#�ޚ*���f�M��3�*�k����%V2��#Rܿ��K��*)e|!�b�CMd��}Ҝ�3����W�W�E9��s�C�Hږ�7�z*�ʃ�V�����[;#>�Ɂ��n+C��ӥƧ����h���t#���������0�:��a����w�t/ZEZ}_��1$ ���0�m�&�-�>����������>���br�}o_��FV��5By�����s�ц-k��J�`�p��ł�-��O}RZ����!8|�J�W�1��OEt�н�r$_�r,��͏�٭���q{�KYs�g�U �h�Ed|'����c��~˿��2���dZ�*��Q��';�E���vT�Т���ò�ն���7��M��T���$u���0s�e�-�`@�#<�D����؉�q�~��@"vJ?2��a}l��§ѷ��@�x��,s����8�q�2�=Im�ʕ���b�$���ْM6"�k���k��W�6("2&�+�a5�Y�p'{-�Nb�I
��{9����q� �Q2lq=(l�8ƀPv�o'I�ͮ�E-�(�z�:t�{v��%CL�{y��b[�o�쀇�[e��9�8H1���SF8&���m��3��(]rg�[�I
�}�:X��[G���'�L����|^��N=����#`)S����3� ȑ�����|3���'�7	�Ab+)#$�5�}��&�0F��Y?}�!߉����L0����{}��{�\�0�����O:�&j�Q�u�k���h+�JL�����V�u�髇!��֌D\�֫�C���|��_�2�����ǌ"��yp�x�dU1�� /]oԺ|�I���
�Egj˔�@�ǚe�mmx�4�t����B��8����,�f�F�)��j|�{�п�7}e���nBѠ�	d�p����N��-§����G���KCU�����s�gx� ʲ=ֵ�P�yLL�7����p�%R���B򆯝B�v�q,W.T��zL����<*�c���ʧ,E[�?}`�l*�}rUA� ��]�{#{B��6��ǻ�(�=$���u�qj��i]hċ��^=!lI��Q�2S�4���%���4������R2U��`;Jg�.�m��5��\S%��t�o�� ���aP�kheBI�A��jc��?6���V?!�2L�>\w�ZYec�Q�h�@W �&��u�-���ϟ��"�(^�[���K+#Qc�ޯ��a%������rC��!�L��=�;B�qw�ʯ���o�l�A�O��-1��^���@G/�k*�U���n�滿��A�6����c+f;�e��1���s����T�d�p%��4-���zâ�)���Jo��1'�ͪ	�+~����$�B�eM��H�5��̓k�0ս�I`��.�^h�u�z�$��>�������-��Ɍ?����;ā^zy�%�o��G��"�k(���tI��+����=�1O�[�oW�������H�� E� �n� �M��;`DK�\�֩�_�ɩ����(�:V��z&�R�?��>�x�Md̹�L���G^M�0���-�?�#/��8C��e͞m�]����!F�%��8��14��X��qX��[�yT-6���un8 �*c*RY�|���7����$�q����v��h�_e+�R�ZzІ��XE�g=ct���0�<���^+cZ�{��>Y�L�Q�8�s�bF���䩃1+���*�%�)�ip���{x�g;��A�!=Ƙ��5+2��fng�<H�;9�Rs8��m���{^�) %S-�1qu)<�_K{Z�̲��l/@	�%+�I�_#N�AI���X��P��>?a���"q��@�7~�
N�F�3^�C�	\��K�_��P��cn���]?+�%	V���p�#�3r������R<�z��p֬7%���n;�0H~(cq>���u$����H�on/�_�sY��3�#	�:��j���v��H��.�B��C��x!9�Y2���t�.H�W��a/����Ƅ;^ >���ЙM��]�*�Jg=�����% ����ù�G���y]0�$p#:�l����B�
�7���t=��e�e$�b7�-��c�/֌�@���U\� � C0��%�[]�>4C?�g#�;je���	}�v)�����,X\5�	aH�BWD��6���4�҉k�d���~~S�&:�a�i��e(��Z�c�l�M4�1ڰ��H����TuZ�c`�j�uܦwNbU3&�s7�?���lڽ� ���Y�Ξ{i9$ya؃1RRVI�q��Az��[c��|(�y����e��D�w�����K.M~%2���B'��~,�-�`�K�_�p}�:���~�\�z��c�;�AF[t9�:[��.G���IDN���֔o�jQ.f$��4�`��CO�{��� %��oǨa���^V�)۽E#�$�[�������y�;z!/[��c�v3��M�8�
_N�)I��rGس�)��_��608�6.'Jڅ(���ݒ؟W�d�2��.��a�:ց�/IF3��I�����zc����\���w����2�x�Z�`��th�\g`�h˻ٮ��_�6��o�]I����w����-�{	{��A�Ӓ!s��m���"��|�m��E(rɜ�@��ɖ���p��r�膡�I?�p��S�ٌ��l4���c��5rTέ]<�O�s��^��O������E,�W_�E�TX���T����7y���Kՙ�����V��}�J}R�y�6��ϝ�����D/_��4h��wv�υ�#�'�D�z ��,�e�q@�pNػ%v��$0b,�1f�1sy���qr~4�z�=f��"^JQ�Y�'��v6�� W4�W뮇_q���&]��>�b͔R����j=
f�[��%����'u�#i진s3��Q; ^IJ�\kMVf>�(�Fh�)�y��+cI"�a3��
p��A_�Sf�r�5YC�9�*\v�f�d���3nkk�2���9���z����K=�Y)��!*��C(P�^}�7D �����QW�.�9Я�̾�H�-�7%�N�e=��C��g:S\>����! ~���C���a�r�}a��Q��#OG@�����h~��UHa�0v��E�wA��/4�ub����U ���lm���(������װ��Źռ�8���B}
��Ao���z��h��!.��L\��w_ƛ#�1���(e�Oص�����!ǜ|F�
�2`X�XoIE��!\_� Z��'o��>K�Y&��&�&�4U��Ah<Nd��ӊ��~Aة�������}Z:<(�L�'w8� �r��u=T�9��}�߿���p3��q7�	+�sOa�a�u����u�ˠ��-tH"@�_@<&C��l���/���_��/�v?5q2K �axT�`��
����,��L��B�������m�;��Z(bM���M���ktZף��5�r�}�Q��taP�Y2/{��N��G
dz;9�Ϗ��p��qX�NEɀ+�ob`��I�E({���l:/�v3{,%i�C'�G{��~�����2���j[ H�9��:1J�S�7�&?��B����Ĝg��oI%.�ܵ��X���G Pȥ��[�Q��4Z�uNX�(�("��S�����b7Ȍ���B�3b� B�	)��+��p�,����+��B��?8�!����%�j0�d��G}CU��WW7���
��&�����A�@+讄��7���5���'���Ȣ�H;6Pw��\6����w�_	���vq������.l���.�Ṵ���#�o/O$�>���!��a�oEMde��gx|�/t(�%�����S�;�pD��A~��dOj_:��Jk7�O^bѻ�0d"��GYωMg-]�ڥ�OjGV�-�����؅��ңBN��;p6=q#~P��L��W�(���ˑ�x��l8K��N�BXOhq'CW�S��5#.��5l<��Ǹi���gT��]}[rS�i;r�}�;()]x83{�#�q��bj�(��N$.���b�q�e�i�o���b^x�y���I�B��?���ف���51��ziM�}ݖ��U$y��RJ"�ֆ�:�5`�S ̬�����Z ������[k#�I*�A�5cڰg6�2��!����t�"w�s�Y��z��Q�h���W;�>�?;�-�����C�"<�1^�vbP[�+�p�c���[��ػ��S��C��!�R�`�;���;�J$��j��c/NO{uN1�Ж�l�E@"��/1�7����@�A���]�<6:u��G%8�y�;CНd�K�����W/_����t��Lhya�Q�e�����ZOoZc�'M(�	��i��z�A�/�Re��,�z�����҇y���r�G����~l��6uu҆�*6�����j)�Hh���'�ך����z��jf�GY�W�&$���T�t��+�oѡ�4�=j�k�VaW�7C��=�^�O"��T��lM���`?��\H2��Z�^>�gyD�RM����R�wW��p+`;#�Ź���L|���"7�B��3��:��/F9ނ�jz���m_�����;�\��%��8{I84��8��$1��e�y�z�x�Ons�*�ɞY�]�n���V��	$<
��ts�X���3e&J��:�Z5�����EwK�c�e*��~���[������{F�Y�\Q?gs���F9`��1&��υ�3���i/&����x���gv�)��/�=����82`(n��+��;Kns@r��,�
���,S��1��)��pKVY���Q.	�zݧ�_�� Ad5����Pkh?�~v����
����
�XNF���`7$�K���AH��^Yu�S�+���	qٲ7aH#�3��ܶi�����uqs�Kk7���l����(>�ʬFu������/��*�����߲�a��#D䅂�ߘ���*��D�#�]&پ�#�S"κu
�1PP�)_?W���H������W� li���{M����%pSg� ;��<t�@��&"6Ô��Ѿ@]�D�p��l	�����F�Rc��N'��޼��aybҸ����/1�����2O\s�����=�?%��ȝ9w?'
���W���yy}f����W��g��5�H�PQD��r��+��OO7��[�q�G~�:{�	i�p ������6b4c~��?7��E���uU-%��Djh�����U�O�s�0�m�u�0 ���3�����iTua�y'�V�V� p,TkAu�߶ܠ�7��y�J[%c���w�w�ՙ[My*��\%�B��q~G9�-�jK]v������ռ]�y`��Ւ-c[��Aam�9.s�[���.�#����I����woaK�QIc��Z�p`ԣ�O''�����%�\��Vdp�V��V��#�y[Y��>f���6���9�;5}�v�|�Q3Z����z¥G��$E��\�G��U)����b��8���'��������Y]��@���_�.ɀ�ݵ���
�53�$��M2��Q���i��3�����ޕhКn���uMg����Rx+X��rf\�W���\�]�e��Twi�e�@��s�����m~�ͥ<m(K�y�|꿧� Ƅɷ1��U���Ǹ9���Er?S�����?"�i��٧9�l�w��?�X5*b�X��O(�����jy��&��أ�xE�6FX��T���z��a[�������ɡ�J�oy��T��w�X^��,�-D����e�Φ�>,,���'�m�z�4��G��e�ʃK���`� 2h�0]wr, ����R�y\q�8��U	f�U�"�6�Q��������(��¾�"l�2��L���vD`]�,���w�Rex��,�l=���[�2G�6�g��7�	9zG}�s�.�QV��I��k(a�>�,�ᕵ)�ZMǆc�.	aN����p]��_��@��
�5T�~ה��*�f�w?W3I��k��[=,���uL�K��L)�s!�;C\pS�P�Ҳd����lWf�69���9z�H���7`g� ��P>�s�ъ�>����tC��0����x9v���4#

������-������%*��Sw��Z/Ё��gQ�ybS �Զ�vvmQ��#��ZՓڒ���K�4ɬ�f���a�}�J#�<�a��ҍ�#9-�<	^�|�Y�Ѕ��Hj�̆��#i�O39wB���<�)|�=0�/�C�E�ai����_I�G�\���]��� ����z$UV�-hֲd2��E	����+�t����䘞$��Z�m҉G1'�5߻����T��XI-�9}�д�+�7@9(�.j�ӈu|?�����ۈ�-P�@�Z<��;�o�����t�㣾?�vz@�2�r�as؉�x�N�=;[��N<,i-���������s��m���?b|ޞ1 �M,/.kO�}��#p�K��Ό�����ak,�Y|c{�.?N��
�-39��}�'wƏǵ�qs@�q��o�����6�E#m:�E�:�nvNo�%�a&CJ|{��?ݘ���L�6 �[�/f9�ֵ1��S�I�&>�$�7��#9��K�gY!I@���0	�XiRuG[��]_#��ɿT�w��INsX|��o��Sa��i-Fȇ��ĝw�3th]� 	�hO+�(���MP�H&Q�&�Z���C?��!�ϴ���0�"!��}�� �RZ�k!��W�&�sP�k�C��K+#3��BC۠{��g&gQ���)l�ÿ+�c�!잒y�s�r�_d%��+���IԌ�2G�{����Ug����8�o��¿}!��XH�;|8�J��I�Ae#��xw�t��}�_�n	��c��R���yj������73Za�>�����d�����@��&-��p����G�%ך���������\�v6.=�nP{�LnL�7���/��b�GN4�% �B�G�q"O�
߯����#< �X�DL`���N�=�}VIv��r�$��V��]��{�^������8N(�a�$��-�to�q�	�iS�܋z-�^���<�WI��4��KT��"��#���/��<��g�1|�U\���<J�բ����5�QpS�8������ ��l��kޠgIEh�A���c���6I��b!򮉿�8Iwl��Y��y�G��hbq�Wv�ʵ� �-֕�U�s"���^������+��c0���ضJ�Ԯ��CPc!�x���v;����z�����e�ꗾ=�O6O31����!�@���/l���û��n������6Uq��¤x��;~Y.��4s��ݮ�M���N������*�fC����F������o��v'��	ǯ�������j�;eD�A�u޻�X��B���ؽ���۳�5�.u�k�P���sV�K�	�c�ɂvo��׾:N�z�8�eWxG����?����t?��J���o�e=c��Q�WBsD�t��&����c󳶈��1�TM)�m`:9�\��z�� ��(�9�����mǖ�4�R �ǁ�«�̭�ý���!SL�i�����}TΏ��5�//������9��+gmڧ1��N�×�4%J?>8v1�4Z�8�g�-���vyJ肛S�Yn�Pb*���Y�����!����z��J$��~��<N������e!�xPZ��4��E�Nc��P�M��r�����#{wiY�"Q���s��Ft9%��1!����⇟�miJ���~�Sx{��g��1�w��=d��v�2:�n�Tb�;�Ys{��գq���'�߲S��1��)2�K1x(B�ڢ��	�����_�m�A�G�NePF2�?׃�X�?Oo����
��F*k�9&���K���_k�Yd���0+Mq	�F��q�#�Sz�ҙ�38��pG&�7�_ ����&�(�m�uAߓ�!J�l�������.�i���<�#@!������������xG��9�m�.C�������d�$��WU��*� +��� �7��:?2M2�� r�g�a@�G�!�[�M�����o����]f��p��ldZ�۸���mR����ӹ�æ۾bm����s /����f��M�,\���ּy�x`�%+�4ک?��^��e� ?�}�'����Ӣ�5��~H�~'DKr�z���j���aF>�L��~ɐm:�i�x��8�Ы���~4�.��矾έ�+R�uP�UǍj#���:�U)��s�iҫ@Z� �c:�ʋD�io�aÃ�y�V��B�ڑAp<��v���,y�{8���´w"2�4 MtO<��?B�)~b�N-y�K8����P8�p��tP�0��c�*A|�9��[��3.��}�~1DWF�`�o�2Qd��Օ'`�sOb�$�E�L%��$�^�/a�V��Ѵ�#���[����������/�A;��[��dYn735�ÔP�@PZ�a���0?GN�_)�vͼ�YQ8��s'��υ^{T��@�`��5.�I��0�9�� �3J�ӕJ,������6�����.�7F�Ć��j4�	���gޢ��8F�є����)��%j�]Z���w�1�:sV�������H�!��m�*���|E2�뻃��Ҧ�������ٶ���r��A��b?}�@��T���l�x��^�דA�5��Sn�O����}Eޅ[��\��!��ͱ�ED�OX��T\��íݡ��	���v�e�Ύ�}J��1y�P����Ho�G��D%����	�8�bᅟH'J��zv�0�b�<e�p��&,y��
��	t0XL�,{�
��ROy4S�qhh�0,�f*�>"�CQ߾��bF|�el?�Ԥ�MHP�uP��D��Q]���B�R ���Gu6= '�[����q`	�]�og�rLs�ϿQqpCI@��k��>X��|�)�[���w�Y�ai=g�|�#p8��_V��R�#5O����!*��f4aI��Z3$M6kOK:��`�෈~���FK�%)��! ؝Cއ�����mA�w�h!gW!��9X�̴aHk��7�1t����}@�������>)W.�E���0C5c}��u��s1���#��91��a���˸��f�����w��-/����v��* ���1J�m�;��	��"��M�&��ů܈�A.#@,}@�-�7��FK��޼��W(���b�9�2E�g���O�������Ws�|<������7YEE�	���_�}��;z�*���Oﵻ܄��z�U�hqh�sd���� .X�����)˞4�_��Zp��B�q'-*2�vɱ��dT�.��3#��t�����{<7��E����7e7u�	�_����-�w�@�u�<�St�*�����4��o.v�k�2��an����7����~�ɶ�,�ը���"�_���m�}��gb�W8�Ls:M��mk*F��ewk���Ji3ĉ�\S�a�jY��{�_�N\`
�c9�=�ׂ�9����q�CD����"o��\�u�EM�w:��-vi��%_�C�Р{*F��3���쑜O[�7(9�ո1�S�{E&y���K ���9�Qg��I[�ܫ6�XD/JG� u��ޢ�9������aN�-�����iS@�ֵ-Ȃ!���t@3�4xcA	,�+�['�����{��!���x?�I�!0+���0� \�}y�g�Mߘ��t.��&�	��Ir�Z2E+^�%��nZ�vS}�g�"�����}�>dm՗��\�ے*F�mu�_�ΈP ��������"���)�U�?��mlo��s�z����6�����%9���3e�S$xrԃtޅ��sJ���D~�f/���� ���jM�ߙ���7�����oo���d�����v���8-�ߥ�[�G{��|���,�X���T��Cw۱�=�^WPv<L]����ٙț��%O�"���`3B�`�q{�e�6ǫ0B���<�6�-�����,�B}Q@�;��r�ƪ�q��]n7{�ꢳ�:�'(�#�$��/��q��vi�ފ�Ud`^��A�xI�<`�Cx�e�Z���/+6������e��@�U���q�J����N�5V/|S�ŋ�%�>�F� �!��rw�k�n`I`��A�/c� �6�}�'�!��*��w'Y�Ua��ah=T{W��ʵu&�-�Nϰԓ"�s�^IF�O+�l�ckZőS�ر��	ȭC�K!�OV��;��:"nʀ�'�`4�lO�H�1���bv�@�e\/�)΍&
�����g���oI6p�n�=D%�wW;�À������D��@��^A��������y��լ�ܚ,o�I'�=�	�9�
�B{��cYe߃�pY:F3������g�=k�ێ~O�yu��(���Oy��N�~ح��A��p-��u��zJ��`hKG B��{����It�R�%}�ߪ*�=�+�L��W���/�t�A4�E���/�l�LM��Z`5��\�	�ːRɩCP}�]�a�˩�+�R�����4�~�~�b��/Lra��زڷ�i�b�0 �/��m�i�����mU�m�����M�%�n8q94��X�"�N�ڵy�u��.ړn�(�*4i`Y��R�$T/�h2T�8+T$2����$y�ο��9edef+c�Z��!�3JEmroc�k�@;�Op�9Ot�-{�
�Y��Q5$,s�V*F�2J���1+b�;:1�Zےie�g��G;xVj�g���'/=cN��p�2���n�5����;�Rs���>h�� y�:��S^LY1)�U�K�;}���=�r	����Z�_T-dA��c����P!�?����vG�p�H< 
G��FE�m��
�-�K4E��w���T���	��+G�	��3-��#��v�R�����k=���7V�U�v���ZK(�ѭ@Mu��y����ϧ��v�(H��L2��#���t���b��͛���ᓕ�ٴ���	���0׊g����W�<�`,=�d\��� �#s�u��M� ���ygN�%�6��v�Q�J ��G��]��p�l����s�ʹ�a��D�Ӕ ��<�b�B��+�/�R��q	8�h�\iY�ر�fǳ� %ƪǝ/]�?ݮ\�l���$�}\����g��ݱ!5R��H���D�
�5}?��ϸ���'*~/?:�2i���&q��﫡���4Y-개�&��w���"�uKբt*wjށ1���XU�Zs�$�{���/ �.��0���K�i�wAa|ª�½|V�~�b�Ak��l/F��vFy��QC����wG���� Mo�����BX��~}�-�߂K�h�!&�����o`��c�˴A���9$~[e�.�ì�f<?2���%�o�6�Q��Pv�`�c�O����<�%�2�ǹ1i�qdV:��L�#f��[ϛ��t������̊:L;�����T��)3+������x��x��G	�)�t@�X$8���'��X�����G�h���c��.�2�ݫ�����3��V��*���@���I�>g�Ȼ�鋎*�������Q����gq�C��a�/�h���d�`��]/��
lIw������̧����#��C�.m^j���I|��x�vav��;��K��}(ʶ!A�ru�c�ꟹ?�Hw������ll�^��QG�Ώ5C5r�N7�O��Ӣ�q"ޠ�g���E�����6E�qX�iT�Ճ�h���ߙ�@��?J�JN�+y�g�G���Q��b7�D�,Z��㖯DeXt�A '� �z1>��}'�e�$��1�ք�h��0SA�,֎]�br�yOjq�ԓv�fe@�"/p�Q�~%�_� z��6ȍ���i�¯��S�]�"��s,R�ø�bb�={��[|Rz������X��0��@sd�6Q�H�I��k��E>����Q�)�|��<��z��a� .���p|_H���|5JsJ�J�*��8fOC�3��Sk�͑��?��+Y�Kn�)� �!��xC���St���������AWܔ�9!�D�/i�HF�Y7�u�6*��ʾ�)�GZ >D�"풗`�5�Cp@ޥ2��nI��b�t#������H��c��������wR�@/F}���c�o� ��l=�m����������Ah�*Q���^>�}۵0�2z�����`��r��rgx���L;���2��pO�����ry�|��������	LoE�x⽍�k_�kc�����E�[�����(!�S��U�oh�i�d�̔ӻr��u�j���yb�����Z1��=[Z'�n/�1�W�'k�T�&�����Aiĕ	�7��������R�ur
6�Z��Q��-E��@Ұ�<7���o�4&�jFP�t��v��2��aiĉ�.�K�����>?,_$��a�w�]HW����m�ND��Gb~S�g��M"��k�z�W�=���a�ߕ��6a�țYr6O{w��NN�z
5��9�����l�=�Cq��4�*�����of��ԇE�����:`�1v��Y%ڰuC�w�{eȞ�΀�����8�[Q_�9�C1���S��&����U��ٓ@����g�f�Iv���&�gX,OGѸ��~���d�
�sJ6�N�"|����s?S{�A��"��}E�S��3��c�Cj	��+���!��~�[�*��S.?i�+!K����0�����!}���H��!���;��&ֿ��a���5��+���x��q�����L��(����֗j쒯�p�h�q_�;���'B���~��G�d]#U�����io@��5]j�
'��17� �30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�$ڜ4qz^��.��?n��!�|,rn:Ѻ���p�Y������:H��{>����,5J,�1��=��u�����k�_Ř��7�7���iF3��p�ӱ�]X�k%6��`� ��}���>j�x�r#����-:-ڥ�|i����r,>N*�~LAׇ���P:e�}��*L_�F�w��Ǔص�i�L�����M}�o��a���"����)9�D&2Q�q-EJC�D��Q풋G�_���gq�J5��qh���G5�=;��Y��K�Ƞ����%��v\
�VHN9�y�x���(�¿E�+/)��qG����e�Y�N[�,������*s��Г.ײg�����˜��PNg��3T�_`6c$h�&����I%뛍={ DL��#�
�4�u8ۼ�)�`�y��ͱǗ:G�V��A�c���C�u{/7:�{G��F_�dO�dٮc�ɋKQy�o�?N��5��+���pm�L��n�QD9���'��f���f����҉�^!�j�j�����m���<�<�Ǹ)t~���� ݬ�_�P�lȐx3�E9�������P`x {��%�"]�����62ZPfK;>�����������R�c�ç�	(JrHZ�2�����lꡣ�����M��]l�g�#�_ٍ��+86vj�8c�B+'����4YFV�FmE.%|�l<��o��_�ǌ�ƺ�qSo hҿ��[�`p\�܄�K��� *�?Q?�h�O	$�*[�~�����Kl��n5��v���h:#��2}�7��Y�Ŕ����5����UV�qG��	q4oh���~��|�'?r���\s��n*�=P��qj��Aa��)������f�U�M$j6����^�C��g.v'����
�,�u.�[)���:J��α�ĉH�v���[MI�T���K�����qX$��&(H{S%@�Ԩ�ȝ���޴=<�ik���5�b�B�s�*'V�w#���b �so��n��
w��?�V�G*O�q�7��<�(zے5�)欥<Rwꆾ|<���'F��}Q���P���)�����(��ނ�F?��-Q�OL�#��V��d�+$, ���������b]�x8��D����+�_��ٲ�}k4�<A����Fv�8	�]3�/��x�)�lT�:*�so��w��Z����p�����N`��6�Jy<���ä�
C�-��
�����ӄ+�R|�1-�pע�� $0z� =�b����~�V]'�FN�b��WŹGΛ�A��ݢ�
��\��W͔殀F��+��X?$w����ڸ�A1ؓR�	�q;��o�IB�m�����E\�v�/�2��Бp�V����_�Amt�2�y?�{>U{nG8�#���k�_x?m�T۫GŻTx�
ue�eG-AL��Y�^�\ؗ�o!�?�t�'T*F�w@��uŕ�����ˋ!��0f��?�r�4���h�<鎮��������c��OIrqI����c���/MSP��>��L��c�-�3ך}̓��Qsb���C�]1�ገ����np���RM���02�b�+�����t5y|Jt���#�ݡ�R���ݴϠ�"�@�ٶ�9hJ_�w�a�a���N�]T-t�U5W�w����"i��v��[�_�ڝ)�c�� dS�*o���L(��G���py���Ec�*蔍y��fqt�=4�k~�+�p���xDy��ga-���T����=��t�F0�nCk�z��k���X�/y����&<{��6$�X�EN��0�6J�iU���hv�i�����$	,�0
y��v`���~P>_�BeO�g6�xP�;�%BRR˝�r�9��~��Oc99�g�&���l����y�=T��rP�*�y�y�k$���氁���.���h�j����3t�2� +њ��l�j�J|w���v�K�,�� �2��+��c�D0�(㞘����g�j�j�������
�y>�Y�3��� �15��7a3��\���G;ˁY���k>�+;2�N�35^4�4-��G������Tk�Z��@�J���38��A�t�Ե�D�D<o�N3�@�L�e�@O�	w�1�,"�+�={�J������DЭ�F���]|ih�d���{��9Q!�՞K�M��U2���i����R��9|�x��C�c7����#�����a��8��e�8yN�tv��lM�2x&��퓪soc�ӛ �!���[N�3P��`�ld���/�I���	�� @���1��:Vu���%p���ͭkX:�,���"ߌS㡅�u���:�,�Gl�F[җO�Ch�� y_��gB:�먄����\eY}�`�O|�;T	#��������)a��h�#\�!�����*��MTc�B�|�,)��n ���dz/@]Zl�}TQ�6[����'�����������KX�����Uۺ���,�if������5J�������j��K2�Pݔ院3yϯƄ��Z����8
�xjjԿϺ��|p���^��!��_��u�Ǽ/ʳ	�6�HJ�ϑ�j�R�!����i�F�V�I�5\O�a���Z�m���"-c�Ɩ�kv�k#jjls����Am�0�;�Oɇx.�{���k��A���m����|��:E��o�Zwx���V<�
��)i�r�ҕ�a�2�E�[�
�,�����:��m��63���7�~n�ey��z	,��M<���'�$ƀq�Ű�����;���,ޥ�Ѧ�i�ܹg���Ԇi+D�|���2<>���˘~J ��\)m�ٱ�-d�k�F!�jI�#K����N�t�1��X���%�uv�L���$����Sz$�!�r�����<:��������r��!~8�������:�b����L���M4�3'���j!��2z���ٹ�[��a�7"��%XG9۹*&�H�c��$�O��Lah��w:#3ȯP�4}�;JB<����T<��K� ��n���H���xTs;�Z	��-�-�LE��*�qVOR�HS�m�ڨ�Y�9�NK�F���d�l�ڲJ:�i�I�������peJ�,W�01��oS8A�b>E��_��B�bA�J|�{ɶ���r����}��%���m'��VP���=�E�N/�l�g,�� �l��LV�b;rxh�A�(��t� Q�'��K(���(�(���}���ql=��q��B�D��<
��Ӹ�}jJ�B��O��7NQߣW����cC�
�&po�bm��߻�RdBB��q�W�L�\)A���-�+�T1���L�d��	��E�p3���u���ZdF�1#5&v�6�w.R����/���l�g.(�bX&������l"͹��y"�ސf��]���9q儐n&�H�5�=�F�KJB	'hrC�S�X��7⵪7�j��s���%����@�[r3M�פP􄛋D#r�K��g���1�䛕�uA�K6P��u���Z���̛�fq 5^�)�=4.v&����]��%D޾7�k�U��)��s�4�t�%�&[WAßd8���W�b���n!&TsZ�t�f�o��nM�nG��=����$:��cqN������Mu�0"�C��}*��'�����3R�� �?��@����D��4s}U24'~��,Fٛyg(ݸ�	��g��Q��4����I^�����rh���1���Fa���BPRt��s�i�ގ�}�s����]�wK=�༉�Ra�T'�`�n�-�s�솿l�����x>�m*рpzN�Fك��B:�#e�e�"�Pz|�`�g�B��v��t��jsB�A�EތTV���L>��޽�Ԧ��ެ�|A�j�( -�i�i*|5MAq5�.�	9��]�W���i��s`�;E�.�RwC�/Dp<(��A[��л��'r�P�M�C���Εv�TT��g�g7^[�,P�!�u����>JAZ���c܋u<q@B��F�D�~����[�x��Q��P�>�Ӽ[�[9���4%�J�� ��"��I޹߈�L��1���JЩEeɖV4�u���^�+�������o��� ���"ds�.����^�B�C���phqϏ�r3���wY��~�G6�0@\f��
��G3o�z�+ƭn���e�y�J����T�����I%����J�V2WMCV7�"_]/Q��w��w���$�4��[�-l5���3�_�&�d9a������][9W�u� �;lY��x��'�uݍ��Ƅ�' o�9Ʀ~��wT�:�;	�V�͐Xƈ!����Rؕ�n��� �NR�ׅ��`�pe=z8$P��폆F.p� ��AEv�u����W��ztw�[��\�ʖ �+�+���k��T��V�H��Oz�l�~����<+�2��_��0J�C��̿�+AjX8(�$bb��� �%y>�fi$E��.���������Ec�J]�s-�סQ{\|#��.�}�5��@3��_8�h^�)\�'{�
D Mǽ�H�<�ȔMUT֖�3�����]W�@	y}'��g=b�FG�U8�&F��'ez7&p��/�/������L�G�B�� ���.<>��]���/u4�s�����N c	b0�ʅ��<XA��bɦ�F��s�kD���	���N˨�"U�Z��㪰���"�?�&{5<��@�ǻ�~�o�1�P�r�{��h��5������ٽ
���D�+��(���ł��@���J� x+w��Ѻ��P�<�}�4���Z-��JQ+�Ѝ\��b�D����Ŕ��F�r�����(�S_q�2�V'���=I�F�6<L)������_I��q�A��_ЇC�H�`-�K��YL S��B.�S��/��X�$��7�Km����/����\	��%p�OfWVIX]��}���H�I8P��a-�W��%c�K�ʝ���}��h���u�����b$���u�cE�V-Y
-��]���D�C�Q��d���w�,YH���[���'T��M�}���f��A��ٓ������*M`��-�����f��BK�v�x�mȗ��K���a�$˳�,[8�#�����t��E5���:e�,8��2R /:��������Y�� �R5r�_;ߒ^�dg�"��cޚ�!"@�^,���˗t��=fg	��l9���0���A���ǧt�;�pL���������/�MA	c�4!�!nJ���ݡMΙT-��D�������(&3���m�X��Qm�:,
!���h6�֡(l'M�q���yw�*��{Q�$�L�6-s�PW٫ń��O�Agg�2�Ht�N��|��B"��v��zy�/�}A�3I��h/�6��Dau��)�3������3���~�(���Z���A��s��mC�,�0�7�6�(Y!M��;��tDň��wc5qr���\Kf�O��Ʈ['����P�L�dE�UA�n��3�����om���#Ͽ��Լ
�!��f`}s��d	2jܒ{܂e��r>nm��M�w�6�l��������{�����F�����036Zc�x�H��2gR����(�1�A�:�����~���_[]�}��{�U�4�]�"0'����<�%;�����]��"���/�).3��7��}�=�@��O�����j�ٝjDH�e3�,7���<����~�ݢ��$����D���5���NY���W���o�����֠V��<{�b?��f��&��+��벰����<��G��3�$���p���=*���א���Nq��'�*�z��_��`-�R���3�S�ťCs�aԗ���'�/�U%� �,�R�A���{d��|^��7Tq�8��"�V�y2%�	��0�}<y�Y�:�������Q�ȵ>�5�L��g���y�&e��ZK�����S��VT�Z8Q#o�t�Kn_�7�!�`�z��.cS�~���|�E��d`��-���n��`�����>%��9�Q�Hp���O�6H-#Tv�59�e&���]G��
���t�����N��k������5\�T� �}Y�S��&��GѢ{�	���.iЦa����5�n�mϸ���b&k���+nT2X�I//�cun���S�》��a���c3i�:��r�@��4�֕�X�ƕ�Vm�B� ȶ(]풜�ZLU�=�"0a��9�ޡZ&��gM�[f`�Jo��u�
1"��}���04$m��|f����oErt�z� =� ��`I��M
��|��/!�,#��N�Zt���%�7QA�I��g���\�ﴚ���#c��$����,��
��q��h~0X�!�@J^#t	S����u�Z4��&�"��>e�0&��U�m�5Ry!Tm�>kg]��m���0-Ϥ��Τ���y��X��3��r��#c�i��;�䥳�������W����ҽJ*��Ӯp��k㞆�Ǧk�$x���B����Ҫ����o��Xmw%t�H�^�ϭv���.,��%)���r�-��u�E:k���}R�q��r�v{Tr�~J�4����iXA:�ܗ�΋L���,N��:���ק�
BΌ^��ً1m8�aKl�"�R���R9��&�\[�x���hO�\�a�jd�	�3�&��F��;X��<B�~����� ڼ��,&H���銗; �+]���(LWj|�V�
H%�xm���Z079���9˃��:_���D���;T#���6�Op�}S����֐����5S��e�Ԡ�W�S����AOAϢ���'������p������!|�m�ԸV"���O3��_�\�P�9�6ӊ��q.����V�;�R�hg�ꇺʹ�FH�Q�����{(Z����SӴ���}�����߰�x�-��BD��2qJ
½n���N}��TBO��O�k�Nc��W%s��"�
��oo8w���2�d�|���W��\��
��#�=��16�/�ކ0d��l	�q ����Շ9侽�AX|1u'(vs%I����zO��?���9�t:Z�d�g�dp�>���gt�̐��`]f�;�'����&��ths=��ت�y�	��^r�S���j�����ZX��8�Ia�@d�yrK�׶$��Ek#�I���Z�4ÿ6/U�s���'P�D���Z)���m�oq*cg^��=Ɲ�&�|W��rO��Ci�P �k�P��;>�s�+�te@&-kl�-�8��W�5����!8e>sU�6�K��AҮ����M,񲎘s��]s�6s�g �q����=���U$MǇ���#��e<�'�.ŨBksڰJ?�������t4�5�U,O�'Ы.,؂�y9S��_)�+��أ4ulJ�X��U�a�t��D����	hF�aӷi\Ru_�]>$��f����ls������\�	Rc�|����E#ۦ|�`�n�-�eS��5����
���}�e5z�H��1'Bz�#w[�t��z��92���M��.��N�B̗��W�T��C��5�r���������b��<ʪ ?�yi^Ԍ*�/���RA��.G'*����/�WW�SiU��N;��d�{C7��Dv�c���嶔���'ΞPĴN�0�-Chg�s�ӕHT���'B1^��aP���u�K��I�lA����3y����N���}V�P_��������xO1��W��Pz����I[��r�u%��8�R)|����I����x)�K�.��H�ԟ�W̒��}�u!x^�O�ٟ9�*������k�"!�s�����x��^�ڀC���p�E�n��{%Y�1����0ҳ��sT��Y�k��ȸ�??ڸQ�M݋��Jc���2��
���%�8	J�(W��VI�_�@�}�S�Zw�A�$#�4��W>l�{ߍ�T�_<j�d������o��9������l+	���y%�����V��'��9p��~z�&��M�:��_"��Z�a������:�H�	 ����|;����e�+$b����.2� a�E�r����)���zF�R[�����������Y,�-h-� ��Hu�z��eߐ����+����������Ǖ,y�Q���@X0>Сv*�b-�{��"yP�\f���E�j�.��폺���%@0�ܡ0s���R�{c��|��$.~m�Gz�@��_��~�:�2)n+�{L� �v��y��p�Ug�!�4\`��Y����z�w�yI�9�c�X�U�7�؅K'7g�&�"E/���*��RIG�l�]�����x<�k]�Y�/_�4Hy���ȍ�`��	�$)�V<*�D�t4��l�{�l�n�="���z	K��N�����WKZ�*,�����{��s{G�ͨ�AN�MH��Ax�b�b�� �h�w"5��7��V��\U`��]s�Ϗ
��T�O�ᥥ*J��U+)��g���b���ڎF���S�3�6�J�,��<�\#�"��m���R�Ŧ	.������i�ݡh(��qa2r�
��&�I	^C6�Eu�˓�Xi�_[�Xq�����l�C�1a�r6�K+zL����v�㷕�s�/x�4X�����2�K��Ы����/\�%�Ayf�֩X/+}��(ؑI��B�po�iY%����\���U���z��7̀�v[�����1��X�2c�N��O-ìl�A�-���Q��W����~�>�<��p���c�s�}y�f�@W���NxThk���M��i�- ��«��/��x1^�E�J��v�Fri� ~��%Aܘ���z�Y�AZ��N;!@0�a�c���ӟ�>
���ǧի�(m�Z+hu���l-D:A�������6}<�*����]��348�1�{�9B�u��AY�(\F0d�%��	��o�-�
U(�]S+Sr�[�"hN[���\�F,�����@� J�?��h���	��o[�Öௐg��lcB�5�Mvu�h=�΍�����Y��������5����gt%.[�h��S��u��F��'"�����s�a�-�=��4�Z�K�a7��������%��w�'�;���!8���wv�N/�ۀ!�o}.p�����:o�ÑU�Ĭd�v^qK[0����f������1q��x�BݵH��i�\lԋ�m�A!��W���l�	�	S?b�����a*��WҎS�,��b�Bo��sn_�aw��p�yg�*��L���<Ȯ��5\-�,	�����w�v�|_�|ɪ��jEMQ����W�\u)�:���KBT���?�OQE�f��6#��̢+N�+�9,#Ҋޡ�����T�4Y�>8����_e+t�����}�q<$��VFF��8w]�Sʽ�|)� ���b�sR��x&������q���߉J�`���̈́m��{�=�CX.�� �oߖ���u{1��p�Q��C��z��Y�e�Ñ&I<~T��]J�sFтȧ�9Ṋ�3��ک��]�
X�� �	/%FU��+ϿX��w3Z����At��e��dc�$��,��m����l����Œ`2G0)����@�<�B�m��N2��$?
�~>���G�̓�F��8i�_[�?#���w�T{��u�g�G��JL�2���*�z��!���>+T-x���څ�\Ÿ�h�aW��K!@G�fG�T�;�r�����_��x����*���G�}۱uqé��9�&��	�?M�� ��Ձ���˼���-�氚@���i�b4�JC�
��$�X���k�q���I�� W0Uy?bZǣڕtxU��w��I�u���B����r@��<�N��Jμdf�a�� NG��-�S���w��ˉeks�5�[���� ��cW�Fd&7-����Q�(-��G8��p|qT���c�2v��4���t��=w�~A\�p�[̕�)P��aP�ʗ�3�s��=��M�FI��ѥN.���Ө2�_:�/\��=u5{_�Y$�CnE�?�LY��i�kB�K���J��\$j�ɓ��hA���B�~��:�%ݛ���B6\u��>G�B}�`���\"@~�oc�d���ǯb�.��f�yQ�P˙c�P�3�����H��܋��Sd��e��'�j����V�)2k!>��
�O��jG �w�O�vA��9 ���2g엄�qDs�l�Aaz������;��Ƅ/��{� \��Y�'�R�##�1�������1@�^�Gu�Y ����+>�ުi1+3ڄg4}`悔�������K�@��n�%�U3�E2�dbs�WեD�T��wNփa@�u�e�d���1�Z����p{d���Qұ/��GLLީ�K� �h ��FA���,�ыK��{�X�Z�3�+��u��9�Tx�zL�����a����1c�����k�eҿCNZ����H��u��1<�����]��Q���NfA	33�)`�W)+ʨ2��IjU���yZ c��"C���{hu�N��Z��*���:��Q���bq����u:�3:�f�Go^�F� YO�>O��s?�hYg%�~.M!�V��\hد}VB�O?GT,��5��̫�)�K���\�5��FK�lKz�p�9��aA_�u)[Z`n�d����z��p�W� T������_�������Gֱ���ǈ�ݳU^���^#ݬVe+��%U5�7�S�
�_j��)K�b��l��d�&y�B���Ia8-�j�}ϝ�b|��{��k��������8ʼRB	��H-蠑�R&��	�(iE;VN�b5:4����!Б�������c������k��l�i�}�$�0 �Ol?�x1S�C�k�U��j��	�.|���E�W�����x� ���
I��iж���|��E�P�
�ʈCh7y�UƋ����h �7������+`,ז7M��2��$骳qi.���J���z���,�O�	�;���x��f��l��_g��u��>8v�˛c�J{� �A������x`k��g���+�ƴ��s?��K6��=+X�V�%%]��/ֽ�g�N�?l/�VkH63NrR�����:�����br�7��U~����FTM�9 :T�2��W�Lzz�=�?�6�����{�/����<G9>�a<��"���(B�9>�&a�z�B�6oO�h^a��V�c-3�쟲�Z;��T<ө��S[��" ˣf��H�I����V;r�^��B6����L(��m6�V�`�HV��m"<���9������1�f�xPE��UL��l���o>陸�p�e����������{S�,m�������4�e*�A��y��!#���]����[��4ڎ���mJ�;Vӭ�� ���P��mG`�j[/$����gz���Vg[�;U%WhX��˕��wu_QP�V�s"R(�͎���.���z}�S��-���FL�~|�B�2C��]
s<��'}��aB`��O���N�YWy$P؆]
{�*o�v)�����dE�Q��W~��\L���3�v���1'tv��UMd�#	�H��3���)�nr_)V1f9Ev/��zOC� #l�[Ч׾���E���U",�uA&o�Ĺ4�_�^�����]Рi�0�Ǻ&�p���4=K�̪�0	Jt�r�#�Sw���z�~���J���n�h����N@��+r���ׇ$!���#,����x�pЛ��UAĢgdW��P������Z:ѯ̞o�q{�{^E��=W�n&z$���뛱�av�k�hR�\se�t���&�3���8���W���L�!�D]s�L1��BS�򻁄�/M玩�Ѐ�����ت-q@�XډHJ����M�>Ŷ�õ��B�'l�^��d>�av6?�����w����4�TU}q�'A,i},y�P���BBҼ`����4����o;���ݥ���c��?��?F-��G�Rir��l�܌c�ALYsv1{�����/�8��M����Z�Pli���mO��+�քk��8S~�TAZN(*��"��[���b�Zh2g�T8f"øo�M���_�"R����y4&�8�R�|���ڶ�oG	#t8�|���� a�I��t
(,|B(I!��f�f��A�u�873^I�P���S�R���z�b�x�1 ���1�he���[qb���%�	f���R��h�I謵�W�уے�\Ep��΢����uYw�^È���o�b7������"Yw����C����^�	�C΢�p�"|��Uv��0Y��ќ�0
����;����G�^�w{⸉a]���J��j�=����?F(�W�\JK��W]]V��~_�i/�%���w�$[���%�l���)�_tKfd(���𧫊9�F����lc����������Wi�Ǝ��'Ji�9�	E~���^8x���rOn��@ƒd��Sd������� ���!?#s����E�eG'�$��+��~.:�Z ���E�앲$�!��z~�7[0�1�T������%�e� �X
HTTz�6��rA�@�5+�j���������]t̉t�,�Xh�衮7�be���*N�y�pf�E�z<.������]G� s���!�\{�w�|���.�<0�@�f�_�S�r��)�={�i� ��R Č߹U��˖l8Q����,��QyG���q��Ð;�U�$�'o�z&��@/:b+�b���I�G�M��)Г�0K<Hn�]2�}/��[4�!Ɓ�wP��H�	�T�O�<b��&8Τ"��Kݖu�\�
	��oN�wa�,�VZ.՟�4�p�$��I2]{����=ǅ�T�ys�?��lh�G�5�f	����������C�	���H��-J�G+ag1��ʉ��{��F�~������v�J�u��j'\[���,
��vE�ޓ��І�����A(9��q��42��դ	�IA�46�Ύ�{��� �_��q�M�)yC��zª0IK>lEL�P��L����H�)/�m�X�I����K������f���\S&}%��f!SXg.�}UX��`�hI�ﲨ춓�ޜ%�)d�����}���f�L�������W��Đ�dc;u7��-��S�y�����Q�G'�I�ٶ��tV�!���E}��WL3}��fH>ǋ��10ܱ.���*�_���x崐�f��eK�
x5���JƋ�ص�a��9�X�����7���y �%u�p��3\�x�e� �`���[ݶ��^�2G)OYn7�q��xuz]�$�I��ܔ�g�(ȶ������ұ��9ך�E�UR�v�ݠh;�ٰ���5!uࢣ?�~�jy>
K�jZ��2ӢJ�1��85��,R���m8�3j������|�L���^�ۛ�6t��,r����	�ӐH�'!�BR�߬��Iti���VB�x5�@��I����� �9c�N��B��k��Jl
��q�l���0���O��9x%6B�W�k����#�ؽ�#�|xtEơنq7x���-�
=�liDY~����E�N�
��B�"
I�$�O���\�7�͕䜳���A,˕WM�R���$]�@q]��qGD��[��$5,�P)�}�K�����q�`��yK����i�P>��eˏ��J���5��p4���9�k8�)��X)�:A��̎�K����Xr�[%ҡ��Q�[De�,�J:���rF��zy":�G�J�VD�r/,�y�c~�T�:d�nH:H�+�RӝLd뱸`�*�M�_��oZߌc��0�����a0/�"r��-�9�-m&U
�`)p�{KO�K�a�BX���X3��=��d;���<GT��GT��H: �����H䜜�O�8;f�v�0!J��mTL��Wa�,VfY�HJ�im��ڿ��9!	2��SI�� |D�+��x��`�����ۅp��I����T�����S4���Y��X�0��٤Atf��b	���[���6���~��V������m�l�V�*����Dj����^2��R����O���QV[��;�t�hL4�?���k �Q�j��g:v(_�5�����?A}�E?��]0���g��PB��)�7��
gժ�*�}�;�B��O���N(YWm�m���*
o�oS�!�&�d9dԅHHiWrȽ\�3o�'���1�_�c"Xd��	k}�'v�ՌȾb'��p�1Z��v��^n^��� `9�D�ށH��Q�I�:��ucYH���[ٮ���q]�t�b���j&���s�=�C���+	��r���S���n}��N�ʷ��ܜ���^8@i�Lr�5
��GI��m8#�������P�����R>K��P���AqZ�ա̒q� ^9�=˱�&n���̙ߕ��ծ�k�� �^sY�tjP�&���8�u2W���G�!��^s��]������%hMm>�l��fͥ��r��q����}Qh��zM�9�=���'`�d�GS�U3x?�v����[�"4�SU�f�'5�1,ݟay��[��I�:Z�h�4�t��dzƺ'��y��|����Fxq5��ƩR�vX��x=� ��5%�s�({��l������k���<P�L�`�*�-2�P�ݼڵ�~��� ��b�Q�z���"�B���#�^˵Y�bz����^����.���'1�t^Bq~X���`T�<�I2���Q�ms��>X������� �piCI*�s�� AH�.�Jr�t1��-6WVEi:g�����;<C9�)�C���D;W�j�*Ѥ�'��P�d���^�Cʹ2�x����@}T3���^rX�P���u����ԦA�>��TC���
fw�R�]���u�A��v�xT�3������ ����[P����%ZS���50��I/IU�ވdf)�0Y,�-ܿ���U���u&դ^0�����=����"�:f���}׃^L>*C�djp�&}��Η���gY��j����0��8����$���z���ڸv�d�P-�J��ܩ7��h�L�e�CAJ� bW�9hVN�_6e��U�|�w�x$�'�rt�l)���g_��d��~�8�!�a�9����7�lP�a���D��$����A'W�y9U��~��K�[�JO��dc���Fū��f��)���7 �W�������阥�e�&�$�ѯ��,�.�"� ��}EM�3�Q�l�{z��[=e���\�Ba���W���ǅ
H!USzcp������:�+mn��3��a��4��V1m���Xu��[�Jb����yӑf \�E��S.7m���p��
��af�s�X��L�{�|�~�.#�����@j�3_h"�_�E)3 {��. �*Ϳ��:9UL�6����Y���ֳK��y2�ޚ�ÝS�Uo>�]i�'\�&&G�s/g�ɰ/4�>1�G�3�B�p�}�<5D ]�'1/Ė�4M̬�O|���	�U#ʜe�<O���9�X��>�qst����a	0�yN4�����Z���a`M����pf{��,�w�������f �'���2Fxh�iy5;�l��z�AŬ�[�M��2��|�������JB��+n�
�L����3���W���^����J�_��֭x\�T�yD\�����k�"������V��S�(F�!qF�*2����"9I��U6�����I���Q_�L�q�WͶv�pC��L�7�RKkY~L��Q��ѹ��e��K?/���XޤH���eK$�Dа�՝&Y\`]�%�/�fn��XT&�}�MX�0(I������ҧ%������y�z~�?6��y$S����E���`��=��c\cv$�-��?��>j�p�Q&���V�	�c���{k���)3���^}~��f��1ǘ�r�ʽ�)����*$I���N�]m)f-��K���x�t1�����žha`􈳅��8?E*�9�(Xэ|����O+�#�����R��б'�^Y�
�^�n�W�nRL�7_2��^�8�g�{Z��M�q�'�o,��ˮy�t��0��Sg���lй��9��5�A�A�Qlt�"Gx[����l΄(_/�LA@�
�K�\B���Y�ίt��LG�-+)�?���s!(&ɤ.�Wz!�="ImM�3,an��`_6��S(c	�M˒3��l9d���c����fe�&�
�Y?#��� �L�P��߂��y����3q'��;����I�6Ԇ�!�Im`�U���4�j�/�܌�M�+j�n���MKi�6𸀗�3��%&���G{�i��L}�'M��N�6d�N�H�Wg�Ð�21Y�������Ո/�	@�]wgf�E�;��ݵgR�"��X�dQ��/�����]"�`"qAu/��.}(�7^^'���߷O��}(���1DR�(e}J7CU�<�Z���֫�'��\����dD��&����ص��YE^����!M�{h�ayw �+u���ۖ�r~9,Uku*&�%��?�$|��2E��`�s�{x�
$��ǝ
��iF8/�Ng���E���
8D-��GȠQ��Ҟ�57|���^���m�,H�M��,X��$_X�q�������7�&�,%4��$��U뛝s*��"�J�U��+b�>�s����Jq�G����r����Sk����cx�<Y���G���DӖXtF�%[;w�%{ԭ:�&���t,czr��|��:RZ�|���
r1X�4~��{����pU�:�zߟ�(�L�ir�v5�ls���=�1qd�e���r�4jza�֝"!a�^ͮ94ր&�ab���l�O~e�aa�3��u�3N����;Z�<Ix�g��ʵ) ��&oH&�(��A;(Ԍ�2����L��#~�Vh��H��m҇ځ;H9#�ŢŪK�\`�� �ˠ5���e�!�]1p�]��)��D��ϩS6�Y�;�b����z����VA�����ɯ�F��")��x�ت��H,*m���V	�l�F�����N�����~���)���pV�k�;K<�h�C�AB7����QF#��)d(a����;��h$}������W-�t��Bki��9k�
����j;}c7�BրSO���N��7W/���3'
�*9o��V߾��(o�d{z*��&�W4w�\º9�i97�;�1����eZ2d=�	�B����3Վx"���G"F1�5v��������",�F1� -~�;.<����q���*���C��2]M�:_��}
�&���=A����	��r��
Sm�o�0E��PH���xC�^e(�p7@k�zr�F��}�����m#����*�H�f�c�]<�%���PP���zMMZ�Y���qq>�^�2}=�f�&�f����1��C����k/�y�p*s�Ntl�+&L��+V8y��WI���o!�is|5��B2�(�@����M�^��n�*�l�}S���q��"ڿW��AMn��;���3�'"O��I��ڗ?���칹׋]�D4J��Us�.'�6,߾�y ���������j��4�DV�e=�|ť{�܎+�Q�L��S�Fz#'���R_�~ۄ+�ѓ�wh9sl�^�V����gf��	�C�A��x�`��-tt�_�j��<���,���5[*P�z�{��ɏB�_#>�I��z�����p���C�K���B�'ҧ{TO��ۜ�"��5n� k`�(f�#Q� J�i��*�.��Sx�A���.n����?�W���i��@���N;~꺫�C^�vD	j[�J"�۬�p�P'�m�P+Ej�wG�C��O�z�=�/r�T����Cg^tXP��uF@[�po�A�1-�����N��9��_K�����i��Բ�xVj��>,~<�TZ�[Ry���
%�al�y$�� �I�>E���b��ȕ�/DW;Ak���˖ϟ
u(n�^rY8���K����Gj�MOy"h����R5^�C]�fpa��������Y� ��sG0�H.�Z��� ��sP���Z��o���ìJ�d�9���7}�Ή,��:�J��W?*�V�F_�>���v�:��w�!$�X$�tF%lH;��84_c��d��˱z)�6-j9P���9�Ml�?-�����E�&�m�=�'�	�9�~���B���h4a��f*��A�D�}�؎��ϯ� 
К�0.�bkΘ�4�e���$)�t�N�.�|U Ȅ0E�z9��.�1�z-��[�����G��D�_�6l�tǼ�G�+H#¯z�}��W�;���s+�]�'����Ǽ���X��α�X������b����Y�y��7f�t�E��.y�0���P�̱��cH�s<{��0��{��i|���.e@(�(@,_,����W)��Z{s4� �B�CL��wJU�o��0j�G�ۭ;LӒy	c� R����U1ζ_�'�Cm&ɋ�/)+Ӱ1�@�
�G����� �	�<w�]A
/��x4Og���w��'>D	[)�ʞ��<�\�K5Γ餭s�$%���&	�piN6��[�SZ=�<�#��(k����{j�9�q���0�������nDh���5}#��g ��]�{�6��v����J�1+��Z�n���uP���3�z����]J�<�X��\ʌ�{��6p����헿�Ӝ�=E���(�G�qg�2��`�8��IP�6����Z��?�o_"^sq��
�x'VC�<�¹�~K-�*L��������~�y�/{/��VX ���K�pвt��h1U\�2q%i�mfp�,X�$�}d��O�UI����Wb�0
`%\ǌ����2���^��;]��a���������p�c^e3f7v-
�E�h!��<Qh;���|��%>Z��_�P�!�TT�F�}�ĳf�z�1Zٌ��+�=���*�������_dufogMK_��x�$���i�gqa⤦�G��8Av� Īyw�>�<�����e�� ��R�#��)kl�����&׍z�RN�_t�x^f��gm�����C���U},��˰�'t������g�kl�8e�{y��X}�A�N]��t�8+ɰ�H�����Ʃ*/�?�A���M�(Z������HvId�R���6/�3���g�(_���&+4�?G~m�U,��-��~�6嫷(���MM��RAI@�Nh�c�Z�F&�(L�Ǜ�L�z�a��oP��r�N���!�	��53s�!�0��5;�_�Ԉ�q!�tk`I�O��8#j����Η���~n��"MM�62��[)x��˨�ߥ�{9����c���_���G6�opJH��Pg)�&s�1�4��ZG���+�ʫc���N]9Q�GՖ�T�����3"|�y�f�'�qW�ˑ�E]�k%"sE�/3�.�4�7 ��	���Y�O��i�?Vc���CD�m�e�|�7��<�qԉ��(ȩ`�����|�D6���p֚�O�[>��0����d=�!V�~U㈁�b��벎����ҞiwV������r��]���a]�5p���=v����rU�^����s0J����Ab�,8 Rd�3�A����%�-�ۗ:���^���
 �CeR�19���Wd5 H�p���f��7@�n�r�EU��U$�0z�+y�r:M�����Q��
>�+��Y�fg\Hyru�TKH dʷ�]S���TY�w����@E�6�7c�`U��RS-����� Fd,�{-���n\��`�rnm�c�Qc���.͛L{-oC�W�����Wʎ�;>��
������N̚3�kZ{K��5(�HBGL�'Y)똺���HO�G�*U���������u�Ȭ�nl�τK��73�&7��w�2�g���o�/�hn@u�SQz���/�-����i��u���U@�e?_�$����2��z����^-Z�ƕ�	n�"|U(�a;�\�Z�.g��f,*.o����d�"UƇ�U�4p0z��6|��Ν䇩o��t�ʽ�lI= kK\I߻
�@|*o!��L���&3��?��7�Iݽ����v��`e�#�7J$v���SP��ѷ��dؕh��0�t���#�6��ku�4�B��n�>1eQ0r��U�-��! P�_z�k3#M�� ��t���:*�pm���A�Xc���:�������;�aS����]V�JvMܨ��) XNh�0��3hKr����3�����v��U�:>�]S�%vǱ���KM�&�]�Y�8�b�,�>��d#�`�Pb�o`����9��ы1�<f��݃c�ei9eT�<�ãܘQ����Z'*��؉��h�<[��/�e��\*w��7�H�6%4%?ߡ����".�W�Oskf��1�L�4m�%�?tR|D����C��A�ъu��A/L��B�7ʙޑ7��3�5������Qx��^~��륑�jɚ��1W�R�B���ŋ"z��߂�,�T ���E7����xt�YE_�Z�*ͩ�A��~ ���%�:����d��qZv<�;$(��ģ��ay͟��B�I��,(�!�Z�Υ��Xl���p���[չ�է0��Ŏ��֍�8���B�δ҈�Y, gF,%�(bo���mV%� ��S�˞ҥ�[���\�`.ҟ��t� �9�?�Ch��b	
Y�[d����z�����lfɟ5oov8[h`e�pn���b Y��©ˣī65r�7��f#�dV�˘�m������鼚'%���%�sF�uPj=6�����a�����d�[���J����F�2� GdvMM���S5��F.3~l��j�:��t���-vc9[3 ^��L觱�g�!�5q>���%=�H�>	fA�ԎBU�����lSЏf����qb�mj���-*Mt��Z��,pb�no���n��cwk�����q*u�ڏ&<+����G��Om��"t�w�og|��M�M��m��QI˥V�g�13�)e�#f�h����ިbO?�DQ� 򖵒.#�Ǣ��+���,f��D1��㶷�tŁ8َ���ƪ+W/�?�
}�0)<'�J">Fm�
8/M�]Pqʠya) ��`�sU�R����7��5V��V���lBr`��pL���Ĥ�CC��5BJ��y�丝�11{zp��?���z`e�숈�����~7�]��Ft�٧����(��^1�Z#
�n�wph�L�~F�܅+�9X�;w��� 6�A�R���(����,m�/�)m_�<�/��>���>V2*'������!��E��m��2k[�?-��>;�1G��<ȉ/��ۗ�_^�@�"%��G?T�c�uK4�G�4eL?,���O�}��!t��� �TP��]z@�x���OI��uI���!��f
�W��rw�@���5��:����&?����@�����{B��		%�L��M8�U�R~���b� �JI-��j�#����)b״5C���Շ����&e��Ц��I��\T0�Q�b��Ǧ��t��U���햂݇�ݯ�yô5
+HwR@�4����J�cZ��S�a�!N*x-�Q�[�Dw�{��f~�ܜC[�^}ڃ�c:�Vdi�;�L���?�(�X�G�>qp�Dop5`c�Z���ֵ�N]t��|=�Q�~�Dp���^4����a���:E!�vIR=e��9�l�
T�������/_�}ܠ<�{"�$�oEE4�����ׇi{�H�N���^�Q�Β$/	���K5	�(��~v>2[��,�v��f�k������*�o�\�ם���b�Ɋo�)�n�8ewR|���c:*K����<��;�?M&�vƥ)�wwC�|i;��"c�U=Q�:��퍄Xw)l�RM�h�U��O�m?.J&Q��Et#�+â�}�+�ZD,-����j���5c�M8 ����~�+>����}8��<�zW��F�)�8V�t] ʇ)�)�.��2	s��7�B]����\��]�:�S�k`�p��J����Cb����--�G��`�o��]1�.�pD޾��pz�˒쯷��
~��]T?�FPs�f��T4�����*�/
♝�^�&��F��+�/�XLG�w=z�'ӐA����߫QՄ��E6���tmƑ�Z|8a�&�̾
��c� K�pe��gp:Vu��;#�*h�
M�<d����Q���(9�"��xF�^d�}pξbA������L܁BC����j
�1�넾l};0B�*)OҦN�UW,���	�
���o��*��A� q�dS�X���wWJ�\���A"h��>�1�@ �=�d�R	�r�����f�ɾ|���}�1���v}�����*s���댾��U����J���{H}.���s^��I]%�)7���U�G&�B���=⾪�Ka	�� r�,�SE$�$'�(��mJ�6��H¢@Chr���U=�l�#c�V���>�g�5���bce�Pm�șRܳZ��7̬�[qI~�^�m�=��"&��X�ox�y*�ޯ�!k�"�Z�s�9*tD�y&���t��8Q{W�bQ���S!W��sT  ��� �s��^M����8�~d�U��f,Fq���ڗe��uu�MF��a�ѩ[�a'��n�!�T�o�?nL!� �5�4"�YUKՠ'���,��y��E�m�t`���B:�4����=���T[G�S�����W��oJ�FR����ņR7Y��\�V���3�O!�sD���.�p�h���	��NۥsU`dE�-LK�7�#�p�x�i�����~�Uz�����v`B�{E#R����zm�,�x����>�C�p�B�蟧�V�T'\�w�G�����=���m������i~ �}�i�_�*m���+=^A�?.FZ�rw���2W�f�iԳD�d��;V����C6�RD�w��"�ۄ�}|c�'c��P���OW�Cg���R"L���T`�����^L�UP�6u��H�_A��Ϫn��&Z.%�75�����(���m�x.����o��g�,�-[*�[�F�%�y��Q'U��n�Iog��)I�ʇD���ũv5`��
-u 4D^Jڠ�x��ѩ��8y�%|f"@ի����Wp�^f��C5�Ip9IC��D"��AY��i����0��^�2�����	�K�ƞ���L�ݪ;�Jb��������-l��YJr��W_�Vh�_�	?�\�(�gwW�S$�ϕ�L��l �N�)0_;�`d�fq�Rbd��f9(��K�lj$�� �x���o?��'��~9��~ٝ�e�l@u9t�>Xj���U��f(=��	X �d/�^$:�ۘ�Fe�0�$��`%�.a. �qE���}���z/#[�l��v��1��,�L�8��#H���z}n-�/�ӌ�'+��'�������yǔ���07���X�#4��Îb��o�1�yokhf��;Em�1.Q_A�Y�u���U�;Zs�<��K{b��|��R.=9���@��_򕿈yz�)�&�{Ko� ����ٓs�y�[U�x�����o��_�ey���������8U	{7�'v�<&�{E/˰	36�X(Gx�!��h"��X�<O�f]bB/^�4'��i�|����	3��v{$<ia�����k��K�m��� �q�#	ʷ�N}�3��Z������ZvE�и{�/�S�Ǭ�����⑁�G�̹qhlP�5U���a�7��u
�5�a�̾𪐂N/l��gJ\�;+Ȭ���}���-�M���e3w�R�3��J�~�0'9\�3$�S| �-��+ԗ����� 霃(��
q�e:2�~��ЪI(/�6�:i�`���_�9�q_�v�PYMCé��	K�L��������Vu���/ׄ�X�E���aFK�>Њ*��@��\���%A��fH�<XnA�}<�|�'z�I���/+��7%4&a�I~�����n8�h�vǱ�_-Y6���'!c6��>-��9�@|�da�Q@����	��L��I3(�Ǳ,־��_}X��f�K_��Q�d2�ܞ�@*~�Ƴ~�r�7��fG�yK7��x|��q'{��;�a���#t8�����Ă�������y�=������Rq�H���s�"������SR&d�_L�^>ͳgE���`���m,}��ˈiZt��}�n9>gZ�0l�E�S��0!�A�m��{Rt�m���s ����VΞ�/[;�A�X�%6T2!���;h�tN��*(ٳ�������{�(7g������[mg�,����[�^6��;(}��M%�p�*P�mȂ&Q�c��>��D� ���s���R�����'P�Y0�&g��@��3Ks^���j�k����`{�!�`!����g�j���ܦ����En���M%L�6
�S�/W��W�?,�J׍Xɤ�2y&S�R����j���w�+�v�s�}� �2)��R<�D�]�a��ǹ���O*���}\�щ�*8BY�c_u5T�1[1f�������l%G���Y��\�4+L��7Y�3h�4Q���Q�˰��%�K�/@����3�q��#��e��D|�$@��N$<v@�7ie����Zj`1�㚼�*{2ȑ�E���U��U<h�w���0ohn�]�T�=���欦�K�\c�f�(iQ�C���
�9��
x����4�ق����}I�ڑq���ie 9Nh���TM4�o����b�����Q�5�g��Nt�3�n`��U	�@Z�I8���Z] �e��0B���\�u�Ķ�O�p��~h:�>�x�p���R�%u�j
:� PG}bF���OP~C�<����[g����&���p\v
e}$�O��Tz�'� ����V,)2P��Y�?\��a�������;�Z���-�)�-n���nz`ץ��6�{��pכ���P�@��c��������ǱUlѰ]�@�:e1yif�_5{c9�=�+X� j��K����e)�$���>���x�a�i8{��j���k�;|A=׹���J�֕��|��u�	P�H�&푟,hRtv�CeiV܋�5�ۓ�{�uN��>�r�y�c��2�� ktm�l�x'�B��{0��O�Egx?#&��kMa{���߽�|u�zE`z��K#]x�-����
�rGi���&����Es!�
߬o�'%�-��)G��v��7To��6���y[�,���Mmj�0/J$7r�qw�\�ˢn�|"���E,�%+��@��-�V�K����K�-(���>��˩�JI#	ӭ��Je�����k��C�;}�O���W�����n]
XLhN%3����r������t��d}���r��o�T�:*�TQ����Pr	�g��#~i���eH'(:b�X���aL�b�t�D,���	���=��J�j�a��"�g�6�I9~&�i:|�)�OV�za9���h#�3ٶ��ef�;WY�<!�_�a|�Ӣeo Y@"��H�A���
; +��
�ύ��L��j���V@�4Hd m���Y�B9�	��o��4�c�=ڣV��zQ��=U�5#�p��%��8u�ʹq�IS���m�vl�RrI��pA�v9���ɇ�w�c�{������ �m�'V������� ��5�x9��<�pj�g��Vu�/;#�h��X�����Q$�j�(9�����^��}p�|�b]�Ӏ��L��BC( ��
�����};��B�FO�B�N�q�W�X��%z
�W�o��-���� �.dSSօ��W��\��A�S��ZA1��B�=ЦdO�	Ŏ.�����f�|�����1�O v}��A��F\�J�-��a�������×�}�?��>s�F��e]%G�7 H�U-&�4��J�=�_���%	��Xr��DSE@���٪(
��	�6�H^C@C��ră��UY<�l��#c̸���>���5���~se��Pm�O�RxZ���̬G�qI�~^�	=��&�SH�o![�y��ޯ�;ko��Z$s��^tD�A&쐫t8Q��W�~ǀ䀍!W�EsT�0��@� G���M����#
�z�U��f�2q��ڗ�u��MF7�}��E[Ԇ'��7�!�0�o]p?nht쑜ǋ514"�'UK�!'ϑ�,�(�y�e��m�#`My�BV�4��A�=�l�T�ǥS�<����W��o��FR���aR7u�\B����#�O��sD�\�.s��h��軀k���ۥ�`daH-L��7�p��iʗ�����Fz�j����B��#n���zm��x����ZR��sp�B��'��rT'���w����&
��YW��	n��'��� ޙ�i���*m�ɜ+�/A�[#.F�Tr�i��'rW���i�Oۮd�=;V�����EC60�D���"��ۄ�|�k'c�aPVp�Os�CgT�R>��/�T`�����^L�wP�H�u��Hn�A���n�w�&vu�O�7Q>���D��	�x.�����,]4[*�5���%����Q�I���zIo���EH��#'�����vQ�����u P(^Jv�x�ѩ�>�T�%<"@�4�?��W��^f�6C5� p9�ݏ�`����Y�O��*]0����2W���Kw�ƞ�L���ݪWJbsv����\��Iۅ��oJrgW�Vh2C_���\�|;?wW�$�k��L��l d��E)_;^}d��!�R����9(e�glj���*U�x�����K�2�'��9�~g~ٹOe�l\&9�>t��sL�U3��f����%n � 	�z1:2���
e��+$;�`�X.aJy ��E����R�+z�F[��(�e����M��L���S�H�z}
-�/�ƌ��c+�R��Ji���ǔz'�0*���X�?���_�b����1��yo��f��\Em�e.Q���Y� ���d�;v�sdb��${bB�|���.=�k���@=�_���y�)�B�{K� �����/�y��U�u�� �XM�����y����\����U	�7'�'v4�&��2/�[�	O��X�OGx�<�����t7<O7�]~�/^�&4'!��il����	3�S�v��<i�P�i�k P�Kʖ�q��q�	�SN*��3�2Z����u&�Z����T�{�K>���Ǭ���������Urhll�5U )�a�½���5�#�h���I�N�H�	�J\`�+�ȣ��XH���K�MQ��eO��Rb��	�J��ͯ0C|\����S�������GE�����I�0(��q��2њe�lDI(K�6����|��6�_�U�q_�նPuC�E4�2KKcL���ӑ��V)��z/נ|X�����}�K��fЊF5�@>�\�ڡ%AX�fH�&Xn�)}<�]�'�I��y�/ǅ�
G%4�S�e���C���u���v㥲_ɍYR?����c6^>��-���@_d}:Q@PP��,���諚�e1(���,�^�}X�yf����8t�d�&�����*~��~a�7��fG,�K7#x|K�qC1���/a�03���8 U�)�Ă1���2����=X4����Rq�u���sk���6���nR&�7_L��^>�gE7��|���6� ,}��ˈ�$t�\��nU�gZzl�"��S�'�0=�A�	�֗xt�	���� Wj�+Ξ&c/[W�Aڹ�%R�2�f��7�hYN�D�*������ٝ�{-�(7���Ɔ���9�mg��,����[A�6��u(}xZM%塺*��艰�&�c���A�� �g�s(&�Ra��XP�ut�&�.��"����%3K�P��8�j�T��}�`��!ש�`!�ǩ��j��=ܦx#���n�a�M%h�6
�ӗ3QN���C�#�{�����҃����ԇ6~�~H�VH�u�g����(1��0�2nx��~բ��c�i]$z�ǐ,�ҵ� '"T?́>���I� �i�F]��L"K��/[�.א�7����m�1��Or$)���}�Dlue�07��<�{ ���ȁ@�v�Қ�CD}���{��r�3�ܞ��F�{�(mV��`ʮb����m���{ǞAl�xQ(�����W��5zę�\��Opd�m=N���{Z~�6��3"�K)�ί�����=R��3j����%-�<ʗ�ז�J�yyc ��R�.g�ZaEd�� �#�[3wͳ�e�F�P�of�-y�0Rs�y��:%����Q��B>�*g�W�1t�g4WZyڴо,��K y�ʏq�S��dT1_u�������(7;ظ`��l�Sc�ز ǥi]qd�-��Dn4��`��T�J����EQ;[��ⓛڛ-G�W�/�A��`>�/F�k2_���M���4�y��r��k2yP��55 �� ��$�Y}p����� J����-Ƅ�����)���.4n�(��\����}&�&�Om�2��d�m�ؼ��n�WS)*A���,� 5��F�ip����G�@q�]������!��8���@����6HZpu�N����n���g��`y���X�ҡ%��b�"h�a�y�z�f��#E�f.�`����o�����k,sD�s�8�e{���|Ě�.mjX^@4��_"y8���)���{{�� �m�	�錩j�U�A����O5��C<���y"s�(���'ngU9��gN�'�A&�J\/1˻�9�=��G��l�6ʓ̆<t6]Ia/��4W�}�����/�#	csʦ�<�j���sΛ���{���,�/��97	��IN>�~�c/!ZE��+1�a]� 
5{�ΨA�i�܌�N����O��.kh�k�5�����ӽ�e���>e' j�~�_�8�J�u�+��d�z ��(�}~�"����Q�h�J��e�`.\� ���#�>&[��Jȗ� ������̔�(�[q��2Bʤ@�=IX~�6�ok�;O�G�_*��q�=�L�C����56K5�L��=�g(ㆤ-�[�/�)X(�4��K��кer�pC�\ꅣ%qi�fx�?X��i}l���W?�I����_��8�%da���y�Đy��}!�C]'��b��.��]�5cf��n�-(�p�'�,Qp�_��g��-����,�X=��\E��N�}���fӬ��"��ٔ��3���*�N��J|�g�fw!�Kg�x�����j7���a��_�O؇8I?{�N�Ĳ�H�F�>��>�m��(�<R�˖�1���~��1_�!�pRV�_|^n�%gu���:��!��,�˸<_t�����g�#�l��߹�S��`��A���t����>P0����/��cA
��Uiyb�l�
�y�b�~ �Z�-��a��	����t�(g0��.��!WS�G��m��O,뎾���f6�@A(�ՔMU�'�Z�ĂVbc	
��N�>�0iǣ��Ƃ>��5MP�4��VF��)no��Y#3{f�\g��<[�G�Ԑ��!f`Q4����j��-��e��}�n�Z�MU��6:�חc�ҩ��]��Z{Aާ��z�����6�.xa�H׶�g&f
�.Q-1��߃b�����M_��ܾ]A�p�O���\[*��#n"����n���y�S˙�]�7y"{��/;q.�7(�ڸM4�af�O���G������D�� e�%7�<�����mȱۃ&x���ٌD>�S�	/�֢6)�c�Ş�W���^E>\V�c��/b΅뺶���Ԟq����LN�����e熙1l��p�H�=~�~�����fa+"��{����يy��4q#R�g3��g��掊5#d�B��������R" �uR�A���[d=��P 
��0 ��.�v�-�M���]�>0�.�y%":U"o��~Q��S>�c��Ta��gdBy
U�\$�KP�xʿt	S�2Ta���1��H�d�R�7k�`���Q$S5�������d4*
-��%nd��`�&�z���&�zQkJ��`�
�-wo��_�t��M��_ّ�+�P   7
  Z  �  r   �(  �1  58  v>  �D  K  �R  ,Y  m_  �e  �k  <r  x  �~  ^�   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl�&X��;O�{�'�jn�!3� ���ٻ�
��3Y�"`�j:.5Z͐�%F!5�̢�(w��p0��?U`���?MR�*\�!��y��F�]O�y��Z�LA6�ݻX��$����*�@� ,��냊�(���*��ea��)CN�!2EcR�b�L�ps��,���A�'���Ё#[�H�2��n�V����O��d�O���O�"��G��"H�J��UP���b��O�����%`D��By"�'�Hp
��O2�'~<��%kJ^�#�A[�>�q�P�'�2�'��'8�;b�'����O��I�{�
U(#�S /� Ҧ�� f`C�I�|��TO��}�N���(�F��O�I<Utȡ��?Ū��"�|�+�C��NȐ2	�O*�d�O���O���O8�D�|�w4cpd�5�Da[�͔�Z���;�v\��h|�V	oZ��dզ���4˛F+eӮ�ğ�����{E�%
�����UEz�ʅN�>Q�ӂ堰�7�J.�N�
�/�3�*�s@\�}r�<�	D�B�oZ7�Mñ�iA���O9�U�N r�
���,��"7D!���X#&d�3�`ӴA�"%���k[iv6���E��E�,@B��ߦ��ٴ-���.K�p��@i��T�n����p��4@���@��v�l�o�M��ׅ9VR���Ɵ%?0�X d�ե!�)���|V,�a`ɟ�<���9q��"k������2��.s��n��>O�$��$;�6�@!Dͨ
��T��&#V�010��$uǂ1[p�	��M�S�HRĸ:��0J_L=a7�N��?�2f��qt��C�I8$�<8 �*��.�B��O(�D[7*"ilk��<ႃ	D�:��!��d��?)O��$�O���z�8� -C�~���x+�ҟ�J��ޗ��)���P�g�t	[��.O�)�Ȕd��=[�m�	8�7��5R����m��j]T�1��@������M�2���O|�6�r�g,ͦ::=J1�9���	П<��f�S�Oޞ��vM
 a6B����U4}-�p���!�,
x��-�We vxxؖ�Ϛ�?	�����\�ݳ"!l0j�E�>��Pq�
AtTB�	;LNtL���ܹl:L�`F�1B<B�8Ic8�ɕH�F
,[ 6�B�ɮT@�x�ݝSN,��-xR
B�2+񐡀"ݾd�M��B��$)�&�J�A�j��<�R�&{����{��"~� Ò�j��p�3H�;K=���&�yƈ)�a3���@��`Spc��y�� =��k&��C��A)a�P>�y�il���ڨ6��<�U�@�yB��S���ӎ�4��|�T�ŧ�y'd9tL�e,"�8�R׎�2��d�+bO�|��٫|��[fiV��Y:m���`�'ަ�#�d�1L�5�	+Zi��'�$9�����_����D�=B1��'r�ɲ���}�h�S�ٮl	j��'	�hBF�|۞�qTkƚlCX�ϓzXu@�i���'���K7!�+c�PXň��R��]:�'�$޸U���'��)�62(Eb$�e���s��O�����?�p�`PF�<��<s��'�E�ׅ�
J�Y�d�X<�&l_�
�29�4� U>H� �ߧZ���a��dӓM���c��o���s�c�j�^͓!8O���s��ty��'��OQ>ŉ	K'��h��g�Q��f9�IB���㟔XKK>es�d��aV&�\ ���O��O�\�g�6JO1��v�IGa[�f�����Ѭ(Į��2D��c$�ۙ� �)%Hѿ~�^��*D��K�� �B�@��ٷT�E��+=D�ӓ�I��r}����."VI �:D� P�쇰;0��qQ*\T0Q3�:D�xzbb�	�>��֋"\�#T����$�r�f��?����@��ey��C�ve�G#Y���	�g�X�6��Y�*Y�J[\7�ު3������|����$���0CN
;�XR!�%@,��]���$!���&�T"1�zVг�'���y����+�����v
4��i<�>����IC�矬��˟�� ��.袸��*Dt���}x��Ɋ��W?DOb�&8jq9s"�(��dBܦy��4���|��'����B 2���9P\rԳq�F=K������xxn���O2���OJ�;�?!����4�݀ ���R5�ȗqZ��+���8-�ba
�'�(s�DU�.Ȱ-�w�V������x��U0,< ���~o1��]�2�������2?n)m�X,Ew&�{�ŉ��yb��O�����
?IlabB!���@��֔|��\��n7�(?��$�2T0$q��lw��5�Č��l�'y��'��l�y:��#���_���;O� d=r���s��yK8߼4���'}����SxRT�%�ĄU��q���=(%. ��&ŏTӆd`q���)�*T�ŎN�'R�����қ��'Q2�FJ]RRd���p`�Ca��'B��'$2��4��=y�8M+G*AqLhT5�_'TV��
�O5�wm�W���T$��I����'E剈\�j��޴�?����)Cg���Dۺ��0#�������6+���d�O��GE�nV�a�h #<Ɇ�I�(����d�?M:����m�V��S,A�x%�R-?QA�
��qRt��z�ܐ!AK�4����`�Mѕ��b�+@�jf�� H'*�Oȍn�/�H���)��N�.�P���& &�9U�6GfC䉃wQ��:T�ƛ�\�bu�A�D�"�?��S�����e8O��(:�Ȋ���4lZ����'�%Q��a�����OB��<��=2c��c� ��茁��+�?���O`�*���B����$�-@ODx!��þn�H���
�?#�\z�B��/�HJE�Ã`�
̀�����	;:�.���"�8�.\�aCR4H�8���O����6���*�<���E,8��l��i�Ǳ\�k+OD���	k̓Hގ�#�M&"\�� ��@��'���C�~I���?qDd��8�O|�a+��ÞGJ����ʜ:��ݺ0�4oZ�G@��'�"T�4%?I!˕�\��MJ �B�PC����J� ��8�,Vx��L,��.J2���#ХB���F|�^4SQb��zV�ݢG.�+@`��I2%`x��\:�8�+w��0��H5��O��d"���O��?�	:uONy����P�0���I�Q�e��;'`DI1	R�-O�c�B���zX%����O�ʓS�i�!���_"w���Ɗ�� m� �*�?�*Ov���O���	W�fC��J7P�p�1�-�)�M����6C�$�X�XK� �q7�A�T��ȁ���{�m��n��H)U`�'^Pm��O��M)B�8EL9ǔ}�r�	':�V���O�X.��L�/Vs0�0��G�JNU'���	X���; �ǲ?%���c�a^J��8�Or@�I�m.�@	g�.4�L�;�e�&:�&��<��N����):-�<�0h��C"�U�.�D��B%N.����O|	�Q�Y�t<��qf@)_�
`��t�O��z�� z{�×"h��m{�O�x�̊4U�BM�����i&x%B߸O:FP�Α5��tP!_*I�L�Od��4�'�b����<�URwH�j�.��De���ce�w�<� ��XQ*X�E��%�r�'�~�}⒨��iش�31J�q'zɳ�ă���<�&�������?����ّ	^�1��oC�IS%͚/M҄�aA%%����b�~E��� �3�	""� 0���
���4�[<;3*�#�Me��4mZ��|��a�~̧���'���F��a�fm KѮ1���x����V�]C��'�ў���H�I���R��59!�K�<AE�M� � � ��B4}A�,Py"�+�S��U�����5TzR�+P�G:M�CA:��U�I��,��쟤���O9Hxs��I.OD�)Ũ.T<���Z7.@\��Mt��eC%�4<O��R&�I� ���h'	A�j �as��Қw�F�	�N�P��0���r�DU�`�		4!��H��E�Z�v���&L&0U`Isfe�O<��!ړ�O�i�A��m�����|�TMpf"On,r5e�nwBU1*\�0�
��P�|�ţ>a�2F��� �-:d�b��:Y:x59��M�y¬̍�-*d�]�HE�B3�_��y���Nr	�"OE�ĳ [)�yb�_����"� ,	ݓ��T'�y�*��:����o�z="}�e����y�&��Q?���4� G���R0�hO�A��S�?<�GcUW긜��.�)
��C�I�*�� ���J&[��x `�zh�C�	�r���X�X������
��C�Ɏu�DY�#������+�"&�C�%�
EG��_���d��*�hC�I'TE�[���r
X-?Q.����"~R%ߥl��l��&<:,Xō���y��+`�P�z��W�l��ĀF��yr� �6>6܂`(����	��yBⁱx�x��(G'����〴�yR�͇G��	9t�>{�� ���'�y�hE�F�fL[ ���n�FaVD%���'}-�|���%�
����h�0�YF)��y
� "���^$/�(�1V�2��P"O�T�UB�F��p@��A	��P"O�(0�`�9 f�)�� ��!{�"O<� �%[�g�-��n�1c����'i	s�'��Y"&�.P�Yr&`Ӡ>�H�#�',Z
	>��b�v�b���MJ,�yB��<a�('W���hB"���y��U~=�d�2��X*���y���|h��ېe�9�$Q����y����r��Ŋ��{�"(�@dC�hO�P���&y�NX�,E?7~,��m+[�|C� N��Y�a-J 	��#�:=z
B�/[� ف1^�7��}���K�N��B�Ibw�%w��2Yݔ5c�f��[R�B�?_9���T"Q>�T�BtI
�}{PC��8l#V�k�m	-<���3UE�<=�>��
)'�"~Z��Ŗ'��$�� <X�Vha��6�yb��%t�p	�3g�FTaD��yB�X�����K `�����y�m+&���W���ܴ�0�S#�y���5rt�ɢ�ᇱ7���Y�yr��SV�݊i}��Eҵ�L�����:��|��k�~����n���L3�y�%��8�TI!m�6c}p����ɔ�y ��>4\�k��52K���)��y��)w��H�`��%�Z����y"#ۗIl������&��,�1n�,��>AƁBS?��L��v���r��{���a� b�<q�O�7!��� g�-vu��	c�ZF�<���Y�g�� ����`��I��A�<)di�<$H��q"L0̴����B�<����&FV��0��d��WlI�<�"�L'�6䅕F���҈�A�'��]3������В��]s$\c�
�#2�!�d�r�FBeH�8�z�R���7P�!򄎓I4Tp#h�3~&���ņ�nj!�d����H�h�%e�()=E!�d��[�^��%$[�:e�9`�-C�<6!���9
���jJ\a\��l*��N��O?AH�g��c�f����Lh�G��m�<a�9|n8�|'��"oAi�<A��K�4tx͙�9w�D�f��M�<� e�{�j��'K7k��PC�G�<��j߅W#b���o���$&HA�<��困S��" B�-)^9��gyB�W?�p>IdV�U�r8�B�C4��Zr��f�<Y�G�3���lI�VxI����Y�<)Ŀ_�cF�ՃK�ͺ��L�<9�JF�I����l?�i��
D�<��&Ƥ��@j  &ڶ�c�&[x�h�Eɹ��R�#�i��yUe�eW���d�,D� ȑi�1&�#�i��~��{U%D�<�C �*	���#��.T ���ċ/D�@;�p> -���Z @���&�-D���W�ժ&*1E��W (8�%*D��H�m��DU�AA��l�.9Zan"�vЬ�D�T�1<H���.�$i�
�,L��yb#fQx����r������yo���D�C6j�X��zCc���y2C:i�.4�5�JMzr��SY��y
�+� ܪ��1���c�@��'�`���۞\��b fY4-��@+�C�NFx��)O�,���B�*b�
�-�7^w2C�Ƀ$eV�aš� /�
�p��M+Eh,C�)� �����j�C��P�@c&IP�"O�A�`H#���v�pX.�s"O���O]:8�.�%��v�0"O�tIVEĺ	��D�T*T��l)£W�$9�,�O�<b �Ο�]��/X�ʼ�S"Op��O�g0$���+{�P���"O����I�LY��H�N^4=�B�
�"O^�����@&1h��P�C��mBw"O��g��[��K��pt�!�1�'���'���0\e}����V�~6�d#'�4D������	M�%���Ԉ)��1�(D�t�r���@��kT�/�8b�'D���tL��"0#&��5d߮�S��&D� :�朩 �����ԣ&Ԏ��0�0D�h�$;;k��!�R�\�l���!-�K%��E�tiۃtE�$�D0E��u�!/��y��ߏf(�E���p�.M��X�y2-J�<�&�B��J�j�(�q�O��y�愰aל��Ei�%fQ�Yk�I��y¢�x�l��Q�5��L�4���y�n@-]yzq����4�^93h
(�?)bH�X����t]��`^�B�2d��	��D�8���<D����(S��c"=d���:Ac?D��Q�G"3�,L���	� �;�h!D�h���6���Cb��4oi�];b�+D��[w��-#���)G�{t��@�(D�k��z
<���C�2�|�1�g�<��d8���6�R>
�x�����_�nijci?D���bN�a�Ҥ����#4�:RM0D�Lr�%żxH��K�.�JD F�.D�H�E�I�fi�`�ը�0�i��+D���):sizhJ�=\j��*5�+�Oj4���O�m��bXvS>���:B_@H"""O���F�D�g�d����>omĵU"O�4[SB	P�I�Ըk�4�t"O&���oӴ�48��
���i��"O��C&z�|���D����׋�y��Q, \�9j�8ِ5*����hO�U����	T`A�B�>>R�`���i� B�ɑh��qHb�"��ɪg��0<�B�	2��T������x�� I3ZB䉥S�x����<�~��!���C�+!u#�I� �l�8p�[+j^�C�I�E{�Ź�B �ZEs1&��veX���#t��"~&�G�A��(�&ϨT��dQ�ψ%�y�֒!��a �'H��`������y��̆!�کz$I�0DV��B� �y��ֺo��|P�C�r��bJ�yB�
5]	`��Dk?�t)GOY�y�+�Y� �Y��ZY��� �F������|bE��9<
0��������I���yE&.�
-r�ڈi�)�"���y"�K�i�ǣS�^|�4a�̃/�y�Q�RSLPa7�� [8=���A2�y"!Mw�|mӆĽO�ƴj0K����>�ǤOp?y�@��(x �G�ON@%�!)�g�<15��6Vr�:�햂X}8���IPx�<���@!(f��Ek8>����1�Z�<9�`Н^���3aJA�$�`��AMT�<��J��-rB鞴[l0��ff�P�<���H5|�Nɀ U�:@Ш��v�''�ۍ�I:X�v�
É�;�� �0ꑧ�!�$����I�z���j��B7w��1�'�q��92��X�A��n(E���� 
	kC�\.*\^}�����o���br"O�Z�����\!��i���"O| �c��/���I�<XpZ}�B�'Ũ� ���/�5q!�1+x��)�->��L�ȓ=�`�%g2	Rp� �c�e�$�ȓ W.���6_E��#g+�*F�؆ȓH/.�' �T�X�R"�
U����~U=b���\b��J=z�d��ȓ$T�I��$�������7]�F1�'m�I!�V,2mX�K����`w�Դ]��ȓ��ĀV��(���[c��5砐��^�i��.m."|K�fC�>��d��D��u�T(���A��V`%�ȓ4*�@SB��2�����gT��	���I)n��q@�U�&Y�TV��l��C䉹 h��q��M�4�H�*�[��B�	�D��`rW�,�X��!�$ UB�ɲA����fA�1����Ro͆Y��C�ɤGX����|t�h��&JQ�C�	��f�3�A��u�����Ԣ=�t�U�O�d�@@��
�:@��(ɮ"��j
�'ȼJ�K�3q�^i���{>Ա�	�'Ҩm���;R��[��#;����'�BY��"--H�Y�ڳM��	
�'yJ�����9�ޅ1׆�8B` %r�'�����d���g�̬Y��~@mGx��I �V�jm*WiZ�c��p�Μ(*�B��5V;���B���*EcP�-�C��9A��#�J�HI0Pq�LT�|B�� QgPD�0��
��Ha���5r2C�ɐ�P��یy��i�a�P�C��"(!�h�P�ǥy�t����
	����Y��yy���:1(c�,)c��#&��ј���!e�N��%���d�O����Oj����^q+��U�%�d��i>i�2OߨX0=�&OW�?�~���$2�e?Mb��4�t}C2�^��MC���"}��t"I	�xYdEs� �W��������Nc2�'�1�H���F�3:�&��S@� ~�@`W������DQ[�/��B�"��qL��A����NRyBgץxP-Q�ꈓQ�m��cS��D܋_|D�o��ؖ'�����I�W� ���Y�\!�r��U<g���	�' pѳ�2D��Qz%o�;�?E�D*G�X�����'5O��`�Iޮ�y��W�
2R�*�B��D�<I�0�i�����鏴5?A
&��}mdP"����@�$Ф`���'��)��9?yD�aM���`�(PU���j��-C!�޺5�ZX���Ӵ2❋����ў�y�����#����P�B�y���t�����<1 ����?!��?!����ԟx��n�L.D�zF�P=��%�򮋛}�x�Dβ]��m��R���3���}�o�;f
�@��(�2����S,�M��)|w��+�$� ���S��'g��"�]1AU�xKV�
W
���O�D��'���	�<1���qx��Z�Γ6c�Y5��g�<�qEʉpLB1+��D3C�
�P��O�`��4�����<�bɄ���9y�FNi��*�`I���2���?����?�)O1�@(*$��9Qn@���.A��UH�&W,g��A� ͸ ds���\x� �C& �8 ��q
�>*�V��U�qst���@�g��i��¦�"`I!�P�ɳf�� c�R:cJA��ƐC4`���E�'��J�h�0*B��$j|F�ۦI?D�{Yyl�ѡă�'I*����^���d��M�	Ky�k�5j�7�M�P�S�~�����XN���pL�,P\��'M"�'�"�\Ix�1'B�N�����O�)\'}��+�愳g�(MS��\8����J�qwHZ�_#��mZ�p%n��ƃrb��	��8f:�B��RF�'�~p`���?q��Aʖ$x�Ó)�4$�Nt���d/�O�C �`�R���� Ӷ�`#�',H˓%�T�2K�ko�$g�D�D[��'�����,|ӆ�!�a�<�)�X�I�O��h<萍qC��vK�E�O����) �Fij6��g����)��|`��B.i�`�R`[/������@�U	�16� a�T(S2�M3�$�[�O��t���-Lw`�T#���П'�v����?��O�OD�)� ����I�&Av ����D�@T��"O���A�!m
��ŀOuD����ȟ�P����/�(�*�/�5����Ǻawd˓Q�zQX��i��4�'t"[����H0���,A.+�( �fT�/�6|�C"��?)0�̹'	��o�n���	cȐ�	&M�i�
0W��'�X�ye�e�2����UP��-�E:ҡ"4�)r�^��
"p*PҊ��i�N�G�P���� �Ik����T	�)>�������*.fH����yB�8D�xtq��W�JD��g r����HO���O�c�`��_�	\�`Ib��vvԥyk�O�a7�' ����$F������a�����'���	4�ť�h99u�I5i��d��'�t1�BK� P
q4e�a����'�l<��茈1�thk�bD�faFI	�'�HR��4�"���i�\���)����#P��n�����	�|*1ƒ?	{�)W�L?a���G�L�<Y�Șҟ��I�ic�"w���(vE�!a�"����|2�:u�J���N5�J�y�cEs�'�h��� g��iEC��F�X-[�栋�JG,>�:�BG/�8g� #1�I�t���d�O����O��22��X��]�`Y�eA�ĉ�dj���O��"~�/�,ʢI؇KKp���7ƀ��$7�S�ԁ�<�� �-8���A�y�XkЅ�oyR�'��5s��'5�O�r����g:��,:�,�H�`�f&O��=��Zy�p)Pbfە��h��Op��O�U&�T�f�'��Ӡ<��� �, �9�8�c����AZE��4�?�3�'�y�H+�?Y�������y�	��C঩�f���v��� 7i�f�a���i�"�^^��<O$ASҟ�^wИ��s(�����5�� ��.q!�T�'��w���o���Iן ��⟀̓��m�	�fQ����O�b�@ٟ��ɖ^�<��	�<	�%�pnz�r����sc���tu����4/u�B��'3�9���?�R�k?�ޟ(���?��ɘ�.��FZR��e@aj,ƄЩ��Mi����ҟ����ݟ�̓P������]��u�φr{:`�"��	��HW*
�M[�'�T�0���?Q��[���'�R�Oh�q�'���r�q:G�A `E��ߵ	��D�%s���'���]��͓1�<�禍:� �?�1Ԥ\:(�T��de�> �� �4�y"E�ϛ�Cf�| ���?����?�!0�чF�� PV�������Ǖ�M��Ц�y����?!��Z���y��Z��ԨC V:���h�8���򵨖�Iy�6N�\�W� �	�b>�I�Y�Ŧ	'Da9�oָ����ȓ:��0�� [��h*D*#$�l�'q��IyB�'�U�P��&�\�`�nU�-�j�p,�I.%!�4�?Q����D	Q����i�ΐ(!>�>aCj�Lf�i����3�S��&�P֌���@�|st�+�/��y��
2R�Е�ټw �ջ�MǱ�y���7���{��V~�af�;�yr퀿X���J-|�h8��Љ�y��ˈ0ٱF�Ǥv�����H�)�y"��+ �̵ѩ�^���fؘ�y2A��4U��gM���xFL��y��"�yr�_ 
�PxN��y�Вs�jA�f��G�(���j��y2�V(t�A��햀S�z������'=�"=���d"wb��"���w.�A@X�"O@���ӭR�%�Ń�71�Q��D i4!p��J�R-�fLT[����GBKR ��i��8ǆ�BuO�9S���p��@^��+3�[/Z�,ȓ��A��@l���V%�I�'o�&��Mj��H�&�f-�f!��r�x�8����e��y��b
*܋�Րԕ�e�Q�+�v��5��F���OԬ��Կ��)A�S�(k�!�G"O.ab�>=�� h��w�H·"On�($�X�p����fIY\�c�"O��0�hYj�&���ŭ_(�S�"O�,�EBƓ�6�H$��-`�xx�"O�pk�FO�9��1�"�V7+�N,u"O�˄�]~�ؠ�6ff~��E"O����1k��yC�	�%|&��3"O̐R���)w1DM�%�==��R"O�1�NQ�Zp��RFC@���"O�P�C�"��i�4�N/뀍3"O,�K���([��t;T$�V��1
�"OFT�i��]r!FT�z���"O� ΁�� �/Z,���� Jd��"O�Ir�-]1&�����B"O�e��*�a#�K�D�:��8x@"OXt�nX(H.,c3�Њ<����"O��q%h�d5��ygJ�BSFt#q"O��#���aж Q�N�_ti
�"O=�����k�-2MPe "O�� �C�I(��Cg�Jj	J`"OԌ����%>:=�e��&3�A�"O
��U�{���R��нl9`�҆"O4��0ؕge����; .��y3"O<�GM�37�L���,X��;�"O8�Ȕ�����r#�5H���"O" �-N9|���)�a�K�Ndʀ"O^� �i@<�q���@
{� ���"O�̡���+8踴����QЦ��u"O���S"M�q��IS�S�Ga����"O�z�l��bZŐ�c��XO|̙�"O��c2Fjr(E*3	D>'&0��"OЁ�S�9z6�(A��N
 c�"OĤ�uc�7���*Tƙ�^"���v"OL� �`�8��#����Bp�"O2�C�ԕh�	�D	�5.��]�T"O*}�@�*oF�����^޴e��"Od	�W�B_8:uqe�\ G"�0{S"O��֢��n�H1!�"=Q�"O������^��d�ՠNB��Rw"O�ب��65i�Y��M-c�|
4"O<��%L-�l傳�v�h�r%"O�	Pĩ]�?v��R��1(���"O��ӣ 7&y,4�&��?����"O^��"C�&���pc�<h�AP"O��s��7sM.`ׯ߄6/Dy+w"O" ��f߻�8�0Ձ�=t�`X�"O��BE�pP�������o���8V"O(�`��Vg����Ɔ�s��Y�U"O��2}�	r���3��!85"O�P�jHh�hB�6~:��"O:(���(za��H�ɇ	rkdY��"Oƨ3�LO�9�4�`UhG�qp���"O����e��|y;"�^Tuc�"O� [d�+S�V!��H�r�2=�a"O�@�&��&oFa�qg8o��1��"O�Yd��!��4s`��3\d�|�"O�������z��A��I'~|ha"OT��U�/Yqr�Yg�˶_(�3"O�|��ēvN&=*d�[**r�"O]�%G��_Vmj։�" �T��"O�����>t�4$	G�h�r�"O����ijdp��jƒW٠=�D"O�P�>�X��I��i�w"O@��J!rO��nw2�"O|p����`��њ��WaJ]�"OL��dךa&�ȢgK�<F�x)"O.����Ǉ=J4��e׽Qb(�'"O��!U�������$�t)��"OZ�!�J�PD�*e���v�"O���P
� ��p� ��|"s"O�� �cڵ5��T�v٧Y� ��"O6��V�A������-[��X"O������_� `����=�l9�"O�e�F'Ӎ�>%�A��*\�dő�"O4(��\�=X�P�$�B�8�"O>�q3�P
���jV��P���8�"O� ������MS(԰3��0�&�
�"O�,a��8 ���Ł<<��C�"O�e��e�F%0��Kl�|qje.�k�<y�G��P�h��)� ��!��c�<��G:���c�?2��g��_�<Yө�n ��&C�t}��QW�<����{�H2��Z��e��#	W�<���D|.-��Iː�V��)O�<&%��[tBhsDM��"c>��.M�<���y}�E��'������J�<��C	���9�Q�9��H�A�E�<���އa��f�:/D� ��\@�<Y�H�tgX\�Բqa��a�Xv�<��h�"&U�ӷ�4p'�T�J�r�<Q�Gx�1�Ԭǅ.m�tˆr�<��e��/v���l��z��7a^�y" ֞6�z��W�8CZ��bTͫ�yr��$t�9Z���@�SW$��y�J�Q��=�' ��ly�e	7ǖ�y҈�=6y�T�4��j �KL��y")�O�e��Ț�v
L���ϴ�y�'	�TK#�Àr:�U���*�y���4=��9qbk�)�n�i4c^��ybɘ*-k(4˰�׻z��Z���4�y2�ֳmQ&�7>+~�q�R��y�*˿Y���p�Ո0�=���]$�yMe1���5�ۻ,��Ca�ʼ�yR\�xb%.K�VcF���ޝ�y��_(����!($��B�䘳�y���N;��Ȋ"�6y^>���ȓ� �c�%��ҢЫ142�|��D�܀0��ƛ1��;�%B�*��e�ȓo|��T�pe�ȱC/�"#�����|�F�pp�Z,c�)t�R�1��Ѕȓ��۰�W6(,q�ܶ:���ȓz���d�{�rE���ޚ]0ꍅȓ>�L��w�K7>[|h����~2��ȓX�����9>��Q�VF�h���#-na��"'w���#B�[j*Յ�C۪ �G㢉{B'�#�@��"���;�8�9��r��@��Ic,��2̛�N����+�G���ȓ9�`Ö�5z�0�E�-.��ȓ5����C-YJ|��6&�y�`؅ȓea�t�4�`����f�z�\@�ȓC�\�C�!�,���թ�? b�(��~V
��(.���T�ۄ_b�i�� 3:�@��J�k��Q��'�>=lFM��)�遠H�?<��(  ��4;����\{�m���%��!(i.,��x����u+O�9�8	*��&6�\�ȓm*�h�+�h�%'�C�`�ȓF�B�S �>m �S�E�%��d�Tչ���>��@j5NSV�a�ȓ	��@2G#֯A0Zp3E�ȲT񺠅�4j�Л����<HjX;�n�-%$��q�pX�)�r���"łħUY ��ȓ+���$��7KbphKaK%g�襆ʓ&O�ca�\)$�f}1��ޚp8C��"D�i�P�YE���`��C�I�Rpx���G�[:HC�	���d�=r\5�c+�+l�NC��:E!�l���D�0�*�$�X�1�2C��-r>ށ���9��Z!Ζ6"�B�)� �u07dLV��\)qgX�c�����"O4%y� �,f7���5�AC�挙�"O���U�Mbi���ˏ��e��"Oh-�q�]�s�؁!�(`��
�"OX��Q��&k��x���>K�"Q"O�l�6��:n#�E����/)��"O���Ӥ�咀̖7�d�25"O�X36�����	�1iZ���"O*�{��
�F���R<.Pę��"O:��p�.��X��9IDh	�W"O�@�ݱT�D�#"τ0B=ڸ��"O�A8�� Py ���#�=��p"O>��EK�r���dd�:dݣ�"O�
V��#}�&A�A��$"O���p##��X#CO y��02�"OF ���/lɹG"���8��"OV��SǘU�@UÔ�M
!���"Oʴ"����>�ZEnQ��!��"Om���y�� �AS)m�*��"O�@�d� a}����F�}qP�{ "O��z�`��:Z1�1�4jq��R�"O�9��^� ���)�,�z^`S�"O���@o��)��8&�,"t1k"O\	jQb4v���t��)Z����"OtQ��F�Oz`���
/(��XD"O ̠U�ך(� 3���1����"O TaQ)<��@$ͨ��0�"O�|�S��3rL���	��a2@"O�m�'���h8�5p�˞<Urp1�#"O�ei��\?5Lf|�e�/6f�1�"OH�6����|C��dY�M��'�vU)"�1Ҷ� ���{�� ;�'��Ms�#��0����&As�� ��'DL0!��8AF���+�B� ���'�6!��Oƻ�:��f49�b�'��I�蕏!jLcG�S^�):�'����9?8������!g�4�P�'��0�g����A���U�+�''&��n@�_IV�"R��#V-��(�'<*��w�� {3:Y��풛U���C�']@�s�C��(�6�6EU6Na��'(����FFC7���f]!t�hr�'ӌ�8a��J��h��e�@�~=�
�'�$�r��"���SQ�/$��	�'ǜ�� �r�0<q��:l�L��	�'{H6��F^�I����Y0
(��'
B<J ��J�:%n�%O);�'���D�t)��J�p:4c�'�t�HGON���;Q&�2V�\I�'3�jJh$�@��(~Bt��'���P�n[8efPiVn��#ߺ�'\.�hd�"�
3 G��t{	�'D��B� E�r�x�%d���!{	�'8lE0�h��Ś��ɨh�U+	�'Q
D���M�@L��	�d�s�'�����6p�b�8i�C�'���0g� ���HI�w���"�{� �+f�����)k�� �4jO����6E��{�>�q nƦMX>E��\�$��#5D��<�2M�+w�`��X�80B1᜘J~�"�� +)�B���y|.L��D!f����R��C�`�� � L�Si�8/�T�p��QU�؄ȓp���	2Q/:�����BZJ�	�ȓ"
�#6ϊ(����N�t��S�? 4�(��M�{����A��U~���"O�x�BCXt@ x4JLZdH[a"O*�PkV�1鵧�Z娄�"O�{�K�N�r S���<�jU�"O��"pcԪL�`-�E��F��12�"O=(�#��r���%�\�'��!k�"O�ZB���6��< ���4)��<@`"OdHJ�%�!z���Q8;*u�s"O����ʦ;t���/8&�)��"O��9���rjVe��4��p��"O��Ig+�Z�48�րj��ٳ"O�л1�S�v^SGB�'�8�%"O�X"EI
[L�P����|���"O8�ru"A'�4���ړeX�"O�Q9 ɕ6Auz��4	F7�ԃ"O>T��<�<x���Ҵ>0܁+�"O��@�������+�� ��:p"On ���»	�V��D�V�<ة�"O��Afޣ:�B�`�B�"����"O@}�Rƌ�,�l�xD�˰HƩ�"O¥��ȳ0A���E��f�p�"Oj�3����^2���t�J��!�"OF<�B�ۡL:��1A�2��D��"Oz��w��L��\��6�B�Ip"O��,8$T�0�J�8X�����"O��ba�6���ȓ�=Ϯ���"O�HvɆ�*��I���Z-�*���"O�d8��ѯ~��
⁚������"O<�eJ
���)��,����"OMq���A:B�i�+�D4u@�"OX��$4K Y%��8�HA��"O�(���.�4c_�mS\��A"O�Л&LBx����G$]�6�@�Z�"O~� BH�
�tʵ���F
$)�"O�8��$ӯ~ۄ@��0y�5�"O<��c��<w�| �C�� �i��"O�1�.��OA4L�RA�5�*U�"OF��s��)Kv��@^�h���"�"O�հ���"ك�mg^y� "O�<����jn�y7��3I�QR�"O�<ZфA�C�> ��!Ɠ�F�P�"O�u"r�U4��< ��
=�4$�"O�	��G�;���g%����e"Or$�s�%�d�j���!n���Z "O�( $�3Y@�K�b��oĚ)۰"O|A����[��	k��F }&~�HC"O�ن��#"Phy�Go@�BkP"O�� �lY�B	�
"O��2{� �"O���@.J���.�����"O�x�S��� ��y⁤?1!jay�"O4�p@�P�D*,���G�bcq"Ob@ABb�G6Z�rhف<���4"Oޑcw�Jr ���W<�P[�"O��҄�F��Z%�
D!�l1"OX��E��}
��',��S�"OP��+
�b�[ �R���"O(�x6HM�>-��ȥ��~�.��w"O`5���ۘ~x�P��� ���$"O���5f��0��5�p�Њ�*��"O�qCo�1@O��^���6"O4���T�[����� e�HY�"O2Ũ�L��pvl��	�1�(�!� �jx�!�I���!��.S�~�!��6�T	ӣ�K>to���t.A�~!�� Lqv��n���c�k
�5� q#�"O��9Q)�s���X=(� �!�"O�)��oZ�=tzl��$��bY9�"O���͛0(G� �aM
�`���"O:|�6lS$w*���G���{�(y��"O�ܛV���[�ͪ�H����"O ���a\�R�x����5,�H��"OZi���^�t�V������s�\)�""O����&R=QqW�G��Y�"Ox����c480!��U#�8�f"Ot]�gU���{���.�(!�5"O������,=�r���R	^圅Q�"O��Yp,��f8F�#a��Q<��0F"OR��Sb�El ��!Һ_#��b"O�t���̔2k��Ӈ��S����"O"��ꑢZ��EI1AЬm��Y(�"O\��R��ed�$@<Q��xAp"O:�U�;=���uL_���`�"O�h�F/�6*�r���ٸ)�z���"O��Z!�BX�����3<�X5�b"O�ə��G�]@ťO�=��H�E"O������ў1��E�&7lƔs "Oj��Dʏ,^���#E�tFR��"O���Ki��.F��U۲"O��30L<�A9�׬�܅ �"OnA3��ň36���Gc�!�
��`"Od1�)��WݤԂ"���b����"Ol�3�N�4��1;@�K=���j#"O8���>h0�yPQ`@<�$P�"OT��- <]���V��@"O=��.W4�\"6f̖yd�"O��D�Kb���N�28�q��"O� K�`��P�( �s����DA�؟H��I��.#���i^D�:�%ԁ��5��'%��0����{�Z)j%a���(����Y���p�&�26��;e(��Y,�!`A��j�<B�Ɋy+�#�JG�A��� #BN.TR`7m7!$^�
3��?V�D�S��M�w�C�F�|DR��W!0.z,��J\k�<��
N��p]k��H��0Q�	^}��J+�򁒀&��:��x��Q�&��Li���w&]�w��0>�7ႜoI��G�q�RlzA��#�Buۂ&��]]�X�&Ն��?�F�C L�x��!��|[6���I�'���3��� ����KTWx�O����ڴ#g�ԛ��[d��@��'��M�B-uʼh6��O�qђ�Ȥh4��P�ě� �h�p��h��$^�v�}��0M;~=�� 
?!���1P��@�G�)����T??�`��,4�pE�6H��>�L����ϨOv}:$#Շf��Yx6f�6$l�� ��'O�Mӂ��T���p@2!W�{ 5ӄ8����Ln� vA�G��~"˅�iv�C G�W����X���'��x��WΦH�AU \^�p�~���K4�.�*����e�a���w�<�eI
�Jq�B�˟iLܡ���і�r���l������:;�J G�T�O��Z���+LO����3[R�9�1"O|:- �-X7@��_Ũ�j���3Qr!F���5�Y�Q��&��<�`D�#���=~a��K�!	�<���,ut�2 ���@A��)��Y1l�����x�Qb&MY�<��q���h��XXԆ����#���Q��1sq�'��&�������O��<��OX}#�O/��$ѷj��e�'�&^���'�D���W�B��ັ�� �l!�O:��ǭe���hi��~r�LM�AQN�؄XE���y�MO:0��͇�%��mh�	��MY��Xl��.C���'�X=:��VZ�xXF�W6\s��#��=b�`���99S i��)V�'xP��
Ԍba���7�f���"��W�4��V*Ž+#$��'�7�"�~DK�@_()%q��-���5�*QW�B]*z��g"O� �-����yYh ��8P&�OT���R;@h��&��}�ԣ�X��1���($�5Q#�	f�<� �ߒIIDH�l���MA�eC���$��jra؀
;<OX�ha+P"Q���Z��h����'������V�M	f����!�� �Vg6J��B�		H�����"VF��pl�8w��B�	�b�h� ;?�ȥy�eՉv�B�ɴ?h����$*G������9bg�C䉓#�b��c�� @��9��N�x��C�	*S*��3J�,2^�����Up�C䉈x��)�qk�"l��逫�m�C�Ɇ�B;s���OH�Q�E�;"�C��G]�qg��v}��0+�5/�\C�	���d��+ �x �!�͋?�B�	EO|���*.��I�X�C�ɤl��	�����T�X����W%BLnB�I�z}�%sC������g��+�B�ɺ$�hq�W+Fy�L�� R�[tC��6n�&仧E���JՉT���~*�C�I&!�4a"�ǆ4�4Yh�j�8M �C�	�Kk�E�ś6��D+q��l��C��3#����r���|�͍${|B�ɵ^'z�1T��*#?*Q*���HB�	d����'Udiq&cɒ��C��/
l�%���M��*�����9I]�C�	�BK�!SO]�/\29z�A�pG�C�I�U	��c`n��]'i���s[C�	�r@h�F�8!�u�S��^��B�(:"��%`��IR�h�%@��C�ɝA���s�+�kJ@,Aw)�6Hk�C䉡p5̑����R�F�\>�C�I�!���pϑ'\x�-*��	-��B�	:)U�   ��@;���ƈ�q�B�?=����A�R{if�CW�F<rC�	�*�xܢ�D�'N�T��Y0�2C�I�U`8���/M�c����;6"C�I�hZV�q��]�E�bYY��EJ
C�	�+Ը�TjJ�x�p�+C�[�K��B�*l�P����U��XE�
hlB�� \�,��%m��=
���FV`B�	;#�^��4�W�Qy��҈{�&B��3I����Ԕ#W�IP��  �B�	�`n&�㵌J; ��@Bf��B�	Dt��# FӔ�^�Hā(K>xC�	1+�h6�R�5����f�"�B�{DR\����дp"�F�lC��8I`	���J���h #�̩za C�I�W
��XD0�ȰKr@J�lZ�C�	�f���H�cD�L�f̓!�(ZݼC�	�Y��D���3'��j���\B�	�̫B��)`���BB vB�30�#���J�-���h�C��#�`� ��(�|�dʇ4��C�9����V���"�VE�5�jB�	�@):h��ĈA�r���@A2Il�B䉈aB�蠅�s��I�2K�oZ�B�Ir�����gN=}`1�����
�hC�I�h�����
�
@�+J�2C�	pO\���
����T�H�U�B�I*��h!$$�Iqԍ��1D��B�IU$Q��a��!�DB��O��d#��ͷ/�J�� �0-~
U
9�DXyѢ��6�֔7��� kƷ �!�d�&d)��@RI�XZ������!��K�m�|��'%E	M9�SSh �T!�� ��%�$��ղg%� :mpI�"O5��ǼJZ,�֭,]bR�"OX�'�	?��L@0_H��V"O�9Ʀ�7�N��
��%.�ə�"O��X�l�1y�Bx�ŊŁ0���{"O20apM1H�بke�7<����"O�  �"T�Zj� O�!s"O���tO�X�r���� -��E"OMkv���6�15N
�l�0=��"O>�H2�E.?ɦ��1H�>{x���']ޱ��% �p9��V�2C���	�' By�rO����(sɟ�}Ī�R�'�4
���R?�����֒`b���'��������2���Pr&P1M�n���'���{'�\Hڝ� �JJnI��'�H0'�M�%֦���Ɣd�c�'�V5
��8P�c2�H��Ͳ
�'~���G�+?���K�d���Z���'�ȴꅄ���ݡ�h�� ��':��q�X�1;�}� m-_t;�'(`�V�)z⑌U)���'���L�PF�X T�U�Gj���'��R�+]4Yy|��scvf�[�'��:CC��#^`�R�ƍ[��8��'gn�q�(ٿr��K�F҂W��
�'S�(����6d��1[�H"d`�'���j�Z�����v��0(��'�*4��o
ryЇKO�K��a�'k$t0�'�>Ph$�LXv���'�X0��ti�� �˗e޽��'Jl���`��f
�}f���'�l�f�D�P �a���W<r/�5c�'J�}�A���b�T����(p_��c	�'�.Hk�
[�_h,�+��&c�L�'~��ӭ�4Pt麤�^^b���'W�zW�<`mR$z$%.S�Z�'��P��¾jX�	t)O?f��#�'��;�G$ p����X��'�vh*�$ƀ6�����ފ@� C�ɴ�v1:�#�Y�lA�k���
B�ɟ8��������=0��Կ%T�C�	7,xYB�%ڋ'�,p�o!GC��&~Ej��e#S�4u�4*L<W�BC��/�nYj��|��9K�"��
�C������&KȞg۰�1�%�7]|�B䉀Ю<0$��#�x�q�S�B�	�,H�J3e�3�J�i���H��C�ɩU�R��pmC,/l���רB��C��f���)� 3���+��U�w�C�I�+���F�(Δ����G�@B�	8c����������PG	�� �ZC�	e�0Ya��#@ƒA"Q��u�C�
e��%i"�ԃ'F\�Pb� S�DB��3m;��Bd|$QQ�c��G0B�,mENݩ��Q�R�=."�z1"OZG�ѐD�䔳
�1<�yp&"O"���ÕM�-���в`u�tz�"O,���đ	q@��	���1~���"Oz�B!�> W�!je`4����S"O�x�Ѯ��= �4�o�6X�Z1�2"O��ѱfF�R��h�7L��0�"O�ب"�X9�.-��Y�:����B"OZM�cB��&�ȇ��Z���f"O��p�Ӌ���3Ai�)V0t�1"O� �<�h�?c�dٺ��Ƀ	(.��"O�UH��W �Ƅ(e���m&�QCW"O4uQ�H�Gˆ܁���=�Z�"OAB�k*9�2H��Sꔱ#"OXTZ�E�&c���H蒷.�j`�"OH`1��z��L�'�G�%nܕ��"OfĹV�ú5���å�Z&�2�� "O�L���mW��6�� �h���"O��@� }9���!�.+��b"O�,�eoJ3u+�-A�AB�Y�a�"OxԨ���9T¸����l��"O��k�mѡi�0��ŏ!f�%��"ON�[v��\~mU�І�!�"O�I�B�4<dh���k(��)�"O�����N�=�^�+�LN���I�R"O���$+Pr�|�Q�GP���5"O�l8`��ƊBt�����"O�*��B�Zz0�	'HĢ"���"On�B��
�`���iS��.�,-�0"O�I�͎!@j�)��EƸ	TPá"OP�b�Ķoj�xR�\>&��Zf"O\�0A��e��]�F��#��t��"O&�@c�N%l��`p�-�7z8��V"O����zJ<���{~]��"O\  1��% ���3���q� x5"O|���EP:"���RĆ�*x�f��"O��P��B�M�D+�+	�yz�<��"OV���홨e��M���+�x���"O�� /e�^�*Á�vvR��"O q)'��6s4py��ߘDt�J�"O����Ɉ�8�ԘY��?v}����"O�ȴ��UP�K��ǺGrLH�"O�RN�.#�F��ƌξg�8�"Ohd��c��[0�k4�^9J� ��"O�4ȕG0m,]���&j�$�"O
Pg���� 7�>M��"O��pH�ivi���ф_I(X�"OlTs�+ɪ��)Jd�M��(�"O�	 0���}��c��-a*l!�"O��Y��#DtͩDDO�DVm��"O���A"
��Ѣ��8E��"O�c��`���+A%I�P�4"Ol|8��L�£��u�8��a"O��J�":`s��5�>�C5"O�E��%�-fF��pCAY{<q� "O��%���=YG��,��4��"Ob�s�F�b��4�N�Bt%�T"O:i×��"�,)Qubߺh�h�1"Ox�+W��50��\Q��5H�S�"OTݘ�Ǐ�	Z �Z�H��s� U"OXȠ�ƷF�$�J��"�<��"O�U�r��W�ځ�#,�#�<�z3"On#1��IBf]#���!1���Y6"Ol8��)��6*|9��\�T�&|��"O�ij7�G	�-�lJ6���XS"O�=�'��?�ȀJ��kr�l��"O�E����$iМkD� ([������ |O�`g̀�PEl�Z��V ���"Olp�CMG�c���*7���0����f"O���r�Ղlx�5	!��l!03"O�A9%�_�3��U���γ�ͫa"OL�ч$��>�z�S�'̓P��4*$"Or]x$�|vPd:F��3/8Y�"OB�`! �%e�UXӄ�+X�X�3"O� ����_O�1A�O�3�6	c"O�ѡ� ����C���:�"O���jS�*��!+�oD�y�n��"O��0ƅ��n�@��q�P/c��|�@"O�!c��o�F����ʡ`f�y��"O�%b��?| �iw��;���C"O�!p�ň&�8T(Cּl޲5�&"O�I�P[�f�~Ax�%�v�Fi"OVi߽sG2��5�Єi����v"O.�f	(n�]ѷ�%*�଩�"O�9��h�E��.Yj���R$*�y���*Ȃ9@�L� ���ɂ���yS�e���
7.�7D�H���y��5k�pv-Y�X�ܼY���,�y2	P�B�	V�Wu�|6AU�y��Z�dZ$�3���I��ϊ�y�'D�3�&�Z�CM�Ph��
2�y�*ǠL���3T�=4�LI�B_�y�T�1쒌)E �.9rΙ(و�y�
\**zH�i4N�/qh�p�f���y�΂GK�т��Ʉ�Y��y�c���\��_�zGй@���y� �^N0H#�(g�,�4m�"�yRjC�b�����2�:m9�@E��y�� �~�����~�0\�����y2�+ ����&I	�h���D�R:�yb���@� |9 �Ӭ^�����yhH` �ɺ[�&9B欋��yRЪ\C�КL"��5�W<�y�È�8ā�F虽I`�R�U�yR��@�,�¥�D�<8����y��1*��y�`eP�A`�@�5�y�L/YZ��b�@B�=�fH�Gh^��y�g�7BtB�
ؼ�"&�ܫ�y�+@"~���B�[~��8��ٗ�y�`@���`3��q`F����y�fI'{BR屗n��(���y�C�K���7e��� H2����y�B�S���2�#� wl՛A�ɹ�y�) �?5Ҥa�Mޘ<C�9�@@ �y2��(�^�ȑC��.��Xea��y�nB�G��#���t[t���y�Iťg���`�#	UV$`c��yb�K�oE���G��v�1�y�f��Z2���-�)��,i֦�(�y�+"h���ԝ-Z�S����y�"P��8h��,О�
Ub��9�y�R4K����,,(��/�y��#7"b8X*1��jT�ʋ�yRL����a��'їv-J���y�����P�GU�FXR�o֩�yR�� Cx �%�U��Q�����y�헐%�dlq@�P(��g�C3�y�'�
$L�� ��F���F$�y�Ď����S���o_T�RB���yb-��4Θ��`�&d߰�iP�@�y�[$"�Lu��OB\�\��M�y��u���!c��-C���M��y"�%0�������0��i�M�3�y���P\��0�%7�a�&��y���l\��f׊(��� ��ʝ�y�)�6�*dI@�L:%�M��T��yB�g�~p;%,M�"���h����y"H��h�-�mS� q��	qnְ�y
� ������~��Q#@��`z "O F�1L�����ϖP�
��1"O�Q`��ڬe�����X#��E��"O���p�DVS42d��h�l��B"O�ly�C�
x�0��e� �"O,�c�ETa�Tj����OaC2"O�DH1��1�Q�X�S��+�"O���KB�`İapMD;@K��""Ox�â�X�ޙ;r�U�>�P0t"O�}�0�n'\9� בj#�Y�"O��U�ELߐ�J��ɓ;���f"O6(�.]��9b��%P�4�"O<,�M�FX�Js(@/x8n��r"O�PV���Dc�d���87$0" "O"���E/] P���tq;�"O��y��<����ƅ�<#�%cb"O&87�Q4�X��e�@��2!"O�!�e�D���'E���j��"O6��e�Z� �2��F)P��9	�"O��ɣ� `�:���ݠ���P"OD��r�ձ�N�9��W*�(�9�"Oҕ���2��qH���%)���:�"O�Uad���"��$=v�R"O&�;�,Ʃy��̀�"o���q"Od�`2,EN�f��ϐ&pZ�Y��"O	f��˒��Mʕ<��d" "Oj��O�K󦁡um���t�*�"O�UQ4B� E~̌��Z�L�Pm��"OjY8e%��+��T2���V)*%"O���&���rVJa`��Ř8$��S�"O��C�R�aU	�h�
i8p�u"O�؃@���y�:C$CJ-�Q�c"O����r9.�$�-*�4�c"O�-��e�0�`�$�ˮ����"OL������c��9G$\'Y�p�A�"O�R�(O�-{h�0QHI#��0�a"O`��Dؓ1F��W�@u���U"O�}���R�~��M�(��p"O2E�[-vI<I���p,��"O�؁�g�"J�4(wlM7c< ��"Or$�W-W\&4X��
7Qb�8�"O¨��3��]��T�?D�+�"O�r��
x���]��\���"O��`���P�m��lY$|q2�"O��:�GY5��[ье ����"O\����|�z���T�h�\r�"O2��we�>G"���R��AI6P�w"O4,��
U�f��Z�Ș^<X�a"O*@J����,�� �ڸcB��I�"O(գ��6x�� ��|7TiRv"O���4���:��gT=O42-��"O���/^F�2��q��Q=0�Q"O��AʤlE<�I�E��3t �"O�䈥hR�X�J�(sfޒG��i�"O�h�Տ�<`��ۇ-(�d��"OtqXSL����ዑ�ֿ|%��`U"O��3�Q�6E���!H�,2,���"O�`���3  ��J�.p�Xb�"OM�`��pk���H�.T���a�"O�03��"[	�	qg�#r�Lr�"O�x��i۽Kz$I�,2ѺUC"O�8������m�#($�*�"O�D�p
��`^j� o� "m@a"O0���!D�Y���e�H��"O� T��6/�n�*{e���S���"O���@BW�d�.0Xd)�1Pf0��"Oj���`�;.d�S�燲p.�c�"O6e*B�6ea� �%f�0#ZD�"O"e�W����Yҡ�tJ���"O�����/1�X�E���
4Y��"O�LH��(s������?X���r"O��I�e�5���
D�H�=�"O(1��� /�n��F2JK����"O�Yӄg�-�B- �0?�T5"O~�;dd	j�b<���ڃ���J"O걪���<-"=�ց���9d"Ob�ؗ@�k�В B,+a�Њe"O�=	e�ս��btN�,�\���"Oֵ�Ł�*�TH��������"O��ɋ9�謰3��(?~|���"O8���e�%J��=�Į;8��`"O�U�B�	9�x�(�N�z���"O����원Q8=h� Q(��jP"O�=��$B�.��}(�9r���U"O~�Y�ޜ(7�[�M�8ek�APG"O�bW�I(�S�A�~W82C"O��"�5��8��<O!��ٴ"Oȥh���6l�T(k��фb`�"O��(�"��?�����q��IY"O>,�G,�)}��D�띄c��3�"O����H�?M[* "��+� �"O�{���u��噠	ݑڤA)e"O,����
N/���7. 7�$�k�"O셋b�Y�nH�����x�"O�0�B�3�auǄ�x��a�"O�Q(�S�hs��"?�Ja�"O��Fc��72���S����"6"O�4��²&5�u�P�=�p��"O������F�Z��׺
�<P0r"Oʀ9�FCw���X��B>a�(ɑV"O�,��+�C��G;%�2 `�"O�t� (ٌ�����Q�:<z�"O.|h���1F̠XAˑ����"O<|��e)'��$s�H٪�޽��"O�D3�B:����6!��� "O�!���˶G�4�3��)>�XKQ"O�q#rW�=�d�J�i�f/y� "Oh%Q#]�-� ��!.�[�"O�����/#��(��(�PX]P�"OۨCO��]�ӂ7Id����"Or�7nO�B��H �k^�f�!��ɮ*�Vx��mZl�{��Y�!�Zd�
�1Ǟerh���f}!��M�.n����&P�N�"��ޝ<�!��P�h4Q�*ԋ	�T`�C� ��!�bX� {a�r]>d��Ğ�!�D�|�cf� HV�C�-#d�!�Q�!v��"��-\���)�!�Sy_�:�'�BU�mjg�ǺL�!�ͩ,t�<�d�X-,õd�-�!�Dʿ���y��$��0­�s�!�V"�������(dw���V��.!�D�^�ب�`o
 \�5�ŊL�?�!�/O4hm�1��[���ELT�!�dC�����D
�`�x`B�*�!��7p�4J"@.I~< � iV�!�ĝ:n���OT( ��зH��!�D��I���r�)|aB���şW�!��  5��ӹDp�mB�&���lإ"O��	pH�-g���r��O��0"�"O�l+�׸���.���=�!�T,="qG��c:�ܲР�9'_!�$��Zۀ���!�,:~4���#\;!򤚶Y#�h*���0br���B(!��/ �h�k���7p` ��!D�W$!�D^;JX-��] 4����!�L�H�!�Խ3z%� bK"��c���!�T%MTV�Q��c��ԑ��h!�ƣt4�׎�l�b���a��!�dŏQ�b8#�
�8	�L��g���X�!�-7r�U�$Í2�PP4��,�!򤘁T@�5�t��B|���9�!���>
�ӱʓ��J ��F�2F�!�����peį���Q �U J!�F15�P���䙍D?05�BQ�~3!�X�Khl��I�+Dժ�G�'!�DΜZ�h1P'E��n �4KE�C�2�!�DR�a:x�SE9���R��=n�!�D�4MV�����^��3Q
��7�!�D�Fp���s�I�b���P2�!��ӿ�n����ԦI�RP�q&�DZ!���-�Qp�O�&����6���/C!�䟊K�V}�F�ٞU����v�ǴL)!�DB�b�c�eA�����F9!��Nޠ$�D�Q�B׬~[�9��"O�����S��17!Jz)�x��"O$�Ac/�0ZKF�0���^mZE�f"O�͉�јBDr����U����"O���B�?$���R8A��i�"O��Xs�[��-I��Y<�P�s"O�E�C�=HR`+b�9I�.�"�"O$���)O�+ǀ8�E^P��,`�"O�q!FI��S |���H"����"O�qe�<3bM�\�*�����"OFHS-�-7E8;㡘�θA��"O�p�`�l~�=�b���2�X�`�"O�(�q�n��1�.��g�l�"O�C���� :28혶j��R�"OT� �'�72�Q�@�o�rdv"O�	��ʞ��^%��#%�*qs�"O­ ��+ui杺�%@�JA)�"OD�Pc�/H�T�R'�&}*MѴ"O^ar��ُv��TbG�3Sf���"O�8����&K7<u+4%��DO2�c"Oz���Ƌ�Ā�.�JD�!�"On�9V�ڂm:b��C,P�"O<=J���9�6�'Z�%Zv"O����oP.Cy$li��S���Up@"Ox�i�	��  +�=b�"O�p�C�(T< �®� Hnb(��"O�q"���,Pޠ@C��&���"O~K�mU#/
��@��:SG�Lq�"O��ӑ/_�maz��eΥ :���"OvL�g�� ��݀L���C"O��H�Q��Y�"��X�ܒR"O�Zp�[�,A�)�g˼s�(!�s"O�0ⴅS!mW�PP���W�f�)%"O�1Ğ�k�"��'�<e���"O`���	��D�T � �Q7"O��"0�L�s[6L��ʛK�ޙ�e"Oȭ+@E�� ��so�p�f���"O�j� I�4F���H�
�:�ʗ"O� �g��.e��R�nM�B�<hʀ"O<T�%ERT��D�Æ�3 =��g"O Q���Ӓ#mҲc�/&�	�2"O��sNFRfN��@�_�)���"O�L��B�w�|z�B��'�壓�	����Q	*>���I\�#�����ń�^9�t'�4_�qO��DZ�y������	�>tN�ٔm<�tE��O��\#B�nD� E�{ A��dʻ;�8�9b��zRb���%)����'OS�0�S��Ok����͝�vҖ�Ez�L�'�?��gg�OU�vȍ�e&�%��m��_ ��Ӫ���$9�)������ª2"�5��K�\��p��$}r'7�#՛gg�v7�\~�F�a�c�4OPI�P�K����0<僧l�՟d���i*��W"E���ұ!�2R=jt��"@~!�&oG�/ B��J�}�aQY_�ʱ�}����M�&@� d@љ�'�9�pl���s�"��1��3	�Ċ2%T��P��k���(�k̗-;ɠ�7�É9��4��a��t��v��?1�/�V�'�?7�,:2��V�ȱ'K`1En���O��=��}�(�.������^'�@�@&Ό�(O2�lZ6�M�K>��'�u��!�L�FlE7^g�1Q&�!w�����YF�i�ay"O�=d�������3zI �� H$8�� aT�ol�);¤� ���)'%����7��h`l��i&
����۵s ��Q�&��9����:*��2�V?1��D۫K���p��lܖ�{c�W Oe����
6�.��I��M{��~�'q�tY��S��@��5�vg�hy��BF%D�Ъ�T�K��C�*L>G��T��-5v���~�V�O���˓2Kd�딄�57�T����I*N��t0���&�vY����?	��?)5È��?i��?9�eI�dGF�B2[�K��R�A�p�p���e��Т�#��شC��*��,Lqfb���r�S$I��YnB����2��0 ˠq�(�/1�:���@�'�%
���Ms6.��� ��0r�И@@��2g��O��D�O��ʧ$t�3l�.�>MpGB:,�eFy��|����"W����"D{��W�����	�M���i��I�fOU�4�?�O|²l
7�j���п38l�{!e}ܓ�?���Q�e<�8!4�*�E�eіd4�=����ᒅ+�Ѝ V�YT(�#=كjɇf�!�sI�F����,L�#��	S�4	A�A�+�9�B�bɑ�C�O %l�/�MS���	p�X��񈘿Y�8��8���Iry�T�"~�	<E�y�ć��Y��u��]�J2���Ӳ!l��] &D"#،[�n�e���Ѫ����S�۵�Mc��?�/�j�q�E�O���t����� �h(���d�a�b�^�x�ʔ�a�V�^l�LA�*9Q05cFٟ�ʧ�"]c�~UZ�MY��~Hӈq$L�2ߴcD~��Ї8�����ȰP�Y�W�s��ht_�p�m��k�,Ȑٲ4/h���k��']Bι<��y��M#��2'<@*��ީ)��W�I?����>a�EҀF}j��Z+���+QC?H>9�i�.7 ��ֺ�uB֜{!�x���d��b5KցZ�'Va{rήY   ��   �  [  �  �  �)  \5  �@  L  hW  �b  �m  �v  V}  +�  [�  ��  �  8�  {�  ��  1�  {�  ��  (�  q�  ��  [�  ��  C�  ��  ��  ��  A � �  O �$ J- R4 �: �@ �F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1��2*Q��'/�ܱ�Dnٲ�0�rG-E�ws���ȓC5p�yaL�!	:Xy���J+K��X�ȓY�h����a�$��'AM�D�d �����f�6n�4�B�j�?���� H,�&��+�b@Q'n�%+Z�Ąȓ6}ܤ�2c��p��������\H���'ba~�a[�:$���Ӧ{�2����y���?Rچ�q%�F�	����?�'�`�)Sn���D$à�S�U[�'Cў�'��^p�A򐡋0+߲5.
�ASl��W��F��6SU�<�L�As�A�'y���OL�=�O��xI#,�(�C����k	�	��'tD;Ue�46�8�q'>jæm��'g�0�¡��kI��0p�ј-�|�+�'��pv�F�m;�y �RuK����'�,d��o��۰�B���sh�0J�O�6M'�S�O�B��t��U��f�����'��p�pL�<`�н�D̑",/�m��'j���7K�7nfpd�5�ƟZo��S	�'���A�/�,;Ϧ�0�V�SFxT	�'q����
:8��R�F0}h��[��HO�8���_>bW��:O���"O����
`�=Un�w�\�#"O$�e��"Z��S��u�4�s�"O4��G�|bI�c��.E���w"O���׫U;�X����,��[�"O¬	b�2x�~!�W p5�R"O�}i� �%z�R�03�� a!�$W,zb��Х�Z",���fI!�D*8v�x���%x������!�D�t��un��u�F��7��7�!�D�sp4�b���B�j���b�!���'7	fE����$���r'KI!�J��H���ӓI� ��$p"ONQ�	����B�Ŗ�j���� "O����KƢp몹���)y�>��"O�(%��z�`Z��S3�D-�""O�!b�-,l��1�^#"�(H"O���b&ܛ.�{ �KX��a"OyqsMZ	r�x&K�9I|�b�"O�x��[)*��z�I�R+�ԩ�"Op�W

�M4�X�T�#�q"O���֣̔T@-�S-[�;���"O�-hf��!"��*��=��"Ob@�&�� ����תJ<Y�T� "O�I��3�.՛0̆0Wڤ��'"O,� �nŦ2��\c��׃w,��T"OΠ�D�X*F>j�!���x!�(�"O"i����a#2����]�#t��"Ol sG�P%�LC����~�,��1"O� �i9���;"mލ؀ҏ3k2�`�*O�9{��5G��� ��D32ޠ)	�'&��S��?��X&�Q0�> (	�'V8�r��R�!�$ޚ)oh��'���N� �|@�C��0�12�'A4Z���rQ���G��5�����'�8�����<1�놦@\4 4��'�
�a��V�M�"��wn�f��A!�'�4�s���BaG ���L��'���KQ��x���п}��L��'*48"6�ř4$��j�xHe*�'hf1*'L�U�H��A�lA 5@
�'s0QR�,�1e)2�3��2!�
�'�,�X��_S�>�E1��I8�'I�̹0L�9|�V�{E&�"\����'"�d��[�n^����^�S��ţ�'܁�E#N -��h0��I	MJ�'t�������\ �a�	�GcT�2�'��mB��Y�N�i�Z�v.��'�25JCHA������ŉ�Z�~ �'4"��b�Q�3����r��D�&���'��臆ֆtaX�s �>;He��'t��b�Ņp���ʂ�Ł%� ��'n��E�V�n�	�)g&P�
�'^�� �O�o����AD�7
bf�3	�'���
��E(���K�J����`�'��C�K�!vDF��O�.ych�i�':D<�'38�8�@� ��-`�'!��"Ǫ߳殩��A�r�"�	�'�A�e#�3��,i����f�ꁱ�'H��Е*ڕY� {g+�]�H��
�'�vM)�敁4߆ȋ�ɋ�����'�h�I�T��I��7ts�T��'Al�*��	/x�؁��ш~�z�j��%��cu����I)t����.�b�<yҰ���%��@ɚ��:��B�I#@e�Z�D��YH���N���B�	WH@)��B����F�-RڐB�	�Z��aD딉?������5Q<C�ɕn�Ҝ)�j�	5�`�z@�A�JB��=3����P���!�#aRU\�C䉹x4�<�`g�%o�@�gH��M��C�|Ѿm�4p���A��	�z��C�	�oI���e�Ӣ���ٶD.,,C�ɰԵ�ӎZ8
/J`�� �N��B�	�Ѡ�0�?m<j���ӄ9�C�	0*�[fN�p*Xy2&荞z��C䉵c,����yCV%�!	�p��C�Ɏy�P�B!�ӸO�huh��H�_>C�ɘ�Υ�f$F���|�w+F�c
nC�	,f�:٢���1r���Ӭ�m�TC��	2t��!P�qO�51dݽF��B�I9	�̼s��A�^�������B��2`nTI��ǚ3��A�g�i�B�I���I{T�ր;H�)�ו\�B�	�m��9�����(��k����B��
|L=*6A_D��`��Qx��B�I7䶁k�o�+9*D��&�<:�^B�I�5M
Kp��$i�\B���&@��B�	���8��)v&���a.�FC��y¬I��˄"�Q�FB�'�`C�)r4�Ɂ5,�51x0����g��B�InZ�0cB/�8ao�kw����B��u��@�M �ϰ\���â5c�B�)� I� ���8"S`m[�"O��8S����E�'P�~��=�a"O�$�G��}݊p�v&T�_�z�;"O���v�אg}@8����=�4��f"O8�BG`Ѯ���+�>�6a��'m2�'���'��'�r�'��'c��N�<V�3����~h�'���'�'g2�'@�'���'���P���%\b$�����p��ԉc�'��'���'�'��'���'����@"�7�h�A j�6Ik��';r�'�"�'nB�'���'�2�'zP����ٖĚ��2ƘTc��'RB�'�2�'	r�'�b�'�B�'\��9' رlP.�p�B�=��9���'��'���'i��'F�'�B�'�����p��bro]*[�*}���'.R�'���'j��'��'��'A
5�dBE/\|x%CR"ʑ+�X�V�')R�'"��'�b�'"�'��'m�ʥI�F���Sd�W�P�8��U�'e��'��'r�'A�'���'k�h��c����6�ܠTV"t�c�'0��'�2�'AR�'�R�'\��'>�I�񯝘3h��"1�P�{d�Y�t�'�R�'��'`R�'^R�'n��'��1��� hT℮N�e����0�'���'���'d��'��'���'���/ˈ<H-0!)P?N���(��'���'�"�'��'��p�n�$�O�����X��>U�uA�fBa��WXyB�'�)�3?��i縬Q5����(v Q�Z4`v$N���d��m�?��<9��g0�a��N��E�����ˮX��{��?qgb_(�M��O��S��J?��r`7R6j�����\�l�"`7�՟h�'��>��U���3x�:�$�� f�Y�Nت�M���IO̓��OV7=�n@jJO��P˲�W�~9&y`��O&�dk��ק�Oδ�ڑ�i,��G�wxh�T���/�>���&E��f�\���*�=ͧ�?YsN
�S_BL1c��c�\m!�-��<1-O��O�m��u�b�|�EaϺJ[�h��Ĵf�
��x�?3Q����Ɵ�̓����8~���
wj�p7�P`C��K���џx 5bF"Q��b>y%�'������!�d=J�ˍpEh��� ��5��'��ş"~�V��QƁI�:�Z( ���  &9�L&�V�ڝ���Ʀe�?ͧt��ز!��9o\<�0bśP����?����?��,���M��O��S���c��P�Θڣ����AW���B��O��|���?���?��J�����A�e"��+1�l����-O0al�45�|Y�I�|�	�?9��ty��<8�J̈խ@�vO�0���v*6ꓞ?y��Of�'	��1��?��ɷLҡl�|u�կmԐU��Y�H�◽7%�u��}y�J�<QXx(���_Gd�U�ۀ9��'�r�'��Oq�	�M��)��?!B���	"2�� .D|\2�c��?�P�i��'F�A�>���?ͻI"VњVI�(jfV�Z�.T�+ф��4 ]#�MK�O�D��Ј��ę��w��]�!�<nhHT����3��tɝ'R�'���'�R�'=񟦴�CQ����5[P�`@ڪ�?���?��i�`�R�O���t�r�O�pb�gP�BJ��Qro�$q��{q�d�O��o��x޴��'-z.��0g҄)
��d�bbj��S;�?���)���<y��?A��?!�A+T*f��'E[�s����1����?���dM¦5�����������O�ډ��߫	��z(W#ի�O(�'�b�'iɧ�I�<X�$4 s�:r8�u�eK+.�f̃�*�ZɌ6M�dy�O.�����;�PؐDG`�:984͔*g��8���?A���?��Ş��妩qԂY�B��[T��FXD����8pq�]�'{7%����D�O�Xƣ��p'z=i�`�<P���O�����7�"?Y0-։TN�i9��*��U�LP���"%s&�hĦ��y�]����ԟ������	ӟ�Oj�X�"HiLY���7���@�a�^�S3M�O<�$�O��>��ئ�]�Z�3��O~�dp#"�1�Ƥ��Y�S�'h��x�޴�y�!��"ClQG�~| �����y"�@uH���I ��'N�I�� �I/ ��	��\+�����Q4t��9��۟�	ݟ��'=v6MI�G��D�O
�d��=L�i��)Q� q�n��"�.�k�O����OΒO:�@1ٟat����Ft%�����������~�o\�'B�.�	ǟh�� J�k��aJ�$�z�� �'����I����I�0F���'�5���V�-�T#�#��aZ��'77Jmaf�֛��4���uL�=hd9PDȅsX,I��3Ot���O��č�'�7�)?!r�A����1�p��#��J�����-μqϚ��H>�*O���O��$�O`���OP8�ub�=c���ڒ{4^,�#��<���i�l���'yb�'l�O{R�O���d�%5{����qo� ����?����S�'E�d���O5Z��$�FI8N�L
"�ļ��|�/O<ѻ2)
��?��6���<�vo���ɸ�!�!��A�֊�#�?a���?���?�'��ā��2̑��@�S�D�b��*��,��ؘ�ʊ֟�޴�䓨?AU\�8���L�I��~��!)��Z�\��3l�:~j��.��M�'Fꐨ�E�?aʤ����� F��g�ߞjnNxR��T�O��L��:O����O`�$�Ol���Od�?��T��+Mv�H��@M���� ؟��Iȟ���4o�+Or�o�[�ɕc������r��U��mn|%��	��0$���l^~b嘳}^�ᄨ5�&�ٶ��3�@MQ!�؟(Q#�|2P����H�	˟H E���&T@��\38�h��V�����PyR�v���1��O����O`ʧ�����l�;+�H=sR�!r�P�'B�듑?�����S�� ؂})����^��}�b�ԂH�-�wAC/K�F�<ͧr��k�t�~��a �,ʵ�2'��{��'�B�'b���OM�I��M�Qg˅<Ch�[ƃT$4����L�6^�X���?���ig�O�8�'�R��L����+ �E����K����'(�H�ix�i���j��?-�W_�`C��ՆѲP׍��J�t��v�l�x�'{b�'���'��'v哗��d(��TV��T�OԾ4�ش�q��?����O%j6=�a�tA�<�v]��@��`S�PH�$�O$�d6��ɇ*0�6�x���ť�I҈�cb��5Zy�����}�ȑd�Ⱥ&�2'HN�{y�OR�X�L�"-����3{�n�+������'3b�'5�ɯ�M�%�ѽ�?����?`�)�^=�H ����C���'�t��?����3�b�dFԅ����͆A"l|�'& �R�DT�'�D��dT��ب`�'Zp��$V�R޺ �M�������'^��'���'E�>u�IA0� ��됉H��,wF���	��M3�$Q��?���4���4�^�0�� �J��'+Q&`��Ѻ�4O����O��U�W	f7-+?Q�	� m�������VgZ�i �3'�&+;��$��'+��'���'���'���2�	�W\ �t[5��8��^��شC�J�)��?�����<)������)-,��Q���h�	����{�)�0T�$���Ц8V8�Yţ�	f��(%��:����	� ��O�9�L>�(Oݘ��Q�C�A�2��:��S �?���?q��?�'������F ៜ��N,��UJ����L9���c����4��'m���?q���?��dS�dRPP
��ؚ6rP��nH
�t<��4��$ʻ	a8��'��O���.w����@V�-��jT�݃�y��'^��'F��'�����A>�$Vڄ#Of�3Iΰs�����O��dM��i`��TyyB�b���O�,��+	=2���ڤ�7�\����*���O��4�Խ�IӀ�(�F���j�)(w
@�6��t�4���hڕu���������4�@���OB��� &�a�&�?�x��CK�]F`�D�O�˓���*И���'B2U>ys4���y8~\�&E8kxmU�&?�]����_�S�T���mt��62\`U ��X;�,���h]�`w�xsGQ���t���]W�}��x�#�"!ʽ���+u#�|��ޟ���ӟ��)�SDy#x��	��G?5��]�A�A��<�Ԍ�?t��O*�oR�� ��	���9PD S�4��!�,r|��f�����O�LdoM~"�2$<T�����6����烋;��hC�ܒ[��<��?����?)���?�-�(�	 #�2\�����"DV�qX��X֦�@�m@������@&?�����M�;Bn4�p��S~ ����#�2] ���?)M>�|�c�
�M�'a4m�n}��q� �P��aX�'����F�\?iO>I+O����OL5�T'\>�h<@$�I(= �j*�O��d�O��$�<it�iCp��v�'W��'�*tţ�(ӠԲ��W0_ڠq��d�Z}��'3�On�0$A�C�ђR���qb}�Ò� �E��=H�v��� 8"ǔ�d �'+/��C���A��b��ʟh���������|E���'����cڂ&����\�	Ӕ�'j�7��5uBH���O��m�X�Ӽ�6���YBn��GF�,|����m��<���?��3���4�����Cč��~�C���Y��=��H��4����݊�䓶��O�d�O��D�O6�d�>l�A����/0��ꃋ|&l˓V���U�'�����'��<j"-������οw��`䩯>9��?�M>�|J֧�c�P���UJ�DC�I��+ ��'��D�&p���)���Oʓ�`��!�Y�z�`�m�"]��4���?q���?1��|�(O|�o��WM��I@d|9��Fr��i��-�����5�Mc�2,�>	���?�;Zup9�|�� ���"h}���X��6m.?1�CL<Pw~�I]���ڿ��bV���02���)9t�r�Ӳ�y"�'6��'�"�''2�IӗA���f_>J���qBȝ�>˓�?�A�i�j��OF���b�O���d$��@(�u�1�ɯ=��E:���O�4�ʱ�0������L��͈�c��X �e��,\H�P�� �t�0��OΓOt��?���?��"~��4�,[.��Юdj�e����?-O6Am.S\p|�'�\>��AȞb5萤���8,�h��??qQY����H�S��c��r�\���,�;��m��Γ/v=Ʊ(�c�=W��U��[�擌���}�I$��q�j�6�yz��]�=��	ϟp�'5���\�#޴8u��3��M6��A�_�(�	����?��Hw�v��\}�'FFA(�m�C|РOU�jh<)c�'�rĀ!rٛ���L�@�М4,�t�~� bQ�P:no~M)����b����5O��?���?Y��?a����=����`�<;m6�+�델N\^$m�I���I矌��^���)�����JU��v�HW�:�B�r�Oň�?y����S�'l�Ta"ٴ�y��/fpaPlR�-���d�&��	r,���'�]'�(�����'�"m3 nƂJ���KG95��,�B�'���'��X��KشiEк���?��`u6�aJG8/I���c�� n�0a�R%�>���?�J>IG��)��5E�C!,�C&Cl~�k�$^
p��4�i;B��4��'��@W1Y+�}��ŝ0Q��V�q�d��Iڟ��������R�O
�E\3i0e+J��R$LT��$;RbDt�p�rB
�<YR�iJ�O�nM-~HPd@�Z�	���b@�S��O��d�O�u�R�hӄ�Ӻ�Bѓ�����0u&��;Vb� F�p9!�0~��O�ʓ�?!���?)���?���i.M��8e�<�xToә^�P�+O2�nڂ!�����؟$��p��؟| tk7���ѱ�I�f���H��ӂ��$�O��b>���)%��	�u��>9A������^)R�k�ryRSpiJ��	�!��'j�ɫ;Ӫ} �˸+�||`�o�-�f���ӟ�����i>!�'Yl7��_2Z�$�)D��bհ�L%��&��$要�?�wZ��Iݟ4��7�حb�(Gw.t�-�H3�B��Y���'L �q���?�}Z��7�
<����e7H\�T�_�d��Γ�?1��?����?����O�9RG��?u׆�����7`��'���'��6��=����O�mZs�	�&%,�*��V�1�������=H�H�'�t����S=u6�	o^~��IK=�`�A9w�]�gF��J�D -��������O��$�Ot��!H��xم�L[Ĩ�Q�I�+sv�$�OTʓ0b�6��s]��'YRS>i�b�%&et��c�K6�N�{�&,?��W�8���X&��=AA8�E_oӂ��GP1x����u���p7m���4��s�� z�OtY��H݇[�H	;Rl�:q��ݰ���Of��O<���O1��ʓtl��.	��li���Y!�`,�0m��3��'9�Cmӄ㟨h�O���� G��3��� .�z�4%Q˓
:F�0ٴ��dM=hl41�'uHʓ��u���1D���E+q+��<�-O���O�D�O:�$�O`�'!��5���yȀ�j3ccZ�иi��E�T�'���'F��y"�l��.�?"v4`1iZ;t��hҖ��&5��d�O��O1�\[��a�~�I�Sb`B��ق6�N�X�銍�f�I!T��mx�'���%�|�'~�'�Z�[���H4�B@��(���#�'���'�Z��3�4n�,%���?��)�ͳQM�K\�D�㘔w�����/�>����?�N>����
� "1�K,�9$�Aw~bbց>5~��KB�+��O"z��Ƀ+�b���EnD����:?R�P��^�!b�'�r�'B��П�xb���$�^]@�,���]:�Iϟ��۴w�$��)OJ mZn�Ӽ�A)	)$�t�eG[�L�rT����<����?��R�pi�4��䓩4Ո����a$���&Y�4�ȃGV��]�pB?�Ģ<�'�?��?i���?�co�2d�X�g`�Cv��a�*��Ϧ����ԟ��Iڟ�'?��ɔi� �Z$��%�"� R�LY��O �$�O �O1�(��%#.I�~���ȟ�c�$�D�\�n�
��D�<i�$�y��D�����Œ,����ڞyD�@E��8� ���O���Od�4��˓g�f˔�v*��םkj�ii��&Б1M�>u�R�~�~㟄��O��d�<i�G�y)�T	^z>pB*��|m�!޴��d���9�'aP�����#���KD�p�S�/��|��d�O���Or���Of�D-���WN���dI���#ư;����� �	+�M�� ��|����V�|�#D�)���rt����ą�&Jݣ;�'�"���$�:d`�6���ݿ)�V�@�12"�ٓA&�[��r7.��8#��|"^���	П�����a"E�e�3p ��.��hq�G�̟��hy��~���!��OF�D�O�ʧg�u��M�Pk���r-�>7HT�'��ꓞ?y���S��gA	T��t35K�~��	%��
M}�AE��.ɛfG�<�'k�~��d�	�S�p�k�x���x�$&&��Iğ ��џT�)��Byrie������M>��⥌����;T��]X�ʓ;�F��O}��'��bS#B�z�H��^D����'=��_1�&�����cC9q�(u�WCJ;IiZ�8�H�[lB0�p6O�ʓ�?�7g&�?����?A��?�'6�����%�U�����ͅG����i�@�
��'"�'i���O���'�:7=�H�ˁϒ�	�\�Y�e��sC��C��O,��$�4�~���O~D˔�l�\�I�p��%f��U�Q�h��,z�'�@Y���䟬���|�X���џ�30��j�r�a���B��sO������ٟ���my��}�F�J��Ol���O]�����s�(��&�G�a���0�1�	&����O���&��.Ѫ�ɤ�����;���2R�	0u*���ɦ9�|�D$����	�,�6�B��ȇ�pA»W\�4����8��ԟ���B�O^���r�i�`�F��4�s�I*^��e`� ��h�O��d��}�?ͻ!}����jE�`�����-e�n���?	��?�F���M��O뎄-o�`���O�? rhb�JL�L**t�@��I��ub�.�$�O��$�OR���O����Ot��eP���v�̂4N�x��'hw�ʓ1��/+ �Ƽ@T�'J�O��������]M��p3�S
��P�Nb�	�X�Ily�S>m�I⟤86	�p> � t$"]z�;uI(*��<GC!?yw�8[Ub�ć�����D@ E2l�`oV?H�}x��M?KB���OH�D�O��4�tʓD%�	I�ROS5��ٚ���$�ɢU���2�~�d�ܛ�O����<Qń�}{`�2����L`BA� �(+޴��$@9����\��^���$<M���eO�7��A��H_���O��$�O�D�O.��5�ӏ�uxiS�8�x�I�E
j$��	ǟ��I��M�BȄ��ݦ�$���@Ѩ0��D��U�#]F�0'�{�I�d�i>��F�릝�'�&�P�J�+�2�Fo�=|��E�A�4�f��ɼh��'��i>��	՟���	KB\b��ي �v!b��7I���i�M++ONTmZ�ks@4��ٟ�	^�$R�N�؝31n]:K=��o��y��'����?����S�$#ї ������uQ��V��4B3}mӑ4�&�<�'b���	T��d��1+3Ꙡk_ĉhd!�EK����柄��՟��)�@yBD~�Z@cv&�
 �*aZčC��Ĭ��$WfH���O(oZZ���I�P����)f����r.X0�Pe �ş��	�U��n�H~B���n�����$�)V1�9�3���-�z�(��C���<����?1��?����?Y/��ģ$�G^/�%�B��c����h���y�������џ�%?�	�M�;d��S��2?.���(�;SF�A��?�K>�|b���M��'�@�ڵE]'M�FVN�(�T��n�hQ7K�:s��"��<�'�?�$�9�̠��:y"��c����?i��?Y����K�I�w$�syR�'  ;��Z�T{4[V���s|TYJR�Mk}��'��O���'Έ)�a����R�R ����tBW�KD�5:� Id��JA� 	�����A�5 ����F�x��]�·�L�Iџ������G���'�U@�%J�=� ��G�?ydF�"��'�6��^�˓ћ��4��Hcզ΁Yu���N[�D�6�h2O����O�����f)N6�<?�-�G8���T����J%6��Y�b@2fY�JH>I-O�)�Ol���O,���O:V�ĢO�Ԙ�%�W��R��<���i��u���'���'l�O�2"�B���0!��9�,�57L��?Q��� ��W,*dxUnu��x�="(�������. 
��� �'J�'���'_�Ի��Sq4���	�5y��:��'���'�����^���ݴ8���Lg����cR�{���U�����R8�&�$�O}"�'
�'nthX��E�:�
(G'�l��p��M����xr��V��4�I��R�BTG�|���w���0�½�;Of���OT���O~���O��?�gLȬp9�5�`8�|5�2��ʟ��	��Qڴvp>u�O,6m)��H�mdX�[����X�@ ��K�6���O@�D�O�)�.��7m*?��@d�=2t/�	b�IP���\��̨�X��?� F6���<����?����?����.PJ�	[��W*>,ZЌF��?y��������FW����	ܟ�O2yBRo]	ġ#�a�$'�,c�O��'�"�'�ɧ�)�3_�ܸ��I��x5��m!L����e�PDy����S %�RBEo�ɺ%�h�K��%K2Hp�%M�	x��(�����������)��y�+n��z�`Ĩ�$������Ԇm���J� �<	��i��O���'�h54��Ը4��J��̈��2<���'8����i;�ɺ>.q�4��H��b1�E�=<}lA�Ń$��<���?���?y���?	(������E13�Y@6Ƌ�Z9��%�æy�aCty�'���mz���TAؑD�����M$E�& �W��ޟ�I}�)�S�B((n��<��eT��B���=0��M�dI�<�AX!qZ@�$ݤ����4��ر
�������#��{0�8,����O���O�ʓ��N��^�	��$��aD1t�n��	P)X�@QU,�B�`��I���Ik�I�R6.y���7��N���=n�%I��$<2�|",�O
��}�9��,�
���ݜ_�л���?����?Q��h�d��Z8q8h8G��.x����T-���MϦ	���Ny�|���杲K�-St�Wx�:hs�(��pԌ��ҟ��'2�	)c�iV��6'����ON����R�l�x;cd^�W��I�[�^y��'�"�'cB�'wbR�5�eRtϜ0n<t$��O&o�	)�M�G���?a���?�O~�a��$s�B���H3���j0
���\����ٟD'�b>E ��V,�����b̌&˔�jP�1v��RK)?�ՠ�h������F6�x�Ж's�p�3�A��%�'k�'�B���DR�Գ�4�������Re�ac���ENR=���)W�F��T}�'���'�3$i�$V$k���Bo�xqW�	�tܛ曟�����D�������I3v�E�X�q���T8TjJ S3OZ�D�O����O���O�?�E�o<�� ��B�CI
��X�Iɟ���4LpM!,Ox�mO�d�������7	8T-"�̗	�JA'����ϟ擔;��AnH~Zw��� �,��"�PO807ʖ''��T���M"�?Q��:���<����?Y���?�W�=s���Z�O�I!�L+����?�����ĎѦ��C���0��矘�O�l4�T�M�(���T�_CF
�O�M�'#"�'�ɧ��U�S�p��PIH�c��
��^e8��\3�$6�cy�O��1����ah�3c�]:s52�,D14y���?���?q�Ş���Ԧi���)$����f'�jMD�2���5�"��'=�7�(�I
����O`����*T�4AǆtA���
�O���Y�! �6m9?i�
���>�ہ䊾8ZL��#�	�|D�4
a��'���'��'R�'���&^$��7� V�"8�t��(�@L��4)�~����?y����<����yg�.Z�58U)�*sv��������'�ɧ�O_dH��i��D��E3`��w P�!n�j�ָ|�DF�V&2��3h�O*��|���ebl�kW�H�P�*�ڴnV�V�����?���?�/O�l�#l�vE����L��+88��yҍJaB*�@f�ʥ8�t��?dW���Iԟ�$�4 �?B�����O�{�l�X�%9?�� �^����۴��O�����?1�J��dzΩ���|�x`�H��?q���?Y��?	��	�O�KQ��">�ຶ"�#8H�����O��n��"�T(���T��4���yW��0-J 0B��?�`�!	��y��'�r�'�NtQ�i���-ldtJ��OI��9�@ԜJH (��l^��BN�^�	�i>��I̟�������8>Tqa��@�]���#U��;1�<U�	�Y�����j��<�������8�M���<��SC���3�-�(�����! �lq���P��?A��?"ɨ�r.�����O�ܛ��Ha���!K/j�,gR��$�@�B�<��D�@�l�D؊����dݢ{y��Sc��1��:	�����O��$�O��4���uv��D�����G�6B)Z������I��;�I���D�O��$�Ov�0�P9t�:1��iȋn�
s#�,!O�7-/?!`��Z-
�|���`1b$�f�.v��H`�� .A�Γ�?����?q��?����On*ٸ@���4��)}Eb�H'H�<��r����X���$�'��7�=�$�|� � !�l�Qi5�\P��O����O�)���6�<?���Y.KB�Tـ�O�2\yIf�ވn&��4d�O�"K>�,O���O&���O$9����@����j���O��d�<17�i��Y��'��'���3
�ҋ�c3fP���@ Q����IП@�Iq�)jd�K�rx�d8�kI����;&˕�G�4�VO��?���*O�iٽ�?Y�!�D�o̅�� �;6*����9�j�d�O<���OB��i�<I�i(��҆�c~ޅ÷�4��Q�D��(i��M��b�>����3�MY�${�Y�@���R��?�E�M�O�R�.y��	���X�F�`!���G�f��4+U�J��d�<q���?���?���?Q/��Pq��_H^h��o1c���@��ۦ(#.I˟��I�P%?�I4�Mϻ"N��C��e>��3��<&��9(���?yN>�|f�.�M#�'(d:AgL�Tm���+�h6h�#�'v�dJ���П��v�|�W��͟|�!�A:_$|)�^� 7���S�D�	ܟ���Ty"�i��-@��O����O�H��8Q��Pڕ-'l� ��gM1�	�����O*��8�Dݪ:�ZQQu*B2\���f�"��Ʉd�Y
�� $O�b>G�'E�����j�ҥ��U�s�LU�%�8z)�M�I�P�IПt��n�O�e z�@�[���򑯆�B����G�6_+]=�I�Mk��wH�$m��Ks��W�\�z��\��'�2�'��n�~�֑��"��^�'��I��!F.��x�2�)����F�O0��|���?)���?���^�������8O��՛'���Ʊ�/O�Qoڤ~ ����l�	f�'�ƽ��l��SŎ���?��p�p\���$�b>���E��q��0��Fϒc7�ea$�� {3H\mZ3��#9�(ܻ�'M�'剬4b���NJ�>�d�x���5w<|�I�������(�0l�|�'Q*6��/l����y��t�A�D�h�M]/����Ǧ�$��ɓ��D�O��o�^�`RA�n��	hw#ٷ&!����M�'��'��t���ӓ%��I�?q��3I�b��BHz�NZ?���П���������I^�'L�ޥ ���@�-I/'d���?��G��R�@����M3L>���Ít!ڭ����
�:� Č^̓�?�,O���Hp� �KT���
�:��D%�4<A��Sj�b�S����$�O8�$�O��V>w�0G`I:d� %D��x�����O>ʓ���a;���'��W>�Jb�Y�B��9/æ_�t`A�E.?�X�`�	���$��2�p�j���l���iF)�
O� ! ���C*��ݴ}��i>A��O��O�qi%���j@(	�	ן5%�h#��O�$�O��d�O1�˓Wf�v`
8;�����(=Zjyx�b�#�z�P��ݴ��'Vj듣?�"G "�\:��ŗ�j �t,ҋ�?�J����4��D�??��%A����S�x��YR�PEDM*1hR+�4�Iey"�'U"�'���'�bP>����5;<��J�g��u�F,��d�M����?����?K~ΓO���w¤�(ݡ=!�&��he#"�'�R�|��'�.˛�<O� ��#ƂY�O� ��B����2O�9�O��?qA9��<ͧ�?Q4k�,�� ���H���sĄ�?����?�����H�u����Vq�f�d�,%�X򐮊�5���g/� t��O���O�O,� G�\�
q�]K3��l�N~r��:Vf���6.Y�ؘOp���ɀX"����<H0!��K�0��FGB�'.��'���Пxxtk<���QIx%��[ş,a�4Rn&<*���?Q��iC�O�������b�U�sj|�x(�m��D�Oʓ@=�y�4��䇏�����'��8(��95�fXA�Os򰸒�'���<����?���?���?I�F\�$�a��,��g`6<�3/ٓ��d������ߟ�IџD'?�I8d�`չ�K�"59��3�Y=b�p�{�O����O��O1����H:8>	�S���kC���Gj#Z".�c ��dQ#�T�F�b@�g�	Uy�߹AT�	�% '&I$N?BB�'B�'��Or�ɕ�MKN��?aV���}	�B�	<L呀��?)�i��Ob`�'�"�'��hV�0L�I��K��^�3`�\��i���*{��l��ԟ쓟�Θ�B#x,1�H��1�DK�d]P��O����O��D�O���6�ӏs"�(�
\*3N���Q
��`���˟��I(�M�$�^�|b��^a���|Ҩ�� I�O�o�<0�&���'������\�L��V��0�D�KŤVA�1���!�=biP2�Rp?�K>1*O����O��$�O�L�C!2;<0ơ;<���j���O����<Q��i�^���'O��'z�Ӭ�,�i0.��T�0H2CԤ���I��������Z�)��dR�F�l�ڛ&踄B�$�.1LNur%�O�����J��@+ǔ|�旣+����|m����'�F�J��?���?��Ş���Gᦗ\�حP�I3.�y�L�4�8ж)�O���ަ��?��W���+'���Z��'�T,@��.!�ּ������ئ�'�V @���i�/O4��#E�*)��p�A�=��I��0O˓�?Y��?!��?�����	�:�\<+���vc�)�fbӧM�f�m��j#v��	��@�Iy�S��<�����!�Y�~��)Qb	ϫO{��[�Θ)�?����Şz+l9�4�y�$�"	眼PjКQ~$�� ]��yb�I U�������?�J�e�y�
�?E�@8�	%O~%oZ(u�R�'��$̹y@`��vg�,W+2�2�,F�O���'�r�')�'����v�*hD*��g�J<n�]!�O�T��݁a�a�� 6�I_�?�� �O����&j�M/>��!��ا�y��|�.�#�� ��}��+Y�w��u��ء��O|���Ӧ	�?ͻ��!��ɉ0��5Q(C�rb��?	��?�oS��M��OB�R%^����-�9�r�RlF�C�L4�V�
k��'��Id�'�&$J�b�[d(���e���On�lZ<_2���	�����Y��&�����J=E��l�S��41ҵxR�(�I̟�%�b>�jT&;\E�Y�&AZ�Bߤ�V�{�"n���D��rؓ�'��'=�I�x/"�J��,��0�ᥓ*F�����S��):��^ڟܛf�Y"A�	����#\0�a'�}��4��'�꓇?q���?�bѲ{������1B����� -��4��ܻ[ \�`�'>�&��v�n+<�[W�I��0�VS���,�O�4AC��t�"$^V�F`HE��O^�d�OB]lڰ,˪�I��&�|��P�Jn(9��W��QQi��iy�'�R�����5�&���9ԭ�d�rHX��V{ZX�5AV�cV��I��Op�O�ʓ�?A���?A��5r��s@ P!]��a dE�/$�:��?�/O�lڱ��U�	�� ��T�����2� �PF#^I�� ����yB�'�n꓄?Y���S��n��lc8xe�'���mR�6���FG7 ���<�'2{��ID�ɛKq��I��OY�P)����&���	ɟ��IƟ�)�SUy£u�e��Ӿ7F�H@f�O�J%v��`���I4�d�O��m�L�	ܟȩ�OH�ğ�,E"�B$֊���oXf�����ğ�B�X���u��H�6�$�^Ny���J	:h�jj_vU��Խ�y�P�x����	ʟ���ߟ�O����h�$})�T��h��{��f�ڈ����O����O���������]	����#�.
R-�w��	7���	Ο�&�b>}� BTզΓM�FL3b��53pr4
�v�̴͓#f�@�#㡟�&���'�R�'��a!���L�
���Ǒ%{��h��'AR�'c�Z�H�ٴ:�<�3���?���S;�1����s��Ս�>8�XM>���9�	Ɵ��n�I�	v���/F<5��Pa���<fV�xjp�	2�I��Mџ�T�ٍ.�|�"l�g�r Vcv���m�3p�H�ࢅ�73e��dͯU�����E�?:rH��Sw^���h�(<��gΦY�:uD�+v9��L�x/��bߓd� 5����/2P�=Z�JH!7BR@���&�zQ��L�*�ܤ�b��4�R�*�l��mBIO/#j�����,S��1kEI���aDѕX�&��&I+WE��p��'jL�)��ı>Q�D�g�-+��b�G֛L�vlKS$�2{
d2�E�<,�e��	"(hd�S)��(Mf��V��M;�� �v�&U���'��|Zc��;�&�倽y���6F%��J�O�14	-�d�O����O�˓-t� .UK@�|��!���:�8-�s$�`��Iy��'��'t��'!:�sw�I�D^�YX���t��̘�DK3�'���'|�U��	�A����͜��2����Jc��x�%�M�.O��� �d�O��D�� Hb�InF��{p
������Ɛ-���?���?a)O~��'�@|���'G�-#�d\4	y����Y1���0��yӘ�D+���O���و��p��RC�y��b�4@ӂ8�2�w��D�OTʓd��Q?�������`�J�N��ԣ�Q��E�J<���?��"��?AH>��O1]sw���PB ���K=��K�4���.6HPnZ��H�Iٟ��������u�c�H�6(H��j*p�F��³i}��'��0�5��/�	9�~�ÕH$_�Ta�shΛ��7�
�d���mZ���	�<��'��İ<q��d��p�EȔ�� �eL܏N��`��O��?��I�d}b�� ��1�@�� �;�`��4�?���?���H���qy��'���%���p6h��Q���0UIÉ"��O�F(�d�Ov���O����`�^Ji���F01�1�/����I�0~���O���?�N>��[P|��'J�Gj0�x��rPv��'�Ҝh�'��ß��I��'�hp�T)��m"WGǷM->4�M�N]����$�O��OX��O
Q!5/��(��ʥ)̓��%��\���O����O(�$�<٣˃�F���q�HDTD�0M(	u`]�H�v^����`�����I�B@��8��-��.K9a�%����	ž��'i�'��]������I�O�-2�(ʇ0E�<�����`�f�Y�A��W���D�	-%�r��=��I��u(�I�W�	;nF��s����	��0�'�&��$��~B��?a�'].�t��K�<<Y:1��L\�#Ŗx��'�2�A�1�ON��
0ʨӲ/�B	:����-�6-�<	�ذ\�6�'5��'����>�1pY� ���Y�b�I��On�dm�ڟT��f$��?����F��;n 4�W�&.��HSj�
�M���F�4�F�'��'��h>�4�����?.�Z�:WaޓF"�鄃Rܦ��I��`�	d�)��?i���?��Hc&��"���6�)i�V�'hr�'O��9L-�4��d��@j�JA�.6q�4  �TH�ȩpb���%�$�~��'�'8�J�1E�0�*�"ϭ9��)�@� iK7��OfEs_����4�'ɧuWl� ����7:{T�a��I����?�*O���O��d�<�f�J�1��0A�?/=�-���̷EE`�'�xB�'���|RS��"Y��3b�7a�|��Y�CHX6��Ov˓�?I���?�-Oҁ�a��|�m��X�q��c�V,�j���~}B�';R�|R\�����x�EL��2r|s"��V���1�H�����O��d�O�ʓC����������v�$���7(�q��'*��7��O�OF��|2����Y�r��Gf��&�\���oF�>�6-�OD��?Ae�,����O���k�֙E�
��GCҽro�eb�'�T��E�(�Ӻ�g$��4(uj�:�Ȥ�D�x}��'���XV�'�2�'s2�O4�i�Պu����ݐ"!ǟOI������$�<��H�p��ħOt`q4E�:�ƙp���;��o��ͤ��I꟔�I�����Xyʟv`yp�Iް�Ƅ��2�M}i��O1���D��Y������A� �0Rql�mZ�����B��7���|*���~Bφ$98��b���}��x:���M����?v�s���������$94N%����\� "R3.��\۴�?�4�U�?����'|ɧu�dѝ��x2S�S�
�v�"���ē�?�L>q����$�O�!��\�.�$ Q ͷ/��� ��SX���?I���'hr�OP��V��\�
��C�Z�x��������O��$�Oh˓S��ɀ8�B�xSH�(b���A,�q�vX���ߟ$$������'D
�#��0H^�딍��mY��(�L�>Q���?Q����dڡW�b|&>����J�v��h���ٵ",�ZReͩ�M�������4����2�D��,٠�Ӕ����� ��Z��M����$�O�غg�|����?���3b���\�L)��f7%���Q�is�����'�zi����Ep�k��QtТ��ЗA_��d�i��;*ܼ(�ڴe���͟������_k4��)�l-�|a��c���v]�d����M|�J~nZ�O8�D�Q	�r����LB�7M;d2`,o�֟��	П��6���|�A$H�7���ۦ*��:*�5�� Λ��'���'�ɧ�9OF��k�Ҕ���4��l�g�_
l��ɰܴ�?���?��O�<e���ty��'��$A�v<�2���K��m��똆U`�F�'$2�'1�1������O�$�OXء&�ܵ*�d�B�,�7{�"!R̎ڦ���8F֒%�O�ʓ�?�*O�����'%F�&����: 8�y��U�����v���ԟ(�	ğ���Qy2�N�/��l�#?.�B�HP@Y�?%n��'�>I.O��d�<A��?)�(������ϴ�yv�K���b���<i���?A��?A���$T09Ejϧ^�"-*a睼-��[Q.ɵx\�nZfyr�'Z�	柸�������i�lZt�C�� ���	X���;-G0�M#��?A���?.O"g��l���'E� Nhʠ)%&X�s�JI� {pt�׺ix�U� ��������q���A�ܴ~I��x���1R��д�Ͼ[nNoZٟ�	qy�*܀$�b�'�?����"��� �J1�Łf�L@.? ��	ʟ0����$�2�~�'C�iP#u
U�S@U�Bjm!�m9s���^�0��d��Mk���?���b�]���� ��5��ܒ�EC�9- oZ��0�� 扤��9O��>�94�ՈmE�lx�*]����Xb�v� 궍VЦ��	��\���?1�O�˓]�^��� �_Sl�����玔ã�i�`Қ'��'s����l@��taF,�Ȣ �X�OK�-l�����ПX�f�
��d�<����~r��> ��xg�� Wb�exp�!�M���?1�7���S���'v��'w�؁D	�5���aV�`��UY�NjӒ�$�����'��	����'�Zcuݩuh�j�E0`�A&tL��O������H��ӟH�	ן0�'�"�C��]�T�Дh�2v�:�Zwn�4w������O���?����?�C��L lP
Cĝ0*�\��©C�ZU����O^�D;�)L�u��x�'H��pC�_OД}�U &�T�nYy��'��Iٟ���꟔ 1�~��߉s �@*B��.(J�4�F����П��ϟД'�h�"f�~���3֮�k D	� ��|N��q$
���@yr�'QR�'���'��s�d�2G �edD�
�JQ�f��D�ik��'@�	PL~��������O��Iʜ]ھ�!e������ 0�}I�4�'���'�����y2�'��	]Z�"�>m�ū� =�X�1������'l���r�����O<�����X֧u���K����Bi��=��c#��M����?q7#��<����?	��ʸO,��P��ʅ8��)
�L[0��	�ٴT�,Y�&�i���'��O,�꓈���_� 9z!$ԟK�ȒPb­t#�n��\�D�Z��`�'�?A�(	�C#��q��@tL��p^�:j���'�'z�ͣ�(�>q(O6�ĳ���E��0"Lx}�U�̒��i���j�O�q�2O�ԟh��Ο�#�Lp�nP��Ɵ8'�P�9��J��M��w�������O�OkL�V���%��{t�a"��H�ɦ:/^���Sy��'���'O�I%+��%J6����@Kam�
E�q�H\��'�|��'�fհ�2�d�U�W���j��u��y��'��'�4k�y��O���Q0��%!2�*��#vayO<������?��s�����0
��#��H����R�BO?���c[�P�Iܟ�	^y�j��?�,���â����zs�΂M7R��0!���1�Iw�	ʟ4�	;O�d���J�䂄�+I3�pq�MF��Ɛ:�4�?1����$��-&>q�I�?M@�k�9��8�ׄjꎜ��Ȅ���?1���}������JY,��� �l5�X )K9�M�-O��%¦݃��H���R,�'�>�`�g�Q�*���K��14���4�?�� �>������O���D�5+X|Kf(K0���)�4�̘��i���'jB�OK�O�������1It�=:)�5
g3\��n�v�*����~��_�X�	4&�4P��!n��\���-J��ݴ�?9��?�oI5>��OB����Hf.��@64I$�̎����f�ēO��K�K�M������	�����ߐdp��U$S21�ԁ��J��M��Z�`����O@�Ok,�5W5ش Í* g��@�E/u.�	�'A��IGy��']r�'剛Q|b(��nG/ObR�_ -��YQ�����?������?����� �b�'0ttfF?�D�$!�<Y*O ���Ox�D�<����<�M(x|�4#�ǌ�S�X#ń�tg�I؟(��^�	؟,���k羡�I<>�µ�I�O��hr�Q��fۯO�D�O���<i� OkN�O,����*��:L����~Ӽ�D!�$�O���E�%b��)}BFݓ^\�*r�Ƅ��HO��M����?	+O^lk��@�S�<�ӗ��I��'7R�dqs�԰N�N�rI<���?��"�;�?�L>)�O���j
�*4o�i��kN90)�9kش��3kr"�m������O��)X~BG���
Y !��)��l!�Ц�M����?A��O�<�L>ɏ�D-Q�c���▭&N�i���>�MӐu�ah� ��O��D�V%���Ɉcs
  � �+m()0r,E�ap �ش�(8
���䓄�O�r��l,4��&�}�j �� W�P��6m�O��D�O��� 
Y쓘?��'|�!�K3[3��[1��'w���J�}R�H:��'�R�'���C��`ԄQ2V�n��P(r*7M�O*H`�
 M�����ID�i�������u��.,��\�"A�>�g��<�/O,���O��D�<I��?��#�B���1��D]�v��U;����O,�O����OV,�Uh�(Z\E1�����!�L'���$�<����?����D
7�y�'J��b�!�<H	�����)�6A�'P2�Dy��'wh�PD��=������M�i���>���?�/O��̎y��$�O��䉜7�ޕX�aӀ/�:�z�lI V��o��,&����cy"���ēQ�(�kr�X']��2��^��h o��<��Cy���:_|����$��#�M��8���I.f�B` ���G��ӟ����iJv#<q�O��<�q���$�"�[9�%��4��"y�$�l����I�O��IH~
� ��!��']��:V		41�h	V�i%��'��Y���8�ӄq���U�XC84�8�C��&&b���f�~q���LR�������h�y!�ʋ�A���VJ7D���+�%K�'�m�� 9S#�(^�z �AHR�nn����
�)�]$) �L��'$�qۀ�y�!�"J�*��FE��.����t�Ņw�J��f@,x2JO�E�t��������G��:��T9���D�p
 �rh|0��k�,��<�A�J�
X@�� ����uxb'�ן��Iğ��I��u��'�7��H���Q:�p��c癅8�p5��FT�M'�2q�["B��P��8��"�X�h��ǃ:k��` ��bp��Y�K]�\s|�#&�ل��L0%�ց#���f�G!X�R�K>�V��L-*��\֌����3n����I�(G{����W�mQb؏C���壃0B�!�d�h��ue�an}A�#��hr1O���'b�I;L]�	�4�?�Rnb���b�E�Th��AU�� P���?�S���?�������?�O>��O�<�F�%��*;T ¨KV8��c�:����D��*Yh��p�)��f�V��dS�d\�.5��8^���́�n�d1��NȐlD!�`_��6�Ӄ<����!�W+!�����}��� W��Jυ**\��6H�g�ɾ>LH����|�����	 7:�Ċ�_��D�i£-� )sui�i����O|��._)`�� ��eĺiԲ���|R)�t���\�^9�E
�嘝~�����>	�d���H�4�ȷe�9r��iV��z]��NY(W[j0)��KO�S��T�I�F��':��0��A3T����b�H�
f�s
�'w\L�F�O�^q�&)��P`�	Ó-����3b��AJ��ׇ�*}_�h��	˸�M����?���#� ��`/ҏ�?����?��Ӽ�HI95
X2��9+�ƅ�����'�5�ϓd�
 �������\3A(P�"����=�.FHx��8�B�^���#@c��ۂݲ�/�K�߂��)�3�d� �,�R���SZj M�4
'!��[$4q2慈�ܾ�[��O���ɮ�HO>ݣ��5q�L�d.,C�5��Ś�3� ��`h�䟐�����I��u��'�b9�@���.o݈�Q*\?R�`"G��l-�����U��?nR��IQ�~p�j!,�h<�9.�
�9�L��se���3l�=
T$��	\��(�cj�C��}��o�f�B�2F<D��IaS$���XA�60���i9�%��'�FlBib�F�$�O�t����}���-�v؂���f����Ol�3
�O8��`>ѩ�H�Ob�Ol�0�*áW�9�J͒4�,E���'���8�BG 8v)�@�޸S�=��eJ��p<�����|$��aa�ϑ�4�1�ұ6����Ł;D�`�!��3"e0B�Ҳ!�T�Jѯ8��c�4v��E8uf�BSB� �HX&SgЄ�<a��8R�v�'��]>y��)���1qkоR�%D��
R$&� ҟl�I�s/I�	B�S��O@��֩ضh! Er@͆#:��Q�>��T���OJX�Ӂ��7W�L��p��D��ոO��2qa�O�c��?��$��	!�%�RJ߸z�X���=D��"fT&Z��z��\��af�=O�,E�D���	v���K�5f��Q��/_�Mu���'Ab�'���R��,b�'�"��yW�)R\���_b�0����>s�1O�����'2]X0�_�51d�х-���2�9�{�-A���<�c�"d:`�����H݊!��.��'ڂ!1�S�g�8kv
q�U��"B���A����|�NC�	��¹DcK�Fc�a�� �5r��"|�ԁ3f��`�t�9IE��y��K<��u�q�6�?)��?��gG�.�O��~>�R�	V�v�{�LH�#>t%p���'GvxC�I�a�2XYЧ�lD���ۆcb�P"��/�Dy��vZeǜ _��,��Eǯi%���4�O�1�v:v@`���a%P��"O�<[�ᑸG�$�BU
��FB�*���XW؞�;��߮0*0�]�6�j؉�f=D���ůףmG<�0 )�?Oh�Ɋt�%D�d�vI�)��:E��0z|� �?D�p�P�گHղd"3�,j��JDo<D�hK�FZ�96���� �1>��[DJ9D�h�A�[�Lq��GH��K������6D��Y�`�� b�y�Ȁ�	�:�l5D�� �Q���қ�r!�$�	=H�T,��"O���֥� |n~�BS)�.F��"O�ăt-��"�q����Lx0̉�"O���#�3u}�1&�ĕf|~1�e"OdA�@M�2�|�@fkw�Qx�"O@��Q�U$FLbx��	��~j��Y "O�u����Ag�9�v��1[�!�`"O��O$P���Yp�y�b8#�"O�ԘA
�U���;�DF�Yo�	K�"OD�ӡĔJQzy��l�5)rX��"O:���
DN5&1h!k�@� �ڰ"OZ	�%��_8��J�5$��8��"O����k�X |'�˚vwA�"O��#�O;?�*��"gX\�v"Oj� 7��	�h�i6N!;�H(b�"O.HZ�$Byz�m��B�S���(�"OL�ۂ)�+E��ZG䒉X��p� "O�В��	�a���6cNeްm�a"O�1��H77�v�Tg� l��<`G"O��I�nƬ+��ȁ���%��"OF�z�/��DJ��Î6>�Mi�"OJ�1A���C$�	+��f%��`"O�d��B�ZY���\@CT��3"O�̙�A�p�hIG-T5��W"O.�@C0?�����f�1%{�"O��b�L�gY`��D�6q-~x�!"O�lǧ1�� �5�^"N�c"O",���[3���c��4Ɖ&"O�+��@DD����K6n�k"O��{�e�Vb�P�'cB.$�$� "O%�)0!$`C:���+�"O����mܣ?��h��n�r�؅"O�Ԫ�
IP!��9�B2&��A`7"O8]!ᏎO|�g�]� |� �"O*q�*��tpu�D�>���"O��wT5Ob$�A ���ڱh�"O|��DK�< ��S����8�2"OV���aӇ-� �@��T��P��"O�!C3��0u�1+ʎzv��1�"O�0rӃ�o���iR��:���"O�X�7�T�}����aɖ�,|z5xv"O��1� #'T�@���W	W̤4Z7"O�@Ӥ B�,�4�� ʖg�F�#&"O���H�Y�0�{��6�*�&"O���-L'Wɒ�r��$4eL�"O�	(����9��x���T�R���7"O��ZEF�mv�W��rr���C]�<Q ĝ�+f���/̷R�N���_M�<�� �*�B˧1���Ӣf\a�<�5&�:����#�N� ��D�[�<��Α%`�m@t�Ӻ=0�H�@�k�<�0G�g�F���H$�X�"���o�<�&��Q��؋7j��
�Ta�t��q�<Q6cݣ-DB�k�b��o�b\�㈙A�<�QNA�$�0�HG�R"B�ލ��ORC�<A ��p�Jq����ZQ�a2H
T�<	�-	I�)г�LYL�2��z�<�e%ۏz�`D�֯J8rp����A�<Y��\<B��t�|^1&
�u�����q���P��0	�͙DR��*���I"4�&�O�����ͩIf>�����($[0		�"O�8����An���h�o�@Z��d�4Y��b>q1�E�RE���b$Q��X���<D�4C�&K򞡀�.��pF-KBBF3pt(`� �)?Y���l�S W���䧀 �@%֨F2��e悠���*T"OB��� �69 [�k|@�ɦ'�]��qk���?����D�,�B���� � 9A�6���c܆d�P�x�'Q6���k̦$~P�z��O@	'$�x��Ș�/�phw�00�b�$��]n�I����	1�5�	��T��SjT]>ƭ�J<Iu�Ĉl:|�Y7��_�<��l�����Feڷ�Ќȥ�42
�p����M۳�`).��>�Q"E�)�>P���є"CTq��@)]�R���/}L+6\��j��v�Ӻ��Kx"��#��RNT��# /��ē/�9��6� I��)I) (Q�$8O�L�3���@�p�C�� Q��A �`ǜU��K@:"�>�E&�}d��sf�",OD|'�\>r{ȁ1��إj�p���G g�ެ��,�>!Z٠��v~�X9� ��E�6-��
��ĻU����=Ig��Gܸ)�2����� U�D $�L���/F!jil8b���b��O�Y�6�O<9:����C$/��90���,C�ő��_�n�<E�����5e?x�<P�A�$�}��Ш���������=1���?�H�<vir	�A�@�m>�����f����>"�,��#
!$�4!��'ĪX�wO4�&ekF��[a�U_p|!�oёj�( �6�π]���ςcU^P�m��A;�X���}�!E�U&1��t	� }�='����KA��ay�G�a$ȱ� N"��d�U��-�*E�ح"t��:`pO�YA��5�.��ܓJS�dQ�P� �'m
A��X���!GÁ$�$}�Ю@�P�89����\�4�뉪3�p$� e�-a�lڧA��s�*�:�W�I�&�����=��D%����k�:k(f��C�2Xz`$�1!D�������bI�����	Y2Y���IX� ��ɕ%R2e�"�ѽS���B�ĿT�B}1�f� T$y(���A���o�)j<��e��P���8�n%A�xp�V䟾x�qY2 .�䗮X�qX0$F�shvQP��.���CD�e���ɈЕ8�
s@ �#�"�<8z�#<�O_�Q�4�)uf\f�A�C@Uh~B%�k?*�8c��f�p�ƤLh}���­s�Щd�7�Ju�@-�7+�ў���Wd*ĲwfA�[z`(+R�1�~DB2�R;������b��"?��烲CJq�eN[T���c 3W�	x��%;&4��$6v�2�r�]�I��	j�=�Baa��$�%W=�)�1"\�wQ���MƖ�7eU%Q|�!+CΘ&T���I$���׌��3�,��IQ�qQ%�8�&�xFf�-��>���9�b�=6��uQ�7����gҨ'���`��'��i��(Y�>qr��$9���,��|"r`��S+2|��R-��I�c � ����Ytl͊U�Af���{$����A�ƌ��"�aT�#���I������7g;�8�f��jmlD��!M 
�xq����-N����v�ӧ��u�%E����^�Ԕ�f�v $9'�/[Zl���<r�xݺ���>���B�E�6:��!c�i7��}[��	���E��&|h>��Dϑ��3���FR���+��1����wx�����S9n!�(ص�D|j3�X:���I�2|�DԗV#ģ�E@�!ۄ,� ȕG�=M��ژ�M�R�#^��Ma��
9{�a#ALd����et�XɧO�9 f���;��I%ǜ-L�(��j�,Bƌ=�e/�����Ĉ��l��!b0����1�L:,����0���m����7}�iF[�����O|���
�}Lqrc��� �%O0h��QA���30�V`x�x�D�2^aX�˕mڊ+�:���4��51�Nx�@�>�؁ȓaº���'F)j������D���K�+��ȓ9k��S�Hv�t�B��������y��c#D�D.�`���I�On]�W �H����JK�K6ph#"O�\�k��kԪݓ�ZRB]rw"Ot�1����s)�c@��a&8�"O�Xb5@F�<<F�G��'s�܉"OT�r"�6B?N��d@� ҈E��"O�p�Wg�43��P Q�a<I�7"Om�֤�G�p��B �?3I����"O,e�R͖�7$�ΐ	-�<Z�"O�4��a��C��=���"OB�Ȁ�Z-C��x�鍑Y�M�0"O
@�)(Y)�p�䧈<	�U�%"O��@J��1f���:��D�1"OL�P���P��Y��DT��<b"OP�(!_7����C�c�"Ot)�Ө.2�(�����]2�â�>Q���'�O���� Gy}�ǡH2��QQ"O�8qϏyب2�/L'L� u���r�N�z	Ó"�@E���=gr��Ə1y�t�}��� ةSɑ�ɜ1G\9W۲��b���5�!�ğ'm|�(N�A�PX@c� k�x��U:]g�L��
:�!�	.pE�aɑD,D��Ð׉(�l��������!S��*}r�VS?4�&N<���T�&���S�G<@,���k�"d!�U`�;%f4vTa�$j��[�HŁI<�I�,k���>�O�!�p�C���c��$�
�s7
O \����0��k�S�#���c��CC�K3)�|��0�7hX;m�ĸ���;I�YA�9O��Sc&�G��O�;s����$d��X�P�F"O�`�@eE�*v�i� ��+�FDh7�>�DA˿^L��P�x���H=B�xxr��4N�"EPI�%�y2`C�V݈�Z�`�I��E��M&4&�d�D��6<
q��'�Xt QǄ�
�U����@Fh��'$*��&ɊA��i"��ʏ6��iY5��zi��X4�<�O�@%��d*�P��0�b�J��'+h��`�`���#}�
����:���]���%�d�<�w���U���rΜ�r���t�V��;U���3�q�)�S6}�T(�'J�t�T)L� �C�I9]�Q�6(�(��x�'MIAqֵ�5�8}O��6���}&� 4����B�S���|�P@j;�,Z�@��8�5H�"L�.@:5�ׯr!�!����[�qO�N⟱O��!(P
�$٤jS Rpl�V���p<!d��I	Xc�d�rfO �(��+Q^�P�j�� ���F�s�qO�>ei�M�l11C���;(f�>}T)('f0�=�"��ɪ�$�N+3��h1��x�D��RnP��
�N��UB0-�f��p���Id���=yQ��&6�r�<�%zΑ� MR'+�\e�`NQ4l�m���&$�`��h�]�,iH�.�T�(�4ڰ 4��l��uW˓����E���7�$eC�V>�1"O��&��^Q�!!ŕ�#)���"O����I�M> [�DD>0�-C�"OZ�8�GC'L"�����A!l$�h)"O�|a�B�9�<�{��&t��mS�"O�I�b'_�P��uʤN�% ��8�"O$��*��6�B�h��qz�Y�`"OLc��G��,�d��0s�cp"O�L���*�"�H�]~�إ"O����ޤdr���L��eZp���"O�) T՜%���Q�J�*>�z�"O��R#�X6�" �bJL���(�"Ol��j�#ht���)�,��"O�%��'�@@5�3Ȝ_�lJ"Oѫå�;rc����խ#`8\�"OY:�3FjȚ�eRҸ��"O�E��/�M�rL
���֨8s�"O�l!���*	��3P`׊w�<0"O��م`�L��U�0��%`PFd�`"O���Ů�e��v�&,�,�"O����S���2#�x�Y�"O�()Vd�3af��pG��.t��!�"OR$�E��-*�h��@7�Du�q"OHP�Gŀ�U� �d`Ȉu��@0�"O. 3cA�S����N֕'l(���"On����ݻw�,�#!��O[�bc"O�,��V�!�浂�-3,R���"O���vB\$X�&�W6#���	�"Ojm���$(���c�KZ��ui%"O�%��N�!&{V;���?nN<ۃ"O����"��P�p�\3WLe��"O�=���]��tYU��DU<��4"O�İ0`1������NZ- �"O�83U�I�ɍj,�m1�j�7J@C�ɰuA����]/-���`� D	3��B�)� �q����M;�K/3bf��"Oֵj��_�IhB��`CG�?��]�%"O&H���?,���`���m�4�E"Ox)��~x"�S�BY9��=��"O�`���K2a�aX#�;*��A"O�YA��S>(�: ����;����"Oօ�m��$��hEH�&��0""O�-��ˀ3�:��7�><0{PÞT�<i�@[*P���fҾ1���5D�V�	{d��#��.�&0Hv��.�Py"A�882�0�g^�2w��"��
}�<�Ogt&h�qC�-?��:C��|�<����g���P�N�uf9�F/[w�<��F�9��̣7��$wN�aG
N|�<9��ȷ4�⭀�AZI�Tq�N{�<YG���Q@�M���_���	#DV|�<ɑ�M- ��� �I������u�<�a�w�8�;#�&P�����\�<� �F�gW
�sd�ދ=�����N�<���pp�xp�`M�f�@�	ǢI�<qEƉE�b46�j��lqD�D�<�c�
4/ސEx�M�K������v�<i��	\%ĐYթ�2�����Np�<���ߔ�
qy3��\n�h6fOd�<IA 6�1���q����bH[�<��@��Mx�iQ�#�
E�P��y��
�usDC�!��0���%A"�y"ǈ)s|��u	�:Į�S��E6�y���`�+"	<,��I5��yRL�7mޜ�A-�@E&�Q!h��y"�&[7*@cÊ®D:@\��4�y�D�9hp�е#��Q$����y�B�v��a���ٌm� �ٷHB0�yAӊ��a�C�#j�ڈ9�%�y��[,q�RC$�F�h�� �f%ʚ�y2�Ʈ{�>]"Ǖ�Z�REOC��ym�
}�|�� ˕Z�6  ���y�n̦�dqq�@=ZB��2"oĖ�y2�CR��&d�9N��9!��:�y����kޠر�\ I��Y#r!���y�L�,�z�x���39��l
���?�y��H�<�h w��F������y��L�<�nxkÂ�%VR��匐-�y��& ><�A�i�4�C��yjC�.̉x����։�2��yR"�>�pѴ�*rc�;RQ$�y҆[�}ژ�# ;j�n��KG��yb� �J��f�D�U��d�D� ��yr��\m�A�gG���l�y��_�U�ɛ�7=��\÷h٨�y�LЈ@����V*�3�B�Y'O���yX$#�xš�I�#P��aGb��y���]�~\ڥM�qV&�aN^�yB���H��!�fa�A(1.@�y�
,9w�u��@��_�t;��^*�y�	N�$��dZ@z�ߨ
��B�\(�y$�΂ub��2��4B�>P�H�zT��vl����n��B�	�b�!
�̓-7��텵Z!�T�.]�gG�>̪u�@l�iC!��(#STXa��W��"�@��6O!�D�r4i�Ο�5�
<Z3*�-H!�d��7&��H򢀹p�T���#W�0�!���z�n@����ԄH��.$2!�� &���Qh y�v� 4��"O lS�Gl-rphV9�dɷ"Ol����6��Y�Xn�,9��"O(r��c��E-Y�p��\"O�m Rft���yc,����J�"O��S�"J�:��iQ;"�nXHb"O<�Am�7)�`X�玀��U	"O���dO8*L�S�+]'G�:��"O\\i�-Hs ��!�ʙ�o��$"O��S�2r��6�XrU٫0"OVE*�g�T,��
A��K<n�"O��a�홝#d��'A]�]	^q�Q"O�A*�L���i� �'a��Y�"O�	�!ك\F0�����E�4�D"O P��Q��V��"�O�s}v-��>���|IŐSJ�\�sϔE4���$l*���/F�_� �B�nT�,��ȓ65 c6+1��lg�A�z"x��Apl��,�7>�}KT���ޔ�ȓ|� S���{W*TsA�\)]����ȓ\NR�r�P�o�n|g`C�6��хȓ�F|[�o	>���b׬�ln�����^��(�� ���
�a���_"��AV�c�`�i�+������:�6�a�ѩ)�bɸ2,8X+|9�ȓ �P�£#�[�����M����ȓr_\����ǗJƦ����]e�8Їȓls�s���|����n�_��<��Rq ���G�>~ܠlҧ�N�I{ҥ��J�5�5(��2�a��
 lU��8�2}ڴ"�/�Yu‾MZ�H�ȓ#8}���Ʀe3�%��˴3���~aZ��`J�9VluB3"Z�f$-�ȓ9�t���ס%<��F�.���+Op�� �1�FH{��� v��8��A�V�h��e8�lIq��8�r���N3t�����?����a��%�Z��`�pM)ǉ�H�>�K �#U�`ȇ�Z��qp����a# ����);� �ȓCr�k��CT'�j��_�l�T��A'���G�A?�������V9�ȓG�$��u��?b��co	�b�`�ȓ3��8��T(^X��s`�D%'�F)��~6<# ����T�v`vE��J@|�=ci��KG8=?��ȓ6*�Q,�
ў�z�� #�H0��#���zD,���	�<���ȓ+l��W�-5B��w���#�ȓ�|`�DI��lR�!{�Z݆ȓ:W�L�g�
�k�x�Е��9ְE��V�RP>�d `� �S<8���,�$�����ĆP�Ko@���+8U��!�a������52��Ez"�~�Ȇb���V�ār*��{Pn�Q�<�VJ\<X6����P۬����@G�<y���P/�a�d�2bi�t�M�B�<���Ⱥi��@a�@��Y����/�d�<��m�6��"U�0�4ܣrËg�<A������j�I�����LY�<����'O^�" '�4�|�p��l�<ْh\�[K�)�+��e9�E{fb	p�<�E��6n���ǛzW��*	x�<����Pp"F� #�`iV�IM�<�V	5;�����dB�PHJ�<� 4	� �!�d���N	f�Q"Or�ՃF�h���%d��#e
h�6"Ob8i��۝
}���ce�	NJd��1"O��Y�t ��9�dL�6B0��"O���)�ы")�{�@�b�"O*�`��)i)���a�9���(C"O����%�^4�Taݲ����4"O:Q����3fh�"6��6�Z�0�"O� �>����i �;ͺq��"O�(zRk�}Nfx:"H�7&�ȵ"Oz�&""R-�&�:'Dv�4�yb�(s
�p�@P�@F���1�y"	��r���Z3;J)�g�֐�y�dN�tD�u̍;9>:��GJ�.�yr���@�(c6#C�5�2Ǝ̎�y�j���l����B�2W��p�H��y��C�ȄBäJ�S?�r���y��F�#�<�����!�ȑ+f�Y��yRn�2��1d�H�	�D��M�y�N��.�N�k$V���fώ�y��2���[7��9g���D̉��y"�Cb�z��1/�����T���y�L#^C0���L̢&�r���gֿ�y��$�$|c���/�2���y"J���T=�e,|�v%��H����x�%u���q�!��� 候�*X��'|�#$�-fl@��F_(��:�l�Q�8�M�"���A �L�m�,�#�=D�` S`�7?��|�`a��k҅±0}BF-�S�''G�ؠC�^^�PI¯N�a��ȓJ�T8�)L+F�����jW�}+�0��} �f!X�*��t��BO�4x^��ȓd4�E�Rm�1lg8�����L���ȓl��,�G�?0K�s�ʔ�>h��ȓp� �Y%L���
����ȓ7�H!e%h���S�k��.��ȓN��-['c4,�Uk#1vܐ�ȓ.���C+W�RL��#{� ԇȓ^�.T#iV��e�	֗Wx�-��G3"yq#�۔\��`��)J�6�DԇȓZ�V�#Uo�0��� �גi;D��{ӄ�Z{��b�?h�Zp�"O;D��+z� "�~�����b�B�ɜ8
�Ps�T�2��$�M��B�ɀu���W�u$��E�ϮgބB�I=�����(]0�J�**.�C�	#-Ը�W�3l���zGI�?l�rC�0kB�uKm `��R �B�	�mX0�і'��@�#�MҔk�B�ɔ!6�4���n�N$"�%I�B�ɏ$�.����&a�T��"l�YbB�ɯa��Y�'ύm�||k�@ʲJ� C�I�P��Ix����`P�8�/
�9B�Dn�A��7|r���4�Tc�$C�	n��-ƃ�r�9I ��3nM�B�*0����#~�^��5�\�z�B䉾�pw��<�8��]�rO�B��X�!��E�5������ϯP��B�I�B���j��*Z�E�$`��/��B��+2 �P���X������Ug �B䉾a����T/�3�f�b�lG;m�|B�I�	]J@;c�ˣ\t��!�ls B�	�4�4�H����_.V��$���Y�$C䉚Eb��dȄt`�d`���+j�C�)� �Q��
�/��K�,^x2�8`v"O~�YƉA�v��P1�k�~K��"O�����s�:�K7k1HI�S"O��9��WH����Z6���""O��#�Zx��1��p��ɐ�"O̙� �@�6AN�9T�6�A�"OJ`�eQ;XD�ISu�7	��P"O���5��0[����Jަ+�
0KE"OzT`�lX"q �t�Ei��![@"O�q�X�x�r�r0fX�K�4�:r"O8��H�0��Ɩ*q����"O^�����U%�P��:)&�i"O��5���m� ����'^5!t"O�]yf�;�l���%���QR�"O*���|굓��<�,���"O|Y�%�
�t8�%��6�6�"O�q8È�j��1DDգ^�\�8�"O2	�#	�83�(�	��8N�^�a"O��)$�H�,����Y��,y�"O���S� C~�����j��V"OZ���/y��$�_�|-�1Q!"O��c&	(7�9a Tz+���"OE#gDUX�c�ڒD2ź�"O~��ࠔ� Z::�O��5��=+�"O���Qv���OM��u3�"O�s�¨5 <�C �[�21g"O��af1PG�0�0����{"O$Q� B�r�^D�R�0DE3"O�h�k��H��@C�ELd��"O��3���bcj�S"�1���"OnM���� &4a��S��=�"O =��nߏG��p2��:�8�b�"O��˧A�ed��DT�nr�4�G"Oz��d
%̦��#C�h$m"O���PEK�.�(����݌F�0A@"O�-	��$..Ա���̊Y����A"O�d�2�N!RrD�X�gC�,�*���"O��(r��$���E�~�2MG"O8������:"�)��C�4I{nA��"O���u&??���-N�G�
�!�$KO��	����T�,R�C�+�!��&'`	Qs�G:��E	��K�J�!�$�%@}�C��O���F<�!򄞹�����A��ԍ�d�N�=!�
���>�JM4h�2}9eJ�"O*���l�p�t`h�lB<N*i"O�����^ق8[�dQ�L
t4��"O��ɢ��40�b������"O��qq��3r��Ф
ɛӸ%(t"O�%����9B��v��(M΂Q�v"OrQC"
GJen���ä�h�"O����B�D-J�
��_�n���"OncD��/?��a� "5����"O���2kY�_O�<{0��d����"O�9�G�ŕ*��F!6�� �"O.��T��&"|Q��?�~�#�"OP D&Ǎl薕9 f�����"OF��&�٫g\���`��A�֥�"O$4���(`Aj�#II"#����7"O��i �PS�LБ���>1�^0t"O�X)�
Nx$��� [;eߚ=J�"Oʔ���kJ!
�Ϙ8)� �x�"O���(W�~�Hr��Ȇs����"O�X0U�|��K�(��>tc�"O� �HR��kEVI 4��K"d 
&"Ot��CE�!�t�Q��P��2�"O�l���*3܂�:��^�m�Sf"O2�
�h�� �ţ*�D��e"O�AB�����t!dE�-�3�"O�P�⅕��p�S��ױ]���"O�x8'"ĩ^B�(�!V&_�b�S�"O����˰�x�G��1�0I"Ob��p-_�Э�3��?%�rp"O�Ah��� 7���L�"��"O�i�F���P�� ��O
~��C"O��k3�V;K	`X)1�#!Da��"O�U�F[���u(�O�k���C"O¡д�W4��X�A��b9R�"O uh��K	
D�tHoŎu���c2"O�5�4#@2P�:� �A:��X1!"O&L�i'�����&S�e+a"O�͑f���%��\�1i�����0#"O6tI��	_�PZ�X9C��i!"O<����_G2��!H���MI��*D��t�%T���Mڴ^��LYFJ'D�PUA�gи3@)�82�E�o"D����g��l����0��5r5("D��C5��x.M�j݄>��be?D��7�Q'�Y�h�� 
���>D�h+�__�m�V�W�����Q�:D�,x�IS�Q��Ai�V!B���a:D�<i��լ[p��S*
7�����=D��@Q�@�8�P8I���;MH�`a�M(D� QP� 2Y��P��=���s��$D�\@!�,fFV�k�kF>X�� "g-D�|c��Z#/�|��b+G�%/\$���6D�|1�h@�x|]�����2:<l�Y�y2a�7ex^��6��/$	ڀ�B,�y�#C��r�Q���а��y���H�$��@�Ͼh#z�x�Iû�yRH
�0�QǞ\0k�%��y��K�A���d�G�*��%���y�-A������n5T�0�S%�yү1R�\����[�w^��0ccR�y2��=	|� ôx���Wk�yD�J�b��:b��:�� �yr��]�.TA��5TFx���o�*�y�S�\Q��[��AI���Xq�M3�y��Fb^�tI!̟US�|�7�	%�yb�U�U�ΘX���S�ZQ!�I֚�yr
�M�����(Bs�ER��E$�y�L�?�����A*��=�y�E�a
]x����.���B�K��y�HP8
}�E�s��)'llMU#��y� h�Q����i>�l�$P�y2���MF����Ua^ Є��:�y"�թyԪ�iUϓ�a�\:uh_��y"I�:f�b`�"JE���㵇Y�ybfM�M�1����+�.H9�o��y��Fd%n�T㎀9�d��C�߃�yR��+&�UY/f�%��A��yB�J�Z�2�x��[(]�P�R�T�y"�� �,(� �Å^0M����yr`*�u��PS�X��҆�yR�ݩ��$ �D/x-�+f�H��y��Ɖ�z@�m��DZ^PB�IB��y�f4<}��x)�:=�V�S�)=�yrE�6u����T��I�Q�QhҌ�y
� މ8���3l���fЌ~�B�"OZ!c�a��0�r�Ȅ�	�|�x�@�"O�%RuG7-G�*�#sڲQK""O�ԉT�E�
��b薔ň�s�"O��1bHS�Sl��*�'�;#�XD�u"O^���Jl4D-&��'�B`�!��U	�ms��۰,\�ȹ���4\!�L�*�tհ6�ޮm�^t��hÈ.��"j�LI���O6HU����.M�;%�B�IP22(2t��✋p�	R�2��d�O����;F䁘P��4 4�D�UnV4��5�����fX	O9�L��Mޯp�ԅ��7	0䢓�A�b��`K�K
A�ȓ��5IS��OJ8l��n[0s�Hq�ȓ}0�a.òU)��ЄM�����za!�c��"����/�=6o⼄�Y`�!#�%��Hl�3=z:�D{���<��H�0���Vm
3j��	���G�	B�D!q�O�h�})��(�A�?D���F�p�\�2��d�����7D�ԣ7�D�$�HY�4�\�RC���4D��86��pԐPT�Y3v�	z�3D���#	ƑQs6��"�D�Eo�E�a�O4�=E��H9\�p�-
 %H�0��1S��� �"����v��cȔ�\�@�=�	ÓMq��3ah�9L��tɄ�!}7�]� o���M.M����r��.�IpwKêT�nІȓ׺�I/g��4�^%A/��ȓL�� ;eA�Z|�(�`�*OqZU�?�ӓ?ޔ�!dL��F ⤤��%L&=��vQt����ǽFi�D��' ��%��b6���@Z�DW`�������H�����_�S�ʹKr.K;��(��\I�<���8'�Hb%[8O��\F�<�Ԃ�7$U�h�c��1�r�W@@h<A�K�^�:R�Oc��i����y"�_&u} u(�-Q\�$2B�ć�y�a�Pu�h2���<I� �$�����d:�g?	�ƌ�m �[l�*6���T�Qq�<�B�ȰF�p�J�K�&���� 'o�<�f�9Ib���Ć	z���e�P�<)4�C ;�N}�5	��X0a�`��O�'�ў��Fa��,{Di�3㘅���H#`�I�<yc��7F�2�F
Eڌ���H�C�<��49�Z�2�l��m�6ԑ��yyr�'&�OQ>5���6W9�Q�� ^n�����?D��s�
ɛ7n����xxy���7D��bрF2rZ̒��W�L�6D��X���+@����耩3�D�h��0D�|�b�%"��BB*�8>�jW +D��#VE�������$>�f1F�,D�,!���gO9��
X I�n%D�$ MR�r����S-T�$�"'D��2`��S�VE���� ,��07�$D���%ϒ�>���s#-Y�n�`��&�'D�X',�>��M�t�׍pl�(���&D��Si։f2HP�,TuJ<����)D�dqdGN,8�P���!�4� ̘Q�<���9}b�e/ɢ"@L8�ÌL�<�v��o�&H�A���"��t��M�O�<a�Ͻ[]M;h�G��x�A��a�<1S�R%W(�Y��� ���ce,XH�<9%��&N�{#(��L���V\x��槀  �[f�gh�	���Zh�ȣ"O����A�=o��(: f(1����"O�Iq�h���)d�^��ed"O
�;�,/1�`K���T��+w"O-q�F�\
`��fϛm��좇"O�%��$C�V�6�,��g�<��1"O�$��A^�����+�� �-q�"Oj !2Y� �P�A+\  R�q"O洃G�8mV�YZ����~8p�"O�Թ�놁4���R � 8/Πd��"OpI�v��$�H��X<�$(�"OR)c�d�%|����QE\��d�	�"OƱ��Ҭm@�� ��9Q��mٓ"O`3�'S�q���j$@@�l�.E�W"Oؽj!I\�t��E1aO�T�9�"O�@8�nN	t�P��?#(�)�"O�(4lɚS�jMIa(O7,�	6"O�)�&�������D(P�PQ"O�D�a�K���X�͒Y��h'"O�h�a[�M6��6hP-���a"O�\����jV�y�Aa=14��;W"O�)�ē/?�[1!߿M\��e"Ot8��@�l)�(㠎ɯs��B�"O��0�K�-b�JR��=�x��V����#��#͚�,��l��o�,��B�#b
���c틶-�`KV
B�[�ZB�IR�
d1���"-�TY�$C;O�B�&bs�S�mH�(/ؐ�/�
��C��9
��H�N%_��ZUH��wbC䉻(��+i��V�h�i��^��dw�4�TU�U�b�Ǝē`1�I�5//D�P:�-hԀa��M�*��	J/ D� 5$\5:�X���'r�U��#D�����O�P�J�#`�;D���i�!w��IP�{�ڼcrM4D�,:4B�9�\=:��ml���4D�P��Hi�]b�ӣ+[r�PO'D�0	�9�|��ê�]�\����#�O�扠 �Œ��R�%B�����V�C��;�6(H�l�2y:��Kٽq��C��"j��!��K�����՞N0�B�I���4x�-ԟvx،�7�ѯJ��B䉟d����D
�M�<3d+U /�NC�|���( BO0Y`�U#�&`0zB䉈v�a�źn�⑩�� -\B�ɋ>hV�w�YH@���F��c+�B�	�oH�l�!�@^��D"�7`bB䉀 TK#��?Z��I3�I3T�rC�Ɋ���{�'X5h��x���
F�C��.ưU;��5N�܉��F%j��B�3g˲$ʒ-�c�s$)� "O"��q"��eX��ȯEx�]�"O�ݣ��Ƣm%Px���۫WszQ��"O�8�fU�1¦�q��Q<4p�"Od�$�6+��h�EֆTl� �"O�	���� � rue��7� �1*Ot �Қ-�TkM�:���K�'�Pl�Q�V���2�AC����'�25Rԫ]4!mҠ�Q�װG���j
�'0���M�(�8�a�i�2��y��Q 9r��O��z5�'��y�]?5$(A����<Mr���yr�E���a�7��<�n`�F'���y����4W"�(��C3���ö�y
� lDC"<+Z�Q�eҞ4ْQ�P"O(	I�d�'Qj�]!�����]�"O ��M΃.&$D��ɞ�p� q"Oؘj�̕Pl)r�9�1�3"O� 2�� :5��>lc��"O�AЦE�y��(g��vb��+�"Oz)�a\�מ�Q��#+U6�)V"O��� 4�����&r6U*�"O\񰀨{E���b�_�u��!��"Oʥ�DL�Yg�	AU��,Z4� �"O�q:���<&�{# JK�Vy��"O��Q!��=�D餅�'�R$ٴ"O�(㢉�P;� r��D(�"O���A��4~�@�▏��L��"O��3�^���JO*pv܈w"Oȵ W�ˠp�bX��.Z�EN�`�""O����r��A��π
�0(8�"O�5�6Ǔ$"�~��uF�}��0"O�X�7��x�����"�2u�G"OƁ�p�ɉq�@1�l����"O,�@�_������L~P��g"OT��T"RLl0q�iڡ(V~q��"OR���Ԁg��m�bϝ<:���"O���c�5,��0�DL�)"�"O�Ap�0]�"ȁ�N�,F1
ę�"O<��抚Gq�n��#%�"O
�u�Y0+�-SuN:W)�s�"O@� �����"�x�mM�\��p"OFQ���يF���[��x��"O�u8㘤��M
�j��E�BIc�"O��s�.	<V(B��qI��A�l�Q"O6��dEI�0%P􊐟?~8�ӕ"O�i�� Fߺ���h0M`�y�B"O���֋�#>�%S4���dBtX�7"O$���AӀp�*����]�F9ҙ�"O�i���&|��j�g�6����"Ovh�pM�C�.�P��$�)�"OJM�`&��u���{���4�V�r�"O\��Pw���f�5�P�I"O��w&��&�e�կq�^���"O��� &=�,����`�RD"O����_F�����J�ot2U�R"O�]A�]X`�@V�,VrA�R"O$�A�Q�I)y���A��)S"OR�Kg�:��T�QC�i�����"O��c�TΦ�k!"�'�"���"Of��bΥY�V�b��ȟ���["O��F�D�3��y9�&2"��3"OR��B�.�T@�%����X�"O8ݚ�̿9'�x�p�G"����$"O�Y6j�W�l��d�Eq����"O���u*p��Ru'?n2�xP@"O�����.��1�&8=*d���"O��B�خR���eT.�`��`"O.\zWB�"�����T	���"O���� �(���(t�R��9��"O�	P���7	�Bէș63����"O�IكEU�>FhQJ� ȧa�d��"Oh��q�Bk���HP��$AZ0�"O���Jn�X�".��D?�%y�"O��+R�Ls8�@�MS�B<�"O!���4{*llԉvݲ"O�h�"H%�r+��\t��"OhIrr�[�Ψՙ��(Y���E"O�  z�	�?F�>����=���@"Ol%(�(�
o�Ř2cU��bs"Ox�X�*��:�6�BT@ �h�z"Oj�&�� Q��q&�'H�$i�G"O޴�@�Y!'j�9!a^*3��q�"O����E��5�jH���d=`P�GZ�<��#X?N�~L3��g����,�Y�<A�%;J�� �/ڵMמ�k!�A�<�t�+QQHaQ���S�N@�<i4���N8􀫆D_�~�U���U~�<y� B5r�%q��G��ʑ�|�<	�a�I���`�/فRmHC�%�z���䓝��S���L��%�=+���`"Opj`G�T޸)zq� �CLq�c"Or=��g�.qU�xn�49�Má�'�z�ųY�8�;�$]�Y�"���'D��)��)uu��RśSG��)c"'D�@z��OU|�	z��5I���)8D�$�E�7�B\����JM��� D��)UL��c�y���H��|D��O`�=E�$�]<g�Tu�D	�
&Ma#�-�!�$X�e�-�3� ����;U��y2ቍG��2����ލ�V�Y�"��B��)�1�'Wj9�d�=L�lB��<x� I���\q"V�i�B䉹L�عI��E�*��|���5'�C�	 ����,@-A���3��F4�C�I�jW��q���+p�Lr�B<D�����?�`83q��0d��s��ħ`�l���OD�S��yǕ�V�~XS���}h���Q���y2 S�b_���ЇHg�\��pJW��y����hP[�DZ�d����	�ymJ7Bpv8C#KگQ�ڑ9� 3�y���`���P�U�FY6!���y�Ĉ�!���`���[2U"E��y�)��˞��%f)Tk���ۉ�y�[ ug�t��CĨM ��!g-[��y@��y[ʄ��IҜ?�
��	��yRh��JSD���Q�:v��f)���y2J'u�Z�4,J�f�D����hO���d¸ �~�r�E̎	�45k�LH1F!��}���1"m�d�T��$f!�p���W<rx�8w �Q92=�'i�@�S�F"�:��V���0r
�':.�i7Dǖk]V��Z���	�'�����o-6TAɵ. T�<�	�'>��:U��(q�m��X {'HUp���)��F1s�|K�K"��]�֭��y�*�����,f��q��N�O@!���A���:��3/ƀ�xUH/@!�Ă^��0b�f�=3��5ʧ	�6_�!�"\N<�ğ�����Ϊ�!�D*h�ne��-ߞL4�q[��-D!򤚱�`}�)��#�4���˓2�!���x"��lM~��!jA&W&w!��F�8\[W��	j��=�U��1�!�䁳%h��ؓFT�`��e� C��|V�y"ቪi'�E�4� �!�����B�	�gN0��B��U��<��a���C�i�	�u�V7h���o
a�QY�'���8t@�Bu6(��բo,���'�B|��L�M�̹y�I�����' ����%sF���
�(�`b�'��jª\�2O,� S�y�b<Y��� <��e��M ر�Sf�F"OT�ф�*<F��X�M
	�ĩ�"O�e��!x'�!;�,ӻaF�ZR"O��j�bbJ�TQ�˔uG�L �"O.��U��'$���(�>ȼeJ'�	U>e�c^2>y��ط/�/�ny�� D��A�k^(%�ֵ�f�%R��xt�*D��$ f�����fל6�����"6D��q��%�T�f��:bu�U�dM3D��	�,��ȣc�5N��E�/D�((�,�3g�!��/�6'`��iW�+D�����A�����݄P�IX�)D�t�p�P>5�,��TJ@�n쬘�%n9D��jq�ѳf�,a��+��N>���I,D��c�m�*!05 bd�}��� 5) D�x�E�;u7*b4m��a�̥��F9D�� Wǖ>�Zh�S-��3
�W�4D�p�ҡ�j���2K�e��]��<D���!�|@��#I�����j6D��30�L,_��M�0���"�z�� b5D��,Ԁ��	Q�}B�(��1D�tT+̛g��i;�
�7�h8Yԅ=D����N��VY1��/e���r`<D�$���ɿ c
�!�X:�j��!�:D��K�Q/u����9B��'5D�4��f��g�=5����i2D��#�kI�F��\�ʋ�A�n�rE�3D��K"�Ǎ'<��0�"�wj�QUl&D����ǎ�(>Y:��T�:1x�%D�p;ĢM�'� ���Ɵ���C�B#D�l0�F�(�,���Q/��""�&D���D{O�O�,�,��赪	�'.������/=+���E�-$���	�'Ö�JS�F�S9tY����8$X��'xfq�,��.$Rש?|��l��'T^ �g�;lcR�bF�%_T��'�҉��;�"�v�Z�!�L��'ɬ��b΍,�D�s��6
�p�8�'= ��wE�D�\�����}�d������,�ZI�'��H���p��k�!�䉎pB�Lyg�6T~h!��(J�n�!�G�*�
s��Xcd�hC�m�!���.P ���@�<1�PQ�HI	`F!�d��O�FT�\�w�8��'>B!���J(uzg��c���2A���#!�$[%[��A�t\�8U����!��,ZD����M�sz�(�I�_�!�[���q��U��D#U�ƣCl!���-)�*� . "�rű`��a!�$�S4lҁ�J���9�+��N�!��t P�*G�z�2c�D�W�!򄕝<�V�iu J�
�&yb��t!��L;i*�I�4O�8x�{எ�eu!�dL4j����N�H�K�5�!�A ����Ú2�
Da�I!Q�!�$D{T�۱�?V�hI���ȬA!�$ֈ9�J�󄭄<(p�ͳ�Y�8!�Ĕ�Z�
L�Fo�)cY�w31C!�IQKRh��D=H�(���&S0!�DP�X���sI�C��p���"r!�d	�;�(v
�\�F���(��A�!�D��]BTI��^&&z�#��F!p!�Q1U)��{R���,�	H2h�5n!���"R5��W�
� ȸ�� ^N!�� �TX �F�cb h�3i:-��4a'"OjA!f�8K�rq���IW�~��"O҉s`����\x H/'Ҕ�(�"O�|�ř7��B�z|�"O�1;�J����g�4�x�y�"O	��̍ ���{mH���"O<�xc �c�p�X�Jݢwp���"O��4�M4�pE;4�B!6���B%"O^��k_ XU��(��S��"O��tV#xT��ˣȕ�f0.���"O��	�b��[�����s� ���"O*�A�b�6�̍��D�;2r
}-�y���G�01�\�D��9o4�y��$�V�۵�G�U���p�\��yRH��0z(c_?Z*L��'fR�y��E�1`�Lڃ��!�
L���Z)�y�a0D2�E�$�,s��1�
�6��=�yR�2R�~����2��$8�mX9�yR�jI:��d���_�.$�aiΨ��:�O����EM0�`Lq��L
9@8H8D"O����h�0%� J�s/����"ObE+��nG<��W��qL^�"O��IWfZ�LE�%j۱t�� �"O�(
�
Q�ab6!z�K�(C��m���D�O������R"[�a�p������L{�Y��"O�|:�V�8!e�`�$SB�p�'���k�	�ct�Q���"�¬J�';2�	��MM�@$�x��{�<��
3!�p�!��r��cJ�p�<�i�*9�NA9c�E9Μ�'��e�<i��u��0H@�=J�g�c�<)�A�q
���!�Z��F�w�<Q4+[O�2	�D��?}�j@��X�<�Ӏ[�Xl��@�߹`���׉T�<����@jt��fՀ3�贀g�Q�<yT�LsƬx ɽ{pxp(姑b�<��9�x���)I:k��X�m�b�<���@�-C^q
���:�v��_^y��'�h�@�%H�P���j\�D��Q��'U,�a2E�A�Z�蒋��}�U��x�j�hf�$i�C�"%��d1����y�I�";p`1��\�	$d�@���y�l�"�Q"ADސK
=S�NJ��y2,�r�ʨZ�K�q�Ti@��y򁇭`,`�kq S�n���+��Y�y"�\�H����T�y��A1ևM'��>��O�=�RgF ��f�6	�T�"O��Y�ᖕ*+��i�k�=�h1�C"O�*���=�<�W��U����"O�2�"]8� k��^mF���"O�� �'����R�HUSN��"O���)	�j[��@M!����a�'�ў"~�dA�'��a؆�:
�H�$�ѳ��?��'�p�y�%�U����eG4G���C
�'�.`�#	�u�t3u�3*��	�'M��2@�K�&'%z��U$�H�<1��ɸK�ĵ ��̡�J"q!�A�<��N~ڼ��n����y�`*{�<�2㞥Bn\Y���_��Lbcw�<YìX����5ř� "r&Uu�<�P��sE0�! � 8�� �!�DN�@ܶ)�T^0m:�:�	�$%!� �H�����_�����Ǻ.)ў��	7|��3�ȵ���#ω�&C�)� �ɉ��l�Ȥǃ-<�<�0r"O���JG�)�Q`� ^ώ�h���{�O��0k ��͘���f
�Zz�ȳ�'y"@��O�kF)(un��z���'��t�W�[Ø��E��&F�t@
�'3h-`֍�[ {u��)%h��R	�'��m	���+c��eK�-�Q����'�Ip-����4��_V:���'e �0n�
ij�l�Ā�Rk.��'���!m�p��቏
PF�y��'0J�B䚛8����Ŕ����)O����ՠH�kקV�oD���r3!�DEj$��`���]�5�Ȭu�!�$��8�pI貅��M'hQK��H�*�!��	(��ܪ��6`|�:�
�2$�!�
=��)����.;`XÀIY�q(!�$QuF�)���L3.X�U"	�<!�D�8V�q`��US}3�j��*qў����<�F1U��u�\C�?_ZxB��e0�hP��6` ��;d��,L.C�	#Y��0%�LCR�*E��pC C�	w:B��)Ț<��(��$�B�I--��A!č�1Ԝ�4l��k�\��!ړ�?9���$���A���4wF �׽pq脹�'����b� ��EJu�hH.�ʏ�$/�o� P0'���
�n��f�1#��� �ژ0�g*X�vL�K-Wc�E�ȓ~�8�&&d~��DBG;���S�D�:A��5+��}١�ۉ���ȓb�ƥ9f�K� ����)�/c��ED"P���|:e��@P�2��d�t����<y�c�T챡���L�:y��`���hO�'�8��wb�����h�%�a��$a�+���(D��n'�Ն�b��K��  X ��T�p��s4:H&C�' W|�Yw!�Ah�܇ȓ<�\��'ሖ;@����4^�F2�'4��)B]�j��C(^Fm���	^j!�Q!#pܠ#�j6A�&p�#!���T��&��gܓ(1�|�U�M�5�\Yw�[9��m��C�(�d�'}v�A�&�qm�8��)Ĉ�`�֭m���E�LgЅ��B�p�X%��2Ȇm*��U�w�v����z4ˑ ^)d)�3�E����ȓoq�P[���Y�t(z�J
�H��a��k`��-@�\1:T�Ո42�?���0<!ao��r��Ї�R�f�,�����l�<1-� _<�)ۆ�ޖK�싒.�k�<d��^�<|ȵ�L�F�`�� 'Cn�<��_^�В�	�%s��a��f�<�͋��z��+����_l�IP���O������Ӳ?հ�#�!��l!�/O��d�+f`X���A�Z$X(��C,=�ў܇ችE�T����
�x�D�J�8��C�	�!����E��-n�0#�!�kR�C�I�J��Y꓆tMV�r��z�\C䉩1)L����
� (9���?�JC�ɏhW�h+�ɂ�\���P�[�c|
B��;mb��S5([�"�9"�Û�u��F{J?�(�̆u�,1bmst��b�;D�H�@j��oq�{cBƓXˠ)�d
8D�ls��4g��aq �;�l]��i#D��r��Jly gd�W�F�j"/"D��`Ղ�)�Iz�,U�ݩF�;D�� hPS&K��(�zV��=Y�h��"O�!BH=��1׮�\q*�"O �b� � &��J�`U=Z�2"O=!uk�ł��i~���O@�cޘ_��a ����B-�CC0D���h��b@����[��<�JQ4D�D��'�oC�RD�6Wj]��N<D����gG�/��0�3l�5�@���=4�(q���!0b����++�i���\x��Ex��	�G)�ƤԪw 0�`�F���?	�����RA0	
$C�n�d��
�,�?	���E�v)ZS�I�f9s'GH%9��`��'��e.�<3>J��ϟ7�	�ȓ9V8�@[@NZ���Q�xj�܆�D�i�� �w�>\ӆ�M1���ȓR#�5��A&x
4%s1�=g0���?�ӓ&K�.�L��e�?�Pi˔�=|Ob����j�(��(	v|���>D��I2���i�bP����eV���F�O8B��Y�XA��.gL�p�$�>SDC�>yL��׻q�(��ט�6C�ɝSE�̛Ѧ�%�D(�Qĉ)(kDC�I�n��Y�3
ݭw�ܨ�Ì�K��C䉞L�~h�bO
�2�c`J }<��?���)Ο5��l�c��:�~HPU� .��'��	y>�"�
]�����4 \�3����$":D���&��&jњA�1�Y u %-2D�h#s"ܔ,��<ȗ ي*����a<D�@ &♤2E�u�&󐁘2g:D��1�W�L�����L Mv��Ɗ�O���G{�O�1�B�y���P�cN�^����!�2B�OύAx�)F`Q�T�@��1�p�'��O�hp���W��UPC��0B�4D��HSÓ�,7��ĥs.틠C%D��*�)�[�
���(cr0qpg"D�@��iP
h��s�b�`� ��K 4��K�bU(N��HՁͰ�(�xg�|�'�a��o�>w�9�#Ɇ'��}1����<a�����-�j%I�$�
6(�`f�$!�d��9�����c�s3� 8�E�Na!�>O�̙�`o�g8�UFH�(K!�DØ�x`���@/}	�p3�,t�!�d��.�ޭ����'�,�N�>;�!�۫�p@�tˁ�7����ӌB�m{!�P�_���$��-wh�
u��d�'fў�<��%H���(�p[�5���~�<A«Y�d'N�)���$/"lĻQi{�<�"��7UlP��ܜu����y�<�6�0s�������J$a �v�<�� �\�*H�`�˯z_Z�P�t�<���Йd���#��--)8��Pb�q�<9q�^�}��H2�H�
��TpS��d��hO�',Y���f�:B̉R1�{�M�'�B��SA�Ta ��W:/�D���*�
C�	9-�U��	}�L�"�,�`C䉹x74X
���K���EHϦ5S�B�I�!�Ft:�'�q��H`V��-���#j�Fp�f�8�ea��6fP���#�dх�о>[���r�4%�b��ȓ�ƀ#q/Q�䡨$�,6,��?9���~:���"ސ\3�dךR��`�T�h�<�e`�a�^5��K��&��)�SO�z�<A�K��O�jw�/e��ɂ�@|�<1�<A���k�ό�E20�e.u�<� �$ �o���.��ïX� ���:B"O����b��IX���12{����"O��s@<�a3#�ˈ;�� �"O�X��F��B#du������"O(�{�H�_xl��V�L�S���r6"O���NڠX.�a膀S aQ3"Ol��D�(Z�츓3Q=Y(���"O �6B<�Trࡑ	I�´��"O&���/Z.���A��"���R�'��O8���%��D�T4j�KX/K��}��C��y�o�J4p�l�#L�0�0����y2����؂��={p�[�	���y�& X�*e��ɀ3�p�Ɇ
L�y�.�"N����Wʝ *G� �v�	�yr���S��Ik��� e��&�2��<��䝱�2ܱCm�).в���5)rў���I:!�+'��#Fv����� b0B�I�_hB�`�D/(�@�� 
4C�� L��D��$��8"���>��C��?T�X#��O_~�����Fg�C�	���p�E��Dr�`I�/��C�	d���% Rj�pt��\�rq�B��P$y��-T�Y2(�"kv4C��\�iY�H��w�$r�L�XB�I%i��Ä�լ)�,I��C��RgB�4^Q�	��35���чW!K`NB�ɝ^dZP�J�=�����hT�B�� +r8�D3%a�A*q�C��93��� �������C�~�B�	�h#���@Z�L~lQ���G��B�I���S���1/F	C2K���B�?,nd�yg@�j�<�r���5MA�C��e��԰E&�BTr�h�a~�C�I�-��ug���yB��u��TC�	e��t�A,J��2B� ��B��m<��B��"6�p��X�m.�B�-gqx@�t�9HP��-A�	k�C�	�O>-����-:Op�c�đ6C�I�'�(Uh��[+bh��k���>1OC�I�Sd�*�S�LPbQ���x��B�l�|`��M.r���R,�B�ɇ#qDl���?�
����f��C�	(~w���dB�`@�����)��C���h�#H<9x��%��>`�C�ɝE;��aE��#f�V�H�jΡ�d��T��uʡ�Y�GQ�D!m�-W!�$��D��%�F#<"���ޠL�!���@N�yb'��DHj�Y �Z([�!�d>Q4�)YblɄ��I���!� ?V����\�[���H�JD!�dO�X�HB�Bۄ+���p�-�+-�!���\G���ݧD�x���>0�!���G���K�%��(�*�1A�!�d[V$6�9
��G�t�[�mp!�$ǐ3uJ�S�̒5
㚴��ӢN2!�d׏	��e�T����-����A%!�D�bJ9����\yT�� ��7)"!�d�s�q�&��tb�U�#�0g!���nG.-yF�ڱ3�(�*���|M!�$W ������M��r��Ғ3!�=>-N勁$�x��Ty�o=�!�ͱZY�#�Q8:�0p:ά	!�$�)\�Q*��7O���T�� p�!��G�0����a�ߕd�p�tŵ�!�� ���!��ڪ�Z0�I�3��(�"O���Js���Ĝ)j�t���"O�eT�$B�p)�e#�VBT�!"O~�)� S����aM�f�Z�h�"O��금&��,n��S�ÑK!�)����-W^��9�G�,o�!�Ē�v�N�Z�F��=I����._�!�$"	�t����]�T.L����[$0>!�+N���\�-�,�1�K,�!��+�)S�	2d�Lä�H�Q�!�B�v@�2'�ŦVBa�3��9�!�DB� ��]"���\HN�S���=!�D��r��A�}B��ro\8~Q!�D��xȍ*�LN4N��'O��!�DP!AؐU7�҇\:x�yÃ���!��H3���u��o2��2��ȃG�!��"뎄o��PB* p�	ڞ	��B��	pZx�:���&�$���05R�C�	�m�LY��Z={ۤ�`&!|zC�I�4�02Wo�('hua�
Q���B�	R����Jp�8��OV��B��-b�L�c�x��k��S:B�*c����_M:��ac~�"B�I���	r! e���@ЍV#@��C�ɴUN
x�uG�n9�1�P	V,j��C��5b1�$���ؠ"��� ��.l�B�I�<��MN�X����bC�I���X�E�EW|��W �'x(C�Ia�Z��RB�h�\�QGb� �8C�I/<
6Yz6&��w#@d�T�<O$�C䉓[�ҝ��X\s�����-jy�C䉼q�v���nS	 �Ơ ��	r¦C�ɸW��Lص�B �p�+�/�2)�hC�I�Q��5��MD�&p�S��̌s&XC�	�t��y	�)��q�vd�T�T�mdjB�	6}��I(Z�/h�� �a#;�C䉫q_��A��0%%���s�Do7�B��M�D��$M2HԾa�g�yHXB�	�)2M�WO�}l	S"�~�NB�'rV�	���5RPa��Z@B�I�m�:o�"`�6�;���`KB�Ie|t�K[�-O����H��"��C䉙r<t��R"�1C�-D��I��C�Ic�Ta����r��O�5�C��!�Z�+�q<�jt�٧"6�C�ɱC:���b��6�X`t���C�ɉB��5
Wć7RV]pv�|�q�"O�0� ��X��xe�˱Tp-`�"OȀ�&�I:za�l@�ܣjp���"O�}	��@��4-@�J�Aaʹs�"O�䊷�P�\#.Y"uh��+�lD��"Ov��uOE�u+��g'H-���j�"O�<�Ћ�p��9�抽[Ffi�"O���ď F��7/(=����"O����֙w�f(���N9{��)�e"O����'[&+��mRDĂ
� 0��"O�X�`J"�*�;���&�Y1"OD"�"�76hЉ�G�+�"psQ"O�H3�Žr_(�!7HB1J�Ρ�!"O���#��Q�\���l��3"O
� DƼBWd5�'�1H��Ȓ�"Of�ٷ�G�7�6�^�y�Ç�!����H��<#��d;���A	!�Dۆ";�}+������r���J�!�� z����&g��L��S81��Ӂ"ODI�W�%o�ZW �?i����&"Ormˣ�� ƬX� ԛmX��&"O�-�eÐ&_>:�$bw�X�`"O��S�iĚk:챓�-�"O�eC��2V��VB��U(�H�"O���� Ц/9^Q��1oJ�4cW"OP�Z!a��B���`M_���\�"O���5��y ���(bv\�3�"O<�*�Iߊr*<�z��G�|RXt"�"O� �£�ay��B�G�E�u3R"OByc�Nޒ ��5�pi�`�,4��"O��	�(G�D��h��"l�<��"OpQ@g�A>a] �摣hF5�"O�@��AL�v= �҄D3mT@H�"O.|� ��'7�쒦BOk8���"O�	��J8&��A��)$�HS%"OȀ�4&V0c�)Y` G��p"O��ǂ�9r1a���#C�	�"O��� V$\nn͸���G�\��"OҤ�dU.��a�
�D$Q�"O�l��&�I�}B�%T�x�d8��"OP�N4.�T�v�V2Ըғ"OL�Yt�S�C
�)#�g%)i*"O �uj�:/���)cg�^�$cp"Ol9r�D�"�h��VA@x�f"O�Pڂ��
L��#��l �"O����#�V��x�Pk߈Z�5"�"O�� �:-5�����Whv9p�"O��WJ��J�2�ަ"�F���f�<��ĝ>�P೎O<^*^�i�<YVm�&�b����$��]A�G�d�<!T 6l�h�$Ɏ#C�U���Y�<)A�;,���+ۊw�p,)5�G{�<Y�.7F��y�k��p�+�~�<q�J��1�R�;�Ȏ�b�������p�<�G)��yh ��S�Y+9uJMP�RS�<��)R�53ṡ&2t���B�Q�<y3,UJ�~)
��O�)�����^K�<I���E��U���������bD�<9����"\\�S��#O�=�� E�<�%�-��A�` E�t1s(WH�<ᐈ^*0��Y�lZ@�tyb��@�<�Bܘ8�[0-����-Ik�|�<��+_?/�Le 5h˫iBn�BAq�<aa�
t�z���U�|1�6͗S�<iDEX���AQ�iA"�t�ȖK�<�WK+\���P��������A�<1S/Q%�Ph�.�:L5�!��|�<9���K4X�c�O�V��mX4��y��`����?��t�	1,�=D�8Y N�R(1�d%I�E�8���<D�Tz&�U�JV���;y���&�=D�@!#�B�:~¹Q��0Z���c=D��R�o
�ik��@1�^M?� S��(D��
c+�-��K
M���D(D����BC�K:���gϝ:%�b|:sk%D�i/.J�����&�3�'�W���'r�J̓��ċ/y �b��	}�����`vLhIN2i�n��dC+P⬄ȓ M��*��ף��q�a�=�r���P�[r�Y /��DJ�@���I����V���IJ'L�D��� ��YsZX�����!�$@�p�C�E8B$�afہa��6�id�"~n:� f�A�0�ٹ�/ŕR� �"O�4Z�,H)j�b4{@O�d�ޱP�"Oā�w��?xi�q7 ��xۈm�d"O����k��t��d�=iɦ��`"O�d�GE�Ng.H�'�X�5䤸��"O�h�ͣw�Mq��=F�N�Z3�'z�ͦO:������8����.ň qs"O<�	�BK�.r\�䏽/D!a�"O>���DM�o|8Q� a�[���B�$0|O2��w�]�2`��D�`t"OڜJM�u�X�'ʸҷ"Oܐ;�eץcR }	>Ha �"O�
�j��>�̐ٱʘ������"O�`�!�5@��Չˌ�̹`w"O�)0E,�7-F��!6H�3( t"O �(�(4��HN�\���"O^ABS�\�w�yap
� s�Y��"O�}�f%Wy״�!���:.�Ya"O�m�V$Z��,�7�,&Ѩ�"O�Q����#30��ڢK%Qh��"O^�q�V�p��H&BFh:c"O`��3�P��4��sf��(���"O�RM�"j���;c%вh���{�"O�@�<;�}H!*M6)�VdB�"Oy��Ly:���/�>�68�U*Onԩc흘0[�q� ��3~���'5�p��E�^�6tc�.L�p�x[
�'4�pk�������SY�G� ���<E��@n�Q���K�<-b���*�&)���y�P�*E�M�+���+���#'#h��V�(h�6e�6fX��8���%�2P�'�ў�|�7��@�L�x�5� ����|�<��N�4 �"%�}�����x�<��2�6Lbu�~�n���`Mi�<�&ElN�=���ѣ�\{���I?y��::H軂����
�Q�h�E��	��=�'e����h
]����&ΣE����%?D�Td'��Bِ��$5��U�U�>�Ic��ħ�T<HeNN�E�8��;�.��ȓ��`+C2abʨi��4@*P�G|��!�^�8taS"p��J���rdB�I�:F���B�^st���@����'���\���'SF��4?��u!�� vnV]��4��}�T?��'��(:����DF�v8B��S&[�Eh����p?)�?*^e�� �9o���a%TFX�ܥO�zFfʞ1z� `�ۘk[ڝ�"O0��G(b�f��`!ɸ3HF��v"Ov�� Hݍ.4�J  �j�J�c"OlT�u��dۀ�@_��d��'��IV��hOl�馪�]z�8YM��=����'�1O"���B|P�m�~��@S�d5|O���FZ�2�DB�*����{��	m�O���S�i�,G%C�oZK(1
�'5��p�N��N��܋q�9pF�r�4�����x�"9o�Z�S��D���С��԰?�H�@}�!���l�@B�+%���X�����b����:�`QG�9t�PC�ɝve�傡HQ�I�b)�@-��Q
C�I$[���� AΜ?x�#/ c��j������!Z��H#4b�,*k蠨��yr�
�']���!)�12G�ep����(O���=H��ଛ�0It�+� �`��z����	�j��v �		. ��Ro�>�!���6��5����#(����fN�nca{�]��է� �P9�.�?��`;�
YKǠH`"O��;�`¸�p|�� ߮����&�S�� `����cɎ��"�����()bB�	�~�b�s�+�6ݺ̨�`W3�C�	�K�ބ����&_�옂qI=�^��$�<���W��v�X P� dZ6iCq�'�a���Ϲ�B<#�G %y^�Pi��ԈO��D�4c �d����焻H����@B�>�yBg�'8d�;�Qr�l�������7�S�O{P�q�<_Uh�0V�F�k��1	�'b�8�d�L�BSJ�ҐCCd�r��H>A
�I%��[sko�"�8��D�,��!�ȓ>ot
Aú2�x���',���>�����Ā��(!3��_���<SAEF3�y"'�yJ��j�Sr^@9r�H��y�K�0m�� �U�L����Ղ�y��`��[D��x� �`6�(�yҤ%p��H1f�t �L�y��D�:���v,�-u�gMW��y�혳~�֜i����q[�G3��'��Il�O��1�eH�m+@A��	W�J|8�'
2��G�S�O'��KI�lg24i �XL\���'�$�c�$����;<���+O"��ā<V~,�bǭGY:��VMa�;\OV��'Cع��MZ��M9w%D8�H4y�"O�q�Oo�)����	��a[�O�C�eP�h�p�C���l��uq��n�<!`�ĉEV*T�7�ʇB��Yq`��m~��i$�O֢|J3.�r���{&�މ_t1��T�<�B!Y�v�(�]��e1�'�L��oӺ#<���Cά@C t1���6π����L�<)�1Y���ɉ������ɦ�&�d�	ӓHy*����@��#�3<8�Ɠ.�jر�'V�TQ���#҃z�<�2 �*$�� ��ըG��X��o̪d1��(��2ғ�hO��2rP�c��`� ��\+@B�(@<�\� ��/K�N�ru/�_�B�u�@����:�#S$Y��C�I!44I
�h�78��摠l��C�	�}K4�2�°r&��I�DC�ɬ^����Ʌ2�ĺEd[�R�0]'�Ȅ�I�&���iUK�+Lt�rr�X<6PC�	����N̵4uTKdm[�g<Z��F�,D�x P"��&:� 灘�@���$(+ʓ�y�ٺK�_? ؼ��aP�s ���L~�<�U%�vq�`P��=7��|[�d�{}r�)�'l�tA�a�֙]-��k�/LaU�<�ȓ��T��F�(m��+*�8� �?!�7��ؠNH��@SQd�D�-�Ɠ'�"�� 8Y����g��75B[�'��i9q`�\�6����%Y�F��'��m�:�:!�CJ(_j��
�'��Dӆ��&��ͫ�ؐKڽ�	�'���� �A<=���: �5A�d�Q	�'t0��$N}�$��J#A���� ���A(�`�0�0C � |�� �ȓu$Wɇ2afA�@�C�=�"!�ȓP~������"�Q��]�?�.A��8|L�%Q�d,��D����m�ȓ~�n���]f֑�c�:'�ę��i���H� �<�~��O8f�V8�ȓK5nP�u�S�xN|�f �	#O�X�ȓ�^���� m>Ehq$�uujɇȓr�[�
�71�d�"�*PB���S�? v�;�mі1C��A�oE�Z� �"Of!��"�	r_N$rn�&f�DM(f"Of�0s#�)xH��T
�)66�}��"O�m��&ޛBZ*�Y�(Ys�4	�$"ODm��f�։	�i���)�yR� A*@�Kڤ�HC'���y�cZ�]�!���ˈ	=F���h�=�y2�P�|KL� �X1o��s�!T��y��/>�6 P��R�4%�ِa�%�y��A7�"�*�n~�W�(��H	�'Ab�@��_�l�2���9��h�'?8� V� m�.��6֋:���'`���皶�F+ߣxp|��'0
yx`�H�<)��E:o�@��'��ԘR)O�uX�"�+S2�ȋ�'��i	�����,GB5z�'/��0�LUtz�2�eH�>��'S�l:���9v�<��éb� ��'��$3�J���>��㟆TɖYj�'���`�(��O�\�r F���Y�'���p�L=5R����F�A3��ӓ._R�q�C#��ԁ��v�T\0��̜~�
�J��\�D��u��:���"��h��Ҷ�L��ȓ"^��`!�G�h����&ʭH���ȓp���K;H-�с����s��a��6���k+��3�Ƭ1p	�'��t�ȓ9� 0Z �W/�쌻cg�4}���ȓuR�� �zG�1Yb��/f"�ن�B�t)�dDhDE[�R�D��C>^�S�Gs� 	x�%W�	x��ȓS�^M(`*�;9�<`#�Z�%i<��T!F�2S�ߨ%��k���[紅�ȓ��ɐ(È.�Z1J����P�5�����C��f��y��>*�z��ȓ.\��fם����V�m�h}�ȓW\X�1��5~,���2.����J�֕�A����"���2;�L��w�
Ii�n�E�
�ɑ.Z^V���B��+]>9J�92�)8j���P�r�R)L�M=^Y�B*	�pv��ȓv�P��@iƏW}n0P����L��Y�$�TM� ��KN,8�\�ȓ]��LƇ�B��`��*�3m�T���N�b��ʹY 'K��4H�ȓ~�(̳��(i\�����^�3�6x�ȓ8��I�s�˹J��I�hCռi��cP�=KdB �)F�䐷�Ҥ/�ɇȓL̎� č�g^1�G�	�'q�9�ȓX	�|�!�!�<h��Чk�l��,t��C*W,9`H�Yh��ȓ#�����)�a�R�#8����Og<�SB�W�����^i�t��/�yK�Ē�ٔX��#��#D�h30�\Bzʈ��
O�Y����s!D�����F dc�a���B����L(D�X�Sg4W� 0�/�;g��Jc%D�D��K�<P���@e��'b���a�#D�����ؔ==|�&,�kHTs4�?D�<����<C��r�"1`�[��!D�$5��Y4$(��։w8$�0D�g��'H:��E����)�q�0D�L���5������ƴ�+�.D�Ի��\0����Qo�� 5��:1,+D�X�egNM��,R1#P%\~d�`�m=D�� T-��.�3FT��s�H�ԡ�"O�4�&��K� �Q'cWS���ۢ"O,�1 Pl����BmD
���E"Ox�Z���Yd8@gN��tJ�"Ol-i�B�.
(�>�8U""O����M�5]gą)�D-�Bq@�"O�-��KH�B)(�#�^{<�B"O����*C�l�V�	Y"4�1�"O��·��.l� �yƀ�Ɖz"O.U�7垚fV�� mS
�!e"O���UeQ�N�D��[��
"OpM��F �b�xjqL�?b�>Yc"O��6d�(><����l�p���"O�%�LZ�G��Q��F*N-�6�0D�DkR�ަ9w2����4>���V�*D���㨏 ���z�㜹 F�P�PD?D���+�>M�40�p㖢i�(P��=D�Dh�ͶxӞ��!��k�P�Rh9D��U?X�<�y֣
�>�"�0D��kR�?(��C��T	���q)/D�{�F�Ge��agP�Y�I�ԃ(D�Tʧ��2d�����#Lј��2@)D�s�#[4@�Z!ꑉF�V�2Ŧ'D�� 4 �Is��!���UT���]�!�DɷR� q5���!"�`�|!��\�9�8=⁩�2�ܡ`wlO�Ql!�$�7������A�N��U�-A&-�!��4\�\�sÓ�M���	�,Q	i�!�d��mid�HbJa� K�5�!��W���A��[^�hh8(��w�!���$LPF�d��m�t۴��*#�!�g�Hᓠ��<n���3(�!��LHRt��R
��v��@�j1!�$V1u�(� ��3|�Z����!�Ĕ�mcH��҈�1��Aˣ/M�!��ݣe�2P�Oف%2���O	:)!�D�1�@��L�p�t��"
u!򄁰P�PbsG�M��<
��I�#�!�$٩d�.��)�<��<SC�/T�!�dԇ;:���KU����X=y�!�dG�!�D�
5[���r��,�!�R�<��	�#D�OD`���q!�䂕ed<����մ\B$h�Lњ*,\QV���p?�B-�}C$q�)68n���#BX�L"�D��ms�`Q��j�-Rb��!���X	K?ޔ"��!D�0���10Zv�(�����: >?1Ah1�		4J�<gז�~�*�<X�Q0_������x�<a�n��;���8�	&vQ��Iw	
�4�l9�3h�ȟdr'şv��'?㞘�$�P�Q�&�9��G\��y�d3�O4��d"i��1��\�K���0���J�q��P�����j*�OX���CI(aۚ ��ŧVD�
��	�IJ�l�y&.�rb�������wuX���D��� ��C&�y�h�00�K�N&v塰�����AmX^hr!k��xeP��U�ȴ�h��]�C-4m�r�Q�@<�v���"O��7��A��t���!��0!��~+&�9d�I� h�)�K��g"�'��'��u�&� m�691A���I�|�������{V��wNL�����T���8��\s#��#'$��OS8hx��=��$
�lA*� e��9i%����W�'O��f���WZD��S�� XΠm������a1cU�R��$���Z74�lJ�"O�12�(_�#�H�)B��E�|�0��Opy�Mg_~�KF��q�7ҧm��Y���
	��(t@�~�4���!�*�23'W%=x�RfΚ+{Q��{"�)7tx5H��W�gἑ���}��'������1eM��(�Lu	�"N�47����o�R`2�٘)����@]:AmIj�J��o)���P�	�>ر3��0lO� �����ͦ/��j��.+K�p��I�+��t�p�
(c���2�I�����;P��s���%�x�i��
|�� ��}��k��Tlm���Q�S�͒��'��pC��MN�>� d?Y��F��T�>��Cf��\�90M��y��� ��TrR��N�-Q��16�11p�%&t�%y�ě� QK|�>1��ޯ`3�j��@�GX�`ik�I���(�+��J@�ISF��^�\�ՎڵG_hL���T7c(}y�E�E����"�16��3o��uS!�H�ԈBƌ=3A@�K�e̹��d�G�~��0�/�|�@
'�y��.BFȌY��4�<���Y���W�#`hQ��2!_z�ʍ�ɒ�p��5P!CDyƌ�й=$!�d�:=px��3.&%
�E�i*����#'?A4��%�Z�>�O
�$�� dd=B関<�-�f
OvP"0�0吭X�5�@Q���q[��Q��ً�0?�5 N5�0��H�Ȥ��v8�|�l�A74�
�b�S��ѡu��U���Y!�W`O:V�!�ă�}s�q0d�1@�1ZeE�]_���b�.<D�Kq��l��/s�O���!�ƽwRƱ�@G�/ܸ�
�'����o8K.�H��"�$j,�-L}�H����.,�PJF���g����(�  /R(@����xj���<��LJyh�">����>>�9C����1�i�Z�գ�Á�	�4�_��$@qC�'?l�v��4c8^\q2$�x=�1p4�[D\#���P�<��d�x����W���.׎o����f	5"" �萝Z���x�H�5L� ���, ��h�)�
z���ϒ3���E&3 ��K�H��@�����H�2\��FI%Eƌ����
E��cU� ,�z/(LR��PBD�ؘ/�1�*��DL;�N�U�CD^&	�?t@܄�KT>Z�0�$哓kG�ϸ'����(�t�2����*�,�Y���U�X�m���B�`+�)�0�e�ݴ,��X�FQ��졧fM3`���N�i[z�!��`�36�/O�X�r�Ϫ^1䔀#mS�I��ܗ+ƂԚ����d��j�@	vV�uB���IM�,b>}(s��`"��qn@IN��B%� �r�,sQ�s��ƼS�
6��5��� }���(����@�q�}�rp 􏒴b���j>�G��I t��p A*`>�!p����݁ F)��D���D]�>�,(0�؎��'�-���o�+c�˽|�.�p�\�+�N���c_��TI8�3�$�4���"�] P�19��F����8���PΈ�}4xN|
uA�p�b��'=.X�g-H�B箐7 F	o����
��,?&L��*WsƄ3v��s Πٵ�&Фz-O� #�֥J�tP��d'>fp�"V(p���Zf��n&ax"�˦�F��'$91B��w�ҥ84d@,K��I��
��\j�;��J؟�#7�+o�-��!̬I^:I�2'!�.��!�Ƅ�2�$�&�tG�6kW ��˗R���"O�
Hܣ[L$�io��8E��Y�8��ؾb �4�>E���[69��" _r�N@�'�C��yrK��V�%k�v�RJ�<���'��rT)�ϸ'p~0)ǂ�`�,�+���Y���
��*upI�+f�6u� h�kD�ā���Z�*#�O~��S�п
�\�bc��8��1xe�ɹA�>@B��Kw0�O��uB$%�`6� z$��X�xh�'w��@3��#�:�s���<_���,O���T�P #�pirL��|�V��=�ĸd�^�ܰ�P_�<DNg�۱�Z��N��A�԰@��\5,�P�c�(��g�(o@11a:yy�!���
�E���(mTqƧ3j�A�������D�ey�8��9�T�I��ȍ\R���DE��F]��	#5v5X��$O�\�qPC�T� ��(U�Pq!�$?2���(��֧K������!h�!�+G��d)$
�$)����A�y�!��ʬi(4�xf��*��BU!�䆘��	��K_��T`��`}!��ؽX� [�&ߒpy���G�i!�d@�<�b�*�Jogx�X ��8+o!򤃇�,��#��1�윹�g�?^A!�׻d���tEL�H���ʆ��6!�xD�����w�<C&

�.!�$C�0A��	7e���sIN�'l!�� ��0��I9�H�!����C"O�,�a�ݰ`nr��"�:�l��$"O��6�H2b�мb�N��V�"O@�
2��5�yi�� �G�R��""O�4��AJ$�|�*'�_*A���"O��@�_<P58�1���39��ĸ�"Oޭ�n�f�������	���s�"O�ܳ6�dW�A�1�
�x~)y�"O�r��yb�r�XCr���"Ob�y�m_�B���f-��b�`�T"O��ǯӿ;�7.�4�4��"O��iA쏅e�b�ᶭ�"O���nG�Z���I�F>Gy؄"O��(	��* ��ˎ)���y�"O���)K#5�(���t���Au"O8)�V��Q�lt94���^���s"O ����V�`�`ܰ����9�,�q�"O�T�&�4ZI�a�@٭��a��"OJ��A	�5��D Y8z�ã"O�(1��׉��@���=��a"O���6���l3�URR��k<�(�"O��:�I�!]nHtj5�� BZ�b5"OZ�#���٪�+r�	 #6�CV"O��(�@��ŀɕyԄaG"O��+g��`��9�_<���"O��F�j�z�xD'V#7��ي "O��C�;(Ez�f��
�,)�f"O�|X���A��9�eN����"O-I�Ô�1z��������xPT"O^ �p	+R�yJ1��?�Z���"O���0��	V�@})Х�!�d��E"Od���ư�a�Ä&5b(�"O��I�I
0����&"H0b�����"O4��2l�-��i�cB�'� �e"O
�3���*4���-7�J��"O­h�N]'H1�5��޲��mkc"O.-����khe�Ag��C	1"O:u�� �A���(.2dS%"OJԂ%��zN����B		�(��c"O≐e��:�j��&DY�T'�Ta�"O����NW���D�5>�LQ �"O`�a�/�%n*-�@�u�FA�"Odz3�N�MI7�W91�:�sP"O��p�V`r&e�1b�#R��h3�"On����aᲙ�!�����2�"O6�iQ懞O����/F-���"Oĝ�d+)wP��B�'!���"O��J�͚eR�h�I�5Tv��:�"O<ȸ1���Ran��r�(8@"O�hz � Z�����5<V�2�"O��	w!�b��rp�8���H0"O̍�@ wgD��%'�U91�P"Ob��6�W�`�'Q� %�"O̤�ԦJ4Pa�XIR�_k>\���"O Q9Ǝìs��3�%�`pn�"O�3c��1����m	�F�H�d"O�Q2�m�>Z���QG��o�;�"O���bÑ6<f����K��(��t*O@l���G�wW��5bW�I����'?�(� 	�wD`�;���~�pJ
�'��(Rn@ytpL;u�X�m�FxH
�'�
�i֦���P�)�@t�X���'�(�+s(CJ��x8�b�n�����'��ea��'}�|
%@S�b����� �(�L�j�H$)�
��0�H�X"O"|�CgO1.�}B!������#"OVt���9lj&Q2�bV�$�N��"O$�U�P�"L��da��4���@�"O�p�uM��c{(�Q�� �~< 2"ON�
��������� ��3"O
D���	?h��ײѡ�"O@�U%�l�!��]�_���"Ohl[��\=a�f�(s�	t���ҷ"O� `#�W"Mɶ���J��>̪��@"O����-±�j�cZ�}L� "O~<��Y�-� ��wo[�C<�"O�0�ɓ:y�	藮�CN�"On�@7e"bZ��1	�U�ɰ"O���W�A{�(�fk
Z��sv"O8�����h�6}{)�)):>uX�"Od�#�jN�E���]v��S�"OxT;Q��[��(��A^��x�B"O��hsD̋[�$̨e@G�E��4�v"O�T���'����0-Nm��Y�s"O����%�d�Ԥ��	
&����r"O$y�Ȏ�!\܈ӵ,��.��Y��"O��bu$� 	��V.O���z"O���fg��Hevu�Y�r�a24"O^ 
g�V�Y�H�Ҧ�:[���"O��e��)&L����ƍ�+�4tJr"O��9ѯ�x��1bŖ���ж"O�-��K�q��H�a��g��M�b"O�$œ�?��ؐ�6}�y��"O@�x�a� ����s(ϥw�ą8�"OzM����8�0�cd�Xɪ��"O�9�O���*-y��H��(�ybŞ_�e�ѩ�?T�`�HMS��yK	��^�pd��N���0��Z,�yBhf(<�*&DU�ALxK�ˆ/�y�׾7�x4�t	�<��Q�b-���y�� J���1�Ꝑ+�h��ɻ�y�M��
E�d���P��  D��yB��-t����#o�@��x�A@�ybJ�(�B�r�vj1�'���y2����Y��E)8�L�Gl���y�ĶEY6��j�1/�B�Z���y2��z/Ĕ�!�"!F�8wK ��y�!��<2�X�Lƒ/�T������y�ȏ*0�x�:')J�x�I[��yRC͖tP
�K@FF5H]�p��(\�yR�A�UA�@h$ B-N@t��Ü��y����m����!l�LA��ט�y�lȲK?�0RE@�u0:D�u�ũ�y�m � �ĩ�e�S�mLڄʍ��y�P�SR��;�E׸c��Ysԉ ��y��.ζ��,�	Z�B���9�y����
U�0��	(l� j��M�y��߽(I��b���c�J9��f��y�o^ ��\�U*-e��$w�&�y����uP�ė]�D$:�D�yr*��7#��q�׈X�E	��C��y��I�t(�(��EE���G�y��M�(�8-�$J�a��YsN;�yOL�N|����by�h���Ӫ�y���#Q\����E�Z�^)����)�y��V�����A�P�d�q����y�I$fʅK��9�.()��'�y�(�(A����fc����Z�"H4�y
� �@K��kf��$g�+9�z%+�"O���Ս�,������	;ېa�"O��Y=
�s6���E�����"O��t�V�?s����& &T|^A0�"O�dY��J��z��1�:]�(�"O��R��H?bԖ�˱�X0���t"O�=rv!)�,P7��S�`��"O��.D��tsЦ޾K�`Pb�"OLY�`�]��Q��
{���"O�ĸ`�${E��C�muv���"O�|�Ε�|�����Ē�m��"O��{����"���!x�5�2�'���2ф�a�	s��;���Y;D`�l> }�C�		h6��1�˘)j@Sa���P�OPܠ�b4+9��O��)(���77BxI���&IfαI�"Oh]�cN�*?��Q*�#��sj���A�>��O���"�3��#xHy�#��:s_�	���T���?�E��E�/H��]��X>"�n)�/�Uh��$~�5���,��ڢ�'�΍���$t�$��+J?yN�d+':Oޔ�w�ѴS�@\�0$�4.=�D	S"O��A��X`��A*��j�y#I�h�,�`�.��B�4L<G�T$Nw&�]�AnB9���Q���ybom� ��ըG|���tcPE����V���c5ʑh, �x��0��ĕ/b(�l3��ԤF�JT`�g��(t1OH\p�'%��O���LīfW@H�B鏡k�jBǖ�	{Ҕ:�E�6)��0�O���p<Asj�i�,�cĬ1����1"_�I��@j�K�hO�� ��-gtz����Ӿ"�Ԥ�Z�� b�-z38��X�� ��:rwb#?J�<D\�Va&���)	lAفN��6�0�h���9�剺O-�ܻ��X�}�L�ʅ$��YR�>	�$�!o�h+"��6#@����j�>�Ā[4ߠ91�-7?�I�#`�c>�!�FP/W�ئ��*a��E�H��qa��A�lz(�*6�Y�7����qO�"A�B=( d�f*C+v�� ���<	������9��DJ[�S�QN�c�io�b�=��	�a_�	Ȑ9k�܌d���A�!e����s�,���Ui�Y1I�&i�f}	% �6l\y	u�^���	( �ܨY�
�2���t�S5f����|��_�x��YABM��L�'����ĐZɐ��'2�`���}|,p�߅/DT-B�%��=��	Y�GG��%�+Gl����gо#/��H���\7����j\&?������\w���T�J��DE���;t���z�" �OY�(�*�:g�����?�h���%"P���{�'A���f��g�g�	���qBƫ�o����(_5^����'��`GO�@���B���_�=��IӭO�R�h�)G�Ht�akElF2����'o�z���
>L��A*�_2ǉB6AO�ٹ�S� [f�$�!G���w���E��փ'�(��$(>  J�O,�HgNɑlGL]�ǫ��@����CaU�(�4��Դ��?at��~2�0'	�q�bH
��D�'R�i�#\9'��]&>]���ɅmbN5W�X�%�8�YBc"D��qA�K�;�N��s%פb���A�(�<)�ϗY��M�SF!}��)�hŎ���EѳH~�iA#G!
�!��,�������0��O�	1��H f4*��qO��)��C�
4Z �U�:<�A�'��y�?��LA愛�i��T��M�l��#)JT؟����I	XO\�2�&P����@aa9�& nK�C|r���0�U^"��e<)�f<�"O�ɸ'�/2v�rF��t~m�[��A ʘ�N���ٕ�>E�D
��(D�F�tH��y��Lz�x�Ś�L�`M�'7�z�'? �6!ZLk�ϸ'��<j2�C$+�|��G�DG�	Q�'��,B�i�-K�1ӢdP$�4˅K��$��M���'��`Yg"G&T��mhg�v)Ç&DH8��ؤj��1O�3u�Ĥ;˄t
�G�"�V0"p"O����	��o*xy��c׾��"O0	p(�E��DW�1��G"O�aba�J6�P�����V�}��"O�8�"��K�'_��V2�"O���Θ�6`��U��o<8E3"OHDQ�b �G����&�c� �p�"O� J(4�A�nu����߶6��|�t"O ���&�#b��Sd�MΈT��"O�4�D���@!�,/�4H�"O��!�ڗWq�y��*rĵQ�"O��!�Gh�V�:��<Di;"O�J0���g�d�XDA�Vɶ��"O��+�e� ab4�*J�,]��"O�U�Q�
	V|��j�K��x�4"OR	s�m� $,�D)�
�
yb"O��PDNS�:@����W2ua�LР"O��q5�]7p�,� �ށe�S"OZ�p�)	Qv���P��;S"Oj0у�8�P���\.COba�"O0<b1Nʷ�T�ѐb�I��"O�I�T&�6�@Ţ�3;��D�"Oؠ�@�Q,S�q��2[�p��`"Oj�����	[�b����U�>�C"O��3�ψ�I�D���◡H��仴"O|c&Aā>APHڲ/I�a-DM�"O&tSL�!�ҙ���C1T����S"Oʙ�Di:]*���,y�*)�#"OܘJE!I�DЩ��_���͓�"Or�#4�Z�}|8��*�tT�H$"O
ꖢ��"P���ç�2`����"O.�)��X� ���d���6��y��](&�n@�B�)��\b���&�yB��9,��P���^���KR���y�	�{�b��E/G:@�6��y���{�&a�G�P:xޢ���0=ـ�ܿh��q�l�R������.y,���O��I<Tt���SQ�<ɱ��K�4As�#	�"(��05oM�<�M̃g�Tx�e�ɍK�<	@RE�<���TM�P��V��� dd�B�<a�A�7<�(����L?8Gr�pb�H{�<�퍹����B�=V���&c�<�cI�&.}P�A[�n���Yt�XdyD_D��چ�� ��Z�12�dH��|��H\M���cJ��!�O�Dn:�fʡ�4J��h�AH��[P��'+�M�4������A?E��b@8��	��C��!x���5��b ���� =���Y}
çe�<a�G�?b^��YąQ)�
��A&��V&�+����LIGH&�Xy ��7a���'�w3������|�'1:��6��� ��O�@�3$�)o���ˋ�
8�8�W+D�C��ɗ	r|yǧM�P��Y��Ea־$	�]�%A����,}HԳ�kN�&����4�IP#��1n]���ːY�����O��I�f_�Ȋ�<�}ʶiݦ)r�.@��Q��@�������$�
V'���h�ӧ��<Q�O	w�iz�Bۉ)��I9#�Sj�<�!�X
I9��U9��ؠ.c�<�7oN���0�� a@&�C���]�<��-`��Df	j� �S�+MV�<1F$�CA��9���. uKc/R�<�$$�G� F�̄�<1[�n�P�<Qu#^�t��UP�ɍ�Ŭ �U�Cw�<�`�$
6�j�e�  �
��[s�<�F���Aӄ�QE.�97���s�b]l�<qT	N� `,�yqJF
J~]��D�e�<	��^�^���2�-�!���6Da�<�r�L$�4#�-�b�-��nIg�<��-E�k{�m�m��R7E`�<�"CӴ`������;�٦�R�<�Q�O�9q�R�.3O��S��P�<1��X�Gr�y�B0}�FA��F�t�<� ���kr%�-5�aC�Op�<��b�
]�hH��B^x�ף
W�<�E��*�3������2&T@��S�? Z�cd�Z�PYy��Y�Q��0�"O�@@F�C�?>����Nu��]��"O:�a ��`t��چ�#��pf"O�$��K�Z�p|�&�R��( "O�9٤��n�0P���QV��z�"O
���2MΤ��܀M<�q�$"O�L
�e�
��W��j "G"Ox��7F^�O����fׂo�L! �"OJQ#�.���l-$g�Ĉ�"O�J��Rǆ}2JU��b�"O�|X�G�'|�ɹaˁ1Z[E��"O���l<� ��C��~&�9�"O���g��4��,ճAr��"O�!; )L 4�� �*H�NQ"�"OFBE*K4���sҮ��Y)�%r�"O����
a"TMW:\��\�"O�9U�@">h�7��e�dMR3"O��+r�;	��� �ՅԞtH�"O�Q6��z8�Q�:B�کH�"O��c�G�>'���)۳,�=�"O.�k���k�l5��h�#����@"O�@8`I����EH��w�B�ru"O�9W�ӡ?RL�j�柭px���"O��R��z%�%^�<�C"Oܼ��"�&=����T�H�s"O�(���*��G�j8�eӕ"Of{��-�ܬp"��V4فA"O^��R�;M�z�B�As�^�Y�"O��C�� nN�0��c[�8�P`R"Oh�E��8��Gc�x|�H��"O$-heA:
��i���7~o���"Olc�J8 7x�k��c��p�"O
�@O��ܔj�ΑbTFQ9�"OB �X^E,�j�h�~����d"O�� �̡hR�D��O�Ҥ���"O�̺�)�+42��։��&ʁ,�y�]�PE�$"'k�M't 1
ڭ�y�Ǫt�����II�l(p�c��y�kR�"��A�4Δ�C삥8K�$�yr�,#ܨHG�4�f�yB!�yB� g���"�ӂ.F�`�F���yb��u����f_�y�Rܸ6d��y�A�g�$��f�3q����P�A��y�a6��iÃJ@�drJ{ ȗ;�ybo�t$�Q8���W]��I�k9�y�o�(w�@�� Z�!q��&����y2j�))$�#���8P`"G͛�yb��)�T��rB2w�TR�"�PyRn�*,$h��<z� #��o�<�R#��9�Z�����G�,�2�n�n�<YǠ\q^=�wO 6��,�֤�O�<�ՠ#Fu)u�5d�i5�J�<����FR8�bQm֘��Q�5DD�<e	�7q̉(6L������u�<��N�u渝y�/�#��2#�s�<yA��J�@�Ȣ35V�Z�F�n�<Q'`�!R	�h�S WM���i �i�<�ui]��0��.YZ�¦a�g�<�0R<$>�w>$P����Hd�<��A+<T����t�I!�{�<駮�u�t�r�iPR"�LCw�R�<іHF+��cbaR�IL��t�O�<9� Ձ<������$�Bb�OB�<�$,U�dà��F"��p¡Bh�<� ���@͕o)Ԕ�2��C2�AK "O
|P���[��X���1��C"O� ��腖h�@�X&+�N�H`j�"O� �d-k:��	�d�+P)@13�"Or]�#��LH�4s5���c�8�I"Op ا���	Z��)&C[�P�0I "O��bDA� PV�|+4��3b#�eb"O�ઐ��~DR���dZ��"OB�ۗ�Ӛrp#��"6 2<Ѓ"O6)i�k�'�.+`M��A��E+w"O�P#D��)*��!��28���"O`�35h��A ��惐�I���cd"O*y��L��S�9�������"ON����E�4�tm)�f�/�xB�"O��#�ܭ/�.��Lȳ~����b"O�h��&��.��0xA�\άdI#"OL)���Swֽs�*�3D"�ڳ"Ov��Ģ�O^� � P�G��"O�PST�0A���h��Gz���v"O�Yx�mM +��=)��
.iøɛa"O�D�U��i�Ea�KX h���"O����T�&���C�jK�A͈�X�"O�%��! �1�,�b�IH�<���q�"O܅���ӂ��Y"�'�����"O\aJ���(]��׬��6%�I�"O�؇��iъ�v�ԷM�Ѳ "OHY�aܚT�0��d@�9�va��"O��1�I��,���N�t�$�w"O,g� �1l������;r���s"Oz�b�H�[F�@����y��t�p"Ox�b�˃$��`	�d��KH���"O���q��)B�zSjT>JH `��"O 0*C&�J��i$k-���E"OF]P%�	
_xS�GyXhf"O��9&�֮k&R\"&
]f�,c"O������$ɴY��D��.fFx��"OX,�m^�t>�D��Α<~w�Qr�"O8��3J�S&v ��D+y`6��"O��;b�S�{v.Y�cA#1�V���"O0`�Ҋ �y�Lp�!�N�x���7"O��+&U�#V�1 �Zh���"O��B%��* 1�lXtN�>n��"O\�(ѨQ�0*1��J�ew�U��"O�Y�6&�)Ax@bK8k�p�q"OHѡ���q�h�Dʆ�\[�T�T"Ol<8S̄
���C��7I�I��"O��*��N8%��H��'=E�l�`"O��K�����1�"��0���F"O��O�+Y�}� `39�z�I�"O�x�'%T{(�DOÿLR��"O��0�A0�6@)���sD��["O���0kނ� p�L�E>P,�"OJ8���=j�U#��EvA�iH5"Oȸ���%c��Z`/�--L��"O��a���6	������#'	f�kB"O�\:k��;�v���P�T&��P�"O�Q{��Շ_�.a9%gD��Y�&"O"��w�� &�H��FB.��T�G"O:��M�n ����r���+�"O|�Q4�$vaH��f�%,��"OJ�b`�2~�v�Q���wL\��"O���q���d��1 F�)U�" "O��Iv�D-m�,��oq $��a"O�t�'��pϰu �G;�	j2"O� q���ǽr����V�3�İ�G"Oz-�ˎ=�,�%`ߐ�bq�"O@��1����k�_r�\�T"O�q� �_� �`�Ĥ][$�K�"O�D�%�
-X<[!^|F����"O��3p`@�I$�p����	8:�`"O>���AQ^N,�#�N�m��UAs"O �P �*[���1�N�!F�E��"O��(�˅�6�	�Y���ht"OV )�ZN �%睳w/����"OڬơN�noX�g�
�2��"O����F��@ ۽-\���"O�jѬ٦I�B�"K1o�Qr�"O�Zw&�f9��KD��h���"O�`�֠�M�d����Ĝ�"O
����
/�d"�H̞J�&�J�"Oƕ�V�P��9��`/Z$2s"O�x���ߦ�v`�0��"��"Or�� ��I)zPQ��0upt�"O��Y�Ι�~!�Ȉ�$�q��"O^���A�B��dX��"Op9x�L@�c����"�>\�Y�V"O�y�5�^�d��#�GXԩz�"O�!I�+�B}s�ыxD�$�G"O�@�dO<X�,��źᠥA�"O�D(� S�B��Y��6$���&"OJ�[��1U�+F�r�{�l���yb��)��3��E5;��0�R$�:�yR�K�;���`�N6���8E�Z�y�C�SZ�+�*��^���ځ���y�%E�7و � J��'��i)1H��y��ٿB���1�I�$�:��c�!�y"oA���w���L�C���y���M��t�4�47�n�!C����y�a�6� �%D�3{�D����-�yR� P����C�5�SO��yb�ےh�V}aMTG`b�!� &�y�E�DDS7FM8��@��΍�y2������`A��nY���%��'����³<����"���y62��'�V��oݳ.��(��º �|!�
�'$�2Ə��-�.��p恸�FAh
�'WNEy��+T��e�g���q���	�'5P��R���E�+hB��	�'��Q���!rj��R%ӵ[TʹA	�'TV���EݔX��-�� ҺTÊ�b�'"@
�蓯6�&x��U�Ju�m��'4Թ����*KC,4{gd�K���'T�35MҾB�Z��ϗ�-
~A��'��XKH"[l���!@-\B,�'���Qө��SN��V�R94�:%��'�����J@� c&��`�'���'�,���"��=�������q�<�q�'����Ȇ��-�%��uj���m�$�T�ѽv��=1��]:��M�ȓ�8UIn�PRr��hS2&�,��r��)����.-�٨tgT*	=:Ć�~,����O��P����E�xd��
��   @�?�   �  ]  �    G*  �5  �@  QL  zW  'c  on  !z  G�  V�  <�  ˜  ��   �  h�  ֻ  �  ]�  ��  �  ��  ]�  ��  �  e�  ��  � : { � � �" ) 2 3; uA WI wR �Y �_ =f dj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�OL ��-ѲS`x�F	�P}�$�ר9D�4���rN ��������$?)��?�S�Or�prI�;�؀7��3�H\��'�����U�7��	SP�fY��?!t�'�6U���ۤ;�t	��1�n,(
�'���f�B�|�+'��+X�U��I�$oB�	2I��u*�	V���#�mI&O�C��:�Dbe���A�p���xǶB�� 
2(C ,_�pN��E��$4N��%�S�O�(�ZG��1���p�-�	���'UV����I�';�9pT�8Ǫ\ZM����I-od⼒�@�O�L����A��B�IަّS"�=�-����#���&�-D��K�U�<��њqI��C~$�B&,D���fB�)-y$�Z%�#�r�re 5D���e��t�����Oɰ�3D��IV�!�XM��I�'���!� 3D��:CD�9CF��"O�&7����.D�p3P����h;��vJb�ꂢ7D��"��.�ɥFK�Z�d䂑�3D�����p����Ȕ>W�����'($��1 ���r��zZm�	�'�>ܪ�`1F q`Q-K,wtҔ�'&.M����w܎4��C��uE��[�'����0�[�^��)��Κx��QQ
�'8��@ ���J��E�dqlm��'�\T3��L�9Cf���X3k��	��� �񰇢�����pl̊^�|Y�"O��Rmń>�ܣ����i�421"Ot]
�n�%�Сf`C�'��Yb"O�lY�H
��6�XQ/��%R���%"O<m�$!�6]h5@qm��zHLL�""O"	�tjDZ��*+\�"O�qQ��D+x���O3#�0"Oxq��BUo�Q"rN�&/!H�w"O@q�%��+���#BJ|�v"OL���#N����՗`�L���"O�`$DHA5�Ţ�΀S���1"Oy1V�K�:�Z���M˷BQ`!Ʌ���HO?�F�@Tř ���e��E!f�!��J+slp�{ҁF�,.L��e�͜vg@L8�8O"�p?���
$�Hh��-7���k7�c�<�4��#8SL$3ĭ'H�ē��_y��'�J��M�n�L}I'֣^*�L�K>q�O��?5�O�D���#H�a��hA��P}ڱR�'���	��^��Ҽ�@CU7z�H@3�'����Ȕua6�{�O�?j�n-q�'�VPa�̃�&l��r.N�ZYF`�
�'�p ��2`�����(�����	�'o*r�凔�<%+�$D>�{	�'vt�C��7*�Prt �1B�ѹ	���?K8H�6���m �
@m�O����ȓ)�� E�����h�6J=Y�$�ȓ/ͪ�yE�/;ԙ���6�-��P��6��1�ISSjױG��A��~�4�+C�G�[ r���c�[a�,�ȓ�Q�lP�L]��	V���ȓa�\h���Ͷ.p�A,�RC�0��1�.b#��A��\��Hڊj����gm	a�D0KM���M	@d���-R&����*t��X�ĒlQ@D��oLؽO�Sߖ����pzt �ȓ
9��ײk������-�$Ԇȓ#����KI�=�p豇/&�P���HR!�K�B���qcM$"��@��;�\L��R�*hea$B�)r=NQ��N�J,cH�M}^pzQ��&j����ȓ{���`Q�gpٛ��,t˦Q�ȓ` <�Ĉ8�4�s��*p�-��Z�&uP��G7�ܜ�G`ƿI(Ј��D� 1�㇣��L�D͕9/����ȓtF���CH�MkH��nR7N!p܆ȓCUf�Am�,�r�#QA~��d�5D�@9�ƖY���`@Z+���0(D�x��@U{7llc��C�n,� �q
&D���Ç�5�\Af��Kӌt1g&#D�ĢS���PДI��m ]���� D��Iq�¥y��)���+@��$a,D�,���25 ��Ӊ^)Cl�	��+D����[gE$����dZ��6D����$��F82��P�+��4D���G+�o����+��g��pQ�7D�8�Z7��<B5�A&	x�V�9D�<���J�O'�1�Ği�NȐ@�+D�L���] ~�V1����t	`�C��(D�@S�C2q���S���c�V0��%D���$�E�r̈�i�%O�F�GH/D�0����,s�*Qh�d�1��0Zq�-D�� �}��1�Q�I�+ ֘`"�+D�\ɱi�4r��DJ�'g�l	�m*D�,ĥѣw����!A>�躄�"D�� Hui�`̎L�`@��/�B�jq"O�G��6��BC��NF���0"O���P.1x,$��� Y��#r"O��!e�3�J���l�#6��1%"Oȕفk�:qVD�1L97
�P�'�r�'���'���'lR�' ��'�z3C�&�l��	S�[4����',R�'��'�b�'���'>R�'"�q�SfVL�k3n�-������'Z�'���'���'zR�'�b�'���(��12�"�1D�U�n��Q���'�R�'oB�'��'�"�'�2�'�V���%.5��L�5C�ɒ�'s"�' �'���'y��'���'}p�����"�Pآ�#P��$�G�'��'�b�'�2�'�r�'���'ؠt�Նm^�X�'$P�Z��H�w�'R2�'yR�'3"�'hB�'���'E�����t���EL�.�<�B��'R�'���'�"�'�b�'���'8�t�_����LU�j1`!3�'��'���'i��'���'r�'��%��� !s�\�цD&4ݒ�Y�M+��?���?���?I���?����?Y�e��[����%)�f������?����?I��?����?q��?���?�᠄����Z�$���b��9����ɟX��ܟ�	ퟌ�I���	ҟ��	
_~�����D7����]>:�J��	����I����Iʟ����ڴ�?y�!��ГH��$���]�n@H������D�OZ�S�g~Bd|�fa!�g߫zgB� �� t�.��b��Dx�	9�M����y��'�)0fLG�p�E��0�ҹ��'���[��֙���'{!�4�~Z�g�#-�и�fw��0)6��B̓�?!.O��}�w���Qب �"G�!�q� �;[�vf]���'��(dlzމ
�+��!V%30CF#
,�� t������	�<��O1��m��n���I+17�-��G-sP{�*J������<� �'���D{�O�R��>`/���7�ӑ
Ŗ�ZqF��y�R�'��۴-$�Q�<9Qi�c�B8�t��Z�Pi�)���'7��?���y�X�@���'o[H�(�Kx	2&�E��	ϟ����V�b>�
��'�D��v��8�B�[*6�� ��佔'I�ߟ"~ΓY�Jh1'��2>�8���I�
#� tϓP`�F�J���$Q��?ͧJ�|94  |����EΓ�?���?y�,�:�M�OF��j�E���"(� �Ҳa�~X
q�H�F�O|��|*��?Q��?���`��F�V^������N4.ű/O�1n�:w�m�I��\�	n�s�t�#��O �X'�ʚ!�V�*$,ǩ�������ڴ[����$�O��陇%"�}�bD�wQ�,�>�4��A�X?h��J !ZH1�Ӊ�r���K�	��$�^-zĈк.;yr3 ��*
�d�OH���O��4�˓p���?�B�D;[0̢���;��= ���yb�c����h�O�o��M�u�i{�+gA��+���'Z�s` ɰ @�:fG��:O�@un	$]> �H�����zI����֝=��[B��2u�0�y�&P�<���?���?I���?���Tşpؚ��J����H@��&Q��'�*jӞ�֤�<���i��'��L����vބm���B�A��)ӁO.���O�7=�X��G�q���|p.�
�D�iCT��ȝ�'��V,�K.��Byr�x�0��?i���?���MӀHK�P�U���@`D�m��	+���?�-O:�nZ�v馽���L��w��jH:)
t�R��gNh����_���DAy��'B�� 7��O��$nI WYLaB�!�W��tG�hՖs�`��kM�6E�<����"���'�����Q���9����H�c���ej�ݟ$��ɟ|��ߟb>�'�7��W��m��ӄI �d8҆�ie��9Я�<���i��O�d�'��6͛��6u��N��<4�p�`l�=P��nZ��Må`W�M��O6}��nJ���U�(�����;4,��5��a� ��T��3�M�*O��D�O���O��d�O�˧&�U�F�!&V��� ��#c<tX��i��2�T��	Q�ƟȈ���[P�	1")0�3���m� �2HʬeԛFe��&�b>��V����=�{��2%��2=���%l�$R`ΓP�`,�����'�7m�<a���?�b��5+˄�b�
蜈[U� .�?����?	���F����mE����	ПD����tN
��a&�U�&��	��MD�i,Obq�焳B���u��,���*���d�G�VU��n�������;�
�����-*���P�7��ԫ �,��@������	�����j�O�$� l�ȉ���7&v�	ؔ��5L��z�:���D�<�3�i��O�P�l�*�XAȝ1$D��5	�]^�ͦ�9޴B.���ӛ撟r�oR�0��	!-��������b>^X�@�@�R�,��R���I���I��I�L�'Z?>�l(g�Ё}���$�@Sy�z�N�#��O��$�O��󤕊�
���Ȯo��l��ɲ.��'�t7���5IN<�|��8:�^d�r��O�x I"gI�y7�`ٴ2剓9⤣�O�ʓ%r��^����@��U�D��E � �D���'Wb�'��O��	��M�%�X��?I��L�R C�/!��QE��<q%�iB�O(�'�6�զ�bڴb4~x��G�A&0���؍o��h2'jͬ�MC�'����
M�n�����d���3�{�? H	{v�71f��s`R %Q����8OH�d�On�d�O ���O.�?]���N�@���0�bYD��Dy2�'�6M��~���O�Em@�	!�<I���%�|��B�Fl�J<a���?�'$� �k�4��D��M�[Qc@���{T�K�)32��uj���~�|�^�<��П��	��h5�ڲbP�q	������ϟX��dy*`ӀXs=O(�D�O��'��`BT�7g��2��6���'U���?q����S���_;rɆЛP�B����S0BЍR�o�u/�uq޴��4���8�'��'���(t����� ,.
�����	�?����?����?�|2*O��ͧD���i�&�������	ٷw-^��A����۴��'����?9�EW�u�����a��>��@gC��?�::0+�4��d�/w>}h���l�w[���������Z����y�U����ן���П ������O�$�1
� _djPs����-�1d��͓�;O����O������睍R���SfmԇA@Z�Qs��'�f��IϟP$�b>= �Ŧ=�p̤��f���@	"tBw�CDS��͓nV��0�࢟$&�����$�'���b%��:(�a�CMÕO��A9�'p��'�RZ��x�4x��)��?���"��m��,N���;�i�#~��b,�<I���M{��xRȝ�1�(��g��ECr-��H����$Ϫ:������(�q�DM���o���|��K�e�<�t��UN��i�R�'B��'�R��h��n͎cD�)���N62�L]�S�՟�eӴ #ug�<Ӵi}�O�N�x�h��T)��Y�����D��Φ9ݴkW�v,��~E���L��bψ��T��.#Qz��K=� ��no���&�����$�'�b�'B�'y�|��ٱ�M�P�m����S�\ߴz�h����?������<��W�	u���$鉄�x�J&OԋL*�	�MKĻi��O1�֙h�/����}�� Ɨ$�$łRKM�e �|����X�ŮV�R�s�	]y�e͘b
�`�oՍpE��ɁL�N��'�"�'*�O�	��M�����?Y�FZ�I%>��Q���*�D<g#O�<)u�i2�O˱>�#�i�h6��ۦ�[��� �<��v�V"���cEj�<��m�x~������kܧ��cA�&"r��s��x��י=��ϓ�?i��?���?1���O�0��T��U1�@�UK�	}���)��'���'��6mSm��)�O�m�|�H��׍� �D!P�n^��A�L<A��?�'}�8��4��B$*If�:S�L�'�TЁ4"��&q�mH#��+�~2�|�R����͟��	ǟT�↖���� ��Y��P�� ������[y"ei���V;O��$�O"ʧ��K�.�:���E�3��d�'O���?����S��fO�f)
�y�@1rė)Rhv)�
�:{�搟擣P�D8���1&�cE�6.e�d��]����O��$�O���<�E�ib���`�5�ڹ�H¨n?��T@��/�M��BH�>)��i�x��v���w�"Э�;�%���wӆUm
�ll�b~r���w�4��[�I��;Rl�3�B��H����k�<�
��H�Q"�<z�J)���L�q�< S�i"����'��'!�Qoz������I����v��Y`���`�	��S�' �J�+ش�y2���B��Wd�=����#���y�)T�~_0�������D�O� 08_�h˖/��\�$�s�H���O���O�ʓ�V��L��	ʟҤ)ߦY���Hҳa����E�c�e���֟��I3�ēEp�
2JH�`6-Z0L�&_���'�|[�*�V+��m8�I��~��'p2�)�G��ΆXX�1��'���'e2�'>�>y��1"��a'��2H%������"e!(���M[�Q��զ��?ͻ`1xI2��9>���t �����?��J�֭ƞi��斟X2P�K�	�	rܬĳ�	^.r��X"$�)�r�O���?)���lZƟ�����H��O�9]��r͖+jn�)��ly2�{�,�f��Ob�D�O~���$Ӵ[�^(V�1C��	�Cف,F�'��'�O1����%���G�Q���7'�֍�!�Ah6m�sy�n��������]�V�QKD�^�T
���݊|�$�O����O��4�D˓H��Ƃ( �2��3O:���7
!Nr:��6&	�y j�T��8�O��d�O��m�e�8Q�'ۭ �*�H�
w�49��Y����'(4�HSYb�O~z��[��`��[<R�U�gAt]��Γ�?����?���?�����ON����܆(d��7�4Х�'��'�7mBR��	�O�Em��H�'��)����Bg��rJ�q�6yAe�9���OX�D��h�zĬa�H�	�|b��V�#�,0&D�5@�H%�'��=@ f\�a�O<�O(˓�?���?	��.�
$��*K-V�%:��I0^�����?1)O�Uo�=x���Iȟ��	l�ĤOj�:�#�-o�X$�F�ܬ���X}B�'�ҏ#�?�In�^]��J���9X�RE@�E�d�&��a@���p-O�)���~r�|2�T�k����T4� K@0����?���?y�Ş��ߦˇ�]�X���L��u�28)fo�!�.�N������z}��'�L�I6%�I(.�3hW/�$���'X���?�&��l	�n�K=q�� l%���ɍ�A��@9?�l�z�=O�ʓ�?����?��?i����5n�������9cPJ�rU�B$��o�����Iȟl�Is�s�������dݐ?�.�H1�@����s(W�?���򉧘O4�)��i����b���`��"*��;8��!40= �'��'��IꟘ�		ISt-zpʍ?]ɞ�F�V�" �	��h�	���'�z6MQ�<N��O�ğ�@U���_���[�ƈ�����A�O����O�O ��� 5����O7T��`��� 	R�Y�`�l�q̧.���	ß��aJ��X���
C[5B��AS�	�����������F�t�'�aq�m�+~I�g�'cg��h��'��7�U1y�Ɏ�M��w�L9k�J��=���l-�+�'/2�'�"ƞ�:����������)�`�h�˳~�}�����X? �O���|J���?���?���i�\�D)\m��8�cO����/O8Io�B�0���h�	v�s��#��P.�r�!5�/P�(MRч�6��$�O��3���I�/���PWb�/y:�ԫ!���>B9ib�gӲ�JB6�9�d���%��'.Bљ#�ې{
� J�%0�]BZ�M[��?q��?ͧ���Ҧ�,	˟��U�ɶ
�����#E�D���f��;ش��'�*�g��6@w���n�1/v�2Al�C�x�5E�8��D����'�����K�?A�}��*Mh��`G� N�P�SA�Y*o3*�̓�?q���?a��?i����Oj¤��-�,�bAӉT{�x ��'I�'YP7m�!!�ʓ��|�-CZ�ٔ�ļ�&I�A:w�0O�Hn���Mc��'���ܴ�y��'�24��� '0Ͷ��ajE�
�$qF`H!zP�I���'�i>���Ο,��6	2�E;�MK#4���c�"նI����	�Ԗ'�B7-S*A��D�O��D�|�Zmm�!:!h	+.��(D�Q���I����Ob�$:��?�����4p��m�	5��=�`(�|�d:��������@j?1I>�@�B7=H�t��4a����?Y���?a���?�|�)O�n�@w�rT,�',7J��k0�6�Р�X`y�MbӐ㟐�O`l��{+�HSc�9�V�Rr���(�ߴ h��ŝ$ܛ��@�hY�9��4�~jc�� ��3�����9���<(O ���O����O����O�'4�Tȑ�J�"�.���'7���s�i� MR�Q���	X���P1����$lY./<iǀҶZ{,Z`����?���w���O�(���i*���<�ys��>R��!Js%$.��7����'��'��I쟠�	�R��a���P���9���1! $�I۟���ݟ��'+<6m�`�����O
�ēH,m���/\H木C��.w�:��@�Olho=�M�c�x�A�&��H��	��QS�"��.L�ps�e�?N�1��t3�D�0����t!~��%$}�D��ፅ �"���O����O���%�'�?ɵ
A�ܮ�!�]5�uH�ʊ��?��i
\	�[��ݴ���y'��N��t‎�*	}��0����~B�'���k���T�v���>X
MhS�⟀tjU+*/�ە�	�3�@�)���������D̛��s4���i��-0��'��6�Meg���?���?���gيm�!&"�Pb�{F��?�*Q���OQn�9`
�I��jƃ�_`�Q(̬pΛ�F�<�"�ÎLbl��v�	gy���'*���-�����34c����'�b�'�O6�	��M�a	�?���1B��Y�d"��:l�p I�<���i��Ou�'�6�R��Ya�4h�<��u�L�g�>�˓Lؗ]/�Z$D�Mk�O~�؁�Y8����4�w�椹U$G:[l�7�"^��@1�'D��'��'��'w�QrEm�7��S�(��R��t�wn�<���el�g\���'A�7�8����P?�dJ�%V�!!�J�nZzt,-&����̟擱��,oZw~bIQ��4�p�-�`2Q�^[��M�s@R?QL>!(O��O��$�O� ��Jۣc���(� ߂���Q��O��<���i��]y��'aR�'u�� ��ŢK���i�W��!��	蟌�����|"�pY��ID��*=��HX0�$dwn�x�%W�Ӝ	�4wC�I�?q���O�Op���"��0[�=��虇�Dyr���O6���O���O1���қ��&C���EB�A�.�c��!����On�L��Z��I��0�T�
f�i1Lή<S0L������( �oy~B�9IX�}�4����p�ې�ܚPDp���W�<I)O`���Ot���Ot���OdʧfAh��c�ػe�FXI�@،6�X4�i���q�'�B�'���yrEc��.F��,���֑L���3h�}����O~�O���O���f��6-|�x���j<0p�D�7w{� �t�o��@����H�$ ��<�'�?�rl\�y�h�#Ak!2��C��?y��?Q����$�ɦIjE���ߟ��5IF�jl������r�(2s��k�Xt�I>�M+ǽil�O��E	ʩq������3���%��S�,�9g��p��'�S�o�ˇٟ@��"�,af�I(v׶��!hF�������(��ʟ�F�d�'F�Ey#�6Ԓ���=7a�����'�X7��s����O��ou�Ӽ�
�K�Lܰ"BޱP[�) %��<��i�@6-U֦pe��Ϧ��'���Q�+Z�?i�� �P��=�lY��0=�\��g/�d�<ͧ�?����?9���?���/2x\�`��V.E�$���D	��uC����۟�k���'ln�3�(*�b0�G�Rm�٠d��>Yt�i�~6�L{�i>y�S�?��c�_��	p����M��s�C�177$1�+'?1��mm`�dW������8p�8��#�6�h���p���d�O0���O��4���53�v�/ED�d^-娅�f��)�Z��Ö�y2�xӺ㟤��O�lZ,�M�#�i�8�۰,TW=ڠ�����G�f�Ap�@J�&����A�N��T����~	Kp�\,z�=���G5Eh��R?O����OX�d�OZ�D�O��?!�ABه��3WoTy�Ԡ!0��l�I�P �4t�\%B,O��o�D�ɟe^�d!��;�*ѐ�iJ��QN<�6�i�6=���ȷ�m���=��U�'��-��8���%1E@�WIQr���č����4�����O�����4kO��y%~d�WХ5�h���O��c��F�E%�y"�'6RX>i��)]Bk\\�E.gd0!�0?i�Z�������%��ǟ<VeճC��ѡD�7^��u
�?`3V���"��y�'���`SJ?	H>�PĄ497:�� 	��>��r��?���?���?�|")O��m�ts���'�E?`B�Q�.��x��Г2-?���i;�O�(�'T�oӢm�>�s�B�
�d������}"�'pN�R�i��D�O�}:��؅��s�(���u�M�ӇU�V���@�L�'-��'g"�'>��'�哜 *2�i�dО#���d,�l>�ИٴT��	����?q����'�?����y�,M�&�8��b�w��k�˓iR�',$O1�"q���iӂ�I�H���"ECE�)��
2|� 扟.4� �O�O���?���x��pѧӋAF�4���A?4�0 ���?���?�+O�<m��~ј�Iߟ��	R
��RPfВl�D�BJ^�X���?94Z�X��ʟ�&�'j�' �ADI�H��RqG%?A�H�<5���z�4�OO����?U(�1֤��c����\�j5�]��?���?)��?���i�O����]�@�9	#C�(����O�o�nw��v��f�4�4���ޱ\l�KāE2!�r\(:O����ON�d˅X�:6M<?!���%��Ә��`q���A^y V���%�p�����'���'"�'�XЊ���e�i%N��LSP��#[� ��4i��a����?!�����?�f
�`�*<�2!T*B�Ă�$�|y�	��	���S�'|S��#�jҀ
q4%部LP�l}��3�8��'�ܱ�䦑ʟL�G�|�V�0�a
�B���Z�o(g	�4I�@�ğd������ڟ��Ny��ӤɈ2��OЀ	TAvC~1d-�=~��1�4�t��4��'�`��?��46a����}�d�Q�	��Ö	[�9yL"�i��I'l��;��Odq���n��Q�u�5$G.��\a�A��P[���O,�$�Oz���O���#��z��P∣g���SP�\)=����	џ��,�M��}�D�{�l�O�y��53��2�� )�B�h ��g�����lz>����ݦ=�'�<9��%�Wt�`m@��@VN�^N��ɒ��'L�i>����T��D�4���Bۋ1e"-[Ӆ�C|��Iߟ�'h7
q���D�O���|j��W`��7��tѱ�~�-�>����?9�xʟ:akS�g�(и��K6K4�[���Ё��	|T�i>��'��p%��+c��r���HJƬx��n��� ��ğ���џb>��'��6m]�s�n! ��Гmc�ؐW&�)�6��ժ�<�B�i��O���'۫�լ���L�&;xݨB�&o2��5�{���mڠ
�0o�r~�/L�&%z���c��R�!�ؼ�@̊�Q>�a�����P���<�ߓ@�Ԑ
����&��"��a뾀:��i�"x��'X��'����oz�S�*C00��QZ����*�#�gP؟���%��Ş9Hb�:ٴ�y�A\� 66�8,�1$[���vݤ�yBcӟS�$�������O\�d��_��"�@�c0⭯?9τ���?���?�*OH�m�g�b�'x�&�# tE�`BĖ
���*i�O 	�'�p7�Ȧ9�K<r%$;<DL���M�%	>����
u~b�ǴDwlXs����OlL��C"IɨD��� NO
:��E��ڐ
���'�2�'�R�s��C@,O�K{b��B�4���;vȟ��p*�4��!+O�il�f�Ӽ���G��A�#k�m�<��p���<y��i�f7�������Ӧa�'۴��U��?)!��ɼT�Rd�U�!%<�-�-�!>X�'9�i>����<��������o�݋�C)d�d��`RN���'��7M�+�&���O��$4�9Otd����>/B��〣��d��p �r}r ��9m����S�'w�d���"G�|iᐣ0��8��OZ�#}���'d�s�`������|�P��y��٫�BI���Ă#evt�G :�O��mZ-f����	���XY`�X�%��P�������	��M���e�>���?!�iڬ�(��b����&�0/~����L������E'̰*8��+�	��ba�5B�8baҷDI mCN}8�5O��d�O����O0�$�O0�?��%�$i�Ɖ�!_�����!
Zy��'�7m�:P�)�O0�lp�I4(���˚L��Q��@e�I<!��?�'-�FEAݴ��D�9� .m�p��4��%��BI� �P��?9�j!�d�<�'�?���?I���u����h��[i�9�@�Y(�?!����D�ɦ��a��<�	�T�O�#�GV�?�a�LZ�Z���8�O*u�'��ir`�O�zS�9s�mR=Y(�ا��g��Ԡ������%B#?�'8%f����LF�x7���o�|�2�kИl,�x���?����?i�S�'���ߦq�V��0���mU�fT��0I-"X�i�'��7�'�I�����Ѧ�1��ԗ(c��@֭��u8@��wK!�M��i�r��d�i���(�ΈHV�O,�'a3�T�Ħ��B���S�+5H�Γ��d�O����Oz�D�O^���|���ܩf�|D؁��2|~ ���,N���ֆ�9�I��l�:��y���	V������d��A�ċx�6�����M<�|�Qω�M�'+�����n��,R���UW\|{�'(��������Ze�|�[��ßd!�n )�Y �,נZ`͈���ߟ��I̟��	Ey2l�"�����<���vu��(�|N՚��/E���+�˳>���i��6�Z`�I̺�Qc�ڽQ:e������y�HuR�]+v ��|���O����+K��AS+{V����Ь vސ���?���?���h������inp2eb�� YΡ��I�R���}�"������M���w��(K����	`B�G�N�"љ�'<7����1��4S�f�ڴ��$�q��I��'`IU�cK�g�"xSr��f�59�0���<�'�?����?9���?i�b��2I�U��Lq�D��4�˜�?�d��a!�3w�����?���0��6^>�	����!K�T��q�E\�4����O�nZ�Mk��x�O�T�O'�Haq��>��¦�I��f0Y�
6�����Or̀�FC�?ѧ4��<���b�m��H#~9-,Z���?���?9��|�)O�Elڗp�����N\�5&�d6�z`gۧD���I(�MӋ�I�>��i?7�禹�!�O�@�j� KD$�)��ځ�l�oZR~�̗=k�`���~�'տÐm®}|�D�u�ODA�!b����<����?���?i��?A���`�waL$��ڃ&d���BߋYB�'��bg��)�#;������$�x�)۠^�zQ`�k��~�;�L�%�ēu#���h��IC�]�7�8?٤gA6o����u�+e�(M�Be����	6�R*Hb��Hy�O�2�'1��U4wڌx�I���`�#�g��B R�'��Ɏ�M�w�щ�?����?�+���U3�����)V�G�y�e���i�OBqmڤ�McE�xʟl�y�#�7f��h*���4�$AZNƞi8T0FϞ�d�i>�h��'�T'�`�� �)p����ʈ�"�����V៌�	�l�	�b>��'ފ7-�
M T���Ȝ4^v�4mծ��i��d�O��D�覉�?�[�4��4�`��Mʋ�4\���	\(�<�g�i��7-E�{{6M;?��-��:�I1����8� |��&Nu�`�i�2�yb^���I�������4�	ڟ��O�L��-{1�:QB�q�4(ԉb��(wO�OF���O���D����]W� 9�+�LvyS�|1C (_ɦ�3�4f����Or,p��i~�� �H��!�9\��}
�g�!H�$đTx����u|T�Op��|"�d��m�g%�{F�XnG������?a��?�/O~�o%\�]������	��r��"ʉ,6J�M�Ɲ�0^��?!0W�8��4	n���3��N"&"�,;���<pɛa�9���D��$c�Ȍ:}r�=�|��(�O�=��*#��24B�9����U��1q��1���?��?����h����	�IY��I1�s��kF포���DЦq���RXyR�i�B��]�K��8Z0	��Ju}`D�5O�\��MB�i�6��I[�6m1?�4@�d����ޝ'�2��s�۽�Dp��#
��t�rJ>�)O1�1O�)J�Έ�k��@�s�U,!�r�A����۴c�֝���?Q���O��\;D��l���逥YQ�����>���?i��x��M�=Y0�ez�hʤrP5�W�Z�t��ӿiS�˓C��Т����$&�\�'O�X	�J��	��v�X�XW��J�P���ØdK��`J$�h|�HEh�m��Bd�b�L��O����O��oڅ,� �� N�9Ú�@�l�-@ PuzRJ�˦9�'� A�@�arM~��;��:u��5v�⌻u�I�����?��?����?I����O�&E�(�r���vjH�)4��'���'��6-��@��i�OP4oZx�I�G�����E�5��FŅ	hx5sL>���MϧcW���4���أH�&$D��eWx��r�̘`=�$Q�����?!v�7��<�'�?Y���?I��F�%�l�b"�I<=(E,Ŏ�?)���d����$��Ay��'��S&�y�%&�L�F��[�v�=^��ll����S����;,�12�E�"���3/)V��ȸ��59PZ���O�I��?I��!�dF7.�u��R4w�T|rd̘"4J4��O|�D�O���	�<��i�����2L�6)��F�\���a�R�y�2�'Z�6�4�	����O��qu1P������e�$p9��O�o�+,:��lP~�显|X`��q�I8&���5'89�]�vX�j�<����?Y��?A��?�.�~�c��ݗJ&���#]�$i�aC _��5Y�ܟ��	���&?���2�M�;u�3,Ї
@��� D���A�iC�7�CP�)�S'h/f�l��<� 8�QD���a��L"c0袰<Ob�ib����?�1&#�D�<�'�?��i'�n)ժ
�,ix��G��#�?a��?����D���P.y����埼��a�P��1#��#,��
k��/��	蟐�II�X��
A-^P)ؖˎ����5��!I� l�ŢuB�����sѡEH�����b��.��1�c]���	ß<�I֟�F�$�'`�%�6���J��`��͕.�0\���'G�6�F0#����M+��wZ�i�b��ज़`(ǻ%�T%��'�2�'��C�V����8ʑhɹU��Iw�\��K0�B$B��2�ƓOJ��|:���?a���?Y�^�Bp��_CZ�YV���0n@�.O��mڗj&f������Im�S��t 僕�;x13b�Kf`�a�)�	����ɦ�ܴ7N���Oz���Fʔ�G��0�'��չ�'��=L���O��sw㌎�?1u�(�d�<�%BWȌ雂V�hY61�C�R�?��?����?�'��D�ڦ��g����/;�\�� ӣ ����X�� �4��'��'C�&�s�Z�mZ�&�x����.UiI�cΓ+L1�`D䦩ϓ�?9se�)ZN����E~"�O��f�Ou.�KQeW?�@��B˖��yB�'jr�'���'Kb�	Ǌ-�©ATC?���S�5�v���O"��F妵��v>��	(�M�I>�ǂ���4az������+f���$�Hش7���O_ji���i>�	<�>�������=g�|1�2/G8r�yڱ�'(�'�h���4�'�R�'sbQ����}�$�%ͳ���Xw�'$�X���ڴ@.�8���?������;�~��&���5�9�DcH=,���%��d����ٴ[*���iTҡ[���H��w���q����Aʴ`�a������h��AII�Ɋt/����M3l����vC�	��T��ӟ���ٟ��)��Qy�f{�6L�B������Gl׶Fc.`��ܘ5����O%oZG�X��ɑ�M#5��!)bF(�L��5VL����l�F��w�q�b�/`p���矐�Oǖ��
<f���J�A&�.U3�'��	��P�I埄�	��Iw�䍌�MI(����A��=y��C5��6-ˌqs�ʓ�?�N~�����w�0�1���P,�ْ��{�t<�r�'��=��� ���6mu�����v�h�F%�`.H�§i��j7���iQ�d#�$�<����?�m|��� k���P/�?���?Q����ɦ墒o���	џd�B#�2F�����t׾�y2��w��!]���	�ē�Ne8�ٝ`{���U����'����A鈍����/����~B�'�<�[eɔ�:���e�T� ��'�R�'���'��>��I%+��(;s� �u~����s�6e�	��M#F����?��WD���4�NPQ�n`p\p�H�H�z��08O���O��n1(�!lZK~BT�T��H��.?�XpM��!1��Ɓf` )�H>�-O*���O ���O����O(��p'V)T F�G!��}\8� �<)��i��I��'���'*�O���ߺuʤ���	��^�z^���>���?�"�x��$�#5���.��j������I�p�\��'"��!�)
K?aO>�,Orl5k��3�r�xQ�8Z�:	`�'ɠ7�ޏU�z���}���b�eN�E-T�r�d���dM���?�2[��	̟��ڴe�T�:ƷdY5��(�D��LB��]l�w~2%V#=���'��'促o\9+� �x��Vm�(I���<�
�2#�Q�OǶy�\D���L?{�H ��?��~���T���)Y���'����Y�Zg�axC	ߕa,���oC��ē�?��|
����M#�O��{�lI�I�t�ڵ��Ptd��Ąޢ���'��'R�	`��B��X�=�|qQ����q�<iGxR�pӦ�Qs��O����O��'5uPu�F�-W� ��:rd�'����?Q�z`������s�����#��n�8��M��L��*��zF�7�Uy�O������"<�H��'D*~��|x�d@�(���j��?����?��Ş��D�æe���B7i��P������s��H�2�(|�'�F6=�	���$�٦%�T���.�<��ƪ��9�0b4E:�M�Ƶi��-���id��4.W<��F�O��'"Då��#1�ԌZdc�A�Μ���D�OZ���O �d�OH�D�|
�gD�i�����?I�}���F�J���	>��D�O��?�r���c�g;� �@	�I��F��?�����Şƈ�ش�y�fG`�� �߷�9�$@կ�y2�B��e������4���$I�TM:4��Cq���Y�����OJ���O@�D�<�i�~��'dB�'���8$���P�`�3���8:�h�G�dF}"�'jB�|R!��dh���}�t��䚊��ė5�Dd#df��c>�&�O(�d��^��0h��n��hw��<�(�d�O���Of��&��#7!�����B�l�@1H��c��?�Ӹi`�R�O�l�\�Ӽ��IW5th��IB�P�#{.��%��<A���?a�=�LKݴ���ɞx82��O*�"U�R,踑��P���|�T���<�	֟��I\�㋆�mn��'%�T:��v�My�y�(���)�Oj�D�OR��h��Ђ{O���G�M��\�0�{�xe�'���'/>O1������ R�l�6���z�y�H��7	]0\=�ɲ��Ո��'�zH$���'�� �"�)s�H��e �qr�D�#�'p��'7���4V���޴`͘ԉ��Il&&'ؘ:(����,��̓z`���\}ls��Ulڥ�M34��Pܞe���%8��<S�a�y5,�	۴��ĕ�0�����O�'�F�v�Z�*� �z���6���y��'.��'f��'�2���'����Mʢ4?���soHBKZ�D�O���ঝ�rMi>-�	��MSL>I�B�D�z�%߆3���Z2*�@(�'Gl7mM��	�ho�y~�HE��r����/z�<��������J���آ��|�Z��ßd���<�$$�(Z*����k���֦��p�	ry�g}Ӭ�� ��O����Ohʧ��F�]��,�`^�1��'�:�!���Ӑ�%��' �T�iLuծ���E��,`��( *րK�t�R�@~�O���� Z�'A4x13BK�T�bȱ'�Qjѹ@�'��'`b���OW���M����}��QC��K:J,���*B�L����?)հi��O>}�'�7��c�b}z�햧�rYfo
�)��nZ��M$CD��MS�Oxu���U'�
N?��E9�bQ��%׀,��< �	q���'��'�R�'8R�'#�+4 �a�'Թ?\X$f�1�@!۴ט���?	����<���yG�)�l9�Ć&��ų�R�|"�'gɧ�O~8���i��D�Q�,�a� ٰ$_`:p�X��RU
�	{�'��'��i>��1#(aqW�Eh���LB�d�����ޟx��ǟ��'=�7�S�j:�d�Oj��ק/���a�cc���f��%�|�p�O��l���Mkb�x�N�5x���هjX�#���� ���հG�˗�
21�8Ћ� 2����1�\���)�.e��0gM�$&\�D�O �D�O��d1ڧ�?4���_�P=��B�IB=��X�?�w�i�t$AY��
޴���yWl�l��8�ߚ0�8�"�+�y�F���o�M��R�M#�O`@��Y�r�����օ��fˮb�"|ö!P*^51b"
ӄ@hTC�H�2f:���&,�h�h%@8N��܃7#U JvѢ���$���K� �+�~��G�-c�|��Q�.8	�so�qe���V���@��3�=!�. ��E�ʁJ� ��i[��ũ@KCW�$X(� ۂ頁�"�(���P�̀�,�]�Џ�m
� 3��K�t�h3ވ��ax6���S�^Y(�*ʘs4�AK#O[�W (�Fl��t�z<�"�:۵�����9�/��g���M^�K'p�Y�Ƈ!8HP��;���Q���+}� �$O[�\�����M����?A���"������
�M�,u���˙L��I�ez�T˓}�(Gx���6�� Z~P�-k����Mc�8�>7m�O��d�O��	g�Iҟ��WNC�T0tx&�U7(�*谵Cʁ�MK2X���D�DW*4&VX8P�^}݌�ks��6z��<oZǟ��	џ���+�ē�?9���~��P�$�8�(��2o�D���S���'�{�y��'�2�'�p+&� ̚ܐ���@d��u�����US��&��	ϟ %����,�&�F�*Q*�R��׻3	��3J ��<)���?I����K�}��Q�Un�!X����7ʃ�q�f�;Í�u�Ɵ��	A��Fyb��"�I9� Lw� �Ζ� ��yb�'0B�'�ӆ0 �e�'Q>�Q�m�����6b�1��'����P�Ly����\�"ü����m�<xc*G0f��IП���՟4�'_Z-�6�"���0x�9C��u	.� C��,\؈�nZߟ���eyRT�����%�'ͬ��0�������ŉOc�)�4�?�����E׮e$>����?}��W�:�,r��&:k̥�G��ē��/�}���	�CĆ��� Ú]q��Ӧ��w��fX�l�f(��M��X?Y���?1S�O�A� 
\��*gڻ&��8Rf�i��� X{P#<�~B�وe�K�~Ɲ1��ej%[�Mk��?�������$; P>t��GYo��(�����F�oڹ} D"<E��'*��R�KϬO�J�`YK~���,�'�Ms���?��f�8A��x��'Lr�O�tc�P;�
}ؓ��&B���5�$�P1O����O���:c�x�m�PV����<���m�џl�Q�����?��������C[�f�Z�;l�B���.Z}���$̘'H��'��'�r���⭐EM�o�1HP��9�_�p������I{�����I�H���إi�����Ԫ��#��mc"D�0"e��?i��?����?�r�����ȼAB�a��>���KT�܋�M����?I�����?A��B7P̓���A�!�݇&�
!���BA��Q��>)��?����?�M���B.�t�$;d���a��J��c��U]J,l�8%���Ijy�/����$N"��F��:�d�F昭��oџH�Iҟ�	�kw�L�OL2�'8�@ն~eYE�M�9y)�2���GM�O��D�<q�U��u^+A���	Ѯ>��z��D��Mc-O�14��q�	Ꟙ���?�z�OkL�$d�X�k���
{��8sᔻ~����'�r�Q�;d�O�>=��f��|>PUau��,��ER��p�t(ȁO����I������?iA�O�˓-3J +8$uq�g��1�hQ�i��L�a�d$���܁�)��m�`�R�>$��}��$��M[��?���_(��W���'>2�O�Dƀ� .���ś#ׄ�0f���e1��O
���O�DC�? bHғOR�q�St��.2NB0���i{�	�tB�����O�ʓ�?�� ��4��U�q�m��O �;HD��'ϖ�Ӳ�|��'�R�'�I�tɖBmL�ರ([�9~&y���K%����<�����?���F�\ʓ��$#N9��`�vjB,a��1���?���?A*OM�DY�|����</��h���$������'�ҝ|B�'����	���(_2�hU�͕} ���E�6G~�I�D�I�<�'����ϯ~Z��_d��­R�Ftb���8Cڜ[��i�b�|��'��'�7u-qOJpc%Ɨg�D��1�Id�5Y��i�"�'>��6f�	��t�$�Ov����,hh��q�����c�T8VW L$���	韔i6"Hl����t���1�.�c0%��v���ǋ���M�.O�P+�F	��m��������?	��Ok)!��$Ⲏ�+d������4ԛ6�']Ҩ[oI��|����r8�D���~HxW\Y˛�e�aHn6��O��d�Ot�	M}�^���o[9cuD��#Y�O�ظ:����M�W�ƪ��'����$�1C#$ۃH�L�u��}>��nן��I���Y��
��d�<����~�(�>$���"]d����#2��'�����|��'���'K��R���P���	�5�,z����F^��9�'���h'��X&?���`��1C4`P
��4���l�D�I>q��?!������P�~�BfB�#�\QXgԩ�$���m}�Z�L�	U�I�H�I���-A�M�W �9RG����b�X���`�I̟��'�:؆�>�wAƔ!�0	���fa�G�p�$��?�L>A���?�%jF��~�K�/�d�FC��q�iA5�����O|�$�O�ʓp]
������˛|���)T��6X���P�fȨQ�7m�OL�O���|����S�w��8>�����-z �4�?)���D"��E'>����?��/�"�� C�C|U�U%C�cN�O��G��L���䧦�)^�n�,q�CҋO��@������O��O��d�O���r�Ӻ����
8�d(��E$X��a�ަ=��ڟ��M�4?�c�b?!�f�Qh��`A��%��X �hi�x`m�ݦi���8�	�?M�K<�'"��az@�S��۷!9S�%�f�i<$����'�rS�0$?���q���}�ԕ!7�X�����i��'����"�)JO�xz4[H ��uA�-�ŨE��'#�q4G:�Sǟ�h�L��4F�V��I��#�y�5oZ��3�uy2��~ڍrj�FnL���`]).Ъ�L؟	n��. 9�o�r~��'B�'�剥V��T3$EW�6Z|9P�.�^��)�dK��ē�?������䖄&l��� J�4�Տ,q�\H��f�O��O����<A�n�n�{�O�9���O<T�B��k��H���4�?	����'�b�'����a�H��M��?V��g\�|,�* ��n}��'���'O�I<��,�H|b�O
hN����K�S���ԧ�.9��'��'s�	����IR�i�5R�(Y!ʸ-
-�QfW\[�V�'<bS��&) �ħ�?�����Gְ~д��U��E�<AB�S�IybD�.���ӟ<W"��3\�����2,M�+�Y�����k+���Iן��I۟H��YyZw�N����%R�������cܴ�?���S��̻ŌGA�S����	a��,C���)&�V�_�:5o���N��4�?���?�'����\c�.x�b�W�Z�Y�-�D�*�Yݴ"���b���?����?��'��I�|"��X�Ni�%IX�i�>Izv
=-���'���'ײ�˱W��'��n��}�u��`�`�� ɞjJ��y�$S�b?��I~?A�@�[�P���O&;R�yQ�����	bN���'��맸�'*��E�P����m�8P�Hd{���>���4�8|�<i���$�O�ps咿bV�S�ΐ&CPX8uj��V,��?����'2�'-�EP�M���T��[6�}bq휛T���+�yR�'��	ٟ�!���u
� 
�&|�ш�6�����-��ǟ��?���?����\3<�oZg��}�G���HtKf[!�>��?����?�,O�ԋg �I�/r�@�!ҝ1m�58��]�;Ċ�ٴ�?�K>).O|Pa+�OL�O+��B$�n��� 	��	��}�޴�?)����;$��`�O�r�'��4j�\��IAT_$aj�DYf��hF���?Y���?!�H�<+��?٫e��v�:!ڦ	JH�����vӢʓj�D�Ӿi���'�2�O���Ӻ��퀝/%4�nJ3޼�㵁���Ɵ�K�N1?!(O��>�p�#Un��� ����Q�2�c�y{�
��!�I�H���?a!�Ob˓��	�`��<����f�$���i��(h�'���'�����O2(@�o� W�zh��5l�Ԩ�LCŦ��I͟x��(Hݖ���Ozʓ�?��'G28��@���U��oJ�Zaش�?�.OT
G<O��˟<���<ؖM��6H�Qo�p�݊�ɧ�M������S�P�'@�\�TZ�wI���L��%�wɂ6-�1m���ɗH|�x������֟���Gy@�P��0�&�kV�y��GCDhUƫ>+OD�Į<��?��
���0���9�td��� Y��<���?��?q���D(6I���g�? 6u�������7]Ntv)��iV�I�<�'W��'��/�.�yB��4�P0��
�=�L��lHv��6M�O.���O��ĸ<i�J�
<��S�֘�
m���Tn�6!��	����7��O0��?Q���?�#���<�,��v� �E:���i	�Y|�m��e���M����?	-O�t�F�b���'r�O�p@e�$��4� "Kj<���>9��?Y��X�.d���	�Oz��!l����抟��	���A�v�7ͺ<!�,�g���'���'��d��>��*ll���3)�5y2A�}U*�m���I'Wx���e�	w�'�0I�ER�d�y"�Y y>dm�&;��ٴ�?1��?���_0��sy"�I<k���Q�#�M����{k�6��y���O�ʓ��OR2	�w��r�E�	��͂���6��O��Ob+�AP}rX�@��G?i�K��F$:d��e��a���j�"�㦁'�̺��o��'�?���?��[&&�ղ#JO��	��U�m���'���`ƴ>�.O����<���sw�	�93�D�֨�t��zC���!���h��(�Iݟ��ǟ(�'�,��%EN5I��)��H0����@Ȃ�\��꓄��Or��?���?I��(;<(0�#@&S�8 aC֊0��0Γ�?!��?a���?q,O�)��"�|�BAҊW��|����y�⨸���i�'|"V�l�Iԟ����E�	���� R�ޛb8�Th�`,xQ��ܴ�?���?����ؿ-Q�9�O�"Hz�v�2�J�tc̴����B6M�Ot˓�?Q���?����<�I�x��L]:j���y��x��a��n�,�D�O�˓Nz�2�^?��	�L��7u�41��g�[���*D��%�X�r�O��O��dW���|Γ��4�ŞCL�1�L<�z����M�+O@	��kB�Y��ܟ��	�?��O뮕#�����Ş:`\@eJ�✘3;�v�'��Y��y�V����pܧz�
%�C�kO�q$>钽lڗ}r�dX�4�?���?���pH�	ly�+Y�%�N�7�E�UaDP)`��>�@6M�����O����O�r픢y���ʗE9fi�
A6�O����O̽y� B}�U���j?9��G�}�:�s�޿mp@�d#�����Gy����yʟ����Ox�Ӡ'[:T
��@�ԡQ�L �7M�OШi HCz}bP�$�IByr�5V�K�n杸�m�EP������Үh+�d�O���Ot�D�O$ʓ$'���A)b����
F�^B<4���ԍa��	ry��'��I�������X"��!-�J$*��G	KjFi�a�#i���?���?Y���D�zn�D�'eEX0��
Ϸa"j�J�l�`��}mIyB�'��Iɟ��I՟p���x��؄*tv<�ĈP���(:��O��6��Od��O��$�<�˚	3w�S���q�:���Q$ȝh�H���(��M�Ȧ��'j��'T���y>y��4+��@k�e�,7�Z���KDϦ��	͟��'�,��o�~J��?��'К$��ܶR��!�Gz`�tQ����ϟ��I6����D�?�Ib�ِb���V��B �8( N`ӎ��@2ַi���'���O>��Ӻ3�i��D���c&n�\��]����	��d2�h������(��ZM>�X���S�4@��쑵fX�7�[�.
��n�� �I֟P��!���<��)C�_�D YFL��
�����&y]��n\��y2�|��i�OΩ�j��cp,(cFC1ö$��RѦ���ǟL�ɤ9�b�1�O,��?��'49�㫍�=��L��i��,���4�?�-O��a%?O��ڟd���<�3d�$�� �0��v;8|�b	[�M�@*�u��^���'�RX���i����W�l�)��
޶�~P���>馅��<���?���?!���䉣:��S�[-}3��`�X�6w�$�s��`}BT�T��gyR�'�B�'��3n�E����ڂ0>���C��y��'�B�'d��'�剷m��p��O	0X� Y�U�`�bA��5�ZT޴��$�O��?���?	�)��<�T���Oz��zCĝ�xu��O����'UB�'��Y�<��n7����Okl�;����#L�d����`�ۇ��v�'��	ş���ş|�t�X�O`MX�+B3q��0�C��!Z[<p���i���'z�I�Y�$ȭ�����O��i�..6��`��G����5��0	r9�'6��'��CH��yB�'��n�!'%��Y�P,��-aW�W릡�'ؐ� me����O���P�ԧug]::H5x�5����0���MC��?��.��<i����?�S�G<޼�u��?��8���N':7-�'�2�l�D��ɟd�S���'8ހ��Z�P̪Š����U�=c��~��0 ��O��O��?��	�k��}[b"КK5"��v�\>`��	�4�?Q���?)�h�?D'vB�'��$�,fᥫ̷ ��)3�ǤK��O����2���Ot��O�,��h�G8郄��M�������		�r<zJ<���?�L>��+�	�C�R�H�b��#'����'I��:��'�������ٟ(�'R�q0�$%<��+�5�B8��ϛ�dc�0�	h��4��	�(�ܷ6,6�! ��?����3���t�'kb�'��]��zDnj�OܩQjG5�h4���N;=;B�AK<a����?i��K����#�m� AQ?֦�+Ю�(e�6U����ן ��uyb��u���*H���9+/���"�3X���@���1�IQ�I�4�	=|YT��	\��\	����n]�p�� �Y��!�ݴ�?����
J$�I&>��I�?!�� ��c�T"E�&�Q���-vp���x��'���>{|؟0E����.aC��  N�Gop0�i��I6	�a�4/�������䁇pG�$"P�I&�"��sE�7d��'Ç��y��|��H���X'fK$�q�EV�\T��͍�+ �6��Oj��O��	�X������W�<ʂ5���DwP���i��I���d(����a���n�0q�/Lv�H�C�:�M����?��O���x��'S"�O��M�/^<y1ah�I�)�P�i�'`��&�8�	�OX�$�Oh�r ^�v����Ii���kZ���IY�8	�J<���?�L>�1C���g��K��%Ya�Y�<c���'�F|[��'����I�8�'LjY��͔=Qq@5�f�ǐ<��4��?&Jc�H��M�I�L��J�r=`�n˷0=
ܲ��.`U(��sC�ßl�'�2�'X�]��£������j;�,a0L�=j�U�����?AI>Q���?�a͜	�~����s�<)��g�� Z�ii!c������O@�d�O��%RvH�'���i�X뷉���L�W.M�mo��o�؟&�p��؟��dy���O�$S��!�ڀ�� :rĘ-X��i4"�'>�	�/���O|�����J v
�k��]+/\ycQ��9p��'��'7�T���'i�'��)�,�z��I*�6����U�TQ�L��M� [?9�I�?M�O��X���`�����!g��55�i*�'H�l��'��'|�Sh?��D�=삙�'�Kz:T���U�S����M����?�����g�x�'��e�#L�/C6��ԉݕ)�HYc���Q$�O<�Of�?��	0���S�^#c H�Q̋�9.myߴ�?a��?��뉥Y쉧�4�>с�:�:�e�ܱ*�������=�?A��4�'\2�'����@FK�~l�SQ ��~��(a���Ĝ]+�-%���i�'u�p�Wʱz��8ȡO��FQ�UyN<�����D�O��O�"6�W��anP�ɑɔ�iC�R�R���'� �	u�'��DI�G��#��01�^p:��R�g����'���|����L�'.��u�v>��ȁ8m��m��Y 6�h+ct�˓�?�/O���OX���*v�=/��0c�4�\y�Aڀe��Pn���4������ISy�A]eF�ꧢ?w� �.�N� ��S�-G"���¬<����'��I����Iϟ�YVn&�s�>�ctj��,n����"ض��зi���'剶'���!��0���O����)B�l��P'j�bB�4I�P�'lB�'��)D4�yBV����jңI�M��}Pɓ($��I��@�m�'0�x�%z�z�d�O�����FIקu'�� <d�h�NӺwH���ߵ�M����?a1)��<��X?�	zܧGp�s�*Z<,�Y+��G)k@��mZ�h�T���4�?����?	�'H���Oyh� NZ4u�P�U(ZҞ��7����6MԜ(��O�ʓ��O��D-b��)��DV1X����Peդ0��6m�O����O�,b��OT�$�|���~b���/>������$UL+���W�f#<Y����'���'7��:�A��]ZĜ2P&
/�x��es�0�D�P:�%����8�Iu�ɂB����3��!�7�\�Q��	�2��b���ן�������I�@R�gޮXϐ [�"FO�P��f�YyB�'[R�'v�'ZB�O����m�1� �cԩ5��<�3�i�NP��OV�d�O��$"?�S����ם�cP��y��@�=�ȃ�^�d�O��d"���O���֓���3'�L��㤏% ݲ�2�O(t���?Y���?��O��PC+�	�	�T��醺5<hYf���H�l�ҟ�$����ҟ��6�.���>�x��-�_J Zo�N�P���)b�>�P�J�m�X�'n��OA�N�M�������d���.���y�̆*��W�,��a��4��x���z����/Z2#����c菀'��	��T$�����l ������!V*���U��;`Ԓ��*lŁ�7�UC�e
����,�#�-t�	�u�[�6�01��I��$� �^5K��l�C.��tYg��zȒ�2�� ����C؅Kk��ao�(8$>�����t�����2_w�u�R�ԹB`�j�,��vv�M�G(W
��*�皭l�����V�o�1�Ru�OT�QR�ҽ 2|�y�^/zVj�pE��5�e!�Ç�2�7D�RԘ! �a�Ծ�qyZ�]�G���3��}��Eە��E��M~�KW��?�'�hO�d��H&�h4D-B/8�ȑ"O��Q�!�Im����N����6�����?��' ��6�� X@��-�b]�Y��H�@~~Q[��'��'�b�qݝ�	���ͧ
��iSc�)^��Q����03�����O<��%Z15i�XS.�6#`�w��P<�����4k�QU�ɤO	�=0*�hӴ�!$�I��`�	q�I��T�	w�_�v,�Dg�.`�"�!T��(E�-�ȓWȘ�:��ѵ��5@���X5�<��_�X�'��kᅯ>q� ~�1�L�;ר�17I�/y*����?�6m��?����aA_���TO��CK����i�r1�F.ؽI���K'V.��X
ǓH�ƀ WH���-)E�/�M�1kB3C�i�NAR��4�@�y8��D��O,�D�<!�n®R	ZA���B�~��㥨u���=� �P9�A��T �YK�/�h��COr�n�$h>�3��#Z��!�oU�<���I|y����w����?Y.����O�O�uâY�`��$��`�+Dh!��-�OZ��L�}$37B��j��pPd���ʧ��i�/�	A���`0գ�$�#��F(�ӤM�	fDy��L��H����u�_�|*ݢ��O�0ޕ���>�u��ןt�IR�Ox�B@�=�`�qG-������y2bV�(�� )u�Z�$�-B��;�0<�2�	�7J� ���>2j��	Q!B2|>, R�4�?���?i��w����ɟ��Işt�iޕ���ތ~�!�l�XŸE�'y�{�`Շ�ɖD����!]?.P,D��̈́P7��؋�D!<Ox�`F@�/&�8�L�YCp��1�%扩[Cx���|�㘻*Qp]��ȫgyH�����y��'Trz ؑD�a6�9)������Vq���𜙷E߶T �䑕A\�;�,A!�O�m���O`���O��ğֺ���?1�ON�@�)�%�`�b^�@���:��[�x�͙>b�F�@SEػ0�`{B+D�kɋh<�v�Dl���� i��`�-i��t��	|�����ML�g	@�	u ��c�H�1��"D�<B�獼������%-�f��CB5�	���'3(Ćd�����OB�ҵ-�5&J�J .I+(���7��Ob�W�����O��&��d(��ǃ|PTbǔ �2CZ�&��x2�]���'��("�)��$ �荱|��u��3pXL�Id�	��Bt�L5L��R�l�6_(C�	KЄ8�-�W���YRd�v��C�ɹ�Mc�S�L��+@M]�U�=�S�G|̓f�v�C�i'"�'*�ӣj���	�0ߐ4��J>����Ӭ�p� ��I����3�Wҟ��<�����Z\rd��ߺt��1xS�ɀ��V���Fx��D����ѫCJ�Z'6L;è�'��I�^�F��3�)��X���O��V��1{���:�TC�	)2�}iG��}܆�8"ΘG����D�'��L rb�2]�0��­iO��ْ�>A���?����J������?	���?�;;���a7��6	kz�ӵ�J�N������\�F�\�8z����]�g�	W�N)z��T,E��y�!.D"t��l@&Mݺ k�	�FU��$��|��.  q�@��0o���Z�E�����$�O� ړzPbP(13�� &; *1��C	���J�`-r�*��'2�
a�'>�#=�O+���ݸE�R�6�Fْq���Y�(��
ׂ�,��I��L�I��̰Yw�R�'��D0f����U�ތX�� ��F�>�n(�M*"M���Y&ޔ�P*�Y�'@��s�>_� ��I�.
u���BfĨ �a���4�\i�!Ł����@;l� �Q$���aE�&p�v�e�'LB�Y�8��̀�q|����� 8�ȓA5r�1��V�1�uhƵH����<1��i��\�������M���?�Eևb��dj1I�
A��fY��?���j#:�H���?Y�O�hԋ���Ab��F���ґ�!&&)�px���8	S��T�T"MR����.V�q�pȩQ�5O:Yɲ�'[�'H��/��lH�i �R�B�4��'2��H�a�7���'
�-�4a�
�'�j7��6)��d���Ku��=+Մ�z]1O A������	ß��O���'��C�F�2�����D��V$1��'�"�C��"�T>�o��9HfE�j}���Al6j��Ot�j1�)���}O*�Q�/��]\V(����V��'���p�����O�8<I�O�#��CR)E#LE��'�a$/Q)dM�b	6E���Óv������-kZ�3# �S2��D���Ms���?���f
��B��	��?	��?��Ӽ��DNbZm{ÇԆ=��Ϝ���'z�$��d؜!�o�"gæ *I�Z�n=�=9g�Wtx����G��M�._.rB� W�H̓qF��)�3��د9*p�$/As�1�U��Q�!򤓯"K,��q���F8� ���$M�ɜ�HO>E�!#
X� I���9]��[s�ѣ^� 
������I�|�	��u��'�R=�����2Jm|�#�cR�w%�I���B�!�$)|��Xq��*9w,w�s���P�O�Hq/\�`c�9R�Q�X��U�y�r�'�za�0Τ%	d�fѦA	�U�	��� (l�0m�C4�m�K',y�dw�d�X� �B}:5�i^��'pkU�E�6��uI6�
:���;g�'uB獪d���'6�)�� ��|�яF��dp�-�-SR9#fL�p<!`G�n�~�v$�ŭ�F8�}�#Ƌ�W�����ɶpF��/�D��i�HC�ٖ&1f��P�+>�!򄁩BX�;��U#OD\��'��B�!�d^֦��u�Y�q}
������%T��!�5�I:=o���ݴ�?����I�z����
rꎕ2�`�9��QfV�[5���OF��j�Odc��g~�揭:p�@� ��#���ɩ=d�#<�B���>P��#�q�X��l�dG9�����̊RT"� ��j ��C�\�v�!������PzAK
'�sN�u�r�'��"=��ѶE�pe� &��}�X��×3^���'C��'���ٟm���'�2��yG/әQ*N�I3�s�H\��.�
b�1O�ਲ�'�����T=o��2�ˤc׮<�{�ߪ��<�cm��Թ��0`��-peL�?��'��-P�S�g�	�u�X��!!�lp�fR�R4�C�ɧ.Ŝ<�׭M�W�<A����(E��GP��"|�fCI4�Z)�l~�&��1N4��3FH���?���?��4�N�OT��`>�;ĊאA
�򆪁4�HtQ�d�*Q�C�	)-��0�$ɕ<�j���+I8f��gD3������/&�T�!�͔R8P��Z�?�
��V�r|r`���x��a�`M˶|*�e�ȓ'��wG;]��Y�p��L|���<y��d��Hl��l��T�I<��e�s�ՑZ�ƉA��Q1=^%�I�* `\ڟl�I�|�d����%�b�b�'$��H��T�j��`(�e5O�,9��d��z%Y�$߾3���Å�MJ��x����?J>�wAѻG�P�)� L� �1�b\c�<)�D����CWg��4��� ��u<�0�i�n=k���V�麳�H����(�yON>4��6��O���|a�[��?�A,JM@�� �,� BaM��?��O8�hr�iA1O�3?�A\7;��B�qV\@�L�Y��
��z��?�{�b�$�^U1�B��+����+}Rl���?)��䧛�'�1[��X*L�Gk�mӸL�<�����<�w+�w��b�@<EJ���D	R�Dh��DO4�rIp��qW�h�C��-eB��l���ן(�M�0	����I�������6&�X�(_���H�$`�rh�<�N�}x���j�.6z��P�АqA�81+�	(V��Y7hx�y���)J� T��)�OF���&?���S��>���O��d�=ukRp"$ ��.@��)G6:^B�	�-���3��Y8U��(�CE\�-*"�U����DC�U
����	!+ml-"���O�!�
/t��YFJXDP,����fy!��d�Ƽ넊F;��1e�P�Py�h�#��Q)&�
p0Y�ҽ�yR��-(9�]� b|�ax�@T�y��K=w
��d�Iz�X�b��y�m�9 49�)A4I���B�y���=Ev�	i%�|��6� ��y2e�0ODq�dI
a4iC�ʵ�yB�
N�v���lCM���@��Ű�y��S2��pb�B�8�"ԩ.�yFE"I��l�<�H�!��Pyr%�"&�dh�1�^�hD���V#L�<9��?ݨ�H%(�a"��H�n�E�<�@���G�БQLΤ!�dY���PV�<���7D6�9 D�ɩH�3ǮR�<�7z���w��"%R���y�<�0lL�C&d�2M�Q2 �r�u�<i�)H(]�N�ê���4�J'�s�<!D�Jc��yZ҂͋D�ȡ�/Iq�<��T��L� 7�Ɇ}B�urXH�ȓo\�48d`��*�� X�c$X^u�ȓ)�� �P@֢m4�}a'H�l� ��S�? z��a�PB$�H��×=�pI�1"Od@*����/�P8��Ƃ�t�+"O�P+��ߩ.��Q�S@=t��x%"O0���fY�+�@B@��1�m��"O���w�\?B��c#M�8E��`"O����Ȑ93�Ā����*ӞU� "ObnsS�k0�H���c"OvD��<�T)Cĥ�e���`7"O�꣪�9!>�$��d �dV4<*U"O x���J�t˞Qr�G�8�|���"Of(�t+��VZp��smʣ'���"OBH��b��h�ԫ)�*�i�"O��Q�]]�@�뛎��m0"OZI�7.�!Cht%��.� 9�"O�p�w"9���* ���a"Oxr�B
b�M����n�ʕ"OP��a��1��tha�O'2NT�"O�Qr��EX&�q[��Ŗ	DTYQ�"Of�[���^��m���G?1H��"OޠQ��M6� d2���>V�:�"OJ�
U��|MvM�4@&SzU�"O��� C]�=�F�)�X�~0�#�"O��`�
�)���'��� �>�)�"O�q��/���*`�`�ժM�]!��'~��_���z2�ݲL@��P�'��@i��Y+�>\Q���RlP9�'c�$�&�ӑIP���J�T�"�'�}i!F�0{E�S�ɍm�p݈�'<�9YE�_]T �
  �<�4̓�'R><!�a�8B<0���=j���'�6�d�*�B�����wNU�
�'.ޝࡉ�WC�)`UGI�P��*	�'`J=i�IK*cff����P�y
�'�@��`+Y�}��j����F��	�'� ���\|�U�U�D =�����'�lX8ԁ�J|�)GL3���'� a��@/J���zWjݬ-�z��'���۔b�;����F��O&��!�'*�,
i
��`xѣI�3V� �'y���
���H��F�D�6�`�' �bě�xIL�cӍ
	DZj���'!�PJ�ě�/&�x�⡑
8��q��'/��s%, ��<��.�7�\+�'q�k�+�!;�8���l��6?Z@�	�'.��T�	H���3V�29��	�'W��s���Z��1��:VŊ�	�'�̅ˠ�S?��13ԛ{Q���'���5$NT#���-"�4�	�'�\m�f���;��/ �H	�'u�����x��e�������'b��r-�t��d+���&F�Tp��'� ��i����#�-r�2P��'q
 �W-е{��x��؉eT��r�'D.���j�#]I�@K�(߱��\0�'�h�ـ(B)Q�V(+Q���$	�'���
���|�!�q�а~�Π��'���#�ށH��I��U5s%����'6@�Eb��>�J�a�L����'��K���B�I�B^h���'�I0c�Վy���A#H�A�x�x�',dtQU@H�dP�hى1��m����Q�IXH�"�9�'N�B��D*ݵ2"�T�t�h����Id�D��T�wNp�9v�X �E�Ɂ>ަPx���"}h�!s���ԥOx�a[w�p�)���'�v��Ь�*+ʢ�q�[�k�8t9�y��Z�o�(Ty�n�IMZ���$j�4�0_>� ��b�AW�\8l@�����&�'��1�̇7����#x��EM?+>��JU/C��_�U\�����H.T�0@!�8 ��O�d0%Z?ט�R)�ѵj�9�(ɹ6�^�F@�B��	��U��G�U<�� ��P�v����D�o���Ac�,`����i�~��i�(�~��g4 {��kF.�����r<0�6K̨�0=�W�
��}ۥf�#P��Y��c�w�&�cG��mf0��`׀}��a9a`�
dLC�j3I�ay���i2Q*�+7m@䵪�l�*��'H���l�(ј\�B(�2:�q� HF�:6����7��裔dԒXY��9!��4U�P�80A�\(<��P�CN����Ԍ��9��zd䁨N���
�I՘:B����H�#�������|�%���ۂ�͚HV��
,V.��p����!�*NH�1�J;��)���O��Qf�M+�0�������1��(FX�q7K9Xs�(�ř�$Ɔ�<`�ѐ1��z���`�%LOx��EN�v�dpR*�v�|#FN�C��؃qc?=ۘ]���$@9�x����5��'�ax�̇-����z��p�L}�<)��q�+��Z�6���)��h4�t��&f>D+�iڬC�(���d��L�m�QZl�����x�A@��%'Һr�� z����9
�BpgO�4� �)���W�ji:�Y; ?�$J�ø������yW�V�l#�4��g�j��X���yB'ݯO5�m���dȲ0�W�a<Bݻַ��٣���]:<��o �07.�j2-��x��%�2?y� 
4�:d�p��u�(I���z��D�Q�ǚ$�y�
ͻF���N]�M ������.�a�CZ!:l���*��1�:����6e�ӭ@R�)�冞W4T�&��+�햾�T��`�F:� ->�Ӭw��,��Տk����K���VC�I�6�� (U2Q���'�gF�bTa�N R$��p�8bun4�|��U�J��6�HWkX��$��!�R��x%j�YҠ�!o��(�2��G<)�i�!�<QrF��6&3O��1/;&� hHq�C�~P�y�'l����)ՙO��@��A 6�j͑4Ã���?:�Ԉ5d8	�<C�I ?֊��K�.V���ː�[}�O�9RC�{7�Y	��J3`pH���:�)U7n��c�]�4Ti�OmV�C�ɗ!5*<�f"��+y.A� �]t|V��-��踖���M�v��n���$ '/i �C&��Er�L�A���7<!�DY6"�����瓴P�P���kԠ:)�d!��~���AJ/�RȆ�	���K I��FYnD�&�~���N�l�"yK��+�(�� GI�
��L0aC�<K;�!�N�fO�4�Tb�d�S��?1sǌ0�2�#�&O�IB��z��T̓	���x��4s��	�u"3ʧ{�(�DN\8,Hv�91D�- u� dĄ��l7�O�p���
8�\Y��[��,�s/=a��7ƅ��~�mɼ��O-����g?Q��<x���y��sJL�F�E�<Q��ԀpC��q��� { �-R8P��Ġ0���s���@� �Q ��?��'#�<%���G�?*DjE��A�%��	._y~���	[�D{��I���C�>/�tJ��ñ&��%�i�H�����_��y�D�X�@m�Cjգ3�|Sc�?���Ċ���(�:?�|����M���d!F +j>0I`��~ݪɘ�D��y���4�֨��Ƀ^Ɲ;�fڠC�A��E
�eD=��m̙�H4L�O���UN$�g?Q�ڍHΪ�"�`�� 'D��#�N<Q��-P���#��ch�(�GD�ި����O�"�:��2<�D����?���ޟ�d��χ��QpҠ�`�n�[��'�Dt�����F�X�r�Κ5�2�۳@ǅo�r�k .ʮF)�D��F��?�b%�[}R.Z/P���[��2�|��Y�b:i�l@7CN����$��$Ƞ.��) �	J�8�Q�Pm�J?�	�dv�KeN��44�3-3AYzQ�EnW�f4ȉE�'2�A4�����K9�&�� (C;��>��w-���2�ę��!q���Z �DJ�^pY�j\�����gL�h����r��$.�hq��#��O�`ֆڥj�I����"O���!
9o�:��"Ł
���1A'=0.�⟄���92^�tx�M�!Y�(LAg�>}�I�T���f��)#o�t�ai�<��D��w'��;�E��s�`PG*�dEQ��b`�˄8@�`���X@�F��M��A�U�6Š�5��Q�&0ZM<Q���W� �fcG&;0�ѷ#O�~�[��|�FX;_t��Vχ=6��T�3k�s섒O�t��k'�ėv!����eOA�]^�h�T6O��(��#أm��z���e���
�`� E�~U���؋[s�ѣq��)A��fI�9_B�'���b�O^ݘg����Mo�̦);�CؑW
t뵡��/���"�f��;����{���=KFXMS��H�M�]�ѧ��)< ��)Κ=~8(y�'ٶG�X��'����썿$[�`qN�D�2t���$N�s�|�I�F�,\���%�
=f�9s�G�T������*�b��ף	�tR�oоQ�vU�"J+/�p<ؕ�[}�	�S�? <)�#�:C�PАN�i1 ��#�OxyVė��ZP#�&w�h�W��o����v�����M�eZ�x�募k�"�h%�!m�������]5�kǦ�,��O���b��vv��s��"2�Ƀa@�
80ZpAŝH�6�RV;0Z�����U��86�%YV+n���1�ϦJ�'�Bلd<�!�)�^�d��.O�x�0� �$Tz�NK'���R2��?(h20� m�����$@S��$�	ڦ!s��˩m̨I 0m�h�"��e�O��<�C'
%vG��2�b�5Y"!�f ���Q`sl_��">��k@& ��I(d�I�um�vMl���Ú=�JŃFN�W6�k���O:�ۗ��?O��OI�T�ʡL�((�C�]�z�\4x�d��GP<F�t@J�b��Ib�hخU�%s�CNt��T����v���SMO��C��_u8�\�C
�
Dﴙk�
.��\�i÷<�p��>��O���b�H˺�qv)\�IW⑀���t���p6&�0 XD��!R~,�0�`��B��F��R�Ӄ/J�h̓*l�)�ɝ�jU><��̛�pu`��Ʈ��>��$��r`> k��U�Ml�Y(p�;D�$A����Zs�Y:b4����LD2T��*�授uך�!F�	JD�>%�̩�,�]�^���m�����/D��:� 3�ٹD��.o�	{�
,D��0�O1%\��`q#�-�l�P�E6D���#)�6$,�9��O��1Dpd�2�7D�L��o�l8"�ȃDܙ
d��3a5D� k�Ǝ7X�)�	ۚ=W*4��&D����a5�f��䋗SU<S�7D�@Y&"�`mJ1;ǉ�#4>T�8D�ԋ��� ��{�ʗ�^� ��m4D�����!m��Y�I�j����?D���À�#F4s���;�����->D��+"&	J3<�EӬof���B0D�<�O�x�LI� *�g:��Y�.D���#ĿS 4!�ņ�/]�ij�+D�X�u�G��%�UA� A͆e�)D����H֒>�d���V(Pup�i;D��HCB�R���	A�
��"-*E�-D�tz1�>g|�92�I�j��|;�j+D��a�j
w��zq���u��16
*D��	�D�_�8��U�p@zHg�=D�H�0����K��"Z�Vx��c0D��1��,z��a��@ ������/D� ����i�*`�� <��T�-D���gd��x�t��bŖ�.�t�P�+=D�H�j�ph6(B&�T�;>`�ᇇ;D�p��D�s�j�J��� �"���H:D�pb�jA(zrV4�a�لA��BP4D�<P��Y�`�8�c]�]3��@�<D�`��&S�S��k��(K�~X��5D�(�b#0j�jq(c ݪi�1���4D��C�d�@1��Z8
{Nq�tD=D��{b �$ݕ&�bX��8 l��yBaE"x�b��:&���yҍ�m*�USD��4��Q�N��y�C�'-�qj%�[�0�^�uo��y�D� w�����{*�d1�ȃ�y�a�9h2e��C�^ڨ�餥@��y⊜�]K&���#��jslXX*Y�y���"�:����	.4sdPʰ,���yR�ɥH�jD�Ꙕ:�l����Y��yBȽQ6�1�&$���xG˃�yR��+*AjA����&�<i�&��(�y�߯I��<#f#a{6nH.�y�e��/Y<��,]�����@P��yb 1_�ŀ�$M�$��!9/	��y��V��� ���]�|���+��y̓�~ ��iǗ��Q���y2�D
r|p�R��qC6$�aͷ�y�L.%��S��)us��c�_��y
� `p��"��m`8�bTMZ�"��|Zu"O$e/�qy�]��������"O���C3_ ��O�7U3x0�"O��YG�˼o5ZT�a�|1Ptӳ"O�sA�V��ru�!C�)b�"O-qB4���h��
��"Ol�Z'l�7c�8�H�KI"��� "O��������Pụ�L�$��;�"O�����9*���)�/��u.����"O�!��$_u�H����	.L��s"O�<R��5��`&�F+���aw"OB}z��՚&�r9Г��z���+�"OV�"�V+n�{����l��a�Q"O� �C&���yb,מJ�X9��"O����ű\�HqZ���Wˎ�h�"O1����nk������� `���"O汪6�Ɵ(B����%:�f�k2"O���֋�!��l1%E����@�"Of��QQ)?~�Z�d_/c��d�1"O�	�EHQX �����I��|i�"O��i�D�����r焸<f6!�0"O�`[儉���� T�S_�E��"O�e�JJ��D40�ٯ`E��ʦ"O. �B	��qt��T��87|$�7"O�5�A�Pd����;��&"OT���a�^ז��N���P�"�"O��H�V�T#.������X��DK�"O�X1�EB�vľ�a�kկJ�:h�"O�(q&ąUK�!Ã%\�]A�"O�Q�蟨1h����ML�EN�E�R"O�� �v%���M��(�$Bt"O����ϝj���Ѐ"։zq*���"O�����b���C2�Ţϲ���"O"e��ܦ5UxD�A�
�~��"O�y�A�F�<�f�QR���q��Ę�"OJ,�6�$g�@��0�^O�N%��"OZ��G�7Ű [0C��T`{�"O֭@i�d����O�z�-�!��Ϲz�)�u�]"9�5�&I�H�!�$̎B�v�à'�Zbx�;�Q� �!�;
(]��.�5.+�p���o~!��U	T ����7)��Z6`W!�D� �d��!�&N��d����
=!��	�D0�A!Z-^ނPp�B��d!�י$%5Kr,K8˂�ѐ���7!�P�~H,���9%�f�چ`	J!������#ݒ.ĶUJC!ǳ|�!�Dۋb#�ix��$K���q�٠C�!��%*wxh�qg	�G҄q�"�&tA!��e�C�Ӥ:��AB%J;!��P�r�2�e��a L�q���8=V!�D��, �j��:( ��2��G�G!򄍨AA���&t�$�	��		!���;>���C	 �{}���N�n�!��6nCj���i�'{ iC�MF;(�!�$V�uk��8$ N���(��Y�$��I\����$H��
>
P�@;�B.{f�@AC"Oځ��$�*�Ruk�'@fXA�"OX� ��I2K��)�) �T�>H��"OT�HN�T�,0"�R�iղ%Z6"OX�y��Ѝр�ґ�׺n� <�"Oƌ;��?>XE��A��c�""O�`Q\8��"�
b�PxD�,Km!�d6s�x��A֮�����ǐ�!�� �I�CS@�IK�yZ)��I���vl(�'#.ؘ�) i�PS�`۾^u�Q�ȓe~� ��Gԡ�^9CRH��Wkv�ҵ�i 0�O>y���O�����L� ��ef�=9�^�kw"On�Cs"S;z1�!"Gř�5�:`!��'P2u���p>�g����܋�;-� Ep��w�<��M�SvP0��D�]�.��/Zo�<�F�ΰ_
ԥ6�N�F}�a��E�<Q���1We6l���	��P���A�<ѡbJ6\�wE^
�X̓���U�<W�GG�]��?q0���'Jv�<�6������kQ��8@7��R�r�<��R�B��ej²�d�u��i�<�%	$n}�AS
Y0|�l�ǆ�]�<�f��m@A�I/��E���V�<A"+]0#ڠXq�a�ɺ���O�<����EzFxѳk��`���Y���J���0=�l��fڜMqMLM,�P@��$T����T�o�
y��� �q�'�Fh< ��'`�6�:sH�n;p҅Q{�<��oÐE�M)�N	xHA�c�x�<�ҧڜo7�x��i���X�i���p�<�&�ԦJsH�0si�-���i�qH<q�)2v�6��ec�"�J�q%K��yQ!�V�B�r��c�)XR� 8�i��F!�#�ݺuN��3"��h
;0&!�T[��q�G4�@��FǾ,y!򤚛#`l�D�S/'�Θ"d`Q�H{!��%cFah��M'*�x���{!��.iWZ��iҶ>�^�[�.��q!�D_?j@n�ZpǑ��&	ao�:v!�d�y}:�S�?P��)ca-�#q!��ʟ)���+��{��E�EM��!�D]�7��Y�k�$f~��X��j�!��ɡ-�T��2bZ�ZڼѰ��f�!�d^7�hcl_�3ʹ���X�!�	
���s�5�H8ۃ�S�}�qOf�=%?��+E�!���ꋁd�L��UN+D��X�CL�1(N�(�bH�G�ҸB�K-D�l@�A�"f���a���}���k,D��a lC?}�H@�A�M�9BPv�(D�@ �Eƴ,ǲ�1��dh���<D����l*a��U1ǊZD�z�"=D����K �:�ʱ&�� D=�[0&<D�P��T-��`
�� ���bv��y�
��wir�Qs��Pn��!달�yB�A-eH���C�����`Y�ye֋=��y`�
	�$�n�i�.� �y"�!<v��M�M{�4��/��y�X/i��7GO�K5H�(6IK��y�H�ĥq��I���elٶ�y�˓(��0�$X� Ⱥa�Ƶ�yA��@�@���cC�P� )����yҀ�+u�ba韢@+1�7�N��yr�^�a��R���5=��m��� 7�y�k>+� �CBN�Κ"����y�c���U� )�{��預�9�yϋ �N��C��|l���K��y"�H>+ǂ��,Jr��S�%-�yB��wh�u�g�/F#���S�p=��}�A"���ҩ'=a�5%aZ��y�	���^m�ej_j�,�Ȅ����y��~T&�J�!�'3���C���yRI�7��EV��1@�\�K$Jׯ�y
� �q��N\�H^戁GU�oD�P&"OTEPd퐡_��*�뚇�d`'"Ox�ZAf�'0Mkfd Y���"OH5����9Z/�T�MJ�=��#"O�f`X�+x:�x֫_�d�lp%"Ox	�U�L|$z9GꙄ�(ؑ"O�u����o9�@��ܷ%+re�"OP5Q��N,P�:���r܀u"O*):�I��Uȱc&$h���"O	��Fגl�꽃#C�%���U"OryC�O������hU���"O.�!�O� .ʥ�w(X(~Kz��"O,��1!B��a(�(H,�U"O�ĳ� ��X���p%^�%p|�"O��x�e׉�� "��Z%��"Ot��ʆ	[ыTA�y��G"O�8�OA��([�MR.A��u�"O^ e��6\!��M��v�V���"O@�8f �|�Xx��B�ya܍J"O���fN��~� ��f��PDb`"O1��\�^�;����/�4��"O���P�Ԙ[V��ԉZ�D��a1�"O"�['b��rbXI�g��4�"O�	OB�K���6��8A<D�b"O�4a5'Y-LҬq��7�6D0�"O�cO$�p���!XӘ���"OB�cT��+ J��[7����y(�"O<mh�����&��ǘl��`)2"O� �ҎN��r�ВJ�4A��\�c"Oly�#�2K��@�/�?�x`:�"O��"�@�1�TY�qER%%��8�"O�TX�!П�Č;Rg�d��!�"O@d�FJ<�H}�P���:�t���"Ot��%ʚ`�|`t�ȳ�����"OF(�ł����� &�D�R�"O(}��"4%�q9��_�0pؕy "O��0!��%��%I�P?}]r�p�"OX�j򆈊|HH����.��!"Of�����,-be��&��(��"O�2׈4����U�%f��Y��"O������ ��AEKۗ{!"h*q"O� ��ᛜ2�p��5�� ��Z�"O��cV!"�ƽ�&O�W��|�"O��  �**�R"�2�L=z�"O��+C��X��&�A���"O^$;�;Rxx������C�>8 "O�R��SB�|`�"�T��5Ӧ"O��P�EI�) ��%�U���T"O~�C��M;rr�=�BMćq	�pГ"OJ �*A�;lx@��>�=��9��x$L�Ð�S.0��j@�de�مȓU��!q��X���  8`*H��{r��W��-�.���d�r%��΀İ����Z�2K�Uj��ȓE�PX�V��SxuҶ���w���ȓX���R`G\�z�l��毞/}��1��kVp�Ո�ₔ����]u�=��S�^]����<�� `�(��8�N��ȓ)��;� <p�ݣ��ȇF�hm��+t��9��P�w�)!'a\�)����ȓ
��xh�J�d|� %���>"��� ���6O��q����I�ȓNJ�m��U%�B40�JJ=\����ȓ=��MS��[�T���:m�`��S�? �t	�e�+o��S�eO�2�ш#"O:x{ԥ��]a,�ؖ��z���"O���Q!ӗv�hT��.�B�f��"Op��Dŷ�\(Q��FI��,��"O� �OE$?��@s�ڶ6��Q�"O|l���b$6�H�k�
{B8�t"Ox����R6Y� �����<*_|u�W"O�Yq¨�"LVm��K^0���`"O�5vi� A��<1�
K����	�"Od1��
bY� ���8 ��"O�[QI�*�%it�[�VGfȸ�"O�c��'�H 3��#.�q9�"O�̓2�-g�!b�K<0 ��F"O�	��F;hx�s��l~�J�"O�Љ�o��"��I[�Ꮯ ��r�"O�t3�j�`���Q/+���P�"O@�ӈ��G�� 
u.#W��1�"Oܵ�$ �P�	(� g�L`ؠ"O���΃!%��i#A�Q}<�d"O��b��A�6?��kV5Jp�0X�"O��S�	�Y-���d�bp]�s"O�d8�@[ 5�,Tˣ�P)TB�s"O楐�k��cd��P,��
1�HS�"O*����ˆQ(@(P,ƀnV,�r"On�+$0p:l����H��$�"O��5�M'�px�D(��0"O��C`L�2�zG[)����"O�%9�)綸�Ak��v����"Oe�!�YD��I/q��;�"O�E[ c:; ���Ѳ0���"O`�����Q��2�Gʌj��"O\�H!͋���@Hǈ�6��9"O�1 �߶rN�٠��)�i1"O|�F_���`b��)uZ��"O���Cl�/ /L�4�<[�"t;F"O482& 0|�f$�戝5|9\�(S"Om���}�����H9i5DyRv"Od�R@�@�Nq�X�g�0d#�5"O�Х���%��CW��$.�,��"O�q6��N����F�1nR��3"O��'#N�7O8�!ģ�T�$Y�f"Ozʆ�CK��=BU����"O~�#/["��كQ�P� ���b"O`$%�O,��(�&C�@�p%�b"OY+Q��B�:���[�	��E!�"O&�J�!)"��ц���U����"O�x)�C��8�z�+ʖp^fu��"Orؑ��D�)�
����ƞoP����"O���`ҝ{^��3#L^*/�l]c�"O��Be6V|���"
;�Z=��"Ot��"0����)�j�Lx�"O���WD����Pibʛ�yU,)�"O�Yj7D�#Jb]1�盭+�F8�"O�-Z�ȫn�z��6k��e�P"Op530��*CM���R�,S+u�"O�e;!�Y�i1t�i�'�
P����0"O�uztO�<Q���;|}�"O�=� V�Z�88�&ްu�^�
"O���l^%����FÈ�*�"O0m;/�OV��aW��)&N�C""O:���h�2�x�{b��-PR�3�"O@e���D�Q��u�� �B @�R�"O4c�ّI:,��o�=�u!1"O�YKp$c>v�Tָ<����"O� ,��'��}�� �L����"O(��fĝ� S� �M�)�QD"O��p@��0!r�� KA�n�Е[�"O�i�4FL�����ۏw��T��"Oj� �4�\�Q+Mm@T!�4"O�\0��ݹ�r�s�̘_#�xYU"Of���ٛS�����̈́;
d�"O���0�V�x�U��O�n��#"O�2�e�8N߲�s�W����'�ek��~* �*Da�:�[�'�vUq҈�Yz�;�j�(���'�\U!$�;�@Z�l_13׀$�'��)�c�6)����ݹ(�荐�'9��MM�1% �3�C��%?�u�
�'�h=Z�U�Q���#���z���	�'��+�Ɔ%$5���B	�}�	�'�{bf�8��pYԊ0L�@Y	�'�4q�(��Y��S�X�<~��	�'��5�@�(�&8� 若3d��'����%�bG���L�%3f<��':�R��١/v�B�� 3fr�'{�@�ǡ�:o, �B�Է����'���� @ <M��#�s��`�'|X��(?\�x�#t��u(q��'�h�tl�O^"D �
;k���
�'od�r"!NwH�S��z�ȸ�'�)�P@��	KaG#l�C�'�ȭ�A��'��|��CkVd ��'�0t��CN/Bv�	���iF:q��'$ȩ��
�"c�e���]�BT��',���IS6D��A�'�V*�eS�'��@5���C{zt#WȘ�a�x���'P\\0�R^�ȈsƊα�P�' ��C�F2t�������*��'}���JZ6���Qŏ�	�x	��'�L��5���j�T	���	Hx<
�'��)�C�I��M��a�<T�rU�	�'7�Dxbד3f�1 ����@�2	�'�����\DT�0�J]�
,��'˶��#�:6�L )c��V!�j�'w����O�1V�A���P&*��'�Q:A�(?�P����@�,�'A�lB�F���� �7�&xH>Q,O��?a�I�<�`�I�4�Bs��A8�i� ��z�<-�8��-�-��#�#�t�C剱uP��趤H;J*l� eÒ8?
ԣ=�q�4��*��p�x���̝p�"���2��Y�rHN6�d@�R��T����R��0SC��_��d*��G����#n��ce�V
�HR5�ǌO�م�	A~�剐@���I
-;͘䢣)�	�y��bW~����p8e�"�J(�y�-[!��zr`A�w�x�9r�Ұ�yҋ#ur\� �F�q�e�$(�2�y�ԅ&�. �IЄ|U�������y�jE?_9 -tB�7 ��\aT*C��y�j!$8�q�@H�q�px��(�7�y��Z.[��21�So3Jti4�	.��d*�O�Ūe�1N6n؃�
�B����"O��F�ϕ$��U�s ��l.��A0"O��GO�	\�	�	�<5F�pU"O��R��Ш^�%qPB�*��Aye"O��؇�.y8�l$�*�J���"O~����+jO<�
d�S6����2�'��)� �T0���7In*�h$.�P�&X�S�h���\�?�}��J�<�ڢh�h��%;T�K�<�����B��1A�vsg�I�<A��ԏN�¼�1A]5^ �r��o�<1��ޱNT6��!Η�42��TG�U�<�1�U���@['S�71�5!DQ�<�ф�K�C+��;����c+Bwx��'axM"��L���{�Ӳ1ahl��'���6�L*?h�Y����-:��+	��'�2�z&��)T��H.@{0�	�'���&�f%��ڤ��ʍ��'�2H�W�ٷ_�d��TC��cB��	�'�.$C�n��`1՞WĂ���'�ԩ����apuB��ǝ{'�e��'~.u� �� �L3�,�X��g�<I�.Ƹ:�}���1ԅ/���?9
ӓD2�[CN�.mTl@�ՠj�ņ�Q�z	b2i[:�уn���ȓz�vЛ�(x�H��It���ȓ5,���E�p���
H���9��̲�'�11�cCav��"���C�6F�0��I5�X���V��B@��OL&���*mQ�ȓz/F�jӢ�<�%$\0@�}�ȓ<�<�ه�uX� ����|��}�ȓJG�P�&�
�yb]�w�֎"�*��|��j�&��0j Hs��S��]��_��n�n�$���k�;�x�ȓ(���X�b�$8��cv��D@хȓE���W�F�<8�YV!����Ņ�z֮٢W��#6�����9L�r$�'�a~�IIa�Ԝ�R��w��E K��yB	==�%P�� �n(x1c�A#�y�� ����m�c��xw�^�y�W 2���"/7]�j���/��$,�S�O��1Jp�!>&dZ�lW�Zex͢�'*���Χ;���tꕵ)����'�.�i�P���F�:3�0ljT�|2�'��\;���v�J�BV/K0o�t�"�'������>P� 	�E*48�d�i
�'��X8NU�H�>Y�R�;45�j�'�D)���+[.e��@ͼ/�0�R�'M�@�Zi��)��#P�0���'D �J<)��@��[�(1��'F�}��c� z
9�FA�y��j�'8 K�,�!o�U�0�@%b
���'D��׮
�@΂��$h�[@�a��'�bi0Aǎ(|��z��^]�&a��'���qىy��j���OA9�'A����Sk� D˺t}z��'��·o��i�f�K�K6hYʸh�'�t��Ud��3Q�Q��hG�W��|h
�'�0�����oL~(K���J44 y�'F��E-N]G4�I�I� ��q�'�Ft���]s9�<�t�Y9\�b�'�>�q��U 8�첓 S������'��]�R��7f��0�V� �����'z�h�J�|�0J�e�X��"O�\�c�B8U�t�%�8f"����"Ob}Fx���Ý<H�apb�A(!�D��^T���؈	�ő�cS�W"!�O����!WW��eTÉ I!�Deh��j�C�j�8���I%H��	yyB�|ʟ�+�` 8q�G�-�0j�nV��x��S�? �i@�T>�̠�%m�� ���5"O��w�ʲAj=ë��재�5"O�U��%����B�&M�����"O않�*����%C�Ԇ&+����"O$�	�y�fD䈡r"O4����C0�z�Z�
��<�l(V�'���hy���{RfQ"�����M:MQqɠk>�y)��hV�Q���E�:D�&
�y©̦1^�� ��4��4w���y��ʠd�J(�s��)'r�K7�J��y��:��r�����$1�T�y� ԎU����VĀ��<*u��2�y�F]� ��֌���	Z/ȕ�?a���<�|�O$�rf��(K�@1����q�
�S�"O���#�Ҵ[2qC��;R�!�vO*�����( �ժ^�t(��t�9D���D���9S9�1�&cӀ�[�#D�|�'i�&�ʙ���Yj��yR�-;D��q�O��S^�xPDX���5B�L=D��ŏ��3��Ń�ռL@����Ox�8G��'���c%��!
mstOR0K���"�'�⡐�j?Q��i��NI'F�t�`
��y��
�7}� z��ϯc"`�3d'A4�y⦖"7LZ�ral]��A�C�Ѥ�y�[�,T�|s���M̬�*FNŻ�y�d�z;L]{E�H,=�6P�f��9�y�e� ��8b���duܘ��"����/�S�OD=��e�t�\�e g ��
L>A���)Մ8�(ݪs&�*7�<�؁Y	F|ўT���1�r�!��ı��@jA"��˓�0?��|E�����a�M����]�<	��˭n��t�b��"T�� �c�VY�<�b�(=�,�C�ƙ�i����V�lx���IP�:�n�����d3�]I����|�ȓ`bB���HW�T�y�5g�s|�'��G{��ԥV�QE��ľ_&C#�ң�yr�ʎGc&1�1�����ò+̲�kM>��C�Y!So�B��ʡ IXX,��8t�1�J+"��
�"q&��IN�pKb ��^��l:DB�����?9���䟑2�xI#��T�3�)`h�?:!�$\�p���Y��|_
�6M	$����ݎ=�avH�ms��z��88Ȣ=ɉ��?����H�vhCt��9%�D" ',�	G��p9��)4n���<\̭��"8D�h��MׂJ6��S��E�f�RE8D��H�2p
5q�!������6������Ɉ�7%XD�l���+!��W�>�luZqf�B
���I�j��r�'�xLqt��0)�ֹ�06V9���'�!�D� N���c&�V�Y���%žr��'��'��đ)�����	�w�j��D�˕l B�(�<��I��fa6xHEɲO��B�	L��(���P��a�CG�,	v��#�nq�їo{���+P�"� \�Ɠ<3ލ�����{k���o�	9����'�x��&m�)/Wh��ѤK�>�5��'�B�x��^���U�@hF�7#b�s��d!��倄
X->�6иŪ��V�4-��"O��!Ҿ0�@Ʉ���5z�-��F!�DP�ND�`�Aݷ3Ӻ�	uBC
S!����=�#M�)-�,@��慰|"�O>����.�������m�1!��K���S��(�Ȝ���U�)B����,C�lp�5	Q"O� РrG��DbL�r0��KHb��"O�A#�v���@@G@jUf]� "O  ��D�L��<B����p�$"ON���9 ��P�	���F�7�'��DN�X��$��(J3�f���R ���d=�g?1�)�*�d�Yɞ�]�8!��GAy��'��OQ>Q�0�ҒRL�+��?W\4}b�O=D��uƕ�f:@*RʍXL(�b"K>D�P胎�uP̥Q!'�ҴAy�<D����ƍF]6`b�X�k6|���9D�\��5Ī�����Y�>�Z��<ɋ��S�!��`�c�y~��;"�Q��(C�	 �n���"���Aǋ� �
C�7�~Ԉ�
�)q�T#���5j��B�I�hA&��g+�6�&���ԑB��B�I7�`�Ə�3���b��S�A�JC䉇a�xlꅏY�t��X�Qo��2�C�I�|~�� h��2�Hȡ���M;�ʓ�?����#RM2���AH�T�s��߬B�	�^���0�OطvB�l	�)���C��#MFZ4x ͌$*��E��"L./'x���;�"]�
4��4<z��Z�~�C�I�\54-��E�%v� �Tf�-w!4B䉹/�,���\���)tN�9>@C�4�JX��CUF���棐d@4�O8���<��x���%n:�Y�p%V%{!��O.M���S�7S,�#Z�e^!�Dڛ!�V�	FCE:`�yS㕾UT�}R�����Ȗ2;|�a�'�F��)D��ڃd��t9� .�7s0�B�&D�TA�]����q��E�g�����l!D���T��*s�H+���.x�hi��!D�0R#�B�b@H���A>E�f��S�>D�\�S��+{������|�>���ǽ<����ӄ�m�g�Ѣa�8W
���C�I� }���#Om����=*���d?�S�Oۨͨt*�@���hA��'S�H�C"Oui���+��;#L=�~�2t"OT��AA�:�X �lжbʨ��*O�u�E�K	L�\��@ׁ"Ԛ��L>9���	��Y7�B�T�Al�ǉ�+"�!�D�{�y�A�S>t�`��d(R1v!�dH&򁻢C�#�u�(�?o��)�'�Ԥ �o;����ǘ�t9C
�'�t�sL�A4�u��8 `
�'�rӰ&���S��<tٜ�++O>��2�O(��C���*����n�;�"Ov���� 6x\�`��5-z�"Of	��`!y�D�4f(���"O�p'j����P���ƫ)@���'�ў"~�%��6�^7*��i�0��y"O�*I΅���3�����dɱ�y�b��n��Bq�ö*W4�qnؠ��'�az�)�
3��ZF�݇:���pЭ���yR��0 f½����8kI���yrb}qj]� � �>����A$ܞ�y�o��ky|��D�=�N�#.ѭ�y�S6cqf�J��،3���	�c��y�
~�}@�"�\ل�eO΁�y�n�<>��[�j��fԹ
�.���0>��߮0�蔺�fɩ-�h�c�K\Y�<IZ*c���1�[�>�*��U�<�'�D	7A���vI�!g�~A�c��Q�<q6��   -�5�HxeM�d�'a��  9#Aפu�D�!�X�>��"O�zPG		�T�,�b����"OҤQ�'RQ������w�N�I�"O�];�� s�gQ�u�
%��"O��`lܧD�&x3$�!;�
�R�"Ob��"W='���&D��0��"OV���
͒����;��cf"Oƽ�'ǡ"� �ٷG_΀(U"O����ɝ#��A�DmM���I	�"Oh�z�ǫ-�֘�G�����"OA#R��%y0 '�U�<���'"O�9�B =窕��$L1G�r���"OV�[B���)�*Զ
�`�YT"ORdᶧR������i�b��X"O�bs� DP�����
f^�8 �"O��#�ׄ��:r�P�lJ6���"O�mIC�J<aˮec�+�-/z�0�"OԱ�p%Q�1.�q��U2H&�'V�	�v�i�QAF������=V/~B�I�mm�E!2-�ʬq�D�fFB�I*O������3oy���R�][��B�	4+4��`���M�����
�k�B�ɕ,��UK��Y�<���Q�����B��J����5GU���4ˁ��lB�ɻ\[Fuۂ�<df���o���*��$"�ɯl�Z����MMn�H�m_�%C䉬Q��d�  X6jV�x� H�^�&C��T�9j�ʈ<
���!	��`��B�	��R�YT��U#�e��'�NEtC�I�s�|Rp�Ov� .]�g�,B�	�E0�p��H�j��Ԙ��*��B�I�?��q"!G�3<������0�C�"Vhye��:Z%tD�E�O�,��=AÓ{O�$A�':aط���W��H��[� ����Q�,�-�t��I��a��Te�Uې�H?z1hD3Q���4�2\�ȓQDN|�o�j�\�f�@�JT��)�n���"ء5���FP$|�8��� 0�	��sn��0�',�����Ҷ�I���Eb��6@ӟOԸ���q;�I(�Mk�́U6��ȓ�`�����kI���Fb��i�\�ȓf�\��iڿ$v`k�j�<~=$��ȓ&�<�3��L��8�7�S5L����ȓ'g�f��D�b�h��ٳ6�Y�ȓY�$���E�T�f1�#A�2z��P�ȓ@_M1��ӄJ�P�v�_�!Ͷ���$���)��^*���H@�_JNP��M��@�$��d��ꃏ�7!���\��{w�L+���a�
�5�Y��$�t-��bK.7#��P��VB\8��T.q���V�{�؃F%J�@kjQ�ȓ���Bd�;0�1 ��	53��X�	}����
9�@ɰZb>V��'T���J��y2��!K�['�R�X�j���yb�2���r���u��-(�n��yrۏJ8��4�'qwl0���&�yfU?��Tж[�L��&�P��y��
2z����X	��u �)?�y��$Sv4Y`g/麥K�L]��?1���S�BkS&f!ۦ"I�^���c�D�<��I��[ffr�Y�#�<!��׃�Z�b�?\8ijf��y�<Y7,�>"Ĵ��3�^�L*"�d��x�<� b��!ʎC�akV`	W�C1"O�[�c4>g���/
07Dpz�"O|-B��9�vn��!72�k�Y��F{��韢7#2���HN�&� `��O�|�!��Ɯ����`�G�^%Ȑ���!��]s6xl�����
�f�a��޿e!򤅚t�N��`��q��Hxr%�	#�!�dlo��U��?�^�锣K�E_!��4C"�����Y��Z�|!�d�VAd�T�ˉ,���jd�!�DZWq��`�%A�pA�N�"m!���rg�D*׭��vKF�1t�[ mM!�d['�i9�g�W/ �l�?G7!�d�.9�"�$O�Z*2�"��ث3!�$���z�[2�99,��:��ƥ�!�d�X�8@S��W "�\�b�H>!���?QH������,S�D�6�!�	)����$� O�"c��(Tl!�$�"k�X�-�b~p��cLF�x�!��)��aǓ>��I��F9KH!�D�%��Zo\�]�VXs��
*cM!��P�E/^lX�����5���(@!�	�H�qT��y��|�� �+xt!���)���I6f[+۔!����3{�!�di�R�Q�m�\U���&�ʤ�'"O��B׍w���CG\>g�TԺd"On�ń֬Q7�)H�刃r�z�"Ozy`�W7J~�|��D_g�P� �"O�h%.���~��C��kfLˇ"O2$��'T8�����hc~-q"O�%+H<�̡CV��v��"O��t��N��R����!P�"O.�S�X�Ȉ��
�7�H���"O-zSLؠ<��i�D�/44@p�"O�W�J9Ұ���N�8Y�"O4x�Q��(gWtd�#ȁ��ʕ�'"O<�SWoKi�v�酇��^�ف�'��>O��e�Ǭ$x�LRf�`�
�Q""O��D�6{(h�%�/=��ˑ"O��9�d�'L&M�@�C�em���"O,� ��ĜKe�`�Jq�Є �"O:]�"Õ�u�rb�f��	�B"O��R�i��掹��Uq��s"O2R�V����1`I2B���B�'jR:O�K��)e��5P�H�c$(<3"O%��矄fZ�H�@;F�ͫ�"O`,b3�U3K�
����c�:�"OH�Z%kE�<'N��4@Ҝ����"OP��dQ�� ��-t�8��@"OƐa4HQ*sט,*� �@���*�"O�� *��C}��yjDJ59�"O��y0"�gA<��jʯ}O
�3���e>��Cݱ''*I���D9f�� �.D��Z39_�l��e�ݥ /����-D�,���Ăs��J7���$����+D����ܲH�j�`Wƞ� �v�b
(D�S�D�%�
��ԍ�(�\���9D�P�e��#y�����c���@@D6D��eI*��e��e��UyX��)��O����3�$h8�$�q�T)�.N'4!�DY'H�Y��.I����̝J�!�Rt���Y⮘,CX�Ѐ��S�!�䅦:!� �U,X�!A*=�ө�g�!�������.�,F"(01�瀑N>!�� DyBd�P�f}QW&\�Z�"};��|2�)��Z����X�t�؁P����u��C�I�-�(��I�aa��piB�	LԐ�;��^��#E�X�B䉧@�zt�q,�0�P�r��Ճv�C�	�F��q���PL��KX~��C䉗0��$2���)Xcz�[Q�V�BvC�	.\����_	` |xA�g3<�C�I:g��i�EG���P8�Q���|��C�M�D;PKA�Y&6@��㍸?��B�	�f��`��+<s��@2�I�TB�I116*���D?]���eȧ{�B�Ihk��QA&��E��J��7�vB�	�����D�^�� Ä�x�C�ɟD�^<�4DN��9���|��C�I7^�f��&���,u�	��CSQ��C�	����0!
��3�3Đ�u�nC�I %1�U8#�K/�$%���*:lC�?8b|��!�?�4H2��M=.B�I"jz�7-K�m,��e���B�I�Y�|u���*�(�`�*�]vB䉝	�L� 6�*�����P��B�I�4T@�r�îy�J��cJ�M�B����,0b��
Lt�H�
B�B�I3S�8s�=,J���-�n�zB�	L����׶87(�q���H�B�I�8�
1J�nU�*�1U��$2��C�	�o�,i��G�?2�ū�D���C�>
���	t��v[@�����2c��B�I&1��Ap���@��A�0�	�O9�C䉆J���D�3%	�{�K�>��C�	)q�FVT�dP��f�>j^f�x�'^��)C'H'A� `��K�c�J�c�'.,�h���������Ҍ07l-�'(�Q���J����w�Ǣ)�1�	�'�f�K�_���2ئ�����hO?	c�e�5_��9Q�%.6(�H0FXB�<�4H��7B����n�C���S�~�<��È�5���)�%�	K�Yr��`�<��	�%�����L�=�,m���]�<�de�,��!(�m�8��@D XB�<�֏Y;�����_9f�@t�R|�<yS	�0 ����`���Cօ��$EC�<����l���ID~=�頤fGA�<� �V�p�ta���K�B1�'�{�<!0�_�d31�u��2���Qp�z�<��엧b�̩#" !)��9!��t�<�����)_�p ���$�AV�Bj�<aSKӗ!�R��KBN>b��4��A�<�A����9u/�b�P�W�~y2�)�'G���r�@ڳ<U�ؑ3�"z�i@�'��s�6i���	amH��k�'�DkS�O���$�B��fFz��
�'#nq��/ѕgL6���&@�(C�	"T�U��C�+��G-Y�Rk�B�ɕt_4���o �� 2e�`[�B��=y:�ҥ� %#��X@A�,i����k����פ))��j�^�4�@<D�\PC� <��k&��R+hh$�8D�
�D�Q5�#�V#J�U	:D��7!٣H ]Q�G��FNh����$D��s�G�(]t��ĥ1�@̃�o!D��z�,"&.hV�X��yu�9D���g�F�k�Z��ejӕH���x�c*D�� `���/D]�\Xx�E(�X,��"O����oQ���yZ`�^'-�|A�"O��вf�2m����E���r��"O�3��T�?e6�ɣE��w�h`{b"O����MP,���h�Ѯs��-SG"O<a('*L��:�>�ĕQ"OĴ`Ǡ�?yfTJ�hڌ<�<`�"O^�j1�,��� �č�(��]:p"Ol%��.!j�j�8��Y$(�dY�"O>�D�	�Ot�kܥ��pڡ�ȓ/%�@���	2T
Ԝ���ɴs�����.���GL�Jc��
G鐳	xن����'!H�Q�#7���
���p�<yΕ*yK|M�1��4Nư:3�j�<	���#m����(��걁b��f�<�V������q���bM!��Yc�<1 熓I*��r!�Ů�Zt�_�<�h�1�|eAՋ��t��e3A��s�<y��R����F�@�`V�Kr�<quMS5M�0��)˲z"��@�c�<���!~��7 \,Ql{���[�<���[�y/Jt �)Tz�$�p�X�<a5�X�l�h��	R?��r�`�W�<���O5$�ȧ�P�y`���A�S�<���˨v�cAF�>��J���t�<���F�W��yS��^�E`�]p�<9���6@���30,q�Y��.l�<T��7$Ә9p!R���%3��f�<Qt��R�>����۪�j���2D�l��.�.��y�􌛱L�6#P	/D���w�  s�]!$%�A^Liku,"D��0BN	�AJ�giұ
��Ȃ�+D��u��A�(^�C��(2�?D�(�r�:[N�0��ݘ���(�)D���O$hu:);�+G�|(��'D��s�F�f��T��目<ߘ����%D��৤�$G 
D;Tn"y��ZA�"D� y"ő�a��s��#B[|���;D��Z���<d��X�l1�;D���R+���)�U���q�8D�P�#�ąA����M:�����7D��CQ%
�q[�^�Bz`5ʡ4D�L��ÿQt�9�qȔ9�(��E�0D����.X�3��!�4S��!�EN0D��𐨉*�����O�Kg��� a(D�����תu���[e掸	|t���a+D����U5b53�.̭{�0Xu�'D�@��NC&Ը鶇K��phʥ'*D�p�C�Ğ~㴙�w�݂8RDJ!N(<Op#<9�皒h�Vh��O1YZ<0u��P�<�AΏ�@9��z�/72����#�K�<��\�{���	�&�n5���\J�<��8&�����N���l�'��m�<�ǅ�Z&���2)	�y��j�<�c�PHU���Ɗ<�&-���A�<9- {������4>0-��Dx�t�	l��l$*�
��i�Ժ$�޻V��ȓ �^Y�T�ƾ)�Q���� �X�ȓ7.$K �$p�u�,��;B�I��pa5�����G��BN�C�I��cW��V!E(%ˈ9:��C䉌.f��T�[�e@��aĉ�HښC�Ɉ#y"��0	\z#�fƺP�^C�ɛj{" ��hn�]X �<Up8C�)� DÆ�������3t���{#"O�Zn�;��aS�
N�<n�"Oz�cB��+՜"c�ͧ4+���T"O�	
����<	Y�GC ]!���&"O������r�@T�F�K��1�"O�6�߼5�֘�`��80e���P"O�p	a���VN�a0e�	/�PZ�"O���#��@��p�Â�)��̉�"Opt���'"��
�+�9�%B"O$�)�=`":�@t+\!+��B�"O$h+�K�BM�Yа`Ә��"O(��⭀7��=����}�Z��"O��r�t.�aӄɎ3�� "Ox !��:W�\�V*ܰ�d\٢"O�4y��]2l���"�"�
d�`�e"O2<�qj_�"v�c��G�)[��v"Oz��c�6�m:#�<qP��C�"O��yR��I��7a�,"m�є"OV1q� ^�n���%�K�8y2���"O�h+�bӄyH���l��m�(�"O\�j϶laP�tIݧ} � ��"O�4�!��'�00�T)�a �qC"O]y��Y"x f�� ��"�"O���d'؁}60L�ժ�8'�`�"O�q��W(2~��;cd��� �"OT��/���P	$��'�l��"OE��C�n)�d"r��<@>`�20�|��)�ӣG�~�(�#� p�4���=3YC�ɼ;V.AC��B}�2�X DS%^CC�ɴh�А�7,O4����
�!�B�	�32�h��C&����A��o�B�I��8]q���l\��f"�|RDB�	7���Y��H�.@k�@#%�|B�	�bs�y�¤�G8C�	�"=�p�3)N��2���/g�B�"nz�;�bQ W�V5s �ыo4ZB䉔2d��U�Dnl#eGK�/*8B�\��]����>��AK5`�Vj,B�I�b���ƹ5I��#��8�<C�I4p����e�k�	����x(C�I%'��;�������-`QNC�Icݚ51.K�f�`���
��
B�[́*���;/�̩��ۻ~��C�	�CMؖ΅���D!#nL89'�C�I"{�|�7�
&$U���3�J2�B�ɲ����H�:q��)�W&*�zB�Id?�M��/
����1A�B�$��IQ��1��	�C���
�BD!X��2r� `5�C�I�8�Z�$h�/4g��{��Y��C��6�B�
��]>ɼ Y#���cZ^B䉆;�DI�T/P�=���d&
q�B�	*�B��rJԲb̦�04�@|�C䉦r�����jK �@��1�]Y��B�	�P�B���"g�-�Oƴ�B䉰o�T��dē"�$��6����C��7J�� �V�C���F��(?|B�	�N�H�X��
)��@��@:8&�C�ɛ	�")���1v���j��f'~B� ��@y�@�Mg��"��Q-Y�VB��!,��A�ч��ԑzf���/@RB�	,N��eb5*C���䃀��#%Z�C�	z���a7��d���R4*��C�I+:)�����M�qXtЀ���g��B�)� @�ҐH2L�\(T�ʃi�5�c"O�9p-���(�4�ׄP��"�"O�Y+u�ʒ`���fR�~U�t��"OQ�u+�H��1���r+8|�"O���c)�#K.�Btk��M�����"O������O��(B�]���"O
���T�,��T.w��a�u"Om����'Đ21�
�2��k�"O𱂑�Ȧ��,�w�?T��ћ�"Op} ����|�I"��n����"O��@�2w���՝e�A"OpD�@o�plX���dɕp>�QV"O�*��. ����B�!Z9��c"O�R�g��Z�zUK���,V��"O��!��ҷ:8`�zBOސ�&��E"O��c�M��14|��q�� �H! �"O>��i\R~��Y��H6�� "O�:�ˈ$*}vX�)�9��"O�ę�`�,H90�h�'C�g��ܰ"OR�:Ej���caċ�l�4 q"O"�����1D�l<�@AF�F�B�u"O������*^���Ê�Q�v��p"O�i`�Ȋ������k�.���9�"O(��T醜1��$Z4h�(+����"Oy�O
8����2n�
=���"O��aU�R�e`�ȣLӶ\��څ"Of�:vO�����+�:EڍpA"O�4(*ՈTb��k��"l�8İt*Or�)t�*a�9���Z�lz�'�Ȱj�:�x\Gd_&�}��'N����Ն��M��-�A���`�'h�8�l�b������3�Z�S�'�\TC�.�����yr��2t4,j�'�l,b%۲�T�9Q�Z,2^L�
�'~bݛU���Y��0/r�	�'P�H�A�� �F`	���8,Y���'���c4+��>{PL�`�M�q�Y 	�'E�P8��@�ц�3$�c�<h�'��`�&�z��Mֆ�')�(��'��	s�3.�J���'̝p�'~�M�ⅈ}�rM�1oJ7#,���'�<� 䔞|�x�!���N�Q�'b��	#�n��q@!��N���!�'&
��I��z@.�A��4L�-��'�x�1`G# �,�i2$��y��(�	�'j��U!��6��`(���aް��'�vy���*� �#"��^k }�'�8l2�3�~u��S�g"�P�'�@=A!��<u<x�sf�_!X$¹��':�M�d+\�+�L�i�o
;ߚ��'�� �ѧ�+`~x0�u���6�L��'�n�R�
>`��˅���&�R%�'��x�@h�u�R��,,!e�c�'>�,��B�J[�$ъ�D��Q��'�H�`�?���h����>�A�'횩s�A o�����˞ o$YX�'D0\��-�Nq���ƧG� �����'?\)F��dD�4/.Ά���'yp���N�z�m
�r$���'��E�#ρ���C��Y�W� �'z&(h@���'��Y��.��P��l��'Б+�g�1q����"P� �	�'�E��f_	q�҉�iʓ�ܩ�'��s����a�'��I0����� d�+��E�Y��|+�ق2�eC�"OH���'y=�UӡaȃB��a�1"O�H`^_��с���lǂ���"Op�c D� ʢ��"$�M�f��4"O:œU1h azU,B?�V�Z�"O�@6O�#�*t��Jd��K�"O��ö*L/'����3$�Y��"O@%��\�\�"�(�����q�"O���G�8� $�j]�]����D"O�e��&L._��Mc4�H;8r��E"Oʈr����ޙ��������"O�1['U�bq�c����&��(�"O>!��A�c��m�dC�u.�0#�"Ol��a�L�Q"� H&m�9A���{G"O���2 K�U1�ِ�⌑���zB"O
��_>�ܨ+u⛴vfAp"O�M3 ��re~���F�7UA��³"O^�# C�PچQs��3m&~1�"O��[E�[�0�2�I����0����"O�(�Cիz�2x���}I�"OR8㍝x�$�C̀�RL�A�e"O�e�� _�'Vb�a��y;���"OfI�e��:��<��M�tR"O&���.ą3s��ƞd`TT��;D��*�8pj��H�7u����4D��9��Ҏ5��a�oO+=�y{�B3D����$Q�l0�[�"�!���12F>D�TI�+��@ޔ�CO��I�ܸHB�<D�\��~\^AX%Ce|���e.D����	(,uh����¡^�M�V-.D� õjG8�����J�u�h�pS�>D�d9V��5؄Y���	�/�J��/D��yf(��1&��!䊇�(ZA`��,D�`��D�2� ����h�:�6/%D�Cr��(yz�=��ݦ*��t #D���C4�BDa٘*��k$"D�,�3�XR^����v`����<D���6iM'_�)C4M%sKb��կ:D�x�w��P����m�T��d�7D�p�
H4.E=Q�J+7�<9�A5T�I�A  8��×��J��D{�"Oe�A�J'mg�B�I�rb�x��*O���#K�:l]�dD�<��ͫ�'���Q晈X$���d
}!�9�'��8���
�w>�9d�E8q ~�K�'��Yq��:��|����
b��}C�'J���
�=���e��D0�'�ܩ*tf��|����(�-rbe��'���0΅�jl����\q}�Y�'$�1Ц�s�@93�@˱z����	�'{Z`���	���7Ȋ�zI4�K�'�� ��	�&������݊C� ��'�N��TkX>C�@g�P�5Q~���' ��� �����ET�(8� K�'%r制���Ԝ���	��1	�'�$]Ӄ�A�,YtADr�T��'L�@`n�Lqɢ��	?����'�����,m��2.�>EXr�'&n�p#�Q;'�B9�m3'�Z���'�6`�v+L�-<j�K k�P,�L�'"�"�ڃ:�� �G�U�T0���'���& �24�M!��V�>��
�'M
s`�A�q�����%�쀉
�'�@{'�i����ث'�\[	��� �8!#��VD�J��cj���b"OH�R� B�57���	Du�"E1�"O&<i��تr�4]Rv��8Gy�s"O��
�Z)_���
��ǻ>F `��"O�t9Sou&l�Q�A���9f"O��R��]�^h��������0"O((D�� ��i�իX�t�-��"O2��6�;<p�9S�F�
LX "O����K9 k���@�F't}���"ORT����*M����P	��]P�g"O�	�Rj��qil�#GH��+F�e�"O�P灋#w
���C-��k8�pd"O@�:"l\�,����CFBDiڵ"O����B�a����f�?(@$��"Ox���LX�t5����̚PD*��0"O�4���K�`)`d³��O`4d�$"O�"�� <b�6��ZP�۵&!D��B��Y�p���*ՌN�juصI !D�h��ꖁj���cč"U�ʽi�?D��0��3h��ɑ��#���9tm*D��"�3CF|$����[u �S2�(D��@un����AFd��2�$dxw%;D�<���<x\�U��@�l���+&D���S��1������+�B(r׏%D�xz$"V�4�̽��I�w.���`$D��q���q�e;� ��=�bL�%E"D����re�B.�b��� 
 D���J���
����A�C)\�ZWl?D���#a�Lz쐫Kޙ�8���7D�<�`�č)閈S7�H'I�\��3D�ԩ�⃤0�F]��'
NPNŨ��O�=E��aI7�Xl��@їAU��z5���!򄞘V�,�ӀS��Rf�M�!�Ď�H�@Y�mPXFT};��P�!���&_�T`@��=8�p�S$� �!�d?|��E?5޼@��?o!�D�JQ>p��F�y,d�)��-rP!�I%�^���N��&yZ�J�.E!�V�1Ӯ5�Hݟ#���H#@5!�X*����F���] ����A�0!��ǊNj�Ă�R�` �Ee� ya��O������[�8����^= M:�"O���瓔Y�pY��"�D���"OĽXG�3)�ЭƱ$��I�"O�r�Ԉ53 Ĩ�
R�{oP��"O��	 ���E�C	]�`$�#E�'�Q��3@�����3����q��8!�<?e�'�~�<s�����T�b��Q�w�Is���OK��	���;Ɍ�۲���$��'N<p�!d�����H�B��q~���Ob��D{��/L��A$ץY�В�Ǿ��Ԇ��f^��\�f ����q�n�����39���	@�S��yR�9t8[�Ϸ@&����߆�y�"҃Y�0���	�5�F �!ƅ�y��'s��c�>@�����!Æ�F���'L�IV�$j��"'d�4� ���'Wr4B�A�:;,�}`g�O�3�ƌR��D!���Qpl�n@Dj��=a�P���'}qO�`�����O��ժ�e\�P��"Of�\�0k��-;"�D8�X�2�O��=%>��/V,)�`��+�i���+ �;D�x�C-_"!#�-���J8D��PBLȤh��u�r� �fU~!���7D�H�w�&)ZF���+݊s�&�,a��G{��� 䵡��C4Oмس��?)����1O����2��0��E��M1 ��L���!���S?���" G#j|�-�vK�!�!�DW,*J,���L�8*U��	$h!�ĝ2�AӪΚ1^�b�\+*��}r���`�ϸ<6�PƆL��&�i5D��@��ݞg�ʵc���U�����2D��{��ß>��X�m�
��l0D�|��HF�2O�ݳ�(��S�>,��j���{B�)�'�\t+�b�K3<Xi�փe.x�ȓ� �����8=hا�Z&�ܦO�К	�0ƕ����;S���A�DI�.�����<��ς:Ɉ]s7)��>����kM�<1��C�ww�h ��-{�(t� � F~�'YL(R蜉(��r�Ŝ^Y�l�ȓq���ܙ.tV<��	/rv�ȓIԠICp-�r`>BT �J�I�ȓ	Ȭ�8p�_�B�^�a'g3uK�х�Iy~b���ɂ����&����UOح�y��)�Sg}R�]�N�|��+�,�5KJ��y�b�4pt-�g�	#�A��yr�74qp��}0�������p<��D�zB!� 'M!\��,�wC�/>���ȓHB�k�mZ�}]�%j$���.�"��O<�c���i�',���0jS~�eY�i+s!�^�_ P1��i��p��f	(���՗xRW��>O��KGmx�cei]vR�)�"O8=zJN$�Z��P��-Xb����O���d�%I��@�F��;B%�V��{��`~2'W�f��$O�8�>�r�-�:7*�C�2�h���/K0{w�aVdȩs����M1a��"� P�&�A#��@��I�`�Φ2�B�(g�� [�_΀�fk_7-��D�D$O 	P�Oh��~҅�:�pӀA�$۞��g����>�U���#&���ԼQ�F�L%�i�pϱ��5"�<)��tGe�+ ��?��Je&(�HO�c� ��t�D�D�l�,Q5P+rd�a���u�v����/�2]e���R"I*q�T�%NL*�hO�O������:m�=h�Z��Z.rnJ8C�U(�x��\��L�%�8˂�b�&���D(�O��Ci��g5H]qe��;>�:e��
O�堔�]'UF%�1eI!Za
8��HO����á,H��n����1$�:V��x��	��� �!�z�3+�l,B�ɗ>GNd��ꌹXLV 8���0���'��I}�)�S�G��\�����RB�H�X#�"O�y�E��QQ�԰'�X/E ����J����2KI8�P;�i�<n��ݸ���y�з3��j��j;HY�>�yBd�3:��,�u�=�=AD����x�	I�1��HS�1<x[V��nI`B䉔^K��@�E����:!ɍ�&�C�	
sqn� M[
�����g�5L�B�I:c�̋Wj�p���=x��B�Iΰ5B!��q�JyÐG8�tB�I�k;J�*�����-{�Mc#�C�	G�6�p��oʍ�d�ZbRfC�	j����df�̲�l��"-VC�I�2�� ��ψ�rr������pB�I�]��d�g�n0i4F%	��B�	#Y����F2[��sa�ޑY�2B�I�~���Y��R�.Х[OR�KG,B�ɺD��㤌E�Q��Ez�*��{��C�	�UB%��-4y��4�N;&�XB�)� 
�xB�P�Q�,����?<^�!)�"O��/\�J�j�ë?3d���"O�8a������Fȇ�bL��'��	�_�4�+��@�̨�F$�G����ĸ<�@KM!H6�if��a����0��O��~��^$��q �. @x������+D�����F�����ʚA��QJš6OlQ���'?�>�g���~튐�FNpa[uAE�<�Ё�(G�k���,�h��Y}�d�)��'w>Q���d�M�0)�1e�P���<D�l��FDy� 
�%{�|���*<��j�t7m0�D�?馟~�h���k+�q�W$�Y�!ɳ"O�����5+�1�sADw=ޔ���|r"U���Oq��1��<�
��k�;dd��}r�)�I53���W�I{J�Y��C�.�!��\��l�q��/l�I:s�ay��ɣ5B�)9C���X��eRĉ�/�"C�ɰ�J�p��!J��9 ���9a�&�	6�HO��=ɳF����Ip�C6{�@d2�K
F8��&�4�$e�D	"�Ǐ\�ٺ�˒�kӈM������$Bc� �4�7�E"� A��">�����y\��ȕb77�J��f@G�bT�ɴG�}2L�9G�X!B˓.So�u��F��HOĢ=�O� Ir4��i���x�H:��(q�|�$��	�3@�5I��G9����� :��b�IV̓�McL|B�)6�h�'�[��xh���d�'���FyʟX� �5��PѤ��-��"O�U��#�0W|�0'dE�~�
���'�1OH	�&�Ѫ|���h�E(E�E�b9D�@Q���*D��`�F0~�~Aq@nv���b%H�'�����V� z�1 �(| -pl:D��Q7IW��is���3�%�U:D� +���)xJ��6�L�;�,0q��9D��*+(f���H�*�(�3��+�O��(.F.�pp����<�6����'������.!��XA��Ȍs��+D�H�k��X��B�%��j�!�9CR����N��D�hg.�+;�!�ā&P�ܵr$K6;$:�x%n�|�!���4Ǣ�6B
-@&��NԴr�!��f����燏�Q&�ݨ׋A� �!�$�<�ܕys�ɤ}�:9U@��!�DF2aȒ���eJ�v��*��X�|�!�$.����#u��kt�j !�u�ԫ4��E��	����,p<!��
}��D�-�B,ڰ�Նl�!��9ix����B�v�$�Y�!��=R:�%"%�ў-���N,M�!�D�6�h�x.ށ#����T��g�!�J���y#ÉN�[�^�j
�5�!�D�+P�0���훌6�d�T�!�$���ܼzf�,2$9c���t�!�DҐ�\���*мt�d�ib	z�!�DB�+	N8S$fQ�&y�Y`Aʚ�:p!�T�c�T���
�S��y�(˙c!����i�L���©u@��gU`!�&x��B�yN�(#����F!�N�{Rd@�qm�6~:*-(B��|E!�^�V��5��6I%���W�&!��+!)d�j��fI��K\�\`0��'��x��V�c�V�)p�ŀ~m�'��SF��T�D�`)��Z��'y��P��1V��`u�T%8&�d��'��A
�q}J��4m� *����� 
icҁIw�h��B�P�O�R�Sa"O���R--�Ub�˔�*3���s"O��$c�?0���J�Ș=,�Y3�"O`��ԦJ�x��e�1�=]*&ЛV"O`�ІOɺ�����h��m<�J�"O�I��!�A��+�	@�{P�R"O܁o�	
�(Lp��V1c���C�"O�(�%���:$�$�\>��XC�"O��2S'N�_�.����6S}R$�"O �R�	ԘU�b(ŀZK^�X�"O�� ��ذ*�iw�W<K���"O�Eo~3r0akɏRfh �s"3D������3$l)P�
5x�="��7D��`�j�`�8y�]4'{���di3D�<��%ְ?�`=�R)��i)��&/D������@�@��ƧO�s�x��*D��""\�L��������N<2-(��+D�Pp�L� /�L����5\��M*D� ��(��<�x]2���q44�Q+D�l0���z\�A9 �	��a���=D�x��"9�깁�={��0&�,D���4�N�hF=�E$A�>-���*D�0lĭ�|@
��Z�ղ�#�*D���`Lůgz8��bj�;@��A%"D���YmN�Mq�mDj�Q� >D��� �;����	B�0g�\;�).D�|kPD@*J��a���LJIaP�,D�@!G�!��j]�%�Tի� -D��#�B$����G��Z���>D�hc�%:�V�{ֈ�4O����@l?D����ND	��D�������` �=D��iQ��bδ�`肘=9�l�� :D�\���� )��i���aVLxC	8D��eNz;�"�2H�j�9D�$��M� [7B�+�kܼMȥ��`5D����"]��)�b'�][
1ڗ�5D��)�8_����-��I��3D�$ӓ��a0� �w�� �J�2D��K��_�*o�]
�f�2l�i�=D�8 G�۹"_mH����a^���@ 9D��:��a�p�a��R8l��W@%D�<��Q�.qkGl��`�{�%D���l�	`�~���Ɍ�8�Di�wH%D�l2�,�rD���	O�akD  D��R0�F���`稅7�#8D�hzT)�E�*=`����|���7D��`��V�4�B�	�1k�P���7D�,R�%G�3�d�����8�(���2D�D�4>��"�j�E��	)�h4D��P�7td�FL�(nX�e�)$D���h"/\���JQ�q�r�1D��z��F�<�2� ��0(麝��#;D�wI  d��PG��#��%�4D�TC�o�1c�9]Iȉ���5D�L����i��̈wmz1b�iC�yR+�.L|C����z�����)P�yr�,r�<=�"�[�M�P����?�L��?��>���V2Z=r��P�Lx^<D� B�<`�T�b���$)N�C��X�o�F�i��t��(�<<Q�T���!Şm�U�=\OB<�r,�0�����9p�Jslʸ
*|�+�3A�!��Y%B^���t@� )�R�t���{R��+u1PІ�>�1���V Ȓ"ԗ>\JC��6�V�A�ƻ[��9D���B>�4Y���� �ħZ�� )L�� ^�:�dX�e��}ȀHU�&n��"O��h���#�D+�`�	K�����I�����OH�`ĭ����9hp��ժ��uj�Y���ͦ��ɲJ۶��OZ����8�8��j�UN���x�qO�hY��Y�<!�a��i��ICQ����q�%9D����'
B��2���ܤY3�Y��@�P�;�O��4@J�.P ��
 ](
pe�'ö���J~�j�y6��	��+vvZ�i�,��yW�l�
�@$
�5'Y�\Eŕ���'g$�����O>�pH^6JD�LR�oS)�`MJ�/'D���#s��!�䂸�Afd�o;�O� E��O4̫����Z�G�DE�.�9�"O<�Q�ʞ�Sς�5B���4�Q �'���3��iX�$��b�P�Lq�	��uR�6ʓ�n-�B��<q�dL	@�<!`E;��Mu�-"$�ه�Վ�*�h�"OZq��A��aJ1i�'>�D��a���*���@){�$I����U8��"����yw@	
%®�!�f��[A4R�\��y"O��;,��p��풥�oi��nٜ�z(Q�($hř���?�qQ-G�t�`��@�N�x���I@�$4�(�,0|OYrc� ��I�2hb`��ؤt��
�l�"QH=�v�V�-H�Uzό!Q��zʐkm`5�s�ߝ-�J�QR�۲��'H`a��ui��斂9��Ⴌ�!��5D��k�MQ�	��4Y���!�D��r�'�n}K��J�O���g�9��	�V���$m�uJ1Г�X�$�~a{�`���䧡yw�T�2@�fL�ߚyQSa�-�yr޺22Ȍ�̂>'�y�2�Wv���c�CM�J�>������)ipe(��37Ƥ�dL�-�'�x���M:���Z�gJ3#�F�Bߓx�c�+E�w�D�	�&1Ψ�R�N�y#>�����j��MBS/��`�WBn��y��Q���`T�.���5d���'>v��%�mJ�CP*/T_��[$��P���v!T�R,Z��rf�.E�`�5�^�%����R�
Q�"*�<Y����&�A`��
P�.����Ū��`V�{�@�>T�q��4x��S�Z��N�..����DXG=,����%�!���%���(�+n�p�R���D� z�H���h�,9D�����?/���'hT�l�d�O~	#F锑sq�4yw(�:=��B��'I�1�nF0�����l&)a"���5'	,TBF@�;Zr\���H�i+2�C'g|<��[�N,9�o�|J��BV�[�BG^��=��홣&(F�
&�I3z�`�k�$��В=rr�,c$��z�MY.d+ �l�n��S�nh<�g�òs�P��M�52Fh���Jy!2$;7�::�qcD��_済��bC3q�V����Mq�w�<����	4ݠe��>A����'ԈY���2Mtи�I�;2'b���r�8�'M
H��C���uGe"��N͊Ș'׸�E��U�<҃��7��� 
��x5�t��ך� Pk���#��0���aSx����cSl�%&
���ɒqB�Xs��T�|D�e�X�	�>)A��3�Bq�nǥXц� ���pB���@�V� ����C@�̚��=D�4��BԑL�L�۶��8��u(��l��_�(.�1���/A�ep�f�O�NX@�CF	t���"�/`�f��y�T m�jh`E&LH��AH	�F�F Vv)I "D�"���L?�Xj�$�6g%��2���P܊(3�*�O�]��d	�:����拰=O�!�5AÖ_ڴ����j����'�Q�է
}UƅS@���T��I���dן+�]���ň>���ܕU;��XE-ԟ�y�e�S��I�cM BM2������y�nʱ-?bIRj;2�<��R�
��y��ƽA�l�[ �U��p�����y�A�.T��=t�Q�`�n���g��y�+w=V 4��g" u��H�yr%Rbh�8���ǤeH��p4	��y�V*N��0!���,/��� cO���y�bٕ�����"&���3/�y����3gM�`,�A�͢n����'V̕�����K�fi�)ڸ
�( �
��MWb˲T\h��aj��K�',�����MX<�t��/,���	�'�L��Q�լf�|J�MP�>����'
f�Z0&Q�@}�%&2J��`�'�^�R��P�� 2!��]�
B*��UfN�kT����'r^M��e�	E����*o=��a�N55)�=���;�Pxr*7��@Xq���"�$����� l��Ş-�'7��s�ı2V�O�'v²-k�	0I���p��)wl���	�6H�]:%n�)3$H�'���K�J��.�T�a���)��� �N�a��H�b�(}��\J��҆q��a��J5V��B��<1��ߍC1&�`QK���" B�<4�,���=�@�*���k.�g�����'d�;��W����c�=<����ٲP�z��Y��i�1/�B̧[��Y��oO�0ƛfN�	s�����Y� ��JU�ϋ��?�7��$T�G�@�3�����.VxY0��ÇzX� ������S���?�뢐>���R#F"1�Ͷ4y�<�����N�(�Ō1�����T?}���{�J��&
�`���vmۖk�T���iԹ��Iv��~¡�$.�,1�Ð�9�倢�X�򄈏@��h�6��1eRd����H,=��a3�
�v�r�dC�2 b�[7�̈1Gk؞(SV-}����F���?@��"H0`}\���'���Ab-��D�O���a2�ՒF�����7�pר�~�����5�򡀖0T����G�KpR�X���VG�)0򠅮h�p�TgIy��H�����=�O@1۱�A� `+�u3�uN��@�z�Tq,O�%R �L:\+6��1��QX��c0"Ot�*��"h���@��X.��`
�(��䞰]�a�d��F���%�=d(65!`jϏ�p=!aO��LO�ҫOD`Q�B��=m&y���40���'o  a1�Z �0ʓ2�͘`�ŦY
�����"^��<��m��\�	
c�:�'&p!����/3���3��:"�ACB�Y�8�	<�vԈs���7!p�S�'0ݾL`E!M�*WĄՂ�k�,Y9�U֐�'�͂U?�9E�2�^��O�qaK�6&=n<IS� ;1�)0��ѝ��a�'a �h)�3}B�H�Nᢁ�ϓ�n���/[/M��,��n��5�,E�v��!)�����>��M4�)�6�8�� ,�P�M<D��1��:�
 �I.�D1�ՃL?A��͓w?��*/]L���OG�5��89���h�䟏+cT�!���� `%E;�jt!�Z�|��(J�X���I,sD���%0��	�p\��Q�Q��|���(���wē�qG& B��P7���-ܒB87���G"D0����V �)�SH��u��/��-n|����n9�����;���GǴ� �Os��t%L�*�*0�'G��Y���|���㷯�bK��@ dZGx�'ǜ,1����$z1N�-����AG9	��X"�S������pv��@-�&g�:-�O��2��4��L�n%�F�NNX�t�Y8)�:��Tn��hO��Y� _Q>�J6nj�$�ӆ�*���2���.%�t�MS9i,�'_B����d�g�
I^�!̎:�P�*��qtc��:����sq�Ё�S�%*���DV+-�6��i��6P���#^:/Ih���'�J�p��x�0�`�'p��!e�V�"�O�)	������D�":�'��a��9|Z��B3s�>A��'��p��ݒmQ��a�aօ0%��YM>i�!V�1'���>	���G�<Q�T��wx�h���$D��"��� $�<%���vJ��ej D������\���c��?(J}��<D�<Y��8O�t���8J�H�ѷ'8D�d	͔%<�6�iԉ�/
�|���3D��0�c���@��Q��>�����1D��+"�2['���� GK^�Y��-D�ܹ�O�o#Virf�G1p ���&�*D�H�g�XV�o���i9dM&D�P��I�/h�$ٖ��9��RTh0D�Ƞ�Mk>)0���V{ʸ���/D�Y���G���guBY;'�!D��1��	$<J�I��L{F9��>D��u.�#���3�tI���N8D�Z���g��A�틷A{����9D�؊#�G,^��uA�o�9�|�вB3D�@�s��.����Ac2#V�m�t;D�V�C�{����@�*F���"�6D�|�ԓk<�!�Q�G�a �]i$�8D��8!��,<;pe ��«s���7D���Q���&Ӹl(`+Ļy���;'7D��&-H�L�ꇁC�X�PV�;D����3:r~����Ě}C���dD8D�� ������9Iml�h��S*'E��D"OJ�xȧ#貔a�
k�0��"Ozh�M��w}+��N�R����"O��bp���{���C�&L��0�K0"O^%2� ���d�
";E9ɵ"O�}c�)bU��k�^�T���"O�M�&W#>Y�8r�%@��:P�"O�@:/L?l�0Ջ@�6�2��p"O��[3ʑ>W*�h�e��>@��}�"O��0��-OZvdI�"V�'�D-r"O:����ɃEm��d#;���Q"O�q[�c	a�p�%,M�@T"OH����8%#ZԲ)ʂcN���"Ol`;�hV~��B�	-��C�"O��Z�F�"�TYd�M*R(4�g"O�(�璘q���"S�Z�x�� R�"O���W	�� ��1i���%�NDR�"O�h���ܥ����C��`��IQ�"OJ����H=X�4�EC��|@i!"O��br#h�&�j��A�����"Or4z��Ju�,�*3�Η,�@���"OX���'��i����$�I�Z�(��0"Oz�JE.�5��nA��*���"O�=�3��?I�X�÷ظZH��Ig"O��c�)�&j�R[�1��`�"O0	c��D8A�z�hEMT?�����"O���B?�� ӅF�Va0s`"O���0���9�6I���0Z�x"O�x��"�/r��dP�K�u���"�"Oδ��㖩'�:i��G2 x��U"O8�ۀ�R.L����XWV���"Om2�
Q�-������O�&8X�sU"O
����\�v��41���<1�H��e"O@�U��Q�D)hu�߾['P��"O̼s��X?�����U�:}�"OtؕK p��	30Y�p�*}�"O�� "�_�P��$r7�#=�¥��"O`�v����#'nW�-�>=4#.D�ȡ��V ��3y�0�@�-D� c��1<pRE�!�	~�*�!,*D�08s�(��ȫ�@�-T"h�*O��ˁ��*���u�$ɲ"O��9'�3m�=&�,c�ԡа"OIq���6�������ڕQ"Of�)"P�9�ΐU��8 C4a��"O�c�&��~Q�b႕	�Z�"O�haB	bྤJKN�h=��"O,0 �HmʁQ�(@n�i��"O2��J*6@Y����u�e��"ONi�"ڞ=�l�Vݺ~z����"O�	/}I�9ⵌɥ����"O�oS,Jr�V$�?(�My7"O������0��ɂ���(s�$�$"O�-3���n&�(���@�nU4��"O�y3�[{�t�b�ę&OP]�"O�]	�o���(�혘?.�irD"O�ӣ�T�K:�%{�b�8@z�9�"O�)A�������1���8��� r"O�L)�'&��	!J�=��h��"O��)+�v�-�F�AE�$ �"O�D*�
̚Vd9cgC�D/�s7"O(�9Q��E]8�Z0e��m(SF"O~��'�03�l��t� �3n��"OV�zƖ�0��}XG"�6��|"5"O� :�y�a�2GoZt��O"Dh��"O�9S��J5:���t�� T�|�"Oh��UK�&�=��E^�	����@"O��K"��1y�}�6�S�fy��"O\����7��5�ת�e��J�"OZ��2�p����l8�d��*O���J�LjX��".n�s	�'�lA'�$S�(�;�MO������'�t�gDW">ʠSף<*�(�'�����*a��qlR�/a�S
�'|V�d�)p\h�V臷"c\�`
�'���II�ֈ�bÀO�f���xuZ(p �V6)~<)HFڜ"2����d�F�����;N��BB�����2���ӍH��{s.�+\�Ġ��xh��@�LF�U�Nɫ�`�ȓZ���wL�!:bء���,W����D)>�8����=�lU�� às\�Ey"��E+:�D�4��z���*Q���;-�	C���!�y��ѓ.ً��e���x���-�b@��I�ɧ���D��`͞��2Û(i��Щ!F�}�!�D��kL�� �Q+F���k�D��d�!)�" ���%��	r۔ْ�-_+
d���Ѱebf���@�
%���pޞ���C�3Q �,(:�%T[9���E�>R~I�G`A�jk�L��&�80��Oܐ+���Jw�䪴o@F��b>]U��<;��� +�-'�PA�+3D�L ��C�&Ǫ��A
K�vIf�⒠��s�&��L����Z�$�ON�}�N�@�� �TU"u����"ap��ȓ�\�8n۞@�^���\��)��q��i���}W��AQ(R��2#S�(cx|���۬F��LZ�&2|O��Z�ML�`f,�R�:/~��eF�D �c�)�*a���7�X�S+��J��d�7��|'�,
���D�F��ՙeE&{O��3"/
�JD�O����ʔ���qFҶ 9 �'� ���oO�/���S$@R�:�TɑJ�)M����҈<@
(�Z�#��F��wo�p���Ə}I؀��ʝ	$�q�')\��gH�.!X������f�z�"�m���2��)"�bI����.��$��W�'4���͍.t�+g��v����
�s����G�"�=p��Օ@��k @3d�~Z����L}9D	!�O���Ed�+m�-v(Ϸ((>��0�	�^C���b��L�B�B�!�I��@�x���i��y�@��A�5M�!�0��ؐ	�;>������l��ćO�٩��&��\Kt�X����h��'��kW(V����[�"O�ј���<`�-�=j�0����o%|�+&�[�3�D��fH�K�g�*�
A� (�(>��u��R�F���I87�|Rĥ_|1� � `G�o��Ѱ��/X=�I�wc��
f\ڶ�'2�
���+>�PP�#���-�zЈ���)e�����E$<�D��rW�����T٦��G��(�x�1��;�y�L
�7��H�&L�&��~rĚ1k��PP�H7[�J�R�"�'{�Z�����+���*C;�l��!�T��
�r$���a���A �E��R���}����kZD��$!c�Q��eȈ���kE&Գa��A�@ð�1�G�=M4%��)��)��z�b{��Bd�|=
�f�F C��0<iūр)�Bb?��G��B�|Y�7/4�.�O>D��	%�\-W�T����dS<�r@=D��@��K0�����CF^Q腠;D�`��*NX�`V�� ��5D���'�22����ֈ.�09��.D��:� ˆ$:��tf�:p7J=	b-D���5�P	��k� /(�X�Q +D����h�J���I��ղ0�4D�$���H$>�D9�@���"��)[�5D�`��NL�yN��������H%@��2D�����#wf����iæx��BǢ-D�� �2���ofV���bF;kH� 
s"O�09�J�_P	���24Kc"O���j��	��`�6"�k\�J"On4 l��q�`�V��K�$Ub'�O��c&#�4�0>�kͪA<���ҋR�`�^�0�O\y� [�J�}�Ή�I�f�-Y�Xf�#�E�u�C�	3�&dxv�ZK�B!����;
�C�/f��͡�Z�,x��	?��&�>��4���gŰ2O^�c���w��-���'*��Q�
�4���v_��jb�K޼��⢏�,H�X`TΎ�%n(�d�.��	]��~2�*!���R�k:�S�o���dQ/:�t+P��>z�����)��@IJX>�i�G�4Sjn�8��'K:4�De�#~�@��I�|6\H�G�#n� ����_��̛��Ä�~"���PzЂ%�)Y�Usd��U����1�r���%Ө-
0�@6C�x	Ŭ-�O�$��� O�t;�D�#C���K��F�iP�J�UDz-"�'h�����OP���O�y�"S�d`�|��BJ$5D(�,]��i2MO	$["I�O��u9f�;�<x�U�¦��8�([�f.!��#}R�܊�ۏ]��4#2���o�:(!0ͯ<1�lH*D��`A�<��#��CF�^Ė5b&�V�,����D�ߟp����eE`�"�'�
��� x@4�o^<e�Q�d|�	0~���@)Z��~������?1�_&v�Hd�V�� >���d�R��,!��'�<�p	݀Y.��7|`TC
C�t����Q��qM�(<qO�5&�,#s!5Cj�dR&W!h^��D��	�rS���0�˓m���G'+���Db_��d��D���ToW7ri����"Y��O 4��AD�|9�'���q�ߩ1,�Qf�S�9����Is��t'N}�<7�ey"�Q&R�U����<iO�&S	�E #Q���2�L7`�[aMđz7��7扑{3�0B W*r?�g)��*��V	��Ds�	$p��`��8O�D�0	�Eٔ\*g��b?y���OgzH�'�±4�B��C�_I���X��<u�� ��iK�.L��?}BB��V�. �VSˮe�TVX# �;��"?�0�ɮ!����W��H�u�<�:�$�0�� �	�6]���C�I�OT^m03ʏ����& ��O�z�I`���j��Dh��W8=��с,���󆎏��(O�Lp`FV;;����lu���0���Щ�����>�j�e�7<�'(�e�u
Jj���*�>e8Qn�,���ʅa�b=3 ��x�-ȓ�7��'�1�S�״��@06�Sc�:x�@��E��){��+<�:�킴���s�i�z�1Ub�]ͶI��O��fQ��Cj�D��ѫ��C�P)���3�}�Z��k�lJd��*=7b %�<?wO75�qi��ũSB�+
$r�Ze#I<qW薕����ě:|{�! ���Fv yҴ [r�p��7�� 7r�It�%K��gL7}�H�ḑZ�(��gۂi�z,B`�D2IO��%�Hy�%D{� ڿ��ጒ�E��D�hD�5.x���0�=��10��>���.p|�>�Ol��A߱Z(2���fќ
����DQ�����JF��H�����\$����{�H�h�̜0W8ĩy�l@��0?Q珹vͤݫ���#a���2T�!ts��{ǜ|B��a�4�^�d�Ŕ>!�B/	|��:�6�A� T�<)ߞ6��\�vN�y�.L)$�|�	�x�*D94��I^�FE��#W m��!�.W!��#wr�R6� oqs"ùQ!�R	�l0�HFVܲ��gs!��;�:e��B��e2�q���NJ!�$���F��u샷|5$)��ȂY!�S�0�\��6�5�ڸ *�h
!򤖢db��� �vg�5���/
!�D�9Y��W�!5&z�j���) !�<r��s�H8y��xbc�!��Iz<���˒	+��2C]=Q!� ?�x�kW(̅i[�T��b�=!��,�r�h���A����I(�!���3cp������i14I�d`�T!��58��8�7	�8适K e!�ę�9�j�I�)<����/dX!򤐨"���3A��\��'`23�!�Ď	�Q�d�������e� %F$!��^9�4UJ�C^ȫ�k�(�!�$����X�d�*)3࠻6i�7X�!�� �ɨ�MȦxI�XHc��_�l��"O�Q94��fR Q�c�ĉpB"O��S@cۉ�6� �HW3N�C5"O��*���p��E!v�m��"O6� �Á"s�%�6M�4m@���"O�Q���.���S-
�)�"OZY��#	�) �:��X BJQs"O΅�W�9J�IX��ï["�"O��95G֊z]��Iq��*���"( !�DF�j\����[P>���>�!���'H���V�+rOLɠ��p!��>dod4��1P�A"�Gmq!�d�0;)��p$���_H� �a1Qn!�Q�wn8 ��&*6�b����8S!�3 �%ѥ�����*O��pK������µxJ6<2�'.�pƇ ���d����"	�'��C � X�>h����^p�'XR�	���6u��
m��
�'�^�B���>�*(15H;�d�
�'����'G�/܄-z4��e �aP�'�0�n�������	G�� �'U \�W�FJ����Fȫ.p<�ۓ{B1O�]"!��*%����A-�<@��@�'��s^�Z�	\���S�O���2@A'6\&%�W%-B�9��vuj�E�<��8�\�S����6�Ld܊t�,)[��տ5jH�'*��L	V>5 тM�T��`+��F�5�6�C&	��Mc����l�ݠ���w��%E�Ԇ�[CZ=y�MW��u'DB,m�U���VN�y��y�� �'ԉ���?��m��!�tS%�B��Ջ�$L�A�$�*O���G���M�����\� �㰯�	G�I(ge��,~B�*F2��a۰ҧ�O���q�K»i��#`L�`��i1J<V�ض�j�r�8�g͇'�����ψ	_CD�a1�>ٖ'��~GN��Iq"|�'���B�?L�J��a��yO�9Iߴ?S�D��t>�ӧȟ$�	��M�85.P��aW��hum�P�� �C�"}��:&��:�����.)�p� �8�Ⅰî�|�ɩp5p�	ç Wp�p,(2�\|zTHS&e(t$�����&M�T� �Ӈ;|�u�&
6 `bL�2��H2x��Q�	C�ԟ@���O��2f�G++����,S~  ���cgz��"��<�%� ���(�!�R ��(O�G�T5"O��р��-:����
�}@t���"O`�ȵ���,-��;_�b"O��� $"��F�c8,��'"OV���iX*M3��֞DH[�"O�y���̠5��B��Z��
Q"O��d��"T����p.$8�n�R�"O�,��!��Ds��!.Ȩu�h,B"O�����)""�(�gQ�T�p�P�"O���ѤU�s�{��b%�EX�"O����"R�b��d�
�V�S"O���W��3Y��Q$P�N�έ��"O��K5��.v6��7�L�Z!��!J��������Y�AKk!�_U�2`�c�K7JR�2V��4_�!��ӢG,R܉Ҏ�3u'�9�3̄a�!� (�E��6$=D�ɷv !�$��Y���#�@^� %��C@�)K(!��?l�D@����P*�hwƙ,G!�Vu쉸�Jܲw4(�䦂
h�!�R� �ȃǺ"r\lrb�F��!���otq�´���+ m�-P!�DY�5V8����1��ab	5k/!���(�����pe����:�!��"����G&H&�\@uG!�!�$�d1��j�)۶}yh�
c��n�!�� ��C`�2�\�p�Cg	B�"O�1b�G�s\̰��.59J
=H�"OlYK�,��"�OĬx-��r7"O�ũ�Q��Q@T��;B+�M��"OR35��-vV�XЗ$�'FA0 "Of��!l˰E�J9
vc�<�p�T"O����Y�2�a(v�5T�,(4"Oj��׮9μ�p`�*&�<�+ "O�\SkX4N[X� �N_~4̴�!"Oba	aܥ�v�Yao��_
.�&"O l�B��4p��\�p �o�!��	�=�a �b�RM�e�!�D Os��X�a<+���%�Q1.k!�D�3_6ΘY�̌�{�0�IŦ�@�!��
5Gw����END���E])C�!�� $����KI���	P��#Ei!򄅻|̄��N˼���{�T�[�!���;p p���׌��؄��y�!�$��o̶	y�L�&"��$Z��H�a�!�D�� &J,gx�*�N�X�!��J�KE ���/�-"H�e�!�d�#
wf�C1Jg��seZ'j!�d@�c8ȡ�&�"Wej�@f
�*!�d��eW8�sSiR�BG(E�I^��!�\�=�`)I��Á=����Z!
!�G����K��u!Xm��䘱]!��g��͠w���H%���x*!��Vݬq���ؔ��I`�[�
!�dJ�*�H�*g�Br).-��A�5 !�{&�(�)L�H)l8p[M�!��_���AP�sD�{t`�6�!�:_�x�%K�o�����F�!�dW�p\�Dz�ːb��dp�M�m!򄉾s	Jh%���'��e1D�^�d!�$�)55zL���~f��C����. !�$��n�(��%E�O�8z�%�"�!�#J��6A�vB�my�N�%�!�D�X,x3���(�T�Em\3+�!��E3��X�K]�nh��a�зe�!��_��ŹQ�A&mX�dۛ&�!�dX4s����mճ
�0� B�#�!򤂂A�>�3�أm�^�B ,�8�!�dM5?pXYrS�e�D`2����C�!�2f�^<���P�:c��y�ʆ!�d΅@�&����G	�Z����[�!���?@�0t�Ìy�A�JDO=!��d�@�s���3��I�1�M�Y3!�D�����Qc�˒�T4S���P!�$Ƌ$�X(��"q��e&C1�!��/��݂�
W�cRdh�e�պ9!��C�L�4�'V�ಘyӮ�3^�!��]�ade��O�8J�&�fD9x�!��)Y��a�1f�-P漌�`D�-;-!��03x��`�S<� ��cʑ+.!��:D�(��.�<*Cv��bJ!�D�� '@}4��s��T鴮K:YM!�),��Iw��"9W�e��
�!��� _X�
G��PKX����%0�!�J5l&���`�� 1�[�!�D�'(b�hDJXz��s��(<�!�$=W��1RǊkvx��3�!�Ė=�@�ˉ"\��M�s�!�D�A�1"���$Y������!��R+b�$Sa�3��}ˣ�Ē_t!�� ��8���}5Ȁ	\,(�b�"O����*٫ �����H��m��3�"O�Y�"���[u��-�	0�"Of�[b��L�
L9bg�.C�@�1A"O`akN�)M���1Kx�4�"OB�A�_a�u�σ�p
4�k!"O
�qF�����,rAԌ'���B�"O�P��¼?��� 
�!�J�� "O�<aCD�m���:c �Ps�"O~�a�M��!�\�.W�Q��z�"OHxѓ�ܵ_-X(+V/�
3pz��"O���'�D�K���W���s"O`�3�V0lpnic#�7�)�"Oΰk�"�Otسl&1܍ҳ"O��å���`�!��+jLQ�&"Oa ��}d:}tD :6|�1"O�d�T��;��(����U�e"O����Q�n
�3dO3q���R"O�0�� �a��,3���C��4"O� ��H�#�����߿]�މ��"O�� IL�6,�H3�%��BI�F"O&}ٱ��?k��@3BK�d��$�7"OP����x��H�w�2g����"O�щ@�L�yy�	Q��C�k�l��"O�
1� �Xz}aã�8LԐy"ON�V��oj\�R��-�PqI@"Ot���L�'>-2���%N{��R�"O�Q��O���EK�o_�4dh�"ȎCb`J�^��2o��(i��#"O�"�h�'LV�� ���@6t���"O	XW#Bc@��3��' 4+�"Od,�a�
�Y�$9yR�A,}ܵ�C"O��%շ:��-�rFʦ;`�E�U"O���G��:]�� �ߡhJ��"O�t8(�-:����mg8 ��"O"UB�,S��	���0(��X�"O�4�,�[�"���J��rĥ	6"O �#��Z�D&��s���9���+G"O�`��hOt�ht	�V(��b"O����攐�k�$w%!
�"OD��+�/WjԹ�gW�
`��U"O��ܒ�p �$&E	�X��"OPh1!� t�$�Y��T�⁺�"Ov��фN�f����AJ]N��%�q"O�h�&D
`-9T��W3�)� "O�J.Ǭ2
hp�c���7��}( "O\�XA�#�t��S��T�YW"O��A���0p�h��":�����"O�$�7c�Zv��S��U���a"O
9	��MP�Tk8w- A"O��p��U2�����Ň�Z̰�"O��Y��)z�8�����r9D}P�"O�E��X��(�d$F�y8*-��"OHۧ�� .2���E�7ƽ+""O�)�#�&dl�{�C�<4�8Zf"O���3	>5�H@�ĳ<h��"O<X��$�w����9R�ƭ�"O�X�cމJUVe#w�?>�&��"O�� �Z�a��� ���"OL���ǝ8�zP�7��:�P��"O��wEʟp�r����;�H�"O\���l��8E� �oE�yB͠"O5�AЄrNh�1�#��bU �"O��#QaB�h�X�ya)��65�"O� ҉���\%�	k�H_�z��I�S"O�4r�����X�Q�й<���Â"O�h�@��H�|�,�4sL�h�"O|��#��H|B�|a�k""Ot�3TK�oJ�|����r�� �"O8�`��P�ln�x�֍�/[�j�"Or4B�Z1�@�#�F~0��@"OҤ�D��b\8S�G�/i\���"O�AC��6��4���
<i@�;�"O�aa�I�H:��Ä�WC�c"OH@�&��*EI8�ś�f,�$�"OXX�JJ
#��x���\�w)���"O~��&��C�Pivb}&u��"O0�S`�цu�(QCF�t�@�*T"O���f$��hDPY�a�:K��#g"Oڨ���Z:iJ��Y6N�<@h�C"O���,�o�ʠhw'��@��)�"O�U O�#Q���RH�Z����"OJhJ������q'4m��1�"O�DKe�X�)�����>�t��B"O��b���uJ0�+b��I�R)9"O���(Ե[���ȳB���ȥ3�"O4E���6w�6�X��G�DZH�"OF�9aB��xN�!�K�a9L�p�"O��/F�Y.�=�`P�;-�)g"Ox|A�H��r�s�
�:�!Q�"O�	�%"�9�(�`��ʊ9�E@"O��ɇ�L� Zt�*� �"O.���l�B�P�'¥h���J�"Op�@���3z��Ҵ�'��)#�"O(x1f�O�a˾q�$Lƥ *]�s"O�x�rƈ!"�$!1
��!�"O�i���-s�T���	X |�Ep4"O��I����Ċ%�I� )o����"O�E·IB}B�� )�3�`�1"O��Wg�E�\���C�z-rL�7"O�e �H������A'�(Ԓ�"O�0�̇XP�D���ֈ��PXD"O���)�%6jd�� ��M{.�R�"O�`IB��#�t�&#�&Cb�d:�"O�:�a�b��|��J�p$c�"O������,�(�æ� -� "O�9�p   �D���A	&�����4(���B�?D��Ce!һd�"�G�U�_��Q(w�0D�d���#���Hս^:`)a�H2D���f��q�(#5�-�,����$D�H)Pa4��@�'�~�A;֊"D�����U5uE�E�e�Q8���B,T�,ٔ� �j�b�R�h_�(��A�"O@����/��%p�肖N�p��"O���w�fR��8dM6`��%P�"O
ͫ�AЃ?���<�"軰"OPZ�b����0Ɏ
b�P��"O���    ��'���{s�R",� �D�8,�f,�'k�T铤�r��*uI��
�'���R�������H7\K<ň	�'sv�1���
6� ���.JBF�@�'94�9�MҫE��jD�ݬU�|�
�'� �J�#΄GU���D#Ve�us	�'�N�;ׅ
��� 0��]��y�'��s�>K��9�g�+W:"*�'o,m���*"x5bp	��T�
%��'���q��ã��:���=K&&��	�'��`�&G�L�1�� ^�F��	�'i��k �w����%b��2 �5�	�'�|����F>n~����䘦D,���'.�T��*=���EÌ�=&�٣�'�@T9�h�s��U�R0��S�'��0`�ʻ )`9��e�5$��'�nT��n�o4��f)܍w�]��'�hu�7� ��hx[F+�5Wz84a
��� �����α�v�˯^����"O��) ��u� �I�M��F�� "OVô�ѽ},��K�Z�x�"O<� 񂔪i����"A�\�H�k�"O*ᲀA��R�>�Y��õ����"O�)8��ƥZ�"TPO%{�nqq5"Oxy�G��8E�p:�o3�����"OȬ����,�~�ӫ�:�Q�Q"O�-�ୌ� �q2�P�O�(X:�"O����H]�p'�YͮD�C"O�����y�|�K�a�����"O9k���ZS�)��@�[��t�F"O��1S��-�|L!ƀ�v�88��"OL-��J$ߜ=�N��/{����"O�0jt*Xz�Hmw,��5
r1�"Ox%:V^Y����5�j)��"O.`�6�Fqp0��"�T���@"O0��ץ��6��RBaC%#}dH��"O��;��̵hZm�f��-ZT"O��鲌̝TfQk���0�8C"O���EM4�`q���ht�w"O����#M�A�� ^&>�0��"OX-��+.6ql���%�5��H[�"O���ƪW�Ҥ�w���p�F�Bd"OB�9V�ݷu=�"0�Ogp��ɠ"O}ӐO��^�dIЀ�>Ki"�04"ObP����"G4�����WH�*�h��*,�=y���OPx��o�@;��]�3^� [w"O� �/X�
�E���:>��Q��i��c���)�|B L�`������#})�p�$�p=q���7tXk$�l��j'�	g�0��G�, �͒;=!�].�����]�-₨R��O- �qOP9�r痂��`1���D�p�b�(��.����
i��qj4�	�A2vx X�9ɦ�� &I2XA�J�ㆴ�}�O�8�M|��%�faDK�O�P�gԁi�P�"�BO�|��"O�Q���O�%M�Ӳn��R����&o��[<�"���/���:5o�l��I�����~���$]�g�D�p��2a�1WC�?�p=!�XG|�����a��9���8=h2�p���
K"��I�.�!.`��ӦS�&�N��X���?�'Clhi��� ' ���'H�uX�e��{2$A;(�&|[��[�Ol�%�r�]h������R;�3"j_#(�F)8�e�����C0<O�84��qJ@ps� .�tx��I�B��\
��>���~�d�ev�-�aB��$ d�֖ũЪD�;���9�[(`�T$��y����%��$v�9�k3\%po�w�PY�$ �;�~�Z��f���ѧ
��u��)�H���A��c�bmxG@�Q�{"lV�v ��'�<�@'P�'9(��d�9x9�C����RӞNs���ǃ0��OD�'9�s )��m~��c�ªrM�h��'�)��ʵz��x��o�1\�k�5r�x�_'�����V�E�4��I�/Iސ*dE�W�qZ��t����gP�Bt�P%m�=��k�4I��b�m�si\�.�$vm����D9$�8����'��#�a��1�U1G�5?9g�C_i�5�N�( �Nh�QD7q&���,��&݊3"ZĨ��ɟ&�\C%"OVt�	��J�ڼ:�ML�=��d�SD�I��9�d)̨f�ʨ�JL%=y�O���$����%Ƅ{#��f���RPB�e��G�);0��ɊD�Ҹ2�f�q�L#	���P�2%�|���I�ayr+]�v<1� �k����VD���On�yPD� Nض2�F�T��*�E�3x��Q��5,��a��9�,��'c�H��d�c�N��i�;��.O���N�'�<4�Z�.Z0��X���O���	Ն��ب40�Z��ܽ��'a���d�@<"���d۫h�p\�d��>H�X�S���H��ꆉF��'	J�ODQ�$֚
$�!ĬS!��T�'�Ld ^"��x���P��ؗG��/�B)�EB�D9�)9u�X�{���DV�%"�1�p��	1.� Ŏ�h��`>T
!�<�/�0�@�� �؅*s�\sWKM���49��G�V�"�+S�4)���n,$���#*#�����_L��y̂oy���:|i>b�0��h!�	�x�:�M��QE�b�� ��A�G�!+&��'��P�)[B�'��q�燿,*�����	'$�q�ǽ t���B�(O��@r!�VLt�  G�//���OD�'�6x��H�<k
��]��0���#f�`�y�5��'	���pn��%r�1���3k}T���1q�a�tVZ!���'��A����P��.�К�0(OZ���θz9T{f� ���O�)����$�D
�a�"=a��ԦT�D
(�Q���dH<�"
z���3�K>�ٻ�+��(��D��h���#L�>�v}�B
���#�>�w�����Ȉ �J�[Q� u�B�y��f���ɦp>����
e�^�{�)�1;ǡ�?YI�@pf�5}b��|��D����d�V�Ƭ���R�U�pq�#c�	�џ�:�N��O_F9�eM�q�.�Χ*?�H��JH�`|l��+�,lڄ�'6���"�W1X��yÙz�4���+�3��0��;��/1¬*P,C2t�t�� �>�S9v4�h(CO�,n�S�`N�|=�q���=!��2:�%2��.=>й�Ċǳ$<ۓᛳ"��$O�r(�0��͑"����Ο�h+���'@6()����kf��a)G�Ch$��Ü�2'hQA�M��j�X$�B/�0>Y�k��DZ�yz#�@5.�*�h�fBF��@0���5ʸ��1O����N������E�A"Ob��`�,�~Mz�&�<p_bأ��D�8-7���q���~"�A�I��y�O��d;AN@�1�LBR��$5�}��'�*<�#�PD�Ī1�O�(��<o��v����ӆ
'$�mG�A~�y ����j��`^�~�4hTj>D���᨝>\�.��BA�&��P
Q�H.�����Қ�~R��qC���n�'xh�r��主lH�X1��',֡�ch�!q�@hhD#=|q��睻?��1R��FX�L��%Ķ]�4�#�F#)A*���-<O� ��iG /K$��O.�*�1z�Bed]�ʰB!"O�1�"W�"T.�#ǡ��r�t���|�K�w�j�Q���c�O���I`f܀p5:	9��e9��	�'�>MQe�P��� 8 ��&\O� �hR�V�
�'��PQ���>qCR�0�`s�p֤�Nh<�#(�"�*9�R��#*���O����p�등-a����֠78�	��ID^>A�U.�&2�y�	|Y0]�nZ[}��I�)�F��D&��~���B��y2���[\DB@$[5P�d�"V*�'Q�t�r�V+f�?���.Y8g�-����6.��)V�8D�,+���.R���*Wm�;IF���X�yJ�xpP�<1G-��!2$�L-uLJ�藨Xn�<�A��F�1	�U�p{�ΐk�<�A�̂#_�r����
��5�g�<)�)�"6�^)�E��*E� +���d�<9�߫@�p�*R� �n'�	{�`e�<�4��_�j4�H"ya�Hj�Yb�<�Q���)ؒ�1 �
V��� l�Y�<�'���qP�D�T���=@�P|�<Y��W0�Ћg,��2�8E�ǈ�q�<��ƈ4R{��I��пRߎ�3a�`�<�`M��=�hP���7G>��(u�Xa�<I�+M�WZ�"痱yS*2R�_�<	�#�9e3�`/d|B!z6AQ�<����)�n����
�:)M�čCT�<��蛧N���{���l
]1�f]�<1�I"o��k"%�:\~�QHL@�<��2nv�q��lU�M�z�P@�f�<!f���+>�8c$�t*����d�<��Ç�/*��#s�Zj��Dc�<�7GB ?��03^�R/tM�f�Q_�<�ISy�ј�eƱv�E�"IAA�<�"]�,%(ոE�ȬdO.�@��Hk�<q���~��m{5k�6�d�HA�	`�<Aϔ�UVh��@�=H���D&�a�<�U�_3T���Ap�,�����aMb�<y6��::�=S`$ۨL�L��4Ze�<���#�갺��O�\Ԫ�᥍y�<� �������=
>��pH<zmx�"3"O>�x�"��VJ���ND�Z5����"O~�eۂl�I��� 2t�r"O�i�bf��{kL��풥l�В�"OT`#���X5�`����<�"ON�	�^k� ���=V����U"O(�	�%"y�Xm�_�p�A"O4�ɱN@��L0��͛[�<IB�"OL�a���0� �wƌ>ab9�"O��1�^�8�r4b�L��W�e�"Oh�2�/Hg��ɝ�^��P�P"O2���ӧ�8=s�Ͱ8.lT�"O4�����0�̊�b�Q�d�d"O��ˁ���(��Tz@M���3�"OV ��� �" �)��� ��P"O<術/�=g7^IR�K�Dװ��p"Ot��]�:�8��-9<�*�"O��m>6b�yR���9����e"O~x��#��"�8�B��r�z�Q'"O���E�7�x�fM8g��)U"O�X҆��'؁�D����.XZB"OF)H�=Z���U��~Cj���"OFPk���n���u��pD�Ug;D�꧃ʯvj��I5c,N_b� @4D�t���)6�X�b�,�,��0D��󵤛�1��ӵĈ#R�&��a/1D��h�dC�8����8Iol@�02D�P4�(M�a�Udƣo�R��0�0D�`�V-��N�}�K�$x��=D�0s��!t)���ȵ�(��K:D��zak��>O��@a��= ���E*D����se�qB�F�>g�-�@+D��c����).�dX�$Ům
c(D��#J�	6pɷN��jXd�c�%D�@S�׭]�,�+	�>`W@q#�>D���W/( a �?�N	�&D�l���ѷd�TX�aW��� �A*'D�lA�DʷQNh��U�m���"%D���`�Yr��s�P�}�|�(5D��p��Re�јªU�]�l��3D��0͚�y=�ČR��\dp(<D�Ps@o�99��d��K�TK>T���6D����
�&Δ;���Y���ȱb4D��1�:nv��p�A�;><�H9D�*�K��d�@�:���Y�^�A0D�0:� $:P|�D�\.��a�#D�<j�x3��HC״����Ư>D�4a��*C�Ұ�0W�	�ҹq�K?D����g$�(�cb�=j�5(�?D���E��e{������:���rT@1D��c���z���@��qA�	,D���Vd@�Zŉ׌fJ��379D��P��;���"�eJ��v�8�/7D�Т5�*iй���y\�53D�\�πg����c���>3�3D��{Gi�z��K��<}Fɋ�:D�\� d���GC�P49�Ǝ8D�P�@�X�qIZ	kJ��A�7D��Q�%������R`�JD>1%�5D�@�bjߩzv�p�dC�i9
����/D�@���۴fW`=��"
�Z���&D�,��,Z,6�h��@ަ72�$�8D�l�A胴eP�㱋�z( e@��;D�C���
J�,HBÅ�+e�X�A�O#D�� F��듽v�0��Ȕ&`d"OnMaԨ�0Z@j�PA��0�x�e"OHaP��13w|�
�J�&�p4��"O�bQ��V�c���8h��`"O��0e��0��m]&vl�"OX,�A/��)�y �jC.Yg�8��"O�)�/��Ң�Ӈ!Lt`z�"O\}:«̪"��)�$Ö��>�Ї"O�`��A�?�M��eL�h3��3"O����YmL�01G�-�cv"O�H�M'�f���w���җ"O$d���P8#�t�Ă
�Q8 "O&��.�
=ߨ%S�N=�p0A�"O�q�Ƭ9�*DC#l�p�&���"O�M�� �R���eғ4�t[�"O��J�G��t#�	ஓ< ��(E"OԐ�s��{��YómĈ1�N���"O��K��s�����@�O�&�Q�"OR�Sse�R}|]�P��N�"���"O@��G��>.�>�h�̆�� Tz�"O���o�e�pջ��(>댬Q "O����B�'� +S�+Ɉ�J�"O�����p��3���f�d%�'"O(m`�����*�&թM}���"OR����rP�!�H�
y�ݒ�"O�]rd(D�%�� @�\��X�"O>��ol���qò�pqB$"O�@!���"�2GH9��,y@"O� k�@�&��uMR%0��e�"O���"ט��8s��miʴB�"O(�A�IL�7FXI �F,�p����e��`�=ي��O*E	���/_�@x��8Z�HX��"O�`�`T*v��4͕!����i��b�NA���|���+X���a`m�k���㵋�p=&@Z;u�v�
��s���s/S��n`��G%lӺ�ӢI/D���䟜- 8`S�B]1F�*��

��0���L�"�?=�A�9B���U���4�1�(D���aᖐ:�t)A̓a"E�H*v!��7}��Q����		G�LRF�;Y2=b�ǘmJ!��9�ܲ��?D��aT��$R#��{�����k�'�,�C曩y�dwa�:Z�Z	�1��uxt��R�ɿ(�D����{�U(�R6\>�I�����S���_���9�T�pډ�$��05�\��h�P��%�"t�:`X�����ط�N���.Թ������<��6��t ��[�8�v	��:NTP�mG�$���OBFʒ.���W�;��R��b@�v��mH<QB��&J���rd
�_a�u$Ŧ1�� Z�H�'�!"I�#.F�>�';�J��5�˸>�R@�'��8�X��I%|p��_�$��K�]r�� R���q�x��ò�����$?�
׫�o�4�?�'�d�{�B��|�!@ɆL��+�'�����>*����@�*�i�ߙ"։���B�#�,`$I��<yF��U:T�`�A�(M(�1SEx8��@�BI�Rp� ��g���)5c�7h8�١�N�-i:���&ԭ8��q�ēh7��PtfW�j� �Y�A�:5�'	d�8�ʌ�!��ezR-�������@6�-\M
��4jK�$6Tp7��;V�C䉄��(�
��
|�q��m��`��i�	Q��`��c�Dɸ)*�I��ēe��XE��G)��%� AS45��ɓg��p�����`�*U�DoG�@?��)g��$_6h[�ҕO�bDs4cp�ayR-�?lb�5 �o��HMzM��ԓ��O���v ���:�e%�PEjd+U"��:�	�,fx�D���-9
�'��U�ȉ4@*���#I�^`8�B-O���(��"n��tK�x�"�͐���O�����$ڻ!�J|��$\�F���'Y��я
�Q�Ӳ�[�\�����Y8��� aN�.���`���',��O}�� J,!���1�^���i���'>e�� 0���#¨v�a�fbS)D�]�%C�,<*�B`�&n#<�aD><O�u&ͮA�9@#�PH����>y�T#/���3k|��(��S���JbG\.�R�C�ַ ~�!hF�UR
m����q�lC��;r��QR0�Ny P���ǘi߄��'4��hՂ@g�m�N�(a� ��~ݡ�G�٦���4*�;�N�P���
#��b�ҁA�R�$�j�и*x��3'ֶR�t@ӵ�R���" �:tha;�	�4\j�G�x���x�?MI�m9�jЕ(T�4���	���O05�7���D_�@K|�P��4fs���ui�^�<=b�@y��l�dţ�(�`X�\B6b�S~�r�(�V��P��<��*١jdB�RC��O���>�!T�_�M�R��%b�K�\�ViQgti����] !�B����82G�.{��9�gC���  ����yB�]�}:��	`.°���xR�Kn��|�1�ލVc ���P�Cs$�&�'�O~$:�)�=GҰ����A�
�9�_:gf��s���.���,@��U2P��aHA�t��E7F�/9ᠨa䇝CDХE2�\}����f�|	a�6��(�Z-6$�����f4�p��L�E�2�l���!5��@�J����1�M�=q�˓Up@0�/G-5����ר���Oz��+�f��f���µ
�]6uA����<�ȓd�S��Q�}5�	�gO�*i6���&L3p���􌸺6�J@�g̓��`��
C����գ���!�Rv�@8�n	�gJ�XsO�<'�bQ�'˃�R�(� E	6����$,pڍ��H30���DE��z�$q�y�!��<!ucLV�6U�rj��@`�M���G�<�ǅN�	�.݃�A!��!��Aܓ`B��#��,v��8R�r�?u�b"�g��x�N�_��	�$%%D�tAB�U)����3`�ܱ���B�&�V�r�O�	��.�<��|BQ1���+�*�~�4���BV�� mH�"O��)
�mM22S��&y���/>m����d�`?� d����4�(�D�0P!n�ky耂��4��+��ܚ2'O%E�%�B�шu0��k��ȯ,y�tbT <�O�y��`׆t~���q�ї^fL����'|�퉱DД[aF��'SP}�d�/�TI�(~mK�'B֙�A�L�B͊�oV����3J>���ֳ���r$=�����eN��ۈ�b0�(%<C䉳g"x��!�u��m	TO<�	�b����	�z9��OI��\�"̸-��L�E��9�OK����<�r%�t��yӄR�G�0�b�3ɜ��� �sԁ	�"ɟ��ą�I�r؝1�≞��	��$�fL�!	�E�&��#��C�"6�@Q!q��<'N���GKI��Fb����	�B,F���ɍr��97j��5������5�y"��5L	�6�Y�'V
y!��3[��Uˌ{�m���ګ�E{r ݣ7)�9@$)ʫ�!��V_��'D�%X��+@�!�D��0�	X�-]"&f&�;ЀW�6�!�D ?o�A	p"���ʠc�K&_�!�P�(�81��ؿdM�ӱ�T���ȓRƄH�	�x��(8�eN�;T,ԅ�a=���C�a��#r�]
�Jy�ȓr��V��L��k�S��� �ȓVRΨ��Κ�`
�8�	��G��U�ȓn���e��8r��@��3����H0�X�r�+F>��i	0O����1��+�n-L���df��j�b,��hp��6�xx�Y	ԟn�� ��Ak �a�,S?�< '&J�c^���%�~u�"N�()&��J �D�&�ȓ,�h�Y=e:���m�0b+.a�ȓ�&�cϓ�3PI�],g��l��l��uK!�
l�^��i�+�b��m��
��Q�3%zM@#�Q8A^لȓd� y�e$/f�d���`N�H�$��ȓH>ʼ��ˬ.@B��եLHDF���!�|���G�6U�lO�8M��8�D|��#�V�x��>3"|ه�S�? ���2��LA!7A�6f��"O��S�
�5����p��	�����"O�-�g�:z���6�$a�d[q"OK��.eT�#G��=}��3EC"�y�+��j�P@M^9Z�9�bƐ�y�ע�y���Y�_���PbNR.�yr�V&���a�C�T��0��(���y(�
�&�����V�8m��GP��yR+[<�L�E�I2xtB" T��yr�Ȯn-�����S�MO�8P�#'�y�+O�s�xA��%�T#���!��yR%E&�x]�rcA�@�Xt;�D��0?1�!�!-&,�P�L�3�<1��+(�d��Ù^�<���^V�����ѱ~�����Z�<�b��G/]�cJ�(X3�I]X�<��Y�6�J"@O#o�-�f���<�Q�]�Y�$�ul��3���<��ȮO��D��ǻ#W0S���~�<yF��=�8���-��4{��o�<)���(�N���e�Y�<5���@�<�c�ІGL��4/�/.DMP5��f�<)g��=Y�@���P�V<s�Ag�<�#.�97�+��ǳ>ː�$y�<aUM&n��)BE��x0�M�7�|�<���!ef��Z���_v~�%`��%�M#V+
���	��uw�7����-0�CҨ��8c2e��B��~��^F�~��	Kw�퓓<�� ��F�~A")|38�c�H2.N8i��7}���_*2��7gR����Tm�?%������
zr���0|2T$܊XB굱&�K�c��h`�J��CD���O(���Պ�&����iS�@�ZE�҂�94DZ��'�\�O�%���qfLM����&H���*OF|�B�F���a' � V8X�X�'b�}*�K4u\�����F��� 	�'�jm !��,��@�Ԉ?�R��'��P��	j���8�� &t� �'&�8+�Xl�԰��5i��(�'�:��wc�<GB�����.��Q�'w�!iQ�˂*�D�B� �~Ġ
�'��pBǙ\,(z�������N��{����%������.3��ȓ�f}��ӳ!w��õ�"ݺ܄ȓB����^&L�<!U�ު��1��_vl����=A�Fl�*_�� ��x�F�2���%j���u <Y�h�ȓ �4�n�6+�`h�S��/ͅ�"z��$@Yd�Bt ��3:����9�2XʂʭP���j��D�x�����~X%'E!A�Vb!���:�q�ȓPCH���X�2d t#ė,"���ȓb>���NԪ_{�0p`��r7�4�ȓ]���r��B&r��}J�/¸;='\��D�/����ȌZ�f	8�	PQ!򄗄3jd��֪H~�Iȇ���!�÷d��e𦭞#wx���AZ�!�D4����&XU�ĊQ�Қ7Y!�d�X�ۥ�B�W��pq�ƘCO!��X�"�H�z� +�͚p�!��*Z���a���,�9�r#�15�!�$�1jQ���I� G@��`	��y�!�$�����'d�c�H��	=�!��'@��Y���ɯl�x�Wg8`�!�$dJ34K��}�^�'�bi!��`-��M�7Akؙq�ȍ�_T!�d=��ъ7���9�r�^�]8!�� ȐY��6IJ�(G�ÿ*�����"O�����$w�qA���2�D�"Od<B���}�Za��ƥ1r|$��"OL((J4������Uʰڰ"O���Ke40�٠d��Z���j�"O��$D�4>���dD`Ty�"O�h�U��)P��4{с?���3�"O�tUfJ�kM��Y���23."O�|9D�;8Q�b߆e#��"O"ٴ�3�4j`L�"�$"OR�V�Cұ�*���pKd"O}{ (ZV-��c7iE�)�D��"OP�K�EUPt\Ec��[��q"OxŃ�M=gV�,{�eM�5�L�[�"O��I��)6Nm��eЁ>�)(0"O�a�X& E\�`�ق0xk�"O<&��_m:|���ԋJ���"O@�v��.`"��TM���
��b"O�i��c9�6 Y�Р�!��(_�l�3��1Ҩ�cΚ��!�:*l����M�N��r,��YO!��I��~,���LD���H��͝HL!�dCq2`z��#v0�j��!�$S�~*�5j���jZ��t��\�!�Ĉ8ܐ4��G�&cE�i6)Q!��Q�~8T	�e��k^�Z���9I!���p� dq#�D� �E�Bq�'�8��ف�d2�lǄ7h�x�'��y�eC9#�d#��@�,�+�'p���ÿg��1�G�ƾ8 ��'���6C�v!�`�N�\*X8r�'�r�3�'��h٫��ٳO|�l�'��P���hm�\(�$^�NG�}c�',���3OA��{q@MR*�b�'e,�U��@�	�
B�.�{	�'J~Ha�a�c��Ɋ�
>$��B�'B�;��*	�E�R��%D�Lk�'� �[�$^.qD}�¬��B����'tV��+E&;��1ڡ�WLH�0x�'�f)r6�^��`kV6���
�'xB���B�d�xu�2'ߌ�����'���:��Y���%$�p�S�'�ʵ����^)���v�V/)�9�'�`�b�O��4�u�Ɯ���H�'3*��[�<��t����A��'�V�a�`�)T�K1"
<�'�`�BA�5{�~��B��t�q�'	�m;��A>@y�у��m$�b�'��(%��9���&�/lg0�
�'F@�U��l%섢7���v�p)�'����u,*��A?��p �'��b�PJ:0�YQ�S�<+��
�'l�p�x{��S���7�B���''d�
�C�Z��K�`|��''��8p)A�Nv�+`㞣+��|P
�'�.y��.("n�I�g5(��H�	�'��]��ț-�\��S�#���K	�'V2�0�%��	��Z�F=!�8�#�'I�,ر烣}ښ��с����\��'p*RlY2F�������L�2`��'vj�r�V	!Ϭ�yUA�*=Ƭ��
�'ZݱR闑*B�h����<e�`�'{6�R�r�X����!H�|�	�''Jly���hzT�4 M�BY�	��� LMc(Z�X���s Ịk�� "O�-��4;���S꘳j��P��"OĜ�ƃ������:���i�"O�h��)�IrHM��Ň<�$�"O�`����0� Qz&D�-�n�F"Ot���n�4U�w�$(n����"O��;gɤj�x#geA=YE&��"O<��b��6x�L2�C��Ө���"OR�i�H��(LXc�(/l�`$��"O*��b��k.�Ag��J3:|S�"O^�` J?�	��+��%�$"Oh���Dr5����V�x�#B"O"E��	v�j$��c�h$��"O���
#�XC���O��d�"O\x���,m˲ ��y��"O0䂂�T�Т��/
HH�0"O$,R�h��8~<�*fk��<Q�hW"O�!!`MR0~rF��%���"@(�"O ���bئjwv�������b"O.IѷoZ���3��,7�ft�7"O$�Y�d�/$9։:���f��1U"O��`�Z��������(�"O
,x�y�x�j��23�"OY[���=<S>��Bq��}�"OtL���^�r�H���/uZ��'"O�$���KJl9P�_b��`"O��a�C8ː�3��S8#PN}C"OZ$ �I3@�ڕq�N��cW���"O$9����1�`�@$	7F԰�"O6Q�rfs�ְj�S#Id%�"O5�.('��a0���Bp9�"ONU2⡍�V
t+'!;��9�"OA@F�ψ:��ҕ�ӘTtI�"O|+���$T���1�#w���T"O�)��Y�P>x#Ў]�I �P"O"����R��Y(BR"�m!�"OX	�1N�:N��($[Ppw"O��yd�@��t�"C�i��ЁQ"OP���;|�>i���0y�ШT"OB����!Wj��Q�܀L�ꜙ�*O��ď9~�T�{'V�fI@T��'#�e	B��$X�� !/� EK�'\�����#������)�Ȝ��'�
�[�i?I'HUz��N�|����'�&���K
7l��@�ǇM{�� h�'h^��Ӣ0�^S�GǶy�@��'/R=�%+
_<��sF���b�p�'���#@�s<��Y����E��	�'G�\{vdI 180�բ�@�H1C�'Q����X�YyF �4�� �'b���-�5m�6c�eܩ	r�i�'u�I�ص	+^�Q7�^�g����'\�x��g� J��X���]��,S�'Y�@CfѶMK&�	|�92�'����\�|�t�4lU���'0\�Ǧ����14���,���'r����D@�u:Cɛ�?!�h�'tlɒhU[�z\�R�̜O\F���'��R����Tg'{�&���"D�$ia��P�rA���I��ܑ��2D�����T����9Wn,�f	�Y�C�In.�=�磑��h L��C�	.G�:�u�e�F0˗I�3�JB��#��B��A5`I2�#sC�+L�C�)� Z�hTbO�vY�)��ˉ=��r"O´�G�R�6|С��_X���"O�\�"�	NP���N�C縕)E"O�T�S��;L5�Z�-9(/���"O8�� �W�rMSS��1yZh�"O�\ف�$B���􄐠w��b"O$�ᇆ�s��� ��x-�A�"O:��w�v��ЄB��P�"O�����|9(���G�0�	�"O�*2���������5.�y"�"O �a��G2И�M
�,lh�"O�P+�!�Cɀ5�M5|��D"O���Qi�����rz��"Oz�9�EÂU�V�K�!̐d��"O����
��hK4!H���2"O���f���q���+��)J��h"�"O(�ɔg��/��Xw�ҡm%h5��"O&)����%k�J��!BԺ!�!0"O�|S��I�u�T���7�z%��"O�+!\�M�iPLҦ:��i�"OR"Ƌ�;.N�P�J5GRXH�"O\UǏT!�	��� I����"O~|�G͍Aƒ0	�'�2C��"O@��^�y/��peW�h;���"O	*tÒ
�$=�p�Hz0z�"O�p��ؠDx�"C"/*�H�"O�\�!��;A��A�K�2L"OD1d�P);�tiP��T�%��IA`"OJl��&�	R�*	*�]+�V< �"OD�p4n�'R�Jq�P�r�ЙJ�"O�������܊ mR%I}��9�"O�<���<H�����ܸfy\$( "O&�S&V%e@��9���!` U��"O�I�����V�B�@CF���"O�0y�&Ogj��#�\$���e"O����-L#`=�{�A&\��"ObHH�� n�i����;�L,��"O���$��sk|ᩖ�ƫ?^�9JD"O`PtO��|'4;�� =cAiu"O��qT'/no��:��(@B� �"O�{#��:��-@��tXf�r'"OA(�   ��   �  >  �  �  8*  �5  $A  �L  X  �c  
o  z  s�  �  8�  #�  l�  ĥ  
�  J�  ��  �  ��  ��  F�  ��  J�  ��  ��  �  `�  ��  � - � � �# q* C3 �: �A �G N R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr�'��'���'�*��@
X�a}�(��MJ��j�Y��'��'�"�')��'k��'�B�'�@i��
�-���Kd�@~�@l�6�'���'���'�2�'��'���'�\��Ǟ3tK��ШV��i��'!��'�"�'k��']��'�b�'a��K2G�3e$���+�d� �c�';��'���'��'R��'��':�x�l`�.=��W�L�p���'�R�';b�'mb�'�b�'��'�R��tOF
z	��
���i��'�B�'U��'���'?��'�B�'�H����ܠ4V�}���
t�>�RW�'���'���'M��'b�'���'��Z��Q bVb���Ȍ�qn�[��'h�'uB�'y��'���'{B�'f��ZE�[�m��12Uf�g`A���'+��'~R�'o��'�2�'j"�'%S��?c�\RtIץp��q
2�'��'�R�'t�'��'���'
��:c�Rє��ɖ1F8aY��'.��'C2�'���'���'L2�' $X����7M�8�cûΜ�0�' �'K"�'�R�'��HcӮ�D�O���!j��EGV$�b�*T!���,F~y��'��)�3?��i��$
�.66�ҍJ��/w#8M��e:����䦉�?��<��:��Q�G 5/����9#�^�����?����M��O�����K?Aj�N"a�PYp����P3��K��1��埬�'��>IS5�>/� ���<3�<)�'%�M�`̓��O!�6=�tip��.�1����t��装M�Oh��~��֧�O�q�d�i��Q�?���z����H:�D�{��Dk��3��J�=ͧ�?�v�Z�8����k�4��q��)U�<�+Oz�Ol�oZ	,�c��r�eW�4�r0�3��[,6��q�Pm�:�I֟0���<��O�p�T/�0Wa�l�%�*|��t����x�I�D�4�`�.�S���'7��	��4(�udV�y2_WZ(�@_�4�'[��9O��õ�N�b��9��4;H8��c0O`�nZv��0���4��բD��!s�	��ъ	^J�%0O��d�O0��OG�73?��O�@��9E�n=BG	����@i(i.�hYL>����?ͧ�?)���?����?�2)
�S7�+�`R��"�Z�i�%���.6BP��k�h���O��oz>��>6��p���_�M`D��3xTx�	�����I4�Mk��i7m� y 4�'�B��yϺ|P�SWp�5k��I�L���,J�K�T%A��S;�p�to_ 9ʺ�\wI^O ��'�:�3D�.	�:��o �����'g2�'�����U�@��4]�D��V��9����V����� �;�0h�@��dE~y��'��j�LL�"n@�v�e��N=%��]��Q�;�>6M!?�w:P�������'��{�F��Vqɤ�ϸ��YQ5��<���?����?����?��T&��=���0⮟�]��L0�f�7Yg��'��eӄ��4;������%'�PB4o����c��U�j
!�n�%�ēԛ��g��IA�3�7:?��(͖R����"��Y���K�i�`��|ɕ��O��O>�-O����O����O��q�摿����7�Hz� E#{"�'��ɒ�M5O��D�O�'B3SB��LI94C6X��'�b�R7�&�o�Ȝ$��
���9T�/FS 13��_�P��`ɚ2i:$�4E ��4�����4ΒO)Ū�6]�`2�#ίd���sB��OP�D�O���O1��ʓe����8�=��e�b;X� �(�&?��ɀ��']��t���`-O�7��$$���8t�>͂Ԫ���l��M�e�^*�M��O(�C��Ը����<y�=4����bJ�)
�����S�<Q+O*��O"�d�O����O�ʧ(/�,A�n
�a�T�.G�o�Pt��i`�|��'�2�'R�O�Bgu��ȉ|��a�̇]}���
�lڨ�M��x����^.%u�v?O�p�Uf�>	�4� 昘5��$=O>�C�ΐ��?q�O"���<���?���1�hzR(ϊ2xZ�kݲ�?����?�������ߦ5�PCELy��'����hReSn�CC�;O��`Rv�|��'��v��6�f�p`$��{a�۝x<��wk��"�0��+?酯�o=������'a>��d��?Q�A��+W����p6���Ȃ��?���?	��?Q����Od)��ۭ^��ȃ�M<1֌B��O8�oZ�P5���џd�4���yG���B���m�*{;ZA����yb�x��inZ��M[��M��Oz�R&����_w���{�R:�M�6O���y��=�Ļ<a��?!���?����?Yf@ႁ�T���R����U� <Y/O�Qo�hk>��'����'.P�¤�.�
Dp0�N,Lg�����>9���?)K>�|j���ki6#�Z�
4�Ӧ!G�ZN��&����1�F1���M|ƒOB˓|h��b%�Y8���E��
趥����?i��?Q��|�+O��n�$>�P��I�k=�"��ҡLY0qb8��ǀ�O<9nZR�����*�M��iV�7M��:�S�
�g��`Z�c����E�k�x�s�
�K��� �H~
�{�? �=`sl�z�v��  �n<�dЃ4Ot���Or���O����O�?�҄��3���C�ޘ%N�)���0�����(�4�O\�7�$��ԡ2��)	�����˧~J�Ot���O�I�U��6-2?��ĩ��BΙtM�h���3��1f�:�?��!�ľ<q��Ϡv��L�kςAW�@�4�O��l/(��	�	�h��A�$Hϯ �2̠�E�26F��fBL1����I}b�'��|ʟ�i1t͉9_w4=ZF N���!�m�n��e�F�ã`xr��|Z���O��K>Yt�U&3N�� �/A%� ��n<i��i�.p�r�D���cq�X=XR��ǲ/S�'��7m'������O�� `G 6�V�i`-Ʉx+��Or���Ԋ�ش����l��F�|$S(O���$�C�)��'-ڋmݺ)09O<���=ie��h���� �WA,x��ԝuț��q��'Q����Φ�9C�xD�4)�.;��5'�L��:ܴX��F�+��)t!�6mb�H�P��Gt�A3!I+њKE�l�@y䎝��B��b�sy��'ar��g��h��O�9 eJ}���̂B���'�b�'k�	��M��lY�?y��?q��*T���ُmހ"�L��'o��j�&K�O�O� QaR	���siU<O� \
s��(�s�%'����fE�ӣ%�fAן�r��ǐ#7,�Krd�l�I������	��IɟPF�D�'�L���[�0ؑU�X	{��
��'6|6�#���$�Opl�O�Ӽ#�DY�n��	Jv+�d(^�/x}ϓ~����vӖ�lZj�oZk~�LEw!D��ӳh9�b��K�V�2S@ҼmT��7�|P��Iޟ��ǟ\�Iן|lD�u�UZ�� )���wy2�d�d�.�O����O �?���_��]�!ږX��yr�����O6��JP�)�Ӽ,&Y�KG)}w<0فc/�HAj��K���?^ԑ
�
�Ot!M>!,Op鹦J��7X!��
#�����O��O��D�O�<�!�'������8B>�R��C��0էܹF9�Q̓VE���ĀS}�'-�ghӀ�X�VA�.,��σ�D���@.PN87m=?G`	9*!���1�S��)��Í2
��PRjX"/��R��w�,��⟬��柠�	����j���|S�U��)n�XmC�	4�?���?�t�'��Dk/O��o�f�y���23.��bd��A�[��y�O<��i�6=��	�rcaӜ�
�}qq��#!]�����R��<����eb��ѥ����4���D�O��d�.V�p�ڗ@�~ĺ-�!��������O��mě6cҾnh�	��|�O���!֢���$L�|�0�@�'&"��>����?!I>�O�ְ�o̚n�!u Kr��*�j�-^���9ׄPlO�i>����'G�$��A�/(>��7�X�)�cER�����ş�����b>��'��6M>�<,��7�.l���Ԫ��i���<��i��O6l�'��6!�
J7�r�I�W��Ӧ��t�6�Gæ�]̦��'<�s��?����I A�%G�1P���,��P4O���?A���?)��?�����I�,X[,���-�$Nz)䋓�/.X���2T�����O ��=�9On�lz�=��M�H䅀m��z\Xu�����@�I���Ş�8�k�4�y��	Gs\3sL�A�N�S�f��y�U'3�0��	>Uj�'��i>�IEJ��R
�<���!N��6P�	ܟ�����'6:�d��<�"�'X��˃v0�����U74�X�Bj�$.�O`�'���'�O��Y�
 A?$٠7����)V��D��j�I�i�,+�S	NR,�ݟxrq떥A5����KYz����I�p��� ����PG��w�İ	s�A�Nq�2��'l�̝c�'��6-�)HQ��i��4���)��>�v��`]�X9�;O����O��d C��7M,?��M]�P��gP��rG$m;���P�3W���*<��<���?���?����?9��hz����@.�4�#�D��Ă��9 ���ޟ��IΟl%?牺w���{��;(�,�W�Gr�!�O�d�OޒO1�f �@�����cSA�q�d�[��)8>�'̣<�q.�~���䟰����d�g=zYbC��#�,��d#�"˸�d�O2�$�O��4��˓(�e�-ەOg�2V'�x�$�zqj�2�y��⟬�O�Ml�!�M���i��\��R�8"���W-<�<Y@�k�*��֐���	",��$�)��֕󆊨v*��رN�:Oy��r3O��$�O��$�OV���Or�?%R��\� �J5LޡbթE�����I� �۴&־�'�?1��i��'�v,F�Ю;l��);*D���M'�$�OF7=�f�tDg�X�i;��2n�;F�ඁ�Kh���F�"�h�Ā�����4���D�O �D�?h�le�!J��3�ư_����O��8��V�Ӣ{��'�2S>�3�b[X�R���#�)h{$9�bC??	�Y���	ӟ�M<�O��Ā0��h�bAX�k�?��Z����l�/և��4������z�ON0�����p˂�+�ʈk|!�ƃ�O��D�O����O1��ʓ0��蛯D@L��ʂ�7HD8��֦�x�C�Q��Kٴ��'DDꓔ?�4c��":1��Y3x����E��?i��ix� +�i=���ǘ%J��O��g�? �a!O�A�����{�@�&>O�ʓ�?a��?���?����:�P0eC�0�B�YS[��T�n!R��|�	ȟT��Y�s�������BO�FtF'�9�d�15�޲�?i����S�';�.=�ܴ�y2�з�<A���m�X�C �yR�M��d��
1M�'�	ӟ`���`����Ƅ8��J8/NB���ʟ���'l���(1R�'k"�^/�xTZV�$�TW�	�:��?�Q���Iş�&����Q���ȓx����1?�IH�53���i<��'>1��$��?�m�0�Z��҃�^
�� c;�?)���?���?)��9煮� * ���,ۧ�ݕx"V[��O�hmZ�q����'�X7�(�i�I�S�T,#����b��#Ev<�3n����џ ��)!`�l�v~Zwvl�C�O�N�ᄥG<�Zl��A�P��n�L�Ry2�'���'s�'
�FҴ;>���V3P$ ����!eH�"�M#E���?i���?qN~b�]�B��f��\T2 ��p���X���4C ��A3���rުH8��K�"��q�c�.�a����*�	l�Y�Fd�ON �J>�.O��b���P�@��X�N��.�O�$�O���O�<!��i�*Q
G�'s�)�7Ƀ4^2�j6õYr��&�'4*6�*��'��$�O�7�������l��x��X�(��ʲ�Z�	��1m�K~+K�k�z��%)�O��F�(!����`G�e��$A3 T	�y��'-2�'%B�'����jب<�/�5ky���%n�n��O��$�� �r>E����MsN>13ER0?�v�!���%j�c�F 2Q�'$r���t��&����� X�d�x���JC�+��`6F-9e��J�h��my2�'w��'�	�`]�Q�DfV3ۮ���)K���'_�ɷ�M;��$�'�RY>�6���I��g5k>(��/1?��Q����ԟH$��&��A��:D�����9�IyB�l@�UPB��'��4��	��.�:�Od��ψ�o	z}s`��  �q�C�O����O ���O1�`�zO����eR��x3Q�F��`�g��J�(-Q�'�B�h�4�<j�O��~�X�ń�)Aڨ bt�^�i@��ͦ�YA��ڦm�'�h�c�T�?���q5�ח/.)i��CSɒغ"5Ox˓�?Y���?����?�������5{J`��D/�,S*�r �£�dnA�����d�	F��_���w:�<#7�)e�=����&HP`���'�r�|��jfD��6OL]S��N(d@ L��`NM�|գ�0O섒�@�?��>���<���?��%��qT!�4�\�4r�����$�?���?�����Ʀ�:��]ܟ\��Οt� �!���%�<O#�-�Og�P���П�n�<��Tڽ���_.ͬ��$$�3%`��'X�1�!³o8�z"��@��z��'�,x0lκ.��}� �b�X{�'���'*��'��>!�	�t6�U�ٳ;T%�5��r�б�I��M�@�ʪ�?���E6�V�4�6����R�r�j�Ҳ��.J�E�E=O�oZ��M����E'��M��O��R�Ę�����M&$5��M�gh�تa�ɷ."h�O�ʓ�?A��?���?y�!Ƣ`霓><�e�qMӏvGX�:+Ov�mڣ!�|���؟���^�؟̛���r`������*�6�z�����Ʀ�ڴW-���O��)�c�"v� ��%��2\*�w)�O��5.���C%\����D�X�O˓s�ℙ�돸��1k�N����L���?��?!��|�+O�n�H$����]����2�@?xϠ\wbʔ,�����M��ϫ>����?���a�0�BU(�4^*r(�Alڍ^����P��?�Ms�O~m���ګ�!�>�	��~$j_
t�
�ٰB�r@�0�;O����O��O�$�Or�?Up�i1�^���Ĵ
���5Zğ�Iߟ`��4�H�s�l�ߴ�������V4�8��sdP�q\ڠ*H>����?�'j60i�4����t���<wW>8�b@�Y3 M�a�ٟ)-$���������OD���O��$
�ϊQV��5�����7V����O,˓$����gWB�'q�P>�S�g�?w�J�M�X�����@.?� ^���4a��f/#�?�Bw��FzM��
ʳ8���D�/t��X��Rm�X��|����OX�pN>�Gn͇�ȱt�T�'"�=�F���?���?����?�|2+Ov�nڀk�ɱB>rO���Q�֯Ae|��%Kџ����M�R�>Y2�i���N�5Bl��`N(a�T���`�z�mZ�L�R(m�o~��ί5Dp�)a��	�Zd�$k&m�u��A�G`�z�	syb�'G"�'���'m"T>�Ed[5F��X�C�T��������M+��Ȝ�?����?q��D�v���tL�eyWBͬЈ��ҿ5k��$�O��&�b>�r�e���]��H�@ȃ
{����	bb`�;0<�G�OƐ(N>	(O�	�O�%c�/��qo�1� ٬<>���m�O��O��<i��i8>Q��'�r�'R|#�+�6+�d�����������zy�'��ƃ>��V E����/ɍ<�P @� ��#��I��(�h���B��'?�p��'G���I�]���d�M.����܌a��Ο�����It��y�Lx6`�a�-c�PɈ��ȻO����b!�w��O���L���?ͻ�$���]�b�D�C�
�ވ�~��VJc�$Yo���L�nZ]~b��t������� ~��s�?tFV!��2U�� �>���<����?q��?����?��H	�u`����?[/`2��P��d�����5$qyr�'R�O��S2��wЀA�6]:�M�yj��3��vLsӾ%�b>Z�k����+A	W!"�0�C	L�H�e��lyrg�0�$u�I�[��'��IJ3~�b�����T����$3$x������ß��i>A�'Ib6�Q�?�$��2p�6� L-ņ
����SҦ1�?�!T�(��ʦ)��4|�Ԑ�åͨ`u]!�����Z #H����;?)!�-v���I,�S��E ���15�$dyC.�< &��-i���ܟD�	ڟ��I�������J2z�t�j�!b^ĚQ`Ƨ�?	��?I�i�Π�dQ�dR�4������S���Aק,}hTi�x��oӴ�mz>Ya����=�'+>�(�}�2WY�t�Pa���)��<�7�'g<�&�(�����'�2�'�`�7���ڶ���ІvdxT0s�'*�_�����iZ��������Y�D-�N��uc�L�x�V�C�nȔ��LX}��'tB�8�?!x���F>��u�$n6��j�	˂*�����_���|�A��O.	�L>��% ��1�Q��D�������?����?i���?�|�-O4�mڐz`ȩ���&aE����sAn�!"Fܟd����M�ҍ�>��7���u5vf��EHX�;Fs�X6��+����̲���:��Ԝ~J&�=P�<���/Hv0���<)-O���O���O���Oʧ)&�<�)��d��@�GZK�����i��I���'���'T��y�`��nֶuy&�ذ�	�hLhb4���9�&io�,�M+��x���c�T���>O`� Ǥբt�ziiS�(��8O\-�ŏ�?���.�$�<�'�?�a�$4�â��S������?����?�����֦%�U �柌�	��am��[�n�ʂ�<��lr���o���˟t�������XB��8����n��%\H`�'sE�͇n�� ���EƟ� ��'�.��1�F��@S��T��M��'��'�b�'��>睷+Jp��sj�܄�$+vi�Omm�
g=�|�	��ڴ���y�K��RI
<FH_�Ș#�@��y��'��'Uv�Ѿi��i��"T��?*�e�e����G���8Zy
4L�0=�':��ğL���(�I����Ii�29��̕&u�HE�&j�޼�'�H7͑dl4���O��3���Q���(d+ݞA�v�N$xǰTC�O�n��M�$�x��Dl��@v�L��#F,��x)��^�� �4Z�t�C�L4zB�z��ty��M�q�E; %�{�����@��R�'n��'u�O/�	�M�7���?��j�0}V��: �K�]�s�&��?�ҵi�O�Y�'�x7��ۦecݴ7��`iB�� `ջ�O0)Ȫ)2�큐�M��O� {�(*����*�����9���/��, A[*`�|�JG=O����O���O��$�O��?i(G��t_TS��<cjSkƟ �I�����4{��iͧ�?��i��'�ޤ�KD)T�41�F��;gy<9B�-�\ݦe���|r���M�O�9;��!P"Pn�(�̈�w�́�B�
�?)�&�D�<����?���?�@��z��ܐ��1i��ʷ-ε�?������W�Dė���������O��`c6&�D>DȦ��R_`�S�O�Q�'�b�ia&�O��U�����^'7DF�u�R�?��X�݋/n-s�[by�O3X��	�o��'XJ�ʗjGl����&�ďRj͠b�'�b�'���O�則�M�`-�
wp�v��t�~�����vBz�`��?q�i�Oʕ�'��6��#�|��D"��1��Vz�lZ��MS�b��M;�O�tՄ͢����<��I�( ��*Y��,Ԉ�K �<1)O�D�O����O���O�˧F>$8���ڍL�L(��݇` Y�i���'�b�'��O�km��nD�:=~*�N�B�c��ÁSd����O�O1�
9��h�0�I�%��+�n�04�J@:b�X��扸r��US3�'���$�X�'<r�'_���`��$Q�0�i� N*5z��'\�'�R�hhڴ Y�`.O�����)���g���{��� ��W���O���p}B�'�ҕ|Ҭ�1P�4Y�ЍB�o�&�B�ρ����9ߘ�;r���?
������?���Ȓ1�R;ab�}���#FJ�!�$���f9KpG�9{��� �ڜ3�Z�d�	�����P����M���w-aL����" J=u8`���'c�i�@6m�7�+?!:3x�ɑ2ˆd��ָ%}�e��;h| zI>�*O\�?��l�G�D�5&T\8h�q��G~��e�0��WN�Of�d�Op�?�d��&V?�uY�$]�zz����#�6��D�O�7MD|�)�)��D�[��\�z�����T²a�a��07M|�|�f�	�O�4�O>9.O0K�b�e�8թc��0N���Q��Od�d�Oz�D�O�<��ih�u�'� �3��
inN`$�%F�P���'X�6�-�ɼ��DH����M�C��DԌ`a"�R���]�5���4���_�2e����$�ғ���ným���5�D4ݨ�Ss�-N�$�O4�D�O����O��d"�S4|��$Ѵ���!���;�U��ӟL��=�M����|r��Y#��|([L��U��f�Nb�y؀/M�-��O��o6�?���F(X�lx~B([4̀ � B�H�w�JP�	�3rJ�TgJ��?��-��<i���?��?�H�&�b���_i�p�(���?�����U���ߟ��I����OI"и��<�fy0d�� s�$+�O���'C"�'"ɧ�i�1!U�Փ�T���5�����SV��X��H���<�'/
�� ��\���{��L�x�28��S�F)hx#���?i��?Y�S�'�������l�>	l2p3��Hq��Il�+Z���'�67m,������O L��� G��c��,�h�Cd�O�$�l�7�=?�;G��[�')��˓
r��`�l:iV�3)�yx̓����O����O����O&�$�|R��dy6) @$��AQʝsr��*F��+
� ��П$'?!��4�M�;���t�rL�!�oP< |����?�I>�|��"�+�Mk�'�^��caW�b�
T83.�?�:xȝ'v�*��ğ@�|�\���I����i" ���C�M�Q��
B�ӟt�	ß��	gy��a�X�C�F�<�?�rtb�&�D����ҧ�#>�p�K>��p��	��MC0�iP�O:쩖�ҤV1�Y!�D1(N y��ZK��tW�|�6e�U��4uPbeǟ,���	�6|z����'j��X�g����d��ϟ������F��w���U�ڸ~Y6�Bq��!E�q8��'�27-Ŭv)f���O��m�d�i>睔�@b��ߟy�H\� �[q<�	ԟ��I՟T2�����A�u��Zv��͇Z�����j�6Ǆ /oFX%��'W��'R�'�2�'��;���V^�Cu������F]�`�ٴ3�di����?1���'�?���n.��p#Z�0Z��F-�t�	�MQ�iЬO1�-��ǛLA��XWJƅ�xE��� _2����â<��Vr�$S�������j�p]��j	�/�p��IH&B{��d�O����O��4� ˓ *�&C*=rb�?!�d3s���V�|���#�y�#g���L��ONem��?1ܴ^��})���y�<� ��B|Ш����M3�O �����:��/���﨡S�'L���	�(��� �c�=O2�$�O���O:���O^�?��qE�uXE���;FYR�s�����T�I矸�4"=���O:67M5��P'V՜`@�a�O�h�@b�}&�T�޴C��O����i3�I�N6�=�thS2]�����T��̐��^�M�b��O�Idy��'#��'����"";��)��Q
SB"����ܫo���'�I��M��T��?1���?A*��Ha@	�;*bpi��95�[��h��O~	o�?�K<�O>��#U�/������F�%��Xʥ��R��H��K�&��i>%K��'"��&��*��
i���³'��//��z�dV��L�����I�b>��'�6M86�P}pG\u,JI��iʼ7PT �!��O��d@��I�?A%]�(��(�0T�C�S)/8�i�f�%1~��ş�BҦ¦��u�S,~(�f�wyB
�z���υs����(�0�y�P���	�8�	ğ�	ٟЖO�vm�A­,�{1dD<@x�P)c�~Ӹ�a���O����OD���dZߦ�]���Ap`��V�s��N!!�`������H<�|b����Mc�'~�@r��R,�VM��`_�}[�xZ�'�.���(��hۧ�|�X���ٟt0�/�!g]�hTh�)��	�E ɟ|�Iϟ�	~y�p�ʼ�& �O���O(�:U��hJm�'��*C���" 2�	�����O���v�	Ez��4+�� ��5� e�����v�["�]%<e�|�.�O"e���.�Ee^�d��˗f�s��)@��?���?����h�`��Cs��(����+�Pi����
$�D�� ���jyR�f�H���?>Gz��v�E�Q�T��阜m��	#�M� �iݨ6]�*7-(?�F�13��	I�I0��kFi�#7v��ǅW�]����L>)/O���O����O6��ON������P����6"� ;�
!�b�<�iri��'���'��O����1 �5�@�8s&q0�7U˓�?�����S�S�]l���3/ͺ��i�� ?�9Q�L�?�*��'|�z7��̫��|rU����#��9���Śt � ��S��I���ǟ�Oyr�t�|:���O�',=���iv>cn.P����O��lZ]�u ����M�q�'F�挞�k�(Ak���6T~Ei��ڍf�(�'�iQ���k��]���O�Z�$?1���v��|ڗ)�7��#��Ү;H�����I��t������C�'AꚈib&��+̘�Ia��"B�P��?���2�F`����'��7�-�dȧ"6,�!��-RI�aS%A�{��t&�d�I���S '��lZM~r��7��联C�$B*^Ay��74M��kJߟX"�|�[����ퟀ�I�d ���,�E�$�(8<�w&�ßX�	Qy� w�\��e��O����O��'oJ����9_ڌ��n��;c���'����?���zA����I�h,�E�v�[<CX��(/��tYĂE�
fչ��S�e���B�#�t�A�
��W|fT�B�7��Q�	۟��	�4�)�cy�i��PpW"H^�0r!�.0澕r��ۖ(�v�;������n}��'2���V#ǻM�����4�$�'�'=p6-̄$�6�"?�֦����*���F:LB���PɁ�Ts1���5�yT���I۟��I؟��ԟ|�OcD(z�'�H�c(�>^�VjW�m�F�
��O ���Oޒ��D��݌NwMq�5�I�&N�<v�������x%�b>ᣀ.��u�S�? n��p�Ⱦ��i�#�A$�d��<O��+e(6�?�g$�d�<��?)��p�~��6��|R�y���?���?A�����^𦑹B`��8�I��p��O��li1AܝO�"�Ұ
�L��	��M���iu:Oʕ�fD�ژ-:��ѽ, <Ԋ��� [�-�40��E��k��57����ɜ,8��5`�� 7���4jRҟ0�	Ο����E���'���HE!1S,���F97?��j��'��6mXh�����Ov�m�s�Ӽ�T)�Y�u����4$�H�JuG�<���?r�iW��i\���2��W����&7>	��.�70�	O� (T1O>�,O��O���O����O���� ӊ`����a;D�"EZ$G�<��iS�}�T�'aB�'��O`�	-�i�t�
h�e*�T' 4V듣?A����S�'m��\W/�,\���`��T��`RWꍾH�v9�/O
HRh�)�?��,7�Ŀ<qF�)Ox�[��9h� ��&O�?9���?q��?�'�����a�3�A�`؇F1Mr�����D��0IvD�Ɵ��ٴ��'�p��?a�	����= p��D��i�DK&�X"��C�i��I�vT8zw�O q�<��B���%��8�B:ъ�$�OJ���O����O���#�ӹc� K��֌+�c��PP&��Iޟ��ɠ�M����D�Te��O�p�ï�-0ڄ]��(�:{�ؠtb�W�I��M[D��i��M��O�p��/ڈu?L��씜CVX�U�
i�� ���ܓO�˓�?9���?a��X#�iWIO8&�$ԋ�	��-W�a���?�*O:dl�t�4��ԟ��	T�����	zv��lѾ���"�����c}�fq�84�	x�)B��\pXI�d�Y�"t��gAR&	�$U�H�vf�%k(O�)��?q��(�$
0����$�Xf�<"�ϛ(0*�d�O��$�O���ɦ<�`�iR��z�ʎ$fd�)z2&�� �V���Y9�R�'��63�ɛ��D��(d�9{i���n�9<��P��M3G�iU�}��i���8z��r�O��-�'i��`�]"\'�չUʠmߒ���'��	şL��ҟ�	��`�	�����P��g�RyrX�5"ՙg�6��:{����O^�d(���O�nz�Y�֖^�*�ЌQ3m�$i�����M�ûi�O1�v���Jl�@牭{x���A�$EU@ KԈQb^�I��=J��'�D�%�4�'ir�'�Lx9B��q�L	ӓB��xaJD��'%�'"U����4 2�����?���	��V(��d�Q�b�1�d����>�B�i�7]K�I�t�(�آn$���P�g��'C�
H�����I�%O���K~"�m�O�����s��Al�#�P�&��NX,����?���?q���h�����7o��<�aE��/tt���%S�@�G�)���Οx�Ɂ�M���wsXZ@ν���A�%ֹf��'��6��զq�ݴ6��Jش��ˬ>��!��I��r$�C!f<�rD�<����"$��<��?Q���?����?y% V�VLؘ5h'rXS�\��^�93G�؟\�Iǟ�&?Y�Id)�U2����œ�A]��˩OҕmZ��M�x����½;�Ѡ��0�*h("�X�J^���Zd�剥c�*	�s�'4�m&� �'G
� ���?\�x����$@SyRR�'|��'�"����T���4m�-)��#�r ��#n�6����w�h!1��#{����\}��kӞAn�M+S�
�z�B��'��
GS���A�PR"�Iܴ��� `����'9d������v4�i��K�^���F�8���O:���O�D�O���3�S8n�E��I]t��	�c�$#Ѝ�'!�i�hh{�>�����˦�$����C/(@`��&[|���\.�䓈?���|z�M���MS�O~���!I1j�b��O�^u� c(؝"֪���)��O���?���?!�k��jvaЫp�Ȩ�F*�?D,a;��?�.Op(l�F�b��I��\�	_��(�#�z C�DP.*��뒍ΰ��$\b}��n���lZ���S���V.��У��p�����\�ڹc�O�� �-@RT��ӹ e� �C�	#F���%$�7K���1�\�Mh�D�I��I� �)�~y�Lx�f��	��R�"�nɂu�|;�fH�j�H���O�lV�#����(g�+
�ȐѰ��W���A"��쟸�I�>��mZg~Zw������O���'�B�2S'��UZ(��&�'m$�B�'v�Iڟ��	�����ğ���X���ĞhC�0�`�Hf>[fG�D��6mD�m��D�O���7�9O��lz�q�C��uڞ�2($ S���uo�ɟ(��n�)��-S��n��<�c�<�:��V�J~hBQ�]�<!��Hd'��d5����$�On�$@���E�/� h�-�M�����O����OʓTn� ��?	���?a��ʕf�������:��܈����'t듖?���>��'�!�1�=j-p��IE�#����O\��%��)SPK��i��?1�,�O�XD+�6*,��ʾ[윍!"O��ū��U�C}��2�b��'��i�"l�r��OP�D���?�;��9@��y���@#I91L�$0��o�.�lZ�
�Pn�\~2�ƴr|�<�4�Z�K���22,n��#)�jl�m���|Y�(G���1�0�#��4�q�f% �����黎Ra՟<�	ğ���b�A�%�^�b�oQ�سԨټ~��	��M'�i�O1�ء	'� b�Ҡ��;Z80�5��9��Mƨv�˓5���L�O4�!L>/Oxu1 ��ӄ٘C�ؑ��HD�'�6��o�p�$�.]����ũ��:�Ҩx��,¤�$��-�?�Z���	ҟ@�	�`�i8�$ՏQ`��Y�_�Sf�p�c��U�'�>$��f��?	Iu����W�U���sad��uM��c6�֌5�`�ȷ	:Rn�&3p������b��p3�g��iu�`���ӆ!�0�6,5�@��ƪ�&��X��b'��!"$Jӥt�V���ʉ# �E3�9�V�0Qj�C47|@��fl��D J"a؎?34Ӄ��{�����:.�Xr F>+D0 �o��5�
�c݄k�T1�؎S2��� �!'|0�n5o���e��ج�#C��N�c��݄O
�x��@0����f�c#Гw�܅�LM{�7��'#�|�۴�?����?��#ܯ$~�On�$�����7m���������b��/�I�M��c�4�	���&�E��@�4ɘ&��^d��A�-��Y���$�f 	N<���?AK>�1')��X�nH�\� }��ђ�:��':��=����?�����ۓX��CՎ�`wl�!O83�]��M��Iڟ��x�	Zy��ƞe�Т��
uT���v~�p��y�'I��'��ɗ%Y:X��O�h ѦI��&5 D�@D�2+�(�O&�$�O֓O$�Eb�'(F�t.��U��,; �]�v���s�O���O2�D??�����ħ��!�bH����Y��.Q؜iKB�i�R�|�T��$�=�I�(zڐ��H�+5��!bU�YI57��O����<��bIn�O���OZ� µ�[� �ґU�7�T}���*��<)���f���)_�R��sV�C$�� �����P��iUGP��M[UZ?1���?��OHMu��"ň!J�W�Ƽ� �i��I	����?�g�%im���O-"���0V6MȒ�Ddo�ן���ş���:�ē�?�CN�A�(2t�ʶ	{�(qc1�v���O>	�	� �K�i�I�`�	㊏�@�$��ߴ�?)���?Q���{��'v��'�����	�v��!�(�&LJ%��ʱO���C�$�O����O$�à��k("��!;���ɦ��	�&��\+�}��'�ɧ5�#S	�����*f܎�h3jE�����(z
1O���O����<���\�ml�nM�g�Bu���� b��񘰐xb�'D2�|r[�ȊF�O\����-B�ĭI�f��&�c� �I��	]y2F�a�����BǗc����eT=G=ɗ#�>���?9K>�(O���\���"���a��"N,̤���>����?��?���t4p���?���@�V�ڤ�	�~�Ƥ�pƙ�Yt:!8`�i�Ҟ|b�'�b��7^�0�N<	�a�,����j='Ęp�զ�	̟�Iӟ��$C����џ<���?BSNG������Xpb�L��h�����?���01�L�I�S�T͞�M��؆�E�>�����ז�M[���?q mڑ�?Y��?	���)Ok�Z +eL����_�u�P�Z;f3�v�'��	8u)$"<%>��p$�:ྡ�'�	b<�0Յe��Q�P��O��$�O���J˓��)B�{�P��\�+6��:����Q�|��*9�S�'�?�0DJ�cTdR��F-}�M!��# ���'��'��I��h�>Y/OZ�������Ă �RU*��A��X��+b�ΓO����VD���<�	�4:a�
�|)FJ�	I�ZE�U�MS��;���qY�Д'�Ҝ|Zc�~@Rvb�0+b�b�V���H�O�msQ�6��O���O������AS*L�R46ϴnh������H��qy��'��'��'D�C��ƺK��A�5	NGw�\a�jv3�^���ៈ��{y��L�FEP擾!�� V�76��%����6M�<9�����?1�y�(�'�Ȉ[��$�����@����O`���O���<A�C͑j���[��6��A4��&`�h9f���M����䓴?��b��쀋{�)Z�t�ܸ���$�˵�
	�M����?Y)Ox���z���'�B�Omҥѳbޙ"�J��p���.����&n�>q��?���90��q)��Ix:�-�#'�0����5U�"���ߦa�'}��ӧ�x�����O����$ק5���8XE�$:�`S�[ބQ��͂�M��?��I���'�q�Ɣ���5Ng�i��) �m�D�R�ig4D���l�@���O����F��'�剳V�@�	(�:�����L��P �4��X�"���OnAx�!E(|~ �e�V�$뮴a��Ʀy�	����3���ڨO"��?��'T$ e)�*r! x�cMUs�a�}J��'�2�'�" �S5X����[obY�	NV�6��O�P[�͛l}2U���I�i�Y�ց��mZH��W�2�`�3�>!F
��䓖?A���?�/Oj����xB�)`b��3ކ��Y�����'��IҟX'��	ҟ���� �u�XQh��2���"ƚi?>@��Ny��'\r�':剤Ob`��O��qBeMG�4 ��K8C^\޴����O��O����O�7F��� �(�_�<Z�#U/�2�>���?Q����PTJ��&>!���{̻���>�6�&K.�M������$��L���D=�Ĩˇ��xk�U�D���
�^�Mk���?!(O@�[����@�s���D!�t�0A"��<d�)(e3�d�<���5�?I~��π <�Sr.�3we) � �4���ٶ�iK�ɝm �޴{��ٟ����d�Z`�`�LA+X�0}��Y9�V[� 3�aPğ|�K|�M~n�t)n=s2��l�h�i�A£1��6-�AO��$�O
�d�O��i�<�O(n���Ә]�v��&�P� 
���0�b���p���.1O?��Ԃ��,o:�Q&�/1�K��ݾ�MS��?9�ꬹ�/O�S^�D��2���ЭII]�A9�k�(4����<�@S�K����䵟0���X�q���-��5(@�\_�&�'�vѸ�U��Z��N�ૣ�Q��k�$��3~F�"�������_1A`
��D�Ob��?�5 vb�Dp���ft��Ic�B�lB��i/O��D�O0㟬�I�أlҾ:b����7cx��JC"z�P�I"?���?����䘄1����'m�]0��ڒ<�����Ε1�~L�'���'u�'��I�0�M�ɸ0@䡝�~�
 �D
[�(?�Eq�O ���O���<c�p��O� ���3dX�G�π!0�z��s� �$#�d�<)� ,�?�H?	IA��X�����o>x���u���$�<��q���.�n���OT��Ɗ)fLO
T+RɈ�V43�6��s�x�'g�K��:r��y���	�$��Y�$�C�j�*���#��i剆j�Bp��4S��S쟨����䕵h�<�kC�~�`���B- ��]�L17�����L|�O~nZJҾ`��!6�25'�]R7�ŗ�]��ԟ@�	�?YIN<�'h_��q2�n�+�N
�7#���i�j h��'h�V�4%?�9Ӹ��L�CA:�H���;*K��Y�i ��'��	&4*�)�N��Ҡ�U<�p-�'��-5D�i�n���':�}�3�.�I�O ��O��JԮ�3d�.*����x��G#�y��)"�U�H<�'�?�����3��YK� �,���(��97�o����IR��p$���	ןt�'�Z�⠥�y��Q	7 ��Y��B���\O.���O`��<����?�f�A�wN�y���$�𑁵�U6�����ON�D�O�˓0�䑁�П�h!@H�,�6�`��ȕl�����4���O�ʓ�?)��?q��<�B�߼}����Ή�1Y���ˀ⛖�'92�'��S�@;��"��)�O�r�ᇦ&2hHd���9���Ȧy��Iy��'���'$��y�}��OJ*�YYP���텂$ZՒ��4�?����D�~"]�O^2�'�����=F�f�����-h�}��Ƒ�skN��?I���?1��h~�V����G"� ���[��ق ���R�lZXyb���P-�7M�O����O,��v}Zw"h@"G�/]��1���j���ش�?���~�t�Fx��)޾-ڸ�'!��$�x�mT�, �f���"6-�O���O���D}"V�h�H�V|��Z6��ծ1��@߬�M����<Q�����*���DhƊ�x�VL�7C�"pyЃ�M;���?��v$�4"4_�L�'�r�OX�C�R/zutA�B+� )ZF�jýig�'�"@����I�OB���O��C�
.J�%�JT,S pJGO�-��Q�@i��O4˓�?I*O6����(���(m0u1s���* ę�X���'l����̟��������IyR!B�[H��4/� MĈ�g�]�V����>)*O�d�<!���?I��T�è�x��|�炏�v��XH�EX�<�/O����OF�D�<��"ǅ`\��8L4��u�4n��9��O�@C�6Y���	uy"�'���'AĐ��'�h��X�<
��ҡ#T�H�m�p.f�<�d�O����O��mm��&Z?��i��˖�P�T�*=��Q
�y��aӐ���<9��?I�u�ϓ�?�����q�(��tѓF670i9��i���'{剃 ��q������O|��W�~tp|�Շ`��Y�M=.���'���'�B*���y�'��TҦ,F�f�̩B�A�h��@��d�ۦ��'��<�obӠ��O����@ԧuw�
�x� �� %�:I�V�ђf��OP��
U���Yy��Ɇ�[.<J������l���7�ˎ$��o�ߟ|�	��������<y��B��L8�lL4I�Ʃk3�W!ϛ���y�Y���a���?	&�V�>:��E���7u��9R�HcR���'���'��a��#�>�-O,����L��_n:L�*�J�� �<���d����<�#L��<�O�B�'	��_�-w��ڇa��v���ä�3.�6��OPA Ů	p}bR�$��Wyr�5F�LL!��ſUn�$qEɇ��$W�4��O<�$�O��d�|�N��vKp�����Cj~D�#����Ny"�'6��Ο�������H;YhS��ү0�&�S�mǢ������������8�'B��1Ff>�S��r��i��"�6KF��'!�]����ퟀ��e}0�I�R�P�aP1��;a��9҂��4�?���?����8bl\��O�Zc����K�%��,�1�ŷ@��]�ٴ�?1-O����O���W&ft�;}�A� Nu�<ɖ��VXc�#G�Mc��?Y)O��(2k�g�4�'�B�O�8�1�M�[��}CW�R������>Q���?���.�j̓�?�)O��?V��CƊѽlV`]�AB��6�<��)A8_!���'��'�dD�>��i���P�˗.hfH���	n�ҟx��0?Z�I��$��˟��}��M6��h���":ܸ�d��;B�>�M��?�����R���'�\@�D���Lk��O�p�)��{�^da�3OڒO��?a�I�� �E��K@��v&�Oʴ1yU�i��'��"�&W������O��ɜR�%
��A?���"�!}K�7��O����OJQk@=O�s9oZ��h�I�dq��d��r7:Л'�]<b&|��4�?�%'��'=��'ɧ5�7
v�
7�G�i}H��������!:�<����?������ΠG��a�"��q[���'�,R8~Xa�W^��?iM>	���?I��I�u���?��tc��n�T����$�O0�d ����9jXΧV�)`��l�(*�
�sC>&�8�It�	�<��c��	#ѐ��giK32�̀d�ܽP����O���OJ�d�<)3U�m��O��)	vf��
�Z��`��� �����Oj��3�$�O��}_�0}�	>V�č ���QVt��.�M���?�(O*�9��k��۟t�:V!(�Ҕ�*Oy��)�P)�U�M<����?�B����?qM>��O�"|1a@�x%����@��YH�m��4��D�#۔�nZ���)�O�I�l~bGL�:�V�j�쇩z�;��6�Mc��?a��N��?�N>9��$�Ȏ"0R��ǜ x�P-��M�$�*w���'�b�'^���.�d�O~q���2 J�<T	�����`7-O'l3�D!��'���|Z��!4��AǄD�f�4�C"��M���?i��x=C��x��'S��O&�9t��Dr�:u*K�s� с�� 5;c1OD���O����h+��!cɷf�(a�\�'��Yn��B2n���'�җ|Zc8	C�K�#�ؘ��Ь/���O8�f��O`��?���?�-Od��2�!�J�0�/ǲM��	頹2�\�H<1��?1H>9���?)�d�-x��Be�5�t���\,y�v-Γ����Ol���O�ʓpi��p<��u��gf���E���D� 8c�Z�,����`&�(����<i�q��:�
�Vh�ы�¼
J����	���D�O��d�OZ�b��E�`��T�1Y4��f!�])�(X�ȋ%:�7�O�O�$�O���!%�I3,�����gX�3��p�3�K�b��6�O��$�<�4�Tu�OgR�O�����%G�6ͻE���p��s�)��O���F'2�$1�Ķ?URj�*CDV�SB� *�p89�f�H˓	_�T���ihj�'�?��E8�I)R~��阂U�4=�ѧ�?jV6m�O>��-T���-��|Z�'KrB�-�(�������;��y�4�AJS�i
��'c"�O�lb�BW�%���1�)��cB���5����M�N�<�N>a��D�'Ӗ�ї.Y�? �9�X��p��}�B���O$��0U�r�'��q�d�|Q�1Rdk��=�@�"�N)ZЛ��dt�Sӟl������0�Q��Cz*��$GL��M���޸�T�x�OuQ��0�m�$Y�\����M�4��i?���O�ʓ�?a���d�OP	A��Z'Jo���#	��9y��P��¼$���D�O&���O���:���O����.�T�趫�3��r��6MDj"��ҟ�����'gz���o>�B�h�:"�4����&�@����.��O��Or�$5�	�V����)�W��C���F����?���?)-O�����p�)vj����'c4�I�i��}lz�4�?aL>����?Y�%�k��@E��CJH�"x�C�E�"1oZ����	DyB/�cH�������`Ey�� 7�����
�,9c�l�	՟\��#:w4#<��Opj�cCHթ�N ���D�ag0��V (}�o�<��Қ��{�\��� �{L�\b��y��>- ř!!�?F}F���CQ$����!�f�Ô旎5!<�1�X6HQ�P�5RU9�RAV*��5@lӘ,_n�k�KЖ�P�b�+��]h�bˣp�,=ٱ!25��j؎ ��6N՜'��`�7���� aH���媃#��$�dJŢn7ء����a����D���{^Tl�Iݟ<��ɟ,�Xw�R�'�IR�"	�@�0�91-��4���ȆG�<C�D���΄�n�!������7ʓPTD�c�M�8�z���-��RT���RCE	��T�Po��_�"| �c�x�7�I��Y#��j��Ɇ�L8D��	�0<����O��=*OJ���� �~ဗ�e[�
C"OR�8�(w86�����/�X����v���I�<	�H\������kKV,+��.O�L�V��n��'r��'��J��'"1�r�2E-���ԍ�	q�v0˶�/u�8�Ӑ��+H���+<O�|rM0X�؜y�bL�6�[�ʕlG��G�nI���?<O̘���'{"��E�n���h��i�JU��JLm&ў�D�C W'�ɛ���gN�] ΂&�yR
�5R��%�^n��l�/�y�j�>i(O���T��B}��'���Z Z��F�B9a�d�
�%Fc��Jb��۟�����DE;��E��Q���2�S�tC[�7vI����)k1蝄�(O~���ֻ'm�ɱ��.���@���Ǘ 4h,9���/ ��2剚 � ���O�?��&�}|�9ʣ �b@��ne����I�1@�Iw@����ūn�*����R�.Y�D�8'i��&�
t�RL��7����*�h�O��d=��@ӟ�����pH��߾Q�����8V,���|�IbVO�1Bk�jd��?�O�1�
� �y�*��G�8�Q�H��8記�� � d7l^u�^=�HG  �&���hE�q�q����4�bH��
�
O����6!��K��'Cҗ�����O�Q��	�"+{�,��f�w���a"OHy��d�� ��S!���n�<���I8�HO�S*@��YbG��hx|�)D�R>P����Iן`3�1v�.��I�4�	�)Xw��'"�է;WܦL2Ԭ�<�8� �'}i�ţ�)Qۤ��$G+O�qۖ�ѻ�LI�&ɞb-�;��O~	����,Y�(�c
�A8��3.ގcO�쫢�N�L�#�ĵ� c���O&�$>ړ��d�*ȶ����\��e�Ƥ֮>�!�݈aD��Q�'�b� ��*.pGzʟ*˓)à�`%�i�^�Uh�PM�	͍���s��'�"�'�"��w���'r��+B�'��H��hA;1n@��T�<��uI�w�<dj�#٭��d��˖�Yz,�r�	/���0�O�D���'��J9�X5��Ȍ.i��z���:m�6��O˓�?i���S�t�jӶ}"�d��,Y�	!W��'�yҥ�mx"	�v�	�R*��A��:�y��mӦ5may䉍~>�7M�O���|:��^�=����#��>`�j|xJU�?*T����?�/����iv�'_哖-6����IX�i��)ha,�:D�<�"e�A��4§)b�k�����C�(�df@Dyr&ā�?���iT�7m�O�˧"$epd�|���ED�-Tn=h�������Ğ�_�@Q�/UJ�.��d�������A{ش�?�a��-O��ed��:�JL�����<����\G
���?+�t}�c�OZ���OdL	�ސ
�i8�k�=��H�H�t�ݨ�Q[�|����Cz.A3A��H�i�!�A!uL�9���/*�|���|���'?�Kq��OH���i��6��l#���r�'���';?�$�4��e�CKP6�ڼ@VD_����O8���s@���x6 	�M��c��J���?�bA�F64Z2����|d|I�S�ݟ4��r���J7������I�h�I�u��'3"��I��X�@L*{F�j�.\�G\t��G.:���F�H&P��y��hO+B�X?,"2d������2����O\�.�� K��p���xh��%�ZID��#|����n�"��c؞d��	E�W�L��::��xs�a$D�,��P>R~��� ��2Q���� �HO�	?���Hh��m�>WjI  cN�c��x`b�H�[`���Iɟ��ß�0u�
������|Z�Eן���2rCx�
��,}��b�aS�[����dQ�{U�I�MB�M�f�[$T������`�������'��t�Ϗ)�$��f���X��'�� �(_֔ �qmǋ�J�I�'r6)rR��7G��pr�Y$�rHk�'�v6�(�S�O}Z$��O�1�T4@��2 
� ��'|<	��`XV��V�H'MF����'%4�)���X�M��ǝ.<ET�i�'gr�AlD&02(K�#�D+P��'J]��
F�&-�T�ٓe� A��'RyY`D4�rs40^ɼl�ʓQ�1���,yT�l� �[0xJ�y��]��@��
���P@�*(|l�ȓtzF�DD��PA�&1��ȓ�  "L�*i��d�4)Pqq�(��;�����0p�n� �	��4o��`r.�KX(����İEN>������@� �	0ѡ��)ȁ��X�t��ch�*�G��}Ot��ȓL��\I� Es�*�á�4d�`U�ȓ"�}�	$��̲B!�<�|��ȓ3��ŌF�\ z����ԅQ�8�ȓ�
H9Pe��)A��� N�>�r1�ȓ&���i�I5d@��.H:l=�p�ȓWb�yӥ#,a�R�Y ���A�e�<a�95��lp
_E���:��N�<�I�:F� Eŉ6��8�Aďn�<)�m��x�dȃCΞ�2ҁ�F�<���H>2����眡� �ab�Y�<a�O�l��N�?�(��oFT�<� �`��X��.���,+lD���"O2���H�7*P)�� xX��"O�d��!֏N�ȁ�Ԋ�| �i*2"Oj�9'"ϣ7�n}rah�$;H*dʁ"O���I�p -��� ,�%��y��)rv�KR	B$5ֲy���	�y��='�V�:�eP.;��7����y���sX�AC�� �腒�M
�y2K�5h�v(�� �E+�B^3�y�䏰r��T�g� +_>�J�և�yҪ�,#�0��@�
6A2�Z����y2ԇ(u�Ū�`b(9��# ;�y��Bk�@�HP	$:��X�M���y�g%��ˠ��|@e����yR�N�B��e�v�,R��\��yD�#��(pdF��PtrW ��y�N� gdQ��`����	��y򧔫v������/K�x�XqN�F�<�NC�DJ� ".�bX`, �Aj�<�'��f�$!�3�ْt���
�Q�<��&-���A��
g��DHp��P�<A��6f\���#b%\{��kgRq�<���F�?�6h���}�ze�j�<񂩀{4T�!i�~%��a��X�<�b�K?�� ␁=f���`D�y�<1 �Z���ʃ� ���qS�_n�<�&
�jf�]vKD�
����D�b�<	��Z�DZ uYi՛Z�V�XQG_`�<�L�,Ω��I�%d�<Y�j�F�<a2�ϾD�)8jM Lj��E�<96H�/_`���GM�6�����l�I�2����9Oba)  �1K_�zT�ͣ4�"��' rAi�`T:S��mc�)O#%:&��X�V�s�O^i��c��v��E����D�	�5�n`��
V̧]�IzqC_�	H\����=(�8�ȓ;L���O�ќYڃ#�4�*4�'�F������|������tw��/ ^,��A	�Y�!��03YD�{�#�'<�@E�7'J-Q��'�Pe�'K/U�ax���N��P�� c����?����l�H�!�z��j��a#p4S�nɄ�x2l�T�3�Ҵ'4,��Ti<�0<��F�e���<y��G�AK����C�h�A�ZU�<Ѫx��}i������UWfS�<�b�#o�R}�� ��t��iC�L�<��@;^�-��n�E��p1�	E�<YG�f�X�Z�� �L`��C\�<񵮞�)�.�Z&;�d�B�P�<ٰ�F�t�	�ufѧ��0`VFPJ�<����$!p��2��!ظ"OI[�<��o�s�`Ճ��[$�BP�Kn�<q�d��]�̈��PI
 BA�<i4		���|�����,�V��x�!�
�d�����+O�'�u��-M!��?!�rt��F�0殽��*-@!�d�Z�D�s�I��9s�IEC4!���|<u٥DF��Z�;��U�2!�d��s�����O�r�8� �ND�!�A ���T���x���*� ~H!���<���f���ju,��D���7!򄊯HZA��(�gfz�y�H�$�!�D�%,� ʅ�ӖlaxTE�5�!��@DV�e`v,Hq1�k�DҧC�!�_�~�D������Q��>p�!�d�#@����!��=:(9�ւ��Qm!�� �}����~�dUD�m0Z4Y�"Od	��8Gv`�͉� �~�`t"O�Y�e^�@E9��M�=�n���"Ox�������$eY�+��*y �K7"OTy�g�10�R��f�B-i9���"O
�pIݴ(�(c'�ʎOD@�ñ"O$���MR.r���0Θ'
���"O�Ic��ՑPZ�P[����!�� Q�b	��Dλ/|I����!�D�eq�PkQ�#j2���DӒ'B!�D�:{Wr��hF�*���-ւn>!�9o7�8�6����y��m��9!���^�~,���	AM�� 3����!�d�?��x��P�F���#�!��G?G�*<�Q�Z>���BG'�!��ȩ
6�T�>�H�1щM�q�!�d��(�0�c��X�x��?�!�d�V_����ϕq�q��F�k�!�D�ѫ3P�l�DQ! �Va!�U1 �1�`E�O�9R�F�+�!��72<x=0�nG��53J�d�!�ŧj"���"�6>�p-�N��P�ĥn2�g"0�9�g?�d ߯K���a�ѹk_�)��p�<�QML�'�rI��!�<�rdZg�ğ�;�)�6hB�p�'o���4��T����m^/L>Y��x��Ղ����yg�6J/68tÐ<�q��M�%�!�Z�'�����}�c�(c��O�Z�W�HG��{��	��P�"�# D�*5���"���	�!�$*���e�dU\l���7��:�HO>�h��Y��b�Ffʼ7�t�ID�rG�5�a�'�=ːN����"��g�1�}���'��Bk�(y6�8*��  ư	�FIS~�$k5I��<�a�G�i���0u팣��`P�]#^&�'��@��LA�O
��i�'�-�e�=0��4N�80��I�'���g.�_�TD����N�1dfA	��DU���Q[�Gn��c&�M����FUt�1�K
Dj� A�`9"ayb��T�EC��>�%`�4SMR	+fJD�BM��)F����f�Y
!EL�jR@Ёi12Ć�Ih��$)���8V�d���� v��1,��
�Al"����L<�N̦Q�\���̎F�ts1m��|��m	�'����b�M:�ܠ0�V)�����}�֌��q6BI'�h�Eﶟz4�~�)�1L��#�L�f�K�zQL �O)�5DQ;_}�2!��;Zt�$y!mֈ �(�O�%{%�O����π)��РO?版"�J5���X誠"�=N�?��"żn�0�a���� V���T"L ���F�g'L>���L����'�� ��'焱��ߨO�>�ya�Q�5��,��'�ꭺ��B�S���C�*g������� �:����5 �(A5OA�R7��{�9%�S
Op�;G�%��
D!T���@��S��R��0�@4����\p�]��S6��4XP����N��Ι&+`xY+�!��鶸�@�фF�a~RhC�h�$yA��=H&�Ȓ��06��!&�%s<���O0L�%O]�����ɐ��p�&դO4ݠcE�z���P�.�e�
�A��������䚦�K�"�(H����-���c��K\���)N�W�P`���Y?�za��mڝ�%{��'Ѣ��o.E�.\�Q��iW�5�'�����Ӈ�<�rMM#Q��c!8�]�W��#����+a*�x��XZ�Vm���	37o�!��2��yC�_ �����G0�p�@�l^�w�������@a9 �v�PG�]T+:�H +�7�DD��O�kz<����}r��Y��'��9�*�? YAS�E����yA!�?f�2�x�&��$�*|1���܃h���&B�&7����'}�+H�]9��;s�Єo�ɻW���Oh%�3#�1=�0ؔ�ڒU �q|�ړm�'s�^��#J�A��Dj3N$f|1��M+}"�1`�\�vc�@��	2�*�I.�)+tn�&H��牪ā����o�l�0`�)BƲ�)�E*Nr�((rb�>1��ӜO����t��&|��Z/D�8���'a:q��OF�<�Ĺe��]������hxd��%MQ�N
��g���$\>I���pTĐ^C`�λ]��%㕧S�a��Ҕ�'�DI�5#S�x��!��H����Q,D�g
H]�2��#��N�0E(#sAӈ�E� *
j��W�>��$X��d��ҒH��b�'W�$K��g5$AdJJ2A��[��Q��� ����� r��\Sbj�>b�h{�f���"�c�e&�|�'.���p<Y7�| jx��
�{K��;�`�͟�������Csg�0g-��fu8�����%�I�W.VݸS	�1u�%��Λ�k�^�z	�'�
��熔��t��� ��(Q�����(9�H��!LF��M3-� �3�6 �Z�Z�p�*�fE(�����I*���o�a� �̾|#����xu$)�N�! ��@����W8�0���(Jgd���P�~���W�'��,���Yn�3��+��T�'%�*<��	M�h��� L@�2@��V�B��&��x�N@A0��!H����ɘn� �	4D��0�VB"~Z���>Ә)������Vc��y���@��!��2,�)[����Hhq	c
r�DQK�>���Q��Wvp���I�G;v��ȓS�I��Ƅ"� �z���%s�D�n�i5ܙrE$�O��xce�<#]�q� C���8Z"O���@�4:,BCG�
I4x��"Oҩ���Z!H���A�l2��
�"O�h*$J�$�ء(�.əC�F�g"OX�b��/9zP;���;z�2���"OJa�'��Rv2�S��V�|�)V"O�-9 ��2��8E+�A�܀�5"O��&��;�8�P`�o���2V"O.(�q�C< �H`a�#H������"O���jM�G�ݐ �ЋT!�ӗ"ON�!@��rT����(; ��б"O������DCBd��΀8W���"O(��)L��� KA]Ӫ	�4"O u�Ƅ�sz^�0@jN#5kz��$"O����-Nf�ɩW�@�!�|�C�"O�����6n�~5#�f��Hp�c�"O>U�`o��p�VEЫd��1"O� �ă�,�#㮒�U�u�s"O�t���E�N�[��4!�@��"O������V4<ȅN38��0qa"Op�k6M�-J� ��B��s�X��7"O��u�@'Gh��r���C�ZMx�"Ory�e��1��5r`]�b�ԡ�"O��b���M�00��$f��p�"O>dK�dNt8���oU.H�<-��"OJ�b)��[�$8� )�PW8�bA"O`ă����
Z�eYg'@�^%�q"O�e����^�������;:
(*�"O��yD��|j���MZ�tZ8��"O�7�٦'2˒,Y�0:�"O�pI�NB,
v �`"��a~rA�"O*VH��������)S!Yk�<q�g�%��%�'X&��{��M�<iD��8I�H�#��D��!�&�M�<��F#(4�ӓ�[vh�K�<I�g�x��t�B �Y<�D��
I�<��T�Ew>\Q'�gDLU�Rl|�<!򧍴A� ��AH�%�&KJ�<��O�T��T�q/�؅���}�<�gN�j�h0���ϸ}��Ia�y�<yu��0(>@Q��>Iծ�aciFu�<�FEQ�Z`�T��g�%I���J�m�<�r,š:��h��CL-j"k�<�F�ܮC�@�����`��{�a�<a��S3�����i5p9[q��_�<��KI�nݦM0e��-6Ūdg�`�<�:p�0uwT� %��Z�<����|�)A���E�`t
��5D����Wh����}��=1�7D���̍;q�����_)���c8D�L:��I��(��#�3�V���*D�� ���L�9\*d��'��(�� ��"O |��Yk�a�`�:^2`�u"O~p���cI,{�oQ=Zt��"O����+G$�P��Ζ�<�,s�"O~$Pd��?���q%MZ�u�� �"O�"gg]b��Qc�MZ��!"Ox5Y��0���Yf�7Qj5{�"O`���=0G0RUi�#U�I��"O��P�H-U�����ǭHA���2"O@��d����H9�nˆd=L�)3"O �y#J��
��ૣ�.k3�(�"O���Dɛ�~�h�GB"w#�]�"O(;c7?��e�w�= �"O,@�B�Qc�H�F���@ɓ�"Op�2lˣU^�� �K�d�2�:S"O�Ȓ֠ۍ{���Be����p��"O@]P劍*p��)ꡪ
�?ڙˠ"Oޱ ��T��Q@Pd�$�"�"O��Ӧ��6s�(ѡ��H���ȅ"O�����N��*����Cy�!�V"O��2̏z�T���Aöwup}�G"OT����:\�%���>id�<��"Of�bA.I��m���H�Mm�\�"O4 ��!��MΨ�U�:iX��у�Op��D G^f\��'�,�c�:z�!�DX(7ᾬKa$�i޼�I��*>!�$�����ϐb�"�G�4!�$�L0�
 ۔4n���P��!�*;'�y�f���0���S��֌%�!�I#9<*�Ҵ�уN�����.�1�!���9�x@��ƻm����tc!�D�� D��Ib鞒���ۑ��(~�!���:>��$�;��ȓ��..�!�D�6��PA	�b�zTi�(jp!�^�\y�Ybs)���>�G_&nY!�$O?�AqRS7f��q�&@�.Y!�AQ"`��`dӳz��9Hp:!��Z��1H��<X�F�A�:!�ˬBx2DX���-`�E���")�!�D��f%���Q
46����]#�!��n���S$w)���S�Ip�!�$Z�:�P%bJM���5à�C�<�!��I(:F�p��P'*�]b��T�
�!�$�)��Q�6f�D9$Cٷ�!��?I�B�qB�|ڲu�)I!�D�;$j(m����<�(i�$"�bN!�D+e%:�#��	�h���bg/!�D�]��\�E�E�q,���&	L!��]=����Q��S&b<Ð���*!�w?��[ ��?h��������G !�Dd)�Uq�c�4� �)�kG�U!�d=��eȨ8�$Z3j�:V!�"�*� ыߩE>EQU(�6_!�Z�_�0�1Nkz�y����r�!���><�ASd�CD6���Ɖ+F!����5�pa��J�<UH$��	@!�dg;����I� �P��QdR/L�!��[��� ��y��h���-.���mݱ��R�OCő!)�9�y��
� z4ږ���TJ-Ʌ��1�yb-��cg���D��*$h��ir���yb���|K����j�$+���K�����y�oؕ`����
,-1F0#�3�y�m��	�\ xâ�2�ݘRb��p=ɏ}
� |�'�ؐ��l#�ٱ
G�!�"O�A8�n��o~$�9&�ɪg��4x�"O�Գ���s�\X��Lt�ł�"Ob�Jd��.2�<9���}g��A�"OZ�u�-�6T��ՀxVyA"O���ǋ
%a�mA���?-�Q��"O�IhY�����L�K��`x"O���e ��K_��R��*P�x9�"O��Q�ԧ�T$�aE9P~6<2F"O�qS4lZ$�~-� fz8\��"O@�I�1�9�v���m>���"O�U(C	)Gńqb����QU�!`S"O���a����A#����ճ�"O��R�hs*8�!i��*���u"O���@��Q���r�ū*bQ��"OFԛ���\�i�dLN�PASE"O.�gNƀfX��F�ϬM���"O$��DbF�=����'ϳ+  ��"O��bG\O�q�D�J�ze��"O@�a-�rvIYb�)����"O��	b�~k X#G��
'ѲY��"O�`�/��T.��8chU�%ꀔ��"O$
թS��>)h�!�,ָi�7���OIJ�*1e�/M�p��;^�Z z�'U���C������P�ң_���:�'N괸D,��q��%˗i�_�~(R��!�S��?�U�I�S�:}j��Y�=1#�	n?��]t��m�$dN�5�ʎ�za��	,�t:r��=�f\�vݳ�^H��CI�E�V�E4�#c����	�'�Ѕ3���MCj8"�X���k	�'�"�`�O},�+�)Z�OU���'��2&LA][L��Ƌ:Ju��:�'�l�p�	�^��;0�̖?�Ý'��R��lR���0��}(�b�1�y� A �t8��AIq���c"��,�y�$��ms�`�㋂o��HQ�`�3�y� �l>�jw Fj�vQ�&]��y��\�][�j¢�a(Ґ�m[�y"թ(p�ģT��-��DY��yb��f�p� ���*���ұ�y��ǇCH$0Q�ϊ3��H�E���y�#�?&k� е�3u�z��菀�y�Q�i�#r�'l �F��y"ԻK���p�b�4t�4QF Η�y��S0?攈ǎ�< ��1cdnF��y2Bc��UK��Y2#�ق��yb N*��y�3.a��#��S�P,�C�ɭ'B��S��C\@<<��oP�i�ZC�I�#h����ȝ����A�6�tC�	"xΥ�G�Jh8y��,�J.B�+]4ReP�b�9�ʀf�Q;"B�	1WvM�5�4��L�Td#J>���r؟�k6j�	C�̠���X�{Hl�$!,D�(H���#�8Q˕�>p�3`�)D��T��e���79��)�1�'D�<�0�����B�"E}��l
0� D�x�q,V�(pI�JĊ+u��95�>��MdJ����R�T�~�y`Gߑΰ��MpЌ���\�����0(ߎ����r�|���C�G+�	*�C_�v�1��dR�r��;%'�e1�X:\}�ȓv ��.�:1�$qQ�
L�\��K�'��I �c^��l���b2S��� (a��f�*k���&$ڱ%�(A"O�s��.$��#�=
:���"O�tX����(���ߗ9���<Oj�=E�dB�g��`	�AD��ٲ�͔�y2φ/]<�0��-1�\e˕����y"`�+B8pH#�0{�$h�@��y�./v%��k���36��#!@��yr�!6ߔ����Y#>���ה�y�o�e�>�z�b�� ��0���y2B]�4{�!��k	�:��a�Z��y��T�L�&<�������fė��y҉�4d����ª�lڤ��@6�y�b3OABd�RB�1j/f5A5���y��Q,ah$�bpa3,Ř		U��y�C�s� 1Y�./f*5�t�H�y¤ƊgGCBg�<+I���JM%�y�lR�S��B����8�!�X��y"N���z8��(L�,��I��y�.O��� �ޚ	Y�������yR`U f&�����*.bi j��y���r
<*TF�Ud����y2��y�L�W�Z�HV �L[�y�-�I�|�
��qDX� b
Ɂ�y�E۬7ꖑ� G��y���ש�y���3(��Y[�BR�4)�J�"�yblw3v�:􉒇>�0��$@��y�A�8s��DTNQ�2���� �>�y��W%=r ��ߛ+68�ŉ��yB���C���(����)�9�y��Cy ��� ��$
�@�T@�&�y��-Wn��C��VlF�� ^!�y�,�1X�@Hc�K
2=�P� ��y҅����u�	�"���*$�� �ybϞ�x�6}��l�>���f[��yRH�%��P���onu9aJ���yR�V~`�&�� /��}X�O]2�y�o��Q^��R�Eֲ:K�\�G��-�y�)	/�����*+�Td��T	�y��A���MSD��)���˰��y��T@��8�'#s�4�:E�]��y⢌�,��.�z��0I�E!�D�����b#�5�$�(��H�!��G#Ĉ��_!�*,��ҩ#�!���t�8]B���j��4+��]|�!���,!u�\r	̍P��b�b��!�Ė�I��i!h:z-N�����!�DW�iO� x��;"?��Y�Y�4!�d�WI6�S�d��J6�(
2���;'!�$�nB�y�1㔼`-D��sb�/!�D�_��)y��v����&˛�?@!��[%�r`��`�8}���	��Ղ9-!���1Z.�5a�!9��i5�ϵW!�Ij�E���3�Rx��CT�!��J$�0y&�G�`}�`���F2�!򤈝"����,L���u$
�d !��Gp#���u��:� �ţ�?�!��i!�Hif�{� �k�]�!��H5���'+��S�0�C��K�!��.�Pk1��.u%8y�_��!�$�?Ä����?����uωT�!�$^�3�V�qI*ц���Qq��,TA� �ʵCx8)PB�zJ���ȓ]r�L��˛A6�!��\ B*.���c�F�`�)�yR؆�ے4Hh��S�? .�5
�t�v���;� ���"On����Ն�ӱ��,��"OTh3c�Q���sV�(s��88a"OnD3����>���U��:D�YJ"O$la!cE�X����Bl�X�b"O�-���6!�d��.�m���"O:�DƗ`x��lJ,h�yq�"OB����[�p����E��=���"O҈��e^ޘ��Þ3���"O�s�KK�{����chP.m�J�`�"Oд��@Vh���sP�;&~��۳"O���g�8����&xc�H��"O^ʧ
�*WJa�Tb�#w-��څ"O�3C�ކu9P""�&exfh�`"On��A�G�q4T�x5a^���"O�<�q�î!�D�B� �Z�(�H�"OM���<�U��Ҁj��)�"O���W�7�E�"�i&����"O��j� �s�H��a�$20�W"Oj�@P
@�)��@W /hi"OX馤G$|D�����V��� "Ol���ò]׈�����
�@4"O{v�_�ML�1�'V�b<�"O�=� �%��P�C����"O>821(U01$��X�����ͺ�"Oh���G��:ULܯ]�>�y "OzɃe�F�?z��P��@/#\>���"O6���NA
;��Eqd�5ϖ�y���s�e�j��B�>��w�V�y��� �"�Ư�:#X8�+�yx~���^ܤ���H��yB�ݍ���Y0��Xd�ћ�N��y"��42z	yVFQ���1f�I��y�lX�&PD����,A��JҀ��y"e�8R�`qf]!K1��H�����y2(;r�ЁH&���I����l�.�y����J�~1��	=�~�����y")���@���H8 _�R���y"�V$s*��df^�r���[��A�y(�P2D�#� T"|@j��P�yfE=_�@���o�+8�B3L�y�A��D�,���ͼ��c���yBk[*t��u ����h21���yr��R����^�t���;�y��X��3�	����h�T0�yRɉ=���7M�t�$�{G���y��'��5��L�m���Hף	��y�����
ͤ\��qh�D;�y�l�;���!�_�<<Փum�y�
��.Q�҂~����3��:�y� �$*~e3�]5j����M��yr΅�,�����;h>�A[����Py�,N4h�:�P� �d,I(&�o�<YW&�v$4	��!YvP��&΍i�<1a憺N��) �N�E�$��Fd�m�<i�'��a� �1��*��N�<YA��F��	q��%��Q%"O���7�Z�hp���Ø0�@ya�"O�M2�a��k�2 z��@$,�@�"O�m+��AmAI�c��q術`"OtY��_��<q"��&u���W"OhQ	�K�XBt�6� p��1"O6X�$�}��5�f�ީ;XD��"O���6@J��HM���$>�ܠ"O� �D��f �-����Ũ\0V P|(2"O8Qs,���&�W�	�� "OB����ݾN(��Ɵ 5S�i��"O"���ŋ�Bv���C�͒4i�h��"O�4�'D�v���`��(0J|�"O,�X��F�,��yh��Zg5�"O�I:��J.�d):6l+o�i�"OvIY:a���
�@�Q��@1�"O���vA�	�4��
*M'�ݲv"O�4�����k8�,�@	T	D�u�V"OB0�kݞZ���:��]S�"�V"O�L�dB�,s�x"��`��Ѥ"O��A�̞�A6���R�ʵGʬ�ӡ"O(��deN�;B	�Q��1Z"�t1�"Or�8���|������P5i�� �"O�`q3�
��`��+d8u"O�|C1ǉ1FC�r��ՉU+�Th�"Ob�"�K� ���Q�,`�����"O�b��]�WĄ�@�R L���{�"O(��+ם[�X)X�Y��)�*O�m� ��|���2ю�,z b�'�H��½1NLȧ���F��'�,��.�!�r��v�)1�X�!�'���%��I0�Ц�ֶZT80
�'��6b�8�Z1v��a>�8	�'� W�0�
��5AF�Qn��'d��	 b#4҆ a��ǘGS����'��xcr�H<.w�L�L�(=� ��'�Lm*���[�BA�bd�$�(щ�'o\uY1i�mmRB'n!s	���y�IL��d@l��j`�2᫝��y�U��am���9�� 0�y2��!|lH���P%Cx!�1!���yb����P����4R��!�1Aϙ�y���rj�c��7��hj�!C��y���������*r�,S�l^��y���.���x��s�F��tbˉ�yRBY�AɃ�Kh�FM0�
���y�b�#���w)%vQ�	5#D/�yBfկ}��,�v��� ����y�h�L�R(a��X��Z��yB�DjT�"�*EF:0�+I��yRg7y���kQ�I4;���p��ybcȓ,d���,/g�3 �_��y��0�&��`7,:���%V
�y�J�C%TQ�3i�/(�(0��mÖ�y"H�<�Q	dˊ6'����9��O�"~
eOǸ�L���CM�8���]q�<y���^��y�ċ�	(��(y�^o�<ɣG�-N���[E	ˊaH��#�t�<aC䒡x^�M��CNRL`ԋ�H�<��?f�"�2�k�sr��%i�<1p�֨S�Dxۘ�(��EE	�y���!�"	idBhI	����y�
Ì)SP5��z�ʬ�d�ژ�y��[4�T��,�jx���)��yB��@�2��S-rs�i��M��y�,PW���4�X'YV`�{�։�y"A�#D���3cڗSO�]�g�G;�ya�e�,�"�i�>A��l&Ģ�yB#޵g������P�7�D #�!0�yn/(Ҩ��D70z�������?�
�',f�!T�Fhޥ%�E<okX�	�'��*��݆%��-JdO�k>��"��� .��Ő4Tr �����16Xc�"Ol�A$a)$�WF!ޥ��"O��R�E�RH�-"� -i��L"O�����B+/}\MÕ�$u�"O�al>gn8�1,��V�h�Ks"O�Py�&	0)�� 0��45j�q"O�ف+І6����Y��4"O���C��'?B00�jE&�8���"O�%�v���qi�g.n�h#"O�*��r�� k�^'�U�"O��!��́L�z���.4G��k�"OP}�smL4qɂp#���28��Z�"O��ӏ�7]� �]�8&��!"O4�p�A���)S�晭Y�����"Ob��N���Ɓ�!,�/9t�"O���rC�w��e��n_L�bB"O��j���V�v=c��Kf)�3"O�y�q�P%V��b��~��Dj�A ��ϟl��	2Fe0����ґE�tyԢQ�hJnB�	�Id�a8"�C�,�3bMZ/A�BB�	�'� &K%e��苲���@�6B�I2���!��=��x���<B@2B䉮0�"���b �=�T�!ˀ�"0B�I�%`�:cA�w� sf �Rb�C�	�O�A�HӞ=�D���h�*��C�	7?ި���ސe(s4㙚NRC�ɼK�����5��ɳ��@2:C�I�)p$3'�ÜX*�9���DQ�rB�	)����'��$�h��V�dB�I;*��r���`�"\*D�;{��B�ɝ0i�Dh�(C��SQ��"(�^B䉘h���PrƐ�����r�+rG`C䉵f��Bf�ͮ[.��d�J��XC�	�;dr033#_�~�d	�%�
~��C�ɦ<@z�R�S*�tiVjJ3��C�I� �@�B$�w�Y�S�M/v[�B������dL�g����熥��B�ɷ	~���Jǩov��Uh�(\AnB�	�K��������V�� ֲ;��C�I%V	h]ؐ�0#���q.�9�\C�+(e2�Jŋa�q��&��e C�2Dl�uE�
��E�"��:(�DB�! ��]�6A�<@�48��b-vB�I<2sBi���x�nh9��Y��B�	�^1�}��o^>&��3��+��B��7p�,�f�H2,��! Q��B�ɂL����2+Ƒ'{�=HW΍oi�B�ɒ<#�E��ļ-��8�.�;]��C�I�y�x�����3���b��)��B��	=���H�ɛ4Z�1�숟.�ZB�	%>K>��f��68ĥ�dAE;C\B�ɨC�XP��H�blv��@��C䉘B����C۲�T$"U[���� �d�]��YBʗS�N ��Ƹ-+bC�ɡ{�����ZH���6�Y-RC!��;����a���?��k%D!�$�n
�X%��&u��pe���!��8s�dL���N�C�U"�_�r!�$�$b[�Hc,c�	���y5!��L�P�f�acÉ<M��@�V� ��:OΥ�@�I� />����Mu�H8R'��F���(@�3�0�sAEn��A��"D��ʤ�ϲ�l�� ߟC�x�V�#D��:qh�<��أ!k]�E�)��3D�� &��C��_܂x�!n�,kS��Xd"O���$EU�F��U�@ tJi�"Ora�Q Y,��Z,ƂuG����'�ў"~��O<ZHDZu$�+Q� ��6����'�az2�H��Fl��G�JT�]s5���y����Ek��%�O�w殜�4hJ��y2��)^����c�{Q�I�åS��y����b9�#��,B\|Ȫ�"͸�y©ZD"�Е��1g�����y�Z�x�v�H*j6�P�F��y�JC�J��Q�Z5��Į�hOB����5�*y�m���A���#a!�{���2��6K��������!�d�>lR�*�h�0X��ƤC�!�$әo��A6[��ڰ�!�dF8#~���DR^���sh�0z�!�DJ2g��⁉V�d��psHFx�ў̆�	-������q���õ'�m�D�d;�S�O�����
�a���(�S�xj�m�"O���Z�r����ˁwX�t���Y�'y�$O�Bo:��DE�����ƣ��-��O셙A��`����+9�d"O2��H��	�
����?40b3"O�	[Mq)���)�� n����D�OJ���Q=A��`�7��E�T٩�۩�!�X�iu�0�!�a �C]�!�@�/g�p`��x\"��wC�,t��7O��@C�:~��8� �I'k3�MS�"O�8�2��r<����,S��۰"Ob-�h�4�i�CKL�"�8���"O���`d����
"�Yc��IJ>#q�)^g$���+��A`��`f	$D�0 ���+�|�T,\�" !F D����G�DJ���r��(\�T���=�O,�d	%,�����֔@��r%X����$#�����[GnUIB�	��p=;w$=D��z�3,�L90 ǻ_j|](w�9D��I�H[�-��!�ɝ�j��t�#D�<14��3w�6}�ר,	�ӂ0ړ�0<��噀V��E�r	�+C^� ��KQ�<A�O�ư���5�TPs(Jy��)�'/Vq� �$�Ḇ�E-��ɇ���ط�~�����i�Lm��&A��j� �,Uw�%@p�H��z�ȓp� 4)�B�#��#�F�_�4Ԇ��^,����Ȣ���Q+ Q(�	ڟ��'���>Q�+:<0�TϘ� J�_�<D���t/\ɩ��2A��w(^y2�)�'7� �q��:�@]Y4�=�Դ��o��I�4&T�p|�\�1I
:���ȓ*�|d��Ձf�>���)�h_Dԅ���q�2��6fV��P���/R@�ȓQ�$;G�_4�:PC%b�:p��'ў�|��
�<m� �!W�u2t1��,�n���0=�D���<n�h�V�ޔ~�:E�1@�l�<�ga�@C,�(s�F�Tٞ���Ng�<�a+ϱ?k"��(݄N�ʅ�c��c�<�7�/K���%oԿ]�ĐS&,H_�<�0���8%�B�&�(�a�FYyr�)ʧ>h�آ-�WҼ����!���$���I�Sܧzk�I�T�-~bLQ�G������4�5a��+.K@i��]�5p�T��^7�1�`j�.u<%� � .��$�ȓs\���.n��ӇU�V��!��S�? �����z�H����7/�xK"O�]q�M�x���5�h��g"O`���6#v%Ӄ���:�0�["Op]BԨҎYk�б6�FB&69�3"O$��bfT�t�x���<�D�IZ�87�&F�oX�vZ���#�R�<��� ==ڸ���`�<t�j�i�<1� \�R�`q���2r����F�^�<��Ƙ�1�z���M�g�ti���YD�<1�lާ5S*�"��#tIҵ;�P~�<Y��7HP䨥��enb�S�B�<��	@E X�q`�M�a���q��d�<A-�
�nEQ�(�V�<����Yl�<i�����0�����w�Q�<�$��,��Bڹc7�	`��N�<���_%B��c֦��	HAb��H�<a�$α8��V
�| \)I�aV�]�ID��t�����Œ���$(;�A��?D��Ղƛ.�l��ʖ/��E��<D�X�V�g�AX��z��A�Q�-D����66-X�K�Bӯf��e��6D� C����y��"5.�!/�!򤉚b�f�J��0m�&Zo0n_�O\�=��:)p�,�/*t���ΒiO��+��'�!�Dh� �d��&u�<�Q�CR�Q!򤂄 �Y�u%�2�r�U�zU!�$��L����)ިXkT���l�7!�$�2(�H(��M!]d���ю�Y2!�˨Qz���Z)K��1�-B��Py"��5[��m!�.�	M ��X��©�y�O9-V� �!M=l��Bϔ �y��Κ\�R1��iK��f\H,�;��'Uaz��	�Z�تtJQ�^-����y�f�F��@�y�pḱ	C��y"K�]�рMѱx�`��e-���y�BM�e��(=T�I6퀗�yb Q��:�a���V��a)v!��y�c�(a�@!�eN;B���O���y��Kg�h��Q�+�zEå�E�y�K�jxE:v�&#� ��3�ԍ�y�C�*O�����֋F����y���H�#��ΏU��qoQ��y�b_D�T����8..$�w�K��y�W�'�vYp���}�(�Rwh���y�b��S�d�u�&t��@��	Z��y��:jؖ��$�Ѻ	xݺ�)���y"�^(a~}�#Ě7a^P�JFC��yB��j�9��C�RInM�RE��yR�Wd�p��k�B��Ep��Ϙ�y�Ѵf�.����A!|1f�\��yrU4�}R���"N��L�@��y� �s�R�ˍ�fY���yb'J9���k� �4XE�[��y"��j�2- �)�>~قс7. ��y��B�t�ԃ@���w�>��՚�y���J�z�����h�F]c����y�$D!��=�#�1HZr�y��b?D��b��ŤX7Rىqi�1/�`�*6 #D�\KI^�,�8]E(0N�BV!>D�D��N���b�Q��LC��dB(D���@�<d
:����3b���j�c�<a���Qh��U�P;^Ul8�Tl�
B�	�U�A����$y>��ȩ)(�C��(�"4�d,]�y����T�4H�C�)� 6媣�ȅ��]�2oZx"�7"O��H�i��Z���M�\���"O�� A�$���J��ؔN�<љQ"O�D(1L�$R4�Ҁ]�"���"O�S��ƕ[&M�L�/�@��"O����ʲH��4K��/�D��"O���A+�?@`�c��A�S��r"Oh���Jʪ)��Ι:+9t$�v"O�Pp��5(q!�MޯyE�$�u�'�Ғ�����2U�����mNqc|$h��-D�$�k���q"���h�P�c-D�`�@�L*Y/& Iec�=8\����+D���a@
�g,�[�Ox���)D�p� $��Z|�[�C��]�Y�L2D�81�]�*�����iq4�.D����b�1+Hl�Ɗ�E༥�j+�Or�q����fj� @�BԢ��7>��%��R,H$P���8zb�J"*��g괄�:̬�5�ч�I:��Y�}�ȓa)@�{d�V)Y���*�{}����Tq���>)���g�!w��l��Qj�Թ7���-��I��*�
!Bh�ȓB�Mp��6N���N]�f���#�>|Rc�	W�Τ:e,�{o¥�ȓ]/Dy$aݩG(Fˤ�R�R�JćȓK��Q0D6g������|����+q<��"�̡v�&|��JQy�d��1�B�c����$UV/��`�2���Z�X�a�ϓwjHb�#ӊy9(M��D��Pp�/~���1y�&��'-D����H�rb��E�'7� ��b)ړ�0|
E�̋M��� ��΀+�2��`bGo�'�axR��@?�0j��7w֜� G�Ö�y"���+Ң`�A��)u|�������y҇�/��AO��y�D�)�y��1/��g�NG�,�u&K��y�ʊ�vQ�NÙ9�U��$��yҬ�!���"�I>@��X��@��yҊ<2�^QsMO�6��������0>a$/D�7䕢����N��$l�T�<�F�	Hd!`#ʜ�Y�|E2��Q�<i�Ȏ�$ $e�u�@�kA�=��C�N�<Y�(^�y@��i��r<��y���Py��' �1qwO3l�a�('8� � �'�8���#H�ŚH�Bh�Uk��D%�N��R/Cn��]�#�/J��L��"O�r�/�3L��aT��z�T�3�"Orػ5H�!0��x0B�U�x �5"O\ի���f�@����E��)q�"O Q�Aa����q"_��c"O�I
�I˄5,��uK�I�K��'O��!3��#Q�f�OV��@Y�+;��Y���� �!j��F�5�3 �v}�C�	�(���C�*B9E�e���=X��C�	<@j!�mWN]N��_>A �C�	�=<� ���2���^�L�rC�ɜF?:ȹ��U�P>q��.�0w�B�I����aVGu��m�4��7a����$0�ɏo�����W0D��Ё�g�
J��B�ɓA�9���RP��#M�
�pB�	|�`YK!D�_�N|�>7pB�I�>C���W6C_:L�e�ШH#�B��-	�tC ,��V�5��/TPC�I4��@���=RS+FM~˓�?q��?YO>I�y
� <�Ia�V�2i��x��E�'��(3-�b*�!��$��1�5�d�Oz��>Q �'�&��d�7�?U{"���OrB�ɢ=�5j���F���4�M<C��69���S�LQp���AaK�?8C�I'�(�P��BK����N	�36��d-?3%�|�ѡ������oJt���?���On������ �I�6���q��3�S�i�	oPl��!皢y����eo�m�O��=��P�!��2��	�Ճ��p�z*r��F�Or�`yv��>�8��!c�7Q��dx	�'�
=���s��)a,X�Yv�1X�'N�dI@ 'U:��� #B:Z`�9��OH�:�
����cfR�k�
!�t�'��[�)�'U~�u�C�=`^Ժ�>�V̑�' )qdN���VȠym����'8 Dyw�zd>�9���p���'�.(����!u���	b�I�'H��x���$pTܐ���2f����'��"�#�5;dx ��	�W ��n���$J����e
 &l����!�5�_�R{as��ܾ'�v��ȓ(�p��߀n38�
�X?�l���/�J���`��	*�;I���$����ɐ|��p��ˇ=��'���H��C�	+�xih����G�U�C�ɀ6�����q�T��JB 5�dC�I�h����c�%ZնxJ2�@���hOQ>�8 �\�[��x�d�J�wI�5�,�OP�	(�<��C(,e�7�Q*��B�p�lm	�'Sɶ`)��B�/p���0?i�N�<$p@����U����?-M.-��4���Ŋ�NR9B�4b�xń�	��m��-�/4~���Aq�.��F|
A����$?�t\)���U��m���+!I<�r�RįW%#�(G{B�'��>��#�W 0��@���V�b��k�<Q���N�𑹳a�㐸���i�<�2䊸N~�bU��TxV�13�\�<�v�U��Lx(�h��^h�p��V�<���Eô ��#[T� 7�V�<��(N=| `\��*qQLu�ALR����<IW\"���B�_\�@f��'Nў�OrDl��
P���G`�5sMs	�'N��M	�s0�xF&:�$ta��D,�'rPșv�	1 �.x�c�t���:�d�!A�&$q��ҴDS�p[f���^���8�kȤZ�|`؃�S�
@�E��A�d��T�����+Q	m�zԄ�	F�'��,Ti˛xf�(y��� ��'��B6�M�{�4�A����~�f X	�'���*̌�բ��d�|Z||��D�O�"|т�rCJi Pg� @
h��Ӭ�B�<�
�=�p���/ʮ�5�_c�<P*�5���Qg�����i*���Y�<���� yL}� � d����/�l�<aV��� ����W%�zn|x@F]h�<��!�"q�B�Z���Q*t�a�<��Q3%I�=���1��1"��D�'a���ܭq^���Hˡ��P��A��yfR�HQlD�M6d�!�D��y�����n�Y���.54D��L��y���9��l�v��5.�2��e���y�_$+���rc��[쐰C�Ȕ��y
� r!� dKm���Іi� ��ٰ�"O�����4"��E;�ιOR4 I`"OPu�� y	�I���)g�D�"O�H8S ۇ%� �C�%Ҙ<W`��"O4ij!��kJ���K�!i���T"OTe�!��:+$�Mz���n��r��k>1�2�F�{'܈��nW�/(v��7D��CG.�}�Li��O�PJ�Y��(D�$�+�+�@�r��L: �j�+ړ�0<q��Wowd[�
��<�y��L�O�<1,߿�P��@��.bN h�m�e�<����	e�U���A�f����Y^�<�K\�fð�% ���&��G_T�''?}�%�xw4y��P+8�� Z�	*D���� A*N�������nu��'D�)2g�-#����$n��tJ�J2�7�SܧM�����2a����2��a�\}��_t����ӛ(tސJ�cXQ̰���ޤru��<LQ�	��[u��Co�����X�<��Rl��s32�&�$G{�����M��aV(E��i��1��x2�3S�KØz�
K4HP�2�J��'�>�!���u9A1A�T�%+�1�)O(�=E�t�	?(�Jq��N�j��`�ݖ�y��j��s�Ƒ��ڳ���y�`�:Jk�tt������y�ȏDJ������?�^��cÕ���'ў�O��T� 
�R��GY�0/D8�����M:�����B�mM�4��\yG!��6��1�)���6DZ� &'5!��/bq��bȃ0w��ը$n�0_D!�d��@�j�����x�Q���y/!��Z?J��KC�h�:p�6E�$!��Ok��eʖj�$QJ�a��af!�D
qjJ(р��LS@0��Һc��'Ja|��O�U�9�'�F��n�n
+�!�D�O�X�pT	�%��ǭY�!򄝖���2Dk�\$(Cc\&}�!��	'���RC)Ս⹨�Gʴ�Py��ۅ~h�A���9RĀ�4/���yB`H:~8,��#=����d�Ȗ�yr�����C×aͺTa��_*�y�C�-$ܠ��o��%�&`��ybj��&�[FȔ;d.�X�H�+�y�$���T�?]xL��UmG��yRğ0Rf�%��E�br ��.@-�y�/��D���(b��*�����y'�;i�N%�C�@7��-d���hO����F7SBdt��gI�z�e�a Ց,!�:|�xcF�^�0Az��J�;m!�ƽ>�����#[REB�O�Df!�Y�'U|������AI���)A�$+!�A�s��@#�BO"|V� ]I!�䇔	H�Ӄ�\MbYk�f�$!�
 D* R��G">$��p���S�2�)�`~�17-*�UHa��"�����'!��j7��42����^F6�
�'mȥZ��
a��:�l�	����'�`�W��n�����*��~�C�'5�г�Eֻv�!zS��r����'c
0�$C�'���'��>�0|�
�'���`�7D����v"��5�d�	�'8�L�梟� ��"��'��e��',�0��"��~���0��#i%�y���� �ѱ�o�)aZ���G%q�v��q"O>3�"œb��-�΀��B��"O�� �Ƚv�$�r�]9L�v�Z "O�y�f�B�4��6�ֻl�>��"O���ƅ�u4�D�ƋwI80����?����CO�9�C�5�b�B5*ȿX�|��ȓ}��ԫ�� �4�x��AO�Z���ȓ3p~Lz�j�->�4�+W�S5J����8��]��c1N���!#�٭!nV)�ȓa�a��%8���2���fp�d��'� ��3b�t��q�U #jh��.�n�S�cH�m���KQ� $��&2�}��ՃDN� ���@ ����|"�1�%{ܽ�'텔h�2,�ȓY'���U�4���Al�R�\)�ȓ �lX�th�)i�È.�­��n��4RK�5�FH3t>�:�ȓ>� �d�
�����QF�lh�ȓa�Α��+B���FC�����'��=+��Z�s�l�H�	Z�}dŢ
�'݂MH6��3-���G�%r�,�h	�'��|����Nnx�r0����	�'�L�wnW3r6�B���T��'A�LCv�;�.݃�c�	O,��'�qp�l �~�ā�& �Q��5�
�'�4�s��N/)L��D�#A��a)
�'p ��*3j͸�%"3t�p	�'�Z�9���4rA�H��mG92)��'Y8 6�I#/_j��s�)��Hcj��x��i�����g*q`\h�˟�yR+%�h�'!�U��ia�M���yBI�T� m*�B����;S�ۡ�y���Tb0)�qOז�¹벌L��y2�W'$�l�j�Oؑ�PU��b��y����OM���G�=	(Z�ࣀ��y"O�S���i�!��^����U���!�O�x@S��I�p��3@�x�0e�"O���p���U�	9�-]�8�Je"Ofx	Pl�rZ��a, ����"O�|Ѣ��'��驅@�̊��"Od��e�J�T����Qo�>q����"O��x@�U�*�����.�&b���"O9���Шc^P�9D8����"O&m0D�G�"��
 ���IQp"Oܰ83nVNЅ�Y.[�n��2"O"삠l����L� Jг�"Orda�+[�'�{���"�x�"O)Q����'���#7��""O�����9R%�0R�~|��"O�(�9{<z��&C"�$�"OԘ{WF_�gy(�P���i��!R"O��R�@�#�Ҁ��d=�d�x4"O�ݑ�l+-����P�m=�ʠ"O:a`  D�0|r� ӏh*@�Г"Or4
�BI� O��['��=wdi�"O�9�����U,�y* �Y�Vt��k#"O����N�� B���sJ��"O�1A��J�o~�ƄR
6�̌��"O��{1+� lQj��s�D�\��ܻ�"O��0 �!B�x�XE�  ���°"O��0�lK�z6��8�G�<xR�: "O���-H�|k��dg�n��i�"Ox	0���?M� �����m��13%"O�9r�G�X�B-z匂�'���"O� !�C�3t��1�O�H�]:�"O0ɛb�U2�j��W�,I<8��"O���ލe�~�:ulv%�d�"OFݘd+�4(i��$�	�Z ��C�"O��p H��n�+��v�	�ǋ9�y���<�<���nޜtW�9�/;�y"FWtYn(�A�:6ذ�Q%Y7�y��T�H����n��4ȮA�э��yçL[r����
y�nU	Do�<�y�iI�aD�i��
�o�49� �J��y�E(kPy�!�7�2%s�c�3�y���6@DuU��j��c���y��L9}�}�ԆG�W<ܫ����yBg��H\���9JF�����yb�Sw�h�Fb�<��`�g��y� G�?9�֎H�5sh���P�y�[?" ��XY�zT���<�y"�
�9Ă����U?O�M��!��y�c)�U�] ��� ���C{^d��+P�bB���u��	�6)��g}��ȓ���"�/a��adm�V30%��3�>�����>1�<���1�q�ȓVd�����[=�,��wo�0�ȓ��]��0J^diks�u����ȓb��4�����%�D�I��ߢɮl�ȓgH����J ��#�j�a� ���3t2�,D!"V$8k ��}t"���<��,SD����0� D4�ȓ=�l�O��2�&��ƒ7i���ȓ8:���q�F @y!�w-�+d���	4��pA���p��H	&B&|���ȓBry�k�y\��(E��
p���u��ٙwg��'"d0���+��h�ȓC#VYj��
�~Q��rCM��K� @�ȓ!=��˴��G��Ы��?1�ņ�ʆ���J���.�%��4��4�ȓ����,�c���!������ ���fJ��4�U(.��\��M}b���+Kp����$%d1���iqe�ǆrT�Y��[�ӆ���*>��޴]�q�	�e�( ��z�B<���	sv�	�0a�g=!��j�>��C�(7rą#ю�:3Q�ȓY�Ȅɰ���uh��Cu�*TSz���M����&�3��#!))����r3��v��u�` �BU&/D�y��A��y:�GH82~,�
�) �e��44��ѧg"Q��իK�!�ȓ\c�A��MZ�>��1ra��Q��l�ȓB���ac$]�	���IFN��=V$�ȓ+Z����H��t���\����8�d�2��Y��ma�Br�0s"O�T�3*S�5�ã^QLĤH"O�9w̕�\ȅSB	� m( *O(ݢ�d�(A����Մ17�,+�'c���$�E7�R`[�!�'�&A��'�8q�oɆh���ТZ%U����'H��Q��"Ӳ�#H�($ �9 �'�آ�аN��x"O^��n��
�'P��)Z�BiI��C����b	�'BTT҃��<`&!B�EC`$p�'K�1��Y��b�P�-w��|��'B�}(�,	�9�Yh!��?���'h����T�N�vPrņ�5y
��� �u�0D� M�� BQ�[�8[l��""Oh���ȓ�,( ���3|Hb�"O���3� �	�3�' "pek�"O����Oէ/ x�G'A2&�("O�m�E�X���D&H����T"O!�E��Q�xu[��)�I�5"O�p� A�8B��`&ܜC�){�"O�`" ��
堡e��S��"�"O�3�ڎb'�i�$�[���(@"O�U97oĜ,�U��˓&B5c"Ob�05�;�ΰ�񃓽d�&]�5"O
�9�E�Ma�%#!$U��p�d"O�4+!(��f�{�#K��2V"O�=R�oD���飔I�P�d=�!"O�%@��'4RɊ2"��	���s"O]ҡf��~���$D���T�!c"O�����E���7M
?�}�"Ovu�T���s3L0~���x�"OP��VRv� �jA�k��Qy0"Ol�D�K1WJ*�H��+4�6-��"O��Kת"S�"FJ��v�ΠA�"O^)��B���~mp�� ɘm�a"O�l����s�m�V��,-Y"O��{�O�/H�s�P�~ق`�"O�3CJ�Yx��5 [:7�Ω��"Ob��0�
�}�vx��(ѕ��ݢ�"O�ղ�e� &�h��!���?�8��q"O���t,�6VKV�S�왊��}Q%"O���D �h{�j���j��P8�"Otty��BE�Dk�J&��b�"O�����b@�����?�H0�"OX�vO�.2*u���״pIz��"O�d C�_ bpV��L&eQ� ��"OD�k��5����.R*�"O��+��T�s�f���)êDG���"OXȳCᒤ#��Ӷ������*�"O0-����0pp��*W��"b⸁�"O4xI�ǘB�U�,F��zs"Oހx�ܪ�(�'�C�o.���"O�H�2�#1�$1���*iR�G�<	'
N-i��@��	'
 �q�n�<� O��#��@�*VrgD`ic��g�<I# X�d��@����K3@����Y�<pCL$:�M���N0�9+��W�<Q@�Ƙ>Y*@�+Ȃd,d C�DQ�<a�W�<�0���$��C��zDA�I�<�t��2=���녷wR���lOD�<���'�2�b@�F-p5��bsf�}�<��N�|�2񋲋�?���"��Fv�<I�+��@5`�:u W	}B���J�<��A�"UИ�0�8pVM
��D�<9�ѫB0��b,�28j �+��~�<��
��h���.hL�SQ�`�<���
�/C���sJԨ(�j��B�<)0kN�HO (A��%����AS�<��ٺc��ᢑ+�#S���(��HO�<�B��]�E��$&c��a�hf�<q#��}�,f�7�~M@f��W�<�LQ�D6=*�m
�@\X�vny�<�:h2�T������9��<i�!��I�i�8����ߐt�p�3ԣ�x�!��L9h��3\�\�r�Y��n�!�S�d��u/۝j�r���Q�i�!�$a�a��,tX0`�~�!�� ��Q J<��2��	�l�B"O��v���mG~m���0M��!Ya"O҄���	�,�)�F�=�~���"O���*�"b��<8�۝h8��"OEAͲ���+Q��4Y�Ey""O�@�Q�GXh��c�.1x�1�"OԠӤk�x�-ђo�	@b 9"Ox�B�^�L�:D#��T�/ű"O.�����(Ya��M��q��"O�yJ�+Θ~ >�rӎR�{�hg"O�ࣷ��+0����˓�s�a�'{��C$�ǺP����M8zߐ��'��TX��ًDQ֔�s
��&V����'a�ebѦ]�d�ִys��"��i�'\�iy�O3�B�	ѓj�H��'���hE��*E���3Č�a�"��
�'����S�ɣ1%2�:'�Wzΐ�
�'�(�fi 3h$C��I����'�Bu�Эژ� ��d�LSBn%��',h���O+
�$�z��,u�q�	�'���Qg �'%����F+m��L��'�J��)��F��a���s�`A�'�p<p��H̒��#Z$��]��'���SQ�Y�DV��r�m5��'�  )��եC�.y`����&�ݺ�'80�# �@��dG���=��'��YPb  ��|у��	�yC�'~������(F*�'��-�X�r�'�L�ӔɄ���1#�Ś(�X-k
�'z� �dŹ}|���1��4��'�zmA��3[���(��$��I�
�'��]��ŝ*]b��d-���I�	�'Pi�+�w5��pdc
5�t��'�L�����j��qz�69��!��'b�!�Qȟ�1u�C�+×)L�� �'φ,���"��y�(y!(h��'�D��fdj��U�s4�̣�'��x�MM$���pUȔ�:��!
�'��䂢iN�q�hq�Sl��㮤��'��c�i�7���#A����'!�[�U�8p����(�:dh��
�'��8��H6}n���� B�0/$�(
�'��=�f��L@@���=-�V�q
�'Xb�p`AG0r�(j��U/"�z�B�'a@�B��P�$�����/*�b
�'g�,�*Z�g����LH�#�j1��' �0��^>y7N��	����@�'`���/���9CW�Fq*	A�'if ҠO�=e��9��g�=<�&�;�'ޔl�@��?�pH�5��
9C��`�'a IA��L��@D+u�<���
�'�0���Q&u:w倲9��s
�'~f1"�Tk�ea�gȲAݬ�0�'��@�1�S(^�A!R&�3��Y3
�'� -B��!vQ&̐B�%"�X
�'�x�'�7<୻����Ot��
�'7`��$ ͗R�.����ŽF����	�'c��aM�66@����G�/8�!:	�'���H�&6=��:�Jȅ7���H�'�9�Q��4aN&�Q��_8*�����'�ĕ���#g>��$h["`�4�'�V���X�L�5���&ȥ8�'�p�B�DJ�ȹ�\<�݃`��{�<�F�W�w�A"�o�*� h���n�<� ��A�\�/#����ƀ#t�V(x6"O������-P�-Y0U�gT긠�"O�i�&�ϕ]�Dm"��M1^?Pٰ"OR�y�	�@f�� S+g*���"O �1ʊ,~ƾ�Xtأ3��!�"Oji҃�+2j���qbϐ1�H��"O��BbZ�����߮���"Of�2��E	�F@dǂa%"O��2eK�}ޱ���Q��V��"O6�:"l�&0���qG��n�dAB"ON�#�Ⱥl�~}s��#Ti|бr"O츑�@_�F IX�K=d�����"O�)c�!h<|]�w)\�L��a�f"O�}��L�<�<��GۍQ�
0a�"OhɲC��}h��H�ѯ%��S "O@r6靻zZ�I���I�x��"O����a�&��Z�)�����"O���BY�{
�4��.D#j��A��"OtA1��9:����G��Ez���7"Od�ir��"@Ȃ��Xit%d"O�1��ڿ.��<i��	%]@��"OT���Hm�2�RQ��
yR	J�"OtԻ�$���hq��.�6ɴ�6"O��q�fL�H�8Ej�o_�Ld!R%"OB��ѰR���Bn�T�At"O��D�(O+4b�MD^��	�"O���A�lW~y�3�
D��9��"O LC�`Ҡkt}kpl��\�z���"O�q0��ßH���*F̏��<c�"O
uk#�p�΍ZAl��o�DX3�"O����l��X2-BCk�o|p"O�"��H�3�xؖ�ߣOr�('"O:��a�] f���*�N���	�"O �#�0u���N�#�`��"O<��Š�
*r0R��M>L�\2"OVt��씅A�l=ZS`ʦ�޽Sw"O��ä�NNq�TQ��I�����"O`HO��U�S�6� ��"OD P��2��풤M�"��=X4��\��I9:�X}ƮۀnmD<�@�P�{�nC�!< �X�4K^�����Ȑ�1�6C�R�� ��$bk�E��2P���D7�0�&�$V���N�(tΨ��2D���Xa����ѮG�CnD���H-D�ds�J�A2X�K0e����/.D��c Ǆpgxu���d�
ٚGH�O�B�I�{��(!a[q頩2B	'i��C�1:1��&K�)Ȧ���m�/J6tC�6J�I�kA7>@|�Bu��(K 0���>�-[&N��р�,�F��CvfDF�<qVł6���*��L	Z�xg(�f�<I�o��m�A�3*�l��Rl�d��hO1���x��@ B܃��=� 8�i+#=E��4I����5t��ز! 	f��'����)�|BD��d?Ry�6)F���d*�<Q�)�O�����
JP�x"c�=�:a�N�M�ax��I4)�T��BN*G\�n�$5�NB�	��m���{ax8S�U�[p>"?�4L�Q>��jЋ:��A�ą�:M��Qg� T�`s ����@�qCa˦37��""Od˄#�%�� B*�@D�Q��"O$aM��eԚ�q4*O�=6t�s��D&lOJ�35,�*�.�Bj�G�|i���������S�
�;!FP�/�X��2-Y&oL���D~�� v��e��'��\)Kݴq&60He"O���c��0PJ���w���-��5���	g�OY�ܠreL�6Y�:�տo�24��'��|І��"g>ZL�#i�!l�T�	�'-<h$N¸��U
��\�Mo`�	�'A؜3��L�4U#!��OF� �Ǔ�HOvQ�kb���2�`[,��DR��'��	�2��|Ze��UfD�j!��6��C�	�Wr�y��h51ҸQ�.�B��#>A���$d����Ƃ2.~�$��.�I��C�I �h��#eQb��$���k_��IJ��h�9�.�?�ɓw�F@DƁ�""Otp��c�CِE�d�;4;��1#�>�	�0�h����aKD,LSm��ȓu,0����K�qy�D˔*��q΄��ȓ.�� {&Eϸ��e�DF]{k� �ȓi��Dۂ银Ft�[�lυ-�v���'3���"+S3��� ����+��<X�' ��r���;fKXU�&'H&&�Vai�'9&A�vL�:Z�.x6�S4 H!��'�ў"~��2�2]����?�$Hٗ`�j�<�1`ϋziD�0#蛰j��!a�+�]�<y�f�(����/��A��	V�'�Q?	�t�K�58���Q!6��#Wn&D��Ҡ�C�E���;��>�H���i�O7�<�S�O��U��Ty�Ić��*�R#c"O������N ����	�]6��7\�����8t�}�sd�
�	��'Ľ: ��$d�d�3Y@�*���䎊^��d�>D��H�kڽ{�`Ԁ�],��qa.<�D��d/>�N3"˼V�� E�A8�!�<OM����D׺d�jq����9��xR�K�'�"d9���9��Ic&㇫y����'	Z�a7�֝2%���Es��z�'L�'��)�!�-ؠ���1����<�����W�DS�dq��� �L�x���?���CA����K-	��\�BD��a��KF�7����$Uv�ڡ*�7�K�.M�>ݺǪ>�S��y⮝�4�����.cY�tB$�
��y“.���H֢]{�8 T���x��'/�S��)5�{��A���*�'�(@���^lDb�d��~of�a�'��qz����K��i�T ͖E��e!��)��<9��H��H�OW�3���١�	a�'�ўʧP̱sS���&�ؙ ����4͓��'�ay�Ē�^e� (���61��U!ӎ��yR��-fi~�Z� O%ㄘ��K�y�F:;��l(�KT�8�Hr��F����hO���d�E�Po��P" h�m��r"O,����N��e*", ϞI"O~�c���6U�&��ɅR���[��Io�OH@�{�ėEW��p�ɑ�D�<�Q��d:Or9Bo��rT��A-�^��`k�"O�Hr �2��8cpΘz��8 �"O��H�.�A�������y2`�UP�p�vOǋF7�`�����y�`F;�v�`��"�RH��yR��24��9DM��Bw�$c��T��yrg�#BZ�(��ӭ�@�@A�8�yBd�<G�p$&��
�J�;Ӯ���y'Z%V��2���|���,¡�yB�	����VM4&�����^��hO����W��P9�c@�2rES!DG�	�!�āi�h���	�*jZ���N�{�!�� >� c!Z-A[,��#f�8۔ȺR"O� P2f�&��A�E�"����q"O��K����3C��PZ7%�\5SОx��)�Qj��S �F�*ĺ��%RN�C�	�|�c�IH�a�$@�����x�B�I
N���i����'��%	�`�.lY�B�	\��m�7e�p��J�k_�l1`B�++�+��B{���� +_6B�I�w
�2�G ά�"��8.���s"O��m�t�@����R�O��Ec�'	���k����7X(]��FQ8�H�C	5}24O���D˝�Z���Q		�d�ZrK��N��	"FS�I1�H��7�`��)peC7�P�b�O^�\S"On���B�}�%�1�G�5��m���'D�ꓑM� ����'�t4�gI:|pN�)�!]�>}��T��f�6�FԣcH�0v�Dp�@G��'!��Iz�`C�Nӝw�:��"hj��rq�6O0�Iu?��'&Lu#��ݠ-��@�U��iM2�Xw�P*r�!�L3x��S��e-J�9�BƸ6��|���?�J��S/U�c>�$Y�3�����:+��A�c�Om!�D���N��n�,3Jy�@�ء	X���,E{��D���
��Α����{ŧ���y�:$�x`�r���4�D�	�򄬟����-G:��#Q�]�,czy�Ơ͸w�>��d�����q��i�mȶ#b����1D�䲤"ԅ&_A��i\�
��%`��/D� h�O��3)�0id@���U�V%-D�A%��/	j� ��	�7�E��.D�XN�.��Y��H*lٺ�A D�@cӣ"CQJ�{�`\<#����Q�<��s� fBR���9�s(��?OR���Ig~b �%FM�)p��٢_�.�!i�4�y�HS�u��P�%)�>Q����fn�1�yBJ��D)2@��I�f50Ƭ�y��B=z)["LӲCr@�B�T��y��
�j��@#3U�p�@� ��y���)�qul�;{��3��X�y�㖢��-`RbɌ�H[6�K��y�,و Z�y�U�ժ.N�Ҵd��yR��?QnxI$D�)�p(�M�=�yb�R����#�hO���ge�,�y�-�?���brEˋ0,�G�Y�ȓn��h�
5	��qPgߍ[J���ȓd�X�[ Q1]~�PCB�<y���
b��T �'X)s�
�!e��e�<YT� �VL��Ȩ,I�E��v�<�bM�%w� ��!��.��YF@�p�<��(>,x ��Ҝ1k�k�<YѰԑa�At�B[$VX�LC�I#e��Qk���8f�*��3@�/�B�Iu�!0�
�s�l�Ā
=�B�ɤ	��xsSdM7C����7K�B�	8hľY�U�ߨ������΁W�B�	��d���{J�`X�lX;��C�	"AF�����$⨤��M̹<�B��TYd	�)ޮ<��L�F�I���C�!C�8���h �)\���� B�IcԽI�ă��N�S����k2
B�	(:�)1UeأZ�jM��=2��C�	�~8q�E�"@	0��eB�L̶C䉗t���J@�F0 �����b�C䉐M�,��E�d'��I��͔v�C�ɏ�J�����8��,��lׯ��C�I�K
f��7M~�f�0�I6W]PC�)� �� �V�,���JS-A_�M� "O<����l�0A!����(�H���"Or\`�E�.��j��	�"�*F�#�Ԣ�␛T�^�	�A��Q�6�ɑ;���'$_	b��`���+2YC�Iq&��$1z1�% QK2�B�ɦ6F��@v��q��\��K/�dB��%�h|��̛{��!��]��C�I�4��M���ȣi8�),Цs �C��BbL�@�M"Ǯ�p���<l�C䉢%���q,HG��9�bT%K�PC�I/0��Pz��Z��N�i�N'8�C�	�}�$Q&�t��f�ѕv��B�>Uq��i��i�^���j�;.~�C�	�l�t�gk]2l�\D S�]�4a�B�ɴn�L�HgA��<`��D =:rB�IR'�m�lB�	�(�.Ao�|B��+*ɨ]�� Z��������5�C�	.)�у�.%��y�gi� Iq�B�	�j�R4��f��t�d!7��i)�B�Oe"�i��	?b���Q�צ,��C�	>�Z� ��B?#����3s��C��C�A�Ƒ��̂#MFj�@C��;z��	����OK�ݡ��ĸ��C�.c�y�HU�Ybb�[�kC�Z�C�()XX(@B�%�z�s��́l��C��5��a��}�"]c��ͻX��B����9`#H|�y�J�;FB��0g�z���#J-B�lk�cȵ8B�ɏ/�p�&k:̠�IՈF�#(B�ɐn���k�M�x��'9�B�	!^�c�/_�a2������ �B�g��11�KJ8|��L۱�ܧd^�B�ɛP"����I6=g���E(�x��B�	�Y�x���F��h�Q��k�C�	�f]���%!�� SbG7B�9Nx�i1E�B�s	΄�	Q(2�C��6: 4e0΄�S �$�!�N���C��F���J /Y�^=r��+B�" �洲���p�(�+���O( B�I�8(��f��12�H�dϑc��B�I'`�*4+uj�|��H�7L؟H�B� 	�FeH���AR�8ХH!@~B�ɋZ).��ō31Y�}�B��`�>B䉪cBQ&��!�`I[!n�u�C䉩r�����%A#Fy�7G�m0B�	8y�v,��L�8����;
�C��.	<(��@b�	�R����L9��C�I�̡B�F� qV�Q *�3Jc�B�I2LOZ<(D+]�Y�A�4n��L>�B�ɘ	�\՛7⁶p�M��ʺZ��C�	&~O��"#�-g)�	����IR�C��W.�*�ʰ*،�SFMD^4�C�	�8��!��f���~�P�D�?����D�;sɓ�%;��4�F$�zT-������x�F��7~=����n��8�����OV�J!C��
�b?5C�n\.-`�����	����&/D�T�d��! wx9�"�zW��� �n� �@ *���g�>E� JcB0X�pD4�d�����(�yB�܇1Jh"N�&�8����/��DD�YE�Y����p<a�G,�Z�x�䙓�.%y�AW��4�P��M1v��K]��6E��DJ45���H��D[�QL��ui�X���Ss'J�Z>�`�F���:Q� �IK$3�B,�R`�?;־0D�1%!�d^�^J�}I�D�>��S����0)�D�@h�c��9��)�g�? ��C�a�`2P��DW�+���9q"OB}ғ@ֻ��a��:~��xʔ�����p�X	Ѵ�'�p���K��|:�E�
��DB�tu(9p�+L&9��ء�GC$98lq�j��{(Ļ�-��*w'F!>�ҁz �4�n��H*�ruj ʃ��(��O�8��SmIl�ՑpD6N�]8�'6V��`��'zVI���ڡ���ҮO<٣��渧H�>�8�i_&!�٘5"ي\��
"O�!�4����[�,�y�%Y Y�!�d�:	���c.M5i<��q���!���1���w�U.�dQ��ȓ'VJ!�B��a�䕡h�*��R��;�qOR`�S�U��0<���dG����%'O��#��h<�	X�[���q3B8&*R�qe�(Z�A��j^���?ɕ�X�\��-r�Thv@-�/�g�'�&pڵ��]��1(+iw�O�~���ش m(Q�b� )�(�i	�'�@�wd�#H�j �bD��2:��OD�sB,)��m2*L0Y��s�?�I���pAb%c��(�S�K�v�<B�	?:��m)peݤk2���p�U�28䳣�Y Q�Q�F�J��@�K#C�Q� ��$��It��iɡO�L����<|O�ʄ�U���5�� �k li[�eى9�rիЍ){J�ئ"ַİ?�t�ƐU�vd�T��qت���LQM��Ӓ�1i"�*Ũ)G;����9Q#@ 
�2[Āܗon���"OV�X�+�H�B�1PĆD���C�� �|�D��TD$I�0F�>�I2e��q�Uc ɺ�0>rH��"OH��-�|U��zQ���R`z���4kވ���%ٯb`����ŧd������yAh�9+n�5@�,O�T��{���eB�	��9s�dK�6�L0�6�X�v��M����2%K����Q�,u�0{@J@��lH�JU�O��O\��	�"_��i����)�@Iɰ�5R�&óa��5K��V�.qp]"�ȓ��!��+`X�š���lW�Q�OY�,�ָ
��
:F��&e�%�h��.�H[ػ���6OE�)��]�'!��25�
���
�G&��q5A�f�=c�@�<'��I4��W �Zv�O��FzBR�"�Ő0l��D������=i�����AR���l� ��	J��-��jih�g�$�Pt��'�����	�-�t���&T��t4��"V�c����ѭ�Y&��S)L�,b��O���V�#]3���M�q�h��'��	���Q��d�h���0 (���x�� �F�I��j�J���|��wQ���!�ڃ͂�ˀ(����'" }�@�C�<����Z"^����Q�^ N Q�N�9�u1�%���U�$�B��:��P5��`�a��=�����@[2@����H�<az�H�-چ��@�M�|�����V�V�a}BE�<Q��⑆J�9��H*���'�D��2mJ�z� E1�cM�U|8i�J~�N�l�\�1�Ɔl+�A:��ڢ�y�`X?d�.L!E��szzPA��^�Q��k�M�S�����F�%��s�AIo�p,FY��ɘ�$�:� &�!D�D;U̎T���@��@�MJ*�`�дR��xI���%�|��D��$<�3ړ[�*�R��؋7�ԕ2'�R7y�����&z~���/��`���ֈ��Q2�G�Ig�PЂOp�Ѡ���A��pR�;"��`�I��y�ʦ'�1�&�YC!��*r�e	��TΑ�7"OT0�q�Q��䈣��z+��ID�O4��Ħ�[x�KI��}Z�*\�u3�<�u�������	R�<������X(��'�8x�p�+�OVO���r�JѺ�H߭�0<�1$HG��pI^;Bi�&*o������F�%o6��� �!xֺ�
T/�J��<ʇi��:!��1GH�h��
N����8�Q�c�@
e��P���]���b)�z'�a�a= {!��!� ٙS�X�\ܥ[�+��.����{���n�B~�-�9��~�ug��x*j1�B��^�Zfai�<��i±+��<#�AQ�<�~�Z�&Ue?����	��m�k�~B�Q����H�@k|��A��d��,*����!�,Y��+�-L%#�\m�$i�1$����m`.��'Kw�-�,�Q���v�Q%D�B�x�dP�,d%��=�O�R��H:|�d)� ��)f�[R� ��%(W����wZ�`U�m(��?�D��ƯH*�d�0@.�0��Ez��͞K'v`�'��Y7X8�~�d@K+0	>T���̀A�-9p'�Q�<��kV-&���@�U�&!h�P���6(�b�Br랪�L�(bB�\mG���{W��q���c	��<�vL��}9����d�=1��BL�F���#ω+��i ڑwQ:<�$��OF{"�V(��j�9w��-
�����=y7�"r]P �����-)�����pi&��z��<`0�,9g���1�'>�d�!��/�<�c��/'����}��("��p�F=_�(���ؿj���BB�"~�Q,@�E�D �$�� �\�!+Q~h<�GK�=\��'A� =�.�CGV�y����u'��x�8���#?phՑ�4y��1��|�n����C�KN��������i.D���`$_ H���@�P�b��h2�JF���O8
�9Aƫ��&��� �_"M�����Q���S&��ȷ�� Q����&��$��Gz�ڄ�#4BT��&B�d�Y�`G�m��d;l��kдq�F���O�^ ��ɋHl�qQ$ϓS�x
S�ҝrD>㞌��O�%�Jd*c쉈$v��
� ��Ms��	Og�}k!j�|b6f�
H�1v�6��x��T 2��C*د'kִ�e˷#�V5Bs��=���"FL9M_�d+���"7�٩j�|ʢhށYt� �8T`�X�Ȇ+v�:�K��<D�4��5sv��� ��(��=0e[���_"<PRH�0[��5�S@7v|�����BC�I�w����	�$n�2���l��.-f���[ :n #C�
Z�.�)򭗽:F0���lI�Qq
�@r̜98�t��#dS
Lΐ�%' �0=�&`�I���b%i�8�� w�Kw�+ �Iӂ��(�#�K%G�X�J?�rSŏ�@CDy�EM[$��Ѳe6D�T�A˚�	>��HҸ.��td(ȅ�u�G�1�d 4���O*�a������h*n�5��"O| �pj�(�v�����ow��f�G@?Q�#�n�Xm��$G0���ɒ(�2����Kߘ�C"B�;Fz����AH���ONl��p�@��U�l@��B�2��l��'���P�ۅ7���a��=ר�����o�ܢ����L�kM�Q�d�(St���Oϭ�y�� 1�d�:�k��I.��J����yr�խa�v�����>G}�dY�(��y�O�%.��]�4~z	 '�'�yR"��v�ҁC�Ñg)�h(@Ł��yr"A�M��������]&�8rg�4�yr`�
8���I�8!TC�b���y�\��}�VF�'0~��$5�y2���t,X�!Y�.&��� D��yB�/:�8 r�NRB8��pd;�y�\V t5[����<z�@�y�7<��@�5���d�x/D�����ǚ9��b�"UZ@ ��5D��s��& =�}�`��4!�ir�2D���S��s2����OV�'�<��PE0D�|����%���Do�v�H�7 D�h���Y�t*���D�T9ZL��"��3D���ꘃf
Lg�ZSi˷�;D�H��d�<D8�􀒥�t�̰�H9D����d+�@��C!P $�q�7D�8S'LS)C7��Y�g&�H�j��?D������7v�\��)Hc
��Ȅ;D�$1�B$�hxQ`�0Y�X�'9�C䉵u�L�P#��>a��S�D�4Q^B�I(m��)s�M�섈�
�Y�B�	�fɰ��3U���M6b�C�ɵ �mc%.��B:\Ȁ M�B��C�	��~`;B�ͻ|e�EA2+��L�C�	�E�>p�R�Y�I$���0"o�B�	�i�&�EiZ2,���� '�B䉶c��k0��*~.D��N��6�0B�	�*�-��@F(�8�u+W8�@C�	�P��DV�sn�a��ۖ-�rB�I�P�:$�&<�A:@?8�BB�)� �1@��#!�6a�ǈɜv�B��`"O~���y�������PZ(�(�"Od�&C�mo��S$nl�\�"Ob%rv�˵OU 'hR�[�,4yg"O�T`�A�3v\���R)c��@�"OD����?E�Vc�����t�@"O��	 �����H*%�W�C��qa�"O̽�q��4~L�	�眷m|� b"O8��F�Ly�I�+��?bz)$"O�����s�(�*�i��LP���"O��P����>�S�fƐ&x��PF"O�r�̥7$2���e#b� �@"Ox`cG���k]���DZ�EaFY@�"OzL����:k@<9S�E�Tl�"Oưz�#�0T��$b�CN�EK��J`"OTl	��
~=�wC[=3 v�c�"Oܪq&ʒ]Q�xi���#a 1"O�|��Q�~��X���:G)���"Op܈`OQ}ZB|s�`�;+����"O(�aB�Ӳ[���3w.�,�t��"ONГ���:{h���Q	e�@��`"O�<0��;�A��-�)X��"O����@_�h�L��I�`g )(�"O�!{�b�o�z���j@J�9�"O�|q��,����c��,�F�S5"O��˃�� �(�h���)�Z��$"O�������d��!̀lҡ��"O^9(�� X��0FT?UB���"O�E���<���s�S�p�i(2"O��;��ŉF�����O
���7"Ox=�$mݞ�*���P�;�z�xW"O��HW��tQuAႁ	�
�"ONyh��
<.%��Q�k��"Xa�"OnQH藩{�U�+Wm�r�X�"O�<pD'��]��}BI�)H���&"O����I�R�0��˗}NxI"S"O@����*͸WnH)|V�D*�"OX�䈐9Qy��Rt-g��)"O,͊3J�:��xږ-��Di<q�"O���o��A�f��T��FtA�"OmՄɠ!��=8�]�l�49�f"O�$���Ӳu�ĭ�2�R�|$��"O ��mN�$���%ظ}�"O��1�� +.��@��:~$Ո$"O���d��LD�U�*6��0"OVcW×?�Б��Cʙ?"�{'"O�e��'@@�+����(�:�yB��za�@Eѽ6�xD0d=�y�bD�?��ڣ!��6��,j`��yBo��{�4��D��r�z`d�,�y��y؁pb58���3w'� �y-�!�8��#L<��3��N��y�ܢ^�V�p	N�F'��&��y/�w�����M�RY�.ɠ�y��"֤�;����O��
`&�:�y�+��h���ꉲC���H��"�yb��$uE������(���m��?)��H�N�qώd1p�.� 9JB�$4�Ѓ�9*�@˦D�����-5�X㨌{1 ���Om�Tz �� J*�}3�-Xj�H��'r�`��a��2�B�ˌ#_eXyq�'2����*7��<�O?�����"7�U��/1B��*w�/D��	���C.�`ˡfW[��؁�J-?�փͬ-��сCe5O(�(�B-lz��hFd��\f(ك�'�����D�� *q�6d�P�V�Ge9p�&���DR�Px(�@�J-����:*�cë
��O�Z���c>��B����R	(�S��2�<S7��y2"�
Ʈ��0�Ͼ"N4]Y�C��yBLJ��{��SU���/K(d2�B�	SRX��l�'P��B�	���S�BVؐ��K�Xb�2��q�!���*����W��-Ȑ#�,FW��t�MT�a~��H+m�2�*�+̒F�6��%�#p
�hS���i��(��@��	����Pt���E}Db�$Y�`�ɗ29��ġQ�L'Z,�d�\F!�䑅3��h
�f�P R�]���GQ4=;��铿q`l0�Lׄ)����,��c�B䉝*���{��s��aq�ܤQͶB�	2j�<,C�E�Dh�հ��G�QvnB�	��$P7�H�+p�
����Z�C�I0a'(�T!�<!�L����8>n��Tڧ�6�axo�*.�.!�G�Gz��=g���x/«,�d�z��-����ǂ�E���2��fx����7T�L�u��+2ޝ���;�(O<���C$7V�T�#�3)0��T��ʙ �@��٬dڨ� g"Oh���+�$��BS�ht�p�y�PX�"�#:' ́p�Ǧ#~Γ~ �=���42�P0@����a:إ��8�������Qr�����ԩSj
_=fya嗿ml� �0���?�>Y�k�,H��8�
��&Ҷ#'Y���HBm3z��q�+�/}�6ِ�`��?l ��E��_�.���)R�Ka�(�`��L��)����A�`�
��'��P=s�����R(h�'>uk����x{��:6��+�u��ݯ�yb��$��z5I��}����M�p��e 2��/T����'iY�2�t���O�9B� �*���1�RG���*"O^(��m�FC~<�#'P�r���;Q��2I��1�dƐ=u��+H�0����Q�q�μ���\3V�BԡJ��y=�{���>���ڷѠs�l(h�a��34a!���U���(�aƃ����Z�)c��!Ƅ�T>Q͘>�O�[���4GU�l9�	N�t:$�:J4���+�,)q.�d�XQ���U�<�r�׺'�����@k꤈���*r�Sr_;�?	�&j�bա��9�65)��ڸ=�X�T���d�p"OR����&�^��E.	k��X	S�E8zY��Z�U�X���f�̔3R��ENl�'� h�`j
��Tpwm�*E���H�vӺ��+ˉw�h��偖_�JKT��{j��Bs�	5]H�%�U�G�<����!`YІAY1A ��Yp�,��O���|IԢ�M�3a�{ H����5j{>Y@�F�J��e�R�	s�!�$�<�&ذ���U�|,7`�+uh4�s��� !Q�n�t���R�Ow�ڿ"H��۰"�E}���V�ho!���4��T��V�]�i��#~��`�	H�v���qR0 ���O��HDz򈑎~�f� ��T�1�t��#Ԗ��=	���91VMɰȑ�P���㜏:��=�"㈗Y��B%�m7�٘�I?�O%XXkN\W2�����fV�O��i�,
!g��J8:�>xJ�˛���IH�a�D�a��/-`Re8'�SGX!�o� ��ǈ�D,�z�"JzqРFOnx�\pD�EE�5�T�7��;��(���V�'Q4����X�<�
-(��I`�E��@uVD�WOH~��Ԃ��Z��9$������g�'G�e�m� >'�="�jC�"Z]���6�	�	�P�! �	X���Ș.;�|vԐ !���.�(��f��Li�nX�5Q��b�"��Wq4�H6�	.#n��xЋN'Q�N�8t
¤*�!��P1'1���dۢAd8�ʕ�B�}���M�&�1BcI���)�'"}�q���^~��"DCL�n���=`�0����x*T1���U92l��OP�Zt'ƨtj��^E^ �ӷu9|��F�/q�=��Iu�h=)�L�9{�� n��vUv���JZ1{W䅓wO�`�O��</�9��$�5e3����I g�����ߒ,N1��\���j>��!qb�N�!��"OhTKA!�e�T�� ��i�R��Ў�$ ) $�"}�W�T,"a�)�WO��3��Z�O�!�� hx�2�Чc���F)� ߘ�ڰ�|RiTݜ����Z���4�� �gI	�fz����'$ҀxC�<�n�o���@�')��@�DH�&��X橗)t�<E��'F,���%��U�L�v��'�FUZ j�"[�p��D�i�\Y�'{N�2�!"j6h�ᓞm�X�(�'�,�y&��1+����C��gm^\i�'zr�{k�$H��mX���Q����'�� �P�m7T٩#bM�M#����'�Li�d-U"Mt�	c��410&��=C�
402$����S�I��&ƭ!'&�q^�1�ȓ.�m+%"�!�Xy�"ٗ!�-�>A֥	vβx����ED	���!�\9X� ""�*9Mn	�.V�a��%��'���P*M�pęa�[	J9fq2S��
����L��n��] t�U's:����y�hʡj�,�-	�.����!D�x���F�kd��xTŗ-J��:�ς�[�n,�FF��AZlź�O����M����&>7M�������9}���k!/�\{�zB�_65�B�ѣW�<�1��7 '����.~�HJ@�V}"Ԛr�]��&����<Q�A�\�%}(�`�D#L�@�]���k>��6퇳!�� �J�G=�RQ��"�$�*׭R(�B�O<��!1�(����fN�/{zq�����']���B�5>/ҝ;����ѝw\���� #/C쨛�f e�h�#�',`�b �L�G� � *��['~<�B+��P�.!��'
p��V��F�O

4�o�g\�����|�|a2�'��i�7ß.\��͓z4-�G�N
%�r��ek�+J��-�'H�� K&�0=	ԩӠ�)J�@�P��x-M�*��U���'Ψ�dʂJ�M0νK�@\ Su�DyD"O~@��,�?=<V=K.�u~Y�Ө��(����=a���Oƕ� Y�"`
�ps�W{PI�"O�ya��GR���A"Q�=���"O|���vx$4��ᘹg�(��"O��U��D PU;���;!�@AC�"OZ���X�|��%�3�ʇe�D�"O�B#-�%�\����=nE�4��"O@)��쎉=h�(�&��3��S�"OpP���J�0��`�%�%=0��Е"O`y˧O�?���Ō�֨ɢ"O�y:��M�A�����2,�y"O��K*wv4ؑIR>A�1"O4��c��5bP�$a�#C
8���"O\E���'n�H��OA�^�܉%"O>��拍	 &}*�����* @"OZP��Ċ�
^ݱC�	�y��Q�S"O(0[$L��nd�A��3Ӹ�X0"O���W��6���D�l�&�Q"O�9�a����y�E�Z�jC"O��pMF����C��/|��r0"Oj,��Ό�=��2�*֡u0�S"Ot}a�,���C�
�2S��m�"O�̳1#�Hɰ%��k��b"O4h����U
�|��Ķ<��D"OH����P�OڰYxwϴYm�@�f"O*�Z���p�h�R�R;f�ܤ��"O�):��O�I�Xer�� �=�f�	"Od���fɔ�t�1�ᄑz��m#�"Oc�®-�\J� K�>y,!sV"Ob���ė�@<�֊�@|�TC�"O�D��%E�A(��jI��	Q��h�"OD9J�5�Y���]?�,��"O�d ���(I�Y��ˏ6q~�j�"O�����N�j.�b�_=n���"O���!a�j<����,c>�d"O������@��R�۠A��H��"O� ���$-�+[���;e�M��`J�"O� ��柨@�a�j�i1����"O�`ֈ���pZ�^��I�d"O�] �B��˖��3�7.�	�"O��3wi_	H�j�)s�٥iX(]k�"Ob�B�Ղe�:a��� X�M�T"Oz���e�2j^�LWH��&ѷP�!�$�qH6��Fc�$98�42WE��!��"E��TpD-A<yS�*��!�ӵ�\�!k��d!jx��*�	;�!򤟋aN 8��j�Q- i��FF�[����,ȇ �D���Jģ*���P�+|�tɳe;��=BB��fxTTA�=D�����J7w�����>UV��=D�l������l��%L�B��s@<D�P�ъR�k�
�����cX�m8D��A�â���y�+�]�PX��7D��ZΌ"9��z�bDv�����*4D���C_1-:V��ՃޯwZ�TY"N2D�؃�+��5��Ж�ɱ(�� i@5D�؉u;l�1��Ҿ6'<���"3D�a0�Z >~���or�q��K$D�$���X�t��!�KK�r[�l+��/D�$�` �
x�v�zv懪B>���!h#D��P�.' =�2G�:nr��"�?D�8�!%�8>���k�G��2����:D��ٳ�Х1B���G�O�؄��K.D��S䝏l�l@�Mð|��x3��-D�z'��8�@sG�.����׭�ON��1���M���:?�O�����n<�uJ�*}��x�Ӂ=[�����T�1�6�ڷ͇>
ջ].�����0|Z��"x�kf!ϡd[�}Ð�� u	N%��	1f�J�E����	Z�������n�V]R!B$>4��2v�W�?�-i�U2!E �K# �c�z!����o>Y��M֢H��R֬��yX`agL�[�f)����ę���%��vǶ��	C�T��j�+�� O�l;Rj�`g2PB��/f����$�6#�xf�~����c�8eR5XE�st��cC �-;�CUUuX��!g��87��
�'Vp �#q�ņ)i�� Vk_qQ�����\h�����.MFD{'���P�%�?�x��tdD1��������2���o�1WN����Ц%�!�D@�&�V2U��9���f���!��or"ٲ�o�4W�M���H�&�!��ĵh�t81�	ȧ
@,x�$��V!��O�"�b%���N8l%�Yp�LN�-&!�ϭvt��3B=jY07��4Q~!��hb�����!O��pp��l�!��|}����Ŏ9���SB�.0!�dU�n�^%�7ᑃ��1B
�I !����Z�뤄Ł ��M��gG�m!��;s"��5l�!�q`$Ǟ�4!��*�jmZ֌��X�U�c��R�!�d�>&�2QF��&��zGhVF�!�DՆ�VZ�Z�B,��
��`r%�ȓw|t0��	��͊��!^i���ȓ]L�E�v�Z:_b��,�$!��^Y��h� ��,���K�ImRE�ȓ7�D��
��
��uK���Q%(8�ȓxb�E_�D�E�
A�豅�"�p�˂�^�YCj��bcQ$z H�ȓe��PCV$���҇G_+m�����g���#��!k�<��
��n>N��ȓ$�{��Q�TQ`��֬��t�vU��Z�:����0�"�ʅjG�/�Y��s5�L�3�ay���t���pz��ȓ�@)2�G�RD��)�!��Fʨ�ȓkȤ���#ܿ,7v-a���mT0��ȓ�<���*'���V�	-ɴ���S�? rڦ���Q1H��GGNp1�"O�i05���X��$��G��Z���"O��BG,X��9ڦ&
�/3VI�"O`�;`�(>�\<`e��,=+����"O����e'�3��f��U!�"O&E��W�%���IC	�Xu�Ż�"Of���UHp䈢#��HB 5"O茻��+*8��y��$
��V"O� !D ��0�j�cs�9t!faڦ"ODa�� �'��-bQM��Z�Hv"Oh���ʐ9Z| qgLy|���"O���VH��� ���Y�R�͈@"Od<br���Td��n�s�(�d"Oa	��ɲH��1b��9--�\b�"O����-��p/P���Y<`��"O&�kҏT�I���+�J�u�"Oj���L��E�8�vˀ� Q0ub�"O�r���#Y�Qp��3#6�H�"O
P7nb��Y��j�*���""O����#�d}6y�2��2��)�g"O�D
a�60;�T°��T�@} "O�0�A��#T�j��%�+���;�"O�Ż��[n�xa�dӫZP�D"O���X� ˄�2 !��V%~y!�"ON��u)��7MH�Hp��03��yp"O`�s�gH>�8TS�C\��5�"Ox%+���#*pN d"ŵx�H	 "O΄ ��i��E#"@ڧcf�"O��a��H�p������I2��"O�\b��R
����& �5�����"O�������������WYN��g"OJM���Ɛ{=��s�iM�g@x���"O��Y�	�
pFҵ���ʹ��hrT"O: ����z��8v/H� ��,��"O�-B���9Jt<x0L�	Q��K�"O�P�����b��$����	<<q)C"O�5"�ψՀ��S�ƌg6��W"O���Öz��a�v$U;��HA�"O�33 �x�P"3Q�hl�!"O���6 c����?Ј�z�^%�yr���0�`<�'�	�2��8RT�.�y"�ʛY�`�C�))N����)�yBe�(*�m��jB"1�9R�O�y�Z��U��L�*f��X�KK*�y�D�5~k�e�3�\� ���
L]�y+S�Q�2��c�
�"��J�L�'�y�aD,O�@ъ�lJ){�gɯ�yrB2^��]��ݨ9P68�5k_�y�cZ�K� ʒA�1�����P�y��&�fXˁ���<[Ih�
�/�y�잙��Aǈ��8�%PAC��yrf��s�tek�iޚg��	k�'��y�K�f9ʅ��'.-]�	���7�yb)�#6-Pp0���"�����y!Q`�0xq�.���h�K�$�y�b�����ab��'��8����y"�Y� 7H�:ׇH�zt2�re��y���7�����tn^x ���:�y�B
�T�j�#"�o��p�BɁ�y⇊8f�yz���:�Q���B�y�k�v#��x��+B6 ���K�yrL��*��D	 �&e�azt����y�J��>�*s`�+�������y)��'F,`cT�?y�h�r ��2�y
� �U�a��2&��4�K!�yR�"O0](�g�d�AX�����"O"
a���q��X@��	3Y�0s"Ot����Z$X�Ġ`0bH�J�yI�"O�)�P�۳'�f���t���"O��΁�\�f��u
�A�R�2F"OF,He��!Z�p)�H_5hؘH�"On`��%$$���RrjX�<���i"O>(c���.�� �镐g���s�"O�ir���~�������U3�"Oƥ���>F+I"o�A��H��"O�����ܨJ�MF�߻ �ThP"O�]���" d4�r�զ��E"O�1p�J�\��1�R���'�j���"O^ͺS��.��]� oT�]����"Ov���팗w4�c���	��t��"O�)���E�J���D��,��"OV�1C�6�<�p�̭"�0�0 "OLq�ċA�ܐ4���0��C "O�4I�N��H&�8q$�_(l:�"O �%� p�dhdN/�8��B"O��1k��_�`��AD��qb"O|�G��"@���S�+7�x%kb"O|���߻<�ƌ֙2��p�"O�Di[=��}�0F��fܨ,2�"O }	��׃p�2���]*=�|j6"O�%����[B�1!ՉE�bD��"O�A��JW`DD��?���"O�T�� �l9��+,D��A2"ORm��	ػAr����M9@�]��"O�p� d�8�4qƦG-.\U�"O^m	D�K�iW�0KFE^d����"O�xH�Β̱4&״vm�1P"OH��J��N��Ukae���8�F"O���Ē*�X�C� g;,���"O���K�["(��#6P貗"O�4��E��`�V�s6��+� �d"Ob���3s�����ƊD���u"O�d(C�F& <�#��1;@ܩ�"O�Ie㐽L��	���B�P7��"O��j� �-����d�`���"O4Da/	59�bb]�'����"O.����ߝ@�:�Z�k��]���e"O�X�K� ��ԃa�)[�a�"O�+7��
!c �y�g��n/����"O���
��E0�@r1��)S�\�"O���BH�_��#�l�&��"O-�%ٻ=u`� !|��H�"O�u�t���p^�$H�%����U"O��l��Z)N��K� &����A"O<���#� <�4k�iI?A`E�"Oⴁ�j����)�����@Q"O���d��4��`Rh�P�"���"O�1���h���!F���!F"O����m�A�
`ْ�0�*5)�"O��
�B݊\�EZ�$M-9�<�:�"O.�R�gVc�D��"��z�ڱ�"O�h� 6Ҍ�t"���$��"O����,B�@�~��@�P"O�X�3BWs$�$\(H�4�p�"OH��䃲⤡�r��Z���˦"O�=�
=D4e"��0[��]A�"O �KQҩu�V�e�q��!�"O�l��Ů��I�'�Lu��{6"O� �-��`V��Z��Qߎ|c�1�t"ON}
wM�i��B#[#D<$0�"O2=婅���c'��Oj���"O��)Â��Y�Rt���ـ"KHI{B"O(I�5��#x�	�c�
20�#"Oڬ��,Ba�Z�C�� f���"Oޅr@�B?����`C)) �i��"O:$4͓1Y��T�w��(
hl��"Oy��E&��X�����L��"O�dA���`;���6q�^��"O�}	s'�'68�Z1�%��mT"O���q$�' nb��%
�v��К"O�����B�S
�r��*d�F%�0"O�(�l�h7+
�=��$��gO�<�G��lr��G̙)��	d,Ge�<Ѱ��?`�Kg%]R۴�@!��]�<!��_�\���25k��9Y�IQ��_�<��`��F�0�`%TDY%˓X�<a��#X��\��&M08r�P���W�<5aٖxʜ�i��M�.�U`pI�V�<9��%I�}��؄ZJH�K�� H�<q��/p��v	�*���@B�h�<�c�ѣ)�ٺFQ%x��?H<C�I���{���`������^�.C�I�IϾ@��LK#�-��L
8^ C�ɚ �x�f�d,h��a����B�	�xx�RLۦu*]r�`���B��!V�bp��`�T�^�y�)�dB�I:��tB�]���B%�^�kSXB�	64���ĵg�x��A&%nC��}��;v�ª-�"�y�,�YExC�ɾ_�ltb�"��DE�����U�SQ"B�	:�j�*���7��
T�@�HRC�l�x��ݧej洡��S�A_C�I=P:��tca���wM�)t��C�ɑ����V�6�l�e@C��B�Ɇ���������ʧ�ոfuzB�I l2�%��_�,�{5,ո*3~B�Ƀ*�@7���=�4=��l]#K9�C�	(n(�&��$��Ө�n`�C�I:;� @  �P   b
  t    �   �(  �2  �8  	?  LE  �K  �Q  X  Z^  �d  �j  &q  nw  �}  9�   `� u�	����Zv)C�'ll\�0"Ez+�D��4��M;�(��<1�Y̟H��Y����4gï���b�愙2A��11��A�"�Sb��{mX���c�u���2��t��?U���C�}����B&PVD�S��(*��P�\��h�'�#4�Ibr�λV��݊Wh���ğ��5�^��@[���m&��P���Z�[/�?���F1���۶��j���Ӕ:o�'��'����ʘd�Z��ܼJ���$��'�Rh0w�mӾʓ�?aŮ�����?i$�^cᔽɇG�8m
.2��?!��?����?��C�%�?�p�G~��O���SQ��=J=��w�Ҧh2L`�"O g��3]B���!"�	8�U��S��Fxr�Oh����H����� 
��=�BZ�vz��MU::�';2�'���'��'3�Sμ��H�w?"A��=�"�A��@�ߴr0�v)|��	�'1�7�IҦ�Bߴ���'6�\�č<���ӤI�&	�=���I�-��>m�#T�&�����"4u�!��L�H���k�]��C'Wv�|lm�+�M[�i3��>�ƙid���X�"�5��9M��)R�܈cP���'S�a�ĨKUf�]ñ���JI
��5O˄M��Y�g���nZ,�M�B��6
ظ@mF�EI�Q���É�jU�2��t(F���ix�7�P�2��>&P�� �
,]N|��JH��la#  &Y��aa�e�a����q ��A���M�Ҳi�86mʱ0e@D�� r8p��eU�LL���e�M�4�3���%v��(bcR̦�aT��&<�pE{0�	#`|K��ݟ��?Î�"Y����eڎY�<<`afO�?)���'�R��,�r7m%��������-H�"�W����\�'�r�'�rD	4�\9��,b$�1m�O6��AĐ�e�X:}�F)�7�ù�0<!� �7�TmR7J&yq���4}w��{�5鰑��Ҵ}�؄(r��cԧ�?����N8'M��i�"ϵZҨ�c�
#q��'<b��S�D���bG��T�v-��,ܦR
>����H�A�	h�x!������,�6,�O���k�l)�'�y�*�Č8��ˬ}VM1��W��yB�V4C=,�X� �A��+���y"�YE��E��<_�Ț��y���FY��{�o�'��2@� �y"�µG_����Z�&�����Z=�y�oU�|
|Q �$��L��H��I��?1P��#<E����"R`�����)y�1i���1{�!���uΈ@�N�[L!2�T)!�!��G�L�uȌ�0�2����!�I*a����i�c�fl�a��*x�!��=<�(�ƚ&z��9`���o�!��ɶL6��3U�C!P�(7Ð�=J��=��|��	�&�^ir�K�����O�I��C��� ����(�����t��C�ɹ+Jс��C*a��0PL�%O_fC��lgȀ��b�Ysf��9n`C�Iv0�z���/c"���l�����dI�a.�m`~�^H�Ȍ�`�/t�f��s�ڙ�?	,O��d�Of�$R���	��Һ8�\�堋������*nXl��"��Jb��S�#O���!Ę�*��]k B�Av�6̀�>�T�	�ش(dɋ�gɢ:�I ��p`F�����UP�4�?ya��.���a�%dbI�Zbd�'�哑}���ʳ��{�Du�4	֨V6���\�t"	�M,�AEҴ	�j�����OV�OB���c�8_m1��|ޕ`ea���Z��I�&���q�<�������YW(��<��Y��s�<�@K�
��)���ݟ���Yv�l�<A�@�0��0�vKA���1fO�j�<9#g�8T�P�ye�[��hC/Fi�<��ȍ�0`��I�q�n\I#� ��M�H>��A������?�����dщe���T�i��i��9�Xo�:��3�iu��+�F_)����'p�Q�j��f�b�1c�[�R��5�Y��R-R� 3�����-�O�^!8�+Aq?�U�\�~����!*z����pC��MSt_��W��O�c>�D�O��D���LB(yN~0��J�Vu`��Di�6�X�z3��	:n����P].H�'��6-զ)%����?ɕ'��H� ��'�<�R'� 76�`�0���	��7��O����O����'9��9uHQ���EZ&愥7����ŧ\0�T�Yҫ=U��C�Y�����=x���p'.�:<Δ�2��@�X;�@�fM�A�0��
�+S��(!�e%�c[V�3DH
�<	*F�Y�5x�Xb��џ���4����O����O4���O$�	��٣�0b�V���ٺm^H����͢,�����

���j"C�	5�M����)Lv���OR���OD�	���Ȑ`����Ëc�B�'���
��'T�>������S��=d"��Q��� `��dI�G8�Ps�HW^����B�' ��a�k
�#��)��~r��׌���=�/�4��@�k�$#?!�Q�P�4%	��@��w�Y8XQ��1f�Ԉ�̒O��7LOp �1�cu� ���2�$%���'����P�2]NI��Y%	Q�8�ꁇ�S�lx����MkO~��O���'\������I��g	��Xl.]@&�'�o�@��Y��֗V�xa�;O>�u�F�'�~u��iO�}Ʋ0��+?q��_�{�R�`��U�DI�گ��q ��6�ԏQ`\y�Pc�6qrd]���䆮mcR�hӼ��O&����I����c oE#m���L7a~��O�d�O��$(�b�Ф�%K��	�"��58џ�q��)̊dК�R�H�C��H�dB�<	�ꓑ��� Y�m����I��8�'Ѯ���D$x�����S����Y�����g*.Ip�O{�i�n;����CGϷo	��{�MU��,l��, ,��^(,��c>-�u�>���"UH�Û7�v� ��ϟd��ş�q�m�ݟ��|�'�B�Y�fmLْ�M�qm����	�V�:">a�y��o�� 3��?7�~ة� R���\P}�[j��'�������鈶Sa����\�DP�HK��[�p��a��惡��؟��	]y2��D�)@p�ٲQ��*��		0��-���~�t���V۴E�@'�6 �ɦfͧM����S ѽ"̤"3�ǁ|<���iP3>q�>	��<D���h'� ��F�Y`�d�	˟L&�h��J��<a��ЧU�v][ŋ�7o��(���y�L�,�����	{�Q�ǂ����	gy⇘50��$}9�oܹ!��S0I�&����C�'�����	џ��E���T�#%��$���g�io��#ɽ>�X(Ԍ��(���	�1*
Y�"���U����7�^���Y���t�(���74����F�5?��>q��Rџ��Ia~�P�_q��s���`���A�!��Oj��d� =7L,��ɓ.*M��R�J,�2��OJ�Ӣ$͑|2H����-tRs@�'�	�r�N�A�O�K���'K~� ���G�Rt�+L� H���'��L�?r��
q�~L�E��h�ʦ#|��V%t#�uaV�]+!���0�h�q~��'a.���f�Q���H�=�]�}z�o�Bl�F�T�p�7��p~2���?����h�����G� ��`�	�O���3w̖`�0C�I �P��T+7J����Po�(0�?��퓌��İ����7�t����Mo@��']�	8c���֟p�I��4�'H�����T�$�H�g>�MD�P�
���F��O�M�u�R?P�1�1OX�EB�0v]+cƆ�W� ʰGI�D4�tAЇ{�>�	��Gs9(b>��P�>��� �h�,@�e_�l���
g����'�B]1��?����ڥ'� 9�@&u��lQ�Jܐf%�C�I�V���y�'t�|eI�P
>|�˓\c������9�t��G�C*dB�)r�<O�"2m�O��O8���<�|jm�)i	�#��-֨ڴ�.`8�+`Ƃ�u�@5 3D��z|�yb#�,A?��Ҁ�!=(]#��P�  
P.������S�]SǴixг���
�r� �H�"�&��s��!e2	hP�'�B�h�'@��I�%O ���`%X49k��R�'p�H
�.�%,a�����RHm:\XJ>W�H�?y#Iz���B#Vm�(8�I�U1���	VR�<��Ài���G��X+�=T�B�	�H;���'�/�`P�%�~B�ɰ��12����xȑ-P^NB�I�:ԌIѽ*��d�)K�W8<B�I�oaB)�ЁK�bѲ���>�Ң=��
�g�O�u����E�"�����s
�'<�D�q`��*Y����싺i�4x	�'����K[9U^�Bƭ�*j2�#	�'���"��%On�j%e_ 	٪<;�'^|� �e�[�b��$dI�Ѡ���'q}����<q7�0Tj�>q|���7�F0Dx��)�p�(lZf���Ur�Բ&��?�(C�	' �D�f��/I��gk�*�
�':�-�p��kv�e�ɣd?jEs�'��(Z��r�~@$.a��л
�'h6j���-t�:�cK]�G��
�'��T��*��h��� f�$C���2)O\0�'�,��BG'5`��gƮ7���3��� L�9bJ.��=� IXW��0�"O8�V���r�
4Q4o��Hʬ��"O\Q�mH<�Ak�'��.1"�"O* Y�D�=�D����P�Pm�Ha�'�n���'� ���޹��<���${�&��'�X�k�MUh�K�L�w��ͪ�'�����0�*�$�Z�v�B���'Hz�/�LTԁA$D6�ٳ�'4IÆʌ*54�$�3 ��D+P���''`h��E�!bY� �7-^����d�g�Q?=që�:A����K#pA�@���(D��J3��r��@K���#V�؜لh'D��P���c�|�B���C*�x0�1D�`9���s����"�2#Q��31e$D��! ����JWo�,t��K�� D��oZR��]��Vԕ����OX(�R�)�iv0��Ø�ef��1H�<p��l8�'*|��c�>������ �n�|�
�'f�!�g��e|�����kEv�Q
�'��8R�mʏ|XPj�0f�Q	�'!b`�¬�1/���Y^�X-)
�'��-J`��)o~P�0�Z'�\1c(OZA��'���Gn��ǂK�&�����'{��ʵ�C�h����e��%�Z1��'">�1�U(r�>t�@�d�R5��'NL�Q��w3d�����X�z��'����a)?ky�	i��;i�ma�D�8���56y+1]�H4�劗��/�~�ȓE���h
8c`ѢD9A74��l�F��f������0o�
qi�Շ�b+��V�U�A���� �!�����>=���FOXA$��bB�pn1��%&��cC䈸K�ڍ�᭎��P�F{2�V����X�I� 0~U��	3E���PC"O:��`΀�+�����#�0����"Ol��� �0��Mi��M>G� QU"O�t�2l?"_�0�jQ0`�Pب�"O���f��M��B��Ψ�2A��"O�-��S*�N̸7g��vm����'B�X���S�i+�DXr�E�x[� "[�-#,��ȓ,|��2$RJ(�9��_�5��$�ȓ^M�l"㥆�'/
8��#	_H��ȓhT�M���Ā#� e��EűWt䰆���]Y H8����F�-������������>?�Y�WP�	���'�{	�[L��Q�;�*uztlB$)4ZՄȓf �ٶiʮh{�����ģV�N��d�p�S.�9"���2-47t��ȓb(HP�'��:�����%M-lTT�ȓ�����)��X������,i�pd��	���	9 *�AЦ��tԺ���OI�d�*B�I�)���b��m�Xh�Q�>jB䉓f*�K �@0�Dp�%�3�B�	\�RL3@��w,0���c��C䉖H�6���oT�={@Q36�]�eƔB�I	Kg���n���k�F��:���=��-f�O�%:�����X�ac��*yp�'!�l�#�ƎP��I���.�p��'���7&r	��$���m�P$a�'Ǻ���:7��
%mȋ2�\���'�4)�ձ�h��쒴9�x�1�'��*�(��^�!.�	}�^4a�]t\Ex����Q�,"�-�0r|;2�R�C��9O�Ȥ�nѬ{�`���ێZ6B�)� >��1 ��L�ZU�$K�11}����"OT�;6��q���y|��9�"O*�j>I��JϿ6��v"O`l���O�H(�ۆم�����Y��Z�$�OJ��pƑ��q�p�%5�|�"O�E���L�	K�c�R# ��%"�"OP(@kX�+7�%��1b�L��!"OL��$�_�x,�<��-�~��"O�K ��-@���cD�E6 ���'���:�'��Ac"��nl\��,G�m��;�'~<e6�֥g�Bic�-T;L�'&�����C#����!�Z'K����ȓO2]��!�~9PD����>�� ��VXԹ����+vT�@��9BK4T�ȓ@ʼmBPO	2M�ջԡY�w �pD{2�O�����t#��	ֶ��胦f�\�I�"Oĸ{GAҚP�mj�	�JOv8�"O��O�J���f�i1��2d"O��h�/D(V��`1��ɵR�ܤ��"OHp��C^�4���uA�!]�b$ V"O�Y�d��?MF��9D@^/Pr�tB��'9V(���
���KAh��A�0���&���%(�R��z�VA #���<���ȓ\��9�凚%`FPP�dP�aZ���qFx]�qN�s�I�Q�0s,���[����-�1? ��!K�,��H����8еO��	z�T��eH�s��u�'i�R�tL�!�цF�`!�`ҥ e�ȓ@�6���% MonP��٬2�0��_��3�h��
+R��ֽG���ȓc^�(q%�Äl\�[ģ�Ec4��ȓ��`�E�	!ۊ��$_�2��Ʌ��*M?T�ɐqu�a�f��<��иg�E�C�$bZ�A !�*�<8�I�$�lC䉵
Yb@�Z�I܍�⫔3*�B�I]a���BW�2e�)���6Z�B�ɱw�f�D�!�ę�f@
���C�I�2Z�)�#(�%/Ӝ�"�h��idz�=�FSi�O��a� ��d�S�M��?���9�'�>�H A?2^\������a�x���'k^q���"����w��'��i�'B$1����%��N�TD�3�'�d���a�*�$Qc'`T�F��pI�'��A�@36���Y�Y�
��=K��K���Dx��	������F� ?�հ��?^�C��*g�@�j���O�u�ר݂_ٮC䉍9�l,K��xD���.]|�8C��kd��A�ԿNuz��r�\$tC��R圝���Շ*�l�-�=#�
C�	����J�o�zq)����ʓW@H��	8k+�̚�E^
K��T�b���;JB�	!�� �	�\�d�#f�Y�-�bC�IE�a�m��~1�d�Y;~�$C�IG}l�����P���R'ͧf�B�	':{��#Vj��*H���IV����Ȼ6����v,�=a��];b����e�i�<9E	;~���b��NeΌ��Nb�<��k�l�����*�x��KY]�<��n�=L��wA��b�W��O�<�3撨�v-s�W!D���0j�L�<a�I$%���K3�V�@�Ry`f��S�'������I�~��Y�l�1	x��R!݂A!�$� H�P@�bƯNzx���.[�i=!�D<g�ȩ��Y%rt�Kկ�q9!�� ����[8nhQzWL�+�h�"O$�+V�R�m�d��&$p��"OJPv�����Ct��'T�֘���'��4S���әf��m��F����x0끕sG��ȓǴ�Y7-_&W,��:w�U�k<���&%��fNu�C�W�@�ȓq[�<�1��xx��
��k�2�ȓ������J��0y���0>�5����H�-�zӦ19�.Q�/E��'��`	���5Qʉ��N�,�c�&%D�`�֫��RJ��B�8��HƧ'D�����D�R4���� �8D���rFAj�r�t��TF���T�6D�,@pM	�3ۂ�cT�T��	��5�O4� ��O��q���(l˳*��A��0ӗ"Oj(p� ]�O8�k'hQ��\�3"O�\8�kA�=S�H*�M(j$���"OTq���E�2ے���K�yK�$S�"O�ဎ�edP���	$�&dh�"O�q�燞,F4��Ek�����I�8�~���ѳ	[D3�"�9
��iv�u�<Y1j���Y�E��#��|�&�n�<���� C��h�"̮?�JpQ ,�h�<9pjA3x����*�;܊��� d�<�g�ܕ
��MC�$�'c���� ]�<���W �ʡyk��<r)P\֟(��E#�S�Oux�HDHԷ��e���H�"O�И���&n�]�CCE�XX��"O��҆J+��i���q�>y��"O��NY�3�E� Q=�*���"O��Bd\�@�a�3�p�CO���.�'  9��ٳL�e�4m�O>�'f$�'�5����� _"U)�$B�#�(��
Ů?��I֟ �	��2�Έ;�ظ��A�:T�z��|��Ft��tj�7[#4���?K��L8���k��u���ȾA�l�m�!�����E�0�DqȤ�T,���`�}�'�ȸ��?���癨?Y����η{���բH:��D*�O�q:�T�7���X4�T
-�NEYA�'[�ʓ
��F�X��У�*R���'e��S�b�R���<a*�r���O2��?�}xp��+�p��!��O��r)�0��$�1��/렌�)�l�<Y�͍�E!ni�t(��r���̓	�4l#��R=x�Rm!d�r|7�͐VQ>ay�`ٌq��Ų��Dsp�{ �h�� �*�O��D!?%?��'{p��4&C,e(R ��A��|:ؐy
�'�>M�����&`��o�b�ۉ��N�O�q�/�5;��}Z�.�X����'�剳2�Q��ן��I��|����k�&O2Z(s3dK�Vy�(��Ё�~ȃW�'h�#fဪh�L=!ʟ����J��4�T(Ǉ#8jp*�vC��l���A���}��4�O���=P#�#.�Q��և_(�I�n�s~���?���hO��	I�!	��<�`(1�����(B�I<:D.1x�ox�!�H�;0�˳�'h�#=�'�?�,OND)@"dm���Җp:���X:B���O*�D�O��Şc�����T�SÒ��d��7�*%�B��^o2P*�~'�D	 �'?��{�쐃I�K�Ńy������.R�ȍiG)�+f:�\�d�iE�l��$ܹ1��oЀT�܅��&�P)�=9qS�|���If�'�65�4�1%�#t(�$8O�X�'<E/�� �J�,Q�M���,O��l�T�'ցp��$��(Gudh"KW-Rm�u�� ����'m��'��Ǜ=pDp�$���e������O�B7<F�q�1��a��,S���@�D��@�b] �]m��
�, �Û�H�
��JG#wnܑz��DN�'C~x����?���4�'����慐 :M��3�Ȇ��:�O����CO������Yf��	s��'0.ʓ)�T���(���-��#_�&\ؖ'�&t���nӠ�d�<+���D�O���!Y�#��5�J
a���i���O�uC1��%f#v<��ׅPa"	�)�6����e�J�E٘Y����7��u�B� w�]�. Ls ��M��KK�O��aaH�*��{�'��YA�a؟'�b�8���?	�O�O��)� 5"�k�`�rM�c��px ��"O�s&d�Yz`y��(��$�퉇�ȟ�4 �k��aeoƖZ��Yh���~=�˓�p�2v�i����'>P��I6 ��Ź5�է1 h�	%e�hv8 ���?�1�H�f>��e�Ji����<P�&1zB��Hr��7�r}JV�~����Y_`0d�b�4b*�ɓZX�T�S`U�x�)�$�ʨ�*�e�D��ٟ���R����$`�61�j 2q�A�/�lq�"���y�b�9{
r�Y�$�����G��?IP�i>U��G���W��`�Q���H�.��5���Dՙr{6`�m�/�j�D(E�n�!�$ʔ[�8H[��M/)D`S�G
�m�!�����*�─����,�!����9�f�W
K��Q�-Ѓ2�!��� ����(�_�"�A ,X�C�џsci� ����O���1��̓#vM�eIC,�|�����D�(���OR��;���9G��B,J�` *�'K��jXw۔$Kt�۠�ܤ2���T!v�+��$S	S���*� �d��I@�hOq����%(��r��x>4�Z�̻#�H�D|����?�5�iVГ�nH�햟fO���'J��*3t��3S�\�	o�𰃫��uqt�;��.w����Rj(�Of�'x��J�x�M*S��>O�Z5S)O`�צE��Q�'���O��h�b�(7�����эssj�#0�'jўq �
�����Y�(�@�)��eO�c>��I�?3���(�+M�$PJ≇9�M��X]�y�'@>�����?����?��'L4�zb�B�+�Hő��W"�)"�l�)x�F�'���Jg�'E�B�6����u��#�1g
l,�T��|�8!�v��.~4�}P�@�O���"m&��Iĺ+��?����?y�'DD0 R�õE��KG���S����D��?��S���+���yrf�5�����S�_?a�"Gs���q#	?�$�����Oxx9��'��HR��~�'�?q�����y8@�y J�1T�H�he��
I�lL���'�d���?�ɇ��?q�'�Z����M��T����Qf���'�ܷ`��I:�!�"��&:O����'�bĔ ��I�O6�$�B�鶄̟{�*����&S#���\"k���	�h}N���O^%���?��'�T�x��M+�gǞKtD�cF��j����*ޑ �n�d�i��$֖9-�7�	��]��;r����f�^6�`
�+|��ic��3c3����9`�DO8;oR�'U�$�'W�$�g���ƮO0ɺ��X�W��ciƅU�L6@�^�����<����?�|�' .�'�,~%h���)e���ئ"O̭	g�V�^��u.��Yny��V�0�'��'�'�2�
�G*n�T�ϳ2k�u/�(2�"=��T?�Y%ˇ�1�4d���[ !��,��+D��`�#�=x�����J��2����)D�|�rH�h��pՅI6"b���)D����	%E:8G%e�A)t�"D��r��Y"L�j5h ��2 ʢ p��?D�ȃc�Q~56�`qAS�m1��ɐ&!D���~1\��u@��%`��Ă�U�!��ϯz9�e[ y�2}��/qy!��X�z�<�!O�Q�谫�B �ip!�$�<�3%�&(��SU�RR!�dֲ�V(r�ΰ;}��d#ð2���E{ʟ�)�L�6t� ��� A��"O`�[S�C*X�u���ŌG���c��D�,/�Py�n+
�x��&	' 6�Rҏ�U����b+�5~�Qc�ʍ*C  ��ō�:��S�2H����D���h�P�.�/+X�"̂4x�)+F���
�j1Ȁ�o p��0���B8X�/Q� �$�ZF�D- ��ہdi���s�̴^J�0Ӄ�ԡ")��z�ݳ9֛��?�$%��m�?2�i 5�Y��D�O�Ո�E�O|c��gy©$�U��V��4h�e�R�hO�)��)�S*a^ő$+���Z`��aVOD����'�1O����W�n�ze�F�ɮ��B"O	�@��|g6f�!�V�c��'u�<�"�/y�$D���*O�f*��?�<7��O��$�O0��E�"�����Oj��O����������Q H�������>N�%Kb�"^
^����
��l���;�����N�*���P��a�v@W7~�l�Y�2QtlǮ�H���F�)Z~��ER��J�I�<$�Zؐǃ	�S�0amZ���$F<�O�����R�J�r������d�Jgゝc�!�䘧*�Ҽ�b�B]Rd�&�շ��c{����Od�!;|��N�8 ł�"v�� L�X���*-�z�bH&Д�"�6f?�܆�S�? �e�֮��`p���� ƈ@ʒ4)�"O>�ҩY�Q�੃����W���"O�C%e	�^/�z@�Ǚ^�(aP"OVXB�&�0	U x �=�� ��"O`Q��JA�r]S�n	2}���a"O�`*���@���Ц-�/���"Oڔ�tK�7�"�����.]��"O��#�S!V��5��Ô1�P��`"O�iXŎ�P֪��(^o���ж"Op���g�<��1 a�0Y8�A0�"OJ��K܃(j�YE/ ,�	�"O6�q�$��gM�d)5d�2}L����"Ol���d
���)%S$��}�G"Oj�3q������bmP9:�аr1"OBԨ�D:���S�$X�|W�R�<�N��W�~<@p�2{@ EHO�<9dmH���(	Yl���tE�<1r��
����P��/�t�Ps�E�<����]zLA����+g1�u�2�W�<��ђn���1U�lSv�r�%�z�<������a�$�$@����#N\�<�'	��S�P`��#�M}�)1�N�[�<��e\�8M�ѡGLP/D Je#�/�Y�<�p��b�gX()����E�q�<���>jE�ԯT2��L8T�n�<鑡F6)���#���/B�1�en�c�<)���9G�P�����S���K�CV�<�S�(\�	��牗,P����BY�<ن@D�PWj����Mva����I�<��.P�_��iyp)ѓRlh�$��A�<�V�'R�Z]��߹]WjLڳ��e�<��h�6�Ass�G�K�n�2�k�<�t��+4����F�M�x\� ͝j�<a�MN�@��@1R�u!~�P@�/T���v�X@|��h%���,�����?D������9nM����4X�:�yK:D��* ��J�(�cb��7;C�9�j2D�@�1��6EህB�i�%���L-D����:0_�����_KՓ��)D��d˜���@0,�"}2��j�'D��8��U�V��b�D�5l[���)/D���!�U�V#�-;�� Y0>���0D�����E�xh!.#1� �:�/1D���񏏓$P�D0�*��RGָ�6*0D��կV��q��,�����p�� D�\JFi׋]� ��%��w�\,�I2D��z.ӆ2�͚�#�:@YQH/D�8���X�`7|���h
*s�����*D��s�.�	T�$���F�\6��ƈ)D��rG�r�t�)�C�6�ڼ� ,(D��� ℐ.�@yɴ�S�\t�X��%D��x�
��"x��!��=�U��c$D��i�!J ?����pʓ�N><�� D�`�"�4jc��a�)~ul�d+>D�Xrrd�4/\r��*�	���tk)D�Ti�'�^Xp@G*��Q� ��ӄ<D�<)���R.<A��! �d:��9D���פ�k��M����ll��^<!�$X<W<μӶ�$sP�4�<!�$�9 A������}bh�8�ʚ�|!�D@��$����3dN-�SZi�!���!ܬ�x��^�XN�<��*�3Y!�䆀[�؍A�h��ND�Y��	FR!� A�b��� M�FP�3G�	
3!�� ���s(Glr*��Bh~��B4"OZ��'҉��i2*�2cz�db"ON���5&c��s�Sc�a��"OT����ג��rH�)q�Iۆ"O�	���^az�Ȓ��I��"O�`�C��+F&-��̐'
L�"O&���,Ӊ.�fi��K�]v]3�"Od��G�N
$ ����"�����T"OPT#��^�IbO�H69"�"O.QJ�.��a=-����R6���"O,�J��@*Plz�m�?*��6"O���0��F�����%O:xQa$"Ol�����"Yb��RC�N
�$X2s"O�a2�F\�SF,J-8�"O����Bˆ5I�9ӗ��<Td�"Oΐx�IW�j`Y�#ś3$�� "O}[���0��倝�Y^4y:t"O^5����U� ɹ�&�=N���"O��X�bW,� �����9�x�"OĹ��(݆-T�a��ak.T��"Oj�M�*�t:�$��k9�i�"O�!ԍ�ql�K��I*/�@Ct"O�h�gS� P�H���zl�$"O�	b�ݱ+$�y �;p��"Ot9�b�s4���)��"���Y�"OЙ0�$�{@D�7OA�tNu��"O��cg�ަ$P�ݪ��i�z���"OJg�2Qt< ���%B�����"OZ8H�	��z�(��=p�� �U"O0)x��-ԂMC��,(��"O���4,�V�1�BնJ�>���"O�1[��ߊ-лu�Y�Y�"a(D�\��j�p�hy���ԲX|�d�WK,D� ���
�v3.�ÄU:-�xT���+D�p8`���9)��2% 3W���c'�%D��!��̒S9�uۓ��*=���a�%D���M�Ov���gn�{!L'D�8#�P�ZI�����A�j��8D����fX�w����kF�<�`��F�6D�X�p��7D�ܼ�ED�Wv��C�3D��ч�P�kv(�g� 6XS�/4D�B�Η�w��Uc��(�'"3D�3���D1~��סU�+�� D1D�l�S�� eB$3�B�?��ɱ&*D���	F�.p�q �`>N�%X�'D��آN΁3@�L�i\e��#D�ĺ��6s�������ra0))e�"D�x�K߄bѺ��u��F5�#.D���`#^,;R���E�V�4�B1�ǋ(D��qu�J�~��<��ϳ{f*m��G4D��!R�&��)pLM�/��k��4D�hhU�8�z 	�Oހ˜æ�$D���葩(�4dqBA].�$U#D�1DKݣj�0y��R�dt��� D�d����Z��Zf�Ց�"D����[�oք}�A��.!
mX�&D�P�29�0
��x����'!$D�(���5z�̩O���Y���!D�� `4��|���	�Uc׀+D�,��
�5N~Z���� K *D��J��Z�(Vu@�ʎ�9���*W�'D���$(�M.���
ɿJ:�I�N'D��s�B7S�T�w�0pp�R��(D�x����JBDH��N�QK�98��'D�� �04�T�L���u�+�xY:�"O��1�
��!���3.	s�yc�"O⼉�擛.��i2�_H\TA��"OZt�4j[7b,�٥��D�Ȅ	�"O�,x�.E	�Xh!�N�s�$�r"ObѸsB_>N�䊲L$�`;c"OJtw\n�PY�Ė�f�*La'"Od}p� ��J)@��Z�N��U"OĀ�� iB=��JO��ܙP�"ODJW�o��M9fI�#b�h8�"O@<zc�l��� �� F[� +B"Od�B W�5���"@�]Y�ع�*O�M��ē[��@z���R�(	��'�^��!���tu#@�0F\��y	�';z�����<8+���嗔S��y��'y"��WO�}I���7�v��'J�����E̑��� /PD]8�'�8	KR�Ϸ4�J��!��4#@�x��'�$ufϘ�a3R@��%��iJ i�'5����d]7��I�` �o�Ă�'�N4���"2��Q��x���'3R��9�1���:s,!�'�fa��9a��D�V���6�Q�	�'�<l��^�2wй:�N��b>�	�'}��珝gyΤh���":HS�'$���棝�c8�P�jǪl�d�
�'������}�r(kC�I/8���
�'�0�`B8CT\��V�,Ǩ4	�'�ج��HP�,0��٥ye���'o�䫑J4^� �'$_-c�\��'��qZq/y������W���@�'e�|�m$E�PC��O����'s,��v�	0�F� Ǝ�1�d��',$�2&T"8\j�ce��/@W�� �'�p��%�b�Z`j��2�>0��'q�PC��YL����遵X�ݩ
�'���x+��}i�����Uo���'z <��H،2�Jd�1��H��'뢡�'Y(~����$Q!z�'R�æ���q�lY́� �,D��'ƶH0n� #����A�!t_l9i�'���k�싲}
������re��3�'���(2*J,�f�p�k	5jI9�y�U.�RBfѨm`�
7č��ybi	�%0���	_����F���y��$_��jT�;Z$�T��ŋ�y��JU��+�I-Y���H�y�΃�ƚ�J�M$;p�2MV��y"�Ǌ����օ�(s��13T
��y�l�;K�a����.���	.�y�nΡ` �Q��%e���cJ ��y�&��P�Q�˓�Z�\���(��y"�E�|�9r�nR|��������y4Tu��b�eFM��P�ٖ�y�iWKU�HV�שBH�|j�
P�y�ʎe�QB����= 0$k�ҹ�y2(�<5yfɍ�`.�Q�f��yb \%0������\h���e�0�yRd�,�0��3h�Z�	#����yFJ�S�@�uHQ��Ɋ��yb-�"7c��!��}� ��4�y�8}�(q��O	�U������y�eFsw�e�}�&@���3�y��H�e�B@����r�̜��L�y
� 4�D�$35p�QM
8Z�h�c"O*1�bT	)��pL��7��=�t"O�M��͈K�:���kWG�~�B�"OtS(`Rr<���Z<Nh�`Z�"O�e�$�MM �S.�=.��'�54��*r��a�V��F�
���M,D��ÅKL�FSq�ŉ�!��)�B8D���c�O�F�T�֢4�r!�a%D�<����~���B֊L�2�F�0D�ȺT�ݑi�񋇡W��,`n+D�����[�?,����XT�X���*D�8i4�E;�e�#��!�7D��T��r�Ri)h����Z��8D�+�Ϟ�bL�=��ᎉ(>�*��&D���T��9e}h��聪�]�6N9D���+�1���3����J��� �&D���f�Z BJ�bD��C
�U� /D��P���"�����bL�b�X<P�J*D�� t�FA�� PF�ưT�̃�j)D�pkU!Q����B�%����"D�h�5aR�U��,�V�љ&� R�<D����B`��Y�P�p��@�%D�H[�eK%��p/�޲��R�&D�L�ÎY�,1�L�p�]�X����$D�t2�'I�z.0�q��}	+�%D�tTF�88j��En6�����$D�8a�&i�5Y�F�f����#D�x9��)��SԄ�.✁ J/D�89��D�[�(��"K����U�0D�0��@�'��kf�����*wI1D�(���-��$@Ư@��J���a;D��K����2������=#W��B�3D��z(O,`ZN|����'%A1�	4D�����8Q���3fAE/H�DQ�`�7D�  g��~��l�֮�31Z��1$b;D���5�آ`ࠤ�S�A�J�6�'D� �d�۬,wЍkP�ҋ!�fqJCj1D��0WE�?�<л� �@&��W�>D�Xi@E��n���$
P����w�9T���4Ù�I�Q�c-M�90�[�"O~5I��Ϊ%��)(DK��\�н84"O���l	Q��)����YA3"OH�,���h�A�j��JP	ק�!��ƙ�:�CQ�=���*�a	5*�!��Ġqx�%����x��Ak7 
.m!�d��
�CC�ŉN5�8��H�z6!��G*%2�	��șW�d��I�:R!��� y[����@�0�4�ZsE�)E@!�DGIGd�*ah�n�ɖ��:�!�$V�y��I2��6>r�8ȱ	R0k�!�D��%t�p�Z6:��+��Ŧu�!���=c�ny��Ŝ��=Ywa F!��h���� ��&Jf9CCaƓ:�!�D޴Q1FLIEHEH�0��D95�!�F%��iX�?��	Hv�ܯ|^!�$�
i�X�X�%҇f�����_1|!�ݷkIB��Ҩ���nlcbƚh!�d̟z�x��p�
�v����o�"8h!�D�9Il��D�ԛ*�dxan%:!�	w�B&-��$X��g�qg!���]�0��G�C|�|�dHK$C{!�E
�`m�&J�h��!U�!�Z ,��'��~~��8�
I�!�Ę�T'�-��d�JSN ����$>Q!�� �k�">�r����!��S�"O
��4͂=y�@�0)� sĜ��"O ɢ0�TR]X���nQ�x��Ӧ"Op`�v
V'�@�����g&	 "O	pU(q�,{vM͂��`F"O�Ɋ�"�.Q�1JS�� �m	3"O��S��+7B���H�	�"Oʡ�u���^��v��0q.�k�"O��(�%~�h�[�"\�2m�4"O���O'KS���!�1c���"OR����9rb�JG S2��"O�M)p�Ӻ,�=Z��Y7~,>�z�"Oʜ�t����H��&>��IY"O�!K�@TkiBY�'*�+'��uS�"O�E1�(�C?bdPfhUr�ƨ	W"O���D��RA�0(\#MժĂ�"O~)k�!�	RN�jǯ�;88��C"O�ɲ�a1�d�so�#<H@"O��zDj�[�(8�gK�y�2<�"O�:._s�:��F���t��-C�"O�@p�&�SI����狵{ÚH1�"ONIq�+Y�iN�!j3'��%���1"O|�����4��t���	)�� 6"O ��A�Q�U�LQjd�^/�0"O�x���5VUX5@Wl�-' �ڇ"O,8i��OgTx6�[���j� 5D�l�7	��k�xD�/ET���'5D�����d

sÚ2T�25SĦ D� ��݇~�@�Z�M'�:Q!9D��(" �ag��D����!�#D��X��Ӊ2��f�1q���㒈'D���@��=-��	�P��\q"�&"D��� O�0i"<���۪,e4�Q��/D��Rce\>LD�C� ��bK�\k�D/D�X����1K�&г㏇��� $�,D�`���>S�Ĵ�SG�Fjh+Ɖ*D��`Pl�!R"(�P׏R�5�\9r�<D�p ��3,\J N_�=�\P�:D�d�E�_7��]B�#߂A,yP�#D���'�L@�ʤ2DK� 3g%���!D�0�@l�4���7���2m2D�L� ț5D5R�Cd/c]�Bd�>D��h#��uWH�`��żSjd,çJ=D�p��B��XYfd�$C�}���a5D��'MA�D�xp��Ǡ�o/D�$��˘�T�2-��M�fUx�:��9D�zV��_�|i�d_A�F��Sn#D�\ڃ���p0����W�5�h� 5D�0z�&�d,���!�H�~=� �Ņ D���+���Vk"n��Hb��,D����F�#8Z���L�����P@�,D���S�|s�Ȩ�n
��q�� 
o�<1֌�,
�N("vHӠ_�J�v�a�<�_L(*��]z�εI�/H\��B䉻s�0�C�ڣ;��H,lY�e�)D�d�.&���J��4�V){u�<D����.����P���-��"�9D��:4'�?�J���ָD�@��d�%D��2bg-�(��mp�r�"D������A��p��E�R`�G�%D�H��EA*Y�<iҭV�k��'*/D�̸���bƐ���iDm�׮9D�@ˣD�V���QA�L��T8�#&D���Bf�=mev�����2R:B�*#D��  �G;/x�|�a�� <��"O�y#%�,!GT���-L ��"O�<�G���WG|��v�B%(*ك1"O`��џ_Gء�a�(lr""O���s��y��KV*&��##"OTt0M
�:s������Lf��g"O*��E��r�4�hRI+�([�"O����]�9�T�t���-t�Lk�"O�I��/?F����)}.9Ȃ"OŐ��L��t��hZ�mv��Z�"O��C�#0ؐ�j�e^�L^tp��"O�ez�O&Px�����N�(U�9�"O��1�<<��Aô��Hg"O���BK��Fd�yq���b��c"OF��!M	����!q�SX�6�@"O(\;@�^%(
������LAV"O�`h�j��8Qp<p�-� ���(�"OpI��g�t"J�[�٘}�Ԙ��"Oz�zU�B�A���3W����@�(�"O����T�x�,�ؤmQ�/�&��v"O�!P���h� r#kM!(/�A�""O���`Y���
���b&���"O@!	lڗ&��9����X���"O�${�䅭/!:��d��? \C�"O���Fa�$[�Z��Z6� �#"O@(��iL8�qi����*x@I02"O<@xA摋,�V 8#��.v��X�"O��K3a
"c�|̱W��0���b"OnY����%��B�fŻK���"O\񋇏��I�4���E�i~^��A"O.����AM�����W�Ka �@"O����%փ'd����Ǯ_F2H�'"O y��S1I<�9y��غS܌�y"O���Ɓ�P*���ǡS�:ݡu"O
 r7�����Z�#8`&�Q�"O0I�
�>�\�v	Y(d�I�"Od����?��aq'��p$@��P"O������!��Hl���z�"O|x�.�!D�t�2䏘.I�DX�"O6�PC�g�԰F샾L�6��"Ot�9Ä	�:��As�M)��J�"O�u �ڵ=�F�Q##S*>A��Y�"O~Q�H���:��,T����Z"O��s뎴�����%)��S�"O�ˁ�#�p�z��[�TjZ8��"OX1��T5���eƘ.U�@�"O�}1W�-_�<��$V6yAlH��"O�ڦ������J�8���"O�S�Uq�Ր��ÏO��"O�4k�ϔ%]"l�7�V/3K�K�"O��a0�� �����¿oPL�e"O\,�E�Q�8#¼I��j�r�"O
 ��	��QV.�6Y�&"OE�7M���ّ�L�I
܁��"O�e���%�fp�0zʑ,�!���e�lX�n��)
�H�c��9%!�W�n�j��E�@"uW�Y�F�*S�!�N1lPD8�CM"]Kz)�ag��I�!�$��'R��R��I���$ �!?!�d��DT�딝v����Ə�i!!��׺.�B�KVe
�(�()˰�@�?!�ė]�1�ҩ��}u�f�� f1!�7w
.��F۳0��Aj��A�!!�R�xn��""B��,d�
�.u!�� lȀF`��fU;��Z�/�T�t"OƼ�Њ��j���\�=�>�c�"O��x��O�r����a��G�N)2�"Ob\[�@�g8��Jv��.A(��"O,Ѡ�iO/��D��"_pԤ �"O��fߡM�f1I��ϳf�)�U"Oj�	D9�~Yb�Q�NJ ���"O�q[ŝ�R�ұѶ�� jEbYj�"OD9��EΉ <.���@ā>	X�p�@<4���+�0$K�%�/YB<|;��$D�d�gJ�Z�>!�q�R�&��%M=D���I�f�a��' o`��¥<D��	P��igR`-�&�D���<D�t0%ビV�2�їhХH�&��CD>D��CG��B
69�L��2��r0�=D�l2�k� 0ä�G��r��8D�t��U�#�0�1�@�$(�$ʲb8D��j�Ǆ2WO��P���x��Q�"D�� �>q��� �_+�N�A!.D���6�H�5�c�R'e�4`:��7D�D��\>l�t� !��
�F�D�8D��K狑�IrԠ�)�!����4D���D��A��8��*q� �Zwo4D�:3�?�&� cD�<�� �c�3D�$j�O�k�H�Bw�uA���U�4D��y�o^	bZ����	�vkG�1D�L��=a�X B-�3�^! #D��*a��BcA��$	�b�;5�=D�h�5j�2$�Zi
���t�x4�C�.D�4����n��噲�M�9CRԛ�d.D�8��nS6.���1k�@2t�A�9D����S(rr
�a�fţ.�*�F2D�P�b�i󠈃e�@ ��%ô�<D���g�]7h9h*"&�Y3��;D�����!Z^d�D� m? A��8D��0#;92r�qfk� ��a��4D��S�*�/!��y�B�f���S�'����+붌�.��]��AJ�'\9�h��1��-�0�,'~�b�'6�P�7-��e�8��u�K :ʝ!�'��BC�z=��+�*OJ0{�'w�H��H�w���`���A��'dQ��j޽�B��!J�\`}��'�^��fC�9*b����OU�})�'���8�\�OxX����S~���'5�t�t�C�	H�u��-��N�ɱ�'����%VW�A�K>`M�'�<)҆�HN�}��*X�K�'�&�QPl�b�(4��/Iu-��'����цۀ?�^�Z���~���'�\��gN�xP�hg��;u�*�'��0IVH�6o�F4��M��}=>,I�'��ق�b���$��>>�K�'��v�L1�����0(�\��	�'k��� �6IѢ9�陰%����'����y >p�dEA����'(��i�@P�6�>������
����'��I�։�2qk�9B*�|s:x�'�,���eГ[ ���-Ӳu���'����U�'���8�L_2uf�@�'B-)�'�I �ؖn/C�V��
�'�F����5ph�c��X0��-k�'���"DŢi��r�O�
H���'\B��f�*��ő���#��
��� ���dH�^��H�dS5�2L "Ot@�Q#ʆq����)l<��Y�"O�I�d��{RR���I�qK�97"Of��N.8�y;�(�MHF�K�"O|q����hI+"��5\�逤"OT���D�_�-�e_�&���P"O�I���w-�L���\�l���"OLX���!J�b!�Vm�><T�p"Od=���U��Zhy2�ƀ@:��u"O��!e0����D&:�P�A"O�M�2BV�m$dp�Ȍ#Ar%"OD$�s��>t^�r��^�j�""OΕQ���Q4� ��8�R�7"OH0)4`O�77`���.�>�P�"O��tCϿHی�A�����Y�"O���cfȫN�6��%*X<	z4�R"O ��1M�7xґ87��^]Ԑ�"OԽ9dB�q!���A�AI� т"O2����J �c5�Tr�4�("Ob�!��	�~��<�E�E��p�'"Ot�f%K<�̰��!�>M�z�ۄ"O~0��$��'<\ �� ��aÎ�z�"OP����ìY,�2���'�jTy&"O)1eg�=�N)��ށ,����"O\�"�@=  B��Mۭ_����"O�)�P"�+v�xy�����j�"O�%���<d=x�kǊP}.�"�"O�2G#�� ��*�� �th�"O�s/
.9r-�_(�%�P�l�!�D��p�$��i@�Qrq���%!�dU(�
=Q�{�Ni¢�> �!�Ė(z<��5����1���U!�)[�Xْ#!=����`��?�!�$�=_��p2J^#Fth\��N�)-6!�7k2]
�ɋ#6�-�pmɣw%!��i.�)�.w"�˳ʖ��!�ש�\a�`+��w-�����x�!�D՝#Hݠ4�J$v,��q�G6-a!�dV�c/PiHБg*:�Rg.�!�45�&�jGϺ[���@,�1�!��2xe�"�L}�AqIM�z�!�E8�v��ɭGo�����62�!��i@��u�W2N	J�{�b���!��X@�&��ԏ�T�x�j�U�>�!�dI�vy�,�)�;&���QfAʱ_�!�$�5i��Y�wO�Y������ƕKO!�$��Q�b�SFE��!%�\8��E4?!�D�'H� �PU�ל�$X/	!!��ЀrABI�E�q��t��nH`�!�$N����
<�v8ӭ	�+!�D�%i��M��۰vʹ4YwG�C�!�$L.!ߠ@H��޺%-	�P�H�!�DԾذ���������'�!�D��9D���lQ�I�� i�?<�!�U/^4�G��Z҅�[X�!��8'�,��R:ޜ����j�!�DO8t͠��s(�$>sg��n!�D/.c�|���W��{bF�Q!��,����g�]8�B���$,H!��(.�;���~�����'-!�ۀ? ��@�/t��YBA��,&!��6m�
�UϚ���IS$��y�!�$A$N5��0h����`��(=�!�D��]��̈@$F%��](�K�
;�!�� ��& [EB|�#V�E���S"Oj3�LM�2?�X��%L�8�L'Oh�D�|T^�QfJ	�b��ZD�T��Py��,b�|�+kEt3�5QԦ���y$]
K��'ʻf��q�F!���yRn�&KjQ�PA����	Pb��y��/�ĉF�ԅ[W���p��8�y�?~��r��M+t>���M��y�M��%	�P�W�?:X��MY��y�aZ�b� �hq��1���0E��y�!�/, Z9�F�^�)�$1[Ѕ	�y���T	1
Y�x�!'�;�y2�I�.�>M3�)θF����fb��y��>=�p�IP�t�
F���y���Yp
8���IK�P�v)^�y�	�.�~��׊oU��z����yr)��E�\�h��C1c�Z��O,�y���8< �Aӓ�l��S`
�y2��0�0��� Xq��Q���y���%T��#����
Ӥ���y�B5��=��
P:M>xmP����y�˛���� S�BY$�(���y��	�ȵ�v�9<  `cL�*�yB�b��9�b�C�/u�jw�ԫ�y��G�}������#=Z"e��A-�y"ߵ$f���׼3��遥���y"a$GZ��͊$~N9��	̈�y�k_�N�"Sc�����7���y"�[�d�|ŚЎ�7t�f�ؖ̒��y�%�+/H"� E�v�\Y�a���yb��`�D�:/ղiZ�] ��ё�yb�8��Pw���L�)X��y��N"9�&�q���' Mb Ѝ�y�ŌBv0��$K �����ɽ�y".њJ~�zDK(b8>z��ܧ�y�)�ti$82�ǻ'Vqs7뎻�y�.��qu.I�UQ�UyL��#��yC��h-h�ٱ$��<!�ջ�y/��t�R@ucÛ�� ��&��ybKA��`D��
j�	�S ��y��N�X�
9�fB�4�Z�2��y��^�o`*��d�۽2�F����yR�I�}Si���,g�]�-Ƃ�y"(��.���z%NϢw� i���ʔ�yªJ�|~�<��Λ{�n��G۹�y2$�!�>4B�%�g�tAZFN��yBɟ�o�v�PѬF�T5�yzf�^%�yrg�r\���덊U�,r���>�yr�L$R��d>��*v�A$�yB��+��� �`&��4�~!�'�ژ�vE��(���>2ҞH�'�z5�u��t��)t
E
#��`"
�'Ў���ώb�l�(�B@*p�صz	�'��U���R ��hU!��hcd���'A\���.n��FW6Z]�}:�'w��˷�	�R� Tn��<d���';��C�`9���aVE2K�J�#�'X���@��8]�(�F������'{�8	� �(��DɁ
i28�8�'��-kV��L�䙢�g�s�'`�A��lǷ8��3��2Z�u�'���E�̩�lH����:��Ĳ
�'����HXC�H�rr��3gt�C�'�f�`��K�wwb�;�@�MR��	��� @���e��a/R�� ��!X~��u"O�,��ݝi.<0�'�/�B���"OJ������B�(���Y ��5"O.�x�N�J��(QD]����"O�mr�Ό�,��q�B��R���T"Ozܢ4��R�H�d������P"O�0��*��S@�a���G}�b2"O��Xi��F6 �B�(?ZE�]�&"O �A�A�<Uh&�E�
�8:lL�"O�i�G]�L�ܕ���B9(�9�"O�#S�$g�	�SxP�:�"O��	��C`!10���q��Ja"O&�[��ƣ)�+)\!D��"
L~�<do�"{����U"?��!�FB�<A�d�M��A{��_��%�fJ@�<I�'�R�,�b�����@�2SNS�<I$�e��d �a��ž��r�Dd�<iB׃w|��3�F?ff�Az�[�<A����YX���l��:�d]�<�@��*0p�2���xA�pB�,Xo�<����_~L�A ԣ1]�)�D��g�<92�Z�<3:��QDݟ?�ڴ��H^`�<Q��S�	�^�C��=�2����\T�<���{ 8
!	�4�RD�r��v�<��;,}���Gµ=����u�<��jA �`*4
�]�"��E�V�<�t����I��̣W��@3eM�<���� �-y��!1��u g��R�<y7�)Ad�R���xL}�CaO�<���7J�XR��@�x���ǒI�<�Gf�{l69hd��N�qr��D�<��W����R�Ĭ��)3Q�h�<I��B��{���+B���"Fd|�<1�&QH�%�@�n{��"��x�<1UCZ&�,Y�O<�:��2��z�<�)Ǣ|��Xq�G�Ctf�j�AK�<a5�G�kC���!��S��1�.r�<)�e\���yy�l�-l���U�h�<a�$�=�|�Rf�փK�bq���d�<��mJ����G�n��JeLA]�<	�L�|��� Q)h��L!���g�8���y���܂9T^�ȓC*�g
��.��J®�[�FH��uXV�I3AѣW�����?D�j!�ȓ$,��`�N~��Z֤��H
���!i\����aJ�A��ش��L�ȓz������4P0�$9�ȳ48L<�ȓCJmj���gcjpH5C^����ȓ4�b�\�#��4�)���ȓc��y�BI����0h�+�f�^���[l8Ӧ�X0Y�x���B&Eb���?��,8��
�2�4�qV�5ܢY�ȓ{,\�@C��@���i��
�Ej��ȓYe 眠38-yA%ܑO-RM��@Rf9@�oO�l��(Z]���ȓy� �BaI��O1~�+��쥄ȓ��`�@^#�PcSK�?(�t��ȓ�3�$_(g�\}�d��mc>��[$$�7J,�ܑ��H8Pp��JR�E�r������`�+!����j0	g�Z�ij<Hv�J*,|����B�~5)��.g���g�){,�	�ȓD���&(2��ѐtjΡ!��(�ȓP�ޔ�2�W8T�6�xa��! �ц�S�? �͖�l>&BP�#>��B"O�e�᥆�b�f}�%��'���"O�	�u��)-�yb���<Դi�"O��(��ж|bR�dB�G�
��"O�As֣�el~���J7m���)@"O��1�(S'L� ��$���+��!�"O���D��H�,�QU��n>�5"O�4c䩀%^z�A��0^̼�W"O��Q$OG,��!B��ZE�Tbr"O��!����T� S3E;_Л"Ob�P�1u{��Y�ڿd����A"O��C�Y�1�M�<� �!�"OD��#e^�fw(�职S%��Z&"O�5�D�
���#��1#"O�hN�:�������X(�"O(P�ݍ �a�� �2�"�@d"O��2�k�:R�ع�<j�LѶ"O�����
;z�"���i\'V�hؓe"O�u�-~��lw:�"O�}qQD2�Ν�!�\Ќ��"O�yvcW�ORp��I�^Q>%�a"O SsJ�����iD��'��E�"O>�Y�a	�"�n}p�(�0�Ձ�"O0آ$��5��Y��D2
�����"O���w�َf� ��L�t�Ɲ�b"OT@%N �}0=��	�l� m`��I�Έ�>m
��߳���3,�*Y� "Odp �,Vc�\�K�4$���"OdU)q"��s���3�Ǻ7z�Q"O�$C�^�h-�T뀁.��"O�ɂBN�u�@$1���T�@c"Oh|#6�
@�)X�(	0�J�H1"Oֹ�@��7g(��#�g�H���9%"O�l[%�+~L>Tk�- |�a(f"O�9r�ㄝ -|��҅�=ʉ� "O�A��l�8?�*�`�$�=Y tt��"O���j5XJ�9�-�z!�"O�=�"_yd]���X%�Ũ0"O��Kb�SQPM"���`��0:�"O��2�f� *D��
�*"���"O�ً���
i�ڜ�D���33����"O��k��vN�x��ȃ�R'q��"O��?G>,�7(�*O���%"O6��B��a �PWg�V��P�a"O��hb��0��7L�Ax��"O�=�1HK=30 ��Mdq��"Oޱx�k�3Y������9Q�`��"OZL� ��H
Z(�r ��;h�A"OF	��b�!�v�sD �+ V�d�"O���1e�Xq�\�%oǫ"b}��"O�iHG��(]l�S,߃J��X+�"ObD�D��Q����<�L�x�"OD!06(ٗ7�p�Z�
�L,�"O�� *�Q�$�;0,T;4Q䍰B"O��Q� ��kE�0	A Qd��3"O"a���#f��#����LiU"O�Br��
a{V�5��@Ր�`"O����"Yz��B���fo��""O �ɂ�(O��g�� S� �:S"O-��#�t�˷OV�9���(f"OhY@�ҧ
9��h#/�-�tX�v"O��R-�<�u�% �6D�!"O�0k� ^�D4�S���_�%Zd"OLh̇�w��}�#DʮK�Zչ"O� \�(�)a�GÖ�7���a�"OPy���
N��2�� =�ƥ��"Od�! Kߵj�½�r�
��i��"O
Az�
X2n1��N���`Z�"OT�i�iD�ȅ˱�RG�����"O ����_�4�mT�7��IR�"O�	K�)�"�v��ĭ]�;��P��"O�C�ς�m��{cMM�\� U�3"OT|k�a���P��k�.~�J49c"O��!��o�0���WJ�i�"O��3u6]��HN2lȊ�;r"O���s��?;vx�v��k��A�"Ol��`�$t�@�υ*�ͯ[�<Qu�ۭJ��p@��X"%�݉��x�<Q�˪!�J r��$j��@ �/s�<9�I�?h�T���E#K��S�T�<��I)(><xZ�$Y��h�E�FO�<9C�ߎg^�e���)QҬ�8"ώd�<�A���������D��AHTdEe�<��v�t����D'i�E�PU�<Q���$d�D(�
��hN�u�EP�<YS���P��)�Dټ)��	���RN�<1�`�"tA���!S<Z�u��F�<���bL�p$�� �� ����@�<q�-S�C�*�#��O�!5�F�<�-ͯ7X@�Y��*g���V��\�ȓ!c�X�`�'�2@�����rYN��ȓl3�0��P�P}:}�D��@I�ć����ȶ���8�����.mWҥ����$��M]�c�NUʆ�L� >9�ȓsh�*��V�?fl��$��] Ȇ�Jv&���R ԘY�pˇ�M����ȓfD�)b���N��1��Y�`4���1�\�r#'��}�D0�w��v��ȓG���!��h��a�/�x�h0�ȓC�6${rOƠ���qaO˖�����0�:p$�ՋD��؆�"pd���ܔUNL��`̳��ȓ��t�d�	#��A� +\$�8��褭���=o����"O&�2���p+ �3&��j1�DY�e���ȓp�q�R*C79��ea�� n̈́ȓ,;�l)D��3�Ae�W��]��D�	��d�/U�Ɉd ���,��%�9�G'�9w����s�U��<��qd�+æ��?���X�P\�,�ȓI!�q0C��&�:�gҺ#�ȓG/�Ya�A�NP�7m�8M���ȓ�6�{k�<����/��H��Z�*L8�A[HK����Ó?H�(�ȓL���c�Η9K���*G�&�8܅��z���HſK'� 2���V�ڤ��c20�ƙ٤`i�
�/!4�ц����̜Tt���a?:-�ȓ/e`� A2���H�,������ȓzq�P�`��r�0[(��I_�(�ȓ[|���Y'WX&���� �h��CS��@��44�4��W�?Xt�Q�ȓ{�$�:w�B1�hYU�o�*��ȓyZ�&FJ=Un@��'Q�(�� � 9&�аW��C�<#<��Vt��Q��$o*H�/��8lx��ȓ	� Yi�/)Y��%e�;��ȓD������ٸj��X���͐��d��S�? ɧ�(�f�ZS�ɖ&;���"O��"�(��		0õ'��!�I�"O����+�|���ږ`��!�"O�� b-Q��$�z�����0"O~Q�Q#\%�y���{���"OH�yR��.��ӕn���n���yBk;+\Dx ��p��Q�reB��y�Ɛ�|Yc�I�d��%X�`	�y��<%��Y0%dJ
�*)��$X8�ybMZ� ����W�|�� ��_9�y2�]'4���eS�w���G�'�y2�N�6�ژB���Y�<�	?�y��7�"�f�R2��l�7�I�y�w((��� ��\dK��y�w�y@"!�3}9�Ix�՟�y���8l�4��q�
�e�Y9�yRLK�u2DY`3K ����jtJ��yB�'�a�6�惡��	6C�\PROE�1�^�p�`��v�8AЂ��J1�,X�i6 aÁ��Z�k)�sj��U��\vn��0�� d8;��i���A�m¥Cs&��@"���I�A�'��d����U1Tx0Wn���4H�O��Q#�O��lZ�c���<�������N�Ókŵ�e2�oߩ	�!��˱�欳b��#��v`ѫp���شT��|r�O��_���%F������?(���!��5J�@�:�ƎJx����5l��5;�#@u:��qB?`��p3�DM�C�.M�jڧ$R�`r5.E�T&��P3�/ܡD��1�IF�I����*��4d��QF+ÀK����,��m؈�d�2Z%��\<����0�ٵwְ{�cOKNrQdm�����<�im�O���'z@��C�΁9Z�\�TK�;y�ȓQc�4�E�=x�~�1E�G����Z����ѳi)剉y-,�j^w7�����~	^,� Oi�~P��ʀ��'>rH'K>��K�MPo�R�Eߨw?�|Χ-��P��"�MՎ�EiZ"<�Dz�a`hhX�<Xg�	�g
5�擮c,)(SKF�#�˞�v#J������|���O�'>�l�%z`�!�"�5Y�bǥ۶\���������:��F$�>z���rD����I���O `lڹ�M�ش;���!c���p 醷$3> a�O�!&"���m�	Nyʟ�O��&Ĕ{�8�sgMT��V��=I2��4�J�
��ׇK"^T`xr�����7`[�s[ū
�2	�P�@�.�M��źh��!�����u���Ug�-�~�|�1+	�d�GJ@"hv޴��,v��o�,�����O:ym���<D��4t�n�A�
H�Qs|,ۢf��p<�}���?	���,��,M�����6l����=}��<)��i��6-4�����(��"ڪ��)�D��C�ax,O|�pȂЦ���&I���T�>~���d�бr�����2u�L� ��s#Uf֦�d�$g�M#�L��jTBRQ5yV^�b���m��VQ4�!4]N�4"3h�[efۜD�F#vk�$�Ji8��'l��I��'!67m�.��Y����h}��_�O#
�@�o�jFƘ1q�V��y�N
+4J��O����,WK�|l���M�K>ͧ�
(O��l.dT
�-}^PEx���D���&<OR��!!�Ea��˼q6Q�*#-�>�S/�DpC3֨��!����OPp�s1�����KB�>f1�S+ V8��A\��P�P� ܜ�G~����?���R/IIX�z1�G�a^��9B/!+߆�"D�i+�\���	iyB���/-�@�NL�H�����,�!�8��`I�A������U8?[�����i0�4�䓌?���ēL��H� @�?   X   Ĵ���	��Z��wI
)ʜ�cd�<��k٥���qe�H�4��6X8$<gT��"�ᔩ^�"u�ǣ)z�4�L��M��i�Z7-�Vx�,a�K�[����݉a8�-q��D�Q_��b�iq��a��	�"��6��Xb>:5H8:�UC��Ǯ���Q�Mx�ݴ��	+hf�(r@[�剟R1Qq�#2�HY���:K�De�R�RT�6�[�;����mbm�cΉ>�l�y�t<�FH6���Z�(8C��<k�H��<������l�����U�l�Hu�O�	I���^���Öo���AB�Oꅡ��N6xP1O��t��	��'�^4��-ԒM��1��Z���'"B�Fxb@�W�'r���O�W�Y��@�+g5�&->�9�Z"<�#G�>Q��d�>x�ÎL�^�q v�FM�d�OM،{���P��rg(Eg��W A�M+v�(aŰ#<3L6��
c%���\�Q��Z��Ȝ�>A>�y(��;J�*#e�}���)t��|��'���Ex��A�����l����kR@J�-�,|�!&�P��#<I��O�x�r��g8�̪P��9L����D���Ot��H<q�C�f�H�"�0��,x��^@?)1�8r%�O,�&B�U�M��4y��	�-J���
��IgˎL9@�$OHi�DQ�O�l���(��S��LB���(t,L�/O��9#F30b�'Vp5�� �ēB,�����u���xS�A;+]$�+��/��$GyB%�M�'�����	�`��xH�&�k��X�'R��:@ ������iC�	9�x��ٴ:z�Sϟ������KfJXYcC�ZO�qy )a˛��'j�R��|B[>	��RL�Y+���<�����o"qG�pn��U��m��4�?��?1��qV�'er��v�"��-�@zX��¥��".7���X��d/��|�'
"-�9HI�@�cD�w�DT��/�W#�6-�O��D�O�Q �j�^��埌��r?!����ۮ�8t�ǀp�A�rm�צ�&�prGN�(�ħ�?���?����6*͚���/Fa��/��
B�V�'��L�v�(�I��&�֘�Sv���N n;�L#4C�'*:N�xP]������O��$�OjʓF��a1h	8� �ŀ��j�.�ZHTj��OT��8���OV�%&{��b � �|>P���OT�rN�g3Oʓ�?���?(O��r���|J�D	    �    �  �  $"  d(  �*   Ĵ���	����Zv)Ú'll\�0R�P����=9pn\�Ёba�#������{�<I�d� �t�Z5$��vT�aN�!@ i®�,]Q�����E���I�A���0�2rTƌ�&���L�/xP�A�^�M� maf�E�m�];g�0'h{G��PZ��xv�Ӳ]m^X�S�a���N�y�D�{�e�>;P`���H�F���_<k��ac5���0$���72>���)�-#��d�O����O�e�;�?����$+H1p��Ւ;o|�ԫ[�gS�	`'&��d���A�4L��HR4rP�шw5�	�6����0'("ݑ�<J"��V.�> �ɕ��<\O����(��@*@9����3|r:�"O���$��A}�@85A�.� ���ie�"=�'��+�B(�4��f�D ��,����4R����%+���?���?�������O6���*!���S�F�j�/[�`��p��l�QЊ�0c��_�Zz���[?Q�4�U&�xUXv�վjxƁ�3�:J��X�t�M�W��Q��`�S�'��QJ��gl6�˰iE�|�2���lB�vT��t�i�07�<�I<�H���LH0Yx�P^� �C��y�&��*8�����ɠ��Ƅ����JM}2P�H��G�6��|`���L8�"nӪ(�6�\�g��t����)w�^�"�"O(���ou�J\(^�12"OJ��g�"L�x�&���{pj���"O`s��]�hZǡ�=
TZ���"O08���̹)�y(�B9M����"O~�����q>� �eI��vr4�"O0]��,�a��ə�\2X���"OX�r��4W��Ҧ��;>H��B"OB���#�m���Ah+ [�"O�H��ݎh��8�t�(�(�"O��*d���l�J�qAhU<3�b�Xv"O^ݣp���[�
�ɣ��S�"OZ��N�e���5�va�Ivl!�dV5��@��� 6�bA���<!�dK�XmD�� ��[N�,ru�ߟ !��G.u��ʷ���a�p�ˎ�*!�$Q�8�ZK�d�h���F��1"O��XD@ l�:��P0���)E"OX�Br�]�f�^���@�~ H(��"Od��o��(��smN�s"O�=2RB_�pʾ̈RΏ"QFڨ��"O(���Ǧ^T.���c��_樘`"O�\S��[�+k�D�0�B�PSt��#"O:L(Ҥ�K^d�z�g�\z��s"O@�tH�V_
�qD���9WؕpA"O�}sr���f�B�\PҍZ�"O<-��X8�$��G�8�.���"O�)#7�ғ|+Ar�%J�Y�p�"Oּ"���-��jZ�u���"O�@��eT�l���Q�)�#�=!�"OH!�d,����I�M�cp5��"O&@�Ť����9��3G�F=@�"O^���`�n`��{6 Ʒ<xn��"O���r.�/5ĩ�&6�� �S"O��4��dP w�� n����3"OD}�ag�[U��ҷ.]�(���ir"O��	3�@�0&$쓒��X7"4�"O� I��ء.��q	vlThB�1�"O����_/��#(:�i2"OB��q
ɢf��D����}nb�Pc"O�(ڇ�#e��}`Ҡؼ4Zڵ:�"O&���k.4^���PO�u{Q"OX��.s�a�T����		C�AK�<Ŋ�;����_\:�5�d�K�<�7��n��)ǊR�H�(�B��Q�<�M� bfŹu�Q�Cm�Ty���s�<�&	+!P��d�@b81��ər�<��LH�0i��js�˘4m�YjW�C�<� :�s-rXEa5e�?�f���"O `0ǆ D�����qH앰�"O  
��9����0��\JJ�J"OΠ�&i��`\�9���$i��l"P"O^�
�$� h���7�"O2��aȭ[�`Q��^/#�~�x�"O���7�3,]�̃��t�P�`�"O������8���ԯj�����"OJŚ�bL7������(@ʕ��"OLY�qf�/-���U�!8MH!32"OL�뢏ɲKg���!$S�;����V"Oz`P���'�U�7�y���"O�H�dFEm�b\�g�� k�p�"O�`` ���m��9Y4��[���11"OV�iQԒ{��`s����D8�"O$��k�v����E����q"O4035��T�r�Q�D�5HF�y�"O0���V<oE��(�˝���"O�(�s���^��Մ�=�ht(�"O�|�qm�!.��E�檐�b��t��"O��Bc[�&A�D�1�#?���"O��´m�1e*�A�'[8w�NU8p"O�]�"@D�hP^p�f��P�,E�F"O�$�֫.�2��֏-���r�"O�a������X󮆩^�.���"O:��m�w�9в�Q=+�|!C7"Ob�r$e��f�Q-�N�r�Q"O�-R�̭t-sFX�d��u
#"O4 ӣ�τC��8BP�P���"O����M�)9�Dd{>Qr"O�`� �3���fĕ2q+��@"O�%*q6�1����0�"O�Q���Km�ő��D�	0���"O�0��
ӐU�4qG.7vd��"O\��nI,2�����?�^�Ia"OL��6�ڨh��摜-�=�S"O�6��?�$��EN�	r$Ð"OxH�Ʈ��z\�kT"�4}�ܔ#�"O����a�H�ٶc�F�90"O�L ��J�h�q���?����!"O�(Yq�1Cю(r�$��h)b"Ovi�Ə˕G!f��j	��d�a�"O���I3���G�@��A�"O:bC�+/z�#F��9_��M�S"O 8:$#����QР��woB�@"O"I���իt9�,�N	&4z죒"OV�sB-E-oF�@��B'j$��37"O�Ib���c�l�3�E��w!,��"OZl����Z��	
"Κ�X�� �6"O�q�BL�~1����/H���@"O�4���H��=s0͖�d�J�0"O����	^Ď�s����.���"O(��j�I)��&�._�،s�"O�$X%�ީ:MNm���%j�~Ő�"O��V`�'XY���b�ΨH𠃃"O�ȇ�&*�XmS$�5,��"O ��P P'\Y�\�$��Xll��'� t���'SN��F�J�i��t0Љ�
��qד�u�eO�"����y���Cf�Vbb]�P�>[!�D�>GҐub�kM�(bN�3�E�_��'�N�1�M�7#��q �r@�����>�x�2���C�	8L�0������%	p��,��n�����{�
˓��D9��L��2��->�����bU9V��t!��0���d�� �z\����t���%��1�	�4��O!��I�I	~؞� ���&G�vXtqr��<\��2�'}�Hb���=@o�q�G��'b����n�zESѩ�c�X��eM6�y�A^L��iu�l5�)�K%���lXj�Q ��.
� jăٳ�(�N��݉��T�#� ,�¤�4"Of�p��̶'��8��w_���n�(G��my�F�#yP�x�]�l1�1OVMS��![1��:R曨؎$���'�VLQ��cǢ�`�
��10�C���0(�l2r$
)6/��)�T�az���&/4�3䞮Vfʉ�A�	��O,�JԈް;:Z�+#f�|���R>{ CF���9ˊh�E�Ĭqu�B�	�&�x�y�E(ҬA��!)���- TI�E
P�q@ê^��dӊ��F G8`b��J�v`F�P���!��21���;U��E"c.�.-�M#�=a,�QkOrfr�PԚ��d	 z��	:��'&���$�w�rh :v�(��M��>��	�Eݎ�@I�"|��ejd��8  �q[��'h$��e^<�AK��$�>M�Óls�آ�J�E^�!K�aC��Y[�)�.\ )�M�o����#�M�<)G�R�}��1ah >b.�y3C�M~bZ�x1G�
�2�.$�$!�'^���(vI�7� ����W�̵�ȓN��a��I�-9�J����C�Wg�H���ݐ��>����O�u��aB�=Ȍe�e�i!�`B"O$��`�1)�"� e�ҷE1hd�Ʒi�:"�F$U �P�
�9�$"r��6Y\A͜�&t̬��+a蠘�Ԍ���yrHG�k�d�����W�F]�U����y��g�ȥ{E�=قT�f�.��'�D���C�F�"~�"�=��M��	n��@�3n�B�<��KmR�a�҃@V��#�W�<Q�U�Ԟ|�GX����R4q���pÓ%�z5�3i��XT!��AՐ Vǒ�ܡ�oL)}�RY!"�a~R�@�����[�6���f�ݩ�yB�]�S�~�H��$\x&l4�y��ɡ�ʈ˰I,X|$���y���U�b����i,��q����y�,�?l�nL ����6T�@�ޠ�yPs^0�(��U ,���y��'A�I���H<B���P�ώ��y�A�X"�`�cY	z{�g�
<�y�G�"Wg\Dx��7t�"���/��y"!�4z��$�n4��9�(F�y� �h ��4 ̄l�
e�R�߻�yRϙ3��j�'ϻi�rJ��y��?3<|FiҮn>�U�P��1�y¥�4�"��6m$9�
������yr��?&��QIŢ]6crrt���T��y�&ʼzĚ<F��"��=�Pb�4�y2j�1sԱ�׺P�կ�4)
�'�@]�v��1��-��Eϖ)4����'S���hX0�L��fK-c$�:�'�l�@��f"��D�%N$ ��'p̉�O�?RLT9�U 2��yA�'�+cN (�`�t�F;0��p�
�'�v�X��=j��hC��R.5�����'J��Qю��dE2�z�L^�;��M)�'o�	��L�=rt���I�$�^(Z�'��!j�Ϸ^*(�� ,H)VE�'�VH��ݮ����q��y:����'��Q򋞷[�m2�fB�r�.3�'c(,Q��Q���;��� �n%��'�F�����f��Qz��Lʶ�k�' &Ы��8�2ё6蒣qߎI�'!�-+u,K5��Щ��Y`��0�'Pt�)���e�4���9N Ti��',&pY5��/���W@��@[r���'���'Y��6�P�l���'�I��-�"N�x�!!F����
��� j�Gܠr|���F�	1lP�Ц"O^RD	�d�UY���u
����"O��P�Ë�#JZ���ɻ-���6"O�ӳ@�\(e��"$�A�q"O�ؒ��Ƨ>_���������Q"O*�S�Z�V�P��@�1`rF��2"O��k����󬑙hvը'�;i!��	���-G�{���W��8~!�� �pP� A.�:~��8��-9`!�D'?'�$11�?q�*pk�J]�nI!�D�.hBJ��r�M0�T=;��W��!��%6���&�V�C*dbQm�3�!�E64K:u��c�8=`��#�Ȟ�!�D�=t=���6U i�N��2����.2��y��R�f|�6�O�y���dU���kX��ָ(�n�=�y� ���O�4[m&��PG�5�yF�4A*Νٕ͈�(&�� ,�y9���I�*�#O�j;�hÇ�y¦�1��a�AHԌ�Уϛ��O�Y7Kb�欙���]��HbѾi5M��m�E1�
�3
͊�X�'�Ԩ��;�)s�Ӆ*oL��'���c�Ͳ,�� ��-}(���'�z��'F�_�*<�2��%�A��'��|ZW��Z��偱CC�[pE��'o���Qň9�x�� '��'�<�
��)tz� P��ˆab	�'Rr��Ǆ�,'�+6-��J�B=��' ����.uE��8v�<<�!Q
�'�R��PkɕU+d��5K�-�~�
�'�l����R�|��e�C3J8S�'!*�c��<�B �-k�j8"	�'Z�Q��
J��VBB;n��x��'������y��d��L=O��x�'�v�q��
 GF�zv�B@P�1@�'h��s��J��N|9�������'v4�PC�n����~A�!��'?��6��u�RQ����}��Q��'�J��tj�Q���o�&���'5�xaF�5b�\(��W���X �'�xu�!��U�B9+c��!<�	�'�~�p鋑{�\$�A킎���ʓ�~� �˃2jՀ0&KR���ȓp�	��6,����E�� ��G�L��� �!i������ȓ{���.L{a#�o�P`�ȓ!G�ja	!xNk�O6j��@� �b��B�`�ڄ������=(��u��)��z'��v����)4:�0��ϑqS����=�ȓj�(uy�c�%�Tm��='P��9�f4�#�U�n>@)��\��vY�ȓoOڴҤ�<ȴ�P�
2R��ȓ$W���	�3]洼(G��]*l�ȓP�X�J�AJ��`Ո�DYFA��}�lȣ�B��j�8��Q�8����ȓ8�p{�N�>0��˕ PA�`���R�\I�%M_�/�jh;�,���}�ȓe���b��OB��mb�mSbOb`�ȓU*T�uȅ�g�Ș�2�kA\�ȓ	6� w*�$H�V�����s��8�ȓV;F��P�hRtax�Ǔ*��5�ȓ�Ve��)�M�E�P�4	�����Z���hǷB�5#ײz�<��S�? v��3�B�ɁA'�d�q"O�@�3
A)/��"!S;JI���r"O�iȆ���/R �aMΤ7���$"O:��,�(p�* F=b��H!�"OP�
pB�جx2%�T�h�.��#"O��؃�F4y^��I����&n(��b"O:��4'��*/�J'��.zp�`�"O�8������#ł+ .d�5"O|����N��i����2�Q0�"O��AN�.r�>x���>���"O�(����|�E�'�q�"O:|�b��Bu�H�1΁%�ޥ�U"O�%�#Y~z\jvL�>ڶ�JV"O"��e� W�~�T+E�@��f"OF]�VJi�U*��	,$����"O�}w���IE
���T��`t"O����<�$!I�,�q��"OD��Γ)O�tq�E�^0�i�"O�5��$��4[��:�Ē�F��PS�"O�A
�fA7�R�1wn��t�� A"O܈d�&�%�DQ�ģ�"O��:�)��L?��q` W�2E0�u"O������h)�Yp�N/l%Ta�"OjBF��+
V Bb�je�b"O2M2�ۼG�<����^0�5�"O0M���35��1�É3zp�h"O�����."0�胠Ə2@|a"O��p��߂xH�e���WRX'"O��h��D&r����u�ǯN�B4"O�d��Gɜ\��1��Kn�6�3"O0�@Dm�(r5^�*2�Rz]�%�A"O]z�N	�8�t�g�kW:pQ"OT4��Ǐ=�f ����	J���"O�= � �n��l#�b��V�t�7��h��D_����`E@!6rAb��@)ny!�䊷9�	i�C�
	�Qc#Z��!�$�5c�AZ���k����Q� i�!��5�u�"�W67�.h	ԋ�%�!�Dʪ\q�13�ᕮ��=
�
D4xG!�כY��ɉ��L���� ��;tW!�$�JP�hA�DG�~�i�R�� 0!��1cm6�"7��u}JY8M8Nr!�d�g&a"�*CRRYH�@�)�!��-��JWc��\;�)jvJ�")�!�$�)�|gI��A�y����!�$]Xn�0��_
4�vfo!�䗯,bZ�j6,�?a�F��^�T�!��V3��5�R�A����s���4D�!�C�mf( �@;���X���1OB!�ڞ`u����II6��ń�94!��ݯ�vC�⓺C1>�@�m̤1!�DE�^�J8��!��J/`u	�m�(b�!�0` *���Ė <Y(�͏�A�!��* p����P.4�,*��[z!�
�"L,hڴ��N�4"����.G!���!�� �Y4	^�IEJ��P>!�Ȫqm�:��7B��B�oݣrN!�	-� )�����]����o;!��N��x��T'*�Hp 0�K_;!���5M;n��k��ȸ��KƯ
	!�$�<��}H��&r�B��k�)\!��Š��FA�T`���e�!�^��\A� $6�蜣��O�>�!�U�.��do�7ڀA���V�DF!�� \Y� #�:d����q�N��e"Oڡ3d�æu)*�G7�
T)�"Oxp+�.�<�`�6���>��=r"O���@ Й`��]��@9]{|i�"O���۟��ժ�V-m&�!�"O�XȢ����Dr��( fܰ�&"OH��vc��C����bMF�y�E�"O�y� ���i;�=p\�{J�a�"Or� �cڣ"X������?:<c'"O����{�l�s,�F2�x�b"OV� /	� :��!���&>��L�f"Oܭ���%�u�ː:h�@e�c"Oڥ��`�1�a�#�ؘ/�H�"O���,q��y����%ea���"O.4�#UrK|� �J ����%"O���3h��VP��h��V�n���!�"O|)1�\���|�ӫD�?���"O�`�b�q���f�V�:E �""O�]��E�(Q�Tj���%`h�"O����!y�`�+|�r"O�dCq ц?K:�J�$>��lQ�"O�R�-ƖK\����t�,)$*O<h1��\�j�:DE��ex"�{	�'�{�lO"	� �#�a���'��٩�G!6ot��A2�5��'�r]� O�A�x�1�9 �'���Kһ*Jhad�Y�\>X�*�'��b`��L��=Hs%]�%�V4��'��x"�]�%�
ăR�%r*�-;�'�p#��2W��� RLg.���
�'��gN	"~|1a�׭Yr.(��'�􌩥 ў4���(S'T6���'10X`�C�	��񪶤֜S�B�K�'jڴIF��
WE����AB!%�X��'���$ڂ��Y�H�z1��'��}���M  rf]r'�JE�^-��' N�� �4lL��0&*/-,���'���L�]qDh;�͐�\��'�T��,�<rЗ��-*�����'zH  !t86����&K�!��'��qЅ4$���I7E4�i�'^��i�bK�&H J�Ϙ	Qh,�'+�I˅m��1O��
r��; 2n�P�'�ҽsTf����ؒٹI�� S
�'���`E�!�l��/ےB+
�'��F���a Pc�4w2��	�'Ӥ��@������GO��].���'	,�:�`CH�� � 
��0dq�'؍ʡ+�6"�&�PCn�,q�EQ�'[�-20�\�6C~A�E
l���q�'6,���@2�AQʖ2�|���'���#/��f�R'�b���+�'��zbIˇ2�f��E�D�]�ԋ�'<��Y�A��C%��$7lT��'�����\�j[�U�TB�2@��'��)(���2�����E�}�0} �'�P�����'�0Q1ġ�.L�C
�'}.�����#���S�öP����	�'���+djL�s(9���������'L*ܙs�_s�b��e��2!��' � �1�@O�!qAOJ�
���'8�=�0"џ_���"b@�O�JB�M@�Q�F-�>͠gC�t� B�I�S�8)Z��5�]��,csZC�)� ~�8gM�1ڂ+�Ɗ�7��PCD"O���e��UFQ`��Md�2"O\hg	O�>�(=p�f��	��Yt"ON�cB��[sl���D��9��)K�"O�2��S!|��
D%�����"Or��bE.V�(s��ʿ�eX�"O�āRD�	"� ���t\^!�"OD�[���'$���E�;=����"OB a�R�� d�<���_�yB�B3F�x�Y3�\�&O�u ��y2�M���U���53���*��y"BD�6����Zﲥ)�ʪ�y'�)H��2���L�F%�y�`ܹn6�dqr��G�H�����:�y"�!�AzS �II���5Ɉ�y����F�h�@"m�E:�)��yIΉ�Fy�`a�-�� �C���yb$�7d���)-{P����Ђ�y�o
�u����$�A�i;��`�cy��Ec����bۊ ~ ۶m]'J���ȓ(�r$U�^- T��Ц&U���ȓj&���b"V�|��H J��d��q�ȓYEqЅ��=4�{�B�ì@���DC��޽|x(i���\j@	��[��X� @�?   X   Ĵ���	��Z��wI�*ʜ�cd�<��k٥���qe�H�4m��_;:<u�i��6���K��=�3g��2�R�9AfN/>��m���M���i�����P�O̚�+������ch�i �o	��M����O���4]�B|S&j��.zU�VnR�q_0��'&Z�Q�����݁-O�p6*�p�6h .O�)�e�Α�Zm���
9HfE��$$�4��4M��!���OZ��E�&�s��i��L�6䨰*�3�R4��GT�+��1�nC�
��ɯAhl��j�th�'�����)�~�f3{��T�u�0Pd����k��~�O�PC��J�yb���GBxx�<ID��%��l¤ �P`���<�%� '��"<���E���˖�f��-�!�U�{P�LɅ�I�)F�ɊE�:�q02�*��En@: ш�'���Gx2j�Hܓs�A��&�.+��{v��4B܁oZ��0���8F�޽�(�(W�б��	+2��%�	�L���f���cq��-Y(ȑz���5��d"q"�<�@
*k�⟬
SB�#y���ї-vhV5�6�0��ܠ��	���k�7<a��n��#�|<K��ܘ'|�Dx��Cp��:-"I�����y�j�'�Hm�f��"u���YT�xB"��P��g))��9�'��L�Y'�O�h�'�NxD�̜P��'���fDM����ݾ_Y2���&ͨJU��3c�$��ę:R �Q��D��j`ԭ�M<�����8�L�q��:�p����J}bh�s�'��Ex��a���0�zpH�Wo���y�@4. d  ��D���<��С�'��(=+��:D�X��F!��,��(ə�DJ*7D�İ�����²BSw�LЇ#D�쓱C���^'!WCF��$� D��P DP9�=�ԅm���s��?D�0�4�,m��S�Nl�~���;D����\,Z��:�=(v����:D�,q嫏	m�� aMF!�r��-D�0�R#�cv u�b��8rԂ���)'D�p�J��e� %*�-�5C�D����%lO���AmB� �T��[�6�ˢ�-D�t�d� D@6��D�e�8EO D�x�@D6r��!�i�<P�Q��#�O������$�&��3����ik�	�ȓ(T�{�jB����tj�-�^��H���B��l0� 0Ɓ�+��u��S�? ����NQ�:q�=�&"C�J��Aq��'����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   b
  V  �  p   �(  �1  �7   >  zD  �J  �P  YW  �]  �c  'j  jp  �v  �|  ƃ   `� u�	����Zv)C�'ll\�0"Ez+⟈mڛX<�	%6��D������&�:)�����B�<5�eO�N`���.��-f�A!)ߓzY��;0ʈS�'"�Ÿ�'x�zikR�1툘��&L�`=�̘c�7<򬃂*�a^4j!��cx������������3R!�0��D�꼑�n��
,�BO�4�����%R7�S��
�ٴFw�(����?���?1�jT6�ZHU1y�*����rn��?��E.-;�Z���ɰL�d�S�P���%��@��K�i�x�مώ�$���Iٟ��	ޟ��Iݟ���k���n��͓thhY�b�1�!��0O�D%����<D"�l�b �T�l\�ڷ
S}��ID?AU�[�K��Bov	��
/+�u��#�&]j�H��ן��	�,�������O��N�4c�F��5�.'�p0����>"�u�f�o�8�M�Ӳie҇u��m��M��iyA��Ol�@#7F�:x�=�G͋�c��"=ɤ炧�����C`قM������H���{#@W�=���T�L�|xh��!~Ӵ�n��M�'�R�&�-'<�"���u2h�(PA"�l!��n�j-8��Q��卂�HQ��KF�H
 ݴ-��fr�(�ّ@��{��8R�C�;�D%��T8����`�lZ�M�c�i
�����ć\x��y"�%*���@ Jém�f	����r�qa枽a(���ǢY�Dq@�wӜ�oZ��M��ᒬ &�<@���B�=(g�׶ �,����
BA��d�A�>a�6�i��d����h����"��LE�d��'�OXօE�_�MqC�4�����b�OX㟜�	�d�D�M�ΟTA0(V�Du�9j�N�2i.��I��'�__�� ���;.69"S���c��
�@Q�s � �U���'<�C����7�!2rGV6!��1r�7=��]I0�Ӵ-�U�@ME �|4Z��0�����P���E>����'�˓p�	O�5T��u
S
A� V}�	ݟ�Ib�Ş�y�剚vzj�&�>z숐�ƈ���?�c�i��i��D�R��q��xBLapw��D�$Pj�D�����oAD�*�j_�n�0 �cڱ�yRKɉe�n�
!�D�h	`a�	��y��έA�PY{����g�La[u!�(�y�,�d�h"�L�ZT`xQr���y"lE�5eJՓ�$MX�ey�)_�y�#�}��(v��H�4p���?!��w������c�H\9I�r!�'oxF��4a;D���`N���aT�
����9D�(�A�-l�|u�6D��l�����8D��i@lӭƅT�r���bV��nRC�IE��HQ��<������`��"O�]�'Ƃ8��!�p�X�pX�Z�]�,Aqc<�O��T��:i���Y�F�6 zq`�"O���nT8|���IF�;X0����"O$�*P�H>9��% 6�0&5�XPa"O�8�`[�[<^���!��p7"ON��QbɲS��DH��	0��S�'��i��dy�>�J�9�H�h�[��G�0 ����UyR�'��'G�#F��F���S�	0�7mDw���$��#�B��ь�?[����DG;�rԸ'Qs�i#f�h�f}0ԋ��/n*P���ϒ���w��y�Q���f�OD(m�+�M3��$�x��	�h����3ǖ�q&l��,O��+�)�'E�ha�P�M����J�>�"q��ɘ�?Y��*�h�%�^���s��⟼%��s�j�b>���[��ƭq�`h�nα`�;�H�w�<��aȊ�6y*��רT��C�a�|�<��I�/s�(�a	��DMz7�t�<A���#?t���R�\�f�!��n�<���&sJju4K�*��Y93�d�<���W"�:*�p��ͫR��Lm�Y�	lM��ܟH�	ßT�'`��
f��"x�b�ѳ�Y8�L\��4Vy.)�T�j��	�!�9'�ʧ�R�yR�G?S��0cV'׶G-��s ��Oe�T֪F�U ��z�ğ='����Ćҥ0Rh��P�ѤMNUk���t�;Z:P�ش	��	�Z���?��O��d�O��X2��S��!VB�%;�t��*<O���?�!A�%q��<҇	�4D����Iy�|Ӟ�mZh�i>��Sfy�MB�/��b	Y���%8th �Lt��Bl�"�$�O��D�<�L~RW'�$����4H�C ����-'OL���)�}��0�$̱�0=yV�U�.mzt3��X�^V�����µp�0���D�.3PD����Uf���`"��<�(Y"p��Q<�aאh�$���͖'�R�'7��'��?�I@Ç�)��蹕��'F}jْc>D�lI�O�{XHK�f^�;��x�K=�����9�	^y�/�7��O^�d�"G�v	���ϬF��9��)̚A���d�O�sM�O��dp>�H�O�c�� $t)p�.I�vOA.+�D���'��0*���
c82)Z''��r�0���Vax��Ѻ�?A�|�bQI/D�k&�J�ufF���B��y��ߥ{����kiy�y2���?��'��%nA�a�Y����8��r�6�Đ.X1(�o��\��x�D`��#��F�;$��@ ̯=n��qA����'D@�P`��@�b/�%��T>��O=�x���Jm���]��q��O����!B$����-�;/�t�}�@�A>^����Q���a��a�A~2��?��i�$"}��'}�Jd��*"p�A�n�0�Xk�'	8ۅ�^����a8BV�����E�O��ܡWM��H�0)R憼q��Ƀ�i���'`�Ϣ(I�M���'�R�'9#��
D�$�
�G���"!�ˎ=�ĩ�V�0�ɐX$�Z�	�G�� PV̝`��ăZ�� �!O�DH$ݐ�O�K�	 %1�1O�D�˝=X��	����0���'��7��O����O(b>˓�?i��.X����-�yT%K&��<��'�O�����G{��n��6����0�� lZ��M�M>as�O'�2.O��c���U�*Lp�C]%-<�x5d�6%�m�r�O��D�O���ʺ����?�O�J���->Wk(�jk�(@sDϋ-O�\xrt�L�Պ��%�'���+��H��2�3t��<jG��!D��XV��^ w�i��'_P�(#g�IK(9�1���Xˠ؉���?Q�i��6M6��!��OHa��K��:H!�M�;�M�
�'{,�mG-_ͺ�Ѳ�6��YSO>)[��'@��0
t����p��!Ĥq�|�T�+�"���}y��'Y�'��͡��ѱ~������!|/�6M��v_Xh�ڲeffK??M��𤈹5�N�0!��0=8I �i�����V����8�.�a����Q�H%�Q��h���Op�D)?A� ̜/Sب{Z�������oN�,�	ܟ���M�S�O��\c���z��E逎�t���'	�&#2:%�م��,30!���?�)OT��d��Ħ1&?��O�� ܱ!���P̍�E�qPr��;��'�z$ȷ�5��,�A�P������4\���"A㛑��hB���Y��
|�G�/|���e	g]h�2�1�+� Mz��X!,?��
c��1���A[~X�	���D��'��MK��O$JR�
�b�L�z�"OV����F�Q��H6I�l�Z��S�	��h�܍�#��)m�y��j�˄����>�)O��� ��d���O��d�<��0I��s�[�L�r��.\ `	�,�Gʓ# h��Θ5'�=
�����Z�>\*`��(� L
Aթv�-����>6x�6-D,�K��1�~U�=�<��"��`6�`�#U�Nh`��	F~Z�
���?I��D#Қ�b���^F0ԁ���=ThC�I���p2nC 0j%�"ď���r�����D��1�#H1w��|�E��;�
=�#��O��d�O8���<�|"􁃥r� ��o� ͫ� �
�jP�g�*g-&���˟�Jf�72O��E��9�~0Õ��1��F	c�0�ĔBY�����3���&�O��"J��be �D�xa0Yb!�D/52�'{ў�Ex"�^HPApf$E"!�Ba�G���yB-�EfT�E�7�2�pMS��H{�IU��~(�H�'�  %��1W`	�([�[I|x��V!~��p‴r�����.
 $�ȓmg���u :d�])�j�N�X�ȓG�R��F�<	$<	��#@���|��䨰��@l�(�f�T�;�U�ȓD�"�󔣎�tJ��>?
�F{��N���.d[cޣ���f"Y#���G"O��SÆ3T!R� ���J�0��"O����ze< {�[A�ݡ"O������B��7g�&
@E��"O `C��0-��%M���Y�"O�8�F M�O������6��A�1�'�,�����e�j`I���*������7x�A��)��9���!36���0Eg� �ȓR$��S�ױGM�8Xf�ݗ!鴀��w�r$e�
���*[��#�1D�x3�.٢M�N�����~�Xp�f/*D�(�c��43��X��ܣ>���Ǧ<၌u8�|ٲʂE��Л�jZ�=MXe�Э$D�� vQ 'D�!	�SE�!T�6uH@"O`��D,�m����æf�̕�$"O����%l@~͛�'�%+��I�s"OY1��H�dT�iܴC
���2�'�Li�'C  �fZ)ޮ})4�!{Jޔ@�'aJ(���߾r�B=�C�YRl��'Z�E���� �T4���4@x<��'[�]�d�ɚY����d��7����'����	� $�W�/�49)�'�,)�n~���u��4$�x�B���
�R�Q?
c����\Seь`,��+pD3D�hB���8y�h�*r��v�^���/2D�0��&��\=L��JK>p2j ���,D�K���*^�-`�`��e�P��6D�c1΂z�j�j����O��ᓓ�5D�$C@�e\�x!g ���xC��O��1�)�{P�H	�j)�j����֡c�M�'�t�a�`�1)�d�p��'�ڹD��\g�L@Pf����{�'� �R��|ļS���=`���
�'��y��$S�5��%�qi�=̼��	�'���cr�E��H�aѶE�Ze)O�i��'���X�����-�pd@�'����.������P3 �&]��'|=�(R����7#��{����
�'ʲH(�Ėf���󠙆x���'q�L��K5R�	�c�w9�� ��z� Vi ��wtRUQ�ؠUo���f{�;�؍A���Ҥta� �ȓkΚL���Z+&�2)�v�C7p�D�ȓ8���ٷ��1_J9�h�G�Ԩ��;�&ԩ�b5K�X�Ȗ��5P����5�\�ߤ��b�^�/7D	G{ң҃��� ģ��+l�Z�$[�t���"O|Db�L�i�:�0V��
s�M	�"O�e����
�J��F�*�( �"OXX���ʘ%���T��� ���"O����( ^���c�aN �f�;"O0\#�cܨ� ���@� m���i��'�8p1����x䶜3��]a~a�Ȑ�7�H��;5�Q�G����yvE�. �ȓY2�Q0���/��8�W9LE�� ���q�+
�MiC)W����ȓ6�����!�N��@�hh(�ȓq$d��ؿI�]��M�_Q$�' ؀��G�I��#1�,,�Kȉ��ȓB(8�C �"X��Ò�
�,b�͆�(�z�RBē$b�C�
�o�m��	���xr��>f�h ��!["iK��ȓ}�Xi!���xvH�e5 ��%��Ɋ_r�I6D��
�ki�̲&f]+V VB�I6Dj������gۘ��Ӊ
A�BB��?p�i9�!Ю/V�Yq�P'&phB�	�5��j��X6����&B[0B�	62)6�I�K��"i�ͅ'P^�C䉬t|~"��޾y,�0� Ǆ{��=����`�O�PPjǋ�_�����/��
� ��'=�P�eڰB�w�]�~�^���'xR�LX�zME ����z\�(9�'���Y� �-S>@Y⯖�ue�И�'}�a��m;j,MY�Nހi��<j�'d�i���pn�y�k��r�Ѫ�9��Fx���ъRX�uh��\8��a�i�{s�B�I�9r��+p�
!�����(W��*B�)� x����B�e%l4��R����"O"Ā�e�k�j�X$.޹($"O�x3TAX?A�*V\$������W�<釮�0 �>zuD�7'S�����Oy�
��p>q�"�Nu\D�����ܭ�b�N�<���  �c �k����F%�J�<�%��>b��×�@=}�:��'�M�<�� YgK"y33�ӯV�n��1jOs�<ك`�R�԰gj�*z�`�'RCx��i�ୟ���ן[��u��j��&���V/!D�����Y�
�:$�6�W�A9��!E�<D�4����7W�.����z�V�b6D��@�it����ӪAuL�@�5D���I[�}�`���V���c��1D��(�bޚn��)(�ᐲZ��ut $�o��UG�t	y��!�q�ҿF`��C ��7�y�B"[����肱C���
�V��yK�C���m�4-䘠$E"�y�.�zg�Y���0#Ą�d��*�y2.�$]�`h�A��y�FӀ�y�	�7 ���ĕ������?���PF���� 0�t!��@���b�5�z2g�,D�l�A@��"�܀��m\;~j���-D�X�D�_��]�t�Ͽxx�E)D��ZTCQ:ITz,Z@ɏL0����*D��D�m�Ҝ�-&	�(��E4D�@`�(N>s]P�b�ˆ�la��<��e�K8�̉�f�,P�Jݛ���{�IA�'D� ���Q/{fH�S�τ�$�T5IӠ$D��	T�q�l�R��U�R9�Vn!D���G��MA`�m���ب)�i:D��!��'e�PqaE�P:Oi����6�O�V�O�	&�� ��P�C�H�<o����"O1VBD*:;���#�C�5��Ȑ"O>5�ƏZ�2Wd����^	~-�x:"OJ���h�:���B�Nŵh�90�"O���#g�~���#mݧI�K�"OF b��Q�*���ˀ�d�x����8n&�~"$([&�H��@\�*X�!��F�< �4���r����\��{�<Y�
0c�@��	�4����2ɐN�<�p�V#3��I�l�iT��AcXK�<a�H�_H�� 2BV�fJ�s&�V|�<�t��H�*�h2�ED$u�š��|sE-�S�O �9�7c��z�&�T�J1��U2�"O~�D�ؽZ����Ui���"�"OL�B���L�|��tJ�a{0��"O�l���4Du�o��hb~�h�"O�k&�ST��йRd��1�*�	�"O�4��$D�( &(�WEѵu>ư�]�|cW�!�O�9����3����	
s2͑�"O�\��K�~��qvC>/�P!+e"O�L��'NBw�� +o���"O^hy!@P)9�i3�F+7/�xw"O�;�!�]&��r�^�"��A�c�'x �9�'H�� �Ų8�"��wL��40\�"
�'bT�)��&�#���3̈!�	�'�V)Qt"B�����M��Y�(��'�L�f�LW^-�C�M@�J�'{�t"IܺA1V|�&�}�}�'�f9�'!�78�PC��v��ē����&1Q?ݠ���4�q��`I�%�d�4#D���7�޳$��(����-"13`F;D��Ё��!L�Z�ɉ�~�=�;D�� �$��tm������-t�m��"O����&T0^�d	�FC��n�	�"O*%�F+X��H�ao�U��	pT�'��Iy�����ȳ� �Q�-���=Q�h��ȓK��!� ��>"5:l�6X2�)��[��Y[�^�G��й��]�م�L�� i˸gJ\)5�ִb�r��ȓu0��F�}HP�Q�ߧY�bi�ȓjW��ҵ�hc�K�)�"?�:d�'�^p��'�,ax�CW*`� Вp��!M8Q��n���0v�D*�}�D��n�D�ȓ:��`C�Eѐ ܅�5a�Kl���ȓ�ze�Gџ2��� ��3_bX�ȓ#�ؕ �Mw�FEA!��y��q��IGv�	�x��i�jÜX�R�Z��P�"�B�I�z_�9i��L�
-���o�:d�B䉮z���x5�� _�����JS�B�	�3�` j�$Oڶ��D�ř@T�C�	A[�l���xr�Ax�m�O'�C䉞h#h�a2	�s�đ�O'|.��=�Q�w�O�������V������0^�N�C�'�ReڕjI�8@7��W�^ur�' �����I�.���d��?~n�P�'����c��84���I�c�>0-t�c�'�h�ل�J�9גu��dV�"bA	�'H�m� �kL��#%��� �S��pGx��)K->��,���ޕIE�� �W�C䉅��t�pj�H42k�63~C�	9�6�� N_�b�4L��C�7	�B�'���" (@�_��"��[�y�B�	�s"fM`���(�-���ڋuTxB�I�{F�
��:=5��rScձ{����_�DUyrOF�c��]�/]N�(c�C��Fe�<%�˓�?q���?i�F
'BX�"���UY~�h@�i��i�.\px�e�`c���Ꚃz���h���57On43�� �J��n��=Jp���Jk��8������g�CV�'��P����?�����6k��x��U!-�:�ӦCԉ��$.�O(�Q�I*���sE�h4��k��'�@ʓ{�F�;�����_�`�Nh�'�0	���x�D�<y/�X�d�O aYOS�$b=I�+ڒ) �Z#��Ou2a���|�h���k�l��O�E�79"D`�%Q����'dp��c�O�Q?R���&�2i�F�ƈ�(�صQ�e Dx��MJ�'��A�E6O\�@�'�Ҝ�����|�:��M�'}�l�SF@>.��ȓ,L�m��.X)���b�� ^<�PG{��4�'M,	x�e�	x4�$Gܔ5y\�Z���D��,��d�O��d�OV�S2s�%�����
���
6hʹ\�hٴH�(L�F�;b�F��͟���s�їm/��@F
2Zx�yA��$	���lZ�9���8�Gϔ�e�Os�U�=G��8�� ��E`n��%�g~bK�'�?����hOX�I=c��`W!]�V`k5��3=�BC�əR�"aʵ�F�"�d��S����'n�"=ͧ�?�*O��V��m<�[�����bܢ�ʜX����O��$�O��Şs2��3$L�8/x����(6���� ^������*\�-��iJaxZ�`h2!o�5<��S��H*D�:�MX&����Á��E�\{�4�^�F}�����?��M\�u6���L=$v�u@E�A��?���d#�m1~�t$W�3vv��iZ w>�E��&����b��5A�1�ɉ�}O<e�'�*7��O�|��)WY?��I�|Z���!(f�s�㊙bPȠ�4^���;�m����	⟔�bAA&�&)B���R<����|�%#o�q0n��`D�L�'���"@�9@�M�х�	{��-�������	����"X^">�������^�'��S���3}��ik�$�)r�L�'�a~2jЖ��	ĩ��]�i�5�_���>I�^�`�j�b����J���\�*Cb:?1dL]����x�OL8c��'��(@�:b�y�uB�+�8u�dLZ<Q�"GV,gNJp�3L_�i�fuZ���O�k�'.�p�B�~y�� BlB1~& �E�Ēt�䶀:#A����UasjZ4�0,(�� �'�z-y4O�IӁ�'����`�S�? >�CĆ.}�$Ղ"��0�"O"�
7��W������m�N�����ȟl��ǁ���5R�:��bG�
��t��~�����p���OD���O��)�O,H���M�[)����ƈ�D`F��٬���I�-^�8�	@P�g�'
�e�K6#�TMk��8:�h`�f�����)����匔���I&6un
��?D�d���M�^���}��I�	�G{�?O"��%��{��Պ�J@8r�!1�"O6L 6�;:���T��p�\M���'l$"=ͧ�?�-OF���R��ظ��TyT8�`o�N��� ��T2$�����O����n�d�O瓕y�x��,��H�h���?:�(�I�M�jƐ�P��k�Fe��ɉ!,�S"��aY�Y;�-G�DL��(	�in��GA.ݮ����hn��Ч#���j�f
$$b�ݚ�%�%J:��.ړ��O��kzn��"C��)�(0c�"OH��B�èk���Ӂ�L�0d�0b�S��Xش�?�+O���t��B��'�鏹��1i�
�:BF���45��F���'�R�G"9�`m[���q#�XAFi�O�)Φ��e�#�"Q:|���Kz��̠���2{�"tWlN�88�O�2(��&Ǜ]��%�����n�����d��R�s��)$?M�lD�'��Z���V����RK�<���0>Icn�o�^|j��ƻr�����Z@x�\(,OT��g��9�hD���"J��A�uX��	��Mc���O{����TM^�o�̤`Wc��X�����d-O�=���%���I�`� ��*]���?��4��>;�c>�)�Z9YP)��g�,BUQ�a;?Y4�OPQY2�>��y�-M�ն5ȷ�@�S���C7@&�>�����(�K����� }��!�)P&$d&�"�uڌ�2��E�
a�M���'�>��K����7S3�R�d�2Ǒ�I�~�'y��'��I8K�\a��r#W��v�� U�I���Bg�'�IO�4���0��
Kd�!q*�>���Cs囉��8����`�OR��OZ�j�>�i.��Z�E�	;���^/���/OT��B�>!��S/{�J\��%��1�|��$�-�~�����|�+KL��'$��Ґ+����C*\8.NĹX���	Y��)v�t���`�D铀spz\��)N,+��1g�ځ{i���G��~���9���?�	6����|"iq�nֱyp*TE"*l���R���?i�*K�R#���R膆\),�9WO�N�<�t��a!�l� ��*T*��-	Ǧ͕'_r�'Hb���'OZc��db�$i�̸�8: ��O6��O����O���<%>)C�Bܰp����xR|���!�d/�S�'x~�x�Wሶ!��ڧ� Cp�e�ȓj��̓���$��oDjcd�ȓ3dHq���M��DH�KT 1�<H�ȓxr,	����)���!��[2:M�ȓ[FZ�Tkܿ�y�E�GKO���xf�����'�V���Ъ|����ȓI�����.� N�\��Ɋ*�t���������CȦ鸲��'R4�M�ȓJ�i(�n�K����#��%\����/	tejFヮ{S�x�JͪI���'J��ccP~Rs�U�w�����n��16i��j��������Er@�?ٖhB�*ڊ9��Ӊ�~��jY�g��Hb,��2��U2�]Rʄ�4hY/���B^ I{��$O=@��U�M���sw�PK:db�oV����S:}���Q�L�5L(�@��h>��<�f���l)#D����Q�n�?T�lLX�*��~Nx��"�|�D��}^��C���p�D%���Ԕ�y2�X%(*�9��׵j,P���ǳ�yҢ��S�4(@T&r�@��ta�8�yb�'?S#��d�"t��kO��y�E��p�)a��`�L��ʐ�y�*?NN�B�F�-`��,�d��)�yR+_�AXY��G�%Eמ���� ��y"��!0����D��ʑhL��yr��?���e��7���K!!�:�y�Q�]�|q�_�2>.]JdH���y�n�>/{��òdٛ$}D��Ӌ� �yr$A�i���!cIKR,Q�􀖴�y��I4c$ti�_�C��S턯�y
� �ف�]+L��2ԦEÜ���"Oڐj��YK�)���7;���A"O�՛��cZh$KŃ�o���P#"O��x����;D�����& �>�ء"O̍ف�A��`Y�ǰQ��T"OZ$d`05fT�A)h֔dc�"O�����lq^10��ԓkHQ��"O�,��A�e�e{��2[OшU"O���E%�(@��ߜ`aPa�"O�Q$��<l��1@�A��a	D"Omc��Բ/��a0È)2Th"O�h 	�^ X��#��K��Q�"O��:�l�2Y���]��I�c"O�8���E��V�A�|�H�(p"O(T�P��26 ���!Wr�>d��"O��3�	
}�� �'�Z�
~��6"O��`GJf���X�IN�~��J�"O����E�IG~%�b�<|ňUj�"OjD��E�
6��[0%y��H)u"O^�p�B %b݂���$X0f4ڶ"O��fi��s$��x����رu"OCa-�b��Eͅ7����U"Of9)��[��
`�P���W��x�"Oj�r���8ceF��'@y���#`"O���W"�J�|��d�S�D�KF"Ov�0�'�n� %C�07�`��"Or����W.���ⅱt>�"Oh��R��?uf�l�P��$<���F"O橊e޾�&-sq�
����"O��x0��N��H����K�yD"O�U�e���T����&;��,�a"OF��j�$]D����Ι-�&��`"O�യ��a�
�r�]!_���#"Oj�
W�:6��,��l<u�4ibw"O�2�*Q�K��{zq�c"O�xZCN�O��%�'���#~B5;�"O�"BM�}��D��f�2Jv�!"O ��޻Aj P�rF�&	n ��t"O݈�0��Qk�+�&tk�I��"O�!
E�O��,R7wDA�"O�}3�b]�(�����Ý�}E*ѹ�"O��H���g
��b �6l\K1"O��:�f�clY�$
^�k���'"O���c-_�Z�� �h
����"O|�Gg�<SFuZ��%o46���"O�xiA�@-@5C��],V�j�"O@d�)O�A@2� Չ9&)�"O��f�V���Xc��7)�$�*t"O\����_9VV�Ԏ_�3��"O���	���P� �g��:�"O$Y �A�a�T�p��$����"OB�����#L�G��2~j�p��"O>	j�����i�ë٘f��av"O���v�%?���jv��</d|�+�"O\�iU�5B���"#��xJ�"O�l���1HMջR� l,�}"O���4-�2��V Z;q��;�"O���"���}#0��;G��ّ"OȰ`ਏ&SV�I4n���x�!�"O��bF��1�D��3�)j�P@ R"ON�v��9*r:q�$��,l��P@"O֕:�JEr�����	]�x��Q۳"O�A��9S��q�I�<�^�z�"O�\����)m������S�.���f"O� ��ĭʩ
F�x��HF�Z�:!p�"O&��Ț|'TP0fB��nb����"Oj|1ai����sϕ�@Y���"O���B#���b'(۸f�)�B"O�TІd�B"@�е`'H�<�"O��@`U�O�D�f���U��# "O<e��/���
b-ƿ|���"O���H	b��yRk��y҂�9"Oh]@�ʟ�6���iF�A�a'j	��"OphДm�el,�P&o�}N5��"O����.�*dU	���7���"OV�J�fԽ2[4=��iU'o�����"OX��-D���Ũ8Q���c"O����Ɯ&l���` (�q*�"OX�[4�˷2	E匪
�0݂�"Od��wR�y)�;��5'^t J�"Onܻ�.�&#��ũgEX�GFX���"O�)B7I�Y��%Ǒi;\��w"OZ%q���<�1QD�>����Q"O.�e�Нm'Ɯ-Ԁ<YQ�7�!��;)x��eǝ(c-�����ŉ�!�d�8�����;^%�A�e)I�!��]�-����EMV0[dŻU0�!��>'�f}`��@/S	��ub�@�!��4ۢ�q�&ґj֖M�B�J�!��3�
i�s��(�ze��Īd�!�d��\:��3�έ@�ꙩ7K�i�!�Ě�@z��a ᐥ\d�DÆ�˝f�!�D�\z���59g���@"^�h�!�����
�k@,��1�Z�	�!�dFB�ʤ ���'��;so!��a`1�#$Dbji��@�`�!��
<�y+�5�~ԋSb� �!�d@QX��*0.[�v�)�׍~�!�?x�����W� y�å�~�!�!�ly�J�7�H0�iFK!�$ҧaj���f��:��h!��~<!��hֶ �! ��7�=�-T1!��¹sۤ0%'�?.l��MI9Tz!�$@�>�ܠ����/qX &��l!�$F1|wZ8�6m5q:�aR���jV!��.���b4�G�$d<����+!��[<,��0@
�e�:����2!�D��"�B�it �O�Hr��4}!�ǧbv֡"D��$W~И�,� i!�a�2��a�6A���X+I+^2!�'d�BĚqQ�8NѰg�ʓ�!���C�@I�b��)&J�C0H|�!�dE((�c�����BT�%s]!�DȒŮ�@�G�n�� Rm��&�!�D���I�1G^*]�8L�`f!�$�?8�0qחָ��W6kM!�D��h�2Y���Y�0�0u����;�!�$.|�� aM+�A!n	�_'!�$H;#���E/$���"mF1m�!�DG3,u`6Ì .�����հF!��L1�b���V����dŇ$i�!�$�,1��Q����v�pm�T%Q9�!��lLM�� �T�v�I�!򤝢$�A: �Oݬ%�2C��R�!���#� �*P)Μ
ٖ$H�B��W�!�B2
��i�E4(�b�E��!�DσF�
��EO\ 0� �YFC!�K�U������>u��ãA$8�!�� X\"�^�2�ص�@�*�y�"O*`I4(�8~@q��N�XC"Ol}c�/Z�!��٣b�{�	��"O�1ҵ�I����6-��*�T��d"O��3\�Ja����k�)�  �4"O��Pb2E#0e�\$O��в6"Ot5ò�� u�h��O�|tf�;�"Oh��Ю�&����%[t�C"O���XQ
l�� /�*X��a!D�x��$��M� +A��c� k!D�h���/H�Тæ�*&����@=D��x�H�"5��Ԩ�F	��h����:D�`�W��6r�t��wE�-e*�de:D��*ѩs�T�5ƅA����<D�Tks��b����N��e�F�8D����\�KK����CO#k��@x2�7D�8�5J�83R���h���܄��(D�x�āX�?9�1��ܑ]�vհ`l#D��`ңK!�%���Z�9}�� D��@�>]�>u2��q��$$�!�H/5$r�$(	9Nbi���S�=�!���G?���$�	@(Dy*c%U�A�!�ͼ~�������ȢB"�!�dL�6஬���F���+!�Ă��@2��$m��( Q&!�D�,|��� �Î+�y�.A-W!�طZh�I�$	6(�x`�p#!��9/XI����(A.��r�!��H\�ʗ�ʿ}��eO�3�!��<3��Q��� �Ν�bl0�!�D\f��T2�dY-L����ȇ8�!�٬�����<V���v��)C�!�D_�1����lFoT�5���I�s!�DI�&���J$��Mf:Q�$���^g!�D�E�.�pA�ϋ5��*�EE�G�!�DI�=����-�Z�����A�7N�!�dM*r���V�
'o]"5Q�� �zQ!��д\>"�5A;]�[D�ߊlO!�..T�y.V�`"P�W�5GK!�$��8!�U�J�J��$9�/��;�!�$T�"lBĪ�d�"�Ι��.��!��R�H(b�E��L	��E&hX!�ĝ�MO��I��1
�`i��0hH!��a�t`S �,���J��ըZ6!��:��u����S��<"V��%_}!�dU5}8<�cc�Z����M!��ޘ t&[�n��k�F��!�D�2A4�����1�S'-��B�!��K���R M��<�0� m�6g�!��/�.sG	�3�6\ل��>A�!��**r�-�p/�Ǧ�ba�� �!�D���j(IW�A!5P�=�����!�M�A���)��2d4���&�}p!���t�f �W%ύ[|8����2x_!�dX,SZh��!J�!Ǽ�pdD�f!�RF@���K:y�GcN� �!��]&}Gp��ؚ�,U�a��Z�;�qO0��)�k���:��F�A�\d��|�-Ce�z�L2Ų�)$  �y ��1^�5S���#.�t�b�N(�y��-(6=����78��4*U/�$�y�� � ���J4�0�JN�y�H��X� ��,V�T���!��y"J�(���0�ć�F=��A��9�yr�<ER��雱.�EjĎ�y
� ���#&Ih�0@30����"O�$:@�ڀ���PQ

/�(���"O�U���� � �`�H�=O�,T�t"O�as#a�)��wh��N�N���"O2���M՞mL$���0�~|��"Or�BEa��L���I�O���M{7"OX�A�gq���3O?�jA��"On񣴢� Af>9��,/.�<c�"OT�;�Ս�P嫒nӟ}���5"O��*A�Ӈid �'ȑ<܂Uy�"Oƈ�r	G�/#<<�U�=7�e��"O�Y ��Q�\�JdI9J�.�9�"O�����ަpjz$;�+^o�~�"7"Or X��<GY�9`ba��Vq4"OJp�Hأ"�8��v� |ծ�XV"OH�;���"-=ȨX5GE�s�iiS"O�U�#KφRKF�e����"O �@��ة^�� R*�;�ڨ�"OⵀëT(L�+ 7}�L�itEJ��y�E�FZ* �#�\6n��0�I���y�ʞ#��2���i��f��y�'��ƚ���,D�N��l��LR �yrL a,&t�����W� �G��yүP�v#��"��â�2�sW��=�y2(	?nҴ��Kµ�j(���#�yR�	9�M��!�?vp�+�A��yBb�lǤ�z��S�B8BF��yB�� ?��*3������@ժW3�yB�6sn���B��6�1�c4�yR�A8^�h�d]3w�$���`�y��Pi��˗Ě%>�N��%�K��yR��:e_�m���֕e�Eq�ET-�y�,U�%�8�!�C%վ�fl���y"�R$g?.i���N�7v�@�B�H=�yrM��S��`���9a��x�����Py��R�zt����ˋ
8Z `���S�<�a̅Q)b�	���Y�I���f�<iq�2I0�{�a�;�XX�C�[�<��ݑl侨[�g!S����)D�DZ�.�?J���C���33�Ĉ��k+D�Ě6�S�l��iٶE�;J�^-�v�*D���Y�%6��EH�^���9P�7D���dU"�Ejp R5'|�e)D�X[p��lH1��'
��š4D�����҃��� ��
�X��+2D�(C�	ތ	�����+�x�$K;D�8��\�b���¡B�'.�(T�%�=D�0s֎�<�nP�v!ں%��S��;D��['ɦ&@�$A].Q#�k�/%D���v`�&!���$&�;l�h kg@?D���t��NLh=�a��b���(��;D�z��V�@а��G�\���q��6D�\p�" T��D��o�h7x��f3D����5v��	ö�	�J�x��<D����	[(	�H�SD5�yCG7D�tc�K�a��Q�C$������)D�(����:w���k�
�6I֩�G6D��i���w�tAe+�uX��-5D�8C��H�:%T)�I�|�Z��7D����Ül�Yp�Gִf�r�
�;D�<ԆF�.� ��!&҈djE>D���V.�d ��X2 ۦIh��td;D�|���Ǎ=�0����,��<��'D�H���H�vxJ ���[�D�H1��%D�� �ءUm�e� #���m����V"O�cuoʸ��]�s䞴T����"O�H�J��䐂t+Bd��J4"O�i��#��<In��P*?a��H@"O޽���	#��Q[	� O+p��"Oj��äH�7*Xs6{�!��"O@0��M�wl$D��'�{\�UC2"O���C��q��=�����Gc�e` "O6��'�J ���F�Y+I�\*�"O����c^=�L �N  q�m	�"O���σ���t U�F;g�@��"O�ei3C� ��HH�BLr���p�"O T���A���I��H�#""O }�g+�'���f�(����"O���Șh12u�8Wގ���"O|m�E.1#P��'�ze�*�"O�h�1�ΰf$1��
'c2�;�"O`=�@=9�¸@㛟)DV��"Ox��g��_�@�p#қ>�� "O8���V
 IB�)�!�}�T���"OHH ���	�*��� C/g���q"OTs�D¯>.��7�! �Y�.D� 2�o_��Z��3/�'�j��a+D��;7����Z�O9q�2P�)%D� �'@��I�b��c'�*T�p#�!D�x�&#�=i@:-(B� $��Hӥ$.D�lѭ��M�4�	4�yK�O*D����mN�BUM������Y�Uo=D����H�sd��a'.�4OS��Ve:D��06���YRQc1�;����#D��"� ]:��C�s�l:��#D�����J�&�,t:� �X��-D��i�j��tD(����z8�\�aA*D���w-^7h�T2����OEB5�.D�<xq�P1k�AJd*X�;&�A�B*D�h3��A�I:7�~Q`�H+D�T����xĹS�ȿ~�@�''$D�����a�4b���2j�@)b.D� �"�i��@�m�,:z>[��8D��٣W�b,	�PB�훵��B�(}�񹰧çW8�a!�c��O�B��5���M�h:x��� c�pC�	VQ�=�4K�u���@
�i�ZC�	��&5D�Y	�d(�J�7�.C�6n���x��GV�*�b���bZC�	�_��0�¢B���4I��T(�C��#xN����N����7d��@/�C�	?)*8\�e�Q�;�NH(f�(l��C��J����ʐ<+�v�i�֦Y�ZC�)�����Ļu�F���`к��B�	!H�*�2��G�W�`a�јC�ɡ1�$8�V���^�-!��\'"YbB�I�<��`�*z#�M�,:�B�98�h؂�Ԯn* �*��2h��C��|� �AO��u�1
��#R5RB��	���Qe�!G�
��uO�>d;�C�ɿE�HB �̜�@�)#ɟ�z��C�I��2�bC�6�U���3��C��6m�V���'@x��ãGE�3g�C�	fK^�
��E4w�8p��D�*�pC�:�N��&b"fٮ@�5�MpC�I!rX��S��R�xH���p�C�	�[�*h��̭�T�p��ՙ\�C�I	D(
C^6s���i��e��C�)� n�	 ȃhEY#�MD(Xz�Ц"O��""�#ⱡ/���'"O�8R�'��Yx2�8y���"OR��(�l�zةVO�.V��J"O�ز�ݽwod0�s��"}d���"O������$�X�$�;F����"Odc��X$%�+w�>�X\�"O�x`�a?^��Ę��A���i�q"Op���!H!R�J)F"����iy�"O���g֘#v|��b^�@)��"O<���V�M!"@ч���d$402s"O�ph�,~N��rN&��a�"O��Jǘ#KlA����سG"O�� c�A�u�B1�g��{���"O��ڂ�C�;.	�0͖�7�rE8E"O�aɣ�ٗ`���jҌ�Dp�q��"O`��NO'b�� �L��Rб�"O�X�d�� XJ��%�Y=�|<Y�"ONك�5@��(��C�$��|��"O��¤-\�m�d�yWe��@� p�"O
�J� O�W�t�C�䎽af\��"OT}S�m�d�ұ�Ƈd�
hSQ"O���"ӾYB�"�ڇu���C"O�Xja*�D�ȅ���;��Y�"O@��#�>.4Y�.S,/��i�"Ob�q�$�4TW�P���T�A"O�a�,�"aPz��T89�a"O
T��!>9�X����P�E(D"OPQk�ť�6�Ԧ��m�dt�B"OT����X��ك@J���e"O*,
3C�1ک;��cJ���"O�P�@�ֿ#�M�w(^�e��Ń""O����p����� >�����"OX03ì1�`Y+�Y
N�H�V"O,*��վ���A�f�c��S2"Or\��.��{t�  kΖ~�<=&"OV�tn���Й"jD8`��KS"Oj��5��:ZO��sR�>T��:@"O�e�J�#W�0)3��=Y��D"OI���M��d��R�]#�"O�a�#A�n�rl����`AJ��"Of�d)�z3�\sI����U"O�z��Ld>��r 	�ʀ�S"O�a��c\�B�P��a�i� �e"OxXDǅ�P�j�Q��֯7��i�"O��P���
�t�֠�-z���"O�6J�8dX��R�F0xf�c&"O�U���9yu�0���]2�B4�"O�����>'����ַ��֋�yr���Y��!�$�z��#P�y��Op��$#�X8���,��y�C 5H^ @EA���\�C ��yb�E�O��p��
��#fI��y��� "�L!dNJ�8��S�*X3�y��	>R�$�a�f�?i�0�U����yҀIv��3(�:��I0�yr��� Z-��O���%�ȓ�y�� �K+x���
�Ȍ�j��a����Q����1��ժP�ȓ,�:�� P�@}�BK�[�
}�ȓE]�݉��� jA-D6E����=�&�2v<�,��F$%^`�2X[�U�Z"�*I"�B����O���B�	%W $�rD |"�%J�B�Ic|q�a�;YVMX���Z�*B�)� $%��	���zWgF�F��i[�"O�$��A�b�28pFF� 1��W"OH��f� <(����H�)�"O��$OS`tD��ؕK��!�"O�l��]rΕɶ��Y����"O�9s�C	@�J�z��y�l��u"O*Ї���5�x�vg]3g����W"O�uB�� l�������(�"O��S��3��KՂ5@�Ypf"O&@H�D�A|Fd�� �8�V��"O\K���Cu`�o�>0f��"O8�*����v���!��
�"O���'��6U��wn�1P	H4�w"O�q�be�����I�F��
��"O����GE� �����p�"O�ȓ��3��`#S$N�l�h:�"O��h���N���tH��?&f��"OX�k�61w�!"ƔZkVXSe"O��(҈ֻ&�v=r"fQ���'"Ob�QW՛P�|�wŕ$!lf�"O����L�^�QD�19��H�"Ol8���:P:p�J�%�=;!����"O|4�,�<e�ݘF*Am���U"O8L�[&3�Z�4��->X܄��"OL��&eZ�0�ԡV"��t�aa#"O�aپV�s%��{��(!"O��j��Ta�m�s�J ��h�"O��	lR�j�Ƒ2c�MQz�F"Od�׃?1?�`b�Ǟ�J�\�u"Oe��e�%z.���U�,��"�"Oژ9Ă_  !&�C�B�x�b)2W"OHq��,�x�#B�?9�V��c"OP]���vn�a&�22f�+�"O�d�� N=i�ȉ�`d f��W"O1!�@�
'Ȧ�Zv��F����"OT����;6����@>\�m��"O\��F�r���ԮA.�6���"O���j��k��|[$ϗ�K�>�2 "Oxa�M���0���`ǌS�`�0D"OT�#$�=�4#�K)�d�(�"O8U!�L��'!����m�o���"O0S�9<�Z�-�ɒ��"OizA�A��~ux�"�(,�V%Ac"O>�87��h,���r��D��"O�H��IЀYg�:%o�� �hY�"OP���oئE�x���Kְp*4���"O��"*��΀��i�6$�ʅ"O` CB�A��`�����	{h� "O�T!�a[�R���d�][΍Q"O�:3L'���P�h~�d�G"O���GC=Jj���ț@��p�"O:�H�@E�wpl�B�Ө92]A�"O1i��@0_YSlS (Rm�"On�1g�_�	&^c��5���"O�(��T�� �;f�]�&q�9!�"O��!��-#���*�Kg��0B"O�d"u���n zC��X^*%t"O.Q�vB�8}*Ę��$]&��H��"O�aCb��<J�J�3����	�v"Ol a펒2��;���:a�|1xe"O09-A<2�l�$/��ʌ0"O2�3�G�	%8�u�7���m��k�"OV\#g&�0Dtջ���?|���q"OP��'*�΄ѢbL-�<ȓ"O� t�����&)�|��"��a�&���"O��K�݊�b�F`G-���""Of�0�(����LE�.-��"Ob��[1�ڽ� �gf5��"Oz��3.X� ��W�M�6`h3�"O^4a��IV��T�V�WP���e"O�8���]w!��H�:?�{T"Of=)%��=7���H(A���!"O�S3 �2o
�Q�`V"���4"Ol���@_Qj��F>ǴA�U"OZ@Qr��1�r��g��4S��2$"OXՃa�.l����j�5%v���"O`i���Ҋa6�#עjo�h(�"OFś���8j�:�!iPeC�"O
�+���q�X2�ye��8!���0������a��a����%[!򤁴Z0J��VcM��xS刐�of!��V6?�`r��.oC�QX�I�,9H!�D ��o��WXxa���DA!�$�<�<)C��˴j��p�'ճ2*!���p#��+�oJ3?��,P5\!�S63�t�r�i>��I��2I`!�J';KT�� �Dؐ7�ތb4!���eCm (@+(��9%�+�!�Ĝ�g��(�hL5����ǆq!���ȁ�M�PAKqלn!��r~�Q/A0��:��"0z!�d��DP+�M�ˈ}xQ�Z�ps!�'w��U �OɖeR�*Eb�6B!�k�mK�j�9�L���^>!�Ҧ1����c�W#
�P����H�!��S�2~\u0E/ o{T���e��!��i��x�B	��3_�ɸV��e!�D��l]�@��ė�g0ZI)ƧL}T!��Ccl���lB�Gz��A%T�)�!��ΌO�H��N�F\BM���
2�!�d�J�[��M lJG����!򤃌f	�U{�75�B#�>Sg!�� s4�@� E�3M��J �'�!�dW�1�,��b�8&��	�쉨C�!�SuR���*Y�h(�I���!�%T#2p��8@�ıX�NYl�!���_�~-cF��_�"9���]�b�!������P���L�`%��#N?(�!�dGev�Crʕ���! �44!��@}���)���_Bа2���=!��?$>H9p���,t��cĐ{�!��s����3�,�����Ud!��3�@�vo
C���&ʆ4bc!�$S�މG��8eKn� ����mb!��Lcnm���,J\�R��o}!�D�
j&͈s�5�	 E��_�!��")n�Q�%#��9C�P�C"p�ax"�	�S�[��<'.eZG&'_5TC�		 *�p�$V�Y�"u1���b}�C�I�Uv(Psuˌ��J5{�HG�E�LC�?��miFJ���C���'� C�I�9�j��*��^J��[�K��I��B��2% �b"F&��҂҅GB�	�U���O�8�*�@+־�6B�Ik�x�
�Qi,��C�5<�LB�2Z��9�A�؟7�������DZRC��F����sKT�Lbt�v�W�n`\B�	�e�2��@*�:�H ��k�0�VB�)� �C��W�N�pL����Xh���"O��b�"\�z|qe'׆i`�I�"O6��Uˢ1�L� ��!z���"O�1�Ʉ6J�@�0��:��9Q"Ob� �?L}ʔ�s*��hԋ�"O��9�b_%XH��k��~۾]�c"O��Bʓ$=]dEWHбo�j���"O���`G�R�br6�S�B����'"O�l�d"�slp�UJA���If"Ozq ������ϟ
j�~��"O���B��K-�,��/�m�,4��"OL$:��)�0T�lP�	���`"O~E�f�;����3���C�-:�"O�P!��G�^��i6��/ 2�s�"O� ��H�oSx]S5�2��9��"O�h��ȭ��
1��"O��JD�PH(�%��"�q)�"O���ċl;�}�wl֜,����F"OF��HV=97�5����9�1��"O�ph#��=qޑ�����:�"O}s�� |V�P0���RAi%"O��@�gP�\> ����$6���"O�t�ch�G��ڒ�/3����"O����/;�V�"b��w��V"O�䪷n	�$�I�Ъ�%(a�DJ�"O�|����4U�ج`U��5BX���"O�ձ�'J�p��=��(s-pp��"ObM���j�N	X��
b:L9�"O0�Y�-B��@*�I	2&���w"OX��GOR�Fn�)��N�t�t�x"Oh�:ԇ�,-:hq�R$[t^�"O
��OɁqe�ݺw�!�-� "O���5-O�j鎈�L�4�Tp"O,�cP �5(�P�R���=Q���s"O6����{2�N�&�|paG/�+�!�CI�:@���ӎ}~����8sf!�*yѮUcWaG8%�p��,��
D!�đ-6���$������,�=9/!�+y�qس�A8f��r��S$!�Ě��}@Wɢ=�6�,�!�D�@$���e��G���jR*w!�C�0	��{�D̓}]j��(Y�
!��=(����L��Mp�T����G�!��w�
��'�E� |͐D
�+�!��J�����˖Fg�I ��]�k�!򤟵~Yh�*K+B���%==P!�䔧]��B˕(8�8��I%{>!�䜗Bx9��c� ��Mʶn6!�䏂zM��A��-,�&e��Ͼ`7!�dݓ0��r����pQ2��1�!�$IE� P�3
�����ǝ�&�!��S�y����E�E�J��H�,`2!�������$2B���jȕG!��GZX@<�E����Ht���&0!�$� (W�)�%@�4�T�ȁ�ƫX�!򄅆x��1S�.���8���֥v�!��;b��a���P��h�^h!���<�����~�`Ţ�L؊= !�$E�/��Lv  O��I �19�!�8l$��@�DE�J8j���*�!��:�
]�g�ڨ[yZ��e%Տ!�!����Me�	��I�;`��0�m�M�!�dC�_X��#
�Zh���șf�!���"~��-Q�N�#�|�� �$D�� ��:�$��1���P)ԇ]���q"O�-h4կz-Z��"T�1���R"O�b�H�P�2#��N��u"OH���J�����L�]C�Ȣ�"O�؂3N׼`6ށIf�[ 89@h+�"O��Y��G�@6}�F��6�A�"O�1��eA<�����ں�p��E"O ��& O�E�4�јw���E"Or8@e�A Ȩ�	�/n}hZD"O�h���ָa��iIs��8�R�� "OP���[IG��hS �D���B�"O��GB�
,�:��R�=jm���p"O0K���|0������ d�K"Od�C����
����N^O�|xf"O`\s�N����ۥ�L�M*�AB�"O��!N�6;� �7�:A����"O�-� B�C���ǡ�H�l�#"Oz=���Q���Pp��.TXٕ"O�a�Kl��HA���*��0`q"O2�.]��}�dJ�fz|�b�Z��y�劎7�vi�"k�_�$�R���;�y��S2 �Jd�"$	,+\��)��N��y2��"o�~�(���>*#d�!׏�#�y�PL:�c���3#�\V���y��6'��X�a�ǘ{�V����P�y2삣z���3�@$zm(T�����y"��-��q핪Gz���X+�y2H�"4�ȋӎ��+�N1�5��;�y��C�s��|@@(7�Xi`J�0�yeT�������07�>LS'Lŏ�y"
F=S���s���$1A��
�A�)�y�˂\�ni
Qj5!�~���E���yf��	�*}d	�;T1H�:�y��J
��3����|ȒT��y2oHG*��Jt��
ꡨ�,[��y	HE2��/H�	pi�ǡB8�y�N��\�ʼ� �-6ɴ����'�yC)$ q��k�2~���t�P�y�L;��4@��T)�:�"c��8�y2�ْZ�ۆ�����1B����yr�V/��z�ɚ�L�����N��y�oS�\s�e_�C���Io���y"$�
1�W�2���H�hW�y�X�V�' �t�r�� N��y��_,�8��ѣ�$<�� �R�Y'�y2�[�;��|��H�iNE�����yRn�Z68��DO�}����y�-P�+<u�%�HF]FI�`��$�ybJS]|.	�P .�� �uƑ��y" ��1[��Q��� !�� �$A�5�yB"x����)媰�I�y�h\+=�8%$߸y��YC����y����6��;C��-���2���y�M�jD`#aL1Ht����y"K	o�j�32�%R��=ۑ ��yRiΊ����� �^�L��\:�y����t4.���dM�\��|8�;�y����rLS�t� ���S��B�	�5��t��|*���jƜj��C�=��jVEP/@�ȝڂECU7B�I�g|ƍ0��Ɩ���f�C��60��<�r��/;k(0���:^��C�ɫX ,ċ6�x��K�Y]B�I�Y���"Ȍ�>ߚx҅�X_��C�)� @�����"3�����Ǖ8�쌊�"O�Y�`!C�PߖTȂ�N�R�TI�g"O	�Vm�5d�M8A �pw�Q��"O�*FO�?d��I:!��"9S$TѦ"O�ei�	�M��4{&�3O�L�P"O�������(`�fF�~<�P�"OJ�(���Ua�H�Gd�@2�\k�"O�pP�N��i�0	6(*9�"O�T�c)C��B�n���"O�l�v��O�����_���q�"O��ʦ�K�wy� S@���!�N��"O�$�GMI�mG|��UM k�`ɘ�"O�Ijvb�+X��܂T���� a�*O T�vǛ�o�Sg-�0ɞ���'sV��%χ?)I��c3}���(�'D`�u�Bq�}��F��͠�'Y�0I"nM�eö�#�_�9�@���'���ifd��U�t�!@��;{֘��'"�����E�+�
H�ᆐ	4��k�'��Yh�͈U�z�01 ܘ0���
�'�`[0JV�NT.d@e-Z�#v��	�'$��ޙ$�� J�@N�#�dh	�'�*�� N�(tu��(ۜ�:Hh	�'�L0��ޥN���c�

.�0���'�D��)R�C�� 0.|س�'�� ���-6�y�ţņ#<|J�'jPLآnȈ&(j�H�Y�aܤ;�'��	p7����x��e�7�X��'���gZ��ՍO���"�'�:��Ƙ6bTX���ۘ�h9�'t�9)�ɳg�,�0 ꛞzb${�'�F$����3����M�����'��╠-?)����CG~>��'g�1��	m���Z��ǯ{Sb�#�'#r�K�ݜC'� + �+h�ްH
�'�j��p�]�<h� �'�/d`u��A����	�l�\�De�.8�N�ȓJ�4�F�(n�
�!I.l�@�ȓA�4���/U_N+MQ�WV؄j�"O�h��,G!ҽ�a��bQF��"O��:�G_�W'�4)���Dx��"O�m���c;�-`�ǅ�$=`U��"ODLr��D�9��ѩ��[E|�m<D���C�ț��I�A�4IV\�C��/D�X�S��9=�f�o�� D8�).D�t ��B-GN��j��1�� ��n-D���U��*��ᓶ���iB�8�
,D�ȳ�H�x�U�R��'X���W�'D�Dj4+ȇe&��#`GJ�g��%�v@'D�0�Nu�H���MH�!�\:Q�/D�����&4��t�6Aٺ:�<8�2�"D��9�d�E��H*w�T.}�$���?D��CW�0�>�f�҅e�"�C�<D���Q!OG@z�F}堣rG��y�M�5u�8p]"?8ά��iY�yRlU�%-���ʂ=7Q��`���yR�[���,8b$Bc6`}�kY��y"Laa�D~��]pV��(%
ޅ�'v�����GGJ�Ds�$Y=���'g�U�Q�ąa3ʱ��ZB�I�;���s�� �F�:��$��uG~B�%j��t�#%�>c�&�J�*%.shB��s<d��!Ѻ2_I�tG?_�`B�	!`P%KNU+2�� �S�հONB�)� �taHϠu�(��`U�a��D�Q"O�!��;CF6����3il�0ˑ"Orm��H�]7$x�`�N��Z�"O�S�IK0Z���UI7��@"O�E��2[C��:� �"OV1X��6j�8��A.>�^�f"O* ��!�A8���l�h,A�"OF�IĢ���.8�������"O�M����3b�`i���.��r"O�P��O�5y�Q��/3���ڷ"O\81��8��R�Jh���w"O���`j�*\��0IJn�`��"O�L��	_8/	L=��)H��X��$"O�x���m���"_��Uap"Ox�@Ĕ7�uRP�I��h�q"O�<�֎��5�Z`���@�`2"O�m:р>��48�U=$<��"O�@��q��$�	!tƤX�"O�:�nD20%V�)��x���˧"O֩p$��h	��r7lA�gMHr�"O��B��P�<��⑋�c.�d�"Ox�y��	�A9�|A��'b�B�"O4����au&�@7���m�"O�EA
Щd�@P��m�zh�@"O�@%c�6L�1Qgɟ8���р"ONu N�\��U�ą��谓P"O6A)U��6dF����D�=�L0w"Otxs n^6
�� �vBʉB
�,;�"O�2窈�W������T���&"O�᥄�~6[ړ`��YJv-��"O]�փ�	j+RAʰ,��h���F"O��񤄼������-;Ѕ�0"O�)�4�E>����E'O
\Uމ�7"O�"�H=w�<A*���@��`"O�)����w���t	L@-�s�"O�-�C��/9ˤ!HW�Ѻ^�|mY�"O� �B�I�V�C>��t"O�yI'��$/K ��BY��a�"O�e��L�N�xRq͑�]����t"O �r�&*W�Qb�l!U�<p�"O���sG��c�2�"���?����"O4�3���:�P� j�q�R��"O��{�f�I|N�c�
C	a^i#�"O����ݡG�ƀr#�)Y{X��C"O��P��S��x���K2=b=�"Ox�U@;c�D-y�0D�r(�"O��
&q<qʠ#9Wܞ
�"Or�y��U(Q�ʜ���k��b"OF� ���&R�z$)`%�=�T�u"O����m�,O�� ��2�\q��"O`��l�)m���F-������"O
L�"��9o�X�Em�����"O�j98�*�Z1�������"O��a7�G� �� �`xX�"O�=[5�
��h��d�ئ!�lqK�"O����K>l�l�����Xp��"O8X��ʇ	�}Rg_�T��]�"O�����_���J4䌋�^���*O�)��40��Kr*�:ߞ��'����ׯ�
>��]1GlP�[����'/�U�g):5D|1�N8��
�'�pLK��Ks���U˛/0���9	�'X �Y� �U�`X5j�� ����'���؁䑃{�8C�&B�0��� ��B1�Ξ�����A�k�@�h�"Oh�!��]3*k0r�gu���T"Ob@�eDC�B}����<E�x�"O��"I?%A�� ���)d�KW"O�X��lH�L���)�$SH ����I��T��]�����U4b����7pt�s'�53�\%3����<�I�+q��e�~h�F�*Em��4HY���i�����à�'�������q��(1�&�\=  �8`�z芝Z��e�==��C�#�v{�Xp���",Q�0�Sb�,Q����mڴ�?٪�����O�r�PLSnG�|EL��$G]ƟD�?E���i��*���� �tCӸ3<���)�2�M��ߟ8ѪU�7��9�$E8�ڕÄ�O\��UOM榉�	dy�Om�<!�ɀ�;�V������ �:����H)������	%X��I`��2z�B��S/^�'��]�{6X{aÉ�j��H9�g�b�`7�ʝ[B���S�_��P�V��0^��ȹ��
����A'�|��>�,	��/�\Q��ѻYRk�iJ�����FjsӬ�d�|���ܴ*N(���F�|��+��.< ���?�	��ay���uD(t��$�!Ӏ�p!�D�Ϧ�ܴ���J\w?V Qc��eo�4���T����<1��ݧ~2���'PS`�ƅ0.��K�s�j`�4��,b���f�ᦕ`��<�4(��*���Ձ�
 �i�%�7*U��1j=��	3�S�zp``�7���)�0����:�t�'�>qP���(#K.�)��\��+1��O��:���O�qn�`%��<ǻi%��8)�����AD�`�0,�D��%V��v��h�n	zV�Ak4��c���h���CW�"�M�v�i��y���dӳ@�	�|�cK�4E�JH:��}��ly���DUj�q��$��<q��D�����N0E1��C�\H��1�<��p�������� ���#?�סΝ>P
���.NR�<�r�Q�L|�	ؤc��30P�x�㇚��WA|_� ��	��|]Ƥ�����a)ڶ@@�̱���`"�H�)��'#B�'K�O�Ӽv�ܹ��[�'8����цw�t�<˓3�ha�C��N�tAEI�)�����{�F�iӼ�\�97�i�b���*�:&-:� Rj��)����E����'��`�c^�9�f�v�v��Tȋc��ͧR,Ԡ��㏌lJ.�a�$��P�Ez�F�4Q�!H+%�����ID8���k�ܠ9�OW"{��H7�չC8�`�%@*��':���O\��㦁�I`���(ܑ���<Y�����#�V��$�)��r�	>�0�JQ�ٷ�If+ͅf�f�����ժ޴�M�uW%*��`d�1 ��(�'��E?awG��z��H���4���oZy≬M��[��ɺ'���Ƞ7=������'Fz��O_>+Ԫ�A�1;"b�>����P�q�[0?�n���kWT8tۢ�i�0�2�]e�y�0���\[p� 
�W��`�7%��s�MR�M�a]�� �cG$Y���{� hӴ%P��'�r6MNcyJ~Z͟����-�4�ᥟ)�BA �L���	}���O�Fm`���'D�	�K�h��<r���榭�ش��O��.Hi�2$��O̶Bpd`#�U�=M��'�����7`� p   �   a   Ĵ���	��Z��wIJ(ʜ�cd�<��k٥���qe�H�4m��_;:<��iF�6��/F]�1hA���>ᜭp'*��,.�n�*�MSַiiD�E���$�j�2��['v���Bf�f���Hy�%{��[�'���nZ�^�=AS�M .�B���i�a����xQ�D}��1�'�6��6�J�X�Ŕ'�h��pE�N�pYⲋO� ���3��=[$�qشHE2���'АQ�_y�5�fT�E
g4�52э׽	b6����(-h��E#'���Uv�� �H���d�3X,D�S�q>i�"�̫2��	�/J� ���������$�
b���EFߤa.1Ol���,(|��)t��(ZflhtOe���2ቾP��ѷ��[FvXҢ�j���p���O�=x��$�3��$���Y�����Ĥ㶁I�\�@"<	Q�=�I�.?$���-(6�(i���}�(6X�OD���D������d��`�pqꖣ�#O�j��$L�O��q�OxE��i'g|�	BD��M��qY_�
��I�A�O�92�×:+���ٰlu �#R퇣�OT����d�
�?�e���+N`���n8[@�s�n��#<)��*�D��fz������U��PȤ,�;����'�OhUK<م�Oth�V9$���Ң.GR��h��'V�ʓn�Iv�_��D�1���|2���<��y ���>T\4`���~y"���R�H>�u�Q8&�bq%��� C<9 ъ�e�*�Դ��d{Ӿ��[�'��EFx��]���af�G5��EbF��y�C�y d  ��%CI��b�0!�Z;[y�a+���:m��8Q���!����x$i+`a<��E�!b�!�'=��iAQ,n
T�wEExA!���!:p1���#[d mJQO"!�d�@����`�
*\�\s��	�Py"j��F�)b��*`HLs ��yB�s�v�Tj2(�p��� S�y"��.fD0�u.����&�D-�y�.G�d��������}~PXG��,�ybI
~3�x��+8��	B����y�'�+�p%��)2n<�/�y2����2�A/lz!��]��y��q)\HS�")�R�nB��y��E�0��❂	<��*C��	�y�-�+#Č��@�2 �써B˜��y"��q����Bu��Qr�:�y��S��t+rhW�P   �	  �  #  �  �'  �/  �5  "<  {B  �H  O  ^U  �[  �a  -h  qn  �t  �z  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈m=�R��/{|@�D R�ؖ�_�}�X�stM�/q�L��J�0����` �{L6J�G��,�;�`y��H���{�')`d�5F�y�x�s��8'2aBLR=�>��"o��7&��Ha��U�ѽ�����:�D��6
���0�AGbTI�ֆG:l}�2���δ��*[����S,	�RLd<��4iq:���?Y���?��w���p�Ν^����1�!~/������?ɏ��'I��S��Ip��L	�.D��Hg���@|�	3���'�R惓B7��^�?)�'��4c�[3�0�5�&F�����-I'�R2O�Բ2KRK���ˠ��
G�V�*Q�xFx"�O�e�G*ɺ���[/��%�D&�1a?��
�JC$)���'y��'���'���'���'��cq�Q 'Ț~�nBb���LY�4z��&%}�NDm@�4SE�VB}��o�Y��ٸ�p���99t�A3�F��x2��.xm��@��=��� �B�0$�키�/x�� �N?��je�Бn�?M�;Y:��i&W�����^�0O�[�.	:wJ�Iݴ���k#k���!�l	)}�9����'+v�pJز���V�ѿ$����''B�'�b����x���T(�2Vsx��D�O ��3�S;-e��y�(@8[41�&�W�0�`ʓ�hO>��	�:v�X��L#-���j2$_ğ D{�'�����Hj�z�'D�$���� ||��K@$A.+�>8�	vy�'��>������P��	��/;��6�9�F���	̓ ��`!���6Oxhjĉ��փC���dCp��Tj��˗Es^0��(�+�ax��R��?Q� �Ij)L�C��p���Q�(�;p��D�O��.�)��<qG�W4F�X��IŰ����'|��<�ߴH�d��T�mk��RBcD�?��1BǾi��O,Lh�3�I�?y���@�r�h�"I{���#�Mk�<�Vm���lU#]��a���\�<����C��x��2G����gRN�<���_�ؓ3S�5��Q�l�J�<�C U�`|�� �+N O�iч@SC�<���X�B��=Qdh�"�^!Ae�ş��'�S�OQ��5NJ�7����%o8t��""O%	Ƌ�~!�`�aeW/r��c"O^���K[;8���mE~� ��"O��	IĈZ����꘿0�@��"OX�⁢�+���o��P�"O�FJ�(9������q
J��S�T���-�O�1��f�����"�#u��� "On�������O��P�"OT�Bb��r�t�;!D�;R��u�W"O�
GoD�6Q�"�ڥv_heI�"O�
[jԡl�_R�=
��'gҌ�r�fӢ� ��A�%זT���UO[���I@y��'52�'"�����58�,ݪ#�֦�N�$G�K��ʒd��@����'-axJލ^�|�E�7�*����'UƩ�%g�r�:tX4�}��d��8jv�I5�M#��ib�<����C�-l~�!sOBy$�	ߟ�?E��F�G���qD�?+��!w@�,��?�G�'����G�P�g���p��DeJ�ő����oJ��a�%�U��<��w�	`�CU��ta� iF�|�	�'~L��L]�1�*��GδJ�P���''b���P'�޸�#�ك?5��9�'�N�{w�]-@��`HâW�0��\9�'�A��^ʔ� 2N��[��<��'����� pu�u��N,G�D� �iw�'��)�1�Oa�'Wr[���2/V4��鍌{$�x��,Q���b�G���M��+�9����,��X�?a�N�B�Q�u�Ѡ(u�<蕆[���!��c���F�](���|�p` �gIf�ɭb�Qc
O	A[������_(�nZ)��<v����'���'�@�,ӪkyZ���̖��aI4�'�R⟔�p�җD�P@L�
:����p��<���i�X6�=�4�v��<�F�U�@����a��P�6��7`2�4�i'2�'�P��$?E��N�94���)�"޳{*�`���N���s�딃a(��4�i��tafͅ|�D;t�ܥ!����@�� g.n�e��gb�S�H�?��"�Z�l�Q���F(��R�q�J��ᾭY�O�TR��A٦��'���'
"�'��?�i6����L�7n��]�C��#�y�C�!��	���K�a�cF����4�f�'��I������4��)�8-r�آ�ѭ6�~��N�kYax���O� ��T��=6Q伹SH׮/b,, &�'�0���DD��q*Bǂ���X@D�UaxbS��?aE�|��
k!$���>a�:��Q�͚�yR���H�N�r��Q�\{&��5��?	��'<�,�r�,]��%���[V�hL>�Ì�_W�&�|2Z>=��y��b�BL(J>8R��%3d�����Ĳ�N9�<�Rѧ� Cf�Z�S�O0�HG�ǌ4���h&�<���+�O%�b.�=uY��ԎH�=��}z�O�u��a�Z�='��1�
�`~R����?Iּi;#}��'K҈C���qJI�'�/[��}��'��£�Ϲ,��o�*u�Ƀ���PA�O��<0����A�����5H�,��i�T�l����M[���?�������L�p*J�YV�[4�G<.2���B�ٓ?�|HlZ=J�A��bJL��.�I)?�l�c�(�,z��ũ�dI�K��0��K&O��T���@*\D�i#�3�	�@�\���b�>.p~�8�K�w[F�D�ۦ��	��Q��Z�gy��'2z��1�B������t�b`p_�����5�X�b'��U�P��qʐ/u�|�M#��i��'r��'��D_��)y�n$D��wP+��1A��Ҧ���ȟ��	Fy��� D�}�v��[-�4I�%$�wvaoӫ0"q��k,|��$0<[���#Ď��t��$ b`�Q3!�bt,�R��_�����ܵ:Px�S�3�Ґ�B��\l� F�'�&7m�ئ]�?�!�	�%%H���)�{�<���$^?d�!�t�
�K'�=C��Se��mu�'�����t]l�T�t���?���@��L�& �1dG=�?q+O(�$�O����33��A�ް	/�ܨ�	�����N̾��5 ��x2�C�+O�T�5�' Qdųg��1����|�fC�I��@��S��
!axr���?�����D�4Rhª� y��5��.�l���'�b��S�n�@@��Ā��SG�ZL����D�ٟ$� O�AW<)�E�٪a�,P��L�O��M�|�PU��'����O���	Ǫ�Lb�غ`�Q���O����'<Vjub��l�X|��.F3�MG��l
�Bb4�r��
-��u(7G����ص,5VUꡨnS^�@�R�O��=CRG�Z�A����=����O�M��'�Sȟ4q�@@	5P@\�@fJqg2q�tBP�<a��Y>��|q�kA��̈�UFAr�'��}:e%MD͘���L�d�{֋#��d�<i�����J��?����$����!jMj#
��c�Ԑw9$``q��(�
��I����/�3�/i]�@�f��Zh��DU�+=(`�W�� �P�I�4���a/�3�ɸf���yт���L �L�8x���<?�0l�ğ���u�'Ԅ�㔁_�g[p�S��O�eV��c"O��u�P�[�J\	��Y�`��fV�TЎ��?y�'����I�]Y Yu�U�yɂ8ʄ�V����'���'9�)�S
s��Ыa�AQ��R2$�/8� 9"�n	
-�ZX!���5"�A�����0���{zd���5wE�e�pT�4VȜ���0���J�7U� ʇJ �X�CAk�e�hmx����H�Iw�'��p)D�W!+ـU[B���[u�y	��7D�,j��#����ܽ6ЂY���7�B}r��G
5r�)٭㔅c􋀊v�~=3����!��*/�	� ��k	<��ř,i}!���-�84�0Ia�ᘒo?����P�M��b�>sY�ܠ��ԌL�z܆��L܈c�8�h��B$f\����g�BE��F�
w����m�*At��F{�%	���x\�3n��%�Q�^���9g"ON����,z8�CfU=�S�"OBLk���
O�@d��@�P���J�"O��Q��yހP� 3$�6Ay%"ONN�J��E`-S�_���`�"OX�S��E�"� J���?�=U�'Ԥ	Ӎ���
Ms:1��.�)ow��
��߀r�RԇȓeT(�f��:�n-3D �:Z�q�ȓ:�.�!�"�Bn��{�L�9f����P�@!�Ū�2(Ű�bTZ(ʰ�����gM�bLܸ�Ua�(
؆ȓ� ��g��p�l�p�P�Fp�t�'<�H�x�1TΝ
y�4*���.��I��S�?  �O
�(,��N}O��`b"O.$XF���2�:�m�Y9��y�"O�F��Y���!�U�-:�e�w"Op��PlE`"����-08~(�#�'ǀ�	�'e���W�R�V4m
A�`�'�z|����4�����F��:���'y
��KA!����fS�4�"�8�'����KA�ؼ���Ɖb&r�'�8 �C+[��5 �@�����K�'���Hǫb�0�H��9�R�(��D� �Q?�K�ǌxhl]Y)�p�C5�+D��iDІd��)�:�*�R�*D�8 �I�;�0���B[<kv�q(��=D�(8��ڐZ��p%�6F�\i�5D���)�:S�|�I@=LĐ�r@b1D��Z d��j �2�ܩ@Z���O�OH�P��)�禙{B���zt����V0X�R"Op���'�$��	VD�}yG"O��0�!�nP|L���H8!C�"Oؘ�r�E�ql4���C[����"O��w��M>dSu$�|Zұ�""O,�6��!/��
#�1$Y�T���3�O耲���Y�`��N�*��"O�JŎ�@��t��Ńy�t��"O��Č�)��(; \�P|�] `"O84��a�73��aI��dvT;'"OX8��/J�?Q�Q�;ezz�h��'��Q��'�d���V[Y9�	ȡ<�& ��'��Q��wi�;�S�I���'�T�%�|� �)�G�z�x	�'���زCP�[�(��tƔ6z�:���'�b��UDϽm�IN�'��#�'�j� 6H6n���3e_7!�
T����e�Q?[U�Q(%�T���(�0E>-U�;D�\ȰP)U��A1�34�;b�8D��2��O�/��mXb�\!#q�(��6D������_*�<
`4����"3D���S��1
�p��զ��(\�|��D1D�\��1j �P@�&�;6pr$j=O.�X��)�'4hP��o��^Х{+�R@|x�'���6�`����
�EuBj
�'��P��>�4�Eiկ=K>X
�'�`�� d^K>���1#ȭ�	�'��M�+6JlxnB�@�i��')r��R
[�A��Ih����y*/O����'ab�y2"C�~��$�D�Ko����'���j��D$-�Q�TI,��1�'���Q4B�
YE�����\�S	�'��=�S�/1�xd*T!4Zp$a�'Xd����:
���c�X/�"x��s@܅�5ݼ�k�j�Ju*��Q�����"��(�Ձ]M�2W(�p.�E��P��5Q�ΟUN��d�wT�5�����Ѫ�$z���VL�u�͇�טy�v���W$x�5�:s���ȓc�����C�rg�ѷ�B

�ʌG{�G�Ѩ��1��'V1ha�խl��j�"OE�B��}f|P������#"O��pSJIH�RM��ĺ1l�G"O�dx��� ��"WN�@��0�$"Ob�zj^-d�	A��[�!Br��T"OTA��李OvU!�A�b�I93�'� s����N���^�.�:�Ir�ZGe�-�ȓ[��P��	�F�@`ͤ;<��j��� �ʁ�ؿ?�����j�pˆ"O����ʜ�u�Ȩ�'/uM0�Xq"O�Htg	y��X[6���G�a
"O>�0�Ƃ�fp�]�g�$FN �2�\�<r�� �O +D�S*_^H�g��0�| Yr"O�@`CA]6���cp��<t1����"O(�@�6��J����)|���"O>�{"+��|]h�&;R+u�p"OF �sA��j*L �fͪ|��us��'r���'	
�c4�L�g����R�;AѺ�@�'� AA&Ϲr�R����Z�:u����'��lїǱ? %3a��2���'r&�Ƃ�7>��0�1/��9q����'XlQ�ɘ$W��S��@1
F��'}fQ��AH���m;��)��`��d� &+Q?��튷0�,�ɶF+
p2�IU�-D����Z7D���[�Zc0
�'1D�8a��A>I�	ū�!b�X#%K/D�ȹf	�(WK��𱪖�K;�c2�8D����]y�J�����#>�(Is�n8D�����S!JJX��shZ�[%D��i�O��YS�)�OHL���2>�B �F�0����'r�ݫv���	)P�Z֯�,u�\���'����5́�B���&a�$pӈ�:�',��B-7���C� X��2�'���`䅕��je�#N�j���x�'��)�#A�)l�z}�&L�2�U�+ONt�'"6�B�/I�5�p�"e��A��  �'v�L�����XįI�b����'�X�r��$[�`��hͥ�����'ώ�6�O�+�G�?U�88�'�1��ɎBlPȑ��)<����Cf��g����%B4�ZV��/!4��U�6m�2�^�Dd�����=?�Lp�ȓG�8hH%d��!��	
��'��u�ȓF��ÇaQ�3cr���.�"Їȓ*�Lx��eH�	(�kg��T�\]��~JH$R�o�; Ԙ���%"�.G{�c@��^|�� �8]=��b�$/��c�"O֩Jѣ��Ќ=�2�3�m2"O�`��CѪFU� ��J6~ 8Ի�"OR��$$ݍ;ՠaj��L�	h�c�"Ozd�a�صf���$��T���"O$�2^�<<N8�r�(bI�lQ�'82���Ӽ6&(��W�XW
�jt�3KYȄ���B�c�#{$��Y�lc2�ĄȓjDn<���!&F$�)+��2�,��ȓ|�ȝbeV$����hV�8�X���^%�C�%���x� 
p��p�ȓS�l��n�5P�	^�Fd�E�'��E	�@��
7�K�US�(���>48���dfxIa��׀/�TA&Ø�Iz���=��!��^e`��yE�E�ȓ<��꠪�D:�ϋ=-�T��Kj��C���2�z�ڣ�@�O|-���0����Nۆ}���x)t�p��բMgjC��+D�����ǏL�tUB"�$m5(C�uo�mq�')ng8�Q�G7� C��8%�жG�V���1�ӧA�C�	oS�P�0�B�S�L(�v	g��B�ɇJ4�5�Ce��4�k��Խ1�Ģ=�N�r�O��,§a�7a!���U-S�(X�'��Epb)D1=�a�F�%K���8�'����ϋ�]'�M�"f�.��EY��� �-�ҫ	�R{��*s��K��H'"O 0p.�	9��}з�/\>@�"O����lǀ}Êu�u�@� Y��'0��#����3�:hp��0
�Ղ�̳%����ȓQ�����#Cb��p�U䖕��ȓLX�u���U�(\�0$�(�`�ȓ�Ru`с�A��[e�_	<t�$���\�0DE�Fx�z�O6 ��ȓAJ����	��xz�?R�@��'��]H�
a� ���ɐ v�dZ�&<k,�ȓ����^� �����^	���ȓ�>Q��H�7��0��
1:�����M��)���|Xn$xD��"g��Ʌ�<h%m�;ej��f� ��ɬ|���I�5�$���@f~�1�9+T�B�2lyJ�Z�ɄT�ld�'h)Cp�C�I)r��cE�tN����y�C�	�9��J�Lk�]d��
��C䉘0������|�v��RJ-�VC�	�`��i$�XVѪ���4�=)���|�OM($�@�fu�����ݷ{5$б�'Ϛ0������*�cwA�,dv�[	�'���U��+Z���s7����'�����y�YaF�6�����'� �j0hR�wJ����\�.˄z	�'mN������e�w��9%��1��^���Fx��I�	Ӑ��эޓ[r�I"���
@�XB䉧Uc�-a�#�3x���#���B�ɮX`q҄� v�\�B��ie�B�	�|j�c��Y'j�^(� g�5T��C��6T&\pU���p
�	y�C�I
����P��0U� lZ%�N!p����b��Mbyr��r`�c����#v�xD3���"j��J�	�����O>�$�O$���4)��q6Lς���i>��SjHL�����B6X��H�`f*����a��Aߌ��ōَ��L�#OJ4�4���;,��F�ͫ'��Qq��O��D$�ӌo ���R�>/,�)'̀�F��˓�0?9t
\��ab�I��8�`
zx���+O~��g㉖b4�3��^<{���]�pX��Z&�M���|����?�R�I�:���h ��4)���.�-�?)co�2M��9�dĺO��}�!���� �����3�D�huy��+�3Ox���Y�F8<��e)!vW΢"�h�-�!!�G����d��<������R~J~��O���i�(��| fb��_ՙ�"O�0�-ڡF8q� 4V3zhZ��I��ȟ���!��?]�X�����?B^H����O$�}�x�p���?���?Y/O�iW?x�) ���rl[��D"e�Eʴ�O�`@B�J�U�d�?#<9uL�ybp�e�&!�����J�c��I���v4��k��Ij�T���O&\�l��8d�Ɵ��T�򶟟��)�O��D9ړ�y�@=`��1�����.1[P)�6�y���,e4��(�U�Q�'�?���i>}�	Hy2��-i�<Ps2�	1g5�e�䆵"�0;p�'�B�')2^�b>͋0j��8�ܰz�h��7�^]�dO�z@�VB�4�Ƭq��X���<��KƆ�4�^"YK����Ń��dt#�G[�~x��vb���<�G[Ɵx��!�'E��R��3`�y�����F{���2sXM-5G��!t� 4OTY��"O4��s+y� $J+oev0	�_���ݴ�?�+O�� %��m�'[7L�AE�:%���բ �#*O��D�O���ʙd5�!RI���1��F�ޟ��	2`a`h�PB����o�p">���H�mLq� H/�*Y�,��0 ��$@^dl#���K..=��������O$b>�I%��&���8F�DtQ���<��gǦy���O�.��$ ��e����I����/��pR�jD>���KԊ�W���3^r���OB˓���O@��-�\���k��R�F���	���'>�|I�&Rf ة𲯑���S'y�!3��~��l� ��	ܨ�Ʉ�r��ĉD�
��SK�~�OMzD*U*�m��H�1��,C6��'�4�����?Y�O�OZ�)� @�� 㚃S��4�r�
�:U(��"Ot��W�T96:L0�a�	<
�#�I��ȟ�Ț�D8��9����)�<:E�J&��⟨�3�`�.I�
�A�԰$��!(C�I��(!�&)v��H�)$\0C��/>圬 ���i�D�LC�	�,������3����i� �>C�.U��[�*��Gv�9�� P:dB�	6n�����]�$Z���]�9*�d7F��~�
�8�8p#���%zl-���$�y� ��"(B�:��E#d�,��T�J?�y�∃^X���C��쉺��S��yr;Q�䃕��#sN�͙�����y2�Мq;�h� Hѵh��@�dS��y���V��M롬��m@� ����y��ψ2d�Z���9`f�MBG*O3�y
��A�R�q�N^Oێ`s6BХ�y�)]�
� ��YE4����y��E>%�2rL�{s��b��/�yB"���=rEɆ�:�)�N����O�d*���P��$,�<0a�JZ��B�ɣ)#HZ�����	 &Ļ)�⟐x'�>�D-�.-����A���g傻EA��!���;E��S��'�t=�'(�4S�h�3����I$a ��'1���)��I3Ӳ�'��>�M�<;	����đm'̘��eS��I�~r�s�x�&J�nU I�	�!Z>@��d��l���'�N�'q�Q�K�X�����3��JJApUG�i��a��'n~(XK�H{ӎ'�'5�Jm�k˨V��Cs;vV=�����p�O�OP�>ᔴiRH�.���`ӀF�fL"q`)O.\��>���S;
n�3�;O��@j�L�)6�vx��'��}RJ���<�Es~b��|h��lަc�l��+�d�ͤO@�"A����5�޺�m�<J.�U�W,6H����~	Ψ���?�,_n�	#!�8����K$hM\-a��Go*�$S���?��l"N��۔'>�%B$�\C�<	��4$�:H1���0���	2����Q�'��'����'�Zc�Aq�Ƣ>�̠���O�6KH��O���O���O���<%>�A$N	-�����a��`�Q�(��,�S�'q@��֋܁7h$�wI��{�T��~P�ɡcX�h�pD[����f�d�ȓ8�v|�sa��L�s�B� ,���ȓ(�80+w�T��0��#TG����p�"AH&d�0v��jG"Q�n����Cm(��$iα&IF�BQ�P���ȓFJ����̚�= �@��� ��ȓF)X�ӳE�"-��aUfFS�$�ȓ7��eP�:�������@L��g?ظ�j� f����R �����	�l���W�JP`� \�
B���ȓ9s�H�J;.n~H� ��Y����?��4Zu��٢�pR¼��c��F=C�͚'9�4q�$˒) ��X����qU!I-_�\yB�8e��թbImaz�01"ƈ`�02�W� �,a0�'D*0�f��l��ԪІ:���+g��;`���@�8F������ Jt�l�Ek�$ v�x�w�|2��hw�Yص(�+&Hi���y�� X�A��o΋d�8�Î�yr�\.p�*ͫ�E��a��=�c��y� �@})��!#��|�h�ya^X ��gc@"!P<iC ��yR&Ҥ[��ܨ��,$à�{�Ë�y�/\f��§I��f�@A͌��y����l80h�A�)~��Y!�
9�yRn������ӂG�԰p�O���y��*���Q�	2K`07�݆�y��Y0P)�ꧠ���$��yҥ�w�#����褰m���yRA�1� �c�͇{�t��J��y
� ~� �d�D�$��v,�8I*��"O\�$��"�KUj.]�*�+"Ob*U�&	 IkT�[�C�,"�"O
u�0�W,N&|c��v�%ѳ"O�T���+b����Y���8�"On��j�MDH�/Ȳ"O� ( GY.I�f탠��*�*8"�"OF�z�̓0ഒVL@0*���"OICjZ�vjn�XA�z���"Ob�c@!@Dz�)'k��$�h!p�"O�E#� nr� 
�n�5+�"O��r�ku_L YpH�$`^�9�"O(uP��
jy��+u�ԤB��qq"O�p�R`�-pD�0�T��b9	�"O��6D���`TӇ���V�(+�"OVHb4��:k.�@S�\r���"O��ZW��.����a�� �깋 "O�(��c��tTn�BתZ�A��;�"O��7/MR��̀�OX�f��\�"O���4`'B�x+`��P��Ⱥ�"O|�W� 1�%p��%;: c"O6!1q��V���P��-/��V"O����!ɔ�8��XdH&���"O�}�L�W�i����&�JLxu"O֔ڕ��25j�-��N��?���0�"O�5�B��wy$�x�nI�L?
$!P"O$H��d� +�l��MA�-,��"O��h!n���E��8`&n��"O<�*���'�Z�4J�-��[�"Oy�&�W�B$Zb��-k�Ɂ�"O\�����o��d�b�3NQz�"O�}q� ;=h�I�OB3�g"O~��)��H��$Kv��*(�ٸ"O  K�A�`�貇	ֽT(=�"OЙq2�(Z�}���K�,�Qw"O��b����M�ᏘmҴ��e"O�%Yǩ�"�*M� n	T1vՃ�"Ov(�B�O� �f�&�ܽ ��]�G"O��%;x����TZ�0��"O���v�N`����'9T_$�3�"O� A�LW6Ĳ�qG�H�P$���"OJ	9�F =6T�P�&�)��Q؇"O���al����i��T���ٕ"O���7c�%sn-K��<��v"O��)��4|��z!�Y�v�@)"OP�A0`�p�v�P�F�5Q	Le�Q"O��h��Xvt��GΏc  Ɂ�"O�e[���I�R�R5�ȑ��x�"O荙���1+u`q�cK�o��Ĳ�"O�)Ң�W�R(���S���6"OP�Y���Z��e(�D-2�&���"Ot�PB�X<}�����h��v6R,B�"O����gȪ$~1���H�+��r�"O\t�q���.��n�?�J�C"O`��	rd�%D���d���"OΠi�� �`t*�䏮,mF�b"O�-����I�LP��_z8J-hA"O`G�F����@�*�|`"O�ٰAhE1H:2��D@X(*	�8yg"O �3cIG
-�r�Y�Q�(\��"O0����H�S����!�BДx�2"O�( �C-�����.'8��"O�T���Y aXx7M�F�d+'"O.	+T��>@�P����A���"O� 2 �Ŏ�]ט�:�m�'_�J�	�"O�	��0
�pE��z���1"O@9��b,O)�T��D�R�Ъ�"O�e	r�̦ k�0a��R��V"O�X�G��FX��'5BX4"OD�i��p�%�&�D^O` qV"O�	�RD�LҎ�!�l��O8b��6"O`�cr��"&����,	0"!�4!�"OL�!�ފP�:��1k�!U2`���"Of�(��1qkR��$@�62xi�"O�e1��D �3�M�!?-�	�f"O���qB00�M����X����"O������Pp3�+Ԡ#d�$Y�"O=q��7<��{�l��SV3�"O�%�A9)(ʂ�F|u��"Ol]3�k֜����� @�6���
 "OzTCR�6j�-YfO� �1�"O����o��'�|��r���
�ڽq"O�a���N'cOX��d�&NՂ���"OF4���(����ɀ,Έ���"OT�	`��� �-;whV��D�"OX1���a��]��������� "O �+f� ]�4���I�+���"Or����5rm��pR�Ûl2���c"O��� !Ԕ�{��J��R"O�غ7��>����.�'qHЁ��"O���@ ��0�7��Vf���"Ov�H�닩mq<}vm��~���"O@Ō1Qtt�R�a�;U�d��G"O4����=_Ք@�EG����̙s"Op|�C�N/2j��'�2�xL� "O�)����QEt-Q�L�{���*q"O����'(3�4�چ�ѵ-��u��"Ox����"��D*pDѤ~��ۓ"O`�ӗ�Y�2u����4w�#�"O��i�K�g?"XAh�9}�Ȁ"O��%"��nf��DGroJ�U"Oi�}<�p��Ƅ|b��F"O�������#� |R��:B]��a�"O�]�F�!��͂�/;<Y��@A"Of��f���h!rp�0C/
�3a"O ��7�$3��U��6s6Q*3"OZ�5HZ�Zw"9�jɏ1��0�d"Ot �CmT P��`��A#
��	��"O �{g��&o�T%�d �o�]�"O(�� [�ٙ&#
 ���"Or�0K��"��Y GB�,�X@��"O�lZ��Xl��1k�q$x���"Oj�
�i[-k�"���KW �,��"OV�֠V�E�.�AӍ[,{$͓�"O����*˪+�NiK�̀���i��"O(D)�ҋL�$t�3,�
��i2�"Oڱ�e�����3FE���c"O��pF遤X�P�tdK,
)$��"O���Sj�?T�������|8F"O���F�?"4�B+��Q�!X�"O�1�ʁ�b�8ax��
�@�|���"O����kZ:9p��8v�&\�J@��"O����ն_G�ũB�K�$P"�"OН�э�!2LS�o�:_�8�7"O�L�C�*{`XC��������"O���ӣ��Ȑ��Oܬ_�@�ٔ"O��S��X345���	�u����"O�l�iձm��b��˦Fb���"O� �YAF
@�i��,ɼ!d�%Zu"O��iPɕ� q�L`���)w1�=sc"O⨣1��7�a�,�
8,t)3"O���J���n(1*��`!�(Hq"Orl��G e���0���9	�@X�"O�Ao��,�d�'P�e�(0"O�"�LL�w��Ȉc���Z�p"OB� ��i��ܫc5��$1"O��ꡀ��y�b�����z).�k�"Oz�``��{���(V��%�PRU"O֙���E#c�bъ�`gT,�2"O*�3eF:0�֌�G(�J7e$D�tvÉ8m�6���Jڧ
�܁��%D��S��C'.���r�C� 2�ٰ�9D�ĊQW��b���@ܘ%4��1�"D��Y���	^:�{���# 1t)1� D�� Lȟ_���)�ՠ���� =D���'�����;��)@�e.D��x6�": �s"AS.r��%��'"D�X2a��h��vL�']Ѭ�BP�!D�8�"��_j�,qvi�bB� � �,D��Ȑ�#0��,cD�� 5~���c+D����W6s ]�1,�1	��*D���CE^UҘ�e�;M���&D���P�*Nw�mI�&�<ה����8D�\"D�M�~�ZT�Ԫ��=�k!�,D��d�ͯ5���`�!uQg(,D����TVب4�'�~���ঠ(D��	3+�L&�)b`?p8�Iz��&D��#F��<�� 5�
u<x���6D�(�!�0�l0g�ْn�Z�36A3D�����1/:D ��W�8T1�J<D�DrjX Mݒ�0���;dp0�7D��y�KGs�X�pl\�t6JțC�9D�x� ,�&U�����"=��0*D�d�B��4�� ӑWv�Ur��:D��4X����&%A$��o#D��邷5�D,��I��ģt�?D���䮃sv�$A�鍐�ڜ1RO(D� �wO��a���u�;cᔩ�D�$D�,s��#H�I����ǅ6�9�ȓ%����Z���D��'��)x�':"�	6��"+]rA�̓�	<�i��',TmQV�#9+̨�u�f��	�'�lYsA��=n}�ɠƌتg�p�+�'��	���3;&�X낟]�N)��' l�s�-y(
iPw@�[�
���'q���-*`邸�mM>Z��1z�'L�X��ÄL��yaB�c_�0�'���2®�E3�@�T�����') ���O�/�����y6\@�'c0I�DH
��5�^k2�s�'L��o�9eKT�2��,[��@�<���.6L<3B��8\?欪`�A{�<�7��j}�4뀫���20E(�p�<ѓ��^��ꑥٯ.��K�!�p�<�t酐i�r՚��ڬ.�B�BU�.���C��koLb���$\��m%��B@���(4"9��X���=D�hj���_��IQO� lQ�l�d<D����B��-R���D�cc �b�C<D����2C�&��,^-�r�n;D���&�/a�(�*�n�T���h0�5D� S���!|������\"!#�5D��	�-Ze �`!�����b�	4D�� ���ɂ�i�H�8ҍ�vZ�l�"O�b&�2~TBH�į$gR��y�"O
�{�%�'���Ir�6P���3"O��[7���X	l ��?n)�+�"O�T+��2\�@8P�W� (�T"O2y�偢,\0��щ�!bi�"O�*�L4
��Zg+ɳU
)E"O$�%T%����i��<�I"O4P�փ L~��Oճ �<a�P"O��X�ɑ�n檬O_ ��B�"O�D����R��b��U��ȫ�"O���Ua�U���G�}�D�(F"O"hPiE�5�(@ ����l`�"O��f��1wF��:��F�Ǡ�JT"O`�J�fD�"�&Ap�LY*�X{0"O�=�U��:I�d�;"�G�~�0�"O���eJS<u%B!�����
�a�"O^U;6c���D�� 6�Yg"O0d�Z�đ!Ĉ\����Ď��!��-zS�H�Zh�!��G�!�ě!v$ٱ��=C b�����)�!�$�#3�����.ر�ʘH�!�dܓY6v�0�.Q�lx ��	�Fw!��&5b�(� F�;���j�敇�!�E	t6�)2 ɀn�רY�*>!���#r�0�+�Cҫ8m"�P��cW!�Ć1l8�����*!z��8�D�w�!�$K�|\�d�BFb����ɫ+�!�W�v'a���]�7i];�ʡZ
!�$D�bY����R:!c0��v���((!����@��]fl��e�R<!� �<���jV���q��TP��J�Pe!��X^0���BQXQF�Y��/QO!�$�	���R3���'��ɩ)�-!�dٳJ�Ơ��x�h�Fjʁw�!�d�(��@�biR�.�.z�/�^�!�ՉJZ����a	�z��/�=!��J5���p�M�%�M��G�%!�d�<&ݖ�)��c��K�
Q!���r��f�F�o�Z�T�S� n!���2x�(P+�͟.(�����Q�!���)pc���s�,�~�QD[�\}!�ĐQ�v�鲍�;*㢙X��Q�1o!�$^7j��1`��2F���aW��V!��Oj�X�筙�h9dmz�g��!�Ցu,�#QB�"EѦLC��\�R!�$U�FE�� Y#w��q�Ĥ$N�!���B~I1d�=3�]H�*	B!�䉓O�$� e"�e�%���_�0�!�ě0�j�SDP5hz<���eJ�!���3!v{ť� Q�,uK�(X�!�$5&] B

&cQ̨ؤ"�L�!�$"-T2բ` ��v�)r�H�T!��~���4��a!n�
��O�	!�D��Wd��K�"m����_��!�	�p�@pkl��j �Ua(m^!�D�	���@��b0Hc�gG)Z!�d��i��
��ñVy�1#�غaQ!�$��f�p���Їt�����S6h!��H���	� t��5A��N#P!�G�~��0K�?t�pȠ���)�!���o�<UЧ��
,�6�e�B�u�!��u-�E���W&x��}���ӕ	�!�dL��i1�b�xО阷��e�!�� ��HC"z�Ld�F�7ow��P"O����+\+B������W�~X��)�"O������A����"�/p@�1+�"O���䝘=XM���W���혅"O�Ջ4A۟R�}Qf\�\ʪĊA"O23��B�44�9��s�z9��"O� ���ا@��鳆��.8��"Ove�cn�VG��v5�:tc�"O� �a�G�4�i��K� ��]s�"O�I��b��P��P�U倸˄yy"O�}ԦlSbE@%�8$�<���"OV�xөF��rdG�{�Ơq�"O�	;�M�Q-���C�ǩ~�~���"O�@*P�U�� �HS� }PE"O�i� .��HNH� ��T��D��"O�ra�E�Rb��X�mT�VH�X�"O�B� ��+���Gb�#7�V�@"Oh��G��6��y;5R�-�<�"O�����
%]�tJ����j��R$"O�G���d1P!@�,A�X��"O,�p@d͢oLL��d $o��t A"OJqG��v����F�
���1"O�8�		5�l�#�U�.�����"Or�q�29�i0EhK6=�"O��+��M�-�>���/�x�@�t"O�iW햙F�y��Y���"Oj,��#����s��5��U�c"O.����7k(�L�>-,X�"O�,j�� $�l�tI;M7
�q�"O���ªB�+i@��T�I�1�de"OzU�F�ؓk2�id�P� �ms�"O0A��Ʌ�JTnX�@ȏQ�\��"O���ポ-�Z��V'�$gn�`8@"O| �2Ն��mʄ��>�Q�"O��qXX!p0*
2H8����"O��(V�ڗ΀|���&m7>,�r"O�)�c*τv��u�@�L��Q"T"O�Cs�^�5Tj`���ӽ|���4"OȠ�L��L���	>Ez��"O�h9&H�uä8+)O
��I�"Od]:��ے:5�,	��^�W! "O0H����KG�����+a��"O���uF!L��f�J0�l҄"O�Y���OF����FB^Ȯh*T"O�ʴ"D�H�8ABt��a3v�s�"O�%��*e_u��_�g���"O�����	%A)�)kp��%l��q2!"O��""��6��m���*3Z �"O��[pD�*/v�Yժ	��^��V"OL�c�%�+�v��4'�*L�ʈ�"O6]�n���E�%��,m0�r"O�Q�F�K�IG�؉���#=U�R�"ONA�J'\ݚ��C� '�z��u"O�T�� ǿZ@<�����<=��B�"O^aHT*6�l��ߊ,���*�"O��
$�ȷL�&��V���@�v�1�"O�H
��4��If.0O���"O��4�Щav~�Ҡ�M0!��Er6"O>�����Z����)8s�f,S�"OfњD�rB��j��l,�"O��r�!~]�@�#Ã�$�b"O�P�M��wh �R�~�>�:1"O(q��l`bd����eB�p"O8s����V֌_arC5"O� �IS�FۤU�X=�EN��'T4á"O�d� �+z�X#�GSO��=�`"OF���	��*(��¢�M�l�δQ�"O>�k��3O��ً%�2}�X��c"OԄʤ��n'���b+����U)�"O�)�� N�6)�
�5E����"O"� !�����)��2-�X�6"O�ð���lY�	+	��k��d"O�1�elF0ۨDHA�gx��J�"ONY�
wOfP0��K6v*Ł!"OhD !k�/�,�V��<lb8�q"O>��vKO#qu 4U�eQ�T��"OT��F �'=�pu�f͐=�l�T"Op����d.��	�F#��;0"O�AvD�D��H��FHH "O��֎U�3̊�*��WR�9��"O:<q7��UI��
ݿ���؃"O&A��
G�LM�]�#i*�*xq6"O�e�C�ќZ��1�-�9�����"OrK�,;P,��#P1#�����"O��!�@�~������L���"OR�����MUz���R�l�B`S&"O�X��͇
uj>�Cv
ΐL�( ��"O�D)�'W?2!�(B�(U�Z���T"O�A��n�0|��}kd� 5DuQ�"O����$�Q?x��	C=E��3"O�}�e���%����,�f"OX�iV�k*0}����X�~R�"O��k�-�
bC��QA2�fUaf"O8��7��;hw����P��iJF"Ob��μ��%e�D����"O��&g�	سM��b���:f"O^8E��2>R�b�q�X���"OέاBC<>"�bJۼ�n��"O�[��5I*Q�A$k8��;3"OL���&Y������D�1�.�J"O�)��e���A��<(zQ)t"OBI�C�ȭͺ���A9]|�� "Ot�#4��fÔ���.�,y�JhHs"O �Q�X�iB0�󣆇A����""O�%�E	5Ԛ$�tDה@��2"O��XӉ	�J��jpi	C���P�"O�c �Љ,��Q�7.ٗ-��� D"O�$i��%>�b�O�%����"Ot�b�5!���� ��)�F�c!"Oz�#� ��Y���;��T�:<,)S�"OQ� ��G�Τ
g�gS&���"OҬ��$��FzЗ�J��J"ORd�g)�M}�����(c��ܓ�"Oi�u��Ir��6�W:	��݊�"O�9�amZ5\��!�5��Z "O\(��.�eg@A�c.�"wP���"O�I:6�ŏv�
d�[�Z ����"O8��=S
��N�`^�<��"O���K>R��Q� /�3D���D"O�́2�;к�Y�`��8�"ON8�S"MLh�q�`�3<�P�"O�	� HǦ,���"�]"5�T2�"O��@\I:�q;j��KF(�{q"O�UWd��ΘB�	��Pa*ᨁ"O����'u���G\+�yQ��$��5�<(���8��B����'��� �>SW@�zA��YfLj�'T �P UM<����_pT��'�<�p4�Ό!'dy��!"i#��I��� �<
�ؽKܼ��b�ډ�N-�"OX��w"W$Բ�2���c��x��"O~P)u,@�9P�T��̛�"O�ɩՃ��Ql�9RbLLk����"O���V��Q&� �U�ΊIL��!"O4  ͨG�\�Z��89j��q"O܈�b券Tv�RU��?�	:6"O�b6M��S6�� ��]/I�P���"O�ġ�EM�C@���&ܭ�,9�r"O}��-M�2ON�SÊG��S"OT9+эҡά���#x��]�7"O$��@(� U��X28K�Fк�"OH�s��	�h��
^�W����"O@]PR�
�,R
�cu��r�P���H�<�f�];+~|$�(E�0�h�2�i�<�/�:0f�ѐ����+�n�i�<�Ǔ+4"�$X��ۘB�(�5%�b�<q�L͌yT8�2�C�F��X���^�<ɧ�ˬ��̻���(:\e��Q�<��ܓy f$P1��;�V0X�ONP�<�ef�l(���8f�.���I�<�wi?(]:���ڱ!I����H�<�7f�?�4�o_-0U��dT|�<Y�/�p*��k�d�,*�,%�7��s�<�m� wg�C ��%��5�\i�<q1eG�i���P��'9vl�Y'CK�<��d�6�z7F�P���E�<I��@�H�8�"@�'�����{�<QfW�>��̛�/�&U/���'� N�<9��*c��)��9^&� �@E�<�V���7�,Ủ�I5��8(�]i�<�5k�9̎y��҆mQ�)R�P�<�U�9$�
����F��\���JN�<�bGǢj�Nyp��J�i�����d�<�p�Y.^n�-�sb	�Z���fC_�<�N�J�T�����?���נ�`�<	" "�:ŋ��
�oK�zSF�Z�<ф)��T�Ƽ���@�M��C�N�<��*Թ1�����H��	���L�<1�BŜ7X%�����,k  _~�<Q�ٛ$_� 	�\����q%Qe�<)�Ƈ�W�̃��
�hQ8�(�X�<�c��V�@;ҏ�>j��a#��W�<�2͓!�(�g��7@Vd��KW�<�Tm�4#�z#A�54<�S�ʑV�<�2	^8\Q�fAJ�Tk�#���T�<!��	�o-ܼsb��q�8��p�UE�<rL�]��(0`�;S3���A��@�<9�JL;��e��7Kk��� �u�<�D�3e���p��	�\:{�� G�<1�FËOW~%S i�2 Bh���m�<�"��'�LR�@��s]�Y�%aMc�<q'�_�y�t���H�.Wu�����c�<�����~ �%����3O
������b�<Yw��=C)5j�i_3[V� 胣�[�<I$-�#lF�!�R��a�TR��SL�<���=|�hyG#��W����XJ�<a��H�Zzh������*D�l � �I�<�抙)`L [& �#=0y`%J�|�<9�(�
�d��	�����sv�<a�צW&DR(�D����Gu�<IKب���5휍���Z�<9��#t�T�ꦡU1"D&��
�o�<AR���{z<��H����(��m�<� ��UOƄi
���C*��#6T��"O�h��֓c�Pq����7,�t�G"OnEg�D9/��"%��9&���"O���A�W}����q�;�"OPV�8L�ƬBu�X+kj9b7"OHx���[�6���@�ߣa���"O����p�(yq3
м=��px�"OV����<&��),�_��\��"O2�)F�^K:ys�ɷgǊiR�"O��Q�H��4�,1a�j��M�L�`"O	�!!5�@���@�[���Z�"Ohx�T��Ap�Qz���B�"Ox0hJ�~��$I�	B�<]���B"O�P��H� &��3���l�=iB"O\10��ٮl|��q&eͳo���j�"O ���.�	�����cF�`�lqP"O������Z����`SA,"O<� �;r�S�d%(|���"O���P�\�����޷��Z`"O�j$E�6�b�IƵT�l!%"O(ECu�S�݊���c��I�"ON0�FK�Z��x��j��E��d�"O꘰&-ګu�6���$��?��`S"O2-�T���$�>�7�ڱS��)�"ON�q���_4d�A m�Ny$)!"O�a�Z��)��M�YLx9���y�-��҉���ā~#���bJX��y�嚺{H���7��#-�¤ꐩ&�y"	
���I���_0�!�a���y��
�&�����!x�)#��H4�y�KӆL�$`C�\3&&2ҥ�y� 2�@:��=�����ņ��y�eM:jiz��[$�VD��@N�y�bGt�\5�C˃NT�����/�y��m%l����½>��9�0%���y� ��P�ڌ�U�0�0:�Ċ7�y��7�� ���ʆ*&N��m��y��_���qR 6�[��ʉ�yb�.W吙�� �E&����yR�;hB�Qm�1�"-��F��yr+�i��i�Q�Q�7/���؅�y������?\jl�$�(�y-ʃ0��IWGD>U'z���#J��yrm�*A-��(�!��;�H
s�+�yB ��n��i�k�8(�Hr)�	�yB�(?O�J�IO�_Eڐi���y"�^?$��,:��*G'�сv� �y/ �D���J��F�u륁@
�y��oU��%J�>S�(���%�y�+�*`�<H�eȰ=�"��3#	�y"������)� � �����y"ËJ	H��[�i�5ц����y�k�	V���Y�4��Kľ�0<����آ�C��>}QՋ��q�!�D��f>��R!�WGj����|�!�[7%��z�/N*[Nٕ�ƺ>�!���,?(U���	�q�� Q�_;�!�DDtNЫ �&�H D�؂9 !�̏Fjp���*�6@@Vl�h!��
�Y*��i�B��	j�X�"�!�D� `D@
"��)@���ԫD~P!��A0>��Qh�i[�S�>��i9E�!�D�&r��):� �}��M	���!@V!��&���s�=diҌ`Ņխ|B!�� .�
�͊�e�2H[���*M�,��"O���U*�!2H����?�0"O>u�t�ܵq��1	:��"O��!�B�V V�Ybf�D�,�c"O"������53�$�q���R"O�l{B�B�mx������
&��y�"O<}���.'|@�"�	5f�"p"OZ]�&O^2F�,�B� .Fߌ�x�"OV9�UHK:b"D0��S���KU"OR�x�oRT8<�Ul�T���i�"O��Z�ʍ�%�=B੗�cM�d�"OpՉ���Z���J*=��"O<9�ǅ�`P�1��ԅ�d��"O"t�'�ZAX�і(X��9��"O\�#�� %P5wh 51%�4qp"OD�i!�O(:H��3Ǜ3?�0�T"OTy����� �T��eޙ0�`�J`"O���0!��k�u���t�6)��"O�����x����OЇ�5ٳ"Of����Z�#��E�dOXT1"O��r/��fЀ�ѶI 5��y
"OV��l�"=�Xe��43��#3"Od ��Ψ�6 �3�""����"Oh�%(^�n2Δ�QG�3~�L��"O��Qf��F�D�%��#]��)7"OXai҃U�V��  �F�H��� Q"O����lI+m.<34��Z�@`�"O����ȃy��R'`_d��9"O�%1�n��1��=;& ߥP�e��"ObM���ߚ���N�-dBN�a�"O���w��jҍ��%��{V"O�����;T ����6OvZ��"OP����>?�Q���fL~@JC"O�qx���Lɘ
^�$�A	"Ov���d]�4K>�0�	�,H�q"O��Z@G�l%a�ۄ:lQp"O,�↩�6�x�aJ�	s6dl "O����	_�A���s�K�/�`�"O��Rfc�W7�|id@�8e5{�"O��{p˚!i>�2��9)ލ�!"OB�rpd��]}za��P$i(��8�"OƄ[cOU����;R��"6� �"OE�r���[��2�G4K��"�"O�亥-Ȇy��+��Y���"O~a��<|
��3�B�z��M�"OT�����N�� R�	�V�p���"O�y���� v�Kc(�
�&	 �"O^�I�--NHS�F~�0=1"O"�	���8=����(�H�K4"O�a`��Ø�F�I0$q�0�e"O*���"'2%�����!�.�*�"O�}�v�(E ��.�8EQ�"O8�"B�9p%�8F�	6��lj�"O�A� bY0vH�T:rdҎzzz,��"Of�Ce��^x�:6��KQ찘v"Oh��ƆG-Mό<$��-C�m��"O$�c#ÜGa��"#T�R��"O�y�d�P�x�4<q"���p���y�"O6�g솧~,X35�;y�ԕz�"O�Q��E�T�!4�@bv�D#q"O~��å��g(|$1蔾�4��"O(hq Cl1nH�� : �Rxk�"O�CT�@9V�|}��4(}Q"O<����Z�ugB�hVL#l��@E"O� `���Nåko�QW�$i�`D(�"O���#8�R݃d������1"O����)�$̪���%Z���f"Ov��%�=*Qv=�ΦN�^40�"Ou����
j�$�dIY�|�b"O�l���(��w珡gE���"O�-�V%^�0�H=@��
5X<�d"OX��W�I ~eB@�#T2A�,��D"O($v̜�{�N�a�a�:sڸq�"O���H^)-f�[C@A�?T����"O�A�czoj��JS�Q(��&"OU��[X�|�f�V3ҝ�4"O��)�Q�<�5��"m#�D{�"O\<�#+ɲ4#8���!=�A�"OP�֥��lz���⥚ gƌl6D�,"5B�	�z�0�fM�p�D�`
)D�Pv���u���"��;���GE#D�<�a��5DlT1c��� -��Ie5D�`[���fPX���BZ�t��3�-D�D�7`��?�p�A4��)
�T�c0D�0idKؠ+F\��.Qp����/D�`z�hZ#- �T��;
,�A@%;D�����
x@P�iX�oW�X	�9D�lHw"�>����W$�x��I8D��� �F�,q6�@��Q�/z�\ۓ'!D�H�hD����a�Ŝ(ٶ � � D�0��*V��� ���#K}|�"�8D�����Z�1Q-�:5Tl�D$D�����u&���I��|i3�=D�<@����q����̓z!�=p�,=D������m`^�8�i�|��a�!:D���`EB"C�{��P�Dgxt��9D��R�DH*�(U��α
�f���!D�tx�)/Kʀk�$�52�dH�"=D�0v�/[5̵ku�ĥU�B���,9D���o��m��1�#)B,60�g�4D��a��,����6�\�C�(D���ҶW���*���>���Qb)D�P�ǂ�AK6	�c
�y�l��h(D�8EH[�d���F�tDTr@'D�ܠ1�K�`l�ł�/8Ay`ef1D�\�q�>(@QoB�����3D��5��%�����:"`1��	2D�t;�)��)��#B� +扫�#D�p��^����Rn͓@�t-�6�5D�8`�F �7[����M�XjM��4D�l;GK��z&�'M_QH�� n1D�(�jY�~i�hx") B�I�$*D� ������&���{V3D�43@��l�r��V�RR�x��1D�@0��{�8H��ґe��
�"D���3�C�B]2�2ЅP�]a$�+�%D����Xe�~5R�INh��1�/D���DG���e�f��6(��8+��/D�ș`e��4hȅ�2M��*�*���-D����H�$,N4���6PE�آ�-D���Ǉ%�l�b�? 1ц�,D���-��h����"ɕ,Lx���f�(D���֌�lZI���++�܅��*D��Qŏ��7A��0�_,Q� ���&D�l���D��)�7��Y{���?D�d�����)��[[���@��0D��q���D�)0L�!9�,�*-D��@��F���턞{ۄ(k�)D�� ,�aag�$y�`�Re`��]=bܛ"OtT�2���p��mؐ8"�"a"OJ	b�.�	i_�(�j�9b ����"OR��7�А]pX$J#�&b�ڜ��"O��C`�Ȃ
����Y�6��"O$d{����ac7dP�{]�8�"O2�#�\�h"�����~\:�QS"O���b!Нe�n5#D�&C�`�Y�"O����g	R� �5C��,�d�"O��g��A\��k�C�}��19�"O���s!ӳP����v#	B��R�"OҐ ���-	�
 0� X>rh�"O ɨł�[o�Mi�쌝 /�@"O�ْT�T�MN֔�O'
h�jd"O�y[A�Z6kp�1�Q*Dj*`��"O>Aj�!nu�b�'�>Vw�A)�"O��P�\�},ܛ��?����u"O.%P�
�/U`)����|n�z�"O��!��M�tzTD- IƵcc"O4x )D�4�i{D$�)G=�"Ot@Q�� Ȟ�bW��"1[@�Q"O:���P�N*zQY�V" ?e�"O&��#�>$��Hr� �\�j�z�"O���SD
4!��� �>TQv"O(��Dc��ow�A:�I#��)JA"O,� �fI�]�Q�7j��"�氻 "O<�0��g@�YkG��	��UC�"OZ�iC���NP
CG(\�\u�"O^̨���)w��@�!�@����"O�����)C�ʟ��0��"O�41�o]>`�TU����$ a�x0�"ON�X��C?�pU�!)��!Dz]�"Op�z%lE<�!�Y+�$q""O�qhւ
Gh0�'
ړ)��B"O�: �o�"`(Ol
�iR�"O<P���/�4QVbǴ	�Y#"O�͋� ��<�n�y���lր��p"O��	f���i2��*:4$�I"O����	ܵK,�S&Hh�"O�@!�T�^��� �
E#X%���2"OP����U<m�H��I�� Raa"OT]�V+�o��sd�H�is�u��"O�ܙUoC�!�)�b	ѩseB���"O���T�]�<@\lz�Ú6*��;b"O��{pl�0]ހy2,J4,̰ "O8A���7x�ȱ�D�{�~2a"O�L�Vd��E�� "U�%���q"O�5�bA�#�y� �V�H��f"Oސ��̛'D�.ajr/ے�l�s"O|��g��5}���N>����`"O���Cˤ7o�����؊U���"O&I�%�����q!ֺV�.qE"O����ρ��Uc�b�}��DC�"OF�bE�ԡ ;@A�%.`JI#�"OD��Њ�<��L@"�Q�A�,[�"O}��}��H��)VV�h��e"Of
p�M�3��Iq�j����"O�m���{��������b�"O�hSg
�h�e�jEz]�Y�p"OF<e����%@G���@U�pA0"O��ڻQԈ�㧅�y�.���"O�d�%�On�@Ĩ���7��=��"O8$"aO��j��cnܣK�*Q�c"O����H=��T)G�.er�j�"O� <}I ��A�j@ �MCfZpq{"OR��k�V�C��3Ei Т"O�|�c甐A5d�fJ]�BX�'"O��0�cD�v;��Ɔ�����hW"O�as Ȯr<|b�O�{u�,��"Ol�SG��5�D!ӄW�_��|YP"O���$��.
\،���_��)�"O���㖾beR�S"�H��0��"O��1hH�y�����AQ�)�:���"O\(�H��c�9�w!��w��Y9�"O~�.�R�r��rA��`�Vݒ"OB�*fg5P[J����Ͽ#�T���"O�@X��cm��r��.@�
���"O��z抝+�=0҄�i{T��"O�̱1ꕝ)�H&�;*yB�e"Ol�aJ˕B�Au�ٚ�6d�!"O@�
t(I&0��`��်u��{�"O*�)E�Sh�*颇��(%_ր!"O.�Z��O?f+(�jI�M����"OX�� ��&��-S��U
���"O�|���(?�J�{ J���"OhВ�͟�b�B���IA�v�4��"OjPA���`t��h�1W�-(&"O6�z��-cS0 ��j˧9:�J�"O�ĳc��+p��"��n|���g"O�"`o�ﾴ�"/V�z���"O
	��k�1��K&l��`n:m��"OpLЄ	�M���5- 6a.  x�"O@i�#G[5X���p��z��"O�p��M���O�-v�,�+d"O����+�(ȩW,ѧ"��L�""O����Q>s�n��R�۵X�*D�$"O* �@�?V��Չ��E�\����"O�:!��+�b`���$(�.���"O�+e�	�
y�lᒎ͏}���"O�y�B(E�T�n��OgR��"O
y��^�(i��!!V�u�E"O�xqĦ�kX�%���ڑZL.��"O�qX���8t�=!��P%s'eJV"O��h-�GW ��T�*�R�"O���V����I\ 6 �E�"ON�*��+7������$���4"O, 
���J�J-0 �Y}bjd"Oeq6��s��tI�C�fz� ��"O6�2"
��I�� �qÂ�~c.���"O���
i��I�a��/xG�`څ"O�}���O�!����D���Ȗ*O��VH��"V	�L� 6�T��'�v�J��Y?P>(@�ߦ�2"O�� �Λp#�I; �6"�Q"OQ�Ug�ݶ�0�O�(�@B�"O�ȅ�U.�� �V4+�*-��"O�`z�oɀiY�+j�9@�U:�"O$��Pk�+�ڱ)��E'0��Aa!"O��s���6N��C���%s���g"O���P̏�����ox
a��"O�ph���al�h���4_k�8�d"O�%B��I1N���M^h�x�"O,�z2���R�ްf��,>`l���"O����ĄC���`��;"�`x�"O
}ɒ��%�@S�M�"�"Ot�R�f�24��cg���@�A�"O<�B-2r��Hi�׫R?`a��"O�i1�O�����!1#,��"O� �`qd�E�|�.��r�Ǣn��22"O�1a-F�>�&��l��=�j��V"O
 ���2^��Q�%e��	#%"O2�J͈R�2ݣ@*W�I�^*'"O�����(b�����5�ai��	�$��/�R̛��	�U�ze U���u��L���(f�Y�ѦWX���l�0 �*��(wF�L�`Xs�����P�sԈ��M.3N�L��F��W���*��ۚ)f��[@���)z�y�j�7������J��#FF.&#(X�'؟,�4��h�m�	�-�:����Y�M|�ܴX�4$�i� �p
u�	�$���'��O�i2ғf��l�B����8�Xr!�)�$���	:�M�U�i�����.#5�Y8���q%/��~�'C%?��6-�O���|�6��>�?����MÀ*��$��5Q�%֙Y�䠢c��2�Z;Qރb/bM��NN7�F�b�qܧ��]cU y$`Q�06�z���H����4N��R�;f�^�ȅN^� tX֝;�́�Z u;B������)F`u�¥�"&�=j�.�¦u2���OL��L�����R��M��>l<��[��'V*���OX���O�ʓ�?q�����v��{姗�@�rlIs(��(Om���MsJ>��Ϯ�uw��ȩ[��(�*A)2�*]g�ʓd�q*��$�?��?���NX�N�~bvÜ(M���%		6���"K�	]S!QbȚV:�(Y�����Haf�OLXDx��NF�L�BQ8!���	�o��'W&��'���sN�J�͒��0�3��\%r�.Xo�����@��'� ��C�D�p��>�6��ןx;ڴ.���'�i�����}Ԕ�� ��5-H��Cܓ�=�q��P��$��=~���q��7MUܦ�'����?��'(\t����
FҔxf!�����i	�A�@�'��'���O;
D���x:�Lͪ�`P�̽w�I�SB�  +F�H�b=)�z��	D��yQ�	:)���E"ޡ
�ޠ�FHA�G��)�"e���+��]�d��B��� ��� ְ	H>������k@��q����!�ʩH��[,V�,S�4�?9)O2�d<�i>oZ5`L���ƀ�88@�BT.U' �C�	�gCjI0���&ts�@ߛ���ɩ�M�'�i��I	D�jش�?iO|�w�s��x r��f$-��FϮ{O62�'�R�'ynP+B޺@�Z�)Q�T�]!ҩ�B�|��)oLԸ�A׵��� a\/�HO�U�R����|ˣIZ�l �Z7-dJD��=�H��~�����
,|o����*��J,|P�j�Ȕn����O�ŉ�c��B���d�N�� ��Of��SG�'*�dQa%F��i��P-Si6@�=����`Ӕ6�E/=
N� �[�g����ÝTv���c�Ro�Ο̗���#�<w)2�'ݛK�6�"M���
#�8��H��1��� �ެX�F0³΍��,�PlЅ��O�����8H1f�v~hTS��vb`��!�i�(8H�]�I0�, `,�a��ڦi�1��#8>���u��T)J�@̍�SB��2�̦�Y���Ov����I�IT��M���0M���*�ԭv$��"���A?a���,,OH��jNx�ҴgJ�]P*TZD�	ݦy��4��F��!�Xw��y��m����*�A#.��&�/�<lO:���  �   `   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4m��_;:<��iF�6�T�T�2Ts�V�Z *��4e/s:l���M&�i����W���DS8Jİ�B)���z��5'S~�As�̦N�Dl��{�i�X�'�4�m�,H�4X�*�"����!	>!;f�?Ǹ J��r��L�'�\\J��$j�l�'pHbVO�y�8sm
9%����C�æg�$�۴~�Eh�',��1O�_yB7�ĥ;�]>/�vq���VI�fhV�łw�v�P�W���dF�	RҹZ�DE;��D�3Wqd���ci>%���5�̴��I����@ໟ�3�hO�nPhb��	&�
8�1O� @C�X�)4�;����<OJA���dY��O�-K MD���I6� "��b���h�'���Fx�eRm}%�:h1�D�蝛���6��	6>w���6��1L�D���?�t�#$�!N��vTw�'9�|Ex.�/j|(�9J@���K��fR$Yَ}�Yk�'UB��'��3'�P??hF�[����df`"-O���D@���'ѠA:�e+P�Tcs.�������[�'m\�Dx¡M��<�g␗s�����oS
��� 2��&����T�xb�/Q��+^*������~���y�'��%����']\�1.X?0L�r��G�dH��c�I5B�R���GQ��5W��X�1%n>��K~%������+s���fn�<�f�".��%��1dF�:6�Onj��](��Q�h�(�$�ǻi�r��"ʓ.��#<��������cV��oX�4�4FLq�<Y 
 2  �s�����xӺ�$�O� Ĥ�Ks����'�����8�Ġ�A�Iz�#Ʈ�z��O����O�EQU�~�A=
��p,����rOЦe�'ъ���K`Ӏ�O���OE�4�����a������(i�<nZ�����#<���Ď�� ۼ����.R;y�R�Џ�M�!��7x�&�'���'��o/�ɷ �i;�'˥^�v3F�+�9�ߴP�րDx����O� s�ϐw�}�g�==lY�K����I������"�tɨO<����?�'��=�e���+����%r�}��6Θ'�b�'��xa����5��Y9p�Ķ-f�7��O��B�f�<a�^?��	j�	��T���ؐ0����%ɉu"��O��ؘ'K��'��V�4�TIW V�P$+S�
P   �	  �  (  �  �'  �/  �5  !<  }B  �H  O  \U  �[  �a  )h  jn  �t  �z  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈m=�R��/{|@�D R�Д㍓QJXAA#fN�3�fIk�A(�n@�(�b�iukѬ6&�;6n.�z��4��p��$�$�Ǿg$��ȗ�*�H�:#%*H1�L�
�I���3H��V� �4�Ic)��E+GWذF`F�U� �)� �٘����~&d4��Nbܝ��B2u�%��49T������?���?���>N]1�-y݈13R͂>i��s��?�bǌ+��*O���F����O��dPN-��e�7T��pK!��wx�dݦ����O��Ę�1� ���+2<Or���7Cn]��A\�d0�`Q�	+iCn���f�S���sP,��4bi�JyXF�>������\�L,\��S!����_�I�0 EL�D}���?���?I���?����?�)�>��f'��ˤ������$
E6_������AJش<���Hy�`����	��4���"o�X��D�:y,��P`��
�a�WZ����ƓQ�Ͱ7d8Z�����[8e�V�"#�є$`���:o5�� �43k���g���I�|{��G����p��7R���B?<����#�q`�b
*I���s�g�R�bD���ş �?� f�9=3:$J/X&�X����?�?���0?�f,��@��8Y���;C��h���i�'���'�1��/<��vÈ}���H1�Ӣ��d6�S�Ot �F�ɐb2��#��3W&�䁕�'�ў���*H��{ڴ���
0X�	A����
1!�@�y�T���Iß�ϧh� b�k�`��<>��lZ>~~q�3� S-,T3�
 Ak~t��IIhF%[b�U " ����,!�N�d��B�H�XA�iR�;O�-���'�B��<��O�i/�T̈)!�j���OY�D�I���?�|j�'�X����_=a��P%��r�&\K����+T�4��\q��
4��y,�T�N7-7�	,F,!�?��'DN�@DlٓUoX,@�hH+pH���'��#gQ��1��-f頶�'aL!��Od����0R���
�'�>,x�V^�lC��K@=��'h�\ѷ�Ud����+P S�'��ir�9H�f�Т �(#�t Z��XBlDx���Ik~]��H�<u���8�ʒ�C�C䉂&�
{ӆNkp�@��4�B�	�'Lq�䏝�n͐��T$��B䉺 NlhH K^��l���B��xj@�ᥬ�L�T����`R�B�	�n)Q��86���COG�t\�0&-��I�z�)Qj\���-C��/*OB�	9��"���Y����Ϗ�B��C�Ɍf7�a	X�)����s��*��C�	�K@:���l��hرq�d��C�ɶW�.TC�
�	�F̻6��<j�����l�J�oZe~Qb\���R'����������?�.OZ���Oh���S�X@�C�)Q���B�ʟ�붎L���0#*Y�g �ː 3Oءg#�C�
4�s/�6���L�B	�ё$�X<y��@��+aax¬�$�?)��i�B6m�O���	˩���k���U�s��<������(��,�Ɍ%�^0�6��r�]��'�N��#H@�E:�	&qB��@ 	�^��|!ɰ��y���'_��z�`#vA�L�5�1<U!�$+"�>��!�
K�Ƅ��ɏ-�!�$�f�`-9A͏���X����8V:!�d ;�`5�7�X�@�&kǈ,�!�d�g�ޥ�D��8B��m�b�RNY��dU�[�>�NÀ^G��0GრP��|�l�=F��t�'���'��ɭT�%�5Z )چ)U/�,5zd���V&�|��|�2���C�?t�L�'��O��S��	0��l
qJ�,#.��+�!�<8	`*��)���Rb�~���4؊ �����s_�(��G*y4��:�%.>�<T0�49/�	1/	f�$'��O~�D�OD��A��"E������?�d��%o&<O"��?�B�x�*5���N�B�h�}y�Dw��ln�M�i>��Cyb!�&S�b��C,CEqz3�x�Q��*D0�6�'p��'��s��:Oڒ�"o��&����R�ԅ3�5�8� �^�H��|���S�>��7nP(Tm(�נA,2���ӫǺ]��� ��Kc��*�/��ܴ�;�(O8mc�(=MO��K���U����o�09y�no�ʓ�?���?9���?�ϟ2�X@AJ<x�.�z�i��R�~A�"O؜)b�8	L���G�O�rH��{P�|�rӒ��<AAj��<��6�?Ugƾh�Z��N�?H� $:Ox9!P�)� |HP(�]��Q�eO�\���'�X+���8]j�HŲI��!;�m���ax"G��?a��|^�	�l8QmM)=,�a'OG5�yR.Q�q�T����>���Z�j�!��?��'X"�2����0�@�Ƞg�Ƶ�O>�`Ϡc�v�|�V>��əa=��S`�D�6�"�Ѐ-5�j����y!�ObDQ2AH��[Sf�k�S�O��b@'�p��(��Z#\���O��('Á�u��w%3T�h�XԳ�M{m5Ɠn�0 ����f~B
��?�7�i"N"}�'l�|5�VEʘ4ф �����H����'��й�_A�(s�N\\)X���w�O������pz��E�$����t�i!�V��B�5�Mk���?y����.lxm�ɲzyc���V���%�ګ'�@�nZ�F/�Aۑ�L��d9�I�>��SfE5.h������5(Vؠ���A!\v����&N��S�!�3�I�N,ى�&մ#���q�C��D�ߦ��ɗ!=N\��H�gy2�'��d�R˰pP��uM�t�d^�l���4(!2���P_|�S̛b͜��M��ie�'�Ҥ�'���I�I�rA�dOÉϴ�ذ̏Lgb�@u/V�]��֟ �	hy����1L�z�ڦ%�Ri$8zd�\&A&,�ó^zz��8sH���(i��0a�2=}�a2�C%>�5��� 搅�PA��GT���D ���sjA�uB�v.�?v}�A�' 6��ʦ��?i���ɹ-�$�����Y��tV嗢D�!��>��q˰�
�%�D��E��8:�'�듫�B�)do�T��'�c�A��Y$B�2�Z�M
�?�.O�D�O$��P%$4b'��L�Dp2 �Ɵ�X��H�@���Y��M�&	�m9p�-O̩���b4q#�E ���3e��X�1nĨJ]�(Po_Sax����?!�����92ђ)��ߕP8�f-I="�'����� e��$��\������&������X`�O��-�J��Ĭרl�=�t*�O��t�H�k�T��'���O�yP
J�Vz4�{�U�\��3���O`�D�/6��e�VI� S@��b-�.�MG�ǮxI��RSk֓���������V�Y�F	�4�Yy��EM�O���2��v����V�o4N�B�O2`+f�'���Sןr��E���r�L�c��q�r+�P�<�'�N�'0���ꆫT(p����3��Dz�>��g���2��6E��;00�3�o�O}\��0�E��?y�I�(�	Hy� F�A��T!Y�)I�����T�]�YFg�y{\�䒁A'���4��=t�x����qjEK�g�7c��Y宋�I� ����>��27��$S�s 2��lM���C"��0�Rm�OH�d$���t96 ��7�i�', 5c��i��'-�P�7)�8z˖�+JX��(O�Gzʟ�ʓ7U&��̱T�����0r} ���?���?!�����)�	���1��ǋHt��j�8��iر��(�$����3!����ɖ#\v`D �0*�c���6����oQq$��rL�&|�%�牚p$��x���@W`�!���:���O��$'ړ�O>`�U+ �Qx�Ȉ�ʖW�p
D"Or��d�P�`��u�A�ř}��٠Ô|�j�>���%A�����5U�8<A�%T�Cm~lN<�y�f��*���Wo�.
�j��"P=�y�/��Md<Dx�B m�J�������y��� N�ֈۗ/�,y�p$� &�,�PyR�X� t��aQɸN�6��HT�<�+�5D�r1XE�ׯT�������Q�'��1��I�tt9rt(A���Ʉ�GZ!�o�*�����=z��Q����=!��I�O%p�IRjN�k�0���NۻP)!�$C�pa��JS�6!�F�R6!��`!Ĕ�*�,�"Uiu���!�d1	���򠮟��֝� �
���D��O?��	�W��
���lK*�ɥf�t�<1�Ֆ��YQp�F#��,�`Ii�<!��A4\wr<2b#�t�ڑ�]�<)u#���L�8F�R�\0l���U]�<�5�U�9�8��gV��m3��`�<ٶ��dN���BRE�ހ����[y��Բ�p>�d��5p�����͟Y�6|)�g�V�<� v5�E%�2S&��FU�N���"O>�RB
U�8���+%dQ�Zy+"OX5!ƌ�<$Ժd�Oh��P"O�5��(TZ��8R��4X����'�&�`�'�5Jg�B%O8Gȁ�/#,yS�'��3t �4�<�[�P:8�}��'}�� ��8�LY��k\?��Y��'tzб�&A�u���uG  �x|:�'��`��Ж+,\��X'w��Q��'ּ9C��8,�Mk��x� �8��G�1Q?a��A���z	�FO�>W�U`G�1D�@b5���Z&�b��c����0D�X3�h�*H�e0��\�Bf ����2D��j�`���u����&=����+0D��Xa�U,q+T �墙�L�y�0�"D������$��5q��8+��d��O⡳��)�'H.0:���*�Wc��0s���f D��K�j}���#�	7P%��k;D�lp�� p� �Ϧ`���;D��p��Ri�0�j@ M�A�y�8D�t2Ӧ�1�R5S�H�_e�]���7D�dqFF�R���#%'L�a���@[�Ʉ	pj����f0�9�E�e����N�s�!���~x@�hJ�v�S���
�!�ĝ�s�Мa�K��x&�ؾ�!�$5�AW@+_�$�aD��vP!��-��}80�[�'��Y ��Eh�}���~Rץ:�����P�-`��+��yr��K,�	����B��J��y� �1{v��W�e�dX�%���yr%��E� !A�.�%M�l{��Y��y�*V&�,9x���dd QO��yB�N�Vm�����0zG�Π�hO�|k���/��h��!E31���J���
�C�ɐ<��'
T�<R��Uh�-��B�=`K�M��D	3�ȃ�jDTC�	�FM~Uö"	�D�C3hد
�"C��+UT*�P�'ۙw��Y�P.W�d�C�O��a���A�f�F�#w����i��"~zp�t�Li����Gց��H�/�y��z)J���T��9��V",���9O��(� ������k=��G�dq�̗��J0��R/{�r\�ȓ�0�`��3-Z�ݩ'�[-I���ȓkq>+fe1��<Kclq�6��';���yXhQ�! L�u	惚0R�⩇�!�@\R4m_�/ Ɲz$�ҫ3�FQ�ȓm���PT�4:@�e�H����ȓk�� �@{���Fm�9Ex���h6ĉ*�N�Xv�pn9@���Ɇ?� �	�{f6�q��0"����#���@nB�I��9r�I]�v��Q&蓯%N�C�Io���� �j�,�K���z�rC�		
Ov�Q ���1��
��B�%�NC䉋B����sDR-Y��uD �+�B�I�N�!�A���!x&K�B@�.��=��A�x�Oʂ�BG�R�3<)[�Ȍ9}r H��'8��K�C+RQsŨӷ|�p�	�'�>�K�S��$jt�p���
�'S��� ي�P���K0`+6aB
�'��Uɑ'�5=p�Sv�ʠh�H
�'��dS��l� L�4�­��N���Fx��I̗�vu�wJ� "$@lP��y��C�I���e�kH�h��l��P�$C�)� \*WI�/\	����BRԎH��"O��3.�B��@���֙d1����"O6�P�*� %�|I K�\�4! "O��VmP"x���JǮ(W��|ڤU��q�"�Oƀ�f��U���ę88��$PU"O���u��'d�( Q&C� =f�s7"O�u��-���z�Z$��*���A5"Of�0!9N�xPB���="��h��"O@( 0��/4�"0C��\��R�'%�(��'�}k��p�ep��X0}2$��'��5�c��%�`����9C��9�'n�<(�b���$ܡ��/#�8��'{���&�N�H��!)M�v��9�'�9��ܖ nL�0Fy�^�!�'<���t�L%x������s.fP���$ɰ�Q?1��C�hj��b�Sx��M3D���Uʘ�i�F����H#[��r�B0D���m�V����P�PI���+�-D��wn���D|���M<����0�?D�0�,�!h`�����JW�y� ��m�L��d�	&���@sf��?�&ik����^��g`V�Kq&�:CF 3�:��;D���B���FX�C�1[�� :�o=D�H��)K!0�������H�=D�3*��F���2�9�Lq��6D���kI�����0;P�N2g�4D������82F���@�8>���N�<�%}8��� ѳL� h�c�J�Qw<�Ɂ=D�(��V&"i�YB�J0�$���9D������(���^10����j9D���#	1�>ѻg���<���xS,4D� �nS��\���E�I��d{t�%�OF����ON��%
 !0�q����WD@{�"Op�$dΝL.Y[DeB�(2E�"O| S�9g{��� ��H��t"O��f@�m=�A1Ď�0A�6��"O��횆4l��lH�Ut�S"O*9� �8��]p3	L�Y]�,!��<u�p�~�\��p1���ФWB:Xy�]X�<q�τH���sV�J��(\J M�Q�<�#��
h.�`��_� >@�C�k�V�<YB�V�U���J3I�2��hc��R�<Q�L�/  f�q₃h�b����J�<	DGA�x-P���aL�E*hP���Ɵ�r �:�S�OItы��1�"l���D:Q$n%�"O<ذ�H�D�(w�ǳpri�"O�$�$lǏd�QZ6lM���Y�"On���D�)�т�1C��@"O&`���:(��u��H�G���"O>)Q�k@륎H92�*���m����ć�]�|�&	�9��E!�
z��4�1L��y��1�Bp��B$0<�9AF���yB��H��{��]�t`� �@�I�<y'J�_���o��^�ȥ1�F@~�<I�HT'�9�A�Ƈ	��,��{x��*�
��$�%딼:�E�7Ȃ�7*.��7D��%��W6� i�g�&'@���5D� ��H�<"$���)eP:����3D�0�`��O���AgJY�Ur��=D�̉��J�4��LA� C�tb֨=D�t�F�	�kؠe;c.,7-,�׏:ړ"D�D�TR/�luD$R y2Zh�"c܆�y�M���D��� U_�miҁB8�y��v��YT�U�F�~B����y
� j��%�E�%����ǨYM�=P�"O���BI�_'<�I6!��!c��21"Ob81�X^8�:@Gh���'LAz����,3��Qh#�� @*��� C 	��%�q�� xX5�h*�����4�T��(+��}U�Ӝq���ȓ=��J��ҁv2���]0 �"-��[�H�2#��WS
8P��^1EL�ȓ]��T���)Fla[u�f)��'�Z�J
�/��bFM�.E��DK1^�l���_;��AؒO�� Y��V+f�*хȓ1L}i�#B={�
=�A�VǄͅ�T�萛����<`�$���уY�-�ȓ3"PU(@�~Sz�K�nG�s(����*t������ �xF� b���R�
0~�~C�	'!���`�!ԿJ!�q�pB��\ZC�h��@�6�\1)�hhq�Y��>C�	?K��� ��48#L�Ls�B��6�,<j�̵_hhyޤE��$�ȓẅI��5K�F9�r�R���G{����˒�ȒY\p�g�m&2P�"O(U�(�b?fY	�`�(L.�*�"O>��F�+4��H�1&��
D`e"O���a���Z`�rV�0�`B`"O���	RH{e(�(G�txI��"O�U�+�.Y����X�YPLѨ6�'O�i����9*���@5~�����7�-��L�#�nX�kJ ����6
^Ć�eL =@���1?v`dʡ�\�>S�-��w4��[d`Y�g�,���)ݣf��	�ȓ/��y�Fd� X�J��44������xq��/�˲X��,<[-����􉑇�ě�Si��>��]�(��FߋQ��0�A�4����'?R�'�Bg�"0�09�eHG Ƽ;���O��
�3���S�I*AR�ur�%Rj�x4��CԥH��ƣxgbؗO��R�߁;k�� R�� ������1qR�'r1��lr'�ʽC�F��ٴ@�B(dT�����u�~�Q�!B3q���/Ԫ�R�&�OT<�'��Y��F�h��e`�f��)O��Iq�������Hy]>���ȟ,Z�B�^��Q�_(wY\A��+AßPi���/��9C��\?���a�S�O��d"`�f���%ǝ�k�Be�'�" (E�Cn���H��?% F�C�x�#V�i�����}�<)�k�O�$??%?!�'Z@i�ƠP�O3,8�T��S� �'` ����R�b�HT T9Q�f������g�O���!�яzĶx�`�h��!7�'��I(�^5�����	�������$!� y"F٣}7�)C^��ca�'2J퓄�F�r��Ο�h2��##P6��#��$<*`F�>U2���ɻHN0��ìO�.N�g�'qlE`����O�Y�E�/:٢=i�O<ܳ��'F����<A�ɻL�b�����Z�耤f}�<9�����M�M5�@*�HKϟ\q��4����<	wh�#W��ժq  �2�X�#���?�r�����?!��?q+O1��4�$
�O���@EO��u=�5jL�:q���9`A�z6�P��y�K��T.�q�M'n���Y�CN�rv5�@�PI�T��Oׄ2^�y�m@��?Y4HT�GW���r�\<���Sb@��?���7�J��|�"EB<sޮ���^���ȓS��0�)C�L�"|�H7[�樗'��6��O��#�n��e�I��3�ؒ⏖�`<�A�jV5����?���?�v��xx[�'�Sq�����T��(������щ`T�)���O
�!�_�Ԓ�z�>���'+4r�pè�[8�u�i4*��F|�F.�?	����O�}��,@&X�m�Ů�XxjA�,O*���������NZ�RF�M"L�Q	�2�剕!��Qh(E��(WÕ�1��&I
����T�'����P�	�{�d���b�\u�fh$�
���w^�%P�ȑ[�&�;���?E�4Ek�Pmh#m�p�LlT�_�y2���:y���r�$!�D���>�ȭ۶��+R�1�&%SD�.�	;l�����OV�S�f~
� �a˄� �:#�+�+a���r"O�� b%V��N�RCDȘS�=i��I��ȟ��r�˞�p�u����[�8I{#d�8C���3���t�׊Ľ@�����`X�H�0م�����?(;&0X-\B�Y�ȓ,~&͚�H�	E�f�� %d]����7��QZS�O���H�H�>F��C�I�p�X����)�|�9`Ώ�*�B�Ɋ=�]Kfo_40����+t��d
	�~B�T/)�45�`�D�A�`��C�B�yb.�:�}Q��e��J��,�yR������$\�ʁ��Ӟ�y�g;�T}��+���Ҷ%���y�'��yC�5Bd��#&Zi��9�y�/H�KMb=���ӭ�V=�F���y�F^�>�0�0��ӽ *�����$�y��	�l!�|hW�ܪu��2Rk(�y��3s�ęw��0szh8P&�V��yBoM�u$@;G惶f �-xBmǗ�y��&[b���ܻ-X�09�+М���O���*��өp�>��W '�v,���h�B��:vȘ�If��Ǫ%�c�F=~������O �D*���!d����S�^ `��oS�9��V=�D9��S��'rp	�$L3T�hy�����o�M��I-��<ͮ�'
d�RJ��8@dȡ�(H	�lB� ��I�~��s��8���?+�͋'������㓆�an��'8�'�x��I�豪���R3A�7����%�6l�^�jd�'�P�L����$��	���e�����+�-����Rn�!�OBͦO�ĝ>�i4,���	)�N��eK�� ��+O :E�>���D^�e��UnR�0�ҢB�LJ��1�'��tkM���<q(
K~��Y�Y���P�fI�I���W���O���6������S����yu�>7Pt�a�=^o|���~������?�I�}����c�x��	O�b4��
*�f�$I���?��ϨS�Dɹp�	/X[�(�v�#D��:���;C��x�"k�>�� �`Ӟ˓�?����?QN~��?���LЛ��D�_�z�aa� X���'.2�'��'*�R���m��FU�YnVuPt�\SR`��x��)���l�
9*����w���a�#	<3�B�II/�)`h�m��IHB��\��B�I>e�v� ���)(�)ª8)RB䉝h�r��Я֙;�r)�'lZ�t��B�I� {��CM�7�>y�-%��B䉁H3"���)a�d$�0�F�o�C��
}>mC�&'mX{����h��C��4Nst��6���9gfϼ\W�C��?+�D�Q"KI,r)�M��΍h,B䉭V��U��A��c�\4�� @B䉹?�d8�m�0
0|1���1�C�	�= =(�ƋA��4��!p�����N9	|$*���,�<`x��HwT��s �B�v�T� �+P�y[��`X1	��W,$����៲� �a��Zʄ5S��1dj&�����\h��He�Z6j@Ƀ�&פK' y+$Iq�
�1a��9rJ=Z����8*J@aĪ *5�M�����x@��zH>IA�U4C�ر#0��P�*ј�l	z�<Y�����Pд�Šj��<���a�<Ie���=���V	�v�y3,R[�<�M^,��%�(�\!���a�<Y%	F����B;�4��`�C�<��	PN�.1�b+���p!7CJ~�<�3����L�0��V	V��(#�G�<�D ��/�T��f��=S��1AUu�<A���"�69�1.P�t)���3�Rn�<i� M�[��C������oA��yBI�+�J-Z�X�m	��t�D4�yr'�"or i�*�id�ad�Ʈ�y�O�&u~u���'�p��S&�y
� v���-_��$���Q�.(�"O�$+��&QXN���.Óg�V���"O���DL��zd�M�{�����"Oz��*I�	���bef�lR�"OH�r���<J$�t�!IsX�}k�"Oƨ#�͕�I�|��Ʀ�oO���"O�Mk��O�H�X��/� Q,1��"Oj�)�Ç�sG�B�	�c�����"O����9sӾi�ՇU�F��"O"�0��@V�=B �1,�XEqC"O김���r.�����1�"O6d���Z�O�e�0#&��"�"O�5j�&�|�'��s�� "Oư[�b�"���W�Z�$�#�"OB(�K�,��(�9�hi��"O��l�%}�J��'SȞL@�"O^-{��Su�va�%i1q�����"O��WD��XS�AeG�����Rp"OLE�����Y�n��,֏)��HR�"O���n��h���$�	�=�"M��"O���1�� T�u�,I�/'�(c%"O�!�W�\����.4��0�@K�!�D�9K�]Q��Ŝ/�hp��?�!�D�E"H��vJG�D��!�P�[�!�P!��`P�� @�����M<�!��0h��Xw�=�fr��W�!��G;o������M� �.�`�S�!򄖳l	Hd;1b�y���4GC�*�!�Q5(h��'ǒ,�B% ��O9!�F49[���+I3���!��(�!�d܄O��x���)0�yxŊ�5#�!�X1GB�����R�%,~A`7�F�!��р#���p6I��R��!���T�(EZg�2b�U�����!���/��yN̎{���%��
�!�� (�3`�E�2ۢl��]�!�Ӈ�6��'�V�T1�V��T�!���	�p#���xٸE��;b�!�dP�ߎ%� ��r���FF�!�$��>䦭��"Q4`�n�p�O$h�!�D�'N��и �ѴKg�D�Q咞?�!�U( �҉S�΂�B�A�L�|�!��i��jtF��ȡ9RA��!�3D��Q�0I��C�p��v�Y+L4!�䇑J-�Ec�.\+W�����9k�!��"��r��Q�8�������!�� *[�q���3�*�ô�'�!�$��y��ѐ$ԩ2��%�ccS�!�/RJ��)Ґh�(`s6O��!�D� "$ ��&G�J�����E;K�!�[�j������W�� �䘐y!��V6�L!�f�<�(�(fd5Ov!��T�y���^�n�3FbM�;!�dA�a'�bV=j��!1m!��G���H#�S%X�� 2�C$<�!��F�F[��pa�(p�p [�l��!���t����OQ_�C$l&(!� �G.���X�=R��i�#M!��e���	�j,q�	H��8pb!�dÕ
��}�e��-T�")NW!��c�x �A1(82���ϴz-!򄈬��!�%
9��f�\�r1!�d�j0���B���J̝m�L��'%n�c��,`�2=��ϰa�:����� �8���7��EIUMG�~X�X�s"Od�Y��Z)ȴUa�E�;0p�b"O\��)��F%���-�:JX"�"O�%{��<\0�qի�1�F�ړ"O:'U�f��0r��<?��@��"OI��GD���P�A�s�i�A"O����H���v��I�	}�~�h�"O��y�����5i��d|��30"O��%�>9}���� Uj<܁$"O��8&�~I���¯ԐQcn�4"O��ڃ)��d��A��$J(��!E"O~�j�g�L�6 c�N�@�D#"O4�9�o�]ɪ��IB�t�"O��.�o��x:�ǲ�<��"O��d�i7��Dkoj�`F"O`@
���~U�L	�ܗd@:�qW"OB�`R�dF��C����e�n�"OTYy���p�F�z'b���"O��DN�=,D��Â
)��i�"O$��mU1gtn�����8!�$���"O�3�g��c��a�b�>T�ȵʃ"O�EȢ
W9g �y��,�6���2�"OL$�A��;����e_�W�T��"O����j�0��I�e�Ü8kB"O��Ä�$PR`�#���-���y�"O�@b�bԛp�J0إ�V�Z�\�2�"O�0�fHN�����H,��is"O���J5f_.5�׉ں=����"O҄A@ ��@��.K�`u�"OXqj�	D�O���ekC�C�ܕq%"O68����S�p��S띌Xφ��"Oz��p ��e��aK�)J�#Y܈("O"X)Ǌ��?6��h��}?(�C�"O�8XAD �������F^��ȓM��X��٠ v��%���OxŇȓ'�,�i�MN6�SI֢.��@�ȓB��]�wJ�1G��\�3��JPr �����㰬P�6�9P�)���Ն�G]��P�B	^���c�j�
H����7;��+4�CP�t�S�d�%��Ї�4��2UM����;)׃0N�ȇȓ2�p �Š��[�J�r#��?n8���3�:)g��{оajw�5e��z�� U�sD��p���2Y��ȓo�2MX��@,\�����9��
�'�.E[��K1T�za��ܹ5�!	�'n�A��OH��Z"�Lzn�q�'Y,Qa�G�^���i��ѱx��X�'�
�x�o�����뷀�G�V�
�'�00p,�]�� �ń�2�����'�����N�������X6��1	�'�0X²D��I��$j4,C������'�#��I!^du��/�GLvb�'x�1[�/0�*�;V >=d��I�'�T�;���,x�ǝ�!����'���	�%ч;
)(u"7,tE�
�'UȜ�A)�.,��x��͗�EF��
�'[�PO�� |�Q��±R�9�'{�I:V��5>��� 5�	��'Ҥر����fz�k�k�L��'5���$�&_��Fhd��'T����'ɭax��8ňV8TU��'��u�t-ë�ȥ���*
�@P`�'���G�R���A "�*d����� �\����]�$�wA�?��S"Oԕ��fր\���ATfɫ:ᮩ�"OF䁳`L=)czei!� = �
9��"O�8��D�:Y$Vm@�
B�y�%Q�"O��(���8yn0�3I��v���"Ory��*��������D��&"Oh�ȂDΛ	���Ie�C1���"O %:BA�"�đ L��@��Ub "OP,s��lL���̪|{�)!�"O����{�(�
�NE0]�@��"O|���lO�j�d�
Ug�3��L�v"O�y*3��	��Ɔǰ0v@���"OM�҉ k%
]�"�ʜ68l�ش"O�
���$e� a� ��z+f�b"O@Z�-�hv0�d���{�"O@p�rF	�$x(zW%=$N|�"Ol(z�Ŝ !�t�%�\���j�"O~�s�ND�U2�ҧ�.��5��"Ox9�ց�;l2���ؖKʹ�Cf"O�e�o|��zRKX�HUK&"O��V$M����� 3\;e"OL4Bv�[�v��P�fB�xJ:�P�"O��J�m�. ;v���)<�� "O�,�B�ĝpi�Q�te�#g&:�P�"O�9�S��/W��MZ�$H9Ф��"O�#ʘ}�<u���%F��M��"OZ�!� 4t�B)�����9�qA�"O�� ���MP�p@b�M�v}NlR5"O*��& �/�29�BJ�h�h��"O�td��<�Q2h��y��\b6"O2 ���K�fh=�q��5|����"O�y�v�H�SX�(Q-U#&�ݻ�"O��Ck�3h]T�5��,2�CQ"O�i"DE�b�I�f����իs"O`��'@.z\3/���@�"O&����Ґ�����А�N\�w"O&�#�Ob�؀���f�Y�"O�����/]�j���zH�y��"O"y;7�Ф4�@L�&�۷\D���"O�D�v��u>YX7��1�P�*�"O�����?C,-��R�8�:U��"Oa�w�>61�i�qh4$�(lS5"OJ]p�.�:8~>L���R9a�Ԝ�"O��r���nv<�0�-?wX�#"O��X�	A�����4MܔL u��"O��ye���� M��l^4
<���"Ov}��.=�(�rq
C�]� ��"ObI��CK�4�۶�\;w}B�"O�8Cԁ�9�"a !���5>�h�"O@[2D$D'����fvK�e��"O,	�&îO�
,P�c �q2B���"OV�*�e�8
��p�s�ۇ6Q(�8�"OF�@��IJ~h�"�8]�PP1�"O� Є��_^�=Ab��0tM�U"O>�"b�ݢ@u�m`� �cj,4"O�0`ūE~��� fȠ��u"O��� T ��=ʓcԷc������ӡ]��Er�A'�z �Y�<��'KJ!�^+mҘ����
	�Y	�':��/�#���E�O��VUI�'�h-8��P��`tdF�j	 ,P�'�$���(N�X|�����c���	�'�����5)'j�q6����I	�'��x��՗\�6���	C�	��a)�'>����U)d^�7f�1,����� �Z��X���do��.�Ҭ��"O��(b������1�~���"O���p'�p�L�8� Ý�����"Op� q�ۼנ�#��ΆH�0���"O��6
�[��8 �*Fv�z�"O��WlZ�ՐTi �Rp�)�c"O���WlL�~��UْTB�e�%"OT�㕤�tC���(�t�K"O���V�WB�ĖO^͛�f �yҪ�9=�&�Җa�K����)Ӥ�y�gA_���/��X�0�e?�y2�Z3�}����|�����	�y��1��ڑeۚ&�����^��yr$8	��|wj��%�jMC�-��y��-�{p�2t����£\%�y�k�!/H�p"R�Z��UW��yR׎����` HP&��y�J�T ��N�3�x���Z.�yh��1�"͎�5o�퐅���yr��:����	�0c�Yڵ��>�yR�^8�>���K���e��gE�y�	��F�F�3�,�>85��C6	ג�y%��*z� r��$>S%�!���y�7jqM;�.�2�ୁ`���y��	���T�;<�i+Qf
��y�Ό:|4[C�
.<X�=� L��y�'��:ZJ|�`�69U�:C΃��yb�˯D>]a��*,d�z���y��Oؐ��$N�!A��Q�CR'�y�d�5B�T�!���<G+�\z����yb�I�3b�cB 	�wF`�C�����y� ��X��|�SKňnK�8�d���y�Hg>ND2W���6��a���y��ҴY��{�b&�i�3��
�y�g˸J�Lm���V`= `s���y�E��`��s&�C�9�a�܋�y���<������P�zu{P��y�%��B��� Xp��S�[��y2�2t�:�򣓞i������yb���S�M,U�]�-��y�V%U�n�!�*BGJ�ⷉG��y2��{�����h.y��=;7���y!�.[\l5��d��!'*���yb�ǹ���+ґ�"��+ĳ�yJMW��p$�֊<����0�1�yB����|����1@i�`g��y���5/�J �5bՙ9<"�k0��+�y���RU�b�1�V`ϐ�y��ϦW�1 )��*����@��yr�:�օZr��0�"<*#뛅�y��5o@�	
 ��0�Rh ��H��y���oj��'぀'�����dȻ�y�� 2+1c�K��:��^�yb�܏Q�xxB��-
Č���l��ybիI\�yJ�Y�Q�dA�J�y���б9����F���-��y�צCp��k�L�6�&�.�J�'y�I��^�lJ�H͖\��'� 5�A#�a����rO�[�DXY�'yT��qM���Ѡ�̂�'��mc�'��>*?�Mrb'_�X�2p��'�Ї#�+�n�;!B��W=6��
�'Bn�)G@�ep0oɁIq( 	�'�0,p"�ܳw�� ��kME$������ b�B��8~w�1��	�=� �˦"Oz�{���,"�j�d��;f���"O2�1�Ʉ=�� ��Z4|�n=h4"O2�k@�*w���hw�͝u=�X��"O���C��(Z{�X��ȟxZP��"O��ҵw�	:`Ņ.�*�)s-�B�<qs @ y��`�0�ݗ-�����V]�<�W$�n��ܙ�O�Q� !x�V�<a�$�7�Ѡ1 ��uX��fU�<	���h�L�5�X�>�PY���OP�<1��	�lA��o�
`��Y���Y>�y�mV�{�6sQ���d�5
�����y� ��n����W���Y@���<�y��--44̡un��x@�4�yB���i@�i����݈D�n
��y���i<Ce�ʙB�a�mH?�y2ʌ��Z�Պ6G6��A	��y��K�r���֧\� |��a��*�yrK�U�6hs�ǡm�]p���y��B���;!.����D� �F��yBkA#m_f�C ����0bʭ�y����=vؒ�C.�$���+�yb-N0���$e'&����v����y�*R�cz���D��/(��a�F@��y"e̲��@Z R1\в!→�y"ޟp���w�A-3����T�ʄ�y���?j�|Miӫ7'����f��+�y���c�=#��F vE��@��y�R�&ъy3��Y�2�����+��y�h��D�岖/�:;���zvd���yү��B�BH�1Ð/,N�yF`5�y�)�o��š�E�P��KQ�	��yb+ -������)X8śƟ��y��^)_����@MO�_��H�����yR��=Y�~����8)�|��e[��yRF�)fu����AÀkb�9Q�Փ�yb�D0��"j+�`0�pB�$�y� ɀpɒa������A�?�yr ɊA�ޔ�M���ajd
���y�(�=�R�;3n��6F�@Ï^9�y"K����J���d6�|�2CJ��y%��#�vѡ%_�ew8�E���y�L0q8����e���J��W��y2$�10h褙T�I�ap�<����y2#�<RXn���	-aN<�qWJ���y��5j-�C��v	 tO�/�y�Ї+��L��$�4(C�!�:�y�(��<�*D�@̀�U�,9	"l��y��v��s��,S*�D`y��a�@����͂��q*@�e�I@�'\q�T��6;�N"$'��K�xj
�'��(g�Nf�`�7�_������'׼�3�jT��l O����-"�'�|��쐙dn�h�!A�3�<��'�5�2�!��H#�ɇ�w�f�{	�'\\��,P�h`��PE���"�k
�'<;�Y)���[%�۱픠#	�'�ڵ�E �*v.�gH� H���'I�m�X�[��U�����9|b%�'����D�=�v�KR+�>p���'.��ɴnQ�`�f�Hr���q�F�)�'��0����rN"tRb��zO��'��$x$'C9y3*=1R�Α&��XK�'���#�^Gni�����Q��a:��� ��9��e'6�4��Q��|�Q"O��Q�ȷh:A��#5�L��"O*�e@���0��f�6�(�x�"O>ԩ�Oi,����R9:���P"O�-RƦ�q�\��_��,݁5"O�X�,�8���#��.q6�� "O�|��'�<r\b�h���?�3"Oz�"���$�>t8�N�"6A1�"Op���M�����:�m�(*���k�"O�$�r��)�	3 ��Y3��"Oxd7���&Z�(�X�#i�b"O��hc]�)`��t
�vg*��"O��(�)�-8-�T`���5d�	P"OPI�e�C<��6)K�.N���"O,l�a�	%:�(`� .�;]HJ%��"O&����:e�|(�+P�y�����"O�i�@��@�
mH0�^&c�D�p'"Of�цM� @��+I�Sa&ٓ3"Oּp�a�:c<d�6�ޗAdT�5"O:��v���_lN�"��+���B�"ON9��*��/��sb@E�~d"�"O�P85NU�E���s"�!<�!"�"O�%0A�H@¥z�@l�D��"O��R	�0S_DHڳ'�/�غ`"OB��_8P0�q����LC l!��=N����AF9��E&�g!򤏸Na�pI �0$E������d^!�=�OR�V����� 7!��*XԀ"�/L;�n���� �!�$͉�΁Hꃫ�n�z�I�'G�!򄏠g�`Q��/�Y��@1H� H�!�$K�6<���E��%�V�ܩh'!�8J�>`��K��Y�6yy�"��q!�d��"�h2�ߕC�P5@�
DK!��"���K��(@��2r	�7H!��qݸ`C� �йS��U3N�!�8����BD%~��,aNXk?!�D_�=���i6#J�'�������!��P�l,��fۭp�0]�����!�x8L��#�zM	��V+�!�d���L� �	L�F���)O�!�dգv'$q��A�=R�������+b!�ȻJV�	&�S��0�� A�c:!�F�#mT�SF�M�;�=0���<�!� !�)�p�q�j��EP?04!���CH$�Cf���S�ͰQ!�Ĉ�K,0�H�Q꾅��CM�^�!�DߛC������.��0�G�ȻD!�$5*����j@Z�b�Jd�!�D�&�Pnʰ#X�y�aD@��B�	�Nd|�&cRrLed��%�C�I/S��x:a�+{&��r�9-�C�I�w(��9V)�	F �$v�B䉀x�^��;jF���}x�B�IK ��b��0�:�RDG�3��B䉘Y��5�
L��F4��e�7w��B�2`�:�rGb��X�8���I�lC䉸�ԡ��/�*:��|�6� 48�fC�	�ZҢ3a&�;7�}�R��J�~C��4)�4�x�\�l��5�bO�\C�	�EA���[=vi�!�X�$���c(S�sC�-���6v�"��O;�D#K������ؘ@�T�9&��&J$!�,rI���OșZ��qqb�#{!�M��c6IU�G�!��[4`�!�� |5�U��#z0fl��M�2t����"OdM*��/6x�y�= ��"O�9@�+R07�Vm�g�� �$��"O渫��G)�}�k�:m����"O��XS�>p����-��QyE"OH���IG�8�}┎6��9r"O�E:�W�]��ec�r�ҹ�"O@ �R##gc"`�WBZ���"O�@D�5c� �D���m�,4"O��#�a� >�$a� �B�A"O�5�4�H�K�vd�S���\"5"O|�[�mS���`k0���Ur*) B"O*�a�sȔd�w��4^I��J�"Om����Qs��4�]�\Y��"One�WOw�*h����!�$� "O�0I���������K_�Az& �R"OqG�D��n��Pk
gZ,�"O�}j���N����Ą�JH�Yw"O�$q4+�,5�|�6���	��<�0"OD��������`4�R�8�0�"O�}�Ɲ=oV�@� ��b֬��'"O�,P�Ayȹ�sb�*H�^@ru"OF�p�D�1 ���h"�x�%�$"OT|�v,\
S��H#a�/���"OH�0����(�k�ŵM�d��"O���SϞ�W�R�$� @���"OB����T0)�@K��� �bl�"O蝪�hŀqQD��-�?_�@���"Op)���9�UB%�@/p�!3�"ON)�+'�4�C�+� ��p:0"O�� �Ѡ4����^&{-�l�"OX|�!E�$>��i�"הQ#�!��"O|�L�[��w4�#"O�Y�3�=����c
9{ <�R�"O�`�7*�Q�ҸH�W&W��)��"O��E F9p��  �,=�4	�"O��Jg�؈Q�"��7!T(&>�U�'"O�0�b��s& (���Y�lDH-h�"O��`�ޛSA�9���!3���)C"ON��O�3D�����J�wm
|��"O�pEb
�ro8�jV�P*^O�I�r"OZE�#��[ezUæ��$Z"��"O�YvOܕ�\AA gݤR���"O�}����\<PA� �/A�V8R"OD��0�cK�0�rF�5z�i;�"O��/G-��h$h�M�&�{q"Oȴ��B��n��ѻH��%�t]�"O�*��y��)[E��j�,��"Of`9eL.w|�A�y&��p1"OPAW�����}��Z�18�ipw"O������#�z�@5@��L�s'"O�p���t�rݰiu.��&�!D��`^B�v�Y��9@pd]Z�=D��į�*2������:v�S�?D���T��b4j��h�/X`qp$ D�l� �!c��R��O0:��t)a�=D��cև���� :�c��/D����mr�y@wD�98*q���'D���" 
L���L<��ؓ/1D��Q�j�\�T��q�Y���N#D��ۤ�؀U���z (� 8�|�6D���h�I�@�VHo��ec$`2D�s��$]�x�+2G��W9(1
�-/D��أ!���9Q��
Vu��d-D�� X�q2([�-E����6i� �Q"O���g%؝3:� fo�>5]�8k�"O@{�HD#X���/�e����p"OFhX��O;M�%E�
�� c�"O�8�l�'Ҙ�����%���"O6�E��4>���C��Dy�C"O2���S ����S ��=Ϥ�W"O8��Ʃܪ_�Y���ˋ@����c"O�ك����8�f��_�0��1"Ob�СV0#�CN�T����"O�5iUAS?iOm��M�5��|Bp"O��,b\�m�%��8K�8|�q"O@鐡��L�|P�"�$�g"Ov8�1`ͽ<����(n���R�"O�u冎 Z|-S��q�
)["Oyp ���mo,y�W	]�bD��(0"O�@ �X9'X��]7
�Q"O$�RO\-,Ր�yQ�I*w,N[�"O�EpUG��u_�ܳã\+�<��"O$d�Q<$��iN䍣�"O�ĳ!+��"I��X�x�("O���W���R��Q��1��͘b"O�tGZ�X�8=���N�Z#J!A"O�ȓS���g�����U�P@�)��"Ol$y��		-����wN�n!�2r"O�X�˕e���$J�Jx��d"OV�J�#�+c~��B�С:�p�C�"OB��!��09�tX:BO	r�(@�g"O�$CDW�S�P�'��S�̉H"O��K�sb.�)���1��i�f"O��+�)
�L��bXk�d�@v"O�4���A�,:B����ۇ"O���BB�>�@밯O~�<��5"O��Q�_�df���,ًl�*��2"O|$01���hx��G��qz$"Ov�z�_�n4��Xtn �^�P	��"O��`�=.�x!���))|l�R"O0<H`	�=�L� Ս�" D�V"O�Ku�Z T��ۣ�I#WB�	`"OF�Ce�خ:���(�+�� �|b�"O��1�l��}�AB2놢�4�b�"Oh��Ѧ1TL,(#dD X��Y��"O��[%L1J�����1(��1�"O��	!�@	`�]����r}�ۀ"O0|3wkģy�ՈEȼ*�B�kU"OnE��I:?�l�z�B J���"O�(9&��Qf��� N�H�)�1"O��d�đltay� 9<��	�"OB*ؔ歈p Ή�r���"O�|��'��`@�L��J �c"O6l�K�v����V:J��B�"O4\b�d�+M�9CE�!�Ҥ��"Oe2"��:Mb�1G|�p!�"O��"Ro�Y�"e�`.h�Iѡ"O���dތHd��z�R�3@]�y�OϏP]D��J^�%bQ�1�\�y�ɉ'�p���+���ʒ����'��{���Vq��Ga�$�Cb�ǹ�y���O���V����`<�r�
�ya��[6@j4��KJ�Rr�M1�y2�=J���ʱ�D>E+ur�HP �y�
<��ȕ
ę<q�eם�y��,����ȍa��3�E	�yB��k��\�a��]��t��H �y
� .�;�fü-4:ݳ`R4TᚌR'"O�$��G�4����� U�Dp��"OZ��U#X�A�TX�f�CUx҂"Oڥ����$b:��PBE@�@�i��"O�2�i�||���%ŝ�I+�!T"ObE�a�P�a�h������u��Y�"O��O(d'Н���5R�h�H�"O�t0�g@�'�z���>,��iQ"O���&�N��H�'АP\<=B�"O�B��Y^���@L�9H���"O�|�⋘�&�l�rƎ�=,L�3�"O��H҃A&�f��5d�9t��`�"O�u�G�\�T��D�ےr��"OP�20�Z"h�p4�!-:I�
�)q"Onً�S6Z���B6��c��ᐑ"Of�HS%\��l���lI�[�*ܢ�"Ov���L8b\|���d	���e�f"Ot�J���<M�%�!dP�5��Ai "O�)1AJ�e�aw��3�Li�5"Op5ð���T @90D�'[�n�"O�`W�ҫv���9b�F�awY��"ODQ�tl�Az<���aB�:�|�"O�E�ҺLp2�9��N�4hQ"On��e�ٹ.mD�{�@b�ȗ����y�",�P�!ibz��6�2�yҍ[�H���2�Ib%<t�ӄ�y���3���s��Z{&p����+�y����n�!�ك>�Ա	�FF�y2�<E��*E���>�:4 $.Ҷ�y��ɟAŴHb�A�$˂%s��*�y�̑�@�B�!v��(��$�FƆ�y2+A�$IR�#'S	%���5h
�yb��t�������qPjĨ�y�&��T�pl_�-�T|y'a���y"gؒ��uȐ��%#�<|"B�D	�y�B�Vr!��.e�n����T��y�%�A%2�
Hd>t��v�^��y�M['!��[��N�l�td2v)ؕ�yg�$+���k��gڤ0��%Z�yR��y#��2�˚[�,ћ�D�?�y�杙!=Bh�T��W\0X`��yr�߸�$�q�n��T���V����yч�H-M�Q@9�U�Ұ�y�`�-b\h@!�	Me��b�� �yG�6��t����FJp�S��y��\؞P"�«D8�$1�-F�y�W �����*;:�pl�W!�]�<����-��� #kSx�sq��!�ļ�d5R��Y99jcf��0e�!�DEu�y��Ϟ0<,e��-��$�!� ��YS[5bt�V��Z�!��\�k��lP$N�B�ѽ<'!��!Dd@�%'��l�&� �<�!�$ɨ~���	d �KҸ��AKzG!�D�4rP�H� �r��c����o6!�	ZtpKWIS�^A8���5c�!�5Y���v�G�W/zU�`�|�!�d
J�vDHd�N,���r��
�!򤘻a,���눟n����'�F�!�@#�L����|�2u��@�:o�!��$+.�xE���t����X�!�0��ě��
 jB+��T�!�d>��Y��F^����:�!��f�q�R畦80"A��"��!�� D����؇A�{�V% %�V"OL���KU��\e���ğG	��#�"O�h[c�S0s�q`���+��xI$"O��'!}h,$�����j\�"Oh1�A0��e��Λ.(��J�"O��PB"�;��X�&T:$Lˆ"O�-c�eD�E�%R��@�K�x�"O�,��N�]�d���ޭ1��J�"O����g
(���ț#��̑G"O�]�')D1%<~�"��@!JP�"O�4�`,�)!&�c�G@����"OPܡ��C,$'@1a쑷~��m �"O �B1�`�,�iL\!Dښ��2"O��:�I�8Z�ƈk�� L����"O$��f��,$�
IpCʄ�I�� �"OJ�D$�x�f��hǂl2��"O.A��b��3�.u��H�-�t��"O��  �Թr�c9<nx�:s"Otdq�j���&�X���"O��QT��OAޅ*��1;,�c7"O$����	T�,s0�߅#P�ӓ"O�|a� �3}�ܑy�K6g

�;1"OР�@cZ���pc��I(.�Re�@"O<�� Mt�5U,
�m�D��"OƁ R��@a�1�d "s#��C"O��A �;Om����r�L���"O^��\�9虈$
pZ��C"Op	���t� �d�ER��ab"O��"����2��HAd�H�!�ΚT%��v	F�����c�(p!�$�p%^!�RNU�c�v��3&<!��
C;VZ6�'K�Eb���!�d�m�c��6iSlu�v�0M�!�DF�RZ�qi7�<� A�4T,5U!�D�?n�I�,�?��p/J�C&!򄔿�<M[�/ڳ${r��u�	�!�dJ==p@Pa"O.Lk����Քu�!�d\L�^���O?Y�5��:�!�DȬ;��������\/���!+D�!��J<�+p�W*�� �M�91t!�d��L��7�H8\�\��#���s!��!/rD�@*=F�&�@ �'S!�DîL� �䩓�d���	�&�!�$�r�T��'��~����p�!��5Q�J8�������%憟	!��fb�]0M��s�Paj�%W?.8!��.��@Nv��$�D%�i!�P_�ԁK�A��0M����D4D�`�GoG^�� ���&���
�)4D���M[6� )�a�<9��@6D�,j#�[�Y��\�4�דf4i�4#3D�@��^+5�ysw�ϛ�Q��0D����B\.]�=���	�-��)��;D�j��M�=,¨󄕖|��\��.D���Y%�`�pk��NނC�G.D� i"�.����T�*Lx���-D��ZQdW�y��	(��U��(l8� -D��ե��`�c�c��j�=D��!�K_,6|ʔ��p��I��$<D��H�AR*_�P{BϢx$I
b/:D�`:O�n��@�/�&+�<���k$T��ȴ��RJ�%@�ߦ^�$!�"O]3FD\9j�Y6�F�$���b�"O��X�eJ T���m�?��z"O� r�ru*�~p��[�y���S"O�,�w����`E{�k�^"���S"Oε�U�K1�@
Fm��6e�1X"OH��%L-P%��Cw���Y%��۱"O�󷬊�9@T)
���{r"On-�7�_�1N~�Ȧ�2x��w"Ob�C�M�a�H�4��\�%B"O$����P[t0�d�H�0q�P"O
��HU#:ư�vc�7�2��c"O&�r%T�]@�b5# �q�"��"O����'T"F����$�
���$"O
�3G�^� �����zu��"O���uA�r�����o��ы�"O��$�F<`�\�����a��v"O
%9e�P���4�E]L��)T"O�Q�D�Zy��A��\��U�%"O�`��V�ט\R�.@Q���(v"O�@���yJ�� n�5�ʔh�"O�칅���L+^8��\6m�Re��"O�9�^"wb-8�薠�&�"�"O�@z�*����� ܬh@x�Zq"O.�{�M��6���"X�V�	$"O2�$��@䚄1T��	��dҥ"O�A�����lvQ�4B�s�N%X0"O���7��X�:�Ӗ�+b�^�1"O]��@�!k�X���­z��"O��H �M��);�L�tDjD�F"ObuY�؄]��H���9J���
�"O�]�u��B|�@DM-$����"O~�B
T�-W��'L��r!�}BG"O�l�2K���X@��G�o taq"O��#	]*DM�k�(ʉx�^�X�"ON�:�b&q<�K��p� y3"O��V�����ר>��=�"O&$�E�N��b%{bD�.�Ԙy%"ONH��K0.�6���F'T}���"O����&�-�V��b��PY��"O�<��o`�-X8�䴻�"OȀ�gH�P{`�03HO>}�8őf"O���DŒ8b�t�K��2vh��3"O|�;Bj�"�=9��\tX��"OhY�T����R��T79�� "O�����Z3:Œ��� ��k��q��"Of<�Q�B�RQ%��
�2B�>aCb"O"���&� ����r(�>V�x��"O���,�Q�v�Ac��&�֩A�"O�tH
�S8�h�h��.��C"O8�Z �
2-ȝCq�V����U"Ox�3q*�t~�	��@4�	u"O�‪	.'>Jy٦Y�xE�"OJ�{F�Z�@\\�Dݨu���"OF��h� NQ���s@��c�6���"O�q�gC0-��H��%��u��"O�1*5�Ч3��e�"�͑��9�A"O��@M�Mˢ\���Rժ�b6"O�pc2��W��k�Iǁ ^�J "O�0�Ũŗc@ �q+�"9�8�"O<h{KM�a��4S�o��^b��`�"O���/ύ(�pX�-X���"Ox��@��r���G��=;TM!%"OLęG���.~8�b�[1M@tp�"OJ���䙄Bv��9�H̋8M��"Od�f΄�G6��bjX�4/�	@"OD�b�I;N�zi�Q �5e��[�"O� ��Kpɚ�U��|�)��@$M�"O�D���N�r�a��(T�>��J6"O~�j��ӻ5�|ɂ�JZ�Eb���"Of����:6�%	F�� o��`�"O� �)��x�aB�	%f2,
�"O|)##�B�x�P��g��tW��r*O�ݘe�s�¡���:"1ʅ�
�'��Dc�On�����+L&�
�'!�yh�GÂ.�"���sV���	�'gjq���X�+eB��&G��6��x	�'�" ��W�K�\����'��$	�'����$�	R��@�R��� ��	�'�� A׿J��4��N��)�	�'e<%C�W#~h,(2 �2#ݬ�b�'�2�jJ�,���9Q��	0����'4�`Y�th<SpH��xf���'��9��T��p��!rZ$ �'��9ń��.����%g��B�'���`�س	��}��O�'��S�'F�s�J�{E2�U}z ��'��-�����D3 @ri�j���'�*��N�M�PB��&]E2Q��'W�}crkۄ��4���MNX��'�&����<��1 aD�F���'y�H�v�Y���"���?\��	�'�d����"<$��C$�b�B���'~�=" j
$A86x3�"O[�Lĉ�'O�	�Ac#+�#��Z�dl;�'���qv�R!�c�S+M����'~$�#īB�HwF��v�SG��lK�'C�1x�.��&'�-c�O�'j<d��'����"�>��آ� Y�5!�'{h0���Z9|��UI��Fcxt�
�'`N9��C�5&�Ԁ��	>0�p	�	�'R�˕dRL-:�3i�* �a�'�Ή;���gѐ<i�H�%�X��'o���ӈ>n�.�;@(ʓ�2��' !P����>=�M�5���'o`ɛ�.Ә���kU�w�U;	�'�xY!��Y/|����)�;F��@Q�'A6�9sۙ{Q���cBѱH�8�'��,����J���=�����'?p�F)S��P��g)�<e��H�'w��P$*I"GW/�< ��'�ʥ����}(�!go/�`0�'LZ��1�ږM�Pm�'<�b+�'e�PJA�Τ :�Lbg��m6�	��'x��#W��|V\��ʛ�~���'���VL�I0���I�P�
���'�!�螖*؅#+�S����'�$9*��gz�%�g��FI���'`�l8�#�"^�<I�jڕ�� �'�.��Dɋ!}�r5�X�Bx�`
�'{����,�
~~���G���Z$
�'���@m��z���!�#�h�� 	
�'�\0@m�Ku��{!әW�$���'��y��S/�5�F�S1M�RJ�'����ǍA�
����!�J�d��'zx�r�<��ꆬ� ��'��u���_�Xtx�G��/C�hK�'�8���!n��(�Anͪ9/~��'�[!�T�u�n� ��e�$��
�'�q���9pf9�b�?^��̀
�'ܲy*FN�0n�
P�Q4��	��� (�� ��Uݐ}# ݃�D��s"O`Kr+D�S�v��¹$d��"O�Y��l�; !�����	�k���'"O����ލ"�5#Sc�E�0i�"O��[E�@.o�0���[V0,c��ǟ�`��%T���	_+>YԠ��5o���JO'!��RGJ��	ƟP@$S0A�0`����*V6�a���O�I�k�T��$m�?���c�*ϺKe��X����aE�2�%�c�!I��-K�Wn�8���`ԇ
Nu`�U�چ+�*\��NR�	�*�$��@Ҧ!I|�ش�]L��o�X�jո�.Q6>R���	E��|���߼/e�,XD���Qq��K��IQ�|��o��Tn���9@iB>^�D��ɮ¦��M��X�2!��M�����4�6=����O.��lӞ��m݃~��G�B���EA��.�
���ڴ{ ��K��WS�vHka�	�v�؇C�f����.BB� ��ٽ�7-�#��I�Oň3�ԺW�U8�u�<v�v���B���Ɛ��L����N�mO�a�#�i��p���?�R�i��sӐl��I�5l\R�(P�#�!@"�O��D�O\�D�<����O�ESQ	J7zkdP(�j��4��(��ʦ��޴��u3�y{\w�ؠ�F�=��� s&�1MH�yu �<!V�ސ4X�5���?��?���P��x %dG�_X�9�@�ޖi��x�N�h*��C�=�L���a���\T��h�CU?;����͞�����ޔ$?�q��&M:�tx��� '�>�4��I�C�F���'b�=R�a��D(��l(���O�lw�'�x6�z�'��I:1��ę��ɤ9
��B��W���➼�퉂�J�XѤ�$~N�2@f՞`��(�&�iS�6�?�4�T�i�<�Y��J���ض<V&]�3��\8���s�)�?I��?I��2A���+����P���SN�*b���gΒ\˸YSU�H���ѨK������V.��O�˥jUP���VfRfjd�GMU�Z|0!D�	B{��c��K��7M��$(S�~�	��8���9�Lx{mݮk�8m�Gߑ	�L��a����	cy��'��O��v����oʺ"a�%��"z챃�"O~0�#��$Y�
L˦�_
y��:��O�n� �M�*O�Mp�����J�r��GGR�zh���F�ri���?����?��
I<]�v�	c琰���z���S�.�paU��?"j�[ejR�OvH#=�Q��h�|
Vύ�'\ =3�����F�Ǎ	4)c�	�J�p�*���(G���2� ���G��$�ɉ�MӀ�i�bR?9�gc߳t�zX��N�=7��xBE��?	��OȰ�G.eј�qs/U�W���`�1�O��n��M�ڴo�`E�T-J�_�"x�*z�,y��ES�	���i�U�擡Cc@�IПoڳ��7��'1�,}{u��d�<cpeQź��� q��˧ �����Q����Ok>rVt�Ҥ\��"��E�F+��:ڤR�D^� �����K/|8�lZ�r#���|�1@�<�+0a�Q�V�A�(JX�l't����O��o�ǟ�F��4ED`(0�F�aL���"D�V���?y+O���D\K
�r���gJj}�!
�l����lZ�ML>y�m�8�u��ۏR�H��*ް �x��N�T(��O����1S 8  �   _   Ĵ���	��Z�ZvI�*ʜ�cd�<������qe�H�4m��_;:<��iF�6�T.T ����A���v�@����:S>�n���M�տid�	]����D��}:�f��U�i�5#��K�x�
D��Dh����{��]�'�r\n�e�8!R��G�&y�lQ�$d��X�d���g����'��`V˄G�d��'tX�c`�\ :���	a�[�V^L��W���0�488Ht��'��tC#by�?��,5PR�8��@ǟ\���8R���:f�I������$W�@+���������й��w>=8��$gA�=cG.B�бǎ��Pq�#÷r	�b�8KS�7�1O�I��c�!oB%��. ���[q4OxH��$��O��҅:'����GA�e�М8@��s�'�h�Ex��R}�N��F�"qa[�O�fU˗m�"��	�`��#a��E�4�|Qc�;Q�+�쒹K��fiXp�'^,�Dx�KB{��U15�L� g�۳�>���}��Y�'!`��'�Z��$CCǦ]rF� B6!,O�c���V��'$�S�n��Z�PF�D"�భG�'�)Dx2mɟ���\ �P�2�'ը^8��6�	�^��X�"�xi�,R���qm��Q
��"ł��~�C�r�'�~t%���'_D%q���C�! �jE�y���+��h��I*Ҫ�	���Q��*�k�y>��H=0�P#���=��K]�	"I��18�$��NM� )���x���>(�p g��~ތ���	�.�M{�͚qQ�P��I�3B�u����6p���2�E QªB�	7XW� �  ���yr
�KO��@��ML
zx�T Q�y�'	�Q��#TA]�[QV�q�α�y���?А$�
Ü~����Ad��y2 ��*�q����}K,es��A��y"��=?�*��DV�z��$�E��#�yr@�����#A�P�;"�H��yb���7��(#�ް-@��f���yl�%u�~$�5�)v�(����*�ynDҒLAe�H$ ��y��+���yb�X
t����;tĀ���Q�y"��?
� ��@�yJ���M7�yϔf!,q���7VH��Z��y�a����6�SN�P�p����y�"͞#�`"֏8:��b���y���>[^T�9�d +0k�x�S�y"ˁ������H5`��ˢ*��yR�y�=����XW&q������yB+�/,�D+��[�$�8a���yb͎�l�{ ��7e���p甈�y�h��r�f���,YP	��
�yRA����u@ �0T	A�����y�,ΊL�0�"β)�Qg ��yb�GBނD
W��f����j��yα%d�<���cM�8��ሬ�y
� ���5!�K>rB G2�@U
!"Ol*���U����C���:]vQb"Oʸ[P�C*"��= ��q%�C�"O�� ��#ߠ�q��c��$:w"OHX��м͘���74ݸ���"O ��A�M���1�D��2#~̨�"O�-���i lH��"@*k&��"O,Ms���F�������OW�T�"O�@�f,ڣVsZ�3��'C8�h�"OP����5,�h��o�v6�	"O�)H����z���n�!'D%��"O��⃇�5#���p.Ez""Ot\�P�� ���Г�T��+ "O��S��f2����&DZ�9�"O.QU��+ީ0�-��C�ً"O�J��1ܸ��2����"O�4�&��63P���0�U��"O2L�iGYl���@�< �X|sg"O,�"c��.W�f�I�΂1�̴$"OP�+��d\TͩӮ��|uqE"O�"e�	�L���F�t��H"Ofi#���5ȝJ nL�>�X,��"O(��BC�F���I.ȑc���j"O�JSkE�.�@(���O��	*�"O։;��'fxBM�����xf*O��o�<8����#
�d�Bu�	�'���0���?T6HY��EE�/�(�
�'F�3 ��X�j �²)����'��Mɂ��{��!��_K�d���'V��N݆f����T?�|�(	�'�H	��]>�	��ڏ5��59�'�H�s��\9�t`aL��)�����'�^ ,;V��1xC�7�����'���1���Vر`P`�1+Z���'�XT*ͅ6=	 �@UȒ�'���'>jA�P����5�բͿur���'g-9',P3*�� +�������'٪��1�I(t{L�H��^p���'K4H ���R��t�ٺ0&D��'��xd�Sі�D�)-1�Щ
�'(R<��KQ!5� �Yd�['�ڼ!�'�v�C�^K�Y�#
��J޼u0�'8��@�����B �3YP�\�'�:Q�R Cc)l�s�eR�~��ah�'�> �v����TB��ݬHh>��'��L�W'̔v	�Y�!-H	B�J�
�'rDY�g�'F�F�"��M?Kz�K�':Jܹg�2P�ƴ�`OT76���'��a �+ؕb�H�{��^� �f�S�'�<����Nz���ÁF"88��'O�XF$�,1��3�ȍh|�	�'W& qqeO�[��a�o�;Y"P	�'ŴP��H�0Y�X,ٵ�O��U��'�T=�t��\~�au,��'c����'I�Dʥ�C�Q(����&����'Ӟ�)'D�j{-���,5hl���#�޸��6.5��i�,�=^26�� �i���M1LuvQ�ĥ:@��g[\�8v	�V���W�^�{W����zy�$bW��1˸0��'̦Bܪ�%��D{��D�@wI���V* �W# ���Y��y�e�S����C��V��Y����'jaz�i�i��(�%h�*R�� )CD��yB�� YJ$1a�0H�r������y
� |���.%F��cǒ�
����Gp������*jÏ�P���.Ӕ��2gO$�yr��/��<x�(ݐ'"T�b�N �~��'Z�T�4Jߙ^�f1���@1F#T<;�'�9(�Au�ؕ#f�[�8@y��'�JIx`���|!!��^#0�dI
�'4V�H2��>|����� �~�(�@�'KrXQ��b�����)V6q1��
�'�2�x��gq�!�6ab��B�'��E�lDJw��#�çZ���R�'7��KS�D�~PX�P袘b�'���w��$3����S&JC�y��'�D��^�]�T\�m�7�]��'ۂ0[4f�>o��zu��DāO���I�S�P2���$��i�L߸B8��􄨟�EZ���FB3t���[κ )|)��=D����*K����x�bO78�Ju�O)D��J�ǁIV��A̻R�>]�` <D�S%5m����oL�4r����,D�D���/�ƌБ��/K�4a�c�.�d5�Sܧr�D�FC�m�=�U�.ڒ��x$����U�i^X�BG	�X=jd�ȓ)n@� �2z�0X��W�4�ȓq��X�s��� � 1�,�
����nZ�)� �~�8�h`�/�h��#�^̚5`@�,$�9c�I���ȓ� �z .���aSJ`�~�Iy����P�Y�!�e�H�B�(�5q�H�X�6D����Ó;<\Աh���O�D�pd7D��#I̩Mͦmy�$	9r�4��Ad5�O"O|��� ]�+�> ��Z�[p:D�g"O��a ���'�!Vj��@�"O�T�t���~�.�pw�9w~^�y�Y�$F{��	��{=0�I��B�Qr����]��ў4�ቌ�Q�s�<[�#�]�#�.��hO�>�5���	f0}��I��~w@�a&�O�B���h���@L�L�}���^�@I��uX�4�<�U":W0���0�o���[��l��P�?��a�
.��ebQ��8_�,��� l�<	v��*��RSh6`=@!�m��hO1�����5,�f��Z)4N$�@"O�-�"V� ��!(�iV�����)4�S��y�AD�{�^�W?�:���j���yBL�n$4G�ˑ@�Ⱥ�-���y� �kI�a��_�=jԑ�4�٦�M��'��H�� K;@o|I�%P+7{J!:�'��ꐨX�.Y@�f��6�0y��dL8�h��<��F5VD�z�%��=d@Q1f"O�P����sĂ4Q�N��4/�y�oi�Fo�dr\��^�/�����Ye��3Rl"LHH���9*e}&���6�'\!�a���&�jb��E�r���X��$;�I���M�O�0⭓�+�iA�Tb���'.�I+���7V�2��? *��{�}�X��+�S�g�X�A�ŀ�2Q4i�qhG�{#=���T?)�L��Q�ₐ	=�BP��Ռ.��$%��)�g~�	�">k����K�g�����ē�p>	V��.7�0��kC,6o:�ôc�i؟\�\�� #�J�)8����&��i�ɇ�Idܓ�MF7�jUa��aJl��b^�'�r���)A9ST@겤�3a�>؋��Eo��	Ex�|�"�(!�аa�Up
`g�r��G{��W�,@C��=z����H�$����$D�(��j�9k��`�D?|�ã<�2
+�O� �y��AXj=���Y���u{"OJ2
�b�� ���;Mh�Pf���G{����'��U�R�/odh��� 턄I
�'K� �\?C~U��K�|@ ��y�'�`��ʅ�;b����0���@
�'>�����֫3N��!'�Ux1ts	�'�8+�"ۂ�5�UJA�jO��y�\��E{�O�-��f�6_V����L�q�z!`H>q�'��iRDh��L��'Xԍ��%�¦��t�)�'�a ��"&T}j�@�&�d$��	u�S�(ScM"w��c�e/SƊI��|��X#�JЗ
bJ��D��+T���Gx��)Zc�_��p�wdY2kΤXr��v�<!�E�-m�0I�U~8� UC��hO?牙nh.dB��� �F��D�D|�p����>�� T.U<a$lX�J;���Ä]�>n!��̋G����R����P,Q=azb�FY�sy�☻#h�0`�6Y�dQ�ȓEŬ0f ��*pNIR
�.-M�9��.x*0�JJ1?�!J��F,R�,�lQ�����v��'N�X���ǿ1G�@�j_+�y^3�:�c�i����E��y���P�bRⅹ;����ޒ�(Or��$ӎy}RI;b�	L�Lhdf[";�!��é:��q3#B�o�dm�gkA2w!��+2z. �C�;�E� k�	rƱO��h�}3Ǎw�D���݄��PZ�	�i�<yv�Ȝ�,�#�B�g_�@����h�<iV�F��1i �QS�Lҗ�^�<qEc7$��kT`�;H�d,{���]~b�o�O�����K�?�4Թ��a��!a
�'̈́�I�D�߮	3�F=]�΄H�'%ў"~��
_�L�.�1�J�-6��B&�L�<�7���xl�g ވ*W��A�RJ�<��EܶH�z�sBsǮH��j�<��eٺb�(�Q,T0 ��˳ɂh�<9�GȐ+㤤�g�5b0l�Ѩ�a}R�'cJ\��
χ-26�{�(�3%����'be�@�Q���+e�D<&���'(|Pv�V�{+L�*�d�9k���,�'z08�	#K���1�߯l<�����`�i�-J��Đ��D*n`�aG{��O���R@ ;r��l�![@Vh��'�v���`%I۠kN�W��\*�K�O
��G��o�6i����Po�l�����&��!�Ĕ4�܍������ڡ%���IS��(��(��i��-�����-�E%�"O�n�|�`aP2  C*�Ԩ`�x�G&�O	�0��+O��Ѓ%A�6��A�'��Γ{�!�U-��F)^P`鎧9�����5>����s��q���&"���Gz�i6f�~�Vo�Y�r�3 ��9��4��	�t�<ᱪS�#��؉FMR�h�G-�?yq��s���
�XA��a&�
:Ѯ@ǥ6D�葂ǂ-G�U�E�0 ���!��4D���W�H:@Z���m�1V��a��%D�ljC�Ub�����͡:PT��
%D��
��_U]"8(��ǜ3�,�X�n0D�T��]�͈e8�̅�U��]x�O0D�0��FB�� a�h�4���h�-D�t�E��_����������R$+D�D���!'պ�!��WPV!I#�'D�(y� �4@�x���M|HK��'D�R�+m�Н� ]6��i���3D�� �A�W��&O@r4r��D�R�5��"O��)B(�V���$�|���"O�L�s�(H � ����0�6"O4��W(Ȅ~�z���OB�R��)�"O�{�$H�W�% ��>�>�"�"O�l� ���keNΎyyX�Y%"O�(q
��C�:iۆ̔�Yh�e��"O�,�PΛ.y��*��/N%�3"Of��R`ސ:��Xg��_�H�"O��Cd <o;�K���b,2=�"O��;���W/�h*�%<P��"Ol:vG+H�p�[+�$ ����"O��n��2���7�IA��"O0��(D�~4�m:�@K�A
d��A"O<L�_����#-�@6"O$���X	dZ�3���7��@"O�Y����Ti�	XV'���e�"O<E@�ا&-�g��-^l-r"Op7��56<�%F�QL��Y�3D�d�B�l�"U���qEn��&%&D��q��Dp���@0u���D�%D�4!4�Ԁ�X�h f��,��!y��$D�Xtg_Ҭ����j��YK�� D��q�m�Z�8�g�\���i`�:D�PH$)�0	X)x��#V�ȹ2D��8��;^��;�"�be>ɡEM<D��`-�%��䲆gI		�;�:D����d0 +���(�+q����;D��c�,�.o�lЉ7$̥0�F�"��9D�D��GN0(̌� ��%��:D���f.Z7}��e��ܕ���1M8D�LZGd�p���e�ڄw�a@g�6D�i��+����%�Y�v���"D���P�������q@,��0$5D�t��19�p�q,��@!�y)�<D� s�IݴW�AH'a�c��)�� D�q3i��Mr9���ߌ^��	�e!D��*��/\Z����J������<D� ��j�����^��r$l:D�Ȓ�z%)P��[�N�Fh��拟�yr��&�v�qd�imr���*�y�#���4=���P�\Z�I����yb*�I�d�@�.W/�U�����y��"{�`	D��6Zq���W��y��x��c!ҩ<]9rl�Z�<ɀG�)֬t���6X�H���M�<qR��J@R8�c��2�"i"�e
E�<@�����ǖ�(�|!��	F�<�AT�}B���'À)�J��N�Y�<���_<��X��ƽ2�� �[W�<�cH�
a�1
���A�4�QPIw�<y���2C��Qpč73�^�A���l�<95��:1 \|�R߬R�H��@n�<i�������Q��/�����!�k�<�`KOܭ�"�M�l뺄�g�W`�<���
��Т`P$y��i�̕b�<�a͝w1�UB$��/��Z��@{�<�]36���³'���� BLs�<a��>Q��₍F&54 Y��EBn�<16� |� Q!�m'i,ܒ1��R�<�we@���L�w#O8r������NT�<&\��!c7%�gʖ��'�W�<a6kǘzzla�G�w��܊@�N�<�F*�;�6����Q�J4��!WH�<� ir���:�-�� �4Ql��1"OJ鵠H�����Zl>L�"O4����r�����R$P�qX"O �b��K�,��K��yD���"O�i@�g�O{��C,#I2�k�"ON`@�AM4��z�@�"z8j�7"Oh��#���p�$D�+���B�"OlpbpG��@���f�ξ�<Hz1"O��j��8 @�ZQb�?�L�;�"O
(�`�,u�����ġ=	�`0"O$YA��)H�k��I+N� }�6�'�舉���g.a|2�M< �����ϵg�`Pb�d ��=��W�Hɒ�! @�O �V@Y/W���I���0��Mz�"O��c^#� �5j�J��a7��%K¬�5�׍�"}*W7$��i�)ɩt�Ti���c8��J�)�S}"�E�A�=�b��I:.}���Q<�H�J��ݑ(�ʓF	��|�'Șk��'M���,G?	��#��ޣy�$�!��iN	a\���+P
9��4jV�K�m��8���"n�����c؞h�`$W�N"���J�5�<���N�Ld����~�����3�$��A���M�����+�r�`7h͌C��tS0�`�<I��D�G��8(#I�X�tT!���<Yt�K 7�,7��)n�m�R��
�S�.|y��"FH:xx���gK�	�P���G�:P�QX�'قY�Oڜp,:����.��jm�H���9��<I�j!�gy��J�X?�`�w'á��	���+�O�I�푔�ȟ��h$]���1�E7������4G�iqh�"RZ��$A3������	?-&��7kE�v]<�
I�S�i�(���rAM��D��#OZ�X5��@B�+َy���S�<9���
�T�Q�퇊	ٴ9��!�D��'W<l�@�I�Y��F�T#Y/C�|���q4�,����'<�!l�J�Ş.|���2O�#����P0�Dp�/� ��9?��ŏ�sX�#}�E�݆�0��$3[���jʣ]��i$���ʊb�g�E�GN�p��ɷo�z�rLڰ��ƢȨ��)�F�ԭPC�~r��:��!!
I0I$��qǄ�+}FEz0'����d�><OBQB@�H��lJ��}ڤ�R�ųb�Yp�O���FEV(�m H<ѷM��,D� `�<��K��rTM�Tq�$�[�'��Xa[�́@�+f��˲C$�8	�P P�� ΋g��'&� j�� ��AF����" �j`;Ed�"(��9�#Z2ʸ'���1�٤a0H2��F��蚜7�5S�
'⦜+�b��I���P�>)DE	����'n�=J���y�h�����0��t����"gq�}�1�Η�yiL����I#fWx�0�oP+7T�]��|������R�' %�C�,�J���W'M�pM8sO6:Ղ��Պ=di�D�x"�w6���)�ny򨍙y%���B�%J>:�S#�R���<�S��'O4.�c��ӟD�ֈ���M�"4����*F�bH �h���ēT�����jP�Rp������$��P�5�L-M���q�ɕ/J�q4LK�9Ⱦ�x�*�5��Ob��c�*Z���x�a�	p	Y�&N?t��/
"�B��x2K�;>�4�%���,81釣
��<T��#��\a���=�h��,O<�I4� ��&Q�)
>}�`C�BF�L"��Ű>�D-ȓd�r%C�E������A=ь)��ְ'V��x�)��m5�'N�I��S$��I%MV��eǂ�%ؽ9���'wf,�󄂷-̕id,V%qj4E0r�Պ)@eJ��U�s�R�\�̠J�E@�ɼ@���Q���I�/rnr�ђ�FF�bC]��'~B�#�����Z'�F(^�1�~�Cs�FDs�i^�6�(�P�a^p�<�ۙJ<�)/֡�xA�g޳n����4@қ$�v�����r�����v��h�BU.D��Ȓ7�^X!�D R�e�B��D�J�9��6�1U!ٶ)^T��W��剋'�Ly�5B�+W�@8��co0��Č�i2����	�Q�H�Q�$J�p��7_�b�j�y�a/$��Ƞ��>e������L�H�PUM+�jX@px���0@��?	��7Q�ıu%C+)�9���"D�<ʳ-λh���R`�܉0����h�OഛF�*ʓO?�ᑉ�+[��8�R55P<l*D�q�'�j�
����{��(Z��US���Z�'�L9����c���iÇ�������'^����(�>Yv�V��:��N�a�<N��q$K�g�\2p�׵yHf�cW�;4�� p��3ǁ|�5��lQ9��d��xB�Y w4��mZ4���IP�� `��Sz��̮4_��b��O�
	{Dt؟��Ff^j� *�KʂpYE��
b0�yz�i�rxi��*�@ؤO?���"W�~&0�h�"=p����`�'�du��a�x��4��Ǖ
FS$�Q���y�|�'(Q�Tƀ�>C�5��	���杼YE�P{���2~+��{�S��e�,?qO�c╻qbX�<��- Q#.]\=��~�l�ɠ�=$�`��EJ�Lߨ���G�D,ҡ��%����F/���E�zU�ԫTm(���?j!$R
^�!�O�n��"@#D��$�zU M����7�:��a �O� ��ES��`���<�O��x⤎�*��r$U� �-�q���>�QDZ�XM��za"ZG��*���	8>np�'�9j$��	�%x@��C�>x�ay��(QD��b2f�zJP��F@��(O`ʃ��)S@ȴz&V�y�@'?�+�,d�:��	ӗF�1�ƚG����O�rXI���N|F�����%4���-j�-k'��h��'���
J����yWF[;G/�}8�	��y�h@@`�χ�yR��G����V��qr,���J���n`�H"'�G�{ʢ$�P�	�`�Ը���~�ء���-�&����
P.�U�Bl�d��負�8oG���WO�5F����&��	������&9���\;�-����d���?�LۢJb40�̆3�z�{@g9�I�52Y�`jF"�# Y��KY�+����y5*a�4Ȓ�[�R�qb"(k��H���J�:��UD�$ ����)Nx7.i�����O"���շL��!ցޖ%\x����'����,J�4T�xR��(�����Ѻ&����pCU�%�Z�J�Y��#BH��[����2v%�n�Q��d��K�P��.�,��0C	���� F�e��ם(Hz8̨���lȼȡ�Y�q�I�U�L�YǊ�9��S�0�Y3���T��H���&<r���UL�*���n�6	=i�c'˸Y�P��r��<�`�P�%;~���%�Վ*���S.`��@!�ν*�,'�<+�P<˧O!����P%�^�1�)S#!
D�aѰd�qj���W�*B��)K��Q&�J��i""X�B!�0�~R�6y.�=1�E� �� �?�p<��$GpR,@9[������3�.��U�&9�HZ�&�!)�N9�q�	\�pI��U�g�<��M�2�Q�ī��>�$kS�ޠs�Z]	aA5}�ؼD���bb*z��̳g�fo��$n��/(8���銽_.�� �2�
�SR�D+/�jܻ��[�
`.��$��!�8
U#�?��ɘ�C`钱9BH�U9�#,��>biyVΘ%�B��A�=��7��,/��睬jd�d��k��ziN*4�'8��B�	53CJ<�QL�Q8Bh��B�p��a�&�ǔ!@%�E#p�p7�]VhF �!��P:Ht�A��u���'U(�q�"ĝ�T��P��/��=�
�;����!г_
�;$勧7�D!W�P�i�lxf :��C#�ԦRu����-�	��J@�'��0�t	��0%������f���N>��ʎ�g��˖늒O���#s�jݡ���Y�3��������$����mB#6R��Ȇ�
BҩR��Na���"�⟔�F=���ߓ+'��Y�Bd�LIqʔ\��9�*@�:�b���@1���?�S��h�PjZ�0�$3��HG+PB��.f�`���9�D(�"B=w7.�䋆Y�x-���iP@���I�2�>O�9;ր����hAحb
A��"OL`Zm؝I�`yn/������>)���^7����ĸԞ� �B�Uc��>gF!�$�|�E���	�X�03��<=!��΁b�lE�Ԅr�"�ґ+��7E!�׾-D�E�P$��>��Թ�X)�!�$��(��ㅤ��2,�P�JרO�!�D�Gf�Aa'R�f|4�܉>�!򤈺�x"�Բh�����i�G�!��>��$�G�}�0U6�!�L=g�ڹ�6�B:dT��	 �V��!��ӁI�4���ê~6Ni�Ě�e�!��6 �^(��j�g�� �6��d�!�����tk��:ٴ1+^��!�d�?^�@�J� �����]�!�d�XW0�1�N���!YP��3�!�݀1�\�"��F���U!�$�,��A�j�2 ��W,�F3!��K�(���x7�	'��H�B�~�!��<!@ �9�bZ5Q�%���֛a!�P�V��Ց$�Y�7��qd J�y	!�� ޕq�E����w/҆ 
��W"OP�A*ֆc�|;���G�|�"O�|���S�bC.Su�C"|4�<C�"O��8����]~��7'��R8B��0"O4I��hA1+*l�������"OP����*l�l ����)>D�����
�=X2Ep��i� �Ά��!�D�?��Q�1�T�d4�x���0�!�ʒ%��� �2!l�C��*�!��H�j vbŕ���1�AN2k�!�$��!dXI� �6��� �Ş]�!�_�/�d���^�P���c�@�<s�!��X/�P���̎P�4US7m�VT!�dƃ,�$p��2R�b�+"��
d3!��ġ����I��[h�0"CD	5!�$O�1�� �C�)W�tDHf��:�!����T
p��R��9����m�!�M�8�̈�քD�8�T�̚$_�!���&NV���.��=�.L��MV�l�!�
|w ��!��?��k�M��
f!�dہo X����E�@��P+�I)l!�d��X�����(tٖ�y��W!��/v��؉�)�\k��a�Ǖ-Z!�*�Z�9��N9�Jd�%�9�!���@���� 
3�d���"�(�!��F�"�K��U�rś�>�!�$�"v*|�8�☟x��=�7���!�$��/L���t���A�rYG�U#N�!�$�/_�0Y�=:��%����!��ۯL�y� $Z� D`b�"�!���!�,ˀ�
�dܹ+$.�+�!�D�n$&���� D����-C�!�ۼ0��9�ĈZ�d�lx���+j!��D"j\�ٱͮv��@Ԃ�.%:!��gɤ�QrDpU­�N֝�!�G�ƨ��E�!�&Q3��|�C��*/��� �O�V��LYH��C�ɠ��8g��h_�4�$��X�&B�	w0v<�ra0}����@k�9�,B�Ig�t��iA�vu�����R��C�	?�NQ����xS�B���%t�C�I/x>T���  �~ȃ��s�bC�I N���t�ѩ`^��"_	:B�O�)����V��w�B�Ia��EOR�S�
�(2b�4s0B�ɤ#��hfH B`�)�Gl�m��C�Ɋ{�B��,��V��A�mK�M	�C�	!�(Q�M^.!��M��ƒ���C��;W�"P�A��}�}�ԁ¹<�C��&'���@#�,?H|sQ'��o��B䉝�"���lE�
�Z��7铩B��B�	�\���fI��=��/�~�fB�Ɋlt�q@���[������,^B�=^>p��s�ܛ^|���4IY/}m<B�	����Ӥ�5޺I���5C��C�	�XzF���l}�숕�T�N9�C��4$(�i�ͿuH��m�$v�C�	�T|��H�!"��ᆪ&^��B�)gޠbeg�aS� W�ވ9)�C�IA� 2���U��$��f��\��B䉿IH�li�n,#`��Ş�`�B�	���ا�'`���ދO��B�X9�0��i�!v"\�E��B�I�V��� �)`��p7��3��B�)� �ZW��<� �3$��m��ti"O$\;�fZj?�AkpVcZ�+�"O�<�š�<�����Գzl��"O*݃�L=4�T��� W�PK"O��_EA�p��#�0��p�K�H�<	d)C���A��؏�t �1 �^�<���P�t�Th0%�ʄ��\�Q�U]�<�Ӭ�6�L�a�Ъs�f	���v�<��'�-m�}Bҧء0����C�q�<�W��.y��&!s����4/�l�<���Jp-h�f#ŀ�H�m�<q�#���xЙSJΕ��@Q�n�<����Ҽmx����H�:�Z��Aj�<���`
��q�6E����`�8C�I;8�$(�.d����+d���@���RV�*�O��JG�P<J����s$�5f�n����'~����,��6R���ɦfdƝ�u�@<l*Ļ��ǎ[޼B�I%07"�#u!ǲ-�4츢E��4�X��b��J�$��A�\i�O#�l`T��d۶��O߇s�HiA�'o�E��h+R�zmY1G��k�n)r&�)�"�U�<���(�gy�jFP�Pݓ�'��(@ �����ybGȻ��02SA�jiVuV��v��S�) 5\ؒ�&5lO�����`�����׸#%<���'1z9��I�HHp�"�i��1[Ȅo ݠ�� ��B	�' Jm� L6�I��IN���p�y�E��}X��T���r��i# Ǫك.� X�n�2��<
p!�D[ <���W菋6-~����*RR�-����x����'�@QE�,O����7_�ɢBN�!�Part"OR�� LARJP����
�0��3Q.E,	�(���I�Ą�	�f�옃1��4H�X+E�	
�����@i��$�Aܹ�?�J�%E�<����`������Wn�<1��.n&�Ca�T�&���n��؈�EhN������c%	�;S�x�
_�T �o3��'<P(�$/]s�ŞɊ@�C b��)a��6F�@�D{����#R��D�4`�bd�HC�
�7e� 5m�D�!N>)�S(����I�K���#GDf�)�E���6m]�Z{�"����$������	U�A��ɇ�3B�n���ɳ�F�:PH	�.؍(s��ViF�i��D�<�J�)��xRh	1)r½@3j�~yB��,h�D�B������G��p>!�ǀPlPqSdKZ�ǈ,&"Q�vm��z�A8_��O�0aU��v�Və��)Y3�(0�C��NNP=Bd��[TqO)�gM��)�ʨ��a���,��VbX�z]��H1c�2�h���J��n ��'$��j�/4�3�D�~�U"���6=�8ҋT}:\��_�Uj�A�3OJ-���>���ӂ<�(Z����S����*��i�2�3� F~���D\�)��q��'[O
���@S@�4��r�ݶ\�dY�5$��~	0O�݊뉁]�t�*O,R�*E.OLDe�D����'N\C���@��=���A#�ua���w�B}��F�)����xR�M'V$����%`�O��|�%R"rvpI9�"樌�H>)�nA 갤�@-62](52w��F� ��tp4爆x���2&��?(�~�:�H(}B��{Z�c?O��pa�Jђ�9�0G�ʰŇ�
�d�ɚ`��s�̊Tp�剄
1#$�	Nlt�v�D~���f�ѲA嶅���'��LJ�#�O���l[�!�(v��61��AY�TĢ��p"QH�D�8��Q{w�$?�&	X�y�D�e M.-x<��֤�tx�L� �,(r,ݺ$��h������X�q�*�MٜO]��ZK�n��'��d��UW�S�'�T�7'Q�Z�1�� &��!�KE|2`��z�U�	յ_��T��e�\rݠҡ�;s!�ĉ�/�V�Jt�5H���A=S���(ԭBF �^Ϧm�'� �g~�N�f�ЕZg'�*�R4�g��>�y�eBڊ�&�9B� ׺iܶH�s�@��ܓ�I��R݅�IKD�h��H'=��3�ڨqh��L�h��M�e'��{��1MO c�pCҠ��{B�cŊ>$�(���J��}ڲ��Bv���,0�f� ���nO�r�<�?�z�c�IJ����ƾ&
p���3D��Xa����%i�%�\�vl�Q��O��Q�ޒW^p�O?=� Z�ag-
�rL�(�c͟0@�ݰ�"O
(Y��m��)y%��	�R9aF�>Y�
�<$����j_(Cc�@>*���2oI�9a~�����@���b��E���w�B:\%�}�'��D�E� l����D�a!�8���$R�!b� XV��~����~��A�Ҋhp`p�!g�<��̕=WTM� ˇ*����(����S�AT��d��>E�d�1ZaHլJ�L�2-�6N"@!�A6��lĴ¼���'�:I�I2�8�v�>�ay�A&)cҹY�H�Yp�=8b���>)2�,�H�B$�����DͺH�0xB�A�B�ɂ(���8��:Y�8ɺ׫ŃXyt�=����.k.V�;�6�S�x�<��kS�|��$�`�%D��g���Uۤ��Q.̕G�PXt��O�h5����LiL�"~�2js��!�L�4�h�e�1�C�I�{YL���)a#��I���˓>�����ǕtXJ��䌑d�ܨ�c�O�^׍�u�a~R��;db�4���ٴ5���1�
���f �f�񤟉'ǜ��f�'<Ƒ�W�,�Q��hR��k>0�DԿHl������17��1�n6D�\#�"���/^Bz��, D�HY�̛�(f��c$�`�bH)�l4D� +G
�&h�ѣ� �|�| �47D�h{��ݭ1(l���<��`���0D��b�E�x�TCI=ʒ���N14����ͮG2�"��^�Ж���n���j��'ZDM��F�	���SZ�5!
˓hZ%U��'��I�c�LĨ�&ہ]M���egB<BJ�B�I}��JV�;(��>4�6��A�>���«o,u"��F�}��Zv�-§5T|���գI�Ƚ��$�H�x�ȓ)능3A�`|pJuI�
Q�|���.غC��)��G T���P%�Fi�g��*��XK�T�� cU�U�TC�t{�	�e�08�\᳁ح�V��"���W���U=���.�XX��A��I�w,��8W��5!��Zag0Oڥ@vc��܊d�����DbC��0=r�ב)\}1c�Ү(�B�IY����2���� De��-U��'���J$]�L�Q��<P�m8��	�>�ݪD��~�,0���8{!��ҙ@�
���?=��=Hm�oF>�)$��\�N̓�ك6�扨���!��W'Q��P�NB�y���"��3d1���(^�)�3�_@n�i��Ijld��_#;�����-��hX�&,O6Kf˸jt�(���W/o��'���yv�î_�(�fB�g���j�X�imP����ϵ^�֔�Ag���x2��;��{���.(�n5{C����(�j=kc�%A��3�8U}\b?S��.��$wB��2p��s� %D�<�Y)�b����@�uݸ!#,���yRj���Jǝ|��I�![򵪇�ܧ�2��!�d�FH�#FD�c����ތi�6�z�	�-$LOf���h߳��-��X<F�i{%"O�	h��B(^�~�ˠ�J5�y��X�er�[�f\%���`g�4�y�(×^������Q*H�0e٢�y�jǺ[��d˂���L,�-�uD��y��0/�)��-B�J�%��HB��yB��~7,@���C��T ���y�k��-�xr1`�F��P��yR�١'�\����+�>Lcᛠ�yrJ�&���W�C���0j�/��yb)���*�&�Ye3���ǆ3�y��%��lw�)Z{\�`ץ.�y�F�<;����GWx�AG��1�yb�֗?���M�05��F�9�y���^�ʸZB,� AJ��y��#�y�Q;�,�9���=���K���yrI
�E"��`�]�J4J����y
� 䤠t�ɜj��x3Ѩ"P�@YC"O��0�ݤ ����/)	��'"OZ�0�L?t��ġ��V�Q��Mڐ"O\���H�Z-���e���0"O\�F [%"N��21�a�c"Ob��ǫ[�gQ����U(bM�5"O��ص�G�P��6J�"���R"Oh"u�LtRdz�ɒ-��0�"O�����x��Fj�<�U"O�P��a��t��'D[e��!�"O ����\ �@�7BFнh�"O:IJ�"��F]@X��C�(M\���v"O���n.2E��k`l�Ix�Z�"O$	�/gA����MU?<ȉ�"O��k����Tb�i �h
�%B6"O(�.8.�B��w����Գ�"OFAh�Axړ��6:u��%"O�D���ɉ��� �O�Z���P�"O����% �Q��عF��@)t"O:��fB�!�b�{J�	�
�"�"O��cb��Ÿ]c�@��h����"O&�zV"[y?��z7�>h��1j�"O,�ڒ����NH�2	���ہ"Oz аJ�M�J�z����\�`�p�"Op�sG�	>$�b�X�Y��y�A"O0����:m�@ŭ3� "O�5ZB���6D��Do^6t�0 $"O�-��M�%��&�RC:4�"O�x����2d���@�O�Q��"O�ѩ�-��e��4A�)�-!T�#�"O 8���S���0(H& Rz7"OXh�2�T:/�D�2e)C7P� �"O�lA$�ќd�yj����.L\9�"O�8���F� *L���O�o��5"Ot�
B��5<��h��x�@�"O�,�k@ &[�l1Ġ��r�8�"OnT��<z���dz�A��"O$0[����kk\�2��>N�Z���"O�QPD�V��l��]B�,��"OP`���ַ!z-�PN�6x��"O>�k#�{*!��F��'�x�'��)�3�?a�bL�.�4;���W�X�3�;�\�/(�<�G<��Iƌed!CR)^4�.8
�b�_1�IJ�(d�x�)ҧW0aU�г3�%Q�"^�D��p】V493!�8}���^�|ң��7���Z�hE�t�Y�吼=��q��<��F�C���>%>��c��g�����z��������Q�*��}��/�u> nF�+h����GX^��B��>I��,?3*�2��x�����f@�QHR="�d���~���(1M�W$#����w���� kq�0=+Bݙ��<yεXPmL2��O�����ʎ����K ^5V%�Q苲hzfe�B�M�#�BS�@�##}*��c>ՠ�� ft�K���m�8,����Yy�r��(�b9��1s�Yk1���)ta�u�'��Gy���%T�2V�7�a��牸i6�T�a/c�"On��(�(��@�91����f��Mղ�:�����O�aCe&2�$Q��ݞ3��}�-\>2��}4j2�$8|e���6H��j��G���|B��͘	; 1�F/�&Y�r�7�ɩ`Ў��C!P3i��i���蟾]��@�$��H���C8O��R�̛���C�	τh�8扡���b>1�ƈ��P�4R�Y�R��`�:D��;�K�6�̑��0�B��Ň8D���W�q~����hB�rZɻ�G5D�h�-LM����,#6�#U�?D���Q鑼&������2�%��!D�$:5Ȟ�;�,iQ�p>��� �9D��B"I6d���!HC�P��c:D�� �
P�+7^��Q��]t<�ȓ]�Z����H�U� �	_Ʈ5�ȓm��RBOM�B9XQ#b	ňiyTl�ȓ}���c�Cz�Wټ\ T"OA�e˃�):صSf�F�uؐh��"O�`���(�j�1�ЉP�<K"Ol�Z�L��:|��0@�b��T9b"O��$� �B]d�/ֆQ�|��"OLЧ*K%o`��PpH�*��PH�"On�:t��/�:)8�'�s���"O��4��rX5��'�%y�Fq�@"O%��NG*��E$0F���"O�퐔�D\y�V��=MV�� "OD(X@K׭L�	���^3�P{`"O��"��$lhu���
��a�f"O��%雀5�6LMTB�hD"OڨP�ZwԴC���(\�YQ�"O�H2�#3��uq`O�X
��"O�}"o�M�֬�&n̾�t��"Oܙ��:t
)�p~���f���y��I�j-��#fP�+H$�#�nU�y��ۭ9��)8BP&%�^ɓU�� �yrfB2[V���.� ��kb`��y�d
�5l���˷j��4#qm@��y򬕽EvP�S"�^"^}R {Њ��y��V��f,#��k�8�i����y��҇6��m��O^,b�Ktퟲ�y����9�@�K���h8����ۗ�y�#[�[��<	"�a}6y��d.�y�g�z	��ʰ��RDV�hrjנ�y��ýw�ك�H�?Kϸ!�a���y2���^�q�$iB/��(#!�A>�yR��4�桀��=�"�
�.���y��`�B��q�}�X�P��0�y�ɯU\����r;<�KЩ�;�yRO(8/�Y���vŃ�Ȗ�y�O�KFb���EѴ��\C�f\��y�o�:ٔ(ȶ�@"���y�I�lq��P�A�2�Ľ�anE�yB��<-�����A6_����1��y"��*yH� K��#]�T8�@��y"GU0i����k\"K���p���y��cA������EpĹ�@ʛ�y2䂙=���(G&��y;7l�y�[�z�!�v��vY@ᚅ P��y��h��=��e@�`�(���L�y� Jm`�,�T.áb��k��ک�y�cBu���*�L_ o;�86!�&�y2�@�<4d�xIE�gdh�pƗ��yBHʻ�M
�iP$x��U��y� Na�(eр�X���I�p옕�yR�0!t���ACzdP�����y��_�L`���>�P ��yB.�6�8t��D�9^���(p�o�<��닮7T-��B�z���$E	a�<��^�}2�I���t����}�<���ٯT<��4��:F�2��Z�<�Ɓ	�`e����- L�
��R�<a3lV�n�z��"��*%�y�<!t�HLF�����34�h �hJw�<����>u���D��E�\`�b�x�<��C��A.P	3%�c<����y�<�Ư���ƥ���%>Q��{�<QJ�;OA��`6iw����Lw�<� �Z�(�D1�5���$"}����"OL�KtDI E,*ez���;.QbD��"O�aQ�`�#8�쭈��ϋY/&�#"O�L)e��R�|�bf��p
j)�'"Op��2/9z=�%�#T�#"O|�cRI�/B�YR.E�~O��"O�{Ã\�_V�L���^�����"O���cFS�g
F-9"*��x�T"OvP2򄃀O:��
�l����b�"O�cC�^*78�m0�M�c����"OkT�@09�����ۛ
�ʑ�"OLui�j��g
���6^�,�"O�9�ۮ`Ңq�Ba�7t��ɒ"O�]��s{du��B��B�b�p"O�T��숼i�(��6���v����"Oȸ�,M���I`@D�"�Z�0v"O ���NN�H!��Ӑ`L�h��Ţ�"O
�+�/�6^oz��`\;\�L�e"O�@I5�W�V���u	�%uM�@�w"O�e8�����A0�Y�GB�h�"O�Ds)3,����ԈW�t76Hh5"O�`d�B����Hګk/R�(�"OJD�O26qH���5;�P30"O��ASe͆]������3"O��Q���(Ҁ{�Hӂ!����"O4H$�>%Ԙ�9q�� @4[�"O,Sdn�8/�2t{�gӜ�ti"O�I@çA9�`@1ᜁVL ���"O��RĊP:z-<� ���0i+0�se"O��N	RЬ�`���@�"O�-aB/DU8��ȡ�C���R"O()YŮZ�'�X��A�B,a:�"O�<豇P�Z]��Z�7J릸�1"O��ե��K�U��:	{ �a"O*e�A�TR�&͛M�6.�Lِ"O�}��ne.D�	;����"OD�{Q�̂L֖;�K̗?��"O��
a\4�hi�C�Ğv����"OJ�0�NF�
�40�]9X��	�"O�`����.6-�)�3f�'s��Z�"Od ���=H��s*@�J��"O*a� �в7!L��6��'�0�a�"O���@N�#��]��)_��p���"O�L{bJ�H�tU(�8G�~a2"O�ACZ<dgB��T��W��{�"O���E.���߹�tZD"O�( �CW]���:bʏ��y�"O4hZ��_2F+Q�ܑ)���"O\d��(IY:�C�+\�vYHe"OD�k���oR�)�½M t(�F"O@�@tk[�N��Pq��m�Ɖ��"Oz@�@\4���A�0	����%"OZ�(e���+��!=}*|Y�"O{��J25ex�x��\A"O���Z}�,Y*GZt=!�"ON@ t!:?���s���!2�P�"O��Ā�gH�t��d߫kBPC"O�1�D��5*֒E"��#r��"O(�G��
��A�,�S9J(b`"O�t��
�t HWa[ ��	G"O4��c�̑,a:Y�Ԁ�A����"O�kr�׳Qz�Sr�d����"O� ��T��bfEG?[����D"O�+�Eےq��i�� N�v�ے"O� �58p�Z�	S�J��ԂZ��s�"O�}�#U/Q��!bDt�pU��"O"�!���
! �F�K��8T�`"O@�˃LTD(��C��H�Rzl5ʰ"OLR���7F�6	�O�h�p�"O-��{
蝉&G�n| P�"Oν����[u��P�K��!�"O�E��叝7s �R��R>,��"O0Y�A@�W�	He
�"P��Lh"O��@U(��iI�Z�ƚ=�l\`'"O����W�W�^H�CE׮Ǻ��g"ON��C���`o��8�G���m��"O���&A�#����c�:]�� ��"O�(��/t~���U�Ͱ_6D�*f"O�q�a��s����*c����"O�*'+�;1UԽ;qj'S~r3"O������S�GK�Rd0��"Ol ���o������ �h֕"Oj� ��!@�P�ǮL
V,C�"O�he듅��MHR��\���"O|0��R�lN����M%I����"O����"V�&X���X</�)P0"O
�%��WƖ��V�.�2 "OPA���9*Rą����*6�"O�8ڣ���gȄ�bdC�	���yE"O�}����gx�=05C�&]:�"ON����r��H�t�W
&�.�q�"O���f�V�`S����F?�R���"O��c����Q��	��6]�2���"O��kt_�V�D-{@�H�ID���"O�����;3�E4��%6RёB"O�i2$�GD�f�:��
>$���"OxAbT��3��݊5*	8"��"Ozh�@O�9%g� kT(�� & }�"O\��1N�&$)i��琶*��X��"OJ����`�h������[6"O4��&��)������-j�ʡ#R"O�E�d���yb BG/�Aʔ"OJ�za�[2.�B�!�7c˺��C"ORM2���!>���!X�,�f���"O��TL�3*6�sw�ǥW�n��"Op]���L�,�,���+AX��q��"O��Bq+�)�B0x�J� %����"O��C�ɨfmDћ�	�C��z�"O8���;��A�JP5���R�"O�t��X�J��� ĢTt�"3�"Odu �� ~�l���+��|[�"O�y���\�*gH[1�[m���Z"O&`���
�&�ʆa
�j=@"O �j��Q����5��b��	;�"O���ϔ�Jɒ����f"O�՚1DX+x%8=�seϊ����"O��H��L�W[��[�D��D���"On�K�@�n����/c� ��"OX!����i4�?�0���CS�<	��
�(���F���t�<�1��-e2��̂��Cʗ7�^C�I0�d�cą~���� �2� C�I57ި{Ud?R�q���[��B�I�(ļ���*Ձ$U �"��Z�F�B�2_�}b�hV>"�'�" /&C䉛ZB�    ��   �  3  v  t  �)  5  U@  qK  �V  b  Ok  �q  Xy  �  ۅ  /�  r�  ��  ��  a�  ��  %�  ��  �  G�  ��  /�  p�  ��  �  ��  <�  ��  � �	 � � 0  �& - R3 ]7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6#\���<4�d5h��'�B�'���'	�'/�'�B�'���$��^] ��/U�Z�3��'m�'�r�'���'K��'r�'cظYA��4Z8�xg&�=�nܳ1�'�r�']�'���'l�'���'��41Cl֝wMƩ���0���4�'��'[��'D��'[b�'���'զ@�R��}�[�&���Ģ��'Z2�'�'���'x��'��'T��s�D
����c̚�	P�'V��'��'2�'��'���'X���EAO91�(��@�{�x=���'+R�'6"�'���'���'�R�'%l$�H^�C

��\�o��ص�'���'@��'���'��'��'��12����4��x�Rk��'n��'�2�'>��'r�'�2�'`P��6�.&M��;�	�:�d2R�'��'���'���'[��'���'��u��Ǎ
���z_��BT垲�?���?Q���?q��?����?���?��O�1^�����*J+Q4	zT#�?���?���?y��?a��?)��?i%��=�61Tg�y����ڟ�?)���?!��?Q��?��Px�V�',rl��~
I�"�m���rR"�U����?a/O1���,�MS�"��#5lQ� A��*���;Մ�!ct<�'�47�4�i>�֟Ђ@0TPq���.UM6E�0��P��-H�\nZT~�=����S���NxP1�u�֓��08)O�1O���<I��	�CV������*rAf-�n	0�m�&Z��b�D����yw���P6n5�
N9Cj� C�oK�/�b�'��d�>�|Re-V+�M��'dl$Pd�Q��H��G�w�̉�'L���ğ z��i>����1n���G^;P��"�'A"(~��~y2�|2�m�:Y� 4�
E3`�Ϗ/<*�i�!��A/��T�O����O ��G}�(��<>:5�Ӂ �E�$Q@���$�O�9FA׻-&1��	1�-&��3�����R+)l�麔��t�����O?�I�n�L�!��A�4�w��Q���I��Ms�,[~��{�����&&�ʥ�C�kxnEҔ��**��Iڟ`�	��ۡ���'��)��?�+W�H�%:^	Q���U�L�p�G�(^t�'��i>��	֟��	˟����~���X1e\�� ������r{D��'J6��U�r���Ob�D*������Uk3> ���h��!����OX�d�O�O1�� Ȧ�f�:U�Ӥ�T<�T�#ݧ� �8敟�t�8O��g�yy���_��'@$@ɦXM�C��']"�'�O�剮�M#Ső��?�ƮZ���@Ж�LK���xǊ��<��i��Op�'���'���C�;�pĨCk_4z�B$�wbӬ~�`0h��i����M��=��ݟ������V�TB�X�1
��v�.� `78���O���O���O���2�S������R+���s�
�$loM�������-�MPEơ��$Aͦ�&��uȇ�[����ʘ�2�X�&�O@�ʟL�i>�@���1�'|]�1E�_N
��!�TF\C�I	�nA�	�	,{�'G�i>U�I�@�IA;|�3� PMiT�M�}���	��'ł7͝�?(���O��d�|����-�L	bm��!���0S[~R��>�������I� 3eTlP�!�&2�؈W��N��R�ûi
�F�<ͧ
�t������1z(CS�^�
	�E�$b�//G�0)��?A��?q�S�'���¦�B���$�@����I����Ĉ�B��\��韈�ٴ��'Fv��?ɲ��U����:\�� �����?��~mc�4��d�9�X`��$oT"gp,�Q$���[��0C	��yRW���������ɟ��I�,�O���m-)�)@�R�Z��0�c�v�R�4��O����O������Iۦ�0-�E�"��;W$Dr�$J?1� �I���'�b>��3F�U��x=��^�;P�̳�n+<,�A͓Ij�1媟�$���'02�'Hy{ �̤;y�x'l�Hy����'+��'��R���ڴrd�����?��rsfq�&kƌD3l���[�iC���r�>����?�N>2��Hڰi�A�Qf���!c~�΃�=��� ��iF��v���'C"��()���� ^�29�yp�i��'0��'kr��՟�����6ly����J �0F����ش+ޕ2)O�Hl�[�ӼSSNQ*�-i��Y�M2�4�Si��<����?���:X���ڴ���� 4hs��� u��b��Q�p�#���� a8�H������O.���O����O���k��7�_SԘ��G�ʌw��ʓZ�F�ʳ*SB�'�r��22~:�: ���tу$�*P�,�'���'�ɧ�O�Az�$]�J���a�C�#���{�"\�w��E�<�ED׃����h��Ny���?�D�8QkQ�l��@��F��	��h�I��cy"�v�b���H�OF�b'̟+���`Tl��O�i�6O��n�X�y�����P��ɟ�Y�?,�J��3�L21��	�C�Aʨo�{~R&eb��jܧ��� |�Rѯ�0,��RE ��;KRJe;O8���O��d�O���O��?�A4랧��dAǃ�^�*lr�Aٟ`��ԟ�8ܴ!��;+O��oO�I3Xe�eK2b�z�z$�D1p�%� �Iԟ��#2�o�}~EV}�	PT��W�|)1��.4���b�^@?�J>�+O���O����O^!���a�h�Cb�"��*P��O �d�<���i,��x#�'��'��S'Cڎu�E�W%�j�e��x�p�E�������Iv�)�0�B�_Kl��������J���K@"?!��4����ߟ�i��|£]>T��h
q��ર�]1�'�B�'����X�й޴tjB ��ZVx��[�(6`�7�B�?y��!�����\b}�'�Q��#� ���-.�ieOÉQ��'u�1ص�ig���d��ן|�]����!	���P��r������D�O��d�O��Ol���|�tMX�b��|��+��@D�x���ץo�#POSb�'[��'��7=�ը它Tg���H>r��j�Oz�$!��i "6�l�x���ī]�Y�_�H�t�Z��U�iD�1��M7��OL��?���^�$�j�	_�RZ�ݚ䈇
�0�����?���?1+O��n��k�lm�Iٟ����VQ��!�p5�	bbC�30��?	!S����ş&����
��
H�cl�4Ry���F�5?I�r3�o��b>�;��'�Τ��:X.�|j@��Kr>q� ��8_�T���Iϟ���r�O��d]1�6l���G�G��ܙFW;,Br.d��@.@2���OڡoZx�Ӽ�p�Ϩ.��*�f�v9���IR�<�����$T&;@6--?i�M�i�.�I�(~b���[�{��e�Sf(Y^
Y�K>�+O����O^���O���OD����G"E7 �h������<AB�i�R�1T�'z�'��y�WH� �&"pKص0��9 u���?Y����S�'G-�TZ��%r��9e*�7@�Ȉ�6�;�y�'�$A�M埘�R�|�]���@<G�.���@�-�4`bu�\ޟt���T����ry�l�.P�p��O�EC� ��;�*�J�,��;P���O�o�E��"��I����	����@�s 
���:.�����@:K<%m�S~2K�
=2 �'��'��#&,��|�����'MJ_���W��<����?	���?����?	��������f#˄^�f9��D ���':�*q�*|�4�<�D�֦�&�|C�dI,E�NlÇ�H{��Ѓ���u�I�P�i>�	2�E�1�'��Y���u�`��'K ����V�e�����>|��'��i>y�����&2��Y�H?*z ���8H���ܟ��'��6\�u�����O�d�|RW�˩N6p)k�b��IrVh� AJ�$+�	����If�)*V���e���I�ć3,�����ڮcEH���EJh��W�� t�|⭛�^]n�XbAI�0{��9뗬���')"�'���T�X:�4#qr����!x�N=�2K�#4@-��-P�������?�2[�X��=n��������Y�GЊg;�]�'�s&�iH���Y_
����O~��'1��X6� 98���х�$4��R�'W�	ן���ݟ�	�<��h��J�7��C�OU�;�hbW!J�a�6-�LI����O2�5�9ObImzޕ�`��:ild��� M�Hw�իU�A��,�IJ�)�S� ��n�<)��N�{�u�N�0;J�	�<���[w���U����4���D�6Q��eR'!�/o� �JuO׮D�\�$�OJ���O˓@��)�?1��?�Emڣ6g�Xk@-�$~�yc �ը��'����?i����]�ԝ����OT�)å�[4b���'�� S���d�F5���ԃ�����'pd��!�)`��Q�Ŵi�H�A6`�O����O����O��}����������v~��a���S�����<'����6R>R�'�>6�/�iޥk%闒��h9�'�8f�zQ�cn�(������	�VZ��nZ]~Zw�z�g�O�~}k>v�b�� �L�@�[+:ɱL>�(O.���O��$�O����Oxd�ł.[F8P��K&Fz����<�³iF2t��'p�'��y��^�3�H\+�#��R nЯf����?Y���S�'oqH�3醉t��`f�ЃOC������2�z��'���i�Ο�`��|�S�L�����(�n����{���;g��џl����L����Fy��yӦ`:��O ���C�9x����U�)�B�O^EmZ`��R������⟼��`BKy��	�)A�2���C�bГ-��m�f~�͇A ,1��\�'���0JɘQi�@�(�%�����@�<��?���?���?!���g�&ṔVb�@O��(�Y�1~"�')"�Ӯ�"!��<	�i�'b�u:���8�����>CtP��|��'#�Ow�h3�i��j����
Zxh�`W;uS05 kѸh*R��G�Iyy�O��'�R��3D�������U��=��ߺ7���'��	*�M�^"�?���?I/�*�ac�M	�hs jY $��ظ5���ˮO���&�)�u�z��a@ۈ��ڗ>]����EĠ<���+O󩞔�?і'��
7f���3�
څ|��"���M����O����O���I�<�`�i ��)��M0s�&!ApF^�B��x��GB��ɳ�Mk��F�>A����D�(|����Y�,�)@Q��O$�$ľ}7�8?�D��$=��i*�� ����e�}*�AR��ٍ����1O2˓�?���?I��?�����iDA��as��qK��
�np��Lmډ"	̱������H��Ow��w��27f��ڪ0Z"��q��hh�'���|����X�v4O�t�� ��r�iI�p����7O)x��Ձ�?Yh!���<Q���?���D�V�%�)l8�h� #��?)��?����𦉣B�T�� ����+c�ߔsP��TE�.w2h�"Ǆ���������	n�Ɉu28�c�a#�����o����	�iB,:�&�XK~����O2���|���RI�C�l��7J��&� *���?���?����h���d�r�(t�� ��pW
�R%�|���ɦegˊ��4�ɉ�M��w���qv�Pe��u·q�B�a�'�R�'������F�����G\'Pj�iǎqʺ�9e�Q�M����o�.8gt�O��|R���?����?a��`��)��ɏ�s
y��������/O^�l+qܲ�������y�':��x��bA�1�KA�[���<ZD���'�R�'dɧ�O�}��(P�S�U���%%/���%����i�O\<�A�
�?��f �Ī<�!
��fY
�9� @�vAz���	�?����?a��?ͧ���ަ��ǄΟ|j�!�7?:<�]P$�0U�@�`b۴��'<���?����?��(W�=���2g�6)�)ȧ��	=�S�4���'6 ��'��O�և��q0$�t)(gGW�)��	ϓ�?���?a��?1����OH�I�e�D�`�g	$̎�*u�'<��'4�6X@����O��nL�I� |�0��X�;8q ��@�b����jy�&`����`��ϼTX�F�R���ʒ�U,\��¯����D�|�_�����������b�Ӫp���8OC�9��8�������IZy"�s�FUJé�O����Ol�'w����V-�7	������J/��=�'�n��?q���S��Mɽ=�
��˽U ^��g��0$ٔ��#�2F���<�'HϘ�IH�IP"M@Aú6u�x�aB�<���	T������)��yy҅b��t�SIB�g�B�ră��*H#��,#�,ʓ�&��D}��'�@����/JaK`���v)R�l���ঝ�'��%a�T�?�i1^�l��G��J�LA���ÚD�����b���'j2�'�b�'���'C哛� �‎�;I��iΠA��h�4	�~ua���?A����O' 7=�Zl�u㉜Yg�U���%MT��JĮ�O��D:��i�#7,6�d�x�SեP�����'=DT�ak{�X�����Mm�.��<�'�?��V4���j��^�$� �.8�?��?)����D	禡��ȟ(��֟�;�m@��TYs��1ꦮZ|���	ߟ���U�	��m� C�ۇ�\6�4�Ӏ�W��M�f��� n?��� ����
�kX�욕��^5����?���?Q���h���N�7�e�b �I�jy�0�p���$�����q�Q쟨�	4�M���w��0sE���o.��)uG��p߲P�'$��'u��	'�F����p˶L��1W�9�pg�
���4@P���4���<1��?9��?i���?��E�|ߚ��pa�1/F�����dJ˦��@ɗ��\�	��L�R��S0�9�&�&C��3�g�I����	\�)�S5lL�����$D�,���œC���Qs��̦��.O
�,̚�~"�|"V��zWG'r#�L�V7.K�5kD�쟰��Ο�	���`y��l��5��F�O�P��ː2��1�JCY����!&�O�m��(C����Iҟ$���C�<\���"�04��f�L/��@m�I~��3�����U�'ſ;���2P��f�v�2	g�D�<	��?���?����?���	�4��`�$��UL�H�/�)���'E��cӬ�+$5�������u$���.�?R�Y����)�b�怈_��ɟ��i>5	�KӦ5�'w8qv��i�:�p$k�8{�����B;�a�	G��'8�i>��	ߟ��I+ig����A4����5��P�.��	��'�67+Bv���OT��|v�Z՚��3X�2��FE~rm�>1��?QH>�O��W���" �뗫P
����Q�qf&�.����4��H�@b�O�!2DҼX{P��&':8�)0i�Ob��O����O1��˓Y�v�Q�S��s5*�{th,���:G��3��'���fӴ����O����@�(���yѲ���ݞ+�J���OƵ���pӀ�2J�}'>�,+�`ڷ�N#1C�%�r��F���	gy��'{��'�2�'Q�T>uY֪̿>��#�i,"w"Q��M{�k�'�?i���?�J~Γ盞w�Ɖ�k���6�����U}H�z��'��|��$�@f �V4O�T��H�I�
��f���k�a�6O ���R�?)��<�$�<ͧ�?9P 4)r�2�[�{&(�#Ì�?1��?�������ĦyJ�������֟�`�R1T;�|:����N�I�4j�N�;��Iџ|�	x�I6B0t�R/�N�D�g��v�,���0(�M�R��tAPE?a��8Mĸʣ� g�b(�&�LQ��?���?9��h�����(��yA�Z	%�X��vN�v3<���Ҧ�B���@�I��M���w�d���'�.���cH5��x��'�2�'7����'ӛ&���rA��&��� x���${��i�B
~��\;��7��<ͧ�?����?)��?wO��*�Ԥz�N�����dP�����ei�����<�I֟�%?-�ɂ2���j��F�%r��d�A&���2�O����O6�O1�44Ȗ/����p��[�S<�
'�7m�ky� �6G�(�����DB�^�t�zp�I��
Ւ�/��N�d�O���Oj�4��|��֠D�rr��&���KDQ;'�ԙ�G&�3u�aiӒ��B�O����O��$G$\Β�K7d�xMʜ+��
(��!�e��t@�������>��]6�6pBW�ܞ����Q�y��I矤���8��Ɵ��	Q�'[y�dB`$�u���ևZ�N\����?a�<s�V��+��	��M�K>I�`��E� �*҈I�.���S������?Q��|² V��M{�O1��S?�$x�G�k��(�]����?A�'���<ͧ�?1��?)[�� ��](�A�y�+��?!*Ot�nZ�x���џ���}�4�� n��ȟ�}�����с���D}�'�b�|ʟ\��H\� j��Cd,0]k"��bk���0��i>���' ��%��BCNؙ"͈�T�=CmJ49օ��0�I՟���ٟb>�'��6��3e�d|�
��RH�([�xiCf�<i��ia�O��'<"��)h��u��^Q����dB�5a���'m��Kt�iP��:v�����O��SXP#�#7.��(��!#�����O���O~�$�O��$�|r� I5;iN�� �dX��Ys�60�f�اu��'`���զ�ݠnnV�7n��Q�&DP@�W�
1j�IM�ŞTi���ߴ�y��Ϧ>?��QeS�n`��4�y��%[d�I\"�'_��ȟh��c�U��`�(��a�$�ȳz�^`��ٟ���ڟ��'.6M7L���$�O����*@��-[�>�.�&N�$�t�X��O*�$�O&�Ot��SIITI1 
2�D��G����bE�5؄s��/�S�5�r���4AR�r��9�D��2cL�j�cܟd��������|D���' ���f�dê��D�#��)��'#7m��D��ʓR�F�4�8�HB�T~�|Z�)O�L�jM)�4Od�$�O���ˤ= �6m)?��a�BE�'�XDA��E��C���� ֎�{��,�$�<!���?i���?i��?a�5D�ё�W�7R&A�į� ��D��]��,矠�	��$?牼���xr�_;B��� �3+i�Yq�O��$�O��O1�r��`�*u�z�6	��Ut�A�L�^Nf�����`
X�%��.o�[y�߮AƖ<��A	��\�%��	}�'^r�'��O��ɻ�MK ����?I #��&B.���٤ tDY��?)�i�O��'��'�c�9A[�)3�˒G�����,U{x�j%�il���T��7�O�q�v�.�����-e���X��&lR��Of�d�O��D�O���+��6P}�T��I�jh�v	şU~`�	���ɤ�M������ĦI&��;�ݘ8�h���>L�Z��N|�	Ο�i>��O̦]�'�N-B�@�!if=x2!�b��AW���I�'�'��i>i��̟d��ks�Ӑ����؂�ɾ��I����'�6mO5`����Oh��|RC�/;���6iG 7�4`��bFT~��>���?�K>�OO�xq��z�8��TÍ*K]@8�Ҥ���t.'|S���|�B��O�M�I>�6�� ��:�@O�o�2�(7E���?���?)��?�|�,O,�o}x�(���ͫ&o\� �D�7?`�������I��M����>������D+� �HVM+�,���?����M��O�)��	W��TT�*lB�K^.�$8�	�oM�Ģ<����?����?���?�+�V�Y��D�W@% ^!`7cԦ�Y��T����蟼$?��ɂ�MϻV;�Q(��TE�|`#��h���?�O>�|BTA���Mӟ'�tk�A�=!D&��''Y�3��:�'�Dݟ�8��|�T����T�E#ݭkzA{T
޶i�v��d��������H��Oyb��O���':r�'JlQk���?m�X�(� �P81@����g}��'d��|"��J@p4b0)�=i��b#��.��$R�S�6i�"�G�X01�m���]0��D�}Ԯ$ &���X����E
Rp��O�d�On��#�'�?Y���F��)�b�.L�ǃ9�?aֹiM�q�U�<Cٴ���yF%H�j�$wn����е�yR�'���'K l���i�����z�8Dݟj�kR��n�Z�@�Ҭ4�p(R�&�Ĳ<�'�?���?���?9��ai���˵|-� PԈ���Kئ5H� ��(���t$?牽=�\ Pv��
��
�6y�H��O(���O$�O1�rF��7:z�0��ˢP(�4��1{Z��)��<��c� z����<�����}QR-"�N.a⒩{��DU�&���O���O�4�"��:�$�Z�R�8�J a�t��E��Lܜ*^ u*�S���D D}"�'��I:!����˯1�qS�L�8�!�N��]�'	0�4��?��r����w&&���ƀ�de�uf�+r�UH�'��'0��'q�'��j�Kdg�&rT\�c�̚y8���O��$�O^DmZ�y�����8��4��M茜�Raȃ)��9Bc) �j�L>A��?�'����4��d:4�� 0l"rK@�E�	JA�	0DCP�s!o���~b�|rQ��ݟ��	˟�#�.��<�X\a҄	�����������Qy�hu�d��h�O���O�˧K�H갉��k���b�N�	�"��'����?I����S�g�&�2�c�曟f�l����!r&i��X���9�O�ɟ1�?�s�?�D&�ȶ�+@�T�ڥ��-q2����O~�$�O���<��i��D��7t/b\³�ҽ?��]Z�nY*@&��4�M�r�>I��{��5H�GC�X:v�Cmě�Ι����?!�P��M+�O��QR���JI?�cQD�?���3R�A�	uTS�mb�T�'X��'���'��'��� e� B7͂�{�<٠S��.#�.���4Hh]����?���䧘?�P��yWl�m#�q2R/�H�� l���2�'�ɧ�O0�BR�i��$��}͠�b��I� Y7�;[l�$),�� q��psz�O���|���8�Р�@�@��mS׆#��51���?����?�*OF�l�)0ߴE��֟��I�x�� F���M��Hd#��G^���?��X����h�a������=�h��䇝Q�j��'z���2���:�4�������ߟ�7�'/z�(�B��j��<k���G������'d�'���'g�>��I���"�78�t@ QJ�3�0���?�M��O����̦��?ͻ+1����'
r��I�(@�-4xd��?!���?I2�<�M��O^)���I����қ4�V5"4-x ���CG�(�O��|R��?���?��!�T[�L� F�ɉ�J�S
�(O��lZ)V���������c�S���{�e��
-asH�?�h 0To���d�O��D!��)�(Dʵ��b��O|U�eD�;.�� ��S�X�ʓ)Z���b�Ov��H>�*Op���B�|�XЉ����`@�O����O��$�O�)�<y$�iE�-9��'r��nH6 J�9B�E-$��� �'O�6M%�ɺ����O,��O�����U�B8Rs���1C��Rd�6m&?)n��g-��|2��q�ֵ"f�*dK�Q�V*�M�Iϓ�?����?���?�����Oۊ� ��D8&7�d���
������'���'�D6mA�N���$�M;L>i�OW7^
���c(V�1���ԋ�r̓�?�)ORY�rJa���uc�@�?g\F@�!eF��҈h�.�q���������Od���O�����s2�p�ˍ�~Bf)�Al�J���fT�hi۴:�<�9��?�����)�0e�l(�"�#f4f<J��$l��I�����OR��/��~j@�ȫS�MGM�!�$���$�<H���IB+O�2�~�|�.ȉ&`�ERv�C��f(������'�B�'<���[����4SVL�a�Õx�*�:SF��.]�o�$�?��d&�f��MI}"�'����[,.*<��i��o�P �7X�li����U�'�]�B��?��^��p䟏�����	4���ԋ`��'%B�'���'
B�'�S�o���q2���T�ܨ���Nr*�(ߴbJ�0s���?9���'�?q���y���!Q6�(���?.���L��;�b�'.ɧ�O�8Daһi��$���)�(L�Q$���@jJYS�Ȟ�� �	�4�O�ʓ�?	��8�aC�-o���k$��D�ʁi���?���?i-O28lZ0y6���	럄�I�/�TDh�̓�}](G�֯�P��?��S�D����&���6I�<Sfj5������".?a4�O=Oe�eڀ�n�'Hd��D���?a��o�ZA�Q<3�h���[��?)���?���?���i�O.��Q���j����ӌ�2g�౹���O��m�b$�ݖ'��7�-�iޅ��Ó	*�$5���-Is0� Mo���I�����gԒxnU~�KRL?BL��N.\K��;�x��W
.�e�L>�/O���O`��O��D�OT�IfM�v�Dl5	 �!�)�3��<Q�i :x(��'<��'!��y�%��3tAiC N�C��S�	՟g����?����ŞN�lI���(�h�(�BX%:��@[Ѡ�y�X5�'v�݀��柘j�|�S��"�A��dTb�O�g:�mb���柄�I��������Xy���j<q'�'���D�P�K9Ȕ�0dr�@�'7�'�	���D�O$��O�0"�ЍQ�<�D��-�0�C]?X�6�9?y��ON.���E����c%�6j��@�f�u�f�h��ɟt���4��������J'td�Bw�_�fЈ��^/�?����?Iõi��T�O?f�ڒO�`9�(�>\��zd��!S�ԁЩ)���O��4�4��h�8�Ӻ��Ȍ?	xA$�\vm�=bB�/�����A^�O����'"�t��!)_Le[�	Խ:1����$�ɉ�Yyr�'<��>�x�1�ۇew��QA��v�J�]��	П��	w�)���i�N!�b����BͻCc�$<���H��;m� �+O��6�?a�'�$��Ь����Q(�,��m$n!�$���9��@<<E\�	Ё�$Bִ���Ø�am
ԗ';7m-��'����O����["$r�"!/�]]ԥ���O���Uq��7�2?�;	Z���X]D�;�.P@��V�@2"�f;$<���D(|OB�ѷ3Z,�8 �I���3k	ަy�&`�dy��'���lz��A7�U�n�`�)��"��5�����t�I]�)�S5t�J!n�<� %:'��j�t��e͏�y�>HB8O�q{�jE��?�'�:�ĥ<�.O��ӉT��d��� �~��z��'�6-R@Y���O
����1#de8!�uB
8y� � 8�⟐گO��$�O�O ���P�d�d�����ʬp����噪v��oZ���]:����t��>(�rHXD�jU��k;D�( %�5+�S/p��d2�����ڴZą����?q5�i �O�ӣ5�d�y�����˒��(x��D�O����O��S�c��F�2� #��?]�&W' �k��T0	�D�c
�G��py��ɍU^Z���E����+2E����F�"����z�Za��XU��Q�c1�B�eB��؟���K�)�S�T��+��iڜ[�LF�)b8��$�CԐ�'���`���ӟ$QӞ|�Q��B���[��Y�n��f�l��*���؟�����Ly��~��u��O*(�A�7"ly�V
/'�$a�E��O`|oo�J��	�����ǟ���ό�sG��&S
�� �ޤ7"�<l�d~B�3{��G�$�w1�8��Z�0l���9~q�y�':b�'���'r�'�����%n�Y�gޠ�x���O���Ox�n��b��'��6m7���n�0E㈑ei����ǝg@��O����O�	�U�6m4?��k^� ��0R��^*����^�VC Hx���T%�8���4�'�r�'���3�?0zڴZV�J�4����':�T����4w�������?����iǤX���P�ߥZ��$��9��	���O��$.��?)��".H,� ��+�!B�ϲ8Q���L����D'Hk?	M>ieR|��Q!��~t�-@��X�?q���?��?�|�.OJ�mڸ)E&EY�+'�ҍI�AZ�P���%A�Ty�Le�~㟠I�O���1�����7+�tK�!��:}<�d�O���u�pӢ�E�~lЭ*�S�C\����Ԏ2ܹCש�"c)��IIy��'�r�'
��'��[>����зZK������cf�iaf����M����?i���?aM~z�ϛ�w�B��6Z*E��=�5K2
�k��'s�|����8- �v2O�����"~f� t
G�@�<�>Oh)��W��~��|�[��S֟��S��a8V`�!���gq�1s���<��럤��^yr ��`+�O�O����O�@�1O-|B"@� T�4ܺH[4)�I����O��$5��߰,m.�P���+[S���í��`����W�� �B.�⦱�|r�弟��	�!�b�!
�O�HHCǫ�'���I������D�	P�O�#W�6� P͖'s���5�B�8k�)d�hI��O����˦E�?ͻ������!��)����'-�&���?��?�ԦG�Mk�O"։�*� ��!{J`�U�%,�y�r��(K��&�|�����'���'���'QXI q�?`$}����h�i�PQ�,A�4�A���?a�����< ���H\�7N-8xH�(�Ss��ߟ��IK�)擂3+r}g(ʴ?tx��b�։>�Fp�5��Ӧm�'&��1�X�40�G*A dLB� �d�'��ex��иhT ��A�S��Ts�FJ XU�A� ;h����ׯ3p� 6��5���T�	�8�a3 
�l�ː�w ����D�=\ RU���_4�����@�(�cE�V� #�Ay��G�\X�?!�摋s���Tp�ɂK� ������!�S�J9�v�w��!�qJ���5��DPS��x���$�K���	�V#)������>G�D:��;J�1���R�'j�W��,�A�tcxӴTb���>f�5r%ЯVg�`:F!զ��' "�|��'���w��U�4,����ՙl� �g�%1��	���I����'P|L9�~:�4|�3�&ِ4� ����5;\�Һi��|�'�C��qOv��L��V��@V��+Τ����i|2�'��ɛt��}����$�O^��B08=�bM�.K=��`U`Ұ	�f4&�T����#�΍g����˒{��` �㇀E�!)D���MS*O���W/��m��ӟd���?�)�Ok�O�f���s� ������V���'q��x�җ|����:?xEQ�ΰ!��p���:>�F(ɐ(�l6��Of���O��iFM}bS���ԩ>��$˓�۸7�$���@2�M;��
���'�����Qy��}肫ߵi[X�qA�itT�n����I�P����8����<����~b�H�,U��a�#e
)b!MH,��'�.4
S�|r�'�2�' ��=X8\
��f�BEKB�p�6�<a��'��I���&�֘���豢��W*�@$�(*��(]�J>����?������Ņp.L1��nK�ú����*6�>�����s}�]�x�IS�I�|��e?��ǔI���lLPjf����IH�I��x��ݟܔ'��U�A(~>i��-��f�h97L�N"���$~Ӳ��?	H>q���?ɂ-�~rf�'F߂�c*���d�c����d�O����O�˓q��1�S?��'F�)��jç
�N��$��*�^��ٴ�?�M>��?�DL#��'��=4��<	jLBf�%�����4�?����Ѓ�N�O�R�'���_E�<H)�H%v��O,���O:�r�e+�	g�B��4��aۦN�?/�D�Ģ����'r���Ohӎ�$�O��D�nէ5V䄤8�.���FC�Ͳ�g�M����?�(4��'q�� ��g��5B�N��F�I����@�i`���s�
���O<���*m�'���1c�ޕ�@,E.@��i��猝<�l��ߴ���������O�bmC0x���	P%T�l4X���D.<��7�O����OP8���y}BU�4��G?�#�M�v2�a/nLH,+aFܦ�$��yw��ħ�?���?q�l���L;Q���/j\C��XD���'����u+-�4�>��6�����e#��|�W�L�T��$����R��ǟ �'���)�Q ��xhڹ�^�F���Z�P����Ɵ��?����~��\Nt�B���9y#f�I�C�M{f$VQ~��',��'��ɴaf�k�OV�ٳj_
8�RG� 5-�X��OP�d�O�OR��|��� {^q��M�G�����֪O�p��xR�'#��\JUT���'�xD��Q�~f!��ʙ�r���f�n�b�\�	ly%F�ēy�ڕʱƖ�HQt;��H���m��ؗ'F2nH=u��ȟ,���?��qR��k$ȉ��]6�š]�O �D�<i��\��u�E)Jr�-q�����,�L�h��'d�Ad,B�'�2�'��R�֝��L�����1+mJ��w%}Z�6��O��T�DxJ|�'��c� e��<�����٦�R@̎�M����?a���f�x�OL֤����#�J�R%�=���"k�v��O��5��?�9"L�DY��a��Đ�2�i���'5r&��^�)2I��!O��R��H��p���9N��O<t&>9����h��<�8�[b�.;!4��*�w-�D�ܴ�?��@�rى���'��'� �e��:�|m���Z�+��0�$�O��O��$�<��oAp8Ef�
ں9A'��w�����ǣ��D�O��$'�	�����\�6И��_�g�x��ɂ�m�e�bc����ky��'4� @ܟt�`�Q��ҕ�Y�w3��s�i���~���?�/O:�*6�iz�͓��*��J֫jdX�O<!����D�Oh�@a�|b��{2R�9e��+A
����,/���D�i��O&��<�Ee�S�ɏ7b\�����V���X��&b&6�O���<ٖ�E-�O�2��56É�7>a�a#[rt��3�oӯ�����O�d.�9O�N@�B��)j֣��~ʜ�J!����	�;�dٟ����$�I�?���u�͜�2m�@J�_� ��d�X�M����$�9��ݙ�ɀ;T/�9Б�*vfT9'�i�0�x�e����O��D��0��'T��*LL����#F�M�L$�.�)�b1ݴoh\��?a���?����'�� (�D#��h�)Ձq��隗`t�����O8�d�;@���'��ꟈ�P.��
� Xn�Jɪ��� /��en��� ������7�}��'�?i���?�V��<���")#B�dQh�M�,u����'\"�h��>/Oz��<��s��X�-Ԍ�{GۡAl|5���^}ң_�y��'���'^>�ɯH0�)W�v����0���I�# ��Ĭ<!������OZ���Ob5ibfM.q�P8�ƞw1��lW/@r���Oj���OH�D�O�ʓq���;�� P5������珵9H��r�i���ן��'���'^BM��yj��I���Vl~g-ۦ��%/k7�O����Ol�D�<�EE�G���؟�X �, h���W�L N6-�O"˓�?	��?!t!\�<)(���չx�6�aTO�O�^a{��U��M��?*OH����|���'���O��yc惛�f۶	��͗-�]j�΢>����?	��y �,���9O��3"�9�V��=Q�B��j�*(6ͻ<��)I2��V�'�B�'���i�>��H�)9��C�
�Bmj�'G��p�o���x�I�V#(�N�hܧ{>B�IE
� pW�ɳ�j����l84�J1 ش�?���?��'z��Zy�	?&p�Cd㗗,��u#�P6�I2��$�Oj�D�O��?=�I�x|�(s��R�x�l�)��3&|@�4�?���?�`&��s�IMy2�'����
F.���2iΜP��X�sQ�֘|�Kʚ�yʟ0�D�O���m�ԕ#gB��i�B2$IJtp�6��O|@#��h}�W�|��Sy���5��P�K�Hɐ%a�*4��%�1녷���S�X{���O���Ov���O�˓@�p�W�B�J�2�`�U<P�0�jG���	Qy��'�Iџ���ޟ��dR�,� 1�H�!�}�ФF�D�	ӟL���p�Iޟ4�'� �a�q>=h#k�	 ��A�g4�p�t˓�?9)Ov��O�d�}��	'@ёF��$=(���2����?���?�.O؀�0 ]d��P�ڼ���A"9[��9��͌gv����4�?�L>9���?a����?�I������k�P���+svI �Gq����Ovʓ{��Xq��$�'�����-D�`!��9�NQ�玓��6O���O�Q��(��`B����j�H�zʠr�����������Z���I�~����j����9QƔ�@/����U�!NP�lb�����O�p�t3O��O��>M�%���FDq0�'��i��PX"�~�>�Ũ_��I�X���?M<��ޚℭ��,^��)�e��Xf��!��i�8����'��'��B�$6Y=�i�e����s�"��vD(Pl�џ����ĊS���ē�?����~R�0r>%@s*�t6�*5
���MN>���OU��'"�� PAl��� 8�ڿcJ��ði�N���O���O�Ok1&�6��v���`ێ�j�$ �E�ɋ4*<�{y��' R�'��	+}"�C��Gv(�Xk��9!�rMa���ē�?������?��#W�#���-�Đ�Sc|�X�c�L&�?!)O����O8���<��O�=b��i��w�D�@g�
V#t�vڭZ��I��4��q�	��0�	�����:elʀ�G�2n���S,_j�Y�O����Oh�Ĩ<Q��V#w�O�꼮@ǒ�I��BL�s�!ȟ�f�'��'0r�'Y���'h�=Z:�iSa�]��ا"^k`t�o�� �	vyҎ�-u���������o��f�%���'��]c�KUb��㟐��Ob��	a��j��l϶7nj`���u<(�X5iۦ�'����d�P��O4��O&F�vN�Jȝ�F���G��f �Im�ɟ���a5t���y�	{ܧ_"����j�"�s�küO� m�)c�e�I�@��ן���ҟ���F�t�V�Zlq�U#B�e��
��/�6-�k��dE�EѦ�
����YD�B�Io/�� ��/D���á+R�%����l˰% v-�OvS��O�9f����p���
�'$p/*�YC�T�:�`拙�zJJ��6!��/0	a��l��)Jg%.d�����_�*Eh�#��%S4��L��D����D9xe2�"�'G�P�<H�5dMm$㖤�+kJ��eN��P t5�0�.W�mp�^�\�>9ѕ�\3�|9B�'�"�'��m��#�R�'��	ۀf�1;��ݎQ��8���dZj埅Q����'�#]���G�{�'��\�FƈO�(0�ʃ�����_�!�D����s���8���K� #?Q
 şT�� ��s�R���%A���.0�E{��5O<�)��چgΜÄ�	(F�B�	�K8��卅4^hf�b��Ԯ2ȼ�"���<�SJ�E��I����OF���w� r��DjΒx���9b�Ֆz"�'�R���/�ը�G9MZ���O�ӎ6��:�A%[a���
�J�T�<!6ϋ:X�D�CF�k(`�I|�2Þ*$���HS�I�'@ڶ�E�'�&X���?ي�$N������B�s�^<w���y��'N���T�5L�p{��K�b�n��z��'"��x�m�Nx���3Ǌ#X�:!��'�f�ȔG�>����ɕ�=c2�'B2�><��	$�3#�mp� ps�]b�΃�P,2Pqa�4��T>�|���������S��x�`��X��"�� y��]�	�.<.ٰ�S��?�a�w�@QQ��Ǒ��t[3[�faz��?��O�O(�'�b�k�]$�B�;
���Y��'�����oI�M�E(�����T�����f�����0�"�@H0�$�ip`�#z"���O�ppf
 �z8�$�O����O�կ;�?���79�!����<?������ZHx� P��mFI�`�#��M���|F|rB_*3��Z+� b+��-@�>H8�����/A�&u����R����O����/�x̓(<S�gO�
Nt4�e�G�.h)������@Y�lu�0���O����O��4�<} 0Γ�/؈+��Z#
�
q"��I�HO��0�t
a��0#1T�Yvբw���4o#��|b��~��y�;M����H����Q4�ٜ�R��ȓc- ��rlWhb�As�̱1�fl��Gǖ08Gʗ�R��!�D(IZL��B=���%�L�Y���M��@��<�,���gN������O�&��ȓr��١��D4EI��;:?�,�ȓ3$�(2���x2(Lbfb� 3�P���\�.Mȶ��.�v����y]���?#��q��ר^)�t�� ������A�й�LZ�f�y�"�9(y�ȓ:R�ͫ` K!V��Ƞ�Q*⨅�b�ܸ01.K�^���H%H.���@Rqqa���`vfG����ȓ�P� �
�2�^T�W
Nv��<��k�La�עȫ"fn$�p�L�N����=�Ze[�,�&��I�%
�a�ʀ�ȓ.͌����z�8���N�H�q�ȓa��p$Ν$\�*@y���ҙ�ȓ5����F�ۜ3ThꐁX�Rt8���V����dcD�G�b����	-c�@]�ȓZu����jĶ) �$&0|��ȓ_�:�bR�"m��ͫ��!l�E��O��H�������) �R�J���U��t{p˓&Z�!R��(��!��S�? *a�A�;0�1�,�:q�"Or`��+*�h�6�O�B�,��"O���⇘9D�
5)�3C��p%"O~բ��BVh@�״f)��r"O���dʺfj �Uȃb%�"O|�b'�ъ=QYQ���%����"O&��'/���d��F�YS�"O!�5���	�.i�6�߭�R�:�"O�hp��^;�|�� C		8�5�Q"O��D)�x}r���Y8?TBQ��"OTX�G]ׂ� @<N24Ӂ"Oڑ�+=~�P�Pn�@<�Z�"O8Ա�Μ	��ИE���/4��"O�c�)G�;�Z�� ̒K�t�"O���BM>���ն
�<��"O�PZ�nפ^�y�����`"O<Ѧ�I?\����&\�tCc"O����,�	~�Μ���ҳn_.�0"O Y��"%p�	�,�z2��Z�<I��1y\2H�����:��XcaH�y�<��+,p�`̊��~��R�s�<I��2��Q2��Πz��H��e�<� �J�J��P��~²QQ���a�<i�O��NTݩ�ʟ�~���!7#�d�<�т \� ���dT�$4֑����d�<r��=̩�F��f�P��_�<�%'T7��L[Nɤ|
^!cuJ\�<�o>��},����BǑ&����p� �i��Do��y���U��'���Z� ߺ��Qa�q3t��T�|DS�d��A����~�Ā�ȓTД�[��Ovꊑ���S��	�ȓ
X�C�Յ�^5��aG���ȓX��:��
8��L��%܅ȓd*�աT�ɯJ* 0f�^)j�ȓe�h���-����g�E	����O��XP攟9w(��FX�\�hͅȓAQ������:��K�1sx��ȓߪ��� >b
r)�sC�i����ȓe����U�ʇv�j�
�'�v�T��qCX+��״t+N8$t�"ل�^N �k�l�j�X��
�2!�vh�ȓ,�vD h	�c��0t�-����ȓkfZ}K"N[+	h���^�<�ȓe��	2�S�X�*�3�N���n���`\����/h-d��e�W�q�����s6Ȕ�/��tA4�[�7�(��ȓ��� d��khDq4K��`h��"J��s�#lC�0c�7Enp�ȓV���+��X1����.Ѫ9 }�ȓ	��e��'n���%�Y&c�$������YS�� ���ԡ] ~l���P~�L@��-,`��萨C6cN�D��?�:,�l�،x��2kxF}�ȓc.^)���@�����,՞��ȓGx�8n�=�Q"��"	�����qWk�9K���֠U	�2)�ȓl�0��剎��l���'�K��0�ȓ?G�Pb�J�q��
Ph��o.|݆ʓ�`�deO�i�(�r+�.%� B�I9M��+%kT>xqtp���;(��C�I}�j�k'o�o|kVi�{,C�	�~Q�lA�����#0�ե�C�I,w���wB�;?v9j�K�8R�C�)� Rm�ϝu�"��B6ӠtP"O�Z�,�-���F�Π���Zt�'>�q���­��
�48&�&a\$�v��d^9R�!�:M+V9#�G�ws���ℏ6�qO�`J��FH �?����('GЍZ���1I�H',0D�L#6�(5�ެq���������6f{0��<�;�gy�*U�md�����xYPwm§�y⮓ z�A�&HV1�֬�V�*)ৡN e�}�Oߊh�^4 S�~��SFl
3�p=���ެcτ1�'֞V̖4F�uJ'(��=^=�c!?D�؋g.��3:�<�F(N�y0��C<�ɾ���a��?�'wi�ԉ�jm�>`c�(]	G\Y��&D�>�	;irI���R;&�K&$ K�� �T?T@a5c3�	��II0^��P=#�k-���9��M��|�;2�M�W�B�I�VHB@sa��I�X�;�i" x�'��j��6�@�J�Y((���|��B�;h<����ӍLR١�M�<���ɼN��Zu���HD�`�=Ξ�9��W�,�]ɖ��|�<)�e'A����)�R�:0(rBK<)�i�.͂��P��69T��gJ��Y�ص�T �j}��*K�=&�����f���h@'	�!l�{�
��1�ax��\3Z���gǙ3����Cm�Bm�U�Q&�}�n}ˠ�٭SH���'�|h�!יc���ۇ�ݣGp֔+�Oܴб	�'O`�j�&�=- �8���[vvM�РD�D���PG�A|!�FUz�����ƺx��ёjY�f��E#k�Il��S��(}iTi@��$N���" �V�<SlH�oD	�!�$V�u�4��TB�v�����+D�z�1�J�	+���)1&�;B��ۓ1�Wa��,.�I� ^x����$��jÄdr�P:dq��Q3G�8J
�qr@ž|�ڴ���V�w �A�"O�tZB�@#6�����]8,��u2����;�Ǎ��\��bO���j��S�y��$��GÆSDl����x�>٧ON�NsQ>Y���*wpL�C�`��~4�j$ܡe��p�T4��i�1M�V�Bb>� m�/����l �V����Op\�H�7㸧���0��+��	QDD�&��*���#��qĀ�0��k� 1lOУ���t]<yƪф!��L�f�>9r�T�K���̶5�~���tq��:��
%;�~��O4��¦�v�z�!�1��\�P�~�<����9���.�Y��a�Sz�'�ܩD�-§g9��@gݹa�@M&{�=�ȓ9�RXjVƄ�<}�`#�(����� ��l�rD5~Rt*�)�s@��ȓPp<]�Bk��� ".-����|E��ʦ�A�i| ؐ N��E.L���rfvaH7�(du(����B.�l��ȓV޼���	�n�,ؗ��
3L��ȓiH�
V$�;]�4�j8Ԩ�ȓj�� Q�B	�xduj\�$�-�ȓ(T$d{#��wB�h�.��Ő�ȓ����(E�'�F98c�n�6�ȓ-���C�V�l�"��L�Ao�y��{��2̑���Y�F݄��\��>؆Yy��Vi��Yj�?M�����3�����B�8s���;Zv�ц�#�B����\ ���5�Y����8��8���O�ѐ�FĜ=����ȓn�n��f$|���E��F�֔�� �����8Xx�M�����vR(|��<����-�u��kK!:E�ȓ	Kf�h��%4:֤k�,���ȅȓ=_�}{�U�?m�����J�H^���ȓ_t�1gOJ(:NH:G�W�"�,�ȓ&�A�Z�a4�	ZQ��=NބP��(~`p&�L\�J$	�R] ���W��� X@� 	 ��0��)��L&��p�XHDSУ�6bɄ�S�? �2bm) � �懰pX8�B�"Oڐ�#@�)�h�ȅcH�1���@"O>� ���O4bL)�ʪ/�Yr"O܉���L�+���1�/���Rt"O�)1`Ə����c��ј��L�"OL%��Ӓ%��-B���\�^H%"O&젲�΂Z�HhȠ�B�J���+0"O|���1G^1����/WxD`6"O~�J&E,p��mЀW<����"O��*�әo�P�P�6.!�A�"OX���Z�vD�7'�*f ;�"O��P�)D�ȅ �CM5��*�"OhH؁�¥*7�]�c�:rSbeR"O*}&�ۣr>�a���CJ�ib"O�	�T�p��Å"�\��:�"O��2T�$6���� ��V���4"O�T���\93�poÚv=�l�"O��c��L�kX,�i�Z<��mCa"O8h���8�����N��5�j��@"OBU�� �!W��+�"`֗?�yr$P�wþ9���$)���� !�|��NLRH҇�P{��U�4-�6�x��H�p,�E@� J.�=� �e�r�ȓ.9���F �$Y2�f؃Tk�4�ȓQi��RF�t�l�8 �PV�݅�i����ƌׅ[Ȫ�{�N'V�ȓj~N�K�--*�A���Ů9���ȓJc&%#��BG�{ͤͲ�F�S�<!v�Ǟ_�|)���,E��) �[M�<����U�T�3�P�)a�[S�<�R�\�,�T|�싊�h����e�<�6ˉ�3�����j$�`qb��]�<Q!@��RQ��șo��0�MZ�<�"/�$/��1C ��;o��� 4Ʌ|�<QF�'A<nt'!�5�Xx�1�Gb�<�!�i�~pІ��O�5x���]�<��P�eԊlH`Bm�ȫ�5T���0c�4�� )��"`/����*D��b���_:��Q��7~u�-��m.D�CP�X�-��4Jg�i`t	�0�*D�0R��	3:��y8�Zr�8�C�b-D��B�ލXX�l8!gra(�3F)D��fg]<Ԥ䳒%��VYfL�a�%D���̍�NNހ���@�n�`Hv(.D��a��F�����&�7�r�w�>D�P*$P4l�}�����Rt Ǐ)D�L�Ħ����J���4U��ѡ(D�H��8� m)��ԔQ^��2�2D���D��=.���Ff'{��5<D�P2!J���۴��?j]0?D�(Sf��$�ƭ ��YE<��ڔ
 D��R�L&R`��Z4n��9�|���1D���eh�]��h# �,\4���'0D��d@4j/~i� ��
g� �a�3D��p�,E9�h�X�A�E��	�b�#D��@� �<
L�	�;�ܡ��6D�tɱǎ!��Q�%�Q0E�l�s��5D�ػ�& �?4�$R��9F4쉰n8D��qw�Ɏ|�]�$#M[.`Ao7D�Ȓ��G  ��1֋
1֕6j4D�D�q�Ohw`��$��4a\��X&�0D���ׇ1�T}S`Ȭx���I3d9D���1I�$dy�r冄>.��� ,D���Z-j� 8���z�<�6�6D�� �@�v*�(fK�)�$B]i��4�"O�:;�D!�@ݢY��b"OL kO&�B �t��,��"O��Hdg��[�t�͗�?��R%"O�8У��0U���̦h��H�"O�DQq����Ex�oʪ�M��"O6+&b�v�Fl�3��'}K4"O���ղ*4�j���`L��!g��p�<Iaj@�/2�I!3�$z��)X��A�<�g�.m:���"�s`�5�d��A�<�
�5��\"7`�;6�{�F[b�<BªIE�U
�F�AO(��gG�<Q`���� (��5P޵��'�E�<鶈�  =��P�3g��BӀ@�<i�l�dD�Yb���Ft���T�<����i��k�
�/'�p���e�<�$�B�X��}.c��a�pMX�<1Eb�]�>�xP$�0a��c�n�<�'�M�����@ܒ��pi�gMC�<�&fX� �f�@�5�,�P�[i�<�!� H� �&/�;o��`lN�<9����pH`\�^Ԅ]�G
d�<Y���#ZXBA�c��.$��7�Yi�<U���a4�4�`+�WX ��B�I�<�C��]I XRhι&8��hSN�<�7&<^fF9ba�0o:������u�<�w�i�.����\d�=Q�KXt�<�����'Ӑ�A�?(�1yBb�D�<����<}A���e_�0i��X�Hv�<�S/�&2��ꂫ� ("�X3eY�<�$�D��$�D�.��T`�D�_�<p!]2��A��&ҡFCz��F�d�<��b� ��E�a���[lމ�b-]w�<�g���,��EM�A���ТJIr�<)4�OV]�)��	A5s�|�P��W�<��k,���5�VSD��*�N�<ǫ��mU�u���Q�<�Z��El	V�<���Q� ���+�O���˕+�N�<q�(��C�g�'$O���1�A�<�d�2�x�Y�%Q�|0A���R�<������=�f�}�䰦A^F�<��_�|êp�"*� �`�z�<ѵ�J=N꘴����*��(���w�<��_�qXU&�"Թ�@�s�<E�-D������ 2c̭���_s�<9 B�2��X@@���9h�I�j^p�<!��K�Q �KR�����D�m�<���1l�����8C��h�<���K�f���h���%~�i��}�<1�Ò�V?�����9������Aw�<a�$�:I܈�"Sh8o���jbh z�<��K�#dzA�/�>="H
c��y�<�ù"v�q&��j����wϕA�<@ O�?�|I����-i��{WM-T�*�
�	g�T�1�I�U���X�;D���l�E�p=)1┉�~mp�J;T��S�,
<9��ʤK�����B"O�h6��5t=ؠ��p��8;�"O���cK
*1��(u P\��<�v"O���GF:�h��`��e�16"O&����4 ��Sa�·\x�i�s"O�Z�bN� p�5�H��2Z6�bs"O�����%�F�Y�;$�Iv"Ol��	Na
9r�ƍ2�\�w"O� ~A!J��P� �1�EU��l�%"O��Q6j��v���*�$2K���F"O:����!	�|(h��ğY`N�A"OFxQA�/�8I�Tj[�:4�Uر"O�l ˲
T|h�i͇�$�@���8LOJ]׎ NC��`�*��n��G"O��Hv��4-0�Lq�ʒ��L4�f"O<HHs��G� -I#ʌ�����d"O8h�᠉6~��M��H�<K�ґ��"OvL��,K���`�Ǌ	<��L�E"O�����bt��Ć�X,+�"O��1��ߵE�����I^�
��"Oh5y��Ή4�d,V�ܕS�^i��"O@qFQ{��G�X�pi�Q"O\r�"��8�ށb��jiU"OZuXtKD:F�(�{�*L?iެ�c7"OޤI�煑� A�ڋ'#ص�"O:�t#P62I)��*���	!"O��!�*9
�I�hW�%���"S"O��:� =s:��@'Q�m��t9"O�p�g����Eܯmd�4�5"O"Ĺ�e�Bh�8�s�lM�y�"O� ap�]$_�J��FC�v8��)�"OX���3�t�f�)*�xX����*�S�S����0�pq�r�Ç�B�	:GA
(е�ʑb����凞�~�B�	
���	CÌ&_�f�B���.O]pB䉊)�*�/�)]t����H�)rB�	����7��$k�~��@6O+ B�
HxIr��C(zlTғ�A:�(C�	'R��x3����-�E+�oӒ"C�ɼ_�>�C�D�P���T
�<+"�B�I�-�����/�3hd��.S�,��B�ɫ�dr헐؁�"�ѳV~B��j�Ұ� A~�D�͕INB�	�>E����:j��LM�8�'ў�?my3�A�[�x%��ʃ%N(�|�Ԣ"D�*�	�=KJ�c��BGB�Y@;D����f��p�Fm!��6Hn�)�E�8D�|�C$E�[�����%厁9��:D�8�wlHH��Z�W60m�����9D�$��FC3K��m C�K/8�H-D�tsbi	�<�`��������"$�*D�x�/���j-0g+8Qh���e3D��*�o��H�n���g*
��;��0D��x��ذ#"v$��4���`O/D�p�HO�X��.h�z�32�-D�p3�������5�780>�X��)D�dz�Ϫ-�.mpe�F��p��=D� �!��+o��l�����wPi D���ƅT".U���'��PR��<D��A �3�0z��%i�Px��l-D� ��_�15����
:h�V,8D�t�#gdL�`�S��F[ �Aee1D�#ƄY�D] h����XI���`�.D��YE�ұT� ���� 1���2D�Ġ
!
l��,�#ua�|c�$=D�����X6��{�
�2��<�dj:��q��|;�F�2����5ݢH����"D�,ѳLM-�VEb��f�� ���4D�����B�24�C�,�,E5���E&D�8)��^�t��R�Xz���I D���3�ۃO�p��7�J)b|��k��0D�$#��B1e���Qo�.����� /D�� ��-"�:]�B��X�m�"O�
`�1��=��n<0<� ��"O=*��Q+N�X-���� $x�e"Oܼ�ԍH��4A�"֝4{ĕ:F"O�)���Y�I�R�`Ýr⥳�"O}�Tl�[���bS"I�W����"O`4hVm^� ��ۅA��J�.5�"OxU���#5Tq{G�3b���"Op�r�ΐ�%��I ���L\p�d"Ot� .��_���aP�
�!�:�(R"Od9�o�-)��h:!ϙ���P��"O~9�1k�mb��5�K�`r��i�"OxD�2���R/pd��M�w��Q��"O.𹤩ӓ�.��P- &�0�"O��k���>�JI���Q8�T��""O�C!�R�[T�=����C�tM[�"O(|�`�
'2om�Rϋ�y�L�a"OD4�*�7ո-��'Y7�ȑ�"OD�r�R���n
0&Xɱ1"O�d�6�G3��)amGt �xR*O�X�'C�Z-.U�fB��:�>�b	�'���rӭE+:�\����b�r��'ۮ�QTd��	�U���	Ä�1
�'zxQ�cMY�D���T�.��'�N,���/~Qr=��(u���'g��(FOĮw�.Y�ƍ�k9�t��'�@�!�%]�!�a�,�4��r�'����d1�e���;���	�'qz�3�E�eb�]IQ+P/{N(���'�>|�G)+Ҳ)X�HTnc �A�'%,���(��[i��sbk�r� �'Z�%�W��#a֒����6����'|.�z��E�aЂ	a��X��'��-XE��A����r�ȧ"��=I�'x<���	o�Z��R�������'� �q"
["�$zbIZ'ı�'�0͐�A8�P]�@]0V�}�
�'�(�A�B\O�<�cA�؅#Q6��'+(��W͐P7h���OY�O`�'V��+r�L������ś��0��'pl �DM�8�jܺ�L�aT�`�'�hP�(� ,�g���'�lz�`ċX[n(B"؛��'��B�b'F�h���X�u�����'�`LKv��[���k�r��hY�'������0>gp�sK�i%�%��'�В��z��ia&��X��m��'%v�J@��<Y��1d@�F�B=�'�J����MT���#�.Y.��(�'h��7B��4���g�ߪ��'=\��� X8]��0�d�V��a.D��Y�+�R �:���Gbv����,D����\gVH��Ζ��9��(D��	��[�:�j�G�т9|��o'D����jǪ�\!y�F
���ԋ?D�x��N�4QpA�A�%~öy�o"D�<�DÉ�H����F#C�4��i�B,D���Q�[��ec&#�!C�
$µ->D���'M�&}>T9�G��Z�����/D���;�(�@��c��%�U +D��9�{��4`r�N)}*��3�'D��Q�S�lel��� �-F��:5k$D����,�����b+Ӻ]�~�`�!D�� P�fdܐ���O)��sg�#D�� �tZf��8�|�7��	�yA"O��ĤCq����Iq*IX"OqHA�Ðl�����*e@�=�0"O��q��
U���A��e�4tS�"O�4�#�H�������	s���d"OD��Fe��,l��ֈQ��yq�"Ox���E�%f����%W��,�"OdС�T�B -*`�
�&@W"O��ru�ڥh��<�RB��C��t�@"O@��b��`��HrJS�kqLT9�"O�<X��� ���`�F6LA^)�"On���%�0L�b��/]=*���"O�D���mܥ;�#ģ]/npq"OvM���c��a��b<(a�"O��1��	v��`���3%��"O�i��'*q�0�hݲs/r|�q"O��sσk$�Щ�'U�- = �"Olak�gK�v۸8X�]Y,bC"O�A�׽_� �kH�-��"O�w�?n2�ĢҪD�r�JtP"OX1�V�����/��0"O.�k���?�
):�̢||Fi�"O*4�RK�q:9r%=:����w"O�(���@,~�f8PA������ "O����ܻ��\�!e�|�nX��"O�+���E��9�e�~��"OQ�P�My�I��" �<��"O�q�+Ցb5`�����?t�ś�"O�I#�.�3NJ�勦�уg�Fey�"OB�E��T���X��նx���E"O�}ppJ�P� A;$)ڿ\��"O� ��!�"l=B��Gg�x�y�"O����.o5��bi[:Nj�˕"O�H���%��h�B+�&d���"O�d�&�O	$d�e	��MoT5"R"O*,;bg��w�j����S�`2���"O�I�FE�,a.�W 
2_W.˂"O 1�v�]1Q[��2��<lL�aB"O�H���-!�4!��-/&�µ"OԬꆇ�<\�d[(+ B���"O�`r��ܺ����m�HS"O8�A�>�B �"��0=���hD"O��'�C�ʼKgXzf�ؖ"O���w��*#���t!�OS;2"OH]�dDڊ9&��Q���:^���5"OZ)��ٖ�p�a 8n?`�A�"O�AC1�X�?�b=ڄ�D4�1�"O��� E7!�� �2k��B2"O��!�����p��aP7E@���"Ov��q�OG����-�g�a�"O~Ȩ��_�D~,AcI>Q���8�"O�!�l�z��ETOQ2��|�F"Ot`겏i��m(�.�&���P"O4\���+,�Yb.3:��"O&��F�˲=[�����v��(�"O���6�ʯ�@���[>k�0X�"O�e�RT8��(ar�_�{�"��A"O�t9!�;O�2�ƨ� T���Z"O���Ø�j�v}�P.Z&�H���"OJ�ʓ�/@��i��¥M����"O�4@��E<M�����բ�B���"ONH��nc�|H3�¢6$��3"O�<3 ��V�
c
����*�"O�9��C��!:ƌrUjݪS�as�"O� 2 �S�~�3ꅅO{�l;"O�MK �Ң��I�i=1BL�[�"O�Q�@Ҩj k1(�a4���"O����ō�^k�(��a�1PA�%"O>頰&Y	Z��ara�<[BTS�"O�k�.�	OD)S��Ұ
̌�T"O%!U�̇[Z�y �Ҁ@���"Ov�!eEG�De���'іr�H�3�"OD��B�]V�-[�f� ���"O���1ȝt�<��S;��;�"Od�%��&7��}bg�;��7"O܈A���^* �2�坃?MD���"O�|p'lãVh�ib'�-?Vr�"O"����X� ���_�D^>8R�"O�}hsX���P[G�Z|I"٘f"OZ�2����Ra�)qcdD�*���"O�D��5mPbV䒮o��`�"O9�!�h��"�T d��a"OX���a��^�XT�F'���ɳ"O$�c`Ƅ=�h0D�V2~�=�R"OfA���� zQ�Ҍ�Tȴ��5"Ol]:6MJC�8�W�W3�^��"O�`�df��jY(bd�F�0�x�"Od�!#�;3Ŭ]�b�(M�r�"OR��f&ϽTD(ys���3.xt`S�"Oج2�`�=r�l�` �nod-�p"O���%��b*Dq�b� iRj�¦"O>�zԫ/	@�����5m68�A�"O�`[b�+d����3�@�M,dq�"O�EZ�(`���R���	p�Q��"O �凇4_I��Ȥ\.�t"O��kdI�Bn�P�	\�N�F P�"ODX0�n	�b������ޔ�`��"Ol�G�V�!��\�w��x��+v"O�	����:��Sw皦PoL��7"O�ٚՌZ'�����4l��(�"O��kLB�l�j1"$R2M>В"O6��D*E�M��A�K=����"O��v�K87p���@Ӫ9�S�"O�T�D��\z��ׁ/\"�!�.�K�<!1�_u��[�J\�[2�I�CfVO�<�d��8�ҝ�%A���ܸZ��BQ�<�$��[⨱�Gƈ0L)iaLL�'a��g�2[�lH��.S�5� ����A-�y�@�oTT#��X�*x����$K�yRA����SK1ܪ��֯KY�<����+�ٸ�G�(c~�e���k�<�̏�P[�eن�E/0Gx]���k�<�%	�p���6Ŋ.1�y*� �d�<)C�Q04�p���莪j�4j��^�'0a�dj�=S��#+O�C���3���yb��z�읐�l�.7������^�yB戊1�ظD�E�"%���Z�y��Ƈvi��`	��oR��M��y��1�lh���ӑf[����@ó�yr�Mof�P�ʔk���`f�͝�y�f�9t:��Sgc����"g�y2�N�*I�gΊ�>4��h��y"n
�e'����"�t�X��F�yrK��J��3��Ghn `��펊�yB ё�F0��+D^��9�ϓ��ybFF�&��Q��g\S3� �%Y�y���S~0ܐG���� ��S+�y��R�^m�aY���Z���g���y
� <��ԆL�������
��%��"O��3�ˀx�6E�!U��N��""O����ԢlOfY�Q`F4��;2"Ol����\�����)�M���"O( ��e���Lt+1��VD�D"O��2dm�f�����] UAZq"O��1!↶�VL��E�M��1`���OT��I[$b9\�Y󋀟dv|T�5Üt�!��J84�q`�,39�]���;Q�!�_���cqg؅MG��xa�Ԯ%a!�G8��q�C��|1�����NpH!��>?D2I�0@��1f�%G�!�Dɢ=�T᪐=|�<���bJ<��}җ�h 5OÕ$�pi���Y4a����5�O���`�i�O6j3d�{D�	-B�9�ȓw��d��%~Fqc�
�=vX�ȓo�T��#B�"?�ӳ�� P�ȓ�D�ס��9:��m�8H��p��-�N}CS�U�o6���&�ٻ	�$�ȓ���I!�ςp��E�bCT6dW|��ȓ�h�ȣLB扲�Ț5���E{�O�\�����>@�:c/#x܄���'7�mB�aΝ=�X�h����:m4��	�'�@��rh��v1�D�Q�93L�1�'t� 앆a-���C53�
)	�'r�Q������l���ù���h�'��js�'<e��r
�]K���'tX5�e-�x'�x�j�Q�޹j���hO?�r`
À���LC��I�TX�<�SmB�`�x�r%$0|y�H
P�<aQ	��x�u�N	{�f��@QJ�<)�J�KC�´�� s� d�5�{�<yQK�,��<��Z���<�f��b�<Y��$2T��C$h�#Jp�%�PG�<�s��=Kt���� 1~Q9UB�B�<���A8*�
]9`F����hqb��{�<aDn|z�Q�d�F,����L�<!���A ł4)C�o:�� �L�<��ib�t}
u�)4��=�IG�<�R�ڦ�21�g�Q���%�D�<�Į@#HQ�\p5kI�\�^�*�hXF�<�pg�j�lK�H�qr�B�Ll�<�S٭z��$L\� ���Bi�<Ԋ�*{L�`��*�Q���KT{�<!U ٍ��̚'�ҎmK�0�x�<����r�b1⣀� CN�ȅn�u�<!�I��I���Һ*,��Ɩ|x�Dx�
�$a)�� ��!��u���O��yBoٍ(�vuPs�ف?�Q�!�C���'�O8�+?�D/F50,�|�B���8 ��)W	G`�<%H�)T<a�ɡ'㒕C�jLP�<5��c]2d��w��Y�E�<y��Ŵ8���E�f0�"E�E�<�s��p��	�MK�1ؔ
��<٧�ɴ&|��JVi۝�^�;�!�|�<�v ��Z�0�s�a��(^�p�B�	�iX�42c�P���i�9�B�	&$+��M̯J.J|��!�=�B䉯C�2LQ�	��U
H��׍�NU�B䉌n���1(ٶT��X��U�K�B�,�Q��Ӻh�����`ӑQ�4C�I�/^*%Y�D�`Τ���ǟI������L����:�(�ɝk'���"!��8+=,5J�A�
z���"O� 68سfԟ'!�l6�
%B� �"O~I��YM(��f
�cf��"O
9Ȣ`�7(�8��*>t��V"O�]ş�]I�<Ht
�)A�ּ1�"OH�A��	&��<�S��"3���W"O
X@��~�� Ҧ��/.�)��P�Ȇ�I?p
L��I�x�+�.��C�	�.�)��c�MʂX3d"�
��C�ɿN�F�8��\�9P��ac��R{�C��;�@i2S7�Nܫ��	:6�C�	� �PȠJҢ[� ����I�	�B�	�R�����f� l��@S$���$�WP\Y��P�>M�� ��N ��Q<� N�=�:psb��i�%b��_�<Q�#��F(�A�!z�Z�٥�D�<��+D6�Е�WL�!��<鐅|������:ʉa�Tz�<i�l�)ZQ`Q�H�8�x��'�u�<y�/�?~������d���BIs�<�gm��.|9���@3�%!D��f�'���_���	[�i���g$\]�B�	�Q�f����{���6�J�_l�B��?�	�FJ�_eP����S~�B�'4�4���"�%C�@2� I!�dE<�(�F2�M
'i�e�!�䁴
2|8��٩A�$�*!�ĂlID��*�68���/I�T�{��|2F*G3ְꤢ�~�2���-	!�d�}=�4Ԡ��Eh�d v�;{�!��W;��0:7*��IR��KT�E�!�<#�vX�t�ؐi_�i(��H6n�!�L52.8j���P|v�z`��8W!��Z�`�t�_�`�qVB�FQ!�d%bB<iY��їR~���aMf�!��fW8�"V�۲FNz�`�`��Y�!�϶y���5D�(9Q\Y;E�؟9Y!��D-7,��&��a^�)a�Ǖ4[V!�D�Qn2��瀟 0���i�;'!��7Z|�ᅉ�#qL<��j˗N|!�D]n�X�g܌�L@`4���y�!��,$ ��7nڿ���@�Ub��R=Ob�b��`ȍR�Fߦp`�}�$"OĥږƆ`�jM�k��u~�\�"O��(6��8-o�8��	ė]~!Z�"O�ѫ���<�6 +�IQ���"O�T�U�ޗ19J̱#�WIBС"O�P#3l�z(a���$l�"��'��D��"[����JJ��!@ܱC�!�ė�b�j�@)?�1���6!���<}er�����mHyk"aJ�.!�D�K�TC�i�9Z-�7�ӽ/!�D�Vw�B��ՓT؊�s'o��H�!�0R����1�M�N�|8(��n�!�$�).ٮlj�L]�	��x8���t�!�$��w7V����ƣ"zf�Y���1�!�ާ��q��:j_��릁��!�P9� $��6[�U�b�	!�_p2����ݤfS��`�!��J�!򤊚[�X��%�]'O5>1_|NX��'��Lz`�++�)�����/mĔ	�'�P]�Vi�Bu��jQ E8\B:�H�'n(�r ��2cՒ؂�AV��t�
�'��0{dFF�\��0k�w@D�	�'~��J�l�}h��w!UuJtY
��� �ڔ�ĳS 섡�͆�r�8(J4"O,�����A��$�d��9�B�KA"O ���@0o�*)CA�9�"�z"O�E�B��0hԾ�G��o���'"O\%{�,ϲJ�AHD/�8n�X���|���3�'%��	p��*~Q+����9�:�����)�iS�9�G˺4��e�ȓD�8�cs���<x�QP�a�~���(Lj=�"L-J"-���ܑ㶀�ȓ`�>��q��;?%p���WP�pE{R�O�����E�!�0<b�C��N)H�	�'���J�jK(Vv%�Ú0YbX	�	�'�ijS C
y^Έ�����!�rɩ�'���c��^+T�,u�b/��&���'���BQ��MT^�p�B<. ��'�1Ҁ� 6Ș#l�2�&��'&=r����az(�Mŕ7��%�N>Y���	�6&���"ֽ� Ş�#!�D�4H����wM�uw#��ff�'x�M���4TS��h�䇭$�6� o�y�DT&˜��"c��
Z������yb�Ǳ}����B��P��A͏�y"��U���A�P���K�1�yB�_�����H�+�h�c�y&�^�b�P;X�� ;R��y��ޅ}�����&��B�Z�s��!�y��6J�B�U�M�A�ܴ���Z�yr�T4p�<��fT<nw���v�&�yC�w�
`aF��;gp�9rw�S��y��Cv?z����k~PpY'.��y���l���雏e�\"kE?�y��J/@��ӄ�[��8 2d@��y��D�b��/O���R����0>�� ж/�.ݑ.���ݨ&�y�<I'��N��eSSg��(� ��j�<i��V�#L���V�� �AD��N�<�!����h���������
K�<���ɉzEnd�#
�q�A�[m�'g?m0��py�!�(ř � �+�@9D��� L#7�5���*��K57D� k���-q*�K?Y���3D����+��Gq�]�R� �V��S�.D�Z����Lpهc�� `��b2D���0Ȕ&t���瑈'�%�Bb6D����N�-�D��@珂3\���a'2D����"H�m�R�	�ID}�!�%D����LC��F�1�'U�^�@a�B��O��=E��A�<g*h�t
+�.�؆X�!�$��T�&/
cdH�*7��U�!�$�2V�����C��N[촀�ꇺs�!��Y6{�j����҄	Ft(*���p�!�dL�w����2O��;FYQ�B����'	ў�>u��o�*f5����C�+*2���#D��W%� �ƅ� �C��4��N�<��N�*�B�d �Ol�t�%	]���b����j�IȜ����6���V� Ո�D�<IZ��E�VIp܇�m�0���eEp&@D�2 P6�v��ȓ_�ɚg�!�ڥ#N41����.�f�X�(�pu��4Cӵ�%���xTkw.�S�P���'�j+@Q��d�m�c?8����ƺ2 ~m�ȓ)�vԊ��F��} @�4X�&���hn��"+7^��f灭/��م�S�? :l3�@x���fY�o����"Ox�&oV�VXXa�eS?<{����"O���FBȖ<�7eKY��E�"O60Z�gޏmڌi�C�+���yR	�:H�Q)�g�ҌX�C�@��yb�ɶ>��{�����cŨ�y�X$;}��)�8�"u��l	3�yrA��1�R
ׯ����x�v��yrkW�8�:hi�͖&~C83Ve�1�y��1�*d׈��`�3 ��y�#�;qMN�82!�Q�.P"
�y���IҚ��5.����w����y�dҽ��y�j��9������y� n�`́e��9w~�`��K�y"Iøk�!r2�"k���P��L�y
�$�ޙ���c���lX��y���1H�J ��B�X�������y�ʊ5 ޖ��w���.�"h��y"�;����%�<$a�ή�y���F����DE�$�RB�-_"�y���C�B0!�`R� @�6�ygI*6[h-��4FQ����&Q��y2����<T�޷ifR����Ȳ�y£�r�"ћ�/JZ���a����y�@7:�37lN=%�D����y2��/�بp+�J4�'ꞁ�yB��'j�(	T�G4s�P��GGC�y�aϐC�n� �7������y`B,IrF�� �
 3��� ,J �yS<cF���N�%��J�
W�yң�9R.���`#s�P�+��8�hO������0G`�xʄsՌ�lM�E�	H�O�:�#dkGhb���B�H�H��'ϒ�A�lT
Mz�UKA��;Հ͘�'d����QQT����֜9����
�'����7J�,!8�ˑ6�\�'��l����&�!c mH4�d��	�'�R�A��������#(6��:I>9���,�� �������bK��Cv�L@��B�I�/����󇆓*�r�9�JՇʾB�Ʉ$��	�B�G	`��i�	�^��B�I�uZ$���P<<�h��>�B�ɝ~��� ��'Xx]z�o�<$�nB�I<7��!kׂ�&d(]��!+�jB�I>��ԋ�H�r���$�I#KJ�D{��d bhΦ�@�'� 25���zgH�E�<Aƞ�Dݔ ��N�|���FLj�<����8���SD��|�a�D_j�<a�N99� ��&�_d��7�O^�<i�E�gI��	�oL�$�T!�P�Y�<��!c'4akЊ��r�8\�� T��hO�'|K���#�?x��8��ťT����	}~�O	�6(���Q�s����ݬ�y"&D�a@(-�D)^g%�݊��?�yrǅ�i�aw)V�dA�]ˠ�ǀ�y�gҤgƆ���5W�J��0�I��y��':�49H�SJ�p`�
Z�y�.T�"�(��D�^����y��B��z�(���;?�0�`ĢM.�y�([���;�C�7 "�q���?����=8���]!F��� "^�|�^1��J�`��
"`b,셠���ȓt~���H
�leް0Ѣ]�Y��m�ȓq������r.��t$�>-�8���S�? &�)��פ4�A��W'"~|I�"O~����ԅ_\4xV'�u&ٰ�"O�쨔"�M�����$'C��iQ$"O<q��d�m��c "�\P�@"O���`S�#�轻�CL"d�N��"O���G��?��dM�'wY.�!"O���"]�%�f9�ʒG>�Jt"O���F�W�h�fA����`9�"OL�Q�&�Z�pc��|�$$#1P�t���z����/�+t�!��<TO��ȓl�N5J# ��l���N��Xz8y�ȓ)���,�:W� Pe!M%=�Ƹ�ȓ>���jq�ƴ'���c �&�ҍ��;ql� $�44�d��a�7�x���,K�$���n(^試Y2y�xL�ȓC��1�(��nrz���K��ч�z��\��՛TQ�xy'*�+m���ȓC24�W���
x���j[�T��ȓH�������o42��)H$n-Z��ȓ~- - d�d��ݹ����j��P�ȓl�N�g�M�Q"���[$kv�E��-����7f���[�$�2ؘ��	w��������b[R�䐓c �7�	�O<D�PqpN��}�X@!�B�.@��8�IM���(�Cn�T��/S`�$U��I8D���Sy��4�R�C���D�7D���5�7 ��q�(PW��"�4D���p+^"� �at
P��^�e+6D�h�@ҬGk�q�O3N2m��d3D�0Z�9\��.!��hhfn2D��Ra
M8a�|P��L;5���{f$>D��
Ƈ�+dr,�Í�}D��:af<D��f�h�XPV�*TJh��n,D�XkՌ>L���0��
�xMHR�6D��j§˼*Cl���g� e !"D�L
��5d8�"�<��d�G�,D����.�A���)�"�t�<Ypj+D�����cXt���h�����&(D����NU�q�&9���A%���#%D�$�O
`��d���56���!D�4�3D�O/ޑ�q��y�b���?D���>c�� q�:BBh����<D�h�T/�[���p�`hpT�<����Ӂl�>	z恁1n�����$TJC��d�~�ztG�݆���fZB�ɿkehU� �X-X���ӊ��3��C�	��plZ4����[V6��C䉠:�:(Jk�J��kH��xŐC�1�$\A�!��K����g&k��C�I<ن|3_�,�5��4�>tbш�<q����]�V���kt�`2������?D�`ȣn��I2N��@�H��`�>���r����Id���X�`"O������!�8ᛥ H�3t�p`"O�s�$�z��&Ɠ<3d"ș"O֬!�J�I���7cնX��1$"Ol=�'�� ;F� ��a��)&"O�m{va�J0J:kBLQ�"O2l�re�:S$�Ю�*6v	�"O&d{1�\hEx��fϟ;u�����"OD"�A�BD����Lj�4�bt"Oޕ[��|�+�MŠ_��\8�"O���%U3퀔k��St�H��"OBx�"�]�0�F8��"P:x4`���"O� 8t��"��p ��4|1�"O���#��7W�Dz�
d��y�"O
�xum��)�,4&�|1X��"O��5')���1c�O�} ��r"O�Hv Q NC|���31���Zr"O������>q���uE\�ui��"O�����=�.�a�Q�!S,��R"O���c���P�1�D=�"O:(��;	Gހ�wm����,zp�d;LO���,@�%����� 
�<%x�"OƉjD��;s�� qŽ+���:�"O>�
�D�
/6!��呬j�dz"O ��%�Z�,����N�Q�f��b"O�T�B�j��Q��M�2vT@FO� #�ݞA�������D��0��5D�����2ab���!��2��x�u�9D�P��!�OP@8c%6�P<փ3D�XkI+r��3Ԫ�ac0`�5I4D�x0�M�o�y���ѡ:2�DR�=D��[�i ��
�˗ � 0����BB=D���dͫ}� 1�̰U<x��R�5D�`��$�;9�Ft��D��r�P��(�Is����ʭ}e@U�ƭ��e���� D�(�BmE-�=�'mN>SpC5&9D��ѭF�c� Ds K�1xF��<�Io���i䣋�
E���
ð��@�Q�5D��*Q���a��ឨgm��s�(D��ō�"i&�9T-�7$Ֆ\c��1D�H3@ץL�Fa�&���V!��1D�d��c�7
hl�^-N�<]��O1D�D(��0	H���-��|A`/D�쨧e�-����k��qq���<��(��D*�d
@��!�qF9tʦ(�ȓ9ȐĎ�(�~	�IS2V��9��Za����,	27�Zq�b�����I��0��b�&�/=1(���C2��ȓg�ȅ���-'hE�%�F�w�^͇ȓLK��07NS��EH��!<���?����~Rt�h���i��ǉT1��٦��h�<!�䇪E>V��sa�'�^u�am�h�<1gGL�|9^�c��&w�XI`dJ�<�����-B E�S�@�<�PhY8�|���	�	^�H�ČZb�<��Գh��d�����|�@M2���\yR�'�i��S8i�n�r�-͌o�
��'p��#UT56�D�%.ǝ_O`�
�'f�։
�%!�`�GX*U�>TR�'��iZ#� $<x��E�#_iv,��'�:h27��](�A����k��9
�'��H���9 X��Mĵr-ZL�	�'>j�
�,ɚ(�j�C��8jL��I>)
�{N��CЧ�.r�X0
��I�f�~܄���h"�CC�]�r�駅�7ذ�ȓ"�9 CH؀	H��b�)/^�Є�|�9�G�RI8�!���U�Q�ńȓk�NAȑI�	Pv�����^qq���)�d���sHl dm�;m!82;�y�iE�tР�s�� �\���OF�y��v����W�О\�଒�@;�yrD�w	l@��c�;>j�����F0�y��:OI\�S��ߏ.��-����?�y"�e�4A7CK֨D�Ĉ͢�yR*�"K`��Pū�*o8����yb愑A��h �؜�¥������0>� ��qF�"����k�@=��q`��]�O�"�z��
�WJԨ�e!�"m([�'|P�b��M��������~����xrjV;.M !�%Hmt���#��y2��aݐ�(���2S�!�����yg�8yf	;���*�r�*�-���y�&���yD�r�4%[VÕ��hOX���N�f�34��g1�}�F)�4$��)�|�4�QN���z�e�:U���'%d|s�kϑN�(��1��sʐ��"O\�k��E�yR�3'��1xD"OT�1c���|�$@�/8W�~8*p"O@U�4lǢS��co�k�xع��'~�0�����a���5c�
�3��;D�x�V
�i���[ 	�6���[h8�IT�ИOh�	�G�O�on�󯐊
N���ϓ�OxA��O����牐H�~%��"O�LJaI=,�XTٮ'��#�"O���r$�YǮ�r��ў: ��� "OV*`!�k39�F�l~���"Ox,��׊���cFسvi�C"OTi�2��`�w��k֘S"OH��p4�pR�D�[|�pӖ|��)6Ha$��.Pe9�@�fB�	X�~d+!H
S�B!�g��W@TB�ɒ2�Й"G�T?�����DI�B�IO�x0�e�\�/�� q� �U��C�I�R�0	�b�E�4wjK��K5��C��"/�@b�
O�(%bgc]�d�C�I�e����"KK/bP���#6vC�	�u9�@�A��^f���Ӂ���0?Qֈ�8�@���_ !4UJ�Ʌ~�<�	Ԛ^�
��_�+ɀeX�N�}�<A%H�_�8U��L
�H��\�FA�}�<	B�Q�R֤�1�E&6���w����<�dB�-s�f
A�08ӄC�rx�Gx+�/  1�Ğ_�N)�4�$�y�C8^�F@0p�
�GR��S ��yR��]ޡ��R�r�tT��D�#�yIS:� y��]�0mIt���y@��0��/ӟF��T�y�o�h�Ľ#��M?Ϯ豳kU�y,�fu�9��Y�PL�c�3���0>Ys��G���ab�� e�th9��_�<	)҄V��5"T����g��[�<���% ��- f��;y���C	Z�<y�`4���%�=V�CP��R�<�vi�Lj.�W-�$��<[VdRO�<YsB�=X`}ҧ.��|���2�fCK�<�G��O�8��r�
, ��'��Jx�<Ex�BÞC��#"�$��8����y�o�/ 
�kQ�M�����y�:i�J���X��vI�EhX��y�FƄ$�2�YEbːY����0�y2 c1�`�cbԇZ����?q��d8�c���ʰ�H#L�2��P-4&�neK
�'3���ۣ(.$���I���̨	�'%�#p��2q�:�ca'C�b���	�':J���Y�yb�%���պG����'(�a��L�;8VxX�W:�ܔ��'�μqd	:ܔ�����5g�����'_����i\���ɜ�Q�"0B�'c������5�b(�WNխ/4���'J�]���":�e`��=F�B�B��� ��p��Ȕ����V퉟7x��� "O�)��l��ۅ*���u;T"O�Sb,N�[{%� �e(t�"O��
��GQS�1�'�rPxD0"O $c��L2�yA��B�\N�TZb"O@� ҇r�t(�ÕGD��BF"O5��&ʲ&�x�(D���e$����U>�z1N[	K}hPї�#j钜��%�IޟD{�OfB4z�Gs�JM�w�ֺj�Ju��'PE2Q�S���X�&�\��a�'N(���@�o�(�b��<�����'��ܛ�G�@�����0z�A
�'�h���փ &D����E`b	��O����'�p;:xV"�&r�5Y@�|��)��{�ִn�z�
��nq��ȓ3pJ��Ł#��]� � �b��7�.pѧ�܅_��0���!|X��~�l�!�: H��®L�D���ȓh���f1Y�N|Ss�)6C�IB��<�F�ؑ6�	��2nR�C䉄W���U�<hc"�?%�N��1�S�'����1Ԧ��o��^܈�N�x�ўX�'�>�����Y M8u�ӯ5�V��QO/D��B��y*�b�$!�H@��/D�õ�r.<�E�O"?vD���k)D�(@ h���Ұ䁍
f�[�d5D�$# j��M�:0 �#i.�ȳ#4�Oh�I)�qcp��*7#��aG�R�"C�	f�L��l��,�5%D�'{C䉑 3R��� 7�적锣E��C�I0Y��}h"R8g{d���S( �C�	� dLĨ�8���`��gC�I(W68��e@�RX��#�	��B�Ivۜ��"��3e�L�(3�͜��B�$�b�"�.9���(V�&��B�,U�܋׮S:�@���OR "��B�I/ע$�s��0?P��c���#�!�DU$ڤĲC��4=5��q����"�!��.ZivI�s
�	&-�������N�!�dhA2�`�/�/
�$+5��3I��'a|��</�D� ��0�6��"Ҵ�y"H �M����0��	��\(�y�C¾�d���C�#�� ��/��yR6_U歑֨ �-�j�����y���R/�hx���<���d#�yO��JJ�]��BC t�f�AU ^'�yI�5�<Ęs솚h%�ykg���y�L�?��25o�_i�Y[�K��y҄��O�Җf]�PӀ���^��?Y���S0��Y��J��ɓ�Y�fm���ȓ6��Ȣ�P'c�Y����J��ɇ�o�4< `F�?�4�ɑ��ZN���9��p�)�"<�dD�GY�j�6���d)��	@��X�Bh*��[3U� ��QC�����$%3���ǣhj�l��Ug��Y�Ih�h�D z�~�%� E{���dزqPt<A᎟
��T�y���&�@HQ�C��hIja�ɢ�y%S?q������Si{,�c]��y��˛E^"�YSab�����	O�y�㙬�z�Q�ֶ}x	C��
�y�猞F��\(R���s�q�2L�9�y�
�=y\A7mˠ>Y�@J��y	_#|ix�lF�/GbE"'@C��y
� ]�TI�OF�\�0���@w�e��"O�U
��Kw����G��-o��"O��!�[���!��ÓQ��a�W"O��A#�8�f�C5C�>W� aa"Oɡd�ߝGтq��3s�f�{D"OL1�c۠
���ŶC��ي"O��*ԝ5�`�xg)��<��#f"O��S'&F"L�)ڞsV����"O>Q��L�aM���N߁w<d@�"O:����]��h��kI�C4]X"OL���͆0ڠ,� ꂴy6��"O���������|�D��.+$�D��"O�I���I�`b��*52�0@"O����EBa�S��A&J��P"O�x�Eh��!t��D�!u�9�u"O.;4�T��0��s�M(%՚���"O�5��ƬA��%9�aֶC�A8"O4컀���<�f��%5��0�B"Oya��t����h�L�p@��"O�q����F]���J��o�ą��"O�����YR�@"g�?{��kd"O�� !��1���z��CP�""O(5�sRш�H�A�]�6��"O���⅚����ȣb�R13"O�0��M�6�.Q�BZP�J�"O��0���0D�Hd�v��0D���"O�Äŵ=j�Ep�aJ�0�݃�"Oz�(׊J���KL�&v��K`"Olj�`��	v����:A��Pka"O, G��G���Tċ�{��d1�"O�-Z��X;@���C`#��ho��G*O��
��B���U"��W12Px�
�'Z�s�ON�6�2h����6��{
�'[�@�gL�X�v`ȂcR0r�RH3
�'�*��B(��*��u�2 C�{��IB�'����b ckT<�QM�=w�<e��'��tJb(A�gǆ Q��x�H��'a䑹4�R�{p��0�O�o����
�'SH,��� �|H@!߸8mj�y��@
I�� �. �{�H��ª��y��!&.0}��μ
!\$xb���y�%��L�6�}�<����y�N״}l����n?Y*�`7�y�
��3D܀9鉈q��Ied��y"�I�+ɚt�i9S{���d�B�y�cZL��d� A���ʀ�y�J�*'[� ��P6@��`��y�B�3 ��'_�8���� �y(��&tS3i��[�q�X��y�g~�p)�R���@9n��T�y��Ս�.ek��ۣ<�yZD�G��y�eD:�h�p��6��|�#�y��4�μ��d@0$|�� &�=�y�N���5�Ga�'�:e��/�y����(ڄ}i��3��	�3ȝ5�y�F^��>�:�f��0�gK��31"OP�Ò(]*]v��[��\yB"OЄ�DOZ��ش ��Sk����Q"O���R>���
��-��]��"Oz](6�	V�dX����-"���&"O������F�$���*� ��"O�a֎$�J!��I��Q��	
�"OB̛5�J�4$yӣ�w���"OH����+U޴�ף�E�%��"O� |u��@K��`T��(tGʰP"O��/ %;�~� ��ݺ="1�D"OS�k� �	t��U��I�"O�P�"�j� �aJ"=at���"OXu�`Hњa@��2D f�d�V"O�))��^�ZV�Yk��ٴ"��U�"Obx�c�S� 4����!]��习"O@�RK�o5�0��ֲeJ%C "O����Ù7)�	6M�`J�`��"O�p &MZ�O�>�87+�5	b�"O�d	�*�2��yq�����:6"O08�#.Vo�]��K7Q��`"O<�y�A5��u!�75X���"O`@�t�TI���N�&�@��ףJ��y��ϊ�4M�LÁ$N�'mG��y"F[;q�T��գӥ!��i����y���f��"����T"�ΐ�y��;�P��o�c*Q!����yR �Rq��st��?;�e���N��yb�Ħ`�e��U;5�|��P/�y�.Za��y��C:`It0��a���yB)ӄ*�ju(�NɠV߼I��,��y���$L�&tГ��K�`pw+�yB�_�
R�܃�b�CeҀ�f\��y�(�O������C�Dh���Ӌ�y�j2El6р�蜪Jx:�a"E�ybA�	�x� ��/��dP1�yr�|��h��@O����:��Ѐ�yR�I�lJ�r&H3r���"�O
��yrd��u\�A1�+F8 C~�)��yB���:�F�6J��r�v�p�눥�y¡��&&�tgʰoLZ���U��y���v�@��@�9l��ͨ%f���yR�8"��i$ɐ�`B>�eb���yB��&��0�7g�)I�����y2!� B�ba(6�ח\��Y�$ D*�y�C�D����֞}�h��/���y�B�('�d���نK�Ɖ;3I���yr�M�HHkK�=&d)k�FU��y�΀ ���	����kP���y��Vu��)bÁ�~jX��W�J��y�D�~����4㙙l���1G���y2fO�9��@��D�\jt����y�A�M4��0Ҋ\'�"`�2�Կ�yB�	�La������Ქ��y�+]T��qT-O�����l+�y�Ě�O^���.@�PBхU��y�HM��|k����k�T���y2fM9]�ɨj=cA��Pa"U��yJD1j¡9��.�������y���1(*�����(� ��n��y�� lS� ��m�jp��ВAL'�y���HWLLz .]]��p�"!�?�y��-�>	zQ��Pq�MP�	�y�f�>��Ei�*ɀM��y!#+�y���iV�z�R�N���cCD��y���^�(��g�'=�Na�B����ybI\�2����mZ	ӌ4
ɋ�y�j�� �hu����b�$��!��,wf&���O�1j�����'�!�����p -[K��Ti�)�(8�!�܆Hrqz�҆J�X��TJ�T�!�d�8s\eI�B���dE�;%�!�djzxp�nE�u�nXCQ h�!�� � �'ㄊ*#x��A2D1r�XP"O,sԈCwWr|(u�X�+�G"O�
q��:R3GBn\H�"O8A�`�T�i��HP�%��,��"O�hb�C�@xa ���m�C"O��X�� 1�L�P��ڃS�4`��"O�#�J�
4�����,B|#"OШK�I�|Y�(����5V� *"O>H�+}�x�7��nT�]��"O��:�n�/��8�%C��E"O^��h�`����74��"O$Ԩ��C���[P#H�`��"O&L*�a���j��I�(�uA"On�xr�גa� ٩�h��u�,AK�"O���c��)v}a�&5m�TÆ"O��2"G��̃x|��XU� �Z%!��3�n`j���y�M@�ʏ�s!���@��σ-[ XC�])�!��Q�B�%��i�t���!k�^�!��r��1f�X�;�d�����'���yc�D�|��`'�ؿpv,<�
�'mA��`�'��@:���jd��	�'��)�
EC�lȥ��2�(���'��c�J<�%���'ì��'Β�1k�(}�����b�&����'��I�&c׹���Uȑ�J�Pu��'���i�k9S���Jd@*Z$2�J�'j�m:�R/D^X7�A�!��-q
�'�x�c��͚
fH2�d�1R����'��e�wD�))�t� �!.�^h2�'����GK�@�!�{��TQ�'��0��j��$ u�7g����'��B��C
|�
���D^�j�)�') ���d�})����AR3Y����
�' 5�D���	���`
��QK����'�LzeC� �L��@M�Qt����'��1�߈���F@
�<��'ưa"��9G^�N	�ԈH�'�����D�1�����	[�,��'�
,�:�r�HF	/�"�	��$5<O�}��o�1D�>����*G��l�"O��Q!AȈ3�
d�����"OH���(�,�w�U>o: ����w�O0>XKĢU��8SB ��{6�I�'��Qrς!J�>���UM:�� �'bў�}zЩ��W<A�&��k��b�"H@����>��&�&�ۃ��r�ё��<)��٣q� ��r�� ~⴯a���d0�h��2w��!�Dm�DFH3 �@�ȓI��:�NȢܰ����_u�lE|b��S�D}����3����풊hT�B�I ]�hL*�
�@�liC$�]�.7��(O?7�1S�<٩�9��9Jh��`�!�Z�"D�������B��bE�֣�!���&�ru� B�4?��Q����!�d�RJ�����@ ���� °;!�
"p�#'��U�x򀀞�}ў<���7=|P���:�p��W@]�o.B��9���ɗ��Pƈ�(��@C�C䉋NIΡ9��1�~�s�)��d]��䋔A)�!2���M���	�lR�!�!�ź0|ܼ�P�)s:9�ԫ�&zU!��ڙH�,4!2�$l,�0K� ��O.q���0���A�ܨ=���V"O� V9����4}4�@�f�ߎ5�}K`"O����4��u��ɜ�t�Ԍx "O����R�~e�`OC��	�"OP�+�!��~A`Ar�m޸ؤ��*O"��H��3��8{'��be	��'^V�pgl�6-膁�_[��'�n��2��T�T���&Y�0��'��#�D�)���͗E����
�',�q�aE�98�ڸS��\C�(��	�'��8�#��"q:ٚd�!A�^���'�j DG5j���Nʙ6#���
�'e0��-��2�(Aa�嘖f���+
�'$Q�ŋ=(?�	�2��<�b�k�G$D�쐔� X. 8b�W&c�,e��7D�`�ufG����:Ø	8�!�F�3D��A#�^�gw��&"Y� x�0E�1D��P��@�V�Y��BY(����`0D���c�=��������2�,D��A"!�Z�@�撪'~�:$- D��
Eg�Y�(R�)~�fԚ��>D��W��(���:�&P;p�����.D�T����T�@9��n�][D�@�c"D���A�8{$1�����0x� !D���C�gD8s������y�>D�� �ք|�����.�9��c!D�0�W��0R6�##"PG��
�N-D��ڤh�
j�!��̨X��X�S�&D���]=6���� �T�,�Τ)��'D��	�Sr�	f��B'��@�L%T���۪K"xyK�n�l1�;�U�D�<����O��pD+�#�^8��K�g=N��&�'���	fڐСf�9�P��B��*2�듍?
�Ӫ�lѢf���b���,��$�I��M�����OIF�����1t`�qל-΢�#
�'��]Z��$HD�b��%Q��$��'=ў"~:���;|]H0�$dJ�bZX��R��m�<)p \=P�JQ�H�<¬�z���eyB�'�2Ux��H�\ڰĒ���ZQ(��'tH�a��]S�l��&GR��p�'�x0��_�Ĉ�υ�w��l�
�'�l��,��9�zP�tB�';S���	�'��e��&��+ZM��B�,��Z)OhEz���[zVıR�7�:�9c�A�:"1O����W1}�hx2��4O���ċ<{�ĩ>���'-	 #�κk��haɢ'=��k�'���g/��kQ����ʄk$���'j��[�l�(��2#l4 �9��hO&��ьx��1��"b��H��"Ox��`�<Ꜽ�p�^�=�΁Y��X���)§1������>`�$m�S�Ĩ��lm�D#|O��jS.��h,����o@�i�d��U"O
�hT��]�hx�o�!(�Lx 
O�6Mݽ%Ö��7KE5K��V��)�1O��D3�)�$!bJ��腪<��ԃ2	�P�B��^<��p���|���a4�
��B�	�-'f�	TGR8��4p6Ϟ��BB�I��>Y�J�sU����/@�➨�����<4+R�b��Q�rɏ�w� B��AZL�hAHݿj�R��c
S
��C�^���Z& )aL�a�d�C�	�J�X���%M@&�i�$L�S�zC�I${��܃GM�#��T�B�	�@�$��'��X����7N��tB�I�CP~���IG7k<�$�G��]��b����)� �����1 �$0��� � %�d��'xqOpB�gֵq�R���D /��ī�"ODy�����v$��I_��ṟ��ITx���U�&=����q�R�:��	�1�O�� M�����G�XXiD�i_ꀆ�`+�@��.��pg�[ j֬F}r��
T�(]Ѐ��>CR�b���B�Ip�HJbm�hV���ͮU���D&��O�1���x�OW�A"�01��g� �"O�q&-��u�6dH�-��c�/O:��Φ��S�'��9O��sr��`v̸!�� �]��"O.���şO��)+q/Y�=疘��"O�y�	�7��A��(�T��g"O�y;&-F�l�:u+A-ܐA����0�'X!�ĊU
QٱF��U�j]��jN1O�"=���Tʕ��b9�$' �����kD�y��Ϳ3�|X�q���X"u��O���$�-4�(��DR�Ƥ[��_�!��� y�*�H�oK"+��d�	�N��'0�|�F�(*��Ɛ�}>d� fl �hO�c�����Y�	�1_GB��.�&d��` "OVY)"��Zb��˷-��ai�4��Iw���	=E�4�;���(.�a1��:1s!�$ގwӮ������ $I�`�!k�'���!�S�t�ҩaG�D{�Q}�V��w�X4��?I�'�&�di�;��x�ƚz� ��
�'��0SeS']��: l�0o�Z��
�'�*@���>?�I��!o�@�S
�'�ū�-I�h6F��ņQ�m���L��F{��t
6_��@���-Xt�@��ޠ�yRM�6-GERp�S�d_��ɥ�͟4�4x%����ok�$:d���T��[�*
�)�v���%�INPlX���dq�Hɇ%� B�I5b��l[�e�3�B��5��	x�C�	�B��b�|�:�{G��
B��4YM�|S�j��:<⡯ߤ��C�Ƀ&:��:�%�4�U�جGG�C䉷9����oU#�]ro��x@�C��+Cy���T�9@έ��J�2֎C��'=��ݓR�~˦�q�8\d~C��:L��p�� Y�d:ĉɔ;�vC�	��rp.�K�t4���Ȩ-�~B�	�^���y�O�[6L�i���k�*B�	/.�EX�ܺ?qH�k�|�B�I$����(�&a��+c���l0B�W�����S;x6z�8W/A97��C�I9U��A���;&И�[%"����B�*�.Uò�H9[.�e0��5l�B䉕�L�Xca��S�$���Ā�F1�B�I2����E,x����ߕZ�C�	�e��(�"��4`��D!�J�PB�bq��b �@##���C��D�u{4B�I�j!�ճ��������ʜJ�.B�I��ɂN��s�:q�/ڜe�B䉮K?`p��<'�x���*R�ZC��:�TA��d{�,#ua�;P�&C�	����*ԋv���V<0Z�B䉼1�V��p�L�&h��ѥ[{�Y�ȓ0�z@��҇� kS$S#H�Ňȓ �$e�8��Ua�+ءU��X�ȓ?ߐ԰�+N��L�s��ׄ��M�ȓ*1�]�g&��R����H�>"�V���o��a��[3Vv
��ƒ2PR�@�ȓ.#���.�P8���.Qº���S�? ��	h80���N܄*��)�"O�P
âD�e��������j�nq��"O��ᣪ�#{]朡qB�9֨��6"O�L���myXm�R�̾)iz����'2T}+���o�*��C�#����Aa�4>|�'�dPCE+8!�Q&�إ(�ʨ1�'� ŻTE%l�2�KJ�z$
��'���J�
�����(Dn���E��'���rjΏ[j���z�B���'��=y���2/�t�0��Ӑ'��)��'[�8�G�����@�� nr�9�'P(I�'/�������'���	�|_t�_���'�BGK��h�7.�
\�r�'k��H`	�5n-�@��MZ�:��0	�'(*�:�eɛ�d�
D�$~�y�'��	�!�$nw���0��3Q<(�'Y�̈u��'_?r�*� [�xcU��'7��PD��'H�WM
�j�&U;�'Ә��QĞ�gI�!��k�NQ��'v��$ W��i�HRH�&��'��t��Q)�@H�Å�*I)�Y��'D�$���<�4u�N7T� �+�'�쉣U��zZ���E{�"��'͌I��d��Rt�@�K�'u~tQ��'�����2h�������)n�4(a�'�"y��L
iR�I��I��		�P 
�'���bF-$r|P�!&��%2��l;
�'�t�P�K_$SxT��5�D% �б��'DB�14�,V�:%���
� �'Ax��Q��j*��)!�ܒ�bi��'��|��m�11�|m��C�����:�'#\�S�E�m AH���(1�'V��P���)h ����̫�'@P��r�A�d6jg�\�-}��'(^��s���"o`|�hؖ|��A�'����%꓇S��i�gJ$��i�'��5�S��~�� �HΓ�<��
�'$L�kEm"9 ���F��@�d�'\���:.�~��Ť�+�Vg1D���v�[�W�h�2�
8.,,����-D�Ъ�ĝ�G��	��Ƙ&!(T��D+D�t�� +~��p��ǉ[��2�3D��գ��R	Ti��n|�s@j3D�
q�ы:wl
��]4=f)�5D����M��U��)�'aZq�Z��-'D��iR�ȃ1�LKy:1��J$D����^H��2�$ͭCP��11"D��H KB�FL�%��
%8d(�ա#D�\��
M*�Q��
�F�xso!D��*Ԁw&�hbm��.Ĝ0���(D��Z���B���d�ҍhɨE��m3D�d ��F,i�x��F2���1@a4D���n_�0�r|�r�O��4��"2D� ��%w�P�Ӵ�
(9,�I+�b1D�\y4�¥6!%1(Ϗ)4leXw0D�p�G�l�cG"�n�x+�o4D�������x�̍r�()�6D��ec� >�bQ!�'Ur�j�8D��	db��'�5��S�lRH zg""D��X�Ϙ�gK�u�S�, ���^C� �:���W���"�ݨ"��C�	7D $i��/�#x��Q)M0F��B�	�2������O18�����ɕ"[�B�)� *�J�� *�嚏2�;�"OMi%Ȟ�w���FO_
���P"O��PъL��ҽ���_�"���E"O�II�J�$�e����;$RA;�"O(���`��:�5!Ư�$��l��"ON,z$�ÒL���CdC�Z���"�"O(�д��o!��e��.4zx��"O��ѢH�sOXa(��~Rx}hG"Olpz"�)C�>=���M�B�Je9Q"O�LY���7�0��@��"���)E"O����B��\���i)"O�d3�M Ec$mT�R*�I�g"OV�	��[�mҬl*���e,f�Ї"O̰��B#�X��%0jP���"O$��4I��z5�S�8+C"O4lj3,1�q�w�OYXu)!"O\����#�����$��B�~��"O����K�\a�lY�-Gk���$"O�d�s�ͺ�xB��&OKn0 "OF=9�h�9oȼC�6^ږɚD"O�ᒅ��d[Fq�$%�?bZ�*1"O�ܚ5��)	v�a�fHLf~ �e"Onb�锊�� �%M����z�"O x�(ٴ-��a�$�=��`ٶ"OȷߧpY豙@��:u
�P�
O��ㅕ)$���Q�F�.	�޸1���'_Z�J
�'l�[D�GP*��PEG�5����f��DV8�d��"+�4�b��+;�E���)X��"Y�@�ݏ�x���'���klϹ��!؀�|�̄C�4{��'�_�8s�p)�ď8��%�}g��\�|�k$g���1�ůM���	�GC$v�z�;U3O�dZ�BC-OP�f�r��*q�&D)6�$Š>j�E G(�(��3��*$�^0y����Jt��=ɓBQ �N�W�7��$�R�w$׫O2r���6lN֐-B��*L4~ ᤊ�vx�Ա�G�56�D�� �
�a`P %�Mt,u[4}�ʟ;��|����*PAc�k���;(r 1�EB'�myu��R���ȓ)}g�}P�\�B�wxd+iK�'�{_�|���4qr9��65}�A�weNe�6kB�١!M��%��P��%&pʱ��ɣ<���ڦ��pn��!
z�lJ��@#�l[�h�$|V0���J&u�(�q���@�P`��U?�kW ��'��1҈VO��A�@�-?b-	�{E��,� mQ�ӭ>
h5Ir�%0Z���ݱ$U2��#���1- ��#D3na�cEÙ9�����'>����	0]���8s�ܗ`:l���8/��	�M�p� I�>qQ,�cvkPl���B,@��r�ǅ���4��G��S��"���l��5(��;�㙤<�̱EN g��	��5�tQ�>Y��Q@�]An\�뗀���uW��D��
Ad�	ƥқ���"���xo���D�,���O�䈲�ђ2��h	E՝v�L
q�N+>1q�I�f^J�	��l�K^���/��̽u(VR��D�&�$���&u�a}���O�ҽ��DO���r��7���0K<}�Րd�*a0A���j��˓N��H��2d.}�sʝ�FfRtGz��'_|��vذ�,����0#�E�0��i!���3�]�>��e♕z����'�-C����}y�-� ��ٟ��&�/�z��7�^ �����o�o��j��	�g
�db��O5^���L�5n��B�Im j�3P�S8�"(�����t����V��� ?"�qiB2Y na(WH�|�4�E'
�`O�ثt�n*�hRm?���'���ء^�fo����'��uPf 2vX�<,���Uf��ht�@W�� e��-�B-,O���"�.uq� �$�OP��q�6|V����B�|�X�I�8DzS�����z�j՝4F!I��Lr��a�'fP��UF��,�P�f�J��2�'�NlA��C�B��'K�v�ʔ�7�\|I���;lXp���}��y+&n-n�!��_�f��	@@��+Ey�`��Y�H���z����@�b�獷����������w�I&_�����/B4X�����,�)/(���R'\���2Q%_�k��E�ǎx|z}xR.�-]����ʏP�p����Gx��e�M{p��+P+�'�N���j+}B�֊<L��'n.̳�%��Y,�<d�L�V\n�����=9����U:,�����b�n,�ēE/R��A I���lۂEHdtS,Ov�{��Ĳm5���Q�uh8r������M���� ��q�`B�&�����M�+萹!��'���A���}w@q(Qa\/A�B����ЀV��,�甆��B���O�
x��'rDu�Ol�'��q�HE"'P��6�I�~Y�M���"��h) ک�ħ\oRY[g.6錩�P�\0]И�':ҸcfnC&w�~I��ɮ}W:����G�=2�����˓{�04�6H�0UoF�c�K?�ӫ7&�	�u���x��[��]�X����)$bfF���O�M!�G��f���	a��U��M�%��`~��`�'�b�	��۷IU�Ua�b���O��R���A�No�横�Ib���DˎQ�XЕFفP4d����5}"epv��[c�E�:�P�O�4@�J�/rt$?5k6&���ţ1E�Q���cSB�'�V�J��G%(T]`bf��O�W$-g����\7���1�V7@��ɹj 8��#�mx����:0��e	����d�T���<�����=M�Q�mSn6*���di�4����lM?��RfVt����NCr�<Qa��n��͙2�6:�J�hf�):2��։^�<�c*�4d��|�<Yv������:�iB�v���:�*JS(<�@�S�(:|��GŚD�Va1&�3ip�*�BC�kpL�q�-5�O���K�{�,�+#����̲��'��b�bG)'���ϓF�(�F$����ф�)(�z��ȓh�ly�CS�0�ْ��j�0��=A�b��[�]kF룟�� &˒7�/݊����:]�\�j�D��C�Ig�l�F̝�!#� �&
��86��Yn�'n��$�7SЙ��.ʧ����,^�0�gưI��g V<1�!�dV /,�9C����XX���[�)�h�Z35�ܭ����Ui��֘#=V�B M��ᝮ��\SC�}h<�jQ����҅_Up��Hc%f����k.���.�)h�Ȋ:�4��77��y�hJ;�,�Iq-�w}��@�Q��d`)0�<�UOʸ�y҇@�*;����дEҼѫE`с��Dײ�˵�PJx""���U� ��`�ĝ^/xȈ��L_�<�@�
�dD*�!�&&�H)5M��(��c��>9�>����I��%��0bX����,J^�ݫ4O�DK���#��d3���e����g�K�'��i��N7��>2ɲ��y ����L�ցi�Bex�|� O�ڕyX��!c�Yv+"�:-��H���yҦ%Z8t��g�1 e%��yBf�� ����Ӆk�l)3㍓�&���R��I��B�	�W�PHF�G�OO�=p�1b�hj�*%�� 0`Q>˓x� Q�#�\D�-[�#!��ȓp�H��b�{(|��%�I�~���R��{�(Ą|���+r�|T@�ȓ{�ۧ�yMP��JϤ��]r�'�Fe����_����.�h�'x�Y´���,��Y�A�`��'�<ō��x�u��Z'V�b @	�'�б�0.�a� 1�ݕ4���	�'s�I��KB��ڡ��[A��
�'� U�T�H�V��L�\VC���'tL��� J�"�fWVƩ��'x �cڪe~��;BַHd�T��'�z%
S�TNj��!���K(���'����R�
�@��g9���'��B�I�&4*!cڠ�P�H
�'�pb��S�����-��\EI�'�����ӑP��pq`,^j�x(�'N�}���wIL�W&�#~?le2�'+�@å�{oZ��'&�t���'�*u�@���f��c���A��p�'����r���8�&ʌ M����'�8\X1���N�֌	�+�r�'�ܹP�@4`S����j�'���PoK*p]�8R��&ddax�'	r���G؊=�~Y9�Wcv�ݡ
�';^�(qʑ�]���P�F.S1�+
�'�d}A��ԅo�
	��DGoԳ	��� ~�Ku"�9[���1����1`��z"O^�cI\mO��U��~sJ�q�"O�(�'�X�[���㳮[&eP�y�"O�$)+T=J��US*��7S�EJ"O������L�xұLM U*<�U"Oz��"�ɿ#�l�:��G�sW�i	"O��*&��t���#�]Gt��@"O(�*3�ӒI��Q��)N��w"OPa� 0/@�(�l	g��	�"O����	�r}��#�֒?�,���"O�k �K%$��(��H�c��ɱS"OBP���%��]b�JH�д	�"O��!��$F4!�-[lz|�g"O��:$]�p�lh��L;�*O�
v��F���y�,aa�'�����=Z���7���{�$�Z�'�а���ox,�Waߐw&��
�'�0������-���sg�K<O�\�
�'����P#��{�t�2�*������'�Fi:�\�v�vIa1�K�jj�[�'䊕�� 2A٬D���P�e���''��*��n���r��-,^ܬ{�'��٨3��	�͸�"J�	��
�'ނe�ʚʞ�#�bE�Uf��B
�'����W��)�����'AT�	�
�'3t�i���{"$�p̛��6��
�'��	)F�E�DWt�`�A3��)��'�0c�N_^ظ���6z2���	�'�aC��A��Q��a&[ภ�'&�p�E&D�D���g�d��L��'OV���^�a��QЖ�S�d�r�j�'�x@�f�3F�(�e�W�I�
�'����V�2��E%̓�A����	�'��I��X����4��'(��K�o5�n��M������'��ᨤ`��v<<��
�b��!�'5@�Q�K�E�F�*�O�f��P��'+�%�@�8��y�	@ب:�'*��(Z�9b\`����<q�'�N���9{�
E���b8*�ʓ"��ɵ�Zrԑ����9G1,��H��y� �*of�Kr&1B�Y�ȓJ�+7%�R�|PKG��/J��D��N�2��H ���@3<"L�ȓ|�:����ֿ��p��ۨZx�ф���`���$6|	b���_��P��R��y "lC�_��$*�ft��h�ȓf}��j����;�z)R��L�pNX�ȓh�Kٍ�8ڠmڹ-=r���'4D�8;w��6v@�R� ��{�R����>D��i��C$N@}�k�&M� ��(D���֋ІX�fq
0����+D��Q���=���矃t�xmz�)D��KE�82a�t��?e��ɚ�o3D�d#"�T�R�N7������3D��yC�S�*Q�=y�)Q�T�)���3D���vO�49PAP��Na�r1+�	-D��24C�S/�����[22�ܢ@6D������ �����
$x���5D��p�D�7l
!�Q�0�"W/$D�l�r��'��ڃ..4Zن�#D��@5��G�Ѐ;�Z=0P�m�G<D��XV��}�\���q���p��:D��۰��C�Nh �[ Bv|h04D�� ��Y&/--vAP�B1s.��"O����F��,Q�`�7 b�i1�"O��W��@��,�f�rY��d"O,���D�5:7�E�Fh��"O��p�KBH�WkC�2Ht��"O��s�w����q)G�I(�1�"Or$��R�� �v�G�Y�:�2"O�)�Ќ�>����g�[�l�R�"OV�;4�;+d�a� ��V�9"O�`��/�/j�D��S(�/�]�"O���1#\�<��B�40M�Q"O0 8�@A�e�A	t��<,,C4"O�ٓr]�A�����!_�h��"O�HB�#ҮJ5��G�]/�̐��"OZ�ꃪ�$OC�s��ɸ���"O�<�2���T6f��foU0<z�2�"O�ɓ�3-�	��P/J`PJ4"OV�X��'��03�� �M�%��"O	���Ӯtn�*�L��wI���"O��xa�[L���Z�,�7�0�R"O e���1T�YA�F�"$t�ؐ"OZA��e�	�05�tF��u.0�	�"O⭃AB��ҐB���q�N�y�"O�q�ԧGu ����-3 �H{u"O�E��GҁQ�.)*��ֆJ/����"O�	�����4R8 ��ӹD�8��$"O8�CUƏO4LٱĎˊ"�P��"O���,q�b�#W�	�t�����"O���i��aY��Ц-��B����"O����B�	L��t  l��)��"OB���B�f�"h+Ҏ�5�^<KP`�nI*P�=!���O48(�m2?�ӗ�4��y�"O�����P�D���'ڣb"��ӹi��@JAʘ)S}�|��V-1D��c���ە&ħo����� Y�1�I0�y���8M�*�)rJ��_k���[��y2.�hj��3\U���eR�ٸ'���iG�u_�LG�D�
#U�8���lF�E�x(�C��y�e�a9T�B�ΞF��i $� IRn z6�U-���,C�Q>˓|L	�DH�M9b����@8[MT��ȓd���Ņ��F �V�:WVذ:a&�ZPF�8AτR�@�\!t��B���~��0�0\O"�(�!��v<�(�'�	��CDA���S�Lvd�A�'#� 
��]�S�OQlMCt����,X����W�~!҈{bHW*F�A��b�O=����xzmPBJ�&(�d�'�����$�L�yK9Kd�1C�b  B���Ꙓn�J��$暳��3$��2�Z��ۭ�&�TnN�sd�ئo��E�F!8�c��Ȑx�H�&z��р׌���U3e���M�d������O�9"7��.w9��=}�OR0j%�V�2�'f��#����p`a(b�>�����0i4*
�)��A�a�CN�|iRp(�@��̱�OZ�8���O~l���*߲��L D;�qOl�3f�/��A�ՙ�x�ɕaCP��A�@�N�!�A u�ay�f�7�����Ԃ)i�=�&��p<yS��;P������yz��9#M(~����S��>g�z �4%ٖ A<���'�&��	� +���\�nHH�O�	86l��6��Ű�HP�W֢ib��@���hp��R�z+�]z���G�݅ȓv/R�	v�I�w�չ+D#�d�9��b�������N(±��X����'Z45��H97+^9QO$W$� ���{^8���եn�|��LX�8&Pܪ�-H�z�Da�&���ϊ}蓂D/I݆���=1�6��@G�9Z� ���}�џH��+� ��8U"� x!��ðͥ\���3�מv�X,`C�6�E�O�H�c"D�-�Ƞ,L)�~��R� 
�&	37U�ĻA�D
/T�Xqg
#0j��>{���#�� Ss�Ջu�Ux"O��7l=r���1���'����� ȡ|�b��J�P^0�(�/�	l
�O[4�$��"W \	C �J�̆���1�<�O΍�@=� ��8��_i������22Aĸu'������[�;<3d,<O��@��8�QTLڟj��=�S�>1���>׼�,���P�#`��T��O)LZ8�F��~��!'қ̾8��o�5"bB�W��=!%���6$��LO.��|�'����D��>����<vE\���`�!���ŦqͻEG�S���w�@T�?>�4��	�DB�A�lE�	a��>�h�*�L�Ӷl�6ĘP\>Qȣ�F�#�Π�ImD�n�I����1��'3[.@�r�"!�f�?���*S��L�@�+�)��V
��su��:�)��&<]�I-,��A�m�ayB`Ġ�8vL�/�B3���򤘰� |@p�5ID*�s�����%&�Ѝ�f��JT�M��Q�lm�dD�{m&h�����@'�+t�Y�P�
��X���_9v��	52V%���
�⩣�']*v�铨ywmлpVT)6G��r�d ⦑��?q"�P�T�����D��r'�؆"R���EZ�Ze��Ato +up��'��h+�U��O�6 ��T1&r����M�>"y3�I3PÈ�!#_7]r:��$dM�|���OB��f�0]n(��`�B~lͳc��@V�',��9��WR�}2�#�6jH��/O^A�)Xoݦ@�o��gi��>���υ27F~�iVB�h��Ċ�+٤O��C�"OLT I�"ؤ,�AgAL�@W�E�G���=Op�dO�s�1�1O$'�	�z5�0%�[9QF
O��q@�8d!���-�t���N�@I �b��
�}y��9d	�:eP*,!4��=�`�뉔MeyBD�,Z>��ƛx����lU�"4e�! I�E&!�5�𱠠gI�,��\���H�bqO��@D�0Z�Y�'����SMC�d�̇_r����+A���S�ˁ��y��%/����(���#C�apL�b˛z?Q�F^�0����)�K2o<����ǂU^��0�|C䉱}�r#�&��e�7�֙
"�S�J�63�a��'��@ ��OU�Ez2i��!,<d�6 q�j$.�$��xĈ~��؄���r�Z�ȍ�	���A�I^Rp��	�ąpVoF0p�x!l� ����$�z ���� ���ױE�Ш�`�;w��a���}�!�Ɩq����A+U)@`�q��C�"#��'b�m�%��!&�`dE�T�V4�X�X�O
�)ր���a��ybH��{��"ۇw�N��D�i�p!�g }R)�<���!�D��ț!4���&ӸKJ�Ɠ)yt�%mC�kR�a�D�<`֧A�]�"D��f5�Ob����>N^ŸgB�,+p�\HW�'OZш�-(u�X�'~�q�范j0�`� �`��)�'��[�%V�o8 �퉡�h�Y�y⭉ �b�I#��7nn i�N�	iJ���Êd�B䉈p�]���Ē6�{T�UR7�:�I)�Q>�#�μjq93����̧��U rHЧ� >B��`�_^�̇�K���k�l?(0��8����ȓe�P����!K�X�  �I@d8��7JdmIbɐ88(�L0cJ�4hР�ȓ��*1�'r�����."Nȇȓd4PEZ�H>�m�Q��y�F���f�晫��)Z�咣�E�F�<9��&}H��"�]){%�	��Qr�<��
�c��� �)S�2��!���Hr�<Q���/`�Hd��O�s@�ћ�/U�<�OJ69�ѕ�E��(��Hz�<��A ��Er��8Dz1d�|�<J#e�d�5��>!�x}Z�)LB�<iW��{��=1�����|-Q�ȓ#L����ÅN*�1�Ũѕ!� �ȓ1�t���h�!i��)A��nILU�ȓ^}�lIAk�-_=�|(�fR�>��H�ȓf:V9{'b�9I�rX��@_�7��h��r4��o̊/��u	�����̄ȓv�8A&�,�d�s�� C`��ȓ�j�hׅ�'Q��j��Q�ȓR�X��h�0����,P���S�? ��%DH�6������!��m٣"O�p���"��d8r#��~��<�"OH�B�ʧJ���{b.a���"O���vGѤ"�jW
�����CO�<�w��k{V,�f�Ça��숇�H�<1ׯ3[�(y$�Q>��]�㦕F�<i���� �)��D�kgȍy�`KB�<9t�	:0�Z��s�Ƶ��ѓ�Lu�<��Ӕ/��t2��3m�bĸF�Jp�<���'lT�s3M��7X�E8�n�q�<��.B�-b��m5l��h�<��j�8]�Աsǎ
�up|�c�-k�����f��P$ڝ�f/�i��7(����ec��0D�|RC4\$�����K�u{��9D�p��Jؾ\��	̕��A��@;D��"q���6���ȾcZ���:D�ܑdb̍=&�hrT��63J�iE�7D��B���/	�pjv"��<�z�k��4D��8D@�nBx����
z�n|Q��&D���e��p㾵ئ��=|��H�Bo(D��c��j���"lA�_H"e���$D��`Ȍ�_�(TaO]
�җ)8D��:tKܤc�t�+��&���G,6D����t�Vu
5l�2a�|�B�8D��u���N@	9s	�)!��{��#�$��1�JMG�Č�; �~:��Jq8%���Ǟ,L>��P�N?��	��F>�`i��'}��IS�**@�j�G�K�`��U�G�D�4���"/}ܸ�>E��N(w�H� ��Hb0����ˍ|z��İ���a���Z;"Vؙ'
�r�f��")n���+J��*E�R��L<%?AKp)c�����E����J�+=|O\ &��m�=6���`�"G}�A� D���a�ВX�-��
ߚ^�4#U� D� ���8.���G�0X�6��b�3D��� S8 �ҍJX�8@��Չ}�rB�I(DT�����K��n��դT|��C�I�<*X��j��q.�I�'#��C�)yT�aH�x���HU
��pC�Ij���+������i���u��C�ɦA�vQ����K��`�.<-	hC�	�|���چb�Mm(�IsM] B�I����0DNC��q�(� Pp�C�	&'��q�f@�]�>�4`]�]�C䉙CO�� �G�&&z�C4 X(c�C�I[��8p#.��)��֦gdzC�	�/\`���l���YS��F/�B�I�7�} �U�(�r]�e�]�JB䉟X|A����\/x�7hDq��B�&��KQO�F��ّD �4Y�xC�	�s�`}+��O�Z����p.�)@C�	&(>�M�F��L65)2gJ�B�C�	2)�<� �E�
u�Di�h�C䉏2�%�e�.e���c"ʇ�B�ɟD�6ȸr��^$�C�#ͺe��B�	*�bfB�=����BƦ�B�	��6�r�j�Miv-J�L�)o�@C�	�D��T�QǰS�E�.ٜ��B�IY�����ߠ(�pI��X�6?�B�ɏw�輑C�JQZn[daە3A�B�ɢ`��s%гCA�1q�� LѨC�I �*$�A� -�8��c�ۿZG�C�F�	a���4[��	g��>��B���
u��'�l�pU��=�B�I3N# �hq�<��f�P�-C�ɵX���VB4b6��#����B�)� ణ7��,`���*��ޝI�zE(r"OV��`IW�1��k! �,�U"O�Hr"��
��\�׏�+1�>Iaf"O\��`E����#�J66�V���"O-��@���%�u�ɉ%���;�"O��iC�ʄsA>U�?�A�"O@�2(Y}j����lL�G(��"O�� �&2�]��+>]�| �%"O�A�����'�<��(D�� ���"O05��@9 ���ӓ���[�"O<)"��V����@�T7�X�"OX�%�P�PS��7�ؽ�	�'�.\YD�B|���"�Gl�ZL��'>z� .b�4���E�{ؐ��'���Y��A]���D 1
֠
�'"E�3�8C������uЪ�K	�'�Z�H���>yT%�"��o�JXs�'�lX��<hk�(���ζ/6^�9�'�nuҡ#ΰp���aB�,/7t�z�'��p��I��.+�Ɉ&� 0#�'\�q���/M����K����'�\��dA O �x���Ozp�'�=;���s�6A��M7c�L�ȓ(��Hsg�4���Cq�������C�dX��@K"���S�	u&Յ�=�%� ͂�9��Y6UTo����,��Lإ(Y�q��Xe�������j��"Ĉ�1��1`WC� |(��D�D=���+���z�GB�d]��N��I���)����(PP�ȓ-$�9����'P޼rU
ŷBlvՄȓ*��a���x�`��!ul���
8�1G�/$H��0t�E�#���ȓʦ��
�&�q e%��DNbԇ� ����Ҋ�9q_x�F�<)���<�b�#i�xwV�7*�;!N��t��|ГiEq�be�&
5[�2��^�d�!�L�T�23m�2?�-���F� ��Ⱦ'RŻ��߷E/d���4��-k�M>ny�a�o��'ɺ��ȓ_7~q)t���N���[��O��za����0;��I�v�H��A���>��^��g�'WeP�;��W����c�<i \<t��h��ݶuqK�,��B�ɪ)o� [�ծu�j���S/n��B�I�&�iq�ۑ@�(}HQɏ5QN�B�	�_�$T�� ׍J�R�[�j��wҴB�I�]�lJ��N��R��D�߱
,�B�	/ �
�{2�?Pxh����I4\
�B�I�Z2�Q�B��%���H�u��B�O��=	.ϰ7*�Ţ�b��4m�B�Iz�H�W�S�UDT�� O�>C�	:�xY
1#�Q$��A�¤_�C�ɥ
�H�2ǋ�4ytJ#-�'4JC�	�@֊���.\��������C�I�B�bJ�`C�y��D7,��C�I�W�ƥ���7��ܢ�ʁ�ZlC�I������嘾-�Z|����4e�RC�-#%.0a���3?���m��<(:C�ɑ?��IC������G?M�C�	G�p�� �ݥ�mS�2��C�I�]��L
�@#Y�,(���
]ބC�	�xn�=Ia�$jVq:U��Z�`C�	�
��'������Q#�B�)� ��z�*:xK�k�.ڟV�l���"O޸��%ĻY�� �tnܦaݎX "O�����%.�#�õ-z\�Bf"O8��d��F> *��֏^[6��W"O�`oԪs�ʐ�ᤞ�sV.!��"OpL"'$ƬK�\����͗<"tЛ�"O"X��܅Gqzv�Q�,6Q:�"O^��NM<!�h���A�� �$�r"O��rA�O�0��r� ��"OD�*"l16}$��*�i�����"O��2tM�OvT �F��ur�"O�!���p0��/G*��"O��JUA�xЉ&Lʬ[]��A�"O�d(�၀F�� Eˇ8X(�q"O�p�K������N�tհu"OfA�Q���)�JxB�R�I�p#_Q�<Y5��}��]�\�[����I�<�,<2r:����J�D��q	�F�<"	'O�����B�=�|#v	�A�<���Eg��t���9ZP���E�<�\y`~��@��>^ಬ���F!�čZ�����M�@��c/T��!򤈳rj�P@�L�T�VM���(Y�!�D� �h� �F:u.p�0�Kȵt!�!��#+��
��(���7n!�C�̌AՏ�]��q�v,U.Z!�$�3h_L��f�����ꖽ�!��׵_����ՇJ�C	�u���b>!�dU�Z�$�2� �(u�!��h��N�!�D؅Czr��22&�1Ƈ3=�!��M�S�x�3G�?O~�K2E?eu!��l΁�4-I�Aa�X8d]�xq!��Y4:Z�}��@��lX����B��=�!�$4&�*dV*��!P�⧢�/�!��N����� <N�$�� A=�!�D�$B��ҍ޺N%@��2l!�d�4A���Dl͎d>$��BE�O�!�ҏC5:p"�� ak�����!�=�&0Yb9}6��t�M�!�ݭ0���#я��I�D$'�!�R�(������y�.0��E�,!�0(N	�v/�J�h�V�ԂD!��_	��Aa@�=���2�4;:!��ƈ;�Z�����H��(c@@0!�d�%:hx[�埦\��Dp��-z*!��QUF�}A��3z�L��.�y!�$B�|�t� �<�r!�0M�9A�!�D
/[Rd�x0	D�&��2Q�Ɲ�!򄃗L�>�D�~���R)�3f�!�D�ia���J>!X���F�_;=o!�ޜlyl�$��5<���2p肬2�!��K�6������
)��9JG�1D!��L~�(�P�u
,i�`�g�!�dE���X��F� {G�أ��$�!�dX4�A{`ĊF$�F.�*�!���%�~�x��@0ta���:e]!�D �GY�飢j�g�lk����/6!�DF�J\d�� A� L�dK�O�!�䗒^��Z�ݔU����q�!�U�:�XPI�ÅgB|��
�$�!�d�s�n��ǀYu#Щ�Y���؋v�L��5�5�ܠ+ ����y�˒�wӪ�ziП3u<ݳ���!�y�ɗ�rQ`��� �)0Z
��S�Ƨ�y
� 쬊�朜Z�r�z��ɚ?
6��V"Op0C����LTyv�)2X
��4"O8�P3 зa]\��r�Ǥy�d-K�"O�$�tF�7;h�q����(M�uZ�"O��cIz�"0�W�o4$��E-*D��5➍B��ӂW��(ɛ��;D�p��V�/0�5�6�ʏNo\�Pd�:D�0G���7�xx��S�JN`��"�5D�P�^04���0ݖ�D��M2D�8(�+I8fk���b�,�&��A�!�dU(�6Y�M@�RO���7�%�!���<O8ِ'FоF۹e�:&�!�DN�C��g�$Q�!��B�V�!�$;Wh�.�|��K� M�!�Dױ�$��6�ݰ~���Ak\�$!�����ؠ��ل�J��O!�Ɛ=V�������$���@�#0!��P`FԿ�L)��f�)wN!�R�6:I��Cэ3͊�
��E7�!�]�}Ѽ�ʤ�����LQRH�b�<Q�IG�N�x��̒Z���@��E�<Q��,����r� +`����Az�<y��6@��d[�iÃAsFe@�F�n�<yg�	����fIV��!r�<yT�F� ~�}5�� BLt��g�U�<qTb�
Sr�����f�X���%�M�<��ߌs��Q��.\9I��Q�&@]T�<���[� m V�Է47����bZY�<iaߺqT�񈗪�U�s��S�<qg�m���`��&Ky]�A)�H�<�VN�+X��(KA�1��ʦ�IH�<�
|}:� V�摈"
G�<��f�Di�C��|�a�kx�<����y��{q��A��ՙ���X�<�愊���!w�O�q0e�Z�<qv�_�	�8���;/D��`aG@�<�F.J&�yɠoB	5�H�*�v�<ї-P 3f�rCK��!����Z�<�1�
:�B	��# bd�z���T�<���4a�\*�#]�r)0��dG�Q�<���S�g�@T�e��Y�LX(�� J�<��4 8  ��I��"y�*4j�
=�`d'?㞨zd#ي�(\*�(x�,�:���m���B��3,_�=س�"'�����M�(?�]�����<��)br�'uDY��GE�l0P�	�+§Q:���<(�p�ъπ�� ��y!H�?��Dz��L=�@��ȓ^���Pэ۴]붹�t[�i9�ɥO�ecU��6��O��p�E�!=��$��B.j����'{T�4�@���r��5Y����
�'*���'EŹ+̀qM0H\��
�'����Ʃ�T�|�kU�K���8%�\�n�nԄ��b+U��뜔>�����N�2a��ቷ_��Dƀm�h͘,j�j����#�K�V�B�,>�{C#D�\������v���Dh�bJ5��ӧ(�� ���2`��
)+g
��}Y�!r#"O�iÇ��!:]6XYC �ZM�Y(�jv�� �&��h��J5���S���I!h@�:c�л9���
�V��H�UML_���Ԥ�}8@ �uǍ[�Ό��I d�-Kp��7H����AE,���?a��A�9�8!r��2��_�M��p';�J��A xT!�D�/��lI1��-R�|p�aI�o^�I�,�\E0�'��S�OaN<C��>~te��
�1P�R��
�'N�0XQܭU�D�Sl��¢�,}�'X�8�9r���{�!M��Tqph[�@j�5k4/K��?YӁ͌��XaDXM�b��J���@���D���d^�1[6����Nle !�.�ax�i�>^U�d:p�|r�=M@<����ӷwʄ�P��y2#�i6Pâ���	���j����	'Dj5r1��ɒH00py�LƻFʑå��7!�@��lDS��H;Q�U)���$�!���0&���\�_�Xy����q!��2NZI����YT(���+п*/!�$"F�&��P��yBP���hZm!�ă+=�n�h��ɤg��)���K�!�D��UV�J?��s0��s!�Z����Ε�	m��RTkV�!� r�8��3��+,B.�j���7A�!��+d��5�nY�9F���FK�_!�D�r�Ly"��:m1��!�lO ?l!�D�<j���Qe�.�P:�l:!��F�V��l8��S�ߺpP&ʙL!򤑸���dAw�V�*���/ !�D۲Y~��
�|���q�υg'!�d�+B��Y1A��a�x�(�,!�ĝ� ����#c�*�2tL�3>�!�d�R$���L�lpj I��X��!�DA-�и�o�BwZ$�� �%1�!�,oHUK�ɚ:H0VX��L�Hr!�$Y*1��pq�䗃h'ʭ��g!��`Ԗl�&��$I�����C�*A!�ˑ@��wO�6�X H��=!��+y<]EI�=�Q��D�F!�	�H�4y�r�"B�1�@KT"!�	���e��*�9�@#�-D!��
F���(u��zߦ��C�L�:D!��S�l:�p���k��#5��<!��HL���R>0�ّ�.>!�$P>+2V4�a�C�?����L>$+!�d;Q��`���ݢ/�B ���6i�!�M�SR\=3@�&̀��5&��]�!�֓��I@��$����E��F�!��SW`p*1�ɱB���
:�!��[
C�E�����(��1�ɂ_h!�d�Ő�	�i�`pV8s1d�#]!���Op6��tE��KJDy�'B�-bi!�䗷^��x�+�>6�qQA@9i#!�dE�M�@���)�+��q���d#!�WD��Т��e�����ơ5!�dM*2��l��m�Qu����a"O��+P�,�
��Uf\�J�r��"Op�(�=��#������T"O����4�0<s���t4�Ч"O����Β]츃g��l�F"C"O2B#
j�A�p�5/�����"O2�FZ�(:L;EL��!�r��"O�@��e&,D� ��L/#�б&"O�40�c�U7j9��kR�H��U�"O$i:��
è�	�&S\<J!�� ��xc	Nn��3M�#`��"O,��D$� y�cfćY@"���"O��{%�ӲP��9A3�͇"O�"OZQ%T��4���U�W��]��"Oι
�*	 �ؼ�	��J�Z�8�"OF�١I)�p![�h��
R�u["O���V��.��@���N
3{Ё�"O0!`E�;��c�*ypΝ "O(�
5�Q�f]H��slЏ � ��"O��H$��R��	�K�-K!|�Ss4O �;�L������(�g��H���AJ�!*8��F"Ox���n^3젤
²X�i �_�LX�#ҫ
�f��I�K���3Ñ�i=�c-�~������<�d��	\?!ApqHƃԋ>�bl
��ڻ3�B�
�'�\�ī�7�2�`Ġ�|r:���аl:A��)
��O�8PRDOۡgH� S�����KBh�<�Ӯ�*`bEZD���	�@��GM�䦝�"EM�N�\H�>E��4�� :R����8�AOէ$���~��{0��:In�42B������'e�U"�E�?RT`���
	#��J�8�� k��#����՘;L�!���!{0d:w�Ć!�ܑ�Wa�d-Ԕ��'^����&{6@˲��(5��D#��dZ�,������Ӽ��OY��B%"P�cK\|�1+T#�T��'�X�!F+$?�I ���P�H��۴�.�EdƳ
>ӧ���F��{��X(�A0E28i�\=�yb��O0����ޘgf�p�W����D�S��c�EK���<0(T/Ki�ȫ ��,,U؛��V~X��gi,
��i�Z�]CďF�T�˧*�`��񤏥�4S'"�D���VQ)P�ў@�#I�5�ЍD�D�ĭPƮ)a�"G���t�Ī@�y�⃿, ��%�y9�@��%Ȩ�y�ˁ]�E�=E��S�t*��E�wq@�0�� �yrc�.��� �� dL�E
"��y��	�k6dxQJ��eV�y2a�D��y�'ˤL&�U u��4\�ތ
LK�y�ҏ:wN��&͔P)r ����1�y�PAFQ#@)7J����t��y�bG�m���-D(�'nƹ�y�-X�9 �&�?�
,�G�.�y�N�Z�Pub��AKz�cX��y��Ѻ<�:�
a@�*>��,qCi���y2	�!� ����42벀�gn@&�y��>��ܛ�F��&#�ia�d�%�y2l�J6�-`@�߻�����ߧ�y��C
j������=A��4�5�U-�yr�ͻ_��)'*<�\0��	� �yeΣ�6���%�(�`��C�=�y"@��Z�qrU�=)�LHHSL���y�B�h��<{����`8b���y�I���B�r�f-l�b�5���y�H
L6�0�p��"�1�R�Px2I�&��402H�d���#�O��� ��"q�pI�ъ?кM��Qo�3�	K��� ,�0g\����F&ː��DO bt�-�R��Ox8y֬ϤM�~�Y�F<+%>�ڰ�,F0�����O6ȓBèپ���@v<�6!Z�!�v$E�a�剄idX@�Ț���]"@B�BG�Y����v��q��$ �nS!<9$�@���r ��+�!��U�7I(�i�W'y��3(8T�TAQ���b�d]҇`��:���C5�ԗ3O ��'���I4E��yG��5;Q��a��S��̑�C!�2"�$nz�m�V��	����P���6�f�1�glN��(��+� �;3�V2~�]�&$�����>Q���AyȀ�@*A�2k���zh��|�AG�?i3���h@aB�"`�)��7(�&�1�eʻg68IQ��.#�����RWV����R��a{2!��}ɨ��A!�-���	���V���,
8�M�2��SF6]�+y����Q!7.�ذidS�R�ݸU$�@���I�9	�<!�'��V���;� ��U��T�	�q3h��bĤ �J%�"(Q�I(xz��\$RdZ�/T�)�U��ყt;d��O�EQ4�[&
�� �����Ӎ&N�a���u���|�kS�FƏ�ZH��̹���7@�(���9ZL@'�
� ��yycD��
T���䁀w��pi�1J� � ����'����G�NXځ �hΥS���c/OGu�4�,OJ5��� �i#,ҕp*���U!+������	m��+��K�.N؁� � ����F���Gr�dۢ�]x؞8"��ә&��`űU�tL*a�R�p�.����,	N$;��� �;שR 
�� ��V�z6mP%��DNOU��!%�մ/���[1����<1u
U�)���;�F��y�kM���G�؉-�p)�@��f��`�����<�"��
j^<r�+G��!ܨP�<�1�rA�#������,Ph$qA�|�\(Z|!�$�2.�K�bU�rq$�	>���!NJU���׭Gd0����>���� f�j�(2��i�,Dz�#��b#���ҏ�6���.�%u=�ʓ�~$��O���`s�	b��'��0�
�2R����+�b<K��Z�A��83��'T��_6���J�&�%�ք��	(��B^+��lz�B�ɼ#SVM�Dú��ɼRϐ �N�p��<+������&9���>1��ưkp�b� �GY�u��e�E��:9��x���J�	D�?I�G,�fǜ�h�,�}5xi��?D��FGɐ[{2�9�A
�Lg8=R�!��ks��O�dB�B}�g�	���#��5?��$´�J.+�C��(���P�B�6~�o�!^�{Eh�  �B��'U�8ɴ��BHB��*�KZI˓���r�Հ4��ʓz
h%f�
�r�p�"��Nu��ȓ� ��Qh�e@h8p�A�k�\x$��X�D�)6�&��p���y
�!/�?&���I�c̀CA$B�Ɇt"�]H�B�4��9e�MIi \W�_E���+��p�~&��V��"�����Ͳi��JG�>$��K�G�)a���b��*(���Q���|~ԵB���(T�}��FL�\h:f	Y,+�6E�p�D�<�Tl�3[QTu� ��<�����g��a��
H��dr�v�<�c �'R� �����}1L������I�|5F��㭎>����<v%�����!��Q�P�;D���N^ ���G^-T��#��[�qOr �1�3?���պB���h�KU!J�2�q�l�o�<��(S�S��q�$��!�P�y�`�c�<r��
(c ɰ�l�M4�1�
Rc�<��$��=;д�UhG�qa�Ei�G�c�<�!�ިG����	H�dE���p�<�7���j�´*�k++�P��jGo�<����"�9�B;!��dB�Mh�<�ae6G�v�bG@�P����	�i�<�B(Ry*��6%q�	V�k�<!�����A��6y`|�2`�O�/S��a %�'2']ÁׯE�<���K�9����vH�ik����I�l,0�\+j�RPAׄݷD�OPXE��O^�+��T�|v5�1��f�.�YC
O��&�~L�b����#Aj p��L�	b���W!D�E� q1
� Jl�ඉ�7�p\ӏ�	~ �I�L<�A�#B�{^X�30�d��F�Ȝw;�	2���v�FE%D�8��@F�;⪔��[��BW�<�r.��7b����\�5Dj$���i�|�
xt$X 14ȃ7k@!��+nj����>>��]p��/K���f��=�B�Z3d�P���{�U�?j��P���e���"@J��?��hջ9���{��n�~�*��=/��PpĬ�8t�f0��Ǯ�0>y�᝼3]逑́�33�\��f�T�'��hd�G5�����ÛGP���"��9�����F�R;!�ā.|+dM�M�629��ycΎp>�ɴ���Ȧ���:<��@�K�J�OW.�r�:$�-s ��e�i�'�d�Q�)��i���C.zs.A�H'����y�2�����gܓe���w�>���NE���%��	�d��h0��/�D�i4���.�	[���4T}���Ga}��T�`�����GY���&��0<a�NH�g;J��H>��K�N�1d�(���#V�g�<�$FŧP��|9��P�<|�ƅ[K���{ �z�{��Ti�1|�"� �8}��8h�-M��y"���,P��	4��t� Pҥn���yB.�1����Gm��k(�� E
��Px��	X�? ��C�A���aw�����%	.8�!�D�#��@��̈́J�����S/ax�#6i,DB�|��[����ǡ�)D�Tܺs��7�y�*P�-�NL��_�2�U�������}/�d`6)J
��)�'Q��SR�"k.���V�N�>e�<��W ��	�f��> �	ׅ�U<S%�>Rn�8�X
N~�=�K-D"��f�C��V#�*���B=[�p5�I��r���@ ��,/���pA *�
|;��Z��*ea,Ɇy�tQ��F�'w�����!�a$>�I��m}V�zd/���Mbt��~�<��Z"[�J�r��:9zx�H�i�]yk��{��رՂIg�哠	�Ś6�@�jo�}�F�޳>2C�	D�a�蟔C�nY�/��J0|�'����7.�|��ϸ'th��'�1)��U��-r^����Ovb��t	]2{�
�qu��
�VAB�i�G��=�g� �O� �	�,&ɑ`�C<c�F�rr�'�b��`��'D��j��)#�\*$!B�X�Y��'����0��$2v�s�bŐkZJ��I��
��E� �qO�&0x���u�dlS Ay���"O�$���%)��Q��\�8mr�!�"O��1��ƸP��Dё�b!�A�!�d�U^H�& K>B��T����/*!�D�,���3̔�7�"�t��{
!���-oR�!��9`�L�x�J(k�!��V sC������ Qݜ�ۂ��48�!���=k�^���!�����f�I�!��WG�rTb4��!�
X�祜�!��s�t��7MI;;��R��H�*w!��N(m��ԠT�5}OPuQRk�0o!�Q+�H����~��ì��H!�d:�~h"��G5P��U)���"1!��Dm��;`��/a���!OY�!�ԯ@Äiq쟼3,M�ĩ D�!�D͖8��͛�"ɚv�@	����L�!�D�l3�q��+z�(�W�!{d!�$�WI�H ��6ib�8Z���#|�!��E�k����dC\ b�*��s�!��]nξ=��D��.��gɏJ!��	�Xm���hȘ4�J��g�ب
�!��+��O(f� K�@ �!�d> ��,�c�88��Uڣ�	�eq!��}ހ�`�*B7%D�Uw�ɥ!��1�h����Q�mȭ
�!�܇:Q
��c�^)_iR���BB�]�!�F�%�6i[f���cNT��!�=[p!���^@ā`Az�Pp���@ ��6�(�\X���'�<q⃄�8�̑Po�69��ڴNB~��ֹ+��ȟj��ဇ{Q��ad՚�H��V=q|��;?���)�F����.tF�!��X��kD~�,Ք'`�[�QP>�� 	מ
�����K@�<���"�	���� hz ғ�L>�ǦܮLåa�0��Q��>a�@Z����A�8�~�'�Z��V�L1j�X�E�p�T���=n�� �F΅P�)�'J��c �I��YCv�T1vlq���[��`[�x�ՙ���:��'	�Zmk'*WqU4��጖��y�@��6v�p�͓�j���o1�������Q���g@�{ʨ9�cJ�|�����|�����?a�D���8���:9#J�5��"H��S�`���#�D�^�x-z�'�BA�7޺&fE�j�^��spT4{��3pB4k��	�E��X�RQ��,�<U��j�z5H�1�U����*��s���G�T�B1�����P�����0��F�]�q0���cI��� A)-o���}<��IzO~���.��xd�O�bUŸ#��M�ӵi!F0��А�8:�1��P���	��%��(iR�^�eL@�UJصY=pʚҧ�6ہ+Uo}��M�i�b��;OP1�Ƈ�*AO���N�"~b��ft+td·Vj�c��@�v�x�qfW1BF�ҧ�g�i>��I5l��*�WW�Р��Y_�0YK<Iu�C����h�g�? �`aΔ�(&���ͮd��Ia�J~b+C]
��;�"���SČ-U�D�sO_'�l��]�l��{�h<yu#7?�|��'�|�0�-�6++�d�&��	V�@�*۴��a�vE�,�F�1��WZd��D�d�]+Y��Y�i�0w`d����ڜ)'ر��jޥ���I�M�ɑ
ç!#����ږk� j"�`*T�ȓH@�eڑˉ:F�!E�F}�̆�E.Q*Tk�(�҈Q�n/�����.2�ޝ؀��Z)� B�>�!��ǣ]Hn�a�G�8L�~�
P�R!�HI�M;V( �}o��`!φ�Y�!��N$��Ey�����^-S�Ά#�!�3V-�,�uG߁o�h���f�!���X041d��&|H� K�%T!)�!�ć�^�䂅 )<$�p�i��o/!��0r��$Ж+G�h<x)�*D�} !�#� e获8D��k�6P7!�DJ�U	���-<%��xd+�BQ!��GApUC�(�2MU�7�K*@!���A�$�#��2�q�	ƍw>!�J�)a&�ӥĊw�t���N��!�$�?l���ro8C� D�J4�!�d*Uwr(&�Ӛ/4�0�h�@J!��W�!+Z='�H!�B>!�<AQf�B�LL<X�a�3m!�$�^dF<;��A�s4���UNJ�P�!��3����֯G�%���u뒹E�!�$��n�.QR�ӆ}�b�+S)!��9T��B�߰@�̸��7�!�d	�b��P�]�}�S��ͤ�!�d��Z�(��e� xleT�Y�7�!�Ą�w�H��"jrx�T��T!���	���3%�1$W\�ٴ�&I!�X (��]Ʉe�).�8��8L!�,^�%*�B	 m�(r��#�!�ڮ"Ĳu sBܪC��P ����2!�I�w�ɲ�!����#<d!�$�'���
�s2L}�f?G!��DL�t"p91�:!�Ao�n>!�� #u�]ّFY�S�����֯dF!���j"�� *.$�"��6C�3!�D�4b@}xGb�&o��h�'#ߙ5(!�dT�@|`@��Ӽxg�i��|!�D�V��R0�1�t샲�J8!�d�4��!o�"�8x �ꒈ�!�$����(������"�Is��=�!��!
¸�o�#~��w���Nb!�2���H�E�$i1ׄX9{�!�\zr�Z��H( ��ܩ�CLl�!��@x�qY� �;��@H�ԪaK!��G�:��`i6�����ђ(�:O�!�$�,S��C��ءB�`19fh�:�!��%Z0�m��j��JN�٩���?^�!�d�m�8[Ɔ;��j�&�+.'!��T��k�==����)�8�	�'�am�>0hd`9�^x�'#�8�C��B��C�U	9�L`1�'�X��u���K��h���"� �c�'C�ĸ!L��8���3��]�-��'I����M� ���r��an�H��' ���GL�@s��3M���	�'M,�x����2)��Ҙ3�|:
�'�@]I�Ώ�6C�1c���!
�'	�=�EfֱV�T��T�(���	�'�^t��(?�p[�Iӱ������ x�@���[a��t��'�%څ"O�MbVDP�Y�ӰKGڎ���"O���Rŏ z&�P`s�Q�|�8���"O��`A

����A�D�	��"O&K��H�"N4B��(t�[�"O4�Pđ4#j�� ��$Z�ؓ"O$J���+Ni���ED`v�bU"O�Yd�ɢV��Q9o�6wRu8G"O��7iS���(p2��)PG�5#�"O��3!�89��n;�$8G"Od��qE��Y��`1D�,TM"$"O�lS@jU�Q��qq
y�^��D"O:�;���KX��)a�R�&U�(��"O�� ��և
�.!���1'[  2�"O�aS��H,����םk��M��"O��h䭁7���Pgǁ5%4<Q�q"OB�k�r��S�Hͷ"+�qs�"O`$�u)��k�*a�B���P�*O\帔hԐ]��Ͳ�M�l�0e�'2:Y`#�M��]آm֜R�$m1�'U��#­�V�"U0e�K;J�] �'"�;f�؟ar��G�.67T���'�J�Q�3a?X�Q��V�|���'�>u�%A�����|>H0
�'�I�B�"mۤ�.=pf��Y�'S�is����F̂�ц��	34)�'4��w��oݞLif��\��*�'<�����N�G�Q;sG��Y�Ց
�'ʞ{���<]�b�#����g?T8`
�'B��	�^F��A!���LPA	�'T2�
�6#�ؑkʴy�	�'�B�Y;#��!h㙆P2u�'s�%��'N�
W�K1`ڐgZ�[
�'��EB�%o�2�p1HӴ
$jTS	�'��	�E��(�� F/ғ}�>�b�'a9Xg�K\}�(�t��q��'v��b@֟l���[��A�e���
�'�,@�m Vz���T�nd
�'7�����H�c�f������o����'���4#)X��� ӬГy��r�'���BG�O2,��2��j\H9
�'��Уbˆw�,�I��˃fU���	�'��[��Ҷ.\���
��
�'b���	�1�|m{d�����!
�'����,ƨ�1�$�0z�X�	�'��8%��Z��$zaN�x/��@�'�+cm���t AP摌C��q�'^d�D�4tY�I��ܜ=�� �'j�����?�$ta��-5��]2
�'�f�3���0T�Z��Y�1�*܂	�'8Z(c�Y3T��scפ^�p��'��l�Ê�YZ#b�X4ܬ��'��hPW�Z�~ @��R�J*O���"�'X��$թ&(0���C�"�k�'Q�)a��\�&�����Lq��''�!!'K��m���x�V,��'�.��'�j�
��t`E�o���"�'��tQ��7w�P �*���VY��'�
=R&ㅿ���;��%v� ��'zNy�/��`0t�R�C�~2e9�'ۢx��O(-&}z��
�Ƽ`S"O
|�EoȩF���YH�9!�T
/�!�d�|�D�"�\� e	�f��>!�D5}�\x�Be��r\�� �fN�-2!�� 4`��Ȋ�?�J4�D�Ì>g���"OB�f���{�Ə�hT�h;""O�4a�ҭ T�AKa�Q�nf1#F"O&H���ğ=٠3��K5rI���"O ���Phy�h2��9*f��"O�,��k�%a�&�l'���"O4��4��#mH ��-�P}	�"Ol�+Q�1��$`��@^�LȠ�"OF䈓ℭ[0x��Q44���"O%ǝ�t�AQd���[�*�i'"O޸(Ӆ��%��	6KФU� �#"O�ti��;}�J�qd�R�H$�"O��K��Č!cJѐ2��!4	�4"O�r�L��:�n\��	-�\	�"O�҃GC:rmz� ���\��a"O��ڒ�J�Ќ��JC�"��"O
�
r��[����ANcn��"O�$�vn���2d����Qav�*#"O�U(�,]?|](d��OA#�\H�"O���T��lBD����-���"O.�ڤ�
Sz��E��"v,l�;�"OJ��f	�3A�K���j���j'"O��p�g��$"⅒qeV>�"��c"O@ � �E5iLԡr�d�]Q��� "O� �V��M���<O�a9�"O�px� 	�|�9�PL�U�R"O8[!��[¬x6M�m�Z��q"O����O�T8�X:�ŉ3�8=�A"Ox���Ll���:p�($x���"O�b�Q�V#Ux1�H#8eb�;b"O�CV�_<޼�+�ǟ!]dĈ�"O��*�苄)��hRF�0hj�*4"O�� Y�7�<)���dF�4�"O���o�~�$��`l�/P�"u"O�M��IF.q� @��l*���T"O�ma�e24^$���\�x�"�I"O­�Sf�f�ʅ���;��:U"O� �!��W�qˣ��62���ȡ"O+O�&D��m��I65� 1�N�<q���" I�4g�����Q�<�&�)|3���c�u�`�RAJI�<���Ր;z�X�A�;.^ �� OC�<�v���2Δ�a >?��#�Kd�<�W��<b���AѨ�8c�� "墍\�<y#B�.)r8 +��A�%h.I9u%�[�<	��Fr�mB��ð2�(`�F̋Y�<u�**�걃�+�+v�x�2w'�I�<��b�LXP�Q
S�0�>ڧ�VO�<��Lzܶ8jTLDB��2�L�q�<1A���gS���'��V�<e�bh�y�<���(
����wN�xZ6Kv�<���ߣ:����'
��<�!`�t�<��A ~0�$#CfJN��6&	w�<J�9�&��%O�uw"��GdH�<�&�U+N�(���>	��d�K�<��h͍tR��F�>Ke��8G��~�<��S��`�Q�,��
�*)�G��w�<Q�+�(&�؀��ش�ڜ��q�<��j�^�l�J��O(�%C�D�<���-٬#&T�1��5��D�<������A��C��}��mB}�<1e��ma���5Δ �P�y�<A�3/ń�I��u�K4�LD��C�	Ql�42�$_�h�D��vC�)� �*�/�,?L�⃄�=���"O�$��Ɣ�K���V♚:�:*c"O����C���!^J��i��"O��2vM7i:į�N�P-ð"O�*0��O�j@�n�0S�h�x�"O�\�' �X�i���6_���a"O�S������K��M8b��,҄"O���b�@�z!Yď� ��@��"O��G   ��   �  B  �  �  *  q5  �@  L  �W  �b  n  �x    �  x�  ��  
�  N�  ��  Ӱ  "�  ~�  ��  ]�  ��  "�  ��  �  N�  ��  ��  ��  w �
 � � �# �, -6 �= D HJ �P �P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'��O��P�]�۴$G��d�q%"O����bN�#K��X	0�O�#�yԮ���v+T�4z��s�����yR"?�EP���2.�R	��%z�=E��\Ȭ i��3Qlh׮�	.���<
�<����$�`�(��@�ȓ|�<��TL
!��qC!o2䭄ȓ~��s�X�\]��9�E���F�<I��^�C�}�R��-�h�J�L}�<�A0ho��+��ݐ%�]bUC�^�<���ɸ{�Z\y���6a.�Qe�Oq�<1t
���A�G��J5�-�3�o�<q��w����EQ�*@�p�S�<Qa�,��ms��Q$i�QzREY�<9�����A�Ђ8�3��R�<nM7w�jǁ\ۦ5#�E�N�<yt�g�zQ�EcKU�Z����q�<sK
 1rT�h�$��B�O�l�<!$�x�Z���U�����M�<�V�h1�\� .jV�S �G�<i��8�V�+s"[,hn��UaE�<��_�P�S��$t`�(;���J�<a�C*!�$�r4�KZt��҃�Q�<eب)����.��{3�����P�<A��]D"A�Di;c��%�ЩCM�<�B�<.�j�D�g���RbaDL�<��!İ<0��i�H�k�x�$�Q�<	�mO�
a2�*kC���[3n�H�<q�M&eP�(Q��^� ��%&͛]�<Aԇgގ�Ƞ��$~�$���s�<!�H�E��q�4�
,g�<	�c�q�<#Դ
���(d*�E�VD�9�!��6x<y�&F�(9&P��G�!�D�;(G�̨#`H�4�=�� �!�� 
%���J�]���"����"��,�u��k�O�m2�gӝY��Y�s��A�h�
�'�0	p�ˊ�F��0a¥�;[`�'Y`!��N<�lh!��5dbh0�'�,P	ĩ�$1:�p�0�Y�'����yB�'S:�H�Ļ9f`	:̘�s�0��'j�)⃬?m�F�h��
�|?V9��'��qz�aT<1��:p�A�CO��	�'�+�Ë�~'�$���;�zL"
�'��Ə�|��L9�H�7n�)	�'|RD1WA˞_@jy2�$�+�Ib�'�n�*̇�<����P�R9!%� q�'q��siW�R��´��Fd����'�i��xg\��4�<@�rl�
�'HQ�Rf}�>L�3BǨJ<��	�'{ȕ`7�W]< �;Cl�����B�'A�	��S1[p�i!F+0B���
�'� Თ�ə	�:��5Kڲqp�]b
�' ��A�(�.l�<m2��:o�0̘�'��`��GP	����B����)�'°HA��E����B�P�|p�y
�'�b�(t�b&]q���C����C(D�ph���jz T�V��pe���2D��q��T�Z��)Β��uaw�1D������v�ز��ˊXkĉ��.D��"�%D�wE���0kɊE�¥�!�'D��sfl�6�Z$��n�c����Ո!D�x��(U�!�2q��͵6�b9Z�#D�t��,ǨSY0�C'�L�P��5D�ș������][�᜴|�!
��3D����_\愚g�*}�*��*O���$�wX����F�.m�rA��"O�'ڱWy8��䯓<tf$�"OP�[��A0r����M^((CA"O|�:�%�4/:y�g��*A����"OZy꣪�2���J7@w@u�"O�x�© ��ic�ݴ>5\0�P"On` 쑺l�Ȅ��eގ,{�)��"O�YbW��g�2K"E�9P�"OX�ɠ���?�p#��Z�iA��"O\L�E���7������ݙa�, ��"O�Y�bEچ)a�)
5/� � �ZT"OD�Qt�Y.m��x�c��?HK��Ѷ"Ox��W��KKp,�Ȅ#8;6M�"O�a���2�64J�E��xB�"OH� �c��5�Ҹ5PĤ<9�"O��	''N�E����	����6"O��p�3��!c�枠E����G"O�uf �F�{���w���"O�,8�37�ڵcg�"rx%3�"O�����Ь��o�4-gP1�"Od4x��L�t��hC)�E��!w"O1rnZ?}y.��0���+�"OЀ��F�zCέ������A�g"O.�Q3��%L���ʒ%�NEҵ"O.��K����M.��pa7"O�h0'×8x�kgiE?���8b"O�����Ɏ/H�� �Ֆ$��S"Of�5cI�p�(T�v�؜^��"Omx����scH�q mA6W��H"O^��@'D-lX,�!�ɡ:\NU�6"O��"��;�}5*ӃA+����"OV�
Ԣѹ���1'!
N�"O��`��#��eۇO@� h�`"O� d����Q:W�ޭx�M[�:P`��"O����1�n�P֬�>r1zB�"O��s���یq؇	3{"~���"Ot�{�J�%��A��zB��"OZ9�&k/u��hZ��J�;� ���'���'���'���'�b�'�B�'�:�+�$&�Q���[1@�����'/��'���'ib�'��'B�'!�`���FH�,@��GJ#w��7C2�'�R�'�B�'�b�'H2�'I�.ٶBc� �"0Z�5$퓇���'7�'���'y��'��'�"G[�g��}y�O�}4�ZJO�I���'���'�b�'���'B��'�bϋ:0+� ZA��+�d�穎����'Y��'���'"�'�B�'���B�*��h��^'
J��j�!6�'B��'��'���'!��'@2O��c-f�RK�5��H+v�(�R�'�2�'�B�'PB�'���'���Y��@IY����F�,:�R�'�"�'1��'0r�'_��'��C�@! ٓU팦n\�0�싗8_��'�r�'���';2�'J��'U�٥K��
�c�'_Q��ka�7\?��'��'���'���'g��'5L�Mx|���
z4`�	T�r�r�'s��'�R�'b��'�'��&��ȴi'Ζ�M�ZG��
�B�'��'���'���'��6��O^���FM4\jb���';"�� +�=�T�'?W�b>�7����-���Hf�
t��P�G�x� Y��O��mZY��|��?q��޴.Ԯ� �2?�(��g�8�?A�����4���h>M2�����M)��c-�9[eH �$�5{y�c���uy��ӠD�������x�������*�4ZE���<����f��.�.�j��CE>Ό�i猈[�����O~�Y}��t�3sy��6O�CdF�}t�Đq�ޜn�X��?O��	��?�&�%��|�Lp�Y���ކ@�Y�4��3i��p����3����E���"�6���ċZ)0���.���pl�?�RS���I���͓��\5h&�[�N��ĉ��+R���p�e#�!4Vc>q�u�'W����xo��b���s��Xf(�/r|�|�'r���"~Γ��H+3��" ܊�A�I�	/�*��/�����dH��}�?�'RpЬ��#=Jq.��秊� ��Γ�?���?�s�^��M��O��,�J��&$^"�s�`�% W Q�� ��PܒO(��|z��?Q���?���7�DZ��W���փ�RiN��+O(9o-�2Y��mޟ��	�?�6
�ԟ��I�~�!�� .���Β� llB�Ox��(�i>�����Õ�@̾�ۡ��x6����Q�_����iy�n>Dz%�	�G��'�	�n��Y�T%��x)�lC�b�
i�t�IƟ�����4�i>Ŕ'��6��ttx�D����ѥI�Bk׿0�C�c�Of�m�R��+q��ޟ`�Iԟ����;V�¹iY�����ކ"�`�[b�����'� �e�?u
g��d�w��P1���"uR�@�P�Z.n�쁙'���'=B�'�R�'J����hVy=���o
9&�Ɛ�B��Od���O� oھL�J�'s����|2 �p6��S�c a ����&U�w�'�����D'�3i�&�� � \�7�|@�cI";E =����Hl�r��'1� &�������'�r�'�ֽ�Ȓ��z<-Sz�h��$)�?����dئ9��c���l�I�d�O�0��n�/�0"r,R<m(���O<y�'-��'�ɧ�I�':�Pmp��/�$t��	=A>fx2�C �6q�����@>�%�D�w�:���.T.`�Z �B?n.���Iߟ������)�sy�`x��Ńs%]5n,�,C�X	��!J���ų�^��Sݴ��'�X��?Մ�6RA@q�u�E��B��$	����3wD�Ѧ�u����+���
iy�h
\�,l8�(K>s]�$��i��y2Z�p�	�,�	�0��ڟ`�OG��9c��5a�q��'WI�hԇl�B��V�q@��D�O�ʧ�?����?ͻ'�&QS1k���ǧ��n:�{��?�I>ͧ�?���=ZP�ܴ�yR͂	nW�p9Ao99�x��d.�yb���T������4�<�z�4���	�hNs'��<$�$�O�4�?�.O�pn��E#Ҹ����4��9��ِ�ؙ8 e���>q��?1�W�����$�l{�F		�4����\44�}
��7?)�CK���9�Ā[�'������?a2��e(�
"�d�����?����?a��?�����O���nG�v��K�E:Y�ĄJ%�O tn4|��'	�7- �i�5Y���'�r ku�F�@<���w@z���	ҟ���7��)l\~r#�g��	�5P��(�%}��s��	���h��|�\��S�x�I����ʟ\J���,n`!���oP^���vy"�y�x)��O����O���󄔷07>���
T�)^N�9��Fd��a�'@r��I*Q��b�n�hR��9A��ɯbGެh)O�a��Ĉ��?Q��,�D�<Y��H���m���[��Y�+S��?I��?���?�'����8��ß�HwMƔpX<�-��Z0�U4�T�������?�^�(�	[y�l�L�@髒��/YNRQ��FH�a!4�i���!��e�O��D%?-�=� n�#�T+�m�E�<*�T�I�;OB���O.���O����O �?��h�`H��Q�B�f�T�qu��Iܟ���4rL��*O��o�K�	%S>u���F��IT�Ӿ-�@c���	ȟ��IGh�lZ�<���6J�|
�>D�|9i��GuN "��,W�P�d������Op���O8��X� q�����5��!�a�I�Q�����>ʓ:%����8���'�RT>��� �Zk0l��k��WN�$� Mc����^y��'R�|�OT�`@�R�T�B��;��� ��tE�(E�./�8�O���L��?�q�!�$_;���i'�]8O2Rm��c_�B���d�O����O���	�<V�i����e)R?ht�(�4"�., G�۪X��I%�Mی�>���>�z� V/R3R(�c�e��n�d���?%�?�M��O�nY3X*��)����$��$�V4��jF,g��4�� Jn�$�<���?���?9��?)*���KC�|��{��Ϝ|Ш(�n�>�<x�	ޟ`�	\�Sޟ������5��
C��<PV�C����:�?1���S�'7[j]��4�y"BQ?�h1���U�ΥUW��ϓ�v-ON�D<�Į<��?a�+�n|(gɔ9�p��MH��?I��?a���d�Φ���˟���⟴�wC�aVplP�"�;G�d���j����I�����z��	l�P�mހ~�q0�@�(� ���0���X�|: +�OLS��ݠɛf���4K��
�c	D�Jh����?a���?i����yŸm���?1�iۜ%�d��d������"ݯ�?�3�ig�u��Q��I\�I՟�]?mn�Z&#҃ZG��
���p��	�������x�a@���̓�?���:=����=�ZX�l�N��l�O��"/��'�x�����'b�'�"�'~����#H�B�i�5�/yd�+�S��P޴	)4����?�����)�Ob�$�36�8�� @ȶk��Œ���9N��?����|����?)%(�'[�dԨC[��R��]8f���0�Gy~�F_�p������rt�'��ɪv�.	�$L�r����Z�w�>��	ş0��� �i>q�'��7�ǛGP�M�7Y��ӷD4
i�-;������������?�R^��	ǟ��I�N$�*`LD�o~�8Z���f�0 ш_����'_��z���I�O#G�S.&��&��;�d�$��.�y��'|��'b�'�2�i�?4�,�J�(	�ʹ(�M�<q�\��O@������qUkp>I�	�M�N>�r[iM(6��5%����!����?���|se ��M3�O�\��A/uX�١�/,rqѳk�Cs����'��'��I���	���I�t�M:S�9)E|�Q�T�U��������'�j6�^3)θ�d�O��D�|�7j�v�PG�*+b
4�Ip~"g�>	��?H>�O�VL�#v44:u��S��M�Gb���Q�醊S���|:���O�5�H>Q#��{�|���"{*$[�._&�?����?���?�|2.O2d�Ӆf< �xW!�4p���+Z�!h�1`҃�<��i��O���'�2�WV���@$-�}td]�qگ`�B�'�F<	�i��iݹAdl�?u��\�����`�P�Y�~�Nؠ�$s���'�B�'���'G��'��Y�������P*̰�� �s>9��4�������?�����O^�7=�`�q�ÞC�| �支v*X��R
�O��b>i"�Eަ��F��c�5{�^9i c�b>p Γ��Q�7N�ÖhL>�/O�d�O
L8ckΏ �$$j��M�v�1���O��d�O �$�<�2�iO"`�@�'���'��ݱk޵P�r[��n���b��{}�'d�O�H���&�������V^�1[�����%f�N�@pb��L�S�O���ޟ�)�Dߒ'1�p�g�^�]M@��_֟��	ޟ��Iȟ\E���'��Q)��t����f����>A�w�'��7m�t֊���O�mo�b�Ӽ{��(+\��CUŁ&s.���D��<���?q��=! u��4���g2(q��b�^�#�I�P���af�\�B�5�Ĥ<�'�?���?����?yV���9" ����2/�P��	U'�����Yá��H�	ޟl'?M�	u�\�ЇS�E!��F�/ ���O(�$�O"�O1��@ #�� pY��P̄'�(��T{o.7-1?� gGU\��Iu��ky�F(L����%��alЁ� �8 Q���?���?i��|B,O�oZ�]��	
ZS��R�ݲ@�DU�V(��f^d�1�M{�"J�>���?a��)2,"���ln.!�]sK�T  �ܱ�M�O�-aQ��"��T�w�Dl�F�:x�ki�0u�����6��O�$�Or��O*�?���8 �𰦊S4G�`U�ܟL�I̟��42�ș�'�?��i��'J���!�>;2��dD�&&Q	��|�'F�Ol�e
�ia�iݕ�1+{���m�� Z`l�Ap�V��ɓ/��'��I� ��џ��Io:��2(Љ	8tHS'95~�������'ތ6Mˠ6r��d�O���|��'s�~i "I� nPhR֍�K~�Ƥ>Q���?!O>�OS�ё��Y�J� x����0J��*&�9�k�i'��|*G��(%�(��I�|�\�KG�Բ)Q'%�ԟl��㟠��ݟb>M�'pd6�M6
�P����WOU40��bn�O��d�����?y�_���+:��%��]G� �	�O�,�Ҹ������̦��'ʸ�y���w�*O� n4:s�3q�$5�` �qq09�5O���?Q���?a��?������m@L���ǃ�J���F܆f�ld���'�Ҕ�t�'�:6=�R�	&/�.).-��,D�cr,���$�O���2��IH06�7�s���U�-Ҥ��W��-��
h��q'�@�b��`�I_y2�'���+�Vl1�|�6D��r�'<��'l�I��M���������O�]a�	��z �ᡲi�H�8����'�D��?a����qu�1��a^-���T
��_��A�'%���C��.g�����~"�'��p�)X��z���-�^
��'�b�'���'��>�	'&��M�CA.s>���A.�@�	��MC%�����Ҧ��?�;Y�bd��"٧v���Sv�\�&�z�Γ�?i��?�Cd��MK�O���U/�?�ڑm��GG" qD�SI���6)ܾ(7$�O���|Z���?)���?I�_�03q�L�S� �3�m��p)������I&�Qyy��'��O�R�C�N��k�ʁatH��B�ߟQ2��?����Ş@t���%�H�l��-۵��+��,�>hR���,Oh�ⰄE��?9;�D�<�)؜L�H��pȔ�3���Q�E3�?����?��?ͧ��$Cͦ�s����s�D��T��P��nMa�H�����ٴ��'�r��?��Ӽk�MMZ~"51@Ύ~�bh���&9:�޴��ē�W�2uk��M�Ғ����Y�����O�s�a� [$���O��$�O��$�O��$%���":(&�X�H�+�v��8g�'��'�r7��W���Ob\na�>� D�6�Kk�l��D,qX�Q$���	ğ�Ӑc��<m�Y~Zw� �����7<�l�ue�('2n5�q�Q�^]b#�d�	Dy2�'���'3���:�:Q���H�nΰa5G�C�'=�I�M�u���?���?�+�&�IvKAmaY#�8u�5b���)�O��d�O�O�Ӷ ��P�ag��^䰹1��ˈ{�eRK�~P��!?ͧ������a� ���,̷�4���Z�$,��?���?)��|�7���?+O�!�S^��Ĉ�mF��@�}ƪ8���O�d�O"���<ͧ���O>����
(����!Rvb���O,��� D �6Mp�|��;�" ��' R��hnn@�"֯	�� �OP�T�I��?����?A#�F;�?a���?���?��->0��Fmǆ�n8K��8*�����$5�h��Y<�?��Q�������Q5F��D�&pΙQ�Z�r�뤂9e����OD�_1Հ�4�����O�	��Lh�l�I0thGH#7�����+K̺�Ɂv�� z�'1��&�����'�(��v�܍omT��Akް'G0U��'>��'�rV�@޴jWj�����?���W�b���q�\����F\
�;���>���?�K>A�K��D�$]�C�U����M~B�;B��PQk!�O��@��#r��%Q�$��� �:98�uXs!B@~��'$��'2��S֟h	�
��.!��LJ;�H���՟,@�4 �Lq���?�q�i	�O�n�7��P��F/P�h�d�dq��O.���O(��"�x�t�/L�׃��Ȩ�af_?"��d��nETa�N������4���D�O���O��d��Z���#�������"vhUh�C�<qf�i����'�B�'���y�#r���8VnR�s��t(��ꓢ?i������Ap��Ш��&��`kf/�3i�����e��ɽh��1r��'��1&�<�'S�蘕N�D�F B� �T@c��'���'����Z���ߴ#Ԏ4��>W��̇'c��lKr���M��ϛ��Jr}��'�b�'���P��P4�L���� `�x iF&8���d����<,*��i��9�onĉA�(��P�\HI�>O�$�O���O��$�O��?�Kp&��6����q珑{TV�'$���,�����޴���/O��l_�I:*����*0��g�0$���'��	���� vQ�oi~Zw�����د\{��rA�e�`��d���~]�M��Nyr�'1��'(�#P���xw�̖T�6hQUY�p��'L��7�MK���?i��?	/��Ӧ�2�t{��ܝ2��x9�O\���Op�O�t�j��n��+��X��@7nAl���mK~�O������W��y�)��WѾ��`@T2?����?���?��S�'��R�9�'N]�kqH�-D��*�@k9��*O�8lP�����T ��R��B6	�}��my��Iݟ�I�?0�l�J~��$6��Y�Sc�)\�W���	p�Ol~�X6 WH�D�<���?!���?����?�/����@�
w�\!`1��h���ÏƦ)��������ҟ<'?����Mϻ4�DI�G�:X��0SI�:�,qK���?�M>�|�����Mc�'A(���C������U%{)� B�'�>�:��
J?K>�-O���O�y5G��(�D�@&O4�YbF�O��O����<�E�i`&���'���'�� s6�G頥��`ǩI��ͺ���s}2�'I�OF�k�nԞOM�����@�ˀ��g��`9Ѩ�p��@���z�q��ϔ�$�VEG/q�:PI�Ce�$8�+�����ߟ���ȟ�G���'u$�ck�e$h4`�f�=3a�����'��7+<-���O"lc�Ӽ��]��Ժ�cb_j��<A����D�bL,6-;?9&f����)]B�? d�H��W�Q ���r���c�0 e/���<����?����?)���?�"�_���M�bā�h�$�� ܫ��$�ڦ%�q�����I͟P%?����p�F �`B�"� g�^�W�T99�O����O~�O1��<�4[?Eâ�u@Z'>t�xZW��
�P7mBFy��Ӫr�f@�����$
J�a�HP�FrP�)��	Y��D�O����O��4�&�U����,U�,�	A����"9���8W%9S�"��L⟘ʯO���<�w�	t4����~
Ҝ���I�8@nu�ܴ���B�=)�C�'m9 ����� O�L R	�X�Ti�%�Z.-����O����O$�$�O���3�S�FlˑL��I��HYg�T��'��xӆ��1�?���4��D�T�[�ֈv�,A�e�P�Z��ThL>����?ͧrh���4��d�7}����	z�f���*V݆P˓JC/�?��I6�ģ<�'�?Y���?15I���(0��C�)�䣂�?�����$�Ħ�Xp�I̟0�IH�O,���2��	 ��/f|�+�O6�'����?�S�,E�c�9EN��W�F�h��L?U�R@��mX?P�8���������p�|�+B����l�r���$��1���'���'���tZ���4�~��w,�]�"YS�O����D΍�?�������H��`���؟��P���YP*��AB�V���n�ȟ��I�R]m�h~rn��J�t��}���[(o�5{��-oЅ9����<�.O��D�O��Oj���O��'�0�*�S�u+��౉�(P�ޔ���i] (���':��'
�O8B�z���(U�
���	�.X���*�2?G����O��O1���(��a�.�%;x1ֆ@8L2$aU<I'���cY�9��'V�'�������'*
h
5�H�H`��P>�<*��'�2�'��Q�B۴A�Y����?��$����"mH�2<X�ԏL�wotT��(�>����?�L>���� ))f��ε�D�N�t~2N�k4�b�i1�zT3�'�r��LPM`�F�%1�X��G߁~Cr�'M�'[�sޡ٠f��=8�I�.4��x���Bٟ[ٴ~;8����?aбi��O���لi�0kG�l�����g���D�O����O�H�-}��Ӻ#����M<<��d��̻U��h�ǁ�J�O��?����?���?a��=�J<@����-8@��*G)�1b6nʓ0����J�'d�$�'UV�Ra�+X"$��i@=?ʡ*��>��?�K>�|zVJ	��D���aT��	���ܚ`.D�۴t�I5��,3!ܟ�$�4�i>�ȖJ;*fP�bk=~�fI�WLğ��Iӟ�P��ٟ�3a��uyz��bk��q{���+<�`Ra�^>�9�c��2�C5�(�4�̩oZџl��蟸�	�J���
QcB�����ı� ,dͦ-��?I�  R��i����d��f����\�^�"�2Y�I)�7S����O���O����Oj�d)���wv9kEaW;{�<����7*�0d����	�M���N�|j��D�V�|���O�dm��L���\���R�'������A�~����l���ӑ>�� [�.`����bROQH1��'2P�&� �����',2�'D�e�(�� m� ��M�*�dA:�'��U�4�ܴ<zX����?������H�,�k� w֠IjQ��&��	����O���'A��#�N.c0̽�e�?v�����W1�p�cܯ��4�F���s�,�Op��rț0�`��C�"/�����O����O����O1���A����G�C�ZI�S� A�c�
kL�0��'�B�`�b�@�O���Q�
��)�rc&z�$B0�ĬV"Z���O:�R�fd���Ӻp㝕�0��<��`�W�����	�bw�#+��<Q-O��D�O��$�O����Odʧ]+0�	E�Ⱥ>��܀��	�lZh`�%�	ޟ���o�s��������ˣ^��i�d蓹F��H���'�?����S�'=�t5��4�yR��&�n�B�2e|=r@�%�y�F%Q89�I!��'>�i>��	#��y��DY�yp3�߮mn
a������Ο��'��6�l�|�D�O*�d\�q ����-�xak�ds{��ܲ�O����O|�O>D �@O���Ί����FMi~¦D�!����:W�OU�=���:"��!$�p�N�/!؉�w��:���'���'�����\{CQ����%��RE����hٴW�<%�)Of�m�f�Ӽk��
�&T�5X�BUt�P��'��<i���?a�s��-��4��ĝ�)�����'.��	�H� u���1�OK�!j2����;�$�<ͧ�?��?����?�b�w���x#e�J)(MiV�#��ߦ@��U	u��t�������kkX���ǟ,�B,ލ��H&��1@%��0�MFyb�'�"�|�O�r�'��fһ(� D�e*��<j������8�&��O���A�?y�2�ĸ<iOG,�BX���d
Q���?9���?���?ͧ���\Φ�(�I�2Ѭ��o��i%��r��,�B�z����4��'Ͼ듡?Y��?��%�\qb#���U��݁1��-d���4��D�k����'R�H��&���t�z	z'�\�<����D��r���O��$�O����O��6���
���0E����]�*���Q���˟\�	 �M+�Lް�?a�!5���|b�_%?�(ȸG�/�Zp���L���'��'��@���8O|��ȿQ~� 0E�W��Sʘ u����p'Ҕ�?�1�%�D�<i��?9���?�w *<S�͉4�Z h7B�{���?�Ԧ��'Uh6��_�l��O����|��U;"�$[pE�v��-A"�I~�&�>A��?aJ>�O���%�yZ�i���3#x|�uJ=^(���%����4�B\��?]��O`��k�?C����7'Q�c�QÅ �O��D�OT���O1�*�E��6�=A�0��0C��9*B��R&E�H�l��'12�t��⟜�O6��Z51?V��cAʇgq� ���|k��$�O�m�2~���Ӻ[a�H����<1d �IW*�`�0_�+�����ey��'E��'�"�'�T>AWɖx�̸���u��CM�MSGCԃ�?	���?yJ~Γq}��w��5� A��3�%�ő�'̸, c�'p�|��t��/I�;O�qj�I�|�≪��V�FHf��7O�DH�n�(�?9�D&���<�'�?�+)7�>lZ��6���ͅ��?i��?�������q�G�M�D���A���uD�x�	�[��(SQ�1c����@��`�I U��Z���c�� !��٣f��3Ǌq%+Ƕ�\JN~���O\�x]TD��� �(��ކK2 �����?����?���h����I�-.��9��G�x�F}�'ʡ-t���Ӧ�C���L�	��Mӎ�wm�HمMB�4�F��"D�j�ٚ'�b�'"���꛶���1ke���J�P0 �/4�"��S�̓O��|���?����?���f�1�Q9��Ż&(�q\�hS*O��n��&���ҟ���^��	�����Z�r�n:f��,b�4��_����0'�b>�Q�7�X��E��-/�����$�o_~B�_�Nrj|��䓻�D��*�1�/Z� ]\33�Jd�.���O�$�O �4��ʓ9��ʕ;CX�M�����τt���ӫ��yB(jӬ㟀��O���O���P�9�ep2J�7�ƥ�  -(���x�m���� ���䟈�>���<�hx�"��]<]R�:2�{�|�	�������I����U�ǸFz�X��ۏF���'M=�?q��?�u�i@���O���g�n�Od�#�&���@�u���0&��O�4��� ��{����x�R V6#xlX���+��d�J��h��p�Gy2�'��'7r�E�)avXx�kC&�2�i���/���'���0�M#����$�O�˧��1��[M��MpsmQ�,z�)�'��드?i���S��Ɩf12���-}U�u���wnly`��A�tQ�9P�O���?!��*�D�S��  $EJ�dJ���;��d�O���O���I�<A��i�y��S5'�V�[B�[�/DJ�iC�4G;��'��7�)�	���$�O�����/���uC��%�b��O>��$�7�-?�ċĠ8v��>��Mŋ�
�IdFaD�Y�`�3�y�[��Iӟ\������	���O��
aЕK8�a
�.ր��@c�}��cI�O����O����ئ睶}��<j�K�xJEy��a������'�b>��5����y͓,e��8KH�c�dBŇ�&Le�}ϓb�$����O<i�L>�.O��O(iҶMUj@BqB�1��,�q��On���O,��<it�i��2!�')�'��9����(Qf�*A䙉n��l�q�|��'����?�����j+h����ߟ�@�� *ƤK�bx�'�	��l1��p����Bӟ�pP�'<~��h�2MB4!z��8h`Mu�'���'���'+�>��ɼ�l|�����o�6��K2��ɘ�M��a������Ŧ��?�;[��r�M^O�k#OL�5��P��?A���?!4�@��M�O�ȓ�6�
4kq�dYP�"�$e�g �<�O.��|���?a��?A��/�����u�A'S<g;�q�+Oxdmڐ��1�Iݟ��	C�s��c�ܟz���$q��@���A���$�Od��2���4� 9#�F��d�¹� ���zz\aA��3���y������'|�$��'O��������� eIB�� �'r��'���4S����4x;�@X��h;>�@vKۃA��Ś� 
5m�V����P������m}2�'Z�w�&� � ��⌶o�Z�*�#�S����k�@G����U���9cWH��a'L���#�/E���!.}�|����@��̟h����B���:��Aj��_�B?`Yڲ!K��?���?�5�i�4Q �Os���~�O ��4
��<�Ƚ��GU�-yV���1�D�O��4��Y�@�n�^�@`n����Le��Q�K��D��y��س^���j�	oy�O�"�'�(�(U��+t�͌]v��`�X���'�	��M���*�?���?(��8#���4q��ԏ3*A*`���ӨO��D�Ox�O��:�(��6hW|��	�bA"d�ܽ���R$>��ioK~�O��D����D�VP!C��7*��Hd	<8�����Y�V�R�3ִ�
�J��`$0w��_���03�'��fӆ�`��OZ��*��\Y��[i#��v��c���$�O.�+Á}���$W�[�Ǻ?��'��q��PY �a���b�r��'N��V���3�jOJ�	
��ɤ=��R���2�M��L2����O��?c���k���@|�����O���%ȁ�?����Şa��Mxߴ�y
� F}AJ^�XD�b ��~R�A"�?O��[Gd��?�'E6���<�-O�� *�,�J�o��v:a��'7��,4��˓�yr���/`0���պk:�DH�
Y���'�V��?��������[�-�{��а+CZbU�'����K��+"0�*P���
^���*��'��퀡[/aT1�n��)�a��'��9�Cm$~W�3Vm\�Y:]���'�6��KǠ��O�o�{�Ӽ�g���-%f��+_-�
��׬�<����?!�-L� �4���@�"!�1��O2*0�ŗ'���������"*��|�P�dE�������]%=_qI�G��d𦝚�Qy��'�I;FjZ�-� &@��N��aCu}2�'�R�|��
]>t�TAb�a޻U����M���sC�&nV剞*6����'��}$���'��T�S#4:�X@Vҥm�5�񉼤M�##�?I�FY�z�f�y��Kr%*e���?��ik�O���'�R�'�RK��8�� (U�J�)2�$�i����Ȅ�Rҟ������S5��Iq��P�$@����%,0�.�O�%*�k�-)@49��#<���X B�O���OV�n�3\F�'?@���|����X`�tC�w�&=
���~��'�����T�X�k��擟,�����D|�P��)��	�䴐�J�<}��B��O~�O^��?Q��?A��)9mhȎ%��	ȺPp���?a)Oj�l�P�4���ʟ(��B��,֌H�P\���Q2�3�瓱��dIL}��'/�'����XR��y���.��y�U�d^�%�X�%�.q���'�������K��|��B�;F��p�ZA%0 �(؆	�'���'���TV���ٴ]��$�� ���aۯ3���;�f �?�<���CD}r�'��T�`�ތ��u�#�Z�^�"P�U��z��Ǧ��''�8 �?��՜?Ѹ`�8d�,;��E�~��\0O�˓�?���?����?����i��7�b}���Ay�d2�Ķ>���lZ�/��4��֟���u�S֟�����1��==���Æ\1@..�S��<�?�����Ş	@`��4�y�ݠ�8W�2,��Y:f�O��y"!�sk"!������4�����E��AiE� �6}9�EQY����O���Od˓^*�f��w��'���'J,��C�&sCR�N�90E�O�'l��'K�'8�<���?����v�N٤O|8�-��x��6�(�Ӄ}��$�O�esv��:-�Ԃ���V�&�����Oh���O����O��}��t���҂���U�* $a^�1��͆*J 2�'�t7,�i�m�7�8�,i��N�r�NT1Gr�\���4���E�nv~¨��Z���,�t����lyJ�$�/>=�J>�*O�i�O��O��d�O��r��è>.l�7�N�dT(I�<iq�i-"xR��'�"�'�O�R�_�
�209��$@d��d�>����?����Şh}�|x!B�8�饬��)���j󋉧�Mr[�HQ��_H��?�$�<��Rb� 4�Y��N|��n�!�?���?A���?ͧ��D��ݱE�ǟ�1j�9h��xqa%�ms(Aٟ��޴���?Q]�P��֟���,;�*�k#$TYE"�+cX0��nɦ��'��a�"�O�J~���:���Ғ꟣P���@Y��ϓ�?i���?����?�����O�H08�`�M�pXƅ��69�$h��'r�'e�7-XD��O��l�Y�I6ҕ25�$Z����LPY�l'���I��S"T\�oZF~ZwX��i�m��#/�@���B�l#�2cꖙ'�R�OF�	Xy��'"�'BR�\�m�L�����Ye`�I��T�b�'>��*�M���6�?���?�,�.)�7G�&u_H���M�Y ��8O��$o}��'���|ʟ����
�� ܓ5�G9� ء��΁"~�H�2n�=\����|j�Od��I>��X�@�RAЫ�i�����l��?���?���?�|�/O�oZ	O��l��"�k��tI��S0N����ן��	��MN>	��(��Iǟ�M����ة�b�(�T�x�Ëɟ��ɞ%�Vl�^~R��06b(��'��$؆k<�\Z�fK�؀���oF+7��<	��?���?I��?	+��qi�	9>���`�ɑ�;���ܦ�µ��џ<�	��,'?�I��M�;we u!��z��*q��,Jp�q��?�O>�|�Bł��M��'�ZX����j�p#�%L�	�'�����N	��W-߭��� R�B�9��A1P��<~�ڍ
�h�4Ȫ|�������@�̊)��C-ɀ͔AKj§6� � �>=��q'O(S���:�(�*f>Z��ǤF��ڲ��<KX8��&�&H��T0&
�<�Z�Q�,��ÁY*n���y!�pM� V�W E�� ���<H6[��/+&tra�K�cir�PB�kDx�P��O<!
V��աXĸ�S֔���F�W�Q�ĉ�G��Z�/��t�ѕЬ�����(G�{�j��!�
j��	�2)Q���@k�)�"2.���c~Ӧ���O8%��D� �N}���f)���^6m�O�O8�D�O��������Ex��c
�Q����ʙ�x���'I"Z�<�Ab�����O<���VM�Ff�*\��,���'v�*��NW�I̟��	)g��IL�I]���lZPac�� ���#��Ц%�'?��%I�.���OX���ק5�@Ò^�Q���ȷMr~ �M���MS���?9��U�'�q�� �CB��I�����hԓ&�8���ix�l��z�>�$�O���,Y�'L�I.E
�C➹�l5�#`����Bش\v�����O��0J��`���!�~���b`��e��ߟ`�� ~u��ʬO�ʓ�?��'�����A�j8�\*��LmvT��}b,]�'�R�'Y�G�D=ԝI&ǐ31�( p�#.�7��Od�5��E}�R����W�i�J�`����a���i L����>�P�����?q���?A+O�)�3��\��BFm�������ݵZ��'���۟8&�d��۟�adAZ�]��D���_�N6�3�	Z&�&��	ڟ��	Dyr��&�n��"x�JН�B؀�nW(>�6͠<�����?��[X��h�'�N�u��k�z�c0`G$Z$�i;�O��d�O��d�<yt�������U(Q�pg�Y�V/��1�� ��M����?	�N��{R�UH25".ׂ)��� O��M����?Q(O�`W�Uj���'���OdT)�u ]��;��,�GY`�'�2�'��$S��?�P@Ɵ	S���T#<H�\�$i��ʓbp-�5�ih�'�R�O~�����"`�z�+���ə��
�M��?A3&�1��'�q��1�v!���ʅ�Rf�2�d+�i,��8w�u�����O����^��'+�I��t �J�;�D�CU��~��ش4˨�`���i�OH6)�l���$)�Q�#o�M���?��J8顴Q��'r�O�I8�+�K�5e�A��	*��'����|b�'�r�'fx5�f'߼K��	y)B��X��� g���ć�N�H$��ߟ�%��]�/3V���)&�Ȁ���X�ZOz���<����?�����d��a#���͆D��`�a\Pq#G���ē�?���������<q��T:�\������z�i2X����ʟ���`y҈�Y���S�q�$�)�C�!O����AC�Xo���?q���䓝�4�����QR�� C��v�E��E�-X�'���'	�Z�x)���ħf20�8�ѽ���!C%�2$��	z��ig|�T��ҟ���L��эE�+��AdO�~�z\��ig��'���1S�m�N|�����1�Y���ěU.������c���%��'���'��yZw��2��+|Y�9�%�Tr���4�����qV�i��'�?a�'�	�Q�}�&l��.1��& �6�<	���?)ї����4@��J9f:Ja�3mDЩmړi�:|�I̟��	����Gyʟ��!cF?[t|����R#J{�Be��V}��
�O>�gF��L��MR�b̊V���b!���Ms���?a� n�k(O�SZ�$�!�� ���4o� 
�N=	T�<Gx�n5�Sݟt�"��+��[�x��$M+�l���X�0N]oy��~��2�X
��U���*I�u8��h9�Ol���O��?��L�=-�	� �;!ܦ(�B�J;-�.��+O���O6�d��F?��"�bE����	_��X����yc�C7�ǟ��'�BNf)�)A�1��!K���7����,� %����'�����O\ʓZ[�m��$ !��:���C׶hN:��?I��?y*O�X���g��(����s�_���ç�Q̌���4�?YH>!/O�)�O��O��(��Fs���jS�նNg̕8�4�?�+O���ݲI}˧�?�������(����r���� 倾/��}'�l��Ay����O�.�W�:����#�B�ҷ-�(��Z���G�U�M�_?��	�?e��O����uJ�0G@�}��Ǵi �I��T�	7�ħ���eX!ᄻ|6�u�D��,����VNfӴ-؅��O��D�O��D���S�4��6�d���' 9&--����)��C�6�Fx��I�, B�0XGA�^1��1v�ǅ�eo͟ ��ӟ�ڡ��byʟ��'~À��Y���S';M�x�/h𱟸�䳟����A�Pg��CA;rή��Vcq�p��9~jʓ���k��_�TzE-�Hܺ�@D�Ro�{w�x��^7����O����OH˓;#|���CL;�<�cd�nT"�!`ٍ8#�'�B�'r�'��i�%�EZ
�)@�M�% �<�Z�N�����<1���?�����O�d
�ϧWVA���J6c R)r�N��}�LL�'T��'I�'U�i>)�	 �69AS��10R�ZS�H;t��O���O��D�<q�a�;7h��؟<A�M�V��˦i'/4�@TF���M�������O6�$�Ox�	=Ot��-�����DoD�y��ti�>���O��#3�	J3V?����8�S$0��y1H(u
����)E��	`�O@���OJ���1���OXʓ��d��p\@h(bDĕ
�x3��9�MK*O���dE�)�IПl���?M3�O��@�H�n+��,�h�ڴ���՛�'D��]��y��'��V�'ff�=h$ӊW��]E��;AfR�o��lt��A�4�?i��?���J+��Ayr�9oT��b(ߖl�|��A�X�7�M�_B�d;��-��Ο�Q�K��r�n|��U�Z�R�SG�'�Mk���?a�X��T"S\�|�'�r�O�)*��FL��$��V=f<�D�i�BR���#�i��?������ �P��, Z�>3�$Vr�\��i��(��b� ����O˓�?��b�48� �N��<�0��UG��%�'��'���ȟ��l�:��a���<5X����*�F��`���ġ<������OV�$�O<�KF�F�
Y��ˀ�F�Uf	! ��<����?�����۠MW@�'�p�(�E��:��Q!HiZMo�Ly��'	�̟L��柠�%�f��X�.S3d�e� �<>�������6��$�O����O��tbf���W?I�	3ˊ���Ȋ�m��(3m�.N� ݴ�?	-O2�$�O��D����Of�
�0�̜0�l�#�F�ydߎf�n!nZџ���Hybj�e�H�'�?����s�6팝�B�I=\�q"b�!%��Iԟ���ӟL�	k�L�IMy�ԟ��m��; �²OőQ�X�#��i剎�e��%��(���?]��O��Ǩ?.+�O�\w�4����6B�Hm�ߟ��I� ��I��9O��>��*M"7d���Z�^�ˢ��f뛶��7��7��O����O��)Jt}�U�HJ�-@�.�f�sEN Do8]�u��1�M�����<������8������"kD0.�e�9S2����#�Mk���?9��A�y��[�d�'DR�O��ZE)C;��M��*̒V��(���i��I���a�j���?����?QE)��:��q7�8,Z5Y�ċ;SěF�'���H��>q-O��d�<y���s+����QBk��(�TS�V}".*�y"T�`�	�����Py�`�������LQ�4�(��!���a����D�>�.O��D�<����?���z���l�f�h�cs�	�KU��N�<!��?���?I����d��B�&��'n>�A���7�M��d܈\leo�Ey��'��ş��	����bn�@`E� Iu�J��D;;&YB�Ç���D�O��$�O�ʓA�(PW?M�� Ie� ���S �މ)㧍=�"��ߴ�?�,O����O����y��d�|n��Z3v�dh��M$h_(3w�7��Ob��<1�i�m�������?��e����m��?/��	�Mƥ��D�O����Oj�#�	eB#^���SFGAe���g+�O�˓�}@ �i���'�2�O�f�Ӻ{чUEg�xj�j�1a
rp
���Ϧ���ٟ$�fa�,'� �}��	�
�d@
+�|YC)�%�C��M;���?����X��' H�H
(�j9(q��ެx�W/pӂH��7O����<����'�D([�AO�2|����_-z̘RS�{�b���Or�e��Kw}�W�$��S?��/ ���D<>5�8CpO��I��@yC�yʟ2���O���9>��;T�r�	aW�(Qr�Ql����@�U���D�<����d�Okl�.<c� O�m3hS�B�.1�6�'��!˙'c�''��'�"V�ذ�/�(X��N���J�ht�3$��YʩO�ʓ�?),O����OX�d�"�r%�e�b7
b#FL(Tx��#9O2ʓ�?I���?�(O�hkQ��|�Bˆ�x�8���5��I��M�)O�D�<����?a��V��`��[cI>DMD���X��tl�������Iџ��Iş��'T�H�B�~���T�t�'��v#L�y2�x��с��i��_���Iğx�IU^
b� �!^[�A G�"�tIT�j�Z�d�O��z-�p�'T?���ȟ��� 9�%�q�4!�VE+��Ҥt��`�O���O$���2���ty�ҟ�5�L�w�,|���gql`h��i��	.3tt��۴W:����@������
�*7b}��*,Ue�<�GQ1�F�'�f^0�r�|���ۋUW��F�
�q�+	*Z�f��!8`�6m�O���O��	Y�I퟼�"�
=?< �k�ᐶF�TC��<�M�@*D�?�N>�/��˓�?�G�n�̅K�C��ns��Z��¸ �F�'���'�fU�>��OD���p�ƃ��lV�C�3v/�!Fo�z�O���$��O��D�OkLO+  2��S��*R| 1 ��t�F�'Pz���**�$�Ob��7�������U+U�]i'dB�WЀ�� U��X�G����'&��'��Z�����l<� EK�V4�┪19���}��'��'���'�.4��G.n�3�a�[
I�R%�>�bP�x��ݟ���Ay2��$,���ӋL&L��4삘N���:5N�+�O4�D>�D�O6�L�$�	b��1NJ6Ww��)3��e�B0�'W��'oR�h��N!�ħz��%��:y�ĉ��(�~�h4���i�2�|B�'��b��y���>9�J&*u�0	��9$�U�%A֦��	ޟ��'?8���K3�I�O���H&s�*�!�FΕ8����F�$<N�i%�(��ʟ�§y��%��'G�ޕ{Ԍe��E�F!�z�o�{y2�B�4}�6�]}���'��T�,?Y�g�;l}�ik��Ɇwj� �P���	�I��H����ڟ'�4�}��,�1<a�m��� /���4e�����M���?9���ⷙx"�'^�!xghܚ��ҍ�D�%�R�|�0��^���|r�i�Ob7�^�{-�p+f�#`��S%h�	�Ms���?Q��]����V�x��'���O��U�]�d\��2 �:(��f���;[�1O��$�O2�DW)	���!=S��v�&P0�o�ן`��@
<��'��|Zc��h���O*7����M8jT�®Oz����O�˓�?q���'9�ΘHphۿ<�1J���"Д  ��x��O��<���O��$4&+��{��+��p�F�/K�(��'�O�ʓ�?���?	*O�8W���|� .H����Px�Ċ�� �6��@�x��'P�'"��'�,@b�O��BS�( �بR�2p�	"dX���	����Iay�bϔ�,���"4,<�]ん�	��r��Ŧ�E{�W�$��z�$р{��0q�'I�b`�p��
*�V�'��S���H��ħ�?�����L0vf�����	�*�X�*J���D�O4���=�v�QGd��@0���f��b7-�O��$��F�h���O����OR�ɤ<��r^�x:�f�.b�R]`f�H1���n�ݟ��'��ub���t(�n��0늲7D� m��M�K(�6�'���'����>�.�u�`�"i����I:s���E�ɦm��Y�'p�'�"`Qk�H���M]0��y��0[.26-�O��D�O~�8w��O��d�|���~�k��na��5�Mnm@� ���
xFx#<������'e��'w�Ձ�,R"ަȢ�Jٟ�
�Y�C`Ӛ��_�Jp�$�Ov�O���|�,�,MM2p����,�B}��]24�'��B�O��d�Ot�$�<)��K
�*��;s��W+W����Q���I����	ߟ��?��aș(�	5"�JlM#FK�:����|��'62�'�R�'�,�(uן(�r��V8J�Q�ȝ�i��Y��i���'2�|��'
�	�k�6-��d���$�͖v<%+QT�|����8�	]y��'d�%��^>��I0Jr -�%S�dC��:��>c֌p�4�?iN>����	pȉ'&,D;�n*GYrH���*��)p޴�?�������.9r�&>����?;%k[V�D9+�	�.} �{�� ����?��a|0�#A�+4̌����0��mZfy2��F�7-�_�d�';��;?y�j�)ZӺ}��.�	�A;S�ڦ��	����#�>���OÞ=gmJ�xbШۏ_��Tz�45�:)Zu�i���'�"�OS(O(�dƸO�� �2��$MtM:󄉫6�F5n�7$��#<����'7 ��fJ�=S�5Y ��	<F| ��m�����O����w�������O���g��p���C�2�10oZ"E���$�[����	�@;-��|i�tAѸ�4�X��M�i��,ZaR��:�����O��'h��%K��R9�@�GD,H0Z|PJ<�N>����?�Ħ���ǟ�Ҁ�� ��ݑw ̪���'I/�I�'<��'"�|��'	��΍X�"�hP�  Z�u#�#G�w~��䋻��"�(�?���<9#&ʟ:�*��V�_��y�"O�,����?Tx�[7� 7]���`��ԮBHJ �gP� <��0�� ����%�c.%����Q�<��(��_D���wg�.|a�q�eI�p���Z�I.8cT��e�칡D.��c<80�`�4H	��f��1<,�yf��~�,��g"l��Lc�#^�i}nhKgj�$UH�P��)u�H�cɩK��0�EE7U����G�������5Ș�2s�K*��'L�jD6#i0ٶ$�G�8n�|2(��� w��V���/
LPT!t�>����Z��AJ- ���P�S4��`8t��;.\�!PN��s��'[�\	��?9��i�OX�����`�4*�c̵z|���"O���k�3׎����-b��'��#=A�f�
b��]	�*ѳ!(X��FY��V�'�2�'(���(Z����'#��yg�G�M������V&��6E��?Ȳ���I5��d�6U:
0�r�|��F�{���g�$���3��71���Iܤz����'Ih`p��L>���
Z���h]6B�F���E�?1�O��8���t�,tg(@"�G�0 ~�����M1NC�	1
n�Q���c80���10 �vő��Sßx�'�-�`B45#�M	�C� 0>~�R���=��P3�'��'��`r݉��ß�ͧF���s�O]�!��D�Vm-L�DJH�0��9+�k�\��x�	ϓ�|��'�U �hZ�E�qs���bH0f�ta���"Z�"ϓe��"��=�ڐ�	�Q��p�a�D���	T�'V�O �����5=4`H.�/�d�@"O�qX��!����B�U�N����������yy��S.T)��'�?)d8��YpFGH)2��y���A��?�o�t�����?��O�2����Z���MW����!db	�J0����3K)�ݻ�9O��S
�	^��%8e)Kp?�0O�8<p$��@�떏Qj8��ؑ��O��<I���a�\���nPt1�j	�H�1O\���P�@9|�b񫎁z�-ȵ�"�!�$����!�]�O�Z$���T�cb:as������'�Yɧ�e����OB�'$�N���G�:!�&�Q4����A.�G������?�����/�Ir�Oԕs��i���ɱ|e���X��Mr-����}�$� ��[,�B��e���S�^���"R�A�xڊ����@8��'����Q����7ҧ�*r(�c��ً'��r&B��h��x�#Әl�|$���-c���l��0<)��,m8*	 �^nP­`b'6�,ͪ�O���d_>$�4�#�U4���ďPb�!�� ��Q$�>-����!hC�1)�"Ou��K������OI�Y�Ez�"O<�c�̷%��ɲ �Ψ\K$Z�"Ohx@��zC��Qd���B�"O M�r�0�zp����0[�Ʃ�#"Ona	/F�7,�{�`�Ff A ""O��� �Nv��W@���C"O��س�H���:o��B�d9ʢ"O�LP��ϵD��cD�����s"O���M���`g�4;:�u[�"Oz�����>Y>Ua���q���"O�l����:WFp�r�2�&�a�"O&c(PK"���T�#�,�2�"O4(;��JvɃE�܏l���a�"O����&u�,���&�*��幅"O�`j�I8.04�A �)��iS"O���r�	a���Q�H	�sv���"O�*B�ܺtA�5�P�À_!P"Ox� �-�Z�BFCȝ`�b�k0"O�݋���_#�P�UKߦS�����"O���@�����ũ������"O�<�P��K�@�TfY�s��A"O�L2��A�U��yಃH�C���"O,%�U�J��8�q�֠A�*$�'"On� 5&˿}�)�P$U�h���V"OD�e΃{�����ȫoW ��e"OdAY���1)S�V�&D�zd"O*����+u(d�Me1V���"O���VdV<c��̫�	�F��9�"O�!��;8ZRՉN�-�f@R�"O�e�� ^��B�.β��I�"O*�'O�B! Dr,Z�S�6x�b"O�pX���l����&k��H��k�"O��j��P=�zUؔF�Q����"O��q�W��5i���4�4{B"Of%����+��鰉�0k�ܵ��"O(**5E	x��UI�i���+"O�\�N^�U~�y�6(�'SBR���"O@���gԌ]��s��#&�"��C"Oܕ�A��n�(X�I"i�B���'f�e3�Kaʽ�C��>{>��\�o��� Kn@8s��&ZA��Ac!�wѾ�F}2��7�>�!���2S��Y� (2�ԧ3D��˃*�9;����MʞF��p&n������Vu�S�O�����Ѝwr ���M1����'3�-1B�V,+�z��F���@�O��P�k؞�#�m�U�,D���/;�6�+9�O�
��iӊ���O�=O��Ÿ��˯2	�(�"O�MC\e|~D�a�1�ܛ���K�'� M�C铫b2��G�N<Ll���\9n�rC�I�.�l� �Ȓw�T���C��:�>�LN��Gx��逭\aL4K�-�'(�M*�Fy�!�$Q�.��AI
�B���!�.Sp!�$҃;�\ͨ�ʐ!? �*3喰KB!��,d�� q��U��u2S�kX!�A�*� q�o�7r�T(u��n�!��@�c+�tA)J�bW�(8pO��!�$W�^0�4�@O<`qՎ$�!�D8QJ�[���(2��b��+p!�DO+.�� \�&���1`��g
!�߈uS����0Ts��W	�!���Qt~��i��lkWs�j���'�V�j¦J�$�⩑��A�c�v���'�"��	�$*o��R�D�H:����� H��~�4kE����"O��륨�\�P���Cݜ��*��'���KM�����آ�����"Ĵn����(D�j�T@qL4�PD	�m�t/:�	�	�dI�y�����)ͷ(	
l�j�j���V��4K�!�$�>{ϠH��t�bf�6jr��s�v�r�r�G��N|��ѵl�j��}u\.A�ұ�t  D��r�ϴTc0!1CY;lH��b�,�.-��MI�n��)��m	����b`z��%EG������
��@�Mm?q0�L3\���O�q�4#RC.�]2f+77�p��'�*82a�'��y���+8�L	1n[(ǜ�ʘ'T�y��Oza{b�G��O�j`yf\?I��Z}ۀy1 J^�3�*�`��?D�X��g%�M7!�*	������(q:R��5��+%���LB8yK����HJ(�x�HI�&ިj3>�C�%��:��}��'�� ��X�+����FP�u��n�	hΤ�1 �p�F�@�BA�mg&̒��-�I�io6"=� -��@���ۥ�Y�Ժ�"MU̓]T��&��a�@Y;r��� ���'�l��V;xU���G�-t�~5�ȓ<�H�Y�$��θhT�Hc���ܭU��{7㔻&�5ϓ��O��5�w�p�Q��A�6��p�дq���c�'Mb�Jb"�?4,|[��T�Ė�B۴|	�������븐�֍��:��ʓ�<ړv�b���	�+�̅��ԬY��I��!�+3g��Z��#"�/��웠�R;��
��C)b�!��ߞI�.����B�j�@V$N�g��9q6��=�qO�9��ܮ$�NQ��B�:=H�ę�Yo��"�>�8��=��!��C�,��B�I�"SpmqRꖻpf]!��B0U��(4	�&Ge��k�%R,Qٴ�(����;Q�p遆f@/j��0⣆�����}���ZԊ@��4�l�?r
���'��g@�+  �1�%�,x'��XІ8ғ_L<[$�� )ʦ� 7�-	�DI��4��)�6�47t��#�#oC��9eV�wt�����_����m��s�f�x3H׬�p>i����$�B,��
XY���ly��c�4Q*dm.+3�jv Q�И���Ô$z�q���/�1H��E��y�H	�h�	��"o��I[�lM�\��@�0���<�O^.ؑ��ɺN9�n�1���A��(aZHu s��J&aR�Ըu�LFB���hz��9Zr��BP�<1��I,fh�ۂQ�S������D�'e��16�ؽq�����f�(%� �����0#w��HFjF����z�LZ�<���g��9ER�)�)�,�`�� F0���W,U�B�|���� ��6F�8Cr�s����d�1,�� .�t��dj	�X���	� c�(�B�#��K�r �f�:Gn!��H�z!7D��~Ԧ�@D.�8-��0��02��Y�C�>%?M���L�1�`�]�d��WŜ=z�>=b��Z�B�I�$st�����
�Q�C�Ơ~��Z�X5��ɫ4` y�hX�o��e��T���\�'�ԭ�a$
?r�.a@^. Ҡ�
�c���1�!zpr �M�#j��b3�ح&ܒ�� �<���Pq$�v��h�%Y���>y�I���<z���r�蓰OU~�d{m>��#i�jo �IE��?�W�R;=���LLe��#�]��܋v�܈��C�* �[�+v�|H���M�>���>r1bS��OȄj`��p��ȅhd��QS�!��lcd@��E?B�����'2�PQ�) *R�	zCH�g�P=���NqF�be���wdxr� �<��o��D{"�'$C�\�n� X�K��0<�$(	�e�|rw�
`ނ�ǘ�U�� ��IJ�f!Pe.��-���Z!� Y�Ն�����`���ۖp��	���S'@|d�'aBP$	� ��P2HM<,��t��iC-@F�	&MI�.fp'�U=n�!�D���P}���V��i�Κ�|AdI���,Pj�'V�	�𙟰� ��
V>(5��9s3rx�E�6D��s"�1H��u�c1g�X��T�Tg�Z���J�&q"�' �ˀdE$uf�hT���v�	ӓz3P5��ӥ%�����M�,���`B�N�v��J�����Н��<�&��&KB�0�������	�<���Q���bR*2$�|"�$�9��]�ա�2z��hH��f�<Y����*�e)�^(���V�B��QJD�4L���O��,���	 y,��y"͞25��s1%	,Mh�B�	+ �>upCr՘�!� Ieވ "3�C'g�8�#S��>"��uS�8,O�\��N!+�:�j���h�hz&�'�i脢*dj��P�������LtA�%d]B.L�@�!��$�nhz�
O� �@x�k�=A4�M��&�9�F����>���]{�:�(#�1Ho|L�#�VѦ�>٫ӎ�"�F����F�8��f) D�D@���&2@Z �?���D$$L^m��(�E� �m��?�>�������f���;b�xèE�w��)�	m�(��q�q����a�d����] t�`����~"�ǽm�I�� �?aa	Ր�(O�5đ)2����c$�+-��6�'&��I����`.���cʸC�DbhK
��-�uDL� 5������/a�7M��E1���������a�)]���S�I�6nO�y)�س�l����	��l��'�>���8����E��q[Dm:B9��j�̼Yc+U�Y\^�ŉ���r�"�ݹq>B������|*�۟���u"W j�ܜAb֬����˃P��(c��w��ز��$$� ��Ӷa�>b R1
DF� 戩*O��
A 91$�'��'r�l����b�p��g\+Mڒ�XS��R���c�!=�I+Osꑒ��>IBj]	6JX�ׇ��4�����ϭ^!���+�-lmnJdm_�k����J�^:B݀V旣�0=���Z�l�҄ˎ�`�R�y��H=���)O�H��$f�佰ROU?4��S��S6���T�N%"�D)���P9>C�	�*Ġ �b�$@�>y3��n�:P)$J(t�6i ��C�wc��֧���?qAЉZj���B�J�*��9�J��R,$���'���R �����@�1s�,b�B�@�뎜%����wp0��:��-�\w�0�8g�Ddb�xz@W-I���2C�$���Ï2�IMKġ��2�S�d��Ǉ��w�t�ؔW5G��X��8!rn����IpTq ����S��'LO��9Q���_�i��<^�a�ܝ�Xb��A�ͿSUH��ɸ6p@��g�u���W$jB�c���0��u��ჵq!��P��]3���:G�0�PsO�R���@�G�B>�q`S+uwԱ*A�-����	�?^�>��uML~M��
�e�9��`��I�e��Y�d�<�� �CI �3peIS��"5J;m�r�2��G� �0�#T��Os]��D	b��Q�EW0NΠY�4�T�/Y�O8�p�JQd��L$��M;I����k�RV�H��Κj%^%`���1�Z���׆d����i�b�C'��:.��ؔD�?� ��G�i:\G�E ����|�q���K�!��_�~��#�"�zK ɲ4��$P�^h��cHb�)ڧ!�:}sN�(>���C��[\����O� b��U�K~�CA�v��&���!��mB ��I0v�nk��)p�ver�H�Z/6��dC6Ynu�ȟ�z:�{��T�.�u�EMS�P���uÆ,)��4aj�q*$�۳5�x��0S�O6h�&ɋ�{��lyuD�6�@��"Oց�Ł��:���+��ΔA��u��"O��Hq�֛���B(�\��ؤ"O�]@@�@H����<Tw�L�T"O,`Q�"ȅD�pE���!6�rh�U"OV�[V����MV��Y�v"O�EEC8M!f�@)K��Ȳs"O�q2���:��55 Zm�H�"O�LJ�m�=}TT��3��xB"O�XIC��#W�ޝ�PnW
x�F� t"O� ���"abt�lS�'���ڷ"O�IPǃ��z�4��-V�1��ʗ"O�0�m
$'����t�V���(�"O݀�eێD���0k�����"Od�`.�?8��4�=dm�;"ON�ЮՁB(x�#L�)qE�c�"O&HxAI�d����(Ӎq�*�1�"O蔈�Wl"&`�H� U�.��G"O��j"�G���Y7��h���[7"O��R5oĩ*���MӉ*�ơp�"O�p��	�op^�P���
��ձ�"OR z��	�k�2�4�̸M���P3"O�"�[�1�f	l<N��4#�"O���/-r�)���B%pP� �"O�TfN :��.��tX�T�"Ot �G_�h�0P@5��X^ܨ�7"OFL*Umm0ii�I]�}(����"O���.ab��vb_�`"�[g"O� @ՠ��C<�6\r�gP�%B\)�"O�H��"l޽sa��jͣ "O"�Q��:��J�%��f� R-7D�8� L�,�Z�ʀ�Բ>�)@��2D�l�%c h@d�z�萁0g2D����-J��hوf��6B��PJ2D�|3��)����☛rn�t��0D�Hn�� ����̘�
�J,J#�$D���OR����ee��[]9W�$D��9�d�N@N���#[ ln�-c��$D��E�G1u�i;-��dL D���A!DP�*č[�Hq��aU D��@���+NX��U�Yum�h�s�8D�l��Ls+�qJ���&v�^`2U� D�p��8}a��QKR�z����?D�x��"�#�՘oΘ{�A�Ԯ<D�L['H�"WF��V&�9;N�y�1�0D�����Z�Z���PŊ�%6��A�C1D��х�������ʊN�R��N3D��5��C���z�쉾Z�B��'3D�����Û���C��@̐�.1D��#ŨW�s��t{E�GF��&�)D�H蓢B�\�h)���4΄q�-&D���VC�;'������h�vX�'�����K%�"ؙ��@�U���'�a����#�d����8N1�
�'֜!�ٓL�(�P�
9N��'^�J����T<`���9���'�@���p�.e�w��@g��@�'Eּr�@�g�R� 뜛29&qK�'!��R ş%\���xK	%P0Q�'��S�-=��*b�ק,�R�y
�'�ZpɆ��|�4:�HG�{5B��	�'b���V'��Ȝ�:��M}�s�'��Eq��|����i�{@�'�^�*�QS f�X��Q4q�Ƞ�
�'�����9
���zc��c<8|@	�'\Y'�H�e�&Q��&QE	�'�<�'	٘)��q�Aא4C�)��'�x5�@c��xF����L�$%.@�H
�'�<8#�ˈ-nc��r�l+=8�
�'�����Ί!Q��;cKOK>��	�'}5Jw�O(k��<Qr.Ԧ{�
�	��x"��� �ҡZ��8�̭�"B��yr�˙�`��!�^�<N8�Q7G�&�yҥcM:�jЅ� hmq��Q��y��	�T��A�/O��𩒢ڪ�yr#�,C��QVI��B�D���>�ybC�p�3�e)x�FB�,�y�N�5V �cb��I&�(&��y�R�/�t�`+�i�ݸ`(��y� ��*er�ɔ�_,��+=�y"��35���ò�G=[\S$ǚ7�y�C�|�b���N�$��h�*Ԟ�y� �s!�l9$F�g&yst�]&�y"CX�	��)�Ӈz��, kY��y"&i��t ��X�jw�(��(֜�y2i>ą�{�Tce`ԑ]6���'�hCn�#�����cޕT*J��	�'r:9Zr/
p����Z9�^��
�'��p*�ɚ��yi��V��y�'&���OL�jT��2�o�@$��'qX����M�T3b�ԝ�f��'����&O2F�a�遠j�
���� ��`a��Z$H�0N� 1���Q"O�}��!�f]v�q�MD8*��@"O4�1�V�oj����1a�p�c"O�����=0�� ic)�#�"O��x�O�3��@gj=
��c"Ov�CtgK&&l(����<O_X�"O\�a��?P�T��׌�ll4�bQ"O@L�0�ݥF2��d���SS�t""O�$���ހ�N30{F4	��̼�yR�"��݃G�1$�� �,H��HO��=�OR�p����.�¤i���l�����'_�\&K�uդ��3d���h�'��<�qE�y���"�K�`<H�'�����٨]�d�=03l�8	�'~ؙ'��/�|�C���-���!�'�&ȃ�,ޮaq(� ��.1�8��'�,x��$�0$��0���٩(d��'�B�:��J5/�����G��ys�'��|"6&�$ODB	3@A��h�r�'"pQ�c��O�D��b ��Bm:
�'9�u��HI���k��,:@q�'����O]�L��{�nT0J��Y	�'/���FD�-�A�)3>����![�����'{����E%2`��ȓ99`�q��]�4��,���!EG�}��+F�B�(�, ���q&�Hs� �ȓ1�jm"vd@=T�,* 
,Q�`���K�"�.ǬC�V�$�����"O0y9t�V�pI�yr'��!Z��R"O��w.I2U
�*���^���"O�@*���q��)E���H ��"O��@'&U���q�P�j�f���"O"�B�aM!d��D�i�l�F"O��q�g��Y��C��w� y��"O��YDMH�py���M�����"O�ۤD4��h�周u����"O��!'��9���!m�` 
�"O��Hkɽ �y�f�5uQKr"O����Bm�T� E�3w\	��"O� ��
X;�MȓD�b$���"Ox��#mO3y��p�E�BgG�8�"O�P�"	�4!�tl2��[3I�497"Obl��H_06��q��=͢���"OV�1OP	p��x�VD�4W�4`$"O4�1���4�� 	�;MU�1�d"Or��-͊�t��"2I����@"O"�S�gк�J�y w��XQF"O���GX�y��%��Z!n�I���`�O�^�06
 2H_��k�O1S��<�'��q	0��,vw~H�a�ހ�4��'c��M��-��0����	)x�1���'�!#�GP�z�]�Z�4���B�<� �A�U�Z-↥�3n��w Ju�<�Ε/=���p�$K�|�hUno�<��n��m�����!":҈����v�'Uў�'N> Yեݞ5d��ѴI�V�Є��c��=PJE�!�q��ɸy��5��G�L���Ɣ�I?�1�R%ò�(���[Cn�*�����U��
L/�rĄ�Ub��+q�O=S{؉���]��(�ȓ ~ W�:9)`��a�N�1=@��ȓ"?t�y�I�I908L�86@\�ȓ��yX���I�i� e۔"���j���8anF�,��ۣ̎����S�? THԧ��o4ȡP�$��B�"OB� ףY"cR��[����
��Z�"O�ѻ��
1�>D@&"ϞH�J��b"Oj%�A <Kb���_	vh�=�"O�Ir6�	�IX6���e�\]�"OlQ����<r��@�Зf����"O
�3B�X
E�f�S�2�v�"OZ��@��}g��r�T�+�60�%"O2�x1
Q�^(��р@����V"Oz�Ɗ�x��,J�'�QqU"O��Y�U�U �q�D��./lT�b"Ox��N��p�5c��$��B�"OH�*�@̦p=�ܛ C����(�"O^���͇\�����ǎ4#���!�"Oƙr�#�8�<���T�d����"O�`z���|��12U��7w�u�v"O��x!
��\��D:#SQ"O*liׯI
gFL���țk�&Xi�"O୲CF;1����"��.�
���"Oh��é��Y
t`)��1gtAPs"O�� �7��rV��j�W"Ob�8`��1���B ��kK����"OrT�]"+�� �T�i�~tiF"OrqPe�H�#�^X���w�а+�"O�g��0����+���� P"O6i2q@��5�9H@U�$���)'"O�!��*��,�g�H����b�"O��I�O��^�|����T-{��=B�"O�D�Ƨ�'z��-��6V�\k�"O4��A.
��-��%7b���"OQ1an �8�`
�+1J��"OH��AgĖk6���w�aN��q�"OD�#̄N�4;0j0L��Q&"O��D�%h4��r1h��1��"O��*�a��[q��3��	!+X;�"O�D�fO�jUh��U�, y�$"O줪 ň8����cZ�:�`)�R"O����C'`�h�#�%
����`"O,�1�N�5x�0�!��۾K����"Op�s'(^U�3�
ͬ4�
�;�"O�-�7(�"7u(�& N����"O�᱕��!H>Y
A��3W�U�"O��y�.<�n�LS�h�� yG"O����M8 ��Z2˒�8X��"O4 ��H4E5 Y�@��-C����"O��q&�-|=Za{v/",�x�"O�̱��.K�ŁQ�1 a��"OZ��EM��(� ,�B���W"O�H��fΝM*�"� -b��X2"O����"�%(����p��E"Ov����ۂ�3���\�#2"O �dD@.l���AFm�@`�f"O�`q��	[7~���@��6��Ы"O``J��I�va�Q�M;*�j�ä"O����ٯ^+��j�gB7/Č��"O�9#���
�^�)q�$DЀMs"O(� �!ϒI���r���z� -�"O�1�@�7 +�m�di���y3"O�}T�Mа��RHF�h8C�"O�x�5��)�����b���"OH��oE�w1�a�ǈ�z�Ԝ��"OL����T�i�N�b2��31|��QE"O��q�i�!�����݉#�0�@W"O�4 ���;@QH�G��j��p�"O� �m+uZ��M����oef��"Ol��!��<5Qb�␄�"j[Ÿ�"O Y@㈀I����DM�!P��"O�9Hr���c�'I�N8��a"O��f �H�ܵ+R` #(ȭ�F"O�4Y��s�2��#AI	"���f"O�Թ���=c���Y����"4,�"ON�[1�Z_zT�,�"2�q"�"O�-z0��A�}���:rP"O��6�٢���>�;�"O�� N[LLI�q�T	Ut��Q"O^5e�Nj�����M\�/*Le"c"O��A4m�+�~{�\ɀ"O�l�e�ڤF�8�yw�S&g�P�"O�H����	'��+��͈Q*���"O�m+ �L��r�Y�|�
t�s"O��$��4�"�	�/��=AVY��"O�!	���m-���
�H	L��"O"m�Wފ<:pq"Wi��EтW"O�rV�H��)�JTk��M8 "O^1��Y�v���L	�v��A"O��P��r�z��B:�b�Ru"OF\x�C��HZ*ܠ�)ѬF8D��"O6CI�y���*W(�,:i�p"OJ��	6<�p�a_;��A�"OZqku$�<#Pe��!� z7<Y�"O��Q�H�|��|1��Z�,��"O8A#��Dh�h��/�7\��$"Oj�2*��	ɺ�PƎߢS f��"ON�����T������Q�o���!"O*T3��a�1u/��$�Y�"O�Z�įUV��*D���0]�"O�M"u�5(�� 4��Uո�"O���3��#w��#�n��)�Xl�"O��'�QD�x@mI�8�,��s"O�ybF(�(�
`+ژOȨy��$%D��[�o\�d��ZF�W�[��E�Ќ8D�0@��' "ֈ��'�	Ŋ0� D����_�}�S�p*�
�?D�x;��PCE�M)�G# 3���;D��)4h�F��L;�$�%%���s,:D��!�K�A��i���Gh��p�4D��jB�W=Yds�ȩi��My�2D���E��P������qN�eC�/2D��� � "$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j���e�{�0ʅ/'D���#��`��`��Gx�q�1�#D�� �uѷgA:R�8%��lБ8��(@�"O��z���|N�!�e��24XR�"O��C�dǗd��F�Z�_b�a�"Ohp��L�PȰ� L�G�
�S$"OZ1�hE.?X����"���P�"O4��e-�8�0k�&(�N�KU"O�QIs��g��5��K�~�@��P"Oh�aЎ�{�|�˓�%,f�� "O\HJa�T���I��*A[��(B"O�9y�� /�l�|P��o���y2o��!u�;��ܨO 0�O��y�U�Fݖ���@��Ze�fS3�y2�G�{Z�eˌ.i�1�D��y�!��fp�h�3��2r�Z7���y�k!Oπ�
�E0V�\顶C��y�����i�/
#8����u�ǎ�y��;m��5K���z�����y�iR#|j���`��%z�� S�$�y���/q�0�+��,�ubҭT��y2�^��pk��"���5K^8�yb��;8px�4�O��43c׀�yB���"��G�8}�"�:"٠�y"M�"	1�1 �n��ph�G�2�yr H�H�xi���5��)����&�y�e�v
zD�� ���D���y�-2P�(јg�����A�6�y2�1N�Q+�(�v�T���'�y"��K��1��l��|�%���yr�G7��Y��H�]��C��,V��PJ3mHai��x5�N�d&�C�I&-��is�ѯ1��$����#��C��1p��ZDo\�S�X����֩3}�C�ɡ"��8aK^P�|��٢�zC�I"s�ԓ��U�ED�u����V_bC�I�8�|��`�Ǆ%z��,<`C�	�(���P�!K�T�jS�ˡ�PC�Ia���"â<j�x4g�7"x�C�Ɋ�`RD�^(`	�
թhٲC䉘*הȰ�-J3���h�'S�ke|C�ID��!��A�	c��p�,F7�@C�	�,�(l�,F���s�D�"C�6&��$L>/)fA�񇆬2�B�	�cƬ���.��3�Fd�"B䉝z���9�*�)*W���CD�%��C��+/ڼ@ҋP�q��;�FC�FnB��<#r�쉐�ز���Ia��}�TB�	'R�8pf�'~�A���g vC��/�����%.�#U�x�r�:D���bƜ"���[3��kS���7D�0AF�E8<��d"��<QڱzF-4D���'�R�M��;�`�Y�Ɓs�e.D�T���+s�R��P�65�i�f�&D�DٶA��5x��BckɷZ�d����"D��S%�yj,ݫ�
�4ْL"D� �)�}��-0�'���{� ?D���D��7�,XZeН:���3��2D�d;D���s���ƍ�8)��r��1D�<��),��{��N�Ovx"�0D�Tb�Nǰ|4�	����ewxx��/D�� �1-�QE�ަ^�(�3��;D�#熋S���;�-ЮyC� �i$D����Rvȹ�PmX�l��UF"T�D*3B�9n�2)#���;��1�&"O�)k����zG�j )�F�vkG"O� 6��Յ�,c���$գ3�=
�"O� rS�>?� ��7�2�\$��"OF����ܕ70��#�C!�%["O�����(
��9b��$VD|�a"O|�#s`@$F4TVB��r]�}�"O�<�� ��b6��cZ�D>F�P�"O��sHK	uz)q����[��0�"O�$�&mY-�>��Kͅb5�tH"O�ٓҦ�(ڂ��J�L�|%�s"O�,[AOߘXr�3	�
^���"Oj��d��;�X��Jey��"OF�z���7��8*����԰d�0"O�]9���g^�0�%_�#� �1"O��Q0"X�2%<Ј�M�=��D"O�z��NM	�܀'-JX�i�"Ol1���,�=��"4Oe��9�b���XF�PeB[�.�,�ȓ%��`6� .%c���?+��h��?9�T�K�c��`�f������ȓ �p�e؝3����`�7�%��L��Urg���Z9��*�6���k��cE��:p�������e*D��ɐ4]���tO<P=����-&D��thͬn�d�+]&+��sTG"ړ���*§ �����ԓ�=ے���_Ghh�ȓ�*��RB�;�n����;5L��Z-��Y�Ā����с��8��+I0ȹ`%}��$��86<�ȓv�\���?+����q�˄p����P�
��ƅA���!��S?!����M]0�%���Vg
8���K�y���ȓ5��9{�.ԏa��|Jc&�h���ȓȑX-@�%�d���C4{��ՇȓFPu�U+^�o��@h�-\R�!�ȓ�r`1�K��d�v�ѯڥQl��ȓ5=��@�F^�L��Pd�7h���K�� ��E�X͈��)�4o r܅�(�z�Y�4o���aB<;3xa�?��N"L�f���[\�tA�g�by�ȓF��a1!��V���[ E�T����u�f���NUij�At��$a�怇ȓO�TE���?W$�t�&C:�>�ȓ'��i׈J�R�b��x��T��۠��cʘm��$/X�,Y|��)O���d����m��
_�+�Ԁa`�ڼk)!�P�e+Bu�r-^�� �H0�>�!��M&b�bAڂ@�>X}��z�I�!/�!�D
�A1��s�eۇ�L���^-'�!��@�`�����j�;S���(����6R!�_�v͑ӅG����#xȆʓ)ciSf�^
�Ű��&lB�	D���h����vp��i��`0���0?ٗ�u��M��m�3�*�����o�<Y�Ȕ:U�&43CksJd���`�<قѤc����A>^�`I�r�<�%�H(���K�$ж���5#@m�< m5rZ6�PU�6��Dذ�q�<Y7�5o��[���K���aJo�<a��؈`ZPp�`0\��r���i�<qd�g�c�k�^}�h�o�[�<��W�sT�SB�\����	D!�Z�<��<��8���j$,=%d�Z�<��!P)DV+0�P|P�C���!��@%"p���%��	|.9eݶ!�� ���Ԋ.�<|��8gly*�"OPi��$T�[���O��~��_�����=p� �zC�N���s�f_8�"B�	AF\���Y<�(�%�-D��C�	�OO<	���՛F�F�rq�,�C�	!8e1!˓�D�I�˕�+n�B�I�.!�$bB�N�T�9w/�,e�|B�I��p5¦JY�Ax%���J:C:B��\X��#bL?t��	��=3Q�C��%H�zɒ�_$l�<xe#P	-վB�ɁUi�H@S���#V渠d,#[XB��<|�n�(��|G�hIs% 0FPB�>�΀��� ?�n��ïC`�C䉜C�����"���w�3nC�IG�	�F��R��T҅���K��B�I�E�R�V�}_DY2h4:�C��9?h�4�2�
(���H�nC��:e��i�J��&N�����R1�~B䉟,���QKF)I>�
��2�C�I	#u�kteV�K�Tu ��k�B��!G�5�r�Ĥ6�f��-��PA��� B��sd��%I.����C=_�!�N�s�&�.Y`��e�!T��O���dB1�ְr1Æ64ڴ ��V��!�d$Qbf�2��
s� �R"	˪%G!���7�j�/%(��0�&�o��q�'{�$ë�>E������Y�z�v`	�'��9X�c�*(@Iʤ��"ۮ���'�HH���J)(���S���|YxO>1�r�I>L�<	�Ǆ��zeX@%�iςB��V�D�pE���y�n���n�XB�	r-P��ب�V�U��C30B�I54�çX��2���W"�C��P9�ؒ	Ɂ7p��g�A&�C�	3v0�K����Z�8"c�Ӆ%��B��
|'fD���+~��7 ��+�B�38 ���ݺ�>��c&"��B�ɨ=��\�0��6 �2\���Ԟ
�B�I3iV�Q���8tt�
�ֺHB�I�GI6�3����"��;�DB�	�'�v��S�Ηq(�Ape�b86B�I�y�0�!�H�j��rL�wJ����h�x
䣞�M��=0�� w��败<�	X�'m�Ɉ)�����Y�Y��EI��C�	�^�&X0���^��X��aA��tC�	 ��QBg�t����b%�V��C�	<tvi�E�\�{��ؒ@e]
��C�I7�8��R�$fa���E���[�FC�&d��@u	�/uL)���8C��8����(��4�pB
�Q'C�IK��kvA��Gd�pR�����B�]u�M�� �7:-)���!�C�I>l����-�X�$\6q�C�I5E�R<9��%	�m:����c_�B�I1�8���/ƞ)-�!!�̋��B�|�|t���O��)H�	�Zl�B�ɖ<�n)�a��t�D���]��ʓ�hO>a�)��Bi�Hڄ����R�v���I�θ P�!W!��Ee�<K^���#�f4xV� +(j8�V�B�qֱ��/ ���_4]3H,cZH���t��ɑ���z�d�+d��>	�J=��h�J�[�˟�i;�*$K�fЅ�e����dվd�4�	g勗qc�E+��� "��7AP2|�.e��
�yB�z�U��G{��C�-[��I���:^�ΨU䁘q�!�Ē/��}Q��S�;��B�!O��!��ĉ!Fu�ҦO:_����dOX��!�䁀}��Ӡ/i��m�L��l�!�Z#ưH��U1T=2�3�j>?�!�dI8�`Iʡ��q'j���)DA�!���*.�Fƈ�9K&t ����u��'��O?�"f�!^��B��CK�*���E^U�<�v��PP�A�Rlހ�n��G�H�<�m�2R0��c��X�H.J��QF�A�<Y���F��Xr����}w�r����<QV�_7@`����%���i��}�<���߀G�Rа���af���z�<�R"X1kc���$�
s��9Q�+\�<G'#�^�;� Z�$ �����p�<��ObA�&S4}֬�j�<q����? �tCNƌy�@3�d����<	�W�&��d���Bz�h��[k�<���׵/D�=q�eJ�HƖ	x��D^�<e(�|��1�$�n�\��Y�<�v�X�H��Mi���	k����%�J�<��'��P����ՠ,wc\D[�a�<9��Td�����\���_�<��&
Q��a���M:�����[��8�I��،�c���xy��%��@����t��CQ^L	�u��0����ȓ_�9#L��:�@q�5ǂ��Z���<X�+@�F��PJ���ȓ#z�Y` ��s��ճCL8 �ȓN��-�ҩ�7�8 ź�G�z�<)q�X�6�*| `������)Ym�E���O����́*[Z9q��?�r�'�T��)J�=����>�0�'���HG2/���ρ5ogL����O0uy�jۖ$���hui��f�>�� �'���|\>c�擪lM�@�G^�|bOG%�6��k�P�Y��Ě@A�!"��j=�ȓb����,=Z֘����	->���ȓIz�1Z� D�Z4B�z�E�C.�u����=��苽UbH�V(�(h���ȓR� ���;+�8Hـ��gO�I�ȓ_�(�hU*�7�‐�E,!?�Gb�'w>	�f��!�EH4e��zhI�� !D� �7$�ř�EL�t�bI�* D�,y0�dD�U U��v�PQBe=4��!4oܩr�@A�g�g[Hx
��x��?!����ɢf�$9��[�n�'"Of(��UjX+��ւ$
�m{B"OԜif��E��tP�	!Q"O��7�	Vp�BbG�{�b`�"O�P+GFB(�vՃ�Il�~ ��"O��3B�T!S$}�#��l�֌�r"O>�ʧc�!��U1�
�F����"Oʉy'�:@�1� GՓr�l���"O�E0��V��r�eШ
�@qb�'w��xbOG�t:sB׳>P�����(D�x:C�2���C� ��%�,�E	%D���w����}�eӯi6J�P�=D�4S�E]s�pA 5j�>gB���E&D�����]�0�
��c�z�ڱRǥ<I��哾,P��#��	$�.��D\P~B�	�
�|�sB�^]40c#NJ�FodB�	I�,K���.9wLa �K� �C�)� ִ�QŔ�m�ĵ9A�ǡ!/�y("O�*�@�n6xKb'Q�}v|�u"O���J6O%`��.G��""O<�P@��
u� h�K���p��P�|��)Z�'GD�K�Γ��v��㬚7N��Ax�'�ґ��G4!���nY�K�J}��'nΑ��O�'ؔ����=�a�'��Y�B��ɖ�]>�3	�'�b�IĂ�l�,���2Z�E��'V��s�䍽_��Y�+Y�3�` ��'�z�*
��1j��~����'ebX�6��z߬�Bb	�~`�"Oʀ��7u����F��sϤ��P"OB��cE��jR�7�@q� "O�)�%k���F �Q��o΀�#�"O�����=
Vv��ǡT�Y��i"O��S�&L�r�B!BL���"O	�� ބ{�]�PAI�-%�!�"O6��4��F^��¡��(-��"O�iK��H>y�BJ�ϑ"$t�"O�X�잠jǆ�A�^�}{�"O4l�~a���8>ձ�oǎF!򄎍g�|:�˓I mRb 
3	;!�dD,12�Y�.E%&� X���U(5!�d%�m�K�6��5�7�̓	!�I�W�|�ݴA�R�Z��_�7R!�Q'Q�̡a��ZXP��u��/S:!��E�I,��R(�c~к��^�>�!��>\&I&�N�敱���j�!�D΄ea6y�I׾R��C��5�!�$O!L�9:0j�kM��`#[�y��y���%U~0Z���N�bp���2�B�I�A��`����SJ=QR >
3PB�I)xt�g�_X*� !�P�'�JB�ɜM��H��WUu��2�-H-/!�S�0���#����bQ-�t�!�d	�9�X����D��!�w�� fA!�d�>�Y��GH�d��IԌ	L,!�D�	x� �Ǒ)P�a����E��h�D�.r�<�w�];"�*l�pc2D��ZF�A�,:���"<�����2D���SB"���l�Ct���#�:D��(׀8g�B�p��V7F�V�
:D� q`⊩Q�zU����@%��6D�d�g�ņ1H�8�0
.249�cA"<O"<�C�֌C3~��֩�z��`#�GV�	o���O=lqaСՄ'a�@�@�]�"��	�'Ͱq*f�ʐ'b�si��]�� (�'jr ��萧~�"�C��]ݖu��'O������â�S�'�8�r�'O��z��)>��s�
�h�I�'dwm�����"�b�c�'�$)�GI_�}�� $`��bd��'�%��,���PS��8�8�'��q��+f�ЃglO=kL���O�Z �'¢�ZGG�0��4�@��uפ�r�'��bG������Lܑ`p�uc
�'����.��R�U���Z�\���'���;c�1=�8�k���YkRE
	�''ĭ�'��:p�p���1"���"O¹�� �����(�h��"O>a� (� usr11�08���1���8LO�܉�B�'q��׭O��j�"O��@D��w��Q����"�z�"O� "�S�I�mQ��	���RR�"O�����z���h��Ǚ&z��R"O�`k��ٿX��}�V-ϡʨ�0"O6l��#t�Q��m�8����"O�"��B�r���R18�����"O�-��	R6eZ�ʓ�ˆD.d�C"O��C,ܷ6,��c�ԴN>��#�"O�$k�M9Vtۦ*�\��"O��0Έ�r�;�� k��A�"O�9�tJ�g`�q�#�L����	}>��1��lt������>�Ќ��$9D�@[��ԆO!EŐ��A8?ɶF�j���ҝ!�:��չVL䁓�4D�\��Y$s����P�S'��q��%D�|ۢ���A���y��Ԍ(�r}{t�7D�� G(��2z�SӠ5'� �ӆ1D��`�b�,�FPq`D�m+DqS��0D��(�I�f���sl� %nF�3��"D���Ѧ�> 4ٺ��X3��%� �+��=�Ol(h��0��h��Q�	
��s7"O����^&�L��M�.�ة�w"O��ÃB�<I�IhUGȣB�*%��"O����!ȼ��,��.����"Of���"-yt����"Fj�_� ��ɂ`\}����}�Hy���D@��C�I�p���ؖ �B���f,�:H��C�	Z2���G+Kh�� R��A�Im�C�	#��b��=e����-�FC��&CR�"����6�@���	�d�NB�	Zh�0t��K�9�N�| RB�	�WKh4��̀��<|�%�ЁW:�B�I�b���aM �E����o����C�ɹU$~p��g�-;�}䚟"��C�ɋ5�a�b:"�5��Z�KO�C�	�H\���%U'P,HKZ�G)6B䉪AM�$�"n֥
��p��Y[�nB�	�J~�H�狚<�\z�B��fN&��'�I�@q�����M�@������z�C�	8<K4��&��(���^�W� C䉋<���%�{�B�1�NڍzOC�ɕGpL�
@�*C�\�JP�ׂ^�C�	�Js�u	t�D*
L�!3G��LݤC�	T�@�[������JʜS$�C�	J�H]sqk	�oz��v(G�Vr,C�G#.=����0 �R)��+�(c�&C�ɭr
̩�靂!e$��gC$�C�I.�`��0�82LO�Ae�B�ɛ(I:pDC?y;�M��LG.kw�B䉈w4v�Yա]�3MN�84��<��C�I�@���� �'J�6([ց�3
�xB�	3�Cԍ\'%����B�P�i�(��$+�ɜb�̸�g��F���P�͇sf���%�ɷ$2���ר_,���yKʉ�XB�Ih�0cw͑�y��u��ʮP;rC�I)5��� ̗�<H4Y����Y�HC�	�?��(�CKI�Vp�X��-aXtB�2��lV��n!� �g� �BB�I�MQ��x� Ěd�-ȡ���B�I;�t��r��*T�e@#��YBB�#Z#��� ��MMR0�VJWz7��ȓzB���A\6���IZ>��(�ȓF$��۱���h)e*������i��e d!�
mT�)��t$�y��{���y����K
��͛�Rժ��S�? lHˢD�,�� W&�}T"O�(�g��?**�ԁA��	�Z���"O�M�O��P.<a�$��@�P@��"O"��S�1t�hg.RU�q�"O&=1vHD3il���#�j��i��"O$(���E3�
0���/j�hH��"O��B#@�P�0�����b24j�"ObYqE "Z(t��T+&��("O�1p1�����TA�W(a�CW�HG{�򉄟e�~u+TmY�04���N7I!�E�D���E�P��2a.�}�!��>+��ٓ��E&p�T�A��^�N�!��(�6�0�@	ӘM:��֫(!�D�Ҙy�S��*ULT!��(N�!�E�r >�)n��d�D6�M(�!�D�<&����nɶL���b�"x��O����;��ʭB�� KaM��>�|D��}��K1�Ý<����gD�|�ȓ<2�`Cv�:��)F"�1r� t�ȓ��ihs��B#8��!%��e�p���d,B��3e�� "���)F����ȓ
}���$�A�HQ�U��LRS�>���zR���

�B�����Ćȓ|\� 0V˃�ĉ���'
z���	Y�? nY�+ҁ�:�y��E�I�ҕ�ȓlR(�Q"�2H�z$�"�ܝH��܄�qۺ�S B�2��5��N�:0��ȓYź�ce@��9� �G�D�wq ��ȓ.MkP��<"%��t�� F#���ȓ+��3�!�)<���B��K�����H~��K�5Ia�At�h)a�3�y��	���gG�e2"dȖO�����d2����
�lS4�b�H,Ò�C�"O����S8g��*�ቪsH�D��"O�T f�	}�^��5�G@�`"O$�i�C��t��d��9GA����"OJ�:U�D�>��z�,�H4�S	�'XD�`�E4;�҈Y�C�zQ�QQ	�'�$:&bБ~���s�H'm.��	�'��@�@V�P]9Uܨk�X��	�'Ȍ���Kâp��0�ԯ��Y:���'���S�D�_�: �� (�����'
��c�vr���Îٝ$(M��'c4h!F��]`bec���ND���'�,݂G�Y[~�M��F߾;�>H��'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\���)Ą@/����f[~b!��/8o\��w�x3�)��GE	#U�O���-�D!�3� 6�yG�A'cR�{��Z�cvYS�'��' ў�OW�I�$��=5��e��B�1����O~���
$���Y�`O�n!��F�IL>�S�͉�6YRP��5���3Q�+D���V�J'FpP�)P�s=�8��3D��0rC�W���S0���|@JgE2D�,�P��I�m�@���\��#�2D�pw��B���"�s�p²C�O�C�I0����dD�aZ���D��:;ɂC�ɚ*��bj�.��̲�X�s��?���ɆK#�P����:��u��A�	�!�C,UA�(�+��5Y�,R�@�"~m!��H�eծ���z+�;��!�DIT��陁#nyԐ ��8�ў4��S�'���
B@3���޻V��C�I8Ơ�$��>�fD T'�.f�xC䉚����1�ɭ{MX�����1}�<�=a�'p�`��ρ@�Z�x��	g���w�Z�C���J[��A��J�
�Ї�<��}���W�D�l�@�N@(<������6&pK� ����PB
��'��U�?����~Z�h�#&�V#1�*i�R�*�[�'aax�Ăx�j��B�NY������y�΀:����eͦ\�20Z���y�HUlp� ��]+S<nt�fnH��y��N�3x`�k]!}�����B��y2�ȫtM��"M�!0��S�2�y��*�"��4��Ƣl(�M��yb��.3�`�q��
^>d�mC+�y�
�HoVq�a�� ��IAU�՝�y��G.YiBQ�r'A'w�������y�j�&���8Ďִk��![W��2�y`�M9X�!�ߕd`�;we��yR�/dŋpm�Ms��Cq'	�yr�K^����c�(2��}Cv����?��'&�{u�0Z���ZBHݰ&�.Y)���'U�8E�E5*����ъJ0���@�'s����>�HH�T�
o ���'8���2�K�5�L�� RA^�k�'�bD`�� �ẶK��B<
���'�Z�x�G?�T�����2��!9�'=�hXg�³c~��6A�4U�\]J�'ޙZEo�6ir�� wg�z�2m��'v��[��2Q���qF#P1~�.}��'���1ׂ_�/	���l�y��b��;����� �S�803jϩ(z9��"O�樑,v��,ie(�9Ng��� "O��a@%��f����ć[d0i�"O>
nŨ	w�%�CH�-��U�V"O|��sEz*P�'�(��"OjI�6*J�o�${f�H�y��"O�=�b�@=�-+���-8�py�"OҰ*HȮ$t�C(F@���J�]� ����Ic�h'�[6~��d�a*�j��C䉝Q��I���G�&L�]���H�M��C䉬2 y�|i�i��Ѳ �C�I*2�ĥI��J.�Vb+�)e���?i���S�OHTj�.B�	*��`��A]�UR�'?f�g�,eD Q�E(1!(�'iĜ�҂F+���1W��.)�-�	�'76������sY�H7�
*�J�'d�9h�3�� &��1AIb�'^9�*�<��;��N$��9��'K�	V���1<,c�IXSZ�a+O�=E�� 46��E�E�L;=���kfV��G{��	�:$���aU�/�����)M�'�ў$�<i㫕/]b�`��I��Ȣ�C�<�W���\�*T��?Jǜ-q%(Ue�<Q&M��� +"��FϚQ�Q	�_�<�`��.	��U��5�b\���R�<-M��S&�¾oq�5;�ԜR��ʓ�?����S�O���AJ�)H��{�*�c��y�
�'����'�x��-zd
a��E��'�\R�],O-^P�#ϜiJ�#
�'Hdp!�hˉaJ6%#��G�.���'\r (F�ƨ.���P�D�����!�'!8pS�HA�Ex4�w��x����'6��A�NM�Xþ)�GҿoL���'_����-g��֦�� ���'Bx��u���2�"
��"�I[�O�H�[׭B1u�L`�%���[�"O�y�$���L�RT)S"���b�e"OR�rΘ;<��̐�o
(��p��"O�\*��K�>b ZNʈ>�\!�2"O�#�ꊕ��mA&�Ѧmˌ��"O^�z�21���4Y,m�D$Y&"OR=H#J��^��䡆�ʎ`I�̀v"O>l��Ǝ6N=��Ҷ�
�g��"O��	3���<�N�P�D;�����"Or4���׬`���b��7K�h�x�"O����ͬ$�J 1�d��UX��"O�p3���;=�(}���9_�=�"O�T���ʆ)l��{q�B+�g�!��u�*@�e��k,�xAm�>c!�Z�b�c�
4I\���e�Ǭ_v!�Ā�_��h�D�8�V9sD��<t!��^ oDlYT�j�.�z	�?7�!���-�h�ѥީ/��|!DH�S�!���O��mIb��6E��H�֍�E֡�$�	f���ԫT52��XAV"���d6�O:9huEiGT��WD�&R�|�OrdS0�[:cD����g��G6�`�H�<�ST���T�'.��a�й=�"!��hP^�`�gI�U���6��17H�ل�G8�m�U�@W�����e���j ��:XL�IE��D�1qbˋ+qތp�ȓq�,�q���l�Z��-�^��ȓ�"�{�Ù�a �8tJ(_�dȄȓ6Ϻ4h�kP��Srj��\Q�̄�f����(3;���F�
>�-��C.�"7�Z� F@%)Q&��a:b���4��b�:a�fͨ7F�z5R���<H�@�!2�T�i&-;����=�9�LC*^V(	֥F�5�����LP�5���zN��< �QA��=D��G'	��@@� ��E}9qƌ=D�����T�`�fL�:�9Y��=D�,�+�n�����4r���a'D��
��P�0Od��*y��a��%D��	��'�~5���H��	���6D�TkW�֖KѪeI�I��n��A�0$(�d8�S�'Gn���V*y� ���(@.P��i�ȓN�B@K2��'>�����Im����<�<%�E�q����"�[!�ȓ9���6d�p0BE Z�h֡�ȓnv�+��g�6��B�0�D�ȓhg�$�쒲~���D36�$x�ȓ$���"Ʋ9nZl���/-�����S�? �Eh�ˍ	�L�9%�nQ�$"OL9���V�+a�%cC�E�h�Ly�"O�x�B�9|��� �o��R刬�A"O��pA�����JD�9R��̣U"O�@)�ヂ*�v<pb�v��Dk%"O|���J��0G����M�2�leH�"O>�+FdS�U_(Ȉq��O�t9�e"OB�ɥ�݌)3r���\<3�d1�B"Odu����1is�d����P�����"O��֭��	;ڹ�ŁR,ib��'"Oh�˗͙�K���'�QdT�@�w"O*PT�dw�\��5TL5h�"O�ؘ�� �zNp|a��õG=,L�!"O����.��Cnm� �9pTv�y�X�LD{�򩃼J��!;NŨ%�����cHD�!�ְ%�\��  ))�"5�#��]�!�S ��ͻ���1v�$��ᆮ}�!�'� 	���J=`e&@HѠZ�!�+o. ��0d[�,�u)"J�!�	j�4�c�.A] ϒ'�!��5f��H8���d��+�HBv�'2ў�>`P"�1m �M ���r���d�,D�d�'�"3ΐ���-�2H`�8D���F
,e�	9�Ϻ��õa7D���r-żM*=h�*�-`��=��B4D��Y�#�y#���2�!��Q��4D��RG�G�P���b
�a$)��2D��������kb��ZА4S�0D��a@�V��6�c!��$=Lȼ*6'9D���
�>f���k3*J���&<D�HYtY�1>0��CC�8h{pn=D�t�0L��90�M���P�>�7�<D�81"�%�%hק�15�xPcFM;D����I�k��8�2AѴe2쪁F8D��Y�ט;�]�,9��&BmM!�d:S?���U�N�]��S Eǀ@!�D��/t����|>���.c4!� vp�(�K�P682CN<I�!�DZ�2.�)�O�o28��׍�!]|!���'�0���I�/��Yy!�gئ�R&B~i:u�I�
r!��ڬ�`t���/�R����O$`!�O�X�Ve��c�`���fh�gw!�D�P�t���+T��Qe�66d!�ď:p��) �޹2�D�wbÞM>!�$[+ ^���'�0���Ѧ"\8i#!�$?�n�WE�i���8bY�0!��LlG͉4aޓ?�]����/~�!��M�Y7�֏U�=�*���'w�!�D��E;�Y� MؼF��u�
c!��Z�Qώ	⥈V��D�B��#�!�r��K���]�m��n 0�!�D${�41���v��͇N�!�Y��1�DM�R�����:!�D\G�
�����g4��i��ă
!�Dշ!n��cr��w9�<��N�Y !�$�& @�B#I"' QY"U�!�$T��(��%M�Q����Q-:e�!򤟸p
���䒊<G�P�J�!�B�"�ڱA �d9ʵK�Ol!�d��2Q��A�Ň,9���`'�3AW!�D�4u(#-^4$D�E�ԀOYJ��� g�,dy�& IJ�� k�yR�ϐ':����J�r��J5�	�y
� ̝H�+�?j:ĝ�FAQ"B���ɰ"OH|�chU0V��W-���%�"O�t�v.Z�-�*Q��K4���`!"OZ�y��L�0֌��$�
�����"O�d�Һ'>�C� V�c���!"Ot
��P� �Be9�F�L��!"O�=�u\)
��B����(�"O�
ՈW;v(i��/=��H�"O�eR�7�H�GN 0��,�&"O�MA�Jx)6p2�˳_�A�"O�t�'fq�Z����P�4Д"O���%P�jU���%$ۋ&���"Ojh��Rh���i�bE�YFlH�"O��{��I/�uh� �2::�ԛ�"O���6L��qגLQ��4����1"O��k%��>~qd�РOQX́#"O�M0�	��r�mr� �/݄�¶"O�Qk&��	vըw �;B�Z���"O��'U
����WO��k��(W"O��z��	a����$ǿ�jY{�"Oġ;�����p&��v��8�"O8�
6Er�r�2BS�*:�Q�"O@)!E�8`� �	��ܑ3(����"Or`z�	�*��%P7�`(V��"O�Q�tW�9s2�(2�θT�phd"OD�q��K
:Ȱ�H�<q�.U�7"OT}@� �pn� {�&��)�֐��"OL�sRm1m��K#�̰c">誠"OD���N��|2ŏ�1�Ru�"O�<R����I0v�@��2-�'"Oj���$z����"Q=�6)�"O&�����/K5��V�3muh'"O$�EҊ	��4hF�O��rT"Oȭ�E�M'@�X��\�MH��"O�Y��ъ#d���!� i�����"O�5Fi�(:z�Af��iW*���"O�\9�F�:��t�O�4>thc"O�uK��Z�('�S9D�""O��!Hv�2P9�L٤:j���"O��⧨�);xpK�i���t"Oڅ�E���E�6� �»d���ð"O6��$�� ����QJ����"O�u2�@U*Ĝ�)@+��R#"O
�2a�ƀ|2�5?,x��"O�x8@a8Z�:�`a�]�?v��x�"Or����W�]!�L1d2Ax!"O`�RӃ¶#��suE�8o�����"O���EF0Y}*-2��Ֆu��1��"Oй!S��}Y�#�A�o}�	Z�"O�����\2xYs�+�>lh�-�$"Obi0�L�p�RP�����(ZlST"O:�2���"#�|EI� żY��a{3"O-�¬�h�`a1D�E�ԁ D"OD��MͰ9�4�S�ܺ%��b�"O���+բ&i�@d�7S�p"Of�;뎚&T��`'��]��v"Oh���X�gF����ʕg�*0��"O����Ѐќ����Q�7�<Z�"O��d��qg� Y�� �Wp�3"O�s�N��Y�l���Y�&ؐ�kv"O���c$գ0����@eGR�ެ�a"Ot<2��Ϧ	�4e�D��"O��(��=BuX��ȌS��ĚQ"O�@�r
�/<Fd5h�V��f�hS"O� `��aĚ��`�ڷ�'d�H��"O�A��qS�8Уe϶/QRa"Oh���.�<���`d�[���p��"O|P@	�*-�&���K��(��"O�՛�%�2��e���rtP"O,�C��؅V�P��Œ22�b�"O�Q��j��T.�i�!$Ac����"O�tR�G.w\��
#��i(0l2G"O�a���E<0z t��$O&G&�E��"O谪a�ΝL�D�10dԡd���"O@�rpG�L�CԿ"�qe"O�ՠtd�Sx$"�������g"O<�ڱ$�4J�r�3�%�8#��x��"O~݀�\6*� ��*���M*�"O\�p�
ZW ��(!���@/�Ã"O�Ea�c�S[h!�
�(�`�"O�!�R�3��I�W�K�-�4"O�|r���+����h[�	�=X "O�))�K�� Y!#.U.�`�"O@�'I�+U�x!���ʨU�T��"O�]�&d"_�Г엇1�2̈@"O-�2䋦GN��)ë��I"OX�R��F�z�d�	2� �0�x�"O�s�A^90Xl��J��g0�eA"O2	�fI�?^�zY�r��&z�c4"O^5�3Myc2@��ş@(�0��"O�@��6����<�t]�D"ONda���Μ$�$AEo&�b1"OD��o�7p��t��o�<b���"O8T���"o�ɢ�m��,��g"O 5���%'6�)CoK�?��P�"O`RaN���Z��^�T� x�"OBPku+�W������2oݾ,��"O��y(I���[��T'̺ݫ�"O�����(WR��p���v��X)�"O���ԥ\q�t`��H�r�v�r�"OJ=��%L=Z�@#�!�W�T���"O2���GIq����E�O�^�ṥ"O6��lѱQ�1�͟Yݲ�j�"Ov$��-��<��eB��f!V"O
hRƚw�`�q�[�yG
("O���ʁ�N_|��1�T4��U��"O�p3Ej՝fB���7�*��r"O�����)�� ����"O�T#qeۉr�2D󲢇.��#�"OB�J��� :�.Y � �=I��	�"O��� � �dW�|�S����t�yG"OR�QaNJ{.����N4��b�"O<x�#�
;�Hi��l$�
�"O �z��z .0���P�?��з"O$8h!�CE*�@ڷ ]�]!�G"Ojly��՚r�0�C�U�k�}Y�"OJ)Ip�U���ӡ��?u����'"O"��#�3Ad:CӦ�IO�,�a"Oh�+��]��2ȣү��-9���q"O���5��!�*8b��P�w2
��`�O~���K�S �X������&���!��P�\a���K�V�����A�!�+d(���AO�f�����~�!�d:,�6t�W(�3M��P�BO���!��з9Yt�� *m�L��/�**�!�$�1x�f�5��h�!w�3y�!�a;�)2�J���تV�C�t�!�Ę�Y�t�P�0{�2�bSBS 3g�|�x
� ̙s�O�B���Hw{�[c"O�4 ���F�R����9^�MC���N�O��mJ�=��S��Z,on��
�'r ����R+� ��c�(,M�9��'�qO��}��-x�c;|� ="��@+XK�|�ȓ~���AMS&�$�q����O$����f-b1�UW�e����2c�cWa~�]�|��F�+,�RŠ�o?02<dSbn;D��藃�*���{V�+4�X�[�O9D��@��/B}��+�>���+6D�H�D�K�DD����V-_7�c�j5D�@�C��'��D8��J>ʹt+��3D��ɕ/�?f�5:5(
�:;��ؑ�2D�����א>����V ��Mr<Z�
0D���B���� Ө|zH0(�/D��#` J(	���E��x9Ь� J+D�x`�mޞg&%���ªl� 0I+D���+�=SN�W��,�v��$D��3ҭ�M�-ď?f���xC�!�O�ʓ:x�=b���(6H�J�MS�R�hD��
�R!q`D@8\{(��TM��BN(��ȓ$���L�#l�BZrH_�<��ȓ"����� hd�m�1��YX(�ȓ}�&a[�K^�)���D.�qZ�ȅȓ:%`��.�#'�0�c���r�;�']4��w�^"���*G�*7V��p�O.��<Q�4|��e�PW�Y�Ir� �1����\��O2N6�H�F
"�ĸyQ%�)4]!��p,L8H���<P/R��N�78�!�B�U^�� ��>�-
����ў�ቯ8��0AU� �;�x�	��"kx��"�ɓ�H��I�v��Xu�4!��h�&�&$�(mS�'%џ {�؊A�G�	�+��2"5|O�b��`v�T�Wf�s�F$%�h�"/�O��ɩfbU�b��5&�6 �w�\)��B�I�O{$�0��D�mHI%��3=�̣=�U�8�ddH��b������٨	�`��IW}R��ӌ�IB�<F�~ �P�m+�w�H�Ity�ȯ>%>-Kɟ�ref�/������;8�@̓s"O@1B� oei��@��p���*���'�bn�M�'��9O�4��LLfh�Ja��?��AK�O�0S��Qo�f��ʶ�&���$_UD�Dy��I�����@��+��)TU�\����*�k�n��w��{��M`�ݩ7�z��e̖�H`�֩�R��M�'��`���iR�����O>�����~B�Ϊ(`N�b�>8k��#���8���/�O�	#�,�>��qLŲ.m|���]��G{��)��1��,	bE�e��5�#OX�n�!�D��mv)[�]�K� t�"$ʁ_��	����'4�x��0A	�tÂh��O�]�c��y�ڼiDb�k��ڈK���x�����M3�W�a~rl���
ds��D�B�N�sw����>�5�����ׁk#���
��"�Y8E"D��S��X��𬂯C��!
p�!������
ç^��z�N�$?���`A�0RӔ��� m ����CHڱ��*X e�	�HO?i�L��M{�|`Ƌ�9L|���#D^�<��!���l�i��EbKZ}"�'Ӭ����9}�Ȍk�eY
����	v��1X⩜�e��+���.H!��hʚ��f�_z$��ʅ�F�(�S�O� Tc���m�b�X���c����'����T���D��TmŶR���r�'�4t��o�rӦ��T,6I|������ (H���V�F�T��CW�i�jЦ��4��I [��(�6%G Q�X� B7f�B�	\��֯�I-Vp#$`:I��B�I�dpj8T��!XF���9ijB�I�-�
}�
��� H9��{�8B���-�
��7� ��0�����Ms2�!D�� "�2��=!��)!7>H�� O��=��-��n�@(ӗ�@�b�zQ�g��<y2+|Q��Ɍ�e�Qp 
=T��F���_���#9F"�/:D�D��K�A!�ʔp��c�M8D������/RуM��&�2�x�E"D�4���>O���3r���"]�-�ҡ~� 6�#�O��b�֙~�D��f*?���2�'Չ'���B�j=zO���W+��{�J�
�'�Ԭ+��[
n�YWmY&'~���d�M���cf�6% ���Y=N�!��S��� �rN�\�e��ўd��I';�$�Dj��Q)�hN1'�HC䉰�|��Ɠ[��sW!�)KFC�	%5<���j+��!��0�B��t�8 ��6@X	#�eɿ%�vB�	S� ��F˶ �hZ9R�ԅ! "O.�q��P�;=� �ѧT1���a"O�\�	����
����Ќ:��'剜	|�@y�!Ӱl��|��̳d�C�$?Ґ��0�T�XLh�"�	IT|7�=�S��M�ԃ��Q�bJPIɽb��*�T�<q�,\�O`���7:R`Q˒&�ş��'��|��G�@��ш�E܂.H�t!C���=!�y�
L {	b�a���'Z X�����y�Җ~t�8�� &="�BFB��'^qO��|:񏂚5D5c�+�k���8ሞz�<�t���#�9j����x�'ўb?��ьϲu�:�x�@F�����:4����*U�"q:���=f�tU�s�qy�)�'&cn��`��c��s3��S�T�?���O�~�������,Q�w��5���Te�D��:5BY�Q[�m֏)���!!2OZb��Γ~�� r��dި8I'N�Ն���O9����#�~!g�r������<ى��S�;��L�a눉{4� ٢�ז�dB�1qN�Y�������I�E�E�VB�I0����#���+:X%q�߻O�6��d8��9K�rQ��Â�$�BIF��Y\O����kx\Pѥ!���0`��1O�=�|�U)��CD�!3��<�|���c�<�ᎸJG��@�/�H^r�+��K^~�L/�S�'D� ���Bˤm��B�̍2*�N �ȓt�d$�pĚ�jnPp�ڢj�1���d#lO��G#�L����G`&���D"O(
 L�%p|zǬ�01��"O�ih/�'r�Ƒ0sfԄ��P˖�$�Şqa��Q1@͜h��Iy�@_����ȓ��dhP���hό<�MGx�'�J$cĜ1dL�	��Y��'?�d��2��a�1`f~d�'�"d�@""���(A��n��t`�'��X��V�Ed\qb� �'f7>(�'�%�c)�<O��8ه��U�����'Z&U	����t\.���&��Lp8��
�'����a[;$^�GB��8��B�	^a~����KP�k��ހsضC�
>$t�ŉ[Mp���� ��C�)� L�Rf+�5���0�,��"O�P�D#�nxh-��$#���+0"OjP0$�%j���w$��	�H1!"O��A#��{�)���W�9K�D"Opu���ľ��P▃\=�L"OP9�!����@�V шL\�x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��   �  g  �    �*  q6  /B  �M  zY   e  p  �{  *�  x�  ��  w�  b�  ��  �  @�  ��  ��  �  ��  �  w�  ��  C�  ��  d�  � 
 G � � $ �+ R5 '< kB K &R Y \_ �e �g  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE��DG{�𩊺9hl(&���洠�H[HGQ� D��݃nĪQ��E;^ҡh�;���0>����t�L���:$�0z�N�A?������Fa��d���<�rf0v
���A��
B�I72���H�A8|�J�8z�'A1O^�=�;c�`гNO���7bێ
ޠ�ȓa�m�'�R�:�,6Ή�aLR|��ē���)	,b�ga\v�P�	E���C��%+�ؠ�U�.���0�ūYLC䉕q�(���#�/�m"2+׵��B�ɝ#��&M^�p<�رo�4�C�o�����-(��qW�R�Qn�C�ɱN�<A�0�ߔJ�H��"қy��B䉈~������Dub�ֶB�	�CcΡ�����	般�
�;o��B�I5�݉B�I�-/��{l�"{L>B�<NQx%��,:Hd@���(r��C�I&yp�	u�E�RI0����Z05�C�IlC$,�'��^b0z��r�~C�,���Ѱˊ�-�Nhir �&e�B��+v�qӁ��2n`�� ����C�ɐY�0Q���@�<�A�#��Q��C�I/'=�d��J�>+�"��9�C�I`|�y�O"H2ΡA5�S3��C�	]}�ѹ��b������10�C��8eJHjfE�p�^���֒h$ C䉌+����3�7J\6`3�Ԧ��C�Ɉ Ta�˜)��ۖH�!h,zC�#7�h����&���^:>C�I BDBuA"��>u%l4��>/0C�ɏs����� 
�>t:-�O��B�I
I�6!�ό�Q��-� Eη��C�I}�������9]��"��ޢG1�C䉩G~�z� ��w( ��pG��C�	OF�)��J�x^H	�H�[|B��E*ޘ��C	[S�UB6��lq�B䉶sE�H�,@$˳G�z,bB�)� 0��F�I$K1�i���?7>$j�"O4�����.:����EB<6�ڗ"O��f�?��X�����^)����"Ot��������� �J,��k�"O�lw���7�� 
��@�P�:��"O�XG�ۅ ��P5i3"�p$ش"Ov�i��ĝ�`"TE�"�isb"OPE��zhr�����rG&hJ�"O 0��-� L4���= 5��P�"O88�G�Oo���QF��v"&�C"O@MB"%b�m	�j�7}f�}��"OE�ƚ0rH�����y�pғ"ODp��܁;�P�ѩĦe�&"Of�9e��,���*	�4,J|�"O¼i"A�|���S��%*q����"O�+���GJX����W�БB�"O�iR�������x7�bD,���"O�e�4']QByS� �"�i��"O@ĐP�!ifl+PZ;!V0,��"Oj��J]1R�*�P��Q!7�y#"O�ݹSF ;�zh�oԶ B`�9t"O<�32L郳��)$ى"OT@;c���g�p���.[q�$ S"OT���&v���A̕�)jDM�f"O���a⑌�Lay4��&}� �E"ON����ȚT�PR��@$G�FŁ�"Oƅ����U�4��c�:m�$d�D"O�����b��8�TɃ�x�4tZ "O�<� �'����ɕ6���@�"O�q��O6�:$�Q6m�vP*�"O��b�-gA*����ԫb�^��E"O����yp44�R擄h�\M:�"O>�2��J�>�N-���_S;V	��"O�tp���vB�͡�
?=�)��"O]�aiW�lsN�#�*�:]lE�"O
����@�9�T�;�cC9G D�"O~1�"�(1�lS(ŗ���X�"O�ᇀ.K}<ݐ��4�ذ��"O@hp�(^�{�r�1�ײf�~��"O�D[f퍛^��C��Ո�40��*O<�7T����z�(O'�ei	�'?,�CVś�>�uHuK�3�x���'L�@��+���ű�1*tm�'-�؛�m��M���
BoŀM�
�'M~��s�Î.��L8�C(��%J�'H)�%��|<�@*Uk��]��'V��z�H��9YT��>u��m{�'����ıYa�u��Dʤf�r���'/|��bO""r"u�HQ)T��	�
�'cn{���$��ts��<t<�
�'x�dqM6��]r��ˣW: �	�'��0�qLB�Tc �y͓�w{�c
�'�(�$�Q�w��4a��k��`�	�'� �;� T�~�,�F��j�ޙp�'�`Z	�ұ��Z0#$�b�'1xR�B��C$�H	-N�/�n�!�'VHI�B�y�F�{"�P)�yҎ�,u�����E�:X��H�hנ�y�@���h�h���R��`21�7�y�ꓼGN��!� W�9�`͒3�yb�M�UZ0z����*\��"��y�a�H�v�B3����(V4�y��0a4t#1�W4��ax��Y�y���7B��x���/8��l��y
� �8���,�B�!$����"O(�h�톤&�jE��Hތ-.J]�C"O�9�se�������*\�"O��S1*��.����˘�|��x�"O8�:&U
RI �e��V�Tm)��'���'��'���'��'��'�<�k� D�s�jm�$jұ�ZE$�'�'���'e�'�B�'���'(4�7�Z��,SҦU�m�����'�'���'���'
B�'Q2�'�@�'
H� 0���P�\, X�P�g�'��'k��'��'&2�'R��'����"��'!�E�/�S�va1��'���'���'���'W��'R�'P 9:�fE� ה�kH�!| ����'���'�R�'�2�'�r�'*��'��D��
Wì�#��ư���'3��'�r�'hb�'���'R�'=t���ˉ�S�t�J<���q�'���'���' "�'�r�'6��'�x���Ӎ^���� �o�&��'2�'�2�'�B�'���'���'�x� �N8-�����P�G2F���'���'Zr�'O��'�r�'���'B�!#D	�1��Cwא#:����'MR�'h��'wr�'(2�'���'EQ�B�8U���b%��Ͳc�'�R�'7"�'��'��'���'�N�C!�B�]��@�1��x���g�'��'���'���'I�'`ӫ�iG�˒:���D8	��Bt�P&W6�ʓ�?Y*O1�����M����Ox�e�X�|�� 0�˞{�
H�'S�7�0�i>��ퟐ��GE4$U��7\�ZqF����	�C�an�P~�2�@���@��ʈ-��%Q!� Luc�L�!�1ON���<�����)Wܠ��&�v���f�g>)n�J�b�P��^g��<�z�ϛ	r�6�[�N�Ŏ���O��y}���ʛ�U8��0O�aD�d�6Tr�cT/o�\�Y�:O��	��?���%��|���]H��؏�*� �/��{d����(�D���CA&�I��
I�p�E&V�T���+	B�6��?�X�H�I���ϓ���q���+tB��sF��rUd�'���lj�j��1�c>mb��'0ޕ�	�Wn����.]� 0���.?����'-��"~�Vd6���3!n� ��L$�P-����j�����@ڦ��?ͧw^4ı��Ԩhz��[�M��?����?A�Ɨ�M��O6�S����W10C���Uz+�|���L~�O���|2��?Y���?�ifm�2 :U��h��|%$�<w�iUR�#P�x��k����SE��L�f1kP��5@V�$J!B�����Q��YB�4A+�����O��Ĉ�8e uR�
S���!A�Ui�І�$��hH� q$�"k�N~�A���$4"�@��e�+��@� 4��O��O��4�:���!����dR�
֎� ��RZrx�G�ϥ�yGyӸ�h;�O4�l��M�i�rY�7b�<9�b੤J��|[D�S1 D�ao��;O&m�R*`�����4�OpF�C!�w�@}�&�Z�Y9�u�t�N:}��ъ�'cR�'d��'���'j�RM��"��!76s�Z5f��x�B�O���O:�oZG�P����b�4��4��1!&�M�p�*���ܷd�"!�x2$}�oz>AI��립�'k8�b���')����3�Ġ�o�8$ˊa�	�A��?�Mk.O�i�OX���O��HcƆ,o��8�&@���F��%e�O�$�<I�i��;��'3��'&�	}�`��-ģG�Q�Fg�#9��������M5�iӰO��韈|RG�J��򁪕��c���K�D�'X�8lcq�(]��I�u� �ʟԊg[��� N"�Pq�CD뮑 ���:�f��Iܟ���ӟ��)�SFy�Ld�|A��+��mI��pdlH8A� ���B�&�dʓr웶��Ix}b}��!�T튬G\ JR,<>�H��cE�q��40����4����jt(:������Z :"��.�����N�8HR�4��D�O��D�O~���Ov���|�p�Z��<�Ǯõ3���A��(���@J>G��	��x�´�yw�I�Q�C��*RNN���R�6�W��)�J<�|���H��Mk�'P6��Pg޽k�$L��fЌ%f3�'r䵺f���X�Q�ؙ�4��4�����3?�,���Ֆ90v�x7c�;���D�O��D�O����Hܸ���'��K��/(�\b"!ן��%PPlϝX��O���'�6M�-�O<Y���M��x!aK��Z(Y⋟Y~�BB�z�z�p���<��d�ĺ����O��R�e^�͐�!/n�j�{��Y�b�l���?)���?���h���$]�� ��B��e��P���I"��d�Ҧi��ݟ����Mӊ�w��@�M	{�8:��5l70ݣ�'H��iad6�Ĩm��7�2?#�����铗v�^L���+lNLp@����"�c/O�=m�cy�O���'���'��H\:�v��ɜ9 l���4$��(��I4�M���%�?���?�L~���E�!�N�[�}'��\�p�شE��$��)����WR�\�ƌ#�֯7y�8Z�ʺ��-_5�a��'�:D�'�~7��<qT��t�@���.!=��*�/��?����?I���?ͧ��d��{Q�����Jܫb^Fyb2F>H,Q��q�8@޴��'��������Ox7�ΧN���PP@ƔWa����!J��m�odӚ�	z�2��Ce�K���yq��ߟ���:(��=� u0GG�V�QY�D֝d�~��:Ov�D�O����O���O��?��������ƫ
�@�%,����������ٴqt��/O�4lZy�)A �e҂	]98� ��K�#�v�
L<b�i$���O����i��	)A:���oǽ�z5iA+�'P��D�P�
���Ay�$sӚ˓�?a��?��5S�l���g���pC��%��)��?,O o�2@E4 �I�L��P����q�-@�ìF�Z��%	����XD}"Mk��5��z�)���V���
Â�/V�bD^A+>P[$Έ�,Lر+O���B�������4�p�a��5l'�9P�ݞL�*�(#�O`���O��D�O1�r˓��ᓭi�$�[fɀRV�ԪN���Ȓ�_�ܳ�4��']��\N�ƭ1MZi���ʇJ�.�2V@�B���u�Ʊ��+s���@�D��Lk,O<ت&�,4Ψr	\<%d��bg���'���'[�'�"�'���"1"1%e��kK� 3gD	�b�ڈI۴/u�(X/O�D$��+�M�;�X��T��8 �� P1�iB�T���'���|J~bdD��M�'��9PECJ`I�<��/ך��ə';�LvDHџ�iAZ�ؐڴ���O��D������Ȓ)U8x4��Vl�p�D�O����O��4O�ƥ��j��'�"S	7ö�Q���\��MQ �/+�OԴ�'�7�B���'�H�PA�$i�8��U�.aN�Bc.?Љ*N�D'��.��纃��Oh����� g\;R#� ��ƛk���
���?���?9���h�"����bBP�p%��	F�(c��͚�<�]Ǧe����_y�cy�����n%��R��D�y�t("��ˬ@��>�M��'Ǜ)�I�ƚ� :V�K.A��LH3��0Ɓ/qb�R(	�E�q�'�J6ͷ<����?����?!��?�A*��}�%ɚAM�8'���9�(������ן�&?���|M�X����7�֌�AlD	<�Ѫ�Ov�m��?�I<�|�D��4bl��'
S�@��	UEN2L�ɓ!�G���$�<����PU��V� �0� �hy�����W� ��4��l���������Suybbp�D���ORu�s&��_�.�6���\�l�"6Op�m�G�	v�I�M���'^��Ԣ$�,lJsF�>� yI���*�"�2�i���$,��1�O�Ҽ�'�
�}�5f��������?t���BM8�y��'�R�'r�'���	Υ�]C"�O>^�J�#t&b#��$�O��$��	FId>��	5�M{O>�E�&Z�ur���08L}��'C>S�'�6��ަ瓿���n�B~��0MV�d[���51<�ST�&sz�7�
��tX×|RW�����X��ڟ(�!��j�#��B�6!�q� _�r�'�I;�M{�j_�?����?y-�F�"�AL>TٌE��f
%(��6����.O��Dv���'�����<�Y�/Y -t4z��D�m��:�ɘ�V0 ��L# ����?�p0�'��$���Qͅ�B4��b�X�ӐbE��	�������b>M�'�"6-4�6�I1�-����g��x�(����O��DK���?�Z��Bܴ"�~�Į�HĊIB�3HP
��i��7�ĝL��7�`����!w�F���Oo�i�'���F�����fa�4�گ�yR^����͟L�I�����L�O��I��`Ga~����H�(��{���ӣ�Ov�D�O�?Ux������$}d��k�āBI.i�mEa����l�L$����?��k�EoZ�<	�(LoLH�`J%K�btoք�y��ͫI7D!���n��'6�	�P�	�n*A��M��8S`���*j��I����柨�'�:6�0Xu>���O��$�'_�l��f X;
taz7�D���<b�O��m��Må�x�etU ���Y&�L%s$��7��O�2��a�n�m�H~�B!�O�m���snڹc�J�`�V��A�&Fu�����?����?����h�����c����C��y�4˴�F[�������9C��џ����M���w^@��L5
L(��	�}ډ:�'x�6�ɦa۴�.��ش��ēq�f�C��o5��z�M�po
i�e��/R���Be'�ĵ<���?���?���?I
"���$U�T#�D��������٦��J����Ο�&?��1h��m#V���~����#�(=Ĳ��.O��Dd�@�%����)����w�� �uTf�RG�I�^[]	W�<��jL-6n��]����D8dhP���=<A�����,CJ���OD��OZ�4�X���V�!�R�5zk�m�$AC>�`��	dd�,y�&⟜!�O�Pm��M3�i����'I5�@a�ѽV����@�ɟ;���Hw/�(z���L�����f���5(�F�œy�
� �~���	ԟ���ǟH��Ɵ���E�8!���L�0���"��/�?���?yñi����OwB�y�ԒOZl�P�Ϥ��HP���@�܁���v�	��Ms���T�7M`�֕��ئ���q�D�i\�Xp��g�I�h���`ι�?�%,�$�<���?����?�` �$a�d��#�ve��CBe>�?����D ަ���J�����	���O�8�`Ӡ�&S?�4;r�P�:� ś�O*�'"7mEǦ=pI<�O~�	g'T^��pG��6��(��Gpp�9�Cʹ��i>EI$�'�VT&�(q��T��a����7�ϟh�	����I��b>A�'H6��o`(�4���kK~D���-Z<^E��f�<�Ĺi��OfD�'o 7���)��I�`��C8c��&*�n��MK���M��O�EB� ����<� R �rN�L�D9�`��;=>��f?O���?��?9��?)����T+`�"3B˚a���-�3?��o�4Dd�I��4�	S�������ˑOM+L�fX��*$e�2�㣭��\����~Ӯ�&�b>M�#���͓ubp�@�8Қx�i���Γ> ]�b��OH	BK>�*O���O\��7���N̺�f˲B
6ɹr��O����O���<y��i,TK3�'���'P�cq.�:N��՚ba���������}}r�@��{�( %�Xw�;9+��B�G/q{����+?�n^�(S���K���'8W��J%�?�sh���J,�7�ܨ3��z���?Y���?����h���䔧$O� ��&NŒ);J fiV�$ ٦	Ō���I��M��wM^̑ԭ�>\a���Uբ�n��<���i�^7�릕����ɦi�'(Xu�����?�Ĩź+�F��Wm�;G�V�{�#��'��	��I�����ܟp��?�����J,Q�(ɢ7	&	��'�+���6âm�����	n�s�����~VTµ
��8�Y�������4*����OY�!ႏ�%���B�NG�'��1�n�W��4Z�l�G(X�Kk�l�{��sy��;�>iJ`���VL��#���Lb�'�r�'��O��I�M���L&�?)�(]�T�>���,�B琥���%�?y�i9�OJ��'e�7�
��YܴpsT�;�b�2��AsvGN�p4�u�X��MC�OT��H؝�"&%����
(��O�v�*�Q��H�p�c7O����O����Or��OR�?1#�O�2
gT�Z�h]�g�R�#�$�I���4^9v��O 6m'���A�4�Ы��,n�\�v�@ �M�N>����l��?)��Ħ���?!D-<6ib��c����K�D�99�ʍ�f�Or�	J>1+O��D�O����O�X2Wk�O��4bĪ�{sm�O0���<�Ľiۊ����'\��'��S23� ���(BD�aʔ+��{]��̟��	M�|
�F�\�M�+���ܑJ��H�am�<�TC����9*O�ɓ�?	��!�$�
J����-�7P�� �D���d�OD�$�O:��)�<�f�iTP�ƥ�(�D48A`Eo���a��jXb�'�L6m4�Ƀ���ަ����<s���3��R���Q�W��?9ߴN&� Zش��޹qz���',��ʓK<p$₉/�~��cJ+bR�8����O<���O����O��Ŀ|r4+�+�P��%m�,X�æ�%b���D�r���'t���Zئ�]70J%aѨ�&��s���*`4y۴-Ҕx���甲䛆?OzxH���m�b�,Z2�&� 0O� m��-�?q3J+�d�<���?�r/�mL�i���O5'p�SD�	=�?	���?����dئM��K͟���ڟt�ud�1)��C�N�)<�$}(�,�W��Z���ԟ$�I^�ɲ���B�ɐ��B��N�A�
�`	`�҆� �t��5L~����O�5S���h@6��u�œ��<��X؟��ןD�	Ο E�$�'�&�9�E�V� X3A.��$hPm�v�'�6m�M'��0��4�4�L�"��yd�	�F��t��6O�!n���Mk"�i��K��i ��Y�}���O9���� �:zfLx1�H7��� ��l�Py"�'���'tb�'�nO-vG�)�FD�'^�����J����
�Ms��_��?���?aK~�����C�Ѷh� 0!WG��^�%T��I��M#s�i��O�)���).c�}�uN=�� X�[9��Ǌߧ_/��c�|�F,�O`��H>.ORݲRL��S�h+��X6�8�c��OJ�$�O�d�O�<)ƽi���8��'#*I�t� �Pd��*Ɂ�*��'P6m9��>����ҦY�ܴ���*�";�ν��)��xE˟ndM��ij�$�Oh�ǍQ��'j�<��ԿSr�`Jx%P��&s��*�T�<m�iy��'v2�'�2�IN�}�๡I�R��I[v��=����?���Y��v��Qr�	��M�M>��"_�$Τh�� �=�x̹�gɤi-�'�r���$(�	؛ƞ�`c1*�![V���e�W�D�����W�,�6Y��'ixA&�L���D�'c��'�D٨�JcЉ���2HG.��'D�U�4��4I�9*O��Ĩ|��#E1>��QbSfɸZ��Lb3$�]~b�>a���?��x�O����4��pi^!�t��N͵/��ؐM���2�O��i��?)d�0�V2_��kb)��z��i�IG##D���O(�D�O���<�W�iX�%ìKn�:P�C��D[�'-Za��'��6-5�I���OH��2c��`:��Q` �2v]���O��m���lZu~��o	������Ovz���%.���,�#r�܁�'��	���ȟ��Iҟ���t����##�n�C#@ ���Z�cT�
��7m��Hi ���Oj�D?�9O&�nz�aq�G+1���#��?�p�2�������}�i>����-����L@ЫK�^�C����7����
��N�O�rK>,O�)�OƀC�C��	PiB�W�,�T��O��$�OD�$�<� �iѶA��'@��'ǂ	ԣ^�@�Q��IH�L��@�D�j}ҍ~Ӏ,nZ�ē2�tp�.m�푦'�L��'ܜ9�C�[�+a�h[���TA�T[@�'t��اh�!��X�&BP6*��PhV�'�r�'
��'\�>����P,.�c�/��c�����ò(lz	�	(�Ms�ŕ3�?Q�R��F�4�\�u@ƾ �rыaKϜ25� :Od�oZ�M��io>(ҵ�i���8m:�J �O�� PiQ���<9t�Y��| k��<��<!���?���?����?1���`��(Q��A*m�d�DM�����I�#K��4�I�%?1�	:t��Y�Q��xN.屔���p)�O�oZ�M�g�x���ɜ�G�TX�6*E�T�0K�o8�J X�@E&�剾i�
��'�,�&���'�Q &i�"-NJ� t,��~n@��'��'�R��D]�(kڴFS��#�mqȨQ��4x�a��<D��ϓI��&�$Gm}��'��'n��n�`�J�*�a��r�(�&b����� ���3 �$�����yp4�͵ ��xs"�G� ˄��0=O��D�O���O��d�O��?ŋ4��5u�nI��Gx���A�|y��'6�\-;��S;�M�H>�`�0,���{�D["Pw��v�ۖ���?��|�4H�>�M�O> �3��~U�9eDB�GS��uK]�1������TF&�O���|����?9��)sbź���~-L�0%'������?�.O��n6u�`=�������E��c���,�����EB�P����@B}҄`ӛ��*�?��&���W\�[v'I� ��B#��*lz�x��Ɨ�ex%����+�ٟ�	D�|n��	������0�d��jZ���'���'���DS��:ٴ�<��1NՄH�Ĝb���-���"�A��?��%p��\_y2�iD�5:�f��
:��qd�)��! 2�zӐo'�f�l��<!�3��Tp�蟘H�'ʸ`�	݁F��]���\�5R����'��	Ɵ�������������Q��G��p'恹#���l�(�@7�	#.�����O��D:�9O�Xoz�i���ҁV�kQ������DA�ޟ���p�)擂y�t�n��<q�N>f�� h��#完2s�\�<q�*�{f��˨�䓌�4�4���^`�3�[�`�P��W��''����O(���O��W��F C�r��'ibn�#JQ�����C� !����>��O��'���')�O^q�G��E��5"��*|�LPz���,k��=*g���&$�9+`�&��� ��36�^�sN4�Șq��G۟�	ޟh��̟�E���'T���r>�AY�7*	���'��7͞`����OP�l�v�Ӽ#��ç�.$�7K֚=9b%AN�<9��?���i�,��a�iW�	�pW�O>Fhݦ$c����:_����$��A�	{y�O���'�2�'Sr��&\l���E�)��}��f�$"��	=�M�����?���?�M~Γ�	�� �aK���aB](f�޽h%P�������L<�'�?��'~�l �F
�<mIU��a�������#m�`�'��ih��H���|"^���� ��hp^AiQ�8�x� 	������ğ��I���Ly�kӚ!��O�1���j���Pǂ�GQ�y�6O�TlZ@��}��%�MC$�i��6-�,Kad� ��q |����pN�Ԣ��v�.�hD�=v��|!K~:��8`�i�qc�(	$XY¢�3M$���?A���?����?9���?a�M�����8�!Eb�'PH���%�	5�������?�ʵrb7:�I�WۄU��`y�͸E#.L�k�,I�� ,�>�6M:_��$�O����h��T�g� �ȟ4h�kQ"�� U��s��@����)F��1B+@�J!2�'���A�'iZw��	��F�$�O0 �B�,<���E2Zx�Z"�O�D��E�<�7�'q����'�?���)O�{��c&���&pgB_�7J��ӟ��'��6-ܦɯO,ʧ�b���+1X�j��يy�"E�k�<H��ݹ%����'z��J���8'�|��֞-�d]����c���# 풔q1��'���'���Y� �ܴ4�ڹ��W5^�h�栁(qZ��á׫�?���9���$�C}��c�ڡ¥��)D�z��2�GH�����I�U#�4U����޴��d)@�<����O�v�hj�PeJL�nX���	$_,@�����O��d�O��D�O�d�|b�&ޢ>�Ьh�hQ%BFVȩsK +3E��� >r�'yr��d�'�t7=��1SAʍXvΠJ�jŗK���ab*�ߦɱٴ7�����O\��]t��6Of�qK��%Z��#Wwt�C�:O"��-���n��~y�Op2K��U�a��3A�B[SK�'K�b�'7R�'��	��M;��� �?���?�*��&Zr(��D�m�^q���̡��';���?�ٴl��'W�E�w���s����"�5���#�O6(7)�F1�xs�f#�	�?	���O�(7/4>����r&��(�8��/�O>���O����Oʢ}b��r�X}qǒ{{Xm9���K�]��$?-$��'O87� �iޅ[s����(��j[�]Op�2��}��شBu��w���i�im���,���0$$��P��Ak�5 ��CQǓ3 �zD�l��䓢�d�O.�D�O��$�O��d�6�^�y��ø�HEEɒ,>�5J��ES�*I��'$�����'�E��'E%-11*��&f�Q�v'�>���?q�x��tAˊD:ƀQ"Q�X�@��Dل�v\JkL������!/p��0�H�O|�M���3
+�ċ�C��5���?���?	��|�)O��lZ�9l�e�ɍE�@�ZT'ÖL7���m��*�D��� �M��j�>���?�i؄l0-��K��R�-�@�zs)��6_��<O\�D(ro�����i�֝���C̖�S��J3A����4�y���	�����ܟ���쟈�:��؉2�铈��p��,�?���?��i���Ocr�p���O�m1N҇!vj���'�13��jǊ�V�I������?�B����Γ�?y��Sx�? :�W�Ԗ9ؘH7;5��Y�鑿�?᳠-�$�<�'�?Y���?A�(f`���C{��zCfJ&�?!���Ҧ�1�(���������O��tQs���\�1�V.؊�i�O�4�'x��'_O�)�OT�@�@"- P쨠솝'Od���̰&D<�����I�?1(��'�$�����щB��ea�ޖUn��0h͟���ן@��ӟb>e�'9�6�C*ڸ�щ�� ��-��� L@�e��O���M�?�X��	�s�l��*�L�Jf�� �ɴ�M����M�O�u�����zK?-���'ut)(AS)�v�襪`�h�'���'�"�'A��'y�@��Hy�j��F0�f���a�K>���	����@�s�h �����:e��)�E_�s���F���0!ҿi�*�O�O����Ǵi�dN��=����<t�Q���Ri6�$߃7*��{��M~.�O���|z��qaf?&�B�C�� 2� ��?1��?a(O��l�B#X�����I�eX��%� 6X���Zb/I/|  �?�P_� �	ޟ�JJ<����o��P�-ŔcB����A�d~�+Z�)l�xpD�5��O~���4-�BAT�vU� Ȟ����acoѺS&��'���'���ş|����t��U!ѧ~)hm"R��ğ *�46
!�,Ojqo�b�Ӽ���8(2�@���]��Ě�<�3�i�86����ApD�ʦ��';�bukH�?%7%�)�F�i��ʤ��9D@G�hR�'��i>e��ן���П��	9(�hy��-�*0b�-A7	O�}�|���9g#<q���� (�(��蟨�I��MS*�D����ܑ7�O*_�\,�A��~��	�'���'��O�i�O���²f�r�"���5*�ɻ5��+�Rq�L����ɻ/���v�'�='���'�������9���	栚UH�E���'_��'3���$W����4yȪ��%�Zͺ�ǣ�8�4Aı�JIS��x�&�d@}�/bӦPn�M��ёyH0y��#�<�DA�i��ȁ�4������2��LF�����_�@&�V��L�w�M�IQ�D�O8���OD���O.�"�S�T˰��vB��5�f�kÊ�6E�μ�I۟��	��M��n����٦�&������a3 ݨVm@�#I����x�I����i>!��!��-�'� =zd@	X\�����d�щ��S�#��I�OX�'�i>����t��N!��Ņ�[d0+�/K#�J���ҟė'�d6m_�&ے���O��d�|�u_�4.ز��0�,�DH�N~�>����?iK>�OX�A��	�m L���.��}y� `����g�D���4��ͫ��7�ғO�p4NB��jue��!x����O��d�O����O1�L��6�O�4��*؍~����%	{�t���^��(ڴ��'��ꓥ?)�d��O'�KՏ�r�2�z�G���?���[zhP��4��$�	.�z�������i�ě�F-P��QF�$pRD�|y��'��'�R�'d2]>��v�w�|���'�&4Cݲ��M#�hگ�?����?�K~Γ;��w	Yy��BG:������o�����'��|��4�
�F��1O|���ቦaæ��!FǺa�f1x�6O���X��'�B�&������'����v�0,�D�gj��P<Y��'R�'�bR�0�شP�*����?��z�|a���e��*�⃥?L��R�>��i�|��%�dPyj�Ȑ��_~@\�5�UO9�ɿ���&i���-'?�ˆ�'��	�I3�\��4��Y�I L�B����	�����͟���f�O���L���!�8[��Y��4Y&��dӂ��OP�Pڦ��?�;n��XQ#�?�h8���Pע<ϓ4�fey�2�m96m��<���jo�ѫU���X��Č;ph�c�G�,t�Yۖ!N�����4���D�O����O��dF�| 2��X��hK�� �T���F���@LuR�'2r���'K�3��g6�؛wOV�dk��in�>����?ӗx�O���O��%����'#�V�����,$��)f�҃ApJDr�O2,�Q�X%�?��;�D�<é�t٫gk�kx�Jr�� �?���?����?ͧ��$Ϧ5zwG؟� ����r���5��Tq$�q�ʟ�A�4��'����?������b*��mד?����AG9�P��d�i��OJ�X"����'D����?m���}Q d΅����ɉ�0>��ן<��⟈�Iǟ��J�'C�H�Aw��|y�-Y(+�f���?���fmߟ���禕$�Q���@?�M�g%�.�&EJ�R��=_�Km��I�"�6-5?)��\���XQ�`3#���&�c��TK��O8�iI>A(OX���O����O�X��H8�a5�i����O��Ĥ<q��i8]�E�'"��'��S�TM
�+ �]�nT�f qb~���	5�M�T�i�O�ӫ!�b���OE<) ,��j[��6���(YGμ��Y@y�O�l5��dJ�'���pڦ	ތ����"|�p�'��'�2�O���>�MSЬ�B��Ћv.T%7�f䒆J,y�����?I��i��O��'2,7�:|,r���.(_����G��oڮ�M�3d��M��Oz���/����<�7�a6���:?�A8f@T�<.O��$�Oj���O��$�O�']9��i���3�\�ÀJ��\��W�iݢ7`�O>��O~��8��QԦ�]&����#>��ف��	0�v��4-`���/��ɐ�W}87mn�� Z!+��͑������b\�"�8O��AN�?Q �<�d�<!��?)c])y����A�-+ӾAQD�N��?9���?����������џ �	ʟD��JUh¬V	cސq"Nf�gC�I��M��i O|9H����`��i����2���#���Ӥ+�?X��d�%G}�7Z��G���h�QZ��k"��G��`�`jП��	�8�	ΟE�$�'�i�+�������n򘙪��'��6͊�0X���Ot�m�|�Ӽ3 ��81$�$��L�<������<q#�i�b6m���Ԯ馭�'�L]2s�W�?	�,�F�T)Pǩ.�+s"��
��'����<����	������c�^��C�v��Q�a��(�@�'	�7�5]��$�O���)�9O�<:B;��hqL˖P����`�`}�`�tem���S�'g5� ���-@�D���JF#\X�j!��	x@�Q.O|u(���?y�'0�Ľ<�1O�#������+)<���E�?���?A���?�'��D@��ݨ L͟��R��,c"dݘ��	A���K6 �ϟTX޴��'������My�x\mZ�n�h���N�Μx�M�3����R ��Γ�?�v�N٪���������h;&5ٗ�D'EJ84��	D�D�O�D�O���Od�$ �S4Z����U��Ye�l`��%&DU����D�I�M;�F��|j�;���|�TQ$������"\�p��Ŧx�JO�mZ��M�'G��ߴ����)l��ciѸ7Dh0�
x����M�;�?�q#-��<A��?q���?A�`!}����,�
�+m�g�j���O�˓0s�֊֘B���'R>)��H�0H㴐
����	zO%?q�X����ڟ(�L<�OV����ؘ Ϻ�����`dfYV%�1P����	��4�� "����O�A��)�3������C�D���*�O���O�D�O1���S<�V�Ih����Q�
�J�8�cIm:u��_���ش��'�8��?�'
�39p*8aǙ62(���sB��y�i����5�i=�	�8���C�Ov�є'�t5#� ��~�̐+�G��u�f�'�Iߟ��	������<�	e��凹}���	$GN&��H(�NְM&6-�%�����O��d+���O��nzޙx�o� 	�Y
�*��-:�9j�	�?�4J�ɧ�'z�e3�4�yr������Q�D/���Pv���y�Kڼ�H��		e<�'��Iϟ����
�\�
�<x ��0�C�mE���	���	��'�7-�8�$�Or�W��b� ��9�Zx��ˆ#a�t�p�O�o��M{��x���:y�������=a�E�5ǁ3���N�z8T�K��`�`��|DA�g���Ē��F���B(l{`�9���-�J���ON���O��$:�'�?)�!�!R>����r!����*�?��i��H��'4�b����];>s�(R$�`*�i�(5h,0bf�o�(C�4/��
m�LSC�h�P�Sh�]x�������T�������������C�����D�OR���O�$�O��$����`"LB"x����`˓x���c�5p�2�'�����'�B`sTg]�aB�i�&�	h@F󱃥>��?!J>�|����3HN�p�ƥ�Ւ�m��0��H���~~��&w0t��)}�'u�	,n�n�tC�;$��Da�H��	����	ԟ��i>��'&6-�v%f�D_?` T`wGs'x���_5d���Ʀ��?�PQ��9۴^כ����8E�J�m.	�"�Ń	
�8�U�*C4�7�|�@�	G��1Q��O�\�'J���w�$D�d!�9T�@0��Qª�9�'��'�r�'�"�'u�Ԙ�B�� |�ڜ��-�q��,�O��$�OxmZ���'�T6m'�DI/g� �x`��_d̠�5��ِ�&��S۴m�f�O��C�i����O��2f�?z�tթ"��l�D���_b_���-rƒO��?����?����
�;�f�Ni �k�e�<Z�f�����?�.O�mo�=#U�A�	�����o��l�8��cV�P7j��ږ�߾���b}���܈oZ����|��'%������ Y@���<U퀭�S��UD⅁b�7������@�ғO��M6n[҄P6� �?�΀�2A�O����O8�D�O1��ʓ��&ܖs�$:�$�68(��2��� ��,0W�'N�Hz�⟐��O.�mZ������þ0����&k�vl���ٴ^���B9ߛ6���`��2���kyy�ň�v'��y`�6 q���5�yRR����͟X��ܟ0��ݟ��O�xe�F�P�P��dITB#[�8�+ rӈy���O��d�O`�����HĦ�%��p˖ʗ&B�-��h0e��i[�4؛��0��	)��6�g�T����	h�s$P�x钕�j�� !A/<Nb.J�Iny��'C�� s$�u��7I�|��Eѷ.6��'���'q��MSr�����Op�y�b��ɠӀַ4F�h*��7�����dMæ����ē:��MR ��-gQ��k���V4�'̢���Y 8 (ғ�te�ܟ(B�'a�[i��^vJh��+��'(�Qp�'��'��'O�>���/#�zu3V!�@Ɯa��B�Z���	%�M#QE�3�?���
K�v�4�Ҩ���¼c�� ��B�Pfh�31Oj�o��?�ش4	�-��4���Prd��'҅Z@���F��|�!�R�LJ� �4�D�<	���?����?A��?�֡�$a�C���0�F���F�-��D���!qj�֟��I̟<'?��	u�����!�%*q��"O�
$R�:�O���{�$%���ٟ��V��� x�J�-ȂK�l��oGr�0����ʓ5�5��$�OP J>�+OJ4yaO��.����C��	�ֵ�BH�O����O����O�ɵ<��i��(t�'��+����u�D��XxR�AQ�'�P7-�O\�Ol��'"�'��Y'�4L��)J�6��ds�7]��i���Of�bܴdX���"?������"cĿv�$�Ц*��:��p�Ԯ��<a���?q���?!���?	���&òq���C&�RG�rec�"n��'�`o�L�p3���W��5$�<��K�-�N����Z�%[�kґ�ē�?I��|"�����M��O�H�	��.���2�i�!P6����J1v�!���T�$�O���|B���?y�<�(=���W�>n�����$�my��?i*O,oڽ����ҟ4��R����{�q�LCɐd�Q<��d�E}b�qӴ�nڇ��S�d�8P��mâǧv\� jt&��బi��6�z@*Q��S�;��DW�	!%Q�]�"g]G�\�+�+{�0|�I�����Οd�)��Cy��lӬ��V�̤BT*UE֎Xi��;����@T��
6�����NyB�iG.Y0@f�%r��
!c��3��Pp�r�� nr<n�k~��r���S�3M�	6s$�%;��Y�"�D� ��8���ry�'j��'�r�'
bT>�椕(k���;��C�6�A�qd�<�M��Dۿ�?���?����cf���/7g�8���$`��y��&�,U��nڳ�M�2�x����G4ٛ�9O<��D�]��$��퉍O�TH�2O�ɐ�H#�?�� ��<!��?I��D>.lµ 7�@64�89�׆� �?9���?�����Ц�SE\y�'�2�C�?��EfC�%� �H���Fc}B�i��o���?�d
_D�xaX�X& �o8?���G�F@^�P6����'TDL�$ނ�?��a�	J�͸M.E�P���<�?Q���?���?a����O��1DHD�YUH�
�N?L\��Վ�O�Dl5Q`ٕ'��6-�i�mk1J�,ɘXC&J֕D�8��z����͟|�ٴ ˰�
�4���%"V��'V4�Xd�ԑ��$�L�V@�]X�k3���<ͧ�?)���?����?�aᒮ?���;�a�w���h�T���Uͦ}z��˟���ܟ�'?�ɠ*. ����E�2�[��B !X��*O�Dq�%���^�I��ؔ�����Q���ERsW�M��LaP��l�㞪�2�HX�	kyB� :UW���(�>���17掖w���'���'~�Ow��<�?q������x��Ũ9�PЙ��M>b�E�ȟ�۴��'��ꓜ?����6o�7s��Ũ磐*$��!���}FP(�i=�I�W	�K��O>q���T�}F������|���
��Y�o��D�O���O����O�<�8	aP��ʘ~Ru��O�R�ލ��ٟ����?�p�}>��I2�M�H>96�֏`n<�R��i��I�V�^�gB�'�7٦�ӵW�]lW~Bl����-�RB�����+�F=����0Qa�|�X�������8���ʐ5� A;�i��q;��ӧ�����	sy�Dj��bRe�<����򩈤��H�ć�F���m.*������d�O
��d�)"T,Z.���H�j2?��E�cV�C�EP��{������͟,�|B��5R)���#��3slɪd�Y*�R�'��'Z��R���ܴJ7&=C�I��[,E+GK� &�L-I4�3��H��?qG[��o�;G���C�NG�z4-C��B`�r�{���M��@)�M��O�%��c�=�d��<��i4icА;��P�B��=<L%���$�Op�D�O*��O����|r�`��Px��h�d�y:U���,"!�V��5i��'RB����'� 6=��eCRÉ}��ZA��h���*��a1���S�'5���۴�yb��,r@�+���-ԑ�pa��y�bE����^�'A��ן��ɉty�d����*d���aE�Z�������Iɟ�'�87mˆ@HB�d�Oh��q��0�Pϛ�)C`��P��x��O4m���?�N<9W�^gYz����HR��� �����
2#&��ϋ;^��:��;���%M����v-��%"*�� \� ����Of���OF��7ڧ�?�@� S�Bhk��:%W��3�$�$�?)��i�>QS��'$2+o���杞~��R׌70�T���Aܻ,b�特�M��'P��IU�e��V����rB\9-h��K^>�Bb��L0$�D��/i]��$�0�'-��'�2�'�"0O&��Q�dr:c�ڟ�R-��T����4+o�q���?����䧥?���R:y(�� fs5N��m��l��矘�����S�'S���7O$���K�p�,M�D�%��p�'����ß�ᔔ|�^�(5I�	�
�I��E:���p��'K��'�R���DQ�h:ݴ"ﶼ��qv>̓��XPP
Pˌ�;�z!�jf�F���Z}�'�r�'�r(�dF�=	� Q�cBWzp4%A@Ñ�X���=O��D����x��~�	�?����l��v�[.-����㙂"R��I�� ��Ο��	ğ0�Iy�'w�����$)$Þ=��b����I��l�	џH+شE���s/O�9oZv�I:o--��C�+�.�+#NV1rT��'����ϟ\��>_Ԛ�m��<)��u��8r �L7�T���"%2-9�D����Ծ����4�$�D�O@��H�Tl�h8�,ʚ|��|���B�2��Oʓ2t��P�6Z��'r2R>𐫀c��4�Q;'����5?	�Y���I��%���ϟ� �Y�v���f�ZY;6�T6�,E@���B� S�j��f����?�	��'�V�&�X�ᩆ�T�q��H:K�&D���L�	ޟ4���b>Y�'� 6�!%���`r
1O�lhs��0R���3�J�<���i��Ot�'�B�L?,��e�g�I�m�D-��"t2�'�~@�i��I�r��IrB�O�!<�����7�|R�d�����d�OT�d�O��d�O����|J�jͣ'Ep����	,Y�@y#'�a���	�7B�'c����'��6=�d{���./"`�SJ d4�!c�+�O�� ��	I�946�n�\s�D�J�@<9s%��J2(a��u�|���3R��RF��Vy�O�2!�B��$g��'�)Ӎ	}4��'q��'��ɸ�M���
�?����?�D΁18�T��o��" �C�d	7��'���(��ӎX$��zN]�P!6Oͱ	���#M ?�BL�C�"�����'S��D�2�?Q+Z�ځ
"`~�a��?9��?i���?9��i�O>��1�T�)�^PX�	9m����k�O�En�%8��(�'��7�=�i�997��B�� �4k�<4�|�cLc���	�����!CC�n{~b&�4���Sܔ\ɤ�@,b,�,P)֣ ��(rѝ|bY��џ��	����p��֗5�Z9*B�A�<�%�v�eyB,m�Jp��m�O �d�O��󤍮AZ����P? �Nd@�K�P[���'�r�'�ɧ�O�x�#Ù�,5N���̈&J` ��A�%����O���t� �?��&���<!�*��p�v�06_	O	U���I��?��?����?�'��d_ɦ�i1��� ƶ:�NQ�@NC�`�X봬r���۴��'����?���?9��̘����dȎ<�7��%)j�%�޴��$ހW�f�@�'��O����n�zV�Y�Q�(*�@۔�y"�'���';B�'����P��B�(4_�E��ǋ�bc��
a��O����O>Xm:mM��'a87�"�d�CZ�d(�σi^و���w�|��'��O.f���i��I ^״HJC�.4l~E*K�=�~�0D�	 4ab�D�ay�O�r�'��cXu�m�G�",u��8����)��'S�I�MK��պ��$�O�ʧT�޵��X�?�4X�U�Hi[Tn!?�V_�h�Iڟ|�O<�O�4 r�F�v�b�#�:9���WH�4GZ�	�a�*��4���+��RD|�O����E��F�>�h�L]"l�H�OR��O��D�O1��ʓ����,Z!��
:�X�����=����W���4��'�X듄?Q��_
J��iF+ە�:M��.��?��h]2��޴��D�+TE�������=$���Z� �xd��n�L���iy��'���'���' 2[>)PӈG	։��`Q3b�� ��$�Mf)���?q��?H~z�u���w@�Y�c�
��8�#��(x��xY�'�B�,��)��,��6mp��q�d�&�1[�͌$��b�t`Bd��D�r-i�	vy�OBr
Q'�*�K���b�!0��֕�b�'Sr�'��	��M[��J1�?���?!Q�������P33O�� EFC+Z��)�h}�`wӎ=o����x�C/L�	��A�B��͓�?�`@ې?����+��$�����C�6�$י��(B��r@ǯ+i�!�ēL���S�)6:�y���Kx$���Ҧ���gyB�c�l�杇�2����G�D���{�����	��M���i�7�_�
�7-z���I;FQ2,{A�O�2x)"B��3�r�3!�!T�����D�ay"�	8`t�b�'MA�X�tG�Uަ�k��fN��B���|�R���5�>���R�	@�bb�&0�����M˳�iPJO1����f��\Q��Ն��::�0��G<}�M��ɲ<�� ��-4��W��䓬��R�z���1�敧`�Ab6�Iefa|b�w��0�t��Oڌ* Ή�5�x�б��8P.�;S6OНn�O�!��I��M[%�io@7MF�8x�!	�n'8�08sӨ�O/,1@6fe�B�Ax.����\�{I~���v��c�پ4���� �M+z����?����E�J�H��
s\H ��/�����O^�m��2!��Qכƚ|�I�|�$4C��(�1��i�>��OЄo��M�'z�ιK۴������P#����B��E����Pڑ�؏�?Q�=���<i�ZE	:���⇙Cc(�Š܆|(�"<�R�i�*e�$R�,�	F�d��=`��<��C�8d0��8��D�Dy��'����)�T>�Z���EEڔOs.�tS�#F�E�����`ۑM�D����������і|��8i���S�);6�R�ccB�:�x�
aӰ@勍l���U�W�@Q�,� 'U����O6�l�U��X-�Ʀs�MO=
� ��D1
KfĲҠ�0�M�g�i/�)!�i��I<�� 0�ODf�'���S�1ng2`S`�ϣ&�� c�'��Q��:��K.|D�򠝥yL0����_��M�S����$�O�?]�����A7�M�%�G�	h��c��%Q��"~�h�%�b>�k��զ��%k�F��,�:s!�PN�J�ɁŠً��'*��%�ܗ'p�	�=�u���<|m�""AH�nBZ�����	B��,�IퟄZ�� z���ȏ�N�vĊP�Si���	��M#a�i<>O� ^�#P1I� ��E�0>͚U���A��K�p�F�ūQY��r�2��˟�ò*�({�t������@�zB�.D������2{�Ƒ�acU�#v�IQ�����4
�̨)Odl`�Ӽ��f��3�|�j�dɜ�,�z��C�<9�iM�6������'L��	�'+�yXŦW�?�Q��S$.�ʄ&�*k����C���'h����Iҟ��ǟ��I�Lj<�c*O�x6����s��'�7�&[�4���O��4�9OjE�B�ʅ��@�t��7��Ȓq�g}��'2�|��� �)�\�K���VWЀ�&��P~�%a1����B+���c�uA8�O�ʓހH��u�1䥃�}��1@��?����?���|*(O��mZ�L���Id,(p�#;T��u3B�k��	��MS�b��>����?I�\�(Q͐�3�j,����9@��H
XRpXo�c~"�[
I��E�cܧݿ��@	63#�4:M,5�8{���<9��?I��?���?!����T|��AB�2N2��0c�4i^�'8Bgz����5��<��ix�'U�p�vL�s��0�l�_Hf��|��'(�O�(�{�in��0�*����1���$)MT�J����W%"�/ZX��ey�O��'�r��9@@=���W3*���;� U���'o剖�M���V �?A��?�(����r�N��^t�bm��h`:�����O(hnZ��M���xʟ�	SoĞ3�t%���-o>���@�4���i�L"k4���|�C��O��pH>Yы�,rR�C
^�<v��¬�?���?����?�|�+O�Dn�+�ƸY#Ϛ�q҈ز�O	�8�xHL[ya{ӆ��.O�7��1�f�yC�˿'8li�Q�`�mZ��M#k̛�M;�On�9S��>��<#bV�P�D���=H�i��C��<-O"�$�O����O����O�˧M+$�z��l����FK�Ĉv�i���p_� ��g�'F��w��X���J�:C� +v�@�x�(oZ"��ŞdGĩX�4�yb˜�*� `��)әKhંA��yR 4��MX7a��#(�0T�҇����r�ށ�H�q�I�p�H��2���Y��	�i�,!����BM5���SE�_����@c�'$xDb�j��j8��+����TY�跅H6����(1�sPU��[W� M��t@�@�RW�Q`��J�� P0�+ON�"�I��@O0��p�B��,}b��4%�
m�a��٬
H��(��t'�����L���J@��� � 	  M�W�&B�Z�Ȓ�(�R��Km��8���)�Ρi(L6^aJ����C)�1��ie��'��Iz��+L��X��E[�5h�%�!j�<�d0�d�O>��Q�ݱOf����H$VѸ�,�9j�<%���i���'V�I]��aட����OR�	ڷ_ؚp���C�ɺ�됦\9^�'����៸b"�S�����͊C�I�C��D_��� �MS)O�����ݦ��˟L���?Ѡ�Ok�ÀD-|�C��&({lL��J�?؛��'I��^��O��>�fUE�ҵ�+��v��$�6G{�`t�(����������	�?K�O�˓,�Ƀt�޻#x1��c_����S�i3�l�f�d2��֟�: bЪؾ�uդ	�Fh:�DU��M{���?��9q�*\��'�b�O&4����+��X�` H.��C���F/1��O\��O^�DD{ޠ:'��*��u%��^��4mZ�����AZ��d�<!�����2嚾f\@�`!;���(��f}hÕ��'�b�'�2_��bЦ�P��:�o1|�����@ ��O���?YN>���?v�E?B��P��R�B�@1��m��U.���?���?Y-O���K�|��Q�����t"U�`�9@Ŧ5�'2�|"�'b��).�b چ�����B<V�hl��cJ!S���?	���?�,O�P�ժ�M���'���r�ߡIF�1k5"77̬ @�c�L��,���ON�D�&q�J�|�p�J�`�l��� ���d�#����d�O�}�hxUU?%�I�H��+��5��)�3Ve�i����oz��O<����?i�O�?��'��i��GN��҉�r�H�d�<E��S���b
��M[��?���"eS������㜔+@����H�:8�7-�Ox��G�S�
��/�d(�ip
�o��B^�"�.)��6M�d�oZΟ��	���������|�S���=a��j�d�.�f��)H�GR���s��'��	^��U�4�I�0Bn��#�[(|��#O��-��4�?	���?i@	��P�����' ��@**Z���Yj�,�b@���O���'R�	:b��x�����O��d�O�dPT!�,
�8�Je���f�w`�˦m�		l���L<�'�?AI>�6k��r�Y�Z}��*4N'c�֥`�Or-����Ob��?���?�-O�(����<&�H Q'Ńai�9���J-^�'�4���$�0��u��bANP�3@=7j<������M������?a*O����4��Ӡ+ot	���ͰXl��q�藕!�6��<i���',�7R|P7-K�_3<���k*6�28�"��6'�	���	ڟ4�'�,XHE�5��wp:(q���8r�w���?6��oZןt%�x�'N.���'��'X����lƄ$֨�fV ;K��o�����Zy�eH5t$d�b��k�%n<��oߢr6�d�4.�,�'��=����	F�V
s�������
 K|��������'EZ��C�t�H��OpR�O�H�=Ѿ�H1.�utԸ+sh��|���o���@���*lq����I�O��I�|n:� ��u�n{���B�3]�F� !�iM�Y���'n�'7��O��)�u���~ߜ˧��1yU�rANJ(D���)��E����y��iطGɚ�",+�ђdcоP[�<o�ޟL�����vJ�]yʟ��'�a2g��k��E �C�W_"�jGO"�I/ׂL�H|����?!��L沄(������\u�X7z���ire�kHhO���O����<!�@ލg�Ȩ����J8,IC���=���'�� ��'��'��'���7,Z�1p.�fc��)q�� ��a��ՠ�ē�?���?*O$�D�O���(L�'0�1�c�Hg$�s�L�D����9���O��Ĺ<�e�2)�)�2S���Yn�PAj�+̌\��������S��zy����҈�<s��|:���2o8$R�o�y���?����?)-O���B��G�S�?`�y���Z���!g�?u��t�۴�?�M>�,O��
���O��O�`�6ʑ.U�h�� �q�!ڴ�?���J�Q1�q'>)�	�?��{kr�
b(��X&Ol�H�0��<aW�¿�?YM~��OI.�w�X��h���1<%\��ش��dI�=�mZ�����O6��^~¤�NI�!�̔�MW<dق�́�M�+O�K$��OX�'>E%?7-�fr6�R�aٞPe�MhT�9P���?X�>6��O�D�O��G�i>=��i�97�����,�"Y|Љ�I��M��@��?9����<���PsO�;8K�u��g	���������M���?���&�|�)O�C�dԀH*p�Y�d��D������1����<�بm\��������2u�%u���BY.D��	|���d�r@ʓB���T�{��yb#5G_���Ť9;^��\��r�ϐY6b�x�IDy�'� xp�lķY�����Œu�^D2p�
�W��	џ ��]���?��'dnL"p��S��/���k�46�P$�'z��'5bU���������\��+�Q�R�t%���d�OJ��(�D�<1�C�?Q@�ӑ#��3��.'h%y�͋=��IП��ɟ�' ڬRC��~��#��`���B� ��6��K��E��iw�P�\��ȟ��I*s2��矄��>U'z�!�ޡ[�\�r�_��u�ܴ�?i���_;9����OR�'���J��_����f�Y&H><��3��A��ꓓ?���?�c�X�<y���?����4KE1n�J��H8D�6|!�����M�(O �äa��]�	Ɵ��	�?M �O�n�/P���w`ݢ`kd#2h[dq���'�b@��y�|"���&_f�M+C�ذEq��86(^;K]���.i֮7m�O����O���u}r\�2�nB�ڽ�$=�(��d���0�>����R�):�<1'B�,% �"�d�N U�i?B�'�/�� [L����O��	�-�rD3G��N�P<;�IP�$6�O�ʓl�:��S���'��ޟ�����ܢN��!�e"�>k��izR
U�$KJꓒ��O���?�1-
й���yѢ8 P�٫r�l��<�Át�����D��ҟ<��qyB�X��0u#S&�!`��&[�����>�(OF��<����?��t�$�1&љlx��Q*}0��P��<����?����?)����D�D �Y�'X����U�ͤ42H��3��\�n�]yR�'���ݟ��	�`c�>���M�J(��ʏa�2�ڑ��馵�	͟��	ПT�'Uh�
⋧~��6�de�כGzP��o�j�����i��Y�P�	֟��=	x��It�Ă�?1�xb�������h�q���'�Q��4��%��I�O��D����X�c�-8\�=X�@=  B�qELJ}r�'�'��q��'�bP���'O8)�D�RS��S֬+gb�lZGy�+�'f��6-�O*�$�O
��
S}Zwy CRI���,����Ȧ�ٴ�?Y�<� ��4�����}���[�C��D�6IКɐ6��˦�Z"mX�M���?y��ʖZ�4�'�j��c�.��Pj����m���i��P��3O��Ļ<�����'{!�oN�J�v`��!&&��ݱ��f�j���O6�$��w��$�x�	����ȼEG�iaw��U�����d�&�O�xI7O��ȟ��I؟\�LY+Q|�p�C3$�x�bK�/�MK����y���x��'RB�|Zc�(U֛z�P�� )&&�A�Od!�?OB˓�?����?-OD�Y���-3㠔�E0��ԥʺ�&����0%���� q`!�o�e�v��-Z��,��G�=GXR�	gy��'���'��ɦ~5�yh�O���Sfk��d 
cІ� ����O~���O��O|���O�M�O�)�g�}�XQ*kۀ6�4�u��g}��'��'�	)�b� H|��a��Z2���]�i���	�"[�f�'S�'�r�'��}�!�'@�H1�����4�Bc[=�| kme� ���Ojʓ���P��D�'��$��*wV��q�`�c<X`*��GEBOz���O`�Q5��O�O���+�n�1R��2�R���m 46�<a�KI����B�~
��z������ß���(b���
_)3�{Ӕ���O
@�0O��O��>��_8?�%��
�CY0�Ġ|�T�A�'�����	֟ ���?��N<i��u�b��raǺu'P��0�Qf�,|K��i�Ҧ���|�(O��D�7+V ɶ �K^�A�	��0)�\n�ğ��	��`"� E,�ē�?���~� }�T�i ��)pq2��̸�M+L>q�+^�p��O��'�H?� �� P�Sv��9��iǢe�ҹi�f2>Vb�<��C�i�����z�
 �0)�8�v����>1DOV��?	-O����O��<�T��;W��b���$��RV��$C)Ҹ�G�x��'�ў��%PuT����"�C�>`e�� D���H�Iߟ<����ty"�T�*��S�B��Y�P��J��҅m��u����?ъ�d�O�0��k�OZ��3�_ ajDx�)H�_�$�y���S}��'k2�'V�I�7�0�2�����_e�5�
�a�"`���Q�>em���L�'���'����yB�>ɗ'��x�XT�r�t���V٦��I矄�'�l�����~R���y��h4�����=��P�`B0.��"QV�����t�I#���	^��''�	�"-�ΰz_qV`p3��,6�*�n�VyEԴHab7��O����O��)�l}Zw�b< ��"S��l���E��
�4�?I�@Fx���֟>&kd̅���(C
�=���a��cO�7��O��d�OH��q}RV�)��?:@HS���& 1b����F�MK�I��<������?��؟H�C�"�*�k���oƞ!�E��0�M��?i�'�U�1V���'���O����l�' �@�X�L�d9�!��i9�IƟ,2� |��'�?���?��LQ�<K��+)C ,�q�*�3���'��1��>!)O8�d�<)��3�^�g�,�Sg�`i�=�4K�B}bK��y��'@��'���'��	%ez�Q���`�ذ�i�4<�&*��G�����<����O��d�O\���B�p���C��o�RMiQK�,p��$�O��d�O���O ʓ�-��;�R<��kI�t�J�R�>9e;�i������'��'���y��W�5� +�O
6y�؈�)��lʶ��?����?Y.O:�2��[��'�8�U�O3�$�Kw+~���Q�z�(�Ĺ<���?��SK���>YĪ��6�XU�@�y���;����E�I�ė'�JykU��~���?I��6��,B�Ծ.V�ʱ�C
]�(��\�0�	Ο����q�8�'���?1�"M3T�栁��ȦF�eB
wӦ�8*0bQ�i���'���OԌ�Ӻ�`Hɹ�,l;�/ԁ岥� ��-��ş�xw�{���IRy"��ެq̞,sF��-J=)��ܵD����S0en7��O�q���m}RX�`c�bA7p`\(�pCF�y5F��d�,�M+&��<A-O@��;�S��'��qMy�1LG�x��ȸ�Σ�M���?��'dnĹc\�x�'SB�OMh�ғX���Q��=���Q\�̖'&��O�	�O4��O���o�.l�p�Z�2y�f�\�R,^7��O�I E�f��������\��5I<% �b#� �E�k��I7��DqX1Od�D�O��D�<	qeǕ$����sh=�p�޻]��X�w�x��'��'���Ɵl�I#L��]�	ŶES�Ěr��8zxa�1�I��p�I��h�'r���a�}>5XU�{
D����/yD�+��>y���?������O���6����Z[J�[iԚs�\�B��xD��?���?!(O���a�NK�S��b�PVe9bȒ�Þ=�ʥyߴ�?������O���ޙr��>�R�
:p@V ��o��p�LJË�����GyR�'W( e�'*��'Mr�OD�1S5�+G��-(�ؤO�0��,���O �$Y�)�X$��T?m��n�.�)Ĥ��'.�#�cl��˓D�F8	'�i	��'�?���q�	�?P �Q�JK�Y@��!.˿2��7-�OP�$MG�b?92
�4~��E	�f�%C�x	 !�O����	\�|��O ; O �@ÆM[�%O2�yr)�2+�"���$R�iԼt�&x��^'L��L���G+3�.��8?5��bU��T�#jѶ`�v�SC�N%	%��nƟF˜���(	S��2�?.�N���M<�z@���K/X-C3l��Z��`i���G���r���:9�z���=n>�x��f)&��Ȣ3$G��R�'r�'�z���T���|����+,�J�V�Q徽+��V�T���S��7�q��V q���1��		�B�2̓�k�Ɋ�,�C�H��3͔�6�.�B���<9t	ɥ��UC/�{DRM'�H[/=dri)we�5\���H_��B�d�O$�=��!؃#��5X���K܈��`fh	��m����W#H*��Ezd�
�" ��<��U��'K�q�%kӌ���OVI��ի4�Q�S�1h��!�O~�D��`%$�D�O2���:xp�w��m�	:@G D�d�	(ywD���N~P��[�:E���X�8���2���UnB�G�0T�P`ڵ--�C��'(<B���?酷i���h��SO�,��)����;$������?E����[F�T��\	 �V`A���K�ў"~P�i�vت���ZG�xar�́*>��G�'副C�
� �O8�Ģ|2aO�8�?a$+��y?��%�Rq�!��P�?���Y2��X�Oi@�����~X*�z˧��`%�T�0'��q�� �O�邆�;��)��$>��"}"u�!.*�J�O�M� (��u��^�4�r�'��>���0�(4!�,�?=4���L_�4H�C�I5��Ջ^�]�@��3�G(o�.��ĂW�'\���+� `��P���&x���>	���?q
!~��t@��?q��?�;0v��p/�cي����SJq gC�=���@��'0d�p�gə����S�? ؼ���)4����`��^���h@K�T�х��x���y�q��'ǚ��D�s�"�BPeZ{(�E�W�'�	57��4���=	����Un�/d���#�G�!�E�U�T$(4m��� :�K%UI�	��HO�Py���={�����C6窭Z�nC Lf0�b�d%-�"�'�b�'���������|B�S�c�r��0j��*���W�%~�B�/�:��͢QK���<���1aP��u���	��ڸj�T�i�0]P#����<QՃ��[V��ԧH�*�vER�ˊJ��X�	���E{��D�y�`�z'F'N��`��@�jO!�&09ba�!�����3�d�471Oj��'��I�M�D���4�?��h��x f
�z�nM�VG�
��+���?i�
Ȥ�?�����$�G�tϛf�$T�B���7�ߢ?��r� *�p<E�9L� �Y�I�4����
cO�(h��B�%p��!�%~��x���?)��i�*7��OUpֳT��g�0]3�p� A
���۟��?E�4��F������;*-feI��7�x�aj�`a饌F�uJH �%��,�h��2O��p�`\r!D��?!����J�~,z�$øP�|�SN�#P��՚��+K(���O�,��� ��!�5%̣f"�裐hE���dY>Y�A�5	�F�
4F�*L@�Q�3�!}RL@)f�d۳aH�1X��t��l��>�'j�*2 B����U�W&e��2}ra�+�?)���?Y����O���4,�l AD�2{��Ĺ�\̓�?9
ϓ 0�%`W�ug�SG�Y#�A��I��HOf��UeL�_xt��&��f(O��D�O�����u�j�`���h�~����?�!�d�0&��84	�1�d�(I�V�!�d��1��1��I]�=�;GO�|�!��߶9��,l�B����	l�!�dH5O�0їOلy2 )��bE�p�!��o���b�J�e?~i�'�"�!��
z��0 ��
(Ă]k�a��t�!��B*0�東��	�5�M��ޡ(�!��7H1���h[�7����3�)=C!�dԼoPp�"p%��=�0�C煛<�!��߸^��ۧ��}�Z�"S�5Sc!�dF%S��["!T���
Ef�kP!�D�b����dN�:������F'<!�d�Lb���,�:}�J�C5!��"|�4�t��8i�2�ʷ��+!��5��y���)�~���!��m�!���v��y{�o�@#"�y�!��� f���.N�f L�k�,o!��Jz��e���04�����/�1W�!�6����!΍�P�����N�!��"�ft�Xh�z�m�*J�Xy*�"O���o�1,jU��B;/l-�"O����	�`|�E���!g�YHg"O*؉�@�zʀe�dG 7fx��"O*uu�TKf<��ĉT:��"O�E������*5o�?8�Ait"O<d� �Р�xa�N�&T�UK�"OR�
�7�'��"��=���ȓO7�YWN�_��Y�/�_Nq��C�R �tI�5`UPn;C�V���UqWϓ�5yj�a��=Qi����Dݲ�C#2��ٷ+� ax�ȓi��h񉅱!,(5�GNP�BO������1S&Ӻn��	�lC�a#rЄ�7@��P�ђc��J� �ޤ�ȓF �z1�f�	c�D]\ค�	�(������ր��^���ȓ&U<XxE�хQ�2�lS�[O��X�|��ԫJ=wn��ي&�����?86����5���0��_�@�m�ȓjr@��D� 	_x�V�lβ��a2��R@�$b��Q"i�mT�|��S�? �t�@�x��I��f�f�ة��"O����^�!(��Z��=a�"OTL�r,�-�H�Dm�"t�Z��w"O��u��:��ĸs�
�f�x2"O2�褨���9��˜�k��ͨe"O�ݸw�ШV���!ԫ�&�|m[�"O�,#��`����,9���"O %��e�"��M*C
ՀR$Np�G"O�1��
�ih�]HƂ81�	�"OV�[%�	%3>�-�֠��L�HS"O2�b��>�`�� Aԝ���B"O^P`So˪f����'��=V���"O;P	/�f=A�y>���"O\���X�,�V�4\��"O��
�ƕ?_n�P�6&��`��"O&�#I�em�ӁC�Boڡ���8�l��)��������#?1�RuV��!��VI��"	ftZ��'\�D*D�>0�>E�$L>h[���u']+2���Y���(�yR�V���� h<"�r`JO����|Lx�h
דj��!��|���� &�= �A��	pX�УnW<��h�H��K|nE����4-!�D�eƺe�B�ܢj���a@�p�Q�L�Z���'�����;JP�x���2Y[���$�I,1��ㄅ.�O�m�4쏮g�r�1��R��to���:&,��'���$&���,k� /ah�U��S�j�Ѷ"O�c���������K�X��^�t2�O��M��]�5��H?��cʁ[z�X�!����D���4�O�XsE��-C�5zC�	�����×<���(�$:}��+q���њ��{R*	AM�H�Bϗ!{��r-�
�0<)�E�j�	�VA (
1�N�$U�yR�����SEĪ��$	��'0QAJ�P������!H�\9��D+R�
�k��M���+��f��,tnz�BƏQ�c��Є#S@�<��˽uF��jN,5�LЗ+@y��^�=��`R�A^�ِw��x�OC�h�C��*�lQ�w� 2R�k�'�4�s���
UI�`��5��r��)s�� ��M#"��fD�c�nU*�1�6��	�'��M��ώ� q�1���5����?���GȜ�%Ϯ RE��!|&h2������8���s�	��9���J��}��=s�e� ��<��Mw#�X℈_�<o��s�cK~��r������0V����fT6�?��&�-"��ɫZ��K*��p�$܃{�L�x�Ol����K$8�@1bK�5kc�m����E�gh4c6���T�����SX�v�I��?Ac5��$�`�Ʌj�*E3 �`[�u;#O�%���JjY�R!N{�6s����YX�33��%	UbT��l�G�xX��S�jX�V)^%;6�O����J�(��Y��ͭtpް2u�'J D#�-�(0�n6�ל7���9��űIՄi(B�z��Q�E��(�G�'Q�L��.\�WZ����-`̍��zm�I�BeH==�����(�McF�m޸-릯��~��O�iP']� ���Ļm��ʣI*H��!�7N�=lB�#��T"���!�޼�D�Ҽ�8�E'Z%F�x9" ��O.�i%㱟0��!�?!�yעٵ�b 9sW��X��p=��OL�@�ċE�&WF�cND! e�!�f� 8�:Q;�e$}"�>f�Q���H�)��!�@�w?Y`A�3-Fʉ��#�@ેe�M��4d���A�d=�f��� �t�H!D>zYXdIדw����F$��}�v-�<�	�(�T�CF��/g@���*ߣ7j��>AƥNhN2�� ��U�
��U ����b,�L2�a[�A� �N�A­^?(�2�<�4���[w�0�dt����g`����8�q�'e�h��M+e9uj'���he�UF��2 ʔ�Pe�@#�rb�!�٫\i�m5A�/J�>���L����$�����	(9O^̐��ϥ�$�����DW�l�'2ړ�$��w��Ic` 35��[@��[�P(�竞�*)D�k$,�!F��L�<i�$��m� ��>>�Ȩ�JD�B�`��	P)�g�� �(���C��6m���æy���t�a��
Ɔ-"1{�(�c:����h @y��8^��q"kP/:�M�
��!����g��#����0�ř�l؇6�P�Y4���_�\!�II�iH����V>�5��Vy6�td�!DhԢ�G@#�@ b��'�@�X���'E<�i����~m`��B^7#�nDAfEذ�x�0>�
�+!M��P�e��m۶���@���D�	>��l�6�O� ��;���� �L2��ُa�bT �cƤm;Fݺ��'O~!�	^�&l�5�ƥ_�&��ED�vA�Ӯ�Q��y�F%
��t���6�����#\O P��d�9Zf�h􁔡w�x3���H��	o��bL$*���9C��O�Y�,�f'��'݊�x�L]�i(�0HA�<�dʝ�/���	b��a�v0�'#&�H��H�`fH0�4F��a�O���n?ͻU������8'fd:�^ h�2X�j@PH "��p	��r�@ߧP<4���d≞!xi#����H��qOPh�a�%u8dr�d�|Ҙ#p�'�J�Kg��1T�t�+V,X8-w*0/�괄�d�Z�"E��	�9�p����&F�P5
�I��Z+0� �N��t�Do(� C<��-O-�M�͜�W2�*����'�B�ɖ1�������>OX`�ƞ�a\�ɟʈq�}��I��p]��3�Bɠ\"��*�K�:
�!��4#�P�C$H�n?�Ȁ�U�i[�']~E�ۓk�JX�tQ�"�b��" ]�?�T���\�4��%d�����SZ8�ȓ2��l�5C]4%�����-�Q�|X�ȓS����WOJ�l�Xa"����7��ȓ�R��Ƃ�i�.t2�؋C z<�ȓw�rYct�E���)��K>G�p���pr�=�@DP�sd1Y���:Xԕ�ȓs�#2�ˡS�D�xᅔ6/�@��	]�QH��s��<��(SN{��������6��N��q�#wd��ȓ~��=���|D��&]�l�=���^��7��3 ^ցӱ���kvrA��WD��K �)?������Y����ȓ,D�eK�,�0�UA�"킼�ȓ�d Fd==(��¢ ���2�E��m�
��t�IV冼��77�Qk�@��D �� �4 BD�ȓ|�|:���<c{��kLk0^ �ȓ'f�$WL�u"͠��#oy�ȓ$@��J󬝊*��7鑤]�����*��bb��'��	��^�m�y�ȓk0�8E�C�<h�%X�EV8�`���f��	����e(�I^�s������\4���]�(�k��Ŝ!�X��%Zm���8� q���t6p��ȓK�ʠ�Z9:����7/�.jj5�ȓ7�Y�dǓ�?x<��DA�ІȓM�B��1�H�|�I�� ����MC�LidBɬY����t��9aD��ȓm|h�U�
~��Y+�ݹ[� ��s�p!����lk�Ặ�ŲI��e��|8�����S-ظ"��+PZ��E6( �Ƃ��>-��� �8�J}�ȓX^Qs!�*�\�a��ρ.�|�ȓ*t��	���Iy@E��r��ȓ+䘀l��]��9��Խ3�̠�ȓJ������R74$I���0����7�y#���m�6�	�wР���R6N(�R�W�r����-Z�^X&]��lC������D��@��OP�hF4��3Y��&�'H7�H3�����ȓ!��Y��<젷��*N!���k#�\��L2NE��͟{���ȓ
�z�B釓?\�hi�����a�ȓ(T���`B�|��Y&aC*
X�ȓw��q��-ϒV;P��@b��;𚕆ȓOG]��پ����gD�'!�����𐨧�O~�!x�h׎
���ȓa�E+��  <d	�E|��Մ�xȘ�갋9C݆e9d&�4,X�y��S�? �5Q�.O�ر3��AF궽H�"O�U���e$^9���=P�p�w"O���� �8y@�"T4��4a�"O�ap��-sF�zR�_?<Ă�"O�M��-D J���H�A��^�F�ʂ"O����&R��z�h0�J���"OM�P`@z"�(I5OU�b$�G"OB��V.�\�F����
�-�@"O�Ĺ��.+����n6_f���"O ��Ĭ�8_���U�fMx�kR"O|��A��}tb�@V�B�@�u+�"O�X'���н9��<t^��t"OrX���V�/~��� �ư]el���"OR3#H����e*SH䅰"O	 �FL#.��a���l�ТD"O6ǂ �	��| ƬP�"O(A��NY`@�i;_�P�{u"O|��I�p�HdP!V�H��"O@�����+��(A�"PRA@`�<I�)׻R����raפ{ | �p��\�<�����b���-R�*e|XQ��V�<�D
�I�81ٓ��)�@�2�
�{�<��(�'~|ز,T"<@"çGt�<����k�\MPӠ��T��
FY�<�F��X��=P��-y�x!��R�<9a��x� �2
A* p��R#�b�<�"���3�\��bݩkY$�3�Pj�<	W�D,h���{�jZ�=�`��φf�<!g(±C�vɣCeU$(Zd�WDh�<ɡ ��U����� ^�8PI!�g�<����9���Cb�DE�bY�6)�K�<Q�f�+R�z��fl�m�0@x��K�<�ć3D�.Õ�̝r*�X��/�]�<�cEJ�S��[���j���t�<��E7bfP�2��
M=���&�{�<�a��,+X4 w�z��4r�%m�<�W�B�x
Y�F�}G6d���X@�<� È@x��*��C�vְ�ҍWw�<��Z�q�"��x�mr���u�<Ƀ�ޒ2r�90"jȭ
����#I�W�<$���&���M�{(*�)T��T�<G�F(C\�`I�f�~�Li;��^F�<����.X1C�Uy5@ ��B�<�%��YG�	��
�(��T�áEz�<���Zt����#iU6�ġ]`�<��(��"����-^6�� -Y�<!��U�wB�!�9{(�k��`�<���N'U�I�(��2+l4�SC�<�@��-���y�
	h�0tf�~�<�b�4u hA���;NqL\��"`�<�IȮKN8��sa�[#�ث��-D����f	��8���g	|d��++D��2�m!h%=�5�ۃoth:��)D�<��7md)*��ÑP�j�I�N)D�,Җ@�6>��7a�S}.(��(D�Ԑ�S�i����T��9a���0e%D����L>�L�j�#� �ʕA��"D�l�ë�*z�H����V;|�fX�!?D���C4�2@u� /��p*N D���0en$i�e���	��J�*D����� ��b7�O�U](I�)�O���N44QB��$ p�$�F��(~m*B�	�W`�:�3|ʰhZG
��8�RB�ɹO,�hC��" ݔ|kf�Q�x�RB�)� DP��� �R� � _/wX�x�"O\���k�PZR�HS��&��XjF"O6�1���,kq���kn���"O.`Z ����+��ӛnf +�"O�Bɚ�Y:)P*7��$(7"O���� �dM��7q�%S"O�D��S�_]n��d�4�d A"Oh,�b��J&v���_u�Q�"Oz�Ae�p�kĎ;0GNh�"O�ݻ���"�R���i=�V"O��B���xh���F��#w �k�"O��8U�
L�ʉ�`\�s��)��"O�	��m8x���eW�R��"O�)�7䔾+����e�$nq:#e"O��mɕzg�X �WHn%��"O|�9���]H�c֥Etk�"Oy��2)bB�B�A	$rCL)��"OB�Ra�����"C�A�iB8(�A"O��I�ԁ(BW��,F9l�"O���$��mN*����G�΅�d"O~�G"��pIF=��L@(yfl���"O��8J]�}c.��t�â%W�D"O����i���(ѱG]=KK�DXu"Ol�A��ې
�^d���9.u3"O��UeĂl������ lH!"O�	�J2u�I��Z�%��y�"O>/�
K�)��&ԓ �,�"O�]��K�>�� �"k_�v8��0"O�lق�F�}�ۗ
�\`]�"O�(2C�
��m��۩i[8̳V"O,83Ae�+���ѦBPߪX7"O��$��9��QKuC6��}( "O���G"�%ULA�ł��*�Y�"O
)�p%�:b�B5"ą֬��"O\�Z���:�*�북��T3�pj�"O���g��!$7�	�%�7\0�yȡ"OX�y���x�樉vF��A-Vy�"O�h��yT+N@-z�Wy�!�d_`0��Db�o�lR� ��!�dʧ�\Q93��1i����@��G�!�$�.T�U *�Xc�nV�\w!��&pD���G�r��)8ጉ�g!�d]d?��W�8�!"B蒩 ���ȓ=#l5��皪y~ʕ���G�tP����1çfR�W�Bi�1n�+8l28�ȓR�p� Tf��A?0�˶�U3R�<чȓ
��L�W��8z��o	��t�ȓ^������g8pЭ�����ȓK��411������>M��ȓ'fP��ahM
T�:0��6�F��MS@L2O�<�V"�
�v9�b�Ph�<a-�j6��bn�]��凊O�<5+8��9B��!~7�1I%��d�<9�-����LQ�e�`N45���_�<q���'���Y��O�!��pR��`�'��?M�6��GJ�,٢B
�{3�Б� D��񧫍'P�p HSM�  �d�D��p����<Np�X��)M�~fLn���8���EN(w��6�͒E�ȓX��E���E��MA��A*	mJz	�'q�����k� �I�7|ژ��'8̝�P�6вY��c�=m.��k�'��@jt�C�u�
+�-�.nY$b�'���UaN5<��S�L Ĕ����� `�'��I)j�ye`ңP�����"O���eƵON<��f��<S�"O�hp!�ԀD&���Ϟ3����"O��ELNЕ(�6DyR�p"O� �@^.�`�!��+i\<��"O���/�[����$��6���"O��J������3.��v�@�P"O`y��'�,i��-��I�Y��"O�`:A.��_�ⅹ�k����=�"O��(s�7��m��/=���)�"O�̑2MH%RxP���]�#�0{�"OP4��L�g�FMK��=a���:�"O��(�jL�zp��d<IF ��"O������o��j�:J״u��"O�U"���b��;�b�m�J �3"ONu�ӢZ�BDkƣ�=}l�Ze"O���ܓj+��DH�s2H�"O
Y�R$݄�C�-�)s��)"O~���ĉ�eU���bl�i���V"O����烺#�1�� %�`�x�"O`E�#N�`=�L&�ۛ#��Ȼd"O���G�1��%���<�"%"O��`���2D4䁅�|��"b"O�:׊Oo��P;$�Оr���iC"O�I����E:4� f�/}|I�"O�PEI�\[�
����W"O��Ǉ8��<��B��.�}Q�"O(0��BܓW�P�xrg�R���"OƵ2gJ�L
���ЀA�� �"O��FM�z�:�F�V�6"O	��� ��|� ���44����W"O.Փ��+Oc�UP@$��.�����"O�Pp�B�H�Ќrb�O�_ctf"O؁�F�z!�T�fL��s��x��"Obu���zPZ���A�8a����e"O��o��ct8�0���?�ܘi�"O�415�I$�~�n>S����t"O���Ǫ��̠ g�{�ԩ�"Of�Sᔆ(�v�4,@�~��b3"O�����Ն4�P�YfO$_j�=;Щ�D�������+Xk����i,��A�I��yC��
�*�Bg�Rwx����ȅ�lu��ք�q�r�q��i��Y�ȓCa0��d9v�Y��Ƃ�Z���!fF!:"or+�u3dO�:��чȓ�	 b&έjh���H�h��ȓ�Cw���T����G�6]���'?ў�|bn?` ���J�HG�P4�NY�<iԉVq(Y�VÑ9� ��b��U�<���Ô}��R�2��x�/�S�<�q��/B�XhA@:Zb�kS��V�<�c���)@��k��u���hR�<���Ͼ������]�b�����#�G�<����,�Z�
e�χ5s�J�m�h�<��(C�N��Ա���Fy �z��I�<���C!� 劕�Y^t�p�nKA�<1�D/M��@��d�*���b��u�<�I��ODF\1�H߆�����F�r�<��JÔ[��P��x�l�4Ho�<A�b�,7`�y׃ �{Y6i+4˖j�<��Ĳj*��0�X�}�T+ �h�<� A,T��ȷ � #k�9��E	h�<����i���Ї�;(��8 �	g�<)p:\��i�1K�`���p�m�]�<� :A�h��8<���C@�q��LP�"O�%��e�2s`d�s��V��`���"Ob���dߞctFI�wF�!|�F	�"O�A��jO3eQ-�BK�x�8�B"Op A��:
�8D�  �,�S�"O$8�U��l�H��W7��Eɇ"Op�B�H_6,ڐ��WF&ŪP"O�Z���+ �h���8�0�"O���e�ц`����םCF�"Ox-���23�DM{��M2���"O�!Ss������u�PX��A0"O<9�E�Q�{��3e����0"OnM1�*��-��4��@ tp�"O��K�"�	>
8:�d+f��b�"O�uh��*�;0��0Ud,�"Ot��u �T\� 1&b�����"Ob)B��0 kz�q�K���	j�"O����:J��Q+�PVt)�"O�YBѯ^�2�����>jG�z�"O~d�&�9l
̴x LǤk4�	�"O�`b�P�^�Fɘ��D�B�
;o#!�D�#50L�E�E��yR�X
!�dZ��5��R���;� ^�{!����	�Ѡ�c�_}�*��>=�!�܇F 9#��YτY��i	�	�!�?
 n����6\!^�q�G�J�!��B>bL8!�� ��v��1�!�-5����d��-S�&�
��O�S�!�ė��]�mB�*�J��"N$<t!��_4
Y��U�ŵB ��P� �!򤛷)B�����*\��6Q0%�!�$\�>j��WFPbD|�b�'���!��#>z�!���'4ly{�L$Z�!򤜛2P�Q��+/��gϵ7	!�Ğ�)/��q�T�N�8���f���!�$�����J�!�'b�0�uH�;m!���:or\3��2���&��02�!�$O6�L��*�=+��E��f�!�;}�V(��`�ML�$S"��0!����bXh%��5R48t�T� 8!�䍹_p��*SF'���Ҭ1R!��4V�؍�M�=m����4��5:3!�]�^��iՃ:u�(BE�.?I!�D�0�Р���Xp2��s�@!�$C �=�!d�+%J +!霂E)!�d��#��0yR�%MI*�ôE��	!�D�X�^m����"�8R��(8�!��~���PjP(B(�g�!�dߨ	�\P����?�{Ĭ��i�!�D�\�X���i�\Yc+^�Dp!�AZ#� U.qߎ%�G+��FP!�D�)l��#J4ܦ�3�(M!�Xd[ziZ�e��rɌ���X-?=!�$]% P���cI��� j��-]%!���BI^ SӇͫv�Aœ~�!���)@Q�wױ��L@s�G^!�]D�&m�Sn�p�
�!%%�5A!�$mǮ19�H�,����7aY�R.!�ē2�Tx�ʓ�e���p��DG�!�D�>(�)8 �_�<����P\�!�Đ25B̙S��(s��y��I�S|!򤒂:ڂ��S�-TF���\�Ni!�ĉ�\���h���TOr�ˁ�<U{!򤇺!q�]��!��LL�X�&�*Z�!�� �"Fg�%/���0�b���,�p�"OJ$�Q!�n���P4�k��!�"O��J���9O��c1a@�j�A�D"O91���sI^��󯖮\p-
�"O �@���:N$$ٴdGxn�Cc"Oڌp�ό'd�|rg�:g���4"O>�XO�-�:�s�j�`1~�	2"OV	�7�ڇt�N]ȥ�!W$�Y�"OvTE�\�/0L�QSe�br��D"O`|�#�޷0�
��ccY�*�� y�"OT1Sb��%P]*t���Q}W�"�"O��B�ȕ#V� �������"OZ�H�"iʬ���3Iv���"OZj��M�-����`�]5p�("O$�5F;S~ܽ��&Wm��@bs"O��1����`r��re��!��Mp�"ORI���u�\4�s�� �P1��"OFh�&!߉6�PZ�/R�ݰ0"O
I�LU�B�!A@� ɲ�8!�DN'+��(юS�x"�y�`
�S!򤁧I&.�+��Ld涸9v��? !��%Tp2�k�� ٺ�xwe ^�!�Ā��zu+t"�- r�jG$�=Q�!�D�S�>T�@OH[x�3@ꊟD�!�$�r�@�3�8Y����(ʕ>l!�DT���H�mX+c�~9C2-��Y!��?V
��hdaJ<~��˵�I7P!�$��~F���A�V�3^���q��8?>!�d�{��E�D#T��I�b�!�ލ��QYg#޻*�&�3��+!�Ѯ7�D�z�H
� �zL;pGF!!
!��9�h�ɟ1�^��l��8�!�D�`(Àk�9d�,٠���!��ʒ$hT���ͧ3����u��m�!��N�Lu�q�F눂y���0��|q!���	m���KuA�fT(Æ�OjY!��ʕ?ϴu�&Z�&-������V�!�D���lL1�K}9����Z�!�D�.0%�Y+�g�+e��q�wn��Yy!��5�8=��B�Mɦ�	҇�,k!��)W̹����x���`&э~c!�d�*��kՀ�,>8��cFZ!�$O�8lJ�� M\��M�É�+{c!�DSO�J9AF�4Ր��r��6gG!��$z%�XP��$%�x\��Θa6!�dY����[�I i����E�$k4!���
M�.8�A�/"5*t�⎝�K�!��U�fA{ϡU�L8���T�+�!����bY�eFp��djs!��_�$�,e��^=O�H��cc�+B[!�$��A��� �cȗm̤���@��!�Dh�P!�fB$�e���Z�M!��H���`�u���2Ei��=e!�$A�5{��ʅ�Ȱ_	�i*6��aP!�D�,+,���FC_-9c�� r'!����d��Ek�%�t5���Si1!�$� ��}�#C�!߾�φ0!�P�1⤼äʞ��,���� c"!�URN�|���-�аM�7!�dF�3�$K�Ǿxn��4͏D!�$M�f�B�τ{kb8�f�X�!�D$]��$jBd�s0ɐ�-��C!��#U�@���h�d�CD̔�o�!�DG�yB��$nʝ�~�h�k�	�!�� "�J�G���Jv���|��L�'"O"���Y�a`6�f
WC��"Ol�·n�+ �:H����8�2�q`"O�hi�
��[f`�c�'Q	9�ri#e"O���F%�,n��U��Į;�nȳ�"Ox�%��*����!��v��q"O��W���T$
�V]eD��0"O�L�WB��4 ��)���"O(�@D숷ͼ����I�
��ur"OJ�ᰬ��L�\®�A�0ؐ"OH4���V@2x=�!�H$>��Y�"O�9`J�$����B+խs��aؑ"O0tc� �4 ʕ9!E��x�rS"O��P�$o�a@��7D�4Y"O�%�S��*'�~y��"M�R �"OT1ye��(L(�E�T�V��"O�tq$[2F��e��Wo��9�"O����=mT�2c��	Z4tЇ"ODe���&W튅�l]2<���2U"Oڔ�dGS�}�0M�Ş�Z���"O^B�#_�.>j,�g��1+�\Y�U"O�X"�G77�LS����]�Đ�A"Ob�qd)ɿJ���JF�-6���yR-$�l���� q&a;r*T�yb�5���s4�
�dt�|��G	�yҁX&�j��2�
���5:t��?�y���CTQ�e�m@
A�6�@��yB��k�I�/�k}�)��k
�y�E]�d{fEe�~�fc�+�y���-���e�aɸ�r�IW#�y��\fl��t�X�T����j��y�.�R/���P�=�j�R�H_��y�X5P��zr��6
�
]��y�
�S�)�E��%��;V���y","{I,\ѦcQB��)S���y��^HT(g������G�y"�LDa�@ a,���9�yb�EX��� ��1e��5���y2�X�"�x�(�&$��U���5�y��@�y6�
L�D��!�yB��#j)���O w��I�!��y�l�7���a突���Y����y�JL9L��\2�	�(H�B����y�i��g&���˨q�JԊ#�>�y���6�Ih ��*!�B��"F�"�y��Z�D_LYr�nѕw� ����y�\�{�xpX���$(��-B��y�/޾/�ơ����m�b�Ig
���yR�i�J  `H�b�J��	K+�yrP�US"�i�^\���w��y-ܪaY��� �)��,P�Z��y��ˤ4:�@�#.���2�ֲ��'J��?):�o���X �Ħf�j(@cJ'D��Д,�*���C��(YĎ�s��#D�H!�釯W>�ڵ�Е$�x���a#D����E\�4�0���B�Z��#�y�,�ak�셏~v@�J�T;�yRm1=߾蓤�nz�%j����yB� h��J�DS�m��q+�<�y�ň�RNFœt͏�3Q���DgY�y�o��.|C��
��L�)�%�ym_'�:Y�qӸ�8�)�� �y�f�
V���ڥ<�h�S��y�;p�`���E�5�xH0����y
� d$QƞP�j !!&̿E�ȉ�"O��S���O�bx[��C;	���p"O�q�R��oWj��ޜwP���|2�IN̓
��|��LD�'W�iP�eԤf섅ȓ�*Ly��8S���)�ͬ{XH�ȓ]��ᨔ� W���"�٨F�8@�ȓ
&z�y"*Շm�>�q%��� T����}�DJQnh��4��($�Ňȓ�༁"��ng���0�Če�f���/�2�IC�m���WƈD��	�'ў�|�e��'m�����m��}��d�Ḡf�<�č�� X� ���pl'��\�<9��	�N��A��$"�R@�CK�\�<)1O]�%Nv����$p�\|87l�U�<Y ��>B��9iB��K$�Ɖm�<1����h���
��)��_�<項X0#� Pr�6"�|����H�	j�S�O��=��cٵ_>>m�1�vY� �"OTQR�'��;���+2��YIn���"O<����=v�Z(!�Iƅ�!��	\�Re*Q�B�/��:)�@�!�dy�R��቞Z���Œh�O������m�z�A��bK�<�a&�#@=!򤄴��qr��
$f9���&��!��0yD�*�$1���!��P�FOj� ���0J"��⫝�F�!�$~3z��T2aPT��CK�%~!򄏤P ��7Iے$N�0j�KE�j�y�ት	����U��!Ԭ�SB�U�K��B�ɲ�R����ðq����FcU*k�zB�I90n�g䑭@CjM�e�T��^B䉁"?�������#x��b&��s��C�Ir�t�����?h���bZ++��C䉄}�i'B�$��!�S��B��&�jF��F��V+Сm�C�ɊX�N$�g��|X|�N�`�O�=�}�a
MO
�����ܘ|=|�i�e���ϓ!��!k�0rCVX`Ƙ���݄U�虥c2L�2�B��@���ȓ�|����Z23잁zw&I�f�����V812�ş�>���z0��2����U�|��&�U�V�tEBq&ݫ�Lц�&�ޙ0F�,.��d"1��'cBDP%���	z�S�'GdZ��40R����u�B#AԈ��yc�QkMX.m�ސbuB�`�詄ȓ�L*r�@1��(��	~U�H��- ���i�}lF�P��X�,��ȓLTm��)�,'p����[/g5r��ȓrn���E��I1��t�	���D��I<���f��Z|:� +<�V�&���	v�Sܧ 7�Qr�/4Vr��bN�.zB8��d�'9DQ�Y1� �kw�����YTC'D�|K��˜n/Ȭ���]�o����M%D� 8��(TŢ)���N23�؁��"D�D�S�&���[��N�K��2("D����n�g�H)�d�� �J�`�O=D�<��^w9�U�@  �.!я0D���n�$>A�m��펏G����+�����p�N\� �Db�n%�śq"O>�+Q��~hR�(S(����"O����"��@؄�tHG�y	N���"O�9#�⅃8��J�I"	�\M�"OH��h�>V>Ap��Ġ(��K�"O�A�s&3+�R��E��)B��"O� �,���S�Md,9#��A`�@�'J�����C����P�Cu㰝HD�?D��3��B
(Բ�ӗ� �'�����=D���Ċ"^�i�*[��L�f�<D���G'݊Y� �x)��a�F:D� K1�W,#��L9/\��R�6D�0�&��:fr�jU�e��Q�,4�O��C?���GKNg}< +u
>z JՖ'6ў�|�VK�t�H@e���&�+�#�q�<�!�H�	s,� ��u n��lk�<I�炒8�^E��GB�X�h���h�<3��f�-�%k�:w�x�PM�I�<#d^�=(�-!�A����@P�<�PA�">��i��	Z�9v�rx�P�'J�܊3(7 �
))��Lq$��	�'x��A���q& �V�ùN���'��ة�h�).V@�,.#<l�A�'}|����ڹ&͠m�5b���*���'K�%0�w&y:��4�ȓ)ބ�G&N�}���R��U�F܆ȓh)����ߦ\ �lG���K$�<�ȓy�lM��G��C���h�5�J-�'�a~r��9@h�e�R�'>��6�֘�y��H04�(gボa�@I� \�y�m��0���/L��i��y�+U{���W"�
G2��X�L��yBcB'ܬ	����34"�� ���y"dܽ0h1����/)�"�	�G=�y���"LyLmE@ͻm��D3�K��y"JQ'~��E�R�҅dD0���A�y2I��z�'���bu"����0�y���!=�B#�	]_(�#�^�y��X'.��MBW��h�������y���	��D9�'Ϩf��xER��y"C�R�D��7,��uz��pc����'az���U� Hx�+L�?u`�@���ybχ���k���G��]�.���6�S�O���-WyG�u tcѭm1���'v�@���J�@ �d�h�U��'N����R F�s ̏�=���y�'�bPJ3���C��0y��Q2�ةH�'(��R�k�*a�4��&�T,Y�����$0O�Y�!�ʓ �q�S�%�h���"OD�Iॊ�o�j|�5�Ơ!T��|��)��E6D11��52�e�vm��mr>C�2A���"� $F&M��d�B�	M��I'`�}�M�s*
�F�C�INX�qY���+_�Bɲ$��>y��B�IC� �i��o0�u�v�����+�d�O��?�'����7}��榋/ n�
����يBQ�a��愵e]v�K������'\ў�<�4�֡Kך�3�k&Z� ��k�<	�l�H��P��^���P���d�<YcDO'oC��H @C�:�= Di�`�<�ǨW�k��3�,�!/r�U!CK_�<Y�(K.ߢh����8@Y��Q^�<	��q�)�n@.k,̚&Ɂsh<��b�.sg�P�cLL?�lYA����?���?�L>1�����bC��V��@�T�q%�r�!���I���9�	�,Pu!���!�d?!d�!�.���5"���PU!�$�L�*})D����Y��$8!�$��q��u��������)��!��D�R)��[��P��8�נO�!�� ��BuC�&hֹ��I��pPҒ�'�!�$��:�PrFN� K�BQ�����0!��J�d#h�c�
�Vu<,�K�!�?S�LV��ZH��pcC�$w|��ȓr����+)��1:�D�
A���@�(�G���p�@5ie����܇�a��1:�ϝ-I:����̂'ˤ��ȓ_�*�m�-�`���=,A���	iy�|ʟqO��z���5A3+K70H0�`�}�<�e�/Z�əƊ� 2=�4�!e�t�<3���V�@�^& �)DIV�<	�AՏ\΢̨�H˗dD�Q�H�Y�<Q��E�^+n$����I�#J�q�<q3�I%(�K��n2�89QN�ph<F%��A��Bĕ24y������'7az¯�K��{K\9t�\�A�(=D�`@���;K�PXs��)9��8i8D�tQ%��E�^��'�9AeVI�SB5D��y�ޏ��1��=0ڱ�F�.D��C�a�5WӀE)��.]J`�P�(*D�� %H9K�ȓ�@� ����=D���q�� +>�%��-�(-pE�:D��zEK@�Z��Ԋ����9gTeb6�:D�89��*%��h���6��H��*D����L]�=�X��L�G��p� $(D��2Q%��v=�� ���) u��"v�&D�d��ĳWs�h�� �:= ԕz��$D��p�B�(R��C*�: ���: �!D�M@]vٻc�]	�܀ d!D�"�I	^���ICƟ2�T���"��?���	�N�!�5F�,7.� ��2~�!�D�I���rQÞ���<Ŝ=�!�d�	� q�e�C8;���;G㇈&y!�ǪQ����.�a���Bh�	!�d�+X�x|���O�ux�I"�� �W!��{��)xS��J����\�i�ȓL��ݰ�CJ�f��y�Ǡ�^�D���l>=@�G �E-Rو���M���� D��Pp�YS]��G�� j��|�j?D��e,��N�B����&�Nd�נ(D�̓TC_!"��y����R,����9D�|���sbh��m�V� �Z$o8D��(@�D�:�x�e�%��aH6D���v(�c*�=�tm�4�ݒ#��x�"<E��'���{��
�ٚ@ɝ�q�2"�'��Dc�k۶�'#��Y��l��'��	�Ũ!l����^�J6R���'�m��Ϥ
X>m�pK.APı�'�:Edaڔ)�δ,T佹����yR�ѓy
�Hf!J+^����w`E<�y��['����_:E�X1�5�?�K>����蟜�1g"�4"���"Ӧ�^d�w�0D�@�mX�/Ӽ�
')�(�l��׈.D�\�AB4:ON�
�`� Y2 +D��H��":�btس�ů�6q�g�4D�,d!�z�z�@��G�i�X����1D�l���L3K����d�"�*�3D��kbj�x���	��T?����2�Iş4��Ӝ$��	�Am�����K�h^$G
C�	 R(��[�Ȕ�B��BS�Z�L�C�	�h�*�tH�|���D`�"i�RB�	:?EI�-�GjԤӷ��E�B�	v3�HEi؊R
�arGAPFC䉹-���q�4z)�ⴭ��qW�C�)� ����G�
e�p9��D'������8�S��djV8!%`W�.�@���͇�/�!�Ď6ӠLk�̇�y�y
���,�!�^Y��Ȉ�7B�z��UG�=&!�@--J(�!A���Db��E=p�!�āXY��0�c��u�|[bݓ(�!��]�T�P�S� x̍�!�3>f!�D �����ĉT�d�ptJ񃉹@F!��6\	J��A׎e��ĐP#P�^�!�A�Cw���Ck<?�����BOD�!�$Wt��"�	ȸX����N
	�!�D�)XPt�f\�>����F)�Vr!��6u�<�Ӓ3�\�	��� :g!�/K5���n�<a�gû�!�ە694���d��Lc"< �d�?!�0[�4��r�R�P�~� C:G�!�DӐ*9�Q�0 �┰�=o�!��Y'hpt�@f��DP !�;'���d�<w�������=���`(��z=HC�I�0 D��a����MJ/��fC�	�@��r��><��q�R�0Y��C�I�R��K�M&$�`��.b��I�"O�-�A	Ћl�v�R�-Q !b(�d"O~�i"��A�H��΅L*@qI�"O�taC��s�̑s���:'� �S�'�R@˩,�i��� �~y�t ��!�DҨ^<��Rō&	̵!A)�0�!��yB)�k�&u��<1@f1P]!�$�a�d�c�GӰx�d(��]�9�!�DP������N,�ƍ3�,�4C�!���Bo&��Ǥ��s�T@#l�� !�ď�%2�(��Ϻ9�2�]����DH��4�f���)��9#�<�C䉆@�����-԰(<U�G-� n|C�ɯ
���Q̓�ĉ��LZ�6�zC䉜1E^�RÄ4��da�L�K�TC�	�:�|��D��J�����*�	9��B�I�E4R aڇNyv�� &�&k�C�!�,��f�]�J�txj$,6�(C�ɓ`�4IG���@���g���B�ɴ�v��&M#)f¬�C�^԰B�	���LA"(�)T�1�_)XӂB�	�q��e��$��p�ٞ���=�	�����ƣR��*)P7�D�4�m�ȓe0�2�DE�~����ȝ9NtU��Sm��7��/h�%�dK�6g:|,��dP���Տ]3%���1��S��\��E@Tu�8��;�ՉV����z����2fI#���(G�$4�����Ը8��,f��e�t�G;�J�Ɠ0䩵7��L�D�?MΕq�'��Xg����24B�0A:&��'��,����]x��	G�"����'Hx��Clc�b��*�\�3	�'�~X8�L�0z��1�R+&]J|��'�����N�P��4�բ:����'���a��Ѻe[@�G��/P�I���?!&�A $���̴f&&�bF��y��&�hh']
a�	r���y���-:���EM�R���������xrE�.(^�HQ�	ښx��ĉ�%G#b��Io���9F��!nv��G��T�t on�<���0�@$I��L
L���O�<���)�l�J�Z��"��՟�G{���1� H\鲅��>� �r�Ȣk���"O�����I&�$��c���Z�"Om��fV!&7�iA��J@rN�sO�xY�D�C�������
4?�j���O
B�	�#v&�E̓i/���DH���C�ɿ%���)�/jؘ]Q��T�v��C�� dj���ŢC�P�ybO��B�$m�6=�3`�!.v�@aV�irȄȓ6����S�zth�6<�9�ȓ�p`���ުDC�EP�%�1�5��Q�w	��&����1�![n#�P��AK��+ϐ
^���Ňу[uF��ȓh��)�GC�71�p+��݀r1�e��	z�'�d��a�_�*p�JR�}� ��'�D���p� ��l�rK�5	�'<t��ٗ��L��Ӆ6��L�'��=as`Z6#z�4�I&&����O氛2fA3*�f\ #�:���)�"O؀���`�p�#o�<9�"O��a$gͨ�ց�#V$=�@U�$�'���:�D@R�|Jt��%�([�4|O|b�,��IR	Wi~M�"���>h�� 4D�@��k�9�Q���]]�8�Q0k3D�D��E6�&�q  �C�6�+�o,�����Jd��I]>)
�� �$�Ի�"O�1��4 bu�� �|��H	"O�M[u�;�r�ه8�X=b"O��c̎&��3�
]>�r���"O����P#��v
�(-�D �"O�"e�x<ssdD!���I""Od���L)1d4�Ӏ�P�YQ.Y��I��@F�� �	'7<��aئm�6�Q3���y��
#/���أ�0zچ5@�I�yҦ�iM�8`�;t���AN]�y���N����C�%m��d1��Q7��'�az��,c�4m #W>X� �%�Ķ�yb`8f���KK}��(�UA���y!ؕ:eb�����u	&���y���X8��B��D&l����	�y�'�"O�h)����6G��IcC���yr%��/��}8V��%#80�ks�@�y���@�.��c����Q����D�O,��-LO ؑ�4K�B�I�ޛ*�PP"O�3 ���1 XA��!P(i
��p�"O,Pñn���A+q�T�@%�8�"Op�JՂU���b oM�1�Ĕ�"Ov���터z,,I�s/�6-�(H{e"ORB�KE)1^U����>P���"O|��#qn䑹���7�
��'"OR�@��Mж�P1��4F�H�a"O���"�PB;��Y�Y���"OF��M�f#@ ,�F��g"Oj5r�A�;.Ad/rQZ����'%!�d6`^��A_�wۨ	P3�@$+�!��'Fn��ĸt��"Q-�.S�!���\v���4�TA8��	�;!��(G��:G�|��LA��d�!���1��Uz�ë^|��8%���5!���+v�"�y��Y�w<����!��D;~���qB`B�S3qB�N��!��FR2|�F�G'ft%�Ҍ�9�!��RS�*qF�Xb*MDZ�!�C+�.8��`�. f�����!�d\8{KxHZ���
��I���s�!�� �1v㇞�x�ʴ�M�fH���"Ov��7�^\��<�h�8GJ�1kG"O=P,�/y�z$1�e^[������'����kC7^�T�&NȜ7�`����<щ���&������IRP�!v E�I��B䉭g՛���!0�;���m}�B�	*�����)O)~T�I�5NB��B�	�]�HP�Bf_yi����@���B�	k*BY�a��"I �%8R�"O�d�mթB��DaP��+i
�7O$M3�C�lp��BEZrX��2�$)�Sܧh�:E��q�8#l�zl�ȓ&浺㏘r��5HQ�ǝtzTtG{��O�h݃W��9B�	ڲ�ބbG�4j�'�P���U��J��2)Z�R`h�'�Ze��A̒|Y@�C��#	���'����?oV��"3Qb���'��E�r��yظ��u�ԑG T�K>����i:z��hZg��u��������_|!�đS�(�C�(#�t� ۿqU�IA��(�x�@��K�G�܄��jF�@���"O��$ڣ#�09*$�V$h�T�g"O�4��j�4,ČsaǱ-�>(9b"O��a앝s���*W	�m�mb�"Oxف�IȉT�u�@�Ї"v��RG"OPx5�[3(Vd�j&�W>J.p@"ORlB'���E"� q)?b:5��'��'�ɧ����R�eQCͨ$YB*G��P�.7D�4H���2�ʌ�Aߠo��`C��7D�P�W"%.H���=)~�!�L(D�l�`�!�$�!Th�)@p�� �:D������9$F��1)�	A��Xօ=��*�S�'P[BPz	_�u<N���f��LA9��~B��i���5:�^�SԈ�"hΔ��۟ ��y�)�=�x��'cASӤ��c�C.�Q	�'�0U�p��$��}@���%�J�'$֜��T�<�j"�B�.R�		�'@6� F�� ܐ�{�f�~uzA��'ڮTjEe�j��2v��{�]�'^���C.8���ɴ&�%��x��xR���_H-�c�ЙnP��T՘��d�O����O����O�[�Pa#�DM<MβU���!��P�0k��BF��)�� V�QP!���v%.�����/)78!�GX�pp��:A$���F�T�s�!�D�j�� QĆ	Ԣ�f>��{2�^��1 2�	�e&I��{��T�j,x��'[.�Hs� ��Oآ=��
ɻE&��<��dŁ�~��:�"OHh7(�*D��1���+���k"O��)F"Y�N^m�R'X� c�"O��bᙼ)�X5��?]�H��"OBA�rIIHu 1��n��&;D��ћ|��'�az򃒝(и���D_��� ����<����'jxr1 �Z⭚d�>�	�b�'�a�t����ЬݽE��A�W!�y�휆<�6�[���;6@��K�M�=�y���g�F`��>x*�m��c��y��@�R v��R���ZLdPe�+�y⯄2E뒅�GcR�U���B���$/��$O�1q��++d�ܚC��x��p1��'"�󐤋=(8E�
��=	��>�	�|��M�O!��j���K.`+�͑h v��
�'�R�(��<�vqz0AƺM�:dr��� l!�a�<a��4re�E�t�y�"OP��Q��:ʤ2F�����ӳ"O�!�U#T�2h�8�$N��>\���"OHxQG��\.����B� ���J��'m1O�k��	$C��qɶ"�lY��"O���R(�N��%*� �{l��"Oh�)��Ūq*$����>V{)�3"OX=C�����S���yc�� ""O�M{Bǚmz�dc	�Ue*%"O���C���H�8<���I-_'�)W"O�ًW��t��3b��(�i��X�����k��hȤə�b� u4I��'�@)!���6��ݙt� ���'� eKC�V&ǖ���΋�}���
���d�2#[z����M�L��5Y#++D� hG�>jV,b���0�� K��'D�8+��[�w/t�z$AIj: �	%�	X�'j�I�m��[��I�g��(&�
�>B�I*n��[��P8 *�y�JBE��C�	3"��$g��-st�B<i�C�	$K~<���ƌ.崕pE�މd�C��<@R飠�2	@�	�cH��>�dC䉢(2�F��7k�ӳ��}�jC� 	�J��@�Q"�
@ U�2U����d�O��mS�T�f��C��ag޻"v�C䉉6��J����o�a�!��ӒB��, &�rc�� '�]����2	0@B�w�DqA*������2"$B��	�(Q�v!�@�¼���P;��C�	7�>e���_+��Z�%����C�9pB�[���/���A$��"���d�O��$�&�N�r�ǜjFB��r,��f2��D$��S�m�<�Ȍ9��\��  :D�<Pe�1,�b��N��h��C8D�
/�>U*СZ�`G6��'5D��`QK��"M:D!Ǩ^�FҰ� 3�4D�����9�$\�����?��m�'�0D�( ��P!�F�acA����j�b-4�2Dn�R���N���<#���ן<���4+68��Z.6��+�*��z�p�����)X�~U&)ɋJ�P ��<D��P�l����p�G	x�L�!/D�0�7������JY�`UM@C�?D� rQlx'���"���x��)D��*e�M>�R@qD(U+9@�;A'�<����/u�vT���y��d
��ݠ��ȓ!�\���lB�c�H�`���)���IaTU�,ۘr�6	�2�$;����d^��/Q<~�f)r5C(��ȓl��t�EG 'pxy:�BͲj����ȓWdi���,����Ĕ9Q�݆ȓh���P#_d:�aen�7DyF��'^ў�Dx"D9-�B�H�J�
�1R֧Y2�yB�.�0YqB@T�v#M�yM��*�P%C0�C�8l,�QC �,�y�������0�����-�y�Q2�����)�hx!��4�y���7FU|YHu���*$ I�7I��y2# )�ܩj��6dw��8�?	���?J>���$9��XB`ϒ�0���Y	�'�x��Ō9v� Pq�M|�l��	�'l���Ҏ�]�Ɲ�EY�pk��'�n0��g��+i��ar�Bb�pв�'��	��`�%Ad�9j���S\H�@��� ��;��[�<��Y�O]96��4pW"O"5�r�M�[X��nC&m_�` �"Od詠R�+�x\P$�=vl�ը�"On�TD@��FC�*;^`�d"O�ұ
�8���h�,^����"O���`��u�u&�N �Au"OQ���$��ô
Q�J.�y�
��:�����!Gf"���
��yBJ�HM�%���j����V����y��	q����b̓e��œ5��yRK��]�yz1*�p�r��H�7�y�Nޢ.��-c��Y5mp���D+�y� �;��q���Ӧ8m���� \��y���Nah�;@dK�|,e��i͈�y�`�/T��؄K,��y$l��y�F��S� �Cd���
B�Ac�M�yR��E��@	cX�1[�	�C̈́�yro̔�2<��n�%r�(��Q��y"l�0w���`.,n�������y2鏦H�6U[Vi=a4���KS��yb�9�T�إ�X]�A�����y�"S� `��;��G���-5Z܅ȓ=\�X
��L�m<Z��Ú+�贅��L0EN��	��c>5J^|��Bs���L4������2iLq�ȓCo��C/�e^!3Ш�F"�ȓ`�"u�Gk�)<&^M+���H��<�`�acF�.hk�;�� �Tj�P�ȓ9葐�  nK�@X��C<����IJ�`>����JĶMsV5P�,֜KɌ<�?�ӓ�b��G��7�q�eM�3���� ���i�K!��24�X�����N��q�х�� \�p�n��9�X���,(��S?f;�أ�&b�x��f��H�3NB�}�:p��fU�x�Xu�ȓM�~���W�r�r}���S!GʼX����${�QW(�Q�Kl�><��P���O�0O�ejUL��$Ėa��g̾)a<8��"O$ �Ҍ:�*�7��#uT�Q�"Oph�E(Z�W�4Lc��6+7� �"O*�@�h��� �&J>�B�"O��a2���+fb} �G�B<��"O��P/�}LrHA��m�]��"O�B�ݞ�0�Ā�*H�lm���'r��'x�dI�vD�A�iɿ}�|�����'�a| ��08$GBA�4�H�vaɡ�y����$-J8@�M@�5h� ՠ(�y�ڳr�h(��"������y��W��}H̓2V�)�iÅ�y�H �pt�**TtJa�W*�y�A�vn�A�C��P������y���:�$�C���I�$��y���h�|*�gO$&�U�dn�#�y�n�	A�pP1fK�� �l\�yB��
q;:zq�$
����FL��y�M���(+e�T({���Z6�D��y4�.�3W/U�y���[6�ߕ�yr���u�eb�Sl~�hxEN�.�y�i��QD��S��*`L(�z��y�KT���c"@ X����j݀�y�Ҏ}��M�sDHKPN�r ���yB��.��@k$"�/��b�թ�y�E16A�2�X�V�&���8�y�n �%t&4 �hY-M���E�B-�y
� ��#� �%�n��c��pŐ�y�"O���2i��C��kdH;5^d�qA"OZ�����2'�=���OEQ����"OP���獧t�PpA�&ǰH�ak�"OV�qĂ�-���x��
�p��B "O2tX��N�%@��3�M51n� 3�"O Ee�FHx����̀y�@4*�"Ov�� �Y�|�*J�#Y�k�ք��"O��CP�
1��<��L]�]��� B"O�5`��;b�&d��
����IR"OL��V�ٸj���S�2O.�A�"OB����:J.@�����2:.|j�"Ot��R�ƒ�J�SLc�a"O3p��g�I�3���(�
5"O"�X��SR���A�U�|��e�B"O���C�Jă��	3V����"O�m�6��|u�7A�&�a"O�q��:	�D����l p2"OB9��,^�Y�t(��/�i� �F"O��Bv`^�X6(���E�d�"O|�4���MlJ�[e�^� �P�"O�rI,6��u�#�`�ш�"O����L�J����`�R�|YV��"O�Lr�Ɗ�?�}��@�Y2
)�1"O�� ��p ��D	/>#v��"O<�{�@ �	��R��Ű	
<��R"Ov��ʃ#�Ι62����`"O��:Q�G� �L�f,0z�U�U"O8Hj�'�/z"�Jk�xy�T�3"O:5��R4�lzD8f1��"O��p�3r�H\��A@�eM��!"O�8��JS����	W*�'�&�2 "O���	��S�(j֩��\��]�"O��[7�	Q�1gnH'p꾔�"O�)�Њ֮�{��C�@ڶ,��"Ob@f�Ȅ@nҜ���!<�-�5"O��:����U��$aRU"O�@���6��ekփ�����jB"O����#˷	,��	����P�b���"O���&l�ߺy�eC5}4ZX�%"O�,
ã��#ⴱ�����<�Y��"Ob��/��b�0��#W��d-�s"O]2F��![��	�e��o�cE"Od�� K�=
�d���K��Vp��"O�MB�ɖje���ͺT���X@"Op��-B�y���ƤI^�u8c"O���5��to,��A�T�8Ke+�"O�]�S� Qt����#�����C"OJ`@�g%��DzA� ���i7"O�TɃ+H%��۷�f�l	��"O�h��L�q)ċگ����B"O�����ѢZ�P,�fMM�8��L(W"O��!�w��h���P�d�L�"O��C��ڴpQ"# �;�($�"O2� �B;hd�DHB����"O��ҐG	���ƣ
1	5d�PA"O@0DK}�ՉrcR;���
a"Ot�هb�o��Ac4���9"O&���Z	V����1☛	����a"O
�X@�s�8�W'�	�r}2�"O�Đ��T PQ�M�p��Tn<qs"O|R2�J�@3���oKtY���P"O���MȩU�҄��\����0"OJ�	q G`�b9�������3"O� TX�pg��I$<spl�5|�(Pxw"O(���T6a��Y�@��� ��c%"O*\�%j>,Hy�Q�K(�����"OH�s��ȐQ�i fI�$��`d"OD��ҨǳfP�H5d�5K�� �"O
�a�Q�����;x����"OF,XQ�&@J�`��_�WPb��&"OFkU,$,�}zd��,1�Ա"O~�@�&�$Q�R�!r�ڽ@!P�30"Oȹ��I�;F�aSCC�.��"O �!5T2qe�p@��l�R�`�"O�����E�j��- 0���H�9"O@��+1����a��)�(p"O�!�F
������֫P3�"O�P
�B�nUDA��`��/(�*�"O:�r��̧l��*�,߱)7��U"O��1w��2<ܘ�CԦB�t���"O.i�#E�[���8��Ȭ{��ak�"O����A��H��0�������1"O:)"�.��1ka\�|�șQ"O~drr	�6�*�a6�	xL*��"O�@"u�;>
�M��]9#V)�f"O(qwJGC�(��-���
a"O$ ��+�-� %V�O�T��"O\h�O,])�ҤӘ�%{ "O`a��46
0X�%��0�����"OF��D$���P#ĺ �JpBP"O�Qu��15M�9VG�6�4%:�"O|�3l�8`tP�#���	|��H؇"O�ia��ڥl�PY�^4���"O�\� ��e������kϐQ"O�t���*u�d�T#!f�q�"O����O�0�0z�!�z����"Ov5�vϭ0��aq��&E��4q�"O\��Q�  N�Q��P#E��P�C"O�*���TX�iïP��Ũ�"Oze2$��;#��run�~�p�7"O������*�;'��bf�h;@"O �r1C�,y���X!�֘c6e��*O�Myvj�n4�zb�ǧ#ޜ��'X�"Si�5�V�;C���M
�'6�ؑR'цh�Er�	XN���
�'~l��%L��jMT��1�P>L�V�9�'��i5�V�L/�@���@�~1��'-*XCP"(Rl��" ��@���'T�P7�
�uD��R���93��a��'��Q��B�q~��dǏ�2��@��'K�h�sϐ�%i�)j�U�,���"�'�� �,țT�H�iTKR�5 ���' ��Ĩ�6f|r �6
"a��<��'��(�Ѡ�T���za/]N��� 
�'#�k�iL*2�@��hH	BU^��'��zvk#~�z��"�ɚ,�A��fź0����vJ��+�=&�N���e�.D�

*y�ѣ:BV&�ȓM�NT�����Z�
8We��ȓb}h�C��!(�>mj���[� m��Xt�E@��/A8��,�3	V5�ȓD�r=�
��(�p�Ï�W�h��ݸM�/�1���E�L�KM֍�ȓ4i��@�7/!�q[g��)(�:���D�`�I�
�fM�(�j<~Jz5�ȓLYԩ3dʣ^��!�)B�+.хȓ#g����;���R�X3p�Zy��S�? Q��u'Ԁ@r�Q�8�\E�q"O� `F��
{}"]:�ژ�����"O m��,��d��� ��+B�k�"OT��n�' �Uڢ�7D�)C"O����]9-@��N\�C%�"OpȫCo�/?�i��_�7��"O�ma����F���q���)수�"O,U	6$F!8In�:��֟UuBȕ"O���6�Y44�\0��7(mĥ	W"OH!��_s�:a�@5lk�ݢ�"OJ����>j��+ں>{�l�$"O����'�tDPU���(�З"O��is��7
n�|"�עu�t��q"Oڰ6a�1o�QP��ϵ<���S$[��D{��IU|�*i���n���J1��$c����W�#�pa:���?<t��	�y���c��ÇC�3I���ծ�y�1.\ع��;i��H�cm�:x��C�I	.�| ���V��
������d)���-q.��f/D�9��ِ��sFB�I2ly@�nH�p�bQ��Zc�B�84.�����Y73�rd��W%~�B�	�4��G�4V ZX2�o��:C�%��7(�	:o>�@e�$��C�ɮ@��`HR79� ���U42�HB�q[��Cp�Em&�9��X��B�I.h��Q s�������B�I"\, (�h4�=01�F�h��B�I�r�i����`�t ��e�V`|6M)�0!K9v$����C��5-��$�%D�D�F��>"v�@#�F��	���>D��A9g�z抁
2׮�(�B*D�s�S7"D~���@y�����&D�8�OE�R����
lq3�$D��2���"�В&֋I�<�!�<�G��>a�(M5�0�۵Ԧ3���@��4D��(�-�LZ�uEL�O�2���o�<��g?�S�Om�Ě�� �0i�ի�HݐP���y2��K��{�('$Od��S�
��O �=�Oj$����[��5b֦�(� R���/��>�k1� #������0�Jb���c�����D�#�t�XÉ8]����Va�'9���˦�Fx��)��`�V���΅-�L(h��ș`�!�ā�H�bШE�ك'���jqň��V��'��gܓZ���K&�]84�E�a%��^8��	�<���B�:���������0��Ay�>i��hO�T`ShXh��Z� a򤨡�A��O��@p�j�OZ�8!��'#���7G8T&��'�L8��N�M�6�T�W�E �'N������qO�a���� �@�ʻL&��"O�,ʥ�X�du��y$����0��x"�iPa{r�]� F��(��~.墠aο�y���r���;�`�3JPH�����>��Op#~B�b�7[�~ȉv�!$���(���V��hO��ŦAE��hʲ�b!O���#�<Ʌ�)�'m�Jtk�&��v88����'*��ȓI��-�s*x{�>X�7���6$�&�$��(/���a�F�x��&��)2C�I��|�0A1^zQ@�ی'G�C�I�!�r�#���ڠ�a�֥}��B�G���*�چ�fQ���g��C��,)�)D�;�<=�W�[8�C�	gBu�$.  6�01X �ܪ!�h��p?�fㅫ��3�KȚ��D;fJ�eX�`�O� LՊ����ɁD��3�h�"O|HQ�O�SF�� MT�G�m+�"O�`��q��i5A������T�HFxb�5~yL�ڠ�W�� h��J=�2Q�ȓ1~�T9RbѲ`�0����g ���ȓl��z`��)�Б�k�-OG��	p�'�"<I�4��(���$�A8��_�r�i�ȓ	1�����+6�B�s���D�'ў"|Z��"qT��g� ��a�#��E�<AV�ǖ+?�Ѵ&M�F��P�dA���xB��b�*� /�,��swρ�hO���I���h���ψ%Kz)����'ݰB㉋i��[E�	��ѡ��ѣo����hOv�<q�+ Y64�Q�cS=2F��Q�a�TX���O4�{�A��d@���V�C��@VS�HmZd8����}�vZ�e����rk&D�8�WA��X�ٓ�-�>:�]n#D��	�.(�2�h⃕Q4��ƫ.�O��5�CBI�^� �Xa, ��m�f�	Z������=����/�haH�(�O��'n�S�3����2ڬ���A1��%^!��МQ�N�B4TF*�B`Í�+S!�DD?؂H9�bT�� HX+m!��]�3eHA7�I�cD`,�%$ہUN!�D Nx;"c�)?��s��E�HC!�$��
2��
s%��o��(2g����!�$��8[��P��w��xp! �C�!�Ă.>2Ŋ�2JX"�j@e!�Ę�I����+�
QJՙw��1da|r�|���`�XRe�� �{��6�y�!��'��T�3�դDn:@��&Z��O"�=�O1<����#TuZt1mM�c�����'�D��0*�f+RY���]���
�'�RTj��R�"�H2Fw����'lA���<s���� �n#���'$��I6��U����a�!^/��J�'<t������h�@G�Qp���'��d��1����#�	�$�/O���N��P\���Q��u���� 	��}�4�pg�5 ��1�/�/:��B��<D��ᣔ8B��ȥhN���9D�8�/ղ	��}ؖ-W4��y��&9�lZ�#}p4�f%��{p��%/ݳR�8C�	?=y��aM�f?<�� A�'Fv���/ғC
1ԭ��J�`q�L�?xv͆ȓ�n] Ԭ�,A�Hl���V�x�'���2�)ҧlmfa��C5N��M��*�X܆ȓb�7�
�[�!�H�0�vYiN<��v=Z�C9H4��qF�rL�=�ȓ� ���F���ܐ�f�A9H|�H����
�V"/Н2q�U�͇�	{�'ϴ�07`�^�!d���dĀ�'�L�R�_ZF:�i�����N��'��C�ER�T9�!,�u�t��',0@�����B���`!�R���y"�)�H4f��$eJW%�t�z�&�� z�'��uY��*�,��ˠeY�D��'���s#�T7b[��A4'��K	8y�	�'n����`�bC���B�<a	�'/��0L��|�{���,=�$�(�'�I���׼V����I�<��$��'t�# LS> ��(i�$@��� �'E��hO�O;���� � \�AP�5��3	㓴����B��8\� Q�r����S�? fX�C!G8^��yhVA��s�"O&���Y(؆�kaȵ"2�a;V"On�@�
�9�xЛ��1#,z#�"OXl����)mJ,zC�1�]�g"O(��桗j�� ITA#m��S�"O�i�,L�H=�' ����qT*O�`s
"%�P�B�n
�(9�'��Ik�)�<Y�\P|`�ʊ9(ҊmC�H�q�<���4L\��aS�[�ut蠴�i
�'{ܼpl��<'�S��ެ\�t�ӟ'�ў擜ٸ'�fd�'E�GLάa%'��.��L��"O�ɫ�C�4m�Q�F�#�9[54O�<)�����"�/j�,��㏏Ad����"O��맫�26Y����6U�K�"O~L����5[6�Z��
n(�� "Oz9B�"0�qI���9_��`d�-|On���шfmЈXj�eL���"O�m���ʩy�8(*1薡��q�A"O��G��l��K���0��l�"O���� �b���E�X|hD"O�@`��ɍ��9�P�K�b��"O��h���4+�A�Z�P&z$$"O��I�	� ��08B�ڠ"O�eR�K"ª���R3m��"O$a�ѭ�2l^��Bhp �"O���1a ,vǼ�5��5�4��`"O0۠�B�� w��7{Mj�"O(�1�N\,�� Jw��6	U���"O�PZ�Qxd�=�C��(��C"O���!N�<ޥ8�"�m�W"O�|;E�L�M�|�I���K��¤"O���nX�j��xpgiΌ*�V|�"O�TXF��3XNb���K=��Ӄ"OJ<� �� H�A�v�ϝy� �#6"O���mP�*)
����і8�"O�5��J��u:���:kĔ�K@"O�-�p#X�M�p]3�EE�'���K"OX�S�l�?�9�#���?`��"O|�Ɖ��A�6�?B	$]j�"O����.[�����=D&�<�P"O�t��K��xE�5�����"O�]y)��J`��x�����"O�@� �I������/�8d!C"Ol�1)D*07d!�1E���a�"O�(A돱R'�<{�����!�Q"O�ͪ��P�&���I6� ��D"OJ�peʃz1Z|��I��O��1�"O���p�<"���a	ޒD�A�`"O�9X1��=c.�}�a�	5lQ��c2"OPP�^�Hzè��d�k�ᔃB����1a#0���0�'�*`˳�C�}#p1B�G�	�!2�'�Zu��/mwDHkTjN�x͠I��'˜`ǡ7�Bmԫ�}�`݋�'���`��V�"�$u��K�8M�D��'mZ` �D�.�f ��&�><���'�����ȋL���9��!bo���'{ �x-�H�,��pH>nD0L8�'�N�W̉�j�b���gY=[���'�􉡀F`:�(�&�]z ���';b��T��F�P �pn���'eZ5ϖP�����-[�o�� �	�'/�L�7��Hhh}a�A�o�� 	�'v��em�;@`����]3f��e��'�I#A���*��q�� f�T2��� �г�+�17��A������"O��iЌ�~��f˅�j(a0�"O�]@b�Z��$�!)�>�%�f"O�����1�N�SΞ�$���B"O�|+��I�]���7"�^˼�!2"O|1��b�3c��\����\��"O���eW�
j�+'�ܕ`�8��"O���-�#���9��=��tZ"O�X�cĞ	R�w�N���9'"O$ �ꃍ^��@O�9L��Q�"O���Gj��E�N@ӲO��a"x�ӣ"O���R�B�i��O	� ��s�"O�ՠ����g�����*J6��"O�T�"
�*s�]���#��1[�"O�����R�48�Т�i\�;��j`"O�9:R.�@?�
�ݍHV�E"OЌ�L�}"@0��l�x���"O��c�.�n�4{�,��R0d"O�9�N
H��ҡI�B��h"Or-�W���*jꔂ��<PM��"OH@8�J��<�2��`��)4�� "O�䠳DիQ��-(#�6z/R���"Oh��.t��wM���0��"Oj)
�e�7e_`��E�1�ܥ��"O��S5爃ij�<ۆ�&(�n(��"O:�0�/ؚ9����,�54�ݹC"O(|r���)+�T�s��V�/y��R�B�V�������,�����C��u�Z-z��4Z(�􄔻R�)�N�T��NL�T��x!�4olB�0��"D��B�!�Oe,M�G�ǀQS
�r�>�	 RY�J5��D���Z���.!�@� ��S�!��pw�@���$Ͱe�R���JH��*�{�������ɶŰ� �̏)4�H�H�_�eTLB�I0AEL�;v���L�`dJ&Z�a��	+��=`$�~/R31)��jS���-RU�Ü�0=i�I|��'���S+T(i��107 ��p��'_f��([~�q&S6m;�p�{�I�7g]�O�Oj��9�MW=F�̢0 
�fB�TR�'g�LcM�2:-� ��Ver��'�4c0��,���',��@z�$�'D�M1��k�B�� Cdz��
�'nt){���!w<�h[�"^���'�����CFB����%��0��'���@֩�"���i`I�L��q�'��a��nQ_ۖڒ�� tp� ��'�d�㦙\%xUё)�
?V"���?W ��f�m�H��nQ��08�6�Z�h
Y;�"O�Hp�	R)l�\�3���/�(Oȩ�F'BO�Ni+���\7H����7@�\��u-�QP!�������[l��a�,��!R��!+�s���H\v?����OL�k���j��@
���`���"O(Ex�I�("Xq!�&V�l�װi.6�{Q�D�)+���
ޖ,��xR��)��0�"��8\C� ��ē_p:� �(!��*�9r`g�	$X94�iI�㍔	C���A-L�b�����Zx��pC��W�K��+S.��V#�\8"o;�	�\&�Ǎ0J��h2�q~�&>IA6��oB�B��:f&I+�!8D�L�/D�
:�S�-�H��w��5b�R�� �8A�ެ0$Q�x�ң|��O�l˵���v�&(p�ōbu���"O����Cy+Fx3 � mkX���?9m�'"E�YT-�ƦQ"���G~��Z��[�,

�F�*G,��0=Y&A�G+X�{��=/��Zq�Q,R2��
���"t+�
� ���'~�1R�8�@iP7�ϕ(�J$Ç�"�X�!~�PI�b9Ӕ,�dB�	U�:�3�ן��ݲ_d���d��1�u�)	��C�	�����Ғiɀ9�$��мy�@�8�&Y28E�P(��m�����;IO�!�'��� xI!pˀm��)�X'�0i�'�}�t��,I^͓AN��DՆx_&��V�� zj"�$�?bI@A�'�S�m<-��� ��O��@u�ԇ~'�)�/Z"?q����d��;R������y�H |����~�x�z����	[����q�p�D$�sG±P@�'HԼ�d�8X8H�Q��X�D4e�#��8@(���'��b�8B�D��[>B�A��ؠF0qțw���FF֮F��T�I��]e����M�p�:�E��hk� [4S��ij�#Q>S-��BNY�
�y+%�''0���[.$㒅A���5V��Y:���~�'��Xr��?�T��L�Pa�xY�j��-n�ѡ��"y���/�=���ْ�J�B	�T�?s���Ң�Ӽss.���eԠ���.��]R�]���$W����7m�6i��D�p�½�' V�6i붊�)L\ @m]	zr}��r���ӗ)K\0��܊|nI����o��E��F��v�r뒟SRn�ď���Px"��}`���R��Qc���r���G!$e��9U7!��$1w@�}X� �[P��yBIL��5V�_?��Ca��wކ�a`/H�	V�����<�5ɑ!�jȑ�HƝ(�>�!Pk��b$�F>�v́"��xi!k�(gܙ�*�4�p���'�00�qB�6N�^��SCؔ�. {�}E��Āؓ����n� ��`Q*���	<
 xt� >}\��X�Ƽg�.�z�+Ƶ:�����$Sh�k��2LO<̉�-L
���cFˀ�f�U"C#C��ڌ�,|��b �ءC�����B�5%~�'/��?D��rk��8��4��֤ ���j�� \+!��,��<y��Be�^��bEۿzl^ɒA�NPb*� 6�+-S����u��#��|���S�T_��  �I���>��G-گGz؆�>�YÅ Z@8���V�št��-- ���g%��Io�x�9O����ɪ|^���Ói�怠B	:,��E-�>"����?�g���r�	A��uZb�O��ب���	!O4X���]a�r0���[�bT�� ��E<1c�J���(�
;cR�k3��3�$���+�i�EIÖA!&��X,��1�B���3T슲b�A�B�Ɍ.~�0Ꚉs��c����k z�1t�;�)�'7p�L
$�Y�B�رB/��:�ȓh���bPo�<�* �����)�HC�IsPP �5yHtԐ����PC�I/ �K � x�ԗ]m.C䉕F����F%S0,��j�ү]8C�I	Z"�����߂$�,|���Q8y�B�	�'6�eX�/�c�8dQ'�-o��P(�év]���>� ��⧛T�<a�f�o�2�S����m�9ÊSm�<��n-L�� Dg��/�@�tk�d�<�x�<8��W�	� o`�<�Wh� �p$�Ɋ.���pUhb�<���#�L��a�Y���sQlW�<� ��1�]��LH�h��9�d��E�<�B%�yD���aBub��U|�<��DM(E#~��I�J�!rmI{�<���@��$��L!o���is�<�ʏ=~���
�L�0URb�i�<єd�oq8���Њ�52La�<� (O�J��q�O u�\���� b�<A����� �ۧ?T���v�������E�I-G���"�*��q33N�;:?�C�I�ʒ�z A�c�q�D��	+Bjc�x�4�)@qO1�ȼ�"�@0x���="�|� ��'T��Q'�w̓x�H`iC+��k9�9�Ǣg���I����YR��|�  I��t[1�� 4����5��D��mjŋ1 :��	��T���3J �3��K6%b��"O��.gH%��[0��#���dc�ԋ����y3��>Y��V(Zy���^}.�猌>0�~��'�*}�F
*��)��L����	��'["e��eB��<�`�%ĥ<?D\:h�O_2��qJ�
F[JD�SE�W�����OQ>;��Ď���
1�_'E_ʡ��(�><�;�E�}���i�Q`��|9J���ɐ�?��K�F��Ӡ>un�7�"��$X�VDԉ��.�<%o�:d�%>�:n���aP�����S�'��B(�j�C٢B^͈�&M�8�`�ě�?��y��)N�)`y�DeC�鴵m�4a�a#��#)��DP�'7��!2���Q��'l2���cO�yʨ��i�1Sp@��'�:ѐa��_���l	?
�ց�G5-� �%-�C������\+u�Y�O�-���S:��k��,����΀('쀷2>��E���\$\X��]1���(���0�� z��$��if��VA�:)�\=�b�G[��wTj�Bpe(��dM�T�������`� �eK<17�I`�di��J�{gj�����#04c>���J�1&H� ����51(�05��H�(K��K��L�%BD7�ʁ��#�XC�UZ'@t{��*����`"]�3F�Sr�DA����#��I��F�<H>���
1c��r"�t31�B/�Q�Z�>6�J���5$��
�r���ӓm�Ɉ`�YS4�59���Z�)��ɕfh@�Ч$�cR��(�7�d�4��y��]k�gB�p�ș�J+D�|#�a�@q�ш� [OPy3�/�$�C����"F&��)A:D�p�賎�qKd	j��++S!�d_�/"%`G*�y���K��ߺt���=��/�:����Ib|9g�R��4�1g$�;�C��$q^���B�){��[�)�=Q8�C�ɖ<�9j�K�2V�X0��G<y�>B�	�!H%p�+����q�sDH�X�B�ɱ&�D��h�h� -��G�XC䉑v^5�FbW,N���� Ӧ@�
C��6&�x�:#n����4�δ"D�B�"�>0k!�.��HP����B�I* ��yK��(A���Wčw6hB�ɽV9��v �h��oK8.B�I�	�<Ȕ�m�|H���>�:B�I�]u�]a� )s8�rEID*�2B�I E���+@�6���c���h/ZB�I\6=����.d�
2(]>I�B�	/h̸gd�!@"����"��C�	�V%����)C�>�m�DZ1C�ɷV�RƧ�=A�xMK7f��T��B䉷b�J����5LJn�xg�$��B�I4�,����N�~WhSG�hC�ɓ"W��X瀂�>�Y"�MsIC�"O��u� �	<��1��_�!����"O��qg���l�ށ�v�H��a�@"O\���@H�e5LHg�XI!"O؀��gX?@��x�@䀱\�R�1#"O� (���p&���柃<���"c"O�Q�4NV�U3p��&h�.�pp"O��p)��}_���% H�i�>-u"O.Ec�
҈0�lA�d�X7.�1�v"O�5`��4HK� ���TF��Q"O��2w���E��P� ���'
����"O�x)�o��<���(K�P���"O>�K�ATT�yXu!�������"O�(aw�H �-!���EӪX�p"O�1�B���I0���0����V"O�ĉ�E�.^�>4�r'šz�I��"O�	+Qb�8*�vA0�H�/Vlz��"O0E �@@�Ga:|��_)3T=d"O~:����X�b40�Fݾ���"OLԹ+m{E���eEؘ},L(F"O�H�gF5A'�y!�O�#��%�0"O6�+��L/6*�����ճe���ȧ"O�ШE���t�\�7#A�r�Z�7"OM�FM�,M��}�򍐙%f��:�"O�2��x ��lE q�d��""OpR�@Z�>�8
�IW
�H�"O&����
��"I���R�	����"O^ܸk/fnU�� <��xU"O��QJ8D�uSEF�>b��T2�"OAS�H�`����� N�g�ZqP�"OLM�$��Ճ�o�,g�X}�"O�qg�	Dp�������)ǔ���"Ox �ƉH�Kθ���;I�����"OΠH�MA�}^�U͇@j< "O� X�+F�;ZP��7LBoFh+V"O.ܨ��V`���c��>����u"ObU)�=Y���,ģ>�ҝr�"O�tr�nA,J�،Q��`�~`�U"O�P;v�͚̄���DEΌ�xs"O��!��	:A�h�B�J_���+"O�S�b�.����vd�zzY��"O2}p�F��CX��"��(
b�C"O�ْ �E�_���Z���$)EL*�"O�ʅ'�"��!�ī\m
q��"O.�q��a�f(�S�ѩdoV�U"O��s)޳S��SjQ�P�0�"OTu��b��%� �㈀4Q<ȩ�%"O:ȱ��>n5r塚�b$�D"O^h�S0n)h`��M5���!"O�ĩw��f>�%'B?��q�"OL(����,^d�K�珗(�"O|��ԤԆt�z�@7� ����"O���b�Q��8�蕃P�Rh�<�y�K�������	��"Q���y��Um�PM��F��H��g��8�yrLQ`�lTF�@�{�(�c�ڴ�y�l��%JUI���|��8�s����y��J�5r3fM�w'���kڷ�y�넨V�B<� "z i�	�yB��bS=�u ֟k�2�څ���y��#}*x�a��1`�L����6�y�ȨO��i�1�B�;z�[̆��y"�Hy#g�=�2�C���y��;`d����B�֑۱��y��U�><���E���Ȱ���y2��/�|L�W ƇF��<x ����y��قP�
���ʃ%������y����X˲iW3�\���ߪ�yG��5�Աq���>L6t���ŕ�y��ʯ��d�B�E�	C��Ò���yR��\��x�iH/�J�A
�y�	��pqд�,β{�Z�2��/�y�One������"�L�t
��y�N��V�V���$�2iJ�����K
�y""�^�D��1�� �SL��y2$�=*�P|q���9��p�����y���f�6D*���]��tC��yb�	 t��Af��rp����y�̓91�(�s��v��H��\��y���$����F*e{F!q���%�y����!��އ$��irȇ��y���]V�\���Մh����O��yL�u������2{d������yr��h��u��ER?����+�y"K%TG
�k� �&R�B����S�y�F�y_
�p�n�M�.-��m4�y���V�`�{��LˠXX'�y���:(xY��ԃs@ � @��yB�D�Z��M�'�y���҄�y�'˚(��"t�I ,�6�sG���y2�  7�|`��1j����DĂ��y()���sPe�:��xb5��	�y�� `�����ϲ�Ќ9��N�y� DІ|�7.�>@����G�yb�94K�Z'�h� 0�L/�y҈���D$�D��j�P0�+�4�y��~�!"E�d��9pGh��y�G0��P��^��ۣ�D��y
� �����VlXy��O�	#o���"Od�Ѵ��I������zY��`q�L��L�=����O�1pӋ�`f. 2�L��T�!0"O��8�`@�Pl �D�Eg�p3Ѹi�@���!��|��݋~�T��� �ky`��H7�p=)�Iڟ@�9��e���BxCz�B�A��f �@��>D���vk�Q��u[3���t�0�ɍŜL�Ԉ��Y!?q3�i�&	5Re��N#��)7� D��K7"0^q�HwD�c5`(!�߹r/:)�EG���!���q��'	Xh9���w�	�@O	�/���Y
�zH,u%o�.�b GEF�T�P�� 7z\���٤u^81T�A�4	��I��j0�F';J:�3���[����7��;v#��pR�NMq�h �B3|�|�[Wb��ph�B5n��3���I3�YS�O&l�!h��KI��ۂ.�l�֍(7�B������پ)��X��k\
w�6t���:IL���*���λ|�~(�r�
rP0=�d���Vi��MF�\�f��)#A?67�D�D�@`��ʑAP0d��C�ź�3�P�t�~x(��L��ɗ(d��qnRk��Q"է��H����DV�I��$�U8-Vܨ@�Q�.T�|I1o�8}G�xc��ӿxY�取񾑓��5"^0��ቀIAt� �!Y :�Ƒ���[�>�nc������,\2�abL�b�#��>n�肅�S�z���E1O�l ��Ι�or��B�M���xҪ�>�}
�K �~ݬ�� ���J�~�S&r��w��*�����ꖃ=�Ajw�@���������" �"ɚ0N7eѼ��rb
n�<a������#Ɯ�!�\,����67
�`��Y>f��Z��3l/y����R���p���B����k��w��� ��ֺ�X}a�2lO<�r���*,J�U��(�5V�����S<ja`3�ҩI�T8��E��y�#�2I<��t�c�1UjԴ8�,�i'�DJ,xc�.�	�k�!"ꔨip�Q���IrCHΑP�H��� G7��q�jű*��0�Q.pB�	�\-<��d(U�<��栈������/J�qO�']����>���:b!��&�6ܰT�M�$���j`"O.D+��Φ8��иC�_Z �P�P��c��!LqOQ>�)A��!��勊 ���)�O1D�y�F��]w<�hԻ�^щЫ1D��ѯV�9r��S5�٥n�
iuJ/D��Z�%�ҡ(1�P�),��0J1D��h�`��4�v`��ѽT$��p�,D�`� ���3��@�f��� 8@��&D��#�!���lèQ���y�Ӆ)D���g,V$ �q��<�h��J;D��4��Wf%�N�y7���J;D��R�a	a���B׉H�s$�!�f9D��&1d�gh\gMXi��ּx�!�_	E�pb�.;na��A_�Z�!����œ1KF%C��D ^� �!�F
5DÇ˞�@�������p=!���"hW���G��ԀA�`*!�DϝaܜM�*����Ta�	!��oG�u�"�C@1�(��L�M<!�d �.��-Q�)>B]t���:(!�dL&i�F`�IȄ}T��:���<!�d�
P>�s�\� ̔��H�^!�I�&̔��S��������!!�D��-j�02�ݤ>
�`�$( 4!�$��T���r7M���<�$∰7!��z�H��F��{�T���b�O�x2�<��}�<A�m�: �(Q⊧1��9b�UkܓX�9Ê5O���jTq�T�ר<=w��+O�\��Z=?uғO1��ɘCꕂn�Bn©d<̚�C2R�T=�
$�O�y�&�*< Qˠ$�(��A:�'�Q�dɾW����,rcǡi��I��IR. W�D���/�u��!aǏZ���i2.��,�1� �s������>M�`B���*�'��>��J��>E��M\��dXj�F�	�����D���Or��)H#W($�K|r&�`nf�:�!L<|h�� ���e��y��4Q��� ��g�GŊ�3�[�<�s���#V��'�P���,��G�NP�O1��-��]-n�b�X���4{P�Q�Э��p��V�ֈ��?� $)�ٴ5H��m�_�M0��#P���6C6L��E�?MSF-F^�q�>���^�Hw0�jV�׀�҃�A ��?��^�M>B��F�I�b�A	V>/D�XGcoL�����<�t�г4}��Z�� ��
�` �B=0L֣?a���l2�	���O�<w�a;3@��.&<5�@�D4c����ONpB�ak����qO|�ZU$�}2���a`p5q2��hq��B
:�>�R�$6�_�^) ��(/�4���
�l�ZaВH� ����
���������sj��Δ� R��hj��ݨ���O]�xZ�V̓O�h��F�O?H2��E���F���z0TD��iI�{��`��j��Cu�K��V������+�O���4	�!S�V̑��M���a�'�H�kA�^ 2��'��=�ڔk���֫ɼ Ę-Ғ"O01�JòvnU�5��	����r�x+�V�둕|���n@̜(���2L�H�(����y2戉}�� Y�M��F� @coϲpa��4��'�x�g�DS}�r�0��z�L�Ҹ:�p��AĄ���,��k`d��^t8t��KT�lX`�Y5V=p�JTƂ;j��ȓi���*`� �	��� �=x.��@������R:��#�+�?f�\نȓ7�j�1�c�v��̃�G�,�N!��6lV�Ʉ3&;z�e�dZ��ȓ$�����;S���X��XXΝ��%�6����Z�&J�@I�le���ȓ[,���BB�Ph*�SӏϘ&<0���D6�єD� Ne\@�ӽ��ф�"�i���[�>�;�N�9I؄�\.���p�% �b�:�/�43��ȓ09�@�{\(�
��Z-w��ʓ ���PG��<���r�'��WL`B�I���	
|����'(�C�+c&�Qq!삓D:�%�Ё@u`C�I18�Q�EΌ3e� �Vd4G�C�ɛ ��TB�H�����c�C�I�NR����J�$I%�A;�C�I3|�p�V��|R'�<	;hC�:N�ұ�c3��4��<A4�C�I3H>��@U�R�$3�H�d�tC�ɗ}�!au��3$DF|� a~C�	1?w�|(���gZl����92C�ɯu�H�z�jD> zPLP��C�ɀ$�H�G`Ҥ2�
�z��\�	�B䉔T�ً��^	=��QHf��?;'�B�I�}�pd"�	8|~��2"\�dC�	..���hQ��oC�� ��۾Q%.C�	6� �9�/2���q�ŢH�B�ɴ#�phr#]D�2A�P�®g�C�I�y#����/B+WN=�"�\�$��C�ɇT�Y�Ɉ�b�\��F!��C䉒�{u��$�p$�a�Y�k,�C�I�@�>Ii�
��/(�G��%t6C�I���{r])XN��Ҭ�2C�Im8m�.�#�V&��T�C�ɂl���P�j�E��؁�G͇O��B�	�ֺ��VOfL��ڕk�F�2C�	�5�D�1M1 �h�f뉾&�JC�I�S�!`,��c8d�B0/lNC�	����&�P�[�R\��I�uN�A���fmY�%��[�Z����2
/�	1��H='����""U��!�I&�6X���Ɯ7�&L�Cg�}$!��yFFT񐫓�&�٢N�T�!�̾VƤ� fG� �䌱'D�=~�!�ė�q6�y����r�!����@3!�<2b�ѓ%m�7<oDԑ�a���!�� � `@H6R!�J��P$U{���p"OX]�O_�"���zQ+ܴu`�[C�����SS��� �����u�.r �V57�hbf�h�TJV��ClQ�`Ø&gt���%d��E�ᓵXd�	�*!��-C���8^}z]�5` ����-��d�
��Ň7�r��#[F&��BM�,N�����=OZ7�_�M�Չ�9����		T��hHa�?E3�-8A�Q�v��D���[$����)�'(^p$s0��$U,բe�,Qi⹊�%�B�BB�m~���u>er1Ύ6?Ӥ�+� �R�����l[�4`���b�aR�^Kt���ӟB�A3 �r��пF���4;i��@£WN�h>�{o[%m���E��;zȢ�:�3����zɠ�2�Z��	9B(a[S�.t��pf\ +��C�I?K}��RUc�$lw�z��-8��|�xB_7y`�h�f�.����ě�y2��kXic�����HAԐ�y��@.eN��P���%�F�%W��y`Ě>��@G�,��;���y�Aɮ���Q��qRP�$��y2��6,�)E	�r���u'�;�y2��6VЈ�P�eɸc����I��yR�2��J��)odH(�@�y�c���� ��Ð(Q�H|Zr	��y�K��ZA��B�HԱQ�4�y"K�%�p ;�/�0/���*��y�n�=���,K�N��aЌ��yZ��y��Qz�$)+����.$�B䉽$g��#W�ϣ*U��[�(@8Hz�B�Ɂh�RL����'Ki&��s	�1&�FB��5v+���J0�*�ddI�h��B�I�EͶ}IE��/L[.��r��+Y��B��#缑(��HFFl(Z�� t�B�I�Q^򄊦�Ɠ$�.��@þ��B�I8n�<�;���t"�YG.�r��B��=ja�T3t�#h�H0���Lx�B�I�=�|�r��F"z
ZyP�Ɯ�+�C�	5ª���Ҝ�`1��h]�dG�B�	�N/��u���^$	�-Z=J��B�I(]5h���и �Y��L$P��B�	- O&l��EF�0������\tB�	�o�&=��B�l݊W��=,DB��MU�!�f�!i�
h�wh]*EBB���@�E�\+'b��#Ƨ�;{�6B�ɪ�<��ˏ�I����3[�B�4_^D��U�`>ʖ�\"I7B�	(
ol�id֖".�RE,� �C�I�a�9���؛|�q+`�
��C�ɼ~Re�b��t��re����C�In�n��Mʶ:��(gEU,B�C�	�H��X��BU �X�o�8X�C�	 [�^hRoW_��0�U�\Z��C䉀���µ`�	&א��u�({C�C�	�o�Ż��Ze�X"��9d{�C�j����$K
=j/jT�(Y5��C�I�[D
|�$�ԣ}�\�	D$ܬsz�C�I�2P{R��C��:�fڄ[HDB�I�z5�}�Ec�T�.qJ"&�(L|C�	�d�ć3z ٢E.��>3tC�#F���s��� �`�+̀LXC�9�8���W>K��؟J�6C�	KKv���(|�@AJ'a�0rV<C�5�X��C�X�9��E�b�C䉲Z6FHxG�G�%Fr	rF-� z�B�	:LIx@�ћuh� �˞�]hB�I�9��jB�0J[<-��]?�jC䉹'0؃�O^���҇�N�l_C�)� N ��bǊSv�kR��$Df|dh�"O��"Eҝo���K�u5�Jd"OVu@wfH�o�le���L�-����"O��愙�"䲔ꁄ%
��"O��W�ݪx�hS���N���V"OX|���f�R�bw��'�r���"O@�R��H�X}��� �$N��"O���U�>Ӫ�{��I�1�� `"O*�1�� $�؝�䨛�(�ԝɃ"O�	��@C8`;��,K��Ad"ONM�6�+3VLᖁ[?�r�q"O
�c� N�/��`� V�� ��"OTh�2��,��4��N�c�����"O���ᨁ�v���-�B��0�"OV�	DD�%� u+qK�8g"�"Ob�ѳ��F�LA�ъ�+`d�"O�E��:s�P���Ӕs\�LK"O:�� �ځX��!�u����0)1"Od�Q֯�<}�(*$
������F"O�Iഭ�9/��	C�#�V�&�z�"OQ��ğ�J ��@�I�x�"O|LzVO|oؘ�j�(}b �6"O���O�k-nLB����N���"O��an��:ghD��$�� �"O<u�ѠΠ>�V��Э�!Xx*"Oޑr��76��b�L�98o0�{�"OTbv�,v�t-��AD�d��@��"Ov�X��ߓ!:Ѥ�[ ��Pr"OJ���m��D�.���Mp��dJV"O�ؙ��׳+�����*b��tb�"O���L9 ��d�V����ڈ��"O>$�*X-�r	�CC��I�i+�"O,�s�	91�6�p��E�i��Ujv"O�L�TG��$���*�Mڝ�<A�"Op9PӁ������1lS�7�2���"OD��B���X{�Yt R�8�`b�"O�U�񬌱=���8V�5�h�{4"O�"N&AĞd�wo@�S�$(��"O��cL#z��)��ǐWَ �7"O����ճ1��I��)H�yo�t�"O(��Ӿq�0Ƞ�Ρ~k>,��"O�բ�n��FX�B��
A�#�"OЄ��[¸�)p��a����"O@�{�)H)0�.�sǮ����=�"O�%�ą+�X�C���|���"O�剧+�{#�4�2�LcM�9�"O���ucI w�� "K�8B���"OF���A�J� �ʐ���L�X;�"O}�t.����B�@(L��� "O"�DP>O�5s���4X܎�rp"ON��"G�OF�t�rC~����"O�8��Ѧ>~�b��I��Qz�"Of���
K�iy��J5z䠫C"O�0�A��cj2H�UO�Y$��8 "Od�Z�+w+�f�dc\�+�S�"Ol=���v�]wDI:��YӴ"O� qd B�&�X8caㇽ!��{�"O�Px�"��)o���FE�8ڠ��"O�4���PZ �LAf+2?�� ��"O��9Ǧޗ1�-���.	�25"O �J�����|`#Dɝ�M�����"O��XF�_�ϼ�+ǈ��2�8=��"O �獝S��(�- 3��`S"O��I������kr�Q >�J��5"O� �H���EVʹ%A"��RX����"OXs��
���1AO?*1D���"O�E��'R	m���I.�4�����"OfM ��]�"�D+#-���T"Op�abgȀ*�p(ҡO$Zb%
v"Or�c��QX���☉BQ���R"O��ԢR5^6BS�.�--���s�"Oh8	�Ǘ�b_�<���H�;���x�"O��"�@3 ��S�ev��P�q"O��K��\�,(蛄cG+d�X�!@"O~��(�"�����
�r��2"O�kk&<�h`��C�K�vM��"OPD!UL_s2~���b�����C"O��1�"�Q����oU	����'"O@R��)�����E+��͢E"O���C��{v�3�� C_x��&"Oҽ�cMS�t���P�E+P��"O�C$.��Ǌy���Ю�aZ�"O$��6g@
k�,�b0̀�cR�*�"OzE�Po�+�����ʉD��у"O�zr��7+Jo�47�V�H�"OV�	�+�"IѴ�S�L�#_���"O��@/���mQT�SGJU��"O(4sk�6m����(�/(� "O���oޢ,�\��ue���W"O�$q��C8qu�d@Z�#U"O�������a`�i�#=h�C"Oj�)U�����$�A��(xQz"O�`�bg:b=!&�O�ƉS"O~����')�]K����F�h�"O�l���1s6��c�	j�}�B"O���k;7��̣��0_@I3�"O��h�*�B��� E9I�My "O�D�g �:BȐR�u)��
�"OVDH�+ɈW��v7n5�"O*\8�G޼�V ����1��"O�D+��W�H�A�J0i���y�"O<`�7�Ď>&�8F�ɤ˲](�"OKW�M:���b�4A���1��y��+W&�}kv�H>��sbֵ�yR$K�$��/����y�톓Oi�4Ұ)�'=}��a�X �yR%Z:�b��I;;{N���ý�y�F�1n$(ʶ� cXvHӃB��y�Q!C���'��*��0�B��y�Ô#J���d��#Ԥ���ױ�y݁M:��F���1��nH��y�'W�{���獟 ��mڷ�_#�y�!X��� sG����Gi���y2獜&�<�K��\�NU���7�y���5���c�FߏR���fȂ�yR
_��!��!ȉEO�l
5J�8�yҢ9R��}@����?��8rCE�'�y�a�?)���΂�>�,Cc`�1�yR��(}�9��/�>r-�B��+�y� ߐK6\Ȱh�jB`1�f�ϝ�y�h��.�*�A�F�bo�y3&M��ybfB&[�
�Ǣ�-S�t;�Ř2�yB�[|4����6[,�{���yr̾)�>�R�^2�y�X-�y"��1>5�iX!nƟV!49�!g�:�y�	�ޡZ1��D���f"���yRm������	 �xY��KV��yBDځ4�� C�� �&%VŲ�y
� ����1!g��Z��"��l�"O̹gL�D���p����씩�"O�y�` #D��1�/�:�P��P"OH@Q��)o>��m�*:�VE�"O�5�V��!�h�3���[eeA0"OnP�0��O�p1��K�TTN!�"O�	X�P/�0��
۞`?�\�"O��p�Lޚ^-���Ɉ;&d1��"OX`R�o*��B��n �D#"O��ą>²�
��T�M��	�s"O�Y5e�&B��:�͕/�␲�"O���e�)Yrp�P1�R��Bw"O
�����y@"��J�hB"Oа:Fn׳G$ �+7�{H,26"O�5qQ G9$2\��C�!2
��c"O�p��I����C��1\�C�"O�H�3�]6"X�d�T�0�3"O�ڧ�P���a"��u��Ru"Oּ0T�س_�	"�N34�X��"O�5��N#{g44��B^�M3�\�"O������5R��"�@~~$�#"O1���\���'X/DH�\cD"O��a!��,ʼY���3�5"O�XbP   �B��1)�͈d%L񺂈H��?)��?A��?Ɋ�)�Or��F�W<^�&L�7G������O�nژ����	���"ٴ���y�M��s�^��@�۾h�@���yR�e�(uo�5�M�i�M�O����ݘ�s��
�KH�tR��aa�
5�(�O�ʓ�?Q��?����?y���j���5'lI��P<p���)O��mZ�]�����Ο��Y��Ο���2�`�h��>����˽��d�����4{��Oql�0�;���C/8/!���@�|� �"\��0$a����nHb�Iqy"���i�!W	&��GDGt%r�'!R�'y�O��	��M��`L:�?�UB˰O֑���okj��æ� �?9�i�O$M�'~��'�2�Z�!���0���)�b��g����i��ɊIp����OB�a%?A�]	׺c�@�p�seoU�V��I����I��T�I؟$�Ie��a\ H�G2���K�JR�/�,<���?I��^�6�
����'�^77��ޑ+H��GE�?Ѝy��&f�O���O�i@8<6M/?��\��\���$R�FLyr�G��?�	8�D�<	���?����?3략��]�u+�'@z���O��?����D�؟h�w�<����=*�~q��O"@	�-	a+I�'�I;��$𦵨ߴ[���i��s|)��g��v����jI����*5' (m��G����7WҎ��ɼV��8Z�%GgRر��� nt�	�|�	ޟ`�)�SQy"�~��8��9^��ꦭ�VP����= (���Ox(mZA��TG�	6�Mkծ��E��S7�ñ'�C��f웖(|Ӷ�y��a�F�F�ͣ��)O�I��mЊh�����/%|qr�7O˓�?)��?����?����)�-gC�T��㖻rw�!����Pr��	�:h��?Y��k~��-e�� mH�~$ ���udp�$�O��&�b>�+�C¦���%b����}#���m�Jq͓9���@��O��N>�(O�I�O���d��v�>PCg��`��G�O:���O^���<aU�idȹ���'B�'�`	���X�P� 5��1u������@y��'���&�D���Ӂ��0��fސ!F�I(�`t2��M�&��K~
T��O����|��H��̨2]��c��=^���?1��?���h�󎒏u[����C0	p,��A�,90�DF���Ο�I��M���w���G{IH�&q��'��<���i	�6��=���צ]�'�]��F��?��� �PKԇ�/6���c��{�%��'�$�<���?����?Y���?��'5���*'�7�����J�8��ʦ}�Ei�eyb�'��O����b��uS񡆡��C�!���'_h6�Ѧ	@K<�|"�E&\6���L�HO�q����_*�����C��d�kSJ�@��E�O@�t~ňee�t�,  v �m���?9���?A��|�,O4`mEѴ��ɿd�^��F���H�F�
�牬�M��r��<���M���i9<�U���M�B��"!��_�����l�1|�Ɵ����V�������(���ɐ 9lx�v%O%y�Z](�8O���O����On���O*�?�(V��-f�4��.T�i�pj5�̟���ߟ�H�4B�Χ�?1�i$�'O��$A�"���eA��^J�bs$>���ަ�Q��|*W�A�M#�O��+5��S���p��K�,�[���#�����0;ʓO���|����?	��PJ�Hґ^hb-J����*��?�,O^(mZ�P�L��	柔��E�t@���u��M�+�Ĩa�+^���d�g}��'�RH:�?��A�G�izBu#E��&p�]㱮���|pK�N8Rۂ��|j�&�O��L>A���`L4y�+���M���G:�?����?���?�|r(O�l�F/�u�!�GS,���R�7�;��WyR�jӨ��ЪOH�Ĕ�~C�c4a��Q��͉Eƣl������%�����M�'�Y���	�?���RU� �@/vn���a�83��c:O��?���?����?Y���i��6��j0��X�kr,G�3�4�lڦ�8�	���Ij�S꟰�����l@"+w`@[�
B�0�A3F͹_ϛf�nӆ�&�b>��va�צΓiD���A�9�  9��}b���~1��O.!�O>1+O��O�CC�J�sJ�+�B�"��1jEM�O����OX��<ٲ�i$��j�Z�8��|���U�OvcT�3�I; ֠�?I�W�X�I��;K<)I�J�8�(U	M����OO~	м��	9v�_���O�����-�©�G���˰'A�zb�X�E`�'*�2�'B��'=r�s�u����5� ,x �OV�~=+pEğ��۴ɥ�Oԟ8�	��M3��w�č2A��U� x�j7.�'2�'��ț��֝!.��S*���1`�X��@�.���h �|�P�������ϟ��I���9@� R���3e�v �x���^WyR�dӈt3���O����O�?��uԵ+4�dB���%N���*��$WҦMY�4"����O����>|�t`�������	B�.`�bS��{�I��	��/H_�	`yB�Di��\S1L�ڀ	RZ�r�'���'��O���>�M��B-�?�CjԞYz-ٖā�a$ѩ@��)�?QE�i��O~d�'�46�N���1�4D�ň�h��L���3��-&7Lp��
�M��O���e����aa:�	�黎�� �'}<`1ئD�!z��$8�<O����O���O����O�?�˶ 'Bq"HZ��N���!'W��l����0޴7h��'�?9`�i=�'{��s��C��cd�h<*��G;��DϦq���|����7�M[�O�`S���0uh	 燚Tm�Ya�������Bp�O�˓�?	���?!��7�p)��I*��ʓ�HyJ��?�-O oZ�bO�(�	�0��N�t+
�~�h���r�8(�%Ԇ���Mdy�'P�� �T>�c�Z~<9�h��(�A��B ?,�83s菂3��!���$���$"6�|B�֗Yd�e��D�Vʾt7ă4Rz"�' "�'e��$^��y�4?Rڵ:vAO[\&��(�
j7I�7f��?�����$b}bKl��+��]�D��x���B�i!���t�I���[ڴ}y|���4��$ݒ	��t��'k!J�'$��� �ꏭk�"Xce@!T���Kyr�'�b�'4��'��[>�k�Şy�\CWm\�k1�@ҷ�^��M[S왐�?����?O~������w�����{ �(h�:��ٖ�'���|��TJҠ���;OJ�cfd�1� ����=9�Ex=O2�����0�?��C5���<Y���?	GC�rZ�l� �F"T.u���^��?����?����D����|,���O��D\1K�d,V?H��o�T|�帥�|��'����?����gz����ԓ(���y��D"Z��'S�j��݅!�D�Xp����ğ�X��'l���CAьj��0�猒O���'��*0��uz��)b�ݷ����B�'��6M��D����O:�o�p�Ӽ{�AҴº�� +�8ظ�@�F|?���M���i��,���i��	m�`�[��O����Sʆa�VH��F�uwL��c�K�	Uy��I�wѠ��r�G�Gm�Ukv�A	9�\�\՛֮_('B�'9"�i��7�2����^/$�x���"�|-�'T�i�b�O�O�*�ȝ-�Դ���$!�(p�.�K���J�\��A�Q==Ab+Ia�I|y�f_�+(zEs�ɏ���P��BT�'�"�'��O��(�MA�!�?9�E�*礜v�A}hX\��@�?Q��i��O���'z�6��lmڞW8ܨ�5���#Jdч�;n~дT�FئM�'��C#F��?o��O��ݻd&�(�ǐ�(|�f	S?�yR�'C��'���'Z���L]��тE�;f�21qU�8W���OB�D�Ŧr��j>����MC�yRe�U��Rj�20h,Z1��~W�'"f6m��iF�Y,6�5?�We	A�? ���c���\NѸ���z��
U�K)�?q��=�$�<y��?����?���L:��HK�$)�mA`�-`4I�����$Ϧ��#��ǟ��П<�S�����޹V\Py�	��i���5-h���	g~��'>�R�ԖO�������ԭ��� %6Q���S�yh��b89�V�\�S <��I�4o�h�6H�|`{W���b,F8���������@�)��wy2�p�2p�`Z>-�-�J��y02��!Ú`����OT,mE��_F�I��xx`��2m�&��1/X�[�B�2c���$��;�mo�Q~Zw�&ɂA�O�B0�'�f$e��,y��a���	f^�@�'���ڟ�����D������	Q�Ԣ>��؀�J�9x� �A�~6m\�$�O.��$�	�O8�lz�����}w. �۩ K����D�����A�)擞k9V�o�<	@���J��7��^�.��f"_�<�wA���:�����O��D�sH*[5��f���W̘)aH0��O��$�O�˓x����"_�	�8�BY�J�M��!�vr�YW��@�	͟�3�ORQn��M��x��{)`�����C(�(�������5���	��8Z�����1�:Z��X�l�ڔs��ҿ5��ɫ�l[_�&���O��D�O��<���k[�x�((H��ٌX�:|��h��?A��i��ēQ�'_��vӀ�O��4�b��BQuI�a��AI0^�fHP�3O��d�O����;]�6m2?�;s�N@h��*���էG�VJ\�11�G 75���9�ħ<y���?���?!���?��E�k���T��M�L�Pi���$���Bf꟨����D&?��I�Pg�Xh���W��� G� �!��b�O��n���M��x��4͌=>ș�FU�f��!��G2x�P]�ƆܨY��ɶS�-[�'�f�&�<�'�z�/
-$w�y0	���(a��'�2�'�����\�t�޴P�:4��U�N R���6����r���0�n�B�:���$�B}��r�B��	�tY2�O݊ٹ�f�7�ŮE{���!��i��ɳ����B�O��5&?����N��B�C�ܠW��-9��	ٟ$�I� ��֟���W��X02dJ���)d��	������?���^<��"R�������&�4ۣGB�k���˔�a�p��ȳ����~����R�\7-8?I^�$����ƕU!�48&
H�R� DH���mkB"�Q��Lyr�'o��'u�/��E�.1q�gә�|�:��߀X���'A���M[F&����d�O�ʧ�$ [����(������;"4��'�"��v��O0O�� xR���s┱"� ���Z�i���M
�2�HM���By�O��(���A�'�Ҹ��K:+�D�3��o��e"��'��'�����O��I��M�ԉ�R����>�[�	���4����?���i��O��'gB 
<�����w�0�)��Odb�'^\鰆�i��i���E��?�)'X��P0*L�
̸�2H��5�Wr��'�r�'��'�2�'��S�6��	4b՛���_�*L���ͦ)QB۟��IƟ$?��	 �Mϻa��z6cabplR���I�|���?Q6�x���a<~��?O*��V��d�`�{.V�~\���q2OLA�.8�?�ǥ(���<�'�?� �D�� )і�Ұ�
�ɢ&Ӆ�?1���?�������-�aI�̟���˟8�p坢7�|�0���7�Ԡs��C��>m��ҟ��ɵ��EQ�-����2 �hY�e_�1����'f ��ҀկD;f-A�����A��'5�3BjV1t�@�q����	��|���'���'R��'�>��I�c�����N(YE�D����9t&��$�M������d�O�)o�d�ӼKK�):�]a1L~�������<���i�6����e2eI����'���qA��?�{����Sq���4���M��nW)�'��i>i������I��	= LR�	�b�K���R�ڂ�<Ӻi�|U���'��'V�O��%ψ7�.���C~�$��P铧l����?�����S�!������K'��ᷧG; ilˡM�l3p�'� �`�G������|"\�T��.��IW.I0a"��5��������Iß �	֟�[y�'f� u�#�O��I"� X��b�m�3S� ��'��O�4n�|��b��ɜ�M�'h�6NV�l���q%��i�py�H��&4hp�i\�I#e����O,v|$?��݉��"�K�:�k�,I�OG
�I��L�	����̟,�Ih��|�B(cO�1w�b�bD/��"T����?�_������d�'{@7�7�dR<t������.��T�	�*�"m%�P�I���S�>���o�}~r)�8:3�i*��Sw2>d��E��c��]矠q��|�R����ן(�	͟Tl�]����n�X�#�P:�?����$
Ʀ�Q�蟈�Iǟ��O�\�)���0۸�PiN�,�,�i�O�D�'��'�^O�S�9��T��(G,#(�1)DI�6�`٘�L�+3O��3rb0?�'_d��Š��Cf`U��Q(D�bzd����?Q���?��Ş���Ϧ����ޑ<���)�ˎ:B܂tUbQ�(|��	ٟ�Iܴ��'�듶?�V V4�B��Yen9ʣiǡ�?qp�i	��վi��I�+Y\zQ�O��"��%l&oABDB�N�!gY���$�O���O<���O���&j�kQ=��b���=��$�6����?�QX�	џ�&?��	7�M�;KiI:��	O�Ȝ{$�W��rD����?�L>�|*���M���� |U�7�5e�>D�bC�TȂ��w<O�X��*�4�?�1�d�<I���?�d�\�X�0�U8:�!NP-�?I���?	������u��ȟ������i�!��N%��ÎS�a��ݘ�#�Y�Q����M�1�i��Oh���K+ze8-!�бU5LM��`Z�K�,�$�0e�_��-�beS͟��^Z�h8c���T�-�͟|�	͟ �	ȟ�D�t�'#�$a�Cڍ}����Y�_,X����'7-��"_��[f���4�ԑd�Z#vt�D%�n�^<Q�5O��D�O�oZ4z�,nZ|~"�ܡV;���#K)�0���p 
B��b�$Hh��|rW������Iϟ ��؟��͑8�@�����;4H!�$�hy�h��y	R��OF���Ox��@�D�\� y�烐
[��HsHA=&�~��'�'ɧ�OQ�@kW���\�\L:ƈ�'���3憶WW(��6_�(�g��bÛn��]y��51��ԋ�h�'����#%�	W%b�'�B�'x�O��I5�M���+�?	���s�ȉ����6JRHi��N��<�3�iY�O�y�'t��')�6�N�r\�%1��+ѐ�

�#h��p���	���O��\�>���o�h�كn�%I�"$��!�p�.��ޟ��I՟��	ʟx��b��?��u����l�B����K������?���(��f��	������M%��`!fb�	�g�	���
����S:��c�O��hܼv�Ɩ��`�n�0]�������%N&�;�D߳6�}��'a�y'�l�'�2�'���'����(@Ȍ\(�m��
�b�B�'�]��Zߴ@�z@��?����IЯ*�$h��<>�����E��I���ĝĦ	�����S��M٘TaX�B��P�B�$R�Zܔ�K5�?2����Q��U�KT�&�4U1���,��𒵧��@R��Iܟ��	���)��|y2�b�X�Av��l�橰d��Q���(���G��D�OX�n�_��\��	��M��i�,\��`×
_<�b1n���y�,	8�jӘ�_��a3����6�2+O�Y�l�d`5��	ӈ2����6O�ʓ�?1��?)��?�����	]�n��q�� !&�&�ŝ���nZ6Nv���埀�	x���������aR�v6�Ꞿ����%�&(��Lc�r�&�b>%в��Ħ��9h��[s@�������#��XΓ7`A�j�O�bH>(O�d�O�$r!	�&�,�C5��g�h��B�Or�$�Ox��<A`�i������'M��'�Ř#�>z��r̉�7�H��S}s�0�nZ1�ē+b^|!iQ�o�=y��ۊX\�'��1yB��:��Ց�������e�'tl�ӗP�$bM\�|qse�'�r�'h��'L�>��	 
������F̤����V�`*1�I�M#�KѴ�?���
�V�4��C�z����7F<>��K�8O��m��M�1�i%%���i���y�
y)��O�����(~��T(�ڬ#!�j�dy��'���'�"�'�R%�>aԜ� ��/[<vE[ӂ�lh�I��M#�蒚�?i���?�O~b��S�c�
*h�b�#kX_!4��Q�@�ܴq���k$���W�>���Y4��b���2/ P�p%+�jGD�ʓ:�t�#�L�O�H>1-O��"ӠJ�jf��S���I��*���O��D�O��D�O�I�<���i2`��'�T���L�������7JL,u£�'��6�>�I����[즱��4\�����2��APbhؖEܵ
ca�=3*r5�i-���Ym�B����9����z�b䄅U\`q0��dN��'6OZ�d�O����O���O�?}5C�9,&B'�C A��T�6�HGy��'6�7�L�G���O"�oL�I�t�Y4�S W[�Pkr,��@���HH>a��M�'��kߴ��$ƂF:��1m�'m���Ɠ*�M�
9�?QҦ(�D�<!���?����?�F)ʬt`�8�0�\?$�|�'���?�����ʦ�)uA�����ܟX�O��!�f��9V��
�ۉz&�=��O��'F�7-ݦ�	H<�Oa�L��)��. �%��/+m� TfJiHF!3���9��i>U��'	��'�X!T<Z�h k���N��mq,�ҟ��I�����ǟb>��'g�7�.`'������*ZQNe�V�2�P<�g"�O��Ŧi�?Q�Q���I�Dp����51�ѺW���H|u��ן��S������u7Ċ06����cy�"�4�p)�&Xnޠm	Ӂ��yb^�|������	����I�l�O���#`�4a�JbC�ʈ6��a)5-z�b7,�O��d�OГ���d����݀`4:P[@e�<E۴�����4�j��	��'�b>i��� ̦I�*��vH]�_.�yD�{ -�j�`Ep�"�O 	�K>Y-O��d�O��� �[� �^�`�!��;������O ���O<���<	��i�.����'�2�'o4�;�,2D� ����3�(T�5��DF}��'}b,#�Ӝq���:��6\G�c�9I��	'l⎀��@�%r�c>�Ғ�'�q���o�����I�5�$T��� MC�	�/������.܌:6��Y+:1����M�͛�?Q��jR�V�4�<���́+@6��һ)Q�d�C8Oܼn�>�M�Ծi����i��ɤvɢ��B�OS���6�y��Ѐ\�N��4�M�	wyr�	"ǒ�qmO��;!�/=��6ěV����'�r�� �X�^Q �_�Z;X�f��R!&E�'�P6������J<�|D�h�? "B$�>�t���o��F@*=3rḵ##V˓[. A�,�O�� O>Y,Oh�q�fS)Q�(��ř'>`����'z6�`��ħol����ӉjJ�h�C�0�N����I�?��[��������I8L��	z cLW���jC"��!(ѺU/W���'8�TO�?���Μ�D�,��6�˃X�f�X�i�:e�`\{gL�:`w�l(��Ӏ3��x����i�|x���̍D�]�k�0q�0�;�I�,L)pщF�Ǡ:Q�QzQ��E�,�!$AP�t��
"�_�ZD0��'�V 9i��N8r��:P���p������2a��`F��� y�V�IT"D��R�K2J�	�ы��dɢ4�eÆ�9d�Ҳ@W���{�F��D�D���ߍL��Q��qC�x�e�� �-�1BR�9�!�wE��P�}A@��/N�K���1����MJ	e��m�dչ�M���?!��h(�z��d�O�I�X��H�?�^=��i�/A�Dc��0��0���X���v��X	�;#�͛,lxq'��M���-��9��x��'�r�|Zc��h��L��hQ�q�'B����h�O���{��'���'�\ʢ��*��yW?-`�BG	Z��ē�?a������Đ%<&v<(�B0!R�H��U�r������O����O"ʓkcv1��3��i�n�8�Di{�Lٞx�E��Y����˟t$�Е'|���O�H�Q�>9�@7 �T^�wY�P������	|yB`� ��l!��>g���&G�S��F���	]�kyr�����'c�}Ӡ S KȽ�Ҡ7b�2|rݴ�?����DR��nd$>u���?��@
��H#W
Ҝ * ��D�����DŤ5K��'�~�0�wV���S��0�2un�oy⅕"�J7�Yg���'��t�4?A�k�<a�"��N]j"'��i�'g�=Z��4��'�����I �'��� MW�D|K
ᦩ�%l@#�M��?���*�xR�':p�+�4{�jxs�� �"\P��nӀ����)�'�?�BN2FK}+�"1�(�c�@�D���'b�'�*p�4�(�d�O��d����P&�(S�B�#䁜��L��+'��;��b��������	�d|(�
�Ŏ�pW4@H�]1z���4�?qE(�lʱO\�?���d����=�Pu�����A�*KuQ���7�>���4�I��'0�T�VɃg�h�1An8��!6�ߠk]:O��d�O��O��~�(p��%�D��j��^�0Ip��A��?����?Y*O��P�$�|�t�UG��|���i`l1�*�k}�'b�|W��
�O�>)D
�3;�Z�ۖ1:.x����i}��'�2�'���'���I��'��'̜����X�2�-*�ȗ� ����2'u�z�D$�D�Ox�$�����xR-R�Y9u�ФHD�q`fG��M{���?���?!k��?9���?���JңC�64�ю�8�����	�0J�'q��'<ܜq��9������-+�.����oy# eɣtHp�yٴ�?���]u�(���?����?����ƺ�ؔ͐��2�J֮ߠC6�Q��i�bR�h�E�3�S�ӣNZ8kꍕ\`����?/]v7�Rd����O��O����<Q(� A���:����@�x1���o}�˛#�O1�x�d� '���0Um�!,
�;u��X�n�n�ݟ\�	�\Zǉ�?��D�<���~R��&h^�}����2i2d��fj���M�O>I �U�E��O�R�'��	��h�'�(%�,�Q$�B�'@7��O�]h�DAE}"R�L�IJ�i����[*af�e�v#α��z���>ч��>�䓘?����?�.OB�ѧ�Ч;�t "cG�-$:��D�͛k��p�'������%�x���� ��X�Q�\�PpD�MfE�� \�=���IRy�'�R�'H�I<x&����O�̅�:tx��!�Ҥ1h��4���O`�O��$�O&8p�뼟L�Iٕy�x)� ��:Z�(���>���?)����Շsa�M�OU�I&eʪ��Ԉ� AsM� �j6m�O\�O��D�Olb�d!�	��9��]$����G/FN6��O�ĵ<�@(����������?�k4�;�8;���5'+5HD. ����O����O2�X�o�|�'�I�2(H4�0�EC��t���zt��R�l�g��M����?�����tV�֘!�&�X�I<L7���t�K76z 7M�O4��J�w�@���}*Enǽ%��t
�͋5+R�᦭�bFR(�M����?i���J�Y� �'
�!�a�F,��"�9r(⇄z�8��gk%��D�'�?9����Y�%jb"Y.���s��^�9ܛF�'I��'N4dC��>a*O����3Qo�R
9 ���"'�&p9�	-�ɪ �t&���I⟸�	������N�*����S���@�ڴ�?Y�c���IEy��'ɧ5&��g���!!��� 7m����^G��O|�$�O��D�<q�f�6���'���8��۠k����f[�,�'Vr�|b�'W")ϮYX����#�m�~Xi6,�=f�aR�'S����D��ٟH�'��m��H|>����D�(P��+R�3�:�tMu�v��?)L>����?A�)C3�~2�U�tȅ��LǏ�R�������d�O���O�ʓ\tn���t"]� �xV��g7�!Q�뇰4��7m�Ol�OB˓Ϊ������D 9"m߮!(����!�=�6��O��$�<��s!�O���5�L�/u̬*u�G�[n�dqcP�����=�&�0�ɯ?� ��SV�Pԛ �*r8c��i��I�^Pe��40X��˟D�S���I�N�ZI�7�Z=��D` T" _��Y��U��˟��J|�K~n�Ld!�f�r�H5_�f�6�Ç ��$�O����O����<�OdPa�P�$Pl�P�Ě^6�I"le�n� ��U��1O?�8�M+[L8y*�&8X�L��/��M���?���e����/O��b�� ��2Ѝ�e���Q��ۧG���<�V�U=8���������/=����0(�<v�J�Ei���DP44� J��p�}YZ��b%i�d��D�p]�$�3T�S�"�Ye�c���	Dy�'���0&�I�T8�w˪�1clb�IџH��a���?1��<��\yw CR�1a�e��m`p�,��	�'�"�')�R����%��t�T�.���Y"O@�p��M�!D5��D�OB�:�d�<AFmZ��?�Ѕ�� ��,��M
�K6�@������	ܟ(�	ҟ��'*����&�i@�c5�t�^H{` h�唘rK�1o��'�T�'�j<���'��'X�d(q���j�S�*�+$ o��t�'����-Y3�SƟ����?�X�MI�,R%EBI��}��k!S	�OZ���O���̖.:U1O���`��$��T$vC����:.d|6�<�`'_R��f§~����b⛟$G˜!J��	�mχ8J�p/p�j�;<x}��m��O���MK���?$h�s�l i�Vp�^ݦ��f��%�M���?������x�Ou�\!щY�H����'�C^�yr�''T�u�'Q�U�x&?�P�X�	7���Xe�3Şpt�i�B�'��]�.��)�K��3g*H$>��5K�b٦G5���%Z���': U��%���O ���ON9#�s��	R��}��|��@��Q�	�V8�J<ͧ�?a����Ě�j��Q� ��e~.t�BE�8%�0Io����a�I�x%�����|�'�6��e�H�!?x��D酵*,~�9��&\ΊO^��O��ħ<q���?���+Aܤ}-e~B��#,5^�ʜ �ś��'���'�2T�T���̳��4'b�[� M�6�Q���M�,Oj���<���?���+�b��HN:��V�����I(���� �i%B�'P��'�I;&�`ʬ�(��
}U���b�D�\���٨c�&�nZ�l�'�"�'��MO��'_F�qDչe�e"ĆD�Q�>�/ F%�I�`�'���~���?i�'<�vq	(7H���Z��LF����]�D��4�	�"(����ħ?-{�D=g[��4� ��%�|�`�paԤ2�i���'f�O� �Ӻ���R�|�aف\sJ,�獌��]�Iџ8ᡪ&�O>�ѴD\NG�I��\#�R�4W"���i_2�'�B�Oz8듥򤈦W�����(	�Y���բy�lZ4u�X�I����'����D�[�B��&!ޗ-�D���◦5���o������|��$��$�<����~�#� s�>��sG
%��`��4�M+L>At��<�O��'�2�܇*% ��:Y"@�&C��v	�7��Ox��� �D}P�t��ly�5���*�Dj�J��7Y��2�습����'���O����O����Oj�J�x5��o��N �Őe�9I����s�3Q���ny��'����L�	ǟ����ʆ6J��5��N���$ƌF���IKy��'v��',�I7'`ls�O ���(��z��� ���R���4���O�˓�?����?AC���<yU��F���G�:p�!:���=O˛��'a��'��Y�`��o������Ok�c��(bL�gO
q��\]��f�'V�̟���韀I��n���I�$3�㙥\ź�y#�&�.��DE��M����?�)O`�1�̏n�T�'��O�r}£m�|�%�4G��*��>���?y���p���?�.O���-b0H	�l�A"��̜WÚ6m�<q�DY�Kf��'k��'N����>��EQ,(��JL�~�,q�/R���)m�ş��I�)j^��2(��A�� �)�� +�-��6M�e�D�l�����	퟈������<4T!��{Ã��C��!��1���ʜ6�y�X���F���?����Fż���hL6>�셺���3:����'���'wYy�(�>�/O,�䳟l[��>T[��D�
L	Fxf�s���$�<��G��<�O���'U��K�̉��^�D:,%B��	��7��O��8�HXe}r^���Ityb��5�ٰc@
�����B׏����Ʒ��D�O��D�O��İ|ΓA��,��/���ua�	��0�T��2|J��oy"�'���������ZBh��(�E�v�هPp�Q��aQV�	֟x�I����Iҟd�'��Q)t>�ɭ7���b7g�u��q�$��?9,O&���O�����3��TrdK���+�h;��G3.�l�����Iğ���ey¥����?�1�d#�ۋL��r�HőL�m�ԟ,�'+��'R"��1�y��>q�K�h2�L�q�\(J ̐�ci�Ǧ���ڟ��'b�Q��~z���?�'Y��M3���pv�T v(��^��@�Q���I���	�q������'��	�)j:ȀEY"x�@���NY�VR�$Z�����M���?����rY��]>nlX��'ҋ{�@�1tP�FЖ6�O��D�����O$���O��>e��D� �>��q�[Gp�Ǣ|�r��@ �a��ӟ��I�?���O��|%���Q�KPx �k%E��o��hp�i_L�x�'��'<�t��MA�? f!�GfW:��@I�*f%�i[B�'��\:d�F���D�OV�P����ak�6e��Pf�,!z7��Oh���O���6O�؟��ן0����[�2�h
XZ �!Ύ�M�6z�L���xr�'Ҟ|Zc���Y�c�輜��m�+�,�p�O���"7OR��?Y���?A-O�]
qmC?s�\�J���x%�A�eB�o����>Y����?Q�{�����]�u��z�Q�1,���%T�<Q/O@���Od��5K��|r���"f,��ha@^Qֹ G�EP�I؟�'���	؟`a��g��Y�g�1F�y�҄dh�C �����d�O����O.�[?d@���4�ѐ$�d$�BÅ Ii ܻ@�IF�7M�OJ�O��d�O*|�=O`�'f�	�Eh[z�5a'�۝g*�i��4�?����䖓L�T�&>����?I���]��!BAE�
&ff�agDի�ē�?���t��t��������y��)4 ŒR]�$K����M�-O�e�&�¦A�������2%�'~�S�D�K��M�$�&����4�?���|��p�������O+>���M�Y��=���6AH��۴A�B�+�i1��'���O�fOL�DE�{CN\�3l�K�Lq�'��	�Ynژ ���Ii�I�'��tG42��E�p�C49|B-h2o@�g�&�'b�'���W�,�d�O������a�l�q��q`�K�+��I��<�ɄvbDb� ��ԟ��I�e) rʜ1*]�3d={�،Bݴ�?q�J�u�O��D%����8Ѓ�`��+]nHU��ظ����"(�H�ĺ<	��?y�����!Ūaa-ռ0���L�27ÚYC��V��矰�	O�矴��̞�p�T*1P\r4�H�R��P8DJ~���'��'�Z��� ?���O0|80l"��N�p�Q)�P����Op��(���Or�DR�C��d>.!HppkG8\�P����Q�]���'=��'�2_�L�"-��'p�27�$���:F�D�5w��hd�i��|��'��.0I�qO�U��#��f����	��PPгõi��'��	�s�(��I|*��2�����ht���H�l�
a��VI�'��',4˜'��'��iX�rt���fи[�*��@̆�3'��_�d��'��M�qR?Q�I�?� �O�)��IN�ɐaJ�J��ic�i�2�'#-r��'i�'3�[?���:'d�a&�7�Y�6!@Ʀ=V�D�M���?���
����:R��1���S�t�ݨ��.g�&�nڼGv �Ir�	���?�`� X�'C7 F�C�C*˛��'��'�J�HE9�4�r�'�n�Zt,����Q[�f�D��-�ݴ��'tz���$�Ox���"op�%s�օ/��Qрg�IVYl����B�����|"���
=��Q�<Wp��Ñ�'	�^����ݟ��'!���:��iZc�_03�8x��:V��	�c�'w�'Y��'��'X��O��$�s����N�;C�Z8XC�i�j�{�O���O��ļ<�L��A��j��][��Kd�ʘ
a�;R��'��|��'�qO�a�D��^θ����,�l�Q�X� �I����jyR#Û7p��N ��[�
�-�������&�ɦ��Ig�	�����I"�c����B���,�k��2@�ӣc�����O`�DJ�*���d�'`��C�-s�@Mz��AO^L���ǞA�O��d�OB<{�t��'�(�kH�5��P٥	�9{�pmp!�ݝ��g�)#��ˣ#�H�HlhQ*�3��Q��~Q�a�+حA�������B��-��Ř�q�����
��g����ߧqqԉy��\$R�Xi�w���Vܦ�zVƟ�`�f�jO�`���� ��3���3�.�jŋZ(��]0qB��T�ֈs�oD�L��u����	|Yp*�<:�L�A �fleJ��H�@8qB� &��@���˼�v�0���?���?YƱ�n�d�O��!��!]el�c#�ݹ=�����"Ux����#��2쓤p.��Zu�'�X���?>"d�R��.kR�Y�H�% � �C���0E6l�4�����2�S���p�֢%�ҽI�a�i*F�� ����Ɵ�G{^� �tG�{�� k�G_�Q9�&�1D���w��m�� 46�$�9�/P��HO��@y���]��6��i��k@��n�֍��)ӄ�>���O:�d�O�8R��O��>͸�C8B������QGa�"���|YrH��v�LIx�P 1o�5?Ri��ܬt�)�r��/��)9�皮>�uC�(]kx�4!��Oj�d�&`D��G0*a8U��>�^�=I��y�B�cD�X�IDi�2	��C��qy��)�G�y�tLB��X��	#��D�<��OPG�������O��Q�ֻz�0(�D���RiV2�'.�,ϊ\���
�&ڳ^�րa��O�Sy/~��T�Xu~��/ʟ-[Ģ<Y@��NA>�"��	h�I�J|�-s�v�jE�{?r�q��[�'�����?���4��	}�I�ޝ��kD�߂�y��'��,��[&Xx$���ĒM��x��Aى'mT�I4@F8ƪ��􅑝H�-p�'\�5@��>����)�HOR�'���3��d�턿,�ڽPנjZ�bb��A��x�`�ѐAc��T>i�|�)� :��%� y���'�,M�:Us���of��ʃ�o�E�wi�0��I&C
;O�q�'$@4%��c')� ��TG�OBHS��'�⒟��>�O�PF��=���IT��-�b���"O���������$KUN��5�6���HO���HL ��,�di��ő�L����px �������	ß`�]w?��'�f,��/�R����kX�ad�y�'�>E#�
�-h����e O��2�I�H0�!��%w�"E�O������_��9���]q8�i�n�+2��qW�S~�@S�����u��Op��<���ɁJ��hu��>8���2�+z�!�ٲ9��#��s^��S!�
i�n�Dzʟ��cB�b��i���r� ��EU����ƃ~���ك�'��'���=�B�'j�(�O,R�'�F��2����X{�$��}�HԨ�IG8�
��"a�h�yV�8 ��&dء=��u0�E=�O���f�'�"�ۚ�<(6�N�a�l+�o؀W>�7��OVʓ�?����S�D!�/[��!�0��ܩ��%���y�"T&S����eBՍE��0�A��y2Mtӄ�nZqy2c�>@�F6m�O���|"��יl��Q�����q��N������?	�GV����i��'�哋Yn�X�L�R�0@C��=r��<�5�(y�!Q@) §{�p�ADf� &�kZ�*D��GyR$��?�T�iaJ6-�O��'m����C/�L��c}�b!��������d�*���D 
�X�8��BS����D��4�?��L�+�L��-��(B��@G�<�1
�a�^�����?I)��%�b��O����O�x�B^A�v���葴|���w$��@ ��ZG�|ҍ���IW���a�����]-w)���D�֤@i��c�|���'���Y���p�x��*�K*�!�!�A��'��'+b�s�(	3�KnCN*�(I�M�r��G3O��$'�Oq"�M>U!楛F��q�!C��	��HO�Sl�<9��T�$�� (֨J 2``��	ğTۤBʮjz� �I����I� ^wr�'̦��0��c�	X�-݈:���!��O�PZ�h�%���������СR��Yh�F=C&h�FMO�i*ց�I!���Cǂ��6쓥ҟў�����Z��taD>6��[r��dH���O~l���/c�u�j0*P*�׻|B�I-8�6��1�7l� �VNV_�(y��4���=�D���,jQ�X�|���Bw�<	��_)0
�yr�F#I(M��q�<yWZ>q�@�q���y�=��l�<I�Ex������@���QWA�g�<�����U	����l	PV�d!��
d�<%L�g��ӄ�0�^5ia�G�<�7aʌ���a&D�!�fQq E�<I� �&j'�+�
����WH�A�<����0����?\�v�Ҡ�B�<�UÂ./��r
[6u䀆o	d�<����G��ӱ������oPZ�<�D����5dZ����ð�	U�<��m$]8�x�Ҁ*��Tː�O�<!w��nn����Z;Wq��:�ɅA�<I�i�:W�l(��D�6csx��Ҁ�F�<a$��BQx|(KY<o���F�@�<gg�B��8M��i�MP���H�<�)�!�>�Q�;t�ҍ���C�<A��i�pib�K�8MQ�3�@H�<i��L�+���G+հ6 �WF�@�<����	
��+t��LHgm�|�<Iפ��/�l��&=f@D�R��u�<��⁑o�$j�!,+��+Fj�<QW��v�\��!��]�}���Q}�<���80�L@��������x�<I�\6��FiϿ[I@�KG#�v�<釂Ƅg�F	�%��t��<���o�<Y5L�\����J�bZa�<�0o x�� ��&߇u�$t"3nO_�<ɐꃾ7��@���,C�@����[W�<	�Nu��c�σN��=���O�<� �l�6��?#:�y�������`�"O�y���DFk��h��K� �R�"O��Q��ɴ�b(BgN�0�8�Q�"Ov���@�P^l��/G�0�kQ"O����e��_�p�O�@9,=;�"Ol������M�BN߂z�0���"O�12�K?-� ]�f�<_�V�X�"ON��fH��h$2��	|�2��"OjX���ޫE?�@s��;ph�	�"O������(O����S�cW�(hC"Ot�[� �'wsxh*��,Fl
�"O�]0��!w��=��T�V8nyb�"O�U@�>xx��W+#rÀ�"O(8��
�R��7�8{-��ذ"O �i6e�:W�j|�3�ˊY<ȲV"O6�+FkS�5��b�±�t"O���b��kҚ5��Og��q�"O8�&�R){n�a��OY�ض2"O���ş� ����F�̣h�(hs"O�`T
A�j@H�@G�c���"O�@:�[�ء�6]�zSv-��"O�y[4aRI��BJE 7_>��G"O荂D�[$4-` �FE��,Cw"O*]�p �9e��y�D�p�B�0"O0�)w�d�������-k���U��ʃ۸h�b��|�#��Qh��{ūƴg�Zq!���k�<��J%lv���/�,*�Vy��*�}�..�FY�5*��4s׎�T�!w,)>��� #8�O�3W���0\@��$"�/7W -�eF3j�*�IC5��Z��&%�,���+��B�:�T�.�>����0�[��O=���0����DT�}$r.-D�;k��-��Q27��hVN�<�7@ňB���zH>E�d��;9t}8ԫK�8ZȘ"p��+�y菘c�F�R�[�/1$y��b���+94Y�gb��0<㫑#Z�`���`J#��SD�a<Qc���5<<%�c톣#4�԰gHβS�ܝC�R`<�G+E�A���pQ���T~�Ժ��T�<��iיswt����W�v�6�z�<�6�	x��A�ǅ�2rйV(�v�<�"A�j�p@ C�:q��Bq�<�����</����^�a����qG�m�<�d��`���8����c�l�<qj[�
b���fT|�����HL�<	��W-(��##!� 0(���B�<T�ԛ:�~�P��X]D�e/�f�<�7n������?H
��@J^�<��S# �����75A,��s�B�<�sMMTY�i�2MX�r,@�<�e})"���O���j�� ]�C�I5n�-�B�)K��e�䋙�}a�C�	�V��iÅ
��&$bC�k������)�rI@`�'#%4C�	�B9���eC�w~���m[�/�C�I�@g6�˅�dB��1Y�DC�	�;�Ց񮓟7��E#B�֦�C䉘7K&�	"oq��0惔�5��B�I.jH-2B�B�L��{B-��5��B�I��\�k��^�yz6��:S!��tP����L�v�Z5#��I�<;!��A�l!�u��n�840-�K!��L�,5Z��#�J1�����D(|!��R�(�S�5(}���&�K�i!�D��nRP���I
�c��;���&!a!�G��"��5
�!%Y��5�to!�� ��!���	v���  :/���I�"OD��ъ�K	򔠡l�#?uvtk�"O��[G��1
�yA	];7X�x�"O��B%��  �<{�2�J��$"O�ؘj�j|�0ځJ\�F=��"O ��s��o�Ɓ�Fʇ)1�@!"O8�؃*G\�E;g��=
���"O`ô��6=��l��9���"O���K�U��h��LP�W�vq��"O��i�M�FĈb�S��<1�"OTc�oI?1'��'.�)'�e�"O�8�k���H��O��LR�"O����+��xŏ�i����"O
��%,D,��:�[�#�D8r�"O��P��P�DP !�#W��@�`"O�I(6��/^X3A �("����D��'.���l�A�c�>��Td��V�uɓ��`�J&��h% 9j��Aw������L�?�x����L���x�ʏA�t�3�֢��[�����o�1�U������]<`��`��S�z��Q��܆>RC�'e�Ɛ����=?�Y���Y�E�N�d\�(��s�N���[��OX�B韽�q$>
��m����/�2Ȍ��'1|O�pi�ٿZp9J�4h��<�s�H�V�`M�9�@E����@���H%+: ��":Fx� �2¥  i�F� �G��0<鐞x�O�+��-��� ���0���y��~�cU	 [�I1"�>���dz�(hI ��&:M8Pk�`�@?�lcF' %m�D��@�'*m�d��af!B��X�Zc��?P,UJ��b2����3�(yG�HbU���[�T�&片1d��"R�aκ�K!`2�Ĭ�3pJ�T�Ou���'��^7@�㐧xx@(�'��xȷhU	F�uB�4'ndi� �g?�t �SҶ3�ci��Y��ú���)����8�4���8GI2u0� H�!�~J��'? ����L�'y*�!���8u8��
�� r{�٪/O��jb#л3��_�J��-c'���O�	`��i�n�3�0�����I�NJ�b��)xn�7�6pM���Os���#��>� �%��+�L{�'������2ؼ�5h�T8��+p(�%-�����	P��7��B�X�f#��?L�bT	(;�0��~&����%QW�)�3��BԸ-��HI�Bቑ�f��C	-'F�	��k �g�O��pf�߰ 0�O��OF}Z0����Y&���rIC�^y$9��'���o��=�Ip��4��������㊨K���Ʈ�����?�D�Z�'�z�{��O|��y�l�)f4tfk�',HI��	��o�X� ���3t����͝�*H|��f�'���0;Z���nxɩ���*�4����2䂆
J��V�	ED�񤏌q�xM Wg@!���^�6���C��&4�6mK���q�	=Z���OW�)@��5^w��A�1)\�M� ���߯d4�i��	t؟�X�2�\�q!��mu�P����-�=�ee�U��i}�p����,_**g��<-'J�m�:"p0��@�i���ɗukX�z���B-��q�Hڋ����3���MI�5J�i��;,����Z�;��� [H�; �ϕR���3�!�i0��>�ᩀ+7 ���V ��p�i��p�- )C��%�`ų�ȓ�_��@ZT�<��b���r%Iθ_2ƨ���WI$����!k��[�x��pH�>�p<�F#ו0�0�ڍw��l�� 	�(��\7,GB��:'��d?���ڪMpR��[��-s�Ń�.[�L�� ���3.��6�/�Ok,� ��t@!�υ1� �Sw ̂��D4�~|YaQ;q����0�A1������ YiL遑f�	wz���㓂1�) ��!OxM���O�__��"�@�B���
7�J�@�B!3�%�<�N1�C��2��IĘ|B��:r���K� c�"��w�������}9�ǅ@��5J�9`6�G�:���g�.y�@m�d-̝k���2$�*=F�%܆i���	�鍲<�}x0+
!Ӹ�3d ֺ �)�'���G3��6���`���߆3T��Q����I�XCխG��|l;EI�(A�X��`ρ7P�z��C�ϦsԴ�Sč����Y��@�Оx�.,°��X���{�� I�a~��w�t�`�b�
���Y�e>0:� J�qOf�*��j���
�G �'�������u��ښbh(��.W>.�xIB��R,'�џx��@�y�m�#E�/y�0���x����Z�=�~)a泼X�D�I���O:Y�@�Y0X+�L�S%߾?�1��>1��(��s�0�B�23��E��(!��ajo�؂�-T���'�аd�?<:rձG��>���z  �.	�@��+G=��G���G��퐄$,O��	#��jd�|F'�s���J����PJ�p��*�' ���:����t�����9���4�Zl>�ٶ&Οz}X\�"O�kq�����'�j8#ԍ�$p��ѻO�07�3���"�I�6������ �S4�P(5n���N̄Tt�g�'���s&�_(�UJB�r �����b�Zgc@�,e��*�H�+=�q��	�z�\�+!��ҥ�u�ͽHZ�"<�E�"`=*��QN�oİ�HW�\�;���k�f8�o�0�~H����7�LB�I�@[�-RDFQ�*��t�+�p����%��!�
�+�lX��W� �Q>��16�*���.X�F�H#���C�B�	��xD�!m�#tͨ�y BZ�c���ĆW4:�=AӀB�g�$$:"$�?�Gz��pZ�[�,̝9�h2pV4�y��$q��б��W2CVJ�:�n��y��˵2�z`(7�·5�6���Dɢ�yBfH��H�E���
L�E�ǻ�y�mF�Ap��?Y\��Dϓ)�yB#�"Ȋ9�A\*ezԸ#�U�y�I�@�U�H�sʜ�S#͉:�yǋ����Ƨ�d��2K]��y����`��C��6�!�T�y�bǹ��y� �[	���f�T��y�[�9!�-���%gv�$z���yr��/.����_��a*ꑕ�y���r�LA�3+��u�i�mI�y�#�#�:-���6d�n���`�%�ybeޜ#C�����J&\� �;"�K��yR���Pqtf"��9C`H��y��8:��12�FD�]��*�yr�A-]� 	���Ý;���s��� �y"S�mT��q6ME� ~�qs1a�yB��a���A#aݣ'��jrCH2�y���1/[d4������]bb�ϵ�y"	j=��O]Z�>��rl���yr�%K0�h��˾OJ�x9�c�7�y�%ϡk�`��G�<Y��Ȑ�ڗ�yB�)�X5�� V��
���yr���AD,��BG�S�|��U�A;�yb� ^��5@&�[�P��m��y�aH7D���Ǩ�AZy9S���yR`�ʀyx��M�<�j�*3�P��y��:Mj�Z� E�:**�J7���y�ކ-#�ɵ��'LhA��ډ�yRn�'*<�G�H+&�z����=�y��3#qİ�7�V+h&�r�+��y��]"g�] ��E�\!@D����y��y
��H� }��������y"�0ڲ�h#+V%z��)!�dݨ�y�c�����lQ�ɩ�K��yr+K�-kr|ؖ�ǥZF�I�Dߦ�y���i�~��ϕ>c�Ȩg)��y���e�Te�׏�x�c����yr�^�Q� ]aV�//�����K6�y2Cې%1*��ܰ� 0R1�O��!��D8�x��w�~T�C�n�!��I�
�d1�	Āp�F�x�.;K!�d=�����̖��qH&X�y�!򄛼T.i�4�S�#�Z�2�AE�!��G�f8J���-�@��D�e6!�o>@ݹ�.T�R���R� O	\�!�dv�}[pH5�!�r�8|�!���RpKU`ݹ�`��S./Y�!�D���pQ��(�d!GgY�B�!��q�$Ä�, �9�t�#F�!�/4Ĝ3򥂀oO�����Ft!�$�+%��c�@G-A*!�U'�9a!�D�D�N �w��A��:�+�3�!�ޫ��£�:A'FYԈW�{�!���P&6�#��ԾX�%��*�%!�� &�#�"ؕ+�$���o��(����"Oƭ��!ɒY(��oZFf88{�"O�Quˋ* Ќ�k�-�8b��L��"O��QGΔ"k����Ӫ|���"O��`�B�Z.�y��X��(\2s"O �y��x�vYI�J(2,<�r"O\)��!^�T����k'�!��"OtU��ɑ�ĝ��Gķ ��*�"O�0!��+(r���)�
Y l�3"O��gɍ�D$��Ȅ|[T��"Oܭ0��IA�h���G	�,Y�"Ofu��N��|P��OX��W"O(1�����}���3&» ��"O�� �I���uR��F>~v��"O�"��<���c_;dh,["O�	��ͼ&�ΐ��Q���%a"OP�*��Q�t����Ѡ��@��]��"OJe�K0D��Q�)߅~�22��y�����杈,��ل���Val|���3�y��39��7��	Yx�@C]��yr��lZ��dJ@5yq@E�X�y�ɞ;>"�`�E5$+� E��y�k��P1��[6�{�l(�y"�Zc� ! gT0���#%��y��M�m4L�����W8$�b���#�y�Ɛ�$c����h�K�6�R蔌�ybƂ�yH��!i�/:�@YAoK#�yA�n�� 9��S�5�p5��� �y�kN�?.U��?b/���ìS��y"�W<#�`��d��_��,j�@���y��
8i,��;r�Q���Kc�2�y�����<�I@M���%+c���y�,ݶz�B=�EB�/�q���=�y���z&��am�{��r6 ��y��M�$5(�a��x��c�e���y� �5M�@�gJ؀p�+%� �|B�	m虪��@U�p�;R��C�	���f�Y4{H�i �-U"^rC䉈BKԁ�uhђG�P����bC��&H��� 0	S$O�`y`�MI��C䉘~f&(p�nJa���C��Y
�B䉌:w��j�*G�c�����˺$��B䉂I����AAPqd�!$�� �\B䉾;�@��&O%H�r%�ͯN�"B�ɘ'�n�Ꮟ''���#��d��B�	�+�^d�ш� �$��f�@C�I�$F��xF������G�C�I�$y���&�����͗D���[�'De&�^�K���ɥiL�hw�}�'@��I�n��q`��(�:b�d	h�'���{Q��o����5o�cg
���'��]�elR���di��r����'kڈ���^�k�h�!� ٍi:�P��'��8{�Ɋ+PE�ӣ��a��}+�'�,�!��qo�AXCʄB~��I
�'��S����A���
cj�,	�'b��� �\`6H�C�p��U�'ʽHe&X<r�JD�$�Z�n7����'�0����t�����Ƨtv6�q��<$�d��O'TԀ}���̓D���9++D��G��t�,)�Q�'�]�q�4D���ag�������X��,2D��hBc�;
�Hh��ģ}޵��#D�\�p�O�S�t���{`M�A# D�� \��b  0�=a7�	#W���I"O�,�T� ��ڳ*O�!X�"O��e�0*�de{u�U%w���ʓ"O
=30`��}J�(D @٨�)�"O,MY�H��E��R�J�B��"OT]��Ƒ�5�B�a`FM�te�b"O2�2���b��� /ӎ}���Z�"O�b�g%2�j�
�$�}���"O.��G�
=	���V����r�"O�h�$O�.�r�fL<x�\ �"O���W鎄y'2)X��Ҁ�3�"O�`�ujU�+$4�ge�kÜ�w"O�J7��A������,_���(t"Oh\3ꈐ�n4�d�R`[@�1�"O�cՍI����%��|X�0��"O~%aF��!���{%�ESL��"O�(p�I��b�@�j�@͵G#2�
'�'��	�WO��! N�*	� �:�)@% ��C�ɗ=xd�� ��+I~,U� 9�tC�I�@��`��ֶh�ڤ�$�P<�<!��T>m�BN8M��h��JK$n��	3�&Ѷ�hO?�$E	m�$!�Gʏq�vIk�-�7!�I�`��၊ZϾ�[Č�20!�G�=����c^3f�N�2+#a!�䈅/��(2�ˁ1��)��	֔{�!�$HBE�t0��N�l�$�X�F.p�!���&10@����(�����1~�!�G�W@���c�)�,�r0��B]��=E��'_\��t��'�@T{��A�BO���'�Dx�d�N��X}�B�/N0@��'
Y�2�T*	c�L�Ώ0/�
Q#�'��	sB��/P|��a�@*+K����'�H��FA����R�߿L�X�'m�U��'f����G�K��h
�'�`�`���(�ې���?�tyr�'���w�	_kT1���\�s��s�'x�K=�<�O�q�mj�'�n��f��(,��$����j_2�j�'2d(����~���#BUY�US�'��س�+e6�8QcIR=CJ�H+�'?�@c1MK�.�X}�CS�<Ɛ�`�'�Iq���U���	s�9]�aq�'��<ZGA�t�@��Ӈy��[�'ˀ퀵mf��և�o�tq�'��\�U-U>I��k�\�bF(=9�'#�`:gl��)ń$R5N
+����'�¸���2 ;�z��W�UR��z�'����&&U�!��oN�?���'>ex��J5��Ё"��'9�b�S�'�p,
�.I�v�d
�]�)X)��'\��ٔ%�� @Rb�N�#����'3&	��Ϗ`�F ѱ�ߦ�p51ܴ�hO?7m��*�83�E�6�����ɯq!��Ԡp��W딱���"��Z!��5_��pg�O
!F\av�]�m!�;Qq
p��ح1
�=�܌6d!�$�6���*Ʊm0�����:t�!�$�O*�h�@�w������x8�p�"O�iG��l	3W�gF*�1G"O�	�dH�\k(��LY6x�K�"O�\H#[�w����D�ҽЬ����J�O�0Ґ#^A���0��-�"ts	�'��\�l&@p�ݳ'rrH��'��Q� ++L����(m��
��� ^��p�;aCp �%����@��"OT�3B������D��t(W"O�|�K��&����8F��9�"Oδ�WjE�wmPI���� y�0I"O,�ۄ7Q,x��1�ʫI��4��"Oj���k�T@�����S� �'"O���M�X@(D��។\|�A
�"O��1���W��� Q�M�)wV, u"O�� ��
#�f�sV��<{{dx�D"OlL�`�>P��bf���9o~�r�"O���֨_���F�|~�!��"O�q $�M8U~�81J��{VQ��"O�]�5�ɠ	��2�h��uqJLI�"O؈�wҾ'�ݠ�͏U��-C�"OR=���؜1V��eb
6$g��F"O�����K��	s��E~T����"O�ds(�0E�*u8���J&�"O�	:�)B@(ڐAІ�� @��:�"Oz�aGI.h�b!��c�5z�bQ"O�M���Y�����0� ;�D��"O��3�H�v���9���Nq��"O��{f�06w֜���݇33��"O����V?�0��F�A1�Q��"O��&E��!�U�r�,��6"OF����5=�$��-�����"O-�T��^��SGC�:	�v8;"O��T���"idQA��&�B�Z�"OT�[��&ex�ZƂ�=�4h�R"Oz�:�Sn��0����"O�����v�2����D�xp�p"OfL�Gm[�W32�Au!S!r��� "O�ӦE@-oJ�z�C�ٔ���"OBDÀ욆�Z�B��D<� 8y�"O�dʑ��G1�ph���-[]�� "O�$�W�Շ*�JT�FMTt�rDQ"O��蔥�j����տd���`"O��D�W/q9���A�l�ȱQ�"O��)�@_�5�� ��^�@A"O$(���U�beP��JӉR���&"Of��`ŉ�זܱE爂&�r!�"O0(�4��?e��p���
�\a� "Of��bH[�D�Y#�DF�	����"O, �Î��;� ��H��=i@l��"O�Ի&dL�[n��"%'��T_HD�"O�(�d�s ��c�)lUnXa�"O�܀s�]�'��qKgcǲx.�H"4"Oby�v�C�E��J1I�58����"O���B��	T������a����"O�dg�7��sKՇi��M��"O����O#&��37�R�H���7"O����ê�9AT�K��m�c"O�u�"d�(V�k$e�2�AU"O(p��I�D ���ڭ@�u��"OP�J��?�(���C�:��i�!"Oj��M�A�I惂x�f��t"O`a) 
B�.Ӻ��F��6��Q�c"O���$�z�X��!�>Z�D��"O@�x���΅���zx)ۑ"OD�R��ץN��w�ɡG��{�"O�l�fo�$_nP� L��E;�T��"O��Y���c�^��sa[!#4ژ��"O��h��M�!b&W̴��A"O��8���;n8����I�9�5"OLQ��Κ
��$�u.Q�$ my�"O� h�N:~�֤��'�3��"Oz�3��_-j*( �&L�7�~ P�"O4(۱66H�Z�)�-`8J7"O�q{g	Ͳ<��JpF�6(��ѣ"O^�ѧPWx��EՂE���%"Oд�6@�d�P�*բ@0�201"O���A�AL;�|���x6��"O½xTϞ#م�C�ଘRT�z���$V�q��84a@� $��Dʅ��y"�ۯu����M ����ˈ�yb���u���I���-�xq"��,�y�b��2�J���F7F6U�q�&�y������  �=,,�A�s�,�y��Z�HTwŋ�)}�!ɦd��y��<M���Gm5s5�C3�y2���Q����*k��]��K$�y�EÈ@�z�|+fFZ$^Mƅ��'� i2�H�">�����l�0ZĀ��'u<��@&u���2Fg�P��m
�'B<�� F�<�
u�uG&;��)�'^�q��	`)^ؐ6&�/<j���'�(-h�I��]�؁��)bB|�r�'\{���=���ɵ��q1���'1N��`��A��`��S�W=$��'��1@e�N8��!��/A�JӂZ�'�b����gdD�b@C�B���"
�'$�y�,_�T��uyS�|�blP�<A[��b� ����	C�C�<G�ӍVؚu[��Fh������\C�<�OܺUN|�!�!W���Ňi�<�&��bYB#�K�h.�Lq7IK�<�KW,4ۤ��u	��w�@�p�R�<鲦��[�8�T䝁C4���b�N�<�R��+V���I�k�j�p#�GN�<5a�.���kDc[_o8<s��o�<���=h�� �,U2`��jk�i�<�&lI�!��s+�т!$Wi�<1W��<#h�Ѓ�疬g�~�R��Sf�<�Dl�4<�DT���F�wM��enb�<���S͊�����)^cZ52��v�<Ѧ&���(2KԺl�0b���W�<��e��肰�:b��#��J�<���!L�,� �8<�ډ{@!�H�<I� Ի_|~�����l��H��Y�<�u� �-��E�G�Q5�����A�n�<qS��L��!�t��)�0�#�F�<i1�\�1h@ږ���r�����_^�<�#9�<�PcZe�:� R�<��oV8��#�f ޲�f��U�<G��=N( )�#	��;��Q�<i3+K�=�6(�W�X���1CuC�I�<Q��|��Yi���&x�Mc�	G�<Aƃͻ9�|��bcM�L��� �A�<�D�ڰr\Ÿw �+ ��qʧON@�<I�mK�M9��a`�<3�q�Sl�{�<�Ǯ��&��a�nڸV?��s��q�<�$Nބ]儽*��A�p�S�i�v�<A�C*젉���]|����UX�<ac"�4^v�� ʃ��8<3�M�<�p&G#���;��Ɏv"[�'�G�<q�f�;1��IHBB����P��,�j�<)f\�mP�m�6DT�RPr}2Q��e�<Ѣ�^m�Ǭ�e�2J �_�<'
�K'`d�� �by���*T�� p�Q�hVͬ�kaO��I�$��"O�8��(r<�����:Z����"O�0�p�ٗ�Q��
>e����"O����)jk���k� j��s"Oh�Hw��2��y��Y�xo 0"On��"�S	��dqpC]�"f��R�"O�<���k�v��+�!ZV��2"O �1o��:e|�Y�jͩaaB�@�"O�\a�I���e[�)
S?>�R�"O�ř��A1!4q�ت^~( �"O�P�K��	j4br�.e$TH3@"O��(��h�����'^�h�"OT52�d&7$�{��Y�[	�1;t"O�e�B��X2"�wʑ�Jn�"O���Qk��<�9
2��9'�&ݒR"O�5���+QF]��>�%�"O�MZ��(I���`��K3K#�i�e"O�MSB$=��Ö�Վeb=
"O�4Ï�]�)1��Y�n�|t��"OT�@I�6�t�0N�u����"Ozq�$�G�H�#�G.Өp��"O�$�8��z��M�l@14"O,��c��P<���
�U�R� &"O��X։L�E�.���� >bX�h�G"OPSą�]v��"׎"=$yU"OH�(PEJ�[Ɯ� BB�o;�;B"O�5��.vQ�ѓ%A�Z�\���"O0�K �Ag�  ��=!~�A�"O�ī��ܓ`K�����bl�"O�!0�BJ��L`���`j�i�"O�������B6��)	�Ds�*O�D��YZ�����؎{�����'���A�	 0��*͞���'`T��f��r�A�\3s�~Ȼ�'���c%�y�x�y&l\�iSf���'\&,J��G�V�b)�)��r�,2�'�2d���L�H��x��i�*"�`�A�'�0=�C(�f�tԫ��$� �'��mz�E0"z C������'��T�RF|�Q�0�ܒ���9�'��c�����ĵ���M ��y�%y����X ,�{��߄�yr���+��q�R'C�t3�xXW��yC�.w�ȜaT���>j�E�6����y£�MeD�pêِ3QmA@���y�o�
�ҝȥŭs���1-"�y�fZ��v�҇ː�8�^'+���y�F�F���T.�3K�uk��޻�y�J�+[�}*�m�5?@ك�.԰�y��I*	M�iQ��پ}i�yhPc��yrʄ�*�eA@٪M
\�� )R!�y���
�i��F�[ͦ��R�J+�y�R?5X�4!�;��՚�՘�y�
pJ@PG�~j�"m��y"f �Ce���q�'~�����A��yZx�ᄄҌJ�q�G��W)n����񳟈դJ@�>$9��]�,qAf�"D��fB����;���g��K��3D�� �?�C���#J�4Z�'5D��	�
�5*�~AP����^�l��e�8D�	����8�P�`H-aL��'"D�\���~�%H��Ȗd01P��%D�T��nA�vc��Rq��E/6����.T�̫ZRdX1��L�x)Z`���y
� x�x� A�,٢���)m�0�"OD\��nհCFf K�`�<K��)�"O�1�Vʂ;	�9SG"[ a=���"O0����_�#x�,ȃ��'38y3r"Or�1��@hTuR��2�*H�7"OnI)�0����l��x��	��"O�L��bڊ̊ [���3���A"O�	�h�9�TsuJ"d�M`"O�ЋJ�)�rK�GC�FU��"Oԙ)�X?8D���eF&V��]c�"O"	3�� $����
P4�>y��"O��kUI�;Z�v�Ӑֱ|�v��%�|�'��Oq�*�듧�!gj
|�Ec\�,�`8Y"O�<xԀ�Y�朰h\4�<u�"OL�d��5S����&&AP�"O\�Ba$JC�ĨVݡ�1س"O��k+:B�e����H��$F"O>��#Q<ltz��̶v��yK'"O��ϓi��|;7c
�n"2�Q�"Ob\����<;^=�� �����"O���ҵ494�2���6��s�"O�8k��!�Dt�t#V�O�X\�W"O��P�7W��ذ��'*z��!�"O��H�B�?OrN���dB]v
��P"O*E�.�?5,�g�N�BZ0y3"O�-���Z.���2$��&XE���"O�ɃC%�!�����xOR�X�"O�@��(hS,(���(%aE"O>�҆�ݟ � p4�õQ�����"O���c�baٰM6cB IHG"O���G��r����rN͓�p"O����7=�~�cь@�Mcv"OZ�Ka��2K��" �d���9�"O��x��כj�>}g���"�qy�"O�,�eO"�v��ꀐ͸��r"O�$�6U�<:`����$�����"O����_M����ªf�vq�"O`9%F�Y�d��Z�m��	�w"O�ʖ��WT>�ҳj'u~&�"O �iA#%ƅ�,����A&�j�!�Λ}M�yPN]�!�����R�.�!��ٺk�K�N
ss�mk����~!��B8.O���0P�)�e�2G�!�D˔Q��m`�g�"(dk���-!��W�`Nf��b��Q  ���!�d�~�b�D�;bo�BCPm!�Ē:6S����as�a[�L��`"!�D�1C��,l�� ɐ \K�����0=�%?s3�LauI�r��%�3�W�<yƠy=�U��[�q�H��}�<��#�U��A��P�b��j*�s�<y���v��;����%�3 8B�ɒk�@�A����-�cR>X�0B�?c]�I�$�4W� 	��S�o�B�I:5L6�"�-�h����/b��O���-�S���; 8P��D-=C�@����%2B!�Z�OS>���ȕ�.�6�Y咏*,!���!!|�%Se+
�]�jE� ϙ6?�!��&<�쵙�T ��%�r�D�gu!�$�;�6E�2�5TkQ �*�Ly!�D�T.f��k�=d�H8�G�):ў ��mg�E �֙Q?��(�K�o֎�OԢ=�}␥:L>��r3fߐ*nB���G�<�0��(VL���t�3�|<�a�[B�<� �����P?L����
�ț�"O~d���	�vg6�1��D)��y�"Ox���'ЄJP\�#���]$v	#"O���ǲF�����N 4x�8�"O���oH�#���y�O�^kI���'�S�	B�0�`��V��i�*���E�(�!����h����N&����Ԛk�!��ځg9��a񫙓)
D��F/�!�d@��T�@�&պo$ �А�B�Q!���S��0�ף�j����h�!dD!�N�X�F4
B�ЊW2����N�p'�O¢=�����f�,V��=�W��5�Ҹӆ�IO>q�cG�`1�Ý����*�,D��Ȗϊ�J�H�A��V�f�xT�.�O��;& Ř �F,ϘA3A���\I$����ϟ���I�BFk2�Y���O=SwZC�I���$�č�<�4��
A
G*NC��#viW+D;|Zh|	!�
�O0��4�)���	<TV0�j�<#�C�Ie��q'Y��:�
V8E�~C�I$5���٦I�PLr�F��P\^C�,"#^���r��dC��5v�6�OD����.t>�J���B,���1�!��.yP*a�G�
����N��ls!���Q�mIvi?)t�x��l��L�}���fn��V�p�aI�I�µڂ+D�(��ܣ[,�ړg��$9N�	�#D� a�WS���FY�0��A''D����lǾC��Y�ք~�p��t�)��O���&O̸P��>>���ǘ�L5:�"O�AgJY��;�*���P
�"O�X���9SV����.�}�P"Ovi��J�R�X��r�=43j����� �S��Z�a T)�[��H�I��RU!�Ĵ7���s�D�qp��S�@ӝ
Aџ�E��N�
��5�3%Ӎ;�^�z�f��y����_p0)���hZ.�fe8�y�%�3Mv��3���'i}�\C�虑�yb��P�j��c�T�4%�A�<ɰN:"V�Q���q��H��'$�'����9X#>�S�#$$b���$C�I�*�,Y
�%߶:� c�V ,��?���	�hFZ�#�
����u�3ꓐq!��@�Q=� d�&-�$M
UOQmX!�{��pyl��J�\hx6@�eX!���E�Vx;D�	!Wp(t�6��F!�G9<����9a~y���A�qџ�F��e���XًT`܎+�<��cd=���hOq�L�Bw�
� }�ƚ�@pH`"O�����[��k�$ɤ ]N��e"OF9�gO�e�i�4΁*��=�2"OH̊dj��$)H�� nE�\�$t��"OD�!gY,Xm���Ш��� B��N�Or���aK��s�ʶ
��7�H�ϓ�?��y�nͦX��I7&��w�t���ϊ��y��!<�DsѠ�w���
RG�y�� =��:Wf�4B3�����\�y��D?�(���A%:2F�9r�G��y"�"~(��]<.IR\���S��y��:j+2QK��#%n&�)�yiӄ,�i�Ǖ�J5�`[d�.�yb���"-����.B ��t����y�H�t5J����e+v,��n���'jў�O��Z�N��A��`���'��Ձ��� �!pǄ�_��uS$Ii��Q)c"O(����U��D+�h٭i��T�"O�-�#�Z�"�@�
S�ry�dR�"O��ê��$�%bW�S�����"O0D��԰8B ��V,r�
�x�"Oj�2���z���0'�ݵ�Ti�"O�T�-�� �L���'�Bu��"Oht�eP:>�t��Ѣ@7�n�r�"O�C���=�U���"4ht`�"O�]ٖ��awFPp$HS���|8U"OFț#B�f�l��X�Y����f�'ў"~���K�F����`� v V���$Zv��`�fTL�����0/�̆�>%
�X�9a���!.:�ȓf�	IG%N'fK~�0�̆2ކͅ�T�| `�n����,,��,��'�n�wm�i�F=��+�*V����Id�v>� ��ˣ\��SdS�H��0G{��'���ə<YU�D�F��:\в�'aHK����j�p&EQ6�r%c�'�����G;;f�)��o�(av1I�'��<%��O �����a 9
�'��P�g����\��������'[J	�kJ�F͜		��^�s�d`�'�L�c�K�������&�>���]�������G݋Fk(=sf�i��D���O`�E�.CB�#A�y�z}��'���ȡ%�=��x� �6A�4�"
�'M<����G�P�N%9u��4x
��'A0���!<dd�`u/̓,�	�'�,�`Q��7
]T����W�FR�P	�'U�p�2��"kt��C�9�N@�'��hc�ȃ1̠��D˂
�L\;�'[�	��L^�?|v1n�+yϖ�"�'f�H�G5[�Z�[æ�ik�D��'-Lm*��ɴ���%i�
��'�L�8�F��y�d�h^2^K�ԫ�'0�L#�E6Y���p��]"T8��X�'Ť�����I�T�7t碰��'�A���ݳ�%�j���+�Ǜz�<9�@ߞ3��|kPov�@���z�<��Eڇ>�����	A�&��gn"T�hR�������0�����Ls(D�T�� �f��,Kp'Z4k��3«:D�l#����F)�s�A�*E¬���A:D�|���ɵL"����̔�{f�<ҁ�2D�tSwF�Y�bDC7�TD~��K�n%D�\2Ձ�{��!�጑�_
VSW�-D���ďG�G�Ld��o�r,�g)!D�<e�Y�3�� �� �xp}ڕC D��#����]1�.S��2e�(D�t��+2D�0q�K_+^� C�1D�@����#o�HҐ�]�s���ۀK"D���� �X�U��$0������|�<�e�[�P�$B�d��D����c�'�?����JԺYHtm�?w��M+D�Lk`eȆ�&1����@��=D�����o�.=���(��ikL1D�X:AA�8�\)1�R�9�fJ +,D����b4N����#!&��.^_!�D��R�fDS5L��7^Q)��Z�0m!�䇸#ۀ�r�$[h)�����7D�!��ǚZdLʾ �肅�XM!��܆gp�4�P�F���Pbf�:~�!�� �̨���3mB�ᅊS3WbR�J"Ob�#ABv�:���r�4W"O�	��Q�^�VآC���;g^!�p"OX�@�J�.����Ff��}6l�8 �'bR�'�Na2���1�&�S�(��F��q 
�'��i[ ��W]�H��H�.����'vHh���X?��`�& J�A�'�>Q�S�[�L!��
;�bU:�'ڈ��׭M�4�(�E�Ε��%��'ff����&X����%���g4�|A	�'�pM��*I���(d���Y��".O���D�!�%�pb��e�!���,e�!�M�p�~�Ғ��/�0"�H
2q�!�]���P���U�z���G7 ]!�V�"�v�{�� :�2HQ�'��M!��<:: ;�5W�DTP���C,!�d�_��p�ǝ%K�@�ag>K!�F�"'ތ a�C<�8�01�R0o!�D�"@,��#�ʒ�_f���BER.c�!���)��]	W$җOZly��,�!�������iI�uP0�B${�!��  ��Aޣ`Eldh��!5@!�$+(�����A $�15��m?!�d�k&�@���.98	b򎓦*?!���i�~����E��;���;'�}b���iV�W,uF:�`ď�2b��葕�#�	_����cAz��0�@�M�-�$�yRE^a�(A�5)���c����y�N\2	>�ta%1��P�d��y��5/E�!�� �Z.rI@�!Z-�y�eؒ���A4��	Zj��٤���y�F�="�䭠0g�%Et~���ʠ�y�aN�]���:�����Ak�
�����!�S�ON�-��a��xV����>�P)��'�|Izg�	�n���Ƣ��(�]�'���( 	�4���"&��+/��j�'<|��b�B�7#�d��,O�0�0�����hO?u�;C���v�ɅRLN��)�i�<��e�0��d�1��%����Ogx��'�.a��Ɋ�,�Ѐ��Ȯu��ݰ�'F���"��2���dəjR�L
�'�b�p�"�_~d	f��1i��I�	�'Yr]�Q�P�)��`z�DO;qK�D��'zҩj������F
k��ز�'J����L�bV���#�PQ�D��'�:����\�Z<bTř0}@~���'1O��ҡ.�2K�A+0�U�-b�)�"O�M���ۏB�$�'n�4K��3�"O����m��p��ՃP�О���"O��A����e�+��<k�!"O�a�\6lT\z�ʕg�n�0"O �SŮFg�ĠA-�p�Bg"O����/B&}�}��C9unU��'�!��W*�p�>V1x��X#w�!��MkE��R4���P�*�!���$����v`�K���4P�!�䘚��!�Оj*����
�]�!�E�Yk��AmB*:GP=PC+�?�BV�P�	xy�O�����"����D�C�[.����$4�)� F��r!F!,\6������Gx����b̓1Ȩ��D?4�PR�i�oJ*<G{��'ھI�6� hXN�(��@% �Q�'�^a��ܫ(�ʙ�b�NZ�$�
�'�T�j���B��Ђ��IJ�` 
��� @hAQ��^�|�cB�m*�S���'��Olb>���N�z��9"iFS֜�Q�2|OTb��D@�I�AB�O�1@�f�
$|O�c�� !�Hm�4��C��7H�)��!"�Or��(7d�U��'�N��b&Z�9@B�	�A��H��`&�: /k�,B�=hF�)���I�j�X*؁1EB�1/8��J���.���Cĩ*�G{Z��F�d�8�z��tȇBB��
.^��yn]�T}pQأ�VAMLU�����yR(��"b�y��E+@8�|2a��yB��gF��%>ր��	��y"oԆ3*��mҮ0�<�H�=�yB�������	R�夔F拤�y���)�Ҍ�5�A�Pa)����y2��b��� .�M��ef�0�yh�eB4$"R�4��Z�a]
�y����E ��&���.� �j]���=�S�O�-�A��nD���d�#@��A��'�b	+dI֭Mg\��7��3��	�'	���%	Nm|��n��^q�E��'D�Ms�*�''�Hsu��#Q�a����*�'���0oK��v ����R�d��ȓxܜ8�r�ZO���
<R�'����	���c����!��0��$5�S�O���E*�;K>�AԃO�Y�x<��"O\�1�)Ѯ� ��Jg�hjd"O�!��D�{�L��r��1kX.�6"O, �&^�ȁ��j
�7Df��p"O���'�L�0g^s�d<˅�'�R=O��V-̇$��Q*d��H�\؛���9LO,�*�/� ��j�O"~Ìi	�"O,��M^���W��zM�#�"O��pSC�5�����،?fd�	u"Ol��6�Q�L5��n�,Y����"O���#�	�*�RA�L�m�C�"O�$� D�T���bJģ��P!��'9�y��$\)�X%��G�r��&8w�!�φ]M���jJ���5E����R;O������:$8}*�ۨ`JR�cd"O�m�I�YR�4q�SF;�!�"O��`��W/h���+���l+hmq�"O��+U�L F%�`���0ذ��O2C�V�}�68z寏"m��`�0D�48$�6si4y��BOg�*د��y���`�8���0-����6��?��M�����H6���7���1�8�'�nl;`�	�4cM��KP�~����'��Q���h���sΚ<[Q��'Y0���E�<�T�^y��K�'P���ǂж �&�y�M�"�)�'젽�@B_����J[��\��'��yŔar@��D	
��:	�����M�(� 0B�,���p��ܟ!��X�N�01c�� o��p��]!�d�9<��)��E�y��Y���,7!�D:+���IBj!O���Ё��S�!�ӑ:T�����lDya�Z8$!�t�TL�4�ΑC�fL�a���!�$׊]f�9�$	�5�XY�̘!�D�0������_iBm���!�!�Ąh�Нh�K�-[��AF^ Dl!�/ڂH�%H\�*���q�û>j!�ՇZ+H)�a\+#�p��t�[< m�}"��� VYSc�07�6]���!.���""O�mj�$VqR���h�%��P�"O@yK%�Ȯ'��1�3��9�*�:��0�S�	J8x�&��Vb�Ih�oG�X!�d�\ߔ�2 =S|)�î�E!��"vTn�w�uK� �,Y%!���k�8�s��P8v��t�2~�B1O�Q��0o�蔫V��Z�1"O���%�LB0xPm�lC�"O^�X6(�H}p�I� ��F�r�'�dq�G�MYiCf ����Y���0D�t�"[uT ��$�>:^�q.!D�����V�nj`p�O����4�2D��E�='�l�T��hiXZS/<O"<0f��?^b�ꗚp,\�����e�<���β�E�3X��駦D��yRoJ�zwN�"q'�0M)nț����O#~:agנ
8��j��#���̌b�<ɧ&͢P	�̹A&��<Bv���
a�<Q K͗[C���\ �t�#F�Y�<)���jkƐQBn�-�����W����<��	bبB�iA�&!r��U��L�<��h����NԎ[�J�qr�QE�<QT��8��X�'�Ow8�)�AA�<y��O/РI���S	����c,�w�<i�׀KӔ���%0��uyS��y�<����f�|�Y��S�Ɏ�2@�p�<�0K�� �x�+N?Qvf�R��q�<�`튲Vf��Sg\%�90��\cy"�)§lPmY�� ].�zl	}�4	Z��d0O��P���$Y&�	p�p��)�"O�PY�#D�B���H�*�06®L�"O�H���AI���Q�ߒ|�X���"O��!n����F�K<B8T�Z�"O�Ї�&�>��t�`)��͒��y�ĕ�^��0A��8�ap�
�y���yH��2w"�2�\����
��y����5d@���4-�<�s4���y���2$H��u�^"'h�];�ǖ��Py�Nv)^��
�n��D�W*Sv�<yVdI�idhc%�Ԓ4,����v�<)& �x��0�E�8Xp��D#�gx���'4L��SM©kPz�yc*�W��ݑ�'� ��ND�Z�~�[���%�̥��'?*TX3+�/m�ؑ� �,���'�V�����H�b��w�R�
�|�@�'I(]8�Tyc`h�9=���'CV��K��(ؠ�����&'����'��U�ʛ�@�����IB��� i��$2�`@��	�:Z�����"̉9��*"O��"dŜ�^��ӢL�@�1yB"O����cQ�Sp( ٠��.9�����"O�(M�@���b�����&"Ob�1e�3��!����+����!"O�L;�i�e/��J�#�W���A"O�<��	^���@mن� u�"Ov�#Pn�-k�-���_���
5"O��ʀ��v-K���c{�cw"O�t�@l�:v�$��C�R"e�j("O֩��J�%m�F��%��<c�"O��7�θc�ip#��[y��@"O�E0�^?�>Y��ō=Y`&m"O�h*�f޾oj�XG��& R,�����D>�� ��>�ء)eDޤH�0`��3D�� ��; a<J3�I�N�C��I�%"O�Q�W(!�p����%Ѫ8��"O�}�gO+ �*YU��>���"O�D�3aƺ�L��L�U�D��1"O|�k���y:���A�0=0�"O|@+7���cf	B��ʫC�~�Z�"O6�!��^.3�T%`I.��ђ�"OB�����C�,�Q�D��"O�l���$H�K�N��!�w"O�5:#ω;9 Z�^�5d����"O�CO��0�j�ޑ~K��h�"O��Y�*ǈcO��
6��J��"O��P�O�0�x1Zc�G�Z<�8Y�"O���%�C�9C�Ӈ4�`}�"O(@�4L��(TBse:p`L�`"O�<���F�R�Rׁ�%,Peja"O�,e-�Ĵ���mT	h|�BD"O吥��#��q�	�I�j!�"ORT�M�>�����^$r�#�"O"�i��.,��ꆂk�D�"O�7�2 �F	5���P"OԽr��=Qi0�q숏_Lx:w"OxhY���[���8b���=���"O<U�#�ţy���*�F:DB�"O���� R�E�w�K �0��"O���E��"����a��.�y6"O�1Dݏ%�����ȯ(,*�"O��
�e�R��8�cY3�ܐC�"O��s�+����'�E���I�"O@4i�M�s%*��Y���֪��y̯�$
�NV����s.Ё�yrH;N�u��oF�5V� ��ơ�y2�
=R����g
�KRx��Y2�y��[$R �	|� �� ��Py��ެx�	�7Q+h$�q��C�<�����F�,�Rp�X����)�}�<���G�\X��(�3p�둣Bc�<uCC-2�{���)g)����J�<��o� ĝ;� �R�^��F%C�<A0���r����W	Ch��a�F�<�옹�z@p4l���L�Q�A�<1���g�h��i��E�V�S�<�!�ljJ�� B�	?A����.ZC�<�TG�!qE�@��;���A�<I��M�����N�g�������~�<��fĳu� ��B~��`u	z�<qD��s�"���/=9Ĝ�G��x�<Y4/^�2��@I�+��b�2��QHZv�<)�KW�*�¥	����X0Ёu�<9�$è":��¬_�^H\ek`�XG�<�gj_#�����  �d���a�W�<���,�tE��c?Gg��]R�<!���	_	�d��|欅Ђ�O�<���4.88�%�BC&��*�VI�<i���9wѾ岕�Y�E�*)I�#�z�<9Ra��}KZ���Ҥ�2�B��k� j@M]��Qh�h�+��B䉮B,����Ï.�\�wȹ���D0r(����Z�1F�X�A)Ub!��6�>��K�N'PL�Z!��<M<P�J�LZ��eȘ	q�!�d�+~d����ډ{6�{���W�!�$��FZ�pz �A�q�0�O�Kj!�D9*�Q��	"L�4�å�$WU!�� ��Y�'��漊��??^�0c"O�A��,C�\p��L�3Y^��2"O0�#�J^'�|���	?}-�yu"O�`��e�I�ժ�
�"O� ��$~�J-)fBP	3g.�Q�"O�=3����n^$�a�JpEvx�U"O��v2�j�3���&Pt��"O�}�ԩ�/]\���,�wL:��C"OLL�v^�/\�I,T%^?�"OJ��H�3��mz4�Ƞ�0���"O�S���4��yx'J�(s�
�0 "O�ɑ�!	�o�[��ڬ7�yi�"O@͐��S��d����)�Z)˲"O��rO�=*ѸQd��}}����"O8�S���ؠ���G~4��"Onq�UlԸF��|��I@��N�<��&_�li
)05EʗK����M�<I�Ŋ7z�K���0i���U�<&A�'a��kEC�<�&u�<���A�r�p��Ū�]Ψ��k J�<�Q&�*\��*�	l���fD�<��O	yn����뉃:�n����~�<Y׋�jJ������Z��u*f�|�<�`N9�$:��K�_�؉���C�<a6θ^U� �F�#C�|����B�<QWL0��)��쇦X>�Y8�J�<1E�;q.����!\�BdIF�X\�<�'(��`<��C�f6�9)&�B�<�C�	5�P�37dA���#�i�<)2n��+H���k�&p~�	��]A�<ٱ�X�b���_ S��B�^z�<��(N�_�Z����]|t� �z�<1�M߰*x���7�B-�8�Z��s�<�/ط!\5C3�Z�I9ڄ���l��1&I+?�q��`�Gˤ:z�hf�<Q!L�5"�&���y��܁U��V�<rfJ�mn.��.�3K�l��oKg�<����xXr�N�X�zLQÄ�y�<�bȉ��%� #:���*V(�TC�I��NQ��'ƶ@Tx�;��#[�!�$E�<���
��H!�4���׾g��}���|�@�(��dT"�25=b�%*D� ɀJ��|��X��)�)8��<r&�'D�p��]�"J���$Q�$D�Z �ª^��d*�K����#D�P(��SRly�1�6a��,��?D����X=��2���D6`��v�=D����Ą/.ٲ �.S'xFF�A:D�,Ɇ�R*���C�۹Z@0�+3l#D����$(K���J��'��icd�-D�8�P�V�#Ƥp�$�֭0Q�8D���I[&���Sa�4&�9�5D��ـ�O�z�����$V�^�I��&D��S$Ŏ,/�I�"�+���S�&D��*0#�6"��룏�A����/D��!K�BTq�閑p��x6�+D�@X�#7���;tI�	wi���A6D��c!�S�5�&I�tNQ��^A���5D� �n����J1��Y�n��P�5D���D69~D�/N� T�3t�1D��r��_�����%3�$��`�0D�d�v��?lh��W�W%Za�,�3�#D�H@1"�V1~5J�������#D��`���IԐth;5/��� D�� ����ȓ�H�0��@�
_(��"OL�óiہ\��1��H��F)��"O�a�ǆ
���7G�#�r1(�"O^�������2�w�ߏqѨ�� "O�a��,/(������F �%�m7D����e��7;�@�!�*u�!� D�0��W>����F�˧W�a2D�*D�4�p��%�<e:%���V�,銇�$D�X�@��5�T�Ơʥw��ZP�/D�L��FVc!~QE��<��P��/D���`O1+
xA��� `���Q�2D��	�hԬJ�ā�N�?n ��2D�������@���^�2`0" ���y��B#2B�@S�Q �]��³�yBi��i��Ĩ�
4N&�x�)L:�y�a��w�b9ۣB��|��P$���y��҉8=�!A7�M�s��ɠ�4�y"�� c��DX�Cȕp�đ��OC��yRK�S����e��eI<�2�З�yb ��R��5�����\5p%@����y��$��d#�o��)��ް�3�'r�\�`D�	u���A����x%4�+�'A��AY R�aEr;�'��X\H�P<�'iϜf�\	��'�\H�䙒yBVi��ZDz�'�d$�L�#t�i����V�"���'�����(�d�� J!�OwTU�
�'�`u��I�O���� !AQ����'F\0r��c�n��捝-���*�'Nl�ƆP�BG�"f#�T��R�'�DA�uڥdXܙ�$�e����'��6LɑBP��K��\V@��ʓ3` x2!.��T�MĒ
���ȓDiP�u��:K�"���eG�sV I�ȓd:R�! �V� ��
����[TNأn�cf�+�H�IP�͆ȓ��	bU$�� ED
d�Z�ȓY1�����x�Z�����
1��)�ȓzl��s�d��]��$��,�p�ȓ�X�Z5o&J�����&}�D�ȓDu0H�O�3ͼ�Y���?Y2�ȓj�^��0��lP�DJT;Qq�х�}"]X��gi4 �5.ޒP�%��q��@g'��Z�p����E�-��I�ȓX"��",�;$ �Iq���K~�L��	�Z�UJ���{�!�p�1�ȓb_��A���\=4#SG�K��9��9'��PѸI����2憚%�~|�ȓ�����ΑS��Y����*�@M��XC�=9�f*: ����O���(�ȓpMfMz!鎲i�qx'��*D��ȓ e��2/�W��و@ �v�0���w�, �H�u�JȘcO�R��P��tR8� �"ͶF"�<3A@H�E*���ȓe�^Dӣ�8-mf�t�̈J��(���X�8ªM�h
V�zp,��'x���ȓU��*���;R�2]s+ ;�.��ȓaR���� ;G��Q��3T�24��OO�!��K�ri��D�o�T4�ȓA���T-��|��T2~���	n<���<
��"�GϠc�T���]�F�h�Ѕ{� �7�	�[�����FӪ%կN�-��4QC�?�\���2�VC��Q_5�Y��a�K���S�? a��LR$eJc��4��x�V"O z@G'��h�Af�k��d� "O.͂���$N5��Xu��;%"O:<x.Z��t cc�|���A�"OX���#;Tl����tt���"O�E���C 6��᦬X�S\� +�"O0(cA(Æ`K����)���P�"O��`Y?S=�"�Sf�����"O��E�0~�utl�*S���E"O�E@�kP%"x��KS;kĶ�2�"O�ā���7�� �q�2�|��"O�����;~�C�d����U0w"O��:�$��gdYb�_�j��X��"Oy[��G�l)e-E4x��&"O\<y�l�9-+�)��fB,�sG"O�E�"�:D�4Q�d.wn=9�"O�8r �I�Rp)�%/�����"O�ɢ����k@xa�	�
���P�"O��@U�M52�� �U'T#
UR3"O0�per-�Ix��P��x�1"O���Dw)q��M�_Dl�W"O�-���<��Y��oL�?�ԍ�A"O�嘗���7�(��+dI�5�3"O���'BA�r�|�dNZ�8V½@�"O|������P��`s�u�Q"O�RP��S"m���X�[�t"O�U����B���={XhA�"OĢ��t�#dӼ;���"O}�I
5�F5����v'�Q0"O�1)�N$�����

�/�
$��"O�pËƊx�8	b�G�1��<
#"O�L鑍�(n�:ѡ�拁{�
�"OZ��eF��r��9�$��o�m��"O�Չ��Q'6`B�CZ6'%\�S�"O�xP@�)e|�q�,��3:���"O4��E�G>�X���+V���2A"Ol1 G(�3��5�f*C��<���"Oʨk5c��E �qcS)��L�v"O��0�\:$>Ai��=I����s"O4���O^7H	� ��nջ8����U"O�욥E`��X�@��-sy����"O\i�1n
�J7dP��&��L���`�"O�Q��A΂J�|���D�O�ZH�1"O���Q�@'J|�B�a�,���"O�D��f�JV|�����ꑃ�"O�L�əp�M��E,n�z�"O:hzR�~���rfG (��e"O��y�OۓQ���T! �cb"O:�@~�{�*B{�`�0q"O�Y0SL�R�2t���1I���"O��8@�3Cx�du�B�4-r�"O�A�A�Ƌn��a�'�A1e�XH��"O�|�"��%z���*Ъ$d�Y*�"O���ôj��(r���+WURaa2"O���l��0�tq�NY@� #b"ON-1�ī}�`!��cJ�u5�YD"Ob�&�ŵ��c$�D��"O��Z��%,�p�P�(u�xr�"OT�9��?A^�A@�߈4\e"O�(��1`�,�'�ˍFZÆ"O ��B�Kq�]J��پ���ӑ"O��Q��H�_������ R�^]s"Od�+�����B�,>ò��f"O�DPp(H/b+V���A\�Pd٠"O� X��a�ڥ?��� �!B.7�Xx"O����kGR�
l���:pIU"OL���:S{�Ř!�,�̜�!"O
�	�֞xD���Pz8L2W�yBi�	����f��~�������y��� 5�{���v4�X��yRd_&O@0FC<u,�V��h��'�z6oFI���(�"QIr!��'b9�E���@�'�EB���'�v�J㈎�4~�Sь�
@����
�'z8	 &�NM`	jPKP�7�|�
�'բq�cBP��ѡ�i��)n�x
�'%�(�G�2%�8ĨT�"���	�'��;�g0}"�04��E�Դ�	�'�J=YcI׶E�j��t������'}X!A�����aP�j_�颹K�'�Ԣ�M�p�$��2�ך\]Ld	�'2lyx3�Xin��+�&���0�')<��f��{,
�:�BC' �le`�'*F,AUfH�	�����,U!�'m�0G�ٶF��� ��)A�'݀�(�!�77�l�FL�`�`�+�'������
�r�����&
>����'�xڇ`]�+����U�řUl�)�'!���f���j)^�U�
�xLR�p
�'Z^�I�-J:W 
t�(ǔ}W�Q 
�'�~�U�hphГ�. 1Ti[�'HșC�i̧ �Ը��)Y�V��`�'"��q�����S-�926!#�'��-	����D0�C�h��w�4��'�4Pk�$�� �	�X��T;�'
���%`��8�
r�+@b֤P�'�2�p��ҕG�@(��E�6	����'7ў"~����� �x9��Jp�a�i�<9�O�mx��D\�^��i�oHj�<p�y���׋�Y�0���j�O�'nax"oE�I-�r��LāEl�s�<�"_-R�b@�D���b��PR%�X�<i�H�l���Q�RW�D�'�_�<�U�7E\f���ȉ(�`�6��E�'raxRJV���K̀�.F� ��
�'�V��" B��Lp����M���
�'p*  p� rb���ԉoRP�'tў"~��J�F0	2aP�(���@k�p�<�1�L�pA�D3���6��2��q�<����='��a ˥J85���V��`�?)f �H�H��@V�W�c��L�'s���ǄJ�<st

"y@�gk��Q1O��'�Q?��kO}P�a 0�Ό7�T��Op0��������s��ϵv���i�N<"�H��d'���	��J�
ĄE:����c߄.�2B�Ƀr��5�k��Xi��<&j���$aӖ�sWE�c��= $S��e���y�@��QQd�+��ةC��# @&�yB��-���8E��>�]�G�I��y�L�>b��(�#�/l�=�tߴ���O���O����/j��L�b�.P���s�'�ў"~RB̠!����� �����ԤE�<!��E�K�!��
�*������	H�	O��
�mޛ"<q�EA�h�}Z�g#�O��ɗ4Dd �d�V�_7J|෇� {!��qڐ��a��.�`�&�iX!��J�3Ĉ0q0OK(s'� ?!� �J\;A�qJ�!Qm�7>��g�� PDH�L�b�<yY�e��` V"Otp`/J� (�cM��7��y�U�$��	/L�4���
]B��;T%�3D6|��d�v}R�)��su���$pr�ST#�y�4���o������?~��>ь��Ӣ<��!���l�U���/W'!��&_\����
0��TYWMь
#�!�S�O[�`8p��@�4=(׆܂f��-`�'�0�	�.�r. �PG�Ӿ_�u

�'�a""@���i�#�lL�h�	�'K��+�7SuJ�j�H_2��䘉�D4<O0PR��)�����"}����"O|D����E\�8��HY�f�>)0"ODd�g̎�6�xth#�H�L��1�P�O;*4QaL٩e��CdA^H����'�a�!��D��#kM�:,x�'Lبe�&dp`Rc��6 ��#���~2H̝K<�郦��_6``�ӯ 7�y�@�/<�J&_�F
����<�hO7M%�~A9���81N�Pq'�c3Z�ȓ|$��P2n�b!�q�g	�/}r�=��U����|��5h�#��0XW.̟+@L�G�0D�D��c��I�0QbKN-wK��pJ.�d(�O�T�W�;wXH�X�#��G�e�!"O�|�Wm��|uP�w�K�n�r�#��$S7�0=9��Swc�8���Q;��g�@t(<��	��T����S'���'��xŖC�ɬQ�F�d��T�ʥ����O~�#>aO>�O~zw�[/;r8���Y֥Qw(m�<)�EZ�/7���@+��ya-Vi�If�'	�	�L�Ԙ������dk�l��f�n8D� ��L�� �K�g�wʴy&�3��*�hO�Ӽ>�l��.]�N�b�����v C�I7u��Pрo�Hi��߅JB�I�*J���V�;��y�4���Fb����ɝT�աB�u4�a�C��E�B�	�E	4UB6�tN�0�B�h�"<9���?�۲�M��p�gcZ�]��(H�,�O�OT4���A�:�}���K��pĨ��(�	}��9O�U1��ĖMSՎ�|wpEr1"OD��fV;(0T-ku+�,J���U"O^�H�뛋���iZlB�q���<����Ap��� �KJ2<��5!�B(I�JpBԁB�G���h���0�!�dȄ^�(m��*	5f�p�Űf��~�Y�$:g�V�t)|p�Udפ�(�jP�9�Is�����F��%`�`yi�NݞB�I)d�\�qV��
�(1�FM�Q9�B䉧S=��x�jԄP���Aj�.�hB��E�4qţO�Y��A਋�}y�B��a�!ѡ�YK�	tBdC�� �A�*��rɊtx��Ɏ+*xB�	,W�f4���'9Œ��e�]�L<:B�7F̠���osz1kT�]��B䉕]bnP2&�y��|r�Z .8B�ɳ!L��cU��,G��1�=gF��/?ɤF�35�T��׎�._>B	I4$F�<��S�Q�j���������B�<A%@U�Z��\a2	��-����%K~�<q����ám��z�r�Q�z�<�M����0Q26 &�8��wX�EyRoӡL�l�uX�$$�?�y�[/q���	a��U_9(e��yR� �)�B���b�
W���T*��y
� �K5
ګ`�2�)P�
*c�x��"O����ۨ+$U�V%K*Y�l�c�"O�hHa� 2C�\�\�\h�"��E��0=ɂ�[��1�E��횡aq�(<	�4cR^��W�
�x#j'�1c B����y��)e���y ��xlIp�-�� Ф�H�'����'��x~X�R�&"]���I��*B�%�8lZ^؞d���wl�d�KA�n�J`.�$IKy���>�I~�OY&�A���2�vTUG���6š�'�^�ea��=�ő�-��#�*��N��At����+��.<2��2��*�v�C c��h��MӰ-�y���X���#SBM�DR����y�aM1ay"�Y:G�|H�T�aҰ�8b/[��(O�������}���{�@͊Ĥτfz��P2g���H�Ɠe@p���C��A�X�Ҧ�Ѳ�hO�r�'P� �׀Dɤ�hS�#T�!�'k�����U1��	2���<	��~���%z��g�Ǿh����fM:��$��B�h1$�-~� ą<_6&����I�I��0�ݓ�hيc4�B�>�E��n��*�&Y���B�	(m���`��0��x�p�8
\�B�I�z�MZ�ˌ�:���B@fJ#�rB�ɭ�섁��N20\t�n�tgF�d<�S�Ov�41�bU
���s�R��P0Z�"O ���O	�Y�� ڪy޽��Q����	�,��Ty�:r�x"��3
B�I)nx���c�� :fQռA�B䉆T����#W
�>({��TW�C�	4!8�Ka�@�|��]��NT�E��C䉎O�lk �ڢb�`�*$Å�H�C�	3ag"�ċ
�x��V�{��B�I�0�tŸ3c�8�Jacd,Ԯqo�B�	d����aj��(�z��#�Әsk~B�ɣM<L�Al̍��P����6+pB���1��i޴��#��̵uzNB�I(c�~\����k�4`p�%V�NB䉪���	tN��T�,�ФEF�B�I
2̾�H��(.��e�dB�"-�B�	��8��F�R61���Q��ř�zB���AElìt�����RB䉴a[����,H�j�j�ˡ�T�9��C�2lQ��u��9�~�җj.^ĶC�	� �0i8MM�f���B%?o�C䉝1(�d�C��3Ub͈�A�"u��B�I�{��0���*-��d�#j�_�B��9w�R��� �RfpX�Zq����	�'^0�!�C\���yrC
5��0�	�'�Q�%<_|v��aC�)�1*	�'f�D��eQ�'��A�kg&U:�'�6���)"E�bp�7u����'����a@�\箌�FW�.��A�'s���$��G� xyf�ֲ�<]�	�'2�h"��ŐF�9@��ņex�		�'�Y:`eB�1Y (�Q�_�����'�fp���cI���W!�Qeh,��'LBH�%�����*7�Ca4��'��`�D�[���e��o�e��'.8J�� ��ɋ��5PU�M��'����7"�8M|H����_:<P�'�<��o,x�c�F�7G�湀�F�B|�)\;eM�}i�F�4�%��W*u�
�'_`���n�Lyp,��C�:�!�'Τ��a��
_^��k�L�1�	��� �Yå�
6t�����{���"O�$��eR=  hY�	�
{E�qJD"O���um��W��Rp�9Wd�"OH���/�2�����(Cj4���"OlX��e�,TD4Q�1���i{�u[4"O�0`��Nw�DI
�eU�Az���"O���tu�`�Dv}n�q�"O�ES�AZW(lš��Mg����"O�U��Ƅ�r��Y`�OY�m�l�"O���� ǕZ�\Y*1�>9����a"O��K��D:E��� R�\�K�0�y�m�+S��`R�h�R�B��V��y�c�&C$��͢b5�]�J��y�'A-�R�/��d���a��W��y2�6xd�J�%H3��v�Q7�yb�Х9v,�;W�S�V׮�jF,ȱ�y� �NHlq�b�/T�6))����y���  �qZ%AK{�pӄ�	��y�	��<V"�x4	�O\ja ��7�yB��6��<x���3n1�dS�ű�y�ʵ0p!��t�|�#�M�y�eE�~["��mA�kF�l�R��+�y�%�,���-�6ԅ�Ha���
�'T�A����%7��04+�+2��,�
�'����wl݄T	�q	
��g	<9
�'���B��˓[9��#6`��	�'=j\�3F�Y�mH4śr��-��'����Po��������t�Y��'��z�`O>8Q<A�`��
��݇ʓ%��:r�	ESl�z�NȀ~oL���U>`�Dfê�88�u'հ�� �ȓ1���↋�$^��(�^�Ą5�ȓyTtt4[�?�8�M�7`u��~�& 	��T�S�h��#ݲkU��ȓ��Qd�V-*g�́D�Cy���ȓO^� �g_�.��M����v�ȩ�ȓ!w�ɳ�d[��V��v��'~�.��ȓ 8��`'D"x�6�I���?)\ą�6����݃)�Z���I,3������yj�g�U�ʘap�T-($���%�֑�F�)3��9�`�p_�-��&�6٢���w?�� c� &��y�ȓ!Z�E8!�qBQpe��Qz%�ȓh���Vl �Z�����]l��ȓ��`E���5c��G4@�Q�ȓB�-�ʈ�n��*�ɋ�M��m�ȓq�M��͢;��٪�H %����1�L��K5-����C�?D
�$��[�gX�{~�y�c�$5��J�i�:D.rX��+�p?�&��<\X0�)`�Ȩ���1n�Kb_��xBG�03%��I�E=,T��vnѲ܈O� ;Fĕ4�`����͎*5��U�$�T9bFCE0�y��Ԭ~��x��ϝ�d�	5a��yB+�n�ȡ���\���";���-'�~P���U��C�4Z���jߚ~���aD$P=[�,�4�$̓�"y����˃-�%@��B�>�(S�@�aa~r�
�5Q \� ��*]� ��*ɜu�x<���W�/�P��{��VnT����4:$�ybT��E�'�6�Y�-ݫ���}�� ��FJ|��@��c����B�<9�E�2m�h݉�$�v1ڡ ��<�fK֟=�:�p�+7}���G5t�J'CC�A$-����`!�7:od�ʂ�a�$�"�l��S���z��U�5����xrF����=�ԩ�o���v��p?��"��;7v�Ha�P6Y b1�2�M+=���)@j�
��x
� ��q��$>�p9�Ĝ2(E\@ ��+q� ����)\4Dzd�q���j(��;@��.�!��Tk�B���.��R��&`�!���b�<�2a�&1
ܲD���!�R�GNP4��S;V2��0�g�!�5-� D
��,�$��t��f �O�h9��&븧�O�^�"N�$c r���^k0�-��'�Uz�l��ޜ$*RK6�m*v�|B��}:���yRh��4m�2�@Р�#|�B�!
�~�����!g܀hPL��u�4AQ�G�(�e��,�	���Q��Wns�:=�p�c���~���Dx¯�7�4�(��,qp��� 5�iO)n��P��tA�$(UF�-�!�d�B����B��T[�|مC�|k2�th

+���u�ɔX?n(˧��  dȜHK��.�t�PW	*D����37�8��c�yN8�sE�	(� C#��2SNK=+����ϨO&=��A���x ��NݎBLq���'���x�A�,!�&�ۈdI�-�1	%:�v�4`�/���^R؟�!�#P<bI@�Y=p��ԘK5��4v��`�!(~��]�x�O�Ҳ��,�")�Mϊ0�qb�<�Hx�8�p�����Zb�^� ��7�en�, �/ܮ$gyD��' :�	ҫ��f�u肯ޅ.�y[�'��հ�l�(}���� *�97��ǹiԔuY�Hm bGF�:�?�q�"�JѹǬ��;ɪ��G�y��,��l�x�愓a���-8��
G�O�� gȔ=Y(Eˢ�ܯq��0��Ɏs���EeS"�IS�b�+<��#<q��U:�����"�L|���E���&�ҥ��۶n�
x) (E�!�� ��ZPcV;3ޝ�P!��
$A@�ϯ0b�3������� �@S�O��.�[� �٦ ����/�.A�!��k+��C�½��!V���j���❐>><�+�b��%A��O)�Ez�%�+$PP��s���,1��8��=��/�6�С+�e�+%1���%�X�>��6�<__��GC�]�����3�ON��q.�%K�,}x6&�.Z���D*����3J��M�P�%*W�Z����cvj�3tEXY�c_S��	"O�����Va��-��cv�����t�A��]2z$���V_���D��;�tla�qبe��|f܂�"O����^���qp���=b�8*��H�}�����c��у ��6A��G�`�'��\�OW	nY�3GA1Ox�	ߓcs�)�� ���T��",D}C�5(4�y��
�FB:0���Tc3���z�h8*RC��to4�󐆓��tBcS���X�0��|��aMg�$C��* �Y(�I�N�
�aU�y��2kfh���k�y��� : �$��!�<-r��m�*�>����'Ԁ��ŏ�S�N�0fG�,h�̕��'��M#�ϳ[�&�#PW�k�b�PH�D'���k���ҁ�'�\)rrWt�Z�`@��_�L�0�3eHHOV� �(1b��;�h_*H���4e/�8����5b�RTe�7ʪ��T(�2�;Ӧ^�FP�c>YH�Aʁ �8-CpgW�n���"D�lXQ��3��)cD��I�d��ﮟ���O%���`ҕ>E������I�I�!�0i�ViD�B��$�v�{�+�n�L�@C$l�'߰�p"� N,Є�	�:�M���x�\\� ^4�p��d��f�,�6��at��*��{�*�aVC�:B&$�'���Z����@�ʥ�&+�&XhN�����T���t-�S���Y�F��|��P�Q��owB�IT�����xk�D�@�λ49�˓6�2�"�)�'~#X���BZ�:�n��L�1��ȓ?�d!��E<a�i�$�3^N��ȓ �� ��1cbH��@�B��a$D��( I�]:� F�X03oJ�#3a"D��s�N�7���* T�e�~Yqp�/D�X�UL���N!�P�X.4�X5"+D��!dMEJM�go�/"%��I,D���V�5Yl��ʜ8��1�-D�h;���2'ߠ���I&Sw���u�)D�� ��SG�U�-#0�C�S�Dt @"O����c�u�Z\@���M;~����'<iIw�EX��H�RqE�#�7⑋��1lO���=p����+2���cfg�M��MݽXSʓlO��Ie��t��y���)ђ@�/K>uJ�,Yrg)��'E�8�Cj�?k�I%>7n���Hs���`S�)ՠ�	U"`����IIf��'�a��ϣjX�:Ac�$�4���s@�,�I�P�C7%��!ԣ�K~��g�=B@���Rˮ���G�/z3Eb�1D�(�T	ܗ {̸ӧ��g������L��y��;{`<�[�O ����r��T$>7�w�HZ.�*Lij" �0𑞌���;s�$C�,	q���	��4 I�^�(С��
���qӎ����΄u4xP��uay�h�i؄��@T,�
,
��ЪA����^Ub`, �i9���#AT�@'>%"���D������ף�Vy�ցH�{���A��84�~C�5&�4�p��.+d���*f�x3�.��e\�@����Ol:İ"�ȴ%�8�P���D�	���������Rf=�j�	 � ��zR [u��b`�� ��*@(��v��<�*��$���VU�A��k��<�q�j��<�q-ԅ6�x!�5.Y�".��r�g��e��G�h�"����I-q�&� �\�Z~�	KZ�&�zpmߞ
�ڸA� S�o�!�#<�d�eH�5U���m�>8�J)���@�[�D{ I�ې�KTc�'%����;׈}�"�Q�y���c��U�-В<��5��!�\�%�8�3��֫{��IPa#��5�	���8'�`���<O�}��ڡ^p��B��Z{�Bt�v�'q�j�NZ��TX��ܥo@y�I��x��*��>��1��T�[�!��!�n9�4�@��}ZUC!i��'�mr5CR#l�V(B���M%d�P�A�,[p��2�Tyc�mN�Z�!�D-[�X��C�C�+���Z�����,T(<B��ADK1s/\��e��%?�Kǫt:"�����%V��k�!�eh<q��R	'`x��p鍙V�r�w��8, �H�Ɔ����	h��|�r]�Ó����A�:�VtRR/�"�Ʌ�I��\h�OK�y���p��;2��Q+�9.�vY �o���|Ӫ]e<	e��?1��`���(B�|�"�Z�C�v�H����V*P�C�h�k\���|�w���ą[�bҦ��}J��z�<q��[�r�y4D�n���ȏ�D���ICK��6�^�p��P���O�)����ɕ�Id0�`�"Oxy:�)�F_Vh��eQ�=?x}��W�a�Nl)d%�jV���p<�R��G��`(��˩5z���`�_���K�e��^|)0��{xl�mX�p��sH��,���S9ѡ��D�7P�a��F���0��Q"YqOHA����/ ��9��}��b?��MH�:�����4�9��(D�`9q�=\h��p&0��9���˖���Նe!�(	����|�'[�4�H�3|���S�W%[�|a�'��T��.7�R$�"T����4��ʥ�Z�Ph���1<OVxP� �8MD�cʓW'���#�'Q��"A��P)8,@��׫g����%L�^5���ʻ�y�X�~��i��>G�Z�ÀM���HO.@T?�h�V���6	r��D�D;�����"O^��\:0 ��s׀��1�	rt"O\�(�\73:��� �B��J��"O�x�7숦^{�U8cMޫItJ��"O�i�e�<z�B=�`���X�n|C"O���!��iε0�B
	�=�A"O��r��Ŏ^�2��a�#;�T��"O��*�E_#�؄�gɜm-6�"u"O����A��9�!^(�ڱ"O��@E�΀Vs�������-qB"Oȅ�cB�{A�}q*������V"O�`�'$�Cs� !7I��z@hI�$"OF9�E�0�~� ��#,L0�W"O�$�  �tL�!�V���yR&"Ob���7S~�x�Aϖl���"Of�ң�\��H<�O�����&"O<� )�(=���UN�;{�xY"On�`&W�p�԰�4�4
��q)"O�)C��+l�Āq���I�ja G"O� ڜ�O2BxVQ;��S�d���"O��Z�'��4��\K��B+v��Kd"OB�I��3ԍzr�R�Y1�HJ�)D�@��>Z�T�c	�h�iBN3D���3�?P����V�s|�c1D�l�]"hɘF,ݝ1~P�Ũ1D��Y��������C �kZ��pe1D�������;P��gZmJ�)D��R-�U�޽��!C2t� e;'&D����R�t)������{v&$D�8��ᐷD��4kw�*B�(��
&D�L��e�pAJ�J��;C�����2D������n c�Ή(#$9a��2D�l����y��y�&�V�Lբ��0D��ۑ	���Y9��_P�j,D�<�&.�#�ڈ딧UD*��K+D�����ݐ$P��Y��
e�p	1TB&D��pJ�q�V���BS�
�X���$D���JR�V�Q��!E��XQ M.D�� 1hS-f�:��G��(Nq̜�W�,D���%��E�^(��Ѵ7<@��#O&D�Tx� Z�4��)���"P��;D�܁ơ]$`2l��3	ɡ"����Uc7D��	��H�x4s�EGl��h� 4D��0�-O�E��}pdH�*:1��5D�ǈ�U�N�A���(�����7D� An�#_C^X�犅CL���p�2D��	D)L�?W2�x�(à<��P���$D��#1a�[8a0A��AՀh �h?D���J^W��L��枔s-vr;D��Z%��,<k�� �\�Ht��SG*D�<ң'�,.���Ђ^�$�&���,/D�0`n�V�u�ٶg��XXW�.D���3jÛg|!�� c�|ps/D�\�`�U�GW  �kB3:@��p�)D��5� ��@ ��|%���`i'D�4�5N�	�&tk3�Y��X@�&D��i�,�:�bL�)�h��|�&D�|3Є�| ��#���]|���,1D�|� ��9Hr���
	+� ����#D�Pp��>VS�t!�d��c|Z�Q�:D�̘�d�1D�$ bVl֏�n-҃@*D�$���͛B����o��s�B혷,=D�x��EO�9�N�8��v���b�%/D�����Yf���>B�2���!D����_&6<�L*�##z��aȆ�3D�t�����|`g"΍,ن�PR
-D�0��H���x�HU�[o\A�cB(D����Z2!�z��T#D~Jc�#D���P�ݫ�⠪�o�9k�"�`�!D���a,�3�xt�2�R+=�x�"��?D�$ Sf�-I��li�h§iK*�Y�8�Q�Nђ\�ϓx�IR I�Pk��#�A;X�����$��g����(��M=A�PY�ʚ 1�>���/�v�+� �[�=)���r�X�F|�咏u���2KTcܧgYh�2֍֯Y�N1��c���6��ȓNF6Ei&.� F�sœ�oB�5ϓg�.-0 !�>tT8ӧ���zg�A&c����B������"O$���C�B��ђ�mȲ:���k�����Uړcy6����'{��X��BV�LU�o� F��`z�JW>�[���;z�8ೡ�^�%$��!I 8ɡ��z��9�,\!�Fd�6���ZW���3O߀4�����iY�x0���A��p�^�`E!nN!�D��q�����"\��pX&W�d �d���(	������)�g�? JM�1�1~�����������"O<��BM�\(|�`#$	�@)Ó��� ����%ҕB��'P�����O��Tqa
B+iˮ� �+6�U�'�ڍL���ʞ�rA���z�Հ	�'���9&�<��L��L*QA��O1(������i �d��5A"7�����#�y�ʞ1؀�R�i�_��B"��y2e��x���)�F��g�p	����y��P.4,�@^+ ��3�ʅ8�y� �xA4�K8[�QbԄӱ��q�����i�"r.�M���
`�s���_!���rb��9�@�9�|�5% �@:n�O�t�e�@�B81�1O4U�taΦb�p�y��D�_�����'lt	��
L�8A�ȎSC(��mB�(2JdR&	�<-���!%�'�T����SѦ$Z#A�+;�B�@������U8+��e	��j�S�X�0!hr�J3�ʠRIY�0rjB�	�訵C��ل�\�"D���Z��n����Y�p�Ȗ*H��+p�%�g?�@$~آ��A��r���4IV\�<qG�\:7ƙ�%�W�������_�u�̭S�a;Yxn� �M�
���3���������G����*(|Oz0Y���]���X�䊀%E����'�t��E�Ж88�a���?ᕩ� ��l�w儖]n�٥$�v�6���6�ҥ8��p��.��������\hѪ�z�䄯���"O�;��)-v� �EF�Y^p��ϺF����'�	A]j����N�>�I��Q�Gɰ
+�d:��"�VB�	�R�N������v����	�j�$nZ)R�j4(pn�{4 ����O�di��]�� Dk�-ݠM٘H6�'����mI�g��`y��:9��1��[�^�����>�D���i�r�a~�,%��R�1X��w�f������LPՖ���c�O���COJ2�ʧa�na+���c�d$��ꝿb�J��ȓȰ� ���V�nP��y��-(�̋�a��qE� tPm��ڃ�Q>)̻9� �1���<3m��� ̛R�p��%�z�� �1!H�u��Ǖ ��R��	��8C"��&{\a!@`��?��`�	�^��!�W�"¤IY�懶Ǵ���&afX�ѬK�_��]9�$�1m Z�����Uk\��@�@FZ)��B��ΰ>i���{1�A�7�sn��E��g��q��Q�$@��.�f@�V��D�� 0�˾~zA��[��sB!_(�ƙ;C#�E�<!��٬�0 *���2�䙺V
��pȈ��1N�! -�#��m���	��ټ�Q`J�B���
��?X܀тE
y�<q7�U�dX&�����%&��1�
r)H�I�e�l��DB�����`��ӛf^��H���3��P A�S	r�c�*|O8�!� 9��@����,+gE��*=S�@ ��\���f��>�(4��3Zdh��2�)e�ѰD�"Ex�(\% c���b�P�Qa�j��`���9b�j�T� A���#nԎs�@B�I�&C�����Y��nq$a� gZ�`䉮[�Mc�	V�EBbF�%����VgXh�e#�
���/!D�����܆r�F��CC�_�:d�E�!}b���]� 
C�����Nՠq�!�,i�:�O^ԋ�bC?Mb� q��ӯpӖ�"'LJ�-�����H�x���j�s�ǅ;%W��{�oW4��O�$����8avR�C��di�ɴu�N���X��!cD��y�bK ?"����վb\hy�#[��~2��&2��@��KS��EAr,��Eoe�AJ"��,NC�ɼ5��`�`�
^��Bv��l�'�|q%�65*І�ɒ@�peâ�W�gz���d+d#��$YDMu�����LRpiC��ǆlp���MЍ!�`���'�4U
 `�g�� ZF��E><����� J)��'0��{7�3�F�l����T!LB�	�%h��� bF"a�r����K�L����ڥ*$�)�'2u�}��������w�˼A�Э��m�FL�g�٘Z�~0r�nA?�n��ȓ�4����چ��IŅ#��C�Ɇ3Ä��K��
�6� N�;��B�U��H8p���E�:%�#r��B�)� ��@0G�}^ ڱnY��(H�"O*%Xf���h�A�n��8��M��"O�	Fʀ&%��$�M�c#�I�4"Oz1�BB��5ꈹ+c�ժ,yD��"O�����8&&��p�,{V���"O(ywMO.?lX	wlL;A�%jg�'������QX������Pp1��%U�� 9��#lO4���&E�	�DB�-��&Q'j����Dۮ�e�L��!"F�f�yrGZ�~Ȕ�p���;�,)z�Z���'��0͚�8�6�'>7�hӨȩ�I�� ��4���12J����oC�cf |�'�`�l�<Sr8��"o	x1��J�"�j�#M�,1da�.E'���Ǫ�g~R(b��
���!d,r!,I�p����=D����$ϞjT�y��|�|����+ZN��6E��Kh���O����8J0��$>7���3�|�uʐ�!��{�FI!��zB�H,� �"(��<�A��`���J;`�Y�P�l}� �Y�-뗍��<����;7�4pt`�;x$ℳv�d�t�qۀ�Sn��搋�ᝦ<���K�6+? 9Fj�1z��r�'K�!�$NJ����@��M)~��0>|���~	�ax�Y���3� $���;����@Oφ<��t��B��j�� ��[���(��/9� �[�n�[!�!�emN�zv�c.�|̓y~�#NB|�'�`�����$x���[�B��7`���<~O\�Y1�FL?�q�28����	
=N=N�y��]f�<�!Z�;����%�9u�|}!�Y�/^3�"���u�A�Ӱ$�Q�$���]�6qY"h�	�����o!2=�ȓ[vpj�ᔏ|ݜ�0͒z;xQ�ȓ�(Ԫ1͎Fz@��\)F�^͇ȓI~`m��D[��h=bD�ˢ@��=��;jj��D@Դӎ����#zBЕ��y-��d֞U�JC`טxl$���R;�l���� t��)c��?	AD5�ȓ?(`�1�(­y��:�E�4x�p��ȓK�>�	�#��i�Lh��gD35_Du�ȓ-0� Z0M!T�L��0���T>�ʓ��Qb�ݞi�T����l*�B�*3�LA���QƬ`��S&sj@B�ɓI���-�
y��٥ �<a4B�	�?ת<�2bݺ#0�ͺ6�$a��C�IlKD�@�K'޵kt�>x��B�,g=�iBv��X����Ɵ0-�`B�I�W)�RL��Y�J�E]
c@B�I
	�>q�'�J�n:"]K'.۫2�ZB�	�x�r�X'/��9DV�8B��T�s���~A4 p�hT�	52C�Ik6P�5KR��%n�:N�C�
V*)Hro�f� �e�VVB�	/��m�mО7�#)�(t�PC�2y��� d2"�� iGEMcj@B�I1r��Ju�ޒLhz�q�I�M�C�#uS��e�B�u| @��x��B�IU���Z��ծ2�$��Ү-.�B�	�j,9*�M��T�p�KC�tR�B�9" Ze�̬zRLt��ˣ^bBC�Ƀk�xM"��8�X�,D��I�a7D�;ٲ!7�Tز��=P՞	�J2D�(��L�j�J���K�|�D���2D�l�ql(�6���o�/G[^��S�7D�l!-ɽ{I����J�>�P�J3D�́�"!G�*S�˦R��z��.D��S��T�5S��p%�6 �"�2�e)D�ԣG���,1��1��Y*ͻ�'D��r'D���p�ʄO^3CRd��.D���1��9&D��0
\�r)n(��G,D���fIL'�U�e�]�yE��B6I-D�� �l����z	Kr��wPZ|zP"O�X׫�!��D�֋��:��}�"OP�
Qʉ�H޺�񇉛&�&p�@"Oμ�!g�(X5���QF��F�Y �"O�l
�'؊;�.@�b CZ���'"�M����8C`,���oj�qv&��G��q2�'&* sL�*J�DJu�
�b`���'�\�+�`��!	Dr���!%�r��'�Lu1gX<�	�0���&D���'ǖ�b�)-2a30�B�Y�؀�'p2|X��N���ht��Dg����'�X����H*n�ṃ�խmn���'�p�x�ӇZ2A[��ݓ��`��'!Pp�A�Ro�|�AA� X6�!�'��e�2��mЁ��ں�zMH�'��5����-�\DHb���^�p@�'�\ӴdͯN���A�eH�]@���'�M�j�O't�{�͓2U��9��'~����I��޼`�f�� 9w�ِ�'�b�Q�o�_��@F�1\�.��yR�_�\�,��=�|b�.�~|�Q�-�iɔ��"�l~���Ґ-�I>��ɐ=KL���@�G��� [2���D�[�usT[�D:t/�O>7-H�B 8��nފ�U87I�*Lw��`H�'���S1C@<
�$Z����@̧ngJ�Y�K�3��2-I�\��f��%�=3�oӤ��+��O҉OL�U�m,<C�V�61\là��a�\�l`��0�O��Ŋ��PW0(�QÇ�a���b/<?���O�^ª	`��/��ͣ�@3#��9hLi�ԋ���əy��IsjS$^��S�O��%�����<ո�)c�Q�i~j<�4$Tqۇ�Z�8d.8�ȟ䍰�ň�t2�%�r%�#�9�Ac��K_�̗'����FM>�"UIؗ��4*�%D^�4�iЪ���� lz��Ї+�0|r���=W�L@T��W7�p��H�<�1�Z�V"���@X�:�6�
�\O�<����g���d*�Kd����I�<yw�`�i�r`��B{�z�F�_�<����$nT681�^�bWl9��R�<�5�S�W�t�[B-˹x��qJG�_Q�<鲫�I�4�WJְF��{���r�<�q,�T�p��EF�,@ ��@�Rc�<�ț&a�0�Hv��5�=i�Z�<YOV-C��ň3K��B�˔[�<�T,G�WDɺ�K�@��iFZ�<Ia탇vD��"��5�ƕ��W�<y��-ê���OB#��Yx�m�U�<Q�C�*+d��1��!-��A��M�<i���Wk^��0F�}�%�k�H�<q��A�L�����푨��6�A�<a�C��n ����-�A��y�<ѡJ�%����D��`�0�Ф�y�<�r��c�i��B+n��А0��<�����F���k�㏧L���	S`�<y��Z�$M�={!�����D�_�<�ů̳.|��r��!.ξæÐX�<	A�C5Y��  ��q�v�˓L*D�D�#h7c� (h�䉈v(ݓ�d3D���ՁL��)�+�a�  Q�,D����@�a�S$&����&D���N87�l#��#S�$[�:D�`�s�٘���@��,7�����;D�DaQJÅygZj��&��qGk:D�0A�U.2���N30o4uE�3D�0��V�����I�bi�S-1D���-�86�V<�sD�6�0���*D�Pp��؍n��䆃��@�q�(D�<��+�F�x�S��4/�l��&D�� �x�Q%����J��mb֘ʰ"Onѓ1�?��A��)
%�ܲ�"O��a�M��QK	� *�d4�`"O�y;R+�ic،�j�#��U	D"O�(�#F�� ���K'	B��ۡ"OԀ����#i�D�6-D *.��6"O�Q��DN����I0��*��"O�{&��8Y�d����_@�|G"Ox�CR�
�%Z���'>�5�"O�� ���O��03����٦"O8IS����E�$0����6�ڹ��"O	���0;
��vI�9GFF���"O�5�,^�2W�Y�3��*.�"O�x�2�=���I	!�́c"O��y�C�>�򠺆�9����"O���ք3$�JQAf����"O��Iek�>.���%&	�`�F��"OX�� h�&�ֆ�+'�vEZF"Od����&�>��a�l�d=�"OxM���ҙAt����S��)�V"OP��!�M)3�6��!ć!h��Z�"O\Ara(�/`,h��Xs�(t�"O�Axc#����41�E�r�yp�"O��H�`�#uT4�%�s`8 V"O�9�����P0�Y�r�I�@G���e"O2ppԣPG0�Z(Ɠ0?\ �"O&y�S�z���5$\52(�9�"Opx�r剿p'��
sB�WC��"6"O�����_G,˵�O#>Ej��v"O��0K^4x�B�2� ��c��P!"O����ч���˒A  c�2Ԡu"ON��i�:s)&��&���yP"ON��T.ޮ]�z�y�e4b����5"O|	ңG!W|��Ę#=�.]c"O@ey�ǂ~H@��Ӣ�'�!C�'��h�a)�L8���5��lZ�'P$S$I�#�����!�9e�XP#�'�l����r���dά��	�'�ly����档��J�U���2�'�6q�r��}|ꐈ5�B(dJ��q�'�&(�S!BS>�s�7�B�'�p�1p�z���/R3y���0�'[�%�DkЬ#x��$�n�*š�'C�(�6��o���ALW��y��'<�d�P��2�%`�#.�'d\LG�>�A��A�)&=*h)�'Z�S�� gy�������h�
�'(^D27���DP�E+!���	�'9ZP�dm\�Y�����"�	E8݆�&z�	j��\()C �M3fU��Ud�(�SLp ��T-�(m_�Ԇ�jh��ʐ*��4� E��F&N삕��v��i3�*�z���[�%�LE"��ȓFG�����/�����h�
����K����.nf�<;T�I�i0 �ȓk��B� *�}��_*LJ8Ņ�_�H�̒�O)ab�A��.�0��ȓ	�x���͆,}��0"�aF�<ˌ��&]�0���2ҮѱsdP+sڞ`�ȓQ�Y!L�<P�����Ѫjz���ȓa����o�7��Q9���3_�d��<���'_��-a`�D
k�j��<�^;��_L ؠT�G�CJ1��Hu�Xp��*n�:pxs��)Tx��S�? �x�!\0\A:ƪB&���""O�$����X��I/��.h��H�"Ob0r��5?��pz�m΍:Vɧ*O����UG�Y�!
<B�E��'��Y���^.]� (%�#�N���'<�p���*H��е�=t~x�'�b�hRFL,hu�� �,ʜ��'����F��U�M���Ny�����'�x�qOGX%��ŭ��i ��8�'D�x*A�wB���4��]���'"0�ұ��9���@�n��e�l	�'���ʰk�q�ހ3�MB��<��'o�%�7Z�?�(�fE w�`��'��q�e(!3�D���쐩a�$#	�'$���6~��[f�
�J�XL��'
^�hё*I&�C��E
t��'z�
��3t��Q&��)f]X�'�:-��O?Š`{��V�3��%k�'��5bG��)�@i���%!HN� �'����NmT��DCM' ׼)�
�'��܋���)2|:I�u�e�

�'[���Di$�|2�h� p��	�'0��$b�M�L��S�b��'(�u�˞m��Q����J�b(x�'2�S��ހ-)���Ё�����'V钤�֎]^+cLH�:�и
�'�0��!h�F�6�5��?����
�'��˗�&����d��5"��x
�'o����T4_и������t��'Ȇ��v��&;ܜE:��Dm�����'�ؚ�	�%wg���`�3_S�l�'�����l�?)�4���oљ $>=*	�'�P�ВeUp��_��qO���y��T�_�@�s�Ԉ!�t�!ԃ�3�y�d��D�`@1b�){�M�TGV��y�m����@Hg�nr�Q����yB�U��y�ːG<���Į�yB��	ZB�2�)F��N�h�	H �yB�՞F@���Եs�`I;�y"+�"�����aK�nb$0���y�"����u���Ղ�+C��yrHE;�l�͝=�(��ER��y���@�2�� ���>㴨�y���^H���l��q$n�2�y�.6����n֘b�T��� Ì�y�O]�i���Цͻ\�4Zr)���y"�E)JH,1�P-�ZG^	"�	?�y�k�2��p�d&=��)�&π�y��P>R�B���&�8C	`��m]�yr/6=ߊQaog�B��f��yW�Z�>ys��>p�� ��H�yR/��|����Bl���;�΂�y",�*�N���"Vhk��Be���y2�X�� Y5�+^��Q�f��y��p%"�ـL�0]�@�C�'�y�Q������3'8�i��B��y`��Y�ȋ�/T�$[*��y2�Z&Q��k��4F8���Ώ�y2i�#S��q�g
�˅L.�
�{�'LNY��
s~H�!�_�,��)��'h�$F�(�X0��H,�f+�'�Jaj�N^�P2��[�hA 
�Y
�'F�Q˵M�d��פ�MnD��'�J��$�'yJ�J7�D>��QA��� ����)*��l;���#!���"O�d�å�_PhS��� z8 3"Ov��$��o'Z��w�Dt9��k&"OfI�*F3s�����y �a��"O�3!Nǩ�Π�����X�b|c"Oqxt�=��!Ӧ�?\m���"O>5KE���S���7��`e���7"ON��0j�*S���
 �ݝ\4�+�"O�̙�D��|�Xȑ%9K�tK"O�񊄮�%���sDN�D9I��"O������^�k��<7^�j�"O:U� ��� �bhC�	"Nx"�"O��b�G��%���  �q�}�"Oz�鳍�[����nŎbT�҆"O�ۄm�R�Ƥ�D�U>t�"O(�H��ظAZ�Ks����a�0 D�p�#ަDe�q#7��u�0L@��#D��00��%��lڤ� ����!D���u�T!0��a���|��U`�O?D�$Qo�@�ʍ�vپtoZ`���<D�@� �	~����'�X�8(���A=D�8�r$J�.e(Y�!�x�21K�<D�<9�)��+M*�TPC���8D�80�!ν,&��g�tϘ�B��4D�@���>~܂9�v�:p]Vp�4D���f�ݠ5@nD��)!'$��-3D���C� r�Z���#~����<D�\P�%L�ryN��mN�) b��1�7D���6Ȉ�Dt�d���*4v"M��;D�<	E�#*x�=ї�V�^E���,D�H�� ��|��D�  ��g�8(��%>D�@	��D?Cv��#�
�\Y���&D�����A2/>Å$[10#�I�dn&D�$��]�;��7�ć_�p�!D�l[��   ��   �  N  �  �  *  H5  �@  L  �W  �b  on  �y  ?�  ɉ  ,�  [�  ��  �  0�  t�  ź  L�  ��   �  ��  �  u�  ��  �  H�  ��  , � 8 2 � �% �, 4 4< �C �I >P JT  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(՘xb�'��O��(⃯"T�����Y3s��eX@"O�-Q3�&&���PFi�&��{W"Oݪo�����XsmF%b�N1��"O�����?l-�pp����k�j�w�"4�L���%U�\�5�Շ<`u!r�!D�����7D=b}�����z@Bm���:D�878B�lq�ɣ%�6o�!��޴%��q���T�D��=��@خ�!�ā%"�na���̥a�A�Ve#�!�X%0��I�3bZ�8u [�6V��}B��ȹ�V��T�S�&����pb:D��1�)\��j�;�lֱx�v���A$�B��?���ӽmTm����X�P���!D�Rl��A�65I�`^0�P,�bƪ>�������B��a�B 	�+��B�	�x���s��q�i�5@T%,BB�)� �}�Q/nI��x2�ݡ ��B��'��'��P��:Ar ��b�-7�\P
�'+(qh���NEV���럢^ti�'?�<�̚
<��$��+F��l	�'� ���J/&���*Ł�1�T�i a%�S��?�«D�5`L�����+Z�d�{�<� �׷,0��0��i ��#�AN�<���׵Y0$�o�a4:�Gtx��Fx�#���I2
�+�`��c�щ�y� :8�8� $ݧ
�z�2#��1�y�n�5"�T�e�ʄ�ba2أ�y�'�BH]��M�>/� ���yr�&^}�M�4�$m��{F���yr+��9=�㭍;kw�rJ�s�!�Ĕ�>Hr���FЉKg��*�DK�!������	*8�r��`+ �!�$��U�@ᆖ�<ڰ�um�r|!��� �4�r�I88�N�-^4F�!��Wdf�H�/ƶ����l��#!�$�*�L%��dԁzh2�¥�t!�ߺW�Y  %�ox(���=2Q!�dϞMj'螁(n�|8��):!��]���l�7�ӏ4��WM߰!��ٛD�6���V� ��*��
�!�ÁOn�X��U�v�����B\)g�!����)�"��i���V�!�d�>H�0XQ#��j��9��OU%I�!�GX�b����ڬm����W�/x�!�^a�@plTR��6ޞ�� "O ��0�	��D�a��Ա>r��W"O�t�3'P,s겱�aIA"��]�""O��A�`�7 R(iUOL5p��!�P"OF���H�<p�1�ED(G��q�2"O"p0"��I�B� C$���3c"O�<I׮�f������9#L�6"OlŢ4e�!"�`K0MS
K0�Y�"O^ Ct�Wk�LۧkS�Jwl�xF"OF0���S5C=�(��oO���"O�����U�L����?>8��"O�����p�<	
%��i6�X�"OxxVD��xt4ahƈ��qs"O64�ǆ�JW*<2Ӧ��]ߚ��"O�m���)Gp�P���o򠹘g"O:4Zg�&<�����
)l���"O��h��O0(|�1aԎR�P1
P"O,�%���r�jƟEY����"Ot@��@� �XR��6K��b�"O<���cU
�^ �1o�?q3���"O�Q$��
W�Q��n۷
�8�`�"O�TD�� ��U�r�3ŚhX�"Oh4�c	 l�Ƽ�k�!��ѐD"Oyx�3���;G`�F@8�;�"O2�q4��7�nb������1"O�	���8~�Ȁ9&-��4��L� "O�����9G0:PA%:��(�"O���Մ_�x�Z� DA��b����g"O�Z�k	a�l���ӼF���*6"O�J���;hfB�!/ݯ6%J�A"O&M)v�1X����͐;��"Od�b@���?@����R��@�'"O����(p�hF�V�6��g"O����)B�a�F擌���"O"��C�čC��}ل�ע_�,��t"O�q�aaW�{�������$���"O� �EQ��šV4���ɪ�l�SU"O�Dr%�8�*ȫE�7%��Ȳ�"O� Yg
W���H��L�8 "O�k��=YYxDC͜&�4���"O���/_���쩀�!$����'zr�'Y�'F��'�B�'���'t*�y��Ջ6��Y	A��{Ĕ����'Z��'��'(��'"��'�R�'T�A���I�6|p\q�+� Q���E�'��'�B�'���'J��'[��'�l�0ҡM3���y ���Vڨ���'��'I2�';r�'�B�'\b�'����ܮcM��:�eQ~�)���'��'%��'�r�';��'t�'��%�T.W/Al�Z֢�&��¶�'���'6��'���'W��'�'�� ��g���Pd���h%�d:��'E2�'��'��'��'/B�'Kؠ����Z=�U��V�R<�a�'�'���'��'+��'CB�'�X,W��������Z=p��)�?���?y���?1���?����?!���?3�ۡW�A�%R:S�TqZI� ���O��$�O����Of���O���O�׀(�x��Ӆ�2@'���6/�z�H�d�Ob�d�O8�d�O�D�O��d�O\���ư���޿?g����D!^;����O��D�O>�$�O��D�O���O��$Y8�H�ŝ�.����8'�d�O&�d�O����O���O�mǟ�I�.��Q���T:]+�,��k�N��*Ov�D�<�|�'l�7���pm����lʉg�f]#PC����Ŗ�L�޴�����'��aԘa�z��4̀�U��P����$O\��'t��K�i��I�|*0�OU�'N�"\�g��:�����F�(+5���<������>ڧ���hWC:o8�d��@"m�y#�i�2A�yB�I���]7r��-ٌ���h͡xlhu�I؟�̓���I{C*7m~�ȹG�ׯ`�6�8G�U�U/f`���a���s��bFf���4�'�a�d16�@m���-h�
�'w�	B��MK��d�n����G|T	Zc�F!R���m�>����?�')�I�O� �,aRҤJ��!0��?�7ɞ�J> |�|�'��O"|���%�@�N@�0��y�Dρ0�R*O���?E��'�����*X���,� j��es�'��6�&?���Mی�O,L!���
i������*^%ز�'���'��P�8�&��Χ��������8h���dh:��_�r��&�����'���'��'V�qQ�@0Z0Je�7��0&Ҩ��R�'9��9S��j�'`R�'δ�T>�I�[�Q� �4x-{`
۶V�fd�-O��`Ӻc��I���$�U�T���_�A����h,=X<Q���q����
?���R�e�'9���]���,��	+������A e�3ʔ?+��I����Iڟ$�i>5�'XV6-� # ����N�S6��4�@���IW�V��dI����?Y�^����4}�&�'�\�+�ǆ�(yB�����F��=�����n�f��<�6K�W��d�~zT��2�*ft���ЙOfJ��@&�/g�d�Ol�d�O0���O�$6���Hpj F�`�tq����Yͪ��I某���?���Ky� d�ؒO�`���B�(��$sH���Wb)�妵���|j�0�Mk�O�``��+��Bo���s��
�J�V$��+�t�)ћ�R����	Ɵ0Vjj0:��R�i`�	��ޟ`��oy�e�O� ���'���'o��7 �A�C�O�D����&>`�R��	��Mc��i�ɧ�	��~��0�/��zNer7Mݕeh	r�R���X	��>^w��d�I�/��i��Z�P�p+�Y!�f�25�fɺm矨�IޟH�I�b>��'��6-��%�-�s,R���e`�y�m1!��<y'�i-�O��'a�6m˵tB�Ó�șn�P��o��]�Mo�ɟ�X�BP���'#�ˢ�L�?ݦ���q嬂4�P�R���H�&Qs�o�ۦY�'���'���'��'���gb��s��#�U����:�$��2Қ��	ğ`��\�s�������$��C��Pa	�|�z�"բɉN�i,1O�O*����i`�d�=p5y�a�++��,I *ƳJ"��!s�Zy�IQ0�I"�M[-O�I�O :��}�B��k�R�,�{"��O����O��<9�i.�����'���'8p��í�*~X�麦���3�LP���K}�i�0YoG�I	Rۈ����$�>��w	ӛM�B�K |��̊1:�@��O�]�e^B�ɟ��E��2!Z1�a� � �w�������(��̟hF�D�'�޽y`�Y�l��=`%$����_�?qC�i��iT�x)ߴ���yg���pDaϪ{F��{'��~��'~��'k��(��iH�	�m@��A�OP�6Jƞ}�H��[Vj�	��Leybn����|R��?���?)��EI`��2f�?cO��+G*r�tɃ-O�Ul��TP����@�Is�s���v��*��1o�8���W��$�̦��ٴ��ŞN=b4���U�O_\u�0O�e�80�Z�&�pI�Oh�r�#������Y�8��4���	>

�8V�O41_���f���	La|��e��Ԉ�D�O��AW�<��$X��z��5=O�=l�F�� �I�t��������@;q]>9넁I01=�%�Wצ�mv~��\��5�'��ܿ� �U�ē�;/<���A����@:O>��D�	 یhqB."(�V�2R��ʓ�?i�'u�M�O(d7�4���2�IfNñkp���WI(t�%'������S�K��9n�M~oY�cV&a�,�nR�CK�&}vLI3���T�Q�|RW����䟔��ԟ�[t��58i"�"��ҍb�'����	cy"�j�8�27O�D�OV˧~	��X��$e�k�@�9x���'���iy��a�@e%��d*����k]�0��� ��s��s�"P9ZM���'kA~�O��L�	;�'�.�ك&�3'O���GY�.:8a�'Sb�'|B�OG剿�M#G%��%��F�UF�ڼ��ܨ�K*O�n�M�@��	��Mf��!q@�.�؀1vŊ-u����4p��:A���h�É��M��4�~¤eԈC*�	��J/O��@���<�/O>�D�O~��O����O�˧j��I3�H���j�'	5HmИ#��i��9�1�'n��'���y�l����<t�S`�˸y��� b+�>w�%m���M��x�����|3��8O�1Z�
7�L@�g��b�إ�U>OڠЦJ� �?��=��<ͧ�?� o�o��pF*V�
�H�8���?����?������u�w�LMy��'�)�Ǉ�^�pi82Eތ������'|�'g���?�ݴ-��'r@h�@@��5J<xn�+��(Q�'+2�Į�\��P	�����쟒�x�%m��DZ�|R@���A���Y��Q�{f�$�OP�$�OT��!�'�?�b)��tl��f(۟G�,��	^�?�i��}��X����4���y�%K�s�k@ˠr� {w��
�V�	��Mu�i��7��e,�64?Q�n���)�9*Q2iX#���p�#���75d�ūJ>,O�I�O�$�O����O=�P��)���E�@�Y�����@�<��i��ŻV_�p�IS��xqU��oDv�� C�z�6T��/��$�O���:����F�>Ia� �
�ՉB���Jw�L��'GX��-�e?II>�.O���P��.?��y�"�Q�[�聚U��Of���O��d�O�)�<���i���#��'���{���w^���&片9CЈh��'�7�+�	<��D�O����OزeZ�y�H
$l۱.`@�$���7�'?������L���)@ J++4ʌ�+��@�����w������@�	Пp�I����z�o_�2	�8��K��=6!7l���?1��?B�i$*�Z�Og��vӔ�O��
�����I(_16D��D�=�$�O�4���-tӎ�Ӻ{���!j���i`h:�q�qMY=%��'��'�����|�I��D��(M�6x��K�a���P��8n��@�I���'�7�AL���OJ�D�|z+Z1 -E��b߷'�(�A�ŗU~�>A���?H>�O�.1Ac�(H�K�,�*1�8 ��(�L��i���|"u"��4'�� v�z�:A,�^�W���S_@���ݟ,�	�x�)�Smy�As�TY��`D�xDH���vTR��]0yN���O�XmO��P\��۟Ċ�adU�Ux��6y��i���R̟l�I*3�o�a~Zw;�ip�՟$˓Cgt�ڗaХh�ℊƁ���͓���O�d�O����O��|Rrc��Z͚�`R��$|�(qX3��=m��e�H��'b2����'��6=P��͊��ˇ(:m�d9��O��0��i/v�6-c�<�ヌ.q^�p�P4^��
ak�4��ᕋG��<�D�<	���?9�e^4���*�憢b!d��U��9�?Q��?����d�����Ug�����ޟ��0d��Ak.�3�"N�`�bb�D�{�2���ɟ(��J�ɴK��űC��2��#w�Q�6�0��'�� ��GQLF�6f3�)΢�~"�'פ�hvC�8"���)݇AjЉ1��'"�'�r�'��>��:2���e?�����D٢
�P,����M�Mѓ���ߦ��?ͻS-��2�'"oV������\�q̓�?!���?)���M#�O�}0alB�7,�<Rfѱ��Ş��P��^7��O���|"���?����?��8;��������R	S&S�8 S+O�nc�0��'B����'<�!j�M��<М��á��=p8�Jŭ�<i��M��|J~�2[�xs,��A���YNޑ!#�G��1�6G j~F8�.9��T<�'��ɓE;:��I��'K���&N�
��Ğ�����ҟ� J��v�@�� /uм:��n�8ߴ��'����?9���'��n��K�J,|ݸW)� //P�Rs�i��ɥhF���ҟN����� [�b�6��*0����	?\��O��O����O���9�|�&���(/� u���X���!�'��byӲY��=�����mK��S�,��+(>u �ؠ!�T� M>1���Mϧ�N�ܴ�����7
� �P/ё)ĀQ�Ǚ?qK.1�`�?�Bl1���<Q���?)���?IfƋ�?dL@$�Fqq���׾�?a���HѦj��˟h����ȕO& �ӷ'��g�d�rwOG�T����O��'�b�'ɧ��Z:T�u"�0m�>�%�Ok���!AeΚ&�~�Ɲ��5H���g�I�	��z��:��J�~�J�з�'���'�"���O��	��M+���2��C�~$$��U�^u�ux���?���i<�O��'=���34�8���p���U#�6�h7��ަ� VA����'0���k�?9��W�� f<R0V0	VY�#J9m��	��>Oh��?����?I���?i����iE�18(3�'0(~5 ��/<94�m5	�`��'l����'�j7=����PՐ�
�V��$�O�d9��ӽ/�v6�n�p�]�+嶨��@�/C"��ݕE[�u��'��'��I� �	�~��g/�+6�ؐ���D�$���쟠��ʟX�'�@7E :}\���O��ѱG���")(Ʋe�2�ֻ\�X)�O��O��O�\���E�F�Bػak�a��"������֤~� mZ���'L����ޟ(�p�N
	�5�îճX���ө�埈�	���IޟG���'���� *�}6`��熠
.$i ��'�7�3v����O��o�d�Ӽ��삌?u,E���- ��ʄ�<���?�'v�9ߴ����:���N�?�9��]�PP���u����T�@M�]yB�'���'j��'(��1a���q� �(z�(���e��	��M;6_�?���?!H~Γ`B�+��5+	~D�V-ЀH_��
�T�X�	�H&�b>��Ǥ�\cv�3���9z�+�⟴B�R�l��D_� ����'��'��ɸ����Q _$��$A�D߱$*��	ٟ��	՟4�i>��'e�7��'4����XH���'��˲�Hw`�Dq���@⦹�?!7X�d��ҟ��:��,ѡ��}�����B; �rH��oOߦI�'�A��{�K~B�;��ۇ�
<�a ���7�2,��?���?����?!����O8­�	=o>��0��D"����S���I��Mk�$�_��M�֓O�̒�$C2�V���!�#)):���l�	㟴lz>�е�e�'@f9{H̱+���0BKŁ�@,�����<�	
#��'��i>��Iן����e��9���-��)1��gA���I��<�'*7��L���O��$�|*S�Ce�L��ǫT$�r1��R~���>��i�H6-j�)�5�j�xSs��0\��RI2 p�	�,Q�׊�����(,��Q�I |�@kfmӏ�"�	WI�b������4�Iڟ��)�Wyo�ܼ(1P�<2����J�: �R 
��I�M;��O�>�&�i2ļ1�gʟ��#3�p9�)�''l��HmZ�)�hl�i~G�
6���T���>��Y��ZK���Eb��o���<y���?���?����?�-������9�4͠`���K�^i�r��Ϧ��3$u�X���%?���M�;b�Q�mV<-Vd�
�7:�ҩ ��i��7mK�)�ӽ>��9mZ�<q5*It�$[�A�'}��B^�<yG�20���ϰ����4���� �Z\�RdՋ#�~̀�!X���D�O$��O�ʓ�f��y��'eBaęV<f$�0A:u��l:R)ޜ9�O���'�d6m����K<y�qS��s�a��Y��@��F~�bçm^��1ŉ&��Ou�%�I%.n2,�6ag�Ѹ��lc�p�qV����'>��'����L�FH�S����J�@��)uk�֟��ߴu�8��'��7�/�i��aãYYdLD�� �"rO�����h�ԛݴw��|�BI� i��C�6���C�f4���1 �����@
)S`8�6c�	����4���D�O ���O���Z�JW�Q�p�@7���^�˓_c�F�@6�yB�'�����'[�����Fp�I�f
<���+�>�r�iA�7m�g�)�Ө{V�CE� s���@u�N$U�T�Q6�24^j�K�����l�O��L>�*Oաև�"D+�����&W&�8�a��O��d�O(�$�O�i�<)�ii2����'F@��J��4xS�u,	�G�'Y�65�I.���Oj���O��T��9���q���B9�r6>?A�J�t0��q�����j�c�t�V�`5b�^f�a�|�,��ǟ`��ԟ��	ڟ���b��t���V\۪�FeM��?i���?a�i����O�b�v��Op��*Ҫg:.�����DK|���b7���O��4��%��u���Ӻ/*3R��&�35�I�C�j[)��{?�K>�)O����O���ORa@V�@�����҆`�A�O,��<���i�"9 Y����q������$�WB�/CA�#�<���x}��'�r�|ʟ��ː�уZ�,�H��D�h�,ZFbL�;�|����z�^����T�TM?1I>ѣ�ζ~p�p�	�0 򮒃�?9���?����?�|*O�@o�>�J=�����*j���GՃ]T�P��ry"�z�⟈��O��d��8���3��4���:G��e�f���O�FbӦ�ӺC�MS���R������9Ҩ�t�ڲB(��щq�̕'���'r�'���'`哗=�v*�[�{�4l�a�!"&8�	ٴ5��pk��?y���'�?1��yGjWRBR���@�[-T�	1�N�~�"�'�ɧ�O��9�i���O^R��"ɘ+-�X�要�!��D������'�'��	Ey���e��Б�U�MU�6���axBeqӲ��)�<��x���t�ك ��&.^=>��E��ɽ>����?�6�x2���kl�23��<������$
	Py��	UM~�hm%?��C�O$�ء0����ņqu��+�p�����O&�D�O��;�'�?��J@�`pD�&��,\A�� ���?�iʾ)�U��0�4���yW "���c�b�;.����L
��y��'�2�j��S�&h���`W����?� ��RO��,��DY0�41�%�7�d�<����?I��?���?1&�H-�CW$3�:�w���$�ǟ��̿<����O�� yc��h��P� ���c����'�>��iR�6�UU�)�S�����na�3R#m�p�&�#��'J���%NΟ���|2^�p�c�ؿBp@0���dLjaA�"N��(�	ҟ�	ǟ�ry2Cr���)�Op%֥�u���Q3��?6ˠ��%�O��m[�L|�I��M�3�i��6M҄-xf�!�cM����t�M�j5��hD�n���4�Јu!Ꟗ�I~��;O6� �&�9���s�:\�4͓�?	��?Q��?�����O��m�	�-Q�*m�@@�6?(�6�'���'3�6��%֮˓)��V�|��F�#V�Y�� �4��g�hO�Xm��Mϧ*/�ߴ���t�C1kW 7�|W�4J��ӢD<�?yp�$���<)��?���?��g�]�I"F�P��$8���?q����Ċɦ51�*�ʟ0�	럸�O����2GV�o{��j�D�i�*�p�O6��'�,6M�֦ŁM<�Oas"L´
�fLhV��y����waP�'s4��!iE��i>I��'�'���'��1Ή��lQ��x-0������	ܟ��	ʟb>}�'��6m����X(b��"uD勷*({f��@#��O|�������?q�_���ɵ09�ͪ��^�D� ���'��I,�Mk��F��M��OfQ�r����d]��A��KD��c��,�rpY�m��'yR�'m��'��'H�Ӎv�(yu�TpϤ��`��G
b��49%��Z���?A�����<!R��y�v�:HZ!)#R찪���@x��c�(�%�����g�zӴ�I�+����^�e�Z���EɈ�F�	
J7�iPV�'N��$�l����',��VhV���"veY�g ( Rq�'�r�'sQ�@J��6�ݕ'*�]/&�l0���11D�����O�8�'u�6M����@H<Q��C ���#GQ'�83��n~C,$b�9@�b~j�O@���~!���#Xl��*sc$T��yj��S.���'��'8��S�h��^`���NXEZX�qnȟ�9ߴY�(Щ��?iv�is�O�N�/�ne�Ǎ7����!�j����Q۴Aj��&�MV�v��R�%����T �p��(�d'lk���g^:Rh��%��'z��'���'���'���Iץ 5�8Y�j����Y���شP���?������?!��M�<�r���
�Ie��2��Iꟼo�*��S�Sz�l���- )4PC����������;��'�
 ْ,R՟��v�|�\�t:�J;;�U��37F� ���T�	֟��	ǟ�~y��g�Ȩy��OF��t)X�I�x�E!޺	J��p1OZ\o�T��f��Iԟ�������4hJ�0�����E�����f��pn�A~b 8���Pܧؿ{��[72ʨB��Lw���I��<)���?Y���?���?я�dH�&x-ʳ�Y���>�b�'w�z� Pstð<�$�i3�'�N�bc�� Sb5�w�+&ӈ�A�|r�'S�O�HIq��i��	�S���z� ���da� �	d ���(�OVf��iy�O{��'�BA� �����կ	4�ݠW���$r�'~�	)�M㓎@��?���?�,�P�0'Ìe+��4A�Dz�P;`���;�O"��O:�O�S!?Сɲ���P�ʽ:aȑ�6}L����L4?ͧ2%�Ę(��Z���y��£e�jXR � S�,����?)���?��Ş��P�Yh�i�0[z���tF�xA$��$�'��7�+�	���	���2��&jCj�P'�K�<�E!�CP5�M�d�iU�e��i��I%k�j�p��O(�;>����ºj@v�� � +���͓���O���Or�D�Od�$�|rcI��U�ʠ�c�L�t�q鎥/̛���p��'?R���'�:7=�9) �Cw<);��Յ$�X�{�6-�ѦiZN<�|2��6�M��'�x�(Y1K�0�4g�;T�h�+�'��屄� ��C5�|�Y��̟�ӁNz¼	҄+Ӏ7�D��u�Y��������Hy��u�4M����OB���OZ �df�-\x�+��1]��ps#�$��,��dB�q��4Ɖ'�����M2x�$I��iG.xd��O^Irs�����h4�	H��?�4��Or
��V�竃M�<q���O���OF���O�}��EHD�bØ7�y�2��8b����7l��lϮOY剿�Mk��wc��SKW�W�����_&o��s�'uv7��Ѧ��ߴ#AdĻٴ��$޿���{��K|M��kB�%Z��fɃ�@�n�P�1���<�'�?���?A���?��M�;.朱��H(wjԀ�M_,����yw ����	ԟD%?�	�N$b-j��4_���uI9[��O`�l��Mw�x��Tm� r/:�gC	;�8hhw�8��k������d%|p 8)��n�O&ʓ%Gnڳ��5A#��S!��US|\���?���?���|*OJ��I�)֒�� T��KQ̊=�U&�<����˦A�?1QR�p޴\��6�b���v
�L��B�D֔O[r���*m�|6�5?鑊K�=|���1���q���ثkH�0b�G�2��8��c�����$�	��@�	� �Z�GF
	�H��!ʊg�t�Y%���d�O�n�=�2�kh��|�#�.zit��h�q�`�' ;0OX�lڋ�Mϧ  Y�4��dG�0� (ҤoEo���� �F�"�3�A!�?Q�)9�D�<�'�?����?1a��8�,XsTf��J ��ӈP9�?	����d���)�C\����I�ܕOs(x0
�X�� B�h�5DL�tz�O�(�'�2�'��O�)�Ob����As�}B��Ym,��tC,,ح��-{�z]�'x�t]M?�N>q� M)u�	Q���^Y�%b�E��?���?����?�|�,O�\m�<b�Ԉ��Ȇ+-b�As��?1Z�J�m�IyrHl��㟜A�O��D� F���R�EX�d����7����brC�֦m�'}v�r�Gm2.O E���KQ���5*K�s��	��2O���?��?i���?A���Ɋ	3���u��>|?�M������m��f�L��I�(�	T��������d���(Y�d"�a�-T��I�K�$�?��C���OL)�1�i��7: �`z�e�x��V�{��D�]p,��'��':�	����0�ipC�Y]?�cY�l�����ʟ�����ؕ'h6��4 ����O���87y.� �d�>X���i �����X1�O��d�O��%�h`o��5:�L��h�M�!�2?�v�ٴj�^8�ܴkI�OΆ���?�㳲XE[�RǄ�"�l�.Ґ���O.�D�O�+ڧ�?ٖ�+ ��σ�0]V)cS.ũ�?�!�i$$�PV��ߴ���y��(k������={��T�I��y��'���nӞ�JD�k�"�=v~Q���?� E�G1ndJU&Cr��Q��_�	Gy��'�b�'R��'1�5�*�#��Lj�E8" �I��M�Qo��$�Oz���D�X��A�`�ž6��
�S�$I�'��7���QzM<�|"%e�*l���R�j>����(5��*4�S@~"�	?Qt���iA�|2W����iٹDb�91��7kl`��Qş��Iӟ��	ʟ�tyҍq�p��Ԩ�O*t�g�57����ԡȊqt���9OvqoZw��-��I����Iğ �a���&�=:R �
Lx�];� ̽[�QmZk~R�@0�hL�Kܧÿ[#F*tlL �!ꉍVh>��ej��<I��?��?1��?����h՞|֑�^^��3�˺���'��v�@��Dc�<��io�'�Z�HQ��D^~_�25��	a��'�2���4a�<?����d{0��6N�.8�7�G���%�pjR�{D�%��'�zp$�8�����'S��'$�m����Hf�4Ut�a9��'�2Y���4%>�S��?�����յO���de�0�b�+I�6�����D�O���0��?Q
#��)�h;"���m��Сo��0b���䌅�#�V��|:�i�O$��H>y ěA�>�q��%h�B=�ը��?����?����?�|J.O|`l������
 �XmY #|02'�Myr+`ӂ�\Y�OX�D3=�Z�IG��&g��[o?Qd�$�O$ЊU�v�n�nr�"�韂�O�����Tx~�cB�vPT��'���ɟ��I���Iӟ��IQ���"7
Q9#,h�آn$a�7��;c�B�d�O���>�9O�oz��J�Q=���k�k�b�Ȣ4��ܟ��I{�)�#I�@o��<�aDV�S�J`mٝ1������X�<)uj�!ל�$I��䓎�4�B�d�=�\@�*�{��Ir@F�:j���Of���O�˓(M���@��I����˜�Xr��Z�-�93, �����j��5���8��x��
[وl�ȃ] �����������;'.� :��|�7��O��R�eA�<B�H* "��gč�l%�Lr��?!��?���h��\��p]S��D?k�nɡƏݸ+���DP㟸�Č�O����Ҧ%�?ͻ'���r��&`"���&єUj��w[�dӶ�m� 6p�lZ~��)�K����ƋEɚ�+�69�p�c�>�䓛�4�`���O�$�O���.s�=2p��"[$����K;1�����_8�?��?����e�W�򩘐$����hC6�/e�2�D��k�v&�b>u���h� ���2,ЩQ�։o�f��An.?�S#�-�j������d&G����v�*��d��c\ �P˓�?���?ͧ��$���R����R�� c�8HW`��@�AA�|��c�4��'��e��He��DmZ�$4��M����0�C#|Кݱ�j�˦��'��b�e��?��~��*oB��D�H�-�N4�w^1_і����4�Iڟ���㟜���Oa$�Sţ	:.�^qJ�m�>�P�O��$��݈�a9?!P�i��'�V�X�U��<�)Y/u\x8�L5�$�����|"�i���M��O����n�>-�@i�J�sF| �n�{�`����f�Ol��|2���?���[��)R�o��:�H��ql]�$��1����?�*O� o�h��Iԟ��IP����>rR����7X�\��h����d�g}�@`�r�oZ���S��ܓ{���٥+K,�xw癡EU�m�&ײM��ł�O�)	��?�A)���B^�p��ڔZ��q)e�A�x���O���O6���<��i���'fa	<�@E	3�8�ȵ��qa�	;�Ms��@�>�W�i�аRpC�w��J���3T����@m�~`ne+�nZH~��w����Z���((�X���͙8���1�TN��D�<���?I��?��?Q,�v0B�/4N�j�'|\�m��N���K���ȟ������$?�����Mϻ}c"Y�3
ͻxvཙ�i��
!���?�O>�|�E ��M{��� ���al�M1�܀�e�"f��'8O� ���~b�|2V���џ��c�d�&���"I�v�n�y �՟���ҟ���Sy�ir�N-p���O����O4x���W��5��j51H"�ɛ����O��d6��D�b�f�:�&��QD���K�V8��mU�"��Lͦ�qK~JT�������L�7��;�|�#��#ڴ��ğ��	� �	V�Ou��ݜ|V�5��һD3���R&�
0��u��i���O��D�����?ͻfp���&͕8e<YZR�޸��̓�?���?����M�O�n�8��S�"�h�	���!mT�P�L�LNl�$�̔'5b�'���'��'<�ԈR%��$D�M8�S��̸uQ����4<V������?�����O*�ȓ��G-pp���S�{����>i��?�N>�|Z��b좬�����a�p�Ы�5�<�B�4V��I�^�=���O��O�t�ġ�m�F0,9��Pj����?9��?Q��|/O֬o�^=����w14����/Cd���H��gF]���MÍb�>���?���-r�H�5ћ=$t5J[�vռ�� A��MC�O�U�a����4����w��E�2m�?"O0�Ex��'���'���'�B�'a��ܰH��?5֥GI�|�0p��o�O����O�lon:���'F6-/���a�`�"�T�H�D���K�AG�)'���4J��O��|���i���:dJ��6.�i�݋#%`�P���ũj�!o�iy��'���'�Ң�o��ucv�`�d	U���'��	��M[SK���?���?I,�^���PSZ	�1+ؐ �`�[�4A�O�o��M�Вxʟ�EhȽ#�:p rN�%<t�H�УѾ�܅I���%�P��|bVf�O��K>����X`���W�K+�^r�!��?����?	���?�|Z(O̔l��W@e �!�0g���w�N(S��H˦!TGyR	~�D��ѯO�lo�*A��$�8"t)�O�7:8�Pk�4	U�&d��
,�֒�P�Rآ2�$OMey�A9]>I��Ŋ�x���%_��y�U����ڟ���ڟ��	�ĕOK
A+�d@�h�2mC�/�Ř��{�x����Ox���O����d����s�����y�b=H��
'w�¸)���M�|J~����M3�'��m�婜�&j ���[`�'��=`�� ϟl��|�T�D�I�\yӭP�j���c��zj��'�şX��џD�Imyr�q�n��"h�Od�D�O\8��G�K�Ub笏,&�*�%���������ܴ<_�'�*D��E�r�:��ǻ1h���O�u�C�ó464��逳�?Y��O�=i��g?dQ�G��%pX˖l�O����O����O�}λ6f21�v�ϛV�����V�{^�
��tMR ,�?!��Fl��4��H����|�H�d�M�z$��8O��m��M33�i�R����i��ɘ!AH`�A�O��-)�aǓb�R�3C��20@�av�R�IKy�O��'m2�'���a�$�	1�_�x����ߨN � �Ms5@܀����Ol��B��аL{��BP)޾� fOJ�)��$�'��7͉��i�J<�|�@+��%%<��N� mFZ�dC�4G��QBQ@~bȆ@u���� ��'p�	�Cf$�5��uRJa���H����	ܟ��	֟<�i>-�'i 6�ǰmR���R�,;�d<(p6a1�e�-jl�$\��?	�\���ڴ����i��ٚ�@R� 	|ȓ�'Բ^DY{��6x�7�)?9emG"�2��*��ߙ(��EҸ�y��� Hsތ�V�p�t��ȟ���ȟp�	��`�z�&�L ��c�I��,A!�7�?����?�!�i���O�R�s�d�O~t��`-_X(q�` �)8�)q��g���M������cI�������4��0�����x�\Y��R=i�B�Ǫ��0:�|�Z��ǟ��	����q���k�ᘩ0�^��#Zǟ���ty��t�j����O��D�O�ʧ_&	� **JH�t���]n�@�'�*ʓ�?�ش�ɧ�i�O���hI�	���h� �,�P1`G��f�8P���S�72�s�	�c:�0��>�<�5�ĳE
���͟���`�)�Soy�s�L��C�k(�3�	l��	��t�Q>���DM}��'��ԃM[��h��Xx�"X��mT��,�I5ކam�U~�`ӂ'-�l��g���uP1g�@�{�>�K@�$���<����?I��?����?�-�4��Q'�fH8`qԪϘS���@�hEͦŲ�+�ǟ��IПl$?�I+�M�;q`��2ǁ�p�b�`�;e�XL���?)O>�|"!��<�M��'I,բ�F��L���#�-e���'m4H���Hߟ�R֑|�Q���ߟԛD�חɖ��Ƌ�3�|aQ�����������	Uy��o������O����O����_�MvʬX����b%��� ��OD}�'�R�'��'�NI땈%Hz��f 8La���O��ґM�5�4,���)���?鑍�O.M�Ҍ�--4Ѐ�`ؼ]��u F�O����O����OZ�}���:J�	IB�R:�ؤrfD��m��9��f$�T��I%�MË�w��*�D�Wؼ���+p�DÛ'���'��G�.��&���+e�
�2��t�Ъ v��t�_�z��H�Ĝ�1��&�蔧�T�'���'Y��'0�����?->ɂB�1��J�P�<��40��ؘ���?�����<�B��� �^�A�@"�wh_>�	����y�)��'��� &U�v�G%[��M����9 Eqr�]k�	�sj,L���'� �$�P�'�xxH��H8 C���-T�֠��'Q��'-"����V�p`�4}�<����v!�hX�Æo�r��dn�)���ΓS2����N}��'3��'!.�y�O�i��qB�ʞ�:�T��oj��V���jPdRm�T����4H�+V�`Ğ1���]0<I9O`���O�d�OB��*�F�I�]�T���}ϲ!QP,P��O�d�ƦaӢ��Jy��g�ГORh��)YZQXe�T�#��)7�%���Od�4�Rt:aAz�����gQ�A9֔�щ��:�I��Y|�$L)����4�"���O.�Ѷ��@�� �T�*�YƌL�G�>���O�˓*��6���y��'�V>9;V �"����B��A�\�!w�5?�U��0�4Gś�(�?m����1�����Y:][0YF�\�}�Սo���|����O�%BO>A$$��ժU.�H�(�3���?Q��?��?�|�-OralZ={�,]��V1*�9�(X6dT�F�2?1Ծi��O̜�'�7���k��h0��@�{��ٴ%�M4��l��MK�
�M��O�l��B���L?���GV(�������g瘝f�n���'��{���D��`γsr䱔V"�J6-S�	���?���Bw��Ε�gb��1�E^{�Q{�IP���D�OZ�O1��)��z� �	�@l�@���q\�@p���%X�z�ɴ�*���O��O�˓�?���}����%�h��)��;cO�%���?I��?�.OPlZ�3� ������I��bu�e*��:�R��	�3r� ��?q�^�t��֟�'��s`�1v\@ � v � +9?��.
z��PBA�c�'s����#�?ATd�z���iD(-J.�}YE��?���?���?)��I�O6���n��#t��:��-�Z�H�O6o�H���==�&�4�AxՃ�>}����qD&]�t��g5O��o��MK��iP�Z�iz���L�4]��O�z� w7�b@�BLS�sŸ���H��Qy�O_��'db�' ����|�� i��'A���q7 ��'�?�M��%��<1��?AN~Γs"@���t��| �K�3t\h8�R���4 ��6�+��:rTp5���d�vPHc�'9�X�PD�	=O&�����'��|%���'�z`�����1� �Z�[�A�b�'7��'iR����W�`aܴ��m�S�2�򰭂?#�V�ӥI!�F�Γ{ћv���v}�gsӔ9nZ+�M�egV6k�.#��1qR�(F�,�I��4�����2�<���'̸O����3A�����3܎�S�oI=�y��'�2�'�b�'����FN����+D�r�1a�B����?	�'��x�O�H71�_�w�zL�A��{��:b(���$� �ݴX8��O�x`1��i����f��"B�?ı� �ܪK�hu�!p�BA�Y��`yb�'�"�'�R�O�0� ���S4p:hc��Ϝz���'�剖�M;r���?I��?	+����&�%]��0�N�#{�f��束�2�O����O��O���my<ɀ��75ݪf����ۖ<d��r�9?ͧq�j��F3��\�<����P$!ꑨ�a�&Xv�y���?i���?I�Ş��Q�Q���*_��щ��/N����u�.,�Iϟh��4��'�j�����;��@y��M6B�ݓ�8�6��Ѧ!�h��U�'���{"l��?����eҳ�'��0H���H��V�d�<���?1���?q��?,�.l�0����]Zc\{ܦ��P�DЦ�3�'R�������T$?��Ɍ�Mϻ^IZ}�AB�^���*7�/����'&�F�4�����1ԛ<O�xj#*�b���@�/��b1Oȝ������?�Q@;�d�<�'�?�u���J�=�D)���4�C�ɂ�?����?�����$P��;��AǟL��蟬���ϸG�Hrw��6H��y��KK�_(�	㟴o�4�ē"��زK1<9HH:�E>-���'}r@���� ]Ѳ�1��Ta⟌1B�'���h� $x �(u��U��A�'���'���'��>���613j�;p�W�P8�!WA�#%�8Y�I��MK��B��?q�h�f�4��p$UW���(OU����Of��f��lmZ�m�vHm@~Bg��*��M�Ӏ#��h���&<�*A������=��|�\����I���	�������?F�]�����\��
ec@Kyb�l��1�P��OV���O���R�Ĝ�� LS�H�^���I�Λ8=�0�'�2�'�ɧ�O�ƥ��G�I�ش��(K,U0֌	�A��]=�F�<���A�"�Ip�IEyr�J:�*�R�@�+I�*X*֍�7:��'r�'��O�剩�MC �ӿ�?A�B��]�*�h�m�$ߢ��0���<���i/�Od��'(��'+���d�ȅ��L-J"�c��8oz�a���i6�I�+��ݸ�۟N��x��Q�j�ɋ��"�^R'اWc�$�O��$�O��$�O��$*�Ӄq�tE��I�)뚽��(ͼ'�,��՟��Ɇ�M�	�|��&Y��|�6i���F��^�*��Q).�'�R�����P˛���֝-iY��I4��(n�0��u+���F[?!M>�*OJ㟤�T��(��}*ă�)!�|�D3�7I��,��h��x�O8��f�(�\�Ï�/o4�X��O��'���'o�O�3� |)qkמ`R���5e�K�����l�6&w�1���Sv?)N>�B�F�0d|@�� �d�.qag�OZ<Y�ib�͈����:@QlJ�%�8�%�Xo�I��MC��l�>��,��)X�iN�X�q�`��##z)���4����՝?������M�[)��<T�݀@a�A��Gu6Te�"
�<,O����ۅB>�ӓ@V�{T��FG�(�5�	�l˓�?���$u��Ŵi���id*�l�!GY�Do���M[��x���KT�%X��4O"�:�Ǎ� ����GFe �A"?O��@�[!Q��<�סŃ��P��� �r�fE����srlH!�	>] @=Z�d�9q�.�b)��  ӋפQɳ�o���o�"��U�R��[���9`�&��J�$TH��!�O����	r8�	xU:9�#��9g,�������! $�$6>2�ӆc�:���! �\�f��A���|��֧���E�V�2Pr9`t��'^��a��Q�Z���C��H�")BU�� �F%��T�"�V��n*a3�����_�t%��΅H��`���6���0�,X� ����������џ �*N�z�.1�K�{@@�`��O$�MC�����O �$�O��T`�O��'&��7�R:@Y�#��~)p`�4�?1����D�&4�
��O���'���D#N�+��̽"_ʁ�g�cO��D�OBS��#�ID�t
ӄN�ԩ�ګ7�0�Pe���e�'�0-H�*f�����O�����ԧ5v��g*�!�@PyD�� D�2�M���?QC��:��'6q�"Y�ѴG��X���C55	��2�i�ް�f�tӜ���O���<��'k�I$,d*�!^��+c�S*(d�Q�4��s������OP��+�Bt�w��L�RKF-47��O����O��V�c}b\����w?A$#�D��e� �� 1Fq5�g�ϖq�L>y���?1�SP�ٴ�[B�TcTXR�Xu�i�r&G�[l�����O�Ok��#%��i�M�2� ���c���+���IPyb�'�R�'@�	�DS�m�3��J`�Σ씬J��N���D�<Q����?Y��B�p�с ��eC"�I�,��a#l��F˕���?y���?Q.O&Q�ƦZ�|�t�Z�^��u�+�:uh1�ӦI�'8"�|��'9��6;��$ʼ��3'&	
YӪ� ��['m�����\�I�l�'���H��~����}s#I��7��U���$F!	W�i�|�'�r�_�h�qO�[��L>@��L�uK
�uh���i���'��I/[b��驟h�D�O��i��O��ZD
ޡL� (2�иJʘ%��	�P�S�T���4'�.�����8�U��a��M�+O(���O|�$�O���������2qs@Q0�F�P�)��
���E�I����`�S�']A���lШKE�L!5e�)�-o?e4�-ݴ�?���?a��Q����Ĥ ��(���k�)�0M��aF�b7�$j!*���O0���<��Y��	�`�&+��Ӣ�ڧ�
3G�i0r�'[RMĘc�O��O��A�%{�H�=�i��}�6��O˓`��1W?��?i�'��1A�*�`�(#���l�d��4�?��	�����X����	�LL�Yj@�'p��V[c�Np��W�t�%@�!��c���	myr�')��{��$2d�1�ĈZv��x���L.�����IO���?��'��� �Cl0&�9�Ʉ2�4垈�'r"�'2�P� +�jH���t	��J�����+��1�ǎV���O����Oʓ�?y/�F�D�5�d��sh{�p�����ZW*��'r�'VBY���I4��'��Y�3��9X� ��]�w�z({��i22�|�X��s��ß�� |8 �[�N�jD��o���G�iHB�'�剓]f<�J|����1A�~t	�(9�DM�q��LJ�m�Oy2�'��kء^R��t��5FEL��#�M�`��i��J��d�O�h�Wh�O��D�O��$��d�Ӻs��ZGf��e�֩V�@����٦5���@شF�a b�b?U�Q� Kx�YЃ�Q�)h���p��1yv��O��O���Ꟍ�S�D�<����n�6u=#���b�6�:2$p+1��z�`MaeШ]������ϚU��iش�?���?o����?	�OP���
���MH�G�a�J-�e��C̓0�<=����O2�ɞC}���	F?t������D�7��Oh�����<�GX?��?�#OE)v������X<8�X�)3�	-�	^�="23?���?Q����(~�\q�f�>l-���`��d��Q@�gU}�W�,�	fy��'-��'5��K1X��H���5	��"��y��'���'���'��	*\��؜O���C@�/��h��ӌ^�b̹�4��d�O@ʓ�?���?�7JB�<!�G�F:lXpE	r�ة���R�@���̟����� �'��!�@�~B��F�$k3@R:-q���DJ�# �q�i�T���ӟ4���X���IP�D��1h��#��F�&�B���p����'d�X�@���Ǣ����O�����Qs�ĸj_0l��MLb6&�"�q}��'c"�'x1�'�s���'X�ր���:�j�Y�#�ɊEm�Zy���b66��O����O��IF}Zw2�)�\/A��ȡ�N��	+�-�ش�?��W�����?I(O��>�ѧ�oD�U%��|�
أ`�m������� �	�?=I�O�˓"=��x���.�h ����f�ib$��'�Q���:��� �5Y�M�x"�%".()����iz�'���ʓs#�ꓔ�$�O`��t���Xc��7����έ,��6��O`�eH$X�S��'��ߟ��B�ԣ1L����y+̑��i	��ɗP@�����O���?�1T�X`���I�@hҭ�ҝY�.��'2�'�R�'B�'�"Y��+s�<�j-P�ӅL&|��&�)
B�ЫO>��?�)O<���OF��29��[�`j�QK �n�X ��n�)��O���O����O��ru��v3� ;�MM�MX~���ʷ{����%�i��ȟ��'���'#��yb�ۤ0�\5	�	��=CF�/�J6M�O����O��$�<�T#�#��S������ݤE{eqq*�pĪh�T�5�M����d�O��d�O�Eh�1O&���O�,��@	g���� ��6j:�)e������8�'w��H j�~2��?��'-h�Y���m@��T�gY����������}���J��'��i��5ܴ��s�ػj�܍Ro4{���V���5J�#�M[��?����S_�֝�&�zzA@ߗ,sz-z�C-07m�O
�d�|����}�u��t"��s�O.Nڬ���ަ�yEj�M���?����bV_�X�'��7
�Mc�[��0U��$b�B���e��j���	_y��i�O���A*])G:q���Ih2�������D�	�7 �<(�Oʓ�?��'x�J�)̌g�P��$L�;=���ݴ�?�)O��Q29O��˟4�IៈJa	�LU@5��b\��ZЬS��M{���t�cg\�H�'D�_�L�i�Ղ�n
e*N�Q���p���>i��<1��?���?)����䄥D�v�擧vJ5#��em��􋘬a��Iky��'��	럼�	������30���q�յ[}~�`�L�<f�Z�I˟X�����Iܟ��'l�՚��y>)R��!m��3��ʈA��wemӪ��?�*O����O����3��d8pRш&�'�p�Jܾ=��5m���	ߟ��xyB$\q����?�1z9ڝ�U�����Q�C<q�<�l�\�'C��'��%Ւ�y��'���D<g�Q�
XDP�G،C^7��O
�$�<y���3}��S֟����?	@�&E����q�J�EG�KUė��$�O����Ot8I0OʒO��ӳ0
I��^�n��ѓ��?CeJ7m�<qR�����f��~"��:F��4zSD��e����C��F�g�hӈ���O�P!s��OJ�Oxʧ�~ \����O��(�����MK�oT�:<�V�'���'a���'�$�O �Ь��4�1����1c���Y�J��}����'������O ��ţH�0�RI3��Y�$����A�צ��	� �	�!��x�J<i���?y�'�L�B�9R}��yԌ�l�&�S�4��M8D���D�'���'��P�b�҄q�����*��}S��eӤ��G v`&�\�	ן�&��X,j_����:5�q	��,�¦x����Dk>��O&˓{ڈ�Tlz9�(g��e��\)�@��5ƱO��D/�d�O��Y�':����<��kvb's,x�2O^˓�?����'5��9�6|�e�~D�Ip�VTP��W���	ڟ�$���Iڟ��"f�ן��2@J�=��к0��l�D ��R���D�O����O@�N��S���hO�S	��1��*���#+�=566�O^�O2�$�OP0R�6Oj�'#:�`�I� -*��֫ыg`d��4�?�������$���'>��	�?�`�@+�ni�M]�`��c3�L����?�e
��`��ܟ
�� DS:Ɋ��Bo�'�i ��?}�H�4]��ş���?��D�%W�T�[RjȢS��YcH��l����'Jb���a��|b��Q2YN525EF�tp�P"^�U��F@\3Fk�6�O����O��i�T�ꟴ��!o��I���(�u�U@�M[�e�(�?)O>),����?��MۻwҶ�!D@�LIġk�(��:����'=��'uD�X��>��O(����0�m ��\H�N٣*vB� }Ӷ�ORIj�`z������Fj�`�$�����6��Ց�����	4 ���M<ͧ�(O��1�h)h�`v��8pX���V��[d�����ş��	����|yb�<(�V� ��8�d
�zݖ�i�o!���O8�=���8`�{7̖$\؁I���"Tr( %Ю�?i-O`���O����<���R��C�]�R��F��8{�v���m�jT�I���F{b�'�6�:��'�Ĺ2@ծ{�$��W��I+jL�aDg� �D�O���O�ʓc~�kМ�\c�|[f"���
\��$��4�hO>�d4O���D+}BNU>�����)��e�&`�q�О�M���?�)O:�(���_��4�s�)T�ߔh��$�W[����$?����;�"���$��'8�r���$5eA@	�?i���n���4j�(�������I���^yZc�<ɂӄ\�i���K~���ݴ�?��QQz16 ]H�S�'Dp<8���ޒq���-�7%<$o��{�4�@�4�?Y���?��zK�	p�$�0�La�QA
'�6LsӇ)#W^7�OQ����}�ןL3�c�T��s� �ߘ�����M����?����V ���?�/������h@O�4A��jU@,�Aa�M1��'��8�m2���Od���O�0T�ȱ �ލ#��8�;3��1�ɷ.f�hڴ�?���?���M��y?��C*"|b���@J$\i́!L�b}����yrX���	����O���:� �x�&��;�d�І�po�����[n�f�'���'=rʭ~�(Ox��L~�鱊Y�,��:u��9&�� C2O���?i���?Y��?a�d��1�&��N!8B��ӾE�����I�@Br7��Ol�$�O�d�OV��?��`��|b�iy0少%QT(�5,�I��6�'��'�"Y��#�.����I�Ok�R��͑@�Q1R+�B�hk8�nZ՟�'��'T��M��y��'ҭ�D��P��U"}�$���+S�Q�$7�OV���O~�d�T�`o�����	�,��m��meR��@t�U�$���4�?Y/O���T*����On��|n�>�u��76�L����v��7��O��� /��]l�䟸��џ���?I�	E�0C���4y'��#&r�����|}2�'��"��'���'Y�b�	�-M?�ݑ�/UW\�"#�	�T�/�&;�&6M�O��D�O��i���D�OP�$�!��ˠ��*9��,ʴ=�l�lڄN��\�IҟL���t����'��] V�O�8�D��MJ�FA�6�fӈ�D�O�����N�V��'��	ӟ��mi} �Z Ŵ`�J��v�tl��T�'�I�����9G�&��'@��HަR#V�A��Z�j��X9�'�f�QF�F�>�)���jU( 8ד{�$i D�	��e�X�yʕ3��:S4 �)�.�N$:�#Z4}B]��D��A�nF�m#�5sg��0C�y�g,����{u%W�I����'�('�h��t!\!o:U;ЧO%D�}� �^;����'Q�b�$�%�$���j��61��aCP���q-
Dô @���t6���	�<�SCKƟ����|"��D�[��q��_DZ4�8�9P�a��$ ;c���DԴn�j5z��	���dh ��5�l�*�m*6��A�U�#�T;@
ݫ �����׏��O���'��S�:��?C�|	�Ђ��N�8���3�Iz��P���x�Ɉ�"�_���0��p�4u%4yv�b|a��h�",�T̓��D]4
�6��'��X>�������|h��J�[B��!�ހiCL��u��ßT�I$3� ������k�p����.�?�O$�S�o<&l��bUUI�!�{���'�LTb��O�=�,Q��˄Z��>�ᶧ'Q�I���5H|��-7}R��?i��h����tUu�ġ%*��`"���I�ȓf40d
�̈́{���GZ:�,���HOD5�s�������
�)7tu�@,Ts}��'kr�ܨFJ�5:��'�r�'W�wy�;Ѭ�
8~��9�����s��65��-���O(��#���(x1��'�ʐ��%���@Q��_ ��$R�o �X<n%���O^�C�H�9����	���!��ř3��ȉ��K,X�� ���dK�X��Obў|2�͜�;Ĵ��fJ%c�f�Rr�1D�x�!φ�D��i$�ɜ+C"��@2?�$�)�-OX��!\mT��f�w��Z���-T]z�f�O����Op�D����?��Oe�!�bώE���8��Nı�у�`(*l '�kA�"�<��<y��(v?~Q(H�_���u$�&`d�cݞa�ԕ����iG�� �A1vQ>�<YW���B��[?Vf(|#K��5�����o���x�+/+��� e�.ȉPm;D��eAщI���"����_g�64�I"��=�T&IR�&9��aɩc�8!x��|�<Y�J�CC9I7	ȡg����CFw�<�Ī�/Θ97n������%�Cp�<)�,�G�n 3��C���iv��s�<�WO��I͒D���9iJ�s�FV�<S,K�>����� HR���V�<q��7qpZ�v�!%Ǣ�7o�I�<���T0Y~�Ɓ!&@B1"G��H�<agAD"_I@uCU�O�'�r鉤
BC�<�Ç�+&�a�̊�+e8�q�$�{�<P��$*<@H�Ќ2}^����{�<�� ס0L\���^ ����'�r�<�7DR/(T�J%��T�1у��b�<��'F�8%2�0O� J̀���C�<	�`�%�:d�u�j�~��U���<�g�)n9��i��H�����)�z�<9�� �Mk��P�A�s�<Q�O��s2�T����J���!p�<B^=�n�a���r!������V�<�M�"�e��T�&pS���O�<���ۤ)�
����@�f&���kJd�<9���7�ʨ�$
ͱ�.X�LR\�<��#X�j�Tj���)S4�����p�<�T� C8�	2ڤ=<J1I�Nn�<� <Kg��6���`D�ǜin��"O\}��K&@���	کh�J��"O�$Iw)L�^�ꩁ�Zk����r"OH�#1���D��&��5�$"O���� @�� ���L�N\�@z�"O4�c�N��[�z�[g�/p>�� "O�A�h]=g�]�@��\X�
�"O�D��� �}��9���2/r(��"OvpWȄ�TXa��ѕU��r2"Ot�y���mzx�m_�Rfp`0�$I�;(� ���e��H�0< z��Q�@�*�B�I
O����rMX Q�t� ,�.Q�ޅ��o
��U�Σ|�'�	8l�V���+�Nؙ~x^PP�'�nyPG
��5�B���P�zԖ���q��Ic.5�O�@@���I.��	�A[$ۜ!;��'nQ��I�4c��ɒ#q�hrǡY�B�D=#���~W�C䉃:���BG�"�Hy�J��ɚ��I�LS�`��E��	%W�򙱗l[${�I�0���y뀙���)$���p�Ĝ2@���t��ip󤄧�(��	�w��D��ݗM.�}��&ާXk�C�I;1q�@�5�ʶ%����f�]&N�C�I?[޶��S ��BA!M��B䉉IG~tٷEÄ9㒱A�핗�ZC䉛@��uq��˺7��9�@�++8C�ɣ"�:d�a.�<R���/>^��C䉶I��܃t�@3^x��A��q}~B�ɺf)0x��怶taēD�n/LB�Ɋz�4*�ދE�2U�w)OZ�B�I�I��AYPO[�>)�1��;-�C�I.17�8�b���Q-�-���!�'������C�m6��q�	)V^$1��'�8��	����JC�@P�'���W�D&uΩ��ν�J�{�'dBJ;2��k��
�] | �'�����E`tK3)�I�'T�d��ˊ�Z��n��sl��"�'�����(��L�L�*U�r���'H��6�V=y&cQ��'d��*�'/Ɣcu��5u��)�h�2��	��'���0��[�����&���XQ��'�´x��К0ּ�����=\���'%�A�玘�%	�1ՁW�3��t��'�j,)��:7�q�F��!#�"
�'d5B!�*�2�4��Y
�'v��B��U�V1�Y��.40���j�'���`"X�>��H���Q��a��'}zf`R��Zci�Z<|80�'>ͪ�.C4 � �� ~~����'�X�k֬�1��YY��b#����'�bM)��L r�Z��A���q��+�'��t{wOȎ8�1��		�lV��R�'Fr(Sܨ;�<p�h�1����'?�`{vGխbʤ�u%L,`��D@�'�$ݣqk�:�L�!F⋌T�Hu{
�'d$P���Kޜp�GS�6�y�'mRA0Ӫ\�HĚ��X=KO�t)
�'���DU&��U@ �ĄF7ƕI�')23C���A�P)zg��;7b��'J�h�ÒH�\�1&jJ�f�(Ik�'j��x@L�"����F͇5����'�0-�n�;n"�ي��_.3Cd��'J��s'­u��aB��2rp�'�u0�C��#� X2SL�u�x�q�' �(�r�M2q����bJ&r��pX��� ��R��ť��(�j�t���N5.^]l�aWRm䧈�rB�(J�8��QP4R��b쏰�y����0ՠ�`(�
K��]�f�թ�yRڀH������',��y��'yE�e��h�9�h�rł�0>��HC�k�\1�Y,nU��E�!U��8J���ʂX���F�{ݤ����#:f�H���+&
�0�G?X.#<���I�t�B�H���c$���+>׾���k��ud�i�pI�2k�!�H�A�VE	� E(��L���{]���`E�@�B��6�ؤ�0�,x�#}�w�Hu aL\}X$�s�&\�@Pb���'brqq�$N�O�6����[}4�4�$.�O����bS+	�4�Ck]��u�͝r�'�X̂�)�x�����Mݕ:��%�ۓt���V��d_Z���Y{V��a�2@�{P�4^���oU�y����Ā�_�QS(T�h$�qc�ڸ(��OXy�2&�	C�}��N]���������:)iC�,Z�@�3����m!��F�e��9!�R&j����%n�l�XƎ32� d�bgO�Q�"��)ʧ.y��[_�� �_�4��EȈ1d!�DZ�Z0��
����Hk��P�,R3�D�I� ����A<LEZ� 1��j�ʊ�����D�f�[�z=:ab��@��{2�ǃS�		@�
�L-px�6*��!�g�V	^%�=A%��.#���%�/�O��B��LA|Т��"O����I�X u�� l��
�ME�<�O��p��" �oٲ�J�mL1�'�B��wG�
�N����|���OK3�����4VN����
Q��hk��9O���Ed�5,�>��g.@8hy*�cG"O� ��Ӕ\�� w�\z��e Ta�|(0L�1C�O�d�EM$���I�n�����@�:^�J�"��8�X����`��7-Fu����ƴ���	b�l%�(׮��+�pmy��'�ؐԏ��YD(J3����	�Ó>T4Ԋ�J@�]V�'B�С.��B�z�P�oɝ~��+�'�rH+���:���PcԆ&1<	*� ��rݠ����.!�VL*�˂��h�J牋|�8
�����f�30�C�I o�T��!�|�~`�P��
�8��Q�(�ry��OE�@���c�9 ���S�	�L@�$�Ʉ;�,5���-/axb
j��{`��Wlx��!�$)�:=3E@Ʈ�$L��]�#Q���d��I#P�p���[5�Z@���)k��H^�ϓ&�`M[7�(8d��� ���|Rw̜/E���Ib��	��B�\U�<���
vW*�:*E�0�n�C�K/8���bs��I}r#
�?�O�@�j.k>I�w#�U���=r����A,�L�8���Q8��2�O�9�ՠ ��S�l�p��ЋY�hu�A��O�9q��+�����F�uW��\�'��L9���Y��݋�:ެ 3���%���q��H�E��)/��I�,��q1�"G7\
���C C��& 7c�r���[-"̭2�ȝ(���$!�CZ��P$��
#�(�f I��R0�=�O��ݎ4*T�AʥZ^$ `Q��h�C䉻;Gx�I�O�'�	ei�[�F��ec�7���J�����6�"}��X�!4���U�YV���4L ��<���L3�)��a� n�\�2l6vK���Q�&D	x�p�Ņaa�l��Yuza@��W+�\���w����*كLab�H�dN�҈��'����ټ&�q���V$y��Q�6�v�1��X>q�%Z ��>L4kGODX�d��/�a��'ɠ7^�:CL��a�V(�vi�L�ў�I6`ӭW'�ͻ}��	�2��9#:�ѳ��o4����ɔ_{@bÌ���{sc�1j��}�.����'�d�I&(�)L�N݁R�ݭ	F��K<�QO�#��p3���sl޹��
�L�'��Ǘ�!�l�a����f��۴,D�q�mH
n��E˵�E���%��J�;gZ����!O�;Z���
c-@���jX���A����R����CJ�b!�}���r��V �	9�P�'-���fصg��� �.��U.B�;�"O֥� ���)�v�2�/!��(��gE�I�<x�fdg�����l=֤�Ӻ+lH->��@R��wށ��]F-��Jr:1��*�O�ig	�.Hf4	�ïWL����d	I�m���BcK� ����f�'�U��`]t6��ţO*,v����{2��t~����S��Ms$HB ��OFT �	Z����v�A�	NH
��'iR��%=mΒM���ξY~ZY!�8�����$�4\y��	�'|��aI��P��-��d�2t ��ZV�
#��"|���"EH*G�|��eA��2�,Ål�<r� �s�ϗ?R��d� �� ���kp*����z�T@a��J�#{pő���0[�� ��E$F^�U9�_y�h	�W�:TAc��Z�c��Ē��� ;UZ�;E�dA��%M�7r�����P�FV"��IKQ�(!"�)$a��)���G�PD0���%I�C�Q�2�,}q�
U$s��Z�L�D��*���7'+qO� :����=�x{"#[�_]�¦�I0#\��_ ��e(��ӣ#�DɧN�4�2a�:�&�E툼v@�}�A�c���'`«T�z��Z�Ȑ$�F����F�	�~�L�1��仵L>Vb�Yb!��?Q�@����b'�V�nނ)�h���G�ɋdk60h!�$�"4�x�r+B.vc�9XAEY��ұ*D�Lw"�`3n��5���g�i����=A錘����R?��*�J��|�\B��!)�C�A��ZҨ@3��[5`�x8�$�
0�$��#�S>T�b����x�H�+r8��ݝ�}Bg���0<�ť��$~�˓�
K5�` ��@|Ta��b�.<��TC�Jqh�O%�����+K=����!�OT��G7?A��[_��a�-��9�^�ya�W6�8�>m+�9��-c�ç}�գ5�4D�`ٓ��y�����ë#�k	�]9\]��勚l�0��Ce� r{c>��G�>y�o�~9��k���~��£��e(<�hW�.t�� ��!����5d���F�R>2za�ߎ ��JެA�7��/t�4M�D��FG�|�ȓsV,c�hGu�j�/.�nȇȓ[^�-�S#M�az��._#-SV��k`�)R4Y�58I3��q?����:�c(�+�����KE�"����܉��X �͐dL�X'>��ȓ"�9a�cB�a�r�k�D�g�h�ȓ@����!�`�
!�� �/P4ۇȓ�pQ2�|�a�!T�ZE��I2D�������*Ia�ǁs/"�2ë0D�h�%�]���(�ǚ�r�U� �;D���U�ۤw�d��/T�P�
�P�9D�h�`�*�0���Ѽ�����M6D��"2�d� �r!��-T�!���2D��B��sf��!B �#f�TH+�n3D��3r�+vm��pi˄�*��/D�@�G��,Yn�A��&hk�,�%�:D��p"��=0!������.�\��c3D��#��\D���B�.J�B�AA$$D���e�ʲa��	0R��
x>�`��4D�@1���:Z3���c�?M���+��6T��"*Q�}v��!��
d�x �"O
�j��:@�<܁�(/6��Qg"O��BcF���p��D���"O�X	��/��+���&X�H�f"O`�'�&b��%��\�p	�� "Ot�1U�'=�(����*'JJĚA"O�${$-Ryz��E�5꼠q"OH1���hn'�0#(�9D"O����ct,�d��F~Iw"O
@ �׃%K�����٥j��mb"O֍S �X�Hq��O >]2��"O@=�.@0?��I ��Ԑ,R��A�"O�!)G�A &"Lzd́9rL�V"OX鋱n�f��2�#Mmy\�Y""OtM��d� v�]#sY:K�ܝ��"OV$��D�5YE�d8�P�lYh*g"OP\HwȄ:Pؔ���Þ�	��� �"O�0ځcǻp���1��u���`w"O�4�$j*x[��eJ_'^��93"OJ�+C�5�&%*Ҩ�N��x�"Op�;��vRਔ&��:�4�"OL�
vcEf�����'����"O���&N�` �8ab�u,	"O�l`��fQ� [� \��"O���9a�!�Վ�9l"Bpk "O�]cG
<���B8cy�"O��ĢT$i���������w"O.��2AG�q8�@Q��S=���9�"O��� 
E�6id$�q`�.��E�P"O� �[���&UD���Dj���It"O��QJ�j�x�V�*r�5�"O�p�&�r�XйP���'k�	�"O��p�ƀ==V|�󠎪Ph�S&"O�5�0�����x��7N
e�A"O�l�R+֣t� HxL"���"OV8Kt��3ɔ)	1@S/S:�4�t"O�i00��+K`1���5��XC�"Ol�A���6�G�N<(���"O��j�԰(��D�B�7Z 0G"O��{3�T�(�P1$�w�D=C�"O����ԸUStA���!�"O�#@fѣz��AV"�U�U��"O�[�JI@�DD,J�1�N2�"O�]1�d\
p�vœ5��8*@�թ�"O�i"AQ�j���,V6\*�Rq"O�x1��3Q�%�F0G20�2"O�A�J����亲��0�m�p"O�-b�i�� ���;7�ݺ.
,��"O��&�����5��͕
8�E"O�J��`9�4�W��:0��I�<�5j��JE�;� ��5��\)� �B�<���ء����'?,@ds4 �W�<1�o��n
�D��&p�F��b��P�<i���r|���ʶL����#D�<��-���,a#fg�j� ��	�j�<�D�j��`AFI�=W�ɢ��d�<yC
����e�4����$����`�<1� ��Ye�PR"ҟ[#j܊�!d�<)'A��bY0��doG�*��G+c�<�� �	���L����`&Jb�<qa��B��X�q�Wp09����]�<�����2�4��)�a�B]�<94gӎ"1v	����(�SPMQ�<�랳i�f���Ϛ�:��*3��d�<�r�C�16`�J����]4��\�<�T�=#"H���¼n����u��X�<1�P'T�1��9Hoॺ�'�N�<�FOů~N؜{�Ѯ�P�5&�L�<�K=��SS�[gXl ���F�<Q�˕�F� �����5y��*�@�<���މ6D�i�Qغ�t���BU�<9�B��|�X�� 8��k �F�<��D�4V
�!`Sh�4�qw#SI�<�'ވB׶	
�D�)���A�<QE�ٕ��L �AʫS244�#'R�<�d#	7l L�a%���@����F��w�<�BDiO�8I'�ۡU�"ف&��Z�<1�CR�[h@h֯9p�v�Y��IU�<�� ѝ.,�-8�O�R���.@x�<a���	3 -�"����T�g,�u�<�G�G�%z2Pq��_)9�f�B$z�<)���0���b��$n]С��k�x�<Q��(q@�pyN�w#�As�p�<Ʉ,ߺ U^|�!�� 墥 VC�P�<���0
�?Qb�*C+�.8�ȓ+)\�[S���E�������J7���ȓ+l���c�H�[m6j�ÀU&���ȓ0Tm�E��{y�@�GSD� ��ȓ=dV������l?f���h�~l�`��N�%��o�Cה�Sv	A�5���ȓA�pF*�z���C���-�lنȓxkN%�AÃ~��K�cOq������� A��d��};0�Ӆ*"���S�? ����uV�Pǋ�?�	2"O丸�Ȃ0�6y��=N���b"O^8
��� ,�A�B"~�3w"O��q�	{�58�HQ�#^pD�"O���w%ά~Cشj�SO��3�"O݉��A�M�F�(ċB�>A�W"O�P1�h�B%���־]�	��"O��r`�ęR���Z�Iʎ=Mp�(v"Oʜ %I.�N��IK�VDK&"O�����
 ��a��B��Р"O`a姈5)r<r*�� ��S"ODl1ҍ�o�R�+��X�N:U��"O��J�g�]�2.:�w"O�T{`��i�V@��N�"�Tb�"On���A��>W����[���,�f"O�!�'���y7���oH�trR"O�T2%�
7ζ �UJ[�1lI1�"O��+�D�FE�w�|#"��"O��`�Ǖ�cF�HbtHA#-c"OV�!A�ˀw�����?Wx�Dʡ"O�!��D?g�x`�"d��w}�i�d"O,y1���u!�}I���lݲ��P�'_���!��Fm\�aT-�`*.D���!�\$A�6V�J���>D�\��]�r�����:�pd1p�;D�Dk�A��LU8��R�ѳ�D	ѡ;D�\���f	��h��M`T���9D��gC/z� ��5$�1s��#1D=D�DR�@Cy$��Cc"g��y{`a D�����b�Nm�����K��݁��O2C��#"	��t��Fm����B�<K�|��ǣ��A�ъ@�0��B�	����H�*�zd�Q�R�n��B�ɚ|J�0���$�B�� `]�!5C�I�Z�8miQ	��HHshَF��C䉟43��V �)��Q"0$Kl(�C�ɜoόUA��A
 h�z�%ʔ2��C�	x��De,Uh��h"jL�I|VC�	r���ȵc(��#'Х,hC�ɺmي%�sJ]�)�Դ�a)F�8C�	�{ V;�ß�,���[Hy�B䉯C��X`Vh�:q���b�B�:,�B�I�L]�lH�dQ"��8�
5�B�I�nV�3��B�~b� R6�	�P��C��!�,:��[=
�XmP��Ϳ+{�C�	5iX�@�� ��Eᴉ�4�����7�I&E��P���\-Y�S%��o��C�ɑ� |Y!�\�8�!���b/XC�I(u�h���*��=~`�-� �fC��iݴ��fV�C�
5�F�����C�	 B�Q�k�P��ȢmA�ʈC�Y��I"��*YJ)*��w�NC�Ʉ6��$*� $~�0yۑ�]<[�<C�	8jU���Ճ=�mbA� �TB<C�	dԐ<P&L�L7�����_EC�=gp�`�F�[�q�ڼ���;��B�	�*g��S�\���cB�^�B�	%&�����ɸAf�KQ����C�R-B<�E�-Ƃ�S�	��x��B䉇"�@Y��H�q�Z�	�B�	�l��C�x*|۲l����ꓞp?�*�[7Tq����
'Z�
�M�<��ز,�2��pmV�>�y�UK�<��G> ��D�%ޒh���#7&]�<� <��@�Z��u��c�I��Pz�"O	#��m�E��Y�x28"O^���!ƺ{(���T�=�����"O�i���.VO~ipuN
�
��"O0�8��?C��cu�Ԛv��� �"OX���&�5#���E�;\���"Ol��&�3U�0�F�#Q�����'L��j��T-uU�%��$��_p�{
�'nu��ک&	>�j��]
 n>q*
�'1"(Yb�-E���p��;}�#�'.:��Lo�h�,�/	���
�']2�qQ�S,7>��R��B#>v5��'-  r�Y�2�����b=��'��T�ER( �c�g�E�����'�8�pG�]$�H�/ډ9���c�'�@ydjրc�5(� 
�6ژ�9�'�����&��{
(1�K�7*p��'�����jx���Ø�!R�I�'A��0e���1�cJܴ^�k
�'�bq���?o��A�/D�	��'#�82�բu��j[��rE��'n���R%�%-8P�S#4��M��'I:肵��`�A���Q����'aЍ�#�J�f�*z��{Ip�j�'������U�a'�89���'�J�pU�ۇ"��͒����Py�'扛�B����0��a��O��k	�'�`����/)8Nu���F�]r�'�x`����&5��8�wi	i��x�'\�IU��,<��
Ga��p�
�'�40��(�欈���-Y�n���"O>� #���\�Z� a�U�N�b�Ѐ"OLA����;<��@U��"���"O�Ex@OۯS���2�	Æ7�p�PQ"Ob!+ Ň�dƼy�7��6v�B&"O��0�͋3E��R��S�?Z.Eq"OT���j�.Q�p�! M�<CF��c"O�$���OV!��-A8VC���"O�ܛU�
h��ׁ܁"�yy�"O������'iی�B�JB�|���"O���JsE:��`ҵb��	�"OVQa!/V3Y���snؐ��D"O�!z2�^�@iA�8�EW"O0��\W���N֣�|�p"O\4�2͊I�PH�͑�2$�y�w"O����kIN�f�K���1"����"O��h��կH�摪�L�"
Z �"Of�0jB�H�BD��1L��"O�ġ5�K�k(|�5�ǯE��"O<�V�ۀ�BL�vhΧ
.�q"O�4XD�Q'F��]�GE>�(<��"O�!:�ER�[k0h��%�h�"O�P؂��}��(�e ��@��"O��ӨD�F�0�;B�!\k\�4"Ob�����g$�ɀ��ƳwbP��"O2��FR�`	��M/ICBp
6"O>�p'��jf<�0����U�v"O���Q��h`������9����"O��bG�Y/R����s�~���"Oz �w)�/�t|� ѣo=�|Q�"OX����Ro��tQp�� 5x ��"O���H܄?���"�܂F�� �"O��Q�kj�4�!ljni��"O>	��Ǘ�$Gd4)!��9�� �"O� xLSv��$m�$`�̌sDmjR"O�Q�ІPA$.U��`�A�� a"O��
ԅY9��I�E��5�F��U"O���p�Ή�$�JG)O 7����"O,��l���@� 7�ڟps��zS"O�m)���i4�٨C��3Pa���w"O@���H
8O`�0����wV|��A"O�!AL�b�2� �#P��"Ol�Ɂ����YeR �����"O ���@�)v�2WŁM�F�b�"O2��j�=$S* �%D�~��p��"Oj�����2��(r`�Q+&|z���"O���nH�}�r�b,>'_f���"O����m��l�Ҹ�0m��cA��I�"O�yآ$�:r���"A�T�W)6Q"O�]�6b�?C�irtj�{��"O�ܓ�g1@Z����;z��	"O�Yp�K]�Al.Xf�Ͷ_l�"O`D�d�A+�X��H�K���F"O2A��@�c����ŝ�G��C "O�mc0����RT9��?�X�W"O�L�� _wP����V�Y��u��"O~���cG��(А>�̨��"O�p"ՋU������E:>���A�"O������~�r��ՌƜ+I�l��"O��B�&Fq�*��K�(�t�s"O����&�:���R��B0@薍�"O��2R
:(��!f\_{B��"O��ZQ�W�5�H�{T��R�F���"O�1��'�(	w*�f^3]��lɔ"ON�	A����\jr(�"w@�8�"OJ��F��7k�6�gE۽\md�J�"OZ�)ićC�� �n�K�"O>�Eh�6����GVN,��"Ot;+ۏm��0�f�mATUR�"O*�	1ћ	��ԉ$D�(~3<2�"OD@�r�V�`P�H ���
}B^A۲"O�ez�Aۆ"��+aD>T�Ա�"O*u��(/r���_;|�,�d"OTdC��	�D۴@�YЊ�G"OL`�l>�����CZŲ�KA"O�lc7�	y���K�!�!HP!�"Oy*�S�{|*u���?)�5�W"O����� �Qs'OA�P���g"Ov,��͚� :�t�1/�T�hq"O��FS1RR���-W����y#"ON��Q�ݹ'��p�;,]�@�B"O�ѵ$��0���b�1��NB��y���*>��P�Mٝ`a��Y#J�?�y�F�9q�K?	:-�b/��y"m�:,�\$B�	�Ȳh�S"�y��Ůk�V8c��-��B��Ұ�y�`V9
��`g�{P�t��?�y⍎���s�M޹pI`@2@X��y��G�0^b��'u0eAp�Ծ�y��E$!���y��I�nC�|`�H_5�y"O���<sEK^"yp�UJ�����y��5K�1�DE*$��܏�y�%����l����D-�y�G�2	�,)S)Z52��M��e���y�nڇe��ԙ�	�&{�y�썷�y�ƅ�r�^X����#ED���N
��y���	c�
����c.��e�H��ybn�2K��(�R�# )*�fB�y
� JT�aC�'��]�$�M��\�"O��Pצ��k.h�'��6�D�"O�@���K���bD�Q�]�4A�"O�*4D�S�P;pe��57��04"OQ0r"۳;�jȺ�Œn8��$"Of@�RDG�  �c�$
;.���#"O��ړe���SR��T#"��c"O�R��M�T+B�۷���v�x�G"O�h3�Ά�< Ό��C	v���a"O�q8У�m���4�ӹ�p�w"O������>m��i�-E2���"OfQ(��H�/
��h��7b
9X4"OJ�ȷn�>����h�*GjFA�!"O@\�p`ۯ'�4L����& �|�K"O�����l\�X"�Q'��A$"O ���i��	>�1sRn@r��3�"O�<�1Zvr$�&�ob$���"Op`"���1?�� ��N�=K2�t"O���"ԓ0����F�U�ڜ7"O���1ŉg��ya+��d�Ρ
4"OQ`�L�$OZeZ��?u�!G"O8�X�j�pit�
���*Z��"O m���"Z����s#�wG^�u"Ofd�A�R�	�����
�& p�0"O^�).�
:s���(A�j. 4�"O�)
�"�V��4��&��t["Oޕ[�@-ztk���X� +Q"O���5E[�B����a���:Yb���"O��B�w����&���4I^H[�"O�({�"EJ��b��ŭ'���3f"ODŒ�o�ʴ
a�	h��ճ5"O�!+Ad�&Tj��BoߗTτMP�"O���[V�l1��ӡF�ȴ�"O0  � �1'f�s�V��&��V"O�}25)-r0b�x���)ax�b�"Oa��B�Tk`��$]���e"Oi�p�34\*�r6�P��L��"O��P)�-`J�y���]�
�I; "Oj�H��9S�i�(]���I�"O~�C$g�?�.�bB�<c�5�"O@���\�e0P����*r��!�"O��
��V>'��E��"3e0z�"O ؉fI56�L�EhB�0Xi:"OL��5 \�"#U�VG�B���"O�)C�D�dh��D�N�v�"Om�3�-4�0
Ձ�2�����"O�l���� w`�3��~��C�"O���'ר]M�X��`Mb<d����U�Oi�5˳M�<*�F0��hY$�� 	�':*(��DW"[`�Ҧ�X��+�'��5R5�"xt <+���m���)�'��$�C��9_��u��I&;ߴ]�^�<���.GĜ�����|�qa	�oS�C�Icl���&�nfn�PW \�C�	&9�!���t�hm1���)tWzC��>�.Qbc${���r��0���O��$؁Uh�h��>��iG�L7&8!���$2�ͩ��F{�	�T��!!�d�j�<9�fIA*LٰV�ʔL!�b�|pX�`�!����-	�W!��q�q(�D�6XAzFB�Y�!�̸u�t�t��/)_��(s��!��n8��$_%ANv !"BO�b�!�B?����g�>Om����C�)��y�)� b���i�
 �l��Ņ�]0�9z"O$��6L �w4X� 7 MA��'�ў"~ւL�Z(�ㆈoM��a"��y2aD~̌aS���3~e������yҏ͆/I4�ɡi�1	�L��8�y2&L�F��hs%�@>~�P��$�9�y"�T���Up��
Ǵ�aL��hO^��-�A���#aQ��8�J��h����Qa��R:Q��A�pm�%��d�'�a~�*S�/Y<��#@�f�pe*�#�yI,A(�qB��@12;���� �5�y�ׄ`,��ţ��M�����y��W��t�֪�"��� #j�y�q�lq4�R&�t��"����䓓��䓧���7��lCS+Mxb��<�!�D�]�^�oQ�[g��)��39!�X�Cx���tEҵ����,P7!�99�:��
4]^j��G!Xw!!��[>Cئ)�D曦L9�h���K�.�28O�L�OD���a��M>d�xP;�Q���ɉ@�
�`���n���c0$�9+m.�O.�d9ړ���\��{�;=��p�G��h���b�"O��9d�u�.xR"�2%�~x�"Of  ��΋j��%B,�Pљ'"O֡�#��S}�p�i�Ao�CE"OT�k��y�d�T� \QB�"OƸ�M�>�ȠZ"/҃PD�"O`����vN�4�_0O�NYI��'�1O>iIԏ)&���R�� h�P�!"O�<�N�5�\��3���2�Z�ju"O��7ȏV`�R)^�}��Љw"O�}Q��#�Z�)ι7����"O��(�FDoK�9�%i��2�rl�d"Oh� Fː�M�	�d�RhH��0^�(�	c�K���0�CV�D VJ���g:�O��9����t�-�WL����Ij�O���v
"?:���n���0���'�z-�ዋ @`�@e��{��A�'�@�"���!s�A:'�:�e��'�"���h� 9��Aʜ���'*T�Z�OЛ]z�M褮'�(%y���?Q���0>���I�&��ۦ�����C��o�<	�L��h}tX�'���#h�<!�H:'��:��."$<����c�<�s�Ƥ��� ��ȫ.�����f�<����k@�ڵ��K?���Ad�<���N�p�5��x��fh<��痳�0lH�B���^ ����"�?	��0?a$B�%p��|I��{?��$�^�<1�AE:w� %����]dyZ���U�<�+\o�D�6�F�S%J*sOƟ�$�h��	b�ܩD���>�䁻�F�2�C�	��>:MZ��p�b���(�C�	�Lɠ�BSN�,��,�G�:��B��BhyڄE[�LZ��c�޿`Z�=��lM6I��\R�����*~��C�I$��U�b_�d>�e��#�:uՠ��5����G��Vi�ь6\�E�&�7D��k��	�1^�Z���l���\C䉿=�@Y��c
8eLq�Pc��h;C�	P2|m�⡇�u����#_,<p�B�I�1�FH"AI�pw��1�����C�	)d���3KC?Z�Pr�/�C�	;Ь\H���
�|K��X
�<B�)� ��2e��T�<QpFI�`��Pj`"O`XK�'G	fA@�R藃�r�ڦ"O��s'mO*+�&tk�[(���E"OZ�� �O�v��zbgDiN�e*g"O�����-���f�?|$n0�"O@�z���:y�x�#�C�Q�LC�"Ov}����"�c�M	"4��f"OX���ڏ7a2�+ ��s"OB���V��\�Bl��#�P�"O��jq���	|�`{�� �r�����"O���Q�85�0���7(�v�����f�O�~U��dO��8���nD+G;>��-OR��^$V�ty���<Y�4:f��#H�!��Р/�����HއXWb���ݢ xџdG��ꗡ0��!�2�)���¶���y�A�I+�5c����x�D�r	�ȓӠQQ�t���7D�e�Rńȓq��q�@-�(1�i�I/��r̔*���o�p�XQ/e�م�	_�en�� �.R��0�Z*t�6y���u��DҒ~eP�P�J?X��̅ȓG��u ��ѢƤ@GB:{	r���gJp��O?�hz��J6n����n�jY ��F"Ph���J9K\���3 �4*���R�Š��M�;�4���3�,��3��>|/԰(S�6p�&����Y̓����AB�r�$�oΜm%\�ȓ,�l4 ��]fJ 3Q/@rZĆȓ'"�1։!DjPyć�=�č�ȓu����ѣ:l>	E^8{�Jx��S�Ĺ��"u!�� Pĉ	.	�E���MP���C�
�pq���2��ȓi]()Ё��M%.�I"O�(6�~���	M̓g�&M�t�D!�Xq)�
v6'���	)�J��V̊<	^ڠ��l��`*�C�Ʉ��)��7�`$�gǧ:G�C�I�^ �m��G��B�G�.�bC�R֜�1rC١Z|L�� L�/]q�C�	� �"�C'A^�aR��9�n <{NC�ɱ;�P
Ї�<4���#�_*P?.���n�'/�D�׍H�V���S�-	�J�XTb�'9��)0�޶*(�lGB�����y�%S�x��	2�m�p4�ks� �y��P�'upq;R,`p�-�"B�yҁD�N^�x��BkX���h��yR�4ma�IQ�'y��Q � @ �yR�P�}�8ip�K��v���YW��?�?a��hO<"<����`J�8Av`�%oL��B�q�<���P$��CH9��]cSY�<��K�= ����w���!m�<��J���˙�;�Xј1��g�<�2/̇a�6�a�? �8���A�g�<Y��BHҽz�;C[��k��Z�<�OT`Y����0����fT�<�78
&����'�:�M�S�<	�H�>n� ���
���2���d�<V�#j"R [��_�y�#jh�<)�����H����]�|��0n�i�<�2�� ��1��䝦3�֥0��N�<�DHD�i,h+�	��"4����Hh<Q��k�tU{���fq����y��5q��M�8Z^���V*��yr?+�x��� V�C�
�W ��y����!���RCY%�8�1�A*�y
� �I� ��;5f`h ܴF��u��"O�帅����Q�2�K"wd��s�"O��{� ��gp`�1��Ή(B(�� �	K�����ڤYyPϞb㖱��V?�?9�'r��B�$تkj�@
�KǇ	�"
�'ݸu�9!EP񒂦ލ}��'��{u��8��$��AƖ�	��'ۦx�n�b�<�����R�d8�'�b�R&1�Jt���Ӟ[��y�'�&���������ᗺU��Q�'��3�n_�q�I
���$Ƞ�8�'� 8r
Ԕ#F��q�ŕ���Y�'j����%�-~���[�ʹc�
�'�VH��)��DTJFeخ	$�2�''r8��jO8WH���B	b`%�	�'�>T!(ty���ۇ`RR<X�'�By1Ɓ�k�� ���Dך�a�'v��!��)+���`@�I���'q| z�G	�6����Gx����'8}C��ȼ8�h��g)D95��y��'��cDJ�JM�I�hD7����'Hm�S@�X��)�� ~��{�'����V&ԉ5�&�W+�/my<\y�']1H��f�T�\�gs� 0�'\ ���<S�5�&`bi恫�'�L;uH�l�$�(sEF�Xo�UC�'	D�����*$:�̀�&N38�h@�'��e���Qro�ec�3���O�<A���+)���dN-�-��Vg�<	��XP=��{aKӑm{ڝC��CO�<��$ֵ�]!�G!��mK6�HM�'k��'
>��E
� pJf�)u����2V�#D��2�D�"X"6�+e*�1�f�""�#D��hb��%�`�#L�'p_��Ct�"D���d암8ԌPP�k�zW|Ce.D����75lD�{p��,+�f�
�,D� Df]*AZ`c3
DB�j��?D��قm��dN=Q��YN�"��?���?��ɍ6]��	#Ouk:��"	X!�$ػq�θa�(�6NV`��Ǐr�!�	�<p��GD'PJXՠ�gǞ_�!��ڱ<P$庖�Q�,2h$:��M�r!��o�<Eɧ�ɉHC� q����!�
�T0i�&�;H��jE��I�!�G��P�ᔨe?4��b&�i!��۱B�� ���!HB|ɒ�'b�}b�',�$�0a�V��h��W��L�N�&�x��D��\@',O�mTT!��n�!
	S� 3D�h!m�.J�H��'��	��%D��;&�Q�#�AY����0#-#D�����G�;Z�����'������-D������2!���%m;cî\��*D�xQ����e:����2�t�;�,(�O"�I�"�.D#��� l�r��A'�/�D�O��$%LO�T�wM̚Y�ar%I�$��"OT�hC�ܷR~U���谡�"OB��g�5k�.�"���4�f���"O�}��� N�����L
:&��t�"O*�C�I�c���l��#�F�	���:<OJ-����>p0�7��;Z���#��)D��X�$�`�����քΜ*�E(D�p�����U�`�H���f���y�o���P�RH�9�&�óg���Py2�&v��\YA��]�~�9/�x�<� ��Ç�f/�(�FYK�9�"O�05n�2����Ǥ/RPj�*@�"LO�-�j%P\Q��M--l �Bc�'�!𤁳����HJ �$���X�!��R�:rb��7�;+�v����ؼ,�!���Թ1�BӰA�����<X
!�$Ɛ+k �q1��=q��d��'K�:�!�d��mp� �Q
M}P�����Ae!�$�<ywr��tcH5���&�IG!��۰����cb��x[���t��_�O�� �b�آ��?'�)�A"O����*@%V������4Iq�)5"Oƴ�J����ׁ�J�6���"OD�K�Fدn��yk���<���`�"OT �&�/�C�j^eB9�$"OP���
^6^|����g�܂A��<���U&w���"BO�Mn�����i8�B䉝E2h��\4� �D�� @B�	�;34�q"!eFpq��ڒ4-�C䉚0l��dH��w�"к��Z�4��C䉓&�n��$V>;^& hq뗊%B�I�LC�=	�c
 �ʋ�mC�C�	>sӞ]1�����B&���>���O"�O:��9�'.c�˅,��iM�)B��8H����J�.�3E�,>�h�a@$�H�%����ɤP0hl*��JNB��g��>R}�B䉯9lt0��m_%�@CUMم+�BC�3/�(��I��`�ħ�3bNC�	�a����Pʐ���%A�n��B�	
�)�Q�K�3��	���R$M_���?���)��6`^P�q��B��L�!�$�"S0��hR+@�/��(
��ɫH�!�D�l>��7��J�v���M�9�!��@�ش����R���:iH(�x�'�2aZ L߸[s�`�l�P���'���ZE�� \jbgݔF;F0*�'2�@x%!ǨuMdb�`��¨�,O�=E�Θ�*X�S�j�b}�@�2�yra̎*�Xk"b�x�����yN�	!#��0��q*������yb�'�����_�lɻ��
��y՜e�� ؐ柸I�8���A��y�M�`4����'W�<�.��dE�yba�=M������D����T�U8�y����ĭ���	97ft��3��<���?�+OrP���j�V��u�JhX0|��8D�`˧$%P(��l�x�@��6�6D����
�.ߦ�c�.�Ȁ`m8D��[���f�^���g��w��c6D��C�(��q(�̅+�5��4D�!A�D 32�H�#`^�MZ�7D�����������&�����p%�(<O��d�O���m��(3$�	���Ǯ,I�ܠ��3D�|�jH�/eRl�'dءb���ئ�5D�, g�Tur�x��#�<j��.D�(	s&�t�~�1�Mx�� �$�'D� Yr��q��5�2.ʲ2�j��s&D��"�K��|�hԊ$EL�D���!#D��Kڍ6�¼����&B hWn4��?i*OX��u>�k�.\��T�J�gir݉�B8|O�c�d�.�;X	FTrgL�8�Q�7D��!H�')���p���P�0D�Ē�+�.|!��E2�q��:D� �U���4�̺u��G<�`9Q#8D�� �4e�J� ��!#R@�	E�t��"O�%�a�6V��#��n�()�p�',��dE�.�B��ד4,�+��C�s��y��'J1Ox���a��Κ�Q�!�G����"O0tE�b�F�H�ש#���u"O^(�S�Z�3�:����4�i�"Olj�L?A�X���/nu���q"O���Аq94��u��+w���	>�r��>+f��a��Q����%�<Q�P9=��K�V��I�Ԣ�-B~)��	]~ra ���TM���c���!�y�#�fmD�@�c;���@�-���y����hW%�`H����B�y�'ɞM���'�|Pqv�I�y��f�H ���X�6���f�+��x2
� ��@P6	�>V^��&������R��'Mm
-I7��I��0�O|�=E���#���S�G���n��6p!�D	8X�q2w��}O�����!�d���8�x�+�;T�j���D�!�$B�f	Z�!���vB�4���ھ.�!�$Cr̀�^QH�T����l�d��ȓi����M�;=�v���^�����b<i&n6U@2�Y�TH-\�b�A�Px��'K�\�(O�\��H˕�4Rծ$K	�'�0���
�O�,,b��	{���"�'~����_�#�\�xQ�ųk��[�'!�Ӧ�4K�VE��%�)1�����'ܠ�D�%���G��V�`��'֎�WMB}�4,���Ք8bh���'�Dq�E�0�\�˗bQ�E���*�'\����R4Y~�
'%P�I��@��'!f��T�
���mӆ�	TZ@�p
�'�ܵb3K�S�tY������'��,�we�%q@��2-Άءr�'�D7a]*mS�K������Mg�<��捭�"��nΣM�(�*�B�dx��FxbeP�Q�*�p�d�C�4��Ь�y���-A暵@�h�K(4���NѠ�y2F���J��t��6B.�qe���y�!t�Tpqu�;���#��R�y�0�J��3d=�''���y򁕾>���6�N�/�"$�Ħ��y��)9\.( �bЦ(���є�J��hO�&�u����¥j�И����(2B}���t��p��K�������N�*!��>�z�0䯇q\,xr��	k�>|��)�65���-5����Q�<��(�ȓf�P7��a�r���_a����C�P�S��U��ń� ���ȓ\��;�"#O"t�8��9]K����s�'~�Tʱ��M���Á9v2	�'��@[���c��P�˞�1�����'=duJ�N�?�d��%�Ȓ(�fԻ�'������
H&�\�6�T�'�
E!C1��M��!ѳ3�~���'�ƀv��j�l�U�2����'��%��~Z�q��Aǐ��'t���p��1F��ܸ�
�p�ԝZ�"�'��l0Wo�	K��R�*�	@U�j�'�TI33 ,���/=� ��'����ը�$8¶H�aS2Q��'�l}�(��A{����F�+)R���'���s�
ѰL�&Ab��7�4!��� Zd���H>��$9�"�8|/�yX'"O�m��O�44@��eb75 2�#"O `�I�<%�B�!�,0�
�R`"O e��+>m-�T8�۰VB���"O�bނ(�~e�1���hD�E:B"O�aq�ᕺ*L c��!L���ac"O��٧�Y>t.HI���d�I�"O�!��F-0�A`v�J�/�d���"O�	�SE�WF $��@ ]ϔlC�"OX�t�:~"^�	���zR�xX�"O�		�Ȕf�I�ą�TD�$"O(ر��'N���h0G�m�V"O&�����3�ތ��'��5��	a"O�-զ�3~���d[>�=��"Orm@0MPT����Ɛ[�8�q��'���'��C�<Q V<���՗.�.�"O&�B4.�"d��]�N5E�\���"O����f-��ԡD�S��<�q"OQ@���-f\���}�=[A"O�ГF�ۃ-�V-1���zv�(�"OHP�E���d�	�}�LP�7"O�j$��9V��	�"������D�'���&3�|Tr��	>g��ŉ5B$k�RB�ɥ5KjarF��7�0��7�ƋME:B��(v��X��ǬUx�	
ʼ/޼B�	
e��]qA��D�l�;��M%2bB�	*JȔ��OܤD[���V�-/�C�	$9�c�a��tU˃�Z��C�I%i��l%�66��t
�c�C�I7P�(�x��1���i�e�(lC�	(z��DA�PY�M+F��s�
C䉳N8� ׏�ID^��4�L<��B��=�(`���!`	�b� c8B�	2ML�X���n��p��˛B�(��� �m�q��I�O\ĲB�I�<����$j��:p)τ&�RB�	�X{@��q���l;����D�JB�	�W%p�p��OW&!�wj��8~C��;/X����V�" ��x�&ݲ)�NC�2Z��Hʤ�29�X��� �>�dB䉄f粍��i_1|@�1��%M�JB�I2@ĈpR�x�`��N���C䉌	��C�㙎_��pG��:�O�!� ,��IZգ�*a�@!�"O,L1��H�L���j������q0"O(-�!� y�t+saU�?�`�"OBT 7A�3�9!ņ��Id���6"O� ې�Z&F�|���j|�c�"O0�+�k ��ؖmC&ji(9�"O�9�t	�%?F޸�wJY�W����"OH�!/��#�����9<�x�
�"O%kѾ�Ҁ�L_�'�B�҆"OP����~1�]rb��6d���c"O<�8�M�frP$b�7��e"1"O���2+)[Iְ�e��F�h�ic"O� ��L[�_o��v�$��y9��O.��)^.�<!��f۬4
��雑G-�'|ў�>MS �,!�<�G��G�ġ��"D�0��U�wg��inȅEx�1�W�"D���F�.5�J�Z���KoF��7 D�
�#�qvҔpAO�0��2Cm1D��a��R�N�0d��d��e:D�\ E 
�2&�ܣAe՜�Ԡ膈9��0|�S,�.p���v��*-��A1��p�<� |a��.� Y�P(m#��_,$QH�"O�e�w��~��A��	��\�X5�"O���OҀzѺ�s�I���|��E"Ou�e��J��AӶg�"�F�v"O�����^<�)�%��Pb�"O����N
�i(�R�f�� g���OȢ}
�'����fV�>v�"c��,F�V��	�'�I�e�%p�\�ڷ��R�NP	�'�`�)�6|D3mZ�S ���'F��D�X�??�$�anS� F�{�'¤Px�օe-���G6��\��'+��#ER���c�]+hh����'clL��N��at�$!�Jh�$�N>����	��}�����R/QT�����]�C�ɠ6e8�u��*'O&�oM1#uC�ɰ�:��隃Z����Ţ�'	,C�I
��$�Ԉåy6ف�1�.B�.����K�����+��� B�	�5�ޝHI8��𺧊���C䉟{/�qp	�� ���.��: C�	�g;rP)GT�<^���C�"��C�I�vH���܀V����.�:�C�	:������ ��u	�G!=��C�I1�F$��A�	\��yITA�	>�pC�		 /y�\8�BAͲ � I�"Ot$;A�Y�(�Ri��� )R�Z4(�"O�8����s��jD��S����"O�j��C��Upc��F�T�¶"Ob$@ņZ�+{���7���s�"O�p8���/�"a��a�~���f"O^ ���Yh����A1�X��"Oz�33�@	?�̨֠Πq���0"O��xe�Ӣ=����[��dH��"O�P�& K6!�f�C���'���"O���RhơD�0�%�Z{�v�r"O&�`���DE�ݐR�W����i5"O��sc��m��`��k�|�a0"O|���oH�#²6�k�V�P4"O��5��,�(Hс��![��jG"O�;�G84[jp#3�(X�Lpx�"Ox:sK[��y�Ҭ˴/���PW"O��ۖ�+He��H&aşB�HI��"O��F��
K��Ja@��-fQI�"O��ɦ��y��m!�	Tj��X�"O��Y�ϋ�7����� 5wm���4"O��J!k�5dP<��6�Ҙ o~X�'"O�����X	l����X�RWּ	e"OV�F(�	l):�yp��o8��"O4��#i� L�!I�R7���"OTܻӌ�o����R�j�"Oθ����O�Tl0E�O3M��$��"OB4y��D�@a��⓭H2]}�5��"O�l{�E�:N��T�
�Ht�"O:p�ᄮz�ֱY��ցzm����"Or|{/0C��Q�`eF�V^��"O�<i&OH�F��l��dM�Zm����"O��S��:VlN(hA�]dy*��B"O$���'?w���7c���S�"O���G��J�{�C9G��pw"O��C�l_�pQ�!E�V8P"O|�4D��1[�m0��>G�l\�"OHL�D�2I0N��e(Z<6����"O"@�I֨0c�0�G�5�2͛�"Oj�Ó�S(_��|�g薌}�j��b"O� ̼ہC��@�����P���5"O�erc+��H,�h��nuf�;"Ob�(G*Z�B�!SG�;v��H�&"O4RB�B�v?xT+wa�)N��E9�"O~]�u��<B �@�B�����e��"O��%�K�J��5�@��s���"OR�ò�ͺ�V#�$ٙ'��T�"O�1p5([F�Q3R���!�bh5"O�8f���v����^�2�fL3B"O�a�$E�u��H��P0c{�9�"OB;�B�I�^ ���A�|n!�`"O�]*&�&W���!�F7|���T"Ot���ڗlT]yJ�	_���"O���`����sv��g~ʈ	!"O,�ꡧX3���`�5fdi!"O��ӡ�<
������0�"OHp�7��,m,��KDa�
2���"OF��%)r� �bn�_!��r"O�Ea2��/���pHѵV<�k�"O��ggĥR�y��T00�8ل"OR��!��uK�aR�2� ��"OLPiG�K/>��1�v��h{1"OZ�+c��(.�x� r ��-��yc"O���׆��tq�H/%i܉B"O,}��O�0��Aݸ:b��"O��&ˇ.**��X�Nx��8
P"O����bP�R��$���9R�[T"O��:$��8�`��nRE&�B�"O���V'��C�vY�6LY/Yjir�"O4p�2�� ���&Ő>�rM��"Oʁ	B��)��f؛�����"O����m�*4%��Qr��D"O`�%��>;�(�)��q|MQC"O�t[��pe�lZ�Bap�b"O��qI)A L�bR�A�5YNpI"O�	�@�Ψ[���p�		�`P�<3"O�4k܄�(�(�M�:$s�"O$�P*ˆ\��#6�;g"�Z7"O��Cb�f�4��)���"Oh]:�bB�u���@��4)z�\��"O�E�iH=(XHXD$�w���"O �Q��ԥ`�d�Z�BWor�3'"O���A9e�(Q��Ã[Eę*�"Or �AJ��xIk2b�>���1"O� K��܊dvFUS���Z�
�Q�"O��{A�G�
�R7 6aXݓc"O�@I�'V�fn8|��h�fCh�Y&"O�i
��̨<��!���'���8E"O.(��ƙ�q	͓t�ZM25mV�<��)Wg�
��'Iy �i*Q�KG�<Y��dۂ�H'̖�`� j�CJ�<	A`ѕ�L��0�{� A!ƌ�I�<	׎�	<�p�Y`J�h���pR�WP�<��j%'F�a���6<�p$�A�c�<��ެ5Ta���ư*Or����^�<���2*�<#��Іq�0���]�<-4D�x������E��>��݅� .�� U��=3��K �=l� }�ȓ9C���p�v ^�'	=*`~���z&���ꀠI�8���T��5��`����F&������1>I�ȓf۬�I�Ý8S�YX�M��3�l̆�4Y5��g�Q�@�U
��P�ȓ^(e��l�>A��K!��|v����S�? H%j�_12��Ǯ=g8<�!"Ova�%.M&QHdm�&~�`�"Of9��$̹n[�[���5&�\4��"O�,!�,��x�\�r��Ou����"Oh���C�+�(1����-Ga��"OĜ�(�3@r\��f!1?,Q��"O�)��S
���B�.k�y� �H>�y� [�i|�@�#�ɳ1 �1(��B��y�-׆"Jv-��&�%#��a�g�$�y��H�9E���=�@�2e ���y��Y�j	��r���&4ZD�4�y��Υ*48���̷M8ӆ����y�� -s��r�Rx����fl*�y�h[@�"��?f=}1�͘��PyҬX��"�/��+v����}�<QcC��v�.}��W �|�7e�<�P�.�LH�aԙ4s��X�z�<�b��@(�5Ca�`�ؼ�0�s�<QFA�f�����4���T�l�<�sc�]�
,�7e�6@Le;"�D�<aר�o�t���/G{����x�<	C�r�0�S�A�)ɨ��o�N�<�-Όa��dإ`�	!^)�w��L�<Ad�U.6C"`r iO,zL��͡"O��K�)��X�T���\�{���;3"O���.8JM�a�QA����4"O@t#6M���e���y㴅3�"O$P qb��d���&g��3�"Ox�"�NXq����c� 8N�`��"O�ع�O�f�V�Iv��:s0N��"OQ�����_� ���4&��@2�"OBb�L��ʎ��s%�y�ДA�"O�AW�K=��$1��V���#u"O~��2�W�$^���*�F])�"O����C&+���x3&�Q���2"O&tBJ�@�\�����d�� "OAc�DS�vD�a�����zYj��"OR����2W,�r6i�6}tŘ�"O��H���;�������/Q��|�6"O�@�e��/d <9PN��W�^%pf"O<{���25�Pa!��+���"O�m��ބQ ݛ���	;@"Oɛ�e�"z��nȳ;$�
.D�L!Rh^�
���J�I���"� *D����N�$V����i�8Y}��R,D�P���?^�$yA�L�YK��i�h/D��q�� ;|P%cPJ�"A|1Bƃ!D��S�"�7ό����
�~䙲!!D���G�R��X��o@�_��P�M2D��)��3bB��:�X�'
��s�<D�4��	��`�=J�.�F����҇0D�h��
�9���0%��f$�jP�:D�l 7i�fY��D'}�"��
8D�x�w
[�9�d�#��V�X��B�2D���%�,.R�9x3���BD�%D��A!F�e8Lm;�ܳNJ�P�*7D��[W��*V]��	?$y�f4D��c����
�h�ԇz�BHS�0D���L�nf��C�)g>0�9D�xI4M�(�ZQ%!4�4Ԡ�);D�L�u�>l=^9�T��<:��=D��ფ��`����參#OV�B��;D���yz��G�+m�P��Z!=�!�AT�n�bA�H�F�`�G�k�!�� l��$8�؀H�I�u
x��G"O�yزl�L�b�2cbŨ\�lXZ�"O�	ڂǐ/5���K�NU�����"ORㆉ
�\�#��9�Zq��"OP�i�Z�N���{fၜ2��8�"O� �reW5d��`�2 ��ə""O�8@���7_����:/n�IQ"O�����I4)s>T��D�Up�"OT�Pb)��p��`s%��).���b�"OZ���^�^A @â��]>µ`�"O��-A7���sdj^�;>.L�#"OZ�x&%ֿ"(�UH�Ց!�u��"O�� r"܋,w�!�b:a2""O���;z��AhC@�+'hHy��"O�	Ñ@H&C���YGl� (7"O��	>Xx�ݩ�
,V�!�"O��@%�}�l�2ǩ�H����%"O2iѓ
�QdrHo� y���"Ohتk���`�Sad�xcB"O�� !��C��=����)y$����"O�1�v��"TO�X�EƟ8���"O��x�O�=P+�-��d�NS��#�"O�K�I�U�Yb��6W�XPA"O�yC�m��}�Y9�C0f�̐�"OP�Mu�.������D�!�O$A��	��=�n�R�=0�!�ćŶl�(=��Lz���c+!�dO�|��0Y��A�\�$�U�ڮ7!�DP�Yf~HYB��L�����*|�!���-ͮ���ڹ5��C7韷4�!�$�#Vޔʶ	@�������q�!�d�9����NE���GXy���ȓk�çG�k���sUF�3~v0��^@� �Қp@��2��N���by����L˽eh���b�t�h�ȓ,2X-���K4�F�t���@W�=�ȓ�x�f%�in�1D1��1�H ��C�MXz0gb����ȓs�����T��s�_:Q�漆ȓ��Q:"�GE&�JSL�Wl�	����9�aBH;�v�j D3uGJl��(3�U���Q(	*ʄ���j'�,�ȓ6�T:�P�v6L�aAD؉�����ma��1��ĥ�L� �⓯k���ȓ3��UYT�E�jr���l"aI�ȓHu�����b�r�@Ճ� An6�ȓ�tC���&��,�6��%����iJ����p����#@�8�ȓ*�{q%�
(�X�Y�,Ҋg��ȓDؔ�fG��9o��	�I�w���ȓ2�L��#"Ҩ]���#� (��1��q�I�b�
�6NZ�]Q��y�H�j�4e
BIX�@��i�%���y��M.bI���IΑ6��l;�MU��y�B�?8��E0��0Y0��_��Py���& ̌�U��!<82d��k�<����t�R\�v���h��H�H�@�<�.��yM(�	$H�f	ԍ����<QD��7d����7](=��MxG��<a�9P���a ��3�XM���<��@�bZ��ڶ�~:� 8�Ib�<��7�f5y"�ʆ�``�w��C�<ك��z���UF_)f�����B�<��OI�S?Ftz�$�����( �<� �2���7"{���-5��ɘD"O�5�%M��yk�Ey�픱}����"Op�XQw���0��7�P�зCK�<� �63&F��+��F�X�+^F�<����6+KP��%ʱv��j��SC�<A���`�ܨP0��-B�Q���x�<yu`ǵ65�8;�k�7ozpr�s�<��բ.�^h:@"��x�z%��F	p�<�N�8#�
�a���qK>P)C�Pl�<qQ
S�&�>���
*(�F(AT��e�<a�䔬h�N,ӲKN�k��5j���x�<YQ◈TvL#vO�0�t���J�<y�hY�0f�0E+?ɰ��s�_�<��":�~y�6jT�9�1c��B�<y�ћ5�����?{�:CD�RI�<Q`�זs09h��ۻc�Z�cJ�<	�)jG(��Ĥ�[`��M�E�<A��^�r%��j�$`̦��
Cx�<�$�P�7�űwGCJ@�	:��t�<qe �>2l�����/j�1!��q�<�b���=�L���F�	æ�I^G�<a��I)pr7j�2C���;"�Hz�<A��� �P!���{@|���y�<Y�/�$ ��Q�((6�p��
Ns�<��`� (����2X؊z�<���ѻ>��� V����A.q�<)�nۚ$�@�#���:3�=�2"Ml�<��J M �K�
�1]j�C%�j�<���04BD��qՑ`��t�w��d8�,Dz��P9S��|:����HMr�Z�D9����]ןlhbH>u�X��Gğ�gL�d�0D���rb	!V��"$H\=+��I�#"����Ԉ�qfVn�8U"7Y���)��d$�S�4m�4�+��м��x��N�Q�&c��:��)�ɞ�T��lK��G�\�\A��Q���	�,�F����������G�18~��=a	ç2kR��Wk�9S�捹��ʖth���In�j\��3���q�u	��N7��X	�'2�-P%bB��Y��/�:�

�'�,%Iu�ݻN �L�pI�,W����'�XC�d��@rXq�w�D5q���'a`,�Q���F�$���D!f�'z�b�6+�����((b��Ó�hO��ە�T�b��z��C����"O�Ԑv���?^��k@�.��䁰�'��O�q�5cW�4�ha���lk'"O���DD�"A��@-��(��L���d#�S�'Or����AŊ+�F����H��@��t�	�v��)��M�=nL�ѪIkQTC�	C�٪j� +���bh�:v�0�Ў}�9O?��@�4<$a: �P0��!���'��|B [�O�$��-]�q��,A�� �M��""�O��ɮu(���q�P%����q�B���B�	�0�VXXbFH�n<����*oK�"<�ϓ|���*�� �A�2�ߓ/tJ�?����~��.0�Z��`��'���ŦJ�<q��a��p҇%�Q,�)C��H�'xa��ۓRt�ؚ�ѧ<��L�%�H��yr���z���g�9��r%㊔����i2�g?ٴLǮ	xP�𓭞�Qr��Lb�<ף�.Z���!U�W�xQ{iߟ���a:
����Qv�`� a�=E�
܅��*Oje����#�%K��(5��"O�����x`f�V�;��h�p��P���� JTa� «A�*h��._T��$��"O8�)Bn�k��4 3��)/��ps"O
%��2E��ё"�H����B"O�I hä{|�k�G�/~Ɯk�"O*��f^j#%�%M�jaV� 4"O���!Ē�A�b�H�!Z�J`~�Cd"O�AC�.���Ph��6cHm�!Z����	�H`��%dM:��E+N3<C�1*�l@Z�c&^��Ȣ��O( C�ɪ%9֙Bs`�f_�l3�D(>��B�I4h�vm3��9,�9Hÿ9T�B�I�d��k�<I����
���B�I!�p9zs%�P��8�C��iТB��3
>>dh��g�֥A�EL�>q,C�	�/��B�L��Y�A�%a�B�I?m�Xӕ��(K�>�1ҍ1�B�Ik0xs����< 0��"�*�B�I�@0���ҫ�vɸU2DJ =+"B�	�I%���W�dӔ���+Ӻ"WVB�ɯT����6���R,4�2B�I:#p�[Ǥ�>T	P'-�F#=q��T?MYЎ�6�`�3�G��j�脋�-3D���B �V>�;eg�2����b0D�� v��I�&iX�)\�%�����-D�l�C�S>
�HVC�#mZճ��,��G�� ����54
5��H�P}���$�p���Do~P�Œ�Y�	H��Q�C�VB�	=k�3�	^2$jr�䏣��B�	+E�� ��% �Lp��K�!e B䉚2�$EK�C]�$��S��h�B�	&FU8,"4���Ph�W	�"��C�Iu ��k����[�f�l���'�b�9 ��L�"=Iq�͐z@�k�'e�Z�����,�`g�M6zAJ0:��d!O�8��Aӕ|Y҅�vh�21�Ri;��'���I-.�� 
�;}<�CЭۃX7�*��T+�'pU��Aa�4v��Ij�,*��m��>��]�jh��I�l�)��#D�8���-{�d�sD�H�c�K�
!�DH9 X$�1�I�C�U ��[Z��p��H�J����N	=a��i�g�-R~MHv"O�Q�ƾ��{�@ç6\�!#�x2�i�'��)��@>C(���'t�9����;�!��ɦ�X�Z��޲�t�L+�Q�Ѕ�I2c����`���Cd�� �nC��#2������Q�vACtc^�Q�6�F{J?p㟅-d�T;��Y5.�pu0D���ɢ ��	�YlY0��*�I�P��}���j�݊��9��D۾vN�㟨���5C��)!�͘5�niY��5N)�O�3eO�R��z�I�&�
����'�
�1�y�b��o���W�̏K�Ȉӥ���y�G18b�K��ՐAxU�t�����hOq�:u��ܽ	�b�q�߾E�Bds�1OX�	X�S�O��s4gHG���7��:d�	�'���SL��e�Ec��+R4]r�y���żE��aR�CA�3Y���g���g�!�D �3�Rܨ�E��iMȭ�vE�&���	�O��?e�vΌ�Y%z ��Ƿk`J�['�+�O Onq�1!�#/z`: ㈅e*�@���LE{���ʵL���`e)�51��c�
�!�D1��|�0��>�ɔB�,[�!�"8���^	5!"h�s G�Q�xD{���'� ���� ��;�`N�0ؐ��� ��ϟ�ٰ΋8�p���OD��d�:U��у5L >b,0������!�Fc�"���
�hd�y$gM�/r!��N�#���gc�el89"�F�$b!��P�Z��w�
Y�DRpD^�8Q!�$P�-����G]�t,�Cs�R.,�!�D��d�xx�%��d��9��`8A"OHm9�&^&|��0!%1w��#�"O�Y�GZ�%V�<��cҡ �-��"OJ`5�,WuF��c��rwĔ���d<|O�T2@��n#��D���ZrL��'|�O�I�q����U挓?tz<��"Oƀ����CJv��*~bD�1A"O�Dj�;{ŸE"OU6�U��"O�A2�ܠ8���dҖ���e�O���$�[����"π�hp6�]�i�!�GCh�RG���H��4�^&Gl�O���d_*N���Zv�7C�n��򩀏Pf�zb�$�~<�*��\����.$k!�$]�8Y���1�&�a!.�h^�'���)�S}C��h��C��>9�W�L�g4ZC�
qc� )ۢ-�(�f�I�NB�u͂4��]fi.0�c'F�U��B�I)N����)J3R�d[IrB�I�dIb����
p����B�Ɋ��}����v�zKJB� SB)r���+1�\��a�8?�C�I�V���⇆Ғ/p�1�>6M�B�I�4���V�@5Y���.B��6�2�S��M����Dհ,��a�# ��rS�l�<��%��G�r�:ѣ؆5�Z�{�FR}"�O ��DQ)E}�$�&��zZ`9d�	B!�nq�A�G��+)���(��L5b$!��}�E�/�@E2�eƁ!�ҖwI�T��E�2��:p��#v!��U�O���XV͑8�
i���0t!�]o��ЄMV�37�$�a�Z(�!�$F=~�]�p+��I�L���
B��!�	7�r@D�͑&��i�ə�!�� 	$�(Y��愪l��@�U)XF�!�C9-�DL���N�Pp�M�#o�|[!�DO�*�I83�6hl���5T�!��S���	C�.M`<����,�!�l����/K"D+�4S�g�B�!��B2u��x�wŃ�I�~�# ݼ!���,J������$k��N�)!�$�M� ��`�޵o�V����f4!�-7IС�F˛�s��\1r$]�^�!�C-�tXk4#�o߼���"�!�$�Ht$�{��C�1k M0 �V�z!�ӕ��5���B�Q�d`�4��=#�!�dҝ(���bۚX�H�1�"O �y��^L
 �2w�M���S"Ot:AN�Z<&�:��ȑx�J�W"OX�A$�M�cBd���%
96�� �"OH�L�=	�|@�d��3�M�d"O�4`#�N�W��\����(Ft��"O`��˪G���wɋ�QZrIX�"O�}R@��[|D�ZD��K��A�"O�Ert%ÜQ����	�&?4�c`"O�j
�Q�<�����X,�"O��ړ�D)J��]��'A&Jx��b�"O4u��D��t�%�p�ƽ\j�ت"O�5 Q��+p��6����0��"O� �h�CBҚ( �Fƞ�A�%�4"O�]�@f8y���ǯ5�D�p"O��Ӎ޼V�P5he�Ѝg�JP�"O@�e��1&,%"  �P6��87�'��y����On�c��Ʈl��2'H�#=[NK������'7a�é� x�m��c��f�!�'�)���;&y80L�a2(�'�\�a��e`d GDƢ��ȡ�'��-b�)F�cfp�v'Z�Elmb
�'�	0�O�f����g�"����'�����IzQA���f��1�'�8a@ ²>�\��%�K�I���'v�Ag͔Z��[P!�:���'����Ed4��ǣa�� ��'�� P�#R���z�*�\�l��'�"I��-�"P�e�V�|Y��'�:�³8U_�Ȑ̍�L�D���')H��<'u�5R��
m���UD>D�@{��p��yk�dB9ʍ0$;D�T�%&Y0��, r��/m��H��
$D��%��
$U=�ue�"f�l0*W�(D�x������&�@WB�=ʈE���'D�z�G8l�����*t�����0D��
%E�X�4�I4(D�J��h1e,D�Hj�HǉfwzTɂ!f�n�0�/D��� �ě��d��C�VFpE���*D�W�,v�2=�p͓�2 H%b�@)D�����
�Y�dU��Q�t�� ��&D���MEa�	I@#et��Ȓ�%<O�Y" �#dv��]�6��O.�pd�'c�:�t���y�y!TT�8
b5y���A�*�$��z��E��(E�1�S�����Cᙃ5<(�B"�^�8�C�I�'2�΂�`#D��k-�����>���������L>Q�NK8_���l���A{�
�(<q��&+S&�;���ZL����h�t�I�%�� \��{%n����\(=H�D�@nA�Y�B��>p������ �l�'߾e��on�P��ׄ"H��r�'�X]p��C�?E�l�7"�U�"��K����/E��,uu�k�OC.�#�!�!�����aˁG�*�'���&��"@����` /'�[���*l':˓ �� C��8�3�S*�H�h=RP|Q  �R��d��Uq�]H���N`D���:�.m��X��
��D$�O��@t�U(a���#0��¥q��'���K�o ,>h�V���o�R�HCP�ϰ?oH���.D�����K[U��c�G<Z��]U#�䐏z��Q�V*����$yaD˓�n4���^<A�D�U"O��`��6c<L��/��y��X��	��'x��H���>1��I�~\��� �:�<����Z�<��՗?� 	�g�N���W��~�<	B�^KD|8֭�DziPK�~�<91�]b�$����E(1�u�<���ݦ��y傄���"�n�<����%��D�D �6d	��n�<�4�ŷV����)R�W��J'��M�<�Z�Q��ZqNH� Mn�
��s�<�EeZ�4g6ѺkߵD[HҡLJp�<��ǵr�\�IvE$R%hرvm�<q��WI���`L�qt�����j�<��ӑ=�!�3"� �2��ЫR}�<���@
��S����wm�[�Hv�<��閜dV��*�L�:��U��[�<�ۂ C������|g��RK�m�<	 �ՉM<� �5�^�@IޜH�
B�<�U�C!#7���4#Y� #�R�<� ŋ����K�� c��D�4f"O�MbPo�5#�8ٙw���&�\��W"O숹u�Ǝ)�D\A�ӎX��e��"O�Q���n,�� �!�:��"O6Y[QHE=󴉱���|r\{�"OƁ��B��P�Bn��TR�"O�ݪ�A�DXh���{�4�"O�I!d*J:O�L��Up��W"O����+I���˓lD�"dh(�"O�DK&��(zhT���ƻ��)v"O�PPk4R�� "J��h3"O-���SqӺ '��"��K��!�DP	P��5(h�b������8�!�DG��h�`5���QةkgFW qs!�M0w-xyr&��w�\Ѫ�e2k!�DY>�8|s�d��\�JE։Olb�{��Ԅa��p�'yJ��F�җ]w�����;�
�B�'%�4C��9�h&�	>=�<Tc�}���҄ ��pR�ؑv��?q��Q���0(��C��
P�j��*U͗U"Dy��$]�S�,�fɀ�S�x1X�Oأ|�'���ǡ>c��2P�ϲP7:���'\t�u!�2
�\� 	̰_XH�ҀE�]f�q# Ȕ	����ŔP8��hv	%b�>�� �M�Rn���f(\O2TR�*�]m�1RB�?[�0��%F{l���� ~���%���x�%(_A���� �NM,�!K�)��' ���%��*vJ�J�Ƶ,�|�|R�c�g�R�ڧ�G!01����ZX�<�� _f��<�F!S�S��ac1CȚ- �16��h*uj�o�61��E�,O8�ACT�p'�����1��C�"O4P.�$1ǈ�0�jT�������2`BӌI��R�R�l�J�axR�E-v�	b&��:�JY�����p<�Y�c�v��R�Z���������'�K�bM.��s��!�����-�P���@�A�����"~i���;?!���G��(���6hpH���67XHT�|Rp�H72�֤��Q�X��E��r�<�1��3r��5��$oj�\xv
H�q�53wk2=�n\چ�J�b����|���
G~,��,���e�Cˀ�2�6�xB�R8+b��g�
|Njt�C��m���Ф��my���5�q�s�'؂v�H"}�:�3L�e�Xm��b@�㥩-?��-i�Z���$H�q��	s&�;KJM�&�%$���Gh�0$��k���SQ��xQ�=?	�Dч���"|ڂI�??����g�DK��\�<iw �8Ze#�n�1ǘٚ��Cܓb�d�j
˓ּ���`u���S�A���0�ȓ:+��h"+�?An�K���1�HŅȓ>n���aP3r2���F�vNɅȓ=5rMB�kw�DIk���>�Z��ȓy%������ ������� 	.h�ȓF���҆�8������T�ҥ��-ƨKd�ܠ�B�7�U�_2�ȓs	����H��@i?
4T���-2N ˑmZ�{��))2h9Jtƈ�ȓ[6�a�C��/�p��)_:��݆�*i"���g�#L���!'�;1�-��(�Q+�Oތ%��Ed�+�T�ȓQ��8 �z�i+Я�c*�Y�ȓeN�H�N:DRx�zC�Ȅ���G}R���%퀥G���ط6ۊ���=/��m �&Է�yr�^�� ��J  	���cT�y���/����|��IΠW�\cĉ¤=�T�F��A�!�d��ɡ���]�޵��ʔ���$�R���S����<�L�}]x����L#�L�bEHqx��BwE�3���1��SӎiPlE����TQ!��~�f�1Q�S�#����Ɇ9[�ўl�2�޸rXȴ��&N ^��P?z���[Q�T�#�!�K-nv`r@fB%v����iټXB���'h8� �^��F�? �qS��&Ͷ˥̟�x����"Ol�A/A<3�����+N���R�l#t�F�y�,I
��'��C�d�9&�V�I%E��:{��a	M�c�wΠ9�t"J�*����W�bИ8��SH<���ɲ���RF��m�&Y�� �|�'�=Y<4����~r�,�91���z�旕@^�p7��W�<)F)�=zV�Zpf_����<у�/b.��M>E�����$����ռ2�b� N
��Py�&B��:���m'|�FAm�d��*�J���,�����vک8Q)K=#n�� ZZ�����J�*ɑB���c���ȓ�ztI�t{��1!);8���'p��a��d�S�O(
`z�DM-�^����̇ct���'���8{=
��N�5��D�O<1VKݧRn\a���=:v#[i�TtRa
6��TG�X�mo�ɖ'��@�Am"�9�D:t�j�͖����Љ�s<�0)G��HW���3�I��_}�9��0n�<�TɃ!Dk0�	0�vڒIi����Q\�P���3a�B䉋?�J�#H0�j���o>����i�zY�f�10����� Q�)�)Xin���O�=���7D#���4��Mbe8��'Fi�VH	= ���@�`�	g[� �e��g* �A�ȉ%B�x���UP�(֢R^���+A��%���B0o�\�*��#�Q��8`ڀZ+$���E�c�6�au��58\b�եY �����6q��e&�l���ɚ����'�S4z2��L����u��6�����aߑeְ�q�d̋^�z�3��)�^��m�g�*)�La���'(�!�����)Z� %"C�R%V�����i�TE�\R�"5�8u"Ř?��RD��Gh0�?fX�"$.L�r��dF�'$�x)���P��ac�U�x�<�����j�ƇDNx��'�By����`kyBD��'�\ѐ�\"l DU�&��&Zd=R��d��'R8xbHڊT^�m��I×[�-X��r�&QD�������7m�4)�'y��R�g^�k?x�A@K���i��%zv��>���Ti�e|��2'_�h;|�>)i�&��.�
Pir�Z�9ޝ*1�@j�<�q��]�\!y���N@��Rh�~P�5�TPu��P`dU�/�|��OIX�Q��Q�	�v��� ��F�J<�Ѫ�$�v���$�x�:'�2r�v�б`�p� RB���@[����8�##�.-(	�c'z�'%�*QV �ǟ1��4G{¬�F�aQp*�Rك�ǌ76����a�O��$a#VY6z�b�3я� ����ē�:�2D�f+�M���c�2��	�RD��+&�6!�=h�.�+}�*�b�D��d)q�r�3�U� ZR1C(�	|<�	P�3D�4a)��6�\\��ƁE�H�v�!��MB3	��[mnt�An||˧U`��`0��*8Z��ċ�,�\�O_	�a~�ψTR�p�B��Pf( ����x����q*�A�f�����P(׊/�y�Y&}��#���[KbY)�߬�O�)��OלPj��2��ɭ)����u��M���5"X�|b��sM�#Q��BU"O,�:�ҥ7���碅'�pe[�O,�Y'��>*�$��*�N#"�P� ��q��6U��S�(�R�<��hő~��"�M�4@�sSBA
H�P���'�QC���5 ����On���3%ʵ�d��;�����'�0��N� )�X��A��|�=�p횱8�4�*�"H)v���	5E��2�4"�t�K�E��-���D��1���"��I/��p�OI<v�zHc���6ZF�C��%S
�I��Qv2���C�<V�DOf83էN�����OV`�8��[�����Y8s݀���'� PQ���;:�\E{W���c�,���'��� %��K���P��!�i
�'!|�A���õl�!v�d�
�'�
5.�V�D����s�`P��G�L@)JA���;s��0���l=�2fnR�5�F<���oG��ȓZv.Q�h
B�,=���V� �ތ�ȓ@J��̛a��q�'�F�S|t��"����gD�Jz���U�RU��ȅȓR�]81+��C(��e�r�݅ȓ.�X�#���e��B�c^�A��S�? "�&ζH��42�*ٽs�`�S"O^�K�ꖋ@ծ@׈	'���Z�"O�����(e��1C&���Je���"Oʼ9��7B|.2g�C�k��)V"O�����8Ya:��KB�+�Ju"O$�Z���3�R,��Q7�n��`"O�2Ɯ�,;P)��?n����"O��8I<?n�DC��@(N:r]*�"O`�b��<�}֊@`�B"O\��B��$�0[�wz2}�%"O^�ae /�R��2g�7We�	�"O~���/Z z~0�f���� �"O�̳Bٜ|ْ02$�2]�F��"O��Y���c��9��AY�U��H�R"Oa:c̀=�����VP�.ě�"O�cC��n\�� ����d"Oީ(�.N�*�8�EI1�;�"O��"p�־Uru*�M	!�T �w"Or`p�K��S�r�����,��0"O�yJ����1E�E��&�u�T��"OU�1�H!~`�M�n��\�A�"OJܚ��
|������7��2'"O��Hah�0j�n˽s���R�"O� 1R"���m���"O��G�:�D�AՎ�:��`Sq"Ol԰-1�^�!��Sac<��"O^���L��l! b�G��0�"O� *��ؤ��^�N��-�p"OF�	۬bZ����3�L�i"O(�r��9s��)%*���a�"O֭rY?\�(��1�l���"O���
��  �'u(��r6"OL� S �0%��0.r��'�  C�1/�I�`r�p�T �:t�R��
V�q�C�0Q�Ц���j:��B�)[�O�|haH�)Q�����*B&@Q�F�*]-�X!���nW!�DY��ȉ �M=6`0��iG,\�9���Hy�쟦�Vl�}&��"��̝����F�,��0T,-��k��GѮ���l�~e5i��ɒY�)��[�+��)��ɚ<"%v�OY����ڀUI�����<|�$�ʊiR�J%<m��Z�8ZM�G�2sG��ȓ#Fܸ�`�̴a� u$E,��<�O6,��j��^=xAA"�(�'a���!�&:^�)ڗ�~<V��P���/G�u�$hۡ��y�v�bu
_�m��		q�i����|���=;�����͗�`�6m��`��PxBg�4���
�+��X��.�7_T�	S�
�;ʼ���'�
 F����|�D�)=�����kl(3�Aד
�����O,L{���3V�D����"(R�0�"O�HƎ�Gx6@j�➡t���xżA&(���GW�OI��bPc�d��)�p�\�,hԅ��'�  k���yn,-[�U"_T�!pH�0��"]P�1��L����K�M<je����g��5�@5D����+')~���`A�{�e)��)D�����S%6��ȱjC+x,��"� &D����߄q���cd�@�T��Q�2D�\�A.� T�po_��=��A.D���� ��q�l��u��	�ѩ/D������-��$��!��-�q/ D�x�h� v?��$��0��S�!D��(�,��N�&�q��4X�I{q<D�t�� �!Dx�ڷ(^)I�f����.D��yV�
)Ł��|.��`)-D��a���)3�L�jE�П7�8��(D���FhS���X�5�+ٴ����&D�� �T�Q�ĝbǄ���'E>K[�U�"OⰘ ��-w(@`:C �h��kb"O敹�ŏ�
��Y��7�zIQ"O.�����'�8����83��8P�"O2�ɐ��f_i�bغ{�@��q"OtIk�͜9�.5Zs�߄��yI#"OF�Ҳ�ǙhI�Q� ��0JтY�"O�@)�D���YX��U }�5SR"O���E����^�Ha�y"OX؁� �Z�IP�j�>]F����"O�pv�H������g[Y�l�"Or�h��'ZD)�a�Q*�	 q"O��Q�W�,b06,H�g��;"O�Qi5+�l�Y��Ał[���j$"Oj��D�
n$.L�1ƒr:�kQ"Ob<�tΜ%��U�҃ rcFh�"O��q��PE" �8,ϳJd
p�7"O!h��]�-pHi�e,E��^���"O<P�B�]�d&L@��Q�c8.<`�"O�P$.��[�LH����o6X����'���F�M}���5^�b�'��Ea�<�y���N~��zRAB��-y�.��'JZ�i�k
NQ?�W�L�� ���Q�-KP��!�He8 2Ԥ_|ڹ�GnX�W��d�$FC#BL�����۟�j��<y�,687�H��.�W�tp���o�<�B��f9��C �SO�QI�m ),Fb� 6c�>@Ȉ��\�v���D�M�~�@��:����=8��z"cC�`r�3��'B89��_3;ת���)|3�� �C]�?�1��g�D������/7�]�G�?̪4�=1i`Z�+u�<9Ϡ\�q�2�Ӯd�>P�g�G�/�䐠P�A�s��B�I�q%������9n�P�W�\,2�mx��j�T�s!F��~���2q�:�gyeN#T����f��;6��
�y��F��A"�kȹO_6���	�U!lQd
�&7����T��V6��J���a��#Y�\&&Ź�n��,uj؅�ɉHt"���q|�[F%Ҿ�zX��B�RB�i�ΟR�6��0O��J3��m�H1c3&��mc����>x�mb�Md���EL�'U���Kr%٠!i�5* 2V��ȓAG�{�F\����s�Ѭy8.�	T��Vj���聙?R��	Z��~r�Y��ic�5f�y���:�y��I�X�,��A�)��ڃ-�8�ē2Q����$�p<)a(R<�R�t�ԕw�胦'R��$9Ah�Qx��ɡ+��Q�&�%/U;�4�O��D�O!"�t5r �&\��0��"O`� ��] ~�`��t�t��"OT� �1c ����̡�"O�,Q��B�n��7�WZ�(d��"OBX�R,T� P�	�b!
��� �"O��2bb�/)H�c�]:�4� "O���@!J� ���:h��!��"O�H%B��j�D8�DBÂya�1%"O:Qs��:7օZBh]*HVvUr"Ob�r��@�PyقJ� Li�@"O^�֫�0���J�B�ձF"O��2�$��I��)BC:���a"OPH�I�*q���υ��5��"O>]r�_�e�t Ë9���if"O���i6FZ$��OL?��X�"O�Th@��l� e�VΖ)\��"O�HYDi��Hx��J(p� t�ɔD�r�P��$}d���� �b��􆕅oZ�B�I"P
-'��0�����ҸRqP�2pv`d!s�a�)�s_�-x��ڑp1��
�`5Jq�ȓR���j�ϔ�7�S���ɗ'Mr(c��L�2���	�?^l��K;�� �f'�v0��d�u8٪w#%� ���f*�4K�M���E+C
�!@YZH<1�e8�DhÏY�ΦQ�JG|�'�Fx��O"����~�t�V!Ӭ��_=�((R�<yѣG9�h ���P�Jކ	؀&����+���I���ĝ>E�Tn@�n�űb��i;�U��FY�G!�ވ��E�C��8;��]��I�_#�2"�I�uWay�J�0a�ZX`�A^*<�lY�ϱ��>IRFϳ}��(#֬ũ6�xt��h�bOҗ*�^B�ɧV-Z�K1��
<���$�Ң=A�	�
�\Tۗ"/�ӳ1~� ��' �c��!�% �N��B��a�\�(���g��- �6 '�扈)jLSJ�b�)�u���d��@-��K�<i9R���GoB-�f��S�܂�%�<~80�O<�%�ˢ�0=	Q�ڄG����?>�k���a�<��mN�{����Z� jR��N�X�<)P�̣$(�Mq*O�B+��r�h�By"���=���=E����4��mҐ�O:Y���	5mM��y�G�xf��c�B�T�J�+T�����4����(��p<��!X�e�3���5:ޱ�r��|�'�y3P�fyb��=�I�g4}�ЁJ6o�$JQ�@a�1BzRE��W�Й�dG	<��2Ӡ�7a�*��'9N���f��L��'v *��N&6�1����(A�m�YaGW �P�"O�C�$7\Zr eL*�j1��O���2㑃,o�X�4+Q��� U�x���� r���2r��PbJJZ�8�P�K/�O��⃈ı6� ���)�,{.�H��Os֥8����~��Җ{.f����EA�$�"E[|� �Kd��9`�����?�,W�}�7�?G�N�IV�X�b-�zČ����1=���e �*4�݀gO���p.�l�Q�aY@"S�Ot�KA�B�a�T��'~���'C	+L4�|�U��s� -�D�֑.����r�~�<��6tȸ�"%��7y��H u�~?I�E�����+V�+P���Oba��G~BH�9J�!���m�21�`�p?�G#p�<e;�O�"���Ȁ�'k��5)fX� ���	���e��I]�c7�x�C�;:�<��B
�R�(�GJ�٨O���((���R~������8z^�1�`�$hb0� �֚T��aÅ�%$��K�jQ���ѯ]�I.���3�>d/�	|��Ez�'zƽhڊE�B��~�h�,� )�u�FN-E�^�<�0�޴A��)�Gf�&\äx���۟D34L�1hbq�5
'@Y��?m��xrdC`�>LR#ǀ�7Ӡ8��g���y�@ϋ`h!�A \%Y�3@2���F�j� ĥ���<�!�]�s�!�c�-�ш¯�}x�ؠ��>n���`�D>N�㥋�BX�@A�G�	�!�&�������;�M2��
6�ў��扆�=�v�HE��ү,���q҂��U�ID�.J�ȓ��)&aǨE�(pOޥ_ ���ɲ`z�b!d����S�O�d* �K75ι�3B��(��l�@"O�IC�"	5>��If��<vR�ݓe��8�l�{�l��	=E�l�K�j��G ����˥
x��������e�,?$�,c��ʑsޮ�S%����y�lG�|���+7�k�y�P��y��e�B�L�l}�3��PyR��R�
��؛k��E����D�<�� պ`EP`�MH{�����DD�<�A��0@X��{�I�b=.�rx�<Q$���1�ؙ*q�҈tMDh���\�<1s)��3f�J�2jP٣�Z�<��AO�x�-A���6�#� �]�<�&�+H�"I�sJTz]4r��LY�<�A�ѱ{`� q�юK-��a���P�<A �ԲR��Ua�ۃ�h�E�Q�<)�OI�?|4����̼\W���@$NS�<ᔣ��Là�;�c�`�@� 1C�N�<�p��{󖉙O�z4
ui�D�<�f��cc���3eC��t�7�I@�<A��1��ƃU�>�~�B���Y�<� �AQ'+�L���k[��T3�"O�c#-��Y��"Ej2X�'"O�"�	�4-U�,�'i�'�ݣ�"O>+�n��+�A��O� ���"O�� �dD6��I�ë�	r�D�)�"O��BK#�9	��5�H��"O�q��'��r�Œ'�$w�J��5"O���qkx�d��T�H!U���!�"O�(cRF�rޢ�ڷC�%%0u"O|Q������\1A#?<,�"O�l6�]�ui�C>#��A"O��1���k������դ]�"0���'���* ��tu�f-O�3�����'Q�
����>J��2�'��J��X�6�N(6`ٝª=�'�h���q-x$"d���"ș�'���Mǟw.*`���>��'9B�- D $k����(��'J�@*Ԍ�������kت��'3z��B��򪃫pH�]a�'���8���>��=�a�Pf���
�'�d��F(z���U.�K#���
�'�4,�����gz��T&� 9�����'T$�ۂ+�!�h܁�FR<
��O:հk�$����)ςq8�$��N2`�dʃ:�K�/N�?.�D@�%RБ� ~p�)�'4
؈s�Ԕsҕ,�>*6:A@���1�LI1�������i8#�uN����$ t��30�5�'ID��ӥ7�ԣcǤ.c�%���Z�es�Yr#!}~EI5r��ć��%�����*GŔ8���5j��'?�-`jk�,�'D�O�� �\<$y{
K1g��Hb�I������ ��سDE	��H�� ��\��x�r�P����)v�ʤWOH���Oͧ)A�0L�bF�Hr�ԋ��OF�ONB�KS��{�� S�_�`�	���84tI���M�U_�a�Nа��i*ʧ)��tO�3���� m�:_:a�B�A�A�&<k�ɏ)�d���S�)��>�x���[1y��$�uUh獓X��k�g�K�<�X��v�:��I_�x�e�4=�T�f�(~�F�����PW.D��h�`Ԍ��O��X��i�}�"��pO�0Xt�̅(�E�G���v�����0|6�f��!Ipbr�Ƙ��C�u?��-	"�K%�����S�}1�d��%ˢ5h ���ٝq�v�#6_�(R��@�����O⡱ �"~,R�A���#T���"OD���! �G�`t�R�F���k�"O�E) JX�_Ye���U7�0A"Oz&фL�UY�H�P	*��W"O^|r�샃-�E��g�b���d"O�� k�%u�^e�c��	�B�S�"O��ʲn�&JL�7�F�FT�"O��k%%�>d������r��X
Q"O��@�8��U���#	w�%��"Ob�8#$1p6��� ��#v8�� "OdA���S�KfTp����:�h"Od=Y�G���:f��|���"�"O��s���T֠�fnE�@`,؃"OX�,�
,����-E��"�"O�kA��j�(3C��9k���
�"O(������tq5��.R���"O �����R�Jyc&g�=�$�s�"O�\Ჩ(_]Jh1aE���P0"O�ѫPcY�]2*y���U�B<�q"O��	���N�:�0cb�\��]C�"O�����zҘ�UÐ'n���d"O�	�	�2j/�(P@c�-���*"OMʒ�8[`�*Qc�Ms�QT"O� @���e�H�0�`�v�T�"O�Hې��8�rT�c���\q��:�"O�Pc�V�C�|���å]��"�"O*�B��*N����=MK��R"O� ԩHG�����	P��l���"O`4��G�>IL�) .C
��g"O�8���UQ&��#	X�8���;�"O�,#�GS1N�9	CG�o~Ԍ��"O�<x#�C�}����%�(s�޼ۄ"Ol�aH]�Ex�5)x>5{�"O���G������CS�~��A�"O4�A7�ř-U��Y���I���a"Od�`�f%K�ĩ�l�K�Z�r�"O$��@ĝl�����)��Ĺ�"O L����nX$�FŔ5H����G"O�L���|��<~�UX�aO�8��[}��*��^�<��r��W����|�����.=������ �s�>����B��U.F>�Ԓ��["�*�ȓ������.��@�h�A.�ȓ� ���g�e!��+�vj���Z�*�j�,L'!b	0��I�Z�@�ȓ��%	k��f��K7훻@�A��R$��p�#'��{���W���5�l����ƒ,��K�]�9S���ȓ`hJ� �+&�p`suR�[
����~k`��E�V���	�CǶa*�ȓC 0JB!_������Z�I¶|�ȓx;�<�3h�  Y	vD7G3���u�|D��F\��z���6^F��ȓ$@��;'N�R�\)q��4e����j�+��-/��9�Ð�v&P݄�n��T�QL�	���ĭ�:4pp�ȓ\�%�p�S&�@�:��TVMFنȓ7E��z7�qF�������A 
�+�����ME�K�^���1ƙ�c	T�T�0�EE�$Jp������0
+1�`����'h��D� �[dhJ�Ff�q�'	�;>�0��{Fh��,T�a'�# [�c�$��7S��ö�O�.�l �� 5g"Q��*SP[�&x괌��Fu� ��m���cHQ5<�^i�D"�y���ȓU�0��Ji�ęP��'��D�ȓ~�W�I�s/PD��L]�\ņȓkQZl#��V2}��4±I߇cu�	�ȓ�Hȁ��9��L�W )U#|�ȓ#)\�K@ܷ:�z,�"���#p|���J��
��2o��	��.b.H4�ȓW��Q�&�F0D�x� �+Pm�1���FѫO��P1��<;�D��W|��h)��P��i�B� �ȓ)�����Gc��u Ȱ�J�ȓ[�F�I2��@	�*v���ȓY&,��޷�
m����${SM�ȓ_E0�H�@��]�����ɦW��p��K��4R��S�P�Z�k�"J�t�ȓ*�2,X��(d��3Co��*C�-I�l��ÆM۬�)�hN+��B�	�_�H-�qiL�l6��!��N�=�B�03���!/R�a�f��`��.bC�I �l��F=/ij�$C]|�>C�	�M�x�g@F�LC�_2��C䉦��kf�M �:��d&I�C�C��$}�,�YVj�Xx�ք5}�C�I�����0�� ^�څ��惦
ȈC䉷+�ڍ��d�V_�堶'T	SZC�ɳW��M珕�sc�����Q�^�.C�)� �`��F�O8�y�vKB;W�^ (2"O�ِ%�O�%�r�ꊬ@⼹��"O&�CB�$`z�"����ji�"O���rL��,���y��D��͋�"O���1��imڧ��%�HI�f"O�Ȋ� R?xBnT(pb����z�"O���9<B0��JF#b��!0"O"���#��0� ��C�<\��*�"OxL�4L��]�LE#���4+E`Q�"Ov���ҷ	���I;"C�R�"O��c��T�Vq�ƧLH���2"O<�v�	�����2k�$;P"O॒��1l�$�)A�<���"O�(��E�	w­;"bés�"O��B �I@�`���٘��"O*��f�)���DNJʀ`��"O���DV?�@��ѭA��c2"O,�k��7~0:���	i���Z�"Ox b��H�yp�x��� 5�fl�C"O�`#�
-rxq��d׌�"O��vS�y �����O�HHV"O~�{$D�h��A�C���"$1s"O�Yh����ap�B+{��t8�"O�}��+�J��ē�;W���"Oy�#ы��l���%E ��R"OQF��Y���-Q�!�U�S"O6��5ۏD��lx��2�0��"O����A�XL��!ơǨ[�0=�U"O�ɐ���0���9��K�Z�bC"O�ղ��T�a|,��!E��<0"O֕1� 1sO�h!�`]�i����"O>-����m��Cp��,��ب�"O:ʥ�F�k��Dk��%n�~���"O|ٲ�A�9:7���%�]�"OV�2g�L:U�&���M�5�Z|
"O>�0����8�Tă�ֈM�����"OĈ1!�/�:1����S���9�"O:]8����J���h�	�";��( P"O��:B�Հf���6�_�Siv`�t"O�����
)2:���E�1pd4E�"O(�#@�F!aC|�QQe5oa�yjB"O6�A��ܪy�~��dCJ�t]�y��"O��K�q
��.=I�*V"O���lDL�t��W��VG���g"O6	�`!�u�.��7φ{%�P�#"O�!1�+W#]�N�$ϐy�,�C"O\���+���8��H�F~�)�w"O�p�v��i��LRb�̖Au��"a"O���H�b�d�!�4ia Ȓ�"OجڠIC�^lv� �9�f��@�!��%�����C�yH�B�E�:�!��G	`�N�h�I]*3�x8E�[!�D�8fȺ�ѧD�>�����n!�Ě	c^j-��'K)v�&����]�oB!�d���}�7��E��a�!�-f)!��ǜ�����aǾz!p�BȀR!��
�w�����������xE�?e�!��-~��bE�֬&�VTY�W�&�!�({\Y���E��	�fD�	J!�ͩPW6y��-�<h!�dB�ě1"!�d�o�d	� �<>Z��tN�!��!m*��b�_�tF�2!��$'�N19���2���Q�E!��U�N�!�g��bݚ�itL���!�� �\��EG$�9�M����Mt"O�D���������.�h���"OLɚ��Z>�y �
�G�2��"O�L�#
�FO�$)�*V� P1"O 5���+m7@m�'�5e�*Y�D"O��k��"��蔌ۜZ�:� "O y�"��Y#Sm�1Iw}r����<!T�;��V(rp���ᇝ�<ޜB�I�r�jh�WɤMV�i�dAl	�B��q��Q���\�qV�����=bB��U�h�B懐�q3.����ݢ�JB�	,��Á��>�^9�7&I7� C�I ��!�[n`E �G�qS�B�$2�t��8&�6�	שƷ�B�	�v��8';B���I�`.|&nC䉾E1j�KC`�4�e�'�<�NC�ɇ_f�{o��Y��� rANC�I*z4�SE*�!:9����$U
PC�IIx���a@xq�ͫ���
&x,C�ɀ.ϖi��P�EQ$A ����(C��2g��a;�)OzZZ����V"Q)�B�	0�*p�d��m�z��h���$B�I 2Tv93�\�b^%c��R�BR$B�	�el���HZ�~���!�iM;�y�$Z1�>�NѶ4��D��y�ǟ�^��X�e�dcD��ဒ�y��پ������4���8�
P�yr� �L�j��p+V*bf�!t�Ȏ�yҌ�}I�`ʜ/��Q�Td���y��Ѽ`l�!��O����#���y)Y�U՞���"MB�lIT�Q��yri?C�*��']-E��:���.�yR@�gDM �G� Tf�p��߫�yr��,�����C�����yr�/�I��H�AN&�9�k��y��
DP\t��k�*O���i����yR��.GDrE�K5N�*��KY��y��G�&��\��"�F�����oF7�yDيlb�I��S5�D8�f��y2��"}r5`��n
Hv��yB�L	(��G� ך]�E�K��y�a�22 `  ��     k  �  �  n*  6  �A  !M  �X  Kd  �o  �z  ��  �  ��  �  ��  W�  ��  J�  ��  ��  2�  v�  ��  �  ��  ! � > �  r! �' . G4 ; B �H �O �Z =b 'i �q :z d� �� � ͐  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�O4����C|���D�4B�nX�lWCh<!�ER��x��ĕ20����,i�'Jayr���<�r�h�7Q�r`�rOF�yR+J?@˸�s����MQȬ���-�O�Y�㝍`x��$l��}AP�$"OPl�`h]�b�t"�!��r�!:��d�U����RA�]�>`S3��5"�B���9�O����J�0�IL�Mg��СϏ�=GxC䉵{��pP�k�2F'��i㇎A,B��ug�`��Hn!AIW�7vJ�prH3D��h��fGF�c���_Z��Z�)�>ٴ�O�>�9�H�h
��WH�Yu�q3D��QB��M�~͸n�&F��@�
#}2�i�V��� �YC nJ�l�X�|q���v"O�h��ɰ>�茹�.�^^���b"O",�P!�ys��I4��RT2ix�"O�p� ��
��eR��9-$�Q�"O� RUe�
��"��	�E8��C"O�c�O�q+���AB�.62(r�"O>���"�E.�Y�3/!(}��"OP�XѬP-"[|:�A����Sc"O:p#d@�*!V�11��r�hv"O�-����(R��6.6��rZ�Gx��S�R��B�$g����脡1�,C�	Up8���J��0��)�W²����H������ VC\ѸX���J��'����P�]�:0�A`�63�	���n��I����?�ƻD�B�8!��4v����K}X�GyB�
�Ax��S�J�mV�8�mT��yr�"i�L��b'�iq�|�Rjз�yB��""ǜ�����0J�ɲ�!�y�盫1L��!�3"� 8��Ƅ*�y�ͯGL��f'�	��-�
�	�y�*�h�H���g\�T�yQS��(�y�bkΰڥdP~�e��k�"�yR�#Nq����E��9!�Aܓ�y��
;��@�` �HtV�+���ybǘ"M��Ub&閬t�ބ�w�T �yRb��l<j\��h2W]fR��)�y�,[�k�N}`�K�G��Kl �y��W�JN����7?3�4cw���y�b�3>tX�`��09��w�Ё�y�g^-4���f-.�� ���N��yB�E&&|5C���Rd��!G@�?�y2iԙ{.NP�rGQwf�5���H��yBɀ�v60���^?!�R�A5ω�y��3}�BYِ	Ϝj���Z��y� �"@p��� M>[�`��J\��y�/ �#�\k%-IW�2���=�y�l�U�Z��ЋX�A� �2��Û�y��6$�Q��H�+ь��7�R�y�	{�\03`E�9��]�eW9�yC����R�^�-�dJ����y�g�Z;�4˧��-(��8�׊G/�y�PCE��!oé	�A��e	�y�S� $��w�C�ⵢ�Gۻ�y�(�sИ�x�T,]���W��yR)��k��3'�&u�C%LE-�y�J�"���%I�#�L�$�V��yBaT� ����N$Ԕ��Z7�y�ģ&Aj0S2i�q�������y�B�!aZ(xSB�g��e���Ӆ�y�aJp�Q;t�e.X�*k���y�n\	L3^�����W��h ���B�#O�x�)�W?l��P�J�'F�C�I�79<��X�L!�G�,ܲC��'^ކ�J"؏h�ț`� >#m�C�-h�ܬ
���-al�c���-3��B�I�v�D��C��Z14�x\�"OH$�E�ި_�ND)ҭK�u��A%"O��Z�挏[K�ȨǏ	�R�:eӔ"Op�� `��<�l��퉹~�z]1�"O�P2q�	Z�͡������"O2Xh�d $N�e�@�u�,��2"Ov)	kIw2�DP�yu"O:հ�C�[$JT2���\��9�"O|��������1NS�"�.���"O� x4i�T*E+.��p��44����@"Oq4o�)�ҥ:&L�V���2�"O���4ĀmhP��J.U�:�3"O8��͜U|$(�dʓ�@�^�q'"O��"�I;a�9��NW��V��F�'�R�'���'�b�'���'���'���%�	�:�3��EN����'E��'f��'��'���'Dr�'K2���[W��H4G�`lp{��'���'�B�'��'�R�'j2�'�P��(���&�a�G�0RR � �'��'`��'���'���'��'.�b!�<9C$�T��+l�rE�'���'��'���'�2�'f��'���e�ԣ;�Z�KF�[c�P�T�'y��'zb�'�r�'�r�'i��'wR�όYu��#d�� e�����'o��'z�'���'Cr�'o��'��ǌ�+
��:e�wK�Iu�'ar�'�'�b�'"�'�r�'�dTZ�BU�'𴹡%I��ti��S��'���'i��'Y�'B�'cB�'۾�Iˎ�y!LQ�&$�/PA�lҲ�'���'YB�'L��'7B�'K�'����  ��"F�����K�@mZ��F�'?��'���'c��'p��'g��'1hH�eE�N�A{��Cn�Ѩ4�'���'&��'���'r��'���'��=�*VQ>�1D$�2|��̡r�'qr�'|��'��'!�gӖ���O�y
g�N�DgҠ�dlC�O�@#A��gy��'��)�3?1��i7� ��]43G�P��M�,Lq.�;s�$��dƦ��?��<9��{���9�0IIB��2���3��?q�\�M��O,�ӡ��N?�p��˙*`�WG�w|��0�>�	ğ�'f�>�KD�7.�>�Y j��Ш��ݶ�McA�G���O��7=��9CEW�	�b�!��K/hO������O���t��֧�O�<0ᒶi󤁾9�t�a"���\xC$�6���v�l��7Dp�=�'�?هm�%bB�$c�m��M2����<).O4�O��m�KP�c�HQ�5-v4�m�'1��p;Df�T��8��	�4���<��OV}۵�Si�>�C��O撈*���L���aF�E�+�aGR��꟠�u�Ɯ5�J ��H�i����aFzy�\���)��<�s�W�A��e�E�S8����#��<ѥ�i��O�Un�n��|����&�,y�׉�o^���
��<1���?��Yh�8�ش���f>����z�0��q捽x*&I+�H�x��� 3��|r+OF��d��'L/�$Us�퀠9CH���1Od��
�H �8C!��ʦc>%���*�C��׊�Bh+�O9��d�O���y��'>i�	���s&���r
LK����Lu2��5#�X�*�@�>�@(��ae���Ҍӧ�'�1��J����fz꽢W	�4	2T��'�'C�7��D%���>{��m���\�݈U�7"[$�$I⦝�?��<!��?�4e
�#�S	O���ZQM)7���G�\7�M��O����ʌ���l��{�J��L��D�$�J"QnV�Z҂c��	DyB[�"~R��q'��a6]�+�Xp��UL�7)��T=��$LȦ�%�X:Gۤ_=!+rB�#���2Q���<�O��d�O�)O'o��7�6?�����@"#���U>����ù��$K ��O�P��4�.��?���,:��*.̋p��)[D��<�K>���iC�y�X>�Y���;�بiKE	y���t�1?9�Q���Iʟ�ϓ��O��E�h�%�(I硔��nEb��'fV�qÏ҄��4�¨��	>�O���mL$V_jĢ��.a3Ԁ#�O���O�d�O1�|˓vB��
@�
����$���Dt��D�5o�a�0�'1uӎ�0ѭO)o�<Xѓ��۵n�l,�`�H�I�MXش�?s���M��O�I�pۘ�).�Dk�6Z�Rq�
�4;��y"Z���I˟���0�I�� �O�XA �GPܼ�"��,BglucfIb�2-����O����OL����D��#4�"�ЁgJ�*�έ01�N:s}@��4k2���|��$�śF=O(�`v��@�M����Oj��3O쭙"^��?I��!��<ͧ�?��b7k��b���,������?	��?q���$�㦹�Qi�ҟ,�	��p��X"%[�Y��d����v�eL�	om�	�k�>�{�Խv(�l[��Q�#�L�~�T��>\G�I�|jbM�O�I���6��[K~�m����,����bK�Oo��?���?���	�O��u-�o��H��K�|<��fc�O�)m�&uD�i�	矘�ߴ���y�FK�%k�MJ�)Q�r^|����ç�y��y�vn�ן�B�o�Ц��'U|M����?�YÇJ!L\�uƉ5�p�u���Z0�'��i>���ԟ���̟��I?bA`<�a&6q˴  ���k3Z)�'�7����O��;�)�O�u�r��9Pr��a��կv��j���C}B�mӚ�n�v�)��#��|��O�������x-�!<1Z����U.�O�(�K>�-OP[��R.`�@��E�J!ڲ-�O����O��D�O�<qV��e����?�sFBX$qj��6����)�<)��i��Oa�'�"7m���޴`2�	'�uli�����:4��d��M۟'�RD� _�T�����?%�=� ft�g��
���eۀB�r}sC;O��$�O����O�$�O��?%�����5h^S.��Ɩ�h���$�ܴ���J.O�nZQ�	5,���CVH�xf�Z&��
6Rbq�J<!��i�6��4��Q)���ҟLÂ)�'u5��0�-�'��Q��w�2!r��'�\$� �'��'k��'c�4 @�_
�Q�B�6fo�aD�'�S�\q�4"@�(OL��쟪�)A�D���*C��vh��D�It�	�����Ob6m�q�韈��6:0��݆8����E#��%��aӱ�W+(��m@S��<A��U���$N���qm�	h��Z21ɞ����Y'����?����?)�S�'��d�Ԧ}��$M6g�-(b�����a[��۔ch��C ���d�D}�j�~�fa�Ξ8  cN!_3бC�KΦ�K�4uJ`� ڴ���\Ϣ(`��S3P˓L�����	S:|u�1�B z���͓���O����OD���O��d�|�#G�k�$$�S-�1�X����*$L�椗'$w��'�����'�7=����X��*�J�	�H���^ȦiشA����O����i���P9#D��B2n��xR�ެ]l�@�{4���-�l�Oʓ�?9��'�S;�X�#�j�����ϟ���Ɵ��	Syi�����O��D�O6��*��<0g^De��@s.�O0�O���'8�6͇Ѧ�3K<ѥΞ@��&KQ�H
@x���<y�K�$q����m�(�/O"��܆�?A�l�O��� �Z��i�P"^}Xj!��O���O���O�}B�'��p��ϛ|'8��T���[�d���� ?��	�����I�MK��wϺXr�E=1��0��ЫJ� Q��'�"7�O٦�ܴ'*�X��4��֠[�p���G�d]�֢MYrZ=�a
%v�N�C�c>��<���?����?����?i���W�p����˾r�D��G� �����Ѧ�;�JDy2�'�>��'�7B*03��5m�"A@u}�OxӺLo�#��Ş��}P0o0]���с�B0-���� B���C�򤋿t�����14v�O�M��l1��-�ѡU"`���2��?9��?���|�.O$�l4q�\e�ɟ�`�" %��b"�Q����~��	�M�ҋ�>� �it6��Φ%���I4E�6����n�E���)�*�o�[~bm� fW8���M<�OA��[<O~��i o�:Lq^���n���y��'���'��'b��i�N�T������&�t���݈i����O�$�ئ�)�%�ry�`Ӏ�Of��^u�d��1@�W膁7,��+�'��7m�����ld~BE3+:R �]�x�mSk�L(ƢL� ���|BR����Ꟁ��Ο�ir��������
3.DHc�֟T�	fy��jӄ)�q��O:��O.�'dLi��)7��rg��)�x��'�J����l�
�&��'@���5�[	NȄDi�H���I$�<JNH�1�lK���4�)A�!���O4l@F� 3�`��N�~;��E��O|���O��d�O1���%����8� �$5F7&��B�թV�m��'Lb)p��올O,�oZ�U��yC��#d�L��>:�dA�4k˛�A\&�F��D[��V$f� �nyb�CKu`H	��(H��ʄF�5�y�W�$�	ҟ��Iן\�Iڟ@�O��txr��:��u��!FA�ư�'�h�N�T��O6�D�Of���dAܦ�ݍ�p�-EN�b���� ���H���M��|J~J�L�M�'�.�:����eK��-v꜓�'�H�q,^��<�r�|�\�����d!RO�yVz�Җ�U�Y��<*lQ؟T���0�IlyҢy��u+���Oj���O&�:CN�]x���h?i�t{�"�I����ަU0ش�'{��H�G)F6��jV�͇c����Ob�	�L�,7�N�)�f'���-�?��F�ON\�B(gFDeٷi�$.�yw��O��$�O��d�O<�}�;w ��P�N�e����DȈ%m��C�뛶m2��I��M��w�҉P�JOXP^X��IH#4���'��6˦]
ڴ7��J�4��R�Ji�%������I ×�Y1j��@�� S�X�A"5���<A��?a��?���?iLܶMV��S�Z!���wb��D���	S6(���P�I͟�%?�	�4�����*�H�@䇈4��eګO�Dm��MS��x��D�űM߸���O�/v��SAB6'����&����V�8W�'#��'��'�h���� $�@ʖ B���5�'���'����dY�BܴZ�����}�*���7%�E��I��T��?�ſi��|���>�b�i��6-���!���
k�ժ��5Ua�1sHڇ,�|�l��<���f>M�����ȫ/OL�I�a���(\f8�!##ੂv;O����O@���O���O�?aJv.T�)�c�5_����$����Iߟ�ܴke�AΧ�?�v�i��'����s��KY( ��9r�5(�	.��KߦI���|f7�M��O"�y��߂z����7c��|��\����`��=��p3��O�˓�?��?����a��ʘ�9����UY6VԂ�K���?I*O(�oZ,ks���	ҟ���i��C�zà�A���l.�Öc���D�p}�i�4Dmڲ��S��LA���3��!w�����.by�����!��y� \�� �rH�`�4Y�}�3�܄F���`��kڔ(��ɟ��	ٟt�)�SVy"qz	�=�h+���(]��-q�K�<D���׫�<9��i��O�-�'��6F�+�C�j[��$ѷ��%��oڃ�M�R�E=�M{�O����X�����<� 2Y1�*(�B,���
�\�92O�ʓ�?y��?q��?�����IF �P���G�+:�x�#�d`k�l�Z7�d�Iϟ��IN�s�X�������H�L�!�2b� )Y��T���Ar�rM$�b>ef�ۦ��w��Q����%Ϩ�
�$q�r0̓+j<���O�A"M>�*OD���O$��@+I��|i�*HG�0����O����O��d�<i��i>M[��'&R�'|�3t	�TSF�*rč0=�p�����j}rabӦ�l���/�R@h�ʕ14�2,`���,͓d�D�霂HV���n�/�?ɮ�0��KOݺ���'�t�7%D�=i��T4<ƴ���'��'���'*�>u��Z$��B�T�>�h0��[�Xy�I��M�Cb�G~��tӰ��*�i�����Ź�e��>���6�M�ǲ�Ųi�B��i6�ɜ:������O?��Z&�M��a�!� %y��`�D'�I`yR�'��'��'��.��~r��S�L"6c�e����I��M� ���<����?�O~��x�̓ ^	�ŀS#�G�x�^�pj�4(1�V(�O�#}��"�+^�X��Vz����rhOw�V�H�%�7���!C0X);�Ÿ'��I�WN�#�A:Kp�]�Í��}p$��I�����P�i>=�'��6�M3t��D�5W�A�-
�Q�0@��!šd�$[Ԧi�?�3T���ܴd���n��q�"/�US��ؤVҵ�w �:U/N6<?y׮�l����������e��/�D00���M�����,�<���?����?���?Y���K�'g�u�\�_d�A�f��'U�q�����<���$����$�H�%c�����c"��M����[4����v�~��	��s;T7�)?���&1�]zCH����f�{�z # c���%��'f��'���'˰u�0��7ÈT{���n>�����'�bX�P�4Br�M����?	���Y4#��0(���
�B�K�B��ɜ���˦1����S�@�$��xs��?e��*�e��^$PIR�ʑGHZ�R��
)H�hY�ɞc��W	�$U�(يhEHQ���I�����h�)�hy2$��8Re��:P1���S&XYY2m��*9��?�e�i��O.Е'���)�>6�ƨ��� ?G4��;	״]��6��ئ�3S�����'����e� ~�.O�b5�30�
A��;���9O�˓�?���?q���?����)ܝU��A���8@z�s�B��%m�
���	�d��z����r����Uk��,zJ܊�G�h�� o^�·i�����<%?�h��	ۦ1Γ%�`dp�h� *�h�P�C4��S�� �� �O< J>�+O����O�آ4*�J7�g����B���?���?�����ę�1@��n����؟�0�*<�NybV,��Lo�y�#�x�����
�M�i6�d�>9���	,X���-�:s�L9��Um~"�)uJ�H(�!� f�O�x��k?ᓉ��6zm�#�OF���SE�?y��?����?����O�h#Da�2�ZH�A����ĩ!�O��lZok��vț6�4���C�	3��x2�jʿ9���v?O.�l�	�M�ҿi��p7�i��I�~�
5�'�OA�x"wo'K�t;t&ҝ!��hs��:�	]y��'���'A��'��Į���#��/�:���i�剢�M�I��<����?�M~�.��]Q0�טF]��3��SH���^����43ܛ�i�O�#}j��V#P�
@ܗ';x�ȗ�>{�x�7b��^�j���Ը'��E+W7
�dY�@�*a�v��d�'r��'<����TS�ܴ'�~T���i�y��չu�ltY��#D�ɒ��l�����_}�ld�����¦QCQ$�*k�vI��]:�Z�X�`T�Ed��m�S~�c��Q�Z(��]��O�� T�X(d����^nR�HvlƘ�y��'J�'��'xB��^;s�x�1��L�RKʲ!����O���N˦y�m`>9�	�M�K>A #Q�k�~�g���*PR���2�'=�7M���ά.�V7-?a #@�!x�YvC�)r�I@������G�O*�K>�*O��D�Op�D�O�-	�� �(|��0肢N�2���n�ON�$�<	�iS��[1�'���'�哉��\�q
�
����F<�Z�j�	'�M3��'4���I�;L�ahr�
@VU���;%̹�P�ܼ/k�y�o�<ͧ|����>��
Ҫ(b�����kT���Ȼ���?���?i�S�'����at���m-�x%$\(Î�ط������Iǟڴ��'*��G$�F�P�Bv��S1LYSprA��L�k�̑1�`Ӵ�9X���VF���(O:�
A ��=KpH��I?���R9O�ʓ�?���?A���?�����۝u�ԌH2��(-�02��5e��%m�2E�����Ɵ��	u�')ƛ�wҪ��-*>�cj�d��yp&�jӜ���u�)��O���n��<iv'�C�6D�U�[�/�+A��<�jRR���Dl-�OB˓�?A���*i��˛PX�4�eN�X�t����?���?!,O��nڧyޘX�I��P��(�~p��4~i�E��DV*<Fm�?!�V���4�2�x�M���5�H
`Ö�{��Y�L&~�͓�?Q4l���Xbf� ����p���_�����zNn,(�ᒴ%?��Fi����O����O��3ڧ�?�P,�??B�S�ޕvP�����S��?�i� ����'���zӌ���T�t)��$	�_5����̋�>����MC�i8�7mT�>I�6�)?�OؗPy��)�n�? ��`� 5�$���-TU�%���'��<����?���?����?�f�9��ԒŪB7h
L䠕b���D���ۡ�`��ޟ��:$a}���c�
ާ"�
���� : �	;�M+��i�VO1�����L fB�X2�*�|"�L��R�o�`6�VMy�e��@�Pm�������,����D����Y���p�<��Or���O6�4�ʓO��^T���<p�h�g�� \[s�S�Tib�k����i�O�	l�)�?y�4'��)�%�ź0��[D
�'��|R F��M��O��:�銿��.%�i�� hR��48�Vh�'�`cq37OJ���O����O6�D�O`�?�ؠԹ����P*<o����	�̟���ٟߴ\�$̧�?�i��' `�"F�а'�~Q3���f���CB6�d���y���?�U���Q�'$`� �I�!i��PX�g��-���G��k�n �Ɇ0�'��I̟l��ڟ4��3]���F�˻AU�X�c���Yv�Q��۟ԗ'7�	�����O:�d�|�C�L5=�RjJ�h��(��Jk~r@�>)��i���'�?����8�$�ipg܄<�Ta���oȚAQŉ�x.l������ܹ֟ �|BN�,l�U�ԃ�	��Ȃ0���j���'q"�'���^�p�ܴf�pQºX,�xT ]�U��ks*[�?������PA}Ҭt�.M�K�1p,�@܈ ��pv�F���l)M:��n~�"�!������I'?͠�k��]�^
�*&�� j���}y�'�b�'�b�'��Y>�i�T�8ȹ�F�G���f�[��M�bQ�?���?�K~
��jɛ�w��5Q�aD.O�r�7H�z7���������n�)����mZ�<1׬0QD��* FSM��Ы�^�<1E��-e*�D=�����OV�$�
\�&e�ԉ(;��PΖ'2Ͷ���O���O�s'�f撻{B�'W�*C��q �	x��ǢQYA�O}�'}6ML�ŻN<��G[�SE(d�i�-n���t�[~BҢvѾx�c�M��O��\��M�b�.O�ΑZŝ6g%���d��D���'B�'r����0���6Y�����۸|�z���ܟp�ڴ\.�|��?���i�O󎝺\k��Nŉ{�4����?G�����)ٴ+N��,�R�����Dq�Y�}��dkM07π1���J�x���Ŗ,ň1&���'�r�'4��'b�'<�Y�)��w_D��FŘ; �(�P����4r��4���?���䧆?	�.�w,j�RU��'>`�u�A�	?f�����M�"�i1O1�*��w�3���R7F�3F��(�<N 8+�Ġ<�G����D�������:q���tC];LZ$��2�K���O����OJ�4���Oݛ�R$%�"��M9~�Ѳ�D�s�4�b�'q��e������O�alچ�?��4/��҆�ŋ[��C�#D`h��#�8�M��O����Ȁ�
��?����,C1�ߋj9��ufI3x)"��6<O���O����OF�d�OD�?�QR���E��˒H�D���Ev���	Ɵ�yݴq��'��7m.���,D�Љp*�'U9F�����`��E쟌�''����4���|p�֜���U�Ѻd+pd[c�'pB�C�*u&<�jv�'EqOZ˓�?����?��M�i
!��/7o�Ъ 	-]|�C��?9*O\�m<c�6�Iџp��D����'n���$�0UT��Ř.��D�f}��xӺ�lZ�?ь�T��5
B��c0K^<:<ѸP͙/,ڭ�@��&��`�S��SU���ĉ�?l�YS��'vW
�;3�Q4-��D�O����O@��I�<�C�iň�T��6���� 6��ŃU扛��������?�D\��[�4@�ƔJ�� Π����2����ib&6M�*��77?Y3A\�#˸�������F����@S�y���S�Q)s��ĭ<���?���?����?-���G#��G��0��)�62�&m�Ϧ5��mt� �	䟈'?�	����w[t5��ͅ.C�|h$���ЍӴ��OT6�ӟ8���'Y���4�y�L�\���_=�)9���y� ��y*��IZ���$�OJ��Q�4�e�sa��Hb�:GD�hl��d�O^�D�O�ʓu'��iG�?!���?i�OB�*�&��&��7Lk�MK��K���'D���?�ٴMj�'O�}I�oK�k=����D>���Op4��B;J��6-�A�v����O����	�d�K� U<�uN��f���'5B�'���s�����W��HC��\�Wp�#�@�����49!�����?��i��O�n��L����g��B�����V�_��ă٦����M����M��O���7��tJL�9�JL�с�!_X�0��5U�V�O��?q��?)��?	��c�|D�� ��$c��w���.Or�nڰF ���?���h�t��Ne)`�v��!iS��ot���f���_�Oc��K�+�~�ġYr�3Z#���E�g�2�@�]��X��9���<i�h8s������b�P�&��?y��?����?�'��H���G'u��!&���2F��?�F�lv�|ٴ��'2`�?z���d�J�l�<C����7��>.x�
�I��'l�hñ������'DJRk��?Ah����p��z �S�n�L���Oٞ~��⇤g����ꟸ�I���	�����I�a�~<�VKX�TI[/��<	��?��is���O��nB�I�X��ʢ�׏z˔�C�k�T�{����!���|��j�4�M��O�5(� TAK��
.v�[u�ǥ
��P�����?��{�^�@�Iܟ�	��
�'mn��	D��h����C����YyBqӢ�Z�=O����O��'p��)x��K�+'�yJ��H�N���'�j�>�� q�H��	M��?���������1e��(`�R�HP��K$28P	�<i�����D,�ɋ0��ɘ!����TB���MmZ���ٟH������)��byr�k�6�H�l�v6����lr�*=�bW$˾��O*Xl�g�\����
�dG�N��d��JU2�Y{!���?�� `�Ul�K~R�Ӏ;�$��Ӹm��	�'���&�V^@�#+�'�2�	@y��'��'D"�'�W>�X�F¾K��s��D6��6$��M�e��!�?����?�I~���`қ�w��<0�"=L��d��"W2�HU���Of6M_^�)���W�7Mt�`�c-E>�p�2`ıM~*����l�@���,�=���<I��?iU�8F�a���T�q�\r3��?����?����D����A~y2�'�䉒f�ˋE�N c���:��M��Āuy��'$�x�鞇b6��WK	 M��
�����$�D�Aӓ�N����� U���6�D*8%��攬��s1JWwi(��Or�d�OH��)�'�?I��&/R�Sq!@�1���։X�?öi�za�q�'�Bhe�����p��C΃u9�i��*ȃ�D���Ms��'����W�X$�Ɯ�x�G"����G;S�8��BDF?s*T9%�<Ɛ&�@�'�2�'���'���'��ىufG,r��A��	���;�^�Ӧ�3W/D矠�	۟'?��	~D�J�`Ҫ��a85'�K�4r�O��l��?�L<�|ʣ��%u?��PP.�)��+7_E���+�C5��$�48,�{��*��O&�g8T͒se�\'�]�1�_�:a������?���?���|j+O(4mZ�e�r(�	�m�dI��%R��[Ct��ǟ�!ܴ��'�,�J���,�O6��&7�5�vi	6!6�����-U���g(���d�Dd"�)쟼]H~���]5	 ��Ndn4��j	1@�,�ϓ�?����?q��?Y���O����dشF��82��T�J9��'K��'2�6�
%Y��)�O4�m�M�I1�ܫUN�p��S�(�ʹiH<�"�i�6=�@$�&Im���4�y��/4Cag��(�TB�ɘ5h�t�IX�uy�'B�'�"��&B���aG0JlXS��2���?)(O��n��gO�$�	��d�	R��� �V�L ��B��;�������P}�'h�l���S�4�
?hK�0��SǣYIf�
t���Cr�lӐ����	S?aN>��CΧi@�A��K	�+Kԅ22v���O�q�����O1���f���K<rJy�ei)n.��fB��Zfڤ�c�'���p�H⟜�,O�6-fB����(@7VH�d�]]��m�?�M��j��M��O��0�7��dZ��9B�^/q�a�U'L+J�nm1^�y2T���Iş��Iß�����Ou���HOhT�h'Nܠh�t���Do�R!I�O����O�����Dʦ�]2F��y��7��Y�S��2�$s���M���|J~�`�(�Mk�'�4�:�MϰQԔ�����-Kz�Y��'��D�l	x?�I>i.Od�$�ON��$?��zeNb�,(9Am�Ov���O��<�i�V�;�'
"�'�͉��U<:v:r�T*��"���P}�u��yn�?	�O@��rჲE� L)f��i�2�㕟d����qg�pEUh�S�skB�O�I�Sg��R��,Y�� _�F܃*�O��$�O&��O��}
�^��y8�$�&
]<!k��JI�9��[v�#ڲ��$���?�;koȈ��B��8��f<�<��F�{�XLoZ'>���n�u~Rb�h��)��Y�yQ���M!*���(̍���ȍy�X�`�I������|�	ݟܣV�� ��a#��R�.43D�VzyNs�ԡ0f1O��$�O����$ͯpU���)ň]�=�c`��ш��'�@6��!���H��+�f�0,���
S9Gu��Cd�\�G�8	+`�<Y�εQ���$�	hy2JI<v����3z���2�� @�R�'��'+�O\�I��M;w�Z�<it�H�F�L�4����9�!�<�D�i��O|�'Z�7��Ʀ�ڴ@���V%;�*���]�"��8�'�5�M�O��Ӄ�!��T�.�Ip�!4j�&o��4��I%([W���y��'_"�'9B�'BB�)��[� I�ݡf/ޥ�UD�9��D�O��d���.��I��M�N>u��6(���F�I�y3 � T�"P�������S�w�l�z~���@��vN�?,p�ИQ(�ͪ�����t�=�-O��$�O��d�O�0xs�L�<��b����xDe�Op���<9��i�Jٳ�[�@��v��/W���	��mruBS����$�Xyr�'R�|*���+�gL0'*��h��]��=��"K�{0�ɓ�R����|���OZ��H>�4Jԋ>!�|"�=z{��B6cۇ�?!���?����?�|B/O@un�wɔ퉋f��kW����C,?)�i��Oе�'4�6�u�R���.��X�T�����#\�1m��Mk��Ը�M[�OV�2���������<�$��t���� %�'g�]��*��<Y/OZ�$�O���O�$�O��'Y�b��g����j9�1@]��2 Q\/᪴������m�'P���w亜{D$�
{�D�r/M��|�F&kӈ�o�4�?A�O1���Eu�@�)� �e�r�?s��pe;:r��2O"\$���?��{�Q���������&�N�)�g.�L����W����I��4��lyht��3Oh��Ol]�h�,�8�$K
"5~9@� 6������O7-�ڟt�'K�\R��A�v� �ʚ1o,Ts�O��V*J0
���2�I)��B1�?)�'����&�;4sP�B��T�%��	�T�'{��'���'��>���.�@䡷D�1!Ԅ1eMɓpw���I�M[��Z~bAaӂ��ݶ-h�ȣ��T(z`"U�f#�扑�M���i�6M�RlJ7� ?�d�O��^�i�<s������Y�"���'^|�.��<�)O��D�O^�D�O���O���`hĨ������#2��dk�<�7�i<���'���'��O�BmPf]̹�D��d.�| �V>y"�j���hm����	d�Oe���d%ԛE��SI\�*�0��A��R���<��i�/���������Ĺ�&Iq@��3uE���tS|v���O���O�4��0˛�@K' bb�$�����!Y,%xc�9
%""b��<�OrIn��M;�i�j�q�P�uH�9��£��x2�,Z9-g������#�\���tgA��>�5�&G��uC��Bv�%� ��0�y��':��'.��'�����u*���Γ��h�W-��As����O&�$��gNn>=���MKJ>�wi� H�L�᫛��6M��C�z��T�$�	����j��n�y~���9�2�p�J��1MJx �@�'M��`0��̟d�|"_��Iş������H��~R��I�b�1]�"q���ɟ�	_yBFe��(I��O��D�O��'f0�҅ν��l#ր,H� ��'�
�8��Ƃf�p-�	a����&�%8�؅0�#Z�c0�@
�,Nqp���O^5��4�lѱ�vՎ�Oz���hA�K3��@"!̌���#�O$�D�O���O1�4��ܴ<�N0iH'��$�C-�y��NH��?a�� �v��L}�}�V����!R�ƅ�w�9�2�9�aUϦ�#ܴX�ܴ���!|Ԗ���'���	�t���&,���7�V�A���	fy��'f�'���'��R>c��Q�`=�	LI�D��
[?�M#��K��?Q���?qN~J��
I��w�-�u(x�1C�	ރL�t�;��O���1����F��m'�63O�)`dmYH��2���o���0O�u����9�?�&H(�$�<���?Y��.#qhuD�-q֠<�W��;�?���?a���DIǦ����������@�1L4C�b�1�LT	[8\�rď�t�
��I,�M�@�i'jO$@0�L
JD��	sI�@�R-av�����R$��=Y2l�W�S,��l�ğD�l̢ 4q�������{6��'��'�r��ğ QA��'r;�5#��3Cjy�e�Zҟ��޴O��'�p6�4�iީSG�T��@]j�bO�b�vm狺��I¦�8�4���s�4���Ǳ��������hk���#! ^dY��T>0�
���<i���?����?���?�3l��N�0�d��	%h ��׾����ܦ�r&(?�����O�� �f���ܑ/
!ؤ
���>�0�iQd7M�۟E��IU�U��e�Q�L���V=~�:&��#��I�Z���e�'yqO���Q���S�i����	��R��?���?Y��|2*O$�m�{�|����:��Js�G[���`�u\f��ɇ�M�"+�>�1�i�7�ݦ��3:��?�8��!R�
�M��O|����!�b��7�I����B�q�4Y��/�:oVLc�H��<���?a���?!���?	���@B6m��ypɀ)�z .f��i���?���E��@_�����':(6m0���4\� =Z���t����ž��@��c}R�`Ӛ�oz>	��L�妁�'��k����c�)��LQ��F����'T"�&�ܕ'���'�R�'�&�q@�5D �d���@���r��'U�S���ݴ|@Ո��?9���)�(L�d<h'Ǆ/%�"�_6D��"��d�OJ7ß��~�F�Ld�����;�p�{v�Jodv<�D�^Z��)O��]�?��.�$B�mT�xC��5휑0`Mԛ
!����O����O ��i�<I�i�v���,$ob`J�� \���q��Q�
]��'�n7�3�I����q�ıB��}J̽@��N�2���B�릵��4���ߴ��dUyK�������j~r��#	Z@��Q�F�N%����d�O����OR�$�Op���|�2+@���j�	֗F�V����7��VmR��y��'����'v>7=�`���ݷ7�.@"�FݼR;��b���֦9��4�"_�b>Ic�AҦ�ΓL��LI�I�Q�H��U��a� HjQ1���O㞔�'	��' �iy�hJ�K�Ny3�\����"�'���'BX��k�4L+��?��Z9�iӑ���kw��`�N�7N�
d����>ѧ�i�6�D����'�&Ap3�МA�`��!X�Y"�� �Of(��V�^�^!�@e;�i^��?��'�tY5�Z�Jt���@\%P�\�t�'Ar�'���'&�>]�ɨA���j��]�O���X7aP- ��	��M�5!�~� r�&��)�|���1j�$u�O;$��ɯ�M3�i�F7�%O�T6m7?Y6J�UM,�	ړ��@Z��
.i�=�Ƭ֘N�"p�<�.O�$�O���O^��OQ#�č=L�� �ď{Z(yC�B�<���i�܍ښ'�r�'���y�J�;]i�@�eM��~] �E����o��jwӦ`�I~�O3|0�� ��6��!|<���A�'o�������|��˓�F R�o�O�㞤�'d�q�ŏ*,�Pd�cE�>*ʉ���';r�'����P��`޴$i��ϓQ��!���&SA|92��/{���ϓK*�&�DN}b�w�l�n��MF���l9��Ä���Z���1C]�9ݴ��D��H���>[��� ��y��X*�-�/`����T(T8�����?���?i���?����O3��2����yʶM����2$�z���'*b�'4�7�ڂ6�	�O�$o�L�	.r���F�Q�mlv��!?pD�B�y�	��M������U������"Wm� ��F�H�N���$
(kvP�6�'`��$��'6��'���'�f�8�N^Lj	@Q��#���"��'�U�0c�47@���?q���iX�P��m:�B̼k&���b#̈́M�ɳ��$QĦ������S�d�οa�¤0�$u�H�zA�=y�����&`�q�p_���&h`2Ƀo�xƠ���ퟪD��1Kr�Ϟwb��	��	쟸�)��yyb�yӎ�Ѳ�F�mzx�R�N	y�j1����I��M��§�>�u�i����Q��q/�|B�k .������Ul60��lmj~r�Bqi�L��.�I� ���bo9{d�����J�9����my2�'�"�'�2�'h�Z>�#���_zȡ�*
W�@Y1��2�M�@a\9�?����?�O~���}��w�F���ѹB��BB럜����t��0���)�S�5���lZ�<�6O��T�E;Ӯ�8[�X��஄�<�G%L�>��d�9����d�O�����~Ea���p�ы��F�CG����Of�D�O�ʓJo��DӒ�y�'�r(��}7p�W�V�4r(8��闔��On��'�6�P������K�ol>���/ѣ[�$�D F)E��	�GڴX�0 ��R�"t%?U���'��� �9�г��9�n����_C��$�O����On��&ڧ�?��]'']J,h��9!���Co*�?�3�iUDu)g�'j��a�����2Go<�q1�Q:j������I�X�-�MK!�'����˩]��������4K���ÒN���8�F�@|0!݃,�f	$�d�'�'���'r�'�v�;� �[�Ɣ"�� i��lP_����4g�~M#��?���'�?�'m��6�V�����
%�ebGh%+��I֟�nڻ��S�6�f1@���gB�J�$�
i=���N��-�-O\H{��ǽ�~�|�S�$E�O,��P�+�O��В�hXwy2�'c����R�l�4z f	k��Fh��@�B�+Z���(1�Bmc�&=���$�K}�Eq�D$nڣ�M��?Y�\#̗:YG01t��e��4Sٴ��d�3FAc�O*�O��
��8q$�ba�u�~p����y�'���'���'c�)擥��<��@щz<Zt��fB�C��I����I(�M�Uk��|B�E�V�|�Bռ|���ɕAC��
��'�m+VOpn���M�'K�4ܴ�������	��東!�r�{s��E��j�L� �~�|^���	�����쟄�b���R���'��r�A�N����	dy��n�@@�?O&���O��'6�.y�'j܀f�����O,R�0�'`�����n{�����y�]3��ؕ�Lqݔe���ӧ9�U�5��'����-];��4�<���'V�\#ՊU��x$��n�Hz��U�'���'�r���O�剛�M�#�'�� F��+Cc��y"A'V���Q��?�iM�O��'�t7MβB��X�r���eJ�a�t����1���VԦ��']@���?1�Q�(�SA7,�P���>��Qy�/d�d�'�b�'���'���'y��)5s�����I�|� �®@�k�|��4Sw�<����?�����'�?�S��y��1WF������6��/���S�i����?�󉘷H��7`�a�ύ#�fqH�B�8�hՉQH{�(�` v "�O�IAy��'��Q�iI V�,rmX<sU	�#jd2�'x��'����M��nE9�?����?�7��>_,�1�w�F�&)�����'���O/�ƍ�OHOۇ��5n�b��&j�7a)�����1E�,�|����R�.�Rƕ�� ����I��0)��v`{G� Ɵ���ɟ0�	⟘E��wܲ�h�R�X�˓kZ�B��4q�'�\7֩<xz���O�,mZm�Ӽ��L8%ݔ�HP(��Gǰ��#��B?����?)޴l�0� ݴ��dQ1hy���'4� S�B�	�	p2D�;js
p�N#��<����?9��?Y��?Y���T����NmK����M ��d����	w������H'?�	�M ֔���R!^kr,�_���I�ON�n��?�M<�|nV+*}�FJ8X��%�bҊ�[W�$�前/�%��'�D�&�,�'�,���".�Dadf�2����'���'/���d[�\�۴x�|���cZP�y6��RN��%i���!+��71�f�D�H}��r�F]nڱ�M#¡�t�4��O=l:�%+6�,>��6�'??i6/�,6v��J��'!k���y�d������X�[+�P��'���'�2�'��'C�&,ۢ�W�;���qmW�~�&PY@��Ov��Omoڻ27*�SPߴ���4��Ѥ�Ec���w��8��ub��x��hӴ�oz>��ʦe�'
�!���`�d����ЄWy��[V��o�~a�������Oj���O��Gq�ʍ�uf���Ve0K^~��$�Of�e�Ƃ��~�"�'�_>�s�F���#hǳzYH)`�7?�&W�(kߴWa�6�1�?� ^�ZWiL�*���K"(��h�E��F�z��f�^P�����b?�J>�b@է%B��ǂK�1�V9z"'ά�?a���?9��?�|r)O��l�&-/&�#ED4K� �A`�$o���B3AB�H�	0�M����>���i�h�b���0 �� k̺2�Y��v���nڏ~�tDlZd~�斐09������dC�q22-Bq'�<�v�#p�x2��<����?����?���?�.��M��g�"U�.��3큥*C@��O\���e��ğ �I�x'?%�I�M�;/�`i��#S��!�D�
]�����'9�FA8���D�A�(��1O��d�@��`�q��ԫ6����3O�֮�~�|�R�@��՟��M��=Bu���ԹC?l�9V�����Iݟ�ITy��h��	�PJ�<���`��|��Y=[����x���%�>��i�7M�P�	.@�`E3�J��\�{.oaM:?�qC۫[�� ���	��'_���9�"�?oH����#|]`�N��x��'���'�R�՟|�B��=��ԁ�H\�k�x����ş�+ڴ.bd�k��?���i��O󎕃��H0
�H�aREM��&o��Ħ���4E���#
�Ƒ�<ʄ�ڶ]I����vY�d(�],e��4�6�ɪ#Y��O���?a��?����?���iP"�7�<rv�	7�6nM�t2.O0mZi��a�'�r��T�'ll�� �S�HXCic�욑��<1���Mc��|J~�t�@�!"�)�����+N`)�ܖ �1#�4Y�	�2�xpP�O �O0ʓE::�y�l,x��$�tfU(-�����?9��?I��|",O ��p�V��O���HDNW�|�#G�0(w�a���O}m�\��M����M��i~d6M�1x�9�g�J�ص;������`W�i�
�h��eL�?m%?���&b@�3j��Ex� �p,Nx��Iğh��ן��	���	i�'<^�z�.1WJ���Ь%����+ON��G��p�t>5�� �M�I>�7�5i���Ǌ�Y�UE��2�'�6m\Ŧ瓳<�Im�v~�oF3 ~�bV�ȍe�e
�A��D�0@9���h?AJ>�(O��$�O���OƥȄ�Y�à|Zc�Z|X\*p��O��Ĩ<���i�0��1�'D��')��;_�������cȤ:��Kwd����I��M{��i�lO�ӸF�<�FWN�b�;��}0�@���`���oZ��4��c�'��'wj����Nc$2a��A~j�s��'j��'x����Oh�ɓ�M�wA�z����!(�"_s����������?��i2�Of��'}"6+g2����瑴Q���O�x�Хn�M�h9�MK�O��电��Ӂ&�ȝYU��xW  �R����c�Е'�2�'R��'
��'��'=M^Q��܉]�^å+_���"�48��ϓ�?�����<����y7ˉ02i&<��EI�b�Xi;�΂�r�6-ĦYA������݃f�6-b�,
���n�E�� �K�}�v���o�I����<����?��J®U}|�� F�@�(}�����?Y��?	���d�Ц�Á��蟼���,1�,�3��Y8"�M/n?��2��Nӟ8'�d��O�l�5�M���x2�O�ٰ��S�R4{B�@�V�y��'R*e�*�0%�j	 �_�P�ӡ�Ҁ���I1�� p7h��Q���"�>����؟D�	̟p��֟�D���')<�=�h|�v��*���t�O��?I��ih�Z��'�B�aӆ�杪�̥JsĜ6(��i����!Z���I��MS&�ie�6�;�6Mb�h��:ސ���O���E�T�&�X����
H�(!S�C�Ky��' r�'��',b���O!�Xd^�J���э,T��I��M�a��?����?iJ~���9PjI�	L�����vO�6	t��&T�|��4=���F!�4��i�h`����Cڈ$c�@ՐD���揎�U���@��<���?*�D�䐋�䓫�D�=}����k��W۶�X@�A�N�R�d�Oz��O��4���`�� ��y���*2yʥz��I�f�T�/_��͓n����Ny}R%u��pm���M{'j���\�Q�GW6=���ٶ
�#g>T�4��Dڪn�R�z��`V��֍�1%ZE"�#�m�֐�Q����͓�?Q���?Y���?�����OL�	@���zd"k�Ț�Uz��'���'��6퍸�)�O�lZv��=D��]ʢ\ ?�Y��g�`��[L>����Mϧi�.e��4��$"A�x�q�K��x�:$P�i�� �X0aA ���?�
*��<���G����FV'I (�{0,���O��lZ���	۟$��r���İ��AZ�q�*X9!�A���py��'��n,�T>u��<)��c�<?g�@�PG�Q�(�a���Ѧ��-O�L��~2�|�n�
)0�Z��~'
Õ�G��x2�q�����%V�:aφ�CW�K&��"[����O.�nb���㦙�5�C�>��B���
G�h4S ��)�M���is(�Ã�i��I6�qba�O�h�'$P1B��?����Ł��D40�'��IW��\;��R����*%s�`��-ӻ�M�q
�?����?ю��q���bZ򸐂��v�j% `bƩE��lZ��Mk�'�)�S�f��nZ�<���)<݊�l�T�m0clM�<��AX�=����ӆ�䓼�D�<A�ψ�,Y��9 gI?QWI�T(y��9۴+q\�3���?)��q��i7���B�E�o$ h�I�8��'��&��&�fӺ��c}
� z���i���l���l�h7�Q`����H�fي);� �[|�S +5��@��=�1#��V�-5��S8D�D@��ˢu���ᖼ`���Ҡ�ǟ���4>}�ز���?ᥱi��O�.R=z9`-ǆK�r�ۦ�
7-�¦e�ش]�V�� '�f���Bw�lT��BB�U����j�ug��q#���%��'Eџ� �E�b@����D��ɂAa;?A��i�p��g�'4�'��}h���
*48۱�@�<� ���MC}B�yӈ�l����Ş]���VF�^��Άf�`%r�"\��McR_� &&Ѥ���7��<y��K^,P@�
[�dt
���o�8rߴ\_(�b�Z�p�Dm]�o�"��������ƛV��u}"�wӶ4l-�Mkf(�WG�9��'GP��c/�D�:0��4�����LC�	��'o������$X	�)�Q���T�J�؟Ia�?�OP�I�Ƅ�=}v�0��2_Mą�ON�D�O�o�*1���'KS�v�|�����D:�k�e����b*�'���O��dx��	�$B*6�'?�ŭ�ae�)�cњT���P'�99Ui�F���'�h�'��O�|���)_���dX�z�ph���	 �M[�摒�?!���?�)�d�k�A�.c��@�8F��\i������OnTm�<�M��xʟ[�g�y���!��q�j��A�P�{�V��&���|J!��O@��H>���<�|������dE�k^~<)�i���j�[53Ԕ��d��(v�����O#&�R�'�\7M8������ߦ�Ro
	u��Cn��u��)� "Ƅ�M;��i�� #��i���uI�ޟʓ0�Ar�J�.��0r�G�o������=|OX��mU�%\:,:B�N-T�rب&��Ҧ-"s�KƟ��	̟���D��y�-ϳ,����1��+>�� ���6��Ԧ��I<�|�4%�M��'j|t�I^��V!j�NH�b���'��}�Hc?�M>I,Or�f\�@��NZ&#8��B�#=.p=��ɫ�M��P�?���?��%�Q�b�E�نY��!"�eV��'i��ΛV�~�bY&��[ƅY�Z���Qe���Zt:?ٓ��:YIrԩ����KM`��	�?��'�m��I�6%V:V,�q�JH�<)�e�$��� hѶ9��Xa�L��?��i8f��v�'M��i����]�~�LL���� g�ܥ�! �"ea\���M��i�`6���Q7M:?y�I���#�D�S�V�]����¢&�$�$��' џ4�U�ҜZ��Ճ�OQL4"' ?i�i]B�p��'���'������D�wr���dƁ$�D�F�k}&|�\]nZ�?q��[/i$�a�B�C�0�H!��K�?��E��o�%P�ʓ+1F�;F	�O�@�H>.O��b�Ώ�@�M�B�O=Q���'D�7�L<<����۟�����!M0>�,�b/L�P���]٦��?rW�X�ߴ�ƍo���i�ŋ7�vA�(�<����B U�(��7-/?��K/gH�	L��䧽�+��©IO���p���:��M�<���?���?����?1���hH#̌L�s��16]T4�p�܆o���'��b��P;�=���DG���%���5mߋ2��P�(�9pJ&�����ēc�F!{���cn*7�??3+�>8��(S�-4Iz���eO��{#I��L$���'��'���'�T�!&��p�u+U�B�W�<t��'�P�\ٴN�����?����I����y0n(h��@�����	���O6�Q\�|�4nP#*�lCFNѸd��ChO$H�4:掅!�M��T���w(�� ���� �tx����!�r8���Q���D�O����O���i�<��iLJՓF&G�*�޽ gP2;�!A�R�i`r�'�"7M&�ɞ��r����m��M��j� e:� � �4��m��4���̰$��J�O�	
b��	��^>&��*Ҫ�=���	Ay��'���'F��'�b]>5{�i�8b���rEj��0��Z�%H��M�T�P4�?I���?)N~B�����w	��`��S�s�N���H��
	:�hz��}n�$��S�'$4��۴�yҊX��T٩p���b��� ����yRI�
hh	�������O��DI��j�`�K��W����ىn�����OR���O��f�E[+���'`�EKb���pc�(k���!A�4V�O~A�'�B�ih�O�(9d*�	S�E�"� ob��a𚟄��(7��lږ��
o���ݟ��B: �܈�A�_Ev��f���$�	��ꟌG��'kҽ Q��0��=��/�<�iq�'^r7���~��c����4��KǸ�;a(�5Z��b��Wy��� ڴp���n�)*������E̍16��d�Q�+O����\�/k䤠��K ��@$���'B�'W�'w��'P�-�7,��%0�n߼-�ta�RW�0��4f��h���?y����'�?�����C2��K,(�"ƆR���	:�M�Ѳi��O1�:$�BDJ��&�P$��{U~�j&�8^�*Q��<�q��-�j�� ����D�y�T����a0*%�b��<LȀ���O����Ol�4��ʓ[7�f��d�B�L&d��Q�/�
�ZL��!_�\���j���:�Oڼl���M�e�� Ҩ� +n��r��Lj��!󊟱m@7M3?Q�`�+%�R�邛�䧶��SO#xKDa+ӆ��!�����<����?��?����?1��4�Ɯ{\Ĉ���&#��(!5!D�20��'��Io�fX@f�<�`�i��'�މ�C���zCrQr�/�%?��t2"�=�D�������|zD,�M��O,�S���U=���C�N
^��T1$�����Tv�Isy��'�b�'�b�K"T��e{��ӫ6�hܙrl0Er�'��ɿ�M�CB����O��'>�4#G,ԙ3�氹e��#���'�>�C�f��O�O��
� עV�{(�Qo_����`�e��D��=�@�Hy�O���0k�'5P�ڡ��?�:H���н|�����'���'�r���O��I�Mc'ʙ�
P6�g�\�B�8`�.�N�|���?1�i��O��'6M		?�����B���@=���	Ȧu� �@Ħ��'�@L{�gE�?�Z�[�\{E��o-��IЀXY��5Kcw��'r�'���'=b�'���p�|�:$ ��u�b}�s	�1ws^��޴-6!���?i���'�?Yÿ�y�G�:Kf�	�(F�P�ұ�d�H@|��Of�O�O#�@��id�L ��xcd>�zd�4(U�[�s&Dm9�0A��ON˓�?	�w�.= Q�PI'�Ȋc\���f��?	���?1���$����A�M���T��䟤#���Iv����%XY��q�Fx��-2�	0�Ms��'��'�Z���� '�Dt��ٵ(d���O��į�T9R�Q��=�)^4�?)���O�tj5�]'qL���Ќ�c=��6��OP���O ���O<�}��R@LI�*ޜk�eɰc��^y��z��Q��v�T,��'	�6-4�i�A{��/��h6Iͷ@�08qF#v� ��4�2�i��m��i
�ɶAJ0\Y��O��-�\;Θ���G�j^�#�G�`��]y2�'�"�'^��'���	�y����B�Ǧ'���^�Ā�4N�8���?�����'�?�`�cҽ۰�œo�.�۵Ã����M��'9���O-����Jך*gJ�� G1�~���Rbt�	�R�L�����N��&�Y��Hy����NAD�Q�ҤD����!�G�b�'��'W�Oa�<�M���#�?itC�ܲ��YV�4�P�ێY��<�	��M����>i��i�b��f�N�)�e�*�r��#�29]�H�I5?f6�,?	#Q'_tT�IK���'ѿ�R�2�2�i@�[�d��r�c��<!���?y��?1��?Y���*L@#b�!�h�6\6dd-�G��'��d��M0�8�@���M#K>15��0����a?I��P2ǋ�S��'�>7͘��)��
6!?5�!U�$ڕ�-O�"���㞝%"�! ��O�ѺN>	(O����O���OF9ؗ T�Yi��K߬:F�2��O�$�<�U�i�H�A �'��'�哷:�|`�+X	,'��e��&�DJ����M�A�'!����2y�&�X@�.wت���D��!�cZ�L�.�
Ǣ�<�'f�,����T����!��q�$H�C�"<B���?����?�S�'��$�˦U��f�+�(�HGGðm�}�Q)�t��I͟���4��'���FϤh1ٸ���6/��IF�ĥ>t���pӤ�KAam�z��|]+%����$c.O�ty�g�Zr��?�l B�`���B�+K�[s��4,�a��D������4�T� r9��[ %G�mJ,1����X!r�O��NJ�x�E��@��	/Ŭ��'B�qr\�Q���je��z��qm�q]Ω��\�/@�ĸ�,��� ��d��(�%XC�J��*Y��o�me�I)r[�;h�dXQ�@�p��	 슩P�Ή��_�#	���ת�<ܖȪ%h�#}��ӣK�d���`Z�y���&i��y"H|
�S2� $-�q��ߛGX�*D��
BnMn�����I������']���)�70��B��,
�)[�Jr�����C�O���O^��3����KU�EH<9pA�yQj� ��D��Mk��?i��/�p����?q*�|�d����Fцk�&Usb���dn�6��'���+��,���O����OJ "".M=`h����c[��´`Ц��	N��������R�D.�MK|:��LG=`Ϙ��햿'����'fF�25+���D�O~��Ol���O
�a�@VSD>=��ל$~�p�do�=@˓�?���?�M>����?���7yO**��]�<�np�&'j��k K�^~��'���'���'6P�dݟ�YӡL3z����2�1T\<4i�i>�'<��|�'=��	!R�H�4��pi �	M�:uK��@q�'*2�'6�'TRFx]��\��V���E� �v�≙D��M���䓪?��JH"u!A�C�I�.��T��b� 
��R�і_ְ7�O2���O�$��]��'�?	���b�&^;�H챕��"�*�Ӧ�	��'D��'�tL��H�6��I��n��$'�x1k��GY���Q��C��&�M�Y?����?���O��P���M��ܡ�g�B��i�5�i+��'D���2�ӕQ%��R�!�.� d�Q��7�\�FKB)n�˟�	��T�S����<��eK�`Y,�*���Ih��T���Oś���[��O��?��ɥ,�DU8E�X�-Â�R�����J⦉�I埨��2\��aR�O ��?��'���GI�?��0��	�:	�~���4��C�f�������'�r�'��Á�����&���R�p�aU�{Ӛ��ӗ���?I��?	M>�1q4��EP�f�]0��D^��'����|��'���'��:oz�P%��3xX4�5I�.	�a�����<�����?��p� $+��,1���*��%�!�Td�$�䓽?���?y(Ov�P���|�3���܈�T` �(E"�;0�@̦�'�"�|��'�%V�T�$�Otę�()��Ǩ]�+�	���	��X�'Pj(�~��Ot��zwk��E2ą�ׅ��;��ǰin�Z���	������iO����y�d�a'�(RÂ۲|s�9"�[���'w�_��ᡢ�
����O�����Ɲ��_o��b��C�2H~�(��d�	ǟ���ck����y�IC25+G*?4!�M��������'��R�+e�>���O���ԧ5��];r��&�Z�#��N��Mc��?���S�'�q��A�b 5��ы��q5V 
u�i[:��,t�.���O@�d���'��*?�Lq��\-����0��%b6�h:ش]�Ve��I�Oظ;�j`R��[Ə+y���a���Q������	#cΐ��O�˓�?9�'��+�Α-R0���fʇ��([�4��C�����D�'���'�
tK�g+e`�IY�<Y~��wf}���¿5*��'b�I䟨$�֘�otIY��
l�*�FZ����P�e�N>���?1������!v�,�p�.��k�	�d��A� ��V̛M}_�D�I�	��@�I�H�
�F�+qp��3E����	�g����' ��'��S� �a��#��Td'QD����93���I��M�,O���"���O��d��+�	�
ʒ!����K����#��y���?����?�(OF$�tiE_�Ӳd��I�]�5�P�Pm�;@�p)�ٴ�?�M>Y.ON`� �O��O¼p�G���Ĵr�)�/Րy[�4�?1�����^��'>����?��a�n�(`1P6yۑg0��O��.*|�b������D�C9����5��YV�����M#*Ot�xEHTԦMث�f�D䟔H�'��az��ʜA�J�{�$�JbLJ޴��dF�^)�w�p%'>�'?7�׸L��D[6�S�qz@��GL>^Y�6솠h8�7m�O����O��	�p�i>m���	(d�ٖ��
I` j�ȋ��ܙ���֟�Iby����'��a�O� *����]'@�"� H.27��O���O$��ɘf�i>I�Iq?�k �g�٦k�*ƬzH˦���Wy_Z�X��<Q��?������o�J�@��ek��iUZ��
"�x�O�"�|Zw���YՉ�,me�$�����KN��ɯO��r&��M�K>������O����uBB�pU(� �v���i��?��˓�?����'���'�.�3���/f�P[�揋5h�h3�+����y��'���ڟ���@oj�+4|��b
;u�u�������D�?���?92Ə�y3$9nZ3}� �wj�����0v�LOV���<Q��_f�ٰ/��$��p�� ���d��G75��mZ^���?���T7B��d��O≥-E~���ךW�t��#D��6��OZ��<�v�͖V<�O9"��5Ƨ�!����v�������䐿�V�=��?-���N�ke68�*��-b�� *gӾ˓}f�� '�i�r꧳?�'1��3oxr�ȆA��lC���.s�6-�<�j�!�?Y�����4Eh� UJ�8s^�9�����>�
1m�&�HE��矸����tyʟ�P�@�R����*܂b7B�##XϦQb�J!��b�"~2ڴ5r�
�1���1�-�5&46-�O���Oq��$�<�O��*�"h�k��0�˲�,K�T P���Y�
Ī�'>i�I��d�	Mh�L��BEzM�py&舝y��Jߴ�?)���Z̉��D�'�rW�H��&�r�ҵI�c�&F`'D�&�M{���������?������,F|�#���b���`��0���	e�Zy�����Iu��AyB�T�|0P���a�p1w�
�QD���d�'.��0�Iꟼ�'����jx>��� �Y����"� 3�N�q�M�>����?q����$�O��DQ�	J���D [#d�(�#�]�U���	o�z��'���'���̟����}�t�'!j(!��9����2�Ǉ ��	�j�P���Iʟ ($�a�|OP��J�5���c!C�1U��ói���'-�I�Y���HM|
����1���a�K�. �6��!T, o�_yb�'�"� �R���D��5��Z�s���٦!Nv@6D��e�%�M(O��ɵ����s�����럘@�'b|C�d��!���q#��9^n�Tܴ���B�O���$�`��^�D�Od�	k�5��5� �O<^����`�i�|h�v{Ӝ���O8�d��>l'��ӨX������	 u���[�G�%�2x�ڴ^N�p���?�(Oh����O6|{���!�fz0cL$'� ��P�\צ���̟��	�5�J<�'�?q�'V��(u�[�6�h�W�ɤk���4�?�*O�ex`*�Ob�O��䳟H��v"���
_��2��6%c��DX�V˓$��N��@��U"#�Ԍm��*vj{n$H0Q���Q��,\N��?���?�/O�I��J�v����I�g[��ٗ���`�t��'D�	����'E��'����:��A`i��d�DI@� 9`�@ژ'���'�b�'��s�p��g "��T̒V��Qq�}������Q��Ms+OZ�$�<y���?a�� ���Γ6�t�k��G?Z�&��ᖐ/�pPBֺi���'hR�'��	�3�P\������٢~2L0R�☖3>P�ᗮm�4l�џP�'���'F"E���yb[>Ic� ~͙�bO��pa�?`?���i�"�' �	q%�lX���$�O��i
p�8�(\?AyP��R!���Fi�'���'���Y�yR^>�	h�s���o�PG �Q (�`U��ƦQ�'�p��dӈ���O���$�ԧuG���V��@*�c��-0 Fյ�M��?Q'N��<�VP?��b�'02D��
�
�p��"<t^J�ov�Z�Hش�?���?��o
�Ify"«�����f
�
�JI���O�4��6��?$��2�$5�S�芲B��lT�d��6F��Yw�[��M����?��1�tk�S�T�'��O��)�$�* �� �#� t�V�i��'�����i�O>�d�O1g�)��;���5�������I�ɇO����O��?�/O���<(�Q)��kN��v�+�[��S|���'��'��R�A���8�j�d��f�2���SF�i��O���?I(O��$�O���3����D�	YԼ��
���q?O&��?����?�(O )��J��|:� W�h�a�e�X+tcz$�t-
ܦ͖'��R���	��IU��Z��D`��n)�x
ԫ�,����'��'rW�	qŬ��)�O�DI�U1���M�j�l� �֦%��fyr�'���'K���'?�I�b��pɕ�*eEZ\)�G��,ڴ�?����$|Ph��O]��'��$וyޭr�F�2K"0�`��>i�<듴?���?Ag��<	+��D�?��4�:����ۊ5L��Ԋq��������i���'���ON�Ӻ�=E�I#�C��l�
�ɴ���������0�9��O��㑉�&a�b�x�N�~7��P�4Y�4�i��'2��O��듳�d�|}�=z���.Ƽ�	�ΰ6��o�\�����ܕ'��z���#,� ��"DԃaX���&�B��Tn�ϟ���ߟ$x�!��D�<A���~��Þ7�<$ ��\�@�T��"eG3�M�����$>�?���柌��C(�q�3lm���r(ɤIː�oZ� �!�����<I����$�Ok�%*�l�CeM�{�̩D�H��ɺ%�t��?i���?����E>�2!���HKrUkb��(,Af�3�*�r}[�H��\y�'�2�'�>h5�R�tF�t��I� v��LQSh��y�T�8���L��Sy�W�5mp擌P�A�pM۴F*�q��Eҥ\�7m�<Y����D�O��D�O�� =O(=����PN�1��O]Q�( ��Ҧ�I矘��ɟ��'8D�UI�~"��d��@HI�5�@����'o2 ��i�W�8�	�����t�|�	ҟx����ɸ�Ʉ��M��_�}<�lZ�����py�Z�Q
b��?�����'CC2� 11���gX6ט%{�HT�''��'�bl�7�yB�'���I4 ��E����%�
�BDP�A�cC��'�|(��oӨ��O����H�էu׎؛~��E��żJH0�J��8�Ms��?� 	�R�'�q���rĢI�Zrx��c_w�,��øiϢ]#$n�T���O�����r��'��-ƚ(�F*k8��Xdk�[��A��4Ò�ϓ���O�?��	%be"sO�%l��8��P<(_�(b�4�?����?IתX9/��ey��'a�D��
�9x#�d3�/G<���'���3G? �)J���?��x��&*Q-�*՚���8 {^t���?��5��Ly2�'x�L��"(Z�k��d��zf���c	Hz}R$��y2�'A��'p��'R�I*6T����ĲNT��Ƨ�5V�X<a�L���d�<q����D�O����O�|i�H�Qہ��0�N��D+h��<����?�����۱M����'VkHxFC�SJ�'f�	\e��nKyB�'x�I˟��Iџ( R�g�����=��*�f7b^��Ё�����O��D�Ov�o���#�V?���=��P���$�z�sw����Bش�?�(O>���Oh�DNLZ��o?�	�#i�,�u�ξr�Z�DH��������ܕ'kN���~���?��'d��Ͳ' äs>1�S΂0S��S�Y����ݟ���3 ��������ϟ$�'j\�|b�)�(��d��$er}n]y��F#&E"7��O��$�OL���d}Zw���yS��_��1�G2V�@��4�?���^�N��'d��CܧzyL8Yamχ�N�s�iH�5�l%nڙY�����4�?Y���?��'.��Py��I,o�0����
�,�z�6���`_�d�O����O���4="9 �eߑ$�:��L��7��O��$�O���)�~�	�d�	D?Q��($d�p��ĤjMpl�����$�x�c�����'#2�'�Zc��\��%�0V`�
�ϋ�p.��4�?Y �Ӵ=��O��D-���ly�c̛h "䢤��^�xPjs]����Ir��'9��'��[�P*��2=�*�ql�:n7�aAC�eψ��K<����?I>���?�F��cO����a�ɒ�GK/�Z�����O��d�O&˓%H�=�e;�B������u֊�kaLI��F� #[���	ӟp$���Iӟ$[w�Fٟ�����i�n�Cd���XrL��c�;��$�O2��O��"t�&��TiZ�}	���/�:�2��0_��6�OV�O��$�O��)34OF�'�X��H$��P�ꘗQ� L��4�?�����G�+�&�$>}���?��ѧ��l��A�↏kf�Pq�����O~�D�O��zb�O��O��	#���'M�?��5�#
��@�h7��<9��\���掶~����:����QȄJz ���v��c5�x��d�O�ѸG��Oj�O�>� L�� �6 �-��_�hq��iv��l`����O���b �>mj�ⱨ
�y����Qi��hQh7-�,wH�2��2��՟8R$��{�4�H�ǩX���s�I�Ms��?1�:�z<I���O0�I�Fe$�rW�U*	�T�@DW�p�7�,�$���?=�I˟d��q"��܈+����q�d4m����F���'�"�|Zc(6F,{�1�N��+Z"��O^�u��O0��?����?�,O��:�DT'5�L!���Ӫ9� %�D�$H�x�>�����?�uG�-���
Al�RTK��,v()�"�<�(Ol�D�Oh��<��ΒF(�i��N�)�smf�f!�7��.e'�'���|R�'�b�Z��d�+yI$`j�@]�5��H���6Z������ԟԖ'E��3h3�i^bJL��a��g�jH"e�ȉx���l�џ$'�@��џb͟�O^D�Ej��>ej<�&Ƈ�"^uԷi���'��	 b T9M|B��jEʇ�)�BEȆf�,��!�� M'Y��'	N!i �'��'��� +BǤp���+��".
)��VX�������M+�Z?M���?��OZM[Ƥ�%�!��X&�N�;�Z���'e�'�ɧ�'�p``����pH%h���l�A�I�޴�?Y��?��'Љ����(�-�7���GY<�c [7L��?����Ş�?E���;(80'���՞g���'���'�|��s�"�4�T�'d�� ��I:d��F5Z�N���4�?QM>i՟���'�r�'<�d�g: Po_�[�6	*�r���D�'c:�'���Z�'�0|rb��)N����ݹ>Yd8sO<����?y���?A��?�-O�E�
e�,�E��\n���v	J!�|%�\�ID�'�Ę'��Lr5nM�X��k��W��'��ٟ`��ߟ�''���j>�D�K?#�$$D�R���PnjӘ˓�?A/O��D�O@�$�kq�dٗJd�D�R�86z��] t���n�П�������IRy�ʺU�ꧠ?��&� pJ犟l�e��I:��lnZܟ�'N��'p"�O/��' ~�20F�ۂ:3HWoԸ���4�?������ϔ+>��O���'����@z��k$��$Q���Z��L�H$@��?����?����<	�����?	Y d����xC��OqVe� bӆ�P�P}���i��'���O'V�Ӻ��CU e����FE����馭�����*!
c��:���d'�ӄ?�X� ��X�R �T㓥G�7�?���l����I� ��)����<I�bJCRj�2Q�v�T
0"���փ��y��'�Ia���?!&e��+��\�(ްl�g�'_қv�'�R�'u"��d$�>/O(�����Y��.O��=AѡW)�~ȓfIm���<���]�<�O'��'���;w��)�s�BM���r��oL���'���"&�>�.O��$�<���[ք��.�(�W�.�L��/Ȧy�ɴ9���Cy��'�b�'�	�}�� �C@�
�N��Q%�0 ��`����d�<�����D�O��D�O�iB�,�Q�T(�ů�~Y\Ԙ'���$�O(���O���OP�+����;�������x�Cg�@1"Y�iR�IƟL�'S��'��yZc���ӧ#!>�yʲB za�ԙܴ�?i���?����䖈4��h�Ob�1Z���cJ��.*��	��&1Kf6��Oj��?Q��?i���<���~2g  W�H"f-�jXv���M��?�(O$�!! �M���'�"�Oh�3eF��@�����@8� �0D��>��?��H��Γ��9O.�ӜW�R���'�����Tz7-�<���-2�f�'���'���ɢ>�;F�P�Cr"�k���� �5hr�5oZ�����0<���{�	cܧ}J��J��)U���*T�H.���nZ-�P�8�4�?a���?���e��	QyB�T�5LJ�P���'v���BƖ�dkB7�\�J^��O�ʓ��ORҠ�_{40v�WD�y�`	��c�67�O����Obe	f}rU����V?�r+ +4|�E	:4�T�H��M���Fyr/1�yʟ��d�O�� A��c�H�FӞ9ۀ*>2��1m�؟(��Mڍ��ļ<Y�����Ok,���
��Ƒ�-Қi� %�5�v�'��Q�'R�'��'x�Q�ѩԉ3A$�n��l�� a�G&H}#�Otʓ�?a.Ov�$�O(��_5D��0nށV�z�*�h�;m!y�8O����O��$�O��d�<1���7K�H-6s�<X���>B�xQ�`�2�FV����JyR�'JB�'�,�K�O����τ[�Lm�wC-w�
}��R�4�	�4��WyrAZ<��'�?�� H	 Db	BE��lh,�Pǖ�4��'��Ɵ��	ȟ`��.`�x�O�[��/Lr�0��?Nh�ъf�i���'���'��b��'�b�'���O�����i
�]�ɒ�œ:(�y�?��ORʓ1�fExZw1��(�m�%T�M8&�I+{��ߴ��䃏1O��lӟ���埼�%����n=2��1ˠ"A,�l*ȅ�3�xr�'�ўd�O���R4Bj
3���#e�"�kR�i������'f�\�d��㟜��ry���Z�$"����'�V!I�΀�Q��J�Fx����'2�piq�O	+�!��hԌr~|��buӤ�D�O���`�С�>1��?��GW��і�՘ ���� ,��'[�9ҍy�'H��'*� �w�ҙg�pX�T��P�5J�W�ܢ�̚ay�R�X��e�	�:�dQ�[��(��fn@�e��hK<qd"~r�'z2�'��I�L�|�s�`G�JK�Ps0���g� �؇�G��ē�?I��?����3}���B$@É �L{ �Xw
�،y2�'��'"�'j lr�П�]3�h��r� �//�,�ѾiB�'a|�'`�0	3P6�0���qZ�
>�2U�G$.��ß�������I؟X1e"�E���'b:����	�*X���TE0NX+�c��)���O�U�~'�@Z�O�z�Q!��;�
����bӊ�D�O�˓_�(�����T�'��N�a��xv&����T��.J26�8�ɀ7:#|J���#΅�R'�$�A��!2N���&a�����OL�C��OZ���<��'��ƨ� ����������!K=�UP��iE�S��vC=�S�<N�дa�@	nؐx�F#��-�87M��-^l������h�ӕ�ē�?م& �0�%ٞ*}���
�\��F�Н�O>��	�L	
v$�,�,@�gIӪKzܴ�?���?�/
�<��'��'i��G$ZhL=h�"�N���Rq��	u�O�l#���O��d�Oj�i��-{�d�
��M`�!�E"����I�_�P�I�}B�'kɧ5&�Wa�7��")��*=v�	l�Pb����ߟ��	dyB T+�Dx�&�
0��]����3�,H5/�D�O�d8�d�O��ŦM, 1�嗰O�}�Q���Q������Ol�d�O|����3>���c���5G����-U�> y0Ӝx�'n�'��'7�lèO�uf���'5��"PN�"Pu��U�<��ϟ���Gy�c��\������,5���936|��� #PզA��}�	��D�ɥT־c��!\�A��H���^�tq�Em�4��O��4J�P6����'x�$\�t��ar!߰�>��`@�� ��O~���O:���~�@��n����%T7#6�R�"�$;z�Q;րA&J���g�5�%	t���0Kx�CF�T|,���,/�8��KWDk�%H���gg ��2 -�Vm�� Y�.����6��#�����ӋW0���s_pP[�	�i�X8��H$����&��	[�tz���U�V�s3i-cw
)x��I�]��X9��C2-�N �7$��cƔ�$�H�m ��'� ]��oe8>��GS�AL�4��]�]��`����?����y������O�eI���	?xd�a5Aަn\���g��d=�`��`�a3:���d\��ND�'>��b��'a�B�li^��j%*l���Ё@4���Ѵ�2����*�vt�V$�If���qB��4���!"P��	��`E{�U� c'�EX�Ĥ�a!��+ P��,D�,��jÛBM�Y��>g���p�	�HO��Sy��2�"6MΦr�>m�A<6�0qr��4p�����O��q����m�ON�db>1`1�<�:�+Vk>Zv�r��K�^R����7�,e�3��qx���B� ���Ӳ�A+dDd@�CĤS�A���X��0#�"�_x�\���O���kߦ��'%=S�vh"���0r���=9���R� �XX���(�
<��O�!D�!�dX�U:F���������Q�P�Mv�v}�_��!#`6����O��'fwz����D��������Ь!����?I��?Y����&�\s�P$*"������K- �G_�3�"��bF%�Q�d)q��6�܀�*���$>mk I��N��T�	�2mV���*4ʓy�B��	����D�����2�Bۤu톘���Z�<�	����肊Z.C<��2関�0X��I��ēDz8Ub'�|���:�A����#֎P��R����m�A-Pw��'�"���iޠ�����*Ⱦm��*	��;u�W +�@,ړ*��_Q��T>��|���>����"�܌XP�0�2h�yh�ȓ&��\ph�p���[xŉ�IY,�"�>���?kp���V���*`
,0���M�W���\��M~J~H>����q�	r�,�!���&0�ц����Ju��7��ъRhÞ4� Dxb)(�S�$'�7Q��JDM�Z<���R�&$��'����Ʉ/u��'�B�'8��ٟ��ɛ!i���#��j���N�"���#(�.�
I�e:@�HǓW��-��S��b�"e������X�z�9�E�{,���'����F£H���R T-{W��c�'E���?����<�3m��j�Z5�N]ݘH�O�H�<�ܓRS<LR��O;O��y�ń^%�����d��v�loڗ/� ��� v���h0��/�@L�������̟�vd>��I�|z��ǈ�M���x��#EHϾ:����k�8��ɸ%�8�BM��A3E
B^���Sh�5M�pK��'�V4��`ћh���h�hތM�X�" Š0��6��O˓�?1�ʟz4:�^%��䪐��
4A�"Ovq�U�O�E&�U���E
a[]�B5O6���'X�	l�vZ��*�d�|��P,�@#��+.��Q9a��H��z��?�������B� c�X
�i��8� ո)�� ���BBP-I��m+�DW;dT�"��I�8J|�A��4Y�z�J��#8���>��ZŒ���*�V���N?�����O>:�:���Ę���H&K���'
�"k�-\5����+[]&��$K]��0>Şx���b��k�	Ls�Z�<�y,F���?*�<�����O���O$`S�� �Aݬ�)ȅ�'��РN��$��x��bь���,]՟ʧ��?Y��;49v�LuP�*1�P�&m���8W�bI!�`K����OB��a �[��P�S��',�XB�'D���D�OP�S�Sݟ�'�vA$.S*}�T c�S(mx0��'���o���n��Ab���q���Hi�'���wwz��@�e,��Q��9��m����?��n[ 
9.����?��?a�������OJ�;�C[��^h9 jEoJ��!E�O��ѵD�	qD\���-jb� q$H-���Z�J@�Pt����%��9�8lO�J刞�k���P`LK�?�n-��OM���'s�{�	�?4aQ`N�]���ǅ��yb*Q1A��3&cәXaV�+�O�6~Y�"=E����
z�7���&��|��M�(���"�,J��$�O����O�ӎ�Ox��b>�	"ŝ��D kC̓&O�K��e���;�4��l�q�'��9��}>���$VQHIM"fP25P���l�.����MV��E�U��8�E"Cm�5����`Ə8�M#�B4��<!�hB�idt�*z�<�7K�C�<�dK�U��dƟ��h�]�<�2_���'���%�|�p���O��'���T��d�
ؙf�W�^Sd�#T��:�?���?iE��!�?Y�y*��a��b�{N �y'G��R�FX"G�I�E��
A���R!v�@ҭQ�X�k��x�'W��+��h�r�@�d�{NPe�,�"�����"Od�[�n��OC౐T($c�E:��'_�O`�����^v���3�@4O��"O�9�e�o����@1o�HH�"O�
�i��	�p���]�n��}��"O�u�����܁�o4q��A#g"O�ۣg��)�r-`SȈ1H��A)�"O��� Br�;���7	b�9D"OH�ڠ.Y?؈�{vIƙb�\�5"OѲ�f�SP�bhQ0A�����"OJ���f��=Bs���t<�ۃ"O�tH��S�2qd�w��x�uk"O\lJ�l�Ԇ�����yj� aF"O�$)��#?���'�
�b � "O��zG��=&V��d�\a^`�`"Ov�sV���;�R0$�<KJR@ "O���T��Hr��
�B�3� �"O�
& �5�[B���Y"�2"O.qegj5��G�9|�����"O�u�Ѫ %E���`�-�:Jٔ��a"O:�wF	��Zy����i�����"O�����-^��|��Ȗ.��Xq�"O���f@ШYWF<qA�rkF6"O̒�gµ.���WF1ax�4"OY�Bj%܈8[��O=3��`��"OЀ�t�R g��(s��B�W����"O��;d�K4-{j��$���MH|P"O[�R,�H`�Վ#=�4�"Ox�X�톻<*lXp+���ș@d"O����H�6Yur�Y��V�E�d��"O�Ż��P�]+�����6�P"O����O�4J�CP�U�j�c"O
��qDCr�J�+��/�%"O�l�E�ƠL����䏚o����"O�i���q�5�Ӂ[l�XzD"Ox�Ei�h^ jr�K-v��E �"ON���k;7� Ʌ�׷�$��"O(��V�H�У�),�%�b"O�e�E�mbej g��>�`Y�"O� �`�BᎧj����7��0C�4��"O&Р��x�Q�0M#:T�R"OVYK��ʊ,�T ����~�TP�"O���Q�&WV��R⋴<��5��"OT�Bv-ߕ
�>��tg� ��a�"OH��U��08�$ժ���T�nIPt"O|iAr�@�d�(�Z�C����W"O`�q#�'�� ��A| ��"O�Hsaɐ2�k��ȇ"f����"O��`5��&0`{e��1fF�؃"O�t��aWv�@x�A�0s6�� "Ob`���1,�]q��mJ��	V"OPy3ÊЊ�V��5�E�R"�%
c"O��B�	�SД&�èT^T "O$-��A1KwbP���F=-ԸeQS"O�ВgG�$R�L�"�D$ǜ��"O��#���3WpXHP��K�Y�!"O,������2F �6�@�#"Oh�Ye(�"V�fQ��K�K����	�Q�	"eo7��Z�#ł]�Q���3#b־��B�I��4��`mٞV⠩Sq�՗1Ӧ��o��R�M<�)ڧgk����A�'[��k�d�H�^)%��+Wd�L�N	9��i�2q�0�u�	�d�;���w�8��Z�ZCx� �U�D;1&Dkc�ر\]���JXX�%�d;�%�j��˧>��M�SK=6��{Ƣ��I2Ԫ�'[�p�d��>8Rd�EAL�m_�2�G�J�#$�)��G[��I��i'V�Ū�o��݅�	�m/F��E��	��D��O�,�ԩt!r��.�ȁ$�O�]�ԊE�g.1O?���pv@K��ǅal�i�"O*����D�D�n��q	�+Cؠ8��x�&S�:�	˓ai;��τ>�|`����8�ZɄȓ ��y�����}Pn� �ַ r����D$�$��e/�e(s�óR�<��ȓ{2�$�� E��w���F���ȓN�l0��/ 6,Q���p�j3K8D� ��
�lVdT��K��Q��p�0�9D��R�.ݹ*p��yʒ#W�z�a�+D��Ӗɋ�&�ܡ鰏�@�f��֥*D�l�r��H�u��1FWH� �,D����у1�� ��� ��$5D���@��`^%W��2�2�pT�6D��	Bm��
��}�e �6��['/:D��!�Kȇ!$�z�g˜Y����8D�(�!�Ec\񵦌9kǔ��S	,D��Gk�� Cw�˕]�px��6D�dY����P�4�y�%˜=�x���?D�(��F2
 ��"n���� 2D� �w
C��X�E�?8�^�1O�8:��[�,j��u*�*;��$�"6!@���}�=�2	��,'!�$�4��Z�l	�f�Z1[�B 4��*Ť�"6N�D`*3 �=� ��$��$)w�.i���fD�! .҅2���*׃|I�X Ƥ@�2}��b�D�G�g̓CN*`���8=�:4[E��L��u���GF:,� A̗oV�)�B��1�j�SE�A�\�� �f"�Ɇ�	�R����1�z�޼j�(���ቹ����3�� ��$�9",�ɁDꕒW���o���"%�G!���)��Yk%n!N�6%+"c�'��*F�2M
�DǸ3F.x���7�9�!���Z�_U,�&��j`�(��FҶ5�q���%7��!T��@���"�mZ��F�(�HD�J�����a�L<��y�B(��_�p9P�H�*A$����}�R�R*3P*�*4�M=���k]0+�R���&��h�>�D��|Z4�*sdƎ�~2$:�nd�u��<h��2�Z��0<��#ڭ_ ���㍕M�*U̓��x����,Q��\�E�a�:�'b�$����)2B6t*�ˋ?�'���o{�Qr�%`��mIC (x�N�b���8T�$8cm�x�'0�p{�a�Z�? �y�CT;�a1�(�� Ⲅ�'��\�:C�K6��$��(��Ɂk+S"�]��`���ٷ��=�6��2!���	$��];��ر�P$�-�iލ�q�@�s�f�;5��$�`���ֈX7�;Cg�S�H���'+r�p��QMn��A�U�Y���A%�'&��d&�{|Ȅۉ}���vp����윙2�N'khl!ق��4�<�b�vHU�#� S���&�%G��� T�<��U �&萢̌�a ��qg�U�AZ����o�5=�P$Ve�.����f���@܂��3�%)�P(uO��)�X�NZf�h��2U[����Zr�O��ZE�ɮ'����`�BV�t��S	�q,��x�ȟI�.%bKןyP���>���?'U"��+� �|����lV��3�%C�<���-Kɰ	���'�2%�'� P9�Dxމ)���/5^n����R�7���9����r��P�햚],�{��X���OԵ�${�ޙ3a�-W�±yG��1�"��s��Wn��p�#������ιs�i&�a����#~�D�_wv��Sc[�bv�l�8)��̞7�Px�Վr��YǢ�v���g[4
�����0���Se�*L1&e�Ů2e���*[OT`�5!���rm$)E6�#�j�')��1�c+�YX��ad�Fs�.l����^ a*�GTx�i@�m�����R�Dd��O�Ʀ�Ҥ�u}�A�J|�'�hm��o�P��5� �� a(�0��(lhlc�06~4�&���|�]��H5+�3o�� G�B�$]-�J1#�/���W���<A�!��&@ e�&K�&̺A��5@��(҅b$0N@�ba۞L^}�{}���l����/�����*!^\�@�W<��D{��T`�a~�*2J�F��6�+{]�sF�\�e|<<��Cܶ�����O�,�����>�6E�֌��|�C��^���'bC�-MH=Ӥ��7 R��8Db�x5(�sD%?�I��\C��[�G,&��S��r<Т��qQIA��^K�N	Q$Ʌ*~����$Y�4��\�p��?��HB��O$N'��q�Y�`�L�N3"��Eꯟ$ۀf"0x�1��������� Z�i�& A���ΓN���/BIttJ����"�:l�f,M"5�`IW�k
�*&�3<O��ӱ�ζ%?������n`M��]�mY�KGO���f
�&��^��)�MأU���l�	��NpC���`�I4�V,Q�f�:�0?9�d�Dxj�A�H�6/�l�7`D^̕�t��> '��j�Z�x0UB��<a�3����'���i��)&�����?nzD���+��P�ۓL��Y�'(����@І0�&�h���O/���Y,��MC�<��&�W�&1T9�)�	���5���$���uȃ#�n=R�Jؿ�axbn����Rq�B?q��s'D0Ja
�~֮���Y�D4:sJ�T&@�c�J�1*iFR��+U"�Sã� ʺq�e���L̰2��t�%�2I�.��e�O:�	�T��OB\,��ƜM��E�rL͡6�*�����wFQ>��t����l�B*
R��0�5�����d�5�P���O$R�c0c��TAtC[��xi�	���y�SH�<�%Af���O����j�1��[��:_J�s"����摔'��}+Eƙ�2�D}�D���F`JϛX�m������\�M$�`�޹uL����Ǘ��sU;h�vt��F(dS\�	���!	GP���`W�	�l��D�e��8u�Z!I��Rt	��|���³�!��&/q���o#Q'�]) � ;"
.@��L?�y�'x����S%�<UѤ��H��QD"���(�~��qᇞI��h'�F<8c�$���_�~雰恫6��Ł�fO�h�~�)�oݾ@Q(�}QжB�W�d-���'o�jt� �����,�S�'-��- Uj�"A��dcǈ�zL�g� V���d^6؀㵥הa��b�b�]���U�Ѽ-;4�#r&��{�����;,OvI���]Ow�D��!]>*<HCJҲ[�X!80"P���`�HˋT$$,�a��C���I!x߶a���߁tɀ�X$O@l�FO� y5@��zXt�* ����9�&	�S����|��EezB)HoN�x�h���F�M�<A`.ǽ|7�9QuZ ?F�vK7@fr��s+�3����kԂi��QC�t�ӈES~H��w�T`
@I�3��qS�T)E�� ��"�@W�����c0���&���M�'�P��-P%P��q���5s�yET%P��TjpQ��X�y�������1eP���,���ه�Z<RNqZ��|���I�=H�����y'KB-hT�w�ڎ+���!-μ�y�$T�:$D��,�^�P��	GRu��J���M�6 a���>,T�V�pS�>q'��+���0��&%�ذ AUF��P(��DE0���4倅��GŪD"�[���#��m�T�H����P>0푟H���To�h��(����>�y[*��F��2֐�Fm�;/X.�o�~
4��&$<�I@��G�I�:A�� �D��MB�'������|Z��.~���'(���"/> J�� �'�D��)&b�~=#'IS5b�䨒�'�](A�*����"��a0��C�'mV��Dh��A�����QH.���'�lm��CϏ3s�%:��J�D%��'�l�{�m�+2@xӑ���5o���
��� 8p2��;?b��B0�Hm]�T3�"OJ�x!��+�n��E�;KB�Ͳw"OV��N3����˶`l�p&"Ot�P�ś��(	���[�Z���s�"O<�`��0^l\��[�N96 � "O(��#M��=�x㠌�R�.��B"OH)CGғ:��<0"J��Vpb"O�LS�p��2��'I���"O�8`d��W~���"�,<��"O����!Ҹd�h�b#����26"O���	�x�aj#T 4��<�"O�I�'I�b����5ȟ��x
�'�p��!��w`�� ��Ts��
�'Q����'�����2�t^���'�z!�+b7���$cd���'2~��d�8r!�"�^?���'�:�2��B+C��y�!�+%�.�*	�'~�q�����~�8�Q�k���'0�̓���L�а���&g�j�	�'%�-���U�4 r��f�����'U\�d 7�Th��`�"���')b�z �.PG��9d.I�$�*�;�'0h48^H�[w55�*�a�n���y�͈�6�z=��jC�1��-(錤�y�XT�A�rOҭ���K4��y�d�1���J2/| r#��y"eϡ?�*��pI"L��C���ybP�Z"��[�c��\\�s�P��ybA�8��5�"kP�����#Y��y�ɕ�A�񐲤�=yجV�Q��yҬ_�	�81����pr�z�T��y���K���q��l�����	_��ybʺNH���-�Q��U��P��yb�J)~dz��ӤPxBk��y�ه	0b��-P~����$�y҃ �&������F�@�x���[��y'A�.����<s���;��#�y�*��m`z�k���+o�
|���y��<r� ��FjL���)b�ߢ�y��oД;A�ňfr�d�֠
��yr,Z�McD`�cA�b���a���0�y� >K* ��O[�d@�j���yba±p���aC��e50dr�m2�ya�8��YJ���Z��e#�bӺ�y��%��Y+ ?�z�ȏ1�yrFQ�F�$SE��,=1 |ђ�Ϩ�yr ��+��@����7k��:w��y� H�*d�D����6��͈��y�ʛ��6��un_�{�2������y�I��24 ��2��'^NQK5�V��y��ȦnS*q���ncB}Q�W�}N!�� c8tA�Wd�r�:��Ƅ�md!�$��Ɛ�sj�4i\�ysC�z!��:<�S Ԣa�q�b��}!��B/��T��m�L�4�)�i	�.k!�dv<-P'���.Ǡ��S�U$-U!�d�LM�A�#�I�\X$kX�z�!��W;{�nR��џt�zQR��K6G!�d��O|.�s"���xċ@g��!�: T�1�fд� ��%a#�!�V�KrĠ<G�TY��7!�b�J�Y�IY _j2�r�j��!�dA&IM�����<RXl2H�<n�!�D*�DP���ݳ����4.�!�� ���W�J3R���a�B�2\����"O�|h��C�4��P��-�4	92"O���W���(�u�@4��YC�"O*d8ň�K�y	���
et�u"OTY���U��tSA���iI���"O�I3�dU#$8�RD�,B5�l��"O� u��h$�L�}2V	f"O2 ��+�ܐ4 �`-��8�"O���G�{�QZ��� $~t��"Ob�`eY6*M�p�΃�t��k�"Ov�`�㝿=�*��4hJ�r�&d"O��;���$�6i�6 �ND4�4"OT�K�-0!�E�E�R�2Ʊ��"OZ}��8g)��A�-�=�ژ9�"O���+P;-0〯ı<e��J"O��P���9.fL\���.4HAq"O�I�W�tJ捈����e�l�;v"OP�q��H<U(pL��J4ւ�a�"O4����q̔&@�F4�""O�i ���2�f���aݳe���"O�9c�MF]Q��F�	����"O�]�5i�~^�S�O׫^8Mh�"O�a��^�X�>X���h ����8�ŞBbx��
�:T�J��)	$ ӌ��h.�`���&:VF���LoaD�ȓ*Wr�Z�#�[�2���K�$n�L��
6������<���yڱ��Y�Lx��2����V�2 f���-��m�g}����R�AE�̅�(8��PU�dl�AC�(T&��ȓST,��N�;��a���J�mӦ͆ȓ���[��1l7��k�D�X݆�L��Q�` ?'*8��FWp�����+����@D?֠����n��ȓ<�����C�AI�Y23b_�RNVA�ȓYJ�)&Dsh 5DEY�a� L�ȓ9�r]���S/J
b�!�	uk`��W�CEc�kc����O�BE��+�؍Ȓ,Y�8~8����T�.��a3,�V�+콐�o�[؂L��,$HA!�Q�Hb`<�ӈI�S"���8�p�����@A�ĺ.� ؄�eV�ѩ��W��ڢiR�A�8���	�b`A�j�q��i�HW0ц�E~�[��I�8X{��K�W¦}�ȓ*��)c�B�9�-���X|��ȓ+�n�2Ȉbzh��B��pՆȓk>tC��s�p�be��tht�ȓ|�бuI����Jf��0c�Ň�|1duC��j9.����W��ȓ&"X��Vj�n^Z��@�G�B��T��F-&��"h�N���)1�
�8���ȓk�l��7�U?P&�8H�^=F�Y��&d&����FX�}Qk6T
�C�I�V���/j�97��24��C䉸b
q�@���G��B Á�)LB�I�.'6�Pc�m��a��O�%C�	!��\iwl�O��B�+||C�I'=~�鳭Θu�E��~�B�	M;U�A7&}X�:F�H�@xC�I1d�.pӱ
G'%�*���%9�4C����4���B>1k�MtB�	g��qk�oC	�(=˔j�@1\B��X�J���ցe!�͢*'�<B�)� V��q�%�8x�(+i!ذa��']��W?����럩*}��b�i��_�C䉄`� p�3#�":�h�������d3��Y
6p�3�C�-2���*�!�d�	W�`ܲ @Ϻ\�� j$o!���)� �j7E�]պM�T��|�!�7=׌�+��Q�N�8��ƀ�z�!�Wh�xK �<w�F41`��6!�$�|��;����EJ5��!�!��9.nr����?Y��Y�C�
�!�đ�=�����ľg�x�!	��X|!�	�r�:���I����{v( c�!�$L3;�%Y��Y5+��X���=�!�
{7څs��P�?������5NT�����	�c��Ԡ!S�$��I�P��<��B�IA��J�D�Y��E�F<4�C�ɽ����>8F�E��FG�}&ܣ=�ç9�̠�w�%V���##�	U���H�>$��ʍ�<��PO�	&��_�сH�_��P�	�x���QP�Pp��R���32l�W�0D�\c���g#�u�/�{�8L���>�'Z�O�O�剤D骱�v�� 24�]�Y��B䉣���ۄ���[�
L��\� b�B��1|Ǽh"�a�?���2��D��.B�0���j�Ǉ�c���[���9v[�B�ɥyՐ�cQB�J���Q�C��rB��b�pK��w��v	�&IlxC䉡�H��eˑ>)��l� @]Vv:C�I�V=R����ؐx�z���$+�@B�ɒ^hl���f�8Q �W��&B�ɪ
1���'�@��j�hǆ�6B�	)$��T@����Ъ�m�h�"Or,�5�/�F �t������"O``D���AB�$�C'�<���R"Or��#N��2�;F 0j�Z-�"O�A���.�R��RN<�*4"O%)�K֤������X�'N�S�"Od��U��7���:�ፃ>�����"OJ}!�)F�����[~p��V"Ot�J8��P@uJ? g܁�p�'nPy�<��"�0|x�lG(ɝk����у�A�<����]KB5�b�Vs�N��� B}����>��`��bl6��S�Ε4���;���o�<��FDsK^���ݘ0ޤ0C��Wf�<i$�K���v�	jS��#\m�<qv�	�	y���w�ƛ!Cz�S��p�<i� B�S]��uL��-��3���p�<Q���?{���Ded`;��h�<�Td@�jl�mC򂎘� �����O�<��;@��D���Γ(�(�z4N`�<s�Cz��
��ؕG ��!�D�$"��8���;C$]��G�e�!���R�E�d�S�3> PuOO3�!�d9��훢n�z72�ӱ-�_!�
g�R����]_0����f�!0�!��#H�x*�N�%�d#�]�x!�$��O��KŎQ/������x>!�D�G�n�k�!�A�)Ƒ�'=!�d��0�p�% �t"@�1ꑦ,!��=�,�U@:P�ԧE!��=}��t��'�p�H֏�I�!�d\g;�e`��4]��݉�W~�!��{2�9���|� (�� 8{�bY��S�? ���5J�>a�$֯V+"�\��p"OP�G-:	P[�#O8Q����&"O��ᚈ(9F�ҧc[^�(��"O���b} H������"O0��	��tO�r�N" i:�C�"OH�K5 	>y&���D6aN�u�"O� ���2+��
E�G�UG^��1"Od�+b	�<UЖiz�gL�50X�rF"O��ӳ�#@h֥P$Y.�hs&"OlO�<���	�%�;z`�I�"OBh���)8�� �JRR��+�"O�r堐��lD���K@��"O��C�\�6�#`�".3E��"O�<��E�Ip<�SDȬm%��""O*9JG��m̈�C�H�}��&"O�-@��[9�it�ʾz	�uQ�"O�I��M̥l��E�g��,� �P"O`��i�1O��#�l#ZѸ��"O*�pjT1pd���d�~���7"O�]�S�6rR�٩U�K��T:�"O*ᒏ��"ulċt�
u`��P"O��o;`��"ǩWx��"O8)��K�b�J��J�(m��!�"Or������z�*�Fi6t�"O�mZ�!˻_=�-+��	c�(�JA"OLc�(�F���SF��% vt@Ye"O�I����A��8AM%B[�� "O��p���"�6��
��\����&"O�\y6��z�6P�P�>P�pT�"OB,�҇
0hI�Uc؀k�t�H"O0Pb��_�ԼRġ��r�BL�3"O�P�@.ڳA��G�M3��A�""O�AAă��L`Bo%	�T8 r"OPВ$ټ&̶d�3��.�R��p"O����l$@Ƞ�^F��H#�"O����ֿa�P��"X7LܼHR"O��c�ުM�2������~�N�0�"O�����ؼi� ���C��F�D%�g"O��a̩X���8�BE6�h3p"O�8�A���%�0��aD��0��q"O����8p�\ �̟7N�yT`7D���D��:�����&$��w�6D��`�.����K�?4^<�
2D�иGf��E��D����a!B�.D�4����
�2(kYF	(=���-D���viH0�<!ѐ�L��Z��N+D�@�*Еzt@�J9�LX2�)D���*H'cЬx#4�C/(B,�E�$D����'̺
v�� �j������C"D�8��ͨvz�
č�* ��i�h5D����?,<&���9#��!@q3D����×,f�p�y�F���	#D����[�L<AH$�@%�!D� �AcH�*�(hˇiĀ:�����:D�TR3'[�"_���T��
s(�	�$D�l��	�/c@�:�B�~a�Y�&D�ؙA��1�p��� p�]�E�!D�PR�+��D��X��=Xth١)?D��:��Ʃa!���%`�S`����=D����ݺ+�q��cB�j!�5D�����h�M�BC��\0�td4D�|(���0c@)���lOȡ�l0D��D��<o�T�Õ�[���A+D�<�t��&\\��Q�9$��d�&D�� ����E�x���;�Aڰ����c"Oݳ���"-YF �$!�&
�l(�"Ohpٓ�7��J%EQ���A3"O�<0��L?,њ4#��S%Ww���"OF����:%�,EzCkׁm� a�u"Or]�A_�Y���+��2i����"O���#-�0B���"#��8V���C"O*����W��D3�٠2h��&"O�%�v�:p���Q�+�]�y�"O0!��#�*Kt ��Y��:p�e"O�٢b͑lc��yw

~��0�V"ON@sG�� X�
W��#�Vdc�"O�)Y"FҰ�;�L�T݄���"O꠲���9pf��똤��XH�"OV9�aţKKF�!A�	���	��"O��a���L�rD�'X�jq�"O���3�.`u�EKăE�x�|A�"O�zv#pg`%80� ����c"O��*��X�"+�=�F&����"Op��6D�Z2r�9���8�½�V"O<P���0bĦ!3�'�>y�"O��p�;z�\{R`�r�R�e"O��+5/�$^�U�g��9-p#a*O���
�W:�@�%�,͎͚�'���ڡ(��F��P�6.ԑG;D���'����r�i��X��lS=DpZ�'���YD
�l�&8��Ǹ7f0<�
�'xĨPWFC,)�I��	6*�*�#
�'d��Æ�pH�ׇ[>$��� �'U���e���p6��H����'���b�̍|��𢦄�h�<�'S�MS���+I��T�F-f����'�z�����uw�ܨ��\d!K�'��!1"Iք_�@!�#e��Y�p�2�' !�3�1�T�COƆ R�q�'�n��t�F#|!�Xbf$G6t<�8��'�<!��Wd�:r�`ݩ����'��8�A��#�ʩq ʃ�u�&qY�'���Y#ā0.�������X�$I9�'�6$0���6~�H�*bвKF��'�@p0��O2�e���8:dŃ�'�L�@��s�6tAh--�bT��'�l� e� �d��`��?��'�Єh�A%R�I0�k��ȕ��'o)���,jE`K������(�'V*���S}W��y�EW'|P��'I>LA)K� b ����ǻo�\!��'Sd�q�_#S����A�7�����'�}��˕�j�m\�D	�	�4"O�2E�*�����R�F�#"O�t�PĂFB>�)WJ�%Aլd��"O��A�_�T��I�#9ú��q"O@�����c'x��ŋZ�`�"O긩u�K�A"j0j@mյo38�"Oj�:�$�0h�Ԫa%�72 �[�"O$��Lۿ1�H Q��m���"O6=�Ũ+b�X�[&��4 �Ѓ�"O�h�J�� @�0an�E�eI�"OB�����]���I4G�U���"O�=!7��*e
(�&%hJ��1�"Ol�I6�ɩc�Le ��>o?�8��"O@�d&w6�2u/��Rݼ{2"O��Gi��jB�R�G�!h�t���"OBi�"HB�]|�D�fԳ}� ��"O� �1`0߮/�X�{�R0y�&A�!"OB��E�]�-G�[6�E}����"O@Lb�)ќ@Y.���[�b�@�"O�(�%�&IT�u��Y��� "OV�T"�!(�����d�PlÁ"O0�r��%� �4![�k�J��"O*48TⓄ\�flJ'���f4ČIt"O�
gkN4:Z�7��B���"O�\��'^�RG �w	̥���{#"O*�AYX�R�K��kh����ݲgY!�N$0�����g:�
��HLM!���*�J(J��U�m��3ӥ��oK!�F�.c 8;pFQh5�gE�J�!�DN���*`��t��A�s@�Zv!�Ā�2V|3�BL�{��y��M\�W`!�Dս%��O��6#E&T/aT!��=w�Ȁu�V  �f��U��>@!��[���#��%a���@�'qO!���A߰Trҏ�f��=����2G!�K�wa��Ӥ�J~���
� C'!�D�2��@��R�e^N�{��l�!�0E֞P�v��Q�(�Pb.�!�=2����M��S�;��_�e�!��i|d�b�ȭ>,H�r��M�!��Q�z��]�'�d=��0ņ�	\!�$ɓdv	P�-N�d�~x�$ĳ!�ĉ)@XB��7�Z�<������Yw�!�$�7!�L���@�[��!م9#{!�ˆ
�h@�"~�r��WC�3w!�D��]�6��hϦ<��+�C]!򤞜yx��`�G�%��8�+� %!���(Z���q ��P}�]���i!� x���Ht�d¥��	�O�!�D�:�x�:uă&]G����H0>�!�#	4�H0�E4!-h�S�xS!�d�4��C��R �h��܎G!�$�u��D��X�__�س�E6!џ(G�$�>\n�iPF��)�Tb2,
���d(�OR����\�L3L)B��S�29<TZ�"O���� �d;��w/A!r���e"O�h�3�ƥ\�6I��+F�y���r"O��ȱ�4ց��kD.s�����ݟxD�l4��|˕��'K�iۢÚ��y��Ň*襃����q3�^�yr/�3gIRY��-�/�x�h"��yb�B�Z\�Ѩ %�"�Z%ѡ�Ϥ�y�H�n� H�(M���!d���ybA.~��@xEG���]! MU��y�D����c' �[]��
j>��O�"~�f�?hI4	�.�'��\I5b�^�<i��C&-P�sJW5'c��NQ�<�B�\)%��M�"b�8B0���O�L�<���/[
^P S��)o���B@�s�{�h��d̜a��+��З�.08.4D�(��N��Kp����H�8i8U�?D��j�G.9�x���?j�H�I��8D�Py��
�.����
9P8H�e1D��I�YRᘑ�ԮhJ���ë1D�L���P>2�t����_2;7r���/D�\rpL�2�xK��R[�R|� )�O(˓��<q�'�tlY�aG�)H@�vJ9��а�'�V<��! ��%�f"�-�D���'O�M���a�8���� �$�	�'�� �f�A>H!6)���gb�U����?�
� ���b����H;d�73���t�'�!��8Z
,ۖ�A�!�4hwk!!��6k&���]� ��W��:��	]��\��*pq�9�k�g}>�#�L8D���3�S�m׮a ��؇2�:ɓ@`4D�$����~mL�)�,I50�1F�>D�l��$�b�R�I+Q\��H��&���O��$� ��H�.Ày�����B�F���O���2�O֡b�L��M+0-�иhc��w"O��X5*K�O{ �[�	;VVX��"O�Bf��T��P��wcڈ� k.D���B�Q�˚����t�>D�8�q�V/?u����X�j��iR
;D�T��j�մ��W��
5Ǟ���9��4�O��`�&_I?��jb�@�u�0Y����d��	f�ޗ|F<�CcmM�%��[�b1D���g)W'(%��捪U����2&.�d�OH˓��S�ɔ�f�θ"ԉ-sD��)"�q!���`\j�1�)�s7�`
c]�Qb!��:�H��È�U5�p!S /!�J�Psq*X�`�4ۀ�àG�����I�|̄m�&Ř.�(2�ТZB��;l���`�����p�#�"�j�*B䉡p��s6E4K��i��Ɩ&���=9ç_s*�D��:14 �U���+�� ��L�TQ�s��V�(��`̇s`��ȓ���Ei�~�� )���6��ȓ��[")�|���м:x-��n�R���?�Ó$v4��@��:l4K�Oȫ\�p��?f���O]��08�ڥw�N��S��B�/�O��9�5�A	9�`���o���	��;'��QևMUf$��_�t����:%�%	7l�\y����@�e�I89�r����~uN��D��M�$�G�
y(���Lb�%�Is����&��8,�Ry�m���T��%D��J� 	+u�.�ؒi��u@xDqr�5D�0��]ڼ�nN�F�>�H7"�OD��<9�����	\�l��_�H0��$+
�B�I�p�t@�cK�W�С�eߓG�C䉍谢4��;V��90c��*Lu��?9����$ �x�*A�z�tĳb	/E���)�' �z�ǃ�-.ZD������<� q��'�=9�P�ue���^9�$ak�'m� �62�l�XU�,���O�����1��DU�&|�� ǯ] b@8�D���!�҉��1�g����Z��{!�d���y��ܮ2B�Cժ��Q�!��'��5 �XA �F�zM!��҅t��QᶂL"$��RG�'�!�� �'�Ru�"iW�~(�葧P�!��P��A���޶H0����'"|"�d&�g?9&J1ey���"փ������]�<I���$�ࠁ�	tN΅�4�D�<���C�8�ѣ�fD�2m�!CD~�<��Ok!2�`䄎|$�Fa�p�<Q��&�@� �&�{.H�w��U�<Q��H��6�rr�a�X�{ebXy�<�����E��|膉^?I*@�{�E@L�<QNQG�4x��ȸ||�T��r�<�qE�tlB��t�*+�����Ke�<��4b�Dqr�C{��}ȲΌc�<9e�0J�hMR��B�f���04�S`�<�ïG!a8�D���]�)в��6�I^�<� j���Dݖ�`�����;2D�������G��N�9pZ�{t�ǼT���{Q��
�y¦کP������^5F�L�	�Gg�y��R/�D�C�EE�)3�/X��y�@S�-��e��@�-)6�%!�;�yB$�)�в @��EX���y�Kޗ����%iT;RA�0"&�y2KEO��)�פ�%y�.q�7����>�*O��Aw�P�Y�,4���޶u��I�3+$D�|Ȓe6�UWcX2s�4x1�dɡ�y�+�S�4`תɔr���k %�4�y�$A�,��j�ꔪ�p|�G*�2�yBE�
I��d	��٣��
�hO������Q;��e	�jl�RS-�f��y��I�K6T��5X�D��U��jձ�h�$D{J?%  �D�y,h̓��]�k��8��3D��CdKP�yO� {�F@�~R9ŀ1D��qЬ�3!d�V'	��Dȉ' 1D� ��jF�C,���%Fi��$���4D�d��dE+${B�q!C�sx\,	��?��7�O�$�V� A����J@�(�X���'�1OV�0��X?)̢� t G&��sp"O�4k�@�t�%Π@�&�³"O2�㖭�7Ed] �"U$m�� "O&�&��5(w�� ��c� ��"OFՀgC2_���� �:aZ���"OD�@Q�&NV
��/�(*��4�'��Oh��Ұi��y&`�P�N�!Ѡ֛?F�}b����'�6.��ŇG��Ӓ�&��#�Sܧ%vQ"�n�(6��0��"6�V��T��9CQk�1l�.ib#�Wb�ꅅȓ]Z\��2Më1���[+pŇ�(�@���H�C�N�Q�!K�-�xU�ȓ�`e�t�Ȼ<�J�� ��#v���ȓ6���$$Ǫ$����EMW}�(��A�@���'�L{lD�BdݕF��ȓTv��Q-'/��,�'oުh����ȓj��NF,��"m�(�,��ȓ)�������;>۰c"�!G��ȓ�H��@�&����I� &���ȓn�dҤ���9����ċ�*PH�ȓ<&4����K�HieE[6&����zs԰b }\]�F2�\	��6�����ϫ ��txW���e���F{R�O�l�>p�0���4��y3�[e�<I��s������&�(p�
LV�<�R��>���b揞1�PQ2t�T�<��9 8~I��eT�>O|�k�"�i�<a��G<N�|��/�6(
p����<9'�C3Th���Aj��N�a�Ew�<1R�A�����sdh`���Nt�<9@-��A���$̪a��鰐��v�<�!d��9w �B�T3�~����Mo�<)��"p�J$ ��6Ze��b��U�<�ab͏R���3�_�d���:�W�<a��6�@�E�N�Mq�鰳c�V�<Q��
�81�]%?��|�F/IU�<��A�p���B3B@�OZ&���LU�<�Ŋ�>=zXJ�X8'f0aAG@�x�<��ǚ,�u@���2n�%��w�<ɥǘ%>+��*�ک"0�p�r�<1&��$�2��$f#.�@�%Tk��L�<a���>L>�!_�cG}P"�4T���GJ �X��-���-6��<�4�.D�� �=P͚)#��4Ð�k�"OzY8��S2'�l����OM��bu"O @&��J�V�I�;О�QG"O$�J"G��p��%���s"Oi�q �7+��7O�Ay���"Oz͚T�D�e�G��Nt���"ON$�D23k�K�Ύ}nB�"O�Y��	�1m�(�`��΂uS���"O�9�q!��0�phĎAu�Ę�"O��'�C)���!�mC���,� "OL$ 4���5yÍ J�dA'"OL��R���^%����j��8S�"O.8��H8�DX�����a�"O�0�c�ύ钀����(�FG"Op��%����#7�n�D"O�1׌Y�Ox	Z����|y��"O��0W�\�z�F!�A�=���g"O�����ܚf��-J���[�"OF�9+ݭy�B�gL�	U��8�T"O�	@�[�|<��*��1���"O�������+Y��cWUy(X#"O�4"�\�4�65����[Y0$3e�'�ў"~�IQJlT���/�	n��F�y2��]<
X�WKN1��5w�Ź�y��	��,�H�JH�u��ac�$�yM�$s:"�		J3g�&��a��#�y�gkG�E�5j
�`��i94aR,�y�d�6`n�8��_�Q�h9#�@��y2�����K$e	-F��5)c�]��?y���4�P����0�d0� `Q%��-�ȓ
0�P�H�a���郃�G'���x�h�yЪέ>����Q+\�T��U�L8�$D@�v.8�+vCϽd����ȓ..�yz�.L�{���K0 ĻV�
�ȓB%�����ET�1��bD
|(e�ȓ:������#KH8A��uX�	@y��'���S�<1G!��^�}buo��Y5v�"��Ur�<��ےr�j��/эhBQ�F�u�<�TA�$A�|Y��2����L�<��dC�Рd3�Z�c��Zӂ�T�<�P#�G�08)�FV4 9v�8�H�R�< %D0$�l��gAI���]yw��g�<Q"lT�9ڂ��4쀩�*|�ߟ|��ԟl�?E�������H{A&U�I7�}��Cѧ��4�Ob�(��_���٣��"��y�)��wEN)6I�D>��ɑ%��y�nL/F�ÍD�C�nh�M����D�OP��0|Ԩ�uR���F�����R�%[�<A�		)Z�J%D�^kv��@Ka�<�]-��	�g�L�Ïxg�	D���JT��9U��|!���'^��q�rJ-D����S����i�3s-n��$�,D�tV�S�k�z�Y�ϟ�g�4�� �5D�d���g~d��*�>F�����4T� Z&̖Q*��Vo	&���$"O�%A �R���!8D��	���"Ol�@V́*��&�Ho�JÙ|"�'&��E�֩?؂�Z�OQ1oC^�a�'�l�S�T����a�_�^?�1�'^n!�«I��	�)�x���OpX�(P�g���V�'?��j��|�|2�I�l����v��<Hn1�4m�9pk:5��0
麰!Ҟk��0@�J5ry�<�ȓ~�գ1�H,.}�Ƨ˳,t�'82^�HE{�π 䰻��I�pU��X��͆wc\$�"OpLYqk'/��p����bXRR"O��3��޳^�ԥ �̃��~)8��'��	<<J/^~c�+e
�K�T�D2��|��$�p�dH���T�������@�!�ưƴ�r�E���@؁$�y2�䕳5E��x�gS�=�lh���y�6ʓ����O��$�d?�` t�6�4m� hr�Ub{�<�`���� ��!�9B�t��0@_�<�pix�)���d<9Kq�J�j!�ć&U�n�"7��Z6��R�^�K!�D[:ߠ̢FoFL*0m�NȮ|I!��ɢ�y���9��vm��G�!��8���4f��oMJ���&��'ў�>-Yg���|S&��k�����1D��2�b4ot�9��"�<Չ֤:D� ���>�)7�W2��k��8D��q͒�S�"%����>J^΀��3��Z����g׼G��uX��	.�fQ;��7D���AEM�3@s� 4�J�rv#D���d#�fDQ��_�V��T;�%=D�T#A
�+B�t�a�	3pě�&/D��jF
��DH��]0�$��i)D�X�rIM40o�h&$�+|��}�)D�<4gs0�䈦c�$1�}z�M'D�����ϙ0\`����b���p0D�����ιl���˶�C�bJ}b�#D�$�uK��/���1U"��4B��G�R��ҎZ�%����8d�lB�1E�$ ��gsʅC���5�(C�.o⠨q�B�|���`w
�(4�B䉧!�|���B^;J��hC�"$��B�ɥ@"�S����0�R\�P�Ф/zB�I�yJ�00aȞ�vt��K�PʰC�	�
��S�H �g@�|�lU� ��C�Ɉ�:Ձ� _�dm8�#�v�C�I�a'��9��Q�/�H)��ιC*TC䉰"*���	^�.�t��2 C��B�ɮx	�� ����l�S�È9>����O����O��D�|R��ܘ'���#�W�!ˮl�Ejи!�t�h�'<�)I+Q�~�Ib(��T���'?~�i�JC>������.1�
�'^8ؒ�B�|��ؚ"	�N�N�	�'�h#���DRu�R��B�pdp�'�xX�d@660��>�B\��'�(�1�lY�R�̤���G6Kd40P���?Q���?	���	�O\b�|�7�׶[T��P5_�ᒅ�-D�<�O�=B��`��
�E<���bo+D���F��%X� ���މ�Ip��*D���aZ���8A���'=�8X[uD&D����ƞ=$qP[1PH��H��yr�F>xb+S�����f��y�a�{c����0�����?���?1���?9*���� �ɿ JT��s�Q92ݒ�:�?erB��)䕂��Ɲkj(����TB�Iz�dxC��#l4�E@5cG�C䉒�xJ����?�b�ˁ��Z��C䉜[`��Ӈ��-Y�N��b#C�C��g���sW����xb��dC��3G�����@�Z��P�1�5M��B�I�M�8�jg��T�.��3��#�6C䉎U_J��`Y�`�!�U5JL�B�I�hǾ��5o�$�dz�E�2NzC�ɿX�U3�G�0����F�Mg�B�)� |)�����#B��(���"O�����Y���c�5.��A2"OPL
0��4=��"�)u�@�"OT�! A�<�D��~�Ci��yB"B�8 �V�Y��¨����y��	�� ��Rl���B-�y��LUy��{���g��b��y�gYz������~ "�����yf�-e�@�����)̍;�yb�D�y76h�a&�M�&�A�Б���0>a���SSh�{�aԑd�*�3%H�<a4!QmF$a���1n�s憗|�<��FŴWS����*s���Ũ�M�<9�.�"^�b���)qJ�����`�<�'[0!=��j��R�u��P�p�<y��M�L�t��vL_��4h:��l�<��]�k�x8B.�*u"D�hBh�<YV��y4�x��33���_�<�dPepU:�g�hŠd`կ�[�'.?-��\!��0�@��Fs�B�	bx���3ڵ^�F	AF�a��B�I�F��e�E`ƫlP}#hB�vB�	}#D)����g-N���LAxdB�ɤY��ej#Ɂ�)C*u1��_�4B�I� ��#��DN~�24��J�LB�I�Vú��#� e��=Q�B��Җ�kn߫%�G)�~�B�*��`fw�\�����B�	��xU(�,G�����ؠ `�B�I�T=>��v�L2E#D ђ�dK�B�	�@1đ�T�i&��Z1�H��B�I@
��A�F�b�%Y��s�VB�In��@a�=|���)�+�3(B��Q�J|Z0!@"�����Q��C�I9z-8��@B�,zy���(1�C�	�YE�����O�B����d����C�I$��5A#�@�HXt��/k�C�ɒEhL�b�W�$;"��$cA�MiRC�Ɂ{6V$�5�('%�-��QAC�I9^���{d䞤��q0�+H�	��B䉖AmIi �î'e��S"ى$J�B�Ɍw,"����-�nl N��`۔�4���$#������ǋXb�Ra�mu.B�ɌUS����Ѓ+����#J�B�I�T��)�������������$'�S�O|���]�LҒ��b
R;{���t"Ov�@/C����C��#�NP�f"O�S�O��Q@"-B�˂�.�8x�"O6���4A�]�-��p����"O�9� �+U@���k#]X�a�"Od��7�ڂ%AV���*��Y���[w"ONyȦ��",K�H#<�(W"O���hX�"OܕqDh몤I�"O�4�Bo�!<@�DǍ�n`�"O\ۗ#�?@�����M7�ܨ["OFɛ�bO�\u�X p�]-c~Ȩc0"O���b�Ź}.luE�Ow�*�"Oz �E
@�F0�⣋8H���"O���f��/)w6MBw�ǘL�\�V���<y��I�=u��)� ��//z-
'c$
{�Ofk�	!&-�I�� ݴ�ux�"ON�U�޺n�Z@� /��z���"O��5��CT��ۏr ��d"Ox�i�����R���R�Ng6 K�"O� ֠0�NLt��(��MnD|-r�"O\�"D)F�G-f��$�U�gs�����|��'="�|�|�#��G�(�0�ƽB�l��t�M�yp!����qz��/����m�"j!��7+����EaF"N(ށ(b-��!��AvNt���XJ�
E�%.ͩ5�!򄀌v���I�DV)K��ԧ��.#!��"b���kuo�C�܅K5!�K�~�*�q@�Y��)�3�_)�O��D,O�K1$� @J�gGO1O(	i�"O\Њ��57rS���Z���"O��P����S-����BQ�m���Y5"Oʔ�P����BDh�jQ0Jڶ�`�"O���ݾ?�(%[����k���Q�"Oz�rA�ʕ#A��������6"O8)!Tgm���6,��}�ŗ|2�|�R�t�|�#k��Vā��
P윒T �]�<I6��),��uH-/����bGZ�<�!�53h�jp��4iLd���(A�<���k�h�s�ԥ.=��A�<�G�П|��5��gȟ5֔x��e�<	F���0��g.����)@C�d�<���I�6����@�(��Ѐ�j�	{���	�O�zfK�Z�H�C�J#Oܠ����4D�(�2�]��V��2�$I�aa��y%�\0@BE+��)��(K$�y2���z��
��]���Y�u�F��y�"���ؓ�(ÑO��͠$H%�y�]�\m!i�Q�"��+�1�y�+$Bj�*�^%�1�F�y�m	+6.� S�Z�4�"������y2�On����".X��*UN�<�y��¤qK��`@���y���<%�̪1d�wl,A���yb#]�J��bb�	Ԧ�@$��$�y�W�WK��"��՛2��pbk�=�y�� ���Å/K�]^����O��y��1M� �fB�d��x���yr`#~��dт�ށE�p�dI��yB��,<��i�O����?�y�v��E�?G�|ذ�����y��[=$�:�9B���}����+�yr��>@읓SC5q�Չ%ʌ��ym�#��ˡ�nBh�{E��yW JQf�{���-U�(iSe����ybf
�j��0V�a�P�Q�fG!�ybIA�|��ȑ�Q�,����]��y.�1%@�AS�ӥu�ąxb��y�Zq�t��IV�p��(1%\�y"d��m��(�FѵjJ�e��ʓ�hO���i�wi����2�H(�5CܢuW!�d6[��r�+	�*�)��1)!�d �m�j@z��i��pJw
ݚ$�!�䚗G�ICʌ�D�K@�A�!�D9iJ�p6o*[���`a�,!�$D�(����u��(a�	>�!�����4�*����c�Iߏ/�!�$���g�?l�zǢ��*��O���r,��g�"�ʂ���n$ ĪQ�&D�,2qG6*$ `d�*k�6졂`1D��� ��d;֌aQ��c�N��0D��Y��Y'nD��A�B�=2�.D�����C�L @���mz����H'D�҆�ڂi�P���('c8��F@2����� 0�h7�L 3���	".��{�*x�U"O ,+�	O�Zo���c�Y�(�z�J�"O�1��I�J�s��#�u"v"O����Q
SF�����I:0�,R�"O<u�dGB"]�:ݘ�f�)�h-1$"O������lh�%�J�� �0"O	�ؖ=_�>Ͳ��5��r�"O��H�-�
h�A������;f"O��{�
J�@U�Y�u�1S����"O��$��%%p�;k_0�❐�"O��Ϟ�7^ �"��į;��X�"O\1A�?� r� !�\c�"OBi�ѫ��22���&Z�q"O�@��&	����+�x�d�[V"O`����ǸN�`��3�A=�<�g"O�iw�\3c6 uk��
�h��l:�_��F{�򩚟4�(�F˃�*FE�@�X1;�!�D��3����E=y�&u��㔯/�!� U<J�b��G�?��IPPb��4O!��ld�c�Hȥ5����o�B�!�D��N���	&,�(����-�� �!������C��)z*!��K�-'a�Ip��x��Ɣ'u� (	q�~n� ��'D�P��	
�~�a@�̙tJ��c �)D��٤#�9?n�R�K-�v�`"2D��x�I���$D�RM�� *2��B�=D����*�7�P�Svp�9wD=D�0�U���.��F��?`}N�H�	=D�4�7��/vNȘshO',0y��'�b���T���ǭN�lX@AM
��O���� ZHȈabi�h�����!�X,C�VdR��toXQ�9\�!�A{��LR(	�bH�`6��U�!����&hѶ#�nĤe>�!�䓅�,Y�%�k$=���$	!��-q�xu�L)h��IX3�G!j�"�)�'w 2�k���LWj%"4��10Q��'�~����1�mht/H�V�r�j�'��y�CѾ;�����N�!C���d�?I����&�ǮM$�8R�H��W�!��U�A�J,���h�4�!��Y�%W��P1��:5�(��&�ɨ�!�
?�D4��ÀwԢ���K��$}!�W���85e?_��`BA��g!�ܻ$p�!��Mº��
Y!�d2�)bEa��_�8���N^Lh!�$�/vT�$Ó}=��C��d[!�Ē�/���9d�ȧQ�b,7,�F!�ʿ*B����ݯ˾IcTM	4!��L�+Bn�8%�(�&0�왶G!�d�|{�0�J�]�J'!��SS!�Ҁ< �e��'?�u�  	�s�!�d��Cx`�r�L�~$��xuH�B�!��*4 �٤�I�<:Z!���b!��Q�v^̘�gEP�aS�a4V�u�!�dR>�:)��V�W4Li�!�E�!���)[��S�N #�*��/�ў�Er*�)h�tá�ڍn4����i(�ў���I�2��D(�DؕM0 တ-"�C�I�s!$I�'�1fF�eb3k�5��C�	�(��U�%��`V.�)$B�B��!) �g�XV�`�y�fB�I�-`R��R�H>MD��
2\edB�ɡ��(c����|}2!��
6���'�	m��ߟ��O�� ��Sc�Ss���W���~hH�d7LO����Z=%"�p�ю�2
���+�"OҰ�OΊ��s�#]eH�#�"O��  ��s� \;��ٺ	H@	��"Oa�V�h*EHR��6B�8�A"OA�Fㇰ%�.U@�(W�`��"O��[D��4#��ZA��Ne�$ۀV�|�I�l�'�ўЁ����bb��m��i��[��E�yb.H�xz�T�,L2���%���y�`��w쀱�)Ђ� �B��y�(]��m��kɏg^�9����yB+�7���P��e��� �I�y�W2~���X�o�[�����yC�;���eG�Ya�L���@	�y��1,�e��(4<�����ԙ�y"#�%
쨬؃	Y�
��� �È�yr�_ e"D0x��ͯ.,mp�ܳ�y���C����5'��&�&�y"%S= ��P[ �ؓlu�t�g�yr�V�[x��i�h��Z�Ŋ��y�䑧.Gl��Ն�5g���FG˾�yB0
y3��Z.X�
9F�y"��D�Ń%͓�O�8�#F�E��y"�% �bR�U�XN��E ��y�g
k�v���N��z�aF!ƶ�y��A5lú�����E&p���E8�y�o2���s�g�9yx�B�bN;�y��J�2�[�	���kӀװ�yBOW�HO�0�t$T#lX�����@�y��҄tCޥQ�Ĥ�vi����<�y�*��D�Y�ga�%�bd�%H:�yR��3\����'��`e�%�!�ݘ�y���V�yt�[�.b��|c�'U�		��Љ*��Es0j@�=�ڵ��'�8�D��[B�
� X���Z�'��P���:�h��W̜�
 ��:�'*b�K`�݌/������}�I �',��I0NmН�"���u�����'G�������u�+��p�)�'�~|���A�4c����cŲ	��'ܾ��0���dm�\l����'<Иe��\���ħD�^�ٙ	�'ٴPҲ�F�h9�	���.E�X��'�T�a낉|�z5��ŏ�=��H�'b���"�32O��a3�K84jԸ�'�D�s�A�]E&� v��.�L��
�'�.)��'�'�D�`��/+p��'Td���e</
8 H�l�B@���ȓ2D�xT>'"�<��������ȓѸm:"�P!/-�( ���Z����v�.\0-w��%'�'�Z�ȓ%[����U8���0F�tP����1j`��!�|�NP���ԧe�d�ȓh��E�5�V@u��s��-��RR�M�2-�x��|𲠐.H���y�`+(�p��� S��ͅȓ9���ue:ghV8c5�F�v�0���q�$8�Ug��M�[�a݊�$�ȓs������6c��Jj�=c0
!�ȓ��Qk�#T�z�bG�_�%��@�ȓB�(�`��X�N!V1"��G41N)��aK@U�� "H *]�����'D�\���dS\m��N�G��@�68D��&��$h)Rᙐ`@3�2#��6D�� ����mŴs$���Z4_��`�"O���aI�13f�;��Y����ʦ"O�ٻ��
k�ڵٷ*�0)J���"Od4�\(J��R�ˍ'?^`�V"O|���LP��|%C�2M���8�"O@aj��T8�}h�K�`M��"O�mz`�X��j����$7 ����"O��áb��:�[u�D(d
�K�"O����\���Q�G�.]߈\{�"OL�9b&�%:H�Qp���k�4�`Q"OXe����m��2ͅF��H	�"O|iҢ��sJ��P���q�ܭc"OV�JR��{*�ii�	�+d�����"O���sJC��N8�vhT��ۡ"O����� �1YF��C)���L˳"O⥺siT�G2�9��Y���U"O��BC��f�JlҶ��'C�$�D"O�����[|lys��*���&"OU��	Q':��r$� �����"OB�����#�*�� d�%�H� �"O��hE��47]�ĩ�ɆE�qE"O�l2��gq�Mb�L�b"^���"O^���
��q}��R�)k��9G"O8y�_�`�9���J!+X�Uu*O`��NތqX�1�ƇK:J(���'Dby���m�r�B�HĎ0$����'��x)�!U��Ѭ�%6(��'E8��G���(���$����Q��'�L-pDKZ��[Azj��k�'�������:�as��p�0k�'7|q��q$6M�ǯ�dJ�z�'.�L�C/Y�+#� +��� k�&��	�'���z�K�$�@�0�)ػg�f�`	�'��l@A#)���4c "\��'�d�� ��1Xolģ�F�W�64��'��(�a�"d��Egk�#:�Lh�'�
�X�&��i[��֥':f����'��� �R6wP��V�K�+��'9|���®��q+�#(	<x��'��A	G%�޸�y K�m��	�'�V4�N����[�+Or���	�'D��$N�;a9Ԭ�@$����b	�'��x�O�$[4E
�K�a�P 	�'Dr�i��"{l��������'��SтG�f���UV�*�p�'�]����� {���>�z�Q�'��`0��[!��}�Ňӟ1[Ԅ0�'��$��	�}�Pѳ���0G�Q��'�>�C`kK�.��S�O)��l 
�'F0���R�p��s���F ��	�'�i3���y���(�HD��p���'$���.��"�b��3�3:�4�r�'��M
�^�i�i��
��;.� J�'ۂ���`Y<M!Z���`�0L��	�'��a��EX/RT����s� �Z
�'���Ŭ�-?5JIp��ϸw���J
�'����bF��j�K�'H:sa�	�'T����6H�L�%+��v/��
�'��c�A�9�IB� �%6���	�'���8 �	~pL��
����Z
�'3ܠ)ѫU�F��1QC,�cth��'{:��r�J.[Vܡ��LS.f\a	�'I���Q�~�>5��F�+���
�'=>��t�ߘe�|a�2D����U���� ����iJ=�b�S�DD�N)�l��"OމaB'T"A:�Y�b��F��[�"O �t�x��-rQBφ*>� "On���C�7��Qu8{"D Ñ"O$���5 ��)��
�Cs�� "Oh8óF�6݉�B��:8h1�"O��S��N&j�3���>��d"O���%��*-�<�����Ck:|��"ONq���
�(�V}�AoT�8f&� �"OD�y����eF�I�c��#"`��"O��mҲf`X|X��O�n6���"O��4jD#'/:�t���9�8+�"O*�*d�ѧ5�`�h��I�Y����"O:�3��X
�
� �����"O��x2E��<�vI�uhބt1�� �"On9U��E6\`�S͜4V�CU"O���2��_I��Ct뎔`&�q7"O���AɝJ]���j�<L
�,w"O����H�"��xP��>*���"O�鳓JȄcޤ|2��l
�1Ӳ"O�)K��E�W �=bчL<�<�K�"Ot��ҁO�#q���U�@�jS4�r"O��i4��y/��h��">d��7"O^q�)�n��IaA��0�m��"O��!�)Ik+H����S�VW���*O�����M5j�`���+�Y��'o~Ee�)��I"}�Q��'��а`.g�F�#��j<��
�'�V@\5.�����	�@�� :
�'7`�H�d�Y�a�@�a*�d�
�'6. �c�ڧ �e�e$��\I����'d(�:1�S=y6J�&g^�`)��'���<p��K���>_�a��'�Px;@˜�gENL�Sǌ;�v@P�'�^��D_T�2A!�%/(��j�'|L1b[��z�tjR�&H��A�'/�S�O�b̔� ���)-���
�'�BQ�#Ħ;���b��J(tb�iK�'�й�e�/~�F����K�q�$3�'�~)0U�<���a�8Y�����'� �����KL��g�D�M�,�y�'���`c+ӓA��1w
ֺy����'B��S�ɬ־��V�T�r�J�A�'7r��թ�-@���ؿe>�x�'�4����O�8Й�#٤�F=�'[�鰂�;�B��n\#J�D��'�� 5
�U���S3�C4~����'h�p����B!*M0��X+@r�z�'����v��)�6QYE�'ER�Pa�'G�;���h�����#ɧ>�r���']�xx0��3.E��""ҵ!HJ��'��C9�h`[d�@��]��'&(c'!��2y�ݢC�Q��>E�'�f���铵
�������=Y�'�.W&U��0qb��|���'ET��,t`.+��7�Z�!�'4
�
h�5Q,J9�!��z��i[�'�m;�L8Y��<q��E 1B�',� J�f (4͐�Bb%��%���'�4t�b�ˏ:䡃닎,� ���'���ˏ/��$�5�m��'�y���8Z~���� 9|�r�'�$ܚ����z��Й1	{�4i��'e"X�e#GY�(��j�/$�j����� ���q�:aXJE��B-n%�g"O������@���kF�*�0:�"O���
�#
��`�l�%v�y"O�0Z�@�5��MٲꚒ	xt���"O�Yp��Ys���h$��i�"O(e�c.:��ʄ�r
Q���(D�����(93.�E�ڨx"#4D�`����9hx��/A�Z^��H�3D�`i�aQ4eY2�3�j�St���u�=D���Z�N:Ѐ.u����h=D��p�"=�
�s�K���t$zC�<D��+���ab��)�~0�c=D��	���q�h(��N7�~�8�f<D�� �b���.�h��C�Ƥ1�C�=D���rO�d��!V��V�8��c�<D��{�K2ŀ���O.��%&D�؀Qf��!S�p�a�$3��*PE(D�X�E�E]ھ*󫐞!3���@:D�P����z=0��̆+8��w(<D�� �`.ݶ�J�+��a��ks)$D�X��X�w09�֝>ڠ�N&D�,[Qj��1�J�+3��k۬�ʒ�9}�1�S��bB�Ȁ�
)KRI�j�\0��ȓ6�Q�U�
!;-l n-cH��=�6�1LO�3F^�t�d`0eV��tm�#O�l���F�:���Y�G��y� L�$4�S�'e�@8�-Ҿ2�Ҙ:�hʕ=|�-�ȓ~�$�3�F�6]'h�S�Maٜ��V����!�R��G��y�yr�i�'��{y2�NHJ��/J*9��8����<���I�@n�Y�FoӅ=G������,q5H�=Q
Ón��x��[�X�&)@�|��m$��E{���CZC�N���*r�X���
��B�	\�����鐝8/2LS��8�Zc��C�<,O��c�]m"���x\.8 6"O�zta�j�dt*OP[�L�@���'��y�lāp*��6O�U�(A�Q���=��y�KH&�~��UP J$xq�X�Cў4o�H�'�yò��*n؅r�II6	�qjv��,�S�)Ŕ�ấ"B4Jx<����=�d6�O�P@�B8�,��+A�.ڎ�"O�	u�_8O��H2�*���9O����ْX}�����C�h��G����I`̓7��V�X��?;r�Z�'t�e�Z�����&|O~��y��vH
�!���?\ܦ�˖�Ԉ�~��IY�O�Z�ٲ턊@��u�ؕUgP-�yR��Q���O.rHSʔ�J�P����F6Nݘ+O��$��l�O*#<��
�3��U�*�+z}<i�tIrX�Ll#a�7��*w�ip�0%p"5�"�λN|C䉖G���A�kڹ(�AHu�̾Iǰ���I�I���x4��.��#|�S�ʬ�I�Ưw0]ѕ`@x�<AF��3�Pљ0o�_D"	wLt�<�կ� T�q��]"	���a��l�< ��}.4zV�Ȝ7�����BR�<�#�
|����.I�tl�t��WP�<Q�W�ik��U�ԅ.���ҵ��I�<�4@�w��1��zPh�!�XB<���3O��;��0�愓5�!%�TD��N������s�Z���;cTd���H�'��@��(�
`��� �=7:laB�'����B-�PX �CRoާ!�z�	�'�� �©:����U��F���' ��jRlՖ���'�\k�u�'�Jtp��:9|���E���
X[��� Da1���i�V�i�("~Oj� �'��'�Z�K��ہ����Ɨ�r��b��hO���%X	3x�E�2'���*E�t"O��[#oQ�����&Ŧ�@s6"OT5	���X%^E���.������x��'����a� �fR�N�h�9�I<ϓE~�E&k��������F�D�3�RH!�H�]Ep\P�`L�B����R�S������� �~�A��!��5#��_�3��z����9�DIț� ��ؐV���jp�$#�S�O�=��X#Ǩ�RF�1�4<)�'�Ԥ�� Ș`�B����)r䲊��!�S��E�#�XӳE�"� E�Al���y��2t&Z���dq�a���'���2�Ol�QhB!6��B�`�*���b���!�d?>�U����]#(	5К!az2G��v�'d h�g$V�E��!��U�$�3D�D�`ab��ؚ���.�L��&�,�Iɟ\�?�|��M��@&�˩|��0*�f�R��%��Ё�̳6"�����l�옐O'�IT؞������Sv��Ќ�6�Ƒ��?�hO��`�Fl�fI��^^�B�,��G<8@�"O��.td��͋�:HI�m��W�!��>0�f�(mΕP�2ti���q�!�4,mJ�a�δ�:��(р�!�?����e�-<����V�I�!�$)t��D	� ��|�&,�1T�D�=E��'���3��,8gf٥�4Fn��
�'L^ �R`H0q�Ȍ��܁;�*t	�'#���' � �X8�E/X�\(�����$�:3NQ�)�!�f����B�d��'}ў"}�����x>z=	')�^0bbXc�<�e�خe-X=� S?�TX� ��a�<����5� 3U�S>**49�^؟8��'@��)?�̜�g�Ҝ���S�'�X�xf�\���v�4m��u���(O��Y��I�7r!h��R�z�,��-��{�$��W <�p AL �J[v�C�B��	P���O��d��A�����߾Z�=��J�0@O!�D-k�d�#A�E���! Y� �!�49��)� �;
 	�C���!�D��hR0buK�@���M�*:!��ٺd[6H �$WHA�M��-�f5!�D�b�(��ϝK!V���,�<!�䝘J��1�Q#؁�.%ax��>��OD�ɱ ɡ)�	��
5��	�ʬ>���S�&���2���|-�ȈР�9��"=��ĵ����ÃJ���T'`	�����*D�Ĉ��V29at��|�8����2?a	�y��T����&"�����.Z�9�q��M�G�
9y�Ha�
[�\1�-+�+IH�'4Q?!෨��,�ĝ��J��l:� #D�`�RΚ�RmZ����	���$`�>D��5��13JbD-&(Р�ێ�(O��'���?�s��H��q �$@>r��٣b�H�<y�\v6Y�h�W�	�5
�9����ȓ8�bS@kʻ�l	ځΞ3 [@�F��~K�X�7/��)K�Lң=��x�,� ���[+t% ��z�(`�'��	G�)ʧI�yF�ɞ�Xe������p@ ���O&���@˧M_�����L�Y��T�t�|"^����/l�m�pl��l8�80�BY")N�I[���Ȇ/N�7~ �@vmZ�,���8�A��y��WF?�Ĭ&��b�'B�xE-Ý���r2�׈O����C�)� ���#D?+����a
�C=��]�4���/
h��馮��~̀��&�f�C��\,�g/��)3f�� M�( ��б�ET���Y��0͒C��/�T8�dn D� �"cyb���X����ɥB=D�țSF��r���{�O�:�3��;��;Q�b>Y�+%UP� k�
Ң=�L � �:�OD�I�<���R�+������Qg��Îxy"�'�A
g&(�)�qA�8Y�xx�'y���&��A�$�0�B+�4���O*�Q �玑�nJ"tT�i��'�qOv�0�P�\^Ug�Ap:(a��"O�탢+c��rs���m(j�x!"Ov5��+c���WlW�-%&�{"O
,j'@�y���1I��@6�D"O���� S���JE.�1 �"O���ҎU�W�:h�PlP�*ErQ�"O�h�s�M�9�@;��D&��p�"O�y���P�A����N#Zĭ3�"O�]�s�?Nt���G�k���R"Oj��#o�
�6]ˡ½Q�x�p�"O$�����ga�A	��.{�P8iC"O�"��H7N�!h3E��"���"O��P�J�%U>]�� �٩q"O<,�M�&JT�Zg�X4I�ZQ��"O�DI���tmB��ţ�ut�$�"OX��C�T�^����bΰ\ZA�#"O&р�/ضk�E2cBG*C���"O���E��a&��G� :g�n;�"O�![�ƙM������j����"OP�zF��e�丐7�
���1"O��QW�ǑD�9�M��$���"O � ��B9�&�r0JK�@�4��C"O,qk0뜏c�Z]����$pvf)�"O���F��N���0o���"O||r!�;�a����=i
�"O�@�$+MR�H�Ɨ=�ZQ�"O�$;Sa
b�NE[Ə�es�"Of�3��SdM�����#o�N��"O��D��^�Fe+�V�A��I#6"Oj�Jq�h���v(�);�b���"O֑2���#u�e�$�V���a"O������@�PRp��7s�H��"O� �a�>s�m����,g� ���"O>�H\��w&��z)&���"OD�x`�w���!�D�J�4R�"OPu��n�-E����G$�;�t�Hs"O8�y��T�cK��������"O�ᓡˀ2�
���ˆ�&�r�1�"OI��SM�`�pƬ�<����p"O6�hu�ƭ(�x]���԰rޖ(��"O̼c���8K�0�ѿ%�"$��"O&���O͒o� �åGA/D�j�%"Ov�2�
��^U�aR3a���X�"O�ɠe_	Rn�Hԭ�zє��"O:u˖b�`^�P�攟\,��0O�|sЊbfPű!S�X$I�f�[7�+���$O�B )�
����C�	8��A�e��k���
0��,RGC�	 >J\���ȇm����6�tU�B�	rdV\�b�	�A�<�b�*(r�B�5kE�왂�,i��q�t�LpR�C�	�l�${������uW�N��C���I�"�#�́��Ƒ*i!�Z����Y�T�d�W#�W!�� *���G��"� �R)�K�j�"O�T	�G�GLزDG�	���U"Oxh��@�+#�J-p�D6;����"O�Tr��C;e����Ck@��ƥ"%"O�tٵΖ�I���kޅs�����"O�@�fO
~PB@"̔�XƦ�S"O��
���<������:�h�B�"OL�
����MR �(L&�%X"O���2��a�m��s**�{�"OX)���u�6����>A�8�sB"O���b^��@}Y0��mp���"O�=Y6�@�Q���H���x0�a"ON0��n�0*ݲ�A�HԵt6]xU"O6܀�J��j<UYp�Ҕ����"O4���_�{� @�A�F�tƺ���"O�8��N��ʁ"�s�P ��"O:�&�L5RN�i�ք4j��0�"O�A�U۰6�X\�q�O�"_��@"O!g҇d�x+���9?RHy�"Or����<8-b� ��W#+D�{�"O�$�v%�7!�*U��9,4��"O�`��ОZ���x@��Hڌ�H�"O<��U�V\j1�߄^�lܩ�"O
y*�J��7(4yC헓s�V�j�"OZe�W��Ddy�-�<c��%��"O�<�F��z�+ʲxV��9P*[r�<Q0��$�f�2��[�^�F$y�F�w�<�P�K�MH� ���l,�͘�)o�<���֝|��0�*���\�)P�<S�S�0=����M_�T�B��i�<q���{tȤ�&P+-�����_�<�������րQ�T�e�/B~�<kP�yLy��A�-���B��R�<�v�;&�Rx��,�6�y�E�<iGk�.�D�A'�ޮ2u�e����C�<�c��Mtnh����Q��PVDx�<Q0A"�TQF�'���&��y�<yФ�����!��S^�(&
r�<Y�̂�Lκ�z�ˌ�O.Q��BNp�<	�A��[
��1#�V"�Ho�<�s�S����*
=:�d�S�N�e8�lrRjè)��&����B k����o�!MЎ��Ԉ7D� Q���B4�{��S�F��d�6?!�,�&|8�ʳ�4}��	�9E鰸����4@s�5�U�ؿX�!�d�2gDvi:k��[rZe0�&5P�9cVT��y�Ĺ��\%?�L#��րO��J�/̰	�c4o(�O�\�ד�,e:b��]h���	{oJ�p�S� "^��āZ>(ȋu��_r���L:R|џ��Po�hSd���O�p�����:��H�!m�A1�EB&gQ��yR��=�6U���90��pak����ď:|�� 6B/z����銳r8���BB�7{V	��J%!P!�ɵ�8�����7j2�(G)�?d�@�PX�����j��%?�H"@eR�xY�ӧCH2����+�O�X�%�`2�,�EQ% D��"�V�_���Q�#� zU��$QZ����bJ�5����'t(џ��K�n�@jKc��B�H�@!�F:[��2���yb���@M(��/�4=�y��HS���d߄k.1� I&��)�'g�ȵ��nl�I@��p���"ڠ����s���і���D��0�|�����@��}&��{�I���<�Kr%��4�1��4D�X�]%�x$)3���IaB�&�p?1�I�Z7��A�ͦQ�\�1 K��ZM��$D�0r�c�;?#��B��-J?P���.?�F�p8[��5��O�6�3�$N�J� ���˟8N\-���� Vy��;^C����ܳ(��*��'�d��Ed�X��9�O?r��ǐh�cAm�=�X5��AF�<Q��]�<#�+��Y���	@}��^��2&Xϰ<����8~iic��.�4<kp*�A8�xàl�Q
4M�V���"d�_H��0	�����ē�Ԩ���zyp�����>}Gy�iS��������.x{��LՐG�Uf���¥BJ68r��
�"O"��fȷ]� )�k�(:{��R![g�L�E���w�|������ P�җ�G�����b�ʽ�y�D(Y��(y�"
�ͦɚr���~r�	
]��8�MW�Iay����qQ~�9��O�mR�S�K֘�p>Y���-_o��D�\�"��uv�Y�/��p� 
�'�R�Q.�3�nhV�)wP%���DU��F�Q���2�fd2f�0�i5�
d)&k�E�(�Q�gB��!�"�l�a�_#z�d!�CvsXM�pB	�a�!�'��56pp7��OZDɗf��E��9��&3z,�a��"O���`i
����p���$$��Q-ڨ��&��&a�;6��g�'[��!N/�<��j��@��1�B��!�E���-a�+ȸaǞ��bl��q�x�U��a���� ��p�LK��b�ܵg�>�=�@Κ�G �ɒ3Vf ���q��	0&=�"�!��,�B� A��?\�����0'>��P�.��<�g�r��'j��D�f ��zQ&L�Q�٢y��ҧ�O��=��ڧr�J}��J��W��5Ӊ�䟃�m
�,Ԧ�Pr͟��څ�^vܠ�5�5��;�
)^{��k7�a��&�3��|�-;P����@���Z�6�Y2����D,CM���A�=�'��I�	����Q�J;�i�tĄ'V��X�L;��>�v��'�vT�	ŜxyM�1�h-s��H�Xܡ�g4 ��O9�T�D���:��ذ�O�I�⬒
B<]ё@ƼRZ��0���T�'1⟔ڒ$� ~�*I1v$�uaI��q�ッ۳sO¼i0E9�Q���284��d,}��C"v�Q��g?a��٨�Da6*9�{$�1�����:��)S%oF%B��;D(�h�[K?6�yA.AۄQ8D�H���/�!È�L�x�D^wѶ����@��a�ȗ'?F�	�-eʼSdJЛE�vu�c�rְb?��C�wh|��$�S"p�Z�H{�>GFVK�8�=����;��`���g2Z��pr��%z�}��1{|�,����#���1b�Zu��&��t4��'�����4J��<�r+O� 0
]r\�tiqO(�Z�n�;��O�����.�!l�`��g ����IJbώ���@�����ɝLl�{�LH*��)��tJn��Ӆ}���R�T>�q��&�	��k�cT�(���[HOa����9��p����F�<���1m�(�%O�z��O �u�3?)�g](z��S@g�	=AXZ�o����o'� �9������5-Ht��I���N9;&�-{�`	K($�G��/4�N��C�\�V
4����=uq��É�#�̱�i.<�J��G�>��
�!L�>��њ#^?}Dybk��U�x�C	M)�q�e��İ>	�j��|���[)��EP%®\�4�e�X�nr���B.��P$��r�>�p%%K�ȝk���:-\dqG{��2*Ri���v�!��.�W�4��10�*e.B�jzR�*�
�p�<�ē�a%�Q
�t����1�L��
v����׫I+vĨ��i�8dV�ɱ�(\����#$�Ir���� ��B�	wº��%'�0�#�8���Qg��t���O?d~�K��uǰ���|��k޵���+Qm�l#�ɀn�x
e�4�O>�*g*ݬR�6l��%	��ə�/�h��p��X��A���ݝh1�D��R<�j��R�v���<)���:H�pH`̐�KxHԂ��g�'�H�����D�Š��m���˙
�~ �.Ƞ�ZH��)��(���PJ��$�!m�߈O:#4�1Љ��Y�:�����P��4h�Z�� C&|F�Ð|r�C$xL� �(qe��ȳ���>�H��F��|� ء׭Ed�'���C2O4)>yCgˏh�{fG^�B���e����	� ��Q��&j��\�a��m"�Z�8��\��H��;oj�qyW�
7|�7���/x�@��M���)�'��d�G�DF�a����d����e8d�;��LC�P1�	�]	��9F�FD��g�dEM��+fe#ZFč�AP��1)�����Q!l.��7��U�6(ׄ�e�'�~�
u�`�\��уU9e'NI@�DG�U�`Q6�D(7H�sV�	3�0�bc+wg$�E�G����"�2���I��3p�2�#L0zǬ�p�i�;���*����3F��O�\��T՘8bQRw·/�(�bN�&A� $` 2ғ�&�[�q��?�J1'ؿw>*�!6C�'��Iy����B �>u; �1&Cҧ��QI�R)w��C�3O mj����Q$ט�a�Vđ�*^��)S!ʌ�/�Z�r���y���<S��� M��'{�^�
SK*�:�c���-��� #k��偔�^Ohe!��WP�Z���Mp?qb���m�,����̭��>� �!1� (!ۦ%9��FJ���\� �Fm�*z8�\��H_c�x@�i؞��'��%j��2��-i��Z*>��Zb"�%Vx.,s`o�k����		Z�L��p�@<{h�����R�ܢ�	�]����f��Ot�1�H�/���e�K�?j�S�Z6	a�˕�0}�d��0
�Xb)܏LЅ��I@e�� PL� �n4�4�Iצ
����A���(,�#��Җ3xq���|%��"�;�"q�AW&����g�ѤV�Ĭ2���D�pc� u�.=���\V���*H��'bov9��$��uT��'	Q�u�,�b��PMx��̊	}As�o�+'(�~b��6��&�����;�ņ����<>��{6���yp���-!���[wយ3ʟ�*D��v�TRsm[I��!��'���6o!"숡��&�(��xz7l��	�*#�n؛9jh����'uŸ���-R0�(�(�'�Ф:�i��f�fD�&��T���0�'���2��R%^�2%�#OS��+ǧ(c[ A������MY�iK���q�'���we\���|��ό*k�.���[�Ƞ����O
���f["G��'סP���R��ve�%A��Q��0?"�V)UBt��+��%{<��k^{8� ��N/s����0��41�`H�D�X�m��=LvxyD#8D��h�/̫0f�y�C.3^�jYX/%}'�c�J�����J>=�/D�����Ԁ�4m�� ��&D�Ty��čV�@i���(��x8�CD�t|J�'R�ٱЂJ�g�Ɂ
���ɷk��`���ʊ[1lB�	}�,R�/�q���'�܊��[����nW�'��Xee��T잵XdF$9���˓?��)C�H���	�Ei��W��tQ�JL,p�
B�	4c�"	Hg�Ki��b�+�3�
�O��r�kI�����O�X�h ��"`�7�;y����'B��SA� �W�#y�����'a��S��Ԃ&$�9GrH����'0\4�e�׶`B �1-,�'v*Uj׋I�>lR竍�"�M)�'�ᓆ�� ��[�^7*��X �'��H`��'$�<ӳŞ�1A����'�j���^p4�"��]�X��'� �j��	�2i��Ѣ�N�p���''���a�E��-8��8���K�'��k1�I�{ �y�f:��'�N���I�Q��5)+p��`�� �콉+�>M6nD��KX+X �ȓ���6��g�Z�9 G¼��	�'����+�=�hr�$�2rW Eq�'�R(��G�d |ԫ���d1�,��'�
���jA3`��M���ҿ!�\�c
�'����Б3��qc�� #�4`
�'jࣔe��e���"R�Y�vn����'p����+y���&ѐn�؍��'3L�BU�el���T�@,R
�'T��ׯ߱4�>UH�!��V�Jd)�',�3ҊD;:��&�Q�LS��'��庑H��NbL-:�1��'l��,7?��� �K�1,�i��'���¢P�)5��G���*50��'<�=��	:Y�Jʿ)&)P�'�ԈXGHڷ"G��qC)�)"�����'�1�g�H%<��a�������'ֲ�RcA��z�
��-H
=��'ޞ�4�[��l%K�Þ1=����'�����iD8���3d�	�'v�={�i��$�mHc��9nD`�'���)Qc��L ��'Pd�'� f��:��I�ŒhU�z�'4M���ޛ������	jw���
�'�H�#	)SD0��Κ�0un��	�'s$�ʇJE�%C�W�7!�,��'�F%� ᚙ4>ڔG�4/�B�p�'Is&폵���b��$�"��
��� �����8-�T�2'ց."&�	7"ODa�Ò�tO�ZF�;�f"O��Q�W�8 ��pf^�pG�w"O�A`�a]-"�&��/H89E"O�1�'NR�H(�f'�^�� P"O41�M�
Q�x�;��P7p�&�k&"O�h`A�ύ���t�\�4��8�"O��q�SK�cV �;K��"O��	�@A�.�RU��i�!"O4H:7���:l^�س��4t(8�"OD ���ֳa�(ABG%O�y<Y�"O.@�6n�*TU�E����_�J|u"O�l8gG�8[�6\�'>����"On��dh��$u����'����0�"Oԩp.�<�P9�/�����2"O�ؙ�.ћ��zW�A��q�7"O�d�EK�3ܖuH�0Q�조�"O��E!I�4}��2�f�b���r�"O���G��A����C�U�)�d�3"OD���)x�0�� ������%"O�,��Xx	��Ӭ��5����g"O4x2�/�!8,�h� ���;"O%K"��I���3o]�&���G"Oj�I�䀟 ���q|"1��"O�a)�LF�"�Di��"ߝ'j"O�ؐ�Y�F ��a�W#O���""O|�RaY$
��(D"�7g
x��"OM�v��Ov< �P�}j��X�"O��j�a;0��Q1,��#JtYa"Ob��Q�!x�l�7At١7"O��۷��J�έ��+>�y�"O�T��@�S��p���	;�5i`"O6��oR)\�t	�F�D\ `"O�Y��-�H�`)Ǭ1�l!0�"O��w$ڨSw���h�6�H$�'"O�l8hT6��1�/���"O�hю��V�N�S�k�l� t"O�I�D)�5��}y�jO[@��T"Ov� �(0B���F��T1""Of8��eع'^D)���j�s"O<� ��n@6��a�6�,��&"O�I�ł\:��C挺kpdu�""OL���ծ.5�)�a�V�fnvp�"Op���BC�P���2�BBx�Ж"OT,��Gί|�B��AfV(A5�(��'���e���X��'� ��k����*C#�����'V�I� hn0T��>`����O$� 0N-�0�K�"|zL��E��prGl�`_���u��[�<�W� v�<�Ƌ�?4g�Tj���{��D�'�Ԉ)#II�h]�ϸ'{�F��3R�B��g��CKj��	��8AF�?7�I�1@˝%���s�F�&>��##Θ��0?���Ǒ=44�ǝL((P&��O�'E�̀��I�{&a���?!��!�^Î���(ͭX�����E%D�!C��N��aɏUwN�g�<�c�9L�Y�Hߠ�0|r���7jʜ�c�mΟH8�@�"�}�<A� -޶��Ӊ#5" ��ʒ7A	z��'B���@$�)M��ϸ'�D�d+��Z�U�����M�2`���}�H�Sd�@mO�ͪPO 9�,ȣC��}�́v�ح�0?��(P�V�,u��|2�d�F�'|^т��G>@��(��?	����#L���eӹ�D��Gl;D�H���Tp��@B�.qN�!"K7?�7�Y��cd6}���?	���6mB�HZ��R�+]�+�!��lN*�S���g��1i���<\�'�4y�腌>q��'��I���$I�N�+'�ʆM������ hd�qD��Lʩ�P�Q�H�Z����'�x�����&� 4���;��ώ�)����ȓ7j�׈�8�a�A�E�l�D|¡F�B���S�	-W�$��6(��|���(�ϢZ-!�2(��	���QHh�9X�IL9?"��
8�����C��ӬbJ,�y��iIv��f(ݜت(���R�'�))h^5v�2f�n��p@�>I�*A�Ą��GX�Q7�»W��d�f�f�p��5�O��3��L<PI����&O��(�Q,g�4�G �z�C�	�L������{���j� ݮY�`�<����I���EbA���Or1
f��2K�m���<`҈	�'�VUsd�_7/y
���.F7b���if,�D,�E�R'���f�S��?���ޢ �^z��]5WHx��s�<y�|E����;I<֬3�d�!��d��-��u�&��%o
����,�8�M��e� �؆��|��CfF0���T��قa���2�"
�D��4[�Oԑ{d��'����`ե|�l��I=�Ĺ+ć&��Ѓ oUe�S<ߜ�Y�A��\	��S�A�}PC�;4��k�MO05������y�Ki�<e��{�k�yn0Mh��!������
 �a�T%K�z���.0D��*Y�fu��ZiR�m����fڲX��7��]�*Y*���d2�`��HO>%k�@$�`9А�@�k�1z��'j�9j�2e��R2o�W0�hR�b�>:<���ʮ � YC5�'"��╉G����	��'8�
���z`���F�2���wr�0@����Q)�ɟJ$L0��0�:#�@զiS����ߘoB|h�O� ��T>4В���'1�P 4�2�\L�qL˘
�^مȓ ��8�U�����wm.��S��L���=-	H����L>і��B��ҁ�Y��D}ɀ�}(<Y�!��z���BK�{&1 �c[�L�����9-�����gRP���'8��<���˛D��L��=NtB�)�4�L�<�ܔ`�j�C�D*$Cu��͆ȓ SA)p$L�*~��Y�,�Ĵ&��`�X�*�Ш"�ӭD2` ��a��)
Y(QAH; 7C��
�v��+p�� *nU%�ALP���ɦV۾��O��!��[�T���8A&��6����ROry�t��(C� : �͏�\�5kȶL��Rt`O���>��dD 	��Q
�/�� Z���fx��1
*��8z�R��Y���X���eIZ�t"�l,D��sv/һO��3.�%b_�X�+4�E�`Y�D"ƋT��ȟ���a�7F¶u��4Y���"OJ�!N3)����`^�8�D��CT����OFɂ�3?ـ��$5�.�S �X>cT"5��S�<�$fۯw����:~�0OЌJc��j��x���S'̖�6�֕��'��J֪%D��	`"��=�ʹsRjMz�����,D�@"Q�\- ��0 �GL5g���)D�)�b��V8Tӡ��F��%j�K&D�X���ݶJXH��j� ,�`�	��:D��iG�F�}�����N�W�J9���5�OH1����M�vJ�p �a.Ŋ9!!�	i�<	�b�!e�����A$�H"��N�'�pTf9���#jN�TrqJ.k<����1�RB�I�8�\`�˥E�Z�0/Qj ���k��w�Dr����@#�<A��șY�eb���5�z�)��d�<Y��S�S����ƃ�&�0�"6��ȉ�?c( ���RM�'Gr�P���&|pHƀ&R�^؉g&��!|�ϓR�T���/+d%��g�!aaT�acƊ�>���竁9FE����d�WqҌ�B�/�'PF���oW�a��Q��T(�u�>�㊑�X>�Y�J�!2�����O�L]�R�˼p��$
�v�CF��7JE��cb+���q��q����V�>E��V&K��(�!|G8���ѷ~�����/H\�ԡ�dS��?�w*
.�<�aEK^�L�D"�,nrV�I�X�J#�4e�>��M b�Vu*�m�>A�'�jk�
�	��d�t�~��d��Ry�pq3e5H��Us�m�N� �q5g
4W�#=�Bl�&Y䲑�f�ݸV���J��UV��ʂ5�ޅ{5@A��Lq�e��5�<�q#��~ru�K(-��9!N�s�̽� |�ፉS�"�#r�Ζ�iP��	�o9���0�(W�8���9	N@ZC�Րy�b�(4��JM����`�$5�\	��@y0	���K8�ybI�|�z�H��� =1� X�Z�����;��[���Φ	�"K'�*J��>�O�c�+N�6J��@Yo���A�w	XA�}c֥	0j��Gs�  ��E�~�n�Rܢ!��G��],�3}�n�!ŤPP�b�_���:�����+��rf�1m*tu1�n ���a�@x�S
�t�$jA/ �J�c KG]E2�!V ���*p?��xr'��I�z��@40��ɰ�(�)M*I�Ӭ� �rdc���8����d��=�~)P���t����%(s�����<I���+s0u+ɾU�*�ZFA�A�'�� @�Y�=�D����w�D$�����]�t��V��}!תE�-�0�5�G-n&<�'�Q�'���"q�].>)��B��Ib����4^&����cZ�ҧ�ʱ/N8���(���
1#�q��u�o�.�:��E�Ṯ����_ĸ����L���Y5�͈|@�#g*�0b�剈7'�I3L\�|ȜQ3V�S7{zR�X#���;w�?ac@�}%���a��\�Q��:�O� �@M��
���c��<�R4�Ǖ+�� �%É�%GT�q��C/D�v@���
�[6Q>%�u3O�z���$+���x5C�#�t8�"O��wb^����SCH��H4ѕ���'�!��
�M1��#�f�ݾ��OR��KN{8T�D����x�'/N�+��H̟��dǋ
������)��l;�
�dv�����Ѽ�a~��u����&
��<q3`G��p<�W�*.tʔI,?y��MM(U��$�X綈A���^�<�%!\�C�E�h�
i�qI�MC�d��ب�2L��0|�V�k��h������Ԉ�Q��<�d W����z�@�0��P@ �P�J z]�O
�� @ӣ����0�RT�1b4�ՂR�M��z���
�C�L�N�Dn �(��ɹ�@�G&¬���$�O�%0P�m��Rw�(&�N�"��'+�t��N�&PM��ò�8S{J��r`si3��!D���*ހ=C�s��&(;Ud!���纉��4�)��=U��[�b��5�|Y��h�2C䉎1I����F�i�xl0`$�>^
�C�	7"����l-�l�q� <A��C�.�F {�#B�K�8����TrC�I?u	
 ��V��eY#�y���'���T�ɦ*q�Q��*|���'�p-�3F�;���.�vv���'�����3QO|l��jR�dp�'ShYx��y�tK���z��e��'�J��Tf52��E�hl`�"�'S��8a ƔyU����Kݜ���#�'���eg�|O��yVe� ���
�'-�q�B\J�a��k����y
�'G�ȋ���?c���Ç��©$D��`�
ԨG$.@b�덭��iy��(D�TS�h�9z;�椟�Kp���'D����) V�:/ݠn
z����#D�t���nrH����X�\z �H�h!D��r*��pY��2�A��>D�`ا��P���
K?"Uc�J?D�بD�jyZY@$�O�j|TASF<D�`�A)JMD��2qj�?*2���?D�3��4O�8A9$����ۄ`:D��	@M� *w��v��Q�$D����E�82g<"&�1_)jP���%D�DaC&^'{��8!�%߇��	�S�1D��2��Y�,Ҕ���s��L�:[��B�	�6��=���-J�ERA ���PB�	��<	�,�9����v���m�C������7W޶I��~K�B�	�fp�Z �g����PBG�8C�Ʉ:��mZFB�yrY�%X�K��B��<���*�Ɲ}4q��*��y0dB�Ɇ�&����0�QY�A�@�^B��Wͺ�XčT=�,����9|�B�	SM�Շ�)&L1��/J�=\r���"��4N�ԈAŐTB#>� r������}�o�S=�i��"O��8����&�uC�^!5�"O��sŠ�Rp�E"�5�Ģ�"O�%pa��=2=��*4!�?�:�"O�!�1J�wy�U�a�j��x�3"O��ЎM�u�ЙRE#�(
~�tj�"O��ѵ�P�U����"��<W�`�"O�y;P�� EH�bdV��P"OER�	/M?:0�p��]��i�"O�г�2�tR��۫o��d�"O���r	�-sT�q2��E�R���d"O2���n��$�Pe�ˬ��hi�D��ē�&��~��m��~�7hњUOnq�p��3k�4X(���q��Q-O1����|�!��o��A�ƫ	��󤥃�����l�����ߧ-f#nZ�Gd��R�����F]`�<Rpp6�L�[k����(M:��������O���[O�9$.l(Ah�;f���QP��<u0�S����Y��0|
gWlŠ��	�A�L=��p�r!�6��
?ꔣ n���өg�x5W�9W�qSB��]��r&��<�c�[�%e�lӵ�?����|�.��i⦡B���U���0K-´@�Gܦn(@� �
����$y��t�O�`���"�L�,�!䍄���c�4V�^ 
��Х3���8�!�8bla��
�.S(P{&ݻ:F�`�נP�)��%�"�B5gsҹ�s�n�P�
�'bu(�-��O�]ig�n���a� X�eCw�S�<�'an��T!�@�(���@'dؘc�>p�5�x�n�01��z�)8(�m�1)̛B�镇���y��N�W��Pℼ@�>}	�F��yR SL`���R6�R��f��yB��"/��*Aњ�~��ѣ�y�J�~�8q���]�b�囡�M��yK��a-p1jQ
�JD񱇧�+�y��6, ��S�=�r��g����y�:� ٵ(1�`���^�y��/���!�D̛6�ĳG����y��M�C2�5����3�8�:��Ӧ�y��C�������T�,vN��"U��y�ZǾH���ԟPFN��P�L5�ya�.TXR9�H^�W�p������yrϙ7���`ǅ�TRj4���yR�H�9�����D3#$\�e���y�W8i)���C��=���T���yR� t�Uq�m��3��2��yB�T�<Rf 3��!��r����y� �*	:�9�B��#\��7N@-�yBjU�^�L��f���Ԡ�wN�/�y� �=!Y�i��1��i:�4�yr�U7f����QR�/6P�GLS��yR�F�E�f���z�t$C�*©�y�,���Tu��°sp�a�f*���y�n^=@DE�&c�o��y��Z��y���G���QdbںNFѻ`��y�M*bЮ�"�ɝ]ڌ��ġم�y���-����DI��VdL��Siɚ�y���8?xx�T�U6H@ޠ#c��9�yr�+'^|�7-�7s�v����=�y2��7��mЄ��f���1ǁˋ�yR�/-ɀ��0F��[ڑ��ُ�yB��'.�恉 eH:K�ҍ�U�ӧ�yr�C�!爸�ek92&Ґ�!�>�yb�Z5�8�7�Ɨ>@(�fH��yB�[���ex�+Z\�P[���yba�KhL��`E�V|Vb�ʳ�yB�oC��� R��aO�+�y�Ɯ�X���-�6Bx�qrp(��yҠJ'#�x�+3��)7�ڰ��(���y�&4]܁�U���欘�o60!�� �q��.Ҍ$B85���gƶI��"Oq!�#�w�>���DE!؄ˢ"O�!��A�����&��h M0`"OdѨׯ�d�z}�t�X�Y���"O���[0?����刮!���"O�:��}���1j�*j�A"O^��PeտK��bp(�&b[��p"O�-	����;�����A�8vnѐ"Od��b[~��zR!��
v\�"O��G�8������4e�Ř�"O~��&Ħ⪱��#D!z_P:�"O���f#2RzPٸt"�'5�Z�q�"O �E�:���s��̶5��#�"O�l*g�W�Y���RAؐf0TI�"O�M�הZ��`sPB�'0����"OX-a�m	�`L|z+A�:	 ��3"O�9JGOOpZ��Ý�)���"O��r�DB�����/�䥱�"OX���҄G'��Z�3a�Tԙ�"O6�hR�s���0eQ(b�Fq�"O���� 6h��;�d��8c�"OxPFI�"�!��߉	��m��"O�9AF�î(�jH�#.��I�"O�xx&,�U�X(3+M)��T��"Ol�&Cõb�� �e�ũe?
1�w"O�1)��@[��Ѧ'�;Z>ف "O� )��H$SC=x6Ŝ�!��s�"O�QJS`Si�IR��f��"O<K�.�&q;�}���B�[D"Oԉ�է;���MR�or�!"Of�4,</��M�	�Y5"O� ��K Gg4kD뛽-ʒ24"O m{�!J-�m�D
�)�\\��"O���K�u b,���(@��	�4"OB!�G'V
�Z��p��m�3W"O�H0�\q �i�׋s�XI�w"Oh��&	����� �2���x�"O\��J�7+ǈ�s��ҩ'�@�z�"O"i"�N;o����#��7-�,{R"O`y���1����_�}��c "O�)���=���8sf�n%�a"On1�E���g�]�P�U$|�"O����/*~���r���+0�H��"O�	##�īu�#d!X�=�F���"O�[񂍹�1���T�R���"O$�q��	Py���F�T"C"O~9��!��A�l�b�Zf��N�<���M ������zV`�I�<��"8\��G���+]���`M[�<��-Cˈ�B���+���pk�V�<3�i2���G@�?��	�-LT�<i0,��rY q�E 4D�f1�Q`G�<A�`R�j�j��ݭq����U�IA�<Ye�
�X���n��zz�-p�T�<Y��ҩ$��R�+�����vH�O�<IV�؞)cJ�
g�� 5�!�W#Iq�<y���9�0�3� �/����Qn�<�b�>Q��<��	>u���,IA�<a��ˈ��"G���� l�<���;�����eN����Go^|�<k��~2�ȷ�Z�&�1����v�<i`J��| C��P
b����Q��J�<1šV.i�$�p�Ø�ceD��ŊL�<Q����
A��;S�MR�4�P�Lr�<� ���&My�6��%,�?:5TZ�"O���JG�B�@l��%���"O�]E$D:!0Ȕ�X�d��d"O09�v�M�5d]À��r��"O�� 0��*z��ʎ[�0��"O��H�$1'M�Q����Dq�"O$�ۂ�R�nyV$�f��06���"O� ��^>q�Lq�ǘT�`	��"O�5��Hd���Zׇ��;"O�m����j��)8G�΢y�j��B"OM;qlU$_��8E�7N���V"O��:灌!_S�����`�n!X�"O��'W�nl�ly���x��ȓ�"O��8��QF,��P��� ��h�"O�]i2�]*=� ���3Tt����"OƠK�V$WmHPk3Ө\�$h�"O���J�F��*�(P3Ix	�G"O*E���۔���A�"�`3XG"OĹaN� �*�Q�=[0T1(�"O�X)�M�8p!ܡU��!B�p�"O�����P M��8;E�SS��%��"O�����|���&?��
"O�hJbK�'A������r�!"�"Ot;�+��JKn��n��XsV"O }�W�>�t� �Ѩ)l�8iE"O%��H͋b��j���N(jV"O��	��ڻT��Q�ļ�1�C���y���0{�6�[�[�X��!�u�0�yB��9Za~쪵G>X�٨�jZ	�y�'�L#X� �󊆧�y!p�H�f�;%�R1xӦȧ�yriS�l�J�A�&�j�Y�
�yRJ� U*��"Hn��1��A�y��ݸJ,�̻��P%7PX�Ҡ�0�y�a�_=��+�B�A4 �!�.�y�/D�����4����5ͅ$�y�8K�yJԡ$P,������y�C�9���3I

f���$
�)�y2G�"9�0���	Ι9�,]:����yr�N�x.�չ�n�%h ���`��y�/�	�$43��[��@��D*�y"�L!y$�7@X�N���_��yR�F3����ǭ�8y-��Kȏ��y�l��:̺a �g�q��(�R����y��_r��J�gT"p��u��e!�yR�DX1
s�i+n��u�a��y�ĳ�����O��k]� Y�DU�yb�[&� ]�$�HeKX\���y�M�t"�����\a!��Ɛ�y2��ba=��ț`�ޔhPC)�y"х2k��@I��#L&���ƞ��ybI���ʴ񐁛��:D�S�L��yb
�2W5������z�����_��y�D�q5|)�C	�4;"Xe�n��y�C��H,<�$-�2,0�ô�8�y�ʛ�s�DP������`M�y2�U ^�x1�iI�e�6�@$�[�y��6bp�L����K����2����y��[�b��i��)Z"r�Z��q"�y�'	�0�Ա�A�ޡ=��T�`�F>�y��s�$�K�	@�98����G�y"I��y�n404�2>�����㑶�yb��xD�͸� �'63��Q7́&�y��@�=�vD��L����%V>�y
� ���$�V�����!J]�h �"O�m��3^� {D���D"�"O���қZ�2S�X�%Ҵ@PT"O�œ�GO�o���1�n� $Pd� "O4��6���`+AȢB��څ"O�ya6��|/�|�Ȕ!�.q�S"O`k�N%�Ze���$"�8j�"O�I��:�Q@ �ΒX�P�k�"Ob	� +��_�n�	 �,Yň�C�"OШ�s��L̠�CG܌u�Rps1"O� 0�]���E	p�x�Ρ{�"O�[LG�Kl<���ٞxx��J�"O�g�E!e�)FF5do�L�"O$ ����^�����b �L� 2"O�����.l�.�Aǡ�T��@�7"O��01cD�Q����$���=���k"O�@ d��!P���ұ1kX�8�"O�@rs��7]xL� �U�/U"�"Ov��6�(��ҊW<mi$�y�"O>���hA�'$֑X��[�%L�,��"O��0v"ζt������/[;���s"O�T��<*�lp�@��$��W"O�aْ�?�6]�u����U��"OVb�(�31��ئ��/�F��"O�0���G2K(�q�t(��H�s�"O��ca�4F�"p#s�9���� "O��bOCH��xb�?X����C"OK�6!,|i�#Ye�DK��ƹ�y��0,.�3�A��z�4e��ܒ�y��
� 0  ��   �  N  �  �  1*  ~5  �@  8L  �W  fc  �n  }z  a�  ��  �  '�  j�  ��  ��  :�  ��   �  ��  �  ��  ��  @�  ��  ��  
�  M�  ��  � 
 R � K% 4, �3 �; C ]I �O R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(՘xb�'��O��(⃯"T�����Y3s��eX@"O�-Q3�&&���PFi�&��{W"Oݪo�����XsmF%b�N1��"O�����?l-�pp����k�j�w�"4�L���%U�\�5�Շ<`u!r�!D�����7D=b}�����z@Bm���:D�878B�lq�ɣ%�6o�!��޴%��q���T�D��=��@خ�!�ā%"�na���̥a�A�Ve#�!�X%0��I�3bZ�8u [�6V��}B��ȹ�V��T�S�&����pb:D��1�)\��j�;�lֱx�v���A$�B��?���ӽmTm����X�P���!D�Rl��A�65I�`^0�P,�bƪ>�������B��a�B 	�+��B�	�x���s��q�i�5@T%,BB�)� �}�Q/nI��x2�ݡ ��B��j���'4�UAW5= �@प
U�=��;�~�D.M�]<�2Bˑ5� ��ȓ�r}���X3O�Z	3fj�h�ȓM���d��a�0�"F��SBB�j��)����V�o�Nur�,��=��5D�X��5{�,�Y��M)%)D� ��N�^$��Nߒi����V�&<O�#<)�F( ����� �+���2�Tq�<A��A<0�s'Γ�N�6Ѻ�
l�'�ў�'X�
 ˑ�I�G?bb̓q7����}�`�S�.'w�h��M�s�dFx"�'L&��ħ�E?�hbl�v��'�\�ehʲ$|Ra���l"�'���K@�`o�T[�*�']a� B
���DB�Y��As��0Zt����l�!�dL�d-j��F��_�~3�iU�vZ!��8�T���	3�MK7뜝xM!�ޛ�	���4t�p��A6!�>Ю̊ �I��R�r��/9!��0K9�E�P!�,Vzډ�sG:�!�
#r]0��)�.=�%���B䉱RR~��E�A/^S�ɇ\��B䉰-dXӌ�<Wy,�x��ɌB䉚��#�]���-��,�>E`B�I�$wD���!ż��9�e�ͣ6�PB��V��`����I�����U{�:B�	�Z�փո;�M[�dA& ��B��,|��1B�	=C!$ccM��B�I�5���̝~�:5c�c!h�`C�ɤ�)*�%�7C�`TI�-�D��C�ɯn�l��3
��2,*к�$8:�XC�I�LP���E�3ZY��q��ϩRd6C�I�U��{��9Eֈx�N�X�$C�ɚa�4d@E�Phu����ό6,#�B�	$Rl�@�d�I�H�j�ba�GhC�	��N�brD�!t�XT��UT�,C�ɖ7>�Y�#Ó�y� ����HB��9?�B�P���?5�q�񥅻b�B�.zY@S@ �*l!�(�1"�B�I�s�X8��`��9�L���J�f`�B�	)PN5c���,[|�jE`D{�B�ɻ}c�PbC�
4 �[ o_� ��B䉀�82�CD���5�W�A�RS�B�IS3JU[FK˫W��M�*L$idC�	����PM��U(�ꊹ'�\C�����'��yM�U ��!>C�I.{��8JF�Z4mq(�@�C7 �|B��z�\$��m�|�J]�5G~C�I{|6<�f��6S4��h�<��B�	����ha΋=�~��`	O�>��C䉂E�4`�R7T� $�L�y��C�	(���F�F(C:<�C��:oF�C��x��Dq���u��g��C�I:sb����;g�} !%�>@BB�� =����
�1!оY^B�ɜJ���"&R�/�d���L�k�&B�
^#�%���H7�vQq�		l%�C�Ig.(���0o�XM ��G(n�~B�I( �Z����IczDq#�#5�|B�	�5��5s�O�{ˎ�	$�UBlB䉮qDؘQ�dqN͙�C���B�I/ôX#U����#p�E���B�	�+aF�r���f"!��=1J&B�)� �q!O��<����*;2Yh�"O���UA^	4 h{���+ �*u"O� ����T�!�kPp����"O���#�Y�9p�0��o� X)Q"O�|���^�w��4p����
��'dR�']r�'��'��'��'j%{p�S!)<]�쇵^�:u���'���'Y��'�B�'�B�'�r�'߀�/	�����%�1�HK��'V"�'c��'2�'���'�"�'X~�8��UxZv ٖQb��R�' r�'���'���'�'h��'�lT�0*� '(x�:�aɨrZ�@���'�R�'a��'k��'^��'Pb�'Ҥ��� �dԼ#0�&u� IYq�'^��'H��'`��'rR�'���'PV�����C�t9��Ň�?��J��'���'d��'Jr�'���'�r�'ܲ�#a�?����Ĭ��@52����'"�'?��'F��'�"�'���' ����H=8�<đB鞡7���r��'���'�2�'%2�'�"�'b�'qrMw�N�M�H�3��y�	SF��?���?���?1���?9���?Y���?���q��e���M�,��UK��5�?���?��?	��?9���?��?�V�K�@6���,ۘ
{i2�G��?����?q��?����?q���?9���?�ԩ�lQt����r��1���?9��?���?1��?I�-��V�'`R��fh�d���jBt�����Y�`��'�U�b>�l��D(1���A?9n p� H�I<\���O��lZC��|��?�)O�F*�YP�T�0��$v&@%�?��VX&�M#�O(瓉�:J?5���[�,�V�b�u�0�Iןؗ'K�>�w��2f)4J�:Q��T�����Ms���l̓��O��7=�^�a�'ˁ3���k�윶w��!r��O2�Dl�`ק�O�nI��i����
�2���ґ}j6Uuk�4+$�b����P���=�'�?A�h�c
�����T	a"���<i)Op�O�\m"��b�����Y��Uʁ*
 ,SX�B�n�Q�s��	ßT�I�<��Onȋc��;�@�%#Ω=|������	�~�.L 7�"�~�"�͟�qeA�g�(��*Q2^�R1�W`YyBV�4�)��< IO8n����C�����o��<ɣ�i$脹�O�n^��|�7�X�`���J�옠b���OR�<	���?���#{���4���{>���c	j�xT·�?k���&�Y�,\��;4�&���<ͧ�?a��?Q��?�gBR���ZJ�2]v�}��eC��?q��,jZ���O�'�?9��?�������Od) ��
o����t���b�2X��jFy�'����O�4�'�n�1�Μ����3EX0Pdn|�@L*̜���'K�)%�Ƌx�\1 ��䬧ON��(O\!��$���	�,�"�����O<�d�O����O�I�<qq�i6�X���'�����J
-U��z�0{T�庀�'��6-7��)��$�֦Q8�4�?�Q�[!D�[ f8`2�;���y��ٴ��d�7�\�����Ӱ�u7�w�x���� (HY��A
Xv�}p�'{��'Vr�'���'�lCbaL�ȼ`"�H��t�5�g��O��D�Od��ɡNg���O(nm�ɊC�Y[Uޯ<����ދH�Ĵ$���ٴw���Oβ���i��ɋ��]�e���QsF�B��$I��I���Z.rf�ny�a���|���?���s��<`�j�$j�&m����2q|n����?9/OX!�I<�d�O>�Ľ|zV��^(P��`,ظ��#Dv~���>���iO�6M7��?�;D��9ur���Sa�.IxWmT�C�YPT�W�M���'��n���?�'�<ͻ�ؙ8VÁ1��Xsb��[L|1��?a��?�Ş��d����r�,P2oad�S@��aL�ś!iU#� -�����޴��'��nB���>s��x� f��bZ���Q�7`�6-�O<��q/mӰ�z^�M�#�����O|�5!%�υU��=���@�!s-*�'|�˓�?���?y��?9����	��sQ�8��&@n�Rpsp#A/h���	!l���O
��5���O��nz�+E��J��H���x��� �1�?�ٴ����{�:�B�4�ymR�C}�Aʀ�6p�����<�~��E��u�7�\ʓ<ɛfR�����	�BJ{�ˀLT�_;�C"+�ԟ��	� �Iuy"t��M*5J�O����O4PY�I�\a24;���g�xa #����DT�eC�4��H��H0������	�q��,�'�,�y�E� ׀1I�\�;R)��D�	�?��
�S�1��Bx ]	��ݭ�?���?����?����O �J ��^;�9Ȗ��c8F�¦��O�`n�3B�����ȟd��4���y�O�=;�,�S���,yN��L���~2�'
���'C�Ur׼i�ɞS@P��O��Ћ�����2Bf$�aU��W}y(y����|���?����?)�\]C��D��ge�9Ѷhz(O�1oZ�o6���Iß���c�ß�h=��p�E�Q����.^������
ݴ��Ş V�6�Q�b�@��:��a�%NQ:z#4!�OR��j���8BD\��Aݴ��$D�� @�N�H�fD��N�a|�t�� �w��O@���k�g�"����В+�4�K�-�O�HoE���	�����蟬 �Ǎyo0����(b�F�{3k��r�`nZ]~��M�]� ����'տ� P�K�
T�ى��K�:����<O���m�`\�A@-sϬLb��K�%� �$�O������7�r�i�'/�TH��4�����M38a@���B)���OD7=��4��b���H8��s&�&��$���O%/sԨɠ���.c���H��䓭��O��D�O��$� i���@
��
tL �����O �z4�fcؓ�yR�'F�[>ɨC�=F��@�@<#�0]��i1?��[�ܚ�4It�֯1�?1Vf'}`41�S�F���-�2a1�qj��?sP���|�� �O���K>��m�o����+�9W�&DAU��>�?)���?a���?�|�,O�o�r�vp��V/-��p�	L��cL�ǟ �I;�M��B��>�Ӷi~�m��x��I��ȉ�(�+��wӨ)l�V�l�V~M��x��i��L�IS�:�>��gʓ3�Z$+��-I��D�<a���?���?���?�)��Q����������C��M��.Ȧ!p0���T�I�� '?]�	��Mϻ(&���A&�;isr����|h(�D�i��6M[\�)擏l�`o��<9�� ?��$r)�iXL���E�<��X"y�v�D������4���D_!i\� ǎ�:#i�W�#_�����O����O$ʓ!��T74,2�'�b�(��uXQ�S�3FX�3D��<�R�|��<����Ms�xҤ�e[ba��@')���릧̳�yB�'���bʍ�LG�l#�O~�I��?yF��OV�ք[]쪩
"�Q��Au��O��$�O~���O�}J��B;����
K��Y��^'tk|K��\���( �3���'�R66�i޵kP,R6�.����o�0�(U"v��ٴۛ&�{Ө�z`kz���ܺ`��埢E�A���X+X�r4g@抴raN������4�����O����O���L>�*ǖ>�Y`P`ŐW'��|N�F�/��'����'|DQ��k�/]\ %��y�Z��S�>y���?qN>�|���<L�ƨP�	ړ>��J�f >�r�9ݴ#b剢6� ݱ��OV�O�ʓ'�°%�v�x�A�ǟYNV0q��?���?!��|�*Op�n:QO�,�I�Va���4 ܛ%A�$#i�g����	�Mc��>I���?ͻC�ٱ��(k0��b�B:ZE�_�M��O��>�����4�w~	�$IR<)츬�K��Φ���'���'���'h"�'���y�!OX1p*����`O.Z�H�嫿<	����搱���'�6�&�� �J�i��b�&L �ʔ�Q��O&���O�	&9��7�2?�;2��h���	��0ж#e���"���&�~�|2V������0�	ޟ{@�իI��<s�f�<r��c�������~yR�hӦ��
�O��d�Op˧8�]� e�{�XY�B]�o�L��'���?����S�dk��t�v����(F�	t��P��pJ�Ɖ$r��š<�'0O ��Q�I�YE�V�j�SuCN';jI��ԟX����)�}yr g�2��Ԋ�+J`P8k���:z�t����ʓ{���D�OH�o�l��~��I��@�gE@"	nR��)(l�Lԟ(�	�8��lZ^~Zwgn,Z�ݟ�˓n� }3�����X!-�e������D�O��$�O��$�O`��|�ƣ�v�@]3���,f4e����*L��� 1k�����\'?i��+�M�;ecp�g����h�akk!6�?�����S�'j�Ep۴�yrEȝR��AE�O1��9�N��y�O�/P���������O��$U7�V\���-���%��S�8�$�O ���O�ʓ?���� ��'�"c̖Q\hTI�˼ e^\���(G5�OBI�'<�'f�'���<mqӢ#H�K&�r�O�0����a��6mg�ӫN����O���f���HB:as6�M�]$��%��ON��O����O�}�;[4��N�$���ht�Q�)������$��N���D�OޙlN�ӼC�m����8h���4M�v��$�\�<����?���~*�qߴ����u*���.(]��/^,=5H�R�ր<�Z(।2��<�'�?����?����?I��=.o�9	��*E@<���׊�����iK���ƟH�	ԟ�%?�I1u���G!UƆ}R ���-�q�/OR�$a�ld$���$�s�H��@��}`tbd�&!�j! �8��OH�B�ty�kR5=���{�
܀���0��T��0>���i�,�ʖ�'ꜰy'�C'	��e�P�>c����'w6-5�������O��$�ӦM)P��0�@�"�	�1�B��qjBf�J�mZs~2oǸ	J�����'����dԖJ��3��9��t��<����?I��?Q���?����) 4�(�I��ֺbȘK�G�g�b�'�Bj�6�s�<�
��R�]%���s�� Dp���׉n������(���?���|��Ɂ��M��ON�q�k�F���&F+��-,VOfaA�ʌ�0��|�Z���	�t���� ��εn��r,�:F�B���J�ş�	dyr�d��Y;d��O.���OT�'؝���0*����%>Y�ִ�'9p��?A����S�ċ��7�^��L�z*D9�
L;a���{S&K5*�d���O�	�?9�� ���r���3a�43��1�f�+a����O��$�O���)�<�3�if� �� �^�H�0$�E{a�Tx��'D7M$����Ā�m��O�^�,�Aj *����s.�&�M�i|.
3�i"�I�_.����O������ |���݀g=.0��g1<��0O�˓�?��?����?����iR@o��@�@�M��=�r��,z��UlڦcL��I�����e����	���s�e��dF�x/������'�?����S�'mq6hq޴�y�he>0���Q�Z�p�A��yb惘b���������Ox�$Z~ZVu�D��;|9Q7�ǹzS:���O����O�ʓ|)�f Ȅ>�2�'����WS^��g�47����A ��Ox�'��'��'u.EI�c�-2�"4��k�);B:���O�E�e�Ea6�BO������O�p��DG�0��RoͺLPdU��f�O����O@���O
�}R��V�N�P#�J%7t�1�cN�
� ��6����fFr�'��7�$�i��[5 #u<0����Y h�D�S�ee�0����ɌLz��nZS~Zw�D�[�՟Jt�QA�&��:!K� o�0(�-�Ī<i��?i��?�����1)L �{g.�Wq�iP2^�$�'.67ҳ|�����V�'a�O���/ � ���1>kL��	\�k���?Y���Şd�V,a%-A5[d�9#.^ߪ���Bл�M��_����c����6�ī<�'�fb�u-A�^$��-�?���?i���?�'��d�S��V�h�b$כ0k�T� T��$�jR����۴��'f���?!���?!5`ֶz�(���(a��|YQ�۰n�JU+�4��EX�V	��O�O�'.ȒGQ�+�{A�qju ��y��'�b�'R�'���	ѽ'��7�'0�dR�G��1���O���C��3[���/�M�H>A�B6��gl�4/߼�����$��'������A�h��曟0�*ۧ;v�ZW&ߪ٢=c���1
O����'q�&������'�"�'���[e�5u��Q�F^�8�z s �'��^��J�4_بΓ�?����	X�k��@ZF�J�O�H�#�/��Ƀ��$�Ŧ@ܴ?�����^�."�-;֋��q�xl��H��!��H0� Z�|�`�����&�2WO��!{�(C7 B*tn>�hT�<_���I��l�IΟ�)�Cy��aӬ�s���T�H��PC�G�֑K�ˆ�Y�����MK�2m�>���i�p!+�K�h��c����%kw�l�o�%dƎplT~k	h,���\��qAk��{<��cgZ� v:O���?���?����?�����ߦ+(�Au�#<r�1�T�Ƨ-0`�n�V5l������	~�s��i�����nZ�1nL �S%{s !�� 	�6�m��P%�b>�c��͓b߸���.4�2�	De�ER�I̓?��TR)�OQL>)*O�I�O���AIԘ;�����K�yb�O�$�O��$�<v�iEl�A�'���'�Ber������X D!�2kѐ ��O�e�'86�	ͦ�M<	rU�m�V���%ɥ)�VԁH�Q~"�KK��DRS
P��O��d��@��Y�6�z��I������Q
^�r�'���' ���c��nx.�(#m#_�n�����ҟ�K�4����'�6�=�i�i�3<pa���<��(v�X:�4n��oӼ�JG�y�z�x��/���J`-��x�a	v���2`b�,��A%�Ȗ��t�'��'B��'T��TGF�:�IQ
	'Arj�@vT� IٴH���?������<���ԧP	h�P�A���=!�-/gI����M��i/�O1���YQ��5���`VK�-O�E���U�����Zs;�{��5�O �L�ޭ�F�~d�8I�Lx`���?1��?��|�(O�nڨ|X�q��(j���;��M�w(D���.��ގ��I��M���>���?�;r.��Tl�7�B��#ˉ�{�(� �T�M��O�M�h݋��t���w7�=�FNR8 c�=�%Dou��B�'��'�b�'+b�'�N��NCH1�(v��<�Ju�wn�O>�D�O�AoZ�X���ǟh�ٴ����C@�Ь)4��㠣ٯ`xɫH>����?ͧ)�bSش�����chϦMx�ͣW�$��R�HY�3���Io��Xy��'l�'G�T�\�i�G1N�����-cR�'��	��M��eB��?����?�(��-J6+͗l$�ib�9a�h3@��,��OF�D�OԒO�S�rG�Q To��b�	J��	S�Y+�B�	wְo�)��4�Z���'��'DM�1���9���󉞼�D��'iB�'�r���O�剂�M��J$���J�Ä�%�| ���<"`@��?�0�i��O�D�'8���;�*!�U�EQ�t��Af�%	��'VN$��iR�iݙ����Xb)O�i�Rd�ܠM*f��5,�
�3ON��?���?��?������e��
�F�٪��!#�oڜ ���'qB����'!Z6=�d��P�T�}ux�E��+�f�A�O���7����-��7�n�$
�!�>Z�x�raڏ-BR=a�Kb��S@�̈́/�� �$�<9(O0�8�f�hB5J��<Z���#�'��6-̯�&���O(��ʗ�n��vQ/k������m����On��O�%��2!��<5�NA�p�0[$2!*��,?�Da�h��h+�4��Oʜ����?a2H f$ "�CP>mL��ʵԶ�?����?)��?�����Oy��/֜�! ���)�@�ë�O� n��-� ���`cܴ���y����R͘�R�OڠH���h4����y��'<"NiӜq!�jӐ�pJ�4��n�?� h��Xn���D���q,���?���<��D� a� x(�7s`^	 p�(+���:�M;,��?����?	��$
�N�H@P#�;%�Y���R�T�1ݛ�q��I'�b>a����|�Ȁ�bn���	h)�0���\>v	��_x���� �O�%I>�*O6�)�"��SqV-�2��b!;���O2���O����O�)�<�D�i�H����'N��ʵ��:5n=���I?\��`i��'��7m&��0���O����O�E� BD 
4�� 4�B]b�/��>Z7�.?uI�?v�8�SS�S��Z��0Ri��Z�K!:��L+�Nj���I;I��B]=5�h-��}h�����������MÒ�P��
o�
�O�hb�M2w4����/��1�"� I��韌�i>-�^Fb7m>?)P"�1}�x!Y���� F�I�oY#Zr��)�� %���'I�OY�A�F%<�X,3q�b ��F�I�M{B���?i���?a(����G�9$\Ī�fĎӘd������O��D�O��'��[��-��HF�a[��yV���m�H����עfm^LJ�4 ��i>Ys��O��O�����D�&#θˢ	�8c��b��O���O"�d�O1�l�Eݛ��Ob6 ��4�&@����L� &�|"&�'@�yӞ����OP���Sֈ`ȑ�ǀV�P嘒� _Gx��HƦ��E���Q�'D2�IF jz)Oise�ւs�"U�HB�=
��3Oh˓�?a��?i���?Q���򉂚P� ,���5Fx܅��M�>.x�xm�`���I�����D����I�������j��x�f�?i�Cq.�|��i�ڒO�O�މ�Ǵi�$� 5vL*E*�8.����k/U��Ǥ�\����v�D�O^��|����`��-X�����'�ב@?6����?��?�-On�o��#ZA�I���	�-
\��K�,-xCi�=TVh�?��V�ܛ�4����-�DU�b�����J�]�.a�CC�px�ɔd2�]�2�H�*�'?թ��'�*����:����ʙy�z-!E;���I�����Ο ��o�O�R�sY�uᘤW�.U�1k�!��v�����O`�������?�;i)*D�-N\�|
S�Ӎd�(ϓ���k��\l�b�j�no~R���E���h�p�rL�&ÜH��#
��țp�|Z���	���������Iៜ����Q�N(a$�M����!cyB�b�P�c��O�d�O�����>s���%Y
����ʬ"���'+��iVb�O�O�<��EGFx��3�ʇ�i���㮒�pd�)#S��k�$��H��L^�Isy"�J�a��kg�
��X�	ŋx���')B�'��Ot剮�M�� <�?W���ʌ"s��0a�C���?�ûio�OX��'���'�2�	�aT�x�����|,"bK{���ųi��	-q@��`�O�q�H�N�Ƽ��, ���J�g��D�O����O���O��d*�S�N?��e]#��L��!_5eL���'�rex�l!�=�V��Ϧu%�d+�C٢+4����ʳhQ�ٺ'�Uw��ӟ��i>u i@æ��'ۊ�Q�9�l�3ǆZ���͒�G��Sȅ��8sm�'�i>���ӟ�	(,��ܱ3�Q����b��V(/�:A�	؟��'��6��Xh���O~�d�|��
�}�Vp�MH��`�H}~�f�>����?�O>�OӠp���Ĝf�Z�@��6M�
�[����Ԩ��4�fm��!r��O�y��E�+07�#��nm�M��O�D�O �d�O1��\j�AM�T��l�C�-�A�`P+]A@�@E�'&R$c��pX�OB�l� 4Q�u��[�1z(�DN8O�>�S۴*��a�!����@�D��3�T�~���҉&����A�6Ge�T�7�X�<q*O���O��O�$�O��'!�֝�lD�mh��&o�=H8M` �i��8���'�b�'E�O�2Bk��.Ѧ[��5�b�!':�`��=hnZ�M#w�x��D)IM3�V6OVb%f��^G�ա�/4bɆXad5On�p�?��L(�d�<�'�?�QޛM�v���tm��raJ�?���?9���D���i�,B�<�	ߟ(kvl�pF]��@>:��a��s�l,���M�#�i��O\�ꀣ�#D�
#˵.��1@V��P	�M^&r[�1b�%��rS���8" oQ�T�|(����"	|(��B���I���I���F���'��@PlǬ�*��p� ��2a��'�6��l���ORAm�c�Ӽ˗b�]Z�<P�lԼQ�LPR���<ѳ�iʘ7�TĦ��%����'�"�@���?]��$�HO���'� w�6|r*X�bN�'��i>��Iן<��矈�����Ik��^ 2�k�@.pjy�'�6��12�t��O��D)�)�O�yU�W�Z�9�VMF<;v0-�֌�T}��iӤ�o'��ŞD~�����/�����B���01G��,,�l�'-\�`���P��|�_�0zv��3l�K�;z�P��A��B9d���O&���O��4���l�/�?�#�_�o0��z�˂�߲-�����?Q$�i+�O���'ü7^��ܴ���WC�'��]:"/�L����B�MC�O:���"?�b����w�~8���T���K1@�)<ԸS�'���'O��'�2�'��*�(W��y?���"��p����Oj�$�Ob�lZ *���'B��v�|�d]gޘb�U�z��D��K$O�$n��M�'�x�	�4��d�$N�� 
-�� ����Eo��brf��a!���?I1N;�d�<�'�?���?ys��=v��pyS��_���	lN��?������������(��쟈�O�$�HS�F� I�\H�,��'��XX�O @�'\��'�hO�i�O�}3�T�:L�i`��q4V4�4A�7?����u�ݖ'����i?�O>��V�n����.� �D}���W�?���?��?�|)Ob�l��:B|i$�E=��T�T듯{��@,�֟ �	0�Mۍ�	�>��~� ����� xY�)!Y�5�������%.x����`h���N�I�<�&�	�<i�nf�q�NV�<�(Oj���O��$�O����O�˧Bb*X)��Ѣ�P���#�*�Zf�i�RŰ��'��'��O�R�}��N' d��mG�u�H��Q����D�Or@$�b>�Q�K���ϓk栵��mR�o��P��U����xخ5 f���H%��'Sr�'��	g��'s����ǫ^�9���I3�'V��'��^�`޴E~�C��?y��sD@�Q� �AT�KQ�њ_]XEY�b�>Q���?YA�x2�A04h��a��hߪ��u�;��DoѰ<21Kd�x�%?a4�Od�V�-	�0c�e.OX�k�
��\6 ���Ov�d�O��2ڧ�?��n̺$@�x CM;&���W���?!@�i�Pj��'��h��杓>h�A0��2 <��͚~�,�I⟬���M�!S�M��OX �dm�?��4��.#�z��d�@/4�ʰ�4˯/Z�'���֟T�Iʟ��	�T�	�:wXlSH�5l@H�O7\נ��''F6�0���d�O���-�9O*�u$�4}!6(�%�0-��ԱÄ�N}�qӘ	o����S�'}���a��]'@�<�B�$k54��V
P�]i���'�j�P�,�⟼��|�\�`���F-6�@V�( "B) �ʟ����H��ڟ��{yfӄXBB�O,��(^�	?v��g�M�܍a��OHnN��~���ҟ8��䟈��±@��H� �6K.p�3]�|qx�nD~��tv���Sgܧ��S�lT j;p��4��8��G7���O@���O����O���7�S��U��!N~�Z�i2X���I䟨�I��MceN�|���P�V�|��љ�y*��S3�����F)�'�����iQ�u!�V���xt�D���L�L^a$R�)3 b����'���$�ĕ����'.2�'����#��(I�2����l2��'0rZ��hٴ,�,đ)Od�$�|�Տֆuxjћ�� Ojl���
y~�h�>���?yO>�OM�Ms �-)�n�c��8YH����d� �p�!�V���4�����qa�OJi�aK�"r\i�C�$]�N�@�O����O����O1��˓u��'B�i�e�$��2�aX~�U���'IBjq�6��ˬOZ�kظ�a����h-x�!4Z����O�0k��x���-f�) t����O�( ��$�
%y��+�L	����'H�I�L�I�X��ҟ\��o�d����� �_�7:��W�
,XP6�ڱu����O2��"���O�mz���Ԭlj�Q8E��RIʹ��П��	D�)�S�yL�Il�<i�A>Ô9хd�m?���ӪC�<�3L��TI|�D�����4�f��W&*���qnl��'�d�O��$�O�ʓb2�v�2?��'��+�f��J0�P�K�ćO��O@��'��'��'�\MSU �7qZ��gcE�f�D�r�O��KA�EH���@5����?5H�Or)&��?�t-@�.�6D��-R!��O����O
�d�OJ�}�;[�)B�@�v���4'z)���3<�f�����;�M3��wC�� ��2sL�s<�@��'�7��¦���4
n���ٴ����v�J���'d�-��H~�D��`�^�.แf;�ģ<ͧ�?���?!��?�I�9ܒH��м���be
����Dڦ����ky��'���c�Oڵ8g�;EM[0{~���d��{}��}�4o����Ş��!��\�<}��'��2+�@�ٶ+XS����'S�QbC��򟜣��|"\�X���ͽ!��=�h��!8�X��L}y��'R���]�,�۴���͓$�|�X�\�T���f�;��H͓S���DLP}RIl�,=n��M���? [��8`a�"�ql<��@޴��$A�Y�<��'��Ͽ�&b���v-�Aƀ*3j5XM��<��?����?�����ɀ%���Q�(��a1*�g'�Iʟ�ڴƦ��'y47m(���=`�\�cvd�6s���A��/
��'�T�ٴ���O�	�#�i�	�{�����-�+��q�$�L���O�"��Yw�Icy�OJ��'��#�9�޴��Ç+8<�+bN�L��'�	*�M�C��<����?/��4��Ɔ�-��Ÿ%�^9C��җ�0�O�o5�M�q�xʟ*ɠ�S�(<"g��-'�\�6M�\��ңu��i>�� �'��U'�4�ì7ybq�(_�{�z��V֟��	�x�	�b>�'C�6�M) �e�4�D����$F�i�Z�ۖ��O��D����?Z�4i�47x��!kVQm��j�J���@r��i6`7�B'�\6�*?��@�]i���<����BO1K��)J�&p�-���y�T�@����I՟����ėO�BB��S}�#��V�k����4�b���`b*�Ov���O���r���Ԧ�L ",Y���&ۖ�����j�@��d&�b>�*�f���S�? �h#7��u��5(��� �°�0O��!Ĉ��~��|]���	ԟ��pd��Ny�m�`��W�ʁb��]�����<��cy2/uӆ��j�O���O�e�PiԜM�Ts��� ��׃=�����d�OT��3�Dx�z�Q��:�pT���֪@D���ub2a2e�̦�PN~�t������i�ޡ�����0Dy���Б~=�!�����I��d�Io�O�"M��M�*A8C+,\t���� J��.tӐ@��OD�d榉�?�;zA�A���:v�(ᄏߒB����?q���?ar���Mk�O�N�C��S�g�0�7#[��T�H��S.l�� &���'�2�'b"�'�b�'�ʄ3"K�Hh��Ч[�w�z�õ^���ٴ6�����?����O���{%�έp��I�p�>C}�LS��>���?�K>�|�2�F�|��Œ0�Z&u[&(V�V�2��4nZ剰"ۚ�h��O&�OP�IV�����O9� ����2*��z��?���?	��|r-O��oZ�`3`Y�ɱ+�����Nֈ��t+<[��I�Mی��>���?1��S���˥e_2a&6٢1A�,
�|ծӸ�M#�O�(��������d�w{�����D<w8�:n�c���p�'�r�'�B�'U��'?�@}Ht�%(+�<q��(uȠ��s��O��d�O\\n1sw���ޟ�ڴ����%�q��|�9;����i �xrbb�>ulz>� ��Kܦ��'	��A����]��Ix��[,g�5��`�	,~��I�g��'�I�@�Iȟ �I�}�z�k@9v"���(/_�����͟4�'�7�������8�Im����Np
9�r#GX��E������J}�	qӲ�l����S��Lli$���lMD���ߌ�,d�T
t�8$�uP���!Rb�S�ɨ+�03�`�Z���X:�2T�I����	ɟ�)�Cy�nlӺ����58a�l�.PX(�� ʊLo����O��nZH�G��I��M�Qc�(~?�8�$nد��[Vj
8_7��g��i��q��|=�=�e.����,O:(§�޹��!�󫄻Z��['?O���?���?��?�����)�lX�(W�o�dAz-��n�lZ�w䨠������^�ퟠ����3ШD] �5@�&�~H��J ��i��O�OV����il�O��~Y`B�yJ���̡R�$GA'J-���i�Z�OB��?)��G� 2�J�A ���eԪS� �����?����?�-On\o��e  ���L�	(p�8�Y7�Y�e����2�� (�|��?�"T�d�Iɟ�'������H�PmJ�gK�w쭃��.?��l�"˪��4��ON�]���?�V�K�_.�9 @�#0i���?����?���h����PWȕ�bO(GL�!��E=t��T���Y��HIy��i�T��^�贂`,۝(Y�U���1��I3�M�0�i]�7-��r�h7-#?�"��Pg��I�G9L1�� �>�2k�*��/��XsL>A-O��O���O����O ���(��9+��Rg*��J$(Sg%�<�5�i��8��'�R�'���yb��1W�&	8e�!B4�`'Ծ7�,�
�& s���&�b>�[w��Fid����l�B�����<k��;?��	$�$�7�䓟򄊁}nq�QÃ�=-�|��e3(���ON���O��4��˓(�f�HWb㟴gA�"�D�A0�q��F4BAcӶ�4A�O�in��M�ѿif��f�@�f^��b�@X�kBz�C���g�����a��[����	��99'h�;h�0��6�"w�V�p4O�$�O�D�Ov�d�OD�?)��lT�r"��>T$+1�_3@^���OR�����9��By�}Ӹ�O���P���O0X�`m����V�L���M�ĳ����3��������@1l0�Q����A�����o��q�Ld��'\5'�p�����'B��'Eb�����IV�J�☪c����'o�V���ݴ\{�Ub��?	���i[�?$�<���ւX.-IBmJ�r�����D�O�6mKc�|�%�2-/|�J��	
ɘ��FAMP�)S �,�-��D�ן [R�|rFҶ0#���MҤlXhz�
�!yQB�'���'����U��0ݴ�,����(�"�طC2F����G(�?��W)�����N}��'�V�qvI�e�����A��N�+&�'�,���f��DGdY�#��d�~BFJ*���;F�ؒ7��'k�<�*O����O����O��$�O�˧d�8e	�[��\�HeJ+~�:��i1��#��'��'��O�R'g���
�r2�1g�����"ȎS,���O�O1��4��z���"J�p=�֏�R� �P��B���I�h�x�)��'?��%�������'윈EM�1� "gC_̞��6�'���' �]����4�@����?y��{e��"sn��@'�ds����B<�F�>!���?QL>��������B#31x<S��t~��F<f6��G���ߘO%���	�_UB��
$�@�p�]����Q�ZQr�'���'���ݟYƉ93�ˡ`@9H�ժ�ARҟ��ڴh�D8��?ᐽi��O�N�wu���SM�"辸x����<I��?���0�
)c�4��$��_���R��ru
��D�o)�:7�
J�X��Ɖ0�$�<ͧ�?i��?���?�G�Zt�P@@ �<�\]CA���̦��bȚ؟��IΟ4$?���8fkvA���"Ep9qc�2����O��d�O�O1���2� ���c׍v���"ō/)g���ǎ�U�	_�(c�'���&�4�'�t�Ői�����E�i�F�'I��'�����tW�D�ݴ4L�l���#�����͐��������2�Uț��d�v}��'�"�'(Y�7+�7���6�݇	=�xt��g+�6���8P��F�������A��Dֳ@��ؔ�Z�E�mQe5Of��O��$�O���O��?��C@̏1UL=pu��>6
�9�*�ܟ��������4@��ͧ�?�»i��'�V���͒�r���$˕u��Y��|"�'��O�^ݑ��i��I�U�d#���o4r�r��:����#�Բb?�#�o�Isy�OJ�'��&2L��� T�;�\��	�B2�'�I�Mۄ�J�<���?�)�l�!!H�.@�#w�|(@ ��X	�O�l���M�g�xʟ�d�ߜ(�R\Q�ex ��&�L�K��Qjӕ2�i>�Z��'
d�'���t��	� m0�_���a���I�����ϟ|���b>!�'�P7��:Qy�Djv�
�sʼ��S�J������8p�4��'W��N)�V�@����Z+Z��a��`ӧI6��h��Цe�'�M�4�Z�?]����qV  �/�~e��ʀ�4�*)؂7Oʓ��=��X3l��CF��3)~-R�
�vn�f�tb�'�r�i����@]�H�6ʞ�0�i�6LP����%�b>u�̦-͓8D켒�^G��q�فj��͓x 4e0�ﾟ%��'E�'��I��hS�Q�|EZ�l��d*&�'�b�'�B[�z�4O-r�`��?����X	!Ԯ�9[�Y�AA<Y��Y+����>!��?)J>��ǒ7a:d�@-�V���F	n~Z0ۺ��V���Oɸ����j�b⛒R�X���h�z�D���ɺh=��'���' ��ɟ�ZЩ��v*���T�_#������t��4GP��'�26;�i�}����&�h���k��>MмH%,h�l�ش��օoӊ1��'h���-|2��J�����3U����HD��ũSFK�h��O���|B���?1���?���/�v�1ԈJ�C��CwC�?���(O��n7{���ğ<�	a�s�\�D18^LS��F��Y������dRʦ�xܴW���O�:A�Q`Q-�>P�ņ=~�����C(�	��O$�y�m ��?ipc7���<���_jҥ�C�C�=���$ؓ�?����?���?ͧ��������i��S��]ƽ���V}�����f��Iݴ��'1v�Z��f�f��-oگ]�9b��DZ,�sA�L�w�,�g���I�'���$I��?e�}��;e�ʽ�����7��Z�g� R�Γ�?���?����?i���O�A�����f�Ed��f�����'X�'�F7픐s��S��M�N>��b�!��"�fS���ӱE�=*�'��7M_֦�7a.�oD~B��+xbqkw.å[bi�ӥS�Z�2h�ƥ���`��|�U�D�	���ß���l�>�܃g@ˏE �,H��۟8��yyR�w�H ���O��d�O��Rt�'� g���rCG�`��	��8�Iv�)JVˍ5�N��6�T�g��Fe��e�|X��%��;X!��t��B�|�j�/m >d����Y�!�.�2���'�R�'����W��;ش}`��5�Ш~PB����&��iY5e՛��d���=�?�Q�,�ڴ y^�Z Kр@��*��C�
x��i`7M:9�7�+?1 �� T��.��+G��DPꥤ��y�´�(���y�X�X��韘�	�L�	��d�O޴��0��!g;�v�r)ae� k��7m���p�D�O��D;�9O�lz�!TD^ز�VJFIl�A��"�?ٴE�ɧ�'+��9i�4�y�Z�l媜)3��X�Lܭ�y�ʴ2ψ��I���'��i>e�	G~Z�j  1p[(�;���)K6}���|������'�r6�*`�˓�?�t�R)~4�`	�m���	�ʚ&��'�~˓�?�޴�'G̐H���^���pb���U��i�Ox��Q!�N1I�R �?���Od�[�c^iݱ@$A�q��!
���O��$�O&�d�OP�}���	�y�ćS�\�� #�/cX\@��jH��Gc剘�M���wt:6E]�c�yQa��i2����'��i>n7�O<7R7M5?�qٴ�P��ұD_�$&��ژ�� �af.�AL>1-O���Oz�$�O����O쉸C`
RR}�r��=6��m`�μ<9��i�4 x��'�"�'��O�R�,7�FeK��HB0���B�?}�$��?���S�'>���!p�ړ1�v�*�D�?TE@``Ʈ�M�R���@,<L�a��J~΢�P%�8���i�e����a"+"GU8]�f�	�t}�t�*0�:q�Ѣ`�����J�(�:�p1-�5h�1;��º_(.8y/�ǟ,Ζ�>R��j_?u���g�.�I0]�*�qTꜯSj�h���:l̼s�.�I����!�}1r!gD�pt��S�J=�	q_'^�)�� G$�\�@>$e����$�21`1eC#\�U�"�ON$�F����A�5s* ���4gx��q�:���2���i.�����,��YR�+�v ��E�(��a���l��CV�L�B6��<�����OB���O�Ģ`l�O�[`��#��Y���;W�}j�,B]}��'%2�'��0r��[��(�$��Br`���� '�:E	���$%�rYm�8$���I��J���gܓJ��
3@����j�+=u��n��4�Iay�L�Ib���?Q��RU�ަJ4d�[����\��\@è���'���'z�P�G�Ĥ?� PY2W(H�I�hʦ��m�����i��I
�J�s۴�?��y�'m�i�-��N�/������%?���)�
q���d�O��Cd�O^�O��>%y��ك#�NE� I]�l��4b�nӞ@�bD 馱���@��?);�O|�g��%1��2t��%ˑ�8a��h��i��T8���$�SǟLH�IОFK�=�2b#[߀�	B˛��M���?i�'_�}�a^�8�'��O�CEN1�N�p�J@(����i��'Ȇ��G	<���O0���O�Pa�S�kO����nޫ[!bT@ek\�q�^���`�O���?�H>��J��0�J��*��C7�� �J��'@�#��|2�'\"�'<��8ϴm�R�ńXŠp�A�_�u�8�diۤ��$�<9����?1����R��J� H���R�O�Z�< vhֹ���?	��?(Oj|���|���	�.����ː�Sf�1�c	��!�'��|��'�֢^��T�d�����ȅo��mRNJ�E���ğ���ן(�'��|�p��~r�d�X!iq��F��q��}�����i�|b�'�ҌX:qO���fd��,xl8 B&����M+���?�*ON=�q�|����y�'Jk T�@�	n��U.Ѿ~�1{��x��'����:.�O�S�`�T�@�i��_���:S�5&�6��<�����c�6��~������X#�ϕ�zw00S���2 <�V��M�/O���O:8'>��O6��;t��$:0j��L%����!ݛ���i�R�'C��O'FO�)�n^�A��ėdS2E�@�Yo�ƁmZ
n��-���8�'�����ڑ4ۘ@�-;.׬��$��2�o���I��w� Cyʟ��'a���B]!>���`�3`&��I"�I$r��9����'<��Ց�0HN�hb$-RV*���'!B�kfP��R���⟠��F�-�	צJ4L&	�����g��'�B�'2T��z�Z&T�~DѲeÙbX�4 .4~���YM<I���?�����O ��2K�b<@si�.y�:��4�����7-�Ot��?����?�-OTaÇ��|2A���7܈�0MޤB1�Px���x}��'���|�V�|R�IܟD�%iI @�xv��T0t�I0�U>��$�O"�d�O�˓"Ѱ���T�,_,�h�F�[s6����Q�b6��O��D�<���?�ˍ��?�I?9���7��$J��C!=�tGw�F���<���?{zUq+�����On��Ƹ��樏U�(��e�t� �xR�'b��'��y��X�C���Y:��Pe���T	0�( ]�������X��՟Ȕ'��tY���P��h8r��2�X�p�^�T�d7��O,�d�$0%f��)��j�<P;nR�yM��𤃓3����K�jHr�'��'���T��'j�*lq� �6a|3v!G���MAйi�<���c������d$���e�b��S��āY�nC˦���Ꞔ���P8�i���i=}"�P&З`�lD̉R1+N,q=�b��ȴ���'�?����?a��յe�L8[��	)Ά bch�~���'���I���>�/O4�$�<���cF�ŬpH��SC�ǭl羉�E������2;�����8��ş�IޟX�'� |B��̡�jś�TT��+�%�ꓤ�$�Ol��?���?9�'	xx�׮�2/� �"TC�^����$�O��D�O��(��qp�<�΁��	��6@�E��(΀}�R1鵱i��	Ɵ��'���'r*��y򭓭^0��RC�=\y�Yi-
�5\���?���?�*O�EJ�+�w�T�'_0�x�� @ s���Gh H��}���d�<1���?��[p\�ϓ��i2����I�ـ��[�:�Y�4�?	����d�����O<B�'3�4B�N"�i�A��%Hu�k�R�<����?����?�i��<1���?���]���`�ٗL���$q� ʓ} `�r�i[��'���O��Ӻ;�h�=
G�|�uM֬@,����Ԧ��	ޟ��A�m��	jy�I/��
A�K��;F,�'6�v��C�&6��O����ON��	D}r\���aO3>��(H4��S |m�Enޢ�M�"��<Q����9�S��S$����R��X�-sR���M����?!��m���6^���'�R�OxLj�Ň<#�,#te�z��ҡ�ih�W��R�@w���?q���?a�L�i�>�	b��#8��c�%��1_�&�'��h��k�>Y+O ���<Q����֌71�U���P6`���Ċh}Ҁ��yr�'���'A��'f�	@���a���Z�(,�󦗆 �������d�<)����D�O6���O�0�eڏ3�r�i�R�h�����_�$�O$�$�OV��O`��1A5�X�2�n�:I�x�����0��)�i����ȕ'�B�'��nZ1�yr.��8T�P�B�j�p�F�#$��7M�O0�$�O����<�CJ�AK�S���P��.[��l��`W�o��C���M����d�O���Od�i48O��禍r�7O*@a��X�ȀU"%�{�F�D�O�ʓ5o�ygR?��I�l�Ӆ?�"@E�.YWҩ��&Q��X�Ov�d�O2��4&����'�f �gӟ#�(�W�V� �fem�Ly�+O*"|,7��Ot�D�O��Pe}Zw\��&��;g���E�شGR$��4�?�C�B���?1,O��>����O9t���Y)���Gք�M+�LW� x���'�"�'���k�>�-Oh�yPA�^�L͂:7����������{���	Uy���O�8� ���!I��+vPc�4v������i��'����>�V듫��O����`��j` *~��u8ӈ�"6o�6-�O�-�D�S���'��'����J5��!��Bk�0l��`l���dÒK2l]�'�ޟ��'Zc�����NM�C��÷�۫|�Ұ3�OF�6OT���O����O��d�<14��/m���Ҁ����+�H����V�ؔ'h�^���Iϟ����T!0��gC
;6eh7�mXi���w���	Ɵ\��۟0��Ny�+́E�~��y��sG���Rz��*V�ץ!8"6-�<�����O*�D�O8�h63O�$�c@�����MR�3�H���æ���ߟ��Iܟ�'��=٦G�~z�x<Y଎�73���7�C�O��[��ij�W�������	���A�D�c��$�~�3&�H&(�n��|�	xyZW��� L|
���vͦ%��E:��^�<�Ͳ��R�
l��џ���͟��.�ҟ%�P�����g��9~���a�hQ o�\pm�|y�e)F^6MW��'��d* ?i"j��vꞍKS�ô9�
��aC�ɦI�����"B�&�t�����,m�ʄڱ�Si�$��6.�4k�v\P�07-�O����O~���f��ȟx��h�,%^%@�I�6Yj�P��J;�M���];�?�N>ً���'G��B5ׄdDH	%m��xxn�b��tӶ���O��*Y�$�&�L�I����eJ.�Pb�"c���n8��oZE�Qg�HqO|R��?1�'��L"*vP����.���c�iV���, ��b����`�i�-�qn!�z4XB�Ń~WI��J�>qb@�<�*O���Ox��R�f�8K�<�;��^L���VH[*l&�'� ���&�$���\1F)9�|��V�v��$dđ)Z���Wy"�'���DJ�P�S�;pP�:�A�
I a��ɋ�Z�듅?A����?I��Df�%Γ;(��AV��Cg��(t��W���Iӟ|��Vy������i"a��1p����ޡl?�Mx��Gͦ}�IJ�	ϟx��
����=Y�j5�����苞H�
�{Q��Ȧi���x�'��b5�:�)�O��i�+V�����{HQc!L�mլa$���	؟\�T(Bꟼ'�\�'O��,�Q�
��Α �!�/BIl�_y �Dp6�D��'���k'?�E��?g0%��G�i��)S�ڦU���4s�,��'���O��D�1:܌�����(�D�Q GEV���&9$�7��O�D�O&�����͟���"ޢ6�t�dH�i,,�2�!	��M��m̀�?�N>Q����'��,���hv ���%00A��p� �$�O���M���&��K�P'�
��4&C�Y$A���%*����'��	�>��L|���?����ԩSP��qr,21%�1*|~,��i�j�EΠO�i=�T#�2�M�!��<1$ ��R7���'�|�[�'��I�l�	ԟ��'� (����<$'NP�d	�=
��)%�B�XdHO�d*��?�6]�����Ǡv���Tm�J �y���?i��?i���?.O"�a���|$)T.~�zE��.Q��H�u}��'�ў����5�Q���\��У�h@�v�Z\xm��*	2ٰ�O&�D�O��<i�%��O��5��'^�h��)V[�\@8�5�d�z�=���V�݃����OxT,�FF��#S����BB�$H6M�O��D�OX��I,D�����O����O��	�
����55P��J��K{�E$�8�I�����n��dc��'R��]��/�(��2m֘E`�aoyyR"�hx�6��O���O��	�X}ZcMx��Ț$Q^�|:c)S�4�u�M<�������'����>�B�m�:A9!�;��B��]�QIƢ��0�	ҟ��	�?��'L�S.Z��Ӧ�*
&��ϟ�E�b�ܴpH���.[\�S�O\BK�e�n�hu�Ȼ	�a���Gؤ6m�O��D�O6X)�DԦi�IΟ ��ޟ��i����YW8�$:4hˠ0�֥ `A}���O ��3O����IJ
b�0g�TؒP	���B��A�Ɍ{�h�@�4�?a���?��H��t?���%;���1G�X<?���Cn}�b��y�T����ٟ��ҟt�I�>��8bu�	�o&X��l�)�t������MK���?���?1�Z?1�'}�Q�|.�hS����n���ؑA4�D��'��' ��'n�Q�$��G�����شBP����/G*.�&�
P�Ŵ�M�.O��$�<���?I��)�����-ՒO�&�C�.9ul�������	ȟH��ݟ��꟨)�*���M����?	�ě�?��l����b�Z�[V�UU���'B�'4��ǟT��c>���j?�L[�b(`S4Ş>c~�6&��)�I՟���ϟ�9.��M����?���RB�Mt�I���A(� �2ě��'��	ٟ�h�dk>y�����Mk
��B&@)4.�Ur ��q�����ğL�hN�M���?����
�'�?����\�A��,�!9���2.]=��	�� �������ny�O��'O�Ȱ2%��i1�6��'�h�n�@	��"�4�?1���?��'%��{yCF
fhMk�c��!� ���b�'v`7�,�$�OPʓ���Q!ӡb%�bQ��[ 퐢㗆g�.�Ɠ��-I�����a�*^RI���	Tp4���9��`��b8�oE�hH�sP+YM���P��<���.���T.�,��5H����i�݁�g��v���jdJ�4��Š��C��hQ``�]�L���-_p�Fdj���!mX�Z�4�C����n4�!�$�f�;� ��� u�I��Z�u���2���Ol���O��I8)����O
�SB�Z�� C�	��tlX�fD�M$^�T��R硇�{�Z�k���Oj�GJ!R�\3�$
K �D�ĦY�7	�0��D�
)P���F$rDmG~�ќ�?��U��i��#�"o$*l����W�N،�3��]6�^�M�f�:2S'�Hp�ȓw�rlx���8^,Q
�Nm�\�H��Ify��9.� ��?�,�^"����)t��T������똇\N���i5���d��\s��Y2˖�����O�S�^����H�� Y�-ʡ'���<�p�i�Pi���Y�<� �`M|�cI�CV<�;D�6BR����q�'̪���?���t��F#.��E.�<������
�yR�'���df]Y��5pV�
O�DHk���'i|\��_���E���DD~X�'����I�>����I�V����O�d�(�64XC��z�CBh�_r��H��T���ˢ�Jt��|:���v��y�VC�@@T�ⰣOq�$a(�*YZX�sgBѾ>U8tad����"�֬G�Ps�gC�%�Xy���qbb�z��'Mr����&�O��� b��Peܵ�`�������"O�����N1	���U-gN�c�	��HO�SZ�t��d�}�Rܻ�fעo�~m������R�O�3�v)��П�����Գ[w���'�jMsꁟ����� �81��J�O�D��486��b�������::r�=3��&?M��PcG%4\0���9x���!�%>^�s�՟%��l���'��j��Ae�"��@�F���'
�(�����=�f�T(^0�
E��Z����S�<�B���4;���r�<m�P	Inґ�"~Γ��kc��� ��q�&�8 �ȓ�88��)K�B��J96�������d�Ԭ;��d��2�z$�ȓF�3"��!I�4�`R�b�=��dk��1�CC,1O�|��E�
���P܎�h�h�j^Mb��ͷf�*��ȓ+�,�҅D8'��l����&��1�ȓ���Yc�F�Nz(qq�U|���}V��{���6XzQ r�JM6	��#�����HI �Z`gS���ȓ!#.T���e��@��?H����DCԹ�S&#�` ��>o�8\��N�}x�	�$R ��S��"{T���J����7B�l��U3PB�7o����_X��rǫ��Y3��jF�@h���h��L��%V����$�U&����2TgW�8����L��f�ȓ��Y!�BJ/�lj⠞*x��ȓ���B���$��{�Ĕ>n�dt�ȓ`�8�`�\�U58�3�⛞T)⩄� >xR����Np��p%�0+���/���Z/r��«�T/�m�ȓ�Ń!�FV$N�`3o�r�$��3<�Pjw�\?v��pD�E�<���A�+�vP��X�V��%�O~�<tA_��АېN�T�p�2�z�<QmISj�iE�����!���A�<)V��A��}r$Z�`o<���z�<�`���Y�̑
FH�?l�I;��Ey�<�TI�Y7���%�Ua�ʖ��o�<��VxD��T(�?�q�t��n�<aK�i���\>ODL�9�g�<��˙�#>D��	����G�a�<!���ݸa�EG�8R�8i��_�'�H �Q�4��OP,yspΔ�6��i�W����UZ�'w�����#�vLS�kH��f���'��<�5c��YKɧh���OH�%���	6�C����"O����D5D*�{�M��/b��4�>1w��.;W�˓l�R��aA�a��e��? Hه�	
V���
�^3�8HP�Y�Ԥ�=v��e�ē����v-֢r���aTbԱ?�D(F}rl�i�rj'�� 
-�JPy��P�Q�g��iQ�"O��S�ДNٲ��ɧI�J��O�T�M\�d@1O�>�rpJ
;%˖�طm�����fH-D������Ai\,)1T�Yt��A��7D����֍3*8�ҹo�حu�*D����8(BP��Q���I)`�5D��H�C�|X��/q���ȴc>D������#U��r���	{Ѻq��E>D�$
DgB�F�kw��]���x�K:D�$��(\{Wb9����bC�ԙv�;D��Jv��3[���s��aѪ|{a";D��ڄ��2q�P�Y�F�P^p��$�;D�4ÉSKZY)���)z�6X�CH9D� �%���'Ϭ����w�����a8D�x� E]�`J �B���:.T��"8D�P ���.I�l ���_; �q⦯(D�����|1a$nʚ)r��U�$D���c���J��aG�@�l8�?D�T8S/͹l^�j&�E�/ʜD1�<D�,�6M�K���c��ǎp(��&D�ps�Ě!@�:���8r���):D���!�MCl�(ӣk5C-J��Q,+D�l�E��nL놌��f�[��>D��h���[��� �/��m��ۀA;D�вKЊ6Bfls���/y�VU�!�8D������m8@	�&@�]O��Ib##D�d�S���Q�$A m��!t#D��qTBBEn�񶀞(�4��$ D�|��'��"��qj�엄��f�(D�t�poC:3�`��I"�:���1D����
V+_yt��	@���F(1D��*P��]��;�(�.[�0��-D��Q��LXs�	�a�u��H��H*D�8x%i���̚�(H2*Rx��,D��q��k�$�!�N�QS<�� +D�HP�͘
V�\JƊ��oE�ڶ,,D��8q�;]
��B��!�̹�!O(D�l�'J��7�x�XW N�-�ܸ+#�#D�Pj���'G��D8��͇B����i>D�83h�8$��E$˳,B��r4=D�\�������8פ�6�6D����` <-�\m��O=�pi�N/D�`rg@�y r,��GO��IR�//D�$�A
�A�:9�t���$���- D�t[f��}hi��m�!'sP���2D������2K5�(p�UWSpEɷ�5D�����7�N�"5H�QO$�Ȗf2D��Af��>�a��
�����*}�"5X��6�8.��?�` �B>`������Ҭ$�6#D�,�c��KZe�GK�${��0:�
�n�&�'촐��\��Ϙ'�������{18,����vGȡ;�' ���^#4������0pc�p�B P@ �4@��N)<F�3.��0=	��#V>����L�}��j\���ޏp��E�s䚥7�`����� y��ȁ�f
V��h)��ܙ���Ɠ4�B�RA�^�_�����U8��H�'Q~X���[/7!��0�)T�p�Q��t��P��@���f1��x�%\�lb�q��X�x�bf��4��� $N�J)������MPv��R���� ��B�S�Y$�'HHiWo«r\���N�o6p��N���fUS���G�
%L�[֪��wuV2�S4���VΌ�m�󄗰���yD��"Q�@X���_�8Y���
�f�*���J�G<����G@� _h�)�!%e��J�$ߖRZ���Oƀ���Q��тΛe�d!x]�� phH�v�^-�#��@	�҉�ئ�?��λ� hѠI�6#���I�8D�8�� ̹!#"�4|��o���@�4n��?A��P8F�x@N>� ��H��ΗfK������ ��C�'��J��ºm��:@L= *
�Z ��:Pߨ��@R�c� ��ȉE�����C�� I�I+��X"�l��m�ax�X27�zXJ��
���lH�)@�:>�#�O�&��K�*ТOpJ���O�92OÝJ*4�zr��9"��0���hj��B��P̔�UÎ��t��j�O�R�Y��Ȋ!�d��C�8����')ҭ�B� �s��*sAO<�<d;P�F,ay3)�v������S��?�F���y�CܭB6.�Qr���b����!Ƥ��O
غ�N�b��'bnxG%��o�D �CS�yJ��ԏ7ԛ���*D�x@�GX0�0=!Ṙy^�YB )Ȯs�~��fkUM?�6��:�q��/2Yl�S�t��-6Q|��Ŭ�-3hA�Uaʻ���#����U�"O,I�C��;3��0�C��?�vH`dɂ�y�@ ?�@ȓ��09�N��]�zi���.I,�"+�L2tE4w�ԁc�?%�����RxX�$�/&8�C��. ��]p6��<kb�I,n; �s��0Ks����Y'v��	I�P�5��/�����$˪o��D|��!J9��Z��<�e���yB�P7�Sg��*}ܼ��n��;t��qKP5l��c��[��0�bK��&cRز�Ks3���SFi��j6.�m[��33+�}�bC#��2FқVR�]@���S�F�X.�������D�;&z�#DlK�~�r�3L�f�$�a�D�O�!��v}r�b3n�,Mf�ݿ�FD��lϦJܘ��WEF��^����#5��<�2ʐ�,n�¶���)?��#�V^��ɞN��@4�xT0 .��?��i�/��/�왳ᒽ.���jSl�:FȢMDy�$�$ob�훷邝n��hWd�H��	/8ՐM�V�� �RrVgʢ��W�,�X�U#� '����$͇e.�B�M�<T����j�Uk�}Zr��
_�A��\,1.6�R��'R�4{�E��Q7j8�c�ƄM�"O���ʍ5/8p��#[�>�nl�@��q*�x�-��,M��������%��!}	>4q�䝄n�Pт�x�t�̐�V��ȐG�06d ����9%v��%�O������/�̈́�#�4l��(�G�%�ݩ<���R��߂E���i�A�
��(;D���PH����E$h��h3?1F�?|B-��$��G��h*A��c�A��/Ăk�{�'����<!�Kα)��-��e�3N��S2>��V�͒zڦ9�3�ԉ� 1���be"l��-Cr�0CTC!��Ɠ2Tx�	uC�_�����m*�}��FG`	pg�U|����+� �ص�lS;m�h!1����������4��MB,�S�&�jr�K@i�:%�a� Kѧ�"�ؑDvP�W��M2|E&���O!jpD�\m l2$��(*(�`�j�)�d� �F�t����"1O��&��N 88P0g�,X� ���.������jT�����M"Q\Ua���-����B�Z�X�%��E5z��G{�f��hn���7������V����+[T!�dM�>���e�m�����}�ў�ANC�O碅�aN�[���ah���s2! �7R��G�~���7�1LO΁!��Bqd���`��I��e��`�e5�5�2�G�VPL����'���RR+M�h|j��N��d���$0>,���&W�^�D��1O^�@�>R?b QT�ӂ|1�lp��$#|�8��d)"x��)h�˅)-[�0�c��:�p?�ҫg�l�+&�&}1��B�3a_(�x��Ɯ�i���p�'B����4��`b�M')�F���="1��s�"O�M�IԵh�6i�1��.�n����ɿ0S�iq%���d�#e�[�[�&��()������Dw��LjE�H�U���$��&��t��
$�DH���D�,�f��IH��͂���?>�f�{��	�f�;����T��O<ɉ6�[F� ��%�Jʘ��s��W%L���bA_�uF@�0��=m1��򢌻"k
+#�Z`˦��6hXJ�z��k2��06�'P��R��I�5�4Y UԠp�M	w��7G�5 ���SA�?E��w�
�QW�&� �`�3H�}j�'��%���J�ך|�V��Y=�?!���u�p���eU���$��e�'Y(�[�Ƌ��r���� ;�L��(��$�lۍl�άb�#]�l1�$rL��>��X�f$�6�Ҕ�Y`G������r�Ї+V1��I�G������4i���P�G�~���@)�O�IN���!BV㍡1�p�ե��>!�բ�f��&+�i��I�F$Z,h�dF�+2����T�២|λ�/ 2n8�Bf+ޝw݈�������˱.��s��]Ք|�e!�.���d�gA��QE�wb���ƄX���j'�S2������7�!��j���;M#p7D��ϋ�'�!��O�X�aJ'�	�z,欨V�E+/!�� �P��|��u�@��h���"O +t��3H�E� �
]#"O(P� �WkZ�2��0�l���"O�e86��$�ST���|M��1 "O��I]�*5<!���x2A[�"O~���h����,*�&I�ލ��)D�8��S�Y�&]:�	�^���T�&D�aCC�&<��aNۡP��%�5E%D�`���W���b�V#"{޽�D�"D��Kd�K=�6�Y�j�m}r��d+D����BD;Bo��J��<w">�K��*D�HPskӾ9�=���φ _"EE#D�\!��2GA��2�BK~��#5�3D�x$Z�R��R��L�U���4D����"M�zr�<��ȋF���d�,D�l��Έ1_�ӕ�ɉJ!��ӂ�=D�L�o�*:��ˣ �.њ�C�(D���g	��Z}�,��.��%(D��Ð���ε�$!�(4��]�*OEOC-[�|Sf_�<5@�"OF�F�9J�6mr����t�"O.y�!�H�`��JT����x u"O�Th�F�1��� �BׅW�F��"OH����u�ʈ��*��%�<1v"Ofp⫉)�6��3O�$Ȋ���"O���!�Oܜ�H
7h���#"O
=�1�1tI�غpgw��xS�'D���pɉ�`?d����+F���`�B D��B�˾ ���ɸiC�Ҷm0D��B�I�6J��ZP��D鰨���.D� x7�5@옔���P�z�+D���Ӯ�gm@)Z�(�*�n0��'D���cK�-;-x��U.�Sml���	1D�e� %�B*��D"53����0D�Dc�X,�гS
Ɵ6�����8D�ܛV6y���p �!J,�8� *6D�,���T-]��3�!Q�/�D��Ն2D��r�* � (p����4z��<D����,B[��UB�I�� �ѭ'D�(�e��L��{DC	���3 �%D���׃C0f�t��f&�d&t0���#D�88���8][N��C��e
��ai,D��[��Ьy$���!k���2d8D�����
5"��X�DT�V��:��2D�px���6b� �rS�n ���0D�Dh� ��*�Q@L�}��o0D�4�V���J�kӏ�r�\}���:D��ر���u�xB��3^�2�7D�h��`��!���M�<�$��%5D�4�*�0�As�)�8a���3D�� ��
�/�Dm�dn�`�ّ�J&D�`qv�9�9"�A�7�I�W!0D�8qAd���}�hU	x�}��,D���',�#�l���@�{����)D�8#�/%�r���D_�ay&1s!�<D��B��E*l�� HcB©F��Kc<D�tq�-�0,VY�6��P�h�S�=D���"i�q*6]�2�%�~���<D��DM��S�`'�аk�F���'.D���%����JŁA�YB.��ю7D�\um\�'�N�J�����5D��{���)�nĚ֣�k��RV�&D�|k�� >���ťO��(�Q6!&D�D�3� �t �kN$������1D�� �����ޯ�Nx�P�^�Hj��"O(q���8z�rz��ܛ!N���"Or0!�*�/,��HԌ�^�v���"O��	+j�@rPP
r�&)��"O�I����g>P��91xlXC"OꀍN[~Z�JT C���u��"O^���í0�h�Q�^�fN���!"Oh���O�4_K�l˜e��'"O��XE�D t,�%�C-��r�"O@ ���Z�t� n�=`oF�[3"O�
����Iܚ�,KV�
�z�"O�� A��4�u�*q$�y�"O�q�D�<r�Zu�FT~DYw"O2bc`B<v�X$;�IcȌ��"O�!���M/#Y�xi�f�5�Ȅ��"O���3���S��4�P&S�p����t"O�hإ��U�F�6�
�{Y"X`�"O(�pH3,�R@ZD��A�xű�"Ot}j�k���l�V�<rz�4f"Or�����z�-k�B����P�$"O %�Z��(р+�5Y�Ĥ��M\�y��_���|��O	�O��`ϐ�y�FT4O�����V�}Nj�c�����y"�� 2~q��jF�rN�B����yrm�`��%�D� ��m��M�
�y���5N������z4akSO���y��?N\|��IM�
�EXSbџ�y�BфM�v�*�����9����y����ig��O���r"+�y2�Y1s���KQ���M���y�m�;K��,�ⅣD�S:/��1+�'tq����!7ݬ�{F�!P�,�'=�̡�*:x����^!����'�t�ç3;W��$�"PF��'l��pQ�$Qw�Q�f��K��i��'�(a�$��B2)v�ԯC[�h��'+x{7��F�4�+�a��&��Y��'&6XC�gɄ�Rt�P4$mHMA�'�y[�)oe�8�Z1���@�'b����J�Z<�]A�����R���'E��K^��4ev�ӯH����'I� ��"� �E����
���'Ǝ]�Wd��*[���Wx4Mi�'��H�cnB*i��Qcʀ^����
�'-&$�BJ�/ �Ԁ,�Hc��
�'�r�#2�R�d�@X�A�<?�}�	�'���RiÈ�Ԭ1�:��:�'�Rp"
 >g�*Ax%�4����
�'�L+�)X3>v��*� Z<.��U3
�'����T��;����3��z�>x�'^�I֡]�w�ҭ�RKֺ^�����'-�e���S&l|>=eD�*p���'zҵ����%^\�a@W8'T 8	�'��U[�-�*��b4���N!q�'� ��&�L)/`$@�#B˦e/���'p8eiƀ��?t�m
�fCW�v�	�':�P�@�G�
�'i� x�� H	�'0|d�� �=�.���������'���;폣x���Rį\��`���' ��#6G�;0j
��C�BҒ9��'ް�P0�̲!A���"	����
�'�Z`��&I(4&]@@	V��	�'�ĩ�B��e��Y��%.N͚�'E\�u
�F��� A�< ���� l�k�CA�<�c5ό���)�"O,Q:!�͜~fn����_0j��Z�"O"�H1,$e�#�Λ]�T�r0"O )C�B�)��))�L�_����"OP}��\$Qd���-υoth��'z��HV*�Z�ț9,��tQ���Pu�C�I<Y��|;�n�1A��ɺ�
)��C�	3|:`��'χ�H�So��C�ɒ�p��@I'a�`��Cµ:��C�ɡ7/���@N&rMP�8F�ñ	R�B�I����l� �Ϣ�X��'�<,�V$�,%�*E  b'#7Ni�
�'��4���/.�@x����) ]J>a�4,�HѫP0<�k6'V%�,���v�i��
c�ݺ��`��M��KLbp��3`'�L�UhK�����������'E�u�`ڱzpL���
�,0I�N��lJ�5@�dQ,�J��'�i!�׈>F^������]�ȓX� i�UM��b9�@��D��K,�����a���K?��b�f�&hR��ȓ �NHkrS	v��,` �λI�NB�	�sPD���W�T�5(��7#t,B�Ʌ*R)��i�%u,��� ��B�	�&��R%ŗ .8̨�M0�B��x�2�k�C�30iޱ��' �c��B�I6S�2�z6I��eqdU�n�=*�B�I�1��|+P)�	,S~d��JT��B�I�4�*	����<rQD@�Ǌ����d�`P�-:D�fY8� �ML��sJ7D���riF�;��AI`�.���J�n5D�@#&) �ԝ����X��@���3D��3��T;N��BDՙ�&p��3D�Ly�K4C�a����"1D���A���X�;�4h��٠�#D���Rd�t�0T�W�l���'>D���0%ܖ>X�
�	\�Nu��E<D�t b��P�^,K���5d��8D��sP��J�q�I�f�8 Z�(�y҃�:��c�M��8F���y���Yfc�o,{@n	�y��w�<�e)O�mo^�����y��I�P��s���]� �A)ݻ�y2�88l��O/&���)4 D���'y�z���qa`E�5��id����?ѐy�E�xYVT*�1E��|Bp+6D���D�>)8��pS&X�=��<*d"6D� r�N]�7��Q��J&���&4D����U�)��j�!E�%լ`q�(1D�l��`ՖF��J�E	a݄�E+D�L�R-�#<R�L�B�Į ]��Sbc=D�j���<*�r�xb�h9���W�9D�0IW���(�04Z0�B�Uc|X�2D�`���Y|� r�F�	C�!�$	1D��&��-��4J�Ćq��cm.D��`��ի)��<���)^��U�H,D�@�E������K/f���(k%D�<J�n؉)!D��Cb[;i����b�!D��c#!<bo�Y3���N��At�?D�l��R�<��=I�GF2"zy��'D�$8׫��A?0͊�i�	l�@�Ǭ$D��B�(=A�wB@����	5D��*�Q�y6�K�K�ĘP)-D���E
*rH�a���O -�H��@%D�� LzE�N;(�T�3投o��͢�"O�s� � (�Z��ɫm�$Y��"O�%Z�G��$���2�	8q�R9��"O8�� π�2��E�1et��"O"q���1�:iɢC_��� �"OB�i�Jزs�p�uț>HR��"Oְ��Ɋ8[>�Ӥ�7s�^iS�"O���Fi=J��X#��Y���(�"O�h`#��6V<a��rV���"O��s��]�M4.X+�@�G�E�c"O���F��RA*1���W�!��"OT��1ϒ 6�zUa# �u�"O�y�4�0	 ������k���W"O2����$le� �7�D��PT"OPJ$�P((�paal�;I�xT��"O��a���ZC�#�$�)S���I "O�1�*>7�jU�2��)Cy�@�B"O�3Eݳ^�~I����!�X��"O`��ڻOZ�X��HV�o����"O�p�"��Vhy#'�A�O�d���"O�A¦��F�X�zB�Ŀ�|�c"O$�8�`ڲ`Zv@s�Q�YR*Hu"Oh-��{lx�3�ͨq"~\BB"O\h�JH�wA�p	�e��c����""O� eo��M�X�r�Ԃ>P�"O�|����j�땉�P(z�"O�E��=��`K&Ґ��"OB� V��g5R!�匓dZ�ĳ"OP�j�B�0�2\�cڅS�%��"Oܸ�s���|y�C�RJ<�"O��s�1�j'X66�`�1D�Ԃ�(-[RtD�W�p&��U�9D� �ؑ2�cG�5#F�Q�g";D�t;��
yf͹�`�+l>�Ѫg�6D�`Q!���e)��K�C�U ��9�K4D�L9QO�v�44�tC�,mV�	Ơ$D��Ip��
����#V��h��v=D��1��%���a�^f�+t	:D��Kq�W�#a��Հ��>慒e%7D��`�ԯJ6��P��d���F�4D��PĤ��6|$ZM[�I�Y��'D��q���&lo~��:a\(���)D����NޏV���@�	��Vر�4D��c!Ս}x�+�D�~)�.D��2PK��]��(�c��O�ލ-D�9��O�hv���v��]X�3P�&D�4�5\<A�p�{�J��G��p�P1D��ZF�ǬRp�e���*6�zUK/D��ba�U(	��m�Wj�!R<�q�K-D������0{����`%�3w��1�5�-D�5��e!x\�����ax��-D�h�3�H)�0�v�Æ`�"V*,D��(Q���V9�  D>L&=Q�c&D���U�àeP	i����,�D[0F#D��"�j)^�$�@��.<}f��, D��YU�٣0�ʅ��̓N(�2�>D��hr�Q�Q�DI�@"0Rn����:D��Y@�B'�s�09	��8D��A� ������3_1F�Vu:�(3D�0sE�P�V �	"&Ș���I�D2D��Q@K�<e���C;[w�};P�0D�DK��)4����L�s�*)�b0D�ذV��/nȽ��Q�T�"ъ(+D��çb���G�P#T��U�C�&D�� �P�c����G� �:أ�"OJ��މm��d���]v�Hi��"OV�E�	J`�h��ON�{�����"Op�� �D)���sS�Ԑ(�&Ļ�"Oh��%V?E��P;de�Q��C"Oृ�H \��P�q&5�:�ʓ"O$����/VM�D��c��h�S"O6iC&$T�NID�i0�ԏQ��X�	�'���b�]�J�Qb��W�_��
�'9��A�gO;:8��ދ��Y�'����c��+�m�b"��~�$Z�'���Mԋq���' L���
�'��h&E8��M�'J; �K
�'P��G�_�c��-�fJ��`@�L����=�J�.4DI��^ ��Ʌ�F����3s�B�ؗ�X[��8��'�lt2�!B�Sb��L} ���96�0c&ҧuP��!��QmK"D�,`��)w��F�H��(L8D�\�3�E�>8b���@ߐ"�Hڗ!!D�D@�Ǆ�B�X����V���d�)D��⦢�m�J�8P��Q�%�&�$D��Y�eA$f��t� �M�kO����4D��
!�ɵr��)	���,�b�)�-D�T����l��5cް!N��2�(D�$1#��-e>µ`'�F� D�g3D����h��Z�P�tŐ�kz�� &*0D���gωe>*�BCȍ�Qa�e�� D��@(W�C��L��+9v �q���>D�\�B�0v��d���D�P`Z�0D�xp�F�*T�8Qą֔>�e�-D�\�6C��C1����,I�� ��&d8D�lp����M��5��L�c��XY0A3D�����n�d��e�ʪhR����E;D� 0�`
���1	jܥ�X\i%�3D��Q���3a/ �h��]�B@aK<D�����A6�����Y8 CD�j��;D���d��`.����Y4
�b��6D���AНa0��IE�	(l-J�фf)D�x����h�@$ ң�	s�R =D�@YF��3\* �[�hE=Bb��b&�;D�<B�JV�,����n�H�d��I&D����8!��8"T�*����"D�x"�֑Mֆ�{�L����.D��'(f�P��B�&b`��,D���H��
P#jN_�v8�)D�<&��_�����	S�A��(#D� Ʉ#r���0��L�t:PX�&/D�����?�$Ջbˈ\���j2D��9�o	�_�Z(�^��� �N/D�l�@O�$Lz�XզݠMn����.D��ԁ�*<�])cb�1x�x��S�+D��h+�v���0�^;>���f7D������BÚ�Ca�]�<:��:á3D�4
�LH�G��8���-���ڡ�/D�\@�狴&��}[EA��8
� � �.D�� !�=(���{�C�$h
d@`�j)D������Pm�I��F�n���c�%D�(P�FQ�K@b�TA����Qc�#D�@�j���Ͱ�e�|���x�>D��bC�Ǔ@��I��I+��ؠ��;D�4�!dFɣ�G	._��49n:D�$����,���7fF?3+�(UL-D� �O# ����dQ�<b!�� ,|����c�"�� �[�<![�"O�<�b%��/ĆY�Ь��P�Q"O��	�'���� Ǧ��|���"O>��Aq �P�O��J�z�"O�X��>�uH5� |����"OU�`�Q���Q� ŤaeX���"OV� ���>�Js�ƁU]m�s"O�����4u�l�RwNK�qK�9�"O:���A�5S�����OJ�ɗ"O���Wk��7�b��UM�=|��"O&���@!N?
�"��R�)��K�"O�0�\�Uz`��@*/p���"O�I�5���-Xz=yP+03���#"Ox4�ǯӂhz�#����*̨�*OT�Q�@�B|y��K�����'﮹WN΂(\�m���O)AP��S�'&谱�M�z�z͢��J5�H8s�'�t ��*ً5+a�f �c�!!D��9!���W@JQ�š����;�O=D� kse�B��*���aF�qr3!D�r�\��4m�s�ط]8ty3�,D��3H�)Q��8�,ՠۜ]�H+D�D�A��*|�2'd,�@��B@)D��;�i�M�MI!(�D�x�"D��[F��T��Q�ԯ�Vu�m���+D�xk� ��	<ɓ$*��9����,*D�x"���&13��x�e^�r�l�s�*D����V!�d��6[	˔tK�D&D���R�f�P�$:/����o"D��RBo�,0^DArO�z�����;D����$'^��˕�>�x{��'|Oc���k^<t�i��b�k�tp)g
2D�����W
�~�S��(#�Z8p�5D����̍3ƆPbt�I���
��>D�����i��j�W�ve�v��<�.O����,V�I��͇g �:U"$!�������l�le`dX�kN;k!�d5l�¡d$��kDd���N�!��.W\K�"Ó*Bv�g�%oў��ቄtƪ��o�L�|��4���C��	t�rB���<� �HC"W�f�C�:`�H�7��j����k�P �C�I�FLn��UDKb��ly#ʉ�O�pC�	lNhpq��O:���*�AFS@lC�	r��*��u�D|��C#[�B䉆Q�t)y!���s�@�J����DB��q}���lȽ[�Pt����9�b��D/?�&h3*���0�	c�ȁ@��^H�<�I ���fɟ�����,A�IQ���OuTT�a`�6Px�� BQvCR���'f��:ՠ^�M/�8`H&pZ���'oHy�V�҄[�����a���'5�cW�T,���ǋV�����'ּC��V;� ��J��9l��h��?��yҮ�sk<B���:��@3
��yBb� أ�,�u�4]�S`��'gaz�!��(&�]z6.Ui��`�u	��y�-Ӌ!�v]�4� e�BL{���yDF0�X\HǇ2����(0�y��ޟ=��T�ń�/C~�s�Q!�yB�.4�DcjҎX�}���ޅ�hO��O��O���7�G�w�Ҽ��*_�W
���8D���H�"���

@��SRJ!D����ʈ�xTz���)�-�p;_�y
� 6Q&"�$6���f�QxI���"O����$UN���7*E ]ո�"O"���k�E�08{7G�.2K��'5�'�az��I;9q.%�"��+�BIX�LM�?��R�s��y��F�|p#F �U�X���HG�<idD��d��&�Y��A��I]k�<	�LO5|�H:��A�t�Q��K�e�<2��2+�pK�4#�]
��_�<�p�J/1x���Eѹ
*�`��DUu�<�vO�:�CB!�Q�6 ��Z�!�D^&M��lЎ���%�S��Z���=O6rCJ���8u	��M��5�"O$��!�)
�(ܒ4�\����r�"O�1CE�5�n|���:.8��"O�� ��	a�q��Ę�SB -�"O<�	U��.Yq��#�c�>F�flQ�"On9�c�ܱ7g��p�$'.�S�d�Ot��͎h�,ɹ�(�m�b����=~���U��\5�%��ɛ��J	�����1�^���c��B�,�@�D�}
�B�Iz��
��]�H�)�0ԗQT�C�I86hp�J�&K�e��(���C�IG�4c��"i!�� 1͑%~�,B�-��9�GlJ.c8��@���0�O����O��𤟬S�re�n�>~�Y@��<�!���]n�eȂ�Z� ��xR�~�!�$
�NӒL=&3z\@�%��G!�ül ���I7H풥��H/!���]b�DY�`C�R�x@�L��l%!�dϒ~�	j�*�>1���1����!���lt�Xv��5h��ĂG��IꟐ��c��S�e��b�*�F+],�ѣ�.=D�x#EȣY#V��`�+3���"gi<D�4Y��\�J�b����
5Pj^���O����S��{r&�W�xq)U�JXR��ۤ�y��:"*��0�+�A����W!�y��2}vIkCC�'5ٶ�y',���y�A^$-hV|r��8*ƌ(�fƔ*��-�O�$"qL�A �a�+d����"O:�� /�vʖ�a�\�)�ȴs��|��'6D��$ڋ	���Ӂ�޷ ax��'��p�7��VO��p� �E����ʓI��ȳqJT%u��T��C�"'`�Ն�>�q�r�$�������z��
/�dұ��1��q)v=dx��v�p�ME6M1�=�d��?�䄅ȓ�
%ab�L�b��:��O ��)��dl�Q��,T" �H�����ȓlҤe2�K�qP��Yul<`L�������Y���&��C�4����"C����*�u����4(�ȓh�P�Ԧ�y��MP�Z2���	O��ea�8)fdH�Mډ3/�����8�5�ђ;36��@+7����l{�bʣ7q��+GJ�'M��i�� �L��"p���ۓn=%�@���GȨ0򪁀L���{E��0"؞���_�E����s:*(�5.	,a�m��Io̓����࣐�[��dS�"�*g��E�?�ӓI��!�d�L��ʨs"N�;DB�ȓM��)�ԃ�?1��x������	\�m�,9u�ä()>z��P_�8��ȓ��Lf�O�N7@<�(K>�Q�ȓ{|:|j��D���)��.F���S�? ) �N�%\:�j�K�8MN(�V"O��  F���D�����>4�����'��d����I��C
m����g�;7!��rj��cȝ�l�> �'�30!�$��]�Z����ڜy��x&J��%L!��<w6$E�w35�|���"1�!�䞾l�p�1U�r�e�� �SV!��!�&��� ytp�1�Ј!�D�_0���� A�O�f9`�]*"��6O�!c���4i��h���\�����"O�������m��y
��$J��!c"O�c��)mx,@+%ڦ։�'"O�PR��Ih�(����-y.�"`"O��j��W4z�VX�D��.2���"O�)t��.�`Pig�ѪB�"OΡ�w���l����NƦ�q�'���6a��=�׬G�����k[�7�ў��ɓqĮ�6�Y8�\uaԮ3��B�71���xF/µd���QҮTel�B��:��|q�,֤B��ku-H�d�C䉄&~܀�1LV�,��=s��I�C��4(��y��5u��E��	�,}�B�	�ro�8[j� 'n�<"D��;�˓��<��O��p�jJ�]X~�r&u�@�"O��j��H+/�r=�D�_�&p�"O>���F�9+v �i�Ɲt�^T�E�'U!�U�+ttiH� �L�"��!���KFZl{�kLu6ȉ��,�+t!��Կ%��x�&�5Q��ܻ2쒳a	!��5F��a�˫zJ�����}��'2��~~���g��@#��*��#���y��ǧW�^��1���̴@8���yB�������b>x8���l�8�yrDѪc���d�ن9���)&���yR�G�U���W�#-v(H��G�;�y� l��đ�Q7#��A�d�B�yRd�	[�P�[���.�)�d��(�y�Q�2b�JB�ѯ9P�M��y��r�$�#���X�UC�BY�y��)e�n)h�ەg���&��y�Q;F����Ə�8Sȁ<�yr��`+��"S-L�|��\2S��yBBɾiJx�5�F4f@���2�§�y�E�e$�oK=P�F�s2�M$��.�O�l�u�P��2��T�44.�K1"O`���&V7�8�&���L����"O��0��ɾw�>PaS�Z�8^H�T"O
B��n��q�V-W�W*J�"O�ZF�ϧW|�����LV
`�`"O�T1�M�]J`�j��6��ђ�'�1Of�K#aAlyV88B��s�z��t�' �	M�hy%(�-W��͐r��O�<��h-D��A���+Q��]�poً~�"=Avo&D�x���
!K����U�¦Y�D�e�"D��C# �;�flPrg LI����'!D�$�lּk�2�qa,^�%Q�u`o=D�P�3!�:��(���]2a�ΩZ�a=D�$(%��y��%[!�H�@k;D��r�AΜ~�5 NسEW��2GJ;D�胂��CMva�����m%|�rg7D�,�Ӡ�!QRܡ���B�\�Y�rC�I�<�"lᑄ�8t���S�H�M�JC��,e�H�1�F�"	�0x�&D�%B9C䉵r�P̢���6-��m�TĦ;�B�)� ��fd�he�艵�\�Avp-r�"Ox%�f��Cd"���L�-� L�F"O���ïҩe�`r���4�N��p"O�10�I��2���}l�أ!"O�Ѣ�K��@~���BO�+Z
�`�"O�� ��;|�Եyb�:e0:��"Omy��C!`�P��CPJ���"O�y9��%�z0�b`J'��l�B"O��s�Öc\<8��Y��9��"OD��w�D�=,P��V�;-��Ac�"O@����ˆ�x1.��O{��"Oڼ��dJ�d����m	�pzyA�"O�X�%� 5��0�*}�G/xY�ȓO��Y���0�L�ɤ��nI�i��	��IR~�Fj����$K&4�6�[�S�y�1h��Ԑ�,G8�����y�lҜ$a~���x�|�@=�y�cIH���(�%��t�l]S �9�y�ː
Q����S�@�8�����y��]�^~>psTk��38ш�aO4�y�Ҏ�0��J�*$�X��5�9��=����D��rc<����/3�)p��'Pp!�d��бD�=T��6��^V!�����z����{�& � 	p8!�D�]�X5	�d�������7�!�Z�Y�����Q&�H����9X!�d1_0!�P���WA����HMU!�bF���(��4�t�tGŉ6\!��Q�ȉW���ۆF�"O@���C$Ѽ��N�g��iˢ�� R'��D>�	ϟ@F|BB[����`	�0}�^�)&3�y�S�%����y��lZBg��y��R�Yq���:X.-���%�yR�S�G���rFI&|D��� �y�Z���F��VTM��g���y⬆�,�� o�+���P�I��y�i\�j 4��Q�U����?)�r�'��y©G����dҷX�Q��<D�l�c�� }�2������r���3��<D����a��.��T��0aV�D0�:D�l�!�DoP=�Ex؈� �7D�h�H�^��e�!1�����(�O�=E�$+].M|�b&��r򼼐�n��%�������4� }�����I�@w���d�-D�4˴�"���;C�F�IXmP�,D���s������oF6i��1���'D�4�����v�R�b�-h��YcH1D��B��Q9v�
��!��
`#�m[��,D��a��moh�-�s�u9���O^�=E��n��D���"�;��-0E�'�a|2���#��]�	.������y���!Ar%�2mI�yfN ����y��/ pi�S�Rs�6��� ć�y�&��T�&�Pa�؀pJ�L��%V.�y�`���=bA��Z��� F���y�ic�|�rd�>f�.� ϝ0�y҄@/�� `v	�B����
���0>�6�[�Y�~E�C`K�4��=�$��o�<aD-]�X���(y4�b�ǐh�<���W"}�r@��D6�,�K�a�<qa�٘ptD����ɇ ����T�<	��{����Gˎ?���2+Wg�<q�nO�[b�H�*���d�#����F{ʟ�b��S���Ls,d�� y��!%?D�� ���3�E��"�9�`� ��RT"O� ���۬VP��B���R��A�"O��kb̀7/9�ܐ��VR�TxJ�"OT�`���#Z�ژ;��ۮ����"O�����R*�T���`��[k�p��"O������.�*0�ѯQ��@Q�Ic�Iܟ@�O�Lrt-K$:I@��Zgʶ�;�'9FI;�bL�NT�
���W*8�ҍ��=O�x�-^�6T$!��
̈+uT9B�"O��H�ԉnR~u{o]�B���"OV}�ª'8FD���(�2�xT3�"OF��uP�
�݋E�T�>��l�B"OD���"C��a4ɇ�-P,00��D�O ��)��7U 2$+��u��2��9!���Wd� p5o־tX���9^$!��f��,��n�|M,���N;S!�dO i
�- ��%LR-�fC�+!�dd���㘸(]|9c !�D�2���gf��Vw�A@ >Lh!�D_g��Q��{c�0�aǓ��O�=��
,Y�J�C�P`4Yp0l)�"O�$Bf!D�Yb���S��5mI��"O��p4�N�z	ČI4E�AO"u��"O|�U�N!������e@TI��"O���F�P�$�c@ɓK�,�ɂ"OX)0�D*fg,��^��!�"�!�S�~�z�Cq���<�6Y��N֩lS!�D\ D=�p����j�dD���/45�}��'=�C�:602�X1(X)krN��|%��j��<�2.���؆�f� ,�d�$D�$Kw�%���T	/V��� �!0D��Wh@4m;������d�v��/D���'�Μn�����>0yl�R�,D��Be�]7`��yb��W�33lѤ6D��qBկ:�`���F�T�2�OT�d�OB��g
.8��DC����G2x)J��O�B�ɔ A��`��:�<�ӌU�=� C�	AhhI���Z@�XA�_�X� C�Ɉ~+V���DI��(�����B�	%a� 3��̀'M�;����B䉬�&��	D��0���({�TC�	#���"�L3&�8�G 2<���O&�-��\���@�,F��`N,�������>��'L����n�w'��;�k\;Hn���'^n	�w��"m����⎎ED�l��'bн�w�kN|԰p���A4>\K�'K̽�rc^�!�Z	�gl��:�l��'� , !�
���\B��H]oȅ�'T^�z���@]���P��x���?ɞ'�P�KB�E}���s���W�t�����ϓq��DX��D�&ڈd�գ��RQ�ȓh�8V�0M�PD�B��LLI�G"O~��%R�$$�,K�ƅ <���"O��
��6X%P����/ �1�b"O�����y�01s�B��N#��'��ɦcO�k4��B ��P
�ds�M:��M��� �L>w疱P@��{y���Ā84�tPB���\͢A$*6�ҷEBq�<��0�6uJ@̀e�ldr&��j�<1���*��%�a&� ��x�%�k�<���U�y
%�a�֔\�����`�<��JM�m	r�kS�*a����T�<Ia�+��Xr�;O��H�i�Py�U�����RM�FL=P�����33<�O��=�}� V0C��^�+�t��lȁ2P!1"O٪�Lݲ,f(X�L�8�b"O��j� �Dw:9��$]��x�@�"O
�0�?����#����#"Oz���Ȩ�
dc��hN�4"O&��UG��چR�'ߊy�pyi�|"�'MJ�PQ���o��Y��j��x	�'B
d����[C��6d��!"Ol(`Q�L	"��	�UB�`#P�""On��g,1z��ª� � u"O
)�N�����1C҂ :<(a"OD]9f�Y5w����S,(��a"O<�`�(C.+\R4���t!�j�"O=Q��� V;�H����IAp�@U"O��1hXQqPtɲ �5nͰ��C"O��9���F��@A%�"�҈��"O������/�@�D��H'��[D"OLM�Sn]4����b� �Er�"O��8���$T�"�p�m��Q)�"O�Dkt;,i�'$(��"W�'��	�<�N���Y��e B瞷O��C�I�N�
E�]�:�j�c@��V��C�	,3qD���j3��T�Uk��<B�	"cx�8Kc��QFB����"+#B�	ql���'�&:�>E8�	Z�y%B��{O��!&k۷WVЕ����>cB�I�K����.QA�Uk7���Jyϓ�?��yJ�;1��ie�á%Td�#4�A��y2��K
���H*,�P1�H���yrɅx	��E � E2rA��y,�?_��mBe��aAh��y���/w�4ВԁV�M4`���O���yBIָ2�N�Ju&ŗC`r-��ڑ�yRlM��J�i��@���d!�&��>�O8uaq�L��r��F��N|J-��"O�����H�����9`X<�%"O���H�)�r�*`8("�-B�"O�9�W�Q-
(̱��G�KplA[�"O���G�&+rP�q+ R�p��"O������b8�6K�4C>�+""O�Ȼo��t���K�)�i?-��"OV WF93*�y���W"�*�@�"OМ���(r���[!OxJ��$"OHy�Ĝ"H����!.q���p"O�5xn�)yL\h�2m�3n���"O���㗢l��1�ҩ�TFt� "O!�!�N�L�X�'	UE�0�R"O2�k�B�I�DXWFW76�hH�'X�����8B -
ӏ^���ͺ�'���h"T'�zlc�i_�5.#�'Ő݋�c�7F��T�Q#͡3���'�(�풺;�ႁ�@3�va�'*XZP+�e3f���ͧ+6̚�'���v�֗G��h�M�8�<ؐ�'�\�֌ �r�b����4\�e)�'
�b�L֑a��*�˕-��)�'&�)ce�������C�('+��j	�'l0�Q��
�zJJi�4�^$�`-`	�'c���Ԍ�,HR��8qA�}q���'4D|@R�K]��ī��C�x���j�'����L��M�X�I�āC�<I��'�J�S%P�/{<�[uI9q����'��bn�.��a�M�2�4pR�':���敋yWDi��D�W�#��� � ������m�-\�9�A"O.Y�Ў�pqZ$Z���w� ]�"O2���ɏ�bk�E{�H�&�.ɘ"O���G$�m���aW��vخ�p�"O�z�M�cH>��(K+44@��"O�����G�Q� �1�Ҡ*y� ��"O8�Q���i�����t��"O��)��\�L+h�Z Z9!����"O�������t \�1#�ԝ4}��Z�"O~i	���@x�3Ų[
��"O�` �f�U��e�߼+�iW"OIz���-4[ �00�|M
5"O��R�@A0AOj1{'��rk�՛�"O���G��"���������8b"Ov! V�ɉj��magd#}<y��"O�l#\1
()GML-V@E��"O����"�Z��0�4�i�"O&�ٖL6�����M�4v�Q��"O�[!e�wD	(���	��|�S"O�rU��)�������4�b5�B"OhT�&��H�F)R�;���8u"O��5@FT���@���]_���"O��2�Ǖ7E�8���}3S"OLm�s!Ɩp����QHae`]�#"O�@Z�GQ�5���%�a�H���"O����M���(���K]�zT"OJi��I�V�4��	�.�(�QC"O�d��GB�C���@�:y�\�Q"O���`o�:qcl��n	IM�L�"OTEK��'r|��x�,Wt]C�"O�y�AIT�}�Ҋў��� t"O���4j�{M�=�	�E�u�v"O���pǒ=��%�TǕ;S'ּS"O�l�1j��x���VeF
ڭ+F"O@��c,N7>��0����S�$���"O��1,M�p�I�B�ڹ�Ƙ��"O�Y�Fn�9j�lH��2�~���"O��Xf*�"$�J$xR��	I����u���1+ٟ1�J�C��܇;�¬G��'Y>�S2G�;g�"@\�|PY{�e!ړ�0|�A��X�09J@ X�A���Z��~�<�,��_.�(Dl�;)&PʂDX}�<	�ߖai&��@�?#�lqPfͅy�<Q��
�N��y�L�:W�0(A�Tt�<iU(ͥ\J�A_9��Y+'�r�<�.�02�z� �)ʊMJMc�^Wx� Dx��B��)��cިA�|8�RI(�yr�M��L�At�K�;C�0�a%���y��[��4��ֆY�8��T1��ˡ�y�ԿAǒ]Af�=+�������y�"�bj$�W	ˁ.Nb��6�y��Pk��q�VS��8���y�;9�༛#��7ER�`�G\���O��$*§J��
.Ϝp��+��U�?��I<�i�����Dl���JgG�ȓ ��R��4K���Ǽ �t���t!2�JR���~�%ꏐsS�,�ȓ[��)�A�$1�\��N��qq�ԅȓ$Z08@v)QE�
n����ȓI�Pp8�Ő�#��)��&Ȕ�E{��O]�eϺJ��P�T�C&�@{*O���B�2�\�O��,r���`惕Ei!��r��'�Z�&-�#��L!�=c�LS�	�3�\�'�Lk`!�� *d�g�R�86ڹa��M�9)|)�"OH B��J%D��9��c�(l�r�"O��C��L1s�
i�����R<Q"O��G%�z�í>$y�"Ov�y3@Ř,&xxq�I�f��(�5"OF���ݑC�TI�c�)��	�P"Ov�zR��=t�h�F�3L�T��c"ON�c�B�g�漉�c� p�J0��"OT-PI_T"����I�T�M�A"O�E�OK�U�&e�v�0oʅ["O��ȵ��C�Hpv'ɮ~�>Y�R"O��	�A�o� �� ���p@�G"OD�hPA�>��fQQL��E"O8y��ôs
��[�#�	(�61J`"Oh�pf��/�tx�R��>��ժ�"O�,:�	��NЪ��Q�^mz��E"O��
�  �<C�����M�2F$�"O���C�^+`W��D�w뎴)�"OniR�S�������85�`�"O�\@�"<�e0�"���N��"O:�!�$LL!&!W5���hB"O� �*h�X��
E��IRr"O�����D1|�H�/��|����"O��;Q��xj��B� S�"OX]kg���Q��;V����"O�`��G�t�(r��	\�d�k�"O��F	rip�h
[<���"O�|Iq�
�$>��[0nM�^���"O�ؒ��K�I4lM���΍��!"O^�c�Mqm",���G�\��\�S"O*`! ��:G�+㌇�`�a�5"O"��R�� �AE⍸-	~�aV"Or�f�[)E��P�Q;,��(�"Oh���$J�rp�y� �F�l�Flp#"OJ�넃C�{Ͼ�8�ʐ1�&u�""O*�� D�	X�0�*�u���1"O�r��@:Go�ːjL�Nu�I�w"O<4���I 5#sf�ӡ2s��s�"O�Ŭ�=��1!)�*\(-�5"O��1ׅاN�b��0�B��!@"O��x�'�]�L8�Gx�Ti�"O&YG<N�Q��,yq���0"O(DY��2��I�D�]v ��	�'�>����N;7!LZk3�ٜ�y)�n�p�d聂�$@$+_�y��ͷ+fp�;�(Td�93�Q��y�Ö��4P��	�FBL�bh���y҈�8?�:�i���@NЙӆȎ*�y"�,%x���>�F4у)�yB�[@�{s�#l�m�s%��y��gx�MB�*1��P����yb��B|�yyQF�!�P,�E&�4�y��ٔcV$tzP��;~ɢ���y�oįK8Ų#�X��*V<�yBΘ�#��W
�@��BF�y2�Z:"ٸU��$2�,���G��yb�H=�Z�ccc�>����)4�|k��,.rf�Y����;>b}ˤm;D����V1p��e�ЁZ�_6$ R�8D�<;e��
���ue�+����,7D���v�m�R5���	����h3D�����V�^�"L��b�J��5��*%D��Ir��]qCj��?�ʥ��/D�l��	6�*�`��iL�r�j)D�� ���"�R�?�I�d��2 ���B�"Oʅ"� ����0cD�$ii\���"O8���A�aў5Ó�:�ᱲ"O�(0��.�ɆC��+L�1j2"O|�2�ʈ(y떅[���<s�N�R""O���ub�~H �������Y��"O�Lٓ#Z;z�)�3���B�(ʔ"O��'�Q�.(a����i͈1�E"O<%��a��!H�����K�bD�"O!ˢ탇~����4
:B���"OH��R��Q�&���xs"O��j��]&[v���M.x�N��f"O�	�r�?�b�	�,Ƒj�(��"O�؃Γ�T܌���Ꚋl�
�U"O(����F@���*��S�F��"O�HS�!�kH2);�H���� �2"O>D�l
�BP|��$.�z�Rp�v"O�"si��sPXA��lP�8�{�"O�)�	C�E����ާǤ=��"O0e���6g��gK��Q"On�;A�$k:n(Hƣ��%1l��"O�X���HC,�TZ0��3	5�)w"OF4c��"G.4 cM��z�xd"Ol���L�m�ꄠc�A33{��"O*�ڡ�ؘ	$\@92�J���Bs"O.$�JZ<7�\���k[7��bV"O0�( A3� �8a͏r��3"O8 �m�<Y�ݻ�@�%!�����"O���Ê� r�	��mX�rQV"O��򷃑<+Z:$��	uA�=�S"O�ᢡ�X�f(*sH�5)$��f"O��X�D�#;��Qe)�8���"O�AR3��F�u��-�>m��M��"O@ #!Q7ꠁP����w5>ҥ"Or�0sgU�Tڐ�S�)cTX}P6"O�%�����@L��ѐ�>y8��1�"O��s�!!�ԛ��G9DL2٨�"O֭��M,{��Ec�(?Jv��"Ox}�s�� !N�<����;E|��"O�ت"�ǰh�JA"�.Y'	A|�!R"O�� qeJLq���E;���"O���噓��!C/�Q0��c"O��Q�f�>j�ibGZ�`ߘɢc"O�E*�ĕH��3��ޠ.����"O�� �	Rt��a��*�&��a�"O��i�!	f�f ��,����"OZ�Q"Z�Sv
15�8'x�"�"OX8�H8L�N��㥆�3*��V"O��z�d[0&����Ą~��8"O�U*`�E��8X��E���`"OT�$IZ w�ε1���Pq!"O&0�u"��C[T�s��-C�v��P"O\��0�ͱ>��rC�<#Pn���"O>�����@u�1;�G��N�����"O��T�y��i⧨D�����"O���F�$5����UH �({�5��"O6�+5�i�"�k��G�[p;�"O��x/؛;�T�b���l���"O�r��F_�:D�S�O�Fh3"O�	Ɇ3쪍�SM\"8�>�"O����ĕ/�����)�	�ؼ�"OR�B�ʙ R��<	��G(/~r��@"O� aA$t�\�s��y$D�"O��3eS4 �yf�,q�%k�"O� 8kACE'3���X�@ :X���"OH�{��й`�~�p�ɖ"��}��"O���R W�q��/����p�"O�;��K����ܒHb�q��"Ot1W�%��X�Ώ/>\��i�"O��i�NR�@d���,g�L}�P"O�5�gM��!�)�o��V�~��G"OʩR3��EȨl��g�"Z`^� �"O�	�]RX	�ܝM����b]��yr�΢E7~�d��;V���1�P��yMǖ9��)�%|�����V��yB��8ym��%.t��$�y��[2d�Ȁ�μ$��a��?�y��%O�X�W�(e�x����y�D/o��@QJ&Np� R���yR��z�Bܻ��MJ=��)T���y�,W�a���@@���V�T'K��yR�"y
p�h� E�[�PtY"ٸ�yBL[�sP0�%O�8O��`�᠔�yA��ez���f��F�B�@�'�y��Q5V�J��*D����ތ�y2�H
kh���Wb:5|����#�yeT'rȉ����3R�1`���y�#ǡse�\B��Z�,Ϥ���B��y���5;@LtѲS�&y�јV�G��y2P�M(���H-g=�����PyR)7%���l�SE�� x�<�Â����$��<2����!XO�<Q�΍~����l�����b�Q�<yĦ�0qn�"7%�s�\��3F�O�<��!T�9W��іCX"�l�EE�a�<�a	�^�1�%�[RZT�h�'H[�<�A��'�N`2��U�TN(=��V�<aA��
�~q�$��##����mP�<9E�:wD�ks�_8x�B]���GP�<YE ]%
�F�����7z�JL��Kc�<��B	�.�btYR�D6r=��YF�b�<�TdE:Հ�`ԣ2 c|*���U�<!��U�Ip�R�A(�d
'@Jj�<�EB�L(B)J%k�`�`�l�<��� �MSt5�W�!Cg|����i�<1�\<Aؽ!	B5`{� �c��<q �ļq1!�		�Y�XK�a�u�<�o�/$Ej1���R�X�� KԎYW�<�	+GR�)�wM�Q�<�w�ݠ��y��C���b)�K�<�w��N�����������lNI�<�hLX����Գ7��QRD	�F�<!V��B�*y����/Z����kP@�<�p��%d}��	�t�\ �Vl@r�<���W�k�zPCGS�=K��aJb�<�r��-(�;������W�<����%1n`(�J�������V�<i◀]K
�*�k\�J3����^P�<1de S�I2��,rS��a�Yv�<9�W�W��X1�H�'b�=���y�<)�$�BBPǉ�n1���I�v�<QdJ�95P�sn��]�tI�h�<Ad��x�y2���=e��1���@c�<Y@�/p�z��%�F�tlĝB���F�<����>.�x�.�n0���U�<ᑦ�]���V�|�lk�G}�<q��#Kq,`:���u���T�LS�<�P��0��p�ЇCv�}�u@DO�<� �dy�B��i�>d�7ӠF�hIS"O���1�|��-2���"OJ]��`�	)�6 ��L�?X�TkF"OKѾ&Xma��2o傰�O��y��!R�I��`���A	�y�&�w����D͖g	�lń�y2��S��yK�J��0��F�y����t�֑��'!�eq�)�*�yB��,�b���0qh�=r�ȩ�yRe�$2!y%&�,m�����y��J%� S���8QX�����y�3if2��!W�*��i$N��ynViK��ban�)"Q��TG�"�y��
�!}�t� ���"��
�yR�7 �(��h��H<SH	>�y"J �ƨ��*�~�x���,�y�F[ ]��}�d��E��܋����yR�X=^H ��!ƚ89����2 5�yB�����%�aE�m(�	��y�cK��z����R��8�����y���<AN�*���K`R��siF�y"ϭn��P���'Js�i ��E�y��X�h�`k�����'��5�y"�ݝP$�Ŝ���*,�yr�	lMޅI��"/����J��y��NN��z���*tw\��`���y"��OvxX�*�s9�Х�;�y*�f���BE�zp~�"N���y�,_��Y�7��H�������y�b�4#~B���k�$U/|]c���y�e�v��[����S�8��QkL��y"�׃G��hEl��T�4-�e���y7?�p��� уL�8���	��y"�[��z`�S�>B���m�yg��KR�I;r�=%�ر������y��Sz2�@�%�"W: �d��y�͑!�rp�`�+�e��Ǔ7�yb�A�aF8�i#+ߘ'�Z�Q!W+�y���uCnh�rɥ!�x40 gJ�y�l���)9��
!� e��N̳�y�855x`���*����I��y��'k'�M�E� ���Dl�y���h�p�*�X��
E��iG��y.�&Q!vɅ�t�a���yB�Ea%raQ!S���Q�ҭ�yҡؖ&�b���3G�hp@�1�y�b:�� B��6NP\p�A�3�yBh�Y��5�r�|������y�ω(f�t����dX�p���H��yB+շO86h��DſUD�1�AP��y�^� �A`C�]N��X��D��y"%��)u0@��IU	:u�P�@��y�kމH=��f/��1���"H��yҮ�1<����R���-{��z���"�y�X<E�=!e 9�
��q�ת�y�X�w������dm�� ��B��Ts�IО �A(��C��B�	�]�����d�!G��)&w��B�I+$���P�3�c��6pB�ɔg�a"�D�#�l�� ��-4��C�I l�H��!鑥hF��UO�~'PC��L�yBA�>]����5� ,�LC�I�c|X�����0�8���	�JC�I� ��i0t:g(ȫ����P10C�)� Lݢ��
�_$ ��N�1U��y�!"O HRKԈ#�`y��u��ň�"O���j�*��=��mc� ��"Oy��! B��� �-�<9Ǵe�a"Ou��j��m����S�u��"O����
Z�V�8���E�0�!)�"O��9!o�+z8r�����Y��Z"O܅3�n�3���U�o���c�"O�}�4Ԉ;D�2T�!����"O x�m�F�M�b�!֦�"O|�S˚�h�]ї	F�:��h�"O40z"k�?tj,���&���e�'щ'��T��w1f �r%M0im�x�M����I�v�,*v�����e�V�a����{��A�ب0� )���ַ�8Q v.-|O�c� ��!�~�A�#ԇ1[(�9e�(��ȟ4 [#� �B�	��F�&����b�I�:}�>m��D0��¤i�<]��L)�F���E{��)6b��9���9����ѦեC'�y��1M`1�#�=-��p���3jb������@�X$V�J����n��1?A�C\6�qS�L�-XAT)"&����B1@tK�ڗ��-	��x�n�ȓ='������<9���P'�kz^������a!���H��e�V�U��ՇȓWD�i�HCʼ����
".7�O�O*0��
k�ȁB ���rGx "O�i���k^�j�A�1O%��G�'E��-�ĀfJX-6��0�DH*{!�C��	D�P)�R��V��P�n��d0,#>���ƻl����fE�6H�]���T�!��O���#)J)n	�A�u�>dƄ���"O� ����" �R98��GM����'�>���.��n�P���6�y��,<��p<�$L�u�p`fJ�	�2��#��r�ɕL�{҂�3p[r����ԧ���#"¡�M��'��;��%T�8�Cʉ2��1�'�ў"~��"��2aׄ\N���"�Li�'�?�P��{v��R�fS������0D�|���2J�J$[ԃ��M=���m9<O�"<��!�,�Pq�1F�\�����l�<�"�"U���4�2�� g�*p��	v��M�?i����<�N�{�,^�� �sf�*P�!��j�J:�R�u����H�~�'�a|�.#A�a�5N� @�ҕ���Px��i��ɗ�(B��Io�k����'C���iC<&����sd�.W�-��(O<�s�����q3'�R�!	�� "O�	q���V�(ysR'�; P`s�"OvG��:Fe��5&�
���W"O���&�Y40X��&@6ۀ;"Oy{�֢Q:����P�tQ"O8�+'��u0�j���B��}KQ"O\Yjw�M
-S��5mB�D�6�R��;\O� �n�p�����i��q��"O�ej0J�V��y��,'w�I0�"Oz=���)�A;A�޳bl�(j"O��q� N?�,H۵(���"O����g26�(����2�$<��"O차�\?o��|2W�E.;ٱ�"O9���]�{���� ^/Q$>�S"O��0Q�Q�<mh���]�ʰ�"O@���>��ԪW�֞}�2}��"O�9�SJ
����mG�^���"O� b��g
��J1���Yv.1�"O��3f�Ӛ0t��b��O�<o�K"O��`$���g�pP�Q��J�$��"O�m��H�p���G�����w�'�Q��u��u^b�1�O
�*>�(	ׂ8D� 1����|���G���Aq�)D��Ye��_U�\B �+/����f,D� #�	�����Ó�'Rw�Ik7cn�ڣ=E�ܴP"p;���aÊ��K_;mb"`��e�j�#G��0q\XakCI��8(:1���?!��6#�r-9��4+ zm1SM[e�<��'��poba� ��g��`p�
K�<Aw�]��A��.�ZY��lI�<Q`��!�|�"�)AJ����F�<��;5�^��â�?L��9�G@�<�샐L(�u�'/.�%b�o�C�<�n�V�u��	;#vy����c}�)�'*G��`�+�Pa,����L��ȓb;a�&���3����EƗ丐l�;��$!�O��Q�0DXM�#�C��\��' ��O:-B�"�tR��+���#����e"O&x!t����yQ#�\�\�*d"Oq�PAV�@h�"������$7�S���}���Qz&`�uET��B䉒Qg"�;@H�y��q�Q��:a*#=��4�䓱��O��t��F��JD����|�<�
�'K�H�	�(���ȿ-2���'1ў�}��'E�l\̀*t'�e�ȃ�Q�<��/N�|GD�K���:EHalVv�'�?��@*�;x�nat��N�N�7D�2�J�,�F83�B�>2,]����O*�$,�)�'+����Z�]�TTƌ���pH���hO?�*� �0Tq�Er�?,(xx�c�n}�(ZTx�PUMӘr�(��t�	�a��1�9�O��?O��I��'UT ,Pv��x]~���"O�x"�if���K�a@"���I|>a�W-	5(�ب ��W�g�~<)T�;�IA?�{����9BĚ����7PI�1�1��9�yR�֍x*F�q@�+F�,YaI�y��6�r�j�D�D9l�1�V\ �X�L���&˩'f��	ވ-���I	��d�<���Nvd@����<�r�k(<q޴R��5�R6L��< ��� C�*�Ex��)Z�Ѳ0��Y8u�9jE�O�W�<�7��J j$��i檀�s��i�<s
U�8�]
�$S�$U`�[%	}�$8�S�'*�:���Q�&��3���?�<��~66��wBW��Z�[ ��-=��=�	�s�QDE�(%�r)۳RB���ȓ�nő��
|L���]�V� ��e�yc"L�Pzؕ�'N���1��aM�t26'�}����(���ɇȓ=����`/���K0�ȩp=$��ȓK| �B��&D�� {R�N 2�P�ȓ[n�O'��z#���F�؆�>B-��kU"B���։��}"px�ȓ�Pzqb�K� ���Ɇ1�2@"���s���A�=I����$��L.�O(�i	r�&�N_^|U��.X�o�༅�g��E�`&���$a`S��>5W�Մ� G�a�$m�/ X�H����=����i�$�E�_�̔�1��2U��H�=qۓ+|dj��1�ԙIEL�$cr�4��)����*��	ڤ�_�v��EnZD������ L� �g��cܺ���G�;!d杺��'-����Ha�c'ڟ,Z.�Z���eC�ɣ^�B<��[1����*Z�q'�#=Yڴ�ȟd49Bc\$֖�HfC��0�)p"Oh��͓ a�����\3X�D�!&"O����+�	ǠaA%�?\�h�@�"OR������aE�v�z��F"O���� ������Ôo��8�"O�<(�%�"�S��Q;���0"O�ۆ�D�ĭ��		4p�q�E"O��k�GY�X���(IOzf��"O�u���  yDXB�%z��a3�x��)�S�sl�������&�Jq� �&(o�B�ɟ��Lh��wp�H��k
`FQ�=	����~�q�FS^"4��ɜ�.\�ȓaw�x �L�s&�a笎3m���ȓ$@��S���C�¤P�@��$�ȓ$�ƭ��N�Q,���@]�;鰐��[Yn x� ��Z�p�X����P��i��P򷃑�D�@����B�� �ȓ ����6������ �k:fE�ȓt�De�Jܿ=�2]PSQ�U~
��ȓI��(��g�+!����F�@Ϯi��*��h*�R}� �!%��91����ȓHz�]��T����WA+bgnU�ȓ'�.��.�F� $��R�p ��ȓ欙���=��X(�h�L��|�ȓc�*�s�QҀ��5�S�Ax,����ė�kh�ӗ�U�K�|�ȓu�0�D�]��(�T#Z��]�ȓ R�xq��A)�u��H"1_���ȓ<���0�������Z5B��h��Dp�;3Cb��VTnm�v%?D�p���ε8���a,D)RN��)D���a��o!�L���\�PF6�`�B5D�Py��ȐU�B����[�zLU��d0D�t!T�;�Q8���5��L���2D����R.�(8 [;ene��I1D��gE^$�r0��EAb�k�:D��ࣄS�j���R�B�S�(��;D�V��U�q�aE�|��"C�\$�y��ٶ-�����M�oD��R _�y���:Y$��%k:g��uR��$�y�X�\�D<h!G�))��2����y�_&����0]�!��k��	>�yD�/�4��Z��E��y�X� ���  ,5z��U�yO�#���c���Jq�,�$C�y )r2��� �N��!�⅔�y��LvUr�L�#9��Q���L�yr#ۉQ2c�N�;93@��M���0?�֥�P�*��
��u0��R _�D�eOQ�<�Nv"� ![0Q��lQԫXy�<��XK[���g��&m�>Ѣ�O{�<�R脪EA���
mP.�#c�r�<6�
O:���fZ�c.�)�fo�<�ǾV\� ����^���I�d�l�<	�c��3��vF�"X
���f�B�<Q��Ɖ:�I�LÊ�AW��v�<#�A�*'ƔHÁ�n�ހ����w�<IV����(RJ����[$L�s�<qU��?p���N�+�|;���f�<�4CFe�faR�i�9^��=���`�<1'mX�a:("�[�,�e��x�<� �)QAR���(
6ʤ����s"O������ 5��X���G"O,�����$�ҕ��<��K�"ObՓa՟D�H@Yj̕K�̱(w"OԠB4 :]�l��ǃ'�Z��5"O�|��)+�.X��4a{`��"O��@wf؁Z�� hP��q{6H$"O�#ՌM�SB5�2)�nj�a"�"Ol`�f�
*6�d�y��V	<\��"O��qGƶBb����"S	�`�"OVdzC�S�HQ`a��9Y<)�s"Oj�RDCO#$hlx!��H�!H�uv�'I�}V��)D5:�R��ANgʭ�� �#(�T"Of9��ɟ�o^F�1�a�1:�>���ɵ9�lʴ��6.���p��c�1i�0}b�B "O\i[T�i�M!@H(V �9�նD�0�����������F�)�й��/Nb������yB���4I����H�1#�yJ�I�<�~"�C2�I���#Oay��U�H2%�B��,ɶ�2c(���p>�+�Vʊ�uȒ!�DaH���+eD�;�ͅ!�2M
�'װEj��^p>K2�-!��yp��߆Dݨy
� X�]u:b?�&D�x��#���#�4T�S0D�T9��F�~�ݢqP�=<�ڶbU�r?d�����.��j)O?�D]�/q�h)PGS�u��1�4`�w)!�؝(���?J�hx"I�"��Ĉ)��y�� �JF��W�d��}K�����tC���w�|�M�#A�u���Y�$p��~�s��R0zT�0X2O�`0�M,UCǋ�mW��Jc�	j�B$�6AI�'���s� ��M�ϓFa�E��"O�)V�Ä}���Ƀ-�%Y ����'�>D�JY�=�ɧ���5�
�%y	"��s���eG���2D�Lb6��	QPe1�̭�� ��c4D���R���L��hJ�^��c!D�|�򪈥7i�� sn��C��%A�0D��QUȕ~6dD��k"�)��n/D���Ҥ�*�Xl�P���ZeH5�-D�
R�* �Dٕ&#-,eY,4D��ӳM��SpiS$�F�!2A?D�8qe�00_�\z0�О/|^��w�:D���CK<Y��͏�B�F� ¦,D��
��M8@�Vy��G�@~28��Mt���gx��kC
�%Z<��A��&`�Ť4|O`����B���$  ^���2,��7#�b!��K/lv���3�!"���ee�O�0�s�M�ȟD`9����1�����\��p��*O��Y���	}�`Y��K�l�S�!�`- ➸G��'A���+_x�r�ۗ_@��	�'Z��W�Z�kA���&WJ�9��2�)�f� �O��AmF�Y�RMK����|�4�a�'����@}򬈢J�(|0��݆w
 ����O��y��Ut+���+_e<\�[�hҀ�OA:�F)��3d�L�N�$��T�A���ȓ5{
@����@+B�zr��pޤЄʓ^��D��-�T�"�xtj�B�B䉵(p�J1�G$&���g�B��
q~�ւ�10��Ha�@�FB�I�(x���b%5/��Б*P�όC�	Q����� 2nT���ĕ0�zC�	n�f@BE�֭E�J�K�ă<zB��|�
2��S���#�.`��C��+P� ����-"�%�.�[ C䉢W�m��đ%���	�呾s�8�g.��E��?E�5�̒l�
 ࣈ͆\��3T�(�O�L��L�L�f�����ۦk�qP ��`�'����Y�� Te*6�<SNa� 	�6Y�p�w�	�h3��2J�D�'i�z@�O�: �Z��!B�=xPHyu�Ǵ|�\�#�Ʌ�#����ٴ~wj%2��2$	��=H,��n
�� @��D��Ir�Lz>��`����h4(�͢�#�>��������M�X�J�dB�I19���(�C6s�b	�B{���]�.�FN�'lq�r�Ԣat���a2O��X�`��.�B1�;_a��	WL]8���N�j$��	>Nh�����\H⑰6j�{���Ab^�uH8��U��k�����;'�1i���9^MF�[�z�1O\Q���!0�<|j�)�pV �p�I�g�(zC�&t�b�Y�`�ś��Øq��C��S�����E耥$���)�j�2f(q���)[�
���N 6K8�qs	�1GZn�:� ��>��Hʖ	��K��ԅ���P�$�d��)�|1��]�p�I"��?���"�J��?K��������$�n,u�S�6iTY����D&���B�Se:�h���Z�F��B�j$2E�ӊ4oDq�eF!�NDQ�D9Ĭ��rtvl"���_�~2��JJQ��`��wk>�2��ĚF� ��U�O�/ !I�&S�ULN�i�P�_�(���S�rg&�b�dD��d�𸳎��+� 5�W�L�>��Gx��O����.ο)�(-���͎:��KpfJk��d���@B��uB�W���F莤,@4hY�gt��xϓk�b�(#
�,�6h§#�.��O�mɖ��mj2 9IX�`�z�	E���i"ѻf&��E��AV��;IRPC��:eU(W���,4��u�j|��J�.��|hD+H�	��q���j����B뉆E��lÐk��p�x\��������y�ƍUP8�A`}�.����T��Ig�I�zj�pe,J�^ʰ����;a����T̨4ɕL��*i�+&h��xEl��uw�|�7D�0�M��Y�D-p���&�O��=�'KԐQ�\�K3R�7�Hm��BV�N��a%�0T,�YC�4LO<!�B�`��}
�&ڲe�|@�'�����X�lÆ�s��@$M��s7��o: (�-͞}�E��mAe�<��#�7��)ɇ�XC�<04-Z��19�mPf���7�x�2�Fz�O�@�CEi
:aHC	Lo3���
�'�����_44'��0r(�v�F�	�Jٞ2�U[C��͟\p�
�����{V0��.��=��`�T�V0z�d��Ɠ�^��/H�.�<�a��O����ǭՀ9��$��/ ������m`���a"U$�(�A�JʫO�z�Ĥiֵ��*��<q���RZ�̓�K]'r^���K�w�<Y�	9E .�K�Q�dϪ��t�t� %��)�'���a �vg8��f�?SJA��$��,9!	�'Y��YF��0�ȓk�,p�Aǣa��E��C?�\Ąȓ���r���~�
����ϙ�����`t��*}P\�[ ��+E֙��I�H�U��P�b�%�䵈a�>A����7k0D�L�נ_#��%�*��$�4(��*�0�tF�T�O�Ι��ɟ���Gh
kӚ=
�'/�1��̕y���a�K�^�^TY��/b��'�L�����>a �
��p`F�� �rLBLh<!p��un��ր[x;Fx�<Ӷ 
W�h	����-��`6k�I>�2��؋@��y�E&�b�-XK}Bm�;'�X= DhW �Μ� ��y2A�'{~���F�"y���e��;��#|���-A�u�#җ38��	�5Dȏ#����gA@x�<a�Fo��L�d�8R�XrP��-@�|x�v�>��@�#����=�:��q$�%,B�x�̖\zC�ɧj4R<k��M�U���4R�,�&#D�!��ye�'�\�� �%;b!ꆫŒ  t�i
ϓ;h9��KE"v�uhY�#ꅠ>�� 3�]�16ԭ�ȓv����#
�p��t(�!�>����<!�������b����.;��1�s�BH�ӒH�5$�!�d�K�����]�mB��D��%F��x���Ē#�(���&'F��rV�H"Hy�a;��J8]��B�ɬDDm�B\�{}��F����B�	��XK&� =E��Y�C�1&����)���],�?%�e�Æ ɔ�HRO��wa���R�+D�,��V;�$04�Vk%�%k��`U��|��&�g}rK��p���vk
no`���A����=��F�XF��ZU"�&�)9<L����بS�����$1h섢��o���(�
�]�T&�14� e��<�I$A�<�Wțc}b)̥gb4)�ԡ��|� ��t��!9�2,�éN� �H!B�"O���p�ŌN���(#E߯8�DpP��8P����Oz�Q�"�SR�a�������Fc��U�~�ӣ��.$���7I�^�<�d�؇ ���C!j�B��,iGLD�M�U��?�>��c'�D" ,CLr�#<�G)Y�$i� ��+Ӽ��D�x������7)(:�$>OV��5B�0Y�T�p!+")�PmU�Y$PPhSE��a|���G�4�i2�B�z�!�N_4��'ɚ�*g�B�"5�Q:�	&�9~�\�S��d�W��I��8�@�-0�ZB�	 ��\h�ᚒ_<�kã���6(��JM�%�O���C�@��n�:���Ǽs��F�{	N�󓃖j�u�A
�C�<Q�◒)Q�%����m��\����w)|%���ܰ-n�͓:���S�b�-[ʣ<��61+֝���Ö?���;R�t�����%�u����#�'ِ�C�>����db�6�R�KY <S��� �X����?c�d�Ǎ�/j���ʧ�:�I�~��}�6���<�e5c���ˇj�~´͋��J!�7ҳT��sA	�s�<Q!�̚?e�U!J]�&%S�	1P̤�s�O6����K�����x�EZ5�
�|˰�c��A�s/0����7D��IDKؘ�\���ؤ�
�2'IX�B��^C�䀪p���?�'�&Aa`�_:��0�â{p�a�'��V)Z,o��crf�F�����ݽd����F�P|X�@c�G^�N�8��N���B��+<O<�+0
��N���O�lS���!?(F���D��Eg"O�|�,�0ZK�q�F�Y��[r�|R��Z��k"	�g�Ow���D{᦬_b�R��
�'�4��4)J@u�ٴ�F*4t\�"�әM��'uX�:���rb��Hȓ�i�.g�����m&D���E��s(�a0F� �~��q!8_�T ��-�O$�@p�K?=�P�-�z��("OV� ���_2h�ڐ,I�
`䘳"O�hС��	��b7KP1���
�'�@���PI�Z�d��a�D�q�'=���fN	V�]P�b�b&\�y�' ä��6B�t���'X��"OD����މ�H�۵C��2@�lr "O$����͗2����#��|`�)F"O�U�F�� %o�4�� w"O:1���SY�QA��	%���b"O��*�OE���t�f�+Z�K�"OȽ,��x^�0*]�?��a�S"O҅±�R
\��Q)֠�:�@�Ғ"OB\��Q�_>�ز!���c�4�p�"O�L��F(d̴(Em<65dH�q"O*]�v��$�eӁM�{+P܂"Oĝ�ŝY�ĸ��P�|���$"O(0K��Щc4���kH9:��"O�' W�s9��k�JK��dғ"OT����	|Zȸ��o�&y��"O"Ԉ�
�+NclP���77��"OFD�M���R5h�ÕZp��yR"OT�S��'� 8s��ÓD(��"O|8�vf��XTʑ��[�/>!b"Oܽ�6�^<>�l�D�Y�X�Nk�"OZݑ�D�X�M0�	Tk�x�P�"Oz��##�[c�	
pΊ�g�v�S�"O:1��J��PQM��OG08`D"O�@��L4+��u@���W��Jq"O��xQB�
�����31��D"Oz	�gjZV>���8/���S�"O�9 ��H�	%~���v"Ob�s��f�Z�YV�J�m{$ᒗ"O��2"�� Ҁ1p��MG�P�+�"O(IRu�m�~;���xCV�+c"O�[@	�V��z����PB�"O�A;fJSM��Q,��I�"O� ���OĬ��M��,�H*0c "O ���L�BX���T�=j�2)`�"O11`��,����FO�\���"O��YAQ\l,����V݈T��"O&���FK-�-YoU'&��j""O��,6��S�,���$y��"O0����r������9_H9��"O�t��eF�أ�	�W\T��"O�%z���L��� ��R�i0�("D"O"�u���p�'�_EF�j�"O��jƓ5c����7���Y7x "O���$�ܾ9�1��
D�I�F"O$��`e�>[� ��P�y#��-�!�9�$�)R��ZA<�P��9�!��D3A�X����
i3X�נ�>s!�D0��aւK����OY�`�}�ىb@	��*>F�,�K��	�(j�@�h�Nd!�D�8/��\���Ē)j� 	VJ���Bb��XE���w���dTʭa6�L�]S��9!oY9�!�d�>0_���Eg��YL�{�l.>�F����(^s�t���py���'r�\qU�Қ7u4�����(z�'�>̪�n�d�:�)B(�s��K�'�f8�u	�G���K��'}l)U�U��
A��;_�h�o9�T�c"LQ�/$|[7�X�YH�0&DL�c#~�:�'��t�Ə�)�ڰ#��� #�H��d�g��H�6_�*��b?�(ǫ�=6Ac΃XY��b��;D����Y�z(:x�c�
w��$�7��I���G"�4:�Ҵ`/O?�DB j�0��Q�3Cr��V�y�!�DؤH�^%�,R.Z0m����"+c�d�c�f���(J&���d�\ڥHiϙ�q˳JZ��|�m�+j2^��-E�~���
�r� �+̡D����7O*���N�X d� �%v$e{��+?����RX-3�n�� j�&r��τ(�a��"OD���A"`����oB 
`���'�,�A�B�|���&!^��M��&��ق��\+0�xC�	�\~�\KT��'���Yu�čz�LC�I `a�Ү]c����Q��D��B�ɏg�<�ː�,(&L�򁖗k<�B�I7b����/S6�:4��W���C�I7{�%r��O&�P����(wsnC� M���EOύENi(���B�It�<	z�iŴq�:�Ə��r��B�I�v�� �q%M'e`���@[;O�dB�I������ƽP��L��ݠTVB�I'p&���7��X{c���B䉾ZG�50��"F�2yB�b
$��B�)@0M�fb@�k���˵7�*B䉇?_:��S�)u�����4h�C�	/Hc�x{�J%>P����=��C�	�f��҅i/Q�� ��� ��C��Z���9_.E������C�	��Z�Qv��by���GG�|}�C��;l�J�D��	7��l���L3X$C�I�{��Uf%���Ƚ�C�	/ ����5�ں�(21�K%�B䉞4(5ic�ܑ"ܜXR��ˍ��B��,]	H�)� U�j��p��I�B�	�LjNXX!$D8�@�:4M-
�B�	�\�\X"�˅:j�~Q�� i�B�I�%�l���M�I��0�bRm�HB�I:������\(�xP����7Mb\B�	��FUɧDS�g[l�"`d�i�8B��)L!*��nV�8�hm(�MO�m��C�!2A�	W�_,N�� �X]\�B�)� �QP�$�01X$���ӃY�t�
�"O �
�/��)�t�T�H�;��Pr"O���3`�=�tX�aE�%�z�p��'�����Q�)&¬�ԫ&9Ā��Q57B1��-`Us�P���!@�MB0x(( E~뚢m�H�kF�韚i�^�)&@�,D��SC�.D!�D�/�!Ѝ��7rڝӵ��O!�$ l�
���N.]�\t�-�'I�4�;3)N�Pnn����H�(��1��c�&8�4��9äq!��ӏF�=��¢O,6-�5-ljP�Q���3�ɣ����ݑ0�(�R��>������"p�H�d��[���e���v��n�CĀ��"k r�`��'ބT�2�Q�g�4�P �u�ܬэ�)�	���
4�	����de� (x��i'l�.�J�S1̇�y"�\�d���Ï})��y�FP�~��H&r���M�3��B�r�O*�uZp	�9 ��MG蛶
�LX3�'�r<�.�����	-*�ɣ�(����΀j���PbR��3�I��<@s�KQ�]I���	BA�����)kt���(x��Dy%{�9�݅X�����ԽNt�����Q�x��l�(kf$���ڒJr�@�"�f�LMs	8TІ|��Y�)ʽn:�6ᙖM���O/!��K�_��z���8 `�Ǝɯ�剪�
���[:%���«�F�O4�)���#n�<��mJ�� �#�'Hȵɲ�B����Mȿ=��$.�:�$�而�Y�0Ɂ��!�$B#�SY�4`P$1D�Tr*��s�,��ズ)i���Ҍ�O`�+���!ΰ>I�ńh��@B�L��b~��&�v�<!� ��(�R��mзak���	i�<���L�LQ�-��ws�EʓM��<9��ƺQ P	ǡJ�H�R���Wa�<1��A4`�$����ސ���[�+Cz�<�5$��K|Y
�x�h��"�R�<���	�bJ���R^�;�I�<9D��T�(̡2���]���D�J�<�C %F=m['&N�M�R(@
_�<�D�X8`7��y�,�6�1���Y�<�'ہ|��@	�MMMZ��O�<Yև��Z���ZFҽ� �@�<ad�ڮB�Լ°OD�Pc1�	�~�<����.<�4��L{���I��u�<�f�ɆH�8QhsCӫD�t�)7/Al�<��L�&Tb�k
�&RʈS�bBi�<Y��Q1F�p����݂c$��A`��hx��A���=�sHG!=�"�Xt���B��B�I+zjU�d��\�5:����b�0*V(X ���F�4�I�1�����ɵ?{�q��)���y��XB�����]#!L�Xi��-��M89}¦W',]��O�n,w.3r���ʝ����ƓD6�`��7? �j���D��`� ��SDDX�C �O�!`�U�pl��V�	�dp��a�'rf肖�aw��'g��Q�?�4��h.6A�@�'�� Q%�%g+�$��T��R8�O>��DԤ�J��+�'���!B?z����鞾1���ȓ �n�Y���S>|q�Qm���>�kЮg��~ dUb��L����肨G;����_�<�r�`�':4�TXˀ1?���uEW�2[� �'����0�#o�^Ua}�Ȕ��S��L�c��@8A
��<Y�g�?`��Xa*�>��l�<-�P��1�6�z�;�e�<鵪��?���q���&h%˄�g�&`1�Ԅ'��걛#E�h��s����l
a"O������>'�()���%^��t���ʩ)qO�P���Y���F �R�	J��Ц�P�C�&D�tX$fwF�X��Q<<Z��kf�$D�tJ���BS�H3r��	��Á�.���p:�����/5��%YS&P�=�89B���#r�C�)� �A���.��'��!j�9�B�^%_�t�H>�b�>�¯�9�J1��3��m9���v���)3	]�R�I���k��7r����Ɉ�@���ѪL8^ndg�(�OȀ�"��cyx,�P$G�D=�T����5&�#n�>I�aH��n�� Iu>)�d���n�����.Ɠk�W�2D���M��ANZ���D� �Y���Q*]ܺ11Ą��T(��S�p�J���)_��y�'3!�6(�Q���x������y`�?kr�X	՘�~l���]F
��㶁։q�\�i�'�8,l��D�Gx҈F	$e|�x�Ip�P�X��S��p=A��-+N����m��r��&�h�� �a�N�CS(v�&�rG����D\��ްz�Փ`<�)���BRqO؀2tN�"/�L���'M��p@�բrHA�'��୕*y8!b@��T��ȓ~lK~����J�f%��%`�=0}V�w��0;G�) k���c�	��yW��9Eq�}�ե�?Q��A��R��y"�J�)ޔ�H%��,U�jĉ�J�#G���"MH�Q�4�B�'� 	"�J�*ր�Dy�eS�B� ��Q�ZA2����p=�"��*UW��	���Om0tJP�`�J*ғe�l�#)I�A�
�2��Z �>�r+�6,����N�
�ꬸ��L�:)&5QT�J-�y⣔<�>���b�R���8IN`��h�K�Dy���Ƣ�y2��&�������.@|2���T��Yy�￟��a"�>�0G�ʼoV�(D����
0�M��y�ǅQ^@�u�M�<�,=֍��bt ��!}"ۦ ��l$܄����)z�(��Nƭ�2�Ɠq��H)���aq*���Eh�8p����B�"F�2�Oe����i�ף�*�XђR�'�q�w�T(�P��'t@I�+Z�nl�Q1��^bdԍ	�'if�1o��"��̠q
	�]�� @N>�Q��.^��8h�F&�'m!�M��FA7L*�8RTGL)���r�`�0+�+w1��I��N�
�J8M�q$��W
*�g~���t��D(�I9&��P��&΋�yb�� �h�@"��{�d�c�R�-F��p���0?�cȟ+L��3��h�,�	��M�<a!/O�i} �*cR�I��a�m�|�<Y'.I.��ҥ@y�%���Q�<Yפ�Q
���9�L����N�<16L�.� X�K�M�<-��·q�<���[dtI�lխ?\��!o�<1� �iጰh��Y�K�k�j�<��&���+�t�HD
�ȓPs����Tg?��$ꙉ>ܩ�ȓa������!R�*a� O�qT$��pP�|/�--2�kҵ*�����
Xi��Ħ�:T�I��v�t0�ȓ��@���׸ tN�*S�­SM�������#`��Zq�&HMA4���E��2&%�:!�Q!��e����2l����̐�{����߼|h��ȓuj�Y�-�aV�놡�7U���ȓ<=��;F��mG�	cn(,�Fh��u��R�LD:-���;WjB|M�ȓt��e ��H>dFTk�'��x�L���$U
�U#w&�-�+Kt��,1�)��$J(N�Vh������9�V�a���A�}z�J�R(:���o�(����uV�����*L��ȓ(��h$��.H����c�b���RI�	�N.D)��@]�?�B��ȓ 1�gkS�s4���恕Y���ȓY8��I�`�.4�@H���'tNم�	�=����M�p��|����8R��)#���6b�B�%z}v��s��D*ve���Z,O�B�	���uB�K,(V$�(V@�B�	*ct��!&ƌ'_�r%��/~B䉼!��=��Ġ0��1$���I`B�)� T`pqbU����B�InЉsG"O^���ċyS�a*�/JFh�]��"O�m�pƚH`��j�m=J]0�"O��
sn�d�
�aE'�Qc"O�P@��+�����I�M	�yz�"O�p)T�
��  ���#�2�
�/OB�qO^��ç�`|����2�6Q�C�u`��(�����En�<�2�'k$ܠ�4�ۓQ�&��oضT���'��IR�	�0m��ᓪC�J=��Oَ\N�4B ��z��I�|�t�zR�Q�@���S�O�"�yt*M�wn��NGKO@����G����a���tP��4O�?)!n]?s����C�{����v*����;GJN�z>v����i�L��Or����J�L���P�'%�U�&H�� �ܴ�V�����8j�� a��>��)���2q�D����.�����*��-j��(��˩�?E��DT��dʕtquQ��>I��IU��0N�^�IG�O��	�'0wH<�'.�R6�QYH�Te�0vJ8�7�[?ys�&*����)EZx��	؅�F��!R�^h�B��7*��Y�LT�a ����O���iF`�)o�����W�}���r-f$�����+^�~1�'̎��0|��&O��$��KG.�V�����Zo@t�4�"{�v�:�I:[޲���S3E)h���U	z)H9c�i]>(�x1[�����Q'u����çz12t���M~>��Bn9F�v�S��x@BJ9I�����OA>A�DD6ސ�2gi!j�+�'�Zp`����7�$�ǅ�f(fh
�'Ǌ���C��p�Ҧ����8K
�'I��!%G&z�0�E�.3=s�'�\����4?ld"Cc��#r����'_B������lh8"ʜ=K�Y��'b�]����'N����镎EW6�c�'����Ū�;&�ˆ��?Bq�(H�'��в�Fr�E3�Ǻ5t��'���*@�$ϾX8��4s����'Î=�I͎10�d	U��ʐ�'�=��\+u�q��ڶj<ة�'���y0�	�_j��2T�Ӥ�`�k�'�d���A�5�t�#"F-0�ܣ
�'r��r�OÀ}�<�#È}3�t��'��Ġ爋�RB�<�aM2t3��[	�'r�D��H\�� ��.�n[0}x�'��]АbZ	R8n�
��˷Y#�=��'��P8�̀>g�2 ����6Mn-�'�l��k�OU�L� F�x7���'@p(�W!?� ��g�@ l����'�0
��S+�h�*�L�&8g�j�'븘��EͻN�;viҶ[��Q�	�'����& �+܎E�UnH[H����'�Fd'����@22�ȶZ*��
�'��@y3K�9�8h�1 ֽB�<���'OR���R���HR&˗<N  ��'I�H���V�%�a��9C4P��'�p��reɉocD�ɑ��=�@5��'����! f��Q�!I��*�j�X�'����gV"m�t����Q$(-�� �'� ��2*Ϋy	~�X!gH�1/T��'vF���b�8#��ː��6)��y�'׆� V%X�o�D	����12�QY�'DsĦʖ}9\BG�As�����'r���&޷|��yS��Q1cp���'G���q�M�r>��Z"+&&�����'?�x�5EZ�Av�Y�d!��2�'���JF�S4xC2��lf�S�'K"��D�Ѽ*���(�,(lČa�'`���g�S�}$�
�i[��Q�'�d4�e��(b�� �a�5MOJY)�'�TT�D� 'Ɋ�CI�<L*���	�'��W	H2/�& QcM�U}j
��� ���]�$]ֹ��g 7*�hy0"Ob�C#�=�Ɛ�fZ�0����2"O\�����(p��Q�BE�?|���p"Op����_ϐ)�ecJ*'2��3�"O���V�Q��	#Bl�@!ʃ"O^]KW���4�H@Rq���"B"Ot��$-IR(b@��ꓠo�b5�G"O0��҅5}�h0�O����7"O)����|Yq0o�	��Mx"On���(ګ&����'P����"O��2e�ܡ�P�Q�n�q�*��U"O �^y�(m0bm� ����"Oơ�㄁5  n|sT�N�U�~�pP"O��+�bةJr@	pN ��d�9 "Od����2
&�E0��G�4� HH�"O"�Q1��B4�-h��&E�pd3%"OL�"#���`?d��A���f��t�!"O�kg�a��IB��9�RdS�"O���0/�#a�����V�_]���"O2��e�H�>�a�G�ʂ}J�� "OleH��@^��܁§�./xh��"O`��ɸ86�Hq�'��4���F"Olv�N�
�q	Y�35J�"O����IH
d�G)�(���"O2 ���V�Y �g �U����"O��JT��bFq %h۷E ��"O�t�'GH�&��0���Ч7F���"O�I�I�y��l�L���I�"O�l��J� �*}:a _TNI�"O����=`���3 N41G`cf"O��d*��9��؆�(*L�+0"O�������F`N�y��"O:uP�ʆp��t���5ɶ�"O��k��_!�!��Nc[�廖"Of�BEf�M�� ��g�<I�)��*O�
P���gj�C(ĬP���'�ޭS�̖+<7��*E�T�h�Ԝ
�'@B`1Q
�����$.��e>ly
�'�&���j�P �7J��(�r�2�'A�<gk�yH-8��� (����'v2i�5C6�{vk:+�Ű
�'#�ЋT�ݮ�V��$H:<�B�ɕ)Ύ$CMQ�
,�DȊ ��B䉅t�S�O�7� "��)G�pC�	��L���.��3�]�(JC�I�^2
��&e�x��o;1xC�"O,�Y:!��dH��e�7�B�	�Ed�l���P�#-����*6>B��O<���ㄓr�6�p�N3	�B�I8�~=�j�+G���C�	�-�Q*%c��4����LwzC�"H�`a[�9�&AnN��zC䉞`�̝
��еK�V��g��>sNC䉿n�P8�-[."�іK6&�(C�ɼ&��  e�F�\c@�"�Aw5C�	�d��(��C�|A�b��^�,A�B�I9m����J�#Zf�p�g! ~��B䉯j}�` nB�����&R(ԦB�396��c5��\Yd)%焐uX^B�I�R%6�[&���G�@i!�aX�n�vB�ɦ+��ʢ�	W�@��$��jb<B�	���r'ҡiD2U��FU!4�HC䉤e��̨���O_���E��	t^C�I�y��&m�01�h��Gg|C�)� ���0�ϴ[��T�7��j�<c"OVq�C�J�[XZq$لܨ��"O�1��_^7��y�I�\�
��"O���,@l�8�"�?7�p�4"O�S"*5^Z�0����t��Q�"O��)��Q�v�|h��"_�K�h�v"O�9���b=:�����v��9��"O�$�RʈB���BH�z�R i�"O����FD�1�Z� `x�"O�*V�̔W���B�e�Ջ�"O���Ta��l��$�Aפ+�Ȉ�"O�<a1�W�5� ��E@V c|P�"�"O���2�_8H�p��mRdal-W"O.�q'��50:š0�ƎvU�-K'"O�⒍C6
�^M��.͘3M����"O�1�R�k���K*Q��X�"O���L_�$���s�P57"h ��"O�9tG�C�>� �'F�\�&��0"O202��.��X��gCu�h�`�"O~�pg���ж�G�
-x ��"O�Lh����j_���s L�w6\�q"OB��RAY�E�4���P8��yA"OͲ!^�,ZqIc�Ĺh��"O�� �F��9PI
2�����"OT\�BU
�u*Diß*�6��"Ol���EhL�S��G�t�[�"O.��'�r�V,b�O���ˢ"O�Հ�P`�XyQBo�*�"O
x�Ed �1��ajg �=%!n���"O�H
S�0U|V���Ů{K܂�y2D��a`)!��6�D�8 ���y��ż%&�8�Vb�0��I�c�L��yb�
��X}�(��)L��hf��?�y��Wb
F�����+�b�9V%^)�y�̟�a���MЖY4� a����y��;��@&°O�5Z �V��yRm>O�h2�	�p�.e"%�y2�
1Q4L���CS!��yċu��\r�IT�A�@Lړ���yb�FY�B��wnK�$�
Q� �1�y�iM�g*Ȱ��ϕ�M� Șv�_��yRI�p�m��E�F�ha���y�I�"&�^A���Fc��[T��y������>�P�y�I�y2N�u�>ܱ �.f�Ȉ�2��yRќ/4���ǗR�0�� �ӿ�y��݈1��(Rs	�)@��]�:�y2M�(�	6 �?(~���U$� �yb�ɗl��Bc�ȞL$�bg^��y2�	10�L)ɣ��K����D��y�	 :x���6K���[��yBiTAy�nB��*��.�<�yR֕4�"x���%{�d,[G�>�y�יTI����Ĺ�F�[:�y҂�e�H���X�MQ�l	�g!�ʘ��iy� C.tdn$�7��f�!���oDųvKt]�YJ"��C�!�d��|�p�%�W�mP��gG9e'!��P7�$�cO#{��h��DS9M!�d�@��ٳǏ6��\; �?!�١c���qA�W ����%r!�$�&r�pr��)|���ҍL �!�D��Ǩx�@Ia��M��B�-�!����Z��$����,QƌD4I!�� �x��~�Nx�
O��2=b�"O@��ffO�ji�`���������"Ob��7L�!� 	�jH	m�t���"O�� sߝX���2�P�<�Y:�"O����R$wپ�
�IT�j��;2"O��[�+�0��ٛ @�2��"�"Ov%b�/l'$4�r�p�"�R�"OBá%�(�թ��@�d��0І"O���d)���Y����#"O�E��윧Y�
��6g� Խ�3"O�t곣��>�����,H�L��"O�J���֙�tj��`�n`��"O4��u-�@N͓fi�=t�P6"O��i�ʩe�d� SG�1rp�@�"O a�G���;n�0"Ve�?T�#�"O<�5������� 4��Ȩ�"O��B2,V$1�Rl�4^�B�	�"OB�y#oP1N5�Ě���U��`	�'�>�"4���k�r٘�	�	;;��q�'��5��!���=җN� ��s�'�<���I�����4@�L��
�'(�����H�����A�����'����i�*Q6����@Y�'�}��'��4S'�GT��ض��wa���'_
�"  ���   �  >  �  �  M*  �5  :A  �L  6X  �c  o  z  �  |�  �  w�    �  ]�  ��  �  J�  ��  +�  ��  &�  ��  ��  �  W�  ��  "�  � p E � $ �* �3 �: �A �G <N Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#����!LO� ��!צ[�n�V��G!��~�҄�b"O�%��$Vݞ�x�` 7${l�"O������$|(�bE� ���`�"O�4;A��c���A1�R9�\+�"O��:�E�M�&���B��C�"O&��T�Z	/ �x O"g�<!z �'3&8lZ"i�L�V�У#��)!%`'VB�I�`$���(E%D���(H0�?�t��E_襲ү� �bEx7�ͣ �B䉙s��u�"ᖵ?�z�P�(c�h�'[ў�?�v�g���ԯ�J��xhsL8D���D�,{�TͣE���&�(��6D�����SƸ�6�f�8H*f2D�l:�ЧZeN9�2@�PpT@0D�n�X�\0*nJ��{�/4�4KbIߤ*�pQ�͔�-K��)�r�<%�1��E�o�%V��n��+�-��&��C��L���5�	-0.24D���%
.�����AG�R���-}A/�S�'}Ѡ(�qk��j�����R	al��d��)��  �d�jDeN�mFM�=��'���i�<�*E��#{N�Q�	�'� �,�x4��`(���^Đ�"OJ-��-��h,ч&�9`�n�¤�'-�O�y�JW�����w�b}PEM�+�y"挤$(��B���p�L1���^��y҆��!}���B�x����mÙ�y���l�f��wpu@�.A��ybD��~`h�� � �څ�F��y�X�\�j��#C�?�ج�Q�R �y�V\QR.�( B�TB.���y�aǟJ��R��#'ABX{��=�yr�L�o�8dpe�;!=�8�3�y�hө&�$�R���zt�����y��J�aA��b�<	u�Lh��H�y�+�9�4��D�X-��\Y6 ��y�)�mv�pr$q�M�U�^�y2d?��̨�G Р�)����y�Ǚ�hV,XLY�Pu2%��/�y�ʊ7S���c���޼)P@���y2��=`di�'MUy�V�ǥY��y�fT<a���Q��� �v���.=�y�J֜'�D�;e�� l�x�����]�<�#�:c���ۓnծI��M���i�<I`!�CC�="� 	4騜���o�<����7)"^�c����8Eok�<It��/NQ;Gi G�Z�k�P�<�hX9
Դ��P.Ż. Yy�#�J�<!�ŋ3��s-Az0�+�^`�<RMڤC|��'Δ ]沬iQI�_�<Y�e\�6�B5�w&�$W�$h����p�<ydiO5�d`VN֕$X��aF�T�<!C��K�fec�A
���AS�Ke�<���@�>���y�b՟P�|��F�F�<����	��������.m�3��w�<���	14��$C�k�2�b�cl�<Q#l,� �P#K�,eV�i�Kd�<v�!}	PV)�Y&�Ih�_�<�KU�3F��9�ޜv`���KL^�<�F�C���ڔ�.]Ʈh��nGZ�<����]��	3�Jۓsq��� �m�<�5 ��7�Nx�&Ï4&��b�Ǖm�<�`":._Zt�"!Ս0cV����o�<�Ɔ�*o'��z�*\/��1׉Ai�<� �	�����iR�JM�1��І"O��8&�?s7�����I��Lx0"O�rt�S Y*P�a��$M�Ms�"OPɘ6���^;d)ې��*Jp\`�"O�e�牂��^5;�I ���)�'��'���'vr_>����,�	!K\j��s(ԛb�SL�D��Iʟ����	ӟ �	ҟ�	ß�ɉr"���bM8����R8,�I埨�	���	�@�I؟�	Ο�ɦX�\`x�aZ!�p}��$Et���IҟX��ӟX�������$�I柨�I�lT �(�P�`뤈�ƆC :�Iޟx��۟����,��ٟ���ß��	�m�R,���1v�\9C�rq���	��d�	ӟ�����D������ʟ����^wp�I"���i=*�:4DZB�p��I՟�	������@�	ҟT��ϟ���IP�]����X�|E�A�	�-~�����I����ٟ����,�	ޟ��	���|�/�̑җo�>8�)���|��ן\�I㟬�	��H�	Ɵ �	��n�`�#÷_8"�����9H����˟�I���	ޟ��I���Iß��I���`ūR�5�v��ՂH�zq���I`���P�	ޟ0��ԟ,�����Ɂ+h��A��'(���DT�Yn��I��	��`�	ޟ��	�������ɨl�49��+]�Y1<�C F: CR��Iܟ`������	ܟ�������۴�?���Y}f�å��/;z<"�b�g^HJ�W���	Jy���Ov�o���,���,`Ԅm���
��N�Y��"?!r�i��O�9OD��H�:D
��Q�^b��P�^���OlM�Q�e�D���d��*�O�^�blG�\m��BR�ӟ�t�yB�'���q�Oi���3N�#�`ґhW#:���b�&��E�-���M�;y����DKӡ �N̨`��D�8���?��'�)擾�IlZ�<��b?*����?%{P��F��<��'{��$U��hO��OHi!�ؚ�
���N�5����v5O�˓��A%�V�\
��'��P#΄82K��ʋ�u^d�b��$o}"�'�;O|�2B<CEfW�Wl>� G�4�~��'�b��` @����d�Zӟ����'��<�&��1Q���dc��d�����Y�@�'���9O6��A�Rv������B��I�:O��&;V i�O5m�S��|z�>���"B��uz5�@"�<����?1��c� �ٴ��De>�@��\���H�B��.&H��2�0�&�>���O2�4�V���O��D�Oh�d� J'(Pz"V;� $�,R2�t���OK�̜&��H����O����A�3?Y�B��~�a G�|���!���?��0���a�f�m�k��D�O���fn�hҢҘS[d59w�ź<�lt��Ǜ�L��Ă�OL��sF7Lx��J�tݱ�M<��^��±D�r,ݐ���`x�@��N�@�Iß���ʟ�Ky"�q���b7��O2M[W�fT`�E�i=F����Oimh��T�	럤o���Mk7	T5 `P�J`I*6@\�5 ��"�Y�ٴ��D� A:�A:���������A9Y�P�Z�����gΈ���$�O:���O����Oh�$7��h��qJ�=Y25���چ4\\A�	ϟP���M[ת��|���Cu���|��D�7(���g҆BcLE"6N�4R(JOƝnژ�Mϧ�Zyc�4���ŉ�� Iʵ>=�p!d���e��P�H�?�?�Ӄ"��<����?����?id�V�*�pQ��:;>Z�R���?����٦Y��.�ly��'���aF@����g�����ڶrm �@����M#$�i�bO��`�5��Ȟ:��};p�Y�1������>�ec��Tey�O3�����S��'�j��?}�t�4̋�[V�8�'���'�"���O��	��M[2a�k�ʕ2G%�,s�J��ʕ��$�����?�3�i��OԵ�'֛��2&�|\�tj�TX�Lq� �.vql7�Ϧ�j�ۦe�'�x4����?YqsT��Ps� �3{� Sn�\%�PRB|�H�'g��')��'��'���B �mZ2�͈�s�ʍ��[޴5��	��?������?)ǰ�y�ˆ�4T�:�i�ҁ�'i�_�n6�ʦuJL<�|B����MK�'R���:t&z��aO
1n[�}��'. �A�×����|�S�D��ҟ8�QN h�NqI��Ą�ȴ�5˟(��ߟ��cy��s�,(Cs�<��yX�d��(D�h �KZDO��O>y�A����M�Q�i�xO"��d&I�4_�� V0��T���*�@���Q�b��v�&�2��D�RiĂ>�x8Ȁȋ�~�� C̟,��˟h�IßDE�d�'�VP���I����SRŤ��7�'�@7-�%VQ����O �nb�Ӽ���o��3��ِW� �i��<�7�i�t6�����Ō���'�&ih3I��?������F�.`�!��ڌ��'c�I����ӟ��������A�ܔ2�O�h�z:�HMn��=�'�>7͝� k���?YM~"�|�����4_6 �h�A���5C_���I��$�b>� ƫ��RKPi�CE�W]B�p�&�(N])�Ty���$�\�ɒo�'��	(u��)��l�Q3W�Y�9�*���ڟl����(�i>A�'�P7M٭@����$�R�`M�/��eBAZ2�h�D�ϦM�?)S���4Y�f#r�҅QP#��H2��K�
Lն�0��V�Zn6�(?����{b������'��� ��{���_4F�
�;<��PW0O���O��d�O���O4�?A���F1W��M3TΒ�L�$}p��ş������޴;��x�OL7�6�D���`M��$V��
#���9���O����O�)��>��6�3?��;���i�%�������|2�i�%ǜ��?�A�6���<��R�D(;���#V΅�_�����U�O��oZ�D*�(�����I@���ѥq��ÇB�P�B!i�c�����S}��'�b�|ʟ�%� @�bΤy��M�)3H:db"�X""fy���]����|"Ł�Ob�L>9�kGQ�|T����	SuC�l�~<	�i�xUj���X�`�����ݒp.�v���'�7m2�I�����OqD�ϸ"Q��� �-t��a��O����R�>7m ?��+
Y���(t�A<ڔr6�ܥ#��Q�ah�\΅���&|Ox�R�L�Tw�ŪP�p~pec�@���)�����<�	���:q��yW��3=�\���l��?:�MS��6S��6-��-�M<�|�	��M��'B<a�#g����03$��&G~$'vֈ��Oɟ|j|�Z�4��ܟdX�*O�A5�@˰�p��#`�ן0�I�q�J0f��zy�$o��X��������Oz�# N�9KjUb��]5;F��/�O�ʓ�?y&_�ě޴�r�xB,B�(Y ���,ߓ��J��9�yb�'���Q,	!�����X�h��7&�B.C���t �F����ĨrVr��n�ܟ��	��\�I��4D���'��p��@2s�x�&�T�Z²@���'��6m��`�d�O(m�}�ӼK�\�Ta��MR/g��R�eI�<I��i��7����A8҉�ݦ��'�<iE��?���FP8�:bR�UKB�kT,"$�'N�Iɟ �I�D������
n���8D
�0œ� �	W4T��'N�6-[.�J�d�OR��!��9d��hW��\����6!��1�O�$�O��$�b>}����r��Ձ�.Q+�]�6��!z��+��3?�&-]3K���'�����Р{Er��f_%$=؀�*��4�L���O~���OZ�4�>�.�VMW�l�o�p{2@�F�gT��D0�y��b����ɨO��d�O��oڐo��щƯyZ�-��� ���	������'�F,�v��?I�}2�;5��9Bǉ�R9�	��A�B��?Q���?���?�����OV"JC�(Ht�`Lq�S�'���'��7m����'�60�$/
�CG�<S.Lba�0LB�&����4'���OX.Y���iY��
^@$@�&&P�Ub�`M¶g��x!�FǑhe�%L�	Qy�O���'���:~��m�:+�|�hT�[����'���<�M����$�O~˧B)�Y��	�48-�R��]H���?��S�l�I���'��K|P�k� ��萰i�W�����G?G̦���JI��4�>9�� M&�OB� ��)E�*��4n) "�OR���O��O1��ʓsf�vJ���)�'#��5b�1?�pI�T���4��'/�˓�M�����)2��p5`Ns�|��!�;���ef���K�At�"�,3>����b�O#\T�w!޾{ Xѡ�C�1���A�'�	ϟ��Iş��ş���f�� Eצ�Q��(�Lԋ� �dO�6��6L��OF��!�9O`9lz�aq!i[�B"	��N�/+6L��d�����Ş7�ڴ�y�@��L��X�D_*|iC�Ї�y�@ț%_���I5D��'Z�i>Q��e�~�SW �c�9�æN�X�>��I��$��ğȗ'�H7-�,�"���O����z��L�Ң��|n�Zш �& �lR�O:���O~�&����.+o�(����K(/�Xg�&?�ס�\|�� .�P̧W~���Đ�?Q��ȯM��9	G�?z��Q��MK��?���?���?��9�0T�F��XG��ܬ*���&��OvTlZ"���'�67-&�i�ը��D޸��١EY� �|���I֟������m�B~ZwN	�p�O{�d�T��'��Eh�!�1!��d�t�D�	qy�'\��'�R�'
�%N8B�z�A�+�(E4��Q�H�^�ɾ�M��D��?����?�M~��L�j�c�:���`s�9�%]�����'�b>%�e��:HN(��� m��#�T�p�� �py2��"~1TA�	(��'4�	��e����$k��y�K9l�\�����H�	̟��i>U�'v�7�ΎJ�v�$�	r6|���M�*+�d��eeV`�f���ڦY�?�EV�HݴId���d�R�ƎW�s5���X�Q�h;CGQ���7M(?ᣭ�^���	=��߱p�$�
��5F(dzdhZ�Ol����ퟀ�����ڟ���v�W0�R���;�����ˋ��?Q��?�Q�i�(ؚO�R�p�`�O����W9a�q�g㗻b �uĈX�����mz>%��$
��'M�,�q�'��eR�!}x��"��KV�}�	,,X�'S�i>���ğ�	�x� d���M�I�.1;��c=�Iҟ�'@7�_u���O��d�|�&�K.p]�r�&a�r0��.H[~�,�>���?1�xʟ<�yS�"�@�� X	
�2�����Ud�0�o�y{�i>�r�'�� '�T�F�B��A	��
5 ?|Q��k����П���˟b>�'�*7�
5eB�����(^n�B+�(q�0�AF�<!źi@�Ov��'���)e6�)�AL�`�P%
A�3�BAs����eӪ��f�y F��π ~p;�H�$L�@䃕.��"��5OR��?!���?)��?����I���YP�K4u��@�'KuNX�m
t�hd��ܟP��[�s�����w�(�<d�%	�R�0`qP)ّ�?�����Ş�z��4�y���2��vM̉0�!��K��y.�7j����� +��'���� ���j\��Hso�*�(@��	~�:H�	ş����ܕ'RN6�ľ9~���O>��X+4 0�8��^
G�U��m����+�Op���O��O٪/ӗ!c�5���I�&�ra��PkB���)������s�S�(�R����W �8��IV�ȓP�Y�������IןxG��w��S�"R07:Zec�G�C�9B'�'f�7M
 )-��(���4��С��K7B��	�ǃ�q��� =O��d�O8�d�H6�7?��\ޡ��'˺�ʑ� p����/l���U�"�Ļ<���?����?a��?)��;+�`�d(_[!�\��)�;����+�ǒߟ��֟x&?��+0�y� �"�^�K���3�r�p�OfmZ5�MCR�x��D���p�X$� AH	+@-��X46cld���7Z�I9bK�����'	�D$���'w�=�WC��G����C$4ڔ��';��'cb��DQ��8�4G�Ha���k���׬Ҫ�bP'��;�Ԭ���4Û6��^syB�'�F�~��q��EvB8����V"K�|QJ�^���6�&?�EiN�t���)�����stk߶Co0*���G�\�% ��<1���?!���?!��?y���aš�%B C��2X�W�X_��'>��jӊ	 �;�8���-%� x �N~A!&���'���t������?���|�7�U:�M��O<�cg�}� ���h׳z�<Q��R>�,�������O*ʓ�?���?)�l�RѪ�j��/oҖ/x_,	��
�����	YyB�bӌ�Q+�<���IJ�&]�Mǻ�B]�C�?n��I�����Ot�$2��?5*F�P8RZI�g	ɟ/���֦Σb9�gD\�z�~ܔ����^ПX��|b����=��F80�C�Ծ8���'iR�'���TW��R�4> ��P��$���BR
V�1���A���?���m�����Hi}��'N�S���c" #f�')"`���'��6M''j6�$?��O�;��	2��fI�~����B#n- H鑭��y[�������������ß�O�.� V%�2M`�(�٬�xٳ,{�zp+W&�O����O �?�y������ȠPc��3��vCp��0A��?	����ŞS��ڴ�yc�;�&��g��;^ɀ���D݉�y"k�}ڡ�ɝl�'�	����	.aGp��Ƀ
6�90��A��d�	ȟ,�	ş�'f66m�+�,���O*�$&l� ���&LȤVE=�㟼�)O��ds�D$��꒦�Y.�(�,�Y�hy%�'?�Q�J>x��d`��Z���'v���DZ�?q�fN.��kC'Z ��֋�?���?���?y����O�}�f��L��څO�nh�Ը�K�O�umڹ:����	ן�ܴ���y��� n�s�n Anp�?�y��v�inڐ�M�r.�2�M��O��0��X����E�-4I6
Z��Q��%�29�̒O˓�?��?����?���>��B� �����FF4U�*O��n�0.��8�	ן���I�Sן8��*��V�\]a׋�G3��kq*S����Z���q�4z/���O�t�J�G_g��d+�(s��e�%���3%�Aɕ[���7L��R%�|�	_yB ��tp(��MB�c�ME��$C��'��'�O6剹�Mkc�?	qB�)ErM����Tۀ͂��Y�?	��i��O��'	�'"�$;��e)֣�V��M�EE��j��1�i���!�)���OS��%?u�]'2����n9�n�H�S	,���I̟���ğ��I���	v�'P3��t��`��9�̓�o7` ���?a��`��6� �剗�M3N>qУ_)�H��Z*_ܴ��'��;���?���|jDHT��M��O��T)T2�H��+j���bSE� k����c�O���L>�-O8���O����O�X ABFWd�O �S�
�	�/�O�D�<b�iI���'�'0��'�ӖM���|��E����m{���OT�'[�6m�榉`O<�Oq�U� ��Z�%��%\_�D4�&��	�d�뚡��4�2����D%��OʠG�6�B�+��_
1�d���k�O����O���O1��˓���̢qyP#\�t�ٳ��
�
�"�x��'4b�x�T�$@�O"AnZ�m9��B�"��6�����%/����4_��v�Z�v���R4+7���wy�I�!p��a�� KDu�ЎU��yRW�(����@��۟ �Iԟ̗O�vݛ���2&@�;!h��u��z&�~�����d�O �$�Ol�?)8������/'	�Ѣ2���a�ʄc�h��?q�.����O*m��i_��3�}Ĵ%8�J�T�D�$��<YFP�X���dN�����4����*d$��*tH��ˁ�D�::���O��$�O��G�&�Q�$R�'��f�!R
��# 9�ysF�S�=h�OvA�'���i;�O��0�ݕ( ���%�0	z���`��f���OF� x�ԟ�YCL̝.j�d��O�|H��'LΟ��	��0����D��w�D�.�9w��k��,H 5�'�>6-�w��$�Of�n�i�Ӽ�P��U\،�T	_+�H��A�<Yֵi�(7��妵j�*N�}�'P.���h��?C� B�P��}IB|�6�˥+-�`��B-���<Y���?!��?Q���?�Pc��u���\,���g�>x�'��6MU>)�˓�?�L~���!4xƎB�W��U!E�
�|��S���ܴp�v�0���4[��k `����"U�_¤u�e�>w�˓V�JK��OܑL>a.O�X�ÊY/2Ά���@ŮY�Tt����O����O ���O�)�<1R�i�����'W����lVb�����N��t�T�']z7m1�������Ov6����*�([�(�l�)�h�iT�x!
�t� 1mZp~�>��<�Sp�'ڿs@�E�$*������}�$s�K�<A���?����?i��?���)ۼE���y#i0�
�����,���'�bji����%�<iP�i��'�8t���3b�(��
W�\�0�#�$��{��|Z�ɜ��M��O�q8���]Zm��ݗ�h��)Ɖ.^�����ؓO���|����?��7��)Q�g������qI��R��?a/OJl����%������Ix�$�P�w�Tqy ���;g�Ѳ�Ρ����V}��'�k5�?9�6?k�i�OC`��8P�^#k9Tc	Wp����|"���O���K>���i@F��qH_�p��v��?I��?����?�|:,Otxl��F.B�j�+3q"�s��J�E�XK���8���MK��Ͻ>��
f&�1�	�Y��W�j�������G�f��6����$�ϩT���~�w֩1��|طn�51\�S�hC�<1+O����O��d�O����O��'�p�{-�R\�O
;Sz�M�C�i�jI��'���'5��y��n��� �*�� b��Ђ!ԈD�1�����H�4{���O��A��i$��#`iA���;]�bJ�eF!>�d�i�����s\d�O���|J�F�t�`�IH�.�Ȉ�V!�Q�@1���?!���?�,O�Uo=0F������I�g�J!&�	l�|�ʡEȄw��	�?a^���	���I<	�N�8�c�-��YRi~ǌ(J�R�Т֩�O�V�	�i��ڋ'��0S%U�Nu9@g�?h��'l��'MB�sޡs��ݫL6዆&2����W����4H|�a���?��i��O��K�x� U�)8D���i�F�2���O����Ol�Gg�"�Ӻ��Ƙ.��g��a��gJZ�W���ե̖jS�O�ʓ�?���?����?)���2�p�T�Q���0��;^D�)O�)o��e����	̟�Ij�'qu����
�%��Y�%��B?�	�W�ؐ�4N��f�'���,�p ���rN��.Q7�!��Z�R�ʓFe�!� �O@q`H>/O�-��g��H�lś��אg�����O���O&��O�	�<�ְi(�ۅ�'�܅���f�h���B���4��'`7�>�� �����5[۴u��̅�@tuJ�Œ�L�P�0��"U��P�4��D@�z�:1K��_�����N�	h:�������#�a��~b�'���'�R�'h2��o��Q��04�� 1@ �M���d�O��Ąæe���w>i����M+I>��(��m���K��H���-=��'�67��˦瓫/��n�q~��nI 	�����z��ژ5�U%�џ�Ё�|rU�d�	�L��ޟ�r���D,Q�ƅ�x��(�c���X�	Zy�fy��d��O��D�O^ʧ�^CfC��f�<��Q:#��D�'RJ��?)�4e4ɧ�)�9�T���R�g�X�x����)m�a���!\^�P�ʼ<�'l�~�䙫��}��"E�H�y>�b��Ԟq�(|���?���?)�S�'��򦹱�H�"�~���V�_H i26!�5I��%��ٟ��4��'�~�K���A��?��
bC�QB.�A�D-_�7-�ݦ��E��˦}�'����?�AsW�X��	I  ]����p�T�k��'���'m��'���'|�+�vTQ���4L;] @��S�ġ3۴Z' P���?Q���䧊?����y���G�(媔��7؈�y��S�^���'�ɧ�O�zH�V�i��dR�>�,i�աGȼ��g�A�󄒖sTlY��y���OR��?)�������I�O���� B`�T���?����?�)O��m�51�j%�'2�-{-<X
�l�>bVp�@�M��'≬>i��?�H>��D@./Ʀ�[7�K�*�5b�!�s~�n��&��5���Þ\P�O��)�I�\�+՟|;H�X�̓%1�D�i�2�y�,�="��@��ھ�X�
.�REu�8����O�����e�?�;a� �t�дAG�,�qG\�����?1ڴu�V�M_����Ĩ�'̊J��	�#�p��uA̖!��� �O�t��m%���'Zџx��mT Ux�$��Ǝo�& �!=?y�iS8�� �'_��'��d���<��p�Ù3/!MS�Ryr�'ϛ�(:���t�J�VP4-F���t���ɬ"�)؅հz��'&)
���'��I'��'J�Xp��<t�h-��KQ���E�'���'���4X�#޴ � �r��W����U�@:D�ѰHK����`��˛F��Vq}�)q������������v�ӓ'A;��Rei��j��xm�@~2J����I�S�:��O��!�0�,�VD�*25�bB��y��'z2�'y��'�2�I��*.��!��K k5���� }s�$�O��d��A��On>!����M�M>Qe$�k���N0����T�UD�'@�7-�ş��Ƅ@|�7�'?qe$�G�? ĩY�KF0,��q��	�|�"��s���?���3�d�<���?����?�EZ�$���"�%
n�jT �7�ZX�����d�Ҧ�@�ޟH��ǟ(�S��M��%�ip���P#h�6���id���I���d�O,�%��O�����#1���g�œ=���L���}�X a0T��S�\?�B��&Uf�����GK>���@�[�I��H������)��yҍ|Ә,�P�
-@D���+Ռ)μ JЏS	J��ʓ=�����L}��'U�AI2Ŋ�P�;%N�>n��.��'��D�e�i��i�KQ@��?��U�D��h�;oB4���������z���'��'���'�'f��=D�h�䐽��]�sH�/;��%��4%���/Od�� ���O^�mzޡK��P̺�H��N%~⪡y��ʟ\��O�)��-oZ�<Q2�%��hÔ�D��J�D��<A"��6G�@�D
,����$�O>�d_�i��X	0.Hp���CߢS޲��O��D�O��?�&cO�8�I����5�� +��9��ʞ�D�p�CTz�	ܟ��O\m<�M���xrC-!�����L8!��ק^���$ߙGp��x,[=B������@��@�l�D��`a�=+�q����=V��$�O��d�OV�d%��S�.DK�(t��D�f>����m���?�&�i*�b��'��+|Ӡ�O�9�*��ł@�[�Uf܌s�B 20O����O��D,Obn6m+?��^�j#�'[,:��%�˨G�NU���%x�H���*�D�<���?���?����?���ȕM����2��B\��C��[���B��1�Ԭ�ҟ����@%?����g���ɗ ^֜B�A4_�,�
�ODlڹ�M�ƛx��$l�nh �$�FCX���� �*�҄�c�F�t��Iڋ��?�n<�d�<1K��.ѷ-˓���$R��?���?a��?�'��D��I�#	�ПH�3�D�x����
;H�Z��Ukk����4��'n��V���J�O�6T����j#C�d?�!
D� KNQy�vӊ�I�L-��N���ȐN~��Fݴ�B+�"`��P�� & ��?���?���?i����O�f|C,[�0����I��C2�'��'�7�(pI���M�L>�ը#{)��MO�,��!r�I^]��'�l7͑��S�+$,<l�y~«�Fy0ɗ�<l�ԵQ@f�A7���<�q�|rV���	֟��Iȟ�p�Q< �,���:�j��ß��	`y�ohӨ���h�O���Ov�'v)^=4j�U���E$\�t-�'4�'��j�OBO��W����i��@�ִ�a�˄s"�xe�O�3r��
��Cyy�O�����1��'�z�Rq�*Qt #k�� ��p��'x��'����O�剭�M;S�Z&>."��m9W_�ݰ����`����?��i~�OF}�'o�*�;qgr�z5�A�g�i��I��R�'�.{t�6����W�8��剏3��u"�s�wB� �N�	fy��'�B�'���'p�[>]b����[��I�۝{^�d{��C4�M�5EP��?����?�L~�#���w��d�4 :R�ر�v��C��'���=��)�<<|6�r��c4���)�԰'��#�.�vh�ěB�	zE��a�IHy�O�Bl��^"9�"�����T�g�!���'���'��I��M�rF�?����?��m�jq ��� D�ˆ��O\��'��'�O���J� @���f"��g�<�#W���Qu��?�΁{�N,�>�BN�ٟ��!&��j�Us���m	�I���I��|F�D�'�l����h\ɳ��YG�$%�Q�' �7�RS���8�f�4���H6�c�U��Uf� �'��<�ѽi|�7M�٦��E����'��x@�$��?�G�*BQ��k�� ��lCSg�S~�'��i>��I����I՟P�	� ���kW��z6�Ջ��K?6pD�'9t7�VT^����O��d/���O�T�pB�rd��흯NC��N&g[�Ɵ��	W�)�iHY��CQt�a�mZ�d���ZW"^�7K�˓k����V��O�,M>�.O������|��xb̒.D��)#W`�O����Ox���O�I�<�G�i^�#��'{йz1h���dz��4t'p���'z6�=�	���ě�����M���,R��)��I�Ą|�c�ɧ*i�H*ٴ�����b��4��'p@�����[��U�ȃ:L��e��k�����Op��Oj�$�O\�D!��� =��`�'��D���A���� ��4�Ms���|Z��MA�v�|bK�����/�3sx-��&Q����Oz�q��)6v��6"?�%�?MvVdTTbU�e)��2M0�
T��OJ�yL>!,O���O���O6�W`W�b�lz�$b�n�׊ß���Fy£w�(�E �O2���O�ʧn3�����N�E<�8���$����'d��?��m;����P`�P�҆V�t#J��蚇[E�TJZ�In3G���Ӱ3���
i�	�E
z��N�*��Lі,N �����՟��ןX�)�Ry�xӾ���fC�H�<�'jķvYP�a�⁕&l0�Xћ����w}��'!D�+a�'3��Hs�(��p���i�'�7��q�6�2?��ȘKF��)=�T��!T�Se8��L�U�
�yrU���I����ݟ�	�ܖOT��R��{aD)s����P��2��|�ʡ�d��O����O4���č��ݡn:!�����E�q�0�	�%�b>��e�⦽�S�? �ih�C�*��!��9�$Y�6OP��CmO��?�S�)�$�<y���?�
�$XRy�'B˹kJ�ygې�?���?1����ċŦ	0��៸������E�	����'́Ih����)KR��?��I�M��i"Ox�`j
�i����U�_oh��T��TQ�ʝe����wI�}�d�"IJ�H����0H� Z�,G':J�Sj�����I�������G�d�'�"�"��+�L���𩅢�2��+�l��L���'>7�.�i��dIH��|a�'ƢBL���a������"�4n�@M0ܴ��!l����LB��3����<���atȚ�u�����,���<ͧ�?����?1���?��¥ ��d���r"�8y�C���P�x����	ß'?�	#&N�� M�mȚ)г�"nM�O��D�O�O1���1��I`|�8)e�C6`�S��ό�Q��<��bG�8�t������1x� �x�h��
c$�u�_�d���OR���O��4��%�FK�w��E�.�bls5�>-�i � �tY�gӞ㟼��O����O�Ll�B��QY�M�3MY6Hy@�S��Wc^����' @$0����?Q�}��;|S��`T"y�
��! ޴$�����?����?a��?)���O�t\�R&�H� z��[�\�Z�s��'dR�'l&7-�y�S��M{K>apĜs�,AR��8fy����*5�'�t6�[����¨>�@6-!?Ap՜F@>\9 �&6�1Y'��cֈD�T�O�`*I>�,OH���O���O����E�i=���c�Y2���b�O,�D�<yҺiq�"�'mr�'�sU�'��.|�6��d`Ƞ]|�d �OZT�'<�6-���'���H�ET'(���"�(B܂��������F����4�D�;��x~�O:��U�W	y[�<�M ��� �O4�D�O���O1�Fʓmk�FMχmB���&>��a��Q�x�|y���'mr!}��� :�O�n���،I��\$|(�1kY�L¤9�ش0+��oʕw�ƛ��Y!�ܣ}/�dk�Zy���h�a���>,���sF�"�y�^���ʟd��蟬�I��O�R��%C-ngR�!c͚:" �x1�lӾu�խ�O����Oܓ����S٦�]�mŞ�����2<hV��b�łq~�t��4F���L/��7-b�0$ڵ	�8��$�zt:�`�&o�L���S�aH�CZ��oy��'���?����	��,Hh��� <��'���'���MGf��?���?���ٮ\l��(t,��o�t�ˆ�ۯ��'FL�m�V�xӺq'�����c�r1K�JiSP�#�<?A��-����CD�$��'#���䕤�?���ܨv���U'�)2(�7�� �?���?Y���?Q��)�ON��]7�6(�$I�*�Z�bQg�OTMn�G�&��	��Zݴ���y���!U��@q� ';'�8ʁ*�'�yBDj�.lZ	�MkV�[5�M��OBࡐÖ���*�Ӳ��O-/�P:#�^�%�<��|_�,���l�I����ޟDk�K_;��!��LQ������	{y2Ba�z�����O����OΒ���<
�U�޾2b`8�g�ˈO��)�'t�7��q	I<�|C��z̚�d�J@fhI����V�>X"�I6����b����&�F�Of�B!�H�L�X�B	i�GQ�*ޞE����?���?!��|
*O��l9� �Ʌ 洸���J/P,��� E�Y�I/�M��"�>	v�i 7����y��o��S������q]�TxDN��a9V,lZN~�1@����'��O\w'�<G<�ÑD�9:��S"��y"�'z��'R�'1��I�?'�|s���rNv�1c�&r�`˓�?ѳ�i���+�OZ��f���O�8c�gշQH@�s&3���Э	s�Iןoz>�r��]�'K�Y�Ce��4��|YU��?��"��V�`H�����U��'J��럈�I����	lþD�#�!p�$�G,�.s������Ė'�P7-a^����O��D�|Z'-L�a��k-��4�^��	�o~"�>��i��7-�n�)��l��n�A�U#n�8���̲L�w�LX�V	a(O�	�?q%�(�d��e��ha�/�6 9F�8�	yT��d�O��d�O���ɷ<�Ŷi[����� ,H`�� 4e2C΋k���'�f6-#�ɞ��d�O�1&�F;e@�BCb��#<�å��On�$7.6m)?�;eh�z��&<z�R��� �8�:� �I�6K~L���$�O�D�O����O>��|�tp��q��̈����7�A3l���N�2�'�"���'i�6=�0�*�n��nx�@�j�#����O��d)�󉏑i�07�w�D"u�� �>��CK^�vX�7mv� �1�<=���UX��}y�'�RHk Ȑ�l��mh����!	���'�r�'k�I��M�tD�6�?i���?�@�Z�fr�����/<X(����'��듖?��8Y�'���k7���>�\D����,9<Uq�O�XR)M^yҒ�醞�?����O�=c�	ð�\�(��@ Hjp(J�"O,А���.kL�Q5i�:l�̹FC�OZ�oڇS�$%��џ$�ٴ���y���g�湠U�^*;�l���@��y2�X�*f�i�h6MX�^<�77?�F�͖	yp�)�3)�l)�)�>R��$��㘓O���H>�+O0�?yf�O\.)�G��37U\I2�`~�Kw�Xz5-�O\�D�O��?�zs䖻U������W���� ������̦�xݴ���O9�B� �A�2A߃�(��P,p�j���i	�,d`˓n� BѮ�O���O>Y)O��*�jJ	!t�%3�ꂿ'r�����'Q`7-�������4ڜ��2���"�qB敥5�~���ۦ��?V�D��۟��I�<[�1�G��2 3RT��cL�}ߖ��R'Sզ�'�Zk�?��%��TꀉT~�z��;d�j!y4M��ar�%x$�ߦy�f��V,�Q��Y���Y�YV��:&�5x����O��uZ��8��԰UmC���B 1���_)\/dL�e�8(-,�uCV�s�!�D #�ͭ��B΅ �>��4�F.x��`�eV ]�dx��j�-^_2T"6
	+@��r�̀
�NlB��A l�����	S*q��q�(�&������<LΔ iFH��o�z�)�<�Dpc���x���[W*�:��iac�2X�Ā)�J[�C�Ψ!�@����q�R^@�us�۶�Mc��?���^��t�����Of�I�@��С�vm�}XSF�o�c�x�&D;��ҟ����QS��2 g`���6a[�`�b�
�MK��Jؑ�x��'�"�|Zc�4��ː |+
�I��)��O��B�{��'�b�'�u=�QJ�� ���T�V�A@\�RfM#���?9������DL:an�(�7[
 ����Ԥ=s�?��'���'y�P��3BN!��t�N�w�LQP�lO��ԧ�>��$�Op��2��<���a}"(�(.�К��+Ae}��M����O:�d�O��
�l91��t��J``Q��L��xz����.чR�6�OؓO�ʓ7�T)�?QcZ�䥘�����)kӤ���O���t�q4��$�'|�d�p�M�� �=`��9#  ����Or˓Io�Gx�����,۔7�5(�!*Az��i�ɮ�jLٴM;�S��ӆ����-����g`�����/V���U��p��p��|&��#��,���1%TX�ԅAFnӂ�Ñ����q���I�?Y@O<�� on�q��(��#n+�$�� �iV�����Ο�pQ��k����EѨ]N̔2��
�M3���?9��r��5ןx"�'e"�O�,q�(4YMXup�d�	&KFTcS���: �1O^�D�O~��#b�$�� 
.�E*@l�T�Ul�՟��d� ��',�|Zc��ic��}b6����)y�۬ON�J��O$�d�O��9��,B��@�	�I*���h�k�F�"P�''��'��'&�I�c�4ڢ "~0�k�0�`L��"�	ß��	���'�1���j>�9�*Ю\�m��� (���>q���?AH>y(O~��'Q� �"O�\+b	����1����7)�>����?q��?��AL |���?��'����Ց`n�u(�nC�TW{ߴ�?�J>��?�e�9q.�'�x���i��E(��\�D���If���$�O6�d�O�<cB�O��ĳ<y�'�lu����?1 ��Q�ϟ�: �C�x��'� �*l�y���a;Po��]@���UG��%�iB�'w
h���'�2P���SzyZc-�����OP2�:��,�ƽ�ߴ�?�+O�����)�ݦg_6d:"�4���2$�Y��CT"L��'C�	�?	�'G�I�/F�FO�f@"�	�n�����O`����)��`�BQ"r\�����D/.� ����\��M����?��@�Μˁ[���'��O���a���6��$�}zm���iS�'X��#!�	�Od��Or؉"��N��P��"%H`��%�֦���;AVĺ�O�ʓ�?�L>�1[��	��b71��"��";W�Q�'�̜Aї|�'���'��	 ���+̍?��,1#�iz�t�`&���ĩ<������?��y�Ĥ��d.zf�%��J��|��T�?�,OH���O��$�<!.ҧ/�	̏+��eZ'P�,+�-H3@���&U�`��R��d�I:Wbx�� .�ͣPJX4�d�@���3Z�.��'���'�bY��8ɔ��I�O���i &t\٣#�PC"�J'�ܦ	��I�	���! @��=I$��<tYft�be\6Ț�Dʎ��	ڟ��'� ��D�~2��?1�'n����j����"C [o>آuZ�P��ş��I	
�@����?����>*S��sӬ��\q�|�pr�ʓ����%�i���'R��Or����᪂3w20dL�pZ����I���Q�	��dA'^����O�,,��H�b���6A��A�ߴ%}�(!t�iTB�'���OL�듸�D�֐l jBv�h�´H�?Xj�lZ�a�4Q�?Y��T�'~6ٱ �'9���/B��(iB`aӸ���O��$��YM�!�'8�	ޟ��QU�\�5Ŋ�U��@���Q�l�,�>�LM��䓪?���?�s��j�@S�B��lR�퓬mP�V�'�Ku��>�.O2��:�����$^�	,�A�)��ԅ�>i�����?	��?/O���1��?������S5m)�B�g�J��'��I�$�(�	⟌�Wj�*�D�Z�Љ� W,j�x=1�h�Ox��?Y��?�-O�Lj�
�|�V~�0�!Wb:�LI�d���Ŗ'
R�|��'�DR��$�W��qxq���t>����(ʺi��I˟H����H�'g��'�U�K�p���lD^�A�  \'��m���'��'՞$��')�'W�6�H�_+L�L�� ���@mZҟd��iy`2j�`����k�WM�E#I�C.��J5��f>�'��3e����C��s� .�� �[�N��cf��?X�� �i剡*����4R���8����D2-,� ��(Rh&,3QB�(|>�VV�p�S�T�I|:M~n�Y�h��5��g����%ć[L6^>?�����O���k��i�<�O�h�����D*}P�����< ��tӶtk�i�p�1O?)�s%L�7���Y�ں	o��Y3e��M�����Tc�)zI� �s��;.(���`B!XH�Ԯ�ǘ'�<��'A0������p�Ud*�F� ��-�"oE�Yo��<	uMCy�ͺ~����
�Nb�Ec'�X�g�L�rύ�rWh�j��ړj��?*O��D� �f���#�nDq�*ðZ��)�2N�<i��?y���'��"��U1
]�e�C~9+��.X,����3=(���?I���?�,O�Q2���|�¥ܸ;᱒c��\l ��Ԣ_G}R�'�2�|BX�,@��H��8w�I>K0�}ai__��!�Š����O���O˓?�������}B���L��*�5J�� 6�OV�O(˓K\T�����7U_ҙ�F�[�]��9�g�D��6-�O�˓�?I6��*��)�O���kܹe9`	�H�.���;�!�>�']b�'���E�ؓޘ���	�J�ђᓪ ��YP�F�FY�,���0�MC^?a���?�(�O�`6AOl|$d	�
�
#���D�i���u�dP�I,��'��禁��0|L�M���Ӧ)���!��Fɗ�|�7m�OP�$�O8���w�i>qk�E5<�B��B"�"t�������M{�)
��?9�����:����Ã� �Xj���j�pTcD���M����?��'A4��(O�e�d�����B�	�c�r8慯Z��d�<A�c8%S�O�"�'���;���[�m��K^���c���7�O��a��_�i>Y�	��'���S��,q�:���0
�n��r�w��d�	C��d$�$�OT�D�<Ab&�'HkzY�&KC&s�n%*��C~}�xb�'���'���ɟ�I���(�J�\I���(�'xl(�b�g ǟ��'�r�'5�R��p�����$�;�p�b`.� ^S
�����)�M3/O��ļ<9��?�f��q�}���[>i ��1(Z.lΕ�a�i���'"�'>�th��l�$җ~ǆ(Sh<|�����ն!�No�ȟ��'�b�'#�C��'�U:�i�#�ڍȗ*�)�����4�?Q����}!��i���'�b�O�NU���N�]Cy�U�[3H
PL�>��?I��u�'f�qs� ����³M������Ŧ%�'��5#0�|�>�$�O��$韖�קuW��
嬄1�nW�N�l���<�MS��?ye�\�'*q�D�0�8?�&JF�%��8yP�i��dרwӢ���O�����'�I�9��`P��A����`��eְ,rڴ�t���?i,O6�?��	�(��%$��0c�J>XB\�Kݴ�?����?	�����ey�'�$�r踨Ck��T����ڪ|ÛƓ|RD��yʟD�d�OV�D�5���e�L`ҹ��ʗ�+F�Ilޟ,��,L���d�<Q���D�OklA��4���<��e4��& �ɭX���4��ɟ���ʟ�'�$Ű�V�$�irÇ�.~��!�&�����O~ʓ�?�(O|���O���[���1��Zְ�q͘�4�l)57O���?���?�/O�����K�|
�+�Z��(L*9��#I�Rʛ&X�L�	Ay2�'Y"�'�@Iۘ'�H����)��G]�4���'oy�B��Or���O�˓H�x���^?��i��L�[�=9�� "�z�Su�B���<1���?�y����?��g�����V���Y3t`�4�`1��i��'�剎�������O��IY�V4`���օ4U���v����:��'�B�'��N���yR�'F�GR��^���a��6E� =a��@�՗'��q{�iӨ���O��$䟌=էu��׃X4�� /�a���9r4�Ms��?y��Bn~�P���}ōM�
Ѱ��oY���A�禽����M����?�����FS��'V��#P"��B&�<o�v�Rdʚ*pQ7�c��$�<����Oh&!7D
A��/9Q�D�@�'Q��6��O����O��S6J�P}�_���IZ?��Ƽ��dQG�̇aVb�s�IK̦���Pyb��8�yʟ��$�O�$�<��Q �/ƈ����`�`�xl����� ��d�<A���D�Ok�R�v�<���;XY2�{0���Q��0 ��ß��	����	y��'U��3�AJ�X�l��K�B�@��&ªs�����O���?1���?Ye�#q!\d��D��dV�C�)|��\Γ�?A��?����?�/O�� d
��|re�!^�����W���$��Ϧ}�'eRT�x�	����I�oe��ICeP]Y��>��(!A������՟X�	�����{yBJ�<7�N�'�~��0:+�cЬ�<IZ]; eN��M������O���O�y�T1O��'�kԲ��b"3���Ǎ�M{��?I,O�����c��'���O�A��nL�D"$�c�H�Mr������>���?����Y�<!����D�?U�5�ڸ]fY���J*1z� y��8CJ�hg�i��'\��O*�Ӻ�Ԧ�= `���"��@�2���EAǦ��I�����~���ϟ0�	a�'j���ǧ��"XDb�@T&ߠel�!��T	ڴ�?Q���?���VB��hy⃆�o#b����;�Dq(kU�&6m��4�$��Οĉ� zAH�l�|$�s�I�  |aſi��'|�·/T�����O���6[ �SCnO��j�{��͐H�6m�O����ORTC�0O��蟤�IƟh���G�o�;�i �W���'� ��M�� 	�ÚxB�'e�|Zcnr�3�IĊ�
E�cs�M��O�`N�<))O��D�O���<��%cX�����&
A��c�D��0��!��O^�O��$�O�]��)ثv�:�)D��2zʦ������<���?IO~��KQ���)��d&bE��B�옊*�g��'��|��'�"b\�y�, 3|���T!N�{�2m���݆up8��?����?�+O:��`o�f�8C�U��i���D'B�qE�D8�4�?I>����?��!��<�I�,��2PMl�[3�޶FAhy�Cm�0�D�ODʓ^u�����'U���]�M( Ă$T����=?�O���O��@�*�OP�O|�SA=��X$%�|���ը)�6��<�jɬa����~��������u�!.�	XF��#lr`4���t���D�O|�	Gi�Op�O*�>� K�,r���R�\�!�N����~��eZ٦-�	�8���?�0K<Y�[Z|h n,l'��W�l��xsv�i�nM9�'��'���S�?E�!W#ƒ��dFv+��o�������HyCNE���?���~2��c��[Q�NG ݺ����'����y��'���'��%��+A�ya@��
��|ZΉ���z�p�$�/Y�,�>A�����a,񰴑p�>V�ڜ(A��q}RbE�/��V��������[y�-¯ r�:����I߼���ÞR���O7�D�O�d=�d�O��:�	�h�rt"�1D�P`��a2OJ��?����?!-OȠ�Ta�|���"F���ڐ =���\}b�'�"�|r�'�R���y"M�5F�y��O���P�����9����?���?�-O8<���J⓼d^�Iud�>=#�Ya$`���Q�M3����?9��bHۍ{R�I2}����ԢT5@�ҥ�׏E��MK���?�.O���$D~�S˟��S6}>R�
��\6|X��g5vW�K<����?qQj�<1J>q�O*8A���<W޹"E��	k��`�ش��I0a��Uo������O��)�u~B�עp�f�YQ�v|%�֏G��MS���?!��9�?�M>�/�p��t��9[�m��4>����K�I�p7�[(H
( o���	�����'��Y+U�W�
��WW9����iv�V� 6O�OH�?��Ɇ^fE3�_q�}yi�`t�$xڴ�?����?�g�pL�����>9�e��B��`��* xq�M���?�����'/��'*<�`�E�qh�qA����brӺ�$G�:5��&��^�'�� F'�z<!�F�5�h9L<������O����<��C���'�Y�$�~��Z�KP5q3n�:�?A���?Y���?�O>Q��~B�F�b�;�@�/�|Z� �M���s~2�'��'��ɝQo��O=��V��(��y���Ҳ
��pcO<����䓑?�{��P�b���;�!!�������O����O�ʓy�x��W���!�),��#��]9#t���+E�,7��O^�O���O݁1�$WIp�v�)K�ԠRH�E_���'�rY���⩋��'�?��'_I�	��U?Y��#�)��rz�ɠ�xR�'����O4��"ऍ��)Y�z7����Æ�]Ubd�I��0���D%?㞄Y'�*C�� ��[vX��9D��sц�Z�WQ�,����U�D�Q��TpV%hb_� <�x���cC"Š&�W�8��������I�4`�Ƃ֒ld�H2�)]'=񸱂��-hP��h��?e��%rS,�Ќ"F�݄@< (�g,X-)����#tc�����i�VD������3�ٰZS(�Ie�
 ���rA�=���'��'��֝��x�ɍiX�Q����=��,i�y\I��ǋ*
�����9b���;���?� ���֌b7���<3th�"$��(`��Y)6��:�uB@e�2R?4�ٟ�hDy"���Z܀��]�	�)�	��~���?���hOP˓:� g�#W�D=A�F�
[����#[^t@A;GE����o�:���E�)�,O2��U�����!��U#�J�Ȁ�8X�L���Mݟ0��ڟ���1^ܐ�	��,�'p򤸚�ǉA?�}qC��Xj���+��f�d)r˘ �L(�ϓN���P��\3���݈��"��j�"5��\��X`�M�rx�:5o�O���84px��(<5^���n����=ъ��M�O�|������d,r&I�]�!�đ�o�t{RL��TOZ��@�w���H}B[�蓁H%���O2�'F�\5i�ٹ!���	� ?g>�-`�K�?����?��ԟr3l����+�|$x����i�t�~�꣬�1O�	�P��}�Q�x�dHCŠ	�"�&>�&>��!NJ���R  ˷y8�`��>ʓU;���(����_�O����X�O�����<���;<���F%g�z�І	�t��	$�����~��a[����SR�����<u��X��П��O$6����?1�a�hm�"�a��|� M�8�ȓvo۫JG� k���9������I8��O� $:��ӻH\H�u�W�0;Z��p�@6�ڂ&=N��i e�#�֔���,<q�w�Q:G�1�J	�_J1����f��s��'�Җ�����OL���$eB̸���©D��)��"OX4Rg^7-/���r���`�Hu�����HO�ӷZ?��Ca`� \�DۥC�k^(8�����k�%�S�0������I��L�Yw�r�'s2�q�J<=�ȑ�nC���5
�'<9xT��,C}2��׊=O����nK�`yxc�ĽDn����O¹
3.N #I"��be}X��8&�8� �����(0��Oȥu�'=�Yy�'�Qq8Q	�h�kׂ��y2������@v6��gZbr���@.�S��V�����:X���(]�]P�(F�'?&9��$ѓzA2�'���'�d���'��'>���V�'L��^+X[��jr)�*&,��0U.L��p>�e%� ��Y�䬚02���+�����-�<E�2��$�P���'���bB4_ ]#7�Q;MF��pp��B�D�<����?�I>�O��h��O/�&`!��Dʆ�
�'К��T�8[��C�O�C��q)�'�7�W����'��M�5i�x�D�O�˧ ��!0���V*x �w�ϕ`z������?��?���Ǖnx���|]>sGS�$��hqU���P�:y�v%�B��ZDF[�>"|jc�СQ���t�1�D�G�' �p���P��Lp����|�r�Q';r���(�6m��L��̚��?A���9O��*"�P)F�6����l��!��.-|O� oZ��M[��,�`}��`�-y��=����:�luϓO2*\B7�݃�?�����iݖ����Or�$���G�	7a  {a�h�m�"�Bn�F�&��'���?���\b<��,�:�Y!7�Q+�9�e�*f�ɧ��R�B� b��X�Ov\���+a* 
r�'���'��OL���IG(@Ud�WYd}�4 c9Oh��%�O $�T	��b�R�qaZ2)iٲ��ɞ�HO���V������h����I�Sot���Q	�(R�)����%JQ��B!��+�t�ѡ"�<[��[e��z"�ц�X&�
�*��͑S�ْ+���r�@��fй<x��) 6Z���ȓ��%H���63�}y�X�Z�<�ȓ�a��i��^��Р�) : y��[��H�T6꩙f�Ġ_bd�ȓ~>��7�� �@�9��	�����
�L�R�ȋP!��95/��8H��r��Zc�ߐ4��t�G�.�j�ȓfn�@��!Y�(���t�X��ȓj׼@!�Kߘ"�r�i�`YLF`��,��� �N� q6��P1H�f�����2C֍��+G�g�n�pӄJ����C�F5+A��b�!�҈һJ��ч�9Y�=��$		%�5�ׅF�<Δ�ȓªX��&0�����^5[��ȓ~�b�R�g�/uz��C�A��4��B,��;�O�l x����S�:�lh���8P���R���� ��'�`H�ȓ;�d	3c���;~�DYE�]�XX�نȓ|D��]�W��`q�oj��m�ȓ����\�
���SS���u��4�ȓ�M�� �uvv����x�'/0D������)r�h4�1j�0?�� 0!g*D��� �8 ]��%��RaR�J��&D����L�-]G���e�O��M2g!$D�(�늦y� �����)p�ps��!D�����
[~>�āݎ���5`4D����O���h �Z>pVr3a�0D��:š&LV"�Y`��\�.��@�:D�D�D/C�%�� ��W�� 8D���D�0$|�
Ԧ�5U�$AX �(D����c�*�L���<Hg��!D��%O�XH���q�84+��1�"D��)ЂΑB�|�����\$�a%%?D�� ~dZ�F�0N�&��j߇I@܋"OHH�%��֌��b�S�|a$"O��Q���>rhy��ǐu��˃"O.�$U�6P�:׏�/,$
`"O��
2�G�#b���V!9+�^x2"O����*Lp����%t��}
`"O��P��81��Ǎ@�L �"O̝RD�!���d��<h�8�6"ORh��$�%;L�ꎕCn�ͻ�"O0��74sF�8��CXiv�y"OP�Qt��>�F�+�
��\ �h�"O�zuIH-����^�r�l��"O�L�f� �:�n�s�?�	�"OD����EN�6�pg܂<�q{'"O���Q�,��@��ݷ�r!��"OR�0��
Q���ے�܋w�d92"O��y��\/w�,�0�Z)G!�9�e"O$�0!�� �M�FH%N$�sF"O�B��ÝW��b3m�O�*ԋ��		|AB�,��2~�Z�������59W4B�	�OE8I�"F�U|�(D`\�{�˓�Fѡ"@���S�O"�=;wLE�j��P�fR3["
x��'�0�أ,�%RS����,]�FP*M>��.Y�VpjÓ?2�M��Đ�Mp i��fI�U8E��I�;:�m�t�D�_�"���)�~�"{��W�H�^D���)[��.�y��8揟'�B�E�Ź$��}:���؆5����� ��
�K!�$F�&*�Q1�,�=	�*�	�	�7�ɱ,�4���'�e�)�'SI�<��*E����fJ�n�l��ȓ=f"a��7'���&Q�^�ܸ�<��P�Z�̘��	�~o���!�֓���V��}��B�I' �i���T:9m��c#�]x	�B�IN��q�i &?�L�X�ZG!��$�����D�.$<b�O�!�$��#��lQ������3w!�d�ji��+��,�X�`�o�,Q!�dۜ�z�A����E���^&HI!�ē ��\�e�0X5z9`'/Db�!��yĆ���iڵ- ���4~!�DH>�q[���G�J�1RMط%f!�DM�[$Z�)���>�>ј��&eB!���|HDr�&V#,�h��E�Q�!��L\���p)�)h���g�4�!�:N<�qH�Zoh0�3�Gr!�+I�bdXr�X�n�F!��@.�!�dۚf{�4�P�D�.�j����!�Dן5m<U�@"�L�feX#KS&*�!�D�@�p�Q/�2c|�h�B	�rz!�Ѫg
���B�3uy���G�:(w!����r�F�zs.�w��7F׭	`!��cJ�!���*+�� E�3]!���@��%�I-��t���T�d&!�dH	p\�2�@�*!��1���t!���']��J��N�4�cƒ�Y9!�d�C���".���aTFI�H!�ݼ&�>��&��=S�B�;Pl���!�$�%�*�#�>~^Dˡ��F�!��Ɉ)rdQ3�Y2l�����Y�e�!��&Jв��Ή\j��&��&7�!�d
88遀��0¤@��U��!�d�2�������3QH��"�n)n�!�Ė#D�!ʵ)?��r̓8`h!�Dt�zy:��ˌY3H`81L�vt!�$A �n`���Q�` vJʴNG!�� ��B��7nD��� 	{����"O����J�d�����N$��5"O�lIS�Z�i��'�[�Z�,�"O��rv��+-|Q&'9D���"O"��E��\&\�FEռ@A�`�F"O
�X��)=$f��U�%E:-�"O6i[��-#yh�Z� ��nԠ]��"O����	�YO�)�d/@)��SA"OP9���62��;s��
`�ִ�R"O��b͗1`��8kQ�%�@�'���т]|��
"�Ly�W��m�F����Y}����<���&�����O�u���U<2���)v�F'v�X�t�d	T�����ة��'V ܻ�%,�>	�% �N20z��aH����������c�Ȑ:�ʘ+T'v��f�Ƀ5X��p���G����O�yed9Pq��ԮR[�4�*Dqb���|���aݸ0:��@c"O�d0�*�Bm���d/f�r#�'�:���"�4�^MB�j��~҉�W����b"���f�N|���(�yaH�� !��	ܦ`G)R}�>p�H�o�,�uG 6��S�8��\��)L�/����|�b)M��~冀N��<Z3�]�8��`����0?�a�Uh�u�듃.��v!V�k�f�aA�":3.J�1��A|v|p��$ �#�uI-/Z��sXY�\4D|��1Lp������H��8��UE@k�n<�pFE�6`:�&Q�U���v�'[�}1I�Y�y��߆f��k�'䁛�Q�7*�ljbDA���S�&�Dٙ�'Ͷ��f@��9U� �1Ȗc��q��cd��a� F�+q�%Fⴵ�ட�Z��[.h��˓� ������@���y�g�1�l{f��i��� T�J �p>A�@�j���L܂S�d�QĄ�
��i���,ry:O�Y׮��,:AA�9̈q�L|Γ_�̱�$�!�fX� N˦Z�R$FxR�M���!�gAY>u´̲"	���?�'E1`8�f�c�9Q�턅�,d�/�� 2�3YNYڤ�2Od4S�
��st�&���tA�BVe.pX8C� �,B\��F�{�J?�O\��kI�%�ҭ:SO�7��O� :!�dYI��O�;����F�_f����,�O��1�A@�-l���֟���sRZ�L8���2�.P���ç�߳LGaybX ���G�#����*���"����E�� �]SZp� B��RXx5nL�w@�	7K����1�m�O��J�B�5��� D[�0 �"�$XA��dHZ�aF�����BӒ��'V��Θ�)���ǌ�_T0�C�����Y9��7�z��a��3O�k��&(k���̋�H[9� A_�_�M�6��U@�Y�4�x�i����x'?��R�v�1x��#;�1���1IjaZc���� ��`*\zr
L&MіeS����#���hR2�"(8?1���+t$eM@�)��1z�h���496�B�'������a8�����ȠJ�i��O�B�X��ŦN�Tth1�G�#\*��V`��M�F_���dY#2��sbR:�:���!Nϖ4�O��q�&Y�\x	��-Ռ5 b"�>��K�Y�jA:�L��v��iCE��F,�r�j���b�W,ڪJ+�� �ʈ��6��V&N�����-@.��J�7
Vtx�!�x��-�rOz.�s��r�M����$����O����h[$c0lX�N�d�<�D�S�d�&C���c�,Q�@�����D��dZ�x/��굨MH�ܭc�K�>y3�^�a%�`�djx��Z��U�0��b04��`�&z�x�p�)U�D��$e��Ӻ����;)z$  G� i˼��RM�$4�}�mH�-)Le���'T}I��֕Y����,����S*Tw.��2,ݶT&����{���)Oٮ�YnۄY��3C΋b��	�-�f4q$�o���0��B�/����iGQ}B`��3^2�ZA��rD�`�I܋�b�Bnțu��8(#H�(&ļ*�!F.hd�x��^0�(A�o�c�2x)�K�\����0`r��s�)�����_0D��X`ːt�S8h_�P�aU�ƬB�K{������'@�l�z䪰 Ih�Z@�[�u[�T�TY &ye���d�� ��)Hl2Jaʇ�H�����C�Q�b��@9p"��R!^��0ǒ�#��x�ЩH�J�z�G�>Ҟ�p��H�4*�-;�L�)`��?h�8I��!�/H_�H��Q:U�-@�ĸB�h��H<)/�H˦�)W�&}�&��"�d�'�R���&O*A�L�W�z�L0�S�R���~�l��s��y�=xІU�<Q���Qfb �q�_���[;E��S�.�\��xt	��%`0��)��R��H�T��j@��E3Qb
}�<���D. X��@�R������P����I�10�*q�m-<�'� �<1ǌ8�.9��+����t'�t���3�͆1��aB.&�L����c���!�ڋ#�l�`6��1j�j�3��'T@J��N7P�;2�M4f�*���DM�BT��8� �_n�Zsl��(L�O���w'S�8�΃VTp �
��� ��;c�B�M��rT��ԉ����s&.5؀b���Q��A��
ٰ�E���BZ��EO%_Fl�g���z�Մ�=z=������Y����Xe��\�U@��v�4B���|����ȓ)�� �Q�C*2�q'�6W�r4��VBHql�®�2��3tHJ���*~8�s�E��~���QҬ]F��i���[w��
�Q
��ݱe���ȓ*x�Lk��}�a�M� 1���ȓ^k�� �G�A�X���D4hȰt�ȓ��y�������X��۷
\d���$���ѕ\q�,u�v�^r�� �ȓTn�8�`��P�n05��m0�=�ȓp�j�1�腴��t�OZ<+�tH�ȓ�@��% �*E�:I�c�� ].��ȓX*,PG�V�2p�S�298@��p�����	ހ6������@��ͅ��`��dA�1(<`8�II)gfI��&�����AN��J	�p�B��ȓ*#F��tOÊW>0�3c��#(# Ɇȓd�H�t���:��n��j% 9��g���D��2���ϛ�R���p�Vmӑ���Q���P�jd�ȓ+��	r�ܺ�@�cኺ;pb���i��L@R&�����"ߤ���kTىgN�G�<��#K�6"�ȅ�n
@JQ׌A��Q;р�(	�d�ȓw�up5�G�:�Qۡ��lXb=��Eb�չ!�ƴwE��ʓk��} l�ȓ8�쥙��#	����.vذ�����9�-=T��bG 	LLh��ȓŎ�I'��5�"!H�"ЇU��чȓ"�e	�]��}9���h��	����Hd2!�(��o��>T$�ȓq��%�̖#������z+d�ȓck0�Sen�;j�Rү�9����ȓ[6(p;��-�D�� 4g�谄ȓT�����c�� � ���X0��p��{rn�@ ԭS����'U�!zхȓ|�̙r�V)|n|�Dj�)k����ȓ ��y�7L�H.�9B�g�A@�Y�ȓVHJ�z���˜�+�)A$ډ�ȓ�a���_���1��<C
�ȓJIJmZ�L

o@2�:P�-�ȓ&���b�:3��(S��h�:P�ȓ@��|��
��Ik2�c۞rb��ȓ}�Y8���8@,F	����w#R��ȓd��c��/OhHY�cO=5ΰ�ȓCO����*0��286 �ȓ4�a؅`B���pjC�[k$��ȓ5� ��,�&L�4ҶY�6#�Q�ȓ>L�T!���9Vr!�βxl��	�Dr�"��	��("�fY�S��	���J�h��\,7n��X�J6�RC��8�0!q�� ���Hم`U�D�C�	sI��{"a��-"P��d�7y�C���I@��~�l�X��Ӷ	dJB�ɋUn����dK`5t5(f��48B�	�=C� �q��7m`h���%>�B�	5P��YxG�R�^L���P)En�B��>�*�m]&�N�x�`ϴt%TB�	
 ƌ h���,%>��F�˥chB�	�'�L2a/%��4��I�I�&C�ɠ,���Q�	
������B�)� �p��޹T�R��2HO0n܄d�%"O�����;�*iȈ	�h�j�"O6咑F�
�c��+i��4B"O�lY��A�C>��@͍c����"O�4[P X/9��bg/��QV��"O X��"P) )Ҭ{#0�x�P'"OX��um�A�W,��H��ݳQ"O�9���>��F�-���"O�Y�f��8e�m��#c�6x;�"Ont����0�H�2��+Zz\�"OL}{b�G�t��"QGG��"O:���+���H;wa�Z8*�j���r����^�"uV-���7 D��%�I�!�ă^P���p����0`�1|!�X�~Xl�K��W N��r��S_!򤃠P�����&\=��`[�r!�)�^�H�M1)v�Ɇ`�:M�!���S;Xt���,&97F��6�!���o���XT����z���04�!��B.r���J8V�zŚ6AV!�d1
�,I&mU�8�ys���H�!�C�#F@��c �":�6�3b)J4v�!򤞋�Nd!�����`�
V�1�!�щI8�aHa��:��dz�*M�!�䖆Tۆ���̐+~� z���'J!򤑬ܬY�O�p4�2�H��J'!�ыu�BIP�ų1���&�F#!���z���)�p�\(p!��g|j��F�.��B�G!��?x)����:>����%X��!���t��2K����r�#Q]}!�R�X(��&�B�9�� �T�	�(A!��\�A�Qq7͚�W�~ ��n�-E=!�$W=d��e;o��S��e��mܘI>!�$э>I6%�$MtFA���G !���	zH\�*֔|�Y2�
G�2!�DQ�Yu��"�`�� i
pP��C!�D�<"f� �q!T�Y�A9���mE!�z@�;��H?k�� �5��A!�C+o|X��TEϯ���R�Mټ(�!��]	 ���kg'O:��TP ��(�!�$�]@��GG҉H̖-���>^�!�dV h �`&�X��`�pѢE9Q�!�Xw�MH� щ+�N�aW!A��!�$ߎ@
$%���]�y�V`c���<s!�dgS@��K�1l�1��iИm)�B�I'K�aiF��3��}cS$ӥ:�fC�	�y3d�S���Fz�i:�QnAC�I�6`1#4Ǘ�x);2aʥ1 C�I�+����� ?[���i�Ǌ0x�B�	�[)��R�G�@}�G��Qu�B�	�-�9x�gD�;�D��+�W~vC�8r�V�i='l-���4N:�<��a[0�C
x���d�T�C�̜�ȓ!�aca�C5�̴�T�\�2�܄�x���j��J$%04�ޏ�谄ȓE�h&���E�`��6'�B�ȓ`����\�|�*�"����Y��8��y��ԧ�b�h�j. ���}߮D���*.N�����7�@��ȓR��U��� ��q�`�Z*g�%��AE���G��u-8dY����x6p͇�Q���OG0?,6��P�8H���ȓb"���%�2��+ܽ�.���S�? �5�����[k@	Y�N�-��X��"O�1Q�o�#e��$ÍU9.��\�3"O��;B�ĀPQ�Pv���v�~,�"O�h�c�8g� ;��T.��i�"O��)�\9z+�G�3]���b�"O��A"d\�O���	�fŐ.�̨��"O6�v,�a�����,7�^@2"O*( fmU�8��
�jT��R݁w"O��FE�Hcn�����L�<H�3"O����F'~���"e	DN���z�"O<p�A�Q�b�`�7�@�ސ(�"O�)8��L'8���6�¹�`��>���Ҷ�G���	���.,Td�� �4A���Ċ#PD�ER
� ��I� Mfx�4
�:i��8��?R��<���T>� %KIC,;4�_
o:���$D��y�ȃ�lȨc�Ɍo'����!D�X�3A�,�c�Bc7�)`�L%D�ء��W�xLl��QN��N�)b`5D�샖kJZ_4��F�g&zdrƆ2D�����-hU�5��E�0���"D�"]�`y���/�y��m6��hO�ӨxA�Yr��-<V8�ȧ�A��B�
7��(�a	=BJ J�ƛXi�B�ɫ<�������~?�U�&KŮN�B�9Qu��at��4�ؙY��<7��C��<`�1Y&��X�ڨ���&�XC�		("�#7�Q�]�� � ��/�BC�	�6_4��0-�6UV%8saWX�LB�I�S�����E��QHԻIBB��b^F���'��y����?,'$B䉎r��"g�գiD��)EГ/L�C�I5l�xRe�i�P�����s�C�	�y����ӋJ�E�8��Bƒ�[mdB�I&� �0�)65�����P&ku�C�	�jY��W�[n��Q�L%<�8C�	�G�4���B�u���@��ֿ5QC�	|f4$���Q�D��wo�B�	!s�\��s��P�kBbֹ|MnB��� !�#�a���#'VS#�B�	�$bT웁�¦uV���'�FB䉛c���h��:^��a��X^B�	�s��*�I�rW�qP.�%S@(B䉬s��{��̻n�^����$�dC��!����VV�%sfQ�`,�*G�2C��B��d�ʲ|�,�'�7>R#=��T?�狞�9Y,4�$��fe5D�<[C��;��Թ��7&�� �ҧ0D��k�O��H��o
0(�P����<D��ca
�0v�4c�ϒ�
Xpk8D����O�!�^����O&^3���5D�tC�� �Hլ����&M��jqi2D�x�@O,C�*bJ�xր�A�C�I�t�^���)K�G�x�a�Á/B�	�R�#o�;rL��ת��G�R��ĵ<��G�1a�qB��ÿa����D�F�<) �:�6�K�gH�\9Υ+��H@�<�2U���sQ`J���@R�<��.Y# @A���z�i"�Ph�<9Ab5Μ� �G
?M@��w�P�<Q�m�'�raj��u?�t��e�<���T�B�B��&D�iq��I]�<aǠ�k����B�e���d�@�<I7�S"=�0�!Ì�:��@B�A�<� �@���>������dC��`U"O8 �D�G��nu�����=6.(q�"OjASFC��Y�0��F!�F��5��"OnTb�M�
I���{ �	0�N��"O$M�g�T>bzmK3�Ñb�� ��"O��9�ašPͨt��fu��P"OHD[6N�>�%i@��;
\r�
�"O�y+%"H!$�x(%A�z{0)Q�"O��h���\�.�hQ*�A�B���"OB��L�*�ڵYgU8l�Qٳ"O������2 |�b�F�%R��٠"OB��WI_�I�I��̩>����"Ob�ۢʑ8mB��M$?�B�i�"O�D� &�B1�"�mK|Q�"O��	G"_~�� go^
R��pV"O�xq���Z(�p�̌=� �c�"O��S����M��lR�I�#�����"OP��Ɉ n��%k%h�
��� �"O8ш��Q�p�^|1�Gݚ~z �y�"O�)r+�cjlX��G9v�8��"O��ٔ��j	C�fH�#p܍�'"O$�":_���E��F��|��"O�H"s�G����OĆZ�f��1"O~��h�1Mh�b�Մ�Jd�G"O� �T�¦)�&�.d$�:p(��!��7`Tc�\T�5!�F_�9�!�J�X���C�m��&�,����5R�!�������ϛ�y�2�1 �BQ!�ںZ6$101
�m� 3�K�r�!���D(��K�]4f�B�1.��!���-�6<&��J�V	���R�?l!�D�� H #U�O������eZ!�$Mf�F�[f�ɧ/�Fl�� -eA!�dř<c�,x��H�]��IUo4~�!�$؄
��uR$�?R�l���GUd!�$�ps�h���ܛ�r4+�L�kS!��0�t�h	d^y�!��,#!�D� ,�  �"�+%bT1��83!�D]�b�l]��hQ�� ��$a�!�B�RUAK������n��ITb�H�'�y���R��,����Cn��:�'[���Sḷt��%z�<a��"aK��^5�h�SJ�s�<iqaB&ֈ�u�;J`��� �d�<�u�T�^dQ�M�:-%�uӃGc�<�M1(E���%��ta	e�b�<a4κ���
�Y�O�b�<���ˈq�Z�����z�Jህ�c�<Qv��V�����T��IPӠ�G�<)"�yC�����^�0�H��N�<��ڃk��mxRg�d8DB�p�<a"�Ųi�Bt�1nԏ^ʂ�����c�<�%L�_���k��KA!�w�<� �F�F�mS��W:X��Bp�<G.ʮ6T��g¨fW�ґ-Fh�<Q&��?s9��j��Z"0�q�?T�x(2�:b�&��--?��c��?D�T���Z�.�r��]��H
�C+D�\Z��ĿMl��1'ѵ+|�)�#D�|IuĐ�h�^[W��d��'"D�D2���-*�"� #D}gb�;��4D�Ӧ��$oT��V�&�DlSa�.D��ib�6��I@�Œ�7�RI�ǈ*D�hG-[d�hQ�&�Q3-~���N#D�� N�b!��=T���Z�%Uu�F� �"O*p;À�4'ܐ쉆�L%b�,��"O�X��G]61��[�/y	��"O��#Vj�g�}�tn��J���
�'�"�;U�,�>Pk�R�"�'�V$r7l\�W:��p2��J����'����� �r���KR�I�=f���'�����8 �$%��g��	�'���H��$v�D�C'b��D1�'�HԒ�^&r���.�e��c
�'�������;rI���\u]�ɩ�'�r!Ru�\"@&�,	��Ա�f�<a��ۯ$�4�
u�ѽ9xz=�6�Bz�<	E �/װ]H�Ը�n�+���{�<��I̲nji�1B��[%ǖx�<a2	R�(3��C�J41ve[�@V@�<�у�Y��J�/	�Lc0�a�<�D�;��� ��'D}�UT+�D�<	� \�v�� �6�RQ�qi�t�<�T��Nnh�#���f�v P���p�<���11�}xG	�Zӎ@Q&�G�<	W�D�Y
�Rp*M���i�<QC$A&1JP,bB@�icb9�!c�z�<��kK "�H�C#�I	'VT"a�x�<�+���"���܍0-H�%��M�<�4��<=�Ƶ B�e�|P���Q�<q��#��dhV�>$����[P�<9�jU�ǀd ƩW�y�踰dHI�<	Я�2�ƀ���4{��@RL	M�<@�>-Ѭ�0	&q��T�pJGL�<	 �ҍ{:�}��̐#& ��RS�D�<	%��`E�y�'O�8\A�S-�w�<A'�[9Q��1gɟi��x�e��X�<�3�ݠC�$��W]�~*ĤBe�V�<a��j,�8����=+H��VLI�<�ƚ#Q�]ydO�>;o c0��F�<��*��MQ�����i���F��\�<)��8n�^q	�����ɐ�[�<y�d��]ú| s�5�	�d`FU�<Q��.N�QíP�n\`��[w�<Y�dh����[M��+T��p�<��̊�Iw��(2cԋv�a�#cT�<��bׂ;�J=IS��� 7�Ԣ)j!�?��X��#�1l����ч�%=;!���2�0��@��U�� {�&�>!�d�E��E8P��A�Rp��T/!�_N�489���7[wHLK��Z�!�$�7 �]�֫cZ"�˔��M�!�D��0(��ቜXv搻B瘸*k!���$R𘱦+�c_�����L!�Ć���R�`��J�>E�֤I4�!�$��p"<�f�� ,Dl�QrCυuq!���D�y�g*Ӱ2���VI1a!���	U���C�mE�O��Y�`C]%!�D@�$0��S�I�ܜ��^�F!��F���s&���p̂w,E/!�d��	S�P�uǕ�N�v`ʔE�6A!���;�@˲�� ���iQ��!��P�Yh«5k��9�e/Ǣ�!��/{���a̵�R�Kc��!��)9��@��-��r�J5��N	!�C�ASx���{��ኧ
�T!��<p62�Cdʣ4����QC�&cC!�����I�L%��j�a@>o*!�� ��4N�:`����U�<����"O�\{Ġ%���R�Ǒ�S��#�"O*-��N�-Sz*憊%w�� "O�5�"���Lvjy��h�4|d�i��"O&�����٬�y����0e�$�C"O�UpcY5Y�4ٚ��:u��9�"O�Q3�F�hL��S����=k�"OZ%�R ��w��g��i$t�F"OdM����=1Z��kA4Pz�4�"O�9KP�X�b.H=e�H$Td���"O�iء�߷�\� E�ӫoL�9��"O��J��ׄi��� $�6/�i�T"Om�����0��\hr�K�V�� b"ON8��,B�a��dh��\�Q"O~`B��#~\͘�G�=�ҡ� "O�\�FI@� �D�[�X@@�"OE�R@ �c�c�7����"O����i��W�Z	���Y�r��G"O>�7�E�/4N�2�=x�Z��s"O�U	A�X�6�z��� �}a9c"O�4��^�\����̬I4(�"O �z#Hү{�<m�b�L<Ұj7D���Ќ�j��$J4�T�pP��2D��ٔ��)
 yGяԜe�U�:D��
%��4��(���2�<��c�+D�3�J��-Ba�9��%Y��-D�ؙ'�L*'�H%斓9���N*D�T&L�7CQ�����V^�p��)D� �>�,x !�� U��:g.'D�Tc�+'[������H���1D�t��,�v�s�6S֙�Wd"D����
����&^$At�� wf!D��� ��!xh�2bN1U�l��f.5D��"Se�:/��I1���b�k��4D�bc�f�z\KqI�`VM
0D�8�u�c�, 	d�W�{� ��1�-��<�O��KS<��ň��K4oq`HX"O��JEh]0"	ș� �+>p�`0�"O:h�/�S~�١��� p�a�b"O@�3s��#j�F	���G*;��"OV��q��$�HQR�O�\6�9�"O��S%Ɣs�Z�a9�^���"O���7�E)	Ml��G��%J���"O�4�
+N�B89�Ä�sq6!�W"O�@afT>�>5Cc�Vfp2"O�	r������5$�薤%ar!��V����h��\xqq1n�e!�Q� .�g�7k��XІJ#U!��C�/����G�ep�EpV&��L!��X�Q�X��)bm|0Z�$/{��O>�=��P��G��*#����k۔Ө-�"O�bG=o�2d����ϴ�"O�A㤚�1Ѝ��gҖ�T"O4�hte�7e��6Aѳ�@�@�"O��B�tRbDˑ��>ZA4l��"O��8� �]�	R3ԜR"�$�q"O|����p&E�rN/�HbB"O0 ɔbX�_�W�%F�$4��"Oh( �9ռ�JS 4�9��"O�$��O�'X�Ī�N�!���	s"O�d�EY�H�����R�S�L�xS"O�| � �>x|}��k�?+�"�0�"O�8q��),�P$r ���9�"O���S*ؖ-���p�`�:ie�Mˆ"O� Z1�d��O.LD 2 Y/eB��"O�!�C�˯.(���@/m�hDAp"O�M2q����M�7��-�y��"OU��M��:�0`�s%�^���"O��f OF�)�j�[�
q"OZ��GL&B�F*�(�pa#�'��Ă�6�N���"N��zA��j�m�!��p�����ϡ+�P�u�ı�!�$2��P K�Sx���ÿ*�!�D؆-�*<�D�X�s�N��!��-�$B'ׄ>�*���/��q�!�$���I��(֧?��Y�aO_'Z.!�䑊U|�����%e����" C!��	xP��F�LGes�J1PG!��,Fe��S�
i������!�$<�А�DdRs��U�+@d�!�� ��m����O�EؠKJ�Q4!���0�Ubf��=	��3�Ō4!�d�'B���+���ę���X�W)!��� �xYS�dQ(������<(!�d�9b8�7�ɿi�\�:7ʂE:!� 	`x��)W
ޞA���,!򤘛L��	��+C5=����͝�	+!�
���$
rN^)L��QY���D
!�dS&&�X�c "KJ\(1�g��[
!��[�E@��?_�,�v(�,!��BiXRU��"������@�/ !�$�1����A@N{L܃wM��%�!��� N���4�Zxph�l�2!��?A	�l���r19�,�!򤖻J�X���g%��Ê¶
!�D}�.�H�Dͽ2��*6�^�b!��.�B;q���<� 窎�N!�d� �Nh2p��tĳvʔ�dd!�ҕ;�����@).�,P���ѕE�!�Dg2 �P�}��7�)C�!���9Y�1"Ħ�a)�;�Zt�!�D��_��Y���+|�����!�����y���]3Q�P+aE[�!��*}M^i"�gR�x`�Y�'�!�ϡF�Es �@	� ��Ϲx!�ě)8Z��g	�P�DUZ�:08�'��D��~b��J�����`q��G$�y��#��Mq!��]�:e`@hH2�yBbR�|*8��u+�&~��D+�bS��y��2,��|zG��)�La `���y�/Njj8�$��'�����iج�y�ꒈ+��x��'�&�f�yr��/A���i��T#6&��F�����!��|
�y�Ò�~��\8��M�lTr#�]��y�k�
Tnu3teH�����G��y�i�%;�h|�%#�BW,��y2Ǌq���+�
Ě z��c�K��y���)$`"��ΜM.>��E]��y���y|��QQ%�!=�R$�G����>�O��Z�mF�C�}{��6k{F���'I�X�����w8��쌝0��L��l$D���'�����"��5U:���P&$D�h�Ă�0+%���e�n���R�� D�h��Hñ`*L"�(LA���:!�#D���A��4�"I�Ӄ֕=��i�CH<D�$�*�"�������0i�1ʐ�8D�L�U��_@�)s���>V�u��5|O�c�������o�"sR��9�(1�3D�� �h*b�ڦv����U*,{�T��"Oti@��SJ�Y��J� UjL;�*Ol��5��Zhz�s���x�'pF�I���8t�eRc��1$%�q��'�F�CW�ϣN���	C�޿ �`�@���'H����M�u��` �i�	Pڡ����$ ;D�)^��mXä%��/�!򄍬n�-k��q'6l�#G�u�!�D��;R����G�k"p"I�l��I䟴��U�Iy�O�,�I��Yx���0eƳ>�����'��`[�(!I�g�P�0іx��'��Ex�Y(y.L	�@�߲��
��?A�yҀ��d�Pa�Y�	Ҕ�K��?�y"���k��U�b����y���yR��k`�����3j�d�sdJL��y"��	=��R���[��	��@J6��3�S�OG�0�`*X�U+�96,T�6[��P�'��d#���5u��IEE��+ڊ�)�'�t9��LT)�#��e4|�
�'e��c�dT�a_Z���aɚO^(`Q)O���䙼{T��Cg��6|�,�h���,
6!�_�|F�Qx���l��M؀�Ey!��*\�|q��¥���8k�	�4��H�)ʧ.���
2��hI��ɱ�^���t���M����A��|����	 �2X�ȓ{Y
�"�B�
u4,с�͇Z;&���)��asOG�JV`�д�	/�����B̓E��Y���� 0�h@���S�Lp��E x�Ð;y*(�3�lčm��Q����<��FZ�0l�+ 2G"��˴��U�<�b��3-�R��ת%9N<P�k�S�<�
2{�<�[�%V$<hǴ��ȓ�����_3c�8y W�[ �n���=��8����v}� �B�!.�>����������$��"uk�.T&P:���8�}�ȓ ��53���=�*�3třk�Tń�	�<�!U��dx(��M;�z��q �q�<�� ��DAX`�OL]La�l�k�<Po��n��`ؘB��i�VAE~�<�JW�,)�i���tLt�P�T�<���p����.".��BIP����F��9j$(\<M��A��p]���	u�'i8�p�fP{2z$nڟyp�Ń
�'�根%#�7A"�t�ւk��X0
�'���qD���)�"@a��Zx�Rd�	�'�����F�m�z� d̕?kS�@r	�'{�lqR&�aD��(�-�8�hp�	���y�N�"*� aC�<�>dR�h���xBa)I.�)�Tŝ�{Nl���燰Y��O8r��۵ ��kT�wk6��P"O*lb�ɃG�Y[Bb��,���x""O�'E�kTH�pNޑy����"On���m;rlP��U�V�%�8�+%"O�]ʁO�u��]�D���H��"O�i���Ψ좥�C �.���(�"O���B��`��3�ݑ\c��Б"O�%z�X��6���ݚ2mR$xD�'�1O��rOݿm_��aoQ�D3$ @�"O�Rvm����yr�rOp=y�"O>��A`4_�x�0�K�*(QR�
#"Ox���ظ]�^1aqj��|5�m��"O����6 ,1ŉ͙J�>���"O�����]�J��T�$�^��"OF|S ǎN�h��g�#'�P$0P"O� (��ń�,�PM	�^�-�����"Oh�R��� P�����!f�:�jf"O�X�c*ƿ�Ƥ��)�B�	�"O�9 %��,, �R �Ic��]��"O����< b�����+[��q��A>��ۦI)0A��"!N�h����"D��@��S,%�0]��)��y4\`2� #D�P��h���AP0o�hӐݚF� D�0��;N؄[�.��%;�� D��rq'ڗ�MQ&	N*C|��l=D��� ,y���
.eɜ���@;D������/����ĝ&nyr��O��O �=��`A��K�'z��J�O�t�����"O�#S�N<�2���c��d�R"OVX 2�
FՊa����<�����"O�m f�w[<���=F�a��"O�x�OG
 ���;$��'VX0�"O]�1	���z�!_�rRHI�0"On�3��14L;vR}+HA"O��%��%V��c���	}@0�T�'���������`V�H�� 9��9D�����e���Q��U�i�v��F<D�0r�� H|̜a�شwb4�#W7D����&�T$�e!$$�K��5D�ࣗm�B,�b �ة:�|�`/D�$����hI˕CY�3��� t�-D��� �/5�p��nˉ���6D�<��,��A����2|~����*D�ıF�=�(0Wㅘ|E��@ӈ)D��yc��?�=K��6k�rh��*O���"A3pN�� �/1���"O��b��c}�����-8k M3�"O�T(S�^�,r�Z4	R��f�#�"O�|T�Gg��r�H�$�i`"Ov���
�㓨���Ib"O
8��I�jM�萀7	
�	w"OL�Y���q|������0�"O*4um�^'��Q�?P��1�"O0lC'���V>,�m��$�dy9T"O�y�N�%8b�ԙDL)٪}x�"Oı��J�kW����?�4��"Of���3R����壕�w�x���"O�X�t�]�n���,�Д�"O���Ԧ�#d�`MyRcU�F�@���"O 8Jլ]����u�G=_�p�@c"O���ʙ%U ��O��M�e�1D��ZC
�-\�te��(8��ׅ%D�d�b�\����� ��YQ4��t�!D�X`�Uw��[Rk�1M\@�&�=�O~�	��xh`�D�x��M*1 �^��C�I# l���@����y�Aߩd��C�/�\ur�dY�nj�5X�I��C�	�N&|���N�2j�x���-ȱ4�tB�ɑX�I��� �	cr���"�XB�	-4���C�Z+V�J�Xǋ��#2,B�?F�0�y��V�*ٰ˙\�B�I%f�tz��Z2��HjP!G2��C䉗;+�h��&��ox��S��	|C�	�j��]��X�a��Z��R�w<C�I�������%gF8�2#/a�B��&����`���S�N�Q~�B�	4F`z�����_-"0���
!h���:�IX��~R��v;�혧B��`P��P��y�jڰ;u��2�Kdx�0�l�y
� ���B��5Q�J q�1v;Ŋ�"O̙�2%Y7z��� FR�6�V�*�"O�x1�gE���poM�
��L��"O@	��s�Yx�Hޜe�0�"O�t�RX�Q�	3��=*� j��'rў"~�����K�xcRmeGZ��Q:�y�L&@�t�S��LC�lJ&i��y��v����I%���c���y�!]��0���B_�ņ�Y�Aи�y�$�QG(� ��}i"�V��y�)_p��y�3A�{�.)��M�y���5c�t[@�zJ2Tpch��y�z4j��0C�t�>}R�,׏�y�	HT;�e#��=��E���y"B��Y�D�PcޅO��,��-��y�FF�s&���]0�ș֪Ȥ�y�)FR%!�cǪ�ceA^	�y��87���e	4b��!J��y�aY�<��Q
1KJ7$
2ՙ��̚�y�"A7.ZX$R�k\�3U�,�s����0����'��HB��<WA��H�HI.�����',R4Id��;1�Rh�7	hd���'��(�Ԍ�/���*��-{"\��'�<mâь����i�|�.xK�'�ހ�p$Ջw��ㆎ�
��pz�'�`�����1��%(s�΢v�䀚	�'m�I�RSN| � �7�x$S��$2�k`�@�C�_���q4)�3W���AD,�H��*6ZiS���V��ȓW����$�Z���]k���{U�5��kL���ܿp���O+w�!D{"�O�T<q���{>j	���@�'v!���M�;y,)��y��T{�' ��B��!��c�B�(le�x�.O�����X��@Gʈ-8�,B�L�!�ęH¬� D$�&�,�'N�%`!�$Q���Ы��n@�[�?2~!�d^I�(����WQ��ɳ��4sf!�D\�s �Չ�NR�|�X+$�+Q!�ښ'Vu@�G��D��Iy����^J�O���$͔Z�ܠ$o�}�V A����>CO�)��<BPjh�b�;"����"Od�"�:py�YYW�]($��"O���l�5e�y���̄e����&"O2�mU�/�`��♲&���yP"Oz%I�� �_�܄�����f��Ȓ"O�t�$�D�, D�(0-�'5������j�@&و �4_^��e3D�j���<@^�@: ��11!�.D��+�GG�p��h�ĕ=b���di1D����ãT��8c��Ba��ۆC0D���.�8����fH�pd~�t�:�����O.��,IɃ�A�w\�e��h�0��q.D��8�g^�I��1A�������-��Fx�$+RE#(�l����[@�h�'fFԟ�&�LE{J?�b�Hmp�L�q&�nf���5D���E�GJ�DA$#9�#��3D����Y�{�Z�Y ��[�f �D1D���e�9{8��hс��"
M�7��O��=�O�1O���ꂅ0���c/�c~���0�'�!�$�<}��(���,M�ш��btBOT0Ӆ��B��Q&9Ip����'�!�$��wwb�b7M�Da�e9�	�'�'Ia|��P�]^n�"&�kXʴR�jʪ�y
� �Q
��� ��@��#%���zD"Oн�efӗA:�D����=�dȃ���2ړ��č�Wd�sb��1�0�[d�/�B䉶z�$�!�F�k,麃�2B�I�[G>PRR(��P� ��eb]�0S.B��<���� {�]�ʙ8b�B��+Ly�(�ȄD�BK�he�C���(i�CKO�8��$ʎ<XB�(`����F��&K�H8U�	�ZB䉼�B07lLw �IyPN�mTB��7��J��]�d��{a�D3�
C�I�~& 	�d�K%b=��� [�Ң?����ɟ/[�u��<`8Cq⇌%�!��M�����̈́�7fr`�W���u�!��.X,�:�Y� ��1��`Q�lk!�d'�x� b�P�z�ָ �aǌpN�R5O
��#�׋J@IyGH�&$sj�"O����(�s�D��M�xo(:AS��D{��	���rbd�?&J�����4�ўP�ᓾlhP�����tct�6�%	grC�	�m�4̑!��:�Ht(��Q��nC�ɩ>�l���A-j���a1o���DC�	[�IK D�V��P��X�pB䉡8H�iB�ϫQ���`���#Q�$B�I�xy"ܚ�n:I��P�gXʓ�?q��D6�I6 ]
�	�É�	�0��b�'^�C�	=�
=�0��!6:�;N�C�C�6K���PE��Ԅ(d!S�"O�m���t���1X�y:��G"O(�ą3p�ڔ�%�̀:�!'"Om!q�h�$Ÿs�S�hj���X��D���7�]"F��Fh@s��O�C�ɣ\H���݁h�N���ĉI��B䉖Tx���m�$ dZ�I�(�p�O@��ē�N��0��,>;U��[2!��A�unlb���X@�J�I�,#!��Gl*��A��Z�Ƚs�.D�l!�D�XسFg������[�1W�O��􄄁9D���̕
k�D����Ψ+-!�d�5_�U���47�-FB�G"O��:�L\�27�5���O�)_�y�|R�'az �;/� �CN<+T(H��I��yB�d�Z�&R��0��$I0,�ȓ2�ꔈ���o�n��F�^h��ȓ(�j��F�H�e���1�h� pR>��ȓ25~�@픬`���V��2]8BI��P�a��,
�L�Ӎ�_`��ȓ�r�K��TZG��Ge&��'~a~b�>]2����_�@������yBOW�$�x�@V�9�\�@�A��yڧ�T~�|a��@;F�r���<D� ����	������@�r�6�Y2�-D�lp��Nn;�0�b�߃^�Z�l'D� �B�փS�\h�D�:2���(�%D�d9`h��	�͈U)�4*Xy$D�,�1'�u�� ���V��A���$D��z4 Æ}(� j$+�'����l D���
-w�X���	Є9Qx\	��2D�!p�O�W(p]�!�a::�[�g�<i�D�R���H�=݀��@��<\`���ȓ5��ؗ�Yu�]�p��y�����J̓l����)F�ĹX�G@>*E�$��\��Y��LٿahƐ��&ɷ�(��ȓa��I�D���ab�շ)4���S�? �qz#,]�����MY?�&��"O ���6����?v�|{e�|r�'
Nl� �;+��BӇ �-Pd q
�'�$(X7̑�1@z�K��Ha
�'�N��dJ/$����wɦ-k�"O��Q%���m�M0��B O�Y%"O0����ȵ
�"��n�Y�G�`�<9t�΄�j\����Ps�P��f�`h<��"��i9�DY��E�ǆŘ�y�\�m�d�IfiM�yd���Q�Ҽ�y��\�X� pš��"8IH�
>��?y�'��H@���+��%y\���'�P��w��\_���q&�
Vui�'>.�b��H�H�{��W:T�\D��'�yB��HԨ��Z֜9H�'T����*_9f~�0�gS����x�@�o�ƌpw�'%¢�zV&L��y�E�Q�����+ �"�����y��D.h��9;��}��8#D3�yR,Ɛ@�h�Ǫΰ7Z�U!�)�y�ϏDH�S'�V(S��DQ��y�dУ�6m��.���\��	�
�y���!�L�3�Y���)����O�"~ʑ պw�ЕA�?j݂U�5�~��hO�L����)5`Dx�(�<\�؇ȓMF��]	t���g虾2D��ȓ1}`��#e�.@6��η!L����}0Q7dіD���@�ʹY����ȓG�dbeִf<��B%PVu�ȓ<�D�!f/��`e"�"V ό	��q��]���)E�}9z���N�l;���ȓ��S�	E+]���26D�[�݄ȓ$�dM0I6��
��ߨB_P�ȓ�Ɯ�0[63J�r���=✔�ȓ(Hlx��ƴJ��b��C3�E�ȓ{���P��I�b�E\~�@}�ȓK���)]�r D���Ǜ�H�'.a~���a5�X�����8� e��y"/�f��2���Ж��d�T��y��U!x|0��Ҿc�A1C	W?�y��D�_�*,�PG�VT�S�"�y�A]���PVbހX@��Sh�9�y��Cc��A��ƈK�@1c�H9��>��O.�ʶǊ���ш�8'j��"O�l�b_'�]� �R/3h����"O�q�E�A�ɸ�-�O0��@ "O�-�'GG�~�=e�Ƀd!�t�B"O�}e� � �
�̃�s0�#"O:Y�%I*"�����*�s��s"O@��d_�dBFM����+px�$�!"O�僧�]rW��M��pI\�z�"Ony$�!��-Q2�z���!�yr�	�:|�uJ�T�� U�С̭�yR'�c;B�����?`���)1�y� �p���AV�ڍ�\)�'%��yB�J@/p�jrO2N�q�E�7�yB'�'G*��mu�f�,Κ��>�O��%j�	������D�}��Lr�"Ov��`ז+�T�s���n�Jt��"OZ�1@$X b}���M�Q6�y��"Oniad�2�rUa$\(#���6"O��x�J��o"�!C�[�eU�}"Oԥb�.�:P0$вۦwI��Q�"O�-b�FZ(�HXV-S�=�\zF"O� �p:�`<!�0��g�I<����"O���uL�	 u��C��K(��"O0P�)��um�(Z�i\�ȳ"OZ�#�lG��L��d�_	T��L�b"O��#���BDT�D�?J�tɣg"O<�&AI1xNh�j���B'T�Xw"O��`�aPEz�����"g>�)� "Oz�"��ǒj��� �T�f�@4"O�D���e���C  x�Ĉ �"O:X#��+�\��s�&i�6tpB"O��� �?A�@ {�H\51�V)��"OJ���&QsI�gσZ��y2"O��'I�&,�ȉ�׆�IJ�Q�"O����)U� t�9}3� �r"O�E�q��:3�p,9���$.�"O��{�eøl�n����4]��X�"O���X�����Դ\�� bV"ON��D%���ٰ�# e�[�"O��1�\>N���'��-�X
�"O�\#,�N*�(B�K�~��z�"O2Q��O�>6��M�aS�J����F"O�$�U�]>[��d�ĝ�u�"OV9(�c�2$v=0��\Q�\ȳ0"O��!`�ڛ'�	
4P�.;�e@�"O�q2ccL7s�V���'�:+$V"O��c��h�  rm>7���"O��Yq)˥����թF�{���;�"O �cc�5$=Zxa��\�sF���!"O���A
�;� 1��Ď79~�F"O\$3�ɪd%"��s�P�(�"ON!�P)�%Z��V��B�Ш#7"O�ɩ�C�G�!������ �"O�Xbpm
�+�xab��#xf$AD"O49����&2 8�K����村�"OH� �mނ<_B��ȜQ̙��"O^	��*�����E��W�*�"OhmBt.F 3��ЂZ4d��#�"O2R��]�/��+�����N��"O���!δ4�b�RãX�zT9�"O�ͪ�락(-$��I�T}2��t"O0�3����3a�ɺ��Q]�p��"O�}��L!g�T�b�O�)�Q "Of�õ��b�~��5�W��"O:eȖ,�.J��7N!H*t�"O��AQ�n[t��N0�2����$��l*�z��#��uh]�&�^�{A��V�<)��Y�F"L�q4R�M�Zqc@XS�<�`�'Ğ�;3��M��k4�IN�<���hi��Ei��3~R�ⷍ�I�<�`�D*a޲���&�e��	٦�k�<A���hh� Te�5���v��f�<9�&��K��	�"Ӿ}�b$��K��0=���7k���CK9	�"���N�H�<a�<�pyCmɫv����f�A�<9���05�<s�)ԿF� Г��I�<9A�F�lƂ�C�:o]xx3���F�<��ē/��9�N�ҁ�6��D�<�v�K�g���q�^1Ew���o}�<	r��&>���GV�	��
��_�<���	�n��T ���W��m-Y�<���-4VjE�rh��v���Q�CW�<YăQ��E��C�N+@d9�O�Q�<��\B�2QSC���&I)�%QM�<�t$��t�tU���� �Xi�6��E�<� yÇ�2'c�=�7�<�ܵX�"Oz�Ԧ�Db�#񧄎/dՙ@"O�lxj�F F�I�~ld �"O��!2�R+�R�s�M�"_��Y�"O�,�F�,�PhA��#5J�I(�"O|-�Q�.I�]
�
/�؄��"O��ӷ�<]1�,�4%G�vp>ͣ"O$�(r!G�OϚa���+4U��Kp"O���*$Q[��_�wb,u�R"O����9�X���nǯNK��)E"OLPP���GQ:�ZŇ�J@B}�"O�H�+D�pg0Ԩ��˞Uf�H "OV�+���z��6f��%^�Q��"OԄ��d��D��Ъm�8	b"O�Y���M7��h�SRFq�"O��[��p���Z�	���p�"O��H��,��x`�޴6Ī �"O��	WϜ��X�c�`Q

$@ݡ2"O:tIG[�X����"-:y0"��2"O�a�$d&�H�a�,#��"O���cERc(�)�2��`�t1��"O��R�|授�M��^����"Ob7H��@���	
 ^6��"O�AA��j�)&�P0^L@ (�"O�͘�"�1't�L,3O>�m�"O�%��
D�V�Bu���ڰe=B(��"O�(k�#ʏ3�h��'�"6#.1+�"O�(�g�0	纀{�'J�F���J�"O���aƀK0Hu�F&�6T�>3�"O��S	����C�%f��5d"O��BÌM��0Q�&p��"O -�U(��wm�|�s
֊id��@"O�x�-��a��d�T��+�)c`"O����l�I�����A���@ �"O@%�֦�C0M 	��Q�.��"ONձ1��LXL�q(�`�֑s"O��c��.Q$�Hbj�/ ��ʲ"O�R����'0�X� ��^y�s�"Oh��*дA��0vϜ o�fU�"O�h��.҄�>��B��e���"O�3�MՕ}�lM '��2v��QW"O�d*�'�r1Ѥj��*fu��"O��z��_'K�H���݀�R�`C"Ov�!riې$�V0�T~
=�"O�9"E,����e3W�U:�"O�X���ѐ\���m	�O�,�g"O� � �8�f��&n'2��}b"O�Ъ�C���a��у_Es�"O�aX���GR,Y�V,؆bpv��"O�`��ۛm8*�p�)ָE�0���"O��k�U�uH�a�7h���c"O��!#��� @2 	<��"O�X`e��Y��a���:��u!t"Od�
�+�%;����$��jВA�A"O
�l�6+�̰E�߶P�"Ot���#i�yP�> y�"O�z�(ɮo@:�0�l�h��h�"Oz����L�g�6�²��CJ��Xg"O���$�Fg��
� ݌4��C"OJ����W��4�1.̖j���g"O��sʗ^r�6)����tH�D�ȓ2��rv�C�.Ve'�6X��T���
�Q

:z��aaA�W��!�ȓ>��
��:�4����y�i��S�? �Q(�CƄ^G�@��D�S~(�(�"O�@h4I	GDL}1�c�Fq�)��"O��K�,L���=��\�eeXEj�"O�� �AXT
X�@W�^�jy2e"OX	�#K�LB��ҨK%ote�"O ��ݯNMt�󆚿+z�s"O��X�&Ѡ`�~A����>g��(%"O�u��"��VLx+5iف$yC�"O�D�(�v�9���ފEp��"O���('!~�S2jW><6��"O ��b�:XDd�!�I̕�4D��"O�Xr��Cz9��.˽U��ŲC"O,��P� vJ��g��w���yS"O\C�*H02x���(hԙ��"O(�ks��2eP�B�hߚRN�a "Ox�c��Э7|�����*pʴ"O$݉�l������@8���"O>�� �5��ɚ&�'F(]�"Ol�-nX�����@FI��"Or��Fw$Hh5���s)�h�"O(��ኼ;��M*��X$���"O���_���ᡥT
�❈g"O��RF�de�f�\r�J""Op��o�11���;��¹ d��0"O@�0Ϝb��T�������"O�E��	V�9t�Q�G��p|z`"O��`WH[�v���cHo�j���"O:�k��L@�Lp���H��"O�u�3dG�������>_��AG"O�A��F�@&�/��+T\ɳ�"O"}Ѝ�;b�Jy�O[8u> y��"Of	jV/�Q�ޜ�7�FV:�
 "O<�(�iR-AΩi��8:Y��"O�d� �S&
���ǒÀ���"O~�on�<�Bs.Vr�� ֆ,D�����wj|9%�{� ��7D�H����t��Ё3��&��27/*D�([�c J��r�'S���(#b(D�h����p!�p !��J�f�&D�T����5>X�U�2� w�/D�0c�I���#��2Y �!QL-D�(x'�	�T�6U� �T:��s��0D�,h��4S+�$yw��;� 
!D�H�1`�
O�����La��Rp`!D��vT�~��]� �L�$����#D�����|n��!j
? ,��a"�5D�,��l�4*�vh�˕�^T��1D���1k�HT�s"Td{کs��/D�h:���{���cH.e�0�:D��Q�J7^ș"1��}(�� 7D��3�	�Cl��9'/�K���F� D�@��*&v�q������A�*>D��S�ж?M�@!�đŜQ�т!D������ I"t�J7(D�y��C!#D�4z�拶U���h0�T �t� 4� D�|�BF�B-H�SR�R�b�����(D�b��k�� ǎҲÆ I�1D���u�	m0pA�T��%R^d�w*<D�#R@թBo�y��DQ�F1J�+��&D��9�(G���rR�Ɋ|&V(��8D���OӼ{16D9�#�
L �1H7D��HB*C`XzmH�JD�0�A�:D���S㍷#J)"vg���Li+��6D��cǌ�� ���ѵa�b�R��3D�� ��W�Җ-y�tr��/�f�0a"O�Ġ�h�ft-@AAV[�ʭ�S"OPu�#K�d�����OĒj[�"O� ��DZ�}
 ;>�|"O��c'*z���Rt.����f"O&|��o��1	�<K"-�}f���"O�(��M�< ��0+O��`�P(""O���sC��0�IE.�e��z�"O�pذnL�q_-���UR�p�"O��!�'�v�l�"Ƙ�`%�I�"O�%��2<ʼ�p��(v.l�a"O<PmӀ_n�S$V�.=�A"OH�x��יmv���*I�b�b�"O��3��ж@�c�m�� 6"O��*ĥ��P i�U����� "O�� �$e�0����[Vu �X�"O�P��:E��Jڠ���q�"O���'&&N6��U���;�&�0"O�Ř�gۇ{m�<�A��!mFV]{�"O,%��Euz`�ұ �,d1����"OF�Fŝ�aҊYY�@��x*�"O��(X�jW�<
A-��,�q�<�&�5�D[��:���+��F�<�D� rz"��S� ;/������x�g�5gf0�*%�Q�#ϔ��$e�͸aB��
��ub���A�T5��p�������'O�,�g9v����ȓHኴ�� L'Rdt1*B�4u �݅�"tHct��4`� @����4L���N:"Ӗ.�/,NtX#A�|����ȓ|� �`��M(}���e��%����ȓ/X�e�r�Ǘ3I>���ū����w�μ�Í�"�2�`�l�,P���ȓoH�S"�V����r&���J��К��cm o��q�H�zR�1�ȓ?�6҅͐�D��$	��CO�2�ȓb:L	!`���a�0�,U�;�$��ȓT �,�v�H0W�~�Є�Ċ?����&����{�X<x2��s�-��mE��c�!
t`��fRr��c �%�`8�,�X�@� �jt��s�XM tEBf�a@����eu��ȓ
h,T��ǌY, D�ʵa6D$�ȓJ�tya�R�N�y�@�43�x���j�@�!/C`F�k���?�����K��m(�FШ/z8���Q-F�y�ȓ�2uWFLb`%+�V-l0�L�ȓ��"j�o�h��� )�$��=0J�:vk�p�D�J�L&N�$\��)�����I�#�Q��#��?�,�ȓ{z�����ӊ@_���R&W�-��Մ����SC��N��c%�O�̙�ȓj�RH3��IN��!B,�<q�ȓ%^*Is��+69�9!������[�N��V��-C!��Hdi��$V؇ȓ!8��TÀ�lD��H��ƥ+�����7��u�������<���"6D��� �B�Y���reZ�m��tKCN1D��0���J��a�Y !:�!SM;D��8��Š`���P�ء_î8!#<D����Qn2IP�*V*qƌ�R�6D�l�P��e�n��6��U�����c(D�ԡd�,v�p���xX�v�3D���2�
>���Z�/�
,�8�0D�<D�� $��!fJ m�-"� �z2}#�"O�Mq5%�p�b��M�2Oa�PH"OPmZ�M�{?�Xs�͗�vH�8�t"O�5���1��pDmͭsF��"OR����y˄�4�ʙ[���Re"O�AB"`)����J�^��1�E"Op<��"U6T��P��4�H���"OPj�1KM�|�#�O�4���"Ot=�B^���L��/�y@�"O� �b�D�}�4fљ%����"OtA�@ꊺLx"��!f�D���"O���J�J�!�o~cƼ�u"O*ܰ�k��8��H�;Zp��a�"O$Hu�  U5D������T�1�"O�1��.K:,Ȳ]�����"O�d������
�QI�j9�"O�MzQ(�	"ԩ�\�Dz��0"O���!�%[�x=0Q��7FuH�"O@#�>=�D0Ps�U,W�e
F"Or|XiJ0K�$����M8?����"O�,�S����H�P��V,8!�Ǖg�J��4�s��Mpt+�?.!�$�1���е���f���jF�!�DЖy�6Q�O��Z��t"�)[�!�Vl�f��V/�2f��"�l�!��Z�i$���s#A�/K�|BAE�)'�!�M$=��	�	::��;e�(5��HE�D��?��t�W �p�a���E'�y��J7O<.�S��T�Rta�D��y2%2:n�8WG��F�n�x����'>ў�O3�{S�ʹ�8m
�o��,8��p�'~8ģ�.%#v��K�!����'�0i#F�� ^��������'�0��By�~5 5�����0Ӎ��)�t��J�(q�bH��c���yU�g`pEMB�E9�8�h���yb�ϤM�"p*�62�X�X�ޥ��O�
 Ǌ�:������"@�`#'�D�<�1�R$O]�A#D�_�h�C��@�<�w��}�DL��F�-x�!'I�u�<9a⬻��8kА��
��p>aa��x)��647>hHb�Y�=U6���	8LO��'���Q9 �X�.�Cʠ�cI�N�ў��e�'�>!�7�/����U�����T�0D�@6E���@1�#LR ��0@h0�	E��$�3���`l� qlܠ�G��qh!򤖻
�9��R�h���i<|��'����!\O����(-,���_3�u��"ObT�#�M�VB~d��Ή�ڨq�"O(���/BȂ�j¨�ɱ�'���[g�P>�p���E'~�Z�%����U!c�J� +h�
Qd�r6�I�<Q��_�{�(Uҷa��M���Q�(D{��鄪]�|���?k�T&fQ�V!��9K�x��%R�%�DY�t�҂!��'�a|b�ɭ<	D4i��D�M���@��y�N \��VhL�[Un��۰�y*҅Y�����P=X��h �T��y�D��f��� �ɾ��ˊ�ָ'ba{��1	6t(�-o�(:2a���?9���>O6��fcX�Le��q���L���ȓz��k �����	��/v��-�'O^����;4Մ���Ϗ� ����\;*��~�[�Ęb�S�Քy���/P�T���<D�� ����--I���ڤY: �#B��B�O6$�y�@-l���
�}�V-q	�')�k�FA�H0��V�H)n/�I�	�']1��/H �=��̫5�V��'�xacQh�KI�\T��=KD��yB�)��DV^���Y�A�p�DMZ��<B��$�H���V(��x�7��XG>B䉜�D��Iٜ2����ۿ\R
���<��/�R� �	�JX���u�<Q�%}	���Q�蕓go�G�<�g
�����yDdӔ	>6�p���i�<	Pi�#�"!ps�K�D���b1Uk��q8�Pi炘')'��S!oƘ��U���>A�4�~�ޤ��a�B¢(�f�#0����yb�֞T������h�Fj���hO���I�K����eމJA1E-A�!�$<����'C�;�Tzu�̸n���@��(��X+	�Y�J�!p醷:T	��"O�Q�kA*%�Ii��ӠcXI�>Q��"�S�'�!�6.��o	%��"(&�1�ȓOp�l�&*63���eg��{j,�=�0�0LO||�!ɓ}9�!`B+�2:G9��'��	9jl��§�Y0H��q�F�E�l�	|���s�H��m��KC�O�X�����n"<O�"<1u/
s+���f�%@�!����<᳂;�O����&l�4�"�� K�fMȗ�|"퉰��"�4�H��Q�.��qX�Y&-��U��Kp�鵀YH
�y�N��&�X�ȓq��dS��l�����'�ў"|�rJX�
�,�㶃N9WOj��R�<A�F�"����-�6@kJm*% |�D$�<q#+�!޺�{w�^���<D�(@���y
�q��D��M����`����&�X�<	��,�3�0��0�	P���Հ�y"IXB��<�v`�9Ř�б�P��ybގl۬���`T�0D��ِE��ېx&[�k���D�b3�8�A��(��B�ɍQ�������Ԣ�#+o�DB�	�uR�a�vkGA��i�.��D��C��?+
�-;�o�`S��Ṙ�JG��'�Q�P�<yU	����ɪFdՅ"Ɋ�(�NYu�<���~��`e�s�X��V�Eu�<qU�%�t�y���]!���@u�<	5��"��� /Q�r��t�<�e'��G���� ����RG�<�o[ <5��FޜC �y�I�B�<i�N�w;,M��.^�_�|٦,�g�<��ҽ[�~�����){�(����J�<��aJ� *8zS��y*̠��H�<�K6q��	ZW�*@�r*�lA�<) P36��A&6|��zy��'ܐ9r�V�6Y�cn%+ĩ	�'st�Q�O)�K�$hPi#p"R�<Q�E�!hz��W�Z;�%���hB�]�� @�@�vL�af�>��C�ɚ5}�A�CװNP�!��P� U��'4��JN�,�r���dU>H��
�'�
�ؠ�S
:lz'ě�8)>(b�'�VYru%�,&yBW�3�$��'۲�9�dvނ��'إ'mb�I
�'Ö�R�� ���E���4j�2��I�̊��)�S�7�~����U:P�
�c�%�3r\B�I�l׌�p%�Vv�)���?u6��'��$2����yuB[�����V�	4�)��'��I1�� ������ri.�#׍^���R�<o�b�'�Q>5*W`L#��H�b���ۤ./��Y�ɺ���>�K�<��U��#@x�[I�'�y�F�)�<@M]�{��ڃdA����j�'ט ��r�a>�S`L*k�|`S�%�~��4�ȓY�&���C��{6�͛s+�����y���9E�DBx�'���b="��h�4���~��h��If?1��ze�\�s*�0?�̃Ǝ9�Jh#�{��N��<�p_���k�m_�V���NYP�'�ў�B
����8U�����Ҿ&�<S	�'1DXd�;�T�95��
H<�0�����XD��[�q�P5X'I��D5��x%f՟�yR�@/=^T!P'	2CԁC��H��d"�S�O��Th@dX^kc�U�R0���
�'��|��J��'��0�IK�D	��'8�PvÃ�\�l�P�1P�*@��'�(��� �^��Ń����P�R�'S�1���z+(=P���#�ny���>�H8�D��TtA`��Y2:\���"O�1���
9H�����P�3��h+��'�ў"~��h�  �#N,�y����y"B�jo4���'��U�7�yrN
�$���ꣀ�<g���׊���y��Y�X�h����W$@�U�L��y�@=��)�⁯M�P�x�lɃ�yr��%J�+�+C� ��!�P
�y� Ś-�����? y�F�?�yr�Ҩ?�>h��CI�14�!�yBLZ�n��0����F]h�h�yr�Z0C� ��M�?/�n��.��y�אd �hW�	8,lv}�b�K��y�m�/���b��2��W�+�y�P"/�������b��(����y���C��(E�Q�l�.��受�y҆Q8Snrk2�!:���9����y�Ҳ��(S��˛,�\����,�yr��*s��Y[�, R�^<�$N��yR�/:��j%JO�:����m��y�
K�w�b����,��h5A��y�[<J6���@ ;,snI�q�(�y�,G9&����C�(_t��>�⤇���" �ЍT)H$i��Y�pم�`(�e�Tk���ȁIO�2��<�ȓu�b��w��4r4�R���v����g�qP6�"`:��@���
;�h�ȓ"�*E+Ո�%g�FABQl�7Q�vy��zQ�u�āԙ5M�ui��B�et��g��*�D�n�F�ag.)�.�ȓm܈RțQ�>����Ndq�܆ȓ�҄�!�̩Mæ]r7#Ă*��؆ȓ �<�y�.�0zs;Sت��&��Բ��T��Q����~�T�ȓ8;�H�c���N��	- �X�ȓt�`#���#���ˋ�C��ȓ0��OJ�*+�ͺ{���)�"O.�!�A�9���C����@X��e��[��'�Ȕ��X�
�Q+<m����'f��!���� .)�mKP�d�<A��E�N�kv`˰D��|S�L�`�<9��ǉ.Hp�q�3m���d�_�<I�`��xM ��m�1>�������V�<Qr��~.F-)�I� JT\	���u�<!򨇇8 �P`VMW�"�Ƭ�&��v�<)�"�6,>œ�H
�6��E�n�<� �m�Ꜽ"����[�y"Op2��V��c[�7�ZT��"O���pB�F"��3b]9�"O YȄ�F�e�2���_,���P"O�@6٢^?`�n�0U��-�"OnQ0����-E�*Ha�A"O��f]NC�PC�j�Q�w"O|D(��<�f�0�»D�"�y�"OHa��K�%%��ԀXn���""O�i�/38$Q�e�آ��"OI�1��2c��2��(�P]��"OL��BO���$Y@��R34$P"O�Piĩ��H;0�KY�����N��y�m��<R�׈	 5��2�yR�.:�9 �f@~֬�؆JK��y�$bq�]�EA���3g�L��y��k���ؕo�
E���v_��y�mW�
|�)���#"�xs��%�yB
��{e�B��<��D����y�/Ƨ]3r��QȄ�B:���k��yr,���z����5�����	l?D��K�+T���'��l����9D����Oĵ�����䎐;�v�"ԅ7D�p� �ۿHA~�I�>X�bQ(��+D��k �U�3v0��T�?�D�0� )D��b���E\���� ��%w
�Sh(D�����"/�b�"!�36�VuHу<D���d��<����a�J�.���&=D��9E������0m����M8D��k����V�Y�]�ܩ�Q�8D�ls7�ܓx��;�)�*	���Z"(D�xr��ƅno0d�"*�4F�@!*D�4��(n��
0g�:�L��m?D���5��T��P!��aj:X[!�Ō88<�TJ��@p~pa��U�x!��R�T�󆁡moDP�F_�r�!�O'HW�����U�`��1S��EE�!�^?A'
x�$�а^����c�/:}!�D� �ʬ�r��:9봉� ���h!����ع*��_׾=�3BK�w8!�ߌp�D%�!m��7�8r'ؐ!��d�4�����-6D�	׍S��	$)Hd�1��Q��H�Ӄ��<2���S&�ZB��<`�J�!R〨 4��Ga��7�J�'@l#a.�'hnay�Y�[߮p# #Nf��L4�	��0?��$�'ʤ�Z���<8�󤉁-=d\`f
�'��B�Ib�
�@� $�,m��d���R#>�L_��40��3�ӡ4��Sr/��L�>%j����N�C�	�+;T4r��Z�g8�0A&Z-(>�ɣE|�5��ƒ�f�S�O�\��0�a��Mpd͉�V89��'�����.�8��ǇAy
�@�O
�I@	N�� �	�^\(;�	I(6wH�r���)��	�z���� X&���  ��PsKM��Py:
O�d�5A �A����EV�Z�`���I�n�6 p��~�q��4#2)a���ί$v��2H��y�ϓ�
�%��[օ)uV+�yr@�nF�\��!X��S!�ީ��Y._{\'-��1�C�	��I��G�%�>y��Զ,���'J�mn��Qٰ��$����\""���+� $4da��̮ �	�+>w���4�0+�p���Qh<y�ܔ��Ԙ���<R̨c��U�<)R�@��EyS"S"98����h�<	7C�'U�P��&aNP0���_�<���Ȼd�T�
��Z����M8��id��*a1O� �u�7I�[�x�@�� �$TF�+�"Oh�3 \P�����fJ8u釚��ӡQȐt&�"|�aǫg�T��&/�5L�h2cGg�<�����S|�@L�)�`*�"�ҁWU�@U����'/>��g�'�K��@Kivt���)<+��I;^���p� �F�*�_������OV"L��� �.��G���
	��C�ĸ�Nޑ1����wW]�a�?��K�O�^�Yg��%oUc�<���.A��%P�RJt�t0�
�0q�!�$�* �R��m�&o�4�)ROB�*�ʴB�j�zݼu�֫��'�.���� ���I�]��9T�W�=����3D���Bɶ:� �)��:z���nۏo(�x�S��$�bd�'�X���	Q.B�8��04��C�HӥIs����ۿw�,a���]R&V�B@hA՜�S%	���q��X+�d�4�¸z ��>c&��Q"�0GT�(0����*d.�Y����~�@(������?t���l܉.�<�3 dI��y��ߚbq�$��G%0���p �U~���y��M�#�zD*��#�������� �hXWbPz�t�2 8D��!�N�B���:��e��eP��Bc��	t�
,P�$Y�h�t�,�i+�>�X��L�J�Аǝ� ?�����9��q�Uߟ��:w���i�h�V( 1���I?KkB�[�h
Yx�<3$���y~������1\�r��)��Q+r$A��&��l��cE�n��R?�
��G3=`0)�&^'^ز�`&D�t S�5d	r����P�C4�3E.K1�Nx�ǩ_=5
�Á=V�d0��ik�����	:hh1Ӑ�ҥ=�)"m4D��k��CryӠ'�pE 
�$��T�ᑤ�4p|9WD�!CFZ��U�HO��XuĚ 7w���H�)Mk�I��'�n��tƘ���XU$�0����b٠SM��"���-JvH��	�J.�����~���#W�7,`8HƏ4h���x�v�[�$�{u��.2hL�P�ޖj��S?
�&�Q���
��1+��� �
�'��}cu�

�n99��U��r}xb��5Sm�@�p���RZRU:mօ%��|j�w��<g��	$��'mY��F8C
�'�4��X�w�h���Q#z���Zb�S��Bl
:m�L���葽d�L1��,&ő��B��Q�Ze�9�M?O����f'�O�q�T͝�79n5k��_K�,�7��u�tH5���
�͑�h��z����=K6�(@hƬP���YEa��UXQ��K�E�<N:�0���Q���IU�?�Y'[,LnP�Cf��1_��(D�0��D��#_������;Wj���"��ٲ�ŷ+m�	�r�>E�d��M���2 JX*/m:-SR��#�y�ę�^��%���n�ZT.M���	�:8��u�P5ax�!h�4��d��o�akdK˒�p?��D�E��%h`��;Jr�m�eb��|8W�� c:C��l��"7���k+B[�I.db:�>�� *t4��b4��^��M�� �36���CE�c��C�?�0�ŭ�3Y�-Y�
 :'@���(l���J�hH3U�S�Os��au���t+��)�@ !,��'����d�o��b�)��u/p�yO�$�����V�R�"��'z.m����9���	D-[�u�Н��3��H�c;���;�a�Ow��h2��{��{�O�l{�D���<qs��&�jD�clU=o~�ʅ%�h�'�<P�1��qy�e�6�|e" '@�c�t�aC>���EK��p ��L��$l�:���p���K~XG{r,S�@"{�mC�k�"&>5K�C�jՉ��Q�Z��H�s*O]�E�R$�4���AX�5U� D�i�lY���v�8���
!�H"nZ,	88�s�*�La���T�s@NB��7R�L͸2�]�ͪen��^�\l;��'�V��Q-Y�a�UM�~Fz"��>X`�@R��j� 
���=�p>1�H�e�.h�0�
����vm٘UFR�h�^z������lՔ��d��t,����0	��5*�j���Q��,?&��#�,�P��UU/����)G�Jx����9h����ׁl�!�ğ%,�@�!Q��.� ��\�u���I���I����B�?ҧ�yG�:$+�q+��:o� 	� gD>�y"�@�	�xI�ஓ:9���OFK�������,�� c��p��\w�"`�ui�J� �$����E�6St8��� O�&���+,\O� �W S2J���R�oJ�_�t�j�⁌A�i�f�
A�4<2�-�*� aDY�i���(�#,O� 4�J�*��\�h�ŬY���!�č�@�n�@"AְQ-ආk*b2���Ȗ�"`	�]�O+�9���F�Q墌���wY�C≙O>-Iƈ�-]�杢��>!�ΰ�1dR�`�N�u�ߪ���+��LD*6�,��	�*�y�皁EƸ,3�"$J���I2�A��y�kZ� ���;�ˆ9_L�+��*���m��| t� "gJ
{)���EW4>(e��"��'x��$��`E�J>�B"<v=�eJ"\O�D/OH`�*��Ն�~L1&镇A�:�"�LB�F���F4f�Ne(�ïq�2�ׄO��ay2	U��&�@�<4���\�k�48ێ{b�T4s�E��Mv�L-�eA��~�DU[�!7J�� 8�A	R����d�ZK�A	q����xr��0U�Hթ�#�%��
A���k%m�i0�a�J* !�P���T�@ٹN?9R 1��`W�ͫAQ�c	���"O�[�h��V�"6"��{���ё���}C���g$~�j��M�N!��D�)��2/(�$�G	�("�4A��	�}��b�N��N�YgN�-1��$U�(��tҶ�w�<�
�a0�O�
��T5L��Ɉu'I�!p|!8��I�=���� e1d�A�����,����pݭ,��BD�L �y"�Q�|����P唹$�Z��ЏZ�yB�Y�VH�SR�9���0wgf�x�a��n�d@�CA/'�bC�ɻm��DӲ#%hHCܿlH�Ol@c�?��<9ń�24^ΑJe&�Fpv�G˚e�<9i�B�zm���� 
�T���b�a�<�PB�.$z(1c���!ZT�cNG�<	��g&1��� W�T#��I|�<)ajG$?��l��$��$h����{�<I6B�%��Hx�NW5�ZӯM^�<!�
�"H�v5"%�
��Y���Y�<� �f��Ss��	$�� �@2T�,����)�]b�='�Vh:�(,D���$\�\�r�U�wY�0�,D��E��n�� A<_E�铴�*D�� ��G�7rfe��&Y��-E`"D��ѣϻf>�\a��+g���&�#D�Dv�oO4��`+��S�.ah�%D�$"H�Xm��&J�0wkD)�F D�`�b�B����6lm:��$D��x%=	��<��j��69�B�$D��:C��f-��9���q�A��9D�CG����(%L�<"���� 6D�4�%�[�j)�I��&qI�4(!D��sQn�,a3ĀP@�\�H�Z��l5D�����5-���+ �I+�o0D�A��O�pnŃa�ٔ/�f�r1�+D��H"fZ�'�%���>�:���k'D�P�ra �I�`tA"��]��m���.D���D.S���G�D+m�t���/D�X��ቁa< ��@VN)���!D��:�H�G�L��S���q�X�S�H"D�0(d#�e�郡��a�����L#D��#щ��~ċdMߢ��I�C�!D���mZ�A@��<��-��<D�le�S�A�3A��`��l�`o;D��He�.P��E;c�V���B�;D�ఇN� �̉Ai�
k��p�9D��І��("��{�m�=w}�@�6D�p �
T�Lu��)Q7e���7�7D��[ �mF2�`��(w�e��6D��;��]м{�Q�I��G�2D�`x���qO��4��&Vv�)�0M"D���h��?��E�e"�)FL~�sT�!D��G�6ޥc�I��;�N%s��-D�LS��1C�\��*j�����<D�ӥ� �Qj�@�Ɯ�Τ��A1D���H��aU� S\�h1�i,D�Pa�V/ R��)�/�ؒ1c�L!�� h�rC��B�hU�$,W�l`$&"O�尃0%�ݨ�̗��$()�"Ol�)v�-k�Fh�u+�T�|�` "O:���K'T�8�@D�5�hY�$"O�I��Z�iԦ)#�כC�r��""OZ��Ĩ)�~����:�R��q"Ob�q+�)�Պ��ʤ`�^��"OHp ��\��1���'.���"�"ON��##�o�^ �����.1!�"OK��NXR0��œ|g����D��y��ez|��$�$!�"\Q1��y"��/jl%*0/��r��V��yBW=�&��@��. ����yb�˄G���a(<i��yWl���yrJ)%G��+d ����#f̍��y�!�5�<ㄩJ��Y26%�	�y2��0�H�J!��.�}!���=�y2�=��0o��W5�qz�)��y����k�����_	G4ب$���y2��S���D�AiJ�iE:�y�(�;>|����8C�t�����yR�ް;�u�7bV?
�L��w����y��U/z6iɧ`�} iS��L=�yB��}����� �~K2<a���=�y2kˮd|";�ԇv��!�Ť�y�%F�N��Ȅ�X?Ѱ�Kd,މ�y­�>JR�XW�+h�K�G�:�yR�Z�j�Dyj�E�1K���EBý�yR��5�1)�"_&�S5N�y�j�6�T�3 Ă�T�p�ā�yrfQ7`�v����Z�p��T��y�oW�-��@���>1`siƗ�yB�X�um>ݑQ�\�A�fۓCЇ�ymJ=o1��{P���	U�u��5�yrʂ�M�$�%: �2�_o�<�0�Т[��Y�Tj�g}���C��q�<��!�9=��`�N
?��,zg�e�<��C�y �`�g9'�J�Ȧbg�<�mG�vF���94F 6bGb�< (ls`c3�ˢ$�Jh�`�e�<Yd�?r4\�G�X�O�X��+Sd�<	�aϭ`�h�ƙ�SB`�5��K�<��jT)w\A�fÊ,*YT/�K�<�a�܋�2i��h*
�59���D�<���S"�Nᑅ,%v���H�A�A�<��o���3����
����V}�/5.T �=E�T�đWzF�{��<����J�y�j��AZ��JuKѳ����F[���ɢf4$+Ao�vX����fث}]�c�Ѯ1���X�$�O`��"_<7�ސ�;�"q�ݠ�sfB���PxrC9q��k�a�x�-rQl���Oj���4xE<����k�84����Th�$�K�LE��y��!%���"Z�~
�ɇä�yr	�E$�U��@Z���9-G\���-\6'd<�Q�ڰ��C�	�DK,D��Wc6(C"�D ����D0v�׷%�D����
P�@t2���m� pfl�+�a~�lE�H�N������]��H��ҹqB��ҦT4T����xl0A�S�ʃU*��a !�+d">F|"�',~~}9���|ܧdɦ]IFFK,H_�!CE��\��u��}��4K�o�cin �d ~�t���,a���K$�ӧ��м�Q�J#xԤ��F�E�^��"O(%�s��3h���i�ESD�p��%�>Q��'6���˓:j����b��2vL>����I!pp�2 @C*����f�H�aA�mH;��� l�C��3)$�M�u'
�Hڦ�	Q"O��rQ�r�`����`��h*2"O��Z��W�zBХ�P���6�ֹ2�"O|;U��C(t�Dp�ƍ�'m
���KPy̓F@|$�3��<k��5�#��p�ȓ ��)�TH�JT���r�ã<.0��'�����E��Fxɧ�4�6�� *,Q1�M:;m@q�"O��1Q$�=j4�2 �E2:#�E�r�ߟس� �(�^0�C"�%)B��I%�:Ց��R�M��Y�i��`����B�M���P$� W�~�3�쁡:Y�8	����N��pe��?7����7w�>�A�BնF��"��(H�TH���(l�Li����k��9�e���EJ�+>��/��y�F�1���y�/�29�P �d-X�K��J�EЃs��	�H"Nӌ]ۄm +[ =(���O�|�� !P��e�#�U\iaV"Od�����4���N���e(��V�>������4�����\�G����������kb�G�N�.5�6s��{BO��T��Pc�
���	+7+�Z��q����}|�)��v��D��	�v�p����g�$RWGG;X����@wk�-���4-ǯ:�4Y���4�F� {��ߠi�Q��!�6�y��	0�������!dK�=�Pd���ԸP��ʪ\�j���
D���*%!7@|Q3���	j<B,'D����I
oǨ��(�%h��S���+o���lڭ-�H�Y�:dɈ�i1����	�ɗbV��4��6�B���ɤH��V"�̟8��[&-R�Y��"S�����ɁRߴq�b��ux��r��:��X��G���:��x�\#t%^�"u(��G�1�h��Q?�Ȅ���qM� �����f;D��Hq�v����v��"jà(9bN��/��0'̿l��8��L�&�L�X��	d�%�O��v�+e�6,� ��G���y�NP�R��2$mc�m��	����Ġ�,S�D�q�6'ظ1���O	^"=16���@����G�V�P��
ZC��̈��}��)��E�*�"t��
-Rx�CͶ
�H!s���E{����'�R�QR
/0���S��8�RJ��r� �tA¢�v��0�J�@���κ�{5��X�I�Ο�y2iLFZD�𨖱�p`bunQ�V�ʤ���D�	�n���$S�Ju),ʧ�y��fF驵��ch�S$����y2�;G "Wʁ�y��[�kȟԆi�s���q�@a��ٹd���!��;E
#=y����P��D�&MΠ2��PK�0y2�ՈN�^,q��δA]b���U�k��bƭ�/8�\��#KZ����^��MS�D'Fdā��IAB�<i0dD_��Uk��ĦDf���'�)j�NG0:���!ÂAʷÜE�<I��]�6�$� �[zl����F?��a�"4��� 3}��I�$N����Ʉ�\�E #j�'6�!����`�I�3i�RXY ����f�&��r��#(���F+~�q�䍎1�DZ� F9��~r�N"�^��@c�'>a�f�'L�Np�֊��	3l���r4� �����~�iҫ_�I��aE}���	gvR��J�Z�'9�T%�w���"�p�� N
�B6��$����2\5Wt��wf�;Zּh��䦙�㌌�0w�ӧh��A�p�P8#��Y3Ã�P�<�`0"Ona�%X�][���Pb��g�*P+��>��D� �fM�v=O��
T��;�a��(�|^��!�'!�YIEʆ5�JI���6E۔q���&�6|H�
O�Rf�Ǻ�X8hd�:
������=�z$s��	�v+��gH;"�T�P���!�d��w�j����N,���L��!�fݸ��I�8"
-X���5~�!�� B�����:@pr�K�?V�!��s-�LZ��N6$�P�H-b!�Ɍ Z69 ��D4̽H��H,h!�D�)s����i��(��	%��<W�!�$���I1֡�V5�}I5��!�0��%�� �s��s��!!��	�:C��!���cw�$����*w�!�d:8��6ȗ�_m�p�%I��z.r����Pܓ�h��� ZD1�Řa=�t*����	z"OX�Y�"�_���i�N�����iJ^X(��\:8r�&���JW�usb>���mTK�A9!f����B1��K���Iu�6?�\��2O��2!�@Obt:d�G6s�!q�W�RbC�a8���PO),O��P�o�s]��s�Ŝ�0�;���X����&���'$�k��ˈ �*`ܠR���0Q��u+�5�B���͐x⧔�O����dhۛ���q'��tR�������37$�*QiUu�}�'jF�g>M3qiM�d�
e�6LظmEBC��95����'�`_Z�Y�!�,�C�i��	�,J�9H�	�f��5�䘖��禑�B�Q�	r`�Ҩ�h�|u*`d3\O� Rg�["Y�ɜ'	E��^0R���v��6Rr(<1�O��zFG�^N���c�'g*)Z�"�g�D�+2O��Hv�{F�%1��y3�QR�Ӥ<��#���+(��s�O�&!F �e$S!l��ĩ
�'�X|�QE���	�U�I����nS��I���'݋>��R�4�*��t�T�e9�I���W�nl�E8�"O452��y_hA�F�g�2=���i@�	cO#�a}��(蜱�O�K��2��}�����A/2<�	���P�QE �Ty2G�B�,B�ɯ+��XS�$/����`�j�B䉿C ��ѣY/ml�u���򄆕2��b����"&t�qC���>v!�C��4��%N(6@�^�dz!��j> ��IN�W(�Qr�cZ'F!�$�8�\=�Q�ʉ*���C�	�!���.l��T��]%���sKO�R�!�W$L��8 ��P�u-*�Q�T'�!�ė�DpN1#��
C���H�f�!�$ѓ=��,���RN���GI<`�!�ʯE�~���T�,&�!SA㞊x!�
�	QFmB���#�l��B�=FI!�$�La�\�6-N!\)N���0b%!�$�|��#��٪D�ؽ�7��<�!�D��#-x� ��r�*�Äb�-@�!�J^*!�\$s�Z��oް\�!�d�5n�M ���"@�Rl�#�R�w�!�ć�Q�,R��>v�u�n[�2|!�$G�h&N"�Ȁ 5{䐃���~f!��[N+�X0C�������ˑ�{!���o�X �A�Z��$�Ѫ��gS!�d͋��@�h�T��I(PC^8YV!���i���a�+�[���@3!��z��8CH��H\�1��3c�!�D�{50A�rMԏ]Vh �`Ȓ|u!�$D�KT��h��_�?��B��[i!���|��("C�7(z`1���
+$!�dX6Q�B��sր&����C�!!�ֻT�~y������c'�(sc!�d�Ǌ���A�:U�.<c��L<mg!�Ę�T*7N�7}������x!�$յP��gH��#~(tC%��Xk!�$	$;���4D�
!,��!dܫ3!!��2�Mr� �LA�͚�!�$�a깩S�b
�h�BK�!�$^�>B�R-�����@K�@g!�.,�����m��ht+��Q��!��"�铧��_b��j��ݜv}!����x�;�f�D��-��,v!�d :���u�X�olJ|�1�A?R!�dć��-�CX����� ~V!�1Wfy����0NF�j�Q�;B!�[D@�������7-��I�!�;bi!�dϻ6=��`Ā�`	ʴ�L9R!�D���nDa�(«-oH��a���Y!�d0ֽʒ\K�0��9S���x�8f�a~
� PQ��*՝4ąV�]�a��Ex�"O��ӕ�լ�wJ@!U�@ �B"O%��O)B�j�t
�-�,�"O�)����>f�`9���t���"OjxN�2d��Y��3\���*�"Oj%"
�(�x��&êK�H�`"O��z��#RV����%��$F�(3"OTE)E�OL��@�J	�� ��"OF�B�\7w'f�X�Q�D���x5"O$IB��ǦkV|3eG��<{|Ēf"OF	�Ϣ&�(;7�)zy�x��"O�)���֖��R��L	S��p�"O̸��GX���n�2[��s"O�L5�U$d�Є�&��)��ZB�'i�A�֩�@�$ӵk���I_��}�U�Ը|X�A�a����S3i����вS�}a7�ʆ,�.�6�K�)'� �Ҁe�ş�ݶB�D�ƸLWRh� �9�vh#4�xb��d��y�L'�Z٘bj2U;N4R'�Ǥq4����͟$[�4�y"��� ^~ם�ӈ����O�	V�@�H���2
�D#!�Џ��Ղ:~�,x�����Ob�q ^*,QY�`�8��eK�OPe�p���:�E�ş�"}jcФ�"ѱ�d�$	
�:Q����:w���4�>E�d��/s�M[w�2���qd���>����"��4u��Q|���OW�D���B¾. ��$IV�@�!�2����'pL�{yA���O�������N����M����'.�p��$�<i�0�_��}��h-[TI!���6���{2 �|�<���D�>l���b�=YĶ��ȓ.)�0rF,O0�Y
'�ٝ!1�u�ȓ�$0p#�G�J��D�$Ohm����0�چ�jخ����J�Τ��`춨��@��f��� 0AK�y�ЅȓD�b��#���5���F�����ȓ
��˄>u�N�`k�*C����ȓ-V��x�n㕓��A��e"O�u�T-W&Y��5o;�h8"O�!Kk�0��0	��0"/�i�*O��I>�t;�c������'g2��Um�}#ZXぇV�ssJHc�'�čaR`Ѱ�FY`���4< �[�'��@yCω�p�a��6.T���'�t�ئ�H�/�RT+&_8-�~Q�'0�$�Z�_E��kU'�	�X8
�'s$���p��1��Lu��
�'�U��R�S�4�6��.l
�'_�����!'�{S�;M|�y�
�'Ě�83(��L\R��"s��0�' qˠ��gB�yC���j����'�hx�f^�w(B����1c�԰��'G�U"�@ڰ&.`;�E�S����'C� ���őg`9ȐK��E��'�h9�^�X` ��J�rp���Qc�<ɷ%ho��s�j��EW�<�Mʼ^V0 Ӷ���pt��O�<Aw�(��(�ܨ;��u��[G�<ٕ��S!}��"�-�D��,�C�<1�m-7�5�!A$��w��@�<1�dX�mJ@����"=�Z�W.Yy�<���#k��k�v�4Ǩ�J�<�a˕v∅��[ �F�*�n�G�<91ʅY��X �i �>H	�� �o�<��� �z�b �eE�$j��u)"I��<���R��Ep��#	� �cs�c�<�5!W�DԮ�7eƥU��p#G�Wa�<1��G� �!U���K^�@��[Y�<I@پ�<��em%%���ZqZ!�� X��b�V!���52P��S�"O�SR�^�7.�8��Gw'vY��"O�Q��ƈf�
����;
");�"O���E�*`���4FD.�윩�"O4M``KәO'P�!&��3c����"Ol`qf�����9���d\I
�"O�)��'XƦ	q�3Pn�}j`"O��q�ߞ3o ��Aa�\Apu�W"OeIh���<I���m]�9��"O��+&nG"G���y�F�T��"OVXi��u���pd�D=�b��e"O�\)e匂g�4��D|�L]�3"OH0[�dЄX+��:P��4���U"OR�9�X[�Xhrd� G����"OrH�hT)zLm�u�S$T�B�"Oز�n?J�F	 ' �\�b�"O����"�A�4�Z�!=~���"OBL1���4����Đ
/2=�'"Oi;`��	l�Ҳ�I�H��"OZt2�J�W�t'���z���!�"O��Wcʊk-�-�F��vZd ˓"O�aK�B�p�|�#%5YG���T"O��A�'7���:B	и6��A�"OԚGh��^���#�� <��	��*O��Kp�h�6��Ƭ��m}���'(iIw �&Qt�j��eB�`��'�f@�%��-�p�u��S>H��TW����yI�Ă�W�1�܄ȓB�dC���h[ԑ��͚;L�x������[)���^8<�f���`��HynH"�r��X1�<�e"O���􂓋D�e�@�{n�!�"O^����+�vQ����8X��1T"O*�֦Ȇ|����$�;�@˰"OT��e�ѡ?|0���^:%4Ҽ�"O�M�`�|Vٻ#�	 ��9Q"O����D�!mj*�d�#qR�*�"O���@�ӛ%�!���
^�D�#"O���jN�mN�"Sd����\�"O���cC!�0y��b�y��1�"O�-�@�n���!���R��"O~i"�'��M(A�����^0Y"O���C�R=I��\a� �g���!"OT��4D�+/
���iZ3g["O�q4Jʐ!�\�1�κ�X��c"OD����A�! �@���"O�Ia@yj@�� ��f.�L�s"O�m�"m��gw��e@6BD�s"O"�:凘�%��/�6/��k"O��`�h�(k�vI��J�,��`"O�|�n�	|��Ǥ�3ks��f"O�Q�%OA)pf1K��$����"O�����0�����4}S�1r�"O���Q@��7NHHgDoL��0"O� �N3S"�L�#�.-x̸�"Or��W-�.c��*dC�<2(X܋�"ODyc�/R!7vTz���'z&���t"OP���D)_@2�c�@\�S� T�"Ox@Qa�4%���Ʉ���8t�G"O�y�� ��ψ��t Y1V�(93"O�h��.d'}r0O^�P:ʥp�"O�,p�ψ!V����Ӕ+�R�E"O��פ��Z�jQɑ��%,��"O�q�� 8�v�8��4#H)��"O� �YSW�Pw�v	�AX;5�8�`"O��;��O�:jE�d.�~��$��"O�t���>P���L��L�\�r"O<`�X"iY�X��J�=ip�"O��x��&l�� ۧ	�|:���"Op�O�9��]��F�:�ҵ"O���V�2E��0CK�x#ơ �"O~� �+�� ��x!u�D�JE��"O����B~�lB4�,=��Z4"O��DZ�+F���A�ųv�~��2"O����&AL�8c@I�!&��9I1"OX��4��6i������7�����"O�p�m	����AjK�Q��"OJ��coD�#�f����)+>nMF"Ony�`�b��h��ɹz+hA+�"O�(�c�H��Y�C��!b\��"O��)+ɤQ�� �	R$�����"Od�挏�dB�`�X�q��8�"OZCO��K�d���n�f���+5"O�k�*�H�R5��c�Ȱ�E"O
��C����ɐp�3z��a"O4��4`��$]����+�!_żA"O�9��)N�f�r J�[�q��"Ol �d�P[V ��Ɨ8sZ����"Od���'N;2�i��Ȃ�4�d]3�"O�Z�%ƍN1`H�v��V� ���"O6��n>K������=Ȁ�C"O�J�BY*W��K��3E��#4"O�I'�	'l���E9[� ��"O�mѶ*�jfUS���B�"O�����)�ۦi	
ead� 5"O� �+�ּ�+�57_*�I�"O��S��^�:���@�	%#\B9:"Od8�v쌵0�z� �&eIRq�"O\��eч�\�p�Ň
P���"O($�b��B�F|�dg$su"OF=��DK�1���# �Z�6�Ұ�U"Or1����23�d�{�D-����R"O~�ѓ�t��� ��d|�U�6"O�,��&�K�`e/�Bl���o�!���5V���d�Z ]Jj(y�f΋ !�7n���@1#7	C��R�C�K!!��O�$(z�H��-/������'�!��9l�\$���8~B�cD��y�!򄈯E8v-yÅ�$8��P$�ݺ$v!�D_bqAba�j�� �O�"!�N�,M��s �=�����2�!�$�j9���P�K�H'�E�e���H�!�d|���Z�f?��S*U�j�!�$N:n̪dy��	;�uH�X/_!��a���0��Z\�+6�G� `!��QdRR�&BR�`�P=�%���w�!�D�9�(`���\�d��OZ5�!�D��C���Y���a�Q�G$ՈSy!��S����
AjP�pȴB\� ;!�4%�,����Ɔ�5���ˉX!�d9�^��Tň�{��xVϕI
!��M��P�0�M�[���i����!�A-2I�	�݃,�R���(˙�!��oY��#E !z�A)CHL�w�!�
��2�[7�[�4zdȐg ,�!� Rfb=x��|� ���hL�p�!��(mfI;�N�Z �p�bGW!�D�Q�C �Շ,=�Ց�$�6B�!�� ~���h�GJ$<�Wb�4V<��{"Of�0�旤r��hXt`��'���"O���'#�-Y���ZQ��,yzݳ"O*��VoPbVF%qeU�<�B ��"O,x�`��;Z���U���\$�yP"O�dZBAY>�tH�ry�6"O���ƕJ����T���_�5!"O���q\R��9�ț�g:P�"O����Q+	�tbČȲ1MLH�"O��FI@/}	p���'zX�� "O���Ac� qHh��+��$W��"O&�YE����f抧%�QyD�k�<�T)�2R������@�E��A�<q�aE?&>� m%)�4do�f�<	d ǭ��ʔ.ϫ,B�;��Xc�<yf��y+�c���vlM˰^�<q"#M���0z��$z�$aYA��W�<y+	�Q�J��@�і;�-IQJ�I�<��%�an(�)a
f?���$�\�<b�!�
�z���=����SY�<Q�]�1[F,��M������T�<iV*�e���c1M�Ue,P��NN�<��o�@�¬Y��>����o�<)tH�?E?� �㋒�|�<ͫ� �o�<�r�á
q��'���1rs��R�<��`�R��q�X8 ���%'�Q�<	ƭ�7=�|�g.{�.�ءN�I�<��h�*]R�m�'��!4gHC�<�4�
�����U[N�����W�<�Ʀ�7   ��   -  �  �  �  }*  >6  6B  gN  �Y  e  �p  �|  y�  ��  (�  ��  \�  ��  �  9�  }�  ��  �  E�  ��  �  ��  R�  ��  @ � � 9 � �! /( �/ �9 n@ (G �O :W �] <d �j �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o7�!Dy�'�L�{�5� p��*кKDX��������8�\�`UBY����Z�h�X�!��oV�y��:�Z��B�%;�!��3$y�TΑ#9LȺD�\1!��	�e���N�dK�ٚA�H8%!�dI.k�e����&,�բ�0!�d@��!���&�fH+I g!�D͋�@�BB�/Y��$��,3!�\
F���+��UN�R#n��V��-�O>԰�H�4U#��C�N��i�B�J�"O,P3�nx�Е ���i�\it"O�$�P���t���4���5"O̤ �&^�$��	�3dD2����"Of�:CH�3K�t�b�����#�"O\����9+Ϛ����@�6�it"Ot���,EMcx񱡡S���8�"Ot��	��K�8-3�ݣ.��i�"O�PAa�;���!aE3rE(�0f^�������L�Ƅ�f��>\�Rrǫ˸C�I��
 �A�K������'F�F�bc���!�X��s��9�����6S���u�'�qO��	dA�i:aB�C~
�s�	(e^���p�4�⌘��h̊"���C�B�:Q�,��Kð=i�����[%M?@��ȓ]V�Ӄ!��P�D�P8`���?�
�j��ү!�ʡ��C-p��r;�L5N�b�ǃ��uW~� �!>D��@B�~�%ic-͍"Sxx�6c�<Y���?a�'I ��n�R�����~A4H�'�$9٠�ޔ-l��t�Ή yVM[���=��eJBӑG^�#&럅n��3�"O� J�D�N�䕐tʔ�.J I�"O�iS`�,�f<x%D����s"O��hQ�T?C��c� �+[�M��"Oʁ�c�נު�P�/G�t����"O�� 	-i�rx�M�Р��2"O<XIaH�2/N�3-�)�vuY��OR�=E��e k)|J�L�i��Y�%զ�y�L�>)<�䃕�.���@���+�OJ4#eC �.6` Z#�F=.�*Oޠ����*��`Z�!@�m6d!�	�'�2U�Q�E�%4<�/��l鄐1
�'�t���B�zSBA� h669	�'����!J�� ��@��e��x�'6�aQ' �T��)B�g�>���'bxY2�X'm��8��[HH:�'�2s�-RM5@���D�:_nl�'�����ʟ!(Е3# #VC,�
�'D�)5�@CLB݃Ir}�	�'eb���ӓr�F�	Ո�4���0	�'��M�����|�qd�a��5�	�'�x���\�c�C�Y�F����'�,<��l� #�d3B��=Y
@	�'�l��ǆ7:�� �r�S�G��p�
�'6θ*��Ť,��x�����;�Н
�'�،�
� 9rAȝ�:�~�	�'H^�2@�/\|Q���(+��(h�'�&�£��3]6�0��
#b�P�U�6�S��?9ҮA.��pt`��9�6쳵͎k�<�"�)b~^��d#Ŋo�%Yg+g�<i��U?�������*Xp�� �\�<�6薰jJdI�Q�w�����WY�<9A�"jС���K��q�HT�<�M"m�b(�#��>z���B�ǂQ�<i�`Q�U���ǎƽ D�-ђ̘W�<��h��<ѐ5��:_��6�Z$�y�g��5y�pc�BM8|�H�8rH��yR	�;CE�Ѫ��֙{�,��.D1��=!�{�	�4*6�:�l��&�!m4�y�!\�){ ����A>�u`@GF8�yrcSv�"ìL*s�0��DL�y�!��T@!��*��XnP��W����� �)�矼҅�B7T�&$١%NY�� ի!D����NT5d�@)�Í͸~W���2<D�t�CbT�i�X� kQ<����©;D��h��J�m=l����J���8��%D���^K��ue7�X7$?D��zso�%4��<9�삚�080T)/D��a���iՠp�!��"¹2�3D�H0!�*UID��Q����h�6D��q!jK�4��q�����c����1D���墓#e �L ͌�K��1C#0D�P�Q'�t���颁��I,�(�G2D�8Ce�,9u�9 ���)4��(#D�x�3�,i�[�!� ���!D�,���/{b^���BG�c���Wf+D���TB�T�@P��.8�Py�E*D�����:R=�&��B��0�7�:D�p�]�sx����(¦�� �P:D�0"t"�>B�tx�1k��؜p��8D���$�	PG�f��?~X��#;D�P�@b�'p��z7hEBuT����8D���o\�F�
$!��C��~�I�K4D��iC�J�$��M�E�B��A*4D��a-�{`����,O%P�4�Fc1D�� l�2��U)Ij)�d&˧"��"5"OT�����pr%M�!6�p�0"O�� �(9߈�ԉdǦ�I%"Odl3�잋�����6X�J�QU"O�� ׈I=mr�@�M� �A	g"O�h�L�l6�A�8->D#�"Or`P�7olA�#���,a�&"O:hٲ˨-�(���<v�:\3A"OIHv�վNjZD�@O1d���iw"O��4"�F0�h)��W(9r�d(�"OE�C
)v��I���h``m�""Oteɇ�
 @^ą"VlXmn q�3"O���7��&;�R�*Ǳ��})�"O�����K� �	�f�A.n�80�V"O|QZ����ܘ���Gk�}[�"O0��A�K�&k���ef	�H�M3r"O���V$�7 !T,�q�Ɣ�D�I%"Oh���N#��x�eY�GFX\�t"O�X�!��DENJŕv��X�%"O❚�`S9�j@�ȏa$Uq"O�0���_�N�%I��`��@5"OYS �B�Rb��J1���:Y���Q"O��`
*������N=P@��"OP��w���*e�e�)�q`�"O�	Sٍ@��d �Ä�'TA{�"OT� ��ȥ=�$�#t,�N耀�d"O��3��r@�եo��Q�"O¹`��5�h�K$�>�"Q�"O�H��D�g]��Z��:؞!P�"O�����Y�K\��B��� �84"Ox�	�#$W��]+e �!�@)&"O���z8^`���B##�XA�,D����8�n�2��
kE���=D�8�I c2ܩ�������f�.D�L�!$�	x�2x��́۠}��-7D��iٶ�y[W.�;�V���5D�L��Ћ0+�ݨ3#?��q�5D�#%��������:Vi�4�B>D����T6o�y!�+�<g
t�ǧ;D��h"�m�� �+9򒨹3b9D���"�@+�:�#qV�?�@}k4H6D� 
`=�4�E��$��T
�/6D��{��ۀa��5�WԸE��PQ�7D�h ��ݒ
��zdD�2lKbx� #*D�X��=^�AJc��Jq`|Z��)D��HOT�]1LI�����V��v�%D��Qv�\69)rU�����60#��$D�Xr���	w"�z"���EB��D�"D���&)�w��� ��G�АC&D���C*S�
�y�T�-�`��W�7D�``q�o��i8��*Kj,hҫ:D����P�:�LѢ��W�J��N9D���"U<t����

;|��y�7D��{��x��e���]"el:D������]��5��j�*[��q�v�#D��0��3�T�`HXOGd��L&D� ���!	�Eyg�U,�(*%�7D����2w��H3�f��@b1C�!6D��S�W�Q"������ �)D�����$��9�+N�J�T�<�Ԍ̹~�b5iӂ2�@s���b�<yŭ�v�� P�e) &+6\�<��nZ+i��"L��q�����`�<�`�A[�V�� �)z�-�£Y�<� ���f��'U������ZF����"O�*a��!!0AY&�çN �"ON�;0d��fOd�)��@:;��f"OV}�aA,P�`�-�Tȉ�"O�l�D��. ��h�H �RT����'B�'��'��'/�'^��' �K�m�]����v,]�;�`��'��'��'|r�'��'�'��Y��U]�z�� *˛j>t4���'E��'���'}�'�b�'4�'��`X���C��{�o�"M'�){U�'�"�'���'l��'m��'-�'s^p�C�3�\�ʢ�ڻ8G��X3�'�2�'���'���'���'M��'�.T�b̨r����ri�.u�$�'6��'�B�'�2�'��'2�'8Z(�A�F�ـ�J�z�t�0`�'k��'���'���'�B�'H��'e���7���1X�
E�S�3FB��P�'�'�2�'��'�"�'L��'Pa
�mPaQ�)g蜛w�B�'"��'}��'���'��'}��',� Ä�ZP8�+�G�7]� d�'��'h�'���'�b�'��'�z��b��zxj�n�*hrt�t�'4R�'+��'���'�"�'Y��'�pP�T��D��A�.�P���U�'R�'���'b��'���'��'
`�BT45^�Xkg�:.`V�:b�'U2�'R�'��'��Lz�@���O.9YV��Vx�Q���֥W;�u����SyR�'��)�3?!p�i���qcJ�B?h�`C��x�  uᏌ���Wꦵ�?��<���P�ĈQ���H�g��9v����?�V�B4�Ms�O�S���H?ё�f��}�L���f�f0{!�ϟ4�'�>�J��M�\����V�v(l��`���M� ��K̓��O�&7=��,� a�~��,� ��$J\��*���O&�dm�D֧�OZ�Y#��i6�Č�t�(�ǋ��&��#��To�s�!��8R��=ͧ�?Y��J  e<d��A;"
��JT�<	*O"�O$mڅ��c��KׇA�B�b1	alP?z�^(��x�b��I��0�	�<	�OL���<>L4)`ԣ.B��a���X���2�>�*�`6�02��`���"��cV���O��8�43�ŖoyBZ�0�)��<у����P��X��1k�L\�<��i���O�-nZU��|r��q�x� 7�6�%3UID�<��?���G?�Cش���n>Y��?�\��L�1��L�s�G_�ޘhrn(��|Z)Ox�������E5~��Ӆ��J��󕚟���4>o�,�<A��� �>L�64�I�q8���@K�t��?����y����'�"ض^DΜ7d�'}`��	&l��[1�����V,Hh es��OΠJ��Y����/�;9*�0�ԋ)�l�����韸�'.�i�	��M�f���<��Աڐ:�V)(�L3��L�<���i��O�9O ���O��Ą���Ȱ�U�@�L2T+e_�!�-h�F�I�j)���4��џ���a]L ��XG� �d�#;P5�C$Hʦ!͓�?i)O"�S�O�P��g�?i�İ���+��9��ybhm��@����3۴��$z����:���@��K��`�'��	ʟ��i>���E�ަ��'E��<)j�!)�)\d�8rk��D������ў�SWy�'IB���	�����W�k�;�'��'!�7-1O��'O�Ha�G�;1�<x"hS��X�'�Hꓼ?����yb���'�"1�� ]$]����3��øo���+bȩ�ON�$���?�S�3���=-�1lڌ@D6@�AS.�j���O�˓�?�|r)O��m�,f����cd�=|�f�bu��(%z��E�yb�q��⟠b�OT�nڞ�] �o�
^X����f�N�2�4�?�vcޒ�M��O8���ۄ��K?�J��Ԉu��
�"5+����e���'���'���'���'�S�(�μ�e�4,�ss#PM�>��۴�*�����?�����'�?����y�%.�"e�a�8u���Y���p6��]$�b>5
�g�٦y͓zaV8@��7�1;3	#�̓�|��b��O�A�H>�*O���O��EӍM�6�0�JєD�I���OR�$�Or���<��i!��`��'���'ʨMJ�&�-C��HE��=+�Y����t}�,h�>0lZy�3�4A��>G�Z��f�5B24�x�7�M�
H�|*V��OdHy��@��l��X�9[�1�Ц� 2bN����?A���?����h��NƒhڡPfQ�f ��Ĕg�t�$��͊�Cy�m�N�杊&�HA��N7GXs��R<C���	��M�u�i��Zd�ƞ���$K� A��%R�`�ؐo�y`tb�g��E��U�|�W���P�	џ��I��D(���;^�YKF[�2̮��G�Iy©l�"exb��OL���O���J�䑑F���C�G@�<��iC"�94���'BX6�ئ�%�b>9S�!��T�,�KT�R�(}2�)qx��I��;?�dl��M�����7�����A���Ls@��O#�* �c*rʓ�?!��?�'�����9�fdEß�`��UĘ���VL�<�2FΟ���4��'98�~+��hj�`<m�!*�.	ر��3r�<Q����<<Q����Ԧ=͓K�8)�'I=LP8�I�y�'ax��s�{�? �qieD�-&]�:P)��&!F�370O����O��d�O��d�O��?�(���&=pX7ҩC�Z{d�ɟ���柄[ݴqO�E#)O0oZ{�	�`����J�`�mVhҷD�:�1I<��i_7=�L��q�hӊ�?%<�B�kP�o���Sb�B\��8���I�����D�Ox�D�O^�$H�c��oT�,�6�ɔ�*]h��D�O"˓G��f.��a�B�'"\>���h��S��,�အT�rU��*?)�[�T��Φ� M>�O=��d�E�����1RrʌP��9A ��E��~9�i>P@�'c��%��Z��S1ڴ鐕���f���cE���	�����֟b>M�'��6�ɾ4=H!B ��7'�\�P�;4��@���Oh���Ħ��?S��lڲi��ơ� ���CW؟NƢ,��4$ћFY�B�����<�F�B����Oy�bF8CD�Z@��5i��U0�JϏ�y�T�����p��ݟ��	�x�O�!1F�}���UoF�*��(1�u�(P����O����Oޓ���� צ��9�̨���wtpq��� ~-Z�4E4�F�=��[�j]�7h����`P�R�p8P�Ö�cr�;�
d��*�*6b!l�	Dy�'Z�Ď�-���Q�}	x��&L'x|��'mR�']�I��M+$�>�?���?�H+��Ix��Z=v`r�'fŬ��'n��l���bg�ȍ%��F�U"3R��8��� �Y�1>?Qq�ڷ9::@C.��2>"�d��?�T��#"�H��2Y��)�$-�?���?)��?q��9��̳WY�&
�]���h^ryQ���OEo�,4m�	��4���yG��x۲�I��'����W��y�Ek��ynZ��M�d "�M��O4C�ß���[P��))�JU.:��a-�&�2�O*��?���?���?y�����CȔ$FJ���$���DJ�(O��mڻV���������b��D�X@���q�T���۰D��8�[����4��H"����Qdb�Ҥ:W�9He��/Y]^I���+-�˓ �Tq�e��O��M>�-O�ea���3�z�$U��� #��<)��?��|�)O��lq����!�BeH3͵.��`�f�3qw���&�M��R!�>ჰi��7�NЦ�:$��>-~�;r��9�.��gn�=8މn�N~��?Y�y�ә9��O����?x�˗�ǥ_��	�&
� �y��'0R�'�r�'@�	ΡEZ��@%-P����)�I����O\����e9#�#bu�i�'qi�7ŖBF�0�ƍI�ڑ9�'1�$\ۦMp��|�2���M��O�(RO�#02�a���r���UH�);�(b��r�
�O���?!��?���R<�d��4r�Ձ`/C������?�)O�nZ�A�0���̟p�IL�l�#J����..�=Ir���ęi}rib�@o���|:�'a�\RV�
3���i�8����l��3�K�r�ܖ'��g؟�Yb�|"�ݥ=��3�cP�Т�s`�I+��'2�'����^���4���5At]:!�S�[2�r����ĞŦ��?�SS�8��4���zq�[�B�\�"oB�h���ihH7�Y*O�6-n�h�	R���0B�O
rȕ'/������o��ʲiƂ $�@�'R��`��ş��	矘�	G�4���T���⢣�32/٣G��t�7�L�]r�d�O��2�I�O�\oz�y`Ɂ@8���̉$*���B���M;R�i O�I�|�i�'հ6Md�ĨE�7i3RuX5�	f�ˁ%x�d��ՂW/�a��@yR�'R�N�`4��^�k�S�j�R�'�b�'y���MC�����$�O�	4bJ3H��2�a	�c�0ɻ�?�����dN��1�ݴ!'�'2��7C�/Z�����#	}ZH���OV�#!]����C�)��_��?YC��O��y�͉�w}����#)������O���O���Oģ}����&��"��/CҘ}�Fr�>���n��MBo��I��M��w� :$���D�,ɐ��H�'�h7M�ئ%S�47GF�:ݴ��ę�-6!���N�&�Bա]7"@pi��N�|��
 J*��<����?����?Y���?f�	2e�����3?�u���/���Ѧ	�g�ȟ�����$?��I9)�JH.D%����'L���Ț��$����4T!���Oz^d㨀^^��i6.�3ؒ��N��
��Q�|K�*�8���W�Gyb&�t�xP��k��4����_�	ៈ�	���|y��vӐi��O������0��U�U�%D[֯�O�\l�W��d4����M;S�i�z6����|�#��e89*�9p���� nc�4���%a��H�K~��;Ob6	�^+��R��L��?����?����?�����O���kȶN6����g��4�UIS�'���'?�7��jh�	�Op�o�M�\�X��EԱw��S��F�vC���M<���i��7M�b�z%�tӖ�I����%�U"U� ��k�a��H�h�)�x|ru�'�FU$�\�'��'���'1<�a��l��3���'T�I=�M���I�?����?�-��a���rph�,�R� 嗟��-Op��k�%��i��HX8�A-K�B�PA $2���Ȳǂ�O��
�m��L2˓�Jë�OT0�N>Im�e׾%� C��J3�y&OO��?����?���?�|j-O�o�}&U�1/B;J�B�C��˽@�r�y�O�埰����M����>¾iĢ;D�Ϝ|�D�&޽-�*4�JzӞ�m�>V�l��<!��}}��� ���m�.O� ؀'(W�{b�5�����鹣3Ob˓�?���?a��?����iۑE7d1vMaD�X���,P7"�m��9@�e�'�����'b 7=廊SSi��+D���=m4h��DN���j�4������O��)�	~�V0O��8'�z�4�X���TV�	f9OҰa�����?�e�1���<Y���?)Ф>:�:��.�9f���x꒍�?a���?�����Ā�=�$����H��̟�{&��[^�$�SGZ�dF���|��:�	7�MKжi���?1�?�\AbM�2\ߞ�wo��<ѱI�O�H)�$g�O�؈���\w�
�I��r݉:��6�bE����N����$�*,*���?���?����h���đ���p�jS�Y�(�cL�T����Ħ�I!@by�gӘ�束~����s�6���� YAL�I�M�i�l6�_�{06�n�t��o�8ۂ� ��k,�95w�Dسț��]@�%�#��I8ʓ�?����?����?a���!� �"8� V a$�H+O��oZ�g� ��۟X��F�s���0�Ȕ��q2�2K�,�(3�����[�!��4d���Ot����e�TA(H�jL�R;�U��Oހ?�P�@X�O��{�-Py2CyӼ�l�m�'΍5Y�"GY�%j�\Y��?����?���|j,O�xmZ�S?� �I�f�Hb��y!�dZvB{+���!�M��� �>� �i��7-�풤�U�BĀ�Æ	+z3�����ȻL��� !*�	�*c�`�T�O\Ą�'K����ߩ0������i�pIZ��zT �	{�l����0�Iן�����,�*D��2VNe1��0k��1�ʛ�?!��?���i��pSZ��h�4��<�҇ᆶ2�>��ˁ�L�����xr�v�n�n�?�#
æ�ϓ�?��E�Q�� %G$X���b+B���� O�OLD�/Ox�n`y�'+��'��NL�R��M�t)�N�x �`nA6D���'��	��M��
��?)��?!/�| ����1��p%��30h��������O��l���MCԖxʟt<#�%F _�R����|X�]��H�3vXhܛ iȮg\ʓ��n�<�?pƭ<�;P��%�C�4]��7"��t8���?���?��Ş��D覥�V��u<�3��&�X0��_�	�|t�'6M#��%��$c�L���V��!�� �, ��@���S�4���޴���B��5��'/׮�[��M�f�v�2=��ʃ�Ax=��i��I��I�h�	�|��t���9���P&�� %
=⡎D��7�@2�@���O���7�9O�lz�#�τ$/}�t��IĽ����aڑ�M�p�i��O1�NA���z�6�	&6�Z|8�@���R%p�bM�Q���	S! ��w�'2�4�'N7-�<a��?aB��!&d��V��&3>�#y�u����ߟЕ'@V6-N�Z�����O"�Q�+6��Hܲ�4xP ���� :�O6n��M��x�
 7Y�b)H����;�2E����?[uPE��*�#)���6�����?a���O��M��{�Y$g�.a3҈��$�OZ���Ox���Or�}���n����X�0��6bΌUG�U�����_#;��ɔ�M��wN܀��&S7�9"'�	N���'^,7���Ձ�4�[�4���+ڴ���Pn�%ɚ�Ѱ���#��A�A�<�g�i%�����	��(����d�Ic��Q��G[��x�{c�ӯk���'ߦ7̓�k�x���O��2���OR8S�E��F6
.`�T	9���Yԛ��b�,-&�b>])�킚3��X�D�$,�Z䢶N7 �t�:#N�Vy�Z.P��T�I;�'��	�yoL��%�2cTtZ�lN^��������Eǟ�R�-+c~�[R�ǪL�$u�����Ԩ۴��'��ʓ�?�ߴ\B����!�=2r����=jt"�T�~HZ��i��O,���Ƨ�Rd�<������f�D<Ky�
���,$ԡ�n�<���?����?���?y�����=�@��r+�4���@�H��_LB�'���z�`Z�;�J�$�ভ&���E�ʁpSNҰy��i"��>���?I��|$i:�M��O����Zd�b�l�B�6$C2�T�"��x���ܓO�˓�?���?���0�L�d#�{�������g�$����?Y.O
}oڽI���	�|�Is��Ɠ�bQ�L+e L�K��7
���'DF�z����O�O�韎�����6��g�Gg`�r���A�t�;�+�v�p��.�O�9�O>�P/�I7��BV��/b�bq�fnF��?�����$�O1���.ٛ�Q*Z) �z�g��TlV�!��ƠA���'z�q�Z⟜Y�OLMoil`	IR+���#*��8Ix Q�M��(m�#� imZ@~BDI�<�~ �S�$t�ɤ[�m�B�
$/��a��ƄQ�P�	fy��'�����Ŝh�t�5��<<~���uӔM�Ob�$�Oh�?������cc�y~ X���V�F��X�m�*4�6�o���&�b>�� ͦ�Γ�h<A�d��/Ɋ�	��X]F��FJ������O���O>�)O���O<�x�&�e�^�!R���v�ӆF���'���'+�	�M�'��?I���?�H
�')XӴ�ގ^��0�uhە��'4H�,���{�|�'��(���o���a&��/bX�-#?�ƌ&�h� Z���5� ��[�?QE�N���#�V�)�����B+�?a���?����?!��)�O����%�"����6�y�2��O��nZ�
��'�>6�-�i�ǢFghƵ"H�
G*pU� .v�dX޴vᛖ�q�N|HA�c������c!��F�� &�zV';g_��9�ÆJ�Blr�;��<����?����?����?Y�͎�AE�xy`o� ����c׼����iP��ݟ��	�($?�I�x��	�3�>7��-�OL�Lh͑.O��DoӂQ$��)����ɃA�f`I��/�XejՎ�1hD�D!��S��ʓM�^9R��OR��I>	*O�]�vhE�7~uj��B���!hi��$�O��D�O�4�6�4���b[:4�2Nܗ$������xB�E�H�<�R�~���,��OD`o�.�?	�4�F�j���X��R��E!+A�R'�/�M��O�`� ��!?����$�b�+i��ؖ�Ai��Ɉg6O��$�O��d�O�D�OJ�?�K�
�+6�f����$c4��$eI�����ȟ|S�4K�(�/OB�oZv�	�j��!�ɋ�s����3��Xt��N<釷i�d7=����D�a�d�r�~�Ñj�T#�����X�uC6�i1!C���D�����4�����Od���%Pf�0��T�$�R��Qq*����O��c��'�%b�'�rX>q+���1yn�����li�VI#?1�U���4^G�&l>�4�,�)�^�9���
9^�&���{�œ%.$\ ��(���KTB!�k�I6%�����C�6s���צ>C�)������Iʟ��)��_y2�`Ӯa#R����ؠ�1�X���1���-���	����pyR�iVpA��� �e���rN�yGw��l�%1��ToZ�<���h-x��(�����'�8�"�ˌ�b�r�R0��A�4��'��П,������X��S��j�`Z���N�v�3�N�.6�0l��D�OZ��5�9O^�nz��)�՞��r���	�Th��)�?1�4R�ɧ�''��1۴�yr�߁wzi�u�.��p� �
�y�g��Z]��2�2 �'YZw��I�O�QS�ދ+�����߃&�T��.��J:�@C���Ov�$�Or�	����0��<����?���
q�0 �	�]�t@�UIJ�?!��?��ثGjZ9Ou�D�i�D���?����Y��IТ|���Ğ#+�9�3ON�D�:�D@��7x���2A��
�u�g�O6M�g��U�r�b§v+~X��E�O���ON���O\���O�h��m�O�� d��O4=�5�!u�A P �(r!�D�O�!n�^V�20�09O>���?�%�їx�ZH��L&;��5g�#�?��iP�7�����
_�]̓�?�CJ�a��1�%"���\�@%Z�	z3II�L�qJ>Y+O���O4�D�Ox�4לּ�	d�`]3v�|hu8��<ѷ�i0N�:`[���In�'Y�*�����Eϰ�Z`��%�(T�[��`޴U囆�0�4���I�.Y+p�ʍ=X�q�G"��ґ���4(T�(�<	G� ��d������Y�&�H����#�0|�ed�'��D�O��OZ�4���	��oʫX�2�	�&jE��>Cv�A��V�y�Nt�㟘	�On�n��M��i��5���+7=���à*��3t/Wi�f��hȂ�P�q���_����E+QcG4�(r'� O#LD`��p�@�I�\��ɟ����t�
��]�D��$G��{�uX���?a��?��i.&ى�O�!j�z��<��c1���ַ���a�(��]���x�)c�l4n��?�)WNFզϓ�?��#�1
aa�?4(�,¢T�\��#���O��+I>	)OH���ON���O,�i%%�%�>�`	܃��|`%��Ol��<�1�iF�q�R�'���'|���O�Rt��[6aي4�Ԩ�!<`���O���'h6�_˦��N<ͧ�z1D�3+ 7�J�P� �# �'#p�P2+O.����?	@i%���eshd� ʆ/|4(;��<*��d�O �d�O>��<鄼i�2<�c�#�r�iF���{Nֵ��/<e��'s�7��O��O���'����
<B�t����d��)�FMNͪ6MԦ�0�̦}��?� �Qn���5����:�� 3Lp��6M��y�P�4�I��,��Ο���ޟ,�O��4�Phc��su�8I�C�kl��I�r��O���O������X���]H���k�c,�0�1^�Y��E2ٴ`>���8�4���i��8�"d�c�d�0�1��4:��m��L�����I�8-�ٳ��'���'�̗'���'��iq�?4V�}�����o�$q�'��'�S��ڴ\O�y����?����� 5��"s]��z��^S�������p�I��M3��i�zO�Ȑ3E�24ll���LoPr���?On��&Bk>�0�ǋM�ʓ��%��O(�*��'���Q�G_�V z�`-�x���O,���O��d�O&�}r��W���ŀ���1�[="�M!�	u�F�<�b�'!v6�"�i���J��S��P�ĉ��F�����z��"�4z��i`�����i
�	Gr��*��O��<K� BV��}��mK6i��iy /�a�	wyr�'4b�'�2�'��D+>�P�e!s�\+が*3��	��Mۓ������O&�?�!�d\��'��A�4З��������4����O������yX��W �uy����v �EQ�|�����c��`WV�	vy�
1���r�R6Dr��Ew�2�'��'��O<�ɍ�M��"̻�?at�ƙ~.DY��UF���&�8�?�ói�O�}�',�7�Cٟ�m�3�`ѻ !Ҡ>�)Ӄ��<R��tmSʦe�'�@��� L�?����T�w��5��j
9w<�Y�J]�:h6�'�"�'�b�'��'�R� ���A+�!p2P4]y@��s��Ob�d�O��oe/,�̟ Y�4��P�څ�D�ˤjV�T˱d\;��8՜x�!i�Ԡo��?Yk7�צu��?!ŬDh�? 6P���C�_��H��ޢ ) 1�����?1�"���<���?y��?���\�*ap�M	4hu��B����?a����D��=�w��I��4�Op�p��v,у�M۳S��p9�O4��'�6֦�H<�'�"$��-w�P�@@�&��B�g2x��'��m �*O���\��?�##�d��=6ZYbԋ�$VTe�d&]h���D�OB��O���<	�i*���VK�:B7J��*;v���DM�j�B�',t6-&�������ڦH�.ؤ��EJ��� @a����bR9�M���iNX,���i��I%f�=RE�Odౕ'��+�Z}'x� ��m���'3����	��x��ş�	I��E�5r�#`��"{Z���CD\�7m�Ud���O���+���O�oz����4PPzm[V%(-@�K��Q��M��iٔO1�2�	iӌ牓s ���4|�zEÅ%�>i
�	=L;^�ӷ�']Ҕ'���'���'`�5��-1�<�4(vbrE%�'u2�'�RR��PڴW8Q���?I��y�l1���
�:7@ܢu�й��RF�>R�i�7�@�	�	ʲՉ���'6�8��R3��7O�m���#O�xt`J~2���Ofth��V��J�H���@��$�����?���?��h�6��_�*��3�O���D�u��	��D����'�V֟��	�M��w�>H���ј�M{�D{4HX8�'h7����4Z��Q۴���H�Q�T����nU�%���[��ݱ�lB?:Ԍ���1�D�<a��?	��?��?Y�Y�%��Y0�e�j��
Th���?��D@:��0BqL�)�?q��?�3�i��s�$�"lS�2��PJN�<�u��IɁ��D�Ŧ5bٴ
s����O!�T%�<h�b+,_8�"R>p��=2��.2��8 ��bv�'���&���'ł��U*�$^XP)rңF1f_@�"��'���'q����^����4.n�:�OA��#�H�)wJ��g���V�E�S��&�Ec}rGp�ZXo�+�M���/D���ڥE3M�l�r��?#���ش�y��'j� �F��?��_�����q;�Q�=���Y��ԪH�*�(��e�P�I֟������	�������wz����$ :*�;�ɉ��?Q��?1b�iS\y��O���}Ӕ�OXh�u��[�zD�#)o��h�6��v�I��M#����O,S������І���b�� *=�<``i۷�f`Iq�/V�%'�p�i�7�O����O:��_�G��RSjZ_h�LIAB�sw
�䜞JZ��d�O$�ʀ�N�n��	�O������3Q{Ҕ+�ˊ0?i�Z��Ul��Iɟt�I�<q��Mg�i=Y2�S>)��F��1��C1^���DTv˘!j�)�mΐ�3��My�OP�C�����%��&��̚���oGw@8�I�+[��蟰�	՟�ǟ ��Dy2+ӊ!U'�!\X
I���3�x9��;{t���O��D�O���|����y��i�p �k�[��d!U� ?ڠ�¥�`�am,F��en��<�޴ ��(����R
Hx�Y� yd,W�,;w���\A ���<Q��?���?���?���?����?���BB��,�)�L;�5R���'R�҉��A��On|����?Q7�i���O��f�O̕I!�Tax=z�m�{��&�Pئ]R�4<��6�;Bf�O��T�O��Mzշi��$E�`X��ďQu��A��<8}�$��Z�f`Uk	ȒOn���V�'i�&
�+`|�e`�c�p�{wa�);^��'3��H %�I�M�Q"�����?�4�!(��&l�08�� I��D��䓸?1-O ilZ��M��^�h�ɳ>8�Pâ%|k�b/m�:��ٟ8aрW�?�j�Ж��cyb�O������9�I<�rr��$Kh8�"tbŹm������h�	៼����ɘ4��ؔO������p�S"-1=d9A
�B6�On��376O����O����O�ܦ� u
J|H�h��Ѣ�D	VޱZ	���	��M�iy�7���7�m�,�Iam䑃e JbH�)�����}���]�I�(
3�O��My��'/R�'�'R$� ���Q�&�h��`�m2j�Ɉ�M+�"��?i���?AK~z�.�&�0�G̘(J��F-���e��]����4���x�O����OsM���՟.���De�<<���Q:\���^�\��/�Dg�i�IUy\
��L�2`̢Bvt�z�ŉ�0>�a�iP�Mh��'�^`朄I|�,X��$k�j�R�'�7�/�	��� 㦹��4h,�&����L���.!�(@!cS"-���P��i��ɎM۰y��OO�1'?��]�r� �W`�EM�(
���>�|�I��L�I�,�������[�'C�b����|	6��7$˃u��A!,O����ۦ�3w+*���i��'|�C&���$@r�� ���	��8�D�ʦŠ��|�*���M��O���Ҧi���c$�&<�zAs%J��,�i��7FP�O��|Z���?��q�t�{q(E
RTJ����'4��J���?Y/O`lZ�r��m�������R�$L0a�d�s�T aS*AP�(�4��d�`}�e�,o���S��玤v��Q ��*尜*�uy�h��H�X��O��Б40���� 0�I(t'V$�r\x���� ��?I���?���|*�T+��K*OplZu�
H3��
�ae�I0IK�(� ty��'Z�'��T�4:ܴNHޔi�ʎk�0zP�J=P���ɣ�i�X7��%�6�w���I+V�l ����*A�� �D���B-�Is�cѴA+ ͓�?I���?���?���?q����* �"B��=2T����g�Zn�t��@Ь��d�I�?��Oy"��y7�Q�"��d�����C�[3�7-���O0�4�*�I��ByI�`r���)� \<9t%�P��������ai��7O��K��?���(���<�'�?A'+�!8��31�P�D�ʕI!��?Q��?i����ŦI���Hjyr�'U,�Z��\�U��xTg�%G��B1�$|}�!|�j��	z�ɦA� 1b�Z�9��Q�@3m{��s�"O�(���N~�p��O���'SBp�����Q3&e�"PZ���?y��?	��h���dA)f�HL��R���!�U ���女#щ�����I!�Ms��w0,4)>%NzIC\��]�֮x����47�»i�U��i��	^�%���Oل��!��2WU>��/ʀ,\pbD��M�IAyb�'�b�' ��'�L��KF�����p�T�D�>�剆�M�d����?���?�J~��<�%R򂖚fKL4pa��[�0��R�4z�47�2�x���,��X<8��Լo�(J %W�W>�T`6���[a剕\�^�2�'Bn�$���'�e��o�g�&�h��Lm^9�@�'�"�'������]��b�4A��e0�j�Ԥ����Z���sa�F��VA�ߛF��}�r�Ƥ�	�!ؓ��'�"�R1hv��7f]�da�InZ�<��
�&�������Ep/O$����\ڀ�O�7f�tHE�5HN�r0>O��D�O.�$�O8�d�O��?���������+�(UV�Sc^����	ٟ�3�4#)�ϧ�?	�i��'��`��-@�8�x�^��j-�$�O��O7����i���)4�h!���^$�B@�@�ۯ�H����B)Dv�ey��'�b�'�"!�. H�h�)Gb�̈7�ۏ1]��'��I�M�NЈ��d�O�'Wt@2�(5�eKCmH a,��'�v�Q/����OO��!����D�m�L�$m��b�N+Z�Y��vy�O�du�I��'��e�+�>N�q�ќL�����'��'�����O��	��M��%��&\��43(
GM�<�����?i�i��O���'X6�٫6�%���ƞ<^|a�m�+3ڱ��¦�`�-�]�'�������?a��R����Q2��P�u�@�-��qd��̔'D��'���'E��'哼~���:��شf�y�z���4~�F�p��?Y���'�?q��yG���*�������]�V�a��֨�����O��O�On�(��io����P^ll[�H��}�<�@�O=(�ƶM��j��h�Oʓ�?1�'�V�AP�
�Ș��)���5����?a��?+Odm�P8NȖ'�$��`LDtBci�����垲yO�O�Q�'�@6�BĦ�BJ<as�D�"�VQKK�b��2V��l~b&��b��lZ5�L���O��L�I�}m"�ƆY�ԕ!��G�TRm�����y|��'��'b�SٟD!R��_��s M�+ �$` ��֟d��4i���k-O��m�V�Ӽ����R�t�����H�QB��<)��i��7���u��-^���'�ف��H�?�,IN��qWbE�G)K��H&�P�'���'/��'���'��x0�&��5��ܙ���&'fBe�P^�`��4Y�T=)+O��$2��hYrdvl�\�N��RM&p�/Oz��~Ӕ<$���望��ҍmO���'��C:�� �(�5�bܠv@�<�ڢ_`��dہ����D�[h�
�F[N�25j ���@J��D�O>���O��4�2�g�����%Y�A�=z��㵎
�P����!ĺ��z���̡�O6%m��M배i�M��Ĥ>"��c$�� �pE!��V3O~���&2��'N}�ʓ���;k�M�1�ʴQ\B��	J�����?����?A���?Q���O�����*�V�H��ĒZ<��8�'�B�'v6�МF�˓!���|�k��.^��$��#vu�4�5m�8l��O�m���M3��� ��4�y2�'����,	�JDּS"b�oJ���*Qd���	8%o�'��۟X������ɵP���P`R�&�bU�p-� �^M�	˟�'HH6m�v�^���O����|Zfm�+�F|���
-b���A�j~�ɱ>��ik�7-�|�i>��S,ݰ��ψ���Ģ�����B�H!�f����Fy��O�lX�ɥ��'��<S��I�GV�ɘ���O2��	�'��6M̴&%3D��F�i�'�M��{r��O��dA�?)�Y�H��4?�p�o\�g�̭J'�9����4�i�7-O�!�6c���	
}+�E���O���'�48��Ϡ<�P����M�XY��'�IK��ܺΎ�H�Uڵm��A��y%@M��MS��Q"���Oj�?=c���SR��%w.���W@�z���b�*�u���e��$��S�?9���y��o��<�6
�1R�.�j���OryB,F�<i��تF}R�Ė�����<-Þ�s%g�D��b��?Z�t��$���:�������ޟ�3q��$4��	PG��)5���@�y�������M��i�rON9i�LK�u(D�zB�: ����e����u�'=�Q����{�Ӄ&4�˅���t��s�*�ك�ޤw���Ӧ� 蟀��ɟ,��韨F��w�޴�@k��h�Ne!�E�('�4���'�N7m?0��˓6L���4��uY�̩l'6|��!9I~�3��OF�d�O�6��%_Ǫ6�$?�rDP�P�`���\�HrgEx�!`e�ƈEO~�*J>Q-O����O��d�O����On��D��0�y��j
6ʢi�<q&�i(�[��'���'��O��O��D8�f�A�vW��W�Z�TT��+	�vO�O�O����i	�2� Ș���^� +~���|I��q�i�	A�|�c$I��O,ٺO>y+Op�r�Q,*ӂ�C0J�M
����O�$�O��d�O�)�<A�i����'/N�S%��0<���AA�)����'׌7�O:�O���'"�'$��(��
�PLBꆗ۰��  [6! %H��i��O�`K!��'�:2��<���ǿ[�>9�`\c ��	N4< �`��<����?Y���?���?ي�$��Bh0��d~G����j�����'F� yӪ�x!2�4�dަ5$������'L��f��R���� ;��_���-�O��N��b�������
��$��G2bT|z��ŦIF0��Q�'5x�$�ȗ'9��'�"�'ǠܳAG�6i|�0��'ʡ\�Z�!��'DRU���4	>V�0���?����iӽT�|�qQ` X
J}�Ō�i��I���� ���4n���)"��Y�W�	J�)�䝪K�:���-O2��8 ���Sd.2A�@�I"J�Y�N~[q�p��?^-<��	П��	˟H�)�SAy2w��@��'�"���3 R$"�!7��� �ʓ	2����SD}��w�	���[�@����@���Y�/��A{�4���1�4�����|�������	"I�Yk� Ԋy���bK&U-��	uy�'���'�R�'�r[>��HځJ�x��r��_.�)�̟��M��oU/�?���?iH~�"ޛ�w���r������b���jQ�IB��x���l�?��Sܧ7� �o�<�Q�̨*{Z� ��h��s�`Γ({" A��O��{I>Q(O�)�O�=��j5d�$�B��e�Z��T��O����O��d�<���i�QB�'���'dL�*g晄��܈�^�]-�id�d�z}b�y�,}mږ�ē/��4����C��j�E:@�`�'��-;��F�V5�I���D�F�����'@����+	�7~��2 ǈ\���'���'$��'�>	�	�{h�b\�\'$ف֣j6��ɨ�M˗�΄�?q�Yԛv�4��@橑�-���1� ;�<��e8OZ�o��r� �¦��� ڦY�'$���?�T���
EiA ْ{�������;d�'��Iٟ(��ԟ�����ݧS���1��[+�]J�k�v4�'�67mM.q9��$�Ov��4�	�Oܡ���8(���2���fq� �r}�J|�Emڮ��ŞI�����	=B�>���Z8R�Ι*l�-'���".OFu�`J��?y«0�d�<g&��!*r����|�U*W���?���?���?ͧ��D���y�	5�'�ؤ�cgI$���eC+�J|+t�'��6m1�I���ĒƦ�9ٴ_o��(G�y4���%�>>ߠb#��h��Hĸi=�I`��I�Q�ON�h$?5�]N�t�"�sb�dZv�H�=�l�	��I�d�I˟p��G�';���H#�^�g�>��p)I�xD����?!��-��V�L�����'A�7-*�$��"KD��4
ߝ��T
�m�<ϒ�'��ܴ���O�`��i���y���P���J�P]bW���sH�7�RDMu�LyB�'8�'s�Å9]��I���X�sܔ-ԅM ie2�'C���M��.�?)���?�*���VD��n�xa��\u�Q%���/O��tӤD&�ʧ ����J�!B��lB��V�T2 
�yT��1n�4��4�2��2�ғO��3�M�\�<C1@7!HPjOdo����h&��B�lJsh�%��0$-LKy�Ai�2�HJ�O�n�
B���`��kL�E�lE�M��,	ܴ�6*�g��6���x�HۑjE��lEby�J�a�t8�왢-�,� ��yb\�����L�	���������O\T��
x����J����b�`�(P���<�����OR�6=�B�bE�b@xٳ��<+���$����4\����O:�J��i�:|�� +L�U����u��G�������!��V�O���?	��>��P-�8Έ��$�G�r���Q���?9��?�.O��oډn�����	�'A�9rAʄ8vu,�ybc�$���?q�V��h�4!��)��݊���`؏2 �� H<I�ɲM < ��(f'?��P�'x�I*�.-���p�0�ȫ|�f�Y!N�������d��ݟ|F��w�pQ�F��	J����Q���b��'JT7�j5zʓ6����4H7o�;A�q��C�6����:Of�o��M3��i%B��i���;l0x�1��O��%�B�L�E��9W��S3JRb�Dy��'or�'r�'��f�)E�"Y����R�6�b!c�%?Y�I��M�q-\�?����?�K~�	~:�r�!��uV�%J�/ǰu��	��U���ڴD����;��	ڄ�xWF (j! GM/5޴z�mӘ�
$�(O��8�
�6�?ِ$*���<Yd�:u���Є�-{b��V�S��?	���?A��?�'��D�Ӧ�A�Pڟ8ZWǒ7g�z�F�I<�p}��&m�piߴ��'Ҝ�$��/v��o#	`�(��Z�^،aѤ�U�`B�c���q��?ya�ϗW?��5�������+��!��̆�s
8�'MZM�$�O��D�Ox���O:�!��8�RT��#��֍{f��5�$������I��Mc����|��:���|����3n<i���g�D�`C -��OX$m�>�M���'��)iܴ�y�'��99S�,2��|�p �/T�|A�Ҥ(����	N�'+��ӟt��ڟ���gZT�R��$=f��s %Ow� �	🨖'g�7ʿ),����O��$�|Z0�G�+c�ۀ!^t(��P���Z~Ri�>Q�i+�7��X�i>��3� VЋg�E�bXe�@�<L I�$�&��W��ʓ�Bw`�OV�3H>9'A�na�l����$���P�A���?��?	��?�|�(OZ�lZu-�-R�K�r�a�%B�{=5����cy�	r���T��OZao��%��Y餇���e�e�ӈ(�H�K�4*��VR�vڛV��@�$���4��Zy��Y
aXXQLG�7�<%����y�U���I�����ٟp��㟄�Oce@�jD6�
�,T!/�����y���S��O��d�OΒ��$T���%fe��Em�2Ȭ@��ɪb�Ph޴2��F�,����__�6-a��37�7��I�fH�4$�[R�d� pcA�#i�B�y�	cy�O�Z�9|fŠ�/�#M�r�1 OL3~�'�b�'��ɂ�Ms@�&�?A��?�Q[�G��ǀ��T��� ӓ��'�D�]E���a�Z�'�p��N��V�<�KG��5*�Ҙ+�/3?��U-S���Q�]t�']���d_��?b.�.3iV�jg�'*�0��-�?����?a��?���	�O���C�2@"N��HW��Uq���O��oګN� a�'��6;�i��i�������ϑ�0�C�e�������!ش���4����%��'>�(���b�?Q�f�Z��Y�^z�"�$�<ͧ�?)���?���?�Z�Y�D� c)\�hP��d���D��u!���ΟP��%?�I,)U��&�)�V�����8J����OH�l��M�x����yq-�&d0��=G�@�pF���ٙ�mKUy2�z D��ɵ-�'%�ɋi����G*�e�Ƹd$� B*������)j�˟��X�B�*�)���tؘ!�6%}��2�4��' 
�3웆�z��lZ�o�*�f˟qy	�d�e�Ua�KЦM�':����?��2����ws>�r�F�^߆<-��a�S�y��'�qqWI��CpV��m����b�'���'w�7�I�VU��?�M�K>�0aY(�2��B�Q��D]K�@��'��7-�æ�S8��nZY~�aP�N��.;/ThD;��/p2hEy2�����ґ|[�p�?�d��(	�80B敟5��m�%,
S�'��7�E�v�d���O����|��([�Q�
���'0�Xk�,H~�-�>i��it7-n�)���ݒo�	�Uj �21\j#��9nlN,�G�S�3�j)O��ݥ�?@�,�䑘!r���s`�Zk���1
�G�B���Oz��?�|�+O�9m�!��<����ny�L�$�Q|fn\Z'�SyB�vӺ�h��O�o�a�P�B�C�w��)���u�Pp ޴Uk��Ϛ+9��f���Z�Ov��D�\y2� e�xX���4y��4�y�X����Ɵ�����I��O2>���R>5�B����3=���gvӾ0�F�<Y����O@6=�6X"��
-\nE:^w-}�bǺ��F��O$O1����` f�F��#r�N�8 ���X��G[
��ɍs�0%(��'�x�$�(�'-��'����t�]�L @��9N�~mS�'���'��^���40��@���?a��{]�% �!?L�HY��B(����B�����M�ưi+O�$��B�=�U+vF��#	K!>O��Y�gE*��0�b���$��OR����@q>��Ɗ��z�
L�ʊ!0���?���?!��h� �Z�W����5G��%p2�"�䚨@K���Ŧ��!NǟP���M��w=��*A�P�b�4���RP�I�'T7��A��4I?���ߴ�y��'�,��aa��?�*��C!HKL����)7y�Pxb���"��'z��蟴�	ڟp�	��i=4����7v �i�b� &���yyR�w�`����OX���O�����\��Y*BD0z���w�_~J�u�'��7M�Ѧ�cJ<�|�W�ŤGL���ŝ	��1�5n.]�J� �d8��׸y�L�b�G�OH�2�hE�%"�/]^��r��H���l���?���?Q��|-O�Xn��h4��ɡB<�U����&�R<��	�MÏ⬷>Q�i��6m�Φ�ya̅*���5�2}k�R�k(�<o�E~bH��u\8��xܧ����([�!���h�����ųu��П�������՟���A��nW��k��]�l�꘻ �	(v����?��/\�F�E> ����M�J>iuK]��J���ʶ5#D����]�V��'�N6M��ə=�V6m2?YuKC:I��Z!�	_J4�홟`�*�p��O���J>A)O���O�$�O$$R��Ȧ2�s�+��4��A�O��Ī<���i��M��'S��'��S% ��j1i�8vyB���U�B�hS�	(�M���'.���	]/��0i�HZ���ڧ8\��RV	� p�$5 �
�<�'���V����� ���E� �ڄ�"^l~�j���?����?��Ş���N���B�:2��7���00�X��(<.d�'��6�'�I���Dߦ��Q�pVf�9��e3�h�H��?�4?&p���4��d�8S3�8����˓<�
3$N�:kjpU@�ADTΘ���$�Ov�$�Of���O4��|J5.ֆ_:�ՠ�j��2t��X�G�qϛ�/;�r�'�������݊k��T�p���R}( ��%l/B,�޴:b�x���/¤j@��6O���p�2J����J�:	P�JT1O<(#�ꞁ�?1 !���<I��?� ��XH �u�J�+!�U�bY��?���?����dȦa�U �ޟ���ҟ� �!�;> p�3�ϱ,���{��AO��1�����M㢷iŰO� �,Z#��$U�)tƍ�K�Bhу�� S���5������A�S�5�(=1 O�~L@�a�)ߞ���4vPZK�K�
D@�nO�~"ԙ�F&Ӻ���z��#�ΤHgß"Z�}�"N�9b��RDB/Gl.� e�?:���V�"\�Ld�ǨO:��3��h������Z "�a���
���Af
V�Ģ�,Br���/��Ddg�F8r����躑[R�JJR���G��G��r�
v�L�9�)ՊR�<]���� 7�PQ��K�	�
H$J�@}�� b���裨��}��ـ� {��W��90��3���6�jR�i�R@Rv��O����O �Ok,�J� pӨѺQHx\�_�5��f�'b�qh�'a��'���'��'l��ϴjȈ�b�E�,i�\@"(�������]���'���|2�'�����\/��R������\�4�I�}dZ��������OR�d�O����O�m��Ϭ?�!��|���oֽr�:�X3�sӚ��?�N>����?�$�>b:�o��h��beB-z�f�@��E�z�v듀?���?����?�wh=�?����?�GK�b�����E�P��)��\"��F�'�'!R�'�f ��e���ēI-8h8�,�eF���0�$]P�nӟ���֟�ɵeZx�O_R�'��@Ö#z�B�&��?ʄ�kP�7�XO<��OF��&��'�1O�$B�|�q���iZ�b��"C`6��O���ԅ$��$�Ov˓����?����Sb�]�3�8���I��B˦I������oX�HH�b�b?�"GGE��Ny3�����b�b������O��d�O��d�8˓��I�
hWJ�Q��̳|Rt��`A�IXH�oڋ�a�a�5�)§�?��gH��(|z'�u���Fa޲-ě��'���'�>�R6�8�I�����r���/S:>R<����i��>Q�aU̓�?����?��F�k��C���A��pC��+g����'�ꐻ��>Y.O`�-��ƒ�+�|� {䖸cY���V"A�	�����Ɵؗ'�@ex1�.�]i��s�^y
�B�����d�O0�O��D�O4��n�Gk6�I��L�#���1ⅉH��O����O��D�<ɴ�ȗ��t#ޫm V�ht��1@�`��⃱�MS���?Y����?Q��pɌtq���|����L���=N���QZ�`��؟���Ny�f©\�d맟?���?(��($,�j@�SB<��'��'��'��j�DB��84�"o�%[،��� n)��'lr[���1�M���i�O����JX��Ӭn,dj`Eɳ)}jF(�B��ҟ�I�,�*��~�$-��	#`Xك#A13ʠ��ڦ�'y�E��k}�z���Ob�$���ק5�,�+H(����,m&�iK��Ս�Ms��?a�b0�?�I>�-���"t$�P�&U "��a�ň�6�
�J��n�͟<��ǟP��2��D�<����z���sÔ�T�`y۰F,H4��F۔UxR�|B�	�O.�q��Ƴ rl��ȂI��oNݦ����L�	K��A�'�r�'��O�����?��X%#M%k�N���i?�'�T�-�i�O���OFm&�ͱ[��QAf��g�8�d)�릱�ɍ"Ɏ���O���?qH>�1F�6]�V�8\4`C��~��'���|��'�b�'��6#1 ��@ԣ�� z@�&�|��#©����<�����?��L��u���Ɂ3"̄R0�h�dǞ���?��?I(OʅX����|
!�R�UJ`h!"\]��$�̦M�'`��|B�'aRA3k=���?��2���n���p��?:���ៜ��̟ԕ'F.q�Sc>�O�p�L`��*�J�k#��=o�8.��'$�	ӟ��Ig�%��e�iX"ؑ�%X�I��aa`��/V�V�'�"Y�pj	���'�?����m@�
���q�R�OJ��xp(�զ	�'��'��y	��'���ԟ,�s��i���$9\`(���"Fu>0mJҦa�'+zmk�cӶ$�OX��O8>�k���!m�Qʘ�)3(�4*�l���h�	2:g�������'�*��Fk�qdH�#'п3�AkG�Ǖ�M���F)*���'�2�'�ċ<�4����ŤU.=����H:�l{#��]�f����L�	֟����?A���].7)���ʇb�&8�C��g��n��\��ş �������|
���?QU*�/>�.�����.x�j��2k��'�2�'kJ��o�~��?��?�#L�.�΄0%��L���w�בE����'&��{>�4���d�O��.�"i��l��VY�d������2�ipRgA�T�RS��SП<�'\��H�74�����$Y�SeD�g�$qSS��'��O��D�OV8؆�޹����@��l������L�`����O|ʓ�?�nF����J%,dj�ZB�;x_ ���� 	�M{��?i��'�� �ۊ�x�4MN��1�ݢ'��u��Һ:��5&���	jy�'� ,�]>������ͨ�+9g��Q���m�֨1�4��'k2�'��i�n����w��Ԑ�c@$V{�R��șZ%oZɟ���By�D^/^�l������klW�rc��(C�5$¦����F^���I��̰p(E�8�O����5�i�a�D��5mF��)"�E
J�7�<!t��/��/�~����ƒ��a3�X"v�a��+�QkB ���j�DʓOЖ�+�
U�O���M�e�C�T�lQPvjI�z��a��������P��<�	��,�	�?�����C���ɪ�K	F�u� ��2���'��������ON��$��$[�U��'��ِ��I������� "H��L<ͧ�?1꧀ ��� �&����2		
���R�i��T���랞��9O����Of�$X�A0�A�0a�t�`e�Je��l��L"�­���|����ӺC3��/c`ЪA  [,R�"D�L}2��1"P���I���@yb�ΙH]@=�����#R��1IT3w�ЀTk4�D�On��6�d�<�*��g�-r��׍t�is���%��A������O ��OH�7��)59��% C�׏J� !�Mě��;����OH�D,���<����?YB/���t�Ɇ(��,Q�a�5	�' �Y�@�ɚ2F��Oq�!Z65S�eyDA�=�H!�򈂫Qi�7M"�	ڟL��#e��t�r�5�_�3uV�C�JQe�Ё��ǫ#�V�']�\���
�#�ħ�?1��S���7jԭ*p�T�o4l�K�cw�Iiy�͋�+���П��!�������[������i��([3�TH�4ao��ɟ��S?��d��r<j���IH��`���蔛!Q�F^���e�ϟ��J|�I~n��`9��I�[�����ҀXK~6�2��uo����ҟ�����|�����@�bhG�d�2�)a+N���i�z��'�BR�($?��ٟ�P��U�G�A`W�]X���Ug�+�M���?�a�ͱ�W�@�'�R�OTX9 �1;��E�g(E�7�e�5�i�',)������Oz���O @�'� 44P@�cUB�$�P٦��:vLq�O˓�?*O���"͂�@nN����k�P�
�S�T�,4�{���	����	˟���iyŁMLj����.�vi��H�`��D˦>Y-O���<Q��?���<P*|[��_�1Д����K>2�r��<��?)��?�����y��Ḩ6���`)�!Y�E*�S>:��mZwyB�'��	����I�l!G�w�֘�\��'j��XG>|1�Ȑ�2n�6��O
�D�O���<a��\�W��ٟ��

ZZ(�Nd<Ti����B6m�O�˓�?���?Y���<�.OJ�x j�O_�1ы�L� �4n�Ŧ����t�'�d��$�~����?���YZ�BL�M�{6iEl~	h�R�l���,�I�N����0�'�i�&���2��L�1�d`��ʏ 8��T�(C/C��M���?9����U���Pұ���Q�xR��Y�J��g�z7-�O���_��D7�$*q�z�s��i�)z��H�-:�7-O&bum�џ��Ο$�?��d�<A�k�Imf)�� X=�f�`#P\I��\��y�'m��'���DU�Cl+�I� �� V�v���b�J�D�O
�DǇa�Q�'���֟h�|� �G���mn � �@�wB֜l�ٟ�'
k���)�OF���O� [���?$�����ab 5�`�æ���

���O���?�-O�����	@g�@�[��@�T�ܹ+��`�P�hY7�z�P�'�2�'�RU������}y�h�S&Qz\�EN�-|4�yïO�ʓ�?i.O����O��$�'>�"�p��%u)Ƽ$�٦s��;:O��?1��?9(O���0��|��X�J��A���g����b����=�'E"_�8�	���'�~扱Pl��ӃD	Y,��s���K�pX�4�?���?Y���%i���O
�..WO��HG�Q^��\ٳjq}�6��O���?����?�BH�<q-��� ��.#�=�� J0lv�z��˅�M���?!+O|���O�W���'���O�����~l�i[&d�n�\X���>i���?Q��
F�=ϓ��9O$�4-��1x1J��T�� J�Mט.�7-�<��O����'�"�'��N�>��v2qP&�4g�Y)$� 5h�5o�P�I�d��I��h��ퟤ�}��F٤NX¤� F�WtX��K򦍹5(�M���?����V��'�&�Q�֎ )��+G�ѿxK��u�<�q5O��D�<1����'}n-8�l�f^� ��a̠��w�����O��d N�R��'^�����?�@�����%��)D	R�A�0=nZi��5���)��?9��P�f=��(�3�>�i��+2
����i�b�Y�;u������O���?�1>�~��N�G
��@䋽Ф��'�Y�'[2�'�'��U������2�Bde�mQyR͕Wv���O���?)O����On���!a��ы�#�fM�`b�j�2h�9O0���O"�D�O.�$�<��FE�x�	�1	ATE���,��e(��U�J���Q����My��'}��'�b�����)�҃�g��p�"-�u��`Z@�i\R�'oB�'
�ɑZB�􊮟���LU+����K|:�ʁ����,��t�i�BX���I����;��IJ�����4��o�+���i��7�V�'�S���Å��)�O0���ޑs���ZV`*�
�w�Ir�h}��'���'�L�ћ'"2�'H۟$����q
h�2�]6#u�TK%�iy�ɿk�U�۴�?���?y��6u�i�Qɡ�Ηa* �@a�m���d q����O��8p8O �O.�>S$�ˆ#y���Sb�d������m�6�)wD���䟨���?I9�O6�\X���f�G.�d�#�<p.�!�iA�aȘ'}�W���j��Vlm9����s�"=z��؎L��i��'No�)������Ol�I�@�bAY� \�4L`!���վ'@�6��Oʓ�.X�S�T�'��'�b�ÎޟR� 8���3@/*A�V)d����]{g°�'����ȕ'�Zc�c�K��mW�4�D}�O<~�$�O����O���O�˓{W����g�K�@!�cA7e?*0bD!��Fy�	{y��'��I��,�	��H:� �e㥌^	/d(;pb<��"w�C�<)(OH�d�O����<i��D+d�I$#H���+�V��)�BH�YX�&R�0��]y2�'=��'Ef�'+F �֥̀$��0i��X��(jת�>���?A����L'>q)�k�D��ݣ`聇hB�� �J��M�����?���1�������I�R���a�D�&O��![��A�L6��O"�D�<�)2I�O2�O��tr3B42;l��`��@Z�����#���O����P.��'��?M(K_%L��6��,`�hŰ6�`�b�k��{q�i
�'�?1��k��	'l����Hs�=�妈	M��7��O���8����}:�gK��f�@D��({��x�����W��<�M��?	��Z�xB�'_�թtF�=���!�L'vK8�-~ӌ����O��O��?Q�I	aLn-��+��EH�(�UJ	���X��4�?����?!�7t�O
�䯟����J�>�A���PN��P qӲ�OFl�ց@b�㟬��ןx���
C�D�P�ֲpQ.0�"�K��Mc����Ԛ!�x��'L"�|Zc�j�ē E<���(q.��O�Y�g��O"��?����?�,O�1if��<�T�'i܎;����ШP<L�h��>!�����?)��#�1)�.S�> ��)��۟tzj$�᫩��'���'��W�D�ɷ�����=0��Rao�&�4hY�$�����?YJ>����?�GM��?�'�1����!�^�fˌN��	���ҟp�'�x�3o?�IL�q�$`U Ȥqļ�����;mX5l�ܟD%����ܟܚCu�|�O�$�`�W����{h�}��j��MS���?Q+ODk��_Q��֟d��#IZ���,Ќ3��$ `���\��H<A���?y���<�I>q�Oe��cn��G���
R�4/��K۴��:|�ڨmڵ��I�O���RZ~b�3�0:��
7��x�r-���Ms��?���P��?�K>Q��t�V���u�V��73/��0��
�Ms� 99Л��'7��'^��h:�$�O~P�n�41�0lcHI0G�M�`dԦ��uaUƟ,%���*�� �F�ڰ/��@Z�d�PZ��铳i��'�Ǖ�0�tO�	&}�N�=y� �� ��&t��"H���Ms/Oz��_�i��E$>%�����=y
������G������"CĤ@��4�?�G�63������7f�<Q����(�v|���D�?���"a������?����?��?A*O��kΗ�2t�҅� k��ɸ�` �<��$�'W�؟T�'V��'cBg��+��Ʀ\�,��)I�K�4�Nr�'i��'�"�'�V�� ����.'�peYf���͡�M�-OX��<���?i���'�^�T�W�o@��{@* �*3~h)�O���O|�d�O����[���$�O���H�p�QS�K�[&��V�<)l�n����&�������s�j;m)�O|��dր@�����X:~A12�i�b�'��	�n�
]@J|���z�d�(ɖ,
pf�:*�T���}��d�F>)�s�h����9��BC�Ҿr��$K�i�2�'� ��G�'A�[�$��yyZc*�:,��z�株¤w�nA{�4�?y�(d�,a R�S�MKt��0*Ķ�LD��آP�f�WB�>ߴ�J-��Cbh����K�?�>9� JF4I��Q� �}�S��l�<9#�\����o���z�ʦ�:����~�����/B�z�2�r�Y��qHl���
$
'�.3�XVBH Env��6�O�UYFQ) b��S1�T�$�ԏbG�Ju�IAᚐIԤ�u�R�sa�L�4�S�yy��O/y��|����6IP%)סS�t'�Q�S��H�vm���?����?����&�d�O��S)EP �uZ�IEL1���^">��tP$&�;n�~���`X�i62������O|͚uѩ���	!�`�idK�({L� D��'5�r(�r���qѴ)��w�}b0�ʛ��'��}�@��(�(D�AƘ�}<$��@��?��hO⟘��^�P.󶣀97�@�Y�J)D�L�M]>B��y���:��&:�ɹ��d�<a�OX�q{�I���&Ez,���'��A��'�0D�b���O(Õ�Or�$j>m�B��*k�ٱ6��(r�~To;.�pf ;A��˳�Q�n�N��ē�;��Ѳ��Êb x�s&hgӲ�R7��(9r:Hcr�æZ��0��'�������?�/O�E����0+������/&��R��%|Of����{��L
�G"���Q�O�Algx�`�66�����~����fyl�9WB���?�/��0a&a�eX�ư��0�T[�?< d��O���3}:f�`�ǐv4��! �d�ʧ���G]@dS��١	@N5a��� 7T�b|^0k3b͵bL �.U�O��0v��n�* Pq-����n�j�D� �rh�E��OZ��B&]2gV�
JK�'���tO"�	��F�Oi��#�N>S%�!��'�L"=��	:8��I��;RhA���yqݴ�?9��?�e*�"}*r���?����?���(����� u	�����'z}�T#VE�$,T�3E�8۔`�.Uu*b>�O��K���W�h�P���:r��*Ԧ4��X�J�ן �`�@+�q��'.�@*���\$��� gςR}��b��'��	���4���=�m�'^
�Re�ھ5:6����T�<� ���6���>���o�1��MӐ��؏��?��'v�a�Ɋ�O�09#��J�;�D�ؐo�j<�U���'vb�'���z�e��ٟ�Χ%�B1��ɺ?��VM]���b`�B)6��ʐM�P�����4t�g�J��$��EǁA@������&d��K0��!�&���`�"��aI�.!��}y�DX֟@��S�'L�O�@�m�u~I���^8C��3�"Ob�ȗg�3+�<��S��t��pT�Di}�Z���'限�M;���?0i��,�N���A�q���F��?I��z���?��,���3��A~�'x��Q*�3Rs�Ur��5�� 
ǓH��y�t�I /��"I�����]%z���a'�c���%+&O����'<�7M馑��X�2�����<6� ��b�.$ i�'"��%�ʡ��B�T���0 ɸ����hO1��Pl�=���2Hܷ!*�� ��#zd���ɔ'�Ը#�a�4���O��';�ɚ��	(�{�.ܐ��@R�C6��H%�?y���0�C�����򙟼��-w��I3�Dώ��E��f>}Rfă�O�I�t!�%Pb �I��2/��A���>��BC�`��� ��A�'2�4��V�=|��Aŏ�'�\M�<q����<9DO�#�@�w�
�$O���+�A����"~,��"�BH��kB��9n��	Zx�H���95��Iӄ��8S����?D��U�ŴC{f�H"�x0ԭ�*:D��!BD�*=(��B��h��+D�8�DO�$� ,R�!4Y���@�*D�P�G+k��`9��Ҳr�8�U(,D�X�A�3�&���^;h\� �5�(D�$+S+�B	�5��2� �	��B��	E����Ԗ_;z��c% �l�B�I4V��`��I	��I6�X>B�C�ɤ5�����[g�2t�BGU%m�B䉇#�`�b#!�
Ai���a��6C�	�$��qbbC��A}� ⤂��a�,C�ɸ*}�I�G'G��� ��ۅ-�B�	�lh�95���q(����� H��B����!֏ӿy����ޛkM�B�	M��r��;`��R�k]���B�	�t�8��L+9Z�J���
76C��T��2��̀f�LY '��:�C䉮!X��1J�v���i�5��B䉅��M�f�$^�s��k�C�ɀx���ps'�	^�4�Q���~�^C�ɍB�eR�I�>�*�)���hC�I
"���Y�c��A�ۦ`rC�A3ppц���)7�� �K܏J� B�"2:8���C�:+!�	���#t$.B�;�^�pgG�(G�}1$�B�n|�C�I�k�$�Č�>����G�-'�B�Ʉ=�j��p`�D���6�ܭE���$'&��8scA$}��ͩ��	I�:i���s�邆퉓5l��`��h����ė+d���Ia�G4N6Г�Թg�1Oҗ�ę'o|�@2#I�T�|E�`[����t�z��G���)�h��6��6˸C�I�|�N�X'G	XU��z$���uY���s�ԬU�r��Q�Y���S��"�m{�)RF刺^3�M:6�Œ5B*�*��;D��7�G�s��j�&S:+kF=���<���i�����k1����GyRL��9�b��5 	�j��qQjS��0=��Y$u{ƹ*��W�",̓eT�NDF @���;k����v@t�@l�A�M���'h}�{�S����k:�(���V��A�P���'���E�@�D�
ٳ��ӭra�jI>���$���{�NL� �jM��㞌t0��K&"�Z�S��y�F��$����6s��6�^59�d0ȴCH��a13�@���S�i��*��V��#)ʝW���R#��y�dR��{	����M@R��kB�s���Gxb�>8�"Y[G��Z$>�;֌�	���?%qS�W�'D��"rJ[��P���3b@f;������b�Is5�M(����,۔:�ay�bػv�PE9A�I�i�z�B�I�+����78>�[��E\JTb��Y��U=�T��&�O�����|�&S�sAJH'h�}�WK�8kx�'��|�SC�+�Hl0�@W$��s�{
� P("-���RN-��Q CF�1 b ��'Jh�ZH>���H���'�5�c�TY�J��*׳o=��y6J#|&H�A��p.r<��I0zm��N,<�b�1��[*.� �Ob�3��+<Oz�   ]�Rq�歖��@qC��*LO^	�RC�,- � Avm!@hr�(�Z":C�`����'C,Z���'äa�����Z�	�$W�/�Z��:h����fLW�~�,ڢ�DG�>,ئJL�%J적��8.F1O�y�Í(DS�,���7Nz)�И|���z(�Ԁϱ�܉@0�ߢ�'v�h5��>�~��򃆢RɎ�bi׬��ad��i�h)(��''���à�>TH>�����
J���u*�>~�*�A���o�
���I�@.���JF@����d��m�"��S����a��.��$�77s�`
w��-����i��!7-
�{� \xf̓Dy�'G�<` �/�8L��y�/W�|� �'�@�=J��.\ꄁ�D�Q��6�*��ٰ�O
 �d�#.8p�F%)Z���&CV�����c¯�Jwx,I�E�� д\'�,K�MѢ@P�]ADf|��p�7�I%[�0�z4��B�ze3���c�u����1*P�G#j�1;2�Zf0�D{rb�=�\���j�I��@!��ϛ6��\��E�J+�a���9lO�X����=T�Nx2�N_��p�pΚ�:��A�'o��#�7Ng�^�x0�F_��P���K���+ ��T��@�P�{���W���As�[�,V�u����_>���d�ٍ?��Y�]z��'�����*��u��×?s�4���?��FcI�S�D@�#
�5S�YrS`�of|�D|�kڹHhzE��n�
�0�Ŝ�?� ��yn��إƁ�U��k��D�R���g"����Y�D�IZwx�
ao'�)��m�� CY���E�Jh�x�F��ȶǟ'm,Q@Wϓ��6�`�O;|yӤź>���9~H]����p����oS�Lx��7֐�ȁ�'�:�#�e�-��h�cj@�"��\3�}��P^L��ض��%�� M����>�u9�(�o����fԪG�Rv"O,R`�ə5�T�D&�W��X����e6�[�E��	������H��Ʌ2����S	� ����b6�B��\�Eb���>�4)��G 7��(�������%"Bpϓ�X��4b�X;�eH�&�/)���퉗L�Х򣩈�$w��(�hLy0ac6�X�$pA��7Q��D���8+'��!`���ñ+�#:��Op����=PJ!�礌���O!�3��Zo�8�&��\�`A�'�@�ᖓE.Z��dˡYWz�bȎ)T�~b�U?��9�g?鴃��=��l���B�#�(�:�́p�<�'
�Ҏdjӊʽ|h"�2 ��a��Kʱ��p�U�]��yB��!acDM�f!�!����۔ϰ=��*T�Cq�Q�t�#����� "���J(s��t	�'34��a��W�L������0��5;���!F60��3Ñy�|Qz�ǜZ�'�)��ŀr��+ �O��4�ȓU�t�I��ҨF) 0�4�T� �SD^�P��)�)�Z�"�ڨQ�d�	�ӪB!0�L>�a��*!�$�R.M�'B�r��e��xi�֊�N�Kq�lF�ɀ�)M�R�p���-r�qZ/мL�Ι�#M97�h��'KWx���B�1o�~�@d��:x�vn#�	�2X��n/Y)�9���)����g���N1.�ipŦ]� �*99��Q�{.B�>#�:50p͚�Z�m��
����sүR߼���I�&- Q)��Kuq�(p�>﮵� ��� ��B�It�&"O�1��ЇS�V8!�ڛ|4�Qd�*g �\{!d�1&���IS-Q���q �хW�F�>iqi�6EF������E��j@o��D��	T@��t��V�OӤPF��}YV�����-8l�
e�!%��ӓiU����҆�'Zt|�vH�������XEP�yB��He%Eƕo�da	 L�^.xc�M$�t}�fN#h���j$[5�JU�w�� �y�d	��|�)���Ut^��(��¨�8[r�L�Cd��|�&�ͳej��~*�ET�����1�(Y���޾���r" �\�<I�� E�|�RD�Q�R.�	2v�ӷPB�)��VTke�#7<|	!�"A�l���0�	�!���f��0B��ʃ)��T���%�PŁoP"h�HU�I4U �	�S�תH����.,r�EQ���x�z�����!�p=���	��h"�`D�m+A�dL�Mk� �9v��"dl��f�x�B̖r����n��� o-�N@�'� cb� T�<ѵ�3U�FږT/:*�BU��Y�`�dŃ)aP���)5X=��t�'P�Hͻ{�~1�T ބk�dh#�J�xn�|�ȓe��Dc�摍<��5���wW�H��^�M�u�:<���9I�h��FF��O���E#�"+�~]q�a���7�'���@���8���� U^p`��3B��ul�@GJH�o�H�RF�9��و��+�0>�gˆ#hl�C���+?��s��K_�7��1�Z=%��Mz�Wd�*��-�?�R7�� ���b��YK4;��A��ΐ� "O� ���/�dm�`k�Xm�ӈ"&��8�&AǔI>�i��дx�!`V�i�
�]�_n���.ٮ-���c
�|��C�	;&馄�ƅ(r�,�`րh�7-ʹ0�عA抣%��e1O��W\�]✵P�g��� d*�'J��T� �%b�)�����C��-ܔ�e�%v.\!)�
ODu�Q�߯E��]h7E�p����$�b��эW)??�hs�������߷H�5��,֙�Py�Z�1с�w�@;��߼Kܠ���1]�@}�'s."}�'��r��cR�c�h\�UҼ��	�'��2  <R��`"EI�Q�HX�C0 �!�@T]��	�
P�� �:S� ��7�$o�1��w��Psf s��B��!����S�u��\�H3�������� ��Q4�t	C��}�:��I-���'{�t0A�R��d�G����#V
� ֩[05�L��,��=s �f��́c�@���. ��8�өǾ��:rlh� L�"~Γ
��Y�m\��$ k�'p��1�?���Z{���Ӝeoz��e���j �L?0��m��!S�`؞dr+ޔ5Ʃ��ӣz���U�I$%���~�$�_�*�2�O�`���J�q�2ՙ2A�P�!�.x�T�k�Y�b��f��g�K�3��'�p��!�\�OA���Hן}�(�I3�<B26$�
�=�1�'�N�Z���^e�� �H1@þ-:�O��(�6�)�'[��̂���$�6��3�R9zX�ȓ�Y w�Ӛ1�d- �J=9�b�����X��)|	�E�T!�o�b$��y3��!$@�k+�̈fKЩA���ȓ	�ࠇ����\�G憼��B�$�"��Y��1�3�^��6��;��I�5���?�L�AM�8T+���ȓWd)fE�9�E!W���a�ȓ2v4�@�
,w@\�I��Cj�ȓ3ID�A��-t��b�ߗv��Ʌ�*���r��W�B!C��^���%� YÇ>\O�]��	(�D�r��hR���'��}[u��*��Â�]5�J�Ç�b�!�D�(_��Pl��!�ʢC�7"�џ0H�#As�OJƉ�#�]޴HZ�APK�	��'�,�b��Il�a2"��E�2�Y,O6���)�)�'=��E���8�ـ��C@3�X��z�~�smAt�����Tigl�%���5�U]���ŉ[�Tƒ,I�i�MҴ��gH,�O��PE��.&Y��z���6� u�V���54�B�	�78`�:3��\5�1�"
�>uwvB�	<?�:�8��Ľ2��V͂�%LB�ɡ����1J�Ғ�1Zm
C�	#e!\%32K�*
��
����1!�B��>~��Q��B��ے��� ��B�ɴB^�xBbw\6Ƞfl��oN�B�|�e��R�%J�鑢�L�h��B��G MB�K�7T�ųt�ʸ%q�C�>�q��G.戱�r��&N
B�N����'�/ ���Nנ)��C�	!dK���V� �~��iħ�3YbB�	<<�a֏Z&c0�3��K���B�I�_ZX�I���H:�E�g`�;U�xB�I%~���Ұ��V }�����Y�bB��.B�0A �Ћl���IU��2��B���(Kq+�s*8�q1�	pD�B�I�=�2lKI��� $kMh��B�	�m�Lа��9d�r��I�.��B�	_L2=x`ː�bTk��2�B��/:B�+�ň�Y�ɉ#�L6^�B�ISul�ST�ڟ7j���6(�;�C�)� 6���*�ثS�Q�6�h�"O��3䙡Dv�h ��� ���"O.}�*�<Y �٣���C���bS"O���V S�PdA3b��\��I4"Oz����mV��+чD�S<S"OJ����1��!� ��}8<D�"Of�	�
	`���)ˎv�Q�"O�]iVAżz�\�S(E~�l��"O#�Ԅw?��z7'�;�ظ�$"Ol-�v	��6���{߰���"O\��F��uY$D�W%*4�]Г"O0�sbk�7V�ݩ�
�P*���"O$ٳ��S�s�Bi�sG�!&|B�"O����"�8���CӅ�6�xL02"O.����
�K(��pb�
�:�;�"Ot\���:Ws�}�Ύ&1��HPA"O�	�d�� xa�\�ez�]��"O��R�FV)�Y��X���@�s"OP���P;��TP��Y�[$ �)`"OĒI��m@�Ȅa@�r�uj�"O\p"i�����CK9VHP�S"OBd���..�в2��j�`H"�"O��1�� #�@�C��<�v�R�"O����:[3\��#�66_��!�"O��P���(Jv�Z�Ē�"Z�|�p"OЀ��Á�-�Z�9���=�����v�<bh�3h ��ëhC�T2���yB�.U��HY��^d1	wč�y��Y�o�Fu�)�(j�x��v�� �y�'�u�������p�tq� 	�yb'\�U@T��F�<�Z�h���9�y��d�l��K*g���AɌ�y��(�޹�ֆ�����x�'߃�yRf���p��=b��<9%\��y��?�����a>����*�y���7�i# V=(����$a[�yR
T$��p����kA �[E��y��'T�p�z�J9dh%���S��y"�~���[�!d�j�2�iD(�y"ā7�=�t��hzI֣��yrώ7C���M %d�j-�� �y���) "�Ez$��2[��ps7���yb�Q si��OY�i���9&�ވ�y��	���� &!�X��ʌ%E�lC䉔/�:��f�@�ee�8�MЇk� B�	�T���P"/�V���G�S�-�2C�I��<��N/V�dX�4��U�B�	�h���y���"�-Թm$�B�I��(�3ތ(1^�Hc@1iӮB� [12	a�M�oL �2��3hl�B�I�B�p�#�8W�d(�g�TւB��������	3e=03���\B�ɲA���#�"S/I�����_�^�*B�	��� ń�kɞq����]��C䉅6_�����9"b;���B�IW�t��"N�#3< bQ�֘B��C�	b4:� .��3JT=L��C�	\��)z���#���[�.�I��C�;z!��B�Q6ID�̪��$_R�%D� 8E�U�@%�"�V��"�<D�����x�Đr�E�a�L��#�?D��a0�M�Y�����R�k��yC"�<D��I���*M�0 �!Z��m6�9D�T@d�rh�+�Ϝ(] �	qԅ8D�� ��5�>��Zd�V�& �V"OfmY@ON�>n^��wLX��x"O�T����Le1�����*t"O�����U�_╰f��=R�V��"O�\Z��n)�q2E�.q���"Ox�z���o�h�(��ط,lN4 G"O$�r%M�\>"d1��Ye8�"OT�R.�lG��zB��} �M�b"O�a[
z��`q�ϙAz-+"Oy&��@��k�SN���"OD��g9�<�R����z�:f"Ol9��
9L�^��G]?c��4"OrHx�G̘>�D���h��u�"O\�+E��83���TG�t���b"O�x03�@'N����'��>����"O
�W.<h\!�7f�!R����"O��ub�'�HիF��/o;�D*"O�� !���E�	��W!P�ɶ"O�8�u!Ϗ5Ѵ�;�[�:r�z�"Oe��!�:!7pLK0��+����"O0D4��+ш��	1c�n%:�"O0 �,�>��	ʔ�>|��t`�"O��8�ME3T	$���.S|4"O>Ũ�NAB���s�X2*����B"O,�CpO��t^�y�R��qx�(�"O^=�'��}�ʔ*��@�c��ps"O�鋃+>'Ԡl�r�E���H0"OV�	���6>ɤ8p,ڋ߂����A�O��d!b��iWNܫ"KC�n���i�'�F��b! �4���@���:9���1�' ͠�AN,ir^5�4׉�:]b�'�d��ǦY�m�l �t����Ƒ��'3�����ǒCoĚ7lL�\P���'��Pce��&�
�1�CG��3�'}4� I	�r.��dW�䲝��'"(U���;Ţ(�F�/[&���'�%�pn�`�:�*��(N�
Mi�'�\MA�	J!��;��7����'��!�Ǯ�h�����'�4O��
�')��Pc(9��\K��Ga�<��'�j!��O��D�(āf ]�ȓ`[>�3�)�*�(���4r����)� ,�$�ʒc�IB��T`*��ȓh����/q�N��!̑�aHe�ȓN��z�O��,��m�#��A�ȓfS���DY�}������ 3�� �ȓno~��6t��śC抙\�4\��3�!`�����&�{�#�W�z�ȓ{�\��P�(H�u�ei�.\��ȓjcz(�BM��M1���c�hL����(��e��0�d΅ �N)�ȓe�� ��̤{z�5�P�Z=�숇�	�С�9[R��z��]�WH���ȓ\���!�( �7�в䢂�6نȓbH[֧����!�.j&�����E�T
L9P�{���;� �"O.��P�%Z���S�g�J�n��0�'1O�-�PBR	}�|�'Q�5��e"O�4 t�K������I��!H'"O��[!�ي;���U�_^�ѡ"Ohi�@�j-��+d���Y�"OH� 7�C�,��� `��H�:$�W"O����w�8	��>hqb���"O��8���m��h`ʗ�VQ��+�"O� VJvŵNh\;3*ĒLP u�p�OL�=E�tG>�L�r᫉�Q$La����yR�*s�}��ƫR��l�dC��y�CȄ4�,�r�"�,D� 0i#�X��yrm�90$ ����Bĕ�"�Q��ybcT�d$�`3��F8"�PG�Q2�y���(#�����A<�'kB)�y2aՎVMF5���GO]h 𱇄��yƎL�D��#ջHҁp�7�y��S��:������%Q�3�yҧ�L!L!��ۇ]�����Z,�yrJ8� �ȖS�>����O�y���u9���C Ɓa���ٖ� �y�(�;H�`���$� �&�
$�y%4O-��o��0���G+�y�Ǟ3,E0��Em&8j�Ö/�yR� �1��I�5k�3Κ� ��ɪ�y��BL���@@��%���+G��y�Kfv4q�gְ+�v�2v.�*�y2���M3��$$*Dc��� �y�dėXv���,��p��'�ل�y�.��I��LI�lN� �����y��'"2([	�PI�����y�*ױw	���D�(G��`�@ǆ�y���,����^/�\�yՆ:�y2��5����#[#R*լ�y��� �h������h�N���y�#	�*7֙)���0�D�.�y����-�2xK���
�|��G��y� ��y�&%��FA8���G�S��y�J��P4p H3�ܫ%)�U;6d��y�T>Nyx�cp��6iQ��i�p<��z��]�A��;C �U��M�!�$��v����������sP�C	a�!�$����+��Ǫ5��@rP�os!��]�'��aF�3�R�Bm�<KV!�����;�ɍ>o��I��+B�!�d�������%�v�TL'HC�H�!���YUʽ	A� ֶ�A�&�!�D�40bL� Ǖ qŮ���A�*_!���L@��x��ȅn��,�E��#Q\ax��k��+�KڪH�����A��qH�B�	�gg�hwLNk��|떆B&.�^B�I<q��걍�'}�x�D�@�Q 0B�ɗ/�-�b�f�hdQ2�;@�.B䉀'(]�GG�,�qc�H�B�	,xP��HI%P�@�?o0�B�	��,aq�J�sB&�����M8RB䉘n�� P�H@Fg�ЧR�-XPB�	��� R�	q���F'N> 5"B䉎 ]�D���5m�}�\��Y+D���ҧ�"�ʰ�v 
<�$�c�-D��ZuNj�5���!�6�Q1
-D�T��T;oX��"�Y�
}3-,D��!@N�j�Y���>%V�|Z
=D�,�$d��I��-:���"��;�<D�0�5�P�(P"�8%����qe8D���q&��O��$�	iɪM��� D�d�BM��F�9����z�l@ǁ�>A�z$�9c�/*@�x��ύZ��\�ȓ-�4�Q�8�F��(����z���:di)+����hM�� Ɇȓ_�V�b2�+�pK$@�_���ȓ?���gՅ!�`ɺ� C�1]T���S�? ��+�LͶ!��{7�ڿ*����"O�I#cFT�X�g)����"O� {6,ԙ�ʭ;ǌVh�ٗ"O2�jUMSQ��b�J�'>Tt��"O�Pq��ĮB�"���	�w1�p��"O����I�b���?`f�C"O5�c�<�r�� X��d� �"OT�����!7&Mi�A���-��"OF52d���:w�5�`�����""O,QQ���	 �Ύ�/��4h�"O����%��3����N�0ʀ"O�H)A��=t����,��iz�"O���`�1o�L��jH-X��L�"O��ș�/y�I��I�?��2"O�P�#D
5���m�4Aڥ9D"O^�AAGH�+:ꥋ�C`�:�"O�d1�	�`���%%U�R�Q�"O��Ѵh҇(�ț��I�
�����"Oֽ���_�Lr���+����"O ���Cʞx�l�Kچk�jl��"O�A
f|Ϙ@J��Z�"�a�"O�	��L�&��; N��q�#"Ob��H� v�m���U#S��M��"O��84�R/on��梇�t�H۴"O��v�Y>�D@�F�P�� �"OnL(Ş1꾥 w&�� �Tͪ"O0����Ĥw�TibF G�Ԉ�b"O���A$�8EF��!Ň�(�����"O��Ұ�X�IK����7��y(`"O�{�mD�'ɨ��"� y�r��B"OJ�ӂe��t[V�ʱaX�w��@"O�xT�T��f�:�Ȃs�&�Q�"O���� ~�S�+�t0��"O�����B>u=.<��k9�`��"O���e��y�J<�E���|����"O�Q�@�N�F{j��$
A���Ʌ"O�}[���
o�A�N�*fK���"O��k�JP���U��i�Q�"O��8TF�3y�a�4��Y�~��"O�x[�d_�:ڄ��$�W&~��MKp"O�1�ʉ�]���T�^$�R��T"O�]Rтʎqa0�04�@�;|��qR"O��X���=XE�]�Iz�(2"O����6�� �ƚ9r�}�"O�4Є�V���@3W�F�P���F"O|�{�i�|�ʡ�$�@4q�""O*xQPn��|��i`�.��6	�T� "O��ߦm~�c�M���X�"Ob=b�)S�l����c	�qլ�Q�"O��E�^��SB�	:G���a"O����=t0,)�U#���8E�"OX8g*�qL0ى���`Q8"Of���.�k���Jŀ�.�HD*�"O�D:��=�ұ*��+L��"O"	�7�_�M{2���l�E4�-��"O��u&\� J,�ABm;�8JR"O�m�*ЁY�T9А��;:xB"O.�k!C;:�s�bY����"O�}��-��c����_��RL�&"O���7ˏ1}Z��ֆѶA�^d�"Ot���o�?o"9��Y�&�De��"Opt��֠�2�SBK���"O��J���<�~���|ޠ�(G"O�9[�$�"�`1��(�;�b�3b"O� ����N��[��a�1��1�"O2���g�2 '��Zbƙ�"�2`��"O8uk�C�tO\�S�C_���Hq"O��"�ӿcKj �'ň�Z}��R�"OFy��蒠�\{a�C�2�l,0d"O�Ej�#_	%��}�t�_�rޒ��#"O�T��]<*�"��#��0�"O����U�s֎}�oO��*�~�<q�V�F��4�e,��8��q@�<��Q�
�xkd���'�je�z�<���ޘrfv��P/L)�H�!co�<�Q��������o��S�b�g�<�����Uӥ�E�f*�3��O�<9��  � #��2W⡹֬�O�<Aԫ��n���'Õ����t:!�$�\�"�қ\,u�УO8E'!��)h���w0h±q㖿!�@��@z��,S$���[[V!��=w/�,� �N�D?�!���ѤwA!�DJ�Q�Ș
a�V	�J �fa�w-!��14@6�SMX�rGT���[�-!�����p��['([ d�A�O!�D�/&=z�@�->H�8ŏ� yy!���(X�I2�G (('V�Q ٓ{o!���H�x��-5��!�GA�3pi!���V�a����W澠ɕ�	�zR!��K
�-��I��x��I�B���!�T<2x*b�W�Y�f<H�%�4�!�䟎QV�B$gA��$���S�!�
!ȪA�A�?n��t�QhƘ/�!��TG�B��*n�0U9�e��7�!�䘷k���Raˏ��b�83n��U�!�d7n;,�*�쒰<���c���!/�!�$�Q�0�rƘ�v@�K��Xj!�d�+}�t�� ��@�i�*͍@�!�������ⓡ��D�2��9�!��?$�P�#B�����D�F!d�!�D9%�8���������Ș	�!�d��w
� e�D�>�D�p���(;2!��]�P	s���K�"�E��*�!򄀽n2����"Z�7@N��$��	 �!��πZ~�Qq�"����!�t!�ą2	�n�zɍ��,�� ��U!��$��5�o�=�4�e
�oP!��B]
�Irk� 	���(ؔ!�D)zyx��C�N�h��	�!�D�1,����vcW�ƒ�Ǡ\�`�!�$�#cS�|�� ��o�Z�!��O�;�<�PaĂ_N�y�h_��!�8AoV����K>M>iF���nu!��D�65�="�O T?�<�䪄D�!��9�� �e�TK X�a6@��!�֦s�|�	6���Zz�!%F\X�!���J�=r`CT "��7e��/�!��өMbr���V��G" ��!��Q[:��0e	�:8�p�꠪X�}�!�dC�"e��͇l�h�Z�j�-*�!�dոq��%�����y� 4�#I��w!���;}@v����%R���J��@Qd!�DU�X. ��5N̳ �R�3QL�6H3!�D��0o�@)���/a���3lT�L	!�������E�\����R_�	�!�D�0=8꽫�&�ܥ���D��!�$�i|� �F��?`��ł,�!�� P쒕iW���\rqm�6;V��"ODܐ�@�)}
�H��.=$zq)6"O� �-8/���YbL�1UB�ib�"OA�4�W"�~��"�L�8���w"Op$�pg�2[� \K��ǌ��4(d"O���T��s��)�)�%4�\�t"O�-E/Κ^�2��Qi��G���7"OH�z���o���KiP�{b5�"O��R�
Qf�*�r��Bi:a��"On Uk$9�>�0���vfɨ�"O6����E}8���i�`j�"O�� .IyX��bK�m�&��"OMZ�N�'[��uAS�Dl���"Ol�˫� �Z⃣N�h��E"O��b�h�`*U+�E��}z�"O�m�"D��S$�d)�v�`�F"O6�;� E�a�L��ݸtl"=rr"O �xC�N����E�rl�Q��"O��[�W/5,���
��'I< �3"O^LشA109��U@Z��`|Cq"O��`2�˴=Xpgώ�Q2����"Ob�a��0M&x(;5n��dKf<��"O�Y����:^t�R�N><�T�B"O����^0�`�җJ�%;�+"O,I(��q�Ve�@LU!Gb���"O�����n-|�8��	���q�"OLp��e�*�Z�I�0n�R�'"O6��Q�)�2R�Y!�H"O*�
�%H%P9j����go:؋&"O��X�&��d�rPB��ufP5�T"O���A�f���u�OxF�X�"OP����Z��+� \�4d�-P�"O�����V $m� �?3XX��"O��!%�:�f,� :QC��%"O ���aߨR�\��m(d0�B�"O�����[�
U�@�˪$�$ %"O�X �XxY�EiAa�,ut���t"O�����&B��܉���+J���"O�3p��Fv�c�t���"O,D�s��P��Y�t�
e�"O �P�O1HM)e,ƴW�P��"O��rQ-ݷ/C.(�P!��Y�B��f"O2��FC_/�ҍ 0]�ZB#"Ox���Fc�^h�p�Vmʲp�*D�{�^=-�0`�g�@�E����u-D�0��bK�`NP)�nߚR�ȹ%J=D����$�y8zX����$�Af�%D�XC���%X$
@��d��g��HL!����� '5٪�g/�m;!��6#jb��J'%�N9�-�,!�$�&ߌ9(�H�#9q��웊1�!��٦by�<Y��(>�Bu��#�!���7v��$⍉1�9	W+�+V�!�DO�*�� �灊$ZI����?t�!�d�LtEc�d�'_�j��񬓬m�!�$ն
�:ڀ���<&8�+��.�!�������)R�Y�ƫR5�!����P��\L蘢�,�LG!�����m�T��"0]�)Sy�!��H(��9qkX��(J0G�!�DM'P���$+�>'`n��H��)�!�^+q��"'��9��Q0�䅍i�!��8oJ���� ,���;�fü7h!���ss&e:�K�9c{~�Гϔ\T!�� �
�"ܛ ^@H��A�v���a"O�i��ǚo��y�&&Ѫ}Q�'�B�P���n�R���Θ�^�Z��'���+���#F�1j���,�p��'Ќ�HeI�I�VbU��6`S�',8ʷ��b��5M�x~q��'/�4Qw��؁QeI��	�'�J��%]�@�R�����L��'Z�a��͉_ բra�'X<h�0�'%@�U�>��c�#÷I�J=r
�'e`m�S$P�+S��hD-��=���[
�'t4QTeŷ`�\شj@�;ߎԪ	�'5�V1es����H�7���'�eN 
];֜HF�1 uPtZ�'��5���0�d9x@���!��$�
�'�=yg��k�Xs�l���
���'����1 J.z>����ο\`P��'�hE9���ڒ��τ�pon8��'>��J� ޷fB>1�Q*�oU�p�'b���F�K �S�"G$Z$60��'���r#lY�*R0�bB�/J�v���'����I��xw.["���
�'.($SU*�Ce��#� L!���
�'�H}���͐\�TT0���7 �Tm)�'2z�c��Zْkv�ʜb�!b�'�ȥ�c�S"|�:2�*ţ
�*H�'Р��g��b�H��E]�y�~�'0L�d�"	�>��LrzZ�S�'��T��M-B�l� �άg�����'+�� �@Y/�����=k�!��'Nf�J2��s����#�?mE�1J�'����ʃ�?k��1P�T�]�ʓ!&�`r%�';�h�S4�Z��ꌅ�D�Р��M�mnHK�&?�ԄȓaU�ݚ��M	'����P!VG���:L����ʡ&�֍(�@!	����|�H]*re@4�P�A&�I``��ȓBY6��J[0�BڕT�X�ȓhM�Tk�h޹2X�K�	Z���{< \�PI�8]����an�H8��@P�=c h�8fv�|�Ɯ�0�݅ȓJ�4)��%8�t�4�$b~������h�LT9��!��O�"Ė��ȓff�(	6H�=�@hň��V ���4z��ꐁԵW�I�P�V�� ��rx.��lX�q��}#2��"=F��ȓ}r����6�`t{�k�\�l1��}��*���
&TK��Ή_����ȓV�8Qt��;Y(Dey���w���ȓ:�ꁺ`D�2td�� o�b`��ȓvd�J�KJ6�|�p��(\p����J�J��$s������Z$l:�i�ȓff�"N�6%�<գ`B$1��ԅȓg��B5�\?u?���JT�\&��G�p"��R�lF�U�A���(\���
�a� �>��d���3d��U��.Nd�#e�Q�(��8Zg`�+
�dH��Et��.[D������#	���ȓS�ZL�f�Y5�\ٱ�L��U�.���1T �l��
x<(� /=/���ȓ.R�Q��� 7.���O�,a9̆ȓVW|�$*צi�f�S暩T8���uq`�MZ#FTV�Z�N�$R�p@��Z��� @�	�"�zCdܙ ��E��S�? �0!�F;��Rh��0M�}C�"O����B���C�֭02&X "On����C��a�)�4��"O8���P��4Rч�0q[TQ�c"O��I$�����u��	�ּ["O��X��ӚV�9�N�0���"O��y�;Mt�ɒ����ʤH�"On�k0��":v�cUdR�BW�i%"O�k ��k�I�!d�9@;�tp�"O*�!��<#���<+���$"O��i$ʇ�g��V�a�8�LD��yB�ߣr^��&��+�p��l���y�D֙w2��2�A�*s��0!�>�y��޻Z�rP�� m˾�2�A��y���#����h8 lb1A�;�yBDM3W#b0��@n���SE��y�C1m�@�
���R?��*#GG��y�� G<�C"��ZD�������y"ҩ�)Fc��(������V�y�	�\+��bw�]�'�()�f��y2"��{[8D�gK�M�� �+�y"�^fO@�
3f
݅ةyC\E�
�'�	����1:TE��'5j�l��	�'<N؀T�Q8e��5� $gf�C
�'D����|D2��`)Ӫ�*,x�'7R�gFG�{�D@�n�*(�r��'b�9�ӊA*{n k'�)+{��B�'+pS��[q
��Qb��rqX�'l���
O.|]2ta�G�]�r�'�,ذl�1+�����<`&���'������ �H~�$c�IW&C�IW�`҂�*R{Ҙ{Fct�<B�I�~��L��
*�XG��C䉴>��Y��)}�Y1!����C�	�}=��1��>��l
�Ѐ{4�B�I-T�Bbu�
>L(�p��3�ZB�	x:���/V�����F@��.���D�5
�r��6b�>M�X��ST�+!��V�)�S�D9�<qɑ��1�!�$��J�(d.O\L�!� 5%�!򤒬�SK]���A .ʐXo!�D����|BF:;˸=���C�!�䊜5��x��k�
ze��P���!�=~R��ʵ�C6�W�]z�!�D<D/<��M��F!�(��[�q�!� 6Ӑm�ң�6	����eϳVv!�֔��qZ��´1�p9B��%E]!�ě�e���.I�Z��0vh��jG!��[P��Ĺ���3���S'�cK!�d S�@3��ܨ��'˒2!����ؼZ�hQ	:�Z�� �ٔs"!��x��I�D�B�+�n$BG�ǥW�!�$��W�M�s�їU J1a#J^�p�!���-�>i�Ơ0Lh�s�N�!�D)6��1)2��9 E���X!�$X,`�����H�7�8�b�F�,!���2+ud6*n�5�cͩ�!��:
Q�C5c�j�+Z�|t!�d�3s�$�R���I��Ꙥgf!�$1O�b�Bg�C�H� 	S$3!򤔣}�j-�`<p���q�K9l�!�Prp����� 0��-�I��!�_�=ӌccBF�!���r�A*?|!������.N��`$�M-ou!�� �K��	���)��ܱ+~$�"O^���ϊFĜ�����{�"O
X�`ɉ��PD��,�'�2Xr�	E>1`A��Uh�y���>�kg�'D�Ӷ��*�d�1��.(Y�Tk'#D�H��I�n�R)T�P��9��5D�D��<y�<��kή�Xn3D�����BvӬ�y����7��F�+D���O�Uv� ��B�f�-z/$D����C��Pa�3�@�V��)�0D��1��o#�(H�g $�`�
S&!D�p+4k��}s �݉xњU�d! D��I��[��p���LҢ[&�<D�D�����W�\���A�g��rc�$D�x9�Dݺ<�!�CJ(�z8+/D�,+T_�"�D�K��H�\J�M���?D�!&�D�Lm���%@�rGF�y�*<D�\����9>���[��Є4D�ph��"X�rۣI#@�����1D���N�vTE��Ά3^\���*D���s\�K.�T��h��@��6D�06/J�V� ��"���(<�s�3D��`B�3�i��F@�K3�\i�G3D�<�󈙯9��N�
+�����;D����&5 i�aV�״
�2�O��d�O���9O�c�,�V�0Yf�Q�e&�[c��)��8D���P��/�(�3'$dPu���"D�٦�-;����B�6��E��� D�X{��Dg����c�"���c�#D���d�:�-�S�R�*Wl�x��?D�|i�	�R#<ɓ�##Y�{U�>4��{d �1h������8��3�.�_y"�'�r�'��	L�'�%���[/h]���#�<fS�-C����'v�>�I0g{��X�I�m�<�M� ,C�I�|��F"y+����5_�C䉺J*$R�'�8_������ UbC�09��E+���%e��%���f<�C�
,d�f�OzǴ���&tR�B�	#$�h�l�9��2�i��gd���2LO����@�6�>�7cж}���"O&Q��(XW�sQ��/P�BP�"O�8 4�:�ȱIp��  �8�"O��rK������0���v"O�˒M!��-;q@]2���"O ������ҁ* �=�,x��"O*A���*G8�X�s!Z�4�d�)E_�ȅ�	�{���8.��L.>`���F�T�C�	D.8Jd��6o��T�QA�4B�	q x�0��_ҹ�T�#G4B� �j�Õ �)l�x�e�_$�C�I3c�4�` f�F F����l��C�ɉD�촃F/�+=_l�q��L&�C�I��l(��A� m�S�o�/W����'�S�D��ѱ'h  �,�:����e5u!�dHP��)1��n�.H������B�ɧh�)C�dd֘J��S�8C䉣�\Y�p�٧h�f�c`�O�tjC�I�q��S4%�2	�!�ś�W��B�I91H&�Qc�*����٢(�ax��o*n��2�$.�z� � �#*x�Ol�=�|��8]��E�d��P��I�7�;�0>��ET~2�W)�X�T�6dܘɐ�U�Py��I� a� �j�J<\�n�c�<!��\�d�I�啑�zq@Hc�<� L��!�ݮ`ǘ1��rʴ]��"O���� �a�̱#d�-p�~�T�	ʟDE����:P���g�:i����%��y"Ǘ�_ ����Ch6��,A��0=�uN_̓S M�mO�?����#ТF��d�ȓy�6��c�U�a��U��늺?T��ȓ(��L��ӆ3쒐1�gU9~�@M�ȓ>���1ע3XdIa�Ʈk�l}�����òGE��IyD��F�RM�?i���0|RgK�]4��r�&�Ś�*�Bx���'���9��)w�T�Q�l�M���00�ץ�O?�ɕI���dM�% �c�ІL�:B��0��Aaf
��sp��d�C��C�*'0�4��ʩ}�l0�倊WN�C䉄Q�>Ԙb'ȠH1��� nI Y��C��;4�H���;|ޮ�UeH/%�F�OR��'LO:�r�X�Ҧ(R5�S	����"OFk�''NVak��Q�Y��܊��'�O�q�!M?�Ӽ�'�,X���
>^p+�)�S�<��`��H�`'JO�E�C�Q�<�����RH8{A B�6%c�e�g�<������nq�%�ʸy��UK�(�X�<q`E٫0I��+�� �3��	Nx���p��B�V�.�%-o�l�ȓE����9��A�V��+��Dx�*I#�0|��b'}FԘ�eE��>:���a�O�<yШQ�`s�X��Mų4������XL�<	�NV�&��`���.H��@[�%�O�<�ş)J��"�P�AP��#�(Pa�<���(f�؂��T'lU���f�\y��'ؤq���A�fK�����4c�|�
ϓ�?���?1��sS&�X�B� &l(�L��`7�����?�
�#�jy8�ʇ�s���1��m�f��ȓaT����
�.�d�W�
�+�@��	�b!ؖ�CR!�',�iT�H��"�d͐4L�?���ڔk��o�Xh�ȓ2����s���ӣd�(9%����ɁC�ȕ��9�4��B���M����d�O�D�O����,2z� �AER�p�`���9$B���Ob���՘��܀��j`���r'ڸB�!���_(�����~NJ3�¯~!�ē1�>��j
�C6-Q�A�+_!�V!Xnt �W�Ə*Qس�`@�hD!�d��X��ӖM�;\�(�/�9!�$�1v��<b#��7�p0�(_�!�y��'��' ��.���&i1�Ą!��D�K�B�'�X���'�I�<����&D�<q�L�2�LI�l��yr�Đ�~m�S��!H��ǭ�!�y���+@�0�띑����gn�?�yb#�!y��k=q�j�n��y�(�1.� ��@*y��@RM�"�y�N�$
��r���@�Ց��'*az�#�����ӯ�'<�	��U,\����y����	�'e~�YHФp�4��GW5G1VC�I�.�
�#AjʗB���#�0`NC�I  Szq@�e������=%��B�I�J��(�Ż���C�Ǟ�>��B�6@����B�3V��!���jB�ɍ'������p�����L3 F"C�	�^0�tA��v����!	�>cG���+�	e��~����9�x�;�a]�B�X7�=�y�BW&I1CM�X��Z%.���y�-�ܜ]Ð([�f%��hŝ�y�IB�Q���(Ӿc܌�!q�У�y
� bd����\��A0%��x�!�S"O2 ��LǠr ��CC�M�N����'1O�����1�R$Ã�L��\�4"O|�ȅc�2�g���ft��"O��:6C	4N��a��
>E��k�"O8eچEB��X���	�zH�"O6|Bu�D�U���ɝc'"\!�"O��B �Ԑ,���
�?i%)��"OT��6W|��[�$��"ON��6�.h�,SrfK*TX"p�'�ў"~�uL�!4�Z�yW�"C�=��` �y�*�Y�\�9�FïG~�Dx��p�
�'F�h3V�\9(��Eb�#��A��'��t��[��R��:Te��'Ƭ�{���-I6�� �M�|�<p��'��!��˔;IN���%�EzR���'���c��z(eK�E�40�
�'��h���;U{P8�#�0ʬa���',���<�����Ɵ(��)�R� C�I	nEV���͸DK�-��e��2C�I`}���7����|5A���,�B䉎i|L݀PƊ1,�Pm���PQ�B��##��Wޢ�T�c�bס�" ��'j6�YS+@�=q~��v,����'Ny���T��� ��pLJ�'�ȭ�� �=o9R��tȉ��F�+�'ۢ�
J>3�*	�E�O�*��'�"�2��ϔ�YАBy/�DZ
�'E8!ICM�rIq,�m-�	�'�n��h	�	��a��g#Bl�	�'�<Y�G�f 
��S ,�h<��'��1�
�J\̲fˈ��P1�'��pP�'\�-����DI��'�����+�U(���B�_"����'d�	�f�Z�2�zr��Qc����'����skÁ~��|��KQ){u���ϓ�O�"��ڤ"�d�B�P��}8"Ox}q�N�H��j�@��
���"O����4u\@����}���A�"O��+1�	�r�n���ҕK�yy5"O:�i�I���Z��B�	�x����d"O�� ��^�v�j$@Q���"O����P]���ƕ(�0y��	̟E���0b9F�Fnm��@��y"��0����lN��zq��@��'�ў�O꺁�&@�)�Lp�g^%�dD�'��=�qJJ2o���/R�!��'� �x�M?X���X��R�f��
�'!l���M�i��\:�m!}]��
�'��T��x=�h;��[=]�qA���'JbI��Z�G����0G�[z���'��	��]_�|Y�@�U!U8�����D'��	�� zx� r�@���8�"�'!�$�[����T��^�Xa��K�^�!�DP{�j"�E�f&�]rW-O�2�!�޲.�Y� �
1&��H�L�X�!�D7Bb��3T��<=���x�W�+��P����I(p!� 
��P�)�� 㔾~t�C�I$O�hTHV��$**>�X��$M`C�I�=�~�Y��OGp$��A �� C�IO{��C�H�n�@C�
T�6B�I"+���@/��XTcՐNh�C�	�H�p�����r��&oH�a�*C�I��l�U��)>$#)%{|(���O���� h3q�H�t��A��!I(tR"O��	5(�3��@밡7?������s�O�졲� �K�L�#ˋ?>0�H�
�';��kK�
*sr(�ҥ�� tJ��
�'n�)�2�$(Ԝ��3��%��K�';��3�F�|��9JÇOJ��'I��{&�����&(f� 0�'ޤ�B�J�h�8��7&N�����hO?]��@݇
�"��`���]P�Q�i�s�<��B$��@�F=<MB!NJ�<	�H1ax�����N�v=¦�l�<��g��S0\�p���*^V�)d�i�<AWD�w3��ADޙbp�YV�_���hO�x���Bƽlծ]��゗~����C���t��  ���b̅�c�ȹ��Y�����JWiU$H���4�ƾ$ִ��@4D���$bŐ_�X�)E�Oo�h�c�4D������xu:ă�gA.!:`���1D����� W�E��L�g��Mk�0D���e'��>"����iG:N~Uh6)D��@H���X�hF1���a�!D�4R�o;@rR����e�H�(�O˓��S�Op!S�°#���&�P<o��;1"O����A�B>4�T�=r4��"O왑.Z7KQ��4B��wZ"@*�"OQ� $U5^���Z=[Z
\A"O��g�ל!�Q
a I!9q6ͪ�"O"y@��-2�u��O�.DV^ D"O��p��)M��I��B�hW,H��"O�`��a1V�*��0$0^��"O��DG.'O:���_N<2#"O����F����bK����"O�p��	�tp����+�:���"O�CԨ�<6΄B!,*m!�t�"O8��S�T����LT������"O|2�<E��"����5�☪�"O|R$O�;A���qI���I�V"O0�:'�W�5��Ye��*p}x|�A"O�����@�*©Z�F"io� ʖ"O$a!)b�M�!����P�"Oxm�7��+n�Ӳ"9�B"O6�[F)@�/�4��w��V'���"O��mII0}���
	}���I��|E���
΁�͒&$��!c�[��yR�V9��� ���:Gn���yRo	�4?vI��
Բ%��Ӄ!�7�y"Ĝ�]n��S ɝ	�:��cR�y��4a9�yj ��9 D� ��̊�y�k��oI�q!V� =ru��WO�y�&R�VL��8�N1n���ևO��y"�E]��%�@b�mkh-`Q���y��hTP���	�d2�����)�y�+�?�^|�"�Z�]i��Jާ�y����00l8��-T/��
�쎊�y��R�N���EυJ��;�+�y��
�Lb�}H�%�Hv�X��]��yB��������&
�N{~P����y���)>6����Pp16g	�y\�}����i��|:dsŉ���y�/�L.
BF
*{��1`��yR>�x}�dz�̥I��ʹ�y�O͛65� sC)] �EXV���y��X�'%��r�$�Z�D����S1�y�j�p��93"͆W�m���y
� ~܂�L�<Q�a8��T�7<�0�"O^u��^,��wN�u$+5"O�m@���J�	#w��;9�~m� "O�ȃgM�BM��J�� $ƺH�#"O�H1B@ R����Gu��uv"O���2D',tՠ�,�*{ަL��"OjP!���(32���_�*��D"O�4��J� u��Q�q��A�]�TD{���?94�K�m9/� �nһSxC�I�o$X��r���6��*eE��R�nC�I��8��VJڒu��]xRk�ITC�	' �P��d.�1�(�1� M�
�6�OZ�$*�)�t���ӫ �-��&
2�C��Ku��3�.F�-X�`��jv��:�S�OZPH4��AHT��*�Έ���|�|�R����x�$��>Nr��7OS�f*�}��E �yҋ�v��q�DΓ3N���4���y&S�w�&��'FZ0��  I�y�j[�;,��,�>�����''2�O���qU�܄�r�s��v4p*�',��;�II�z��gEU���`�'�A�6�B�$�Ժ�ؙa�*���Z���	؟@$�d� &
�h�j��e�%Y�j�h�\�<i���[m���֪��?A�e81��Y�<�u��Zɖ5��^�
0���Z�<y7�0F�bD�F��0\zp�f.X�<1$��o��1�Jh��]���U�<�Enŧ#��a�e�B�>C��Ii�<YD^:-�r4�����uA�H�Zx���'{�I�o.�8 U%�"8{\![	�-m�B��$|��ta�I��jV���S�[. ��C�I�p�y;Bm�q��2C��Dx�C��#x�h�j��P�^�����?F��C�Ƀ=�ܬ����c}�����ۄ%�C�	�cw��	���3dw�E)�Aĸ��B�O��XY�֍X�tI��D j��B�I�.� �E @���H�L�#�BC�ɤI�1�̹`f%��S�C�
#���;eJ�r�^���'N0C�ɵw�$�����:;4�[q-E"��B䉭j�j<��Z����C��.be�B�I�k�H�=Y��Pؖ��8�BB�I�fʡp(��*Ġuc���p�NB䉽	����� !JY�qۗ��M�.B�	�S^�A)I�&+t�"T�ݗ| B���Y��$lbp��H�.1��C��<b���h�>�c��8Q��C�Ɍ�"�(Ad|(%��.#D�C�I�'����#� c)����Nҡn��C䉅>8s�Ο֤51�]��C�I�}���cI3n�4Ճ���6B�C��0�L���H�v�q:F�׫,O�B�	<S((��-�o)�i����d�hB����E(��
�n��I�����e{B�/Lr�k��w�^%�vk�	��C�I�T;��:Aн^�*�XT!�	�C�I�*�ؙa�f_�mT���ԭ[���=�Ój�����:QnM�섑0�J݆ȓZ-�hS`ۦ�Pi�lBJ����>�����&E�h��bN ����A-&U��d��W�����Қ@�⸆ȓ/�\��ʍ6D݂�pub^�*�Q�ȓ"|$�E!�jx682M
S�F{b�'�ᓻO�RȰ��k��̓�
	�MW��<1+O�qO� ��S�E�!�.$K&��4�b<�A�'4�'��)�3�ڕM�T���/'V���&Ԅ�y"�΁	0�xD�D�'j�3�"���y��ngl\����(+؅0�⊗�y��q�`�xF�K�\��8�y�I4OҌ+LVxQh�O��hO����O
�x�TBۣ9�¢�A' ����4"�ҟ���M�IO��O�l^�C�<�&8
Qd� ;䰖'��'��>��:YZ9Z #]�uZ2E�QFLi^"B�	y�Q�G�>�ix�m�5.B�I�z�b�0�J[�6;�R�'w��C�I�+a� IS���I8�K!n�1��B�I�ii�d��E~!"��Z$����d2?q�K��~,*����@�$!�Gy��'��h(�"@	%�0E'��Z��e`�'�$T��)��8��$�E��;����'�x� 㓢}y�ƣ�8G3��8�'�ԩƯ��$�Fb�CU\���''�������TC�jԌJn6d�
�'�Y�>5�P�k%Äݾ,�ʓ�ؕ��,�',Y,��RiƀQ���ȓmmrH�F�ߤ2u���r�9i���ȓS�-�cT������%���X�ȓ挡�Gg:�Z�G�e�ScXI�<y��L�kO����#[�cQhEr�E_�<��T
A�Ђ1G���}Qr��yrkā�@Jf�S*)}�	�1$ڕ��>)�Ot��÷��!N
`$�5�V"O��w��MJ�Űĭ�18;F���'+ ���� 3��V]+^�n���'��\KP��(�lȲ�l�X�tq��'�D�� ˄[����c��!U-��'螺��䒓�6)т	Y7M���	ߓ�'�����S%���b'�1S�r<3	��'�<�I�T�o8��Mts
�'3$[C
ŕG����
� qu��	�'L������Hy`(i���a�ҥ0	�'N���G��g���ӭܴjy��	�'J����J9{ؖ�k�˖�c�Q��'Ռ`�v�ԧ/���bǀ7m�p��'&�����dN�|�#��c�HL`���O�"|��#0y|8�4�`��Iч�^F�<	񮒜�^�I���A���I�<�&��9R�4�ѭ��
�R}�V�P�<���0 m)B��3j
8Y(D�g�<I��_����f��.-x�{�L�H�<q�\�1pL��.�&1h��KR�QE�<!��1�r�*��b7���T�]g�<��*ϋ�ni��\��c�y�<Y�@��0�H��(PT64hH���x�<a,:p�Mj��Y{`��dr�<��Δ�q�`�93-
R%z�*��n�<��"T�~EZ�ǈ9Mz�8a�Kc�<!�*M�!d��� ڌa�:��f�\�<I0�Ur6aqƇ	N%�f�L�<��J��_�A� � {l�AY��E�<A��9a��X�C&s� ����y��;{~9c5o�3�8��#�y�$(_ �:��$zx�y�d�;#�0`�ce�'j<�l҃�Ԣ�y��5�Ԡ�� &`2�e�v��y��ҺB�P�*A�H�%�N��F���yRM��#1�����s�����O��yR�2'����hI�W[Tp)��6�y
� MAfaG���Ay��WM�q��"Oԙ��o/t@�v�O�.�R8�"O���a]5AX!P��ҳ"j��!6"O 1��Y���ؙ�گLJd9��"O��0���0���[�e�:l$���"O`��q���U0<9���/a;4���"O0t�����$��p"�˄:����e"O6�U@�T����N�s|��r�"OQ"&h�	07���P��Kg�Y;�"OR8hC/փzj��p�˗AqXpv*O6(��@�.h��x%��/�z� �'1�d�S�Rg�xuH� �:'��2�'D]�!CCC�Ӣ����'���%��&U��(�Ad�=���H|�"2&.��p�5��<ÐI�ȓ`��y�N�$P=¬��K6����l��@M62��M�]����ȓ5���2�k˝W!�m�T��*c$���>J���3�Lk�t0o牜u���j��E-y�`y� �jM�� �ހ�
��2)FU�� ���\��2i��:��K0yR�c����*C�T��"`�@����8����T�k~z��ȓn�H��VN�*3��35`8x���ȓp�Ҝ;ԉ:'	�H3����]�ȓ.�� V�M�p���
2ތp��$3:� #a	7�Z�BTMP�+En���Ѡٲ7BH;jކ����i�f(��s�L٠���{z-��F�?:t�ȓ[5lrr,у|�L<�b��v��ȓs�^�1	V��1h oԍ+M`L�ȓGh�s�D �@&��3�����[]�!S�H���8�B*F*yf݇ȓ(����t���y�ハ� Ү5��d2��;���Lư���R�W�(�ȓD���R�KP�(Ҁ���x��L�I;���&�f��b�[�k��9�ح�7�ڧ)aN�0���q��ȓb5\�b�O���I��8h����
�!rw!�]��v�O(���W&����]5��;�E#UeNy��E�j�ɠ��!W�ZM���Һ:4��\>h�ː��0!<�*f�ҶkR��ȓ8�|�Cǯ^��1єh��<���z�����%3�Q0%σ4M*�ȓ3J4䰱h�_s̈Q�יzl,��G�Li��v����(B�`���ȓմ�����h�`C�ﶍ��-F���0%%}��!��׸_y���f�R���D���R>��-�ȓrX��Ə ��ݨ�e�1KD����5�2�"�oñr���x�Z�fT�=��&��i$���( �U�$��f�����l�P��j"^E*���C#]�ƙ�ȓr#،+�ԥ<����%I9bt,y��h؀8K"oD�:�@X*u�ĠP0��f<\�R�f8f�"�ȓ�<�(%lXEd���`'�5S��L�ȓp��Pg�/!0-H�H7�|d��G�:	�F S"_�0�B�{����vy�5���X�r�� �Uh0�!�ȓ]^`�U��y)K
?)M��?�m���#X���@�,�vi��|�ٳ卝�a���-�0T`Մ�S�? �@�-�p�)�)�Z��G"Ot�䊙�g��I��-�^��X��"Oh�)l�7oq�s�Ѱs���CR"O�KU]#����fƌgd�a"O�#G�
�*<\MЅ�� f"O �3�b
{٣�Ŀ	!J���"O��lœ*io:YS�$֢Xj��W"O�q2���#�ܰZ�P�iR �t"Ofܘ�@���ʂ��#�bI��"O�I�u � i@�,�fl
���"O����N 2��[��;Jxy�"O���ai� ��AB��
-D �"OJ���o��D��	�(��"O��DW
}lyӤ��
	�J,"O�ms3#�eBE�
UH��bU"O�Q��)3XM<� mBoUJ0 "O���	�%5<!:s�:s9Vhy`"OH݃�Hm�����&$	a2"O����暤?�������Kg"OX8��E:>�>�2pj{qI�g"O���c��V����
� �@��"OFe)BKT�tE�q	b�%�$ę�"O2��cH�F�6��B�RN�A��"OB���'R%'\^=�@�!^��E��"O.A)��4
R��Tl�e���R"O��@RJ�c�pM5>�^"O�u����	X �VV�s�ܤ���R{�<�4�C�|[У�v��9�⭘u�<����;׈�$��=;X���Ko�<��M4h�2���偔�^�
�� n�<�&�6(lm���v�%��c�N�<��枏Q��ik�G��|�\yC��<!`'�.(��3�/V�^��}C��Kw�<I5������*Uj�XФ�s�<�C�*2�j�`Q0є�����r�<��̋r,�=x7�ɺ�� �C��s�<�c���c��Y��ӹ> �3��U�<�+C	K��h�F��;��S�@Q�<�"��2:,F���З5<�h���w�<�Յ[�\�D�FfNI�,�&Gt�<aK�O5>�ٓ@N�q�*�xq��l�<�Q@Z�'�6	Z6�
$�2�ԊO�<y��Ɔk�\ubT��[��X@"�Td�<q�A��s6-BF����i�6�_�<�P�OKt�����#�N�R#��r�<�m�x��B	 M�ag�s�<qbƇ�D|�Q�;>�\�Df�<�4F�F��4V�@6p�&cf#^�<�@�Wi��(B�M.(�}�P��A�<)��S(E�rM��G�$�ze�X�<�`��.~���eT-Q��뗮�n�<qnߤ������#�]�+t�T�ȓH��M(�W{�ma�׺����ȓeN8�2�j\
L(}�7�¸fmJ��ȓ<����� �$<��y�]�+��E��	���t�
8Hy�%������ȓ"��ǏƭX(xyҁ�ה�l�ȓ6�|�R�hN���ha��[M�D��xP%(`�]�嘘�'��]���eZn���kZ�Ji����ȁ\%����W�V�S��
!n�xq�çK��\�ȓ�����"�����ũ,p��ȓj��3��3� ]�cU�]6���)N���T�58�X��@�y$]��S�? Hi��A�KH�AIs���5�B"O�L*�K�8o�����ET�ԙ"O�h�4�ņ4��`��:�R[S"O�h�w��1W�R1�����\}�3"O.#&=���������˄"O=0 � ��t��E�?�xܚ�"On�3�̎0��kp'֪=rf��@"O ���● ���'�L!XXrT���'!�޹<��i�EG��PY��w)w'!�Dηy��t�L"�t5(Ĥ��!��
0i*`��
S�j� �"
)3]!��L\
2&��2z��cA�ȓ�!���;�.l3�@�tC� S%�M�(�!�X���rn��<M~˅ �5Ka~bS�����<��٦KG=S��Pb)?q��uT�-C�xu�`E�I�v��Ixy��F�����eO����x���yR/�	���� d^�
d��$a@��y�a'@K����Ĕ� ��|ـI���y���gux89g�=K�,aB�*��hO:��DR2^�H� y�=���t�!��~��}�Ƃ��BZ�M��N��&��O@��5�W�O�2T��c�;�����	D�����N����uc��C:�ha���%$!�dE�U3F��nG�Y+J���j[�@��=E��4k3Vu
Ch�� p�\�b0w�:4� �D��4� ��@�
�z+���@$O���*-�ɸ�t"P�ӹg�p�pMЕf�B��7lk���5��Id,(7o�59_��'`���3��~���S�Čm1tQ:QC��>�K��'$��:@��%#�07]>Q�7��Q��O���R�_�Iͬy����q]
�C��[R����:�	�!$b���ΓE�R"�h�(4I�C�IJ������@�l���B��M�˓�~���~��Z���5t}L�೩�	P�B�	�(f�J�ٗwW� W�Vp�p�O&��d�/.e�c,��^-�x� ;)!��bF�A��c*
�*�/F�+!��1��L��e��!��m�ю٫f���`��:�L�^�b�s@��^�VȠ�\�ȇ�	�>C���e��1<��ER㖶_a�C�	�%��P�`�K�aک05o�W�C�	:A@��ę��|��WԻ]G:B��6?:��!��5�@�D�7"�C䉣J������Y�|y7�,0��$G	X\kBJ˧yh���t&T<1�a~�R������yo�e	��J*{�T1�DL>D��򅏨(x���ʇq2M���9���ny�h��r�ؐ�jR56r	��"O��(.�7��D!5�_�\�Ȉ�7"O&��0�C�erf��)�,�����"O�ЫT��q� -�D���&�d���"O�*e��ǒ�:'��g�LQ��x"�'t>y�w���Xy��#&�U/uXv%�	�'!�9+pC�0S��"aD�d7�A��'�M�7�ی<4�Y{�:ː��	�'���Pѯ5hj��őx��(���hO?U��o�>#������:��3�`�K؟���Ew��X�v���+�K3q��=��"O2Ҵ��Sh�͠��n�.�sr��4MY?�*��¦q3�$��Ȫ?���B7D�\���%FC�}��/G��U���k���S��|,�R	ŕ\�vPJ��<C�	8X���(�F7[S�C�� T:C�)� V�2�"_�����M�&c��x%�	F�O7j�9 �Z� ��X��T�o� x��'\����.L�xr���U%�k������d;�Q0��0�6��,}}!�d��X���䁯k6(�"�
�~o�I~��H�)�0'
��-A�J*.<�آ"O��2ņ*����G�e'2�63O���g8����&W"q��Cg�"�z��)D�H���T���⢈�3 0"@�<D�\�Ѣ�A?�4�A��t��鄂;D�`Q�Y�"Fb�)�d ��8D��:��Yq�6x��jW*I5
���7D�t3���H���:�*;&pYB* $�,��E���LH(�>9p���E�y�	?�V�a�0Ԟ�@��yo�,(�"Y�#*2�4��(�MC
�'I�����?n[Ru�Q�I�Ap(}��0�S�'���E�[�p�� �G'L�C$�3bX!���JjD ���S:�@u�M�In��6�I��HO��]�~��\��Ս��<���,o�!�$�,��0�Ah�4&��Ma�Nٙ�!�Dz��0�����8*4�C�!��Cb2�;�aZ1{�&���.�y�!��'+�r����	�d�F���g���[�����`رe߆�Rrh� U�����I%�O����OPH0
;7R����D,;��Ti ��L���=��I	��2L������j#>9W�i*�>���*D-���6O�'h���r� D��`��9D��H���j����\F{��i["vJ9���'/T��� !�$#
��I��&-f�`��d9�A�	Q����ˣT�<� L<hzVչE�"/!�dL�s��Di�3^��bUC٤~.�FY��'���<�! ���	�6\wH�`� 1�8���^}���7T��.��>ș0#I�MsO��O�Ϙ'Cj�АiT?��M�����c�|���$Y�O�>�*��
7��-�pk�'g;���'���� 	5%��!Cό6[b�����x2*�{/f�F%�>^��`eE��d6�Ș'�!�קd���V���I�l��'�=�!)A�r4(X 1��	v��Ɂ�r�x���?g�ڹ�6�E�Z_|�s�e���C�I�h�����Y�T�P�C$O�^�
6M�<�M>E�ܴ2~hB&i�v�xX:$bK�(l}��U�@�h�M�r5h1�5���`9D����R�1�c��mL�Ѣ�Q6����@y��E&A���H�&M<q�4�'�ў�u�I�E\���2�%D�T|!�Ă`_�B�	�=�Z���2�tP��;(�@�O2��D�)4~��$BI�V
���"Oa��O��%�'"�!���#s"O�����=jf������?o��Pv�	V�O���ƫ�:l>����+d4��'��q�J�f\(�#q�U(*��D-OmDz���I�dh�a���F�$��B�Y:��|�g }�+��o��!p�IH�΀���E��yb�K'3�`��N�t����Ԧ�OT��D�Oz��b�ɕ�uJ�S���3p�#�'͎�p�ٙa	�(��R�{i�̃\�����i���*!�g��*F�*���yR�Qq3�Y�pGC	,���$�*���䓕hO�nA��θ8ң�@�MjwN�T�!��G;8� ��@�i��ȓ��uߺ!���'�ў"~"����A����,�c�#4�y
� �@h�o�Y-�����B�]�l��i���26IB#1T���CJ3[!�D�J
��o8>�yA�"�!�Y5s^)�O*L`p#O�!��Nl�xx6	A�Jhi��,m�!�䟨=k�4�鑵|���+Ǣ��I�!�ĞPd�����]�`K�!��!3��3�h�p�������={�'��|2�:*)\���5m@�X��<�?A㓁�dՄid�1
�ڷRij�s�-]�`�!���RI��jTL��5C^���<���9�ɫ���(�ωR�B����J�JQ�B�I�<���[R��(/�(���
�a�n⟈D{J?�#�O.,�ݱ�-�+<a��P�%D�@�b���@�K��[��j����$D��Ha��%�<(ۂ -\�&eh�`-D����i�=#+�5 �\6�d97.!D� �/S5L�,qE%>T8��:D�1�aQ3K�*m��n<6��<D�X�@�Č:^����$0��-:D� ��� �R�JPL�0���P�6D��!i�.u��������� p�/D���w�S9U��Ux-�0��S�+D�d#� K�>@i��[�p '.D���(i�<86cG� �1�'.D��qq So������lK4�X6N>D���SZ�-���¦�Eol�r�O.D���Q�K� !���!/>���'D����qo�h`d�@/y�D%��K�<������9x���E�&"|��:�%p"�Y!_`p��$��Rx�ȓL	zmq1�D�
Ոfo��d���ȓJ���I���`��9��8fl�9�ȓ"b⼳Iݦ.�����09� \��w�� ��
%8@��E-%�B<���<�!�a��^��˲�Q�6@ꕅȓDM.�[�.7c���A���ȅȓ\�Ȕ	��]#���`H�z��h�ȓ_z�P��ԃ�)�.��H��ZK.���! )|�yr3�Kx�l��ȓipp���!v�-*���&ń�%�����(e^�!F�� ���	|�Hv!��Yyּ��S�0�ȓ"���]i�����G�@&��0�6)�Ɩ�S��P�g��k�}�ȓhp�|��ƇE�h,�D�:	�Ԅȓ �"��4�D�T���#˕�
/��p�Ƀ�IT�3u���e�BU��	�OhVi��o�7Ѻy�dB׎1�C�	�6*AD�g�pY��p��C��^X�]3B�4�I�lC䉐G԰�s'L�!�`���� N�C��v�Ջ!@U=~lQ�j@�Ww�C�	�!�N���Y�`[4X���@�8�C�	�q�~Qu�4G�0l2�⒡P��C��xw�,��ˋ�+��x�W��`C��1@����ң�v����w+�QdxC�I�-N���j�!������nEDC�ɛn:l��?9Id���EV}zRC�ia���_3�`в`W9{�j��S�2D�T�K%nԼ�b�#��6�����6D��k֋�do�K�G\�=q�HЃ2D��`��=��M��N�!��ie�7D�xr��C	1�4<����y0l����4D�t�1'�z���91;�9��'<D�� tH���П-B��B����SÚQ��"O,�{G�ڨi�"�b���JAX��W"O�5#�M�d�^���mC��"O�u�N��HC�<��@�Z ��hq"OND*���o1(*v��1Y�r��C"O������"戳#��
ɶ|�"O��P\
`9A��x�L)�E��y�KO35RX�ӂ��f\Ĉ;e+�<�yR�Z>c��CUoX'R�
�`T�,�y"NR ��UJu%�>�����y�a\&Nj�8rF'(j�P[󮛮�yRH؎=����"�'p�#2��6�yR�ٿ;r��@J9��G�yR���1���?��,;A���y"�N,L�\�)�c߽ZoN�Z&��y2`ыj�z���G��^�B�������y�I�xL)���7]'T� F�(�yb ^�iC:�ɣ��%B��j�LA��y�\5}�AE�:E2�І��y�I���Cd�4D
@[�A
�y"�W�Aj}��_! ��){��B�y�ޒ/̺���G\(t���QS�%�yf�.z��f+I�Ƣ��[��yB�#�@�"�	?'n\����0<7H(rH���)];]�rP'ˁ�'�3�(D���,A�|O:x���_y��(���<��)�|6���K>E��"	���}��mn�a�@c@.�y2+�H٦T��� �7n|d� +�50��5j�А�!אhe���'��\J6(.+M���!%Y�O�D8�	 �]�$�Ǔ^�b�s��x�� ��W��d��I6�O��Y@Έ&�����!G�c��!+��ɃqM*h��=�O�,l�Ѥ˳>�j�� Ǜ�^�֨#�'�:���5Rl�i�OA�H����O�ɒ��{�YjL�"}:篑:_Lx���Dݱy`X�Àz�<	�՗3S61;cKީu�d*�N�7��I<P�,����.��g�'Z�KvJ)8'���Tv!^|`��J-$]уԩ��S���q["&�&��`��K�T�*��� #�o"[ �A!������)�a�!P��� ��O�Ll{#��RL�Q@Eݾ*:d=)�'Y�̃-ǥP�(�1'�E0|&���'�N	�ɼk��M����s|e��'���Ї���WW����/�#t�y	�'8�lr�0YVj�:�+�36�	�37�
�coӞѱ�/�R������CdH��"O�Ppp�C�QS�!��E#���	�9�\h@�ëPR>�� ���q�:`����>A�X ��� D�Й��D$B�H�e�	]y̹U�K��LT��5!_����'^�>�	CiR�j� ��T̈Eh�*FآC䉈|eޱ� ɿg��Ш�7�L�wl5�GB�qf���<O�p$��F�(*�/�=Ox��r��'$�5���Ͼ\	V�9��J�`!$�C�V.��e`��
��5
O4 Z2�ük�ޠ�t��l3��j2�ă6Nx-�%ѐu�E�f�&�O�"�It(�gN�������
�')��:p���sh�S� �"��J��.!kw��;FhH���*�(��	�]BRMp�V2J	�q�m�&6%2B��#$p,�+
	%*�T�A>-�m r�G#	�����R#���<.�iD2��-.��ak݀p�č�(���0=��� 9o�T  T��t.�Hidi��iXx(ۤ��uKP��E����Q�,�Dgǌe484��!­Q�D�<����,R�hsUӏFb�`�3��+�H�����f����%l�搅�W���A�b�(1�(@�҄*�`I�/	"��rs��Ct$A����Uyr�.�Xpg^T`e���,�y���7X<�<�r���uH�D�T���Κm��cI�.�A1G$�6N��1��Its��A��4(�|�!�L*n�j��dڔE;ܰ�F4E9��3� ��)��x�nX�@h��2�����dFKhP�# ��3x�EçI�bL���> �nZ�i�>��@�B-�� �`��[d�4ϧ:杷rVeb���)��Z���2C�		�R�"�[�fߚ�gkӭ��P��e������s�2ݪ�@N	�X�
V�[*dڐ�wk3?�p
�)~�Ĺ���V e�Xx���B�:�Z4��
���r�`� 	2t*ׂ5����b�'��ღv%pӑ�K+��ɵ"�� � (hvB<)4K��RyВOF,��Wq�|{�J	2��6펈%�l� %�ϛhCB��&ʛW��L2��ŏm!f�0���nk�B��n��2`�[�6��Bs�*����V�/��M1�/54@�Bi��l�� ꛖ7�7�F�	S ��;q�H����!66�&��8U��y��I=N�"�����But�1�E�%eo����L9[�Y�GF�bR
i"F��.�?��ePDzl�	f�P&ce�O�����6 E��	�EM	,��]"��Ɂi�Du; DN�W̤���&Ds���hF��b�'�5F���ؤȭiR�_8x��=⇥F��0=�D��<d02���g��4y���'�U?��Ǭ:)���S��?D}�L��!0x�'?�ѩ��n���`�@�~�L0넄[�N�5I�F,D�T���C��8y��c��,s� C��$*6��j�i>����犐3���O�x�<�cRd����m�0f���4
�_���*�'N}D]pE�4G��B�"�>U�#�eU�\S�O �&���#
�a��=���=���$��EY�xG}��w�ӁZ.HO6�y��7`��Y?~d^�( ��H��H� ���D�!�D[���IsCF�'�*��悓Z���1��9��M6�x���M����|$��b�^��i��^���%"O�c�Ď#s�̛� S�'��k`Ł 9�X� ���H
>y@r푾W�g�=��\ ��]�EJ�%:0�u/t���."~���b�&��	2��;0�9�@�.+2oڶB�x3�'����DA�B2B<��˂�_�tђ������ ��
Mj��5+~>�x���!��y1���8t@�A�)D���-d2*��	��~���)#ʓ�<�+T� �d�1�rț�Ԃ�hűW��C�$�
��%+�I1v�X���zI�6-�2�`�#\�-��'��Y3��/��q)1��!N�0�(D�DAV��X-����3�u�[��j��1�|b�;�g}�ڥ"TZ����֡~��d���7c��Y�=aC�q���	P5��2���/�������ЕcX�0���2�'1���T��;(p��D�����m*K  ɠ����C�P���?M��D���Sǅ��Zȸ�E�jgay��K+|��!��^y� ��x JM#5�ͻW�䰸��W���'pR@8'�]���G�4@��0�2a���E����E� �ē(��AV����
Î6��ibFcD�%�����	��5��1#f��S��(��	FLଋ­��T���v��-�11��Nz���4X0&��~&�T�3��(3�E��
�=���]%=��R���6=�������C�R��IlIr$J_!s��d���1��@��ā,J�P�{����y2�P&SN�Ћb�
;f0M
�����<�G%�z�H�Df�<�O]/d���ǧ�\�؝��[ܓO�Ę�s-z�x#~B����Z<�6m��x�"��p��_�I�_��u2��=��?ʓ)I/p�c�H�$��y���O!>��4��|��/�g}ҡ��5�"�ׄ�^S�A*��B�*^Dp#�>��Ç<Y���'����So�M f�C�E �:@� ��?�R��$@&�O��	�ḑbxHa"�� ��"�W�#E�Tz�@�%��>�phȈH���{�ɵ��P�ƮvX�,���h
����]�,q5�o�� ��((l��A�8D���!�e�5CGK�	Q�� sf�3�dW	S��4SF�3��['ˀ�V0��ëX*�Љ��"O�b�A�aZ���UȚƈ%P�Eo��=)� �V���d	E��!w��^���۳��0YP��9	V���I����Q���6�p`�� ���d� Rq��k�'��Ij ��X�)���&��@��'��z�*���I0�VA�p�J>A��@�t����!��'9��n�e���=	����5�̠%�Z��$� �CU��"��D�1i�:A�=�Q%S8V�@�S�IOeܓk'�>���^Q&�3c��6�j��w G�Q�x�E��0qLp�I��@`4��P�:X�l�;���٦a��P�}|d�a)ИQ2 A�hZ�o�@�J�ʬ¡!	�G��ҧ�i�51���'��#���5���b%��{Ԥb��� \�b�)ϤlX��W��e7x8e�>��O�.�v� ꘊP�ODϧ~���e�B�&(*�Y�y�Ɇ��~��[� �<o��2שANax1�� Z���fOJ�i �ۢ�Y��&H�\������IU���	PZl1��<��Ш��P@$#E/W�,QҦ"OZeх�H�*��E�v%��g5 ���O�E��l÷.�,�I��}�Z�9ܘD+Jp�`�&'g�<Y����bm�$�7ǙR�hA��c�D����̏��0<���^����1�Ow�,e�KS؟tyB�ߦN��R+G#B��
�华P���A	�{(<���@�Z"bU1� G�\8�(�F�'ln��u��B�'�FQ�A�X�Bܢ��V#D�������{�ң�lJ�J<��(�ȓQX&�r �Q�J�3c,3�쌄�Q(�m��H;�`KB�.�&,��nd��F�\�Lؚ�,��B�����~��H����#x�pb���	r����ȓ;���"c��:`�u����&�"y�ȓ&r(��+�c
l�x��?cs���� �P�4�^d3� D�8'�ܬ��X>j���n�E�xxA��;��=�ȓ:��I$��I��A�	ּ��o��;�-J, �]�Gt�5�ȓ#U��A��٘2<܈a���N�h,����Z���$n��la3�ƿ?�-��|=�@�W�K=w�� G�J��0��ȓ[
����C04����1e·@���,��9�%L�1i��!�u�խb�ڌ�ȓ�>�ۣ(�U�֙�'C�w��Մ�E�F�	ef�:��i�a�^`U@��Q���BS�L�pL��.�/2�؅ȓ)�X�S!"id�������'}hm�ȓU7����]VILUI�ϩ-�1�ȓm�n%cA�Dx~�PM�'n�H�ȓZ
6	�Ɛ�LQ!�wJt%���g6�`��F�Z���J�dl�ȓo_�=��BX3l9�U���l��ȓc
psdӞ�L9樑�x��T�ȓO��cr%��r�&�bU�=~f��A  �4˜�)��<���2Q�*��ȓ{�$}�vB�1����&���F�V��^��@Kp�_�H"�p"���A'����!��L��.ɠي�J�"����q��QeB"s�zt�ggA�,Xąȓ[j�L�Tg�%Q�z� �Q p�&!�ȓz���)�����
�Paߠa+̥�ȓ ��,�`�ŸS� 00�ݛ%}ĩ��qA��b$���-��;Egؐ&8�ȓZ$��h$钟'�蝃1�KkB1�ȓf���)V炋N���H�WՇȓk0�q�bӯyB`��J;c�T��lFީ�'�_[��L�*v��P3�q��dD/V0�A���B]d<�ȓf�1�"x�6�'���+Ԝ�ȓf'���`�=6�̊uf��n2>���;)e����}6؄��a����ȓ#�@�QT?$�V�+�jܻq��ȓ&��%ʃ	�� ��u�N�0n�ȓb�Nx3��ʅ![��!D��.5�.9��:�XB��7U�I!��і��a�ȓw�PP�EFƒwdJ�O���Y�5D���a=6��X�ů� ?YD���0D�([��V���3� ���.]��#D��+�+͸xv�U`�/	 m:�D�V�:D�� �a���إ��@�%�B"O��Pa�), �K�O+:�Y@�"OHQЁ�:ZĨ1��º*T00"O�H��nj>���呜����E"O��Б�X$4��qz�@�RRȴ�T"O�D��Ga)E�q�W�8���"OjQQGԵ��h���V�zL��"O�:W���*Jf^ .�*���"O�#%�M#68
���
=�U"Ov�H�'�+e�&TR�/0q�f��"O�,�ѩG�V�|]b�,;�j]Y"OIDX�0�R� ��@s܁�"OF�[���,�B�B�>
~�'"O�=�� `��CX�R�Y"O5�6a�0��K�+��W�(U�"O�q�"RDP�� �gA� ���2"O؄���m3�@�f��=�xm�v"O���m@��
����R�*l�"OB%+0O�tE����M�� f�I�"O���Y�Q�E ����l��1J""OFp�'͡5m(ԪC�-9��f"O�i2�AZ�Hr8�j���8 �숙"O�5��Bҟ_�(!"��\���C�"O�xk�EJ)"�h�� 	%Ҙ�#"O���pf��ʒU�D d|���[�<y"�ړR���q6څ]�p��'�V�<1CT26(&@��CtkECFP�<�P�Ԁr��Љah^Kw��aE�D�����N�B�qO�]�7>�^Ͳ�		�����"O���"�!1NaZ�ѰuD����Q�d���E��%��|jg�(u�,T���ȓl���ȓ�C�ǉ��%!�'\�%A�$(I��c2h��@��aH|�>�s*�daZ�`�@�N���g��e؟x�4��� �bЂ�4�吅*�;/@��B �.�2�E�nZ��C��d���'���O�h�"�_��9;H~b����Jn:Ո%ʞP<"]xG.WE�<���/%x�a��K<��M1 �T|}�k�:T�mD��@�铍6=Ҡ�����0 0�)�v�C�ɱ	�(�`#@�aԔ:WSR�O<�y���1��4&>c�\p���0o;� i��K�I�x�$�/�O 큐B��*|4Yq�3L��p�Fחv���� ���?�"	(��< P�,لm��HLH�'�R���@�^21�"<�#�Q�0�!��x��"Op-��)
�@� �A�G�k�(�"O�����,��k��.�.���"O�@�󊐘C,�( �4���P"O���a�J&jXƌ�G X�v!H�"O$dqe���*�C ���-hX��u"O�̉���>K�r�Q���8���T"O�4a�l�7�Ԃ�aD�1)��9d"Ot�{��D�LMj)bsb�y��R"Ov���i��l�̩ڴ �*=�nx�"O��t��K���@�n:�69k'"OR�Ƀ�	4�D�0�-�Q�`4�G"O18#`����Ӆ.�8i��-�"O"��&b�k��Y�a'#� �
�"O���&��.�q��&��
�f0G"O�ɠ��ćNfmSq�]�b�!s"O��yGL�!|�Q��2(����"Oj�RW ��_��	����r�ܩ+s"O萺P��+?=�0�Ѫw"�!�"O�A�`� W�� �F�^�{&t|��"O���#�Ϻ\�h5��JJȣf"O�4�4-��w]V)���]4�:���"O� qp��:xYF�XB��f`2���"O셂�K�c���p�`�'Ͳ��p"O�b���q[��#!��!�6��"O-@�n�=XR\��ɧt��}�d"O�ay�f�r[*�19Ħ䐣"O̝��:>}����o�8^_%�8���&��I�a�Q>˓W)�xhrɌ��� ҲlI6bxX�ȓm����W��,x�!�uDL1v�"P�&��;}2 ��'[�^E���d��G��ӑ�Ctaʁb��UNx����*��wfƕR���"����q�� hu�;iG��^ R4J�I�<�r@F3M�����㛰hD~�IW��E�	�jBn���W�+p�t�]o�O�n�C&�-�l��N�=m/�1a�'��q ��� 5���B��Z��u����#�=2���*�1�e�ޅ��'��'�	 u�+<J��Q���
�B^$h;P*�"7�\�04��r�؝rp�߈Ah5"�)	F4|�Y���azB��n��d��F7S��ٛ&#Q?רO�&N�7Cf\S��?j8
��OP�oc�cFi��9��=�wKYZ4��'�4a�)�	D�1+�i��H��yB�'[F�`r�سH��mB�̒�o�$P��eH�O���V�?�N4�է�7F�$�C�'F�r�f]���Eٖ`ݙ4��9a�Яun����ț�nέ)c�����6*�1O��y�B֍{�`ű3)Џwn$iPC�'�L+R��"����c��:�"ѱ0�Ԏ òT{2����EN3Jq$!דBƖ��`��,�6x � ��4G}B��.:��R���Š	0	;t��>EP�&�<?�����P3hp�d��"O�|i���\Tð�Q�{�d�k��O2��d⛄(��L��}�#�|�JY�N�d�� O�<q��
14���ޏXK�)����a�d�=��kp#���0<�P�@�))�#�HG�[�d�S��v؟�6 F�V!s��=L���	�v��[�*Ur(<��M�B��8 DM�2�v�׫�n�'�J��@P�$<�5P�$[�y�(ё��^
q+Nć��T�
T�S��X
��
(�Xl��.����^�)�H��Q,�=Vm�ȓ	�9Q�l:M��@�̕#���?�R�Y!;�#r%'VSW4����Rrzju�3(�l�<�p`�.{T�2�iڼ;r��F����ʒg5���a���dˑ�d��P�bH`ѐ#��'v��{�S���	18R�0!��u�6��т��P��Ӈ��ն�p�M3|OZ1s��no0	��'M24I�ǒ1)��&3�q�]��B�Wx(�I$pcF`!t�7��*���򤝻@��8�e�ʽ��D��A�����C���!2@RqO$�/`�ڌ�	
�`0 �M=U{�5��D%C�'���+�L�N$�HE��j
�{�8�3�	U#>d6D���W�����gj�?��	/N,Q>�;��*u�IDl<��&��|4���S _���ɶs�|P��L<�C��:�H�A�(D�(�<�� Y�:&�U�c�1�H,���7H� ���ś�`P��2�(�;g�8���NA
S�%#&�	3P �(G���1X��W=��
�V\�z��F)3ay2��2#�0�����MyH�p|MڒΘ:=��%Z5�$��'��*��E�G��B��B���|���^(R
H�I<�EY�V�,���%��`� ��e�7"��ti�� �(�c_ԒO�D��O��ʣ)R�~Q��@��A'r8f�8�.?�&�'�zЀ��#�3�$��>�ʭ۵͟
UY��	b/W���\�\�����ɟD�.�)��ԏK�JE�ݡG�f냚�\�d�'b
la�HJq�� ȃJ�n�+˓�4ڄc���E	�����ƹ/������'����ȓ@=��&ON�=j��ه&���'���ǧC������S%6`	��G�x��\�Fˊ=�B��!re�E�$���Ƞ30kJ�+�2G�\j>�o�\��+
0Z�)�f�,�J�ȓ4��t�kC���sf@?v�ȓ]�k�f�0��s\<Y��i�ȓ:B�u` ċ Y��˸M��%�	4�K�Lay�H�s��S�.��3fhș��?1�C�3n���j�(e�1WɁ0#���ѶbƟ�Px
� $�SՇ�r��Rc��cB ��9Tx4��QGO(4�1��k�J��2ߨ��t�~nDQF"O�hb�l���@a�c�=K� 2�O�|��J�&�I:M��}r���mG��s�b]��5�Pe�I�<�΋�s����#E�gD�ɳ¢�K�dŐx��e$�0<A�/�kܜ-Z�7Μ����p?�%᝘{v��(�BJ �2H)�'ѬkU�A��X
A,�B��%,&�y`��ǏLL�qB�a�6�>�2�@�f��$.�/��T�*I��H8F�I�HC�	�8:r��OCGܙ��6-i���}:�@��""�S�O�����&J]�X����f:YC�'L����cE;Vޑ`�"P��"N��3w �F���[U�'Iĕ�'��<_
����їK�,��ߚ�5�
�L@ǨңC�x��v��R�����'R ��a,ɞ��xAb�^n���;����%yr�:������AY������k�R��L-�y��Ja��SHLT`y���ވ�y�!�2�a�Q�T�H�Ĥ�i��y�Bɦ` ��%,��K � �䑻�y��A"f�`�� E��'[(�yBa��4��x�'M��B�"�$T��y��P�w"��R���&zSdИ��y	k�t�c��B!i���f���yb�,/L���ީ?N����yBA	�\��Q&���d 	��"ڙ�y�!S�oLY�2�'Z��p;eC/�yr�'��es�`U8ڠ�`%�ܶ�yr!�(f���E�Ȅ?֦�g�̘�y�<�ހ*g@E�y����Ǝ��y2HLX��̳Ņ�8uLc�O
��yN�(I�/=P��vnWPN��'aNpy���(t �uc�PH���'�P���ީ(X6��KM*-��'*z�A1�f�� �S�Ah
Ȓ�'�V�k>��=�Æ�nL2���'hd����?�v�RO �r�~X
�'5|�j�'� �$a��G�C˚�

�'z��!e� >�H��A��D.@�	�'�>����8�%A�qdj5��N�<���ǄO�L(���U���N�#	�'�z�F��s��U�b�{�"�Q�']"1*3�KAd ��wa�6&j\�
�'�B@�`�ЁV�����/A���	�'`�p�B�-���'<2pe�	�'��m2��I�c�}�uL�L|	�'���c�F�s	iƅ�9*�-	�'M���%��LP��`X�>����	�'B�Y!d�oLa�sEF(-�xS	�',�#���������*Vb���'�^���gF3eJ�]�U�'=�C�'D50`g�}�����!J��'�!Y�˳ϐ��d�#|�8���'0zT��Ą0����F.�-1��(�'e��A��M��| �MQ� ɣ�'��l)E�9q�v�A��8�B�*�
�U��cשFS���������o];N4��z�&�_�4%��8]3`�J�K��b�ٖ]RP4Q��OXX2��U��ᓺ!x���b� ����0�	@D����2 x���Ѹ��Oy�(�3G�)5V
lCC�[(B�2��� c��Zs���4eqO?yBt�ز%+�ћ�+[����ŢħD��)S���O�4\�#�_1� ���Iع:�"�k���'�*�'@�`�����������
�V�d��<��*��V�f��(6�'<�)z3�&\�(:`������'�4劐e��kF\츴l=�'u9z�[��І<���g� �S�θr�-����F���y��;��*xz6�Hr�UNc��v �)<���	C�0tc,�)�'�� �0p�-O���G�h�|*�H� �X��/��)�^%c�$ �D�U2R� _�:�(���fJ OFqrA�)���`3��+��th�@'�b�H�|�# �'�`�@�O^B�x#d�%C��I� M�/l����+Oɺ6�ô!���n�h��򩔫�dd��� �I�'�F=xRH�"pm`h^��'�|�����zW��q�X�0G��!�� d�+w$�y�'�NвG�к'������S�F�D2��WdM�^�$I�ҝ>�Ï�$�M�<����9w���(�0<@T��J<G��I�D ���}����h�tM��j�,b9 �cծ��y�m����O��'�ZXb���Pk.KR�ʃmX$��'���`�OG$�h�C�!��Ԇȓ0ؒYSS��-
J�6͔" � !��'��5��R�7~�AoJ�m;tP��'����.��1��,1���������'�f8�ԃz���宜"�:P8�'>�&�7e$$`HUk��4���'���#b�,CuޕB�
̴e��B�'Ԛh�̙�N��ġ�叉}�.8��'��e����2hP�@�n��'B(ikD�X�8�2[��=u��8�'5n� �/'�l�U��*|P�9�'yQ[&Ȋ����+u@`�'��T%L����BN� h4D��'��DH�eӁw|��Z����J���!D����,� ��c2�F�f��@�"D��[p' 2� 4ir'ڳz���9�!D�p�&�Y3$r��%��.Ӗ��4K3D� !4��=&Q~L���
gq�(���2D�TH�l��
Q���6k��.Ԥ��5�:D��[�*/#,��dG�=��k�"9D�dZ�(8|�i
E5\�Zؐ��9D��kW	�k16���&3�0�6�;D�$�$�"���#�
%�^�x�,8D�,Ǟ.9\I�q��������4D�4�׏�,V2Iɒ�gM�(k��5D�ದl@Kii!G��Ul��{I D�\�%�ж���B��8t�8��d>D�@�H�:$���Q����YW�1D���4�*��0 �⍸r^f�a@�.D����
S,��­
<q>42.D�`9��x�ث�d�	B
�q`0D��0U!7�hiI�ON�HՐ�.D��1��;C��P�m�t^�my@k-D����q�"a9��N�QC�+*D�H�ڂ�C����R+�,b�x�Al:D�(�S��F�>��$#K�r�~��7D��n${������
<f�� �S�5D� f#ɩ]�|�r.J!l*�5D��(�ϙ�}�lpQ��E%,���ц D��bc��[1|y1t+N�O��:1�!D���b�8ab����M��xc��,D��2�P�?g�݋���8jn"')D����,��ī�̏'w4h�@G'D�!mM"}j	{�J�(t���e'D�4�%3�VP��
˧,Z�Qb��&D�@B��]w����	5��a&)D�ܺ��'�%���I�cո�Jg�'D��:�)N�qO��q���0bZ�81V�&D��+f��y��٢����>fV�ɴ/*T�x��dE`���ڋM8B��v"Ov���-2~���) ����"O�J������������5�2"O��j6��`qp ���5p�"O�@�׏�%b��xx��B-2��Z�"O� �1��c^�zQ
s0m��k"O���Q˗�j0��-��AI Qї"O��[��ļ$��`�,�ҵ7"O䴫���{�n����G��0��"O\@�F�ԓc-.8 a7*uv�s"O-B�k6غT�����PjN�8�"O���a�	����²MƆ�Z�"O&E"�!Ι)F*!j`��S�DL�"O.�S�M�v��"��
�J�Nu�"OJ��k�x�l�9�K�(I���y�"OdyC^9a)J�caAϺ]�|��"O(%oC7A��݉�����"OV���G�4HPލ`B`X��0�"O�]x�Nɔ_�N�(p(� e�x�a"O>āt�P�g��5�T�P�.r�٫4"O��� [	��p3��Q6O�B1"O��U�F+M�b �e_�'�pt��"O�U�&��{М���CF���q�s"O&��8A3z�0p�ќ#���"OVuj�\�$H��H��V(�"O�����j6d܁�Aȑ=�d��"O�جkc��wk��r"O�H#�fR�.c���O�74f� `"O�|��FR�9g��u$�f"OT���\�L���3/J�X�
 T"OPDS}_��mܔ���a"O�����4t�A��:K��"O�+��3bD�p,�����"O�	����2��S�гsd52�"O��ɦ!�$U�,8D*ٽd^v��P"O$	��_6Ea�ٺI�8Q�c"O�@����Lp IH��7,�^�t"O^�:v�¿3�R���O$3��YK�"O�yc%/��(��9`��Z�]��tr�"O���A��63�LA��ÝAQp��D"O���v�K�l��ܡtOG<H���"Oީ�"�_n��R��2j�&L(@"O^�K���X=
l�2�@\�-�F"OF�I�?)�V�c�;iߒ�§"O���A�+Tv��[�*�;0�(@s�"O�8)��R�^5R�pʅ 5`�]��"O��k�jȺf��'�c3�9� "O\=9�$�d#��q��4[���"O�@�2#�%V'�A�+ߜ-�셈�"O6����`��B��V�w�.AÑ"Od-ˀ���UE��c4n/9pJ-�P"O�T�3�N3��L`�"*n��*�"O@���'Y���]����-jڽ9E"O��P/d�aA��\,]�B"O�����lX�Y�Î�W�T��"O�B��7�T���`\\���"O�����-\��#ρ"3��@"O�p���*|�BXq�����թ�"O�1���;��5"�8�"���"O�EPq�N�=��l���º����t"ON���b!h���{�#X�Ζ4��"O�g"�	���X2cJ:-�	$"ONuaV�X	���a�>q�Ѐ�"O��@��P/5�L��A�ƢRV�%��"Of��2�� �HEH�.�QR�4��"Oj�q@'[�)g x�a�tH�(p"OX�1D���)�x���cB�)�U"F"OBD8s�[$Z���#ޖ6�२""Op����A�N*��eI8�"O� dys�)�Y�Z�[u�=E䀲u"Ol���
X%E�H��NW+�A��"O6mp CR�CQ�$�P�M� �(P�"Oq�&��� =���%mJ<(	<1P�"ONh�ǌ_2uP�X�ɫ�� "O�]����/Ov>��f�4$����"OfU1���
Q�"���A?e'��"O�ES� :j�85��+K.�L�� "ObĘՉIw�xE���)�Nt�b"Oh�O^5O�n �w)R;3���1P"O.����I�k�aQ���}xV"O2=z����ZH�"�I}&8�7"O60��k�[s��I'��N�<�"O�HD[�}��0Aԗ8�֐�3"O�`cdk1	T�=87`������"Od�D�e��բ�.�L<R5"OJP�Qʒ�2��yd�Q�d�!RF"O���vD� �~��4/� ]
�"O@���f�"(�!HU�"�TP"O��+�>L�ћr̃:MlZY��"OZ�PG�I��dH��L��S�ّC"O��P���.Ana�k���5"O�t�FoS�O01XcoYb�<�a"O�y$��:y$(�� ę9,t(�ٶ"OԴ��a�N����� L>9"O�q{��X#/���˕(D.8x`96"O�������/N*�Z��A�R��2"Orx��ե=�$\�&,@��0q"O<�E���p��EJ��5�����"O�Z��\�d��xxt�X�u��kw"O�� Ώls|t��(�3v�"=��"O&��U䋜2fx�*�d�����$D��k�ͷv�>�H��_$��$�#D����K��R#p-F6C4��i�d-D��j�K��F��5��DB87� ���7D������ ?�e���	$Xŉ�� D����l�B�V127�;nvu�Q�#D���Rd�2Xa�ܠ�/`�F)� #D��0�IN*s��0	B�^�U%�HRà-D�4���.B{J�8qϻ"렘X��7D��z��PGl��t�O�X��
3�4D�<����c��۠�N�h�ŸqL1D�H���źA>��8s�0%-zep�C.D��Ib�V"*�I�ToH�E���c��-D��;��F�T̤�Hr��Xuf��E�&D��+���5^d��P$�8w@���1D�sd�ҹ_�z��N�R"��� 0D��҆,�,� Mh��K e���.D�$�fi�<s#���$�]�N�X�@ D���Tk��IC���Bg�>��1R�,#D���K�,��� Q�U����B5D���#�Т#J4He�� P�s�k3D�� �^Qr4Q����&�%3��1D�� g/B��!N:[%2Pe<D�|9� T�T�*�˶Q�~Ж 3�4D��ӆ"ϯQ5"DzB���h��2D��` c�1*�x9��K�U�<Bq�/D��Jp�L�Y��pˤ=K���A-(D��t��m���P���~��:T�3D� ��\)2�8 g��`8�+�n4D�����'m���q����X��@K3D�x٧'F�g�����"9b��rE&3D�<����.��H�RŖ.&����$D������H�f<�u��=�%H# D�� :�Ivn��m뒽y�ʔ���}�"O���c�ǧ�fx��	�(� 1�"O��j .�&$��$��L�Y��"O�`{���^`Di�r�G>+�$h(�"O���
l������&�H��"O>�1U*�.(#�X
dS�8$X�"O��Y��W�f\
�d��*F@�۵"O�h"'J�%�j�F�" S�"O��0��W�O����:{�D�F"O�����L�
�����P��0t"OZԓ�JS(�a�E����"O� %l��T��"�`�+%x���"O���j_6hra@*u���?D��ò��;�^ �Rh�	=8m9��0D�l; fO�*���;� �/R��B�0D��B�k*L�5NU�M4�20D� 0!�_'`�`�FU�=�LCsi,D���"�dN�0�����g�&D����ΌDƪ%����J�j4�sb?D�p{,��Y�J��=%;�tV	=D��S�C   ��   �  f  �  �  *  h5  �@  �K  WW  �b  �m  �u  �}  Ć  n�  ��  ��  N�  ��  �  D�  ��  ۿ  2�  ~�  ��  |�  �  U�  ��  ��  ��  P  �  W � #$ �, �3 �9 B@ D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1��2*Q��'/�ܱ�Dnٲ�0�rG-E�ws���ȓC5p�yaL�!	:Xy���J+K��X���N}BI$�dH�ѮI�4�S�[��yb�_"`3�a1�$�H��5p�+Ϝ�O�"rl�$RB&��JW�z����y�<!�c��rrY��/�t/�u�e#Cny"M+�S�O�t$8��:���ӇԢYӮyz�')�T���܂f�l�Ë�Oې�s���x§�)9��Ź�.
r}\�K7)��y��)�N>�͍�_B�FG�>S	���r�<!���5k��y�h݈��`Hqy¿i���&�S�D�ˑ>�����F6!�ѩ�+�yB��$�xRP�K.~Z�CK;�yfΥK��p�&
�ۼ�� K	��y�ggd"|�ãY�V@�P�Z��y���� Vb��aӐD��Q�������c��"<E�D'S!&��L����
Is�UAO��yrkǴ�;���/���tH��y�:~ls�	R�(���)�N��yRG��U�X,�d�!�*}�Pf��yr�gq@=)���LÞ4��G �p<���8����ԓ�f�	6 
T�!�$�9-"�"P�3��D�ׁ��$�!��B/�haB�88�L��A=gU!���21܅%�O��l �7P!���J鸜@��%��@��	��w4!�Ěe:b��p��{�,�I�D2w!�d[�-N��AҖ_KtP)2'�h�!�d
-r�ZP���0I��9��Z�!��H�s �^�v ¦	�!�D�Җ��S%O�`�9�V�Ҩ?!�D��\��i3�O�Ih؂����_�!��U%0����HAzTXȐ0aP,R�!�D�~�$0�%��|K4Qj�@��!�A��4�Jt�"3� x)�O�!���b�ѡ[ t��{g>�!�Q4 �F�"wőjrN\���R��!���V<�
c�[C���P�J=Kw!�Dξ9W�Q��E�|������W��!�X"M���[�sHȄzDG*T�!�V�@uمʇ*�m!F+�!��V;������e��"J�_!�d��)�j0�V��QВ�
�˵q�!�B:�nQ�Q�̇D�T���MZ(}!���t�}Y��[�:���Ǳ}n!�dE�1���l�>E��#0tW!�$ �GҼ���HU�̘0b221!�dY�b��
�,�!�ڜ���9�!�^�:�D|JT��K�m3�@�g^!��>[h�QsG�e���p{�!�� ���ր�$OK�]Z�hB�1*Q"O��@�08��ȓ#K5����"O.4Be<* �7�Ȫ�n9�0"O��SD�I�#��;��=ڄ�s�"O� r�xu|�[�/K�*ר�ف"O<@�VV8y�P��$y��HzF"O(�x�Ō2gd@���V�3�v`+�"O�V�E&\h����8|~֠��"O ш�C�NX�����e�}�"O�Y�wm�*H���C�ei��[%"O��Bb�  �M��C\&VP�P@"O���ŋ7lP̢1�O�$�|��"O�<�+ �}�^�i�`��*9K�"OTR������G���Y���$"O��{����d�͌]���@�"OX�Kŏ�56��A�D�0�&l8�"Orܪ��έb��%�S���iia"O�ᆎ&7�|��Qܨ� "O��P���_�D���=n]-S�"ONP�t�\-6�=HR�#Hĭ!3"O�[��קBy�a��`��)84��"O�,�6i�v��������"O0��A��"P�a�� ϗ �r<�#"ON��D��ą�����T�W"Od�hG�^b��C��.L���"Obh����n�$��R-�.wb1�G"O8uA�,̎k�D�%��ro<]��"O�)�T+J:Y1:����ªT�[�"Op�K#�׾4\ʔ��8HB� �"O���S��'7��Rtm�^�j�;0"ON̡�o��%Ⱥ��&�N�h�Q°"O
�B����qZxl#�k��KA�31"O���d�ȎR2�1�,�%	�y�+��X "N "�B���yB��=hq`D�[(K~nQ{��9�y��$e v�a��2Q�0qi��ybc�2N4��cF�$�Z��aR��y�	�;�� ֬�%D��b�g��y)\��lt3s��a���X��y��S�4hA'MG:z�@��5�ybJ�?Q ��o21Ëն�y�U�/t�٣`�Qo;�4;��]��yr%6c$c��d_q�A�B�y�Cr���D	�Vy8�"N<�y2,:p82� g��*�֝B�C1�y��9fkL|���Ͼh�>��⮔��y�g	�Ґ�Y#����@���yR@<O���7��+5x�X�F��yI�
k(��^���J���7�y��(vH��`�I�Y��d�`�&�yZ�1���%F�K5�u�T$٨�yr��)Ph$\���=2��h��;�y��/�H8s��ߕ'���`�щ�y�-����P�%>"�z���Ԥ�y�ͅR��%�)�`D�����yR̎Q�Z|84��k	}K�˲�y2�.  9��+�c�}��E���yb�L�@�T\��7b���ɖ��yR�
�t�E��"�6������yB�W� ��A�5oFz��˰��y�B$h��f"�%��1�L��y��'=�v%zt &�R,@0)Z��y�+�6Ы��U�R(q'!B��y2j�!
w�eZ��D��zq�ݿ�y
� @k�N��:*�1�Aͩj �-� "O��CE��7!�VLbb�ǿ�"Ud"O���#� h6��!`�+s�yH�"O$ȡ`�@<'U��d���'Fm�"OjL)!k3+6�쀡HY�C��ت��'���'���'nZ>�	柌�I6:w�M����i����?+�n��I���I����Ο��I͟4�I����ɨd%��7�J�s�2!{A
1sib �����������՟���ڟ����(���m����f�
��jQ�>[�\�������I���Iȟ���ϟ��������)4�HP
����0�h�Q��%AI(�����\����H�I럸�	ǟ��I矀���������T\�t���]�fW�a��˟�����矨��,����H�Ʌw1tc�bN��2�vM�[s�����p�	ϟ���Ο���ҟ��	���	(E��p�Ŧl��k��$DX����ß��I�� ��ڟ����T�I����1ް�M��>����r�,m��ޟL�I՟��	���	�`��ʟD�	�!a�((���n~��P��"'�Y�Iş�	֟4�I�@��T����p�Ɇ\�D�a�9I�z\�Œ3=�¬��џd�	۟,�	�������	��InpM���s��Yd,��S�Fu�	�d�Iܟ|��֟$�����	��\��0�:i��Iܲ bD�"�#o6���Iɟ���ڟ$�	ߟ��Iݟ���4�?���s1B)�� ů�X�B���I�d�S�l��wy���O4n!���``��X>�Q��G��qc��)?Y5�i8�O�9O8��E�DD�$1eiſ(��ck����O�\��`xӄ�����O;�e��X�"�|�P+�1��}��yB�'��	D�O�  !T�G�8I��p��׆%5��8#�e�:� �$9�S<�M�;r����$I �$��Hc���*� #��?�'��)�ӆ,x��m��<��Y�qVf���υV6��0�+��<y�'�^�d���hO��O�y�AJ4�kQ��L*��bB:O�˓��uV�&D ʘ'�h20,�F�@���B�����$�V}2�'��8O��"Ş!�O��j�D��Pr����'�reǒ	�X���tE�ҟ�A�'f3��ѩ$����B�λ
���Q��'��9Ot}��j�5���AK��(�`��0O��nZ�j�?���4�.�ˆ��"&�x ��/w���K�0O(���O��
#%�6m#?��O�P�	2\�\��DI�M��k��OT���M>y-O�I�Oh��Ob���O��A�eX2*JH�ɑ-�		���׫�<�Դi>��2�'v��'��$'[;.w�ɘ&�VH�KA&t����@��]�d�P�O���2�i>u��Ο�e��+F�� 	H��=I'�8���[��Ny�$��Z"a�'+��%���'h�Q��Yl��bm�6Y-�ak'�';r�'�2���TW�0;ܴq�(�;�(8x��e���Ū@g��(�E���U�Ɛ|�O��ꓪ?���?Q�>X���U,a�����ȟ.Pyfd�4���#_�|e��O��O���J������hϤ{���PЂ�yr�'�r�'`��'�����r�Qz�k� �"e��B=�4��Op��U��8�q>I�ɽ�M[M>�"$�A\�B��]2X9H2h�]̓�?I.O��KŬ{���-B��A`H
T#����!�'3A�P(֢S��������$�OZ���O�扅	PDE��^��i�'!�`��$�O�˓%,��ɗ(�r�'�W>5����$I0�P�@!=_����>?a7Z���I�D&��'�"��0�S�K�A3EC;�Ƭs�/)Ԑ��ڴ��i>����ON�O�h�6�4�2�� U��e0Th�O �$�O����O1�4˓ ��Fb�M�z��' e��x�
���d��X��@�4��'����?�E+["
ӚA�%ñrX�pRn̼�?��640R�4��D´NPR��'���w����Tꝩ�h9+s
��F^��IMy��'���'2�'��Y>�"g�N n�"$T,D>pL�Λ�g'ܴ�v�d�O0�$5�I�O�$lzޱ����p8\��� ��dY��)��@�?�|���9�MS�'�8%��i��1Z|a��9Y�z�'���c�W��ԙ�|U�D��럼�gSht�P��D��в�K矤��p�I`y2��)�Q��O���O\	�a�C�d����̫>`b51��5�I����O���-�J�Y��|�Df�LB,p���r����+�d:&�����|�d,��D�	�Z!���ɒq�*��r���%8���ǟ(�	ݟ\��j�O�Mԣc��p�W ��{<�����ۖ�ҫoӚXJeϧ<���i��O���^�0YI�·�C�:9�@��,��O<�$�O�9�2�~ӎ�MC�-����lQ���	5
�ŋ�ȡ$��a�����䓦�4���D�O��$�O��D�/uq"�Ѓl�|Z�@a��*��˓d(��E��{���'�����'����;S�[���oR�䫵��>���?�J>�|Q�@�  ����И�Di��tF��������$j�% ���O��2���x思�S� ��Z��p�����?I��?���|�.O�nZO;@��ɾx~F�VG�1s��A��ĹQf�����McN>���e��	����	��s��
����$�3F�<�zG����@n�V~r띋s����S�D#�O�� $u²(�$;�±*���Dn�5 >O0�D�O����O�d�O��?�S/Y&���#�Rc���NX��(�I۟�@ܴ�ϧ�?)5�i,�'��-�CT+ !��*V"��d�|�'��O<�x÷i��)a 1�%�+N0>ıĉ+���ϕ�ZF��\��@y�O���',"�$aFfQB@�Kpp���ᘩP!��'��ɉ�M�Չ�0�?1���?�(��8�d�� �,��F�M�@�zD��Hq�O��D�OғO�/������JNk�l��G�7nք���$UF�lZ���4���'�'4��1ů6&�}J%gD5BIŠ"�'���'�OE��M��ڠ>�f�)%��
&(H��D�^��	���?���i��On��'���29��Ъ�@��z�%D˱Mx��'�(E���is�iݹ���?��P�yPfM*GU�D�`�!�Hl��Gr���'Z��'T��'���'�S�/� }@f�a�8�pÕ|m�۴'X��y���?����O�|6=�����&V�  !T2�@F�O<�� ���b��6Mv���`c$T��hU��3T)�]��e�DB傈V�2�E��Ny�O��BA2�U��K[	!r��e��1�r�'�r�'��I�M��*��?���?1�GԦaY�$����K��-+�ş���'��ꓡ?������.�����=e��S#'?�o�;|ca(3�z�'{b�����?�5ȏ�A0��4�ы5��Q8�]�?���?����?��i�O���b�5ep�D�%aA�7><)��O��o�E�&8�'4�7M?�iށ��ΩK������ C�.t	��p����˟�I0b�	m�h~2�P�I���'p�B��,A6K}��&�l28�IM>�)OP���O��D�O��$�O��2�h�A1.A�m�e��5�Ƚ<iŷi�0���'���'���yc��d��7⋙2����r	��t��?�����S�'r�9�n�!Hՠm#�I�0@  S��"Q�'2� R� Ɵl��|bW����"]PT�P�ۺE���ƀΟd�I�����py�)bӾDXR�O���*4R�h7n���=�b9O�doZp��Z���؟������;fr`��͎�L�����#l.(n�z~R�_2�p(�[�'¿+25rZ��A/�?F��r#�Z�<���?i���?���?A��d�YJ:|1DJ���(����"�'�"Lm��DA�¶<3�i��'th��eό�+F��i��ƾFr�d��|��'�OUzH[2�i����f�C&�f*CƐ%�Zd�ĈL�L2i�a��ey�O��'��
KyA�x��K�B|hP�n�0���'��ɵ�M���ʼ�?q���?A/�R��r%�nG��e�ƥQ�)[a�����O��$!�)R��ʰd]a���s`��5��[7�&��x-O�	\�?a�<���@>��c��7�e
𢊆���d�O����O��	�<��iw�E`hq���d��o���؀,�D]����س޴��'2���?   !�ՈfO3+��Ԁ%o_�?��Ww���4���FE5��s�O��I� :D�`���t�-���r�IPy��'��'2�'rP>�"� �����QΙ����f��$�Mc����?9��?M~2�9ʛ�wa��'+ئ�b�:��M;?ɼt��'�r�|��D�L!
��8O��%��<`uNƸ  �X�A4O@XC ��~b�|�Q�\�	�`BQ�ɍ��ip��\&��9xã�� �Iӟ���Wy"#`�:�rDN�O����O�l9#�o�z��s�U�C�t�0J/��?��$�O��@�Ac��#o:�H¬���0C�+?y�D_�0[f�Rc&R#��7Yl��R��?����8NN}��Qv�ڠzO���?����?Q��?1����O^p��'X�;M���cǅE��黑E�O��oZ)/wz��I񟬫ڴ���y���;Ȳ��ƹ,"-�����y��'���'��1��i��i�E����?���вN�~(�U�\� 52��Ʈ�G�'1�I��X��џ(�����	�Z��H�#"ƭ��FO���T�'�6m��{���d�O>��7�9ORh�$H�iz�\˧n�����4��T}2�'�|���k�)�������l���ö�@);�1Q�.IfG�I��\����'3�9$���'=�r��U�54^PisF����]���'���'F"����_����4[ۨm���=N))��P��x�GJ�]�h�����V��d}��'{�w2��a�$[<k�:�(1a�
"�Ȭq�͗&�V���#Å�bu���Za����uؕl)~CxQ B�9*E�V�y���I̟��	ݟ4�	�����F�$ZI�)2隩���W��?Y���?�R�i��ȣ�O
� iӼ�OxɂX��q�a¯v4%�L��'S���$���R��擟����	-�P�BDg��{�-	���?����"�O�Of��?i���?��x7�r�.J�0;�ol�D ��?!)O�Un?r���'l�]>EۦFS�mdz8#Q���'�ޠp��)?Q�R���IT�S���ёz�5����aҩ�!'��iy�(N=g](���L�$��4����HRS�	�Dh��#��Ei��aѯ�"wg�����x�'����R�x+ݴYt�kc�D>/kB����[�nD(��>�?�������$�c}2�'
&�yG!�	KEnX"A�(i�ȣ�'�'�*6}�&��t�1��[�d�~� ��I�nNP�L���+E�f�R�5O�ʓ�?����?����?)����6U?�4� l��Й2΂�5ݾ�o.1l�Iݟh��x��ݟH���s �Y. zb}٥P�X���	�?����ŞT3Njڴ�y���`Ą#Y�\a3�]�^�\̓FL@1��H�OΕ�H>�-O�i�O��bP�ϖ� ���+�<� a�On���O���<ip�i�J����'Kr�'�D1�䛣)�V�� Dn�� s�Ds}�'�"�|�#���1��h�A8�[cM���$� �$���t�J�%?	" �O|��щbz��E"�Q��`Kݼ�\���O2���O���9�'�?�a��8U0�a�R��vs%�S��?I��i�&]��P���ڴ���yׅ��b<�zi�V�T�Jѝ�y��'��'�4�x��i�i�q��?�(��O�hH�.!Fl�� ���99�'�	Ο������	�T�I�2!��¶$Y���cĈ�61@���'w 6M�Dݼ�D�OB�)�i�OL<���*]1�Eم��C�T��D�q}2�'��O1��;�'D:T0��u��x�,@�1�F�VB��k5�<� %�(�P��8�䓟�Ĕm�vds�`�&�H�)ŨB�t�f�d�OL�$�O��4�XʓE^���l��f�>b�`�H���~�������yr%g���L��O���O��D�&D�<ZQ�̘<}���2��=�|t�"Nn��O�V43���B�>���MW|���F.���
'l��h'j�I���	�����Ɵ���J��cLH�"4A%
TQ����ߦ�����c�4e���Χ�?1²i��'�0� ㏓�FT�$�� �>Y�ğ|��'��Om���s�i���?�$D�w������r� �هbN�{���$���<)��?A���?1�͠��"6��\J���"�?	���d٦�³FP�� ��͟��O}L�`χ_h�dҠ�R=6�l��OX�'T��'�ɧ�	��rS.i���K�n/�X�T�צCodX�5e��2QV��Ư�<ͧ&����?��I���dD jv� �
8�X����?A���?I�Ş��G٦��$G��V�={�\6_�<��j͕"v�����X�ݴ��'�|��?y�
ޱ��ܱ6.C�&E�$����d��L�6M ?�ѫ�n�8��R���dɏ
���x�tsN7 @pI͓����O����OT���O����|��^�g�����s���J`k�5Q=�N��R�'���'�~7=�IZ�![�x�jQ����2Q�\u{ n�O���6����	��7-f�,���ٚ3��p�F=��C���$�%a�@ ��6t��O���?��P�`� ׻E>�H���A<������?Y���?�.O>xmڧ1�V�����D�I8|�1p���k�(	�o_��*��?	#Q�0���%�!�x8�dZ�a�m�6�1p$?ٴ&Ș^�b��`�ϼ��'U�l���<�?!���V�hj�������7���?���?���?��	�O� �G�/L��K�e�[`(��M�O&Mn�n���'��72�i�a �h�-����Uig8�QR�w�0��ʟ����M�x�mR~�C�f����M!�-�' ɔ5�<S�O���e[�|�_��ȟ��I����I���� ��&�x�0+ҨM����ƩTMyg���"O�Oh���O��|���x3N� ��Zr�`8�>8��}�'�"�'rɧ�O�\�� ,��:Űq(g�0_�8�p�E�Pzb@3�X�tiCeC4V��q��ty¡_4i�4@�2�Lb� ˀ�>"2�'��'��O���MӲ�F�?��e���)7O�<\_��	`�M��?)�i��O��'X^�h��*[&��� �E[�δ{P��1�F�mZI~��������7{u�O���?�n��v�KR���1NȽ�y"�'���'���'�����0{�xpSH��@�\KQ��)?}R���O�����ԇo>�����M�I>91��9�&��s�טUs8�cr�����?a��|����M��O��(���I�҃Q8X�4S��(R��U���z�IQy��'vR�'a�c�G2���.�?�&D�үM4ob�'��ɱ�M������?���?�/�t)rk\2&���Hu�	�}��tJS����On�D�OO��<Fql�(��?*��F'�C�L�c�ƙpY8�oZ���4����'��'ݔ�#�䜞y��p%���pܑ�'2�'c���O.��9�M{p�� b�8�@ԟX�T[g��#XDL���?�i��Ot	�'��(�����Ҟ.���zadj�'پ�P�i�	<}�>������j��Ǽ.dL�c7l�%'I��<9��"hb٪��?A��?���|z�̊�/՞����O�v�$be���֊�uj��'���Ou���'�n��N��_F�yѬ���L���
�,.����Oj�O��O�$�Eq�7������* v�q����#߸Hb*e�� �[
�R�KA��Ty�O��2DH�82è�|w�$3�ɚ��b�'���'��	��MC�I>��D�O� 9�$M��SF�ThlT�� (��<���OJ��5�$X�}�E�+���Ʀ0j �I�b�"�:7m>擮)w��O8@b��7�(@��$NE���$O�OZ���ON�$�O��}J�*Ia� NF�D����cb!I�i%�F�_�"�R�'�>6�:�i�q�R�L�E�.,4�H����a��������8N�Lxl�m~Zw�꽳e�O?�� ���'o։yf���N�TD���	0�Ĥ<	��?i���?	��?��[\C�=�Cc�3DS�(��点���	Ʀa�Ce	ݟ��I��%?����N�����h�Lp�d�C3����O0���O��O1�D]3G-�(��q���|�8�0���kV�ےC�<��|y��$J�����D�1,4����4z�f�᭔!Q/b���Of��Od�4�V�雦��)�r�C�g,�Er�J�� Q���1+�\V2�|�^㟜`�O"�d�<A���.*7�}��F��6�8k��)QȪ���4���	�4�Dd��'rߴ��Z��S����WN�:��P($�X���O����O����Ol��!��/�[L�>Q�آc#֏(]�d�'�Rk�n��G4���$ݦ1&���ª�"�CC��)F�� %�H���t�i>-� �ߦ��'*�`�1��;���#��L;Cv`��i�Z=Z��r�~�OX��|J���?��%�j@"���C���a��̓_�6E"���?I.O
�n�Qy"��'��[>��C.�>$F�p��A.^`��7�o���������O�$6��?`A��_�)k�F�w ���FH 4���ƌ�ݦ�k*O��G4�~B�|�\�b��A+!�j�`��r�c��'��'`���X��Y�43Ū!k���Vbũ�A*6���)S2�?i��^��$�F}��'B���
�
�4h0@đB���� �'�ïf��H�B�$	���<y�lG"1ҭ봀ξ^X��t�H�<q)Ox�D�Op�d�O��$�O��'�Hh	�*��<X}2o_|8� ��i�&��W����C��П�������DڿLAR�J��6V��cp`��?�����S�',��a#ܴ�y"j�������R�2�����y�`�:��M�����4�6��>*� .������7� �f@����O.���O��o�� ш_K��ڟ�e�1YI����*�c�K��������џ��?i3-$U�"� K[3. �Ek���U~b�f��|G�$B%�O��h�I%Bl�ݦEAr% U��c��A�u	7;�B�'��'S�����#��E-U�Tmy��v#�
 ��� 2ܴA��.O^4l�c�Ӽ;V��,�v<s��-S���@��<���?�k�8i�4���7Td�8x��#V�P��9G��=�K�HBJm�VD%��<�'�?Q��?���?�qޅv�`�yAM_.Y�J	��B�����jXƟ������$?��	�HNP����*)AJ7�T?&����O�&�)����:�g�9�D����~�tO��cй�'9 0�������Aw�|�T�P "�pN(zv�.}��*��͟��I矌�I��Ny�n�Ѡ��O���.�:ap��4�J�9��@�S*�OB�o�o��r��I����IП����]2q��$8�GX2ʨ��2�Q�5��me~��%Gf���oܧ��d��0#�r0o��ھ�Ab)��<Y���?	���?���?���T�[(����!-0ƍ�	%���'�b�yӂ�ڱ�?i��4��u� :V��; $�����F�AO>����?�'e����4���� B%�0�4����!�JPP��S���������O����Ox�Ę�3�;�OI�M�T�K@ ��D�OʓT���Gg�ɟ��Od���C��G�x�*�`Py� 8K�'����>A��?�N>�O&�x����Y"r%��A�x�$�b�gB��l$a��i�.��|�t���x'���fiP���hF�N���)�⟨�I���	��b>y�'��7m�}�U�3�U=tp�Z�ѯ&���b�g�O^��^��?��Z�����D�2�z�����3Ј�`����I!Z4�}n�n~��]�aJ��}�uHL"T0K�pP�95�L�<	)O���O��$�O|���O�˧�� �mG�-�ݸB�KP�&�Hn<W� a��՟8��N�'#d��w@92���{i��Å�
+U�=��'�|��+��Vc��:O�E!Aʙ4�@�w���A�n�@�<O��YFL��?I��6���<�'�?i�S>\����I�B�jȫ�?A��?����D�ĦA����I����B:}V�\�S��>��D�5ʞn��
��I�\��W��B*0Hs��٢V�ы���3,�|�E��q3@��/X��|ZP(�O���Q ��h��>?�ޙ	�d��u�:�*���?����?a��h�@�ę�Ŷ��,~R�(U��Z���Ħa�Oky��m����].`$���U'Ç_���eſxچ��ȟ|�'?�1��i��	�^ Pԛ��O!����֐BtL(��`���4�iV�IK�	wy��'Zb�'�B�'5���|�~@�M2b:���r�����9�M������?���?�N~ΓL�P:1��8,�"��-[SG
(�WT�`�I���&�b>�H�f]�m�!�.O�(q�:NH|�`�ض�+?t�5�v�$���䓴��(v*����蒜R}�š��_0<v�$�O����On�4���s]�v��'�ƘH�xP�w�ӀF3��c��y�f����O����Ot��SYl�D���o�(�4k�)��cCdӎ�0df���>���7�qX�h_�4L&�� $�Iǟ���� ��֟�Is��H��d�a.T`��C�n-�XU����?)��(ƛf$�+j��	��M�J>���R��*�Ⲃ��L�N�Ҥ�4���?���|r�޴�MK�O��YE�? ��t#MH�H$`e�
3wh�`J]��?�$�-�d�<a���?���?�5��B�(��u��,~n.��*�$�?�����$U�!�C�����	��h�O���g��=|񰄉�5榁C�O���'�2�'�ɧ�i�/W��XǗ:]F� #��5C�0�pE �m%P6�My�O|����b���R$��PNxd��Ō�'R����?���?��Ş��ğ䦵�E-^*& "̃a���	�L�<N�I�����Z�4��'u�듀?� ���Y>�YP��B�<ٛ�ݭ�?���V�z��ش��D��x�����e	�@CjDIvY�� 02��T7�yT���	�L�	ޟ �����O1��������<�l\4}
��u� �f�O���Ov������?���JB�צ4H��M�v������$�b>� �MD�a�y�Qh��
b���˛�@P�̓m�q����O�iAH>�(O�i�O��U�ܳ����%cO�&�3F �O\���O���<�4�i:D����'���'����,���#��n��pP���S}�'l��|��:"i� D�:-G&X#1�M.��d��bZ���Bs��c>H1�O����~��5�ťZ�`Gl� @��,s����O��$�OH�:ڧ�?Ɂ$ �U�D#"�^ �t��ƴ�?���i�� ���'��/h�z��]�mg��pREu9h����2qB�ٟ`�I˟�Xw'���',hy���L�?��R!!��1 �% >H���CL�'?�i>=�I��I��,�I�v�x|8�(J.5�=�a$U8��'��6�Qeq*ʓ�?�M~r�bRI�b�D�T����k��We�%��V�\�Iş�&�b>ɢ�'�;{�� ;��C$G u飦�O�`m%��KE0|*�'��'則-]�x��C�e��+��Dd0��I�h���l�i>��'�6mU:��ɒ
Ǽ=�t��98S��f�1���$���?��\��	���I�Dd��S��s�f$�3안+�=8��'#6�&�Q�O�KF�9e��{��3A)
��1�yB�']��'���'V����')�&�1'G�'"nޱd�Ԗs}���O������X��o>I����M�N>��F�RS��
�
ޜ^^y9�㚘�䓎?9��|� f�"�M�O�a!P��S�vxH$$�bV�qW�L)�����AB`�O���|���?i������Z�7�����8��TJ���?)O��nZyhjE�	ȟ\��]�ă�=@�(!*`�
Z��<�+���D�W}�'�B�|ʟ>)z�B@��4=)�DÒT5j=if���*+x�I'�������|b���OJd�H>Yh ��Q �O	Z�ΥxM��?i���?1��?�|�,O��nZ�>�j���� :o��t ���;J!x4ò�V^yB-a���@ �O��DW?�F����{�^�Q��S|t�$�O�p8�v���Ӻ[�%���Q�<�#��(�1 �P���pP�<�*OL�D�Od���O��D�OZ�'�5 1��]h�1�t`�=;�`���i�dс�'���'��y"�~��7)�������U��q�h��n�
�D�O�O1�f̑lg���/|�~�ٲm�w����jOz�R�ɜ-��y�'��@$����4�'�a  F��`�Ʃ��.Y��(0�'|R�'BW�qܴR.Zq#��?y��I�� ӂ�R�k��Ց�J*� �ی�m�>����?�I>a�a[�k�\S`�L�$!k�k�C~���.��P�`W�O����nMb�A\���
� X]h3O��l���'���'�"����ؙs�*����#��&`����Sߟ���4~ML����?���i%�O����x4��ꪉ`wZ�Um��O����OD���w��n"�����?i��Օq�p�7-*t�
���
�V�Ijy�OJ��'���'G�E>q���Y6AR"+FUР���X�I
�M#�/ˆ�?����?���4��v�Y �$req��$Z���?���S�'Q#-X�G�U���B!l¨Q�A"�a,�M[0^��ʕ��D5��<�C�ݢ)�hI�6(G�w@D���ڑ�?I���?��G�R�������֦rҌ��	�!Rĸ0� T���#)��+$T���M�I>������џ��'ʰ�����/�p[F��Z��{g �>N��8O�z�i���'_�˓�B��Uj2��e	����ҨV?��	��?����?����?���O�DY����*���1��q��%�'9�'}@6M�q��˓����|�R
<���!�߱cА�1f�ј'P2^��RbDѦQ�'� }�3� ~H��z�JYFx� �8(��	�7��')������I̟�ɀL��bJ�c���p���(�ԟ0��Ay"irӔK� �O ���OZ˧7���pF�ӂa���F*Yw��'f��?y���S����W^f��@K� Uf4��0JI����Wt�9 �iy\��|�G���%�du-�.�l̫Ҏ@�q�6D��ȟ������I�b>��'#7M�=���u�![�Jq��oªz��i� �<iS�i�ORq�'r�E*Dmh�猼_����ٮG��'�ʤ�F�i����CKڥ1s�O��'n�n1рh�l���Qk�>sn8=Γ���OL���O���O����|BJ�E��-SR�����A�*�)�����%eHr�'�B���'lB7=����R�T��1�"cP9�'�O��d!��U
f 6-u�� (��^��@|��Aӣt$���t7O�U���?G�:���<ͧ�?q��֙:����E6��x2���?����?����˦�	��Eȟ���ş�����0
"	ބ� 42f�J��$���柰��E�I�=-�H�E�@dʶ�T�B=����4mCd��Jz��|�t�O���DrH<�ˆ�$���NT
H�P����?���?i���h�����
J&л�M����2�䁂z�
��������Rٟ4��2�MK��wh�Xq�i֊q�(2u�ߵ!�Ԭ	�';�S�<������'���R��?Mq�L�1MK�@'L�}�n����H	$��'��I�T�����	��l�	����t���	a�WJ�'06�}�t��?QI~r��$MptK�m��Jki��bn��GT���I۟'�b>��1,X�Q�zO��{��� K�&��m��dx��4Y�'��'F�I9��8;w�*]bn�q �!63�������ӟ\�i>��'uD6퉍?�����MY^��t�ȴt�|z��������Φ	�?%S����ן�9K�¼��`F�=+���'�W�L%h@����'	^2%��f�M~:�;,��	� B�õ)�!VHΓ�?A��?q��?���O���I�4[�(k��B�JJfyR��'�r�'wp6MZ:i+���O>9m�\��G��͢�a*4Җ�j�'�t���$�8�����|��lF~bÑ�v�X�c�n��
լ��R��$5��UR�Ez?�L>�-O:�D�O����O�]٣b
�'�:\��̌m0��p"�O���<��iAN\[qV���	@���J��(���hz �(F�����Mu}B�'�r�|ʟK��#�F�p�@��Ji�5˃��Xx:bC;��xc�O�	��?�Ƭ>���]E�de՛-^�$l܏D|���I䟸��ğ��)�By��o��qz�II�gs��/�h���J p�����O���_ئ9�?��V���	�^aM�D.�(pBt!:pdԗE����Iğ��
�ɦ��'8��a+�Q�(O�����<)�W,��8�{P:Op��?���?����?����5F�|�A��X�Th��6,-mZ90�
��'U����'��7=��-���"=ހ�pi�H%"�K0`�O��,��)��{B6z��ؗK7H|s��>&����k��q#��W;�0��<�O�$���b�x�T��5f���	Ó
7�F/��I��0+@A�_�1���N�	�P��%�s�3�	ݟ0��M�Ʌ� ��5j\>XxH��f�'%��}������ON^��J~r�l�OJ���i����"h؃Y)f81�/V�D��P�ޑ�7
��S�����U
��b�b��vB,P�	��Mk��w/�E�t��`l�{k���ĸ�'GR�'�R�ӆ��֔��Z�� �<5���.c)
l�dj��w��r�8l���O����O��������2����68��������4[�x��+O �"���D��̒֫�+ (|sd�M ���O����O�O1�@��c�G���I H��%��.S�7�RKyR��?)_t���䓭�D\��A`�� ꀉ#b��a|��y�lDY���O�l!R�%g�0$����^r�Q�6O�yn�F����	ޟ���ҟx�1��qc4�IS��	z��j��?lb��mZr~R���'
p��S#�O'�(0� ���+�#Y^p�a����yb�'�`Qs��^�$L��־NH��]� ��;�Ms�O�_���`�ΓO*�����&+p��"p͘� ���6�"���O�4��a�~��
�4y��(�N!��JEN_4g���2�Ib��9�eR1K���EO^B�xU���}GedhS�Hؼ�P��B�I�@2�W���U*R��&�n1 ���_�ո�W6�^!SPJ��ejʄ0�0э�D0]����W�S�����$�k6	���J
�.30�Y�:^�0ya䑵V����m�5	?�5ɢ��zf��D��N$�xDJ�*j$ ����)�|��Ì�}��\C�N&'��,�s��1&�x9�L�0^|�����?'�@��"�	�t����F�G�6��U6�d(�!o� NنȷK33ƪ�`gB��K���'�r�'���Eތ��"l�9hN^���N�>BLO����O���b�1�	C�F�\" �fQ����?3*T�Zu+����'}�xRq/u���D�Od���~�֧5���5g%hE	LT}��U{Tȅ��M���?��O���'Vq�^ZW�A�lL�kp�}�$��!�ik:�k��iӄ���Oj�d럮1�'�剶RU���b����1��;WX���ݴm+��Ӌr���O6x�G � [�jBjL�rl�x��覹�I쟈���N��X�Oh˓�?��'����˹1FUy���:x�@ћ�}��Q�@��'eR�'��'7%:���224����c9P7��O�؁A��_}�S����w�i���Dm�F͢�ۃO���	�/�>y��Ѓ�?1+O��$�O���<!3��4V�]	�ԁ&^�8a䫔�.M#Z� �'�r�|��'�b/M	}'Ȋ�
��J�ӥϕ�!��(1G�|��'���'��"�0�O�j���gK/x���c�J����z�4����O��Ox���O2�+�[�8�e��BuFL� A�)|��Yef�>)���?�����ئ5��Ocr��^���3�Ȯm���"��=i�7M�O �O��d�OzMrG-�p���T痾&�np�'h�0>�
6��O��Ľ<�K8*������	�?q�� z��!@Iv�B�bҗO �8"��x��'�LE�{=��|rԟD�v�T�PH�dp�/�?o�r���i��!	�xߴ�?���?���g��i�-� l�)�pA劚�	�QӢwӆ�d�O��#��#�Ik�'ug���S���aI�0c2D�D��nD�
|�ٴ�?����?!��2��|yRƱtzB@��Y#q��ј"��	8x�6�X�� ���B��!�ؑ����ZC��D���e��iH��'����L�f����Or�	�G_�[2K7Z/���uKևOFFb�|�w�YQ��ǟ���ߟx1'�z���D.�x�8G�*�M+�X!�a��R���'12�|Zc��|@���"�ΡQE�7vºӪO�����5���O����O�˓W��pX�K�Q\���#����#�-�a��IoyR�'��'B�'� ��>�|���I?��Z�eE�13�'>�',"Z�|�PeA-���O]7"l �p���Z�P�2����$�O��$4��<�'�?���غ1�šU�Ο�����`_~���P����d�'��(���7��C�m�ͻUęE��}'���b�`lZ�4'�Ĕ����'(�'d���Ъ� 
PMz	�/.�zyoϟ�Ijy�ɒK��"����kX�2E���B%�#+��qC��Z7}ʉ'W�I��$��\�s���?�"EhaG�d�g ùs��6-�<�߾Q��̪~���Z����3 �)A��R�C3\t�-J�Ji���?��@J�O���M#'٨ΰР���,�+ae��[��Y��M[���?	���C�x�O�F!�P�]Ƅ 3@-��ؽ�`�q�,��O���1��?�	��y��
.D���{G�(��iY�MK��?)�u=�,�U�x�O���O�	:�
T�x(�� �*ID�8�i�|��~�'��O@؀gm�j����=~0�i���K�w��	����!�I<kO����*15.%�B@�'i��J<��j_q̓�?�)O��DF5�����HU�b����t%hEɓ�<Y���?��b�'��$��
��E*�HƵ�A�b��7�����'\Z���I!/}��'vS,���79�H\Y�Ξ!�Ql�ğ��IY��?!+O,����i� �av��"d��y��(
�88�O�d�O0�Ĩ<Y��0[P�Or�UK��M'+a�\3���Y�u� �{���D,�d�<ͧ�?�K?}����Ҁb��[�xzf�l� ���O�˓S-��7���'��\cf�]��Iqc�d�T'R#'�hK<�.O�d�O����'�_��R�ɇG `�U���ɫg���	ן���̟���oyZw�����)[<z����Y�4h@ڴ�?)-O�0�S�)��7$(�$�֢%vıp�٦E;����$\6��O^�D�O�)^K�i>%AD��OE@hx*B.7u�̹
�M���?����S��'y���;o���⨌4���h䕜o37��O�D�O@�c�m�c�i>��	v?���^_�t��G�_N H�όƦ}��n�������	G?y�$�2c~�Yn#4T���΂Ħ���	c�i�'$�'��'�,x��(�WHt\��дF���hZ\�'q����O�$�OR�d�<aiE�G�"`��e�?$h�-��C�8N��;S�x��'1B�|�]��ݞ5g ��u/�%�|��J�U��7-�O�˓�?����?�.O�ax�J��|b��Y2{N!���Zj� "(Tv}R�'|b�|BZ���㟈K&O_�[��(��	^L\H������d�O����OF�]�6Y�Q?��	�[K2�yDJ�*��Tج�{���M��jyr�'�"�'j��	�'^��'v=�1�2F,�@��J��1sg&�����O�˓Wߒ���Q?��	����0,��*��p��DJ�,�i�Ҡ�OL��O�$�?r��|Γ��4̘#S)X �`(8������.�M{,O�X���\즩����I�?y��O��#�L��@�����R��զ��	П$������zy���׺p��U�『�CL��`��؋b���S5j�6��O���Op��C}�\�d�ŏZ�w�h� �2ox2���.Đ�M#@L��<I�����,��ޟ ygi�\�2ɱ��lOR�B�G0�M���?I�*v��ȱ^�ȕ'5��Or�*$Eʸ<u����Я|��i��W����Ov��?���?!$�D�V����&M�8S�* y�+V�/����'J���%�>�*OV���<����i��@�s֧ [���z�&�h}��t?�/O�D�OL�����#%SW"Phy�_0�S%��<S�x�'�џȕ'��'G��߭[��$�UgEbw�P9�m\1H�"qП'wb�'���'�bW��(6,���Ċ��X�BlJ�Q�>�v��M�.O���<���?��g�܁�h�4�EÌ �D�� X�#P�W�����T�IpyB�G(8��?	EC6�S$��� c��H�s��v�'��I˟���ٟ4js���	��8���#J{�1���M�N�
�ZcL޷�M����?a,O:u+Q��e�t�'�R�O�(I�Bmߤ�8�`�!֭,����Ʃ>���?��q��P�'��[2����K~R���ߩa�a�5�Ϧq�'7{�cs�r���OP�����a֧u�O�U�$Ft�� j��7��O��d>!�D=�D"�S++a@��c�F���̀"jL7�!x]��m՟H��ڟ��S���D�<�� ĨR�� !S���%�^S� �iM����'�[�$����pR�[��8�f`⒇�4$|�`�a�ii"�']�M˙,�j���$�O����s�b��,F�f�,	CPbPn%�6m�O��%�<�S��'b�'�bKM7!��h�aP�n1�1�kӠ�D�*,��'���ޟȗ'�Zc�!;�-إ{^uS��z��� �OX�{�<O2��O����O2��<���-8��)�r�-�@��db���ġ<������O��$�OؘIS��v�(�r�ԏ4�(��Ӫ�u���OL�d�O�d�O�AG�*�6��A��E���0��ۃ1Nν�Զi`�����'a��'��#����	ϩE�H�J#F�[9�(��;��ԟt��ßܔ'�E��E�~��E��H�m
��%��L� -�8��i�BQ� �	՟$�I�V��IA��|b�$�Q�@j'f� ̐uJ�F�'R]�8�v!���'�?q�'tb<�ql҉+ȡ����:kQ�I�xR�'�B׀59�|�П R+�4L�bÀ�1Z�$k��iE�I�J�b��ڴZO�S��������W\z�y�ݽ<.�Bu/��gg���'�B'M�O��>�#,
H�^@Rs�%W�A`�k����˦��	ß�I�?={�}B,��F  M���V����͖�O��6�T
���3�$ ��ៀ�dI��@�L�KfiI�`3 %Ƒ�M{��?	��v����xB�'y��O�y:t�S8�9s��\Y"$��i��'�ެ�	,�i�O��D�Oݰ)ԛ>�f8�%<_��A1�Ԧ��ɼiK����}"�'�ɧ5&�_F��0y����֣�3��D��]�<A���?�����y1z�#ۑ0�LQE��r?~I��d(��c���It�ϟ��	�k��(q-ӊ+���'^�,�|�X�g���'���'�R�!F�0��d&W#����K��w��I���'��$�O�d�<a��?Q�>Pt��E
䪰bņ�*#@��\���UU���ӟ�	lyB�*^��(l�����Ҷ�7NUس�,�ۦ�	P�	�� �ɌC���@��Ap-~m�D�e�i�nG�l����4�?Y����Ḏ2�$>����?�k�"�+P�\((a���["h�A��	�ē�?���-=8Γ�䓒�4B������`�b�U�ֹ�M�+O
�K������������'�x7��I=P��ǿQ;x� ۴�?)��eKT̓����O\�a�1�F& @���1#H5��xH�43uܠ1�iG��'��ÒO>���c�V�aeK�����ʓ{�Hnڨym�e��q�J�'�?q`��9���c�$:��T'-$t�F�'���'�hP��.�������m[�5���u��T`"���L��Hl�@�	�f�<��H|���?���;��0�H;XI3�O��-��}9��i�CO�i��O �d�O^�Okl�>P��]xb��0�Pd�EI��;���.b0���myb�'���'��	6{K��A/�X
S)�A{�y��>�ē�?����?�s�� t�%O:�x�^n}��؜M����fy��'I"�'���'[v�mO*RD�Q�Ӫ��,2ҋ���q�O\�D�O��O^�d�O�4�T��O�Ĩ2��s��%r��H;��1 F�`}��'x��'c�ɚtC2�rI|j #�B3��J$� K3�Lp>T�V�'��'}B�'s0��S��V��pa� �46�Z8JV�V'����'��V�$CV/Q�ħ�?I��^����d�1�93�ϩb��t ��x"�'�R놁�yr�|֟>	�%�T�s�����ǂ�t�;a�i��<Q��ߴ��͟H�S��$T�3邵+�N�R�$��hK��f�'���4e_��|2��QYƄi`ʫkD�*Eƀ@l�v&�0�*6��OH�$�O��i�E�i>Y��j�q	�(�DÙ0�>�h�bT&����O��b>i�ɱq}FP@7�,(8*l�I�yg�(��4�?���?	��?�J~��~Z/��9���Ԭ!@�K*̄4ʜ��d�f�Sߟ��	��0zW%��.���Z�Ix�Aq��M���h)L]��x��'�"�|Zc:0X���ҎK��L�#/[��h���O�m�d�O����O��Cr���G�ϰ^��u�è��_
���$S
�'��'�'��']ʰ*��"���!e=0[sJ����'sb]�dA��̢}Z���@x�Q�#��V8�A�5�JL�<�5%��b
�����~�� �OH�J�؀焬-��83��Քgi����dv�zB�Hl�A��$;s+�%ؔ#X�c��taF��'RZ���Z�{UZ��u�G
X����a"!OSx�$W�W�@� ���W���H�V��a�v��?20��e�݈jtX��0hY!eX�E26D̀g�4�i���3�jͱ�%"h��L�	z�B��3'�>a�J��E״K�rA��🨓)�'74��G�^M�B��0�ޠV��I�|.��p�%�O�X�����6h��Oı��훳$��g� .� 0��͛�ڦ����!Nl֝�G�©ŉ��|,���ф_�N���'�^4���?a��	�ODh�@��.y�R�p��ѣN��"O4�g�;U�T�aF��Q׺�2��'h&"=YD/Z�2�*�@��&���4oռDu���',b�'&*�7���|o��'-b�y�\+m�����͝ %0�G-�y�1O����'�́I2,S�$�\���	B��8Q�{�	:��<� (ze�Z�_KJj2�t�*�$�3�ɒv�"���|�D�O��L�T�n�t8��ڬ�y��ە(�2�#Κ˨�͟���CJ���Xd3�c]�r`j�0Q7�HI��X<`7��� ��O\��O��D]ٺ���?�O�^7a��a�$�^F�j����D|:ə���/%��',�h��ý!Al]	Dۡs^�]b�'�82�\cq��R l�K��'�\+�,���q��.u�~��Ƥ¼�?1���hOx#<V�ϔy0F�zg�1%���PK*D��$5{\�`1��S@&p��#��)��ļ<����Rٛv�'��)�+z��,�צ��~G����V��'������'6r<�*���'M�'�,����,ZP���w���rH�I�	�,ܰ��?!��;l���Z�5`;
]��FF8�"���O��O\)�0�	��-��+� �"O�����R�k"��'���FO
=oڑ<���(�OG>y�$��ǀ�nc�@�����Mc��?-�LqRs��Ofy���F42��ؖGV�8���V+�O���Z��D0�|�'�~qxaըL����$�v�[L�TPGa%�S�',ZbA	PG̹h���P �;!J4�O��)��'G1O�1�� .r�Xx��o��cu.��"O���dZ5YK<e���}�鳄�',T"=ѳ@S�U����!l�S%d�ӅA�.<���'��'���'hW�>�"�'��y�AY�j�0�
�;+���D�O21Ov4��'Ɏ�S���F$X�f�ͣO�x�ۈ{��<��<�&b�dh�tI���81QX,f���'VP,1�S�g�+��l��F�f��	j����7�$B�I�:���) @�Q����K�1��X]��"|B'N��*��Y(���2pZNt��%�<P00zU��?����?���+5���O���i>�9��)F�X�E]5v�~(
ud�vB�I2*�A�nO�U���,!/N��<�ˆ�X�^@Y)���?�B���gC�2����1�OZ��
�0��!�1&ˈ|B\�"O�X ���;�� b��Sh�YH��di�J��V�i�"�'�r$�!APU9�x�D�,"6�� t�'�^�.K��'��c���|A�*[��86�G,P��3�@�p<�d�m��}���1�iW!����� �*�9��I�_q��.��6e+�h��/D�QZ�d�.�!�ĉ f�)[��σ%P�����Q!�$V�-!C;l�.�épg\��$�(D�8�ks��2E�X<a\T��s"D�����	��2���!�1{p
 D��j1�%kl�yX��}�U�un2D��+�D	\�<��v�
�&��	��,D��!f��D݀�9��I�:�(�r�l D��は�8���J�B�U<�
�)D���d	'v�65����d�C� (D��+ �X���H9`%�6*�؅�%D��)1,�u8����@7H"`�S�!D�ؑ��+j{v���(��0�⽀��;D�pK7@ߗ1?�h(�H�{vD��I;D��w�J�W^@���I�7&2)
@�:D�Ġ�	�<�8��.B�c<�\���4D�,���!n?♈3n���@�P��3D��چk��w�:1���܏$�4T���1D�LP�'Ģ}�8�*�-�R��j��+D��Ѕ� q&������&��9�#>D�dqO�a~RL�E(I;OH$,��k<D����O'Hv���f�ڋf4� %�:D���d�Gc���-T�5�R1�6D�Ѓ��ų��d 0!T/-eT��%�'D��k7�׫XǶ4i� 7����I+D��*�j�X��Pr/�z�ڈ���>D��P�}e�]��)�^�f�1�=D�,�b��9(��X�J��xi��!:D��d�vZl� �(W$�ʹ�c�6D�� VmYa��VVh�ak�B�l�)�"O@��&�\R
NI1�㊇HА��'��E��bL�T�XK�Y�Y32�)�'��D� ��(7	B�V#���
�'��٫#?;j���pb��E�	�'��� w�8�0n��-��e*�'�(�a����\�"���ې��'��M��A;2W�8�C�Z��ɓ�'�����ʀv��|���q�r���'���(6@��*� �"�a�P$
�'e��\�6.��"�;'s�t�' ��	�FB�{O�u*�Hq��pP�'����)�$l��������,h�'�j���'�8?�Xy�gW��4y�'�p(��ޞCSf�v��,��'�!
뒝s�ݒp
���"�'��zM��3�0ys�ix�B�y2,�3=Jvu��C�t�lL���ƭ�y"�]�4jH0t���rv~�K�#,�y"��:J0-�R�U�@�Z�vK���ybb��m[uJ�=f ���֭��y��"FGz��և5�(Df��7�y�fE�j0z-b*�4CT��Մ��y� �[�4\p�T83�j�rEg�y���*[���j["&���Ǧ���yb� 8dY�P��}�f��ɟ��yb�Ӗ6�yz���f���[��Z�y�R	v�Lq���@^%��qr���y�耀YY�H1�k�$F�݁�ǂ�y�O�Hb>�*��H9Tø�
 ʗ�yb��5u��V�J Hlb��V��y�	C�Q�l�;�Ɯ�V���s��>�y�B�"Tk^�8��$��q@Ci	-�y2J�*��h�0��1Ǵ��R���ybk�(7����2lۢ�Y��yJ��	�>�9Q'!yπ��2��.�y@�/#HHX�B��pO�4���?�y"�P��� �;*��C�͞��y��HZ\�Pp'��16ȃ��-�p=	ec<扻=���U�NBq��Qu�R�<�HC�I���kլ76�.}c�m��g�L➰�2A5�S�S1W��m@Ӣ�v�L�
�/O	4�HB�	�U4�1�@@((&(àZp!�?AD�B����	bf�*�|���JP�!�dD�U���!�R�7c�ػ�Ğ�K�F�Y��?| �z7�'��x����~r�ئ
7�l��h�,@�H�@�d���{0i 8�$h"V�۟�IqڤGh�E˒�2gD(�3&'�T��L�=��>Y6N�W���d-F1dɂ�Q䡓h�I$I��S੃�%c�=�L~d������	<B�<�q��Xp޹	WkH���C��'v�}rFĺb���a��U��9�v�B�D�)�Y86 ��Q�k$�x�bL���N���i޹Pt��8P�U�&��,��p{a� $��"b'U?}��9BRJ����qX�(�'����T?	z�I�1��*d/E=W�����p�����0�q��W`���^�C�&�0�Z�=��  ��%�~@)t�
���MQ1������Q׺|��j�7V��p��l�=LMt�L<)V�YO{ܱȢL����YS�Y}�A����
�:E
5I�a�Vٔ扨A�:�ѠX�dF�@���c�b�i̦k�KHC� ��Ԅ�A�
��0n�}ay
ʨ5:�U���!�������� ��X�I�{�*���'��xҘU�T���m?�O(�i�D�>f7�-kr�ݪ%�����*�O�i�`"@��	z�jK�R�IF��$f���䐰7�6�(Rȟ�AH?mW"�pI(p{��T�b����P��%�(��k �o.p�Y�'˔�TF�A(���o�{p&բd��w{���7���<R��
�	������j�/7�ƵЗCR�<A�`�C��9N/v�p�cL+=��'"�"s!��	��2��G���K<�7mL{�x!�R�.ZT*Q�\�F����'��E!C
�2>��ѫC%Q�F�"�*WF�)���Q=P=:Ue�rQaz�gX�Pj�"@�sʾphF-����{���6�5;��{�(���^0Y�Ң�<�'��� ����M�	4�7Sl�	SpOި�0���9Ju�"AJ�>ؤ��Α�-�Z�+��\�&Ih+O�Iuݕ�$M��V��H1���u�����'�t�`p��,�-j4���g��c��0	w�
-$d�{� �l����d�;9��5X��) ER�8C^����ɺO� *���92���K6ʍ,0���=�r&;O��뷯J�s� �# Rܓ�M�'�h���`(��>{��8�Y��!���>�.��f ��h�Y`�J�ZQ̓*��Ȉ�I�%&.43d��~H.�E|r�&ţV��H�
�h0��B���cf�A*�l삐���FJy"Ó�>�貦��!j�`F;l2}���n��i�q��f��K��`��!�YM�y�)	z8�@
E�ş4��5ﬨ�`��F�J��qM�;D#hx0`�'WD�A0��'CƬ��d�_����{�`Y-*�)���Q�qO�3sb�O�Z��EKziS� _w������'�x�i���%F�`�  ��2cb|��}��ȥX��D�1��&7d����ē�A�1e�"H)��V�ָnSv��P�'��-���>-�n��m�Om�@���.�("��쒔3�E�v��D�2��2�&Y�Dk�y���ص&�PTx�+V�+�HpĞ�h��|)� T�W:b��dC�H^]�Dfч(��a7k_1F6�����E�dƞ"��ԟ.d�G�f<�V�_�~X��Y|1$�t�c8�Ē�g��K���,�%<�Jɬ(jĨ�|"]��X�hT�'�"\��ñ���Ě������5�A�&H쉓�@+8�laa *ړh�r�s�2;b�$R��~Γ������(�Kȓ�=��n�6�� ��*�8�xP��L6�>�3ғ+9�8�C��� ��b��\(�RD�'��(��.���6曞�?Q�*µ\���4��);2�C@ȅk�ĠEa��q��+�Yx���֫Aj���@uB�=755�r�7��7�4�v��:)=����.�T��'nW��Q*� ���'��p��Xd�����hZ����FT���5{��[-8�Э���<O�DD*�bH�7�Ԁ�ͪ�ȟ��M���R�AB�<Ȁl!��X�y20̈́yIr��w��u[�
0s0��dw�1{�O�%���,�Q���bȔv���DK8ή�� 1D�9U�)��������a��o*D���r��%op�3���|$���*D���Bԏo6�+�$U�q�M:D��&b��c� 0���-b��Bb�8D��V�@
F�"��F@�[|]Ʌm8D�d( ��+ Z���&
��D*d�:D���)К��f��q|�0:D�4�R*�,��5KD�7����5D���D� #�y�#tVvdA� D�h2��˻_�.H3fE\S�F8��1D��0�،{�N�b��5Mu��ys�1D��Ԩ��2g4��$!n�K�/D�{�%A����g��<��(�	?D�`ôD^-ihTًCh0���1��!�	V��8Ǔ�VA�EΏ�a��8FA�2'�H��z���F�˽j�ZeC2�\��#o�B�	zw��U���[��`�J�M�\��V�j�~uJ�yRfO>p����Ŗr�b9�A�P�y��VF t#���?�2ь���	/w�aC�}���b�R���SѠ׍����5KZ��ybG�*5���&�o"����$14~d�&�$i��Hf`q��'_V� O�S�ИfH�@$���
�'�R�)�BS!d 6u� BL�hu¸�Ӕ%$5�b2�O�9�p��;a�$@�
��ZRM !�'�uӀ!�(D�"�'Þ�*��=ZT "u�&��Y�',@X�h��F|ܐ1�ラ$8�LqH��a��WA`�J<����έ�v�*֨ʮei~�WL�j�<��0w�iB��.y�Xma�J��O����$̸��Ҿ��� 5{�v�*� 'Q=���mWX�����K�l����T�cd�`�)�U����4�':vh��@�=��)H�H�/Y"l�y�x�' � !��_�(Y@s�8J%��13��z�(��z�x;*�(e�Aq�ceYA3!2}�c0F�0���O�����gUQ�����r���A-.D����7}` ��R�_�	j���N��'��RT�s�g�	&8p��P��c�"�#��B+�bC�	0� �E!�	]3v�-#�@ִAor����^&��3��'�
�y0&<=�:�KdK��8�DYǓx�� ��.�/z��m��ѻ�ΓJ�ҬyG�GT����r��p���S�~���� N�hP�0E�D��'ٰ�!�	H�S��W�Ab�h/YvQ�R�	���\�O����O�0=C	F2Қ�"s�G�h@f�Ltܓ'D$ ��&;��?�ᄣB8?�"u����>y�Xې���~��Bቝa� �##"�M�x(��	�|��)u
A:6*Q��)�I�>�����s>���M�-�xQ�v2,OlIW�@̓eRz�I�F��R���;P�F!r�p�'�T�rd�<�)ҧn!JD�tAZl�^�ه7z�؅�W.�ݣ��\�jmc�B�}v0��"����k����H�Ԅ�"Їȓf���K'!&��\􌕀m�:��ȓ	gvՓ�脵9f���$ͼ��8�ȓ,+�E��N:$K�Y0'YaɌ���h>���s+C V��F�Dz�=�ȓH�(��](W�)��C�yWTT��j�@����ɤf4�@`fb�F��!�ȓ^W�P����N�{ �UL�@��&�F,���&G�ZW������ȓG����S�O�B�j6햞n�|���]�乂�Z��<QR%�D2{朄ȓ(�t(b��2:I�A��G'99.��T�f��4!�����N�إ��^�6UQ�c�8Q^Tx����w-��ȓ7��T�$[4�$�:�胝0"��ȓ<[$٪�N��{R0�ӎ	��J-�ȓ4x,�&��H�v
�D� ��5�ȓW���E��� ��0K��z���>��P���ɂwy(83��4`�|��Z�[S��jƌD�A�Y
�2�ȓ\�����N$NL�% �&�eL�(�ȓnTc�o��T��q��,D�3��x��$R���+J�pc����%�0�M��JZ<=�cʮK_bH�󦖍-:�]��g������,]}y�I�4�dP�ȓuj����̦9��0i0g�0;���nTU�A�ɒ:�2�F����ԅ�=V0��+�}|���$ƋK�
��ȓH;���� �b��|�(��2(B؅ȓu�x�gA*�.��V�؄3��@��:;8[cf�K���e�U6�(�ʓ>�:<)N�;(��c�#�;�B�	�>��
Q��RE��(��Dn�C�	E��+�g�8�5�E.xC�ɑ?G`����-�����Lܹ+bC�	,��=[G��|E��9�EY�Js(C�ɹV�Ԝ�w�՚� �0�Q��B�	m�8}�d�'��Ҕ�6;��B�I�q��QÇ��W��D���ކ+��B�ɸ~L��H@L��}�	r��^+� B�I��$���
,A�`���׈Bb<C�1wP8��,�?0�`2�Ԯz C�S!Z�PC��5h
(�B-�d�B�I^x��P
,�8��ץ�.=��B�I�S�4��(єc�ƌ���N�m��B�>ؾ@j�}�\5��!��bB�Ii��D��> �V�"��c"*B�ə;d��a�30�V�IV�6�*C��<m���1�@M�R!���
D� C��!#��Q�D�.ɻ�D }_�B��1-Z��@ƅ\�<���`03m�B�	�nq���BE'e�A���jϚB�)� ��gO�%^Ͳ�d�V~�QB�"O�����7}RN�X�&d��"O2�Y�E<+T��ƍ�'K�x��"O���.�M�|�JvŽu�X��"O��!�b�Ɣ�9 �'-�J��"O6�y,�8of�i�*�#MD�x2"O�	
�H"8t���է̵(���"Oxt�T��!h�d���eҩ�pl8`"O|�*ĘP�%�&�هX���"O4%qC��Cr����h]�w��"O^�SױT�
���=/`ayW%K�y��A�	��l� ��3�|�w@C0�y2N
�?_�(�!F�ܕ���T��C�	�LOVE���96��;fO��z|�C�	�QT�%�2�łȈ�K�	!N� C䉘7��8��OM��<�Õ�m��B��:/�))�G��0������3p��B�	,H�A��)M@���7N��EO�C�+�Љ�mO������2iT�C�I�'xډp́ S^<`�3'N�RC�	�:�T��hK>)D.���Y%vB䉨ap��%.Z�p�E`բɡaSC䉄;�]���D������4B��0�qs+��0�<�+�� |�TC�ɴn�be�H@sk�]�%�N�C�ɫ���b ��-g(	ԅ،2��B�It­�E�N�`���e�Q;*^�B�'%� ��U��]@��9�+\5�nB�0l��p����1V�!��%,B��>:\"P�����4�'��G'�C�Ic1~�a�P m���+!�K��C�/a?��:%�9)48�3.گ�4B䉆0C��0�
��n�Vl�p��o�$B䉀?�2@j��ʜK8�K��L��C�ɯj�,$z���h2f��f�T�a3�C�	�Ne��Ą.
�8�'678����#�	9��m�*��3�h2��	��C�I��Ę�Da"��A��^�fKLC�	4��� ��?jz�(Q��\�,C�I�:��1���@|\��a��?�C�	}\|!ٖ��f�8��$`ǻ:�*B�I*;YΈI�<$���+i�.C䉎ԞU����Sܥ�"
�v{C䉔:����K�4-n�0`D��R|DB�I�2�@]���ƽN��D�r�P�C�	j)Rwf�YG�����F4�B�ɦd����A��Y���zЭC�4�C��6j炍3�9fF�Un�S��C�	9��PR���_;d���Z��dC�6v�ts�K}��� w�p�)D��@ ��`H2@I&Ñ��~�Y��(D�ܑw%
�e��&�z~e��*D���"o[6f����Q�'���r�-+D�4
��ӢC[���#��H1\�t+*D�����(��A)v� �9t�<A1+(D��xw�&���E4�:����(D��)ªԄ*w�Ua�Z7m(�\c�h2D��Z�`��e� @͍�e�l0 5&=D�ܩK�DQ~��v�K2�,̳Ѐ<D�8q�7��iQ#_;^��`F�:D���C�G�U�V�Vn��~��ճbN7D�L3�-Є�nU!eM����-K'A+D�`C7쌖t`LGł�H�x���/+D�dq�G�4u�Y���6g��5b��4D�� pȹ���<J�l�#��]9q�$��2"O�X�)ޟj1��Ԫ�8h�"O�X�,R�I�z���:�<$�"O���t��.U\ C��J=���(7"Otd*���fXm�MI"C0��d"O�9�D�4��X��P�;�a �"O�aQ���:�ūP���5"O��{��F�u�ej��e� )�R"O�M��E�n��Æ����"OJX����tul] �FW\��e�"OxH��P�J�L��8|PQY'"OP�pb��JU��q�)�#UF��"O
l�l�d3����ǊLZxʓ"O���3$J(�$@C�'=[�j5�%"O"��1i��:e1�<q90�H�"O"���"ð}h����

S�`E�c"O���4���U�����4���g"O�����#NƼ��� �lM"O��b��Iz��a%"]�w��y��"O�!�@(	_Ա�a�-u�U��"O�t\��gLN��h(�G�y��o�������z_&��B��y!�:1� 1�%scz�8����y2)�"a��C�e�=c�BIi0�H��y2��I�2�s�̌�_u���
�<�yb�&&��Z�.`:1C�L��yb�NL�܌&�X�����ɿ�y����F�h��0�C9!�(@�%և�y�h��V�h��*�vU)�(��y��@�-,����+�j�H�A��yB��]\�JL�#X8��$_�y�H�9�bI��̟�ȖDSNI��yb�H0G�a�����yRE���yR�K��x���	�%$)-��dl�Q�����&K�(8#6�8����y2���5Gnh�W$J�Y�8;4X��y�.�M�̩��D�W1@�"�i�:�yr��V~\-c���Q�4`0A�
!�y"闍qM�81O3	` 90�֢�yr�d�+�N� t5�O��y�^�s%����^�x�ndY�d��yBd̵c 8���R�@,.q	f-צ�y��V�I��OR�1���[lҽ�yh��KU�թ� O	&l�@�  �y�ǋp��|x`�,#2q��H���y�jT�_26Rpo΀�����y¤\�$Š^/���	p���yRʙ�8^�-��X;q�\ى����y�DD�r:�qO1xz���#JC/�y�O�� �%!GoЖ�KçZ��y­�$V
����Ѱn7��HS�D��y�A11�r\1+@ j�6��"!���y� )C��x�S7Z��@��^�yb#H�o��]�f�\�T�&2r ؟�y"����(�)i �M��H!���y�ņ\Ѡ�zR΃n]f|�a���y��ŭun�U����{i�-��N�/�y� ұR��Z���'��"�����y�F9��4�f)���I�I�y�⒮kft�S��̔	UxS���y�g�%��S��=0.ty�s`��!�;�,}v-�=', ��F%o�!��H%���ۥH�<TY�pm��Z�!��?~^	h�@6IXM/T�!�� ����� +�pCpޏ"��a�"O�ܲ�̊<�X��#�
nL�PS"O�rFX�t���'Ϙ!U^��R7"OnS��O�N�V��Ut���"OL��B�8�:!b��R�
�"O��p�Eܿ#o��륅��;"Z���':�F�D��L}��O�4"����a�`�!��\ n���	�'"i����F��x����?��R��Swu���B�&D�x�b?D�PH@�8l�`dJ��d���A	#�I,�p=�`V,$�(]���� �Z!i���I�<����$Ai� �e�;J>Ƞ5F�]�<�eHݒ�M/T8F�em�S�<i�L�d���� �(Q�H�MPO�<Y�g��ؐ�"P&[�I3&$�E�<9q-��d�>X®��(����~�<ѧ�:/(=��/��\AՇ
F�<�5{[6��(,omT�2i[�<�e��#e�X�k�!T$_K�(s*�n�<1��7ߺ:P/�!-d�}h`��@�<Q�Ꮔ;lflڤ���0���[� �t�<� G*y�zy���X3@��8�p�r�<�s��\B@��hJ��sISq�<aF,SV� u ��F�,�Z�9'Dn�<1q"u����Kƫ3�
���k�<��(B�� P��C�%}P �&�q�<�����{_\��8�u�T�@m�<�?O��SU���ڔף�B�<�TDG(�\�����;J�XH��Oj�<��(�U��9sf�lܜq�[N�<�*Y�l�跧6�T4��H�<��L�1�f(b��݋v1(��[B�<�b�\��>Ժ�AR��Q@�A�<!PM�/]�FQ� �=q�"Ys��E�<�#)֓pv̐�\�m����paf�<�+�/<�<(P�4.x��G WF�<	�O]"d�7��.lm���RF�<���#D" @��&\�>H�5�A�<���F[�\�&��!86�Ѱa�|�<�0��%*"D!�6�Ȉ��u�<���=x$j�+��0���i�<�E'E�TƝ�C�:t�A���h�<��G1?ј�U�0qg&-re{�<q�
.[{Fd)A$ϭY���� '�{�<�"�J"F>�"�a'D;Bp�U/�y�<�gF�iDF	��+��1R�(m�I�<��N! �E�d��쎏m"DQ�ȓp�d�:���=ҀS�,H�7����ȓ&��$U�L�e����"]�g8�܇ȓ@�K��ߜRp�J��T�-�ȓ>E�Y���p�4�bs�3r���X}@�+��!_e�mڄ��$8���QZ�L��A_܊(��J�z��a�ȓ��c'\�4��ɅƔ8�ȓs�����?h	� �	"8\����<>
E�soѕ(�n9c�J�)X"8q�ȓ ,�v��'F�b����������A�CJ
(�
�@֩o
���4�P}sG"]�l��Y�w�I�-��,�R4 G�ޢ(��D�goéOqH$��e�"YS§��`�D�6BX�+gD��p@B��S�'݊|[w@D�EDr��ȓ9Kz���LO5r�ܥ
�`̚W���������"j�0�)rB�Yf����S�? ��s/ȴ.�x�C��{�<K�"O����m�c$'
�9�@hT"OJ�2�/#�@1�r�\��<e�p"OP�;�%[S�
[bL�v	\�{W"O��;�
m*̙��̕�S"���"O@���̅�R)�d�_�K���D"OD`�/Ǒk�Ơ�w!�F�("O�Iq�H�u���J�Z"W>^�`t"OLLq�F��T��Acdo�x��Qz�"O��2�oߒe��[@n�m2���"O ����r���"��V3<	:"O�i��B��LӔ�A�S�Z,�ђ�"OdiA�ÕH�J�1B��e!�)+�"O�� �m��/�ʸcT!y�B$"O��ZqjD[���Xv�J�+�`��"OH�� �ʴ*E^�p ��}YXa��"O�Bu�L� �c�j�bGpB�"OFa�­	m�\ #	LQ@r���"ODŻGźj�A@ S��	�"O�IC�S�^X`Z�|�X���"O\1��_&ex	�]>`��U�"OhI�`8Y�Q�`�B�v��%"OtePc��{{r=j�e��m�w�!���'j��eE�4�ţy�!���_-v)�œ1܌�w�]�1�!�	N����*V+-B���@�)r!�D�k���f�S(6P�0�ؠ�!��
�IP�x�Ӫ��#1��UYy�!�JGn�b/�*"�1q�g!��ٟ4aJ��Q�I�V^��t�Q�!D!�$�0W�]0�B�6���3(^"xB!�$�R�tԓ�	11��5�&�[9!�d��O�Q�a̫���f��#t!�d��XG�(ba%֮u�P��N��!���e���Hp두ej��7.K�q\!�D<�n�����z.L�:��߫�!�D́
��,�0�C��`�4���8!�$	|xnQ�7�'mЌp��ɀX !��ډ:G�E�Ԣ�R��2���Q)!�dα�P(Y�C�[g�Ċ�	��!;!�5/�~���ɸ^�2��BbN!�DZo��a�����iY�M?!�$F9 vd��&��"03�e��M�
"!�/+�\	'�A�App/>ܔDR�'����q���g��9��X;�'Q�@���7i���W��/�����'&�xҋ ��ua�,Ϧ/�����'X��B�*�f>h#M͓:�� �'�8��%�I�_
d��qAŎ{�0���'��m����%�����<w���	�'�~9���Õ?r��*P#|4�
	�')��C�X�%�L��0��)��'N漑��B�D#ΐ:@*�Um:���'�v|�@Aɹ��$�g�ߚ�p�	�'��Ha��s_.�`�ƈVz�A�':@h�E(�T��w�G���8��'f�%*�ޔW�V�3O�z�z���'uzp��Y�Jδq� %b���'�Z ��)j���B�$(X�'�-�*Ϧn��	1S���Р�
�'��`r0�� Fwh0�a��9�e��'��"a'�fR������{	pEB	�'��P#[�Mʖ�����]�P<:�'���E�� ?�� �������� �y@(�t��k�-��'��u2"OJ=�(ѢY��[��P�f����"Ov��fl�R�� ��I�SW��i�"O�\@�/S�oW`hi�<s>�I�"O�1��Μn�N��� ėq2�8�"O,t�PdD�m� �q��@'�@q"O��Ha��C2���g�!?"<�:2"OF����Q��D�Dy��KQ�9D��ط�>&�(:um�}[	���=D�8��(�+L�k��ƞ@_�@1��=D��q��BR愡�P#J��"�$;D���k�yN2M�F��;vPS�M3D�l���G)��@Sc���>��Q��6D�`��(�5/�*8˖ ǒ��l4D�P��f�3[�!�T��#bA��`-D�|���3� )��V�l'6[�-+D��p��y��DA-�"N�rţv�'D���3%�>q2p�c�R�I�"UQ�%D��gH@,@tܛ�&�;3LtU�#D�`[�a��f��!�"
J>]&"���N'D����h����DJ3$��j5)!D����)��y��ć�s�¸���<D��`*F*w���S�hZ�jǞ�Se)/D�(!4ߑ4,M�WK42�T��&h9D�d��#�.B�<D��[�7)(�j@6D�P�wDߪpI؜"�S[� 졇K(D�`�!�\i����$��8�Lܹǋ%D�\����h������,�2�&D�����I""��q�&���(D�z �˽1�����G�\dI�&D��a����8kրh��E�� !a&D���wnj�����ę���FJ���y�&�9�>��aҒ[�Փ�
��y"`��ϖ}��7������y2"W~©c`KJ-$o���p��y�o�����.�!�"�:��ɳ�y��U5����������u��&�y��N/kVrH�WΆ,	���j��׌�y!��>$��$S�x� �9Ū�yB�P�3�k�Jt4�r3�[��y��� 7"q��1p���T-ݦ�y��fK<�x��� >�l�J�"�7�y��FNx`�)��a�@�cN	;�y2DD XP�������S�,�yr���2�<�r�aV�7��Eł_'�y�I�Safh�1�W/9�.iä`[!�y2�A.JxF��W�M3�\@X����y��l{�� �ᘔL�`5�����y�K��$b�'"
B�Ჲ@�<ABA��/3���j�P��a@Qf�<��X7]���r�!�H�r�+D�g�<��$������Y�UTDB �Wj�<yV�ϋ���>F���Ŏfx��Gx��1��0�smO�~�z��C-���y�`8�Q����wm��x�����'���O�H1�wI�b���v��)BSP��
�'V�����D�+�\*gGՖ=h���'�l*� E"e��!�х�4�	�'�X�(p��t~����K�RgTmK	�'�np���[�LEr醀ϢP�&Q��'�D)t�	>c�tM _�O�b���'����CE��];j����uڹz���hO@⟼�;S�<��#(u��f^7Ay�P�ȓ��f�U�NCD"���'IVą�S�? �͊�Dڼ8&`��F(����P"O֔X�oO�M6��1�	(sx"�{'"O�\�DM	
t�@Y3,!pzE"O��'i!��i2�����[�T�p��I�\lɒ�֏�<e8$�ҕ>1���$7K��}����r�T����+��t��A<�@�N�M���z�L_�jQ��a�̐}�<��È(?3N�rd��t��e�dOT�<YC�t ��h��om��@� �P�<!�`K%DAĹ*D��;���ȴ�Kh<Q��G#LW��Dd�?-�z4��I>�y2�Ց6X���&��%�0�D��yBC�0[o�1R��P8*��E*��!�䞅cvh����+~Lι��ϛ�Y�!���� �q�J\h0�ဥ�Q�!�6Sr�1�%F�h�a�%]q!�M�~�pH�&�¶>M<�I���Vf�yB�	�������ӆ����	-Q C��.�~(F �v�09s#����B�	.@��Bd�>k�����M	)��:��/LO��rTF�Vx�0�� kdAس"O*	�6��~��ɪ�F���޴�t"OX���U�W n;�E�!����"OvUE�¶^�Ȟa��D`�P��E{�I�gC�� �N�8z2����"|7B��f�BQ��ޚ?(00�
�=H� C�	;uo�ie�.}zdK:1!��O��.LO(u��m��N����AE�FS�x%"O��pCT=e�pȋ�ǋ�YH¡�"O )�ɋ��HE&�y�mA"O r�E�	`�<+�?��q�"O��ЩԱAښcЯ�]ָ���"OK���\A����T?ǲ�G"O��Y�'�05  l�A(I�?���d"O��2��]�����B�z:!�s�<Q��W$l<�ܙ���.@��|p3��q�<��΁Q݌4" &ޫr�~=�@ F�<I�[A�0KΠN)PH�<�tI%6<&��#2��`T�<�dhMt���{G�H	u�ڄ�bYu�<y�G)E��+�M� �kP��n�<��̋����Dj�2,^-��O�<Qoų	Q��=
�L<�-�N�<�a엖]�|�'/�7�����M�<A7O5%�"�y����S��`�J�'ka�Th�0S<�"��--��u��G̵�y�B��/Zt�]9�� �
�V�lB�	3c��8[�@ĿT����8��B�9'�z@�"G	b�6�����tAdB�	�=0�ե��(Jfl�bIA�BB��yCL衇܅)�LЉV ?�tB��b��)�̜�&��*�4��	(����k���S`_"�젆�9�L����,��ȡN�{6�I�ȓ`%p��ϝ9	�v�٣끍Zk ԅȓ
<�Hs6/�;x�`�� �ȓ�|x�&�Cv^�)��:�`��5L�$j�ް'>Ht�3eŬb�`X��4M>11�-�xW2����$@l�M�ȓ4|� bҠ�1��*�N��l&�l��F�z����E��a���O�m���_�6�P	��^����i����J��xۂ�ԐP����EǏ�
܄�f�\1r	W
Y�i*D�/�⁄�S�? �PI"-��L[ ��L�#?	�"O4��`@�#b��+�c0 ��`"O�T�-��*[ڼ��l�9"6�bG"O��"���8p�����Z�s�5���'���b�8xZD՚G#"���9}�hC�ɄE���@@�N�Zi�+�G	%2}4C�-tZ U��.]�H{�ʇ�T�TB��.�ȠK���0����W-�6l�8B�ɝ8.�p)�0&��o�&e�C䉼=]�񀆪������D�%�B�	�z!8����Y	~��8!�CE��?A��IA�x�T"���bF�����%!�ӟM��ū�M����उ��EX!�$Sr�Шa �V%ڈ���ޮ�!���k�����J�����6�?
�!��?b��ڀ�.���"�D�%6�!���Z�\��B�����W䀃/U!�䇿>;�0	%#��S��)����k!���	���[r�r`ĒË,Vџ�F������i��*1���H��Ղ�y�C_�p�9�*�4X #�ѯ�y⬒8s�Z�[vk9v�H`�2d�	�y�?n� ��1�6_s� ����y�ܒIA�L[Ã�b��8!w.Y��y�f��qm9��1Pޑ�ևٙ�y�D�#Ll��ڻ*�p}�����y����
p-��"Ɠ\z����yB��:r!Rĭӝjr��@LO��y�o�/���s�&�#"��*����y�Dn�����!{Z\`@LL!�y"�B"?	2�����(H�C�,�y��#JG:�S5EV�XJ�rB&ѻ�y�HݖrΎ��#��+��Rq�׭�yb.��FԒp��Q�w��p��K��yb��6s��"I=[�^�Ď�y"GA%v�0�Qn\(���Ǥ�yk+\����"� �)���y��E,eTfHi���3����G��y2l��4�6Ș�}��ڡ.�5�yb
_�J��(1lؖ?�S!)�;�yBɈ�[�r�$�2�� ����yb��'I�q3`V�"|�30�y�B�q>��b4�J�wr�qc���y⍑�z���a�W�@�D#��N��y��!�$*"`I�>�4Y������yĈ�F�`l;�'�5�%Ð����y"��kb�]�L��$�Bu�ؠ�yRi�2�z�)#�� ��$)$$[)�yr�:P(Lq��I� ���p)��y�%Bp+`�Ӓ)��bQ�BH���y�Y�(�Đʴ�+�|+l�"�y�#ڔ<�R�Pf+���[���y�A֓1P�K��)�lP����y���RPX�Um�,�E�GC��y2�S�lq�f"N�4e0Th�h6�y+;<<Vt@�nзƚq���״�y�M b;.������4b�e	<�y�m֨ �����
.~D0��ō�y�,�&9�	���̧|u���3/_��ybn�?Yڹ�p ��+�bȹ� ��y"���h��V<�]20B���yŜ�PB`�j��*��u�B㍧�y"@N�9� jӂ<_f��O˕�y�h�9_��U��!B�`H�aD���y
� r�[�g��Hbpa��-�!�ȁ"Oԁ�B�ڐ�d�l��~��d��"O��F� n�x�bJ
���t�"O�uF�ϨS�<�)��� 8䈀�"O�go��Q�(Ps�V&a���c"OH��F��,`�]؇�\�	ǰq9T"O��A!KC�U��D#@ν��=�T"O
U�#�%�@Q��oE�3@��R"O��+����M�1�!U�g�S�"Odi�d֪w��'�\Sv�Ip"O��+�#@:o�D�TA��f4n|��"O퉵L���ybA!��v,\�
'"Ot��WpfQK�mF�����e"O`ma��<02Tұm��^�(10s"O$8�l�#~iHmA1���<rV���"OT��wg�&HV���2D�H�pG"On$Sētݸ��
�Vo`�r"O�=Y2�ڋM���K$�"g��:@"O��֫�3K �D*�5b�ؤ"O�L�C�_6r��醈#,w�%"Oda�G+ч+k���F��
���"O$��萵��eJpc��T�2"O��r�l]>T������/;ޙ:�"O�h��D��jh��ʶ#r;e"O~�p��5���@5���J�"OZ��T� %�$�	�	4�R��A"O:]Y�-Z�al��A���a���pW"OHȇ�\E��z�%�m���X�"O|1�B�$0h�ϱM����u"O�`P���;[��KV�I �8�31"O��c��E�Q���[*S�,t�P"O`�eVy�6��Tf���V�ۑ"O���.ZBI6o�,Lf��JS"O����ٜD���V
UJfx'"O��C�[�p[a)� �Ԙˑ"O�z������A�E��c��A"OA�q�Շm�&��gS*%��	�"ON��e�#(L�F��S�P�U"O�P��'��3� ���e�Ay���"Of	��dy�ICW�
�(N���d"O8�I%*Z�X;:��t��p���e"O
����ǐ71��@�.l��:�"O���R�$`��JA�A�2X��H�"O�u�$S7u��
��XVP"O>|h��u���Zf�Ɋg�x@"O���C��(L�-%Vو�"O�L8�1W�h��[x�;S"OD�9E$Y/���L\����'>أ�C�rl*��`$�<EF`�'FFmɆ��1f��Y��쏞"�n<�
�'(<�ֈ�w]$�	g��(i2�X	�'���yCEP��6���E�����'�hQ�!n�J�p��-����'�$�õ�*,8z�АP0�m��'�<�N��8����'�+KB���'��Xy#��:��a1�ɢ4�*���'���Ai�sLx=��6'�-�N>9,O�}�\���5��.c����d�	E"���N���HM��wq ��}*���
$��=Z�pG�K�Y�@D�3D�9���v��p�B��4�����5D��b�H˫/|�:���7�MIW-/D������X��q�3E�3u����/D�h0BD�S��i���X�#ך��Ћ.D�� %�'��C˘��cḽ1�>��V���I9�C �H�ry�"dŔ�oJ�B�	�~`�85��T���'�� ӐB�ɛ�*��a�N�Z!37�E�;*|B���ppG�)�"��!%@�ifB�	l3�M6@�/k�P���B�2B�&(â�Pc�ğL��p�Q�t0�C�ɏ>���VFM1Q25
�b��i��C�I�_��P!w �\�e�Q��h��C�M�z�Is��ܲ�!B�QRC�	�P#�Q'K�R���׭[<bfC�	$��9��.�)W��P�f˙�	�B�		MBv�[GO �e�ls�j�B�	�xq�Uy`�?z���A�F?�$B�I&l�`P������8cP�B�I�'���3a��>�i`B��C�5u����X�53ޜk6b�:g��C䉑S��們�S
Cj����O��C�l������]�����k��B�	�p]!�G�1�m�u�J�dMxB�	�Dh!B��{�TMA�����b�D0�X@��K��}B�ΕH���)2j#D��J��ܙ3�lz%NӢ`l�-R�K!D� ��̎�J�v�K�i�(M�����*-D��F�؛/�|�s��)�Dk�o)D�`��b7z�2|�g�*a�`���&D�D�&΅W*���ğ�9�
�� �%D�H���Q1'�-)�@]�I'���)��0<q��ʤMcJy�ˆ�.�j`��^s�<i1jr�"d�	�6ܾ����W�<9�؆'�� cnժd!F�˲��M�<i���07�J�SQ-Ҍ
�"�K5HDM�<I��
�N`|��P��Ft;WQJ�<�!�E2�c�i!�pCO�H�<I3FΛSj0��Yc���e�A�<I ��.o�����_�h×S}�<ar-�4p�p"�g[��];O�|�<�G�~z��G��@��}�d�{�	j���Of&�ss����	��d�8��'�Ș��G�� Ƥ=�g�υs�A��'Ƽ-�ɒq����Ԧ̭6y��'�ٰ��S�A���{Tŝh#��I�'���g��$�قS�O�
6�x��'��q��DF�0ZIK 1 p��'.x�����,�(�'6{.R�'�����i�0�x����ib��
�'Ix���?[�ɷ"[1K�(A�
�'�6 ���*� �P�i���
�'e4�K#(�aP�	÷A�b��a�'�α��`�� X��U���9��hO?�#��F��ljA���M�SMV{�<��Jֲ
D���ቤM���SMAx�<i��W4)q�ޟ1���Y�`�~�<Q�k�.SA��s� � C3m�{�<�Ƥ��܉�KNY�]V
}�<������u��}i��8���N�<���̊3�`P$	ז#�)Aլ�A�<��ɛ�(��`���D�����e�h�<IW͈�L������mw\��f`�x�<�4e�Hd��J�LM(φ9�PE^�<14`2 ��E�X�	��ы@ș�<�p�$e/�8��LڠT��l��LU�<�`F�%n�dxF%ހ)�tY�gZG�<їn�u����"L?��M��W�<� d�z.��?}��p#N�9b����#"OИ�S��:R�@"�n��6Ɯ�#�"O��A��e���qH�0��ѫf"O��ؖM�e��H�'U=	��i"Ox!�e��R�� �"�U&�,��"Ol᳃Ze�u�f��6�i�"Oph��V�`�,���Ԩ��|S6"Op�U�	��%��v&T!�"O�	�EG���0��ЫFm����"OT��ϛ���5�t.��7<�0�G"OXI�U�W"Z���#n�C;T�R�"O�} 4��4pQ��H7|&N�X�"O��I�G��O�x�r�+���"O�P�a��o��SK�6���yrF�<cd�ܛT!S�Yr4
M��y�Y($��֯�4� \��'���1��DY�V��@ ��?��pi�'G��0�iD�=Ֆ���^�� 4@�'�������z� ���QЊ%��'���:��G1>������ "0���d0�48�4/P�Cz,T��$
&i3���%"O9A��;kڜ@��"V�FG��"ODݨ���=�l@;��ؑ>;��e"Ob(k��,Yl�0�"D"��1"O
P��G������ąZ�*��"#"O4��]$J	h@�9�����"O���p��r����@C�7n�ت1"O0h����>b�=��Ģj���"O8P����'�jMC�IB@����"Ol9�snΏ{;������v���@"O�E�&#΂�n��p&r�0�"O<���ݸ{����
L �L�" "O0����<u�mY��A��Eaf"O&��mB�b�(hp���+��"O�����d�+�F[� �ѓ�"O  	��ʬ
��|���[��j%��"Or5��d�<8�P�ϻ(���"O%I�ǷdB�STN�'3	چ"O��12d�H����A>bU0G"Ox������,yDlR�Zn��V"O��S��$}�̥¡P�2��C�"O�����-s�6���E?�x`�"O�Mb��՚x�b����ő;���B"Or Gʗ�C�����@�@�|��"OH�ۢo�������K>lN�#"O�] ��Ҟd!.�#B�3��"O��A����LT�;�/J�*~Z�"O�I���$<����L
P�8$"O��D�_1
7Pi*'M�/Q԰�B2"OpTŦR.��d��V��"O�c��:K<��.BxY,�y��Vl��v�ŇWFK��q/@��ȓ�vx�N�&ޭ�lRm�.��ȓ%�&Л�'��|�&ac"�a��i���F��%
s�pvlN,�te�ȓW�$��b�Z/s�h
vD� g��0�����Gi�%\�]���
27�dŇȓ��0Rt͜2s�B�ər�`Q�ȓ^AL����
(:�/�x�B��ȓvg��@g��5*��Q�K�[�=�ȓP����߹Us,y�g�K~h���4�E�3�T�u����`�isXi�?���~r�B�Q�"�	�b]�)�dl���zx�T�'Q�{����t�hƥ�eNhл	��� �XR�֋�I9�
9�d�"O�ys��@n#��!Ɛw[8p�"OS�`�)&�񦭖 B3��+�"O4Ӧ^�i���JD-G' /�""O����ܺ_O�<ZÂ5vs6�(��'+�	^y���au��#q��ŐoWe����'D���.������V,��@X�$D�`�Ce�"{f)3&�WJ�Xb*O�Z�M�&��'�V;tZ�r"O����oB�5��A�S(�
*Y��2"O����*H�j�8E�T�ʔN���K""O�z�eG좁�C�^���"O��R�f�T�N0��e�3U2��"O^��Ն��4!x�qd�	4*2��"O��	������Z���
 ����"O�� ��aK��2��÷m�iB"O� aA��0
���b�3f��\S�"Oz�y�,��Th��@Y�+��(p7�'��	w�ʱ�UR�m���X4�XE��C�+yа���;Kzr��w	�=@ ����0�IFZLp���Ƴp��0���\��B�	�6xjL�uNlc��cV�ۗ)�B�I%vcш�a��k�L%��^���B�	�n΍��V�� }A2͜���B�� 9��"ЎN�&Q@
�;!�B�I�+�r����~��U����0Y�B�I�=Ғ(��&:P��MF�!�P�=�	ç8�x��Am�꘳&E�SU���*uРRw��J����C�w��_�L�"`�D3M��e���N�z�����j&�y��k�%":5�E�ݾ*였�ȓm��+���6�&�⤠�>8�r��ȓ 
��2J׈*�dy�"�>}U���'oa~��JE ��į��C2;�e���O�#~ڃFÐ9��X�Aɝ7�B�@��Kb�<�A�Ȁ='�=&#��sI�ehUKDS�<�t(��v>:$� K�s��#�t�<����S����/��a� ���Lf�<�����45a���:��Ԙ��c�<��hD5=Jeq+Đ|<(A��Ib�<����"o�h[�YK5z��h	E�<��F�\��0G�]bDD��g]B�<�w�bd�m2dlO	�Z��r�LB�<�W<~��
�Cٞn0�#��ӟx��!I !���U�}�Vܹ��r��t�ȓ>�lP��R<�&Щ�F�>���ȓ�Йö"�)dj BG�5f��'�ў�|r��N$6s���$��%7����K�o�<	s��7{4�$B&&��8�	!��g�<������

)��	#�X_�<��� =:xL���"��(����c�<!� �,6\�3/ĆBM����A`�<������8�d�:Gj��(Gp�<�BL#z�t��➒0OP=ɠRC�<	��[�?KB����mRذr���Tx���'a"�3�=�� ��mD
I>�(
�'�b]1#bZ�*�@X׃4D{�e�
�'��c����LhRР��:�6ٱ
�'�n����V�w?��Smĳ4p�	�'�İrW�Z�*�����:Uh~0�	�'B6�taX����L�8I7�
	�'��<�D��I��9��e�;d]	�'}`)ɱ��$x���C7-ֿ4y�p����hO?����6��=�k��3���Yf)��<� ��G� Ab4����@Yl�,�D"O�9��4i��D5e�#�"O1K�mށ �̠����R[�p�"O�Z�E�{.���G\�i۪!�T�X��ğ�&��D�4e	�l���`�<Zᇜ�y���&2Ҹ���X������d9�S�O`
����N�(��8 ���'"O�̪��M�w���0c˫,����A"O�h����XED���J��T�b,S"Ojj���#H(M��`	��$0�"O2���%�.rD�p� ��7]���3�S���'�ɧ(�荨��ʥB�"q�� o��Y�"O��0V��/0��!�V�-4���$��H��� "
X���b���|ږ"D���N\�AP����S�2��=��d;D�t�2.�*@aJ�mS���҄8D� �&��R�@v�S =�-��0D�,Qa�N)V�����g�#�H�dk�<����?�I>E�4B�<v�՚#*�mO����y�D��@ip=y�ϋ�x~��X�l����&�O�(�!��)h�lifQ�͈��!"O��Q$ԯ0N��bP#�?Gg��X�"O�|)�	$���1r�5 gX �3"O�����>O�~��ASǆ��F"O��Z�=�hȊ���+����E"Oz�*�k�x\(#&Ǣ*���UO���aL��7ˤ�d��#�-	��mJ<!n�6R�NQj�ψ z��ec E]�<ɕbȑv �'$%�x� ��X�<I��57�p5�Fo�h�/XE�ȓ;\,���n'�|�ã�y��Ԅ�؀��+�H+tep�-{�$�?����-?��KB'��x���Č�XQ!o�<Aq���I�
��V���$�Q��ԇ��^�X���G{�z,XE�,/(,��W�He�@��x�C5��V�zl�ȓo�"� VC�)mR���)�&fIZ��ȓy?�Ր�Iʷ	�p[�+�W&х�
{�\� %T��)�EX� �$!�ȓ5�BT��M�;o�V9@�M9
��D{R�'-��֏@>=S�4�g�8fB�H!�'��չuGT3	Y7J�V\J@A�'�b-`P�S�@Ӟ�q֩T8h:`�
�'�\��G��<|E�ty�/����
�'�̽�G��hv�d�� *���
�'F��C!��7��d�q��=)���)
�'Ap����2=���X��?���0	�'kRPz���r����X���\3�'˼����,�`�p�	̺Q�`�ϓ�O�K
�e�e��Y!V��yP�"OP]�V��=b`��Ѓ{�2hj@"O��v��E��Q���b.��"O���pmђ��Y�Sˀ�6,���'���e�Ǯc���A�`$�0��M-�d6�Sܧ?�\Jp��~�0�˓fS�5����?!��0<��@
��~qc5.�#\M�UQ4�X}yr�',�	����J=Y#kE�:����'�V)ӷ�Ǎ1w�hFm�,L��;�'+1!7j'E>�}'ߠ4&��P	�' ~�eK�g�<�R��(��c�'�h�E��,f@�
���qFzm��"O&H��J[�tV@���ؑ�<���D9�S�I�ɒ���' @6�dthMR6�{r�W�� ��1��'`x9���		2�!�� �m�PƋ-+�F���m�1kDH�`"O��&ld��1�©3l X@�"OŒS,�7bծHysD[7Uj��"O�D2�GWPx��Ȑ��iEz�rg"O|���-�}%�X(�]�#BPd�5P��D{��	@-u[.,��X8�Fq��.��Wc|�\�b>�'2>l�� `�Ѝ���5�NA�
�'���*"A)x��Ô�Տ.��C
�'�D�j�	B1:\���\+�Zp�	�'���SŁ[�JB���'��uؾ1�	�ј'E�8���4�T���'T�=�@t���hO?��G�!� X��,�'{� ��� iy��|��OK^�� �G'4ҥ�S�PĜ����'�ў���X�����aM+Fs��8C`0>�B�	�*��iRA�N�r(X��%�1�B�ɄVK,!��)��4����ϦH"�C䉟`FFp���9��}ذ�S5����d)(�r;$o�d���F�7VZLL��~�������
� ��qRoD�N�Y��m8�'�S�' l��K�-P�H�hb��f�t���'���y$�J�<�4�x'	^(5�لȓp̮urE�\Pt�` &o�*~��U��\��EC�*B4�Z!��"1��y�ȓ&1��)���2a�=ZU ˜|�"��ȓMNa��*H�s��`x@�"���I�<Q"kD� t`9��J,X�a�B���hO�U�hl��l
pE��Ι)$�6]�ȓ.�P��^4Z$��$gG=3�L=��A�ʘwE���$C���a��q�ȓP4z��$�@�Q���>��)���|���A��!�,�B���k&���>� �'HY�@�����f��ʓs�����0Ml�2o�����=��Z0Ұ�u��":����@�H@'�l��Q��@���2�`M�Dm
��e� ;D�L�Ę	"A�5�2I�x=R�g�7D�̫�#�#j�P��ҰP�����8D�T�Cc�=O��L3�9Jގl�l5�d+�Sܧ%��su�B�m� ��T�<mp�ȓ6��aA`��g|N�!��ʋR�=�ȓ)�x�(��ͺ0�(pt'R�ɼ�D{�'�|E����0b����gL!``(���'��|���PƩs�n[��@�s�'�l��G�W[���e(���D��'���SS�g�`�����=�����'�Đ�ņ
�V%d��@���;@�L��'�x�� �<U0@�[�2'�|�
�'X*����O;:�J|h"I�)~���c
�'�詑�.Q@&�����$o(@ٻ�'{�4Y͙�gzTq���f��'-=�h��ˮe01$�.���	�'�4m��h_>0S���@E�V��'�J99ЮN4y��[G��U��
�'b�L`���4	8���%bLʤ����?Y���	�W�>���Y�U�\�F��e��C�� �>yq�ٹ!��(�J�E�HC�	�>�@K��3}�h�7�l�xB�	"^�� ��?Ϯ�"Q���b��C�ɚdl}�&�υi+T-{�C���C�	�iv.�:�_�-�D�rb%ӈaK@�O�=�}▊�&k�L�@em�&[4�"���`�����Ȼ�+C-1IĈ��{�$�ȓWPl�(�/�~D���B��H8�ȓ�����B�0E�ܐ�g��-t+0̈́�S�? jY#��λ'����Q�]b�ɚ�"O��S�X$|�uPEb�'�ҙR�"OB3�d��d ń9���E"Od`�g^�1i�5�V�S�v�-y�"O��
��#v��Q�@Z<���"O�1�B�Q��͚ "��T��"O��y1d��H�H�(��	&xy�!"Ob����&�
E�e���)�"O�c�.A�{�@���P�-T��KS"O��Xd�*�8A:��<gA}1s"O���Ʈ�=BF���B�7$��I%"O" C�I&����I[�#�%z�"O���	;�����E$�	�"O����*��U�k*j��q@4"O��W���2$��Q	S^��}�"ODP�6��@��Y#\�(, �"Ox��i�7�8|#��Q�Bwġ�""O�aD'�DXj �@C
�k�"O,���] �\�P0kI6[$\��"O�8���D�3�ŕ5C�4&�A"O*xC�&�|�9����-Pd"O �а*p p�Ӂ �n�.�J$"O���匦. r��Ntn�
3"O��aB
�5i>иC/:;sp4��"O�4��%	@t��x��V:$>����"O�!�T��-*��p"A�� Z���F"O>E{5��!*h@�!u�͔|=tR�"O�( у�%8�z�g@�=��u"OPE�B�	�n��j�H]3)Z �G"O���D��&x��1��]B�I0"Oԑ��ש0��%�-�4 1"O��1���@�N�)�'�1>:�k�"O�$aK�$rH��c���@�H�B�"O�yY��ZA����j�(a�qb�"O�yc��N���{�&Dz	� "OR`3rF�>�x��6��_?�u�d"O*��3�
�ye,X��!L�ڠ"O��2���(]]l��fiXp9�Q"Ozm���: UX�S�9TaJ�KQ"O�uz��'��!B��ں0��<�"Or\��nШT�p��H̥3��\q�"Ob�*�	
c `�e'ڀ0�q)�"O�]!G˒H��i�å�@�D傐"Of���N�[A2\�F��+,�$��"O�����^�u12�j Ý�Q�\t�E"Op,��$�52�ʩ*�a�4Y��i��"OLĊba�d�\Ju��Z|�
"O���j�<�t�X�ꀪ^M��d"O�5�3$�"�TX��W98E��C"Op	��J��j��\�%a^�Y��z�"O��L�|��Y鵈��|YprX<C�I<C��$cAkU:.��yx��f)C�	�?�r�X�$O�н���N�X�B�Ʉw\ε;��ۡ3pqcg	_�:g�B�ɔ3���p ��g� u���G�pӦB�I5w�4�Э��-�&�B��! M�C�=>{� �BϘ{�H�!P���tN�C�ɋE�ݩ���I�֘�0,ٺ1B��'r�-��
�ĕ%�9_�rл�'����V��/c��1��[R�V9�'�}��I!+��	�f Q�K2ĝ��'�lh@�L�R��y��l۝0���Z�'t��C��5���
�e��,ؖ�a
�'��8�Re	u,�P#Am��*�m���� ���_/w���r�
�D�A3"OR�
��"0W�0����96Tk�"O�8�t��6S�3���l�z�YU"ObI��F� ނ�R�j�2�"O���(G+0JE�d�yn���"O�9bS��y j� G.J^뤅�#"O�	�Ƥ:X����/r�Tx3�"O�D�E&ʝ|���4�Ǚ7�] �"O�8���.}��(&��78̨F"O����U�D��'�� �\H"OZ�Z�mM�kvf��^�
��"ON��K7wVt%I�k�{��y��"O��F,,�$�Qp�M�����"O��WJV�i��RTj1p�*=a�"O��	���!Z͘th�
�����"O>a�W�5P$x�J�g 3�F�k"O�a��AT4_4!pe����""O�5@C=7x�dö��l��u`#"O̥�R�J+kUt)���'�8�x�"O�p
3
�bվ�*!Ϟ-�@���"O�����=a6���mP�N�b��"O�eA7�ѨUF���v�5*��Y��"O���2M�6<�*�;VPz���"OV�	p�m>�U����S����"O6	�$ȅy���b��͞�@p"O�� $�դ�8UIq6����U"O�B�I�RIHi�IT�C�"��$"OJ,1�ۢ?�Y`Gj�� �*�ID"O�3c��~�֔�AI�g���+�"O��� �!�M�������"O0{��?fBRyc��-_��C�"O�(b���v~�\�g*�d$l(X�"OTPp�Ύ�R�p��ƨ
���a"O^hj�AύX�ai�Ȕ#z��"O|RT��4:�Nl�P��\]{�"O H�@(H�%m��x�G�+�Hu�"O ;r��51>Z<�3�';�EC�"O��BA�^�D�ZR6�Ҝ6���q"O&����Y�+"��0_b3�0�a"O��X�n�+n�<�چ�]qK�%��"O^�2,�g��@��A.B��Y�"O&`���¨00r�4��P7��""OJ����@�Y��Q�;Q&����"O^}q��,@�͚3�	�
��`�"O�3s�1rq�,�c@�F����E���"も7�"ła/� R̈́ȓq��ī�iضk:	��9XF>y��i�BJF֏KU�ݱp���iML=��nF4�,īQ �ܹ�HE6R�A�ȓ8x�� �	+���aF��8]䱄ȓW;.�9��!|�A��߭D\5��9�T��Ŏ�#��s#k��B�B�<i7&M):4E�%f5\�~�yD�H�<�&���&�Z!)B.>	�c�YZ�<y��e]Z4X��J�#�����T�<��u@أ�&HԛVcGu�<9��?�����%]R��I@s�<Q���'8B%�`J��5���1��Tp�<� '�%[�8��V�ћDb�P��p�<�0�3#���a�*��:3p��'F�<yGb����b��ʠZ-T�b�Eh�<�t�j���ف&D�Z��A���`�<��B��[�9%�ܤ$���э�\�<YS@�%���-��N|Q�A�Z�<� ��� �: ���(2`(���	4"Ol�P�S�s���JD�C�(m�ɹ�"O��yvh+�}� .^�S�g �y"$�I���kG�bIf����yr�L��3�@V�����&�y@W���q2KW=J�ļ�%����y��R�H��5��T-�yRN�i�r�#��#�8%:Dm�<�yB�Ȑ*C(u��-ƣc)�D��(J��y�)��? H�҇ =è��y�	65�J(X0C4\�y�k���y� �t��[��X�� V�
��y�E�:ц����ا<�\����y��N
��{��\>1��A�bV�y�ɺ-#�p���0�ʉ*��	�ydֻM�<X�bE�+j������yRBD`p��7�'R霁3a�W��ybJ z���W�D�,}2��>�y��*�d1+A" ���y�π��y���������>c 6�[�+��y�iZ�;���!��X�lTI
?�y�s� ��o�>g�eKv�/�yr���.��
!Gȇ^�Aڥ�F7�y.� 84A�P��PfpUz�̂��y��0E3���P �
3�m��ў�y�M.[���S�#�������=�y�B����<B4	7w��iC��ֱ�y�A\F�A���twb��H���y�@�_��`�� )h}١ī�9�y�؎�ؠ��i?L!2�+T���?1�'4HD���C�^��26�]#�	 	�'ՐL��jˊ][���e%O	��	�'yx��"Z2TYd ;�D�H����'�UҶ$ǈQ�|��Dd�'mc�k�'�h��A��>f0�b�
E$3Kl���'q�<KQ�[�^B6���ˌ�(ǒ,:�'�N��2��u��2%�xV\Բ	�'/v�@���r�����Q
p��@`	�'\�I�������� "��]�2*���;,O|���$��"H�a�7�P3 ��3�"O�Mp��ҰK��4���
t�\�c"O�4iS�	k��r�f�34nBuX��'��O��k �޲xE�ŝ�KT0�Ǵi�ў"~n�e���{D-�nC�P��5��B�ɗb9��@`�ˆ&�5 3C�" ����M�O�YHHE�Ϙ���Ѷx$�ȓ9��j��Ʊzv]�e���&͊̈́ȓ"�9�a�O%�-��)��iy\���+EL���Y,��YŭS5��X��)&D�$��<
/�m�EGމG)�ȓvTf�sMF��r��n�Gx��B���	I:~<�y0�̓�r��"G��!�M�`6,x�i_�sR!:`��- !���O����N����������"O�j���#{����·m3��X�"O�)�ĉ?�LH�BW�,0:���"O��0 �Y�F\|-�X$j��"O�%�� K8n� J#\�HD� �"O��#�rS�tpfh>��8�2"O��wF\�+��ip(��8`��"O|)`3��4!:�K �ř?�lH"Oixq$$�J� -��&�M��"O��k"� ���ul� l�j�"O�\H��ؕW��!8���0"O� ���s��kY$ձ�C
j�F"O(��L޸M �p�bɟV�  R"O�U�C)@�!8>��p�'�5h�"O�,���]���!��6� S"O< ����͆����H�G�5"O
y��AX�lUX�ۋ1���p�"O�(S��$���ɷ�R�*6�G"O�l�猈�)����'	L��1��"O�󱪊�Av<9�(J�t�~�Y2�O�O ��䑄x���תz�	��Ưf�!�ă�=��y `X
}j" ╏�<.�!�$C1�V� bᗼ$n��-� 8�'ua|�ń�!�>a���5nD�H���yb�^�RC>�.C�t	�Q:s����y��Q3�^���06n�;�.M�p>)L<�`x�M��!��Z�أ��V�<YQ&��np��ɚ�XK>@`�F�W��M��O��|����99�A3��3M-d�P��P�<ɣ��i?
8��e2M��2$��H�'$�xB�[�aT�-� ���a�0��Z�'g���j�u�훥$K&�"t�'�ў"~��J7_�ʕ�2�Ҳ6�n��H�|�<y��P*��У���a���6��'�a{R���=�̐�'/�L��g�/��$����I�����d���!5�T�&(S>�m�t��;M!�$0Tm�W� �k��
fFX9xa��,F{�����'F
���RY"�u���Ȝ�yb��:-��� 
�h7$Ix�˕4�y"e��е�f��3e}X�Kbo����=�O�Ʌ>��kՁ�1f6Y��"ǬYm����>����u������&
�b�
DY��hO���O�fNëZ����C�/F5v���"O(���54|͉R�F!�8hG8O��=E�4�O
re�qЕc�u��ga���xR��"J(��{����rv��|��p?����=b�0��"A:���B�RK�'M"W����0h4�J�T)@�&��'(�X5"O����Kf9Y�d��hQ[�"O�Mi���bV99Ј̦i�ԪAO<���7]<��P�Ӷ$,|���o��OQ����I�_�$4nXl�*����9o�C��?�:�pE톥(>	P +�I}���
�'�|h��u�%(C)O|2���{r�)�)��AQ��jG�="kz�z��V5!�$R���
1gܬ�E�31�Oz꓿ȟ\U�P�ۦ���d%R�(v��0"O��%K��;���c��2�"�je��v8��Q6L�1=������%� !�2;D�`��H����IAB�5K뾽Z�&D�`����3�0� E/ٛZXf���	#���2�GH]%-K��h$b

 �ܑ���'�ў"~"��U(?"0�5�� q�̑ 	���I��HO?)�g�Ѣ�v}��lޢI�D(���-D���K�5��ه��;5XD�x�!,�d-�OX�q��H�7��e,FZ��]ڢ�'�d�`� M���J(g���@憋,!��7��yH��7�x���F �
 !���{�b}!#�" �p��r��T����H>J9��蜗.e湐sK�;v��B��&F�����h��-���j �Y�8F�B�ɭ)f����]��'B3�B�	)O*8�
K�*�:! �i^8��B�ɾ~>�m�U�3ng��/	��B�0>�P+g	�:	��$n�$qo�B�)� ���bjN�&6���3��P 6O2�O�S�g~Ҧ]�L�dZ�J��������d�C?qӓN�1IӠ��^LR�n�v�<��IP~R�P�h8r	 �^+:Z`����2�p>�J<�el�U��� u�D�V5K���M�'`����ؑ7DRal�!&��� 0B�"O�Ms�/ (�B�w�Q�P�����'�Q��ɷ�ݠ:^ �2!F�?㞝a5�:D�L�!��BXjR�	�|�CB�9�d�M��}R�ēB���!aO�n�����@]F�!�dDG"V�2�%�	��J�o_�fyqO�7�3<Ohh�i���=1�h˞Z�dM���'`�'0���3�S+�Z��$��5�f�Dm+D�Hy�B� *���s�,R'�3<O��}2`�El��n�;�J����y��LA(r-���	�	6�Zr�ܠ�M���sӮ0�d��}���� �K'@���"O�09�����s���&X�P�"O�uUt��1D� 
>��w"O$���B�1{l1���]/P� �"O��#Ύ���0��N~�F����'
�'c��N%���s��	*SPl�"e ��y��Ɲ3�P�у7YghYKN�
�0<q����&G��Ɉ�K.M�"l���#!�r�V|u�T��r������8�̓�HOz#}*�iJV����4,7V����{�<Y�B�b]�l��N�>�`�ia�L�	B8�t	�D�V Q��FU�j�`���$4����'E-힕k �������V�\�<�O��y��ඥV	��БT�Bx��Exb�Ɍm@z�%@/�~�C�M��y2�+i��!S%�<Q*H�l���yDŲ)Al�j�AN+g>V転��y2LҚq�8����D b��y��-���y�o�1x�س���]�aBLS��y�`��GN�j&(�IP�h��c�;�y���	ox>i�,q��� -��y��.�X0[&C�q�*D�� @��yB�!b�� �Q�T>e��rƐ��y2(՟~T�q����K��`R�j�%�y��.M�9&`V-B�x���#�y��=�֍��
A6p�����y�aNB#��Ɂ��Dd"���.��y�.��:p,��IƯ5��̋'�B+�y"�Ԭ��hQ�d��1��G+�yb��8Na��p%$O>cZ����T.�y���#GS�Qm�=.h��рM���y���*;O�	�O�,�~,YPb\��y���^o�p�b��TJ�J�%�2�yR��2B�2�� ����<	�F� �yҧ�����sf�,�LX e!���yª��\����f�1!��J��-�yr۸X��=�d�+w�|�0���yҌ�57�raY� ��D�fica���y�L�$�������Abd�@����y�-��b�V�k��%A��ER؆ȓ.°5K�'�$-3��x�)�?Rzb)�ȓN����[�F��*����5f"$�ȓ��	фM��_�N܊���U �ȓ<��([�{�FLP�f����'G�mb��6Q��A�[��j|�'�֑�d���P�y�����O�}��'�H��B��,Z�t��P
$݉�':���'�oH��y��O@.Ĉ��� ]�#e��	_����@�$g�p��"O��J�)�MF����A�,G>� ��N�xH �x�.#�,p���Yl1O>�#f+�r�ԕ�!�7���7"O�E;�	�)y�0u`��ܼ`����"O ԀTN�8s����T白ln����"OƝ�v�&|��� f��-+��i�"OD�BT�y"�C�HW�D�H)�"O�a����L�'_�P�"O��& �0R��ph5�R�	*'"O��P4 �:z�b4BaΎ`��8kT"O��q��ڋU��H�a�91�D8u"O�̋�EO�5L��A���!`$���"O��"�H�����#�r"Ob<�k��.�@Yphؚ��%٦*O�yB���|A�S�]8`Wt���'G@��2,N�J.��i�(����(�'N�h� U	}8r�&�K?q�9(�'�Q�#��>th�@B\]A�'�������m�����J�J�yy�'�J]!d�(��ؐ��ѵ�r8	�'��������0�m�Ђ���rA��'Š��'�͢'��� ��]n�
�'T����_> ��C�'n��
�'$I2��
'}6=S3�����	
�'�a*5��;P�0���O�1xʰ)r�'� ��'��=�@�I��&xѠT�
�'x`�b�ǋ�d|tiw��NI}�
�'詩�f�0>1,uQV.S
��4[�',�%��$���{���5F���'������ 3��8S� 9:�p��'3b�Cf/ �-�.pV눀;�D�	�'x���4��Y�G]Y-��'��:�Gŉ|�:%i�˕���A)	�'"�Ui�1KVC�2~�V]b	�'��ۤ�0$��XA$iu���`	�'�����MՇ�zhC�Q�a��%Z�'V���G$SV�-���mW�س	�'Z-��ܲ/�pp�1�њ)A�4H	�'�>u���N�P����!�'.Cnk�'H�$�o�/8̒u���loX���'sny���1��Ŕb�^��a�TF�<�wB�� P2J$�27I�}�<�G�F�&��ԣF�U�a�vM�Ԫ�w�<�7��"'��Lr�`F&A0B���p�<�*Ԑ��0�b��"D��P��Hn�<�6oԶa���Rvl�XX��s3Ac�<��!� ? �J`��$�x�c��KQ�<��M
J54qA�O�������R�<I�ϊ�/�pH�B�j���t`QL�<q�M7Z�ad爞X���C�U�<i	Iy-pS���$�>��A�k�<qB�^�d��㓓C�4)3F�o�<)�&�.N��*pW���A�A�<��㏮p�ƠK�"�6}XTJFˉ~�<�3��W�5�� ��U�ƍiю�|�<ɠi@#�bB�0D��kQt�<Q��I4<2�剴��4���C�OH�<��$�`E�a��ϽY�����`�S�<���P�8x
��?�	�Pl�S�<���"?|b��5�N�*��}G�K�<)��N�N\��!O�N6�\���O�<���זb+dq���ɮ/�F�r5�Fx��z%�X]<�����g�p��/A�Wp��jU�
%�y��E��\����N��=���'�(Oy▢D��T���� �50�	ǝV*8�k!g�R�\0d"O�ٻҫ/X��E�S���	w�=*���5��$>wʄ��h���	2?�dA�Ԉ@�^bv\z�H�!�Dڥ?dhܸ��_�� �cj�{�������TH�kћpJ�qc�'�Ā�C�<&96�1 �Z��u�3lO���6�`d����J�4ir�f='l�SUN��0� ��i3��5�R!b�<�0h��� '$5��JA��#�
ޯ5�S�aE�@r1��!��#K�<�R,\�PS$᪂"O:��$&*��������H��	/r@`H�Bi��}�l�4�ފ]�Q>�w�"���3{��T��C���ȓx���3��oX�)�$�$ƪ��-�8䎉�����w@TB1�
;��O�¢����l����3V*�Q���'I0ES#�X)�0�;6�Q1�t�pFT
̞T!2�H��,Q�D�W�f��R��Q��ڰTd&48����'e $`č?y��xe٭	\J�Q���F����sS��f�Ja�ᅣ�yb�].����#&�[�*0��e�;q̭�"�.9nT��";[�G��U�u�Y1g{�]	���*����r�%D�Ӷ��T���P�w�	@GΔ�l�f\+��^>!�+P�v�JG�՟1=��C�@"%�(l��U�0=�S��V��)A�'2��9V���p�D�� ُe, �٦ �`%��yCdE���/_ܬ�U�W�aTfT�<�u��bSvpɇ$�&	5���M���'Y�4{�ke)`�9K9��;C�6D���U(8��ңgѢ-�v�#×�X����m�.9}9�"-�;1tc?A��O�R���?<�(�(�4Q��}�"O�<ҔF�28|$ٰ퀒yB��Ώ#Lj<<�c�F�	�4)��k�axr-��$h�&Q�u��z��Ұ=!�n:A	p]�2*ڏ>1a �o<RFPa��n��{����ц�Px�ɖ&��&�*`���QE��'�rX�ǡN�Yo��Z`�Z�b�q��=�#�;6DrЬ�,0�P0"OLsJ�g�| u��5or���T�V�L=P�M �SnY��h����8F�c��1G�my���z�!�dޝ������w�X @�����DFA'Z���B��0=�'��p>�9��
0@���SE��mx��[U��-{�ƣ܋8��|�⍚4��l:�〛�y�)؉u���b7�I<5�E�e-�+�yb�H9.�0E���&$h���a -�y��'<�51���ؘ�j]�y2�O��`x2�["g� ����V��ygL<|"h��V���V���y���Z�]qf(Q�Q@Ż�D���yBoȼV� Y���`txx�%�*�y�l�?Ay��Pc@["Vd�tF�:�yB致H�XHl�H�^���ڂ�yr��!@T��e Q�B(0I���y�̗�:g��I��:� 48$
�y���3$�9��)92�K�'�yr�4z��x�CR�P��yY���y�¼	��� �ōK���(B��y�&��Q���(@�|)C㑻�y2.I�Y!�@+D��s��1Cd���y�G�?2$+�Y��rhiS/A�y2�����$@C���r�V��y�a+8�Q�G��i����%���i����9�)�S)Q�>�p�T��̰!n�K\�B�	 S{�Cg���E�`����.� ��|��2+�c?O=�1K<kc�ay��,@R(i�s
O�0��§ǨЙ��T;$n
Mhe��J� `�,��0?�3$C7�,�r�Ռ�L��qF�D8����DJ�R9r����Tq�τn!n�e��^�$	b�f%D�th�h�]��C�,-��(�� }2'
TB��!�����E�4	ԩ0̭*f&_*'����e��y"�Q$_�̹g���%�ܝz�'�Q��ϝz�"��(Tp: ���y���EΊa�s��/J��dʛ���?a�a�F����V�B $��`Pf��Js�� �[.k�&xR��g���䗷]�� �@jp��mS�I�D�XP��р5e�$��O�A�"-�9l��1�J�5��܁\w�vhjSK
S�L���+J�h�j����-+QF���>�/J�ᒆ�	�\�!���S��'	|]Ġ�8BUX �x��#}�K��v��A]�+Ӕ\�A��a}�@��A���JN��G�
����!^M��W�47f$�I�+���դ�x�tæ"���,�|}ba�	,fwJ�f
3���X�ℨ���b4����q#��+WGʶE�
`����:{������,XV>�;���'-
X��	�ckaxҡ�Y&���Ӆ+e�1�Be��Z����VB�,?�:U�'�n=��/[l���)B�6ьl���R�C^�MK��ߺ�Q��?���*�`S�i�P�:��r�'4��e/T���D�'�l �1��N�P(�A��Y`  �I�4���nK�BpL�����PX��O�ȅ�ei�E`�%pR ��m�|���O9:c���kbx3�ObI��(�s�K|bEG��TJt����1�����VvLc!ė�?�lͬS����|�<�IQ7,G��'���Zz�@�p�8�p�j�z��ī�<�N|�5�B�R�q��&Dߒ���KX�O\<a4B�E�03n��h��1꤁EG"ay2&�2�xEZq�P! ��D�sO �Z�Z�ۤ"
�' 2<�
ա�,�D~2E\"�[��<x�p��ǯ#��OrM���U2���fVɡ%�L"f:�)��F�g��C�C Z��Z��.�O�l"��bm@�H�6�*����Z�c���6�t�j��
�ǉOG<i3�Q�cK^p"gg�a�ap�'��C�L5Q��,���H)^��!X,OF�j�Z�!�r�zO��|�ƥ�+5^0��2Gα9O��<2��B�I�$��XSuÒ-�j	�͒��bD[J��2�g'x3��$?����,N�V���JU�0��z��$�OH�e���z2x�)�D�\��%kJ?��X���߰?� (��)����Q휢:$�d�S�'d��*f*F�v��$>��T�:�Vu�"<dRT�Q�%D�jf`Sm��k��iX^�Z�c�<Ab���'n�IA�+=}���{#$<0Qb�6yhиf`1!�$��J���k�_��b���4�!�O|�Bc!��lJ��qOR����3����*�%&�����'�V��K.q+6�R�l@|ef�sC��[���"�"�j؟ �1��%x����:�
�j��5O �3'�d�ҒO��S���s��-k�ǆ/��TzC"Ob(�N��]ɼM`�+F��h@c�>���׌E)���?��EB�m�dA����"�!.D�\i�HM�8�td��r���z�/D�`�1f��J���Cg����`�"�A*D�̙��P/Rd�2�$��؈�+D���$ʸ.�l�al�D��}��(D���D�N�t�p�sDE�u����g(D��VG�J�ͩÇÕJ�|�pF2D� ����ڄQ�����w�1D��!�$�D��p���΅JӐ�B��=D��;���T!-:q�"�3<D����b��"䚄�6��xX�(D��&�	;�9A�P�e\蕘7C)D����*6.��
�B}h}�'&D�dv朁#��%�a.�J|�0�AI$D��+fCV"*Π�d�H&at��"D���4�J���|���6�ʘ2�<D�$�ō޿@C��G9��h���&D�#����K�`(*3��H�@pAE3D��ĕZfr-*���h4<XA"?D���A�2h�x��s�K�%tFq��*6D�p�a�&Ą�W�E�JR �4D��؅��bm��b��
�&�y�B4D�T(�EYi������J@Fa���3D�8�t
��K��T�p�d1a!.D���W.�1���Éܙ�R-��/ D��� M�;<`}�3�֙���b�+ D���� 	�l��3񋋯)J�5�",D��q�AJ4�l�x!AF���g*D��(���> �ջ����iHZ��Q:D�h�u`d�C� P�E���@!L,D�� ��㣪,.��1@g@�1�ҵ��"O�@R�Ƅ/]h2P���|��Y�"ORe3��A�fZP2*R�('�25"O�PJ�MC33U�) $� >8O�qrr"O<��A��p��Q3�N�D>I�""OL�P�F��@��s:̅rU"O�P����k���beKC"bk�"Oz� ���$�, ���7�Q�"Ol˳+;rԬ��%"[�F����#"O @S���4��(�e�G&��Q"O��+զ�0��a�<�F�*V"O����J��n!�98��l�d@U"O@Pئ J��P��9P��B�"O���aݜp��9�/�)f��4["O�bVFթC4��1�[�tv��� "O ��!o�b94$�".�2d�k"O,��R�?%@�D�Ӎٌ;��M��"O�q+�Ċ5'؈y字�5{V���"O93+�}�UB�GǶ1Ujؘ�"O�З��'�5ñ � O��Q�"O��{���C���(B��%���y2-жhqn�C1E�!b~�sf����yb#ʽ{X8l�A�E�Q�N��%��y�� E�S�Kك8�D}ᅊ�y��>��q��M�e؅.�*�y�F�A�\((C�H�sS�,Rd��yҨ�*8�A��G�:hr�u�B�L��y->�@�ōՊh�8��#�y¤ظ<>`	�鍕b�����C��y��;5���V�Ϲe��a�	Š�y��Я)�} ��	!U�LL� ���y"lКM���Bi�&H�������y2e�"d�X3`��8N�̰!��ݼ�y��B���E#��H�ȁy���)�y�`�-95ƕ�D�E�
�Q�'���yRE�,p���JZ���鈟�yBF	)����6����	M��y �_����/����A$O�yZ�
��D��}��3t*�+v�"e���&ucf�ʄAϚ��<.T�$��RT�u�h��͡¥��1�݅ȓ8ĺ(�ڨ= �t2�H=?.1�ȓ� a	��ˬe���1�i^�Q��)�ȓ3��x���*,�V�A'�N�krv�ȓRSBHiWA���	�,^�Ƥ��s�`�Jգ5޸�����[`��Tђ��b��	�$z�c�a����ȓ'F
ň����R6��jƈ �&X�ȓ>LJ Y�%��)kR/���`��}��L�Ɏ7+�Nj�D�#}˶,�ȓg��(��O�/�M���GW��ȓ#.��s�ۘM��YU��
!�����*.6�V�Q [�l�9%[fS�-��y+�œ�iA |�QV&�2�m�ȓwC���)аO�@�'���``(��\gvs�bŰ"�
���k�G�(��ȓw�\��j\"`ߊ��R�
�ZU����faQc��Q+,�ӷ�Ͱ!>y��;�^�ۥ���'j���,HI��#�ܰ��U�s, S獷2��ȓ&Rx��Ɔ�t�-0�lʭX��h��!�.t��j�1c�(- �	ѫ��I��2�X�B��Ɍ*F��kR�A�搅ȓE3�  ��Sɔ��*H�����S�? X����1���1hs>�"O�=.���QcWj9���{T"O��!��&^��0��{f��"w"O�����lm���5���4���S"O�����#;j�Pc�ƍdި��"O���/8|�I���@(9�H�7"OB��)2/ X���Fi�Δ	e"O��HG*����QS��."�"L�"O���GQ��	��H��U���"O����8}�ޑ�@Te x�4"O�i��ý�x���aŲt,lL{�"O��c�CZ�9�|��@ɴ7��T"O����%��LES�)¬9�,}��"O�1J"M�=%�m9�M90�����"O�A��;w;��bB,,I����Q"OR1��m$l�t�˄&[�8ш�w"O<܋ר"N2��fkݳp"��p�"O�8���?K^�����5	����"O
�j���]ٺP��AH�=�r��r"Oj��u��cL<i��� J�[�"OtY��С8��4��F�� ��"O���� ��3e� #勵���Y�"O\�i�� �/��d�P�9G"O2���^28��xS�� R�a�"OR�9��8'}b�9gFU�a���Z�"OpQ`���1$� ���>�H	'"O�R�
'oV�I!鍫lxf}X�"O�aD-�N�-�� �H찲�"O�*�' �
X�M#s���j�"OH�F��t0f�3&oCn{�8� "O��kdə�~���[�l1F0X�"O �ôN�*k�T�9 �K^)Ba�B"O�D�g�D�X��0bD
� {�i�b"OX��� U��HD�/�X(�P"Ob}z�/Q�?k��ȗ3���"O�4�'���S�n}Q��RP<􄂶"O�L�O���S�O�aJ ��E"O��� �M+�R �Rw#r���"O�Q�E�9�R4����]M�p�"O ���d�=Mt�z6�ޙJ4�	�"O`a1�(�ZZ	Y��"'���1e"Oh0��Bߏb�2h@�N�.�a"Ort0��S�h��u���?���)"O�Xrt"G�}�������"O��ۥ���nS�as ���<ѱ�"O"U!�nؤO�M!b]+b90��"OL����1$Z"�Pv�:#$�i$"O��r�7k��e��DL��μC�"O�!)�ӄb��!y�#O�o�,�B�"O��1��d�� 1˃��F��"O� �a�_vĘ�rJ�(m�@���"O2Q���*]��s��y�x�t"O�tH ��oL��I@c�l<$
E"O`I�t��>g�� صi�3�<p�!"O���a�
B�S�����n���!��],[K*��aM
:z���"���!�$ܴD6	�ƞ e�:3@�?I��'d�* ��SܧZ��6��<{�έ�`>~7�}��'n�lҶ&ݽ�ʨ���H>r��QR�f+���>p��E�~&�|�AJ��	����$B���p�0��0u�Xo��%���$�U"d�kj�y�F�P�[�a~B�Ln�Q��եY:Eƈ�p<q$��S�r�hTa8?y���m�6L�7��R�R����I�<yq��:5�<@D�K%�6h���TI��ZI$�]�Iɨ-j9P��� 0�3��W�-&Tا/�7�v�Zc"O����C!��]�vG+2��;��[�N<��0bk�O��
���81�1O:��F���B���S�Aǥ,ђ���'>��6���b�Z��uii�b,�l�n ��j�� a�F�VX��P�#;3k�-*�%�>�R�E�=T��#��I�G#����l���JR.Hԙ��j/�Y%�?Klj��'*0��9F$�-�&�����&Z���1�+�d�V�s��;��I..e�:����x�,<�u��(?w�>y�%M�F���b�K(�����>It���_�N1h��-}���7A	���l�{~X�JR�_#PmCT��,�l���'U�!y�ua2���{r �u��SV*�8.c�M���T�	�qZ�x�g8��Oᰔ�)�O\	pa��,���ո$�pL���Y)y,����ΚvF�+��0<qA��
y8�V��YK8�(����j�3�� n0��v�:t�N��M�!��� �n�y�NT��ԩ�#�`�	�GO^�
wdA^1*E@*:��"?�w�V��\2�ʱ>,��z��PB$J ��K���q��`a�'F0�$�:G��R0'��0|R�nL"(%��
�oSY����Rm�P}�̕9{�����L�W}���`��ٛ4Ŗo�ӻ^����#��=xCHȆBLz�+�E��(�����6��x ��'�3�Ʉ:�4P3�C
{�q����6�tD�'X�K����f����4��&l��*�:�H�V�YDyNh1��Q� ��3@jǞeI��R(���D �
Ҁ!#�яF�z�q�b�,�V� ��Zc��`�O`= �ǳ
�����W��[�
,{���*��Ō[
џT g�ͺ(�荖'$+�!V"b T���L�
�.I��OF-{z�pR��U؟�ce�[�Y�`���6W���n#?y�D�"o��o�j�G�G2��Y�q)�6M��p�mF�2ea"O4a���1<��mY�X�SAR�0�d�Z6fRjta4�>E�+L�l��(g�Q��f��33\*B�	� u�Tee0,��o�2 �H�hx��^8.|$?��ۄ�`Eܝ����&HۚT�ǈ,�O���$����Z�!��cK���$�h�hZ�KU���?!��ƹ �x��Rj�=B�q3S/�h�'����J�`��'>Y{Qa�/0.�9
v�\l�d�pE�1D��ʑD�\�l����0�zݐ7(�<���9m[ظ�%>}���ܔ`�^��Rk/ݰM[#jԘc!��*h��5���]1�
!�P��O�����.J��qO�z�ɔx����l�b���pU�'t�J�I �/-V���F�uκlb�Fmf
�ɂ"Ux؟\KG͕%]P�A'��$�zPcG@9O ���O;3�f�O昪�M3C��Rb!L)�l["O�M�V
@tT���= ��ƛ>��e�;wy��?qhd`i�\x&F�r��㵋8D�@�А��T��B΄i���z74D����l��/�>�!��+8θ\��(4D�����9iL��2d��t���8�5D�d��'��tP��qt!Ǥf���"`�,D�`hB�O>V����Dov[��	`g>D�D�K��&���m��d���1D��iV�a�H�!Ɓ�:�l ځ�8D�$"�-Ʈ&���31�\iTD2�9D�{2��\h�%�ݶ�+"B�y2�D/�&=£N}�Q���:�y�kD6|f~��� �.~�A�A�/�yB�ۻ%&�QX�G̦�dt��b��y�9>|X���(DFxs��ȣ�yR�Z_?L!�Ǡ!=+��C�����yb��d��䫷�	(�z�ȶIǀ�yr/Gll����K�
#��ؗe_4�y���H���ZWFK%���/Φ�y��)[�,�)TnV�.ܴdղ�y��<Pmz�����|��Ceá�yj�Vt�1�`��`�c�D��y�G
�� 2a*E��qflE��ybL��8�l"1�R7	_^<*�m�yb�G�8|[����	 D
���y���O�~E����k�R���4�yҢu1Xو @��`p��1���)�y
� �p:�)�zH���@˄�7bT1"Oh*"�R�+h�d�a�ʦ~�IH�"O�U�$W+*�� �Åu���J�"O��㷂�Y�={RK�V�@�S�"O� �N�3�EGi�'k��s"O��:ԍ� 'o�l�g�[�_%�1"O��
%�8N������13�x�"O��׃������Ks,@��"O8\�Q��*U�\�p�G39e��r0"O.Ps��ѶfղdCK=T�	 q󤊾[�5x�ö `Q�͊5g?1O���斖"�^}�b� �#HP��$"O��x#n�,��C���|��TA�"OH���jf𬴁��
�.��@�0"O�}Qe��.>^��J!c��A�� �t"O.$�$ ��n�qC� N���"O�Ei�H�Q\���$�#�����'����'� �*�)�0T����%� K�(�J>��ԠJ�,�O� �t�qx
��2E͓Na�4j�=*X�ߴsV�	�F���)��{V���<삢7M&Р�GT�!�A�Aa?a"�F�=�l� ,A�����O�����b=yF-N�u?f�2#��T�� Ϊ�!�·;B�)ڧDH�ez2�X2J�5𠎅�BK��K�D&'B�!)����Z�	b�O=&���39���[�w���C���4�����h�7�П�?�韠-���� ;�z�� Y:X�<�
w&��y���s�7?q�,�������sN��Q�	�*�<	�фY)8�,�'����4@S>�
����9�h�A4j��I �R��,��$�蟄&h�u���:���O�S�>�,�ȧ�ثL� ��U�p���J�$T+�8�g�)�iW�9�¥q��S�r t0�Pk1!�d���*dcK��M LR���{!!�����0�'��~��!��!��K�;���mI;h����f��+(!��2���)�l�rdi���=j!�D�-�ʕ�S慠R��!J@/J!�_)+T5����$&�~�$kI!�@jG\y�7��ٸ�:�*(I`!���:,�!�HD�d$0���)ea!�K1V��mp�H�-�tMi*̸EE!�	�6 �#L�T��jc��.V8!�ޝe`~=Q��;H� J�k�1!���Y9 }�'&@��MҢ�C%l�!��(�Bb$Bާ+���YG�9�!��C�L-f�A䧗8t�h((�E �!�$�y��96��(�=�u��,!�d	8('�b��(_����)	i%!���0~��ّ g��ĭSB�F�/!�d��`�PI�J15�%����A4!򄔰\�t����">Ƽ�%(ɝb!�d��s`DJ�kO	 �©׵ �!��,��`�@3|z� �emS��!�P�?
B�����u[��xr+9l�!�$��6h��#ǀ U�顩��j�!�$Րs*�"� WC��+��#�!���+�x�A��&:�%@+�(�!�䝩N���2v��p�|����Q!�d2v�V���@�xiT$�F��W#!�$Ӻ?Bi���2cp�2��]�h!��6of��Ҏͨ6���.W�)!�$|�#wN�t�>1�$�
!�ąGbX�a���:���D�A�!��$��r��� �dd!��ع�!�3A�D3ĭU�g�^�:��.�!�dG;Ҏ��1O�-P��L	2FU	
�!���4o�)7�S�yy �	 k�n[!���s�i@���JB̽�@
��a2!򄔯VO�sӨ
$s'�H�	�=gM!�� ��!Ȑ� n 0H�ǚ2�\ "OR��[�wEB���Ϗ
P��A�"Od`hS
�{OD��D�K� d �"O��ehД?)n�{G&H�N��"O���q�ʝK� ̢�<��s�"O6����Z�R��FD_N��u"O��Z�ā�d�xtH�
�N�S"O�=y���d�0�R�AI=����b"OlpP�.0�H�#fp؛�"O�]p������؈�E��_f(92"O�@S�0/,�zs��wep ��"O@�[��{+�ᴃ��n�����"O~�(T`A��L���8�NUh�"ON	ۑ+Oez��A�՜}��i7"O�mq(��6aV��@�4-��0s"O��R�KȐF7�� b��c���#"O���Qor2fq4�ACMP9I@"O^@�sC�U�B2��>fQ@P�"O�Q��;*� �Z6O� *J�p�#"O�8�$ą���زK�<v���"O���g��U����@ s6$�4"O\��§+5��4*%�R`9R�"O�9�f�!A�>�X���'��p3&"O�d(�(�,: ~�$]�N^Ԁ#�"O��r��J�_�d���e��iS�]�"OJ�"!��+ר �d��	rr���"O�r�M;9�t���C��#���D"Ojq#R���-|d���<���c�"O���V��8�d�3VBX�K��yc "O`���M��w��wA�PwH�K�"O�hz��ͯ���P �	�9Ӂ"O��c%B�C�	�#oN�BF�"OQ[֧ŸR���G� oTI�S"O���a���%��-M��̺W���y�̚�[��UK ��n^�y����yB����0�E�4iBl�ɓ��y��0�pt!@	���(���*ժ�yB�R�h�9&���.���4�yD�/���㌕� *���9�yB�[hq������Cc��y�jP ����a���]��@׃�y�FX9d�L�P��Ź}��${��H��y��!R�^աV+W(w� a[�Ť�y�n��l�T[6FE�%r��hu�:�yR Yj���RA�34	��&��ybC��e��ӥ'l�����yb��.���à��^	s��T/�y�(Z� E:yy�.����$��y"�T�1W�����I�X�3D� ��y�M�-�tђ�G�6�F����y�lU�0f��J� �)�9�����y2OD�,F��U $�S���yrD�b�e[��ׂ�tP2�l�/�y�+���3Ɵ4H,Ԕ�"�_��y�� ;M�R�����FXf�B�eÈ�y�$�	EPȤ�0�E��L�Q�C��y�G_���7N<hY�!���y⇝L�&��2J�iYj�"��T6�y��,(Ѷ�� �݆g�
u���$�y�AZqm��� H#6�$`a�m���y"�ުH�̜��J�* �d���dΟ�y"(V%x*E����szQ��˅�y�M],i$ꑹ�EDR��$l�-�y2� _F��q*,k���n]��y
� ���.�&Z��Ƞ�bYY�҂"O�����3)�Pq�#l��� "OLt�0��\ �X9��25_,ĉa"Op��tg�.�$���=N�|�1"O�;q�M�+�H��7쌹�"O$+��$�����#�#2D�R"O���Ǭ�e)�TV��S�}"O� ���KQj )���G d	8�"OD(�/�|�Kw��n�byJ%"O.��0
F�.�r�oQ�_���"O  P��!����a+B+�V"O�Ut�х�N��I�gΉK�"Oh�{�K�>2ς�b�"Y~��4"O�$�al�W��듍�F<��Ӑ"O�l��sZ����>/�jd��"O���L2f�()x�hR�g*$"�"O���h�A��i$
^�+٠Ec"Op �R��E����'<��U"OL�P���)�b�Zw��Z	a�"OHqc���a"�aQ�5]��"Ojx[�����va��J���]rS"O����@�R3Yt��� ��V"O"���X7O<D���A�c�Np� "O���%C hY�C��Zo((�"O
�GK��@0�%��4z�*C"O�ɐ�i�J�����&[�q�"O���dT�Y�$�W�>��8��"O�	[��q�Z@ފ�Q���_�!�d�=F�&�A�G����kɖ�>�!�ȿZ����Z�'�*q饂��/�!�B*�BLI)���b	[��F��!�$� e���^'T� �Qqh�;{1!�Ǎ�0Q����-`Ď��P��?I%!�d�0f$D����G%e^��JdJ�'$>!�^�TG��!H]�IM"�# oQ@C!��N���u�#_C6�����ѓt,!�$D�Z���Z�J��p�BW�[+!򄟇WHPp�iX�lp�{��@"�!��	m>��gႬbR2D��QV�!�S�#j�Tj�Y(O�!;'�Ce�!�DK9#K��Pm�<==����&�/�!�DA�$`���- +�nl��k�)�!�C�7ʴ`SE�����&�O$%!�أd�*�!�Ǎvr&ly$cÇYl!�D�""��83á�*g�%�U�P�`^!��#_V��0b(��S�
j�?D!�$I'M�*D`FǞ�X]�E�ɿ�!��_h���+\�sR��EfH�Q�!�dճA���"�d$�pEݝH�!��� 5jT)��R���A��=Q�!�dS)e��a�c�=p�L���9!�$�z��4{u���fX��6�L!T!�dU��6��P�	�?�X�*�GŐx
!��UޢmpD��H��@$̘?�!�d�&k.Ԥs�K~�cM\�Hg!�Ӂp�*}ӔfO�&�� ��o�!�ĉ=&��9� ��*�s�	�s!��Q~
�I��-P�	W�����L�!�D^����p�;X<��iuBW2o!�䍩[����w&�=[Ϥ-�!��d!��oalݫ`�S��H��*�D!��F)SI�)�#�OA�,Ʌ��0V�!�D٣3)N%�2�]�WD�i�!�d��O�xZw�	(?:���8n0!�� �y9�EQ9�|����zG��e"OP�!��NUu�a����v	�0T"O�̊F,/xw��P֥N�0Z�ؠ"O��C�f�lՂ���$� ��(u"Op��qBF�(@��$�,,�pX�#"O~Ѫ��X�s"��Yai����� �"OИ����>����Y�)?A��"Od� ���	*���pG�'J^�)4"O����!�sD�)C񣅃V8���"O�aA$K��:T.`��%�D= �S"OB��4�ޟnהD�A_�q�J��"O`��6M	TЁ�a��	U:�"O��z� Ӑ5b�2�*��V�0�"O"��&�'QtH�"	�>�Ν�"Oti(M�;>���`A��'|�4��"O���'k��r��W�1eh��G"O2E�0f��&�$�/�-R>@y�"O��!(X4� ��smӦ��@ T"Ov�9��)XN�[N��*��(#�"O~�Uj��7r���bf@�x�t"O �!T/�1f���sǮ18�@X�"O�����O<}�,h%-�<�Bř�"O�)hq/ϧ�H)��W`��\�d"O�!4h^�|u����C�(����"O�T#T"��A��i����8\i �1�"Or�q�&�;)?�u��`RM� ��"O�X���#}��l���J&M.!"G"O��Q�ቾ\�<�$�]X���"O�Lq�F?�|2s%�4j�\@�"O��8T	 TӶ�@�
�qo��t"O� S��::B�a��A0dY�D�7"O����K�^��QI�aLJ4	�V"OHU�Sy9�iRT ��>B~Ey�"O����C�Z�#��ەq1V��"O\X8"��&vn�0%m�("/�	�p"O�� �E��Z���-�=  ��1"O�P�QH,�TPJ��o���"'"OᘕI!��r�훑�4r"OP���mR�p�v	+q/ظJ���Q"O���
   �