MPQ    U�    h�  h                                                                                 oRB=���	����y�o�7�?I*A��KL�aUp��;�O�3���xa��
��@/3G�O�
1�T�8F�P�P]�˫����eYE�@�BZ(-k�P��E*��cY��=�/�����Q�1{9�SY�X13ŬJ�U����~�Z��2�pU�?0���m��y�e�̝��%MA��+�举��ڴz��� �q�h�V^�r���Lf��$8n�J�0z���C�g&�h�L�je��)!�Z�=�x �F+���8�W����7+o)T�>�|�>�[SVHi8�:���%e4���2��TJ�M/�r���*�[8�z�
�h��@�x�B�=G�|�8�{����4V�g*Wx#���OG	�8�0T������.T�Aa�xO}
�5!>�
ܭ�"�d ��W��S3������@�~����}2H��#i�x�����܎�*�P**Y�[xS��ۍ�,��΄���h8_9PNUt;|�Ų�����<��<�'�/E#��'ZИu^���
0��UA,�P[���^-�f�23(D:���O��$8���!9��\�δރZ�糨-�S��r�e�c���y;4U$���{��2�3X�>W����-ʴ\Z}5�z��(o�*��>$�| f�sa��إ'��i܆L�47������Aj`���'J���:t���5���l���߻���
�~m����|��\�jU����� Ž�~�!{s�؏��Kr�����Cv����gK�����,���cl䜻j市�ć���g��{ٔ����@x�ʙz�L-�=��;؅:�V�6S��k�����#߱B��N�5w�:���0�f�-��4��k�9D�i]BkJ�Zx�W�=�Ϗ�\�ka���ix��#P �R�&46��2F�N}�.�Ҫ�(�?�����S]�W�*X&Bd�u�Q�'>C��q�ʙ��?�vH��j2۶�t�=�gQrC���o�P�(%�*�U����y)u����	���u`=ڢ��*�/�/�Ա	<�ɔz�6��IQ�Ee���J�!�B��
F��L�|�?��7�&j�j�(�r� R!kL�H���<QGC�`���ޝ�>v�LY8����U�d( ���-��
l�����!&�=9��'��ʺ��⸽�$� �[;�����B � �y؆k��E�~0�)mc�8�����bNu-�ه��z�O+î��KD����&N=����6�A�:�3/��d�`���Mˆ�'�gأ���O"����eQ{y���$���h�&�՛�2@�[wOm�a�=��ć�<%���H�ѽa피v|�W3z�(���b�B�2Ǆ�f�:;�U����₈���~�=,bJ��ʍ�-,f��;�z����Y]3�ݏ�Z�^p�W����m�)v�Iթ��S�N��T�x6RRB�jA汬(Zh�%�H{��Tʌ�ӈ�t�`Uf!b���}��B����l>�͇�	߻��k����g��)6��Dt�a̾f�NR���=w�V,�;�*�d.B�[5��Zw��S��p��
k`�V8�dR:����c�TF����ٺ�oBpp
�e!??�8��<LIP_���&��sYr�uڔ��8��ao��\�O��+�D�zޣ8�K�%�q+��na��;p��������?(�H��,�b���@�8�>$���|x~�Ah�1iy�M��!��@�1���s[4
�C'8��Z5�Ra� %���k?��ػ���9�ՁHƝ��(_^�y li'�ן����������KT����u�	h79%�GW�A%��WʼDs�U�����5E*����V���K
ªr�u��PVb �D��\�;6�q���OOk�W�FnЖ�?��R�,RL��Q���n�T�g��.|����9�o����Z��@��|E������M�u��׫M�����m��9v�%�L2�Ї'BCi!\��q�nI���e��`��%��}�p�Q~�dSQbY'�z*l�3���L}��}KØ�f�pʚ�rҟ�%��)'�(IN�e��
{ܨ!��>�kw`�F�lf�֮��K�^��㑔8�Cg1<�XC:!8R��t�Qی�kN�c�>���&Kp�9HO�J�be�"�晟1��Yn�&(�Y���Ѐ�	g�KO�ѽ']\�]���k�6%�i�ߜ�=�/�)�#*��lw_Lފ;��݊c2|Hn*� ��K"�?�E�q����Z�{;@���XmD<��ڙ'^���)=4z	l�e�'ъ�A���]?���\��Ȧ�ّD��F75���=<b�� �mS�p���I:�p�aI�=�X�����  nwuZ0�"���Q�����$Z�XJ2d���z�	�q5Ix��6��¨|r�ek�ۃ&I�0a:i9l�)}��Yҁ~	��W!1o�0^î;͸FV��D {����-(���6��=��<���@���?*/[���Ic��%V�H1U�u����9<�d�Г�>���N���]�ހ��ݓm��8=����:�Sޖ��ŕh~BW`�+��H�̖���~�$�t��t�2)r�9ي3�:�^���|�4�� ����_��	�5!�o�d!^��V^�{�+�1�dI�+�~|�e~V�SX�!{���8�n���ņ����4L5ީJxPob&�������(��sX�:�-~�5�X?	ZYͪl�٩
� �& 6�L��"9q�6	�8(_z&.���l �ı]�F���y�i����$��"x�:!��|��o9$jK�Υ�ԧDXNc0�g2�n���������+%&�!"%hC�]z7� �+AFD%��r���j�Qk�Fm�S�����
$1�T`bGR6w#�#Ur���0��<�

	j�4�Yn�}h 1��m~(�g@��޳!��u
���aA3I�t;��c��)�1vE,�3�{\�ҏ�_�.�,���s����J:��"��b�p�xW�|O"1,bc@y���:k�V7,��^��FC��4�[�����H=�L@^�O�1�rnɽ���[���e�AYU4-z��ܔ�7�'"���i�7ź��m�		�7����.N}l���ucs5����[���f��$�ۦC��ٟ�����ʄ}]�Ǹ��\+JܩB	�̠��������Xϐ��`M�EZ��p4����nzm#mv����;����I�f&�J���%�ŧ~?L���$�	��\
�Z�Y<r��'͹�{ȃ���Ҏⓐ��h�9j�$��Ɋ��'��#%F&1Sޓ���M��"o�/[>�,�|�w�Ԯ��VC�1���7�cq*4��]2&�J�C[��d=F�[3���e~Mh���@�&�Bh��W�ɑss������/���gxӄ��)(�G�P��i
T�Oᬟ�E.OGta:�}Š<�	
W��"ݹ|d;��W��3�&�D�@n���U��r��,�iY�xM���5���A�P�,��v�lD����,.���ܨc>9���U/ɟ���}▟����<��/�}D]�Z+0w&�׶/�=��u�|AG*P�{]�Y��f8˥(��؛˦��[��ơ�t��\����~��Bwo-��U�����|��Zroi�9��vʏ2"n����܉x�/q}�F=�(�u/�%֧>�� !0�s(=p�So���4��vU4��>��h����e��Bɒ.�t���K�%Bߙ�[���
�R��[:��.��׷?U���:Uz `�~�\t�U:�J��K�-��Sv�U��!�o���Z��Tqݜ�l�$�j�p���گ���$����v�b������x�=�z��@-^�*�@r~� �1V����$���|3#�k[2�N��/�u����$f2<�6{��&~DĲ#B�#ZS�ԜxC�s�IkMx��fx�d�PO�R?�9�J�N����Fs.��eƃ Z����n|�Wk-�&��d���췺>>a�q�̍��U�R�NP�2���t6�Ag�QC��}�%bPqR	(@�m*���˶Yyd����(c��Q���`��z��
�/�����<IF}�i`�7�I�0�eRi �e�����
!�L�5?m��2�)j<�L(cQr m���pK����Q�X`� >ޘ��vY�8Bq�pSf��'�ʁ	�f�lF�j��L7!s��=� ��B(��5�~⓼�$����\:��}B[ ]�Oء~�ږ�2�Y�g)�HZ8tf����N�L5��X���?���4����<��D�u�!9��Af��Qˤ'������/����o�Y<ˁ���fy�^�/�އf�n/�e,&��(]����v&Ov�����[�r���箆�p���f�}���-��O�|f�z=Ը����}>��գ53~�)�h��#��N�a=j���M<�f�q7���_�O��3/y�2�I^Kg�P���
jv��$��ۘ�	~�T	H R���j�+�c�"���J{�G���N�zה`p jb6�'�)��I���F�j>�P�d����Y�ԙ6gr� 6��t�j,�Y!�NM���
�ˉ�,�t*e��B�^фQ�vwi�'S���&�`��8��y:&�/�����o��GjA�^����>p+���l�?��L�Į����&�0qY�Qlu�����w#J��\G��OXB+�~�zmW�8��"a�1���]Ga�9*pP~V��󯆚��H�|�5��
��=Z$*�+|J��<8:1�HVMg���ڬ���w44E!='�R�U�wR��V���<��y�¥93��Ha���#h>^A�E ':x��T�a�ܾf�V��V�T|�����,	Ç�%A�^�,�\E�ʗJgKI���{��0�*@�����	@�%��uŁ��ݵ z�V�WS�6�X����k� B��:y����ԍ��,�
U�Lp�ɦG�"�3�I��Ÿ�J��X���\j���)rJ�K>�ha֚5:MЉx�����΂v�Mf�Yj�B:/C���)Tn$��K]�f`.��t��=��Kdn��b��zt�n���-��� ����Ȍ����p���rM��%�U��d5���oN����e#��;mY��w��F������#2^|L���έ���<�n�:���R���������c�]P�G%Ap�y�HjJm����}��`a��r&#�L�,!�~^��57OA�l\ߗ��o��6 G�i4B���� `l��*��\l�Kt_���;�J#���qH)�1 ���"���� �qX�-5'�v������X(:����'��v�|�14�d� U�̠�A5�`]�Lp��^�CB�f��D��7��x��b=q �y����� ߭KB�Iޮ�Xn�r�ҬNnҠ^0�f��K����������d�����d*�5�I�Q�a�#�'�@wa
�v ��q&:ĺ��侚�(�,��EE�~�!l0�7��6�1F�z��|{��ר:����[�xUX<:^��;����X)��c9���#>�S��繁&���Sg��N��� ��<�]������ǆ��H�ԗ�US��c�@��~�!�f���/r���1���A�/ut��r�wI�Ѳ̙����z/�/��飹���w�z����9�5�rџ�>�`�^����Fr��4+�/���R�V����\Z��4n˝N� `��Q��LPzJ�o�b���sė��'sSU΀:�X/�kZ�7^G;��E�8���66�|��}h���#h�A_�/n.[)lZ ��LeF���yo��{(O$�@"��:��e|=ƖoԖDK�Κ/-�X�~�0쯿2,Y/噇��א*e��F�|�Wh�����78�c��D`3>��>{ƗQƞem���!���ȱ�A%T�-GG��#�J6rީ�0F���
�5,���Y�}h�O��~�P@�Xͳ<wM���޸�Hn��t�R��^Y�)%�;E�u�Ԗ;�
Z��	�,Bg�$���J�4ؔ@�}����d��W�1g��@�5�zV���\"�a�B�'��s&�􃠑L�
 �J{�}�)Rج�Ǫ"NE�l)o���6��2|�"T�q!r�R��cm�tD	-0��>��Ѽ&.��8��q�c����w@�6X̡
:$����>t�����r�����߂B=a�7?���Ѥ�g�~'�� 8��Ő/���uE5����
��s#nu��*�Ȃ/;�(��Gd|f���a6�`�<~:,U�q����m�\%/qZj� rZs�b}M��2҃ҩ���鐽5�hGj[����D����ȮENF!�����.f o+>ԗ#|�= �IVbV>�&��;ե�s4���2�l�J�Y��5|���[.�Ϊ�	�ho��@�iB�@"�2f?��O#�GNr��E�w8x���D�G�,��մT+7٬:v:.J�aw5}���Wf�
�܀"���dv�*W*R3������@)����ys�(ͽ�i��x�$���m�TyjP�O3ÑLr���G�,i劄3�!^�9��U�v��\������ <.�/{���*KZ�������B�
���P�cA�H�P�a �T?�f���(��"���K��A��|����\4P��y��Z�-\ј����Yf"�5����T�[��q�_2u0D��S���ʪ��}�c�x&(B�˦ ��>�- ܔ<sC9��΄"�o'X����4=:���-��;��TI�]�X������q�Oz+�4�o��`
l}XȆ��g�R��U����u�� �lR~��))���vK��#��b�vjŉ�RLNB
��7���9(�W�&l��jB������[8����q�,�j��`�x�,z�@-9�)�{�Uػk�VЎ�����7�#���s$Nm����� �f mf������2��6�D�2BaC�Z.	"���܏:Mk���q�DxB!_P6�}R����u���Vݰ�0m.�����t�q$�����W�O&xUAd�����>9I!qHy�s��|�ɽ�2��ntq��g�e�C�9��t�P,�Q([�*z�}ݦ~y�v�US��iv�E�}`����]/�����w�<������}�;I��e݊���8#�
���L7�?�-Ij�qN(P� ���B
z�i[�Q��`.l�ޓ�v���8������ɩ֥���UPl�n�����!��0=�C�]Ԋʰo�nۊ$�_��3�Г�B�V ��ؼ0�y��4�)�M8��� wN+��O���p��E�R��g��waD���D����RY��B�	�0Ӻ�No�����!��|�U����#԰�ߒ��he�N5$�ߏ���&�6訷�[����u�[��e���ψ[)ݞx ��sQ�
Jk|/��z��u�l�hԸO�ǺO|�0j�����#��>�[���I=��Y�F9���j�f�s��0A��
:3J}Q��Ix^&�f��8����"v���RH���u�T$7RRH�"j�	�����[��{��m�B��5Zu`��Zb��3������}��K!>�s�ֿC��tg��^�g�_�6aft!�K���NH&��9����"�,!|�*��B��݄�^w9�S�|Ƣ�{`O7h8�z�:��R��w���j����"�V��p�L���m?5i#��uL�X��M�7&���Y(��uP��&���2%խ\�%�O���+|�nz��.8q��=���Ţ,a�p�o�������H`[ϻPЏ����$e@�|����7(W18M"_/�2L �'~��ǜ=4��j'n�P�R���l��Y��9C��u9nLeH������^�r �*-����ܴ��AY��-�T)ֻ��	�s%��G�כ��rp��*��.��+-�*n�?������ ��u�R<�ɽ \�R:g6Kވ�kSk�ɽ�<'n���ȶ�,��u�GƬ�$��ݿd�d�኏���%�]䓘������V�� ��懘� ����M�[�1���5��v����r��l@C�#���|n�����uz���+�3�g���Td��bO8z������p��A^����3f��H�p ;�r�F�%�(���c��^��Nҗ�������ytpw�hFjHa�L܁��^w��J����<���:��R�#���Cq���nc�>��C�p�ciH�/�J��O��Q��ߨ���&ٛ��VQ�9���PC�O��$��\�
�C6/ii�煳����3�<*nl��_�ײ;���Q�H�� v�"�A��nSq�q��Ȭ��q�VyCX�O,�5U�'��W	v4�����7��wA��G]��5�'����wA�D�m7k���b�&� >�g�����?'�&_I@9X	LF��x�n-�0�ڣ"���� E��;��bd4F�z�����5�۳�l\�)���Q��\P���G:\'�����CYh�w-�Y�g!��[0R1��1'FGBO�{gt�#m��e���<���6�&�����:k������ 5��j�vv�TQ��[����	kϨ�%����U]�n��<da��r��4[�!���S����~�<S���D~���0��4Y����t	�rv�Ŋ����ԇ��U���*C�DG��{�}���s���a5�Ks������-6^����s��\O+�[GV�;Ք�Y�.�n�W�{Y"��dLk6�Jn�Ob���"~��^K�sN�}��,��tmXJmVZO"+��܄�\u6��=�ط1��^�&=_b.6��l� ��%F��Pyʑ@�6�I$нl"n#�:��|x�oo)�KzzӚ��'Xwϫ0`2����tbJ�.ԍ��b-gc�ע
h����:��7�m�,�D�tx��a�vBgQ!�$mh��<7t�uʄ�rXT�y�G���#��Sr9Ъ0���<�
�:���_Y�hPh6�B� ~�m@h՟�W�okXޓO@���tq���Y6�)�
E�}Ա:.҅<��&�,<�?��
��UJ���'���sR�n��2�A1�2v@��!�01�V�Rz�|�q�*���N����#�LB�y�EI2�zP��V�.`�����m�)���g��-�y"�3��,U��mT$�ލ(m�R	h��0��̐X.��C0�c�Az�򙹎���ܮ�$�Ǧ9>�U���-}��?����s����y�y���u�]�Σ��Jw�VXE�.�5���tnp��#���=�Z;����f���'[��`�~5,��̻��X�\@q�Z�D�r5;��M�;
���t�D��x�h/t�j֥��iN���I�OF=��I:L�?/M �o�F�>�"|0$����V9,�K���hA4ՌS2�NJ`�c�#'O|	[)�"��`h*@�[B^�Q�Ge��K��ѓй��xM�xI�l�_��Gz)��a/Tf>���d�.E��a�x};�rr*�
M$�"�!d���W�d3� ���:�@�E�\&�k͘бi��x��(���ώ��P[��ì�}b�1�l�R,�7��SYA09auU�D��� �Ц��;�<Ga�/����Z�@o���w<�E�+��A��P,g��O��f�[(u��=��Q ��W�)�\����t��]�-@���Km��o������zo7��lHl2�^��o�����%�9}�GN�c(�⿦�E>5�= �hs^U@�I$B�J�k�7+l4��+��#�nZ�d��x�p�$��[8���(�����F�
�,~�Aq͠���Uie��5� ���~�2���;���2K��d�I��vEUv�����4Z��}�=??�Jl5��j|�肮0@�8�8B��l����B-�G_x4��z}�L-��ɶ���V4�V�j�����#0,4QհNH����<K�4�f�_��g����RD���B��&Z	E?���بk����8x���PQmR5���\����:�.�)P�9���,� ���Wa��&S��dQ}�"��>4QSq����.�����DK82l|t�fwg"E9C�Y�ۦ_P�-�(vD�*�~ ݁fy�Y����w��T�`n�V�!+�/y���e
�<�A�K��x�Ib!�e�p�������
�!Lr3?�i(7�j�$�(�n~ �����ԵDDBQ��`���ގ��v��8�5����A��wր�V5e�l|e����!)�K=jJ��x���+[��Iq$@, ���(<BK� �X����^ڌ����)s�8��%���kN��
M�3���{�����<:D�,��o���Z����]����?|�Ď>���~��wy�8���ԃܰX��de��aL{�����K�&��c��[�ڷ�T�����8!���k�s�Y��#`���[|J�z3�^�Gt��p�U3[�+���fﵰއ��Y��D4~=��ف�I胹bf��C�����ş~3e�'�(�^V�ƪ��>]Svװ8���#���T?F,Rù>j�KP��qӟ��{��ʝ�\���y`���b,5���G��z;�|ۏ>���&�/�,
D�gh�6<�ut\q�̏��NCt`��D�Aۻ,<L*[/Be�Y���w��`S��k��S�`
{�8�5�:���͊��ۘ}�4�\��9p�x㶘P?��Z1�L�j���&�n Y�NuBdA����� _\��OP�+wR�z#�D8,�cX9��}�aS��p��>��]��Pu�H�&�k7� Hs��P�$�u|I#R�281zG�M�Yl�M��ڢ���v4���'	:KfqRr8�V�s輖,�9�xe19�7UH�5����^�p� �;F�(���W�0��1�M#�T��xֶh	y��%����b�Rc�M���+p�ɬJ�&i�*ɖi�&�)�#�Wu{C:�y ����MAW6��y�&,k�Ƿ3��w�z��Z,#��B�E������y����
T�� /��κג�
�f(]*�������/�+_�M�M��l!���W,v��@]�и�uC����Qn�&r���@�����^"��BCՂ��d���b�p>z��F����c����gڎ#@�A�p��rC�a%�p�ڱj����N�`�����R	�v�w�k�FE�6��Z���^rT]���ܭt�q<���:� �R~l*���<��c��h���mpMm�H�p�Jc07��E�P2�*[&G��a��g�koUO����/\Ul���P26�i�<��n�+�b�*Ia�l(6o_+;檂�t�H��� -x<"�)E��c�q���cD��l|z��cX��
�PB0'��/�2�
4+{�6:S�,4A�͎]p�_�B�:�9�Z�DVI�7}m�@b�f� ��7��ip��M���IT�nX�$2��d n�WG0P���=�����εܾ	$d�Y��u?�7d5z=�ć��Rw����y������U�:zU�Zx��^���4�4��!⅏0�Je�,T�Fg3�
L�{2�{מ��@�����k<pG$�1�&�P��=ќ��ݚ�&�ٷ4��^E��@��	��	������k��2w^]of�wWF>O����IN����$LS/ǥ�6�U~����܅������ɏ���F�t)$�r�TN��LS��6��ݛ%]��
��6
(���c�z�R5�D}����ɡ^�d�<4��.+4�Ň�[{Vn�˔�x����:n�1��r-����L�J�bb�Eޤ]� ���
sIY�>qn��D�Xe4�Z�li�l����Ql6�<��3'g��A�l_~�.S&l�`zĂ� F��y%,��ӈ$�Z�"�c:�:|�<o
܁Ku����)X2@�0"��2"Pv�O]�i*��`��8|�2�=hA�i�UVs7.D���bD��F�C�[q�RQ|��m#���W������;T�-G#��#���r�10�����
���Y��h����2�~9��@#rV�r����(�n�'�o�t���T3�)ۦ�E]����Y�� ?��xC,w<,DԈ���JK��N�I�}����(��1��M@J/�+��VH�������h�8x�)Vd���xL����@��B�O��9�I@W������!����l���(�"
|�����`�Y��mxPj	����� �Ǆ�._w���Zc��p�m���N�s�$�/�4��ٰ!���z����p�8����%�ZPXϝd7�t�Вc���_�e����E�_�p�J�S��nk�~����;��
�=�`f�)e�=����O~0LǱ'ۅ�:c8\[�)Z`��r���=����_�ҟaV�3A�hJ�njQ��fi��F�����(F��ޤ���O�6Xwo�Y>��n|k*���QV4���\����4��2�Y�J;�?�^8�MR[$��v��h�:�@7�uB�í��G;�$h��}u���%��Cxj��z�>G�EezT�eE�ps,.@�4a->�}�&��$
ȋ/"n^[d��@W`�03��C�U��@�},+[i<:�s�Vi
D(x���=Y�
H�P���Ǡ1��\�G��,�U�ik<T�C9��U`2��1���I����<���/�M�&�Z<�a�T�(� �y���A��Pǌ.�JщfIT�(0�B��h���v�2�7%��\jQ&�o*jS��-���ޱj�O�J��� fU
3��g��2+�0�*���-
ʠn�}�K����(xI�$>� > R�wsy�D���͞%eo�r��4s�ֶ�(�� L����&�����6���ń:�j&`��\
"����+͠:��HX�UDj����k 1��~������{,3K��m�ăv ���T��G����D��d���zlP}�j��{���0�s���ӿ�gݴ� �5�֢qxOW�z��d-����U����V�f~�5����k�#K���ViN#9y�&	*䜇�f�&ЙG��W��DN'BW��Z�,�)i:�D�\k��'
�x��*Pl��R����c!���D��c�.��Ɣ����{����W���&.��d�j��>/y!q��%�����0���2Gj�t�^`g�DAC��`�6�eP�ˮ(���*pw��\nSy]������S���`)�Z�<k�/��k�@��<�Q�扭sr�I�ɻe�$,�����. �
��L�!?>`�#��jM�1(��� ���8�[�M�Q3%`d��މ��vj�\8s�f�����[=�p��l|��!�G=%�̓��ʦʓ�$yG${I�ǁ����UBl�� �8T����C�ꗒ)Y��8E�X�� �N�j��r��NԀ�;���~����GDP�s��]�R���!�x5A�&���]�Pn��WA�r����؏I�/�ߡ�e�����x.z��,G&`g���[��k;ن����s�%�:�n8��)O�W�|eP�z�t�"x/�.(���6r�&8���E������t6�����=�ѩټ'��(%f��S��#	��L�3��e���^��5�=z��6�vҽ���i�:ŐTZu�R>��j����ʟ���{�o���tʈ���`�5b��P{�7��"-���>���u(����%Iog�O6�&t�$��*�N>���2���P,W<L*�r]B@'F���w:$�S���7��`�ފ8!:�߼�e�-�@k�����
����p\
���^[?+\�Z�nL5�դ�a�&�=�Y���uƻ�\=bv�3�|�\��iO�Kw+r�Wz~�:8�s���/��X*ra���p!�f���Ɔ�y�H�Z�����{���
$�
8|�s�-he1�v�M�t��ha���}F�4��b'�	�Fa�R͒y�5���"���Su39�B�H2���Z^R�� XlÓC ��+����G��9�TM��ֱ�z	�8�%rv��}M!�ͨ��(��L��d���!ŕ*$r3�Bb+�D�8�uVT�B� KS�Hh�6�*����k���2`<�Ro��>�,���=�:���`�SYs���Ê�˾�ە��	���-�S�������|�{���(��!�Ma_O�n2�kLev�������s2�CՉ�����n����;7ֆѱ���^�=�4d�e�bE�Fz�KZ�j�������� *����p6[�r�m%t.o� LД+�N�I��vܧ���w
Z,F ����Ӻܷ�O^m�� T�/"�<�p�::0RY�q�=,&�׼�c�zϲX�p��H��J޴j��Y����X�ňS&MN�=IR��󆻍O�O<�H�\���@2�6&9i�2�)8�!Ftݵ�*$˗lc�
_�P;;ኜ���HZ�� H��"��ձx[q	�������g'�nXY�,�kO�'`>�i�4f6f��\g���AF6]+���]}��ԝ�ĒD�e7�
��TbN�� �\���LR�5���#�I��8X?6��p�n��+0�!�XU4��#�ΐ�_D��dj���pu��55��Ģ�Q.��Zq�`�������:��b��L�y��m\���!x�0����'��F�?x���{Me�2o�~:�)�<�˾,��G�G`[��q��|[Ĳ�$��gH�P*��kd.���p�п��3]J~x��j��Q�������]SJ#��#}~����d��3��B�꩚�`
�tD_�rl�⊟�{�J�l��ٛ �������Xv���{���o5�]7�P2�1�E^�����P��+OćQ�;VI����p�d�n�+~�1���U%L��Jd��b��,���<��N�sDD�վ�k4#X��ZE7��(���fY��Nk6��^Ύ�r�"4C\�~_�N.��l�!�<�F�k�y�����$l"d�x:���|o���Kp�q�@}�X�Є0=HY2����*xP���V���)�����h��~�p�+7�:����DW��ޒl�ZQ���m�.��r��k-��4�TLr/G���#�Br�|w0w���C
�z;���YZwshlk�撄>~�pI@�.��a�e�I���t����OP)6c�E�����{a����,��,�(���g{J�l�	��Χ��dM��"1�Y@��n�&w�V����P���'� ��=�4�jLx*��;%5�ծZ���d@{���l­dF ���s��#��"e�����
���
�mSnU	�[�f�*�.�
^��c�͏�謀��R{�RWo$Q���/������@��%���c��:ܕ?p�8;M�o���+|I�D������LKbEƽ�᫙����gnf����ȳ�;���s�f��8�x��1�=~+�j�������\vUZۯ�r��NA�q@��j:���l����he.�j̦hA�R��Ԛ�m�Fɱ��D%���GQ�o���>e�<|�PY���V/N���O�h4�i2 2J[���i����[��k�h��@R�BT�5��h��_��9��.Z+x�K���Gp��@ٔTܬ���).;��a��}��e��
C)"IՅd'*�W�w�3��Z���@Z{G���N�iE��x�Қ���~�eߓP�w���z�X�3�"N�,�+���O�9�DU@��LL�₁����<�'�/L(�T�Z��B,�C���{K���øA3c�Pbҹ�E�}f�lq(��7S�G�d���`!\�j�����-�};��7���� �ƕw[���N8�bF92�G��7��H�u��}|o�)�[(а�~T>� �ks���?�Ş 4cܭ_S4����<��Lץ�W��m9���E� :`��<���
}�)ȷ�U7L���LU���&�$ �c�~刲:�=�6�wK��>�?Dv��?� �z���iK��݈:lk�`jr���d�Į~+�n]p�b.s�{���xjJFzsC�-ʺ��,7U،%�V����4��hrz#fȝG�MN�	�a���7��f�ϙ�ԅ��7D0BҨZZ��d`���uhk�Tn���xsgP�_�R+��}���:�f�U�+.�+���ň�����8WWw�&	k8d�wϼX��>*��qY�؍������:�s2"�&t"w}gXdC�%��k�P]��(�o*���7��yP��&�p���Vo�`���W��/oY	��<5?Ք��n!I�e>�B������
��eL�Z�?��_�Nj��(O ������u�QnX|`�n�ބ�vŤ�8.���>�6��6����l��&v!�T"=�d̮���!Z����$��Fb#�����B�G I8���Tڂ�a���k)��8��#���(N<
w��уi��߶���Y�.�(��D����%������Ƥ���� 3�zn�������#g�m�B�{��J��J���Z]e���g��h㎄-�&�7Z���[�>K��A�����Į#R,�Оiiф�^�;)|��/z)Z������i�sǋZ��!����B�T�#���ۊ:M�=s�	���@蹶?f�9��A��;�3�I���^���<�D�t0v��<�cM����Tu�xR��j�/��O�ԟ,_C{�g��SlX�f��`�Hb"aVX�5�R��Z�>�\���JP��P�@ng^YW6�'t�����K<N9p?�J����I,rLd*Q�wB���=�qw��yS�'���$�`�b�81i:>�@	a�{Ty����.0�g`pp���D�?�N5��Lp�����&�,�Y9˚u�U�w;�&� 2\3��O�29+m�Vz�|8�é��
o(�3Yaɢmp���Gq���H�
⻡e��<���h$ ||-�(�V10�MS�R܃��ژ���X�y41�,'?1�A|[R(��];��p��	;��.��9n1H�:D�@U^��7 ���^h�M�5�҉���oT��P֬��	/	%-R����4�H_R���7�f��]�A�*m������_B��:*u1�F}N �&��C��6\���ȓk#��ǭ��-K��y\C,YE�8���5,���P���P� c��D_��P3� ���5�7���ԝ��!WM<���ە�a6v-�7L�.�LC�s�� n���7~iҞӆ�$��DǺ���
d�:Jb�Azqӽ�Z�񯙡�����D�s�yr}pQfr91�%Oa��P���/��N�R���ۨ�J�Ŭ3w�h�F�����ll�Rf4^h�:�[rk����<�:���R4^i�x��r�c�r��^�p��oH�R�JYY��i�
��]S�`�&�����"�j���'.O�>�n'\�����3x6[�iz�؅��<��X�}*�Tvl���_S��;܊R�*�H�0 c�z"�PՌ�'qD���Ӊ�b�M�g�FXQ�ˆ|�'}0��H$4�7�l�S�8AA�X=]���x���/��O�D���7<�B��b�G� o�d��O<���?��YIʳ�X�5R־�"n>��0�<�sC��հ�k~��IdA��k���5�`�Ľ���+�ڬ�hm-q����:0 Q�б�ДE���m��)�!X��0#�)�"N�Fl���{h#ה�|��_��d
�<���'q���>�	�
#��8����?��%�F�������:t'�9UP�(��]%�>��td������i�A�Se���,��~����R�"O�����c�E����t_��r籃�zH4̅7�&}�Es�U�����h����p��5h��ы����`!^&���?���7+j4
���GV$�)�H���Y�n�EF���=�[L�*�J�-�bmCk��\M�/ �s?)���Y�&D�X�"GZ�!��b�1��-k6~|���eC���)w�8_tEF.���lFA�ĸ��F��Qy��c�g��$!�"�D�:h:�|)3�o@�Kk�
���MX���0X�2�m�����6i��u:����#h��ۋ��7$Qwr~FDL���y[�gv~Q2L"m��b������k�T��GY�]#�&rJ~02�x
x'.�`�Y�.�h
��X~�!�@�p���Fܟ�$��Z�EtB�:�J�)�?RE�T�������I�u|�,�Az�M��o�Jt�ğ�������I��?Z1S[�@�Ω�!JmV��P������ɇ��f�om�Lu��6À�2n�+�`�����[����(��`W"�l(�]�����Oylm.��	U�m��̖.���t,|c��ֿcf���;X̍[�$�&O�*���f�8�^�G��"�.��������N\��1��j������ቐ�{ �ǚ�E��������9�na�4<��nns;/E��3vfm���6B��f�~&쩱�y�Ͱ�B\���ZV�krƙ�N~��Q*���k�UVÐ�̷h���jG���L����dF�o�Z���p�Zl(�oYJ>@�z|�TԵ�!V*Չ\�K�
��4&V2�ƵJ��Ժ@M-[Ȫ,w�h[@mm"B��������� 䠳I�^�����xzM��G�޾�T���~.6��a���}l ��6>
���"$l�db�'W�1�3~����@-}b)]_|�)6�i��xT���|�@����P����t��7���:�,UFt��j7Jj�9r�@U�mO�g1"��	��^�m<���/�"���Z�=��g�^�������`AnXP�7=�@�mf��d(��r�R����^��|#��\����e�c	(�-HL��ݺEL#ҡ.���&@���]��2��\�c)ʖ��}W�rdA�(�v����>FS� �gCs�i�Ϻ�)��"G��)�4�������駻K�S����钕��쥫�;�ߠ�����
����r9�p���>c~U���av gK%~�cX�9��� Kا�$�v���>?��Z��.�N��C^l��j�	f�?�a��t�	ӓ]�-�֓ƠL�"x�]�z-� ��g8}�'N	V�����#��#�Ǝ¹^N�����Ҏ�f�
���!��=PDK =BM�fZ��w��w�zt�k�&R��|x.T�P�3�R�S�X��u}��.��R�J�]�|����W�&�\ d����>%)�q�V��_P.e���2���t]��g�yC}E����2Pg(ǣ�*f�����y��҈�=�����,`�n��rKR/�ܒ����<p�͔��i�eIsz�e�����s��$�
h�fL#��?tA���j��(
�� �E.��վxQ���`�Zd�Yyv ��8��4��X�
�����R�lM	���l!:��=������ʜ	i�ږ�$�������B"�� X�(������U)Ϣ�8{��{`�N��W;�ʃ����1삮4{��c��D��
������E����@�U��Ƅ��&��hJI�r�fN�e�U��8es\;��d�D�Ni&x��&�[��ah��_}Y����˧�d���N���|���z��"�ؙ�Ԥ��&�H��S�wR��M]��HA��	�=NI:�2�z�Te�f����������3�����k^��Ŝw��J�v�7���9�Ű��T�3�R4Q�jc�������={��ʮ��!�``���b��1j��pӬ�MJ,>�??�+�a�`�[�}g�A+6ͅxt��`��N4y���q�rŦ,�|d*̹}B�Lo�x��wp��S��C��`;�8L'�:��W�W$��]��NW�rĮ�#�p�G��K�?!�	�(L��ɤ�xA&�;�Y��u<���[l�e��S\n�AO!9S+h��z4��8]#�m������a� pWv��없a��HL�E��,�q��Z��$QU�|Y�#(�1�5>M
�ܞTb��6�3pC4l"+'�xd<��R��&�C��h�{�	�'9Z�Hh��
F�^a� �-�y���"�������ŽT�֧߰{F	���%�MA��P��5���G�r�������*ڈ��O"�z��[�u�T��� ���>�6�7��W��k>.~�(;�G�Դ�u,��j�3�8ᐝ'��r���E�{������y�c�����9�{����Ｒ���M���i����vz�n����w�C~���b�nk��r�m>��Ƿ*���Vճ%d�/�b;ڻzL{q����4�A��Unڟ�4;kpl�r�&%*����\k����N�{��,M������w�w � F��8&���F1^c�ӑ��"���v<"�3:5R�����4�c��P��Pp~J�H��}J���D�N�-"���L&
Aq��Ӏ%���6OxNI&s\�a�vU�6�3iչ~��MW��J*��dlم~_�I$;ת���HЊ� ~>"��W�g$qr��4���]�Q����X��=ˡ��'� ���H�4�\���A�ͤ]��5����+t��3D�,7ׅ��c�b�� *���s.�+�v���IňXun�ֹ��n�Y�0�8���Q����F��kd���f$~+�5�"�؀�G)ڇ��=�����f:�!����Я)g�cƅŀ\!���0�W@���Fx��;s�{����w��a��G�<A��"���a��ܜ%�A�r6�j^��z��������kS���a"�T�����A] U�(������>_�N��.�S�֯�*�~d�z��@U�7��ԦɠzV���tz5�rb�0�U�|��l�������gV��}$���-5C����0�g\5^��j�M����c+����GY�V������+���n�j��~���~vL�f+JZ�!bH��Q���cs:.��O�_��s�X�IRZ;,����lq~�ȧ16yL��D54���4�Ś_��.�#l���Sk�F���y6��"E�$<�"Z�:C�J|d�!o۳2KfR����oXcR�0s��2��������1���j��C$�hrX5ۦo�7��ZM��D��*�D�br�Q��amTܑ��o��a�FvT��NG�K#��!r��D0�c8!
��l�;{�Y��h�Ȭ戈�~J��@Tӳ�	W�#������t���E�)�;E���w��qP�P.�,(�j2��՗J\�)���\��Z�\����1�S@Μ�=�VY:>1Ë�a���������pJL����1��S����:���{��_y�c����N�=�����"��d]��@D��Fm	
�	TnT�Aǖ� 9.p���/kc�E��?��}D���$��A�%�������x��g����~�R�~�nH��ey��᮵��6���g֒B
E|[��!���$��n\�9����)N�;Jؗ���fH���{��gS�~!l��8��kC�\���Zњ�r�Nz���=���̃��XҰ Z�d�#h�h�j�'�(���jsȵ��F�	޵�~�+r����o���>�(|���P�}V%𶉷�i��נ4A٠2�EJ̦5�,d趾[�����h��@�۴BJ���y
ޑ�|��N K��8���x5o���^'Gf[
��:TR��A_,.1�1a>bE}'���z�
9�`"�"�d�.�W1�3y���f,t@�d�}X*�����i��px�;m�we��n�PG����=N����G�,����:IE�9;|U���6h�x���9[I<3n�/�=���ZM6����yw7�q���iwA��[P����;ZfZ��(aTQ�m�P�=:e�Ê�֎�\;�x�`�
d�:-;��/�S���Q�|��т���X��2<X��[��~�$��8}2� �(I=���>�,� �l�s���5����1�#4D򧶄����}� ��["�����_"�v��;����Fh
3*V�-�������\U�8��v2 Sf~�^��@ج��K/|9�5%`v��I�yU?�������\��L�l���jhU��\��$�g���-�X0��1DO�v�x��*ziP�-�f�ɢY9�IV��F�����#��=��N���-��mBf�;��X�}��-Df	�B��Zut՜ڮ����k���8>�x鰋P�'<R!�:38i��a����X.�]�ƥj��k��EWM��&�n�d=�o����> �4qޟ�Ò3/�0�_2�@�t�Tg��Cx��G��P�d�(�X *� ���Ey�&ވ\����
�`Z��Ӎ�/e��ѕ�<��9��ʳdͦI΂Ue�������K
CY�L^-\?�G�j^2�(�)H �������'�Q�@G`5f�z�*v{A�8�B��Z�����!�~l���(�!�Gy=V]������u�Uk$,�O��󷼋B}\� ��}�C�j�x�A�{uN)
H8R��v@VN�X�r烟ڪ߬Q�����=�D!K��[��c�- tݤ��p��A�0Μ�@��(I��c�-�����F簀x
�P4�eN�8���c��z��&q���O�U[4�ܷܮp�:�k�$�gbĖ�_���:���ۆ|�ZGz]���Z���\G���]���а��Z���0�H=)�:�m}���3}f�]���g���z3�q��϶^m�u��������vä1�F;�k,�T���R��'j>�Z�Ŧ&�b��{ӷ��	�Ԉ���`�bk��(���:��Y{>�Bpֆﲘ��v�gTJ�6��tH���� �N/쎁 {A�-�g,��L*GpB������wusS�9٢Hu�`��8gb:[����w��g��m=��t�Jp���"ql?�����L�R�T4�&�jPY��2u�������lhE\�!lO�_�+czhz��\8m��i� NO��a?�p���ٱ:��F�Hʭ��<챵�5�P$���|�Ui��1�ęMɄ�ܹ&�ڎ�M�5=4��]'u��76R�a�BI�(˶���	��d9�$^H��l�^cF� ��������C�꾈�)�9<�T	֢l�	�	I%�ia�Φs�>,rʹ��p��5�0��9*5�Q�s�������u�F�Fs .��9�p6���kY�bǣ����b&��j|,�"D�. B��.[��/���(����l�
亃���[����������
�C�)=M�T��X��<�vu�G��}ФJ�C&���^nF����b����jP���2�nn�dE�b��(z'Cu��S����V���(��X(��#�p���r/�%'��*��e��N�Į懵��>r�b�w{�F��.�s��܈GF^^䈑yz�`��<=��:~��R��h��x����`cַk�i��p9�HH��JO��Uc�<Ũ��M&댾N�d���r��_�O�}�$E�\A�1���6%�i0�$�Z��r�QN�*��cl�V_���;�ꒊ�M�H�� ��Y"w�BwPq��V����X��M�X��,˼6�'s13��h~4(Ռ����ľAWcl]\���%��%����,DB"?7rs���b_�� �_��-�(��'��m%�I@�X��ִT�n�D�0<�\������*�!�b�O@d;���a[����5fE�������b^�x֗c�g��T:�b��Fk��-��ޒ�����!��0Y�ή�6F�$J�j{���׊I<�����ڤ�<ܙS��@�%x�Ҝ@���S��E+���?��[?���M�u5аoa�o�ɪY{]ۅ��cd#��t��ڝ�����}S���"�{~?�ܼȾ���������t��t�Хrݎ�0�U�����\�[����X�":���f�5h���J�x�^�#:������=R+��n���DVڮǔ�5G�5Ghn���B��CuL��J���b#���I�J�e�qs5S�ª°���RXѐ�Z�Vi6��&/�c�6t<�Ο$E�Sdc���_j;.}&�l��P��2�F�<�y�ջ�ݪ-$W�"եS:�|���ov�Ka�њQ��XC�0� 2�廈��U���6(������
h-����b�7�I(�jDI��L�]�Q�bAm�d��M��ܱ9!G�T��lG���#��kr p�0��S�`
n�����Y��h=���:�~��#@%���3�����'и�tx,]�@g|)GX�EI���8�����+ n,c����r����J��:�����U�y[1�k�@��G�P�V���������Ƕ�5���8LIj��,_��M�&��� X����>}T��]�������"vݹ��7�􋠺E�+m�w	��_7�9����.˄$���.c0ݿY9v�Xm"���$"�l� z�ې��a��:��$��YV��FͰ�	��`���<�;�u�D��s���EWڄ�\H�\�nW�����MC;e��)��f#�)�@�`�~����s�&��\Ǜ|ZL��r|#��>
�B '��K��0���h�5�j=�)Ҩ1�2�]�P��F��Ż����xEo��>��F|W����G�V ���4\|H2|��J�|R�J��oh[�m���h�U�@�ioB�I��T�t����C��l��?]�x�D��ׯG������T�B���1.,U�a��}� ���
�i�"���d���W��3t�����d@�����UF����i�xx����r]��ve�P�$�3ɑ���t�,˶����@��9(��UL)�[v��z��3u<nA�/x��XZ��QM�𔇺��%��r��A��P3c,�6uBf�u�(س������wƞ�Ox�\���[���Nb-�I��J��;��W�vw�va��S�/2�&���ș�hʌ��}���(�#��L>�% >��s��fϰ!6��`��^U4�C3�k�]�8����㒋ͪ�9��J��Xb�ϖ�
�y��V5����4��U��x�ז� �z_~�y�K"�g��KJ�b��E�v�Ǵ�A1�ѓ�����:Tݹ��l�]j�� ��6S�_�3�?���S��X��Q�x��z�?-[���ݚ��]��V��k����F�#�"���N�<}�z���f߂4��癵C�D�2sBC.cZPP�珰ќk�*.����x�-tP�;4R�b5����Å�&J#.�:� ���r��+�1WȾc&���dx_^�)�d>Ysqj����UNk��W2��t�g)��Csڒ�� P���(�-%*\�D��ͬy�=������_�g�`�TӨ��/�Cj��ȗ<��R �_��I)�3eo3��"�����
7L�Ƙ?���Rj��z(��T *R,$C0���Q�`Б��uwvֿa8_f�-;U ����LQ\�l��m!���=2���|�ʒ���4$gr�3����B�09 z���^@B����V�W)EO8���q@WNM�y�](��	�'�#��ă���D�"���%@�����N��)������<�Ëd�^'��w�{G䰛����Oe)RRs�����u�{&�X4�
9[O�1�Wf���_�P�ܝ�Z(�ѕ<�l�|�Hz����;��Y?�\���T��-߶��p���䊫��=A٨�j�"�f�.�Ri,�l?33�5p��n^H����]�E�Pv�1�tr��&�T�qhR*V juE� �m��L�{�\�dÈ�
�`-��b�H��cٱ������>�e]��qD��YL���g�r76��
t�1�̖�N*ڀ�[(q��V�,�<*NB��X����w�z�S��j��M�`��8��q:�#��R[�,м���;�ZA�x
�pH�=�?���L!r����&���YJ�u����Avb&�GL\�jOW��+^�{z�(�8���߅:{��ĥwaz�cp����ԖY���H����*g�d�2�$�|Pr��h�1AtM�����	���g4��'h2�=R9<��n��C���z\����\9Я�H��-� �m^�K^ Do���`�ﾙ'�c���t҄T�zY֝}	@:'%^���Y���Bʔ���/��W��u�*���.������u�ׁ.� �a�4D�6m$p��]�kt ��Rj�����*"W,*�u�)���F�n�?B��h�q��Gq���E%י������j]�ht��%[]��k�M����8��^:vp�$�F�_=�CA�:��]�n!���-����=2�U�N�)�%d+z�b1kaz+ɼ7h�j!D��q��U����,sp�r�;�%���[� B�N�-���=u����n@w�SEF��Ԅ����#hs^YZ�l,r�ݮ<X�o:�_�RŸp�)}�C+cѶ²ę�p�}[H'�J�2���G�w+<�1��& ����Հ�/��+�On�|���\|������6��i�˅w"�bV�_�*��rlO�B_$�m;�J�;��HF � �bE"�dk��q��E�j��S��x׊XEr_���"'�ar�y��4Rc��=')���A��]R�ɝ���c��D}h�7�G��.b��� �K�H+�!��H��I{G)X�?7֯�nOP�0�c��͘�u������0��d֋9�\���P5!H��-�q�=J��=k����ܿ�:A�[��]��QW�Y:��{��!	��0��ծ�F.����{���<Ś�"}<w�[�9M�e�3+�[�w�h��� ����]�������\����k�䨊�����]�r����E�0�(��8�r��S��)���S~] W��� �V��LYct���rX������6���������f������7�m��{�5� �<C���^��E��:�<�+����=�5V��Δ��6���On�Sǡ�ц�n(XL?BJP�b��Ǥ�[7� ��s0�����W3�X�� Z1��DТ������X6oL���3v�_��IW_�7.Xkl���ĉF|�y�ȕ�0�$rL�"P��:��
|ڔ�o9�K\~���R�X�S�0�(-2��K�#����Y�g�u�,���$�h�o���u_7�TE��D����Ju�XʒQC�m�	���KB�Ws�7�T8�>G*S�#���r[V0c��n��
��ν�YF�hإ��~�~ �,@�aE����MF�޵��Lt�"�;�)���EL.�S���g+��`,���K����GJJ�7Y�:���PC��T�#1��@Q-����V?%��F�l����p}�� �zL��']�	�F���Ѐ�F6�p9��s	��["��B��+%�����m�%�	� ��"Ė�(�.&�Q�H�cKf���R �3��>(�$��Ϧm:�w]��k��U�ɂ�\��4J�܁<Ϥ��[����a��0@x�쟺�8I�E2yf��,�Z�nR�wE��ȟm�;�*����0f�Z)�df�����~���W���x�\��Z�3rWδ��
�ݷ9���g�f�G���h�"j�(�H�m����F�`��k�X�����P}o|�>��|�)�Ԇ�Vo�m^&�;O�4w?�2�ىJ�r���ngH*[oj�=Y�h�,�@�RB@��/,��K������#r����x���q�G\���H!T�	Ԭw��.'��a��l}���cr
/qH"��d�(Wg3o���U@F4��]Иyͺ��i1V�x%%��mu.��|7P� �N#�D�I��d,���pٔ;��9�#�U�P丠L�ncj��*�<�4�/��k�L�Z�k�s�%�gYV�M��A��P�(��1�&f?(�{������3��y>L��\q��V>�*-yxc�e����H3�2��G�'���N¤2�"��^�ȴ���� }�>�?�(*���%�>W?b ��#s �s�+�ޞl��ܙH�4z�6�z��(>�b���+��.�}3@��N��q5���}
��ȣ���?Z���U�bm�� 8�~Ѵ���C�"i2Ke�T�+��vgT��������_���t#l��ij^L0��1tĚt��̓N�E���}M�x�V/z_ݓ-6����m���V�2����ͰT�#ҀR3��Nj���M��	�f��#�.v��3D�{zB��SZ+L�P}��K0	k�\&�� �x_�@P�o�R��e��&Fx��f.�7��[�3����F��WC�[&u�d��`��ܸ>!Nq�L獐�i#�&<�2��t�g�"3Cn����tGPI��(#�*�1�ݣu�y<M���}[���$�`�hM�Ë�/['����<!8o�핐Z�I��e*���=u����
�4�L�i?E�n
6j��(;� E�����fY�QZ��`k��p6Bv1^�8Ш�Hܗ{��֢���`^l�d�x!K�P=�&_�	)����k3�$�L)��'�FB3%� 5wX�y���nRR�1�q)��8LKA�l`�N�Ǻlh���~ߢ|�������DW�����9Fv��vy��2�歬�w��^��Y݈Z���6hE���,�F�?e����5�9�pq�&'�'��ɠ[j��қg��@Ě�����Ut�����')u|�V�z�s�i<*�Uu���(/�k��]�@2����"�&��=���� �%1f|�����'��3��
~�^#H��(����VRv���Ͼ��ỶT�@sR�ej�v@�;ɟ�1�{ɇ{ʿ�шRm�`HqTbF\���!L���A>���<��GR�BpgJ�o6^-Lt��[�1vN%�N��� ���,���*=B��u�)R�wA�MS�����E�`l�i8�8�:���� ωg9��oR��)��-�p���X�?��E�f�L\�~���&�(�Y�D�um�*�oݚ�"P�\ =O��+Y��zE�)8�������&şT�a��p(�9�ϛ�ro�H}	��B�⦟��y$�4|��851�C�M?����*�ڄ4����4�^'�-(R�6����^����������9[�H9�+��.^q+ �?��HP�9�P�>5F����TT��֘�Z	���%.�-Ӳ4y��o�K#�D�k@��q3*뚆�����z���[u���i�� R���/�6�����ϔk��Ǚt�����e�,���$$iᡱb����!1��� �"x��0(i�47c��@�Jg��#�$�@����SM��������r�kvkt0�P�C\\�nn�s�#�,>����0й�P���dFςb�cfz�2m�F:���	��/2ڰ3]�eU�p�[rr%7%�l��<'�Л�N��w�=樨�Y?1��wq��Fg9���ܾ��^TlG���	��A<s�I:t9R��(�d������c��U���p�G2HB��JE+��՜���Z��̹W&��ؾ�&�V�{��O�<���'\�魴Gz�6�n�i�Vq��V��9�D�*k��l��B_��v;��C��,�Hkq �$�"mjw���9q0i�rn�N^ƖӁ�X h���px'i�}�T4��Ì��u�ЬA�]�Ґ��5��� >�nD�ο7���̦[b�� [W��c�5���b�#q�I���XFس֪��n�{0����;����T��A�k(dq�&�W)r<]�5�'�),���\��V����k@��E:�E������ �k��X�VE-!D�0��T��nF�]�l�&{��׀N,�b'��P��<����r<���+�v�������$�+pe�~���s�+���&뫨��c��R]��x�٪��ņz��p�=�-YoSч/��~�P�>��܂��Xɱ#1��Lt�f�r���濷�qh)��+�����>ʨ��RoN�\�5Թ+�w��8�^�^9|��}+�8�vrV�V��4���k��n������ҽ)-L(��J��bپƤ�E���s+���`�R��1X�Z���D��̸�P6j|��Ucǐ�y-㻱_`[�.3��l2�t�$"?Fw�yGj�S֘$���"ˆ7:Թb|�3o��|KWD	��X��{0�p&25n�q�	���<�һ�T��h�+����@7�L�U�D8�C���S&'Q���m�P���i���T�HTs�G�<#��r�\0�����
d��N
Y�KKhsę�y�[~['@��T���Ƚ�ސHF�t�`�6��)��jE�3��n�������d,�+^�����JmѤ����UZ��P��/s1?��@�ƾ�!Vj�o��9!��k8�K�*�[:L�r�"{Hd�,��� ɪ��v��G���?��
D�",�K�I?O�*�q�;sm��^	z2m�f����.���`�qcf܃�O�����y��$X�j��6��w��J��pG��Y�^�ܼ�U�?L�V�d�������Ȓ�`E88��\6����nM�P�M��Z�#;�an��1f��M����8��~���I7�͜C	\��ZBkxr2-��:?�xo����������c h�/Gj3٦�W��</Ȇ��F�� ��V�\���H�o��=>�n�|����!CcVSE�Ⱦĥ��S4�"�2r >J]�<��?G�@[{�����hG#^@��\B�Ls�
�������h����xf���*�Gא���LT�l�kE."ylaO��}X��/T
��^"�ldN�fWX3j{�w�F@̮Υ�K�͕}�ilSnx���h�`�,��Px�@�i�2�m}�i.,A�����6�%9ޅ�U�d������k���B�<�G�/SM��>Z^~���?��y���(R^AZ�Pi��,�fk�2(�?��:������Tt����\U��Q��u��-4�Ǽ����12������:��g�I�U2M#���8��ϣ�ʂ�V}�P~�(Q���>�x� �:�s��Ϧ �G8�Ԓ�4G��u�t����Rm�5������XM��'�J�2t�Ŗ�
Dx	�^, �B�*��Uf'��M7� �)z~�Ic���n�K�S����vBı�*�s&W-���Q���c�/��l�j��K��L�Ս(�uQ�I���B�8i�x��z���-Xd�S}�ؓ0�V���W#�t #�����ZNE����r)�>�f�pO�i���D\D���B9'�ZhϜ�6���kծz�I��x��P�\R��n�,"�a�^�\� .�T�ƶ?O�I��a4�W���&Pd�d�w�_1�>	�q 4;�Kۘ�M���L2i7tI�g_�CiQ��X��P)(38�*R���~=�yw��-( xَ�b�`�Q��ދ�/�*��b�<\8��+sUHRI�[pe��r�X`��-
�R
LY�?��n#6jo��(��Z `��V#�A"cQ���`Iu�k�v��8�Y�c�"�lm�} �O�l��P���!���=�;�5�ʈ%�FR $�F�i+��B�9� ��ؔN����,�s�)�� 8���g�-N'��� ��Bu����O�D�1�����t��15��䩢p��ͬ��1���p��T� �&���
�� ����We��)��Y��{�k&���耕�[�N��MBu�˔����3n��P���K�L���|�z�ё�D]Ԑ�Kǒ얣�k���İ����;@=������_�fwD������Q3"f��!^��&�cJ��{��v��é*+Ŝ��T�/R �UjϘK�v^8�36{�7�! ���`cK�b�c���ʱ\���H�>�l֗�'�LU���g�#t69��t����P�N ����^h,�|v*���Bb�d��w��S�Ă�Y^�`'�U8��J:y���҉��#�����.�.qAp�B��s��?5�|��L�z#�%'�&���Y �7u(6%��X/[�s�\Z��O��,+T(�z�;`8I[�Wq���z#a�vp�|2�����3�H8Y��(��]�f��&$=jp|���(31�2mM��
�
]F�����CK4Xc-'F׮(�R�P�sV�y�S�p�E�ut�9F&H������^t�X �0��P�ﴐe�����^T��֓��	��c%�|ڴ ���|�JQ^���I����*F6褪���X1�x!�uxYo��Q �(l�*�z6#��Ca�k����ʖtv�Ԡ��,`^�ֆ���6��%�<�+�g82�����k*��π�����?�ޣ��[y(��P�M�j��	޴��5vfUt�[9�Ղ�Cw惟|��n��׬^�_�����C*��G՟G7daDb'|7z�Za��]�������ч� �30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮs�
օ8�9�$���q�|:]���;~"喢z��l��&[@	Z�H�đel+R�U��]��iu�V�>�5S���f{SN�:D֙��c0���k:�lj���n���L0T��O@�x�8���k�m��?"�]V0|{��E&쥆��kx���?)
�Wi�x�l:R���E9�	
e}AbP71��xS����Ҽ�S7Z������Q�,+��3�4dԦtrTF1%�ߓ�O�e�����`D��hG� �����Ğ�.:�Ij��*�V���n��b������Br�O��F㝰rr �.���Ca�����q2*p��h=\�J�I���I�@��Y>��f�{`��RDR���38��WMf�SU(� &�������� �!R�Ho�(�Pd��.npu�i��́�6���3�k��;�J0 �ya�:s�߬�UQlq�>R�| D�?��g�yh�,�z�K.F��]��SR{T���`����� �,7��8`� $:{�S�Yg� �J�w/nd��-Zs�n�;�`�"h��d��Q�K������5-���}a����8��~���K���ĺ���i{� ��k����Je5� ��"r$mY�ט`�H��8�mt];y7�����ą��n��a�*o����&]��]NE2z�d���ؼU��n&B�S���=��S��VRi>s��$R@��a�f�ʦ��_�Y�4ϖ��,��'Z�-%�/�@"b./�W�¿�Zdgެf҂�oZe���"��I�A4��9���|��;��&�o�nSt誹�R.� ��Il��
؟�|�{!E��E|Q�L���%)�7ê�ICz���^�;��e#��$����9Aw�w�W�ʚ��_0� /Ѳn#&�0��@u��43���Ԃ�>W:0X�tUa���o!FH؊Ew�kټ��ϱ�"���:,�j)�+�,X��ϊͽ��ԝ��;��e��G����װe�� �)a�h1VK��B�r�����Y �v�QaUc>����ቱX���q:��ie��+��R��>���#h�Pȅ�o88���9�-��7���9�i�0�a�e��ܦ�z�71�-�*A�ĉ�}��]�әme헽*��h7�lM6��p?m�a��~���WW*�J�^k�WML���mSi?��D%&p�);��
7�J���L�#Q���m����Y�Ǧ̝�D�޳9^��h�G@jo���v�xq[�����j��5�c�RW �������xdx�P_EE�T�v��!�a �k�%j9��
����Z\��;�	��*�E��\���g��b���(�'�Z��׿B-�l���*OD��Z��_8�se��Z���ް8B�D	jB������PY��dFy�%�H�Uo,���~}�F�%S{���K)m[y�\��/*�nh h<?�>?h�@�	���[���������l	5�P�v^��hFK>� �CZ�Y)wI�N�j1'5��8���K}Џ���@k̐$0b�ϫ�'˂Aԋ8sl(�6\I=�?}}�P"__a�i�2v���b��N0�<�6NƮj;V�&}�v3H�ׄ�
�8��.YW���h�:�X��ڑ�*�v��v[ٽK�`����_3��uq��-ËRH<LH��4&A�
<�@���up��2�Rb�t��z{*3�{����Eb�F�o�B�n�i�w��?��7@*[�r��s�<���9��5�*��F�w��|���3R#mQ�5G|H6��*)}������ގ��?M%Q���=#�1��T;�+$̾,����*��É��0zB68�6�وk|+�S5�e(�}w[�<͞����F���8{P]�:X��%)F�R�F�~s��Z�y���"�
)��!��҇�`��V8��+����CA!$�o~%�T��\��U18mpc��"�z����nH�O�3~�Cp]���FZ(����c�S����r
�q<��Ǡ�r �Fޥ1+��^XK��w�	��A����^�"4�k�����mœ��UiH�$�Ż̚2�������������,Um�A&2���?ǆ>�}�GD`[ȯ������_�j�΅�Ӏ�T��;u�N�G9�qLe���j�5�#�b!�ǘ�  �T6�)��T��a��!r�����.̀!	��f0Gw�S&r�f�%��"���:����ݿ�fo1~�5�!/��o�߀r5�M
�N"��J�g�8b���-(2e�����"#{b���CL�s����= �zΦ5�%��0���b�z��L+KtA�v��ü��-�D��[
<.|�@T�h��YJ���m['a(&N�6- nA>wFc��.C��[���)X
c��+d�T��]Z�:m�(�:2G!n�p�X��&c��*� [����t6m�=@:�~*��p�;�����a��q� b|�=��\6��R�����w�ɘ<�
��o�/ʖ�16{H&r$��E�$8<7h�{gia��:6�ĿӲET$5ɼ4A���-�Nb~\�{�����&l6E\��G�B�H�˩����U
~���c����sq��KtF��#�yz X�ↃP?����J܎���+��<������P�{j��ɿ�W2��(]�G��dj0��w��3v.�)8�4 +6�2�r�-$D<���*����Wέ�������|S�6��%Y�Q��g�,Đ1���C���"���aG�#�Y�+���+GO	���3#Š4l���&ˋ���`!��!�@���N~l3D�'������DW5-{�N�2�@��e����16V��7C�{��_^Қ�"�P�?��ϯ�i�h�Z���"}�����8K})��a���K��O��ެ�9ox�&R�om�J(���i�5��D�@e;��N㳞�/�}�>�ZO���Xx�C������F�N��3ܨ�`��6���;�I���I ���������u�j���ب��9��:����}��-
�u�7:u)Gx�F�|O���W�Bk �gΊ�
��?>�\q,S}�O�~T�����e��u�)m�)��lj\���5L����٩.�N��#)$��n�+����z��mf��	v��B�ɛ���ȋm��j�;���GĩW��:��U�YZ8k�u�^dF�]>5�p���s�bj��K�8�ݠǟ����Wz�k;��r8�a�jv��F��||�r�\������9L�������	��>Hֿ�����RY��in��V���5�l�*0zP�ȑyS֮�c�;�����k/Rxl����0�IROUWx:hl�gkь�O��X�|P?0E�O���x� ���
�m>i9�ҡ����2sE�
z��J`aU��נD�����7/_�qkM��p,��\M����?$R��q�
7��=���,����,���2�_�� �f���u¥�nf�>�_>!�LˤU�J�ެ�h��ec�9Gzkm���v�����^?� �3�)�XgQ%��\��g�0�(s	�_Oc_��r��>�o�:�f"/�w�+�r�Q�2:~�X�����c�:�)���xL�9W�&I��?��y�����Xȣ������a
�"��x�1�9g��&�GU�0bCO1�at"��`3Դ@��#�;�G<<aH����}Xx ��Iz5�H�
��Ƿ;���%SX�9�(L�y�6��V�}�H_�~mKM�i�9`�����	u�A�>Bn�u��易��,�p�'�8�/P����US�������՚�!��E:A	&I������T1��Id�� �{1��'m�2}V\�����7�hbVȧ�s�fM���+����OV��l;���h!7ć������Qy�^���i(T���4��9 �}�M_��_Q��֨է�B���,��
����_%�}vH�BI�wO�c4Nݱ6W�����M
~6o����2���edN?w���gWǼ�\���/0���1���=d	 %d�|�Ձ���I/�� 1/ivZ���ՂI�7[9�ʾsiG���,����^�>x�]�S.2����]����a�
l&����b�=tݪW�E	�	yrOfpS ���C�b������w��S��+@^ɱr?l�0Q܄��,#�&6��,��)�������PHgk��v�Z#��̧�eq�2^���=�3n&�
�Jom���F�J#k����s��t_�+&gZ�O�8���Wy-�ߏ�!��sv�� ���{[ɄZ�jM气��*3���å��:![q��2�aY�P��M�au�����Q'�UJ�<i���v?Ib/�����ߑ4 �U�`,'���,��Yys[[�H�<����ݝ�4�п٘C�����nSR�~�r�24��1
F��H��g'R�:������r���H�s���iɟ���Q��v��`�`��-Ǌ������'�S,�*�]�zZ����BF9*#�y�.�z�w�s�<�J�R���|�h#B��n2TboF�0���X��"�y���ޔ֫�v�� �@�i~*�0�&�oA��b.����i*W���i݁��۵;Q�7�ޠ�C��'D��,�����_�^���'�b&P����e�C"���m3���ǝT;���94^���P�iuy��79A��ժ�i�ɣL`H���L�ǫ�N���g]�xIg�����g�[ŷA��N%	2�����@kI�|����>���EXq�����b7u�^�:C�S���q<�ã ��"����:4"�rq^᝿C��pt��h�v���YO	īS�p0�Q~����ӻZ��\��9J���Q�wjJ~�,��^�&���%J��W� V�|�_i;��w	�+Uw2��$�f���lԍk�__�~�dźʱ�9���Ge9ck���4zleA��l�3T����Ɛ�8'�'X9*��~t�`g���'�F5Y��ƔD�04#ء�O�B�� ���cp��󵘚�leI��$�����.�X ��NE@%��f��vz�2�~.?/�{ف��RiH�h�9����l��4���������^ƙ�'�`�9s�~���{�p�����B6�ƝuǫY����wE��Ij f������Ș�\�eR�$R����.e2K $��E�t�o3��u�z�U�[�c��N	� o+��y_�P��ǣ�*H�!�z���3V�C=+�x[ԃ���������4��*�~XӢɡy#�b��`ԵX�ys��f>�mEq}�.�Qُ]��(���?n>s�\��ē{�k�|�E8.�ol���@��_�m���R�)�/{�x< ����]�}�Uj�K���Ȉ���J�i��y��4�|����E�U�|=;k�'��X&���/���������G|&��`��|G<�?]��/��4+���*���	��zc\<�I�����O0���`��u͒	N�N�۷"�ZN��7F�^��T��{�����:ǰ�
�V@��sS�P[�hp"�5ٖ{�eFd�_9��9�2𒀶��~��#ሃ�J�B+�Ӎ�j�s�Ů�ѭ@�i<̗��)�GpJ(���43\&[�W8A��i>��������	�� bO(�z�qd��2�����P�I,��6���B����_���q��<�T��CGnG�K���L��?�W\]�ZD��/یdX|N���z^KBOYЎ�{��L�\���%�fLm,X��}@����JI�������%����k�8������)�z�/��_R]���[4c:K+��j-�M��ā�h,Q�*u��W�فtq��a���0�ٞ��}\TWf'��'!��q���F�*���SV�;)fˎvK;�@x ��uǇ�c�Va��:����8� �Ć����ߓ��/���I��vR����OT�U���qG�u aR*�}_�7�^Bg��(���O�x���,afˌU�ta-��r6�g�{�l�T����4 �A-��+�t3��A�����c�"ݙ/_��A^!ņ)�a�]�ޠu���R�ή�ó��3�]Ix�I�(������u����m���,��=��0�6��(YYM)�|��������o[c�����t5�f���L/�V���j�<P�{オg~���C� �3O��pP�nRY�g��da�![��`%����j����*%M��'�n?�M)�6��G�7pL�C���{������E������6��Li�H+�hg�����8�1��у��1��d�&���gx-]����#{��VK�ŉ�"��E�B�x��j�m=�]@bF"O/�2.���7|�������OvS����қ�ХD�6e�A�7a�<��i�N�kȅ3Xz�4Ҟv�D�����P����ѵ7�y�i���}����V����R�b�H�'/��e�Ŗԃ|�_�h��䣅��F��z!�gM|phW�=�j����ź��C���9��ՊqV��Ra�&3n��M��	L��7��������� �;oR1%��^(�d�Zj$�+���qͷ���ʲS�!i���0V�yW�:)7�i�Q�]>H8M�j��g8��y^�I�0�~K��ʓ�gSH2T5�}�~e��E�7?�i`ajwpmS��:ضf���c�d��-P��n8�0`_�p�NK}�z��Q?��d-���6�-ˉ��3 ��M��3ë�O����L�x�ش��k6�N?��5A��(��Y�O!����͹�#���:�����	�&���vnp?�`���M�&]��%>2��x��pe��n���S-�Y�3�Z�	�$�xC�it_�ul@uu�yJ(� n��UTk��;��^0��:��Z�樹�;"�����,���Z���g���f�%oPR��@�g"x����4̺dӸ�q|&���D2o�S�t�.i��(U GpIbI
�r|hW�!{��;�����֛9�7���I9���e��s��<ZF#��$R&�֯g9���^��6�D��0 r���b#cϨ�#�ut��4iaL�ʴ�>��0΃nU�Z7����!�#y���sk^�������W�L��L���!��X?Ǔ�C&8�K5��;�߷�M�����צv5܄��)|�7hg����6�rheC䏉ۉ�Ev�P�U�@�>7���%�N��'���s93[�����0�>3��#��P���o�1����9ͱ���b�B'��_ϜA01e�^-���ᘭ<?�c/*7Bˉ�]��4���e��*S�|7��6%�?c����b�~��W`Nu�@�.L�?m�2*?���D۱��P��[�-�ڲ��L'qn��4��{���>�B��z�����^ZYE���j�����.���&F<��g��+�0�(� _O��!��n�xP�^E�� �z���u��< ���%��1� �.�x�~Z��1; �u� �W�=+A�K�,�%�9��F(�a'Z*
?�x�l�a��s���Օ6�i����� �2e�8���:�Bm	´.�.Y��Fo]%��u�xob킁�����S�ҁ�D[��\�1&����o 	�`?�e�h6>�	�a;[����*.���lB�d5��vE�h�^�L���9#�Y�^l�aΣ�ޢ5�)*���g��%�[6ʒ��m��E��'Zԁ�`s"Q���T=n�s�)��Va6t��h���⯪�����r�lRǮ`�w��f�v�h�׺ھ�.��.,s�PԞ:�2��в���i*v]�[���VK������}$q��Á	nH��'��ji� U_��QR����hb�b�ճ��f�*�c�5���b�bbso
�n�Űwǣ���y�*�#W���3<��y��e��F��x3w��|~j�ɩ�[I�MQ�9�2ˌ���Q)A�%(�j���&�?�C�Q+p���m# !��+q�,B�Zޠ��ÿo�`�6785<�پ�+��3�}�+<~�d�FIV�8��]�����R)�����#s1X�y�Rʜ�ב;(�2�����+`�$���4"�a+a���LC�QZ��z[����YD���1�J�p�p����z<G��䥡����~��l]i}}F�P���u�I6Z��\��_�
�Sc���(h*FT�+���XAn�w�
�\�RA�S��TEb�L��Ӥ��m��߮�㠚����Z;2��l���~�?a)�!�]mv!F2G�?�|>�cG:K��e��7s�_:7\�D����GT��u'��G/%�L(��Q��Yb�!���ⶪ�T�x��9� ��x��g	��d�!�j�f�'��K�rS����Ѩ�~nˮw�d�p����2�����W���e���(�
M��+�	�@`�>�i��-^Ă�v���Fb3��C�����v�a L��R��k�֯Y}0t�0bwǂ�_t7��0J�Ihf���f�]���A,	�b�	/�mb�7�I�%H��3EEٱ�N�b#]Ɠ$��ցB޻���C֤0�eE��|�#n�u�5^ uFK�4{�����>���0�) U���/6�!��w��Hk!wQ�gҫ�j|�0��^��s:�X��v���VZ�cVk;=�K������<6�9�)N��hy�i���sr����aE ��Nv.I�UcC�>	�n��Q������1�T�7K[����.���>��#��bP��o��јɵ�9��Z�߾����ݱ��S�e�D�1qߘ��u;*��@����������ye5K�*��7��6#�?����?Z�P��Wr�ڐ���!L�K6m�"?"�7Dm�-�q��	d̺�D�L�X��%���?�㽡|ͦ7S�v�&�<^� ���D3j����P�����x5��ܸ}�AךA� 1���3^i����x�p�E�� ����WS"4u ��C%�o��R���
�VZ�r
;$a�r���(͟i8�7a��f��(ػZ�Rb���l>'r�'��w�է�Q�����3ӣ�`�8
5恌��B��� �sY_�F�h6%PUy�%zot4ǁ:�Ǝ��S�R�ғ�[I��\W��\@���g [�"?%+�h��	���[��`i�ػ�lT�5��v�|�h��w�^�`��	FYq}��#�����5 ��)j��յ�b��∐l����'����ns�l�~)�=$�1��j�
a�!�z���	��)$dx �~����Bh�nm�v{A�������_.�+X�"�#:�^�"a4�]��v/�[!���Ҙ��(�O�q,�����HO����L�|�\�R�ވ5�н]��zrb5��G�u*{R����=N�b�r�o��8n���w�\�*H*��v��G<ٝ�f-�} ��m�w>�k|���{30[w�Q���K�_�)S��η��d'��*�?��7QV�_�#�M#�>Ƣ��+lKX,�j�rG��ђ��e��T�8����+�ݰ�X�}��z<C�IyF��8]3]���N�$)��3���~sC�Z����.���coX�D0��_8`Y�L���s���N�C�����Bm���'���&�41_ɖp���T%uz�,"�=���Q�~�#]��F�����ٹ��&����1]8
�׹�%�ʔ�82F&Ǥ+�6X�M�wd�ܠ.�MA����}|�s�Z���%�m�0��-W�lXh��k2�I��DYi��j�3�m�d�2�Zy?[�j>)<<G����5��	l�_LJ4�ƫ�T̞du9� G��FL�������kg�!"{��H<,T~<��K)��&yj�ir/����v�x!QD�fx+E����re�>�N���S�I�������0!	߮�Ʒܩi|��1)���GMf���PՒ�CЬ���-p�����j{�b�C�Ly�5VΚ�y���ކ�}�دm!�0��b壍ǔ}:t�VP�м���uƣ�JH���AvmF@����_*�J3�k���ap$@N��
-H����*w�E��vn�J��[ 
&�q]c��d�����&���(>.$Gi�p�=�^T�c9W��h����.rt~�-=���~r�p��ҕLa(;��a���hsr�d=�=a~���B�[��������0I/M���N|�{��M$�R�E"���>
i��\�<j�Ӏ����$]:A��`��iC��}&~�V���_�|6���Ï�NB���m�~.~�)c��X��=���U�D��y�>[�*��P������ֵ���t���:y5����j�B��2<u[�yҥ`%Mjx.�w�#�vvt0�) s��2��D�u��D��=�rm�
E�>C�-"������L�eME�Y*�XV�tyD1	����T2��/��Gf�Y�s�?��+�̡��2Q3k�M4���S�����A��tB.�@,ʸ�l�3�vS����(n�D���!�N��@
�eUM��]�1~�"��P{U�oC���pߘ�6�N��7�hъ��\��<��)�~K�=�������F_H�&�L9`p�x�P���K�������}*소�7e���N+}��w�����b�p���U7|�T�՜�ΎN7�3$c`��8����]I�}�]�" q��aZ��tu6���S��IJ�́�:'l�d�f3��uT;uKZ�:� �G�>[F/�8OSw,П���	gg�@?f���\�yS}��O�=XT�TX��)���)����<��\��b�����0�!����pPt�)lu�n�J�ݤ`z���#Q�����ț�=��� ���K,_��M�����nU/c
���ݽs6\H���5��@�J��jVk:K3���
¢���W�:����d�8���j���ώ��|��^����8���3���]X�t\	��HJJ�"�iRW���Z��i���V�<50�5rY���p�����#�c-�y�?�(kwQlG�	N�p�0�oO�#�x�����kP���`����|�!�E�zކ.4�x1��*��
��Bi�l��"��݈E���
���_/k��F�
����d�9�(7w�:�&[�\�5,(D�M&�3_�$���q:ư�w����ĺ�x`,2��z���0Y�����Ppq����>i!��J��Ӱ�Nԭ�'���Rk�U���2y��^�)d��HF��q�@X��I%�F� �}�x��p�����r�	4ѷ+:�dw���s�)r�#Y��C~�2�מ[���:%#����L���n����\(��c�������/��aM=P"�C`�y6�9�b&��E��w�x�?Oy�Ea�(�K2$3�p���;Z!(<��4�$Q���җ �QX�a�HA���L%;F��mc���^L��~eV#r6H�-0m�?.�\X�9^8��`j:�W�a��چ�t��������8�up9�:��F��s���uS���V���O�U�l���AQ�q��U�
8;�F���0�(�S�;�#J�m�b V���Zh�a���y���{�Bd�s�¤ʆ"V8מ;Frhi�{���f��qQ��w�(����|n����}�پE�����wBF�:�te
D:�ߓ}�K;B� �OYN%PhW
{H�79`
Lגo��:�o���d��n�E�VW�_\��U�Q���E�18,t� dX�o	hSY���I�ɓ��?3e�1wr��&gM���}E��F�C���˞@Uo�WZR���c�S��ʋ�6~�"��p���=Mt��ZҖ��CG�8�ʈg-�P�,7�#E�R�-3Ih�ň�V嗑QV�*X����7 �W0R��f�9�7d����2�ڰ?�)>���.�5A�1�-[�"m�;q�_
��j��ן��`q�����(|�ݥ	M��i{K�9���'b�Ш�d���l�?�d*��%=���W4�%U���'7��,��y`]��ݣȾ�ª��4�٥��Ƽ�n��H��k��￰��?�F���^�3R�5 ����Be�����s�x����}����#�É��C���`��3-�cr쟮4�ب��� ��)��jT\z��\��B3�#~�ӵ[�}z�A-�࢛�WӅ��d�Q�B���^ߙT�������e�/��@wS�U���cm� F�[iEݯ*�Ⳝ��[A
��.�K�ڕ�VwmW�$i<�̝�;�}��	CC�mzDI~�������{䰿'ˡ+Pkv�>C�y;Ⱥ��oN�T��0�^���PYܪu����{�A3�ªֲ�j0y3i�����N�[-���Bx�>��~�>W�����[�m�F%f���H��UI�ڽ�&
��2u��ox}{�W��	P�luh�z^�5���H���O����K~"������E���^�5�C�L3p�c�5�9�"�EY\�� ��0u���޼`�1���9��q������QJ��P�y����V��9��J�$�W�VЊ�_��ʾz��w�F/$
E�ô�l�7��x��_��5d}㱺E�vѷ9�&��yU�l�{k#S�����fn��}ay'�9W(�~A�t;̊�l��-��>�Ɓ���7i��UV�� J�I�pr��7�爼e6�$i'��:>.�� ��E�߲S�0��zm�K[�\��tA��Qh�v�8����Ǉ(Hc�xz�ٶߗs����+G��g���D�6��79̘�XN1X7�С]��b�>ԙ�,y��f"AiE�9.��ď�N`���棼As|w?�p;�{��|�%D.�\�NNx@l>H_Z�ň�X)��b{��� &�K�A����[UN�;��$Ĉ�;t�{	�M_;yV�`��_}UqzK�%�'���&	�/i�c�qA����~G�T�D���I[�<��]���/��14��f�ѓ�g�	�U���ez<ј���>��5ƭ���d�1��
j	2�����f�jH��̧@:����t�����II�F�ώ���6/��A��U��M
2��I���u��3Γ�ҳ���]T�D�U( Q�������`*�mМ�,D���v6�7R(f��M.�P�S541�0��`cb����27����\(��[4�:�P�����m��|��;3]3oy��w}�s�4�5�ԩ39!@�%`��U�1'�jIj�܏*���`n�1BMn=�6s����&�h�%�u�{�K������Q���6����J�HP��g�	���g�1����[p��ط�y��]�*���t�9���T"}Z���~��u���t]e1"HM/�p�.�c�7!��*'ꚃ�O�SE�����F�DU�!e��h7�<�m.�3N��
��0��c�CD�D���@D֛���|�X�NaH��\�_%V����Ik�b�	���ພ�YB�셰��	ϩ�������ԥ��p�F=�B��nn��T�Me�4|:�_�����Mx�RF��3���rC���˗����ʟ�C� �*R'���f�d�i�t��D8�ͼ�ߟo���f���ʭ0���y|SQ:���Δ3Q���>�&6��p�bg�N�y������K	0�ʘ�S��]Tz"޿���;S�7�J`ƕru��S.����y�ҹad��-u �n�k�`�b�Sd�I�Q�A̺I�*�c��-�Aq��ܑ�r���8�}����A����<U�##k�Z���~5	RcI
�m�Yj�.�F���/��腎����Yڦ�����nU����p���&����8:M2�Uj��2��P��n��aS�p��X�"��,����iy�ϻ��@���^�̅��z�{֯����n~�?�DZ�R��*z�"���D�i�ݹ�Z�RdgZ˴f�o����N�"]�����4�Ŕ�}X�|s��Ź~o�i�t�����;L ̅II�eP
Sse|�T?!�K"��1�G��րa87~�LI^5�*>��)C�A9#���$��4֔���2�h��@A	2�0e����"#��&��L�uY�4�����Z>��03@nU��.=�!A�f��0k����:Kc�ϱ)-�Q4H���$X��Ɋ(�0�<D=�6�;p���w�t|�K�6��0 )ap�h�Pб���r-����h�� av�9GU>�>'��gO�s�g��Z��c>PM�9~͌M��>ce###
P�o�> �\;�9�΋2�������/֜��eջ'�d�'�wE�h��*ܩI�ǹ���b�T��e��*��7y]�6�t?(�����c��W儠�Gw���Lbzom�#g?uwD �P��"6�|GpR]O�wdCL�j��Aޒb*�T��'�S�{��r�^/9�f9%j�:B�2�_�s�^�e����P�����s �rȡ&(����x���E�3��*MsgO� b��%�|	��7�� \Z�>�;�r�E:|�����>�*�t����(��Z�R�� �lg��贁��՚e	��a������8}	D�__�B2���%0Y5-F��%tO�o�˟�����USV��҆�[���\
 �o���S� .�T?X�\h���	�/�[e�������v�l�(�5�g�v�� h!�D�Q���ކ�Y$7��Ạ%�\5��#�\3�X�C�D2�Q��y�*��'��gԦ�$s�8�%=�����ca���6&��:ê\�2ּ�q�O���!�v����?�"�SV�.�}P��^&:�	h�uj?�5vBO[��e�{MާR���!�q�z�&��H���ޅ��%�~޻�\�P��m�Ib�7D���@*��66q�1b'NKoo9{n�;Xwl�5�݄�*��U�~� <���ۙ��%�$_w�o|��JɎin�o�Qʏ���o���)F��g����o���:?��Q)�:�V��#�)��.�+�&�,�[�ޅC��D��8`W�;�8�ٶ��i�+X�`�n}��<�B�˹FP�8��0]�CBʡ�P)A�㒡`8s��L��a�Z��{�76Q�m#N`���&���Y!�!�C�5���`�g�zc���/t1rQ�pT@�'� z I�I����ݣ~8��]�0F�l.�@`�n߻�H*0�ę�
���x�O�m�LF9
+eEXfl�w�����A��>���E/���mV�����m�0�Щ��Z@��D2+=������$��ۦ��m���2Z�?���>�GG�}Ȫ�0��n_��CB~�NW�T_gu,��G�,TL`$ҙ����ރ�!�%t�{AT�T�>G��yU��ٙ��"���!$?f���sOrXV������TǮ\dݓ�L�����&JY)e�\��
T��m2My��	J��e�M;�-c���$җ��bu�CuR��̚&�V�U�p�&����0�Mb�l�i�t\��Q�Ἦ���h3*����Vh���@���2��JfꚼH�#acԑN+��-�@Y��Ww�P�I��}4�[��Y�dc;d�d�H:�Ю��K�(�pG��p`xQ��c�K��_��t�֎=[�?~��Cpn��?�M�H�a�..�{+ʫ��=�iB��-�N5z��}�7&C�Cd�/�I8�!�{Àr$n��E
������i�9P��E���!L����$����$��L��Ic~�7�߉����sF6�L�"}B�C��D����X~���cf����y�Ư$��ΐy���}T?P:A"��0�I?���N�淃h��q���+jg@Rɺ!2O��B�3 �j�c�wt�Qvi��5� &M�2�hz���DWɂ��Q��a�1ԉ��^��_W���Y�5n�R=�1��n��ω�B֙G���Y�⧞r��+"Q���I63���4g>��f�&�F,��{ۚal@�1��Ɣ3�Y��Gs�;g�D#e���N:{�@�Y�eH�ҰY�11d`��C{�����K��+�N�.��[h�3ƚ*���ݳ����K�"�<-9�1g��x��P�9s��x@�%������Q���p����ıe65`N>=����Y����}��\�*����N��}�NJ3�MS`�&�k�]���I�iЛ�	 ��$����J"�uۑj�,*Ũ���tK:j4u���F�����u�v:�YJGS�[F"]IO�'K�Ry���g��Nﳺ�E\L��}���O#�T�j���r�0�9)��G�oXE\��U��P|S���8��[*�-~)?]o+�Ϧh��x8㲮���1L����-_r�՛䜔|L�]Jo�x�W��.x�Z`v"�����B�{˂V�]���"���/�^.py�7��;����*o�O��K�P	����D�(�ep��7�g#<`�����eȚ֔/���2�D���rv3�+kh����l6��eN��V�N�پ�b|n]�Cd��I�:�
���a�Rg�9j���׊�p*����p=@�=Gn#���o��K�����8gEO�����7R�c�3�;��#�^౗���d8��2k	 i.?R�rP�s$WdF�yֲ�����L�e���E��`��&��0k?ySI:~|�^�)Q7!Y>}nC�'*��gM,�y-*��,hK��3�(+&S}��T
� n�H�1�X�r/7���`V��a�S���؋m�bE�d��-�n�P`T6}��]�@nQ+��ٳ��-���l���Ț�$Ԉ��_�����r�̫�k�x4�Q5����!W��3Y�q���
�Y�?�x�9�=��kO��>cp�y��n��u���H�\&h���M52E�T�&jƼ��n�HSB>a��,O�^���m��i	�n�O�y@J���	�=�
Ŷ�?×�S����I(Z)�����b"Ma���ŕmY�Z#�qg�tf�@|o�z��(2"���<�4����z�|⶝U�o"�6tsb�=�= \�nI%
�$|]8�!�3p�m������7�.I�+���h����#@$'d��$`R�����u 5�O0���}��#Q �xfu�[o4~�����>bPU0��*U,�}���!�k��0k$�:��J��-F�AM������V,X������!��Ɓ�; ���B�������a��Y��)�k�h|�бD��r����H|�$��v�zU��D>����el�$�|���wr
Ε΋�uw�݋n>�~k#���Ps�oCp����9b�Ë�|jr��T�ƜVee���T+��j����*l���W��T���A�e���*�+7	�Q6��?��T�����Wu��|7��b��L� m�?D�D�!��~F������ֈL��.��"*���B���Ŏ��o���^�0_��lj:������#˦��Z�����3��]�
 T61��]`󣋗x%]�E0(s�Nͺ|��p| �6%5B�5���Mj�ZG��;�p�������#�@�[��O�I(a��Z��׿���l��C5_0�l�*Kh��'��vx:���O87���>�B�y�#)CY���F�$|%��v3fow��~/��Q|�S�,$��[,��\��"�s���P� ��?��fh+	{�A[����[�{�lWm5���viDkh�H�����n^�Y�  �z=֣�I�5�����D��O��kjm��#º!�'���6�JswZ��u=� 8��g��Ua��Ϡ}�8�lz'��$�9/����0����v4��r��%�.d?ݻERK:co+��oĠhvҊ�[$B���o��"��r�q���ö=TH�Q�7�$��/�����Ko����S��(�boQ��&�*p�>|���/b��o��nSQ�w����m>�*F���I�<<���)����X�����w!s�|S4���^]�QZ/a�w���ߩ)�,���i�?��yϣ?�&Q����#}7���+O�,�M��1��f���M�i8*�}�S�=+� !��=}b�<�[	F��l8�<*]�)j�1�u)�{��1�sF�._����׆7�ǫ���J`�K�Ar��v���,GCL�������H�
��i٬1-p��I���Sz���ٺ��s�~���]>j�FE�&��=
��n}�ث#�TM_
L̾�|n��YFF�=+���X���w'�ՠQ�gAh�m��5K�C���Ḥ �Jmp��`K���.9ņ]W2�4	�������/�6+3m+	�2��=?~%�>���Go��:����_O������T�Z�u�_GdDmL�-�U��n1R!��n��GT�ke��<�	�8Ŭrή��ry�!�(f;� �c�r藛�1���S~���?��0�����q���̪�����р���M	�P��������<DF�-�dؚ�)���4�b��"C�b�՘,ᚶ���٨� �9�PqM0I�b�x�Ǘ�ut���᱊�>������-���і57@�����f�J��Լؑ�a�)�N���-�:1,�.w�T��]��vG[#^�����c���d�������y�(�ПG,�p�����csq�3����dt��t=�J�~5�p�"����� �aD�o�A�gEj=vi�A������w�./��_����/P'�ܱ72{S�$�r�E�/\g�Me�iL5��?���oA��P�E$��*ɇ�|��Qޕ�a~G������n#>6P��ò�Bq�p���W�P�[~�c�C��鯯V�"�g2UyE��ܪPʺ�p:���\��P��GE�]e�n�j�WT�J+U2ߺ��s��_*j;�nw�v���c�� ���2�4k�x#�D���5��-��Y�	τ#����P��Y��>����1��1n�5���h���OGYPYt��]+��ת]�=3N�4��������o�{�@O�)��p3o���X!3��r]D���&ۋNʜ@-�.eد��@�X1���"��{X�����ҥ�a߻�gޝ���;h-���F��{����K�I�̠�N!�)xo�i�V9N�x��w�cJ�U#���� ��o�Ne�N�N�M¯zd��j�%%R�!�\��p�7`�*iN��3'��`i&������1I^�w�@b� W�Ϭ��'uk!����ʨl�K�E�:�f��_��z�x2u��(:�k@G�F�
O6�"���|V�BgΏ��O�J��\ܯ"}J�O���T �v�����K')������\A��������dT�9�SK�)�,�n�#{� ��z����� �{:�-e���gZ�6�m�uƔn��������U����G� � ͨ5�ͺ�#�����j��+K	��K�x�ʡ��z�6=�Gҳ8!x6ja�0ϑ�G|'u}�)�[�=����ڇ�F�{	z\�H!�����R�h�}�i9��V��5s9�����F�$�Gֹ9;cP�h��U�kZ4�l�A�$� �0tI�O`LVx���70�k3���ѝ�},|��YEF�a��o�x;�<����
�E�i���Ҍ0D�	��EY�Q
�?��Vw+��Ɇ��ϼf���i7z���ރ40,K�M���$�-�q�C����bM����,U�������ԝ��`���S+���[>,��JoIӓ�s���$�k�c!�!���	�LW�˝�TΑX���%���#���l��3e��ʂ�*9�rƄ4���::�Woz�b����r��8��~����L��@`:�Փ���L����1�q��=���OV���K��}�ٰ`2K�a��3"�*�����92�&��e�!����O|dMak%�,�3?����0G;=h<��x��ܽ���q ?Rr�n2HdeV��n+;����U�$v�L�;V摦H�E�m\%�?�9����s�Z���[�I1^�����cq��Ĕp|�5�#��lôW&�S��Q�y�`�N}�8�R�Y�A��'�⡛�m�	��SG��֎����m>eYVG3\����ĒuaH ��z��T�V4���V��;I�h�܀��J���1QDCs��"(�����%��WO}Vn��&�9�$�r�B)g[�� >
�]��w�}!�BT�{O8��N�1�W팿�z��
��o���I��Q�d���ȠpW�0�\@����ZJ��1�*R��ڟd{��	�ڔ��^��8��/��1�#�v#��Y�ࡈ�:��^
x�9�q��@n�i.��!�(�Y�א}��]���]{��;�&���6=?���J�	>or:}�Sk�[��%���@Է��"�\u�.G�@�~r*>{�{`ۄR�#	56�h���d�:�*�Ė� �C P��~�8�&Z.����qo��^��2=K�&�􇕴�_���U��km�����s�P�t��m&R]R�d�87)W��J�!}v�s:�t����fc��<M������P�h���{��LODq4D��ٛ��vM,�9�Cj7�x��
'��<��K���;�?�l�w�����4�1�Uq��'�$�,]�y^J���jF����74=X�c=X�:&���]�i���},U�F��3�\oR]���B�v܀f[����sj�a�`����!4��A�ۋ4�`
#|-����]��V�"���'H�(��z��ٚ�B1�#<�ҵ�U]zn ��VԆՏLm�B�ϧ¸T,��������>���C��5��a ��iõ�*�#����Aȓ�.,3Nm��T6�W�]}i��T�
��;������(C�D��`����۪i�bŁ'	F0Pi-�u7�CM�������mI�T�K5��^�YPW&�uDN��.=�Aq�����L������_��������^�xԍN�|�K���[�+���%ګM�7�.�9��I�/����Ѱ+����y�1��-^���u�͠^������я��56���"f���e&ì�O0^��eC[�pϼ�s�̸ �3Y}��~��0W������!�1��D*�����Ѕ�JHf]����V��3����J��W}�V�&�_��N�x�Gw}�0$����l�q�6��_!]�dP^�N_�4��9gt���	l��i᪜�^-�ݤ�s�{��'���9�~>\�4����f��<���{v�L���M�o H D�.�� ��%��e4/$'��FU�.[V 3ME����00n�zk3[����,�����tx'�r[����H�M�z�xi�U�mcu+����e|b�f��z�2�֩~X�@ѡۅ�b2��ԗ�y���f�D7E��.�u!��X��0���3sz�m�.��{Hqb|:��.�Ugf@�n�_� ���Y)��
{1�� d#%�?����R�U��\�9������9/O�<�y����^#���PU���!�'܃y&��/�r�,�9G�����ד��F<���]?�m/D�H4�Da��P�%s�	�j��<�Xb�ϥ�Q�%��kY�b]s=�j$�k��eЮgA��vB�x�#��c�zVzԂ���F�P|�"y�W�sBR�����T�=����&���ս�ߺ7��s'��� ���id�:*�A��r�Aɾ�.M��Y\���VWW! i[�O�ˋ@;�+��s�C=�D�S���CX�+Y
C'�PJ4�vD�CnJ��9�u����T��-8�^��lP8h+uE̐�O{pA����5���9����➚��������-�xAݪ�ڰ��ļ�,[��8��!%�`�X���z&%I6��ew	�Q��n1�Z����L����u��^fZ����0��N8�l��"g�F�����>�^-U�C�W&p�y��4��s�Y0����k0�[����ʼ�h��Ңb�Z�����ѩ�Ji
l��+cIў�MW��%��J��W^{pV���_�S��C'�ن�w���$)�mó>�lg;��7J_B#�d��r�!���9�U��xh�l���!+��U���{��+�'X�9v�~@2��������@�%����C-������W�� )���/�FA<N�f!e�t�$����v�.Ȱe �@GEκ'��:��mz�I&[>���"_����U�=�s�n�&�H�LzD`f���*��I+F]��F,V�$Ǜ���Zm�4XvC�|�yb��xܙy���f�METc.��� ?�+��梸as[�^�/3�{i��|{	�.���@���_Yk����()��P{R�� ���͠ቌ �;UmT���>��f���:���zy�F��Þt�U����n'��&ȴ]/t��QA��GHp�cr?�H��<�"�]@�x/e��4��0�r���<	�����,�<�?Ẓ_�r�2��d���	Q��Nu6�z+Z<oA�}E�Az���9�{��ר�!��)���q쑨���shSK�5܅�4��b�s�����U���U ��k�`J#�R+o���m��(D���﹎��m�Y��o�XJk����z\)ǝ���̤U�2��咗��t�v�c`(GAXqg�628��W�[IO �6�P��7��M�_�f�q汜��K+C
�Z¸�-KܿLx�����f���.7�/>�X?܃��K�Y+�q3\aY	%ȫ
f��hX�.�}cb"�.�4IrOE��cœ�?z%����"��������;	���]z�&=e ?�^Esc��Q��`-	�|�GFK�Q���W��ل����o��S��%b�}?{�fj	KǙ����}rj���	��*�!ó�|��j�f%�K�#Kx�u��Z��&�a�ɳ&�,8 s�c���)�l��e��1v7���Q���Rx�V���:>�_��x�JR���_�]�^e�ZgL����HR���,�����t$fl���ga�]l�z��i��*A��=��t�i��'��m^3�eRu/�'Aa�R����yt���o�\5)���ճ.��`n-��Q(~I�%�s����ufm.\�,b����I6$"�(�ݖML�j�1��Ͻ��흃c�����?"�g�bǺ�z�yPM���P�����(�砣C�>~3�ջ�3���U���~A�G�i!�g`��0Rj玠���݁���n�y�M��6�ȷ��?��F��X�{X���҃͡������6E��+�H.�hg]���E�1�p�9��m�
�i�#�
.]�O��%:�sM���X�"[�=�%�f����]C""�d^/R!�.��7�EŸ�bv��2nO�,�������%D�#�e���7�M�<ngq��{d�(�i}-x�:�DU�x� y��y�D��R��y�"���Z.V!�㧕�b
��&��UI����A��k�V�G͝�|�-������FpKz=��"�ŽK�Y ������Qϊ����i�R��O3�Q�P8��l�ؗY�����~��w3 wĪRt�.�v d�\������Z���Y�M���%^����0�>|yZD�:�,+�,5�Q�7;>�Vh�����g���ya���u�KgN�ʶ��S�9Tc<�����@�7�`$2<���S�Pؙ�`�0U>d��~-S�.n��`"}օq~���r4Q"�8���#��C�-�*�����:�ViSr����ev�_�nZ�8��	k����5'42'0��"Y��:�9�碆�tN>��y ���Յ��n�|��p*��&v7��L2ӳE�tTҼ�?%nߴ�SЭ�6�ßl)��;}�i�����+�@X�����̣9�X���M|��!}�]~�Zwp���S�"�^b�E���'Z1�g�W2f+#�oӮ-�#��"�!��"�4Ϡ���|јߝ��op�ht�Nq�Ea ��Ie>�
�g}|+�U!��	��������7�a�I<Վ��n60�_�#���$5�����PEq��`���0���3/#�A���Zu��|4߄����>p�0�B�U����`O0!����1�k�Ζ���;�����o�פ��X"�݊�!��Z�����;����Y?��)���g��)�m"h
�屒a{r����R���Bv_EIU���>z����N��Q�(��A4�E��\�K������->v\#AH�P�v�oQ#����(9��G��c%���"�!��_�e��.�T1����p�ɣ.;Zck��	���(Ɩ^�{4�P��&�zfv�\��:M�� h:�5����$����Y{��>aH�\��Ro�J��+����i��o��ۇ莳Wo�`t0V]GJ2^�~�&\�8��!#⤜���������[I��*�D(��Mq��2�����'Iv/ 6�D�h����__H��qmQl���CQ����$K��L_&�ai'���mq/��X�Љ�3>�K�{�XRg���\�%Oyf �X�y�}�	�5�IY�������V�\%Bꉖ��"����&Y�!*T�D���F�e��@gc2�̘A-0}�NlJ2S�Q��`�������ir��6S�zj��,��}&��f1%��@(r�r����/�Ps�*̱������f��K�o�x����?,��m�`a���-�@8�L*æ����$�jΘ����N�FR����2��a�p�����R�D_�	�^��gSqn��D�?d�,���V8�tki�����gh��lx�Թ�A,�~R*A��J�8�t=�^�/.���Tg��,xa/�ژA�߆����%/�(��v�)bθ�ҳ՗#��\�I�i(�u�L� �b��l�m�/�,	l�i��6�4(=�Ms;��8�����HWc'�H�,�������$Ơ�-���Pq������G^��M3���z����������.�T!ea�`obϩ�֑jN��4G��ӊ�n��M�S�6�����h٩��1�Fh{�=7��Ŕ�Ϫ��a�6���H��g�同.]1]�@t�TY��0�ڔ�ĥ]�4��͐�����"bsk��O��[˷3�]�!�"�/��.%�74A��p꿾�O��M�%�қK��D�:�e%��7�R�<U��Xު��}|^��h{6D�_1�'�Uր�ѵ ��sF���qn#"hV��d��Z�b1���Y�韞ϓȃ�jӰ��Ϯ�Y�øo�%.o��i�p2�=������DA������.������Rk��3�v����K�Ӽ���}����� ^=�R;`p���td���W���{��V�T���딒�X�0�D�y���:�7S�s��Q츓>����kf�
g��Ry��о���K�J�ݧS��NT�`0�g�fU_�(7	�`kX���6S�:؀���F�dR�-�jan#�`i�����~�^Q	�nz�(%�-UA��������}��y���|�]�&/>q�̀�Pk |�I"c5N��.I���uY�p���V�.Y���m��T� E禓��n��nz�^Ϫv@��z&݃˳�%2����{�)��gen��=Swk� ����Ȃ�.i������@?�����J�m�ߝ�ִ�5�h��Z~����i"���	�+�B7�Z�|2g�5HfR��o�:4�
��"��m�ɘ4V��ӂ�i|�v�
�Xow&�thR���ŏ �T�I��
X�|ri�!��zų��� ֥@b7C��I�q4�/�}⚆W�#�n�$�1ֹؐ��L��J�0�0
XH�2�[#����mŴu~�4����Tzf>�!>0��-U���gN�!�ﻊ�kYD��F�¢wO�V�Ζ�׫
yX	���M�%��؜���;u���Wl7g��0�0�N�A)��@h��ձ�gr2Zg�~��g9vf�,U��3>A{�K��؉���!�����,'���ңG>=�g#�RPH�ko�za��f9UN�oD����朋h3e:�v�iS��߽�|�*�8��L%������em�*Zq7�b6K1?��*�w����LW���QV���L�ym�Ӹ?Z��D��ϑ����A��� #�|t�L1{%�]>��w0;���L��Ļ�^��^$t���j�ԭ��>���0���H򖸵a;��l i-��k7�����xxEš�ԮL͏��l�� C�%� #��DI�B��Z��;J�ͪ1�Ě�Uk��o�\���(VO�Z4����4�lv��6��&2����d���*�k|�<v�8B��Ā?B7�7�84bYR�F�H�%�<I��Fo��-�Sv�ƝYS�|S���8[�0-\�����z��� ��?]��h@��	0��[J����O��l�C5UH{vޯ�h�"����j���Y���ޣ긩5XM�aU��'�y�����W��O�B'K�����s���3x=\��i���a@࠲�U�A��ao�����߮�r����v�_���{鸊.�>ǻZ@u: ��ZI�ĕ�~vg{�[YE��[�W�3Ї؂qdF����H�($�_oԴ-ѝ�
����v��Gy����bm@��"�*���ɝub,��o�jn�3wQ��b_�*��C{o<
%۞ <��Z��HjwvN�|Hz�ɳ���Q/����&�)�VsLN��4����?��Q����[��#*	Т�G+���,U�ުm��	�2�H�o�8?���+=�s��O�}�rM<M�q0�|F�8�R:]?}ʆp�)�Uǒ�4�s{*���fn�כa2�|i��R�W`�X��O������áC�P�$G'���_U�^��1�ϵp�幌�nz(J����~{�]3��F�?��������Mg'�iw�
9��]\����F^=�+*F�X�1�w�?D�fY�A���޽��֍���U_mE���P2����;��2B��|X�I�T�k��m ��26 ?��>a��Gė��/�P�A
�_���l��Sh~T�!uq]G�[+L�/���R;أ�!Z?b �T��.��"�^�oš�خ����!��Nf�.�+�r�b����H�H�l���1��7[�hU���������v=�����\M�!��)��ʉ� �$�8-��C�	U����)b=E9C�Ij�m�ޚ+����pQ��d���!x0>��b�F��2t���V�)�S�;ݭW¯��8�۱I�F@�]~��> Jkn0��ia�m�NIl-�?k�U�w�j܉�:�΂�4[8Ęک'c ;�d��[����(v��G��cp���Scq7�蠂ߵ��t�t�=�1~��p#���}sI�a9L=ʠ�����d=KU!�[D���z����������h��/�ѹ܆(�{�u$��EZ���B#�iᱜ�t¨�D7���|�$����<|��1*��D|~���N�C�C�6�C�����B&��);�E��~?c+���D���W�|{)y�Ga�b��P��e����%#I��u�r�]�оjL�r�?}@2tK&����i&j���wV1v������ �]�2$����+�D��S㪓B�B/k�vt�ez3�$�ф���R�Yb�u�R7��M1A�������I��g�}GG+:YI��w�+�&e��3�|P4�mh拢��Q����^f��@d�n���R3��ָM,��`�9D�<���(N?Q@Bٟe�^�ҕV�1��嚷�{{���V�����(z�R5��'�h	�{�O:�E���a0�K�5��V��`�~��^TW9�x�~��*�ʏ��3 c��c��� �e��#Nc�w���y�����6ē60o����$���No%
3\0G`>b�p~ը�r[I'қ��B L���+ ���u@b��1Ө�d_͹QD:O����m�kG�㭑u�>�:�kSG��Fg�O�����U�7!gN�@w��%�\�j}�޲O6:TTy��i��t)�9��t�s\+��|M�56��Yџ��"p��|)��Cn,����z;V��C�����E��[���q��Z$�ޅ��J�����ӎUgq/�r������K�15�5V82�xi?�l�j�1�K>��� ?X�?�X���.��Tz���8�j�"���_|��!�q��p��k����;�s	Q�HVGr�ZX�R���ĒI�i�؉V�5h�d�G�Й~��J}�.ce��wT�k�	�l�����Mq�0I�Oվ�x��D��k���v�pa|�FEG��f�xP��b�'
%�i����!9��>��E.y�
�����q�|�ī"�q��7�f��b���,`n�MH��k�A$�Ayqr�g�&���7����,j�Ѳ�hUD���D��ٵ�uy����>��?�$-�f��N!�����tu�R�ރ��k[���.�;sG��t��&@�H��8��W��8�8*!+us��C��ǲ�T�фSd�M���ҀV�?�)j0��qba���V�I�5M����d%�/�'N��������#!?B�=��GË	�4v`�U�/'#�T,��yL@m�A���� o4zz��ƨ@˥'*��W���+�?ù^F&O.�JZ�Rx�۰��ܮ�`����s���Z#�<��j�������`8��-�ʯ����z��=0K�����jz������BB#��A�G��zA�؇�˾���ox�D�B�¦��{wT{-�K_F�o轛���,�������OX� �6�i13*A�`�5�AvB
.��F��B�+W���i(���8]s;�*��WT�C��D���v8�X�0�^'7�PWڡ�#��C�=��&R�[��T4=�	=^ ��PE��u�f��k�A��1��M>��be9H��G��J��{E� �x�6�jO=Ù߼���[��-��%�`����s�gZ�I��ڈ�Z���˒ۓNg�L�J�Ֆ��QuԳ^�TP�LEc��e���ܣy 3"��ӌ��+�u^��QC	�yp��~��"̸�&Yț�싁0�f���]޼����b��rG���T�~r�J��@�����v$�z�����\JF��Wk8V<�_/��0lRfi�w+�0$�~� 2;lt�w��s_��d~���@���)%9|����x�l�5����Yu��g��i�9'��r9C��~�_��{ފ@�#��r���mݽ�)�qغu�{_� 6u��x��S�e"K<$Ճ;�$�.5� ���E{���?e��{zY]�[ke����$�b骾 �}�sTH�?DzѰ��(��Nq+���S����������<�P�X�D �I��b`E�ԅh�yC�`f�AEA;�.��͏-[���7���esh<��ܝ{�e|h�.���s@X�_�cP��3)a��{�\> �M�-&�M��U:�:�gT��sX�����9g�y�"��L����'�U]�c�'�Hu&u6�/U+�����(GL�9�0;���<�_$]�/�E�4�X;���l��Jv	���J��<�9��gεο�5��c�P���E3	�N�
ۇ�(Z���O+��.�?�$�i{��e.\ǀ�W���'�U�,� �h@`�5��F�58��/e+�	h��b���I킢�\�X�gJ��/+��4�:��$C���m�9f���Sb\%�J�G���&\�J��'~`�biFř���Ŝa�u����(t��q4��2�N�d <I���6��n��k�Q_�ޘq�/�$��Cu�e��KYx�Le���'d��*F��1�/�B�XL�D����K��^�C��$�\���%�#"f�nX��x}��{k�I_�в�����N]%��2�/��G+�m
�gm#�Jw�����-+g�+�c
q����-�'#����8�Q�r����]�Q��     i  �  �  [*  �5  A  WL  X  c  �n  �y  =�  M�  ߖ  0�  y�  ĩ  �  J�  ��  ��  B�  ��  �  w�  ��  G�  ��  ��  8�  � �	 J � t  �' ?. 
7 �> �F �L 7S 2V  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�=A!L&�S�ӰS�����<l༛L��5_�C�I
/y$Ցr�C	ʔ3d�O��"<yϓ|���q"��L��aрFF�1����`�^h�Q��hPN�}�d�ȓ!��x!D�<Tt
iz��ޭL�e��~��TbԀ�.͒��G+/���ȓr�]2)��ԭ��
�Vلȓz�<���!�P��fͬ3���(�����w���t,\�H���K�D��`���58�Y"���)A��=�����v}��B"���sΝ���l�{��ı;X�C���zC:T��'�J�x5��+s(T���	ف����ȓE��G���V󨤢�.�=x�i�ȓ�P��dC)'�l1�c��
Ѱ����`��C�
iv�@1
N ��Xpz��)k�<Bd
�>r���ȓ��
�h��l�R�ѻ�����)�J�0���Rn
顂�T/��A��L���S�)	�T\J�c��>�r��ȓ|6`IV�5^���Y4��E�P�ȓ�b�෠�3%�`��/@�J���NQ
\K�HJ'�]	��Fp/��� ���b�BA�;�:��L��K��@��}vMc��O'�=���4��9�ȓX,,����W�Δ[���L�&���T���'-JH
��ZT��,Z
�'	�p3Bl�v�`CRCς\Z�'��$B���q�(����"M����'���Z�Cq��%��K	=d���'�~�:�K
�gM+t"ݚ8�4����� �����H	��hT	�&`M�jY��HO?���<���K��ˉ�a�ʇ�<�!�.
��9����"�!�D��?�!�$ݨR)Ҙ��F�3\}� �)�i�!�d�%�����d�	�� ���/!�,��e�J���H�G��Y!�D��� 	҇��Q��U�Ɓ��B�!�
Xۄ0��݁�L5b��ՙ%�!��!��)�wI��'��L	"'_�z!�X�`�┥�6>��pQ#DG�!��͉să��w�e��ˤJ�!���6L\I*��n�����'JB!�ۂ�|�b�RS9��JC�s8Q��D�t���I��D�&�S EN	��n��ybh6S���HO#<����gR��~"�)ڧ
�~m��%��>��%�\\m��!�L��Yq����6ō��R��ȓ2�|�0s��+vS򹫑!<6J��ȓx�<y��'C9Y�D�3`Ν0{$�ȓs��MXIE=)�����*oHd��]�hX�Se�;�̵qEg��l��C�����8��1�e�^�F�dQ�ȓIȐ���C�k� 1ӱ�2(����u����呼	vzQ�jTl���ȓ>ܒ���!}[� �0�V�fxh4�ȓiw�0����)��0�%*D�|��ȓ*������J����\k<��ȓ1JX��i�,*����C�Ϩ���<2��(��6Q�6|�Gl,^�hx�ȓ�z�yqC�i�Eˡ��+���ȓ"�qy&��k������Q����[g(�(c�\�j�a��_6�M��A�Z���/t"@�A� 
�%�ȓN=�)�����jF.��+<@�ȓmTY�D)@)X�HARd��e��X�ȓ��u��%J�=��eb�K�N��Ćȓ������Ƅm�`�V� �Ƹ����i���Bvu`"Ԧ͖��X���ޱ0��:)VE�RR,HЅȓN��ra���R��hg�-n`(��F�D F�'`�,����G$�]��|�J�:���(��	>� �� ��"���*k56�MC��G{r�'��A��� W��9��J|HYY
�'F�z�*�*`Q9�%ARC6������x�,8/�V���L� W���c#%Ư�p=a5 9扡{�*`l�q��Ff�4��B�I�q�|���	,}�x�NU�b�E{J|juG�7`��H�G_�N(p�VL�<)Clə	d��)H�hlT�#��^�<���9)�����j4R��;֬v�<�ǒ���@R	��5�(�Cd�L�<�G���;��@��"ƪx�Z ��AF�<�0�X�%jFL��r��	p��B�<9�˙9[�$8dOH'��X!����<���)4���� �;j�ny�g�x�<���\0(}�1K�-�<�*�LWq�'@axb�H��H�2$�k��\�j�<�y"�.m��A6. ]�P�s"���y�N�61��#c�V�AB��y�Ά5xr�A��W�Trt����y����0h�J��R�P�^�21�ʂ�y��ۨ1*��I�I����ע�y�n��P9,]P��4Bfh��ɣ�y���� ؍��C�W�rAWF,|��Q
��'ԉ'W���\;����R��7x�Z�Q�'V����y�e�"�J=��
�{2��L����$��f����`�ѰZ���"O|�P���9Ct���
'� D����O�㟐&�L�,�GG��#�kA/(Ѭ�*7g)4���`��.f�Q�&)V/\=��h]n%!�$P~�i��M3LWF��4�Y0w-�y��I 
��A���`)�ep�!P�mښC�ɛ9(R(ɰ��S!~��M
�dC�ɏ"��Y�h��:�(兌!K��C�	�}!H�K�G���&���L�L�*B�0g2H5����h�6h{$B�&c�B�	�:X����3V��=�a̳.�DB䉜_��V�pU^@�vE�1�.B��(8�U �"��21\���N��r���d*�Ĺ�
�-�������SVν	bi:\Odc�@���*�`��7O�v��"�%D�����
囗b�4�M��N�40Q��>��ŌÊ)j�G�4.:%o%D���D�R����+�e��6���)s�!D���N�1:����}]��D�%D�p�ǡ��Ez�����]�1D�H�Ç���L���'o�����k"D���CĘN�p�kD�%~�Ci?D�t -��H�t��"��]U��aE�)D�|�Ѓ�.�qIW��TeU�2D��Ņ_���1�M�-�)�Af/D���4eտ;���r�g�Si(�K4�:D��s��/a��I��zl��m9D���榇�2͒�
1�P�C��<D�l��d�f h�hN�FI,m�Q*O:,P3�>0���(��'��x"O�倎+@ܨ�pE�9Hz�c"OD��,ܲ?�:� �$Q�o�1`!"O �����*mL��m�=M#w"O�����ӽCE�����/$쭙�"O�+�DN)ܦ����1Չ�"O`H��/ZF�� hb��2��u�3"O8�A�7q !fe�
pt�0IQ"O�����+A��:	�Y��"O���� L�Q����cT6�i"O��'�Y2!����߼GN��{�"O�H9�74�X
3kT�#N�Q"O.��ckN-E�|��WI�'?��9"O2��K��z��!)R�v�|@�"O��A�lM�/��������B�X�
 "O"Ԉ��?EE�`��.;� �8�"O�}�J,Զ�avj�#w�� �"O>�[WLPj���A)��v��� "O�1� ��b|f9�?�JM#%"OZQA�C�'8x�p"��a��`:"O h��P+x�lJ��,*���a4"O\���],|�>�I��Y=f��0�"O�G �(rޙ#��Ʋk�	�Q"O �RvfB�v�,�zF�:)�^�+!"Oĝ�@��pH|�P6�[h�*�"O@�G,�(v{&A�����^ѸG"O�8�r.V�p�
w'���r�"O8r��V�NeaElU$u�ڢ"O��ƑR]*=��k�*W�0}A�"O��p���DE��+�/d�|"OZtk3�S	�D�KS/i�u��"O��!�%z�^�9K�3s�*u0�"O� �- R����W�D�<оy��"O���ǙR.±r�
��L!�"O�E�a��4+�ֱ�B� >6	2��1"O��f *~��;d�Ԓ@�j�ȗ"O���f!�`�J�*�^�>��xs��'|�'�2�'��'E��'#�'�I+�A^$ܴ��P��E[6�{��'�B�'���'+�'_2�'Qb�'�{`�˾RO��A���'|�x JT�'���'~��'���'<��'���'�R'�X*J��l1� 84���'���'�R�'���'F2�'�'�P�._�Bi4q���H@�h��'FB�'�R�'j�'r�'}��'W��s&�y��E#uÏ�#���(&�'M��',��'Z��'���'��'oh�Ȕ�F�O�͛r��|��l���'m"�'o��'��'L�'���'���8�͙\E
%���D�4�v��@�'���']2�']��'=�'���'���p�� -��)���1`�'O2�'���'s��'��'��'�V8Ir�ߘH�2%B%*Y�`��=�G�'��'���'�R�'���'�2�'�b�fҲC�`�ZU%����q9�'B�'�2�'v��'��'���'��3C��xz�A3���k�e��',r�'x��'��'lR�'a"�'"8@�"$N�I�mY�	��N��g�'=��'�B�'A��'lr"`Ӣ���O��ac"�>1T����
y��*Q�Xy�'
�)�3?y�i�8p�aa��0f�'`�~4́���$�ڦ��?��<��4>عR�Q�gjH��'
�(*�K��?i��ʡ�Mk�O��S��
H?	P��ǡ`ʄ�����%�>Q���4�T�'��>���f�-$��(�6n�U�Τ�Іܹ�M;���Z���OV6=��|K爎�A<N-��K��6���L�Oh�Dv�`ק�O[�ysr�i"�� <�0ň��'f�z�����'6��r�tj�{+̢=�'�?���$C�`X��8�� �G�<9,O��O�qoږqwRc�xX6B�"�&��ݹ{�6�a��G��="�������<�ON���b+�N��Z��s������U^̡�3)�+U_"�韬��$Q�}�<쑦a��?�$YŌ�Zy�W� �)��<�j
:zⰅ���£G�6mY�$V�<��i+�9q�O��n�n��|�RN�%1�
�'Kغhi��AC�<��?!�na@���4��y>m����(���CB���E��*i�0�2�$�<�'�?����?���?��l�Z������ܰoon����O!��Ď����0/�]y��'2�����̇�ln$���.��ݹ��I_}"Iu�<�m�9��Ş��,�.\0A�u����,��,G�n�	2�u]҉�pMУ�j4�^w��O��'� �ppj�=�شΆ L[hĻ��'���'�����X�"�4|�@Y��_oB�O�b`}2�9'g�d̓�&�Q}b$j����'+`��ރ ��8���]\^X��߿X���>O�pC�˫4B�J��\?J���]�2��`Z��܏�":	Y��I�D����`�	����Y��5����$��4�A���p��{+O�������%|>}�I��M�K>QSOA gNT��D7T(���k�4�'�$6�R��v��$n�L~⦞�@�>�CPh�0~����e+��=B�����w�|�_���?G�Y�1����)ҳy�&<���	L�'06mN>s�����O���|�n�:}0��"��9���hT�U`~B��>i@�iz�7_L�)b��.�ڸ�C�dB,�7�%4�p��@#H1^<,O��H��?Q�9���u0��1A׺����� b���D�O(���O���<���i�v��NZ�b8xR%��"{�M�D������'��6�/�4�>�'��/T��Ф��&9��d�	�9r�'����i1�i������?M�]�T���������w~}s�}�Ȕ'Ur�'>��'���'����X���Ҁ��@c��5Y���j�4�zX�(O��$��.���OB�d��6��*��L�_ ��ꔖH9�pi��M;Ǜ|�'�r�'p{���4�y�$ŗhh�qcq�A}��P���-�y�:x0�IE��Iڟ��'���'A��c���%��iR�?~��'���'��U�kܴB4@,O����;���h�69�lm�&�>ƪ�Oz���y}��'S�|b��AKP}�R
Ի���0��Y����Z'��K���ɼ����s���.�DX)sxq���6:�Ի�G��3�!�DD�J2�!�B���,�w�U�uv^��ަ�	!�Qڟ��I'�Mی�wT��`�'㨘x�) �0P�8�'��6mDզqشHafߴ�� <a��9��[D̓�@NԴ#"d�,5a�i�'d-�ĥ<Q��?��?)��?�m�=��*���P$L��Nġ��dU���0Ilyr�'��O�R&��Hd��'D�%���x�aAR�l��?���S�'%DJ<{Pቓ%e�1	gAύ]�-pToM'i��(Orq�� �=�?yJ)�D�<Iw��A���n�cg.t�6i���?Q��?���?�'��Wզa�hP��L�bş�b�:t��O'E|��×A֟L��4���|Q\�p@ܴ>�����q�V��P�ɲ@�2[����_ ��qog~RD^�~���S�9&�O� �p@
J��y���4t!�!8OB��O����O\���O��?E���'#�ȕ($mǕ)>ӗMUy��'�6-C3&i��O*inZF�	�:�����e�]a�d(1 wX�h&���	͟�S0�nZm~Zw��P�#W�+6��#�.[�$���A�:7£�m�	Pyr�'�2�'[2'~69h�(�+ )��@�rZ"�'���M6$F?�?)��?9*���!�
E<.
�sc���Ұ������O��d/�)�K?]I@��udL1N����I!��+!.^pG̨�.O�8�?��3�D�S����+_�z������@6 ��D�O����O^��<�&�i��{3j
�'����d�¨
��Y{#@�+7���'r66�I3��D�O��S�-!b>Yc#�6	�p�4�<1j���ic����EGL%ji��&�Oy���K�R�Iԧ�������y^����ݟ(�I��p���(�O� �E
��2���h�3y��Y��m�r�3O���O���d����)f�t����/9��4c@l��5�f��	���&��ן�I�6�l�<�7G�Qz�V#"���6K��<�g/x4.�Iw�I}yʟ�A�ц�=T�(��+lp���'��6T�[o����O��բ,�����ȴ-9h�*FGI���RϨ>���?�M>� AD�@��`$��c�AJ~�*�>T��(R�Vc��OE����c��/Li�j��B�I-�I)�E�4g���'�r�'q��S��|&o�&������l��yā����۴F�PC��?��i<�O�N�5I��)) ���i���>:d�d�O��$�O�=	�l���ӺC����´@�@l��##̓�'�ŢALD9d�O��?���?I��?)� /�r��({�ܸ�1i�iv���(Op�oU4X��ğ��}�ğJ3�*��5a���0��%^����O�$/��I�`��b��"4`��j�$>憱
��A/cN�˓@�L�����O�9�M>�.O���AAW�D�x���%�"!8�m�O����O����O�i�<�a�i�b�ʖ�'H��iWA9N�8E*a�`��cKr�u�D�`��OL���O����%V�H "F�M��5�>`�h�S��b���ޟ���	ԊM��D�nyB�O:��C�GYb$���O*2�P�4"�#�y��'��'��'v��)z���`2��W�X�s���C�����O������� �Rvy2�a�P���<Q��O�B #��N `0���V����?I���?�҈ȫ�M��'5��.kK�шUʔ����pf���QZ�9���OX�K>.O��d�O����OY�IЀd_NP���E1E�d�c�O^�d�<���i��´�'g�'U��*b�5�eX�P)x�e숯!�J�}���ߟ���S�i>M�	�h�,t娂�W����gT�����¼=���{5�@oy��O��4�I"��'U�2���qaA⴪ʧ}� 0��'���'�"���O����M��&@�-�XŪ㒇@�0�{t�>cݠ����?���i��O�'f"�ِ2ԞD�R��_��8'G��	���'�����i�D�O�=9�����qN�<�Œ�Xiʄ���D�6�U+&G�<�-O�$�O����O����O�ʧ`9��9�uy˵M�
,-pE�vmۣ�M[�-$�?A��?QN~�Ǜ�w� �� 폠:t�l �&�GR�ؖ�'2�O���O���D�.��6�f����N9k9
q[S�Z1N����Ix������4"�b�uy��'Z���& ^(���KD>@�!�S�U2�'��'(�I��M�Ca�%�?q��?1V D�d��pʴ�"#���@4��>��'7�ꓤ?ɈB�C(W9�� O��!����)����$�R'��;wIX�g�ؒ����e�J�D��_�)�3��15��HV� ���O���O�$5�'�?��'��S�� ��	��X#AH^��?��ihB�2��'%�`l����ݲ1MD`:��[z2��E��i��	ޟt�'���HW�i����^�8�V�OHD�j�`�3Chʉ���P�L��z��Vy���X�Laq`�M�(]z���0�,�c�v@�r:f��O��?Y����d���kJ4m�0ت4�R:���CΦ���4Z����O�fa����q?� ��g��j�i`aύ�xapW�����<>��O�	ByҨ��Q��x+e/��,җ���0>at�i�Zd���'J��B�\ x��Hk��k��:��'��7�4����$�榽Yܴ%ϛ�j��-H#��.ܤj&������Q�i����7Pv̂�OR�%?��� V�d���M?,	�.��`3O����Od�$�O�d�O��?Iȱ���[)(� �?vtrC�ş���ϟ��شL�8ļ�?i��ir�'9��� Z�1�na��>;t�᷃)�G֦m���|�r�˃�M��Oz4i2��NR^��C�*���"��*W@��8��O��?1��?���r�M�D-̅� ����$�u����?)OPo�n���'m2T>���U�͆x����&TO4�q�%?	%R����4)Z�6'�?ɩ�]�I�EI��p7�H"�蘝z):�I�#�\�JȖ��TG�̟P*��|�o�BKqCQ�=\�dX�3^�"�'�B�'&���P�Ȋ�4&B�KT@��z�ܤJQ�K�5�5KA���d��y�	m�	������8jWl{W*J�O[�I>�������ٴm0��4�y��'mr�����?HrU�� �@rk\�b
D�r7A�i���=O�˓�?����?a��?A����0Jtt�F��<'TIA`疟.DIm�f���	���	y�s� ���c���/N:!�4��!��i��	�?1����Ş� <Hܴ�y�P
�w�H.0���!�b���yR� 4qp�������4���dH �̩
��� v#��9a� ����O��$�O��A�����<��?ac� ~Bvđ�y����$k�O$!�'\"�'��'H�j���vVՒ���	��O ��&/�8~?�7M?�S�q���O�K4O
�n�A����(�Zp"O޹�a����.ś2�ډc��huB�O|�m�.x�I����@��4���yW(ڲ4�@ �-+��t�U�y2@dӸ	o���M�c
��M3�O��k$(�+�r�揃t���3��,NZd&�עs�l�OPʓ�?���?����?!�I�tUض�3=F��b��	zm��*-Oh�m��L��I�X��]�s�,� JU4}�a*Q�M�5m8����OR��!����<�&��3�K��l� �L�@���>L,ʓ3MJ�5b�O�0�J>�-O�����D�s��re	%/dN�Pw��O���O����O�)�<Qa�io �e�'h���gH�g�3(���iR�'6� �4�dq�'v�7���1pشr�p�r���>��D���%U=�(�@�E2�M��O\���d_��ڲ�(�)���d�&�Y	�<��la��>O����O��d�OL���O��?5( `A�)��Y��MܑJY�<�	8?����vl���$M�%$���Df\/LqX� ��[�@U�2@h�����i>��1,�����'�"	7��d�
)�t@ӓp+z�	NT*B^Y�����4�6�D�O`��5������O�̱��I����$�O>˓ۛ��ȗB�����0�O���S�[�B��!���!B��p��'.�>1���?aI>�OM��yFE��S�*�p �U9j�2t���
�g�E95���p��i>�"d�'<��&��ڲ,��%%�9�!$���J"l�� �	֟��	��b>�'��6�Ϙ-�*��$ɞ,D�a�ؤjhq�(�O���٦1�?y�W��I�e�m�"a���P�%����I����'� ɦy�u�d�����%by2l�c�z���O�u��X��H^��yBX��I�����@�I�ЖO������,PHǍ<FaC#�k��9*��<�����?�Ż�yW�A�'���S���!#f� !�/UR�4��$�O^� 4�a�b��xƖ��7'ÌW�hl�T�L>"�D�I?}E2�h�'P��&��'�r4�p��\�k��݃6��1HVihp�'�2�'�W���޴n^Eϓ�?q���t��!�Af@O� $
h���k�>���?YJ>y�K�^�9�dd����� ��<�dFJq��Ϟ�M��O��)?�~��'�(D��\��}�ׇߔ��� �'4��'(��'��>�]�M�h�+���µ��B�%tJ���I-�M x~�p�d��]��\1h �?*z�Qc�	hr�	۟���ʟ�Pv�����?i������?mxj��t`B�.�r��ҁ�:KlD�'�������'���'���'b`���$X�J�:
vb j7�h6U��zٴw�jT����?����<�R��*u��T��G��2�����)s��	ǟ��Ie�)擡kn�9 ��#��k�"��cf�y�����8�'���p������s�|�V�8Y�l.9L�q��"�$��U�T�ן��	� �I��jy�`ӂ���G�OT��� ��`d�<h׶�S�&�O��m�C�i>��O �d�OP��Ӎ[�T=��!Pbȉ�G�/_ށ��oӾ�I
|QT��0��J~���UPT
 EQ5^� ���0 ��L���?91�ǌ'���weO3
���4�ܗ�?a���?�r�i\�͟� m�V�	!6Rd��T�P�"\Ȑ���w�v�I<���i��7=�*�,}���@<����]+T�b4�o�n{F 2N,����F3�䓮�$�O��$�O��G!��� ���;ĝ�p/�BN ���O�ʓc�F��PR��'��X>�[5�˝`h����K^���z3l=?�`P����ڟ�%���Z h"�**P�p0o�;ľq��� K2�ѧB�4��4� e��T��ObLtЀ9���xPm��2��(����O���O��$�O��
?FK�<��iO||#�
�]/��YVi�U���v���B��I2�M�J>a�O���ݟ���7��������U�8A1h���I:USlDn�<a��oT	�թ񟠜1(O������I���s�0��W;O�˓�?9��?)���?�����V�cv�s��v�B��fk
�F��m�F�RI�	�`���?A���ş��ɞ�Mϻ4��r�a��P&��r�
&<^(�H�����T�'��o(��=O `'��x{,�@ʟ�p5��h3O��8�'��?!W�4���<!��?Q'I_�����VH� �Rg���?A���?�����Ĝ˦C�������C�#܏;��9�V�̹2ǲ��Èx��ea���8�Iy�#=�dR��5 Ą��JՔg��j�������~�<ВN~� �O(���p0-5c���X��%i!�i����?���?I���h�V��D�dV���+�5uv�2�%p�K��'��6��"t�	&�M���w����gGa4	��(�gn}қ'�r�'�rlށߛv1O���P/1����π ̙*�dún\(������B�<�d�<ͧ�?����?9��?	�_@_�Q%� �ݓb�U����5e͞՟��I㟼&?��S�N�[U)Y"�)*Ş��5B-�>�`�i��7l�)��G#8�p C�w�y����2����A�5z�'�����i�ş��1�|�Y��;`��S���S�*L�S�`� �o��l���(������IyB��O&����' �\����
U3[�M��D�'47�8�ɢ��d�O:�k�(<@d��3���dH�7P{�Ea ��M�'��nO�(ܜE��g@��?U����$)�F 2|��!�d��[ˠ�	ҟp�I���֟p�Ia��}C6�kbǉ51*e�3�ƪ5+.�/O��F���3��h>��,�M�I>���P�~���ʀC+2꒸��
z��'D�7��ަ�S�*=o�P~"ѓ����K	u�a����d�
1������0��|�[�������������5CI��(`Ȓ)nta ̟ϟ���By��gӼ�<O�d�O��'KMX�����	U�82�N�+Y�R8�'���?������|
�`�<�u��r�G�+]��;�c�LlA�4������'��'�9�pD�0>Tz�Z���d����'{��'hR���OS�ɓ�M#���1�%+�G��1|^�KZ',x��'��6�,�����O`�C'�lh���� ?�U����O���W�W�66�e��I8�д{��~�*���H'eŠm� 9CQ+Q������$�Oj��O����Oz���|�Q���u0$9Q�	�F��<x���9ߴN=q.O���&���Oмoz�A�ŌX��`�j�c_��4���H��V�)�S�ve��o�<�v�$4�e��;c��4ۓ�<�1 I�W����J3����d�O����$v���u�ƌt��2L�o����O���O��[��HT��y��'MY'Vt��v��p)	5���|��Ox��'�r�'��'�ŀ���/kl����'�m�����O��!t��/a�x7�>�S_����O$�`"h��|��{�h��C':y �O���O<���O�}��DW�t�Hf�a��!�Ca8��%ӛFj˶,�R�'7�6�)�i�E�E��KQ��1���<6%��h����wy��A)6o�����c#�Ѱ[��̌#J�E�#��Kׂ�zt��<\+'���'�2�'�R�'�B�'��`�B-�$���d�L�p���Z��R�4u����,O���?�)�O���f�ɚ-�@&/ �P���+c��n}B�'��O�)�O��e<~}�"�ϗ=y����'ؠ��Eؗ.Mjʓk�`�"��O�4�K>�*O�t8��J�'��qx�c�9T�����O��d�O���O�)�<�P�i ��C��'fr|8W�	�Q������
R��Zp�'�6m?������O���de��B8~�=�S�S#qi�!��	�M{�Oƥa��ų���6����~�k��3�E�d�N��s�0O���O����O�D�O��?͂���5C
�%�r�P�>�P��H�my"�'��6�G4l��O�m��I"&�8b��B�Q���/�6�c��	Qybg#"ԛf��0 ��$!dL�	��K��������~l�'���%�d�'nb�'�r�'�X�	C��=�r%	�G3QH���'��[�h�ش8�H�q��?�����iC�t�F�('��4��y�i�=n%�	���d�O6���ʟ���\��슆d��DRސ��,�=@���`�O�hM�y�'���Eџ �v�|�o�dB���0b�	�c<�b�'���'���Y�ȊشrR�$�U�÷|�& #�ᓦ5*�5��b~"�`���4٨O��D6 *�ɰ�Er�2a�I��o����O���Oc���Ni�lr C<Cf���a�]��r�D+��V���|yb�'U�'�"�'U�Q>1tNշ��p�-T6[��:,�0�M�$��?���?A����9O�lzމ4��
R��j���6g���!ʜ��,�?ͧ�?i��S��۴�y�o�.+!��KF��!Z��{��ѣ�yB��d�H�I�'�'��	ş���e�]X�%H�DG"�!uf%\���	��D��ܟ`�'Jr6- 	6���?�u�4WFT%��l�=e"��Ȧ����?ISZ��#ڴ̛6l$��0&����� ����9�+�:\Q�	1#���W�6u�|�$?���'�|��	>���w'�+{�!S�QV���IƟ��	����	S�x���'+НÓhՉ���0����@�T���'�27���2'���O��o�q��李���Ӵ�T�\�n��'I�K��	ޟ4�I�,��(�IΓ�?yu���6����U�J&\��K#���XԂɟ2%�(�N>I,O���OZ���O��D�Od���ڞdUfM��"[;��d��Ƞ<��i��y��'��'��OK��.�� �O��Z��Pr�"Z�>j��?���O�r�'f��2��# ��Y��5 �4� -��AT<(ze\�@�ǂ����c�	vy�&B�[NXmٲ�؎{���7��ct�'�2�'u�OU�I��M˥e�1�?	�ć�-���7��&i����2�?y_����?��Z���	Fy�F#Rf�P�!Բ@�|��� �'d��TK��i�����A�O.�M%?���LN�+$o�
`ɘ1_%~X�����	����ܟ���B��	�x��G����ZM�lKΌf~B�'�6-X���$�M�H>��ʝ ]��NbQ:�������?a��?�d"��M�'�%F��� D �a��Xo24Se$G�r�@��~��|P��S����IƟ(�5M_>S��x���j� ��w �ڟ$��Gyr�xӼ�X�?O<�d�O�ʧ|�ޔC�26�����=�F��'�4��?�����S���Z$Ms����@ڝVs���'R�
���Dk�5u��&����$-��D.���Uq���S(C�^�p,A�k ����O�$�OP��<��i���
 �ӥO�H�2͚2c=3��:���L��?�f]�8��&	��в�C	/�ll#@+ɛH h������`Ԧ��'�,aQ��`ܧ>+�z����zP����Jg�e̓��d�O ���O>���O����|"�j@�)���;A����\(`�F���m�&�y�'���'�26=��P��څ^Hn�)U��-̀R���Oh��'��i��o�7�v��:�#Ҿfi�5��.e�0!)D-k����f/X��$)�$�<�Oڲm1�VC.5`��E�D�Q
Ó��&�fT��'���%P����M�Y��x"4���\�OX��'��'��'���IA�I�x�(��(G�����O�Qx�	�jk@S=�)��?!�Oz	����L��l�iA�i�h�rR"O��R�G(���.vHe�F/�O��m3�q���L[ߴ���y�M�/C�Qa�r|f�b@��y�'��'-�1饱ii�i��c FI�?�2�B��&���b)�9<�ʁB�j�ma�'��	X�'޸!����.^�ĂS�Ǫg_bl��O �mZ5H��m�I����V�'J�f9x!�G�J�8B���X?�Za_�T0�4��6�'��ɗYz�$ �n��u�T<�dF���͙�U�b��c�nd�G�O��I>�,Oz��*T�tIЄ+�@��2S*�O���O<��O�<���i\.M!��'��ի&�W���pґb<�vp�1�'�@7�3�ɓ��$�O"�$�Od a Ɓ45{6�aa�)z@��D�H?<7�r�,��yٚ�P��O`�L�'t�t�w�:LQ���-AKx�`@���#�Լ��'I2�'���'��'�2��ƏM�n� ����؂p{7��O����O&alZr�d�S۟���4��N�в���C�R���M�w�Dp�L>����?��?{���ش�y�ԟD�O�#@�P) �]���FT?9����䓻��OP���O���ˑ�0=I������J��=y����O��uśf��P���'C�Z>������_��A�b�J�@�̝��O<?y#T����`$��\����r�C���R�ٸD��|���+i\y��/��4��H��%h��O��RD%�46�t(�^,/>t����O��D�O,���O1���	���ˁw�J��&���)���0aF�[��p�[�48۴��'��ʓ�M��G<h�J��T'g�z�NZ�q��&�r���f�n�"�k���ad�p�K.O��d��?2�@�1Gē)sEz�#0O^ʓ�?Q���?����?A���I�:r�^L�A�_C�m�ࡕ
�x`o�~i`%����	\���H����{��@>Rz@ ��^��lug*��G��j�Ĩ$�b> ��զ�͓<]���1%ɒt�,�&DV�qK�ϓS-����On�SM>�/OV�d�OR���:AK1DZ:8������O��D�O���<��i�����'Y��'P>��F�2����Կms��`��'i�'����?���6Z�@Kr/	�a� X��y��'��x�dZ(dD0u�X���Ӑh��a\�Q1���Nq��)�M� u�y�4�Dܟ��	ڟ������E���'P�a@�)-;���4.��g��8��'**6�0V�����O��o�K�ӼC��	(a` ���%80��(�<����d�(�<79?�c�E�/�h�iщ_Xp9�dI؜G2��b$E�L���O>�*O����O~�$�O���Ol%�ta�@��$!c	P�Pk�4��<���i�~�S#�'���'T�0x�]	%�����)ǛXXM�E�D}��'��O�	�O4�D@"�	[��H:U���"T)�KJ�s�E�0��jt,a�n�O�;J>y-OL<RGm^'o���I��8L����'06�̰yD�DJ4�X����V�y��H�ʶb��ăȦ��?	�S����4{ڛ6d�V ��ŗKP����P�e�j9 �t=�7�7?��U����I��䧔���l���U�*ޗY&t(Ee�<��?y���?Q��?�O~f�I�c�la#�b �\����N� ������?���or��-��s���M�N>�$�?��eԦ7�n�%�Ox̓�?����?Y��&�M��'"D�%+��`��}�=�����|X�,�&����|R� �?YS)�	\tq��k�7+:�Tb�u�'�:6mv,�D�O���|Z�2����5���u>*����q~R��>	�i�D7��)��N�H�|���N�d �\�%��!�6J&B��h,O�)��?��9�$�j~��h��ڰ�KY.y9*��O����O���i�<yV�irzTz��"Y:��]�F��e!� (g���'��7�8�ɐ��D�O"�RE&׷jf�y	u�R|�u�� �Ov��H�6m2?��Gf�q1�'W||˓
j\E��N o2��{Wc�"Ex������O^�d�O��O��Ĩ|�����
=���ʤq$�T�#T�]]�V��
uR�Iޟ��OV�'�d6=����D��l\�r�̈W�5Z�L�O�������I�ҘDm��<� Zp�a��(� 3���I*�r�;O��1s`���?���'��<����?��`��a ��@`eЫ oD�c ���?Y��?I����Ħ)���U˟�����X��!��_���
�L�
�"�L@g����"�M��i)O�EE��1�� f� 4P�	唟dA��T�SN�|
C*TL�1RG*ޟD���h�&��!&fytSDm������ڟT���pE��wR{�D �BŞ��#�T���h���'`6��8'x��d�O�EnZA�i>��;,�h����Qu��6ʽ�6�I�M��i��7��($t6m+?i�m�t>���-O�`�Y�ሃk�(@*���4Bf��N>1.O��d�O����O����O�My�&�x����mC�͘���<9��i_L���'�B�'d�O��a�)6�Aj� :V�p�T�Z����f�`�Ɯ&�b>5w�y8lԚ��o��r�e�0_+����#[yR�]��z��	�l��'�剰]�	��׌D����3D�'l�D�IΟ���؟D�i>ݕ'-�6-H�M����!_g�,�V�ҥb;|e��` �D����զU&��S�����k�4w���"��N�0�g��h�"�!�G��fQ�1�e�i����P��O7��&?����l~�hb
؇W�p����Ѥn���l����\�I�|�	S�'x��؉�-�$�����Yr�����?)��S��l���d�'��7�?��V*Lb��0��/w�Š���(7}j�Op���O���]5�63?�;abHc�O��(P��A!8mH��e��?�q�+��<����L�j����Z�<�(S�X3�O��oZ�x2!�	��I`���T[6� �Od�.ܙ��@����X}��`�ޑn���S� R�9����A.�>ٜ%c�b1"��c(�[�y�Y���&qz�ev�	9��[F��3�ؔ���O�09�����	���)�by��eӞ}ٲ A�4��U
�:{p܁a<8
�q?�F��H}�K~Ӑy �_1#�h���c�Bڧצ�#�4U��M��4��D1v#���,�<�ӥ��,z1�O5{>��do��<�*O����O\�d�O$���O�˧"������PVǬ񚒫��4pXоi�F��'V"�'L�OU�q��.�}zP!9��U�0�eH�?ݲIo
�M���x��d�[v�&3O��If�C�ca�A`��n��<O64x��҆�?10�?�D�<�/OXiP���+'<�r"��],t�A�'{�7�ȣ=�����OB�R�vt�S2
��<����UW�"�(�P�O4��O��O�"m��^��X�$0a��a����CeI�(�x�c�j�ӕ)��\�����K��b�x�/͑]G� Ӳ������؟L�	���'?E"�kt>��I:(�>Ȁ�k�y��L�:E�a+!�'}�7̀1n��R�Ɨ|b��y�!�5"V �(E`�:�"��_'�yb�'���'@�c�i���O��EFJ?��FD-g��tjQ� L�ꥠe��cf�O���?���?���?���2S4P���-7�Q6��
'����*O*l�*i�T�I՟h��V�s����O���S�À�D�cҨJ%���O<��>���I1m���R�&	2!��	�R��	{,\�bD~��;���a��� %�Ԕ'Ɍ�{�B8q��Ve=�<ɐ��'>��'v2����P���ݴI���y�∘��/;����F�_Lل4̓2#�6�DO}��'��'HZU)�`F.tl:��e�V�*��!�iȤ��v���#���VSQ>5�ݲ+	&�q�K�R����.D���Iݟ��	���I����IV����D-S+y�ޥ�#*K������?��<�fM������'MR7M/�D��K�s�\�-�ĉ��̌m���O����O�	Or��6�/?��f�&�B�
=�`�XԨAqb�C5G@��?��)/��<���?Y��?�I[)VK�x�JU�+ 98��^��?I����$��},j����O��D�|:#�0%�1�C��n����jG~�l�>����?�I>�OtptH�\��j`MT-$*�Q���G�0�+���"q��i>1"')�	�4���G�Ue��G�
2�K4�g4�9�Iȶ-��H�@Z�^��������;�L��u���Kl$�PrOŬ�,��bG��,"�9�kՈ�j��fB�8+s��9��p���
u�zAaB�9"P	�iQ��:=��g�� ��>Ŕ�Q�-��%�@骷���C����8Ê��p?�	a@��4�$��(��	ؐI�4�<�B��Ȑ�C�f�
Q"�I
��1gȰDWy��营
���u"�g�|�����W����Ӥ�f`��S���� w/��:�>$�%(:�f� b��r� ��C��'��|�P��KҊ�?vL���G��P8 �#���b���Iϟ4��ny�ɓ�8��~���n�O�X���J�[ .��?	�����d��c���u��az���95��xqP�ՉE2��?����?!*O2�{�&�[�S�e��,{T��,U����&�J��Qܴ�?�L>�+Oj� ��d�0@���A�C)�����C&>N�f�'rP�,��)W��ħ�?��� @�(
�[������F T����a�x�Y�(( ?�S�T�V�_�Y�/�*�"m1�.0�M�,O�)	P٦�3����������'�p�R�ĭf܈PB�����Hٴ��䄱��b?]�#O�'�����+w��e��duӞ!��#٦=����,���?8�}�NX�u]V�Ѥ®W����Td�+h7��'��"|��5�X�[��W"�h�J\3`="�"a�i���'��ַQ�
c���	���� 6�����,8U�2,ρz����@�1O��D�O�����5!`DRgC�?Kbu�J�j���m�̟�CI�ē�?������s���5��l��F�EJ �A -�W}�,���'��'��h{t�Uo
��!��4@��1I��`V̨%�����%���';^�pg ˟@�$l��jƼh�f���յ�'���'12Z�@��+@,���d��f��ԛTJ� VP��f�����?�O>�/Ob�]��SF�{Dy�T�js#囫��$�O@���O^˓]kM귖�tF��#�ʸ� �]]��"�gK&s��6��O��On˓�l��>�5�Ѵ5�)����;�ư0�)�ߦ��I��ܗ'*n�C:�	�O����4u����M�м@ǁ�{.i&����t�X�g*�1YNLpe-Ջ�7ͱ<�WD�(��&�'�r�'��s��X�!���&hP8�촁�딎"p�6��O��K��f��!�$8��"vN�����;�I��I?&�7�^$M�<o�ҟl��ɟ���1��ĳ<�#�~����"5����#��(}�+P���On�?��	�B�:�`��5gjY��d�7' ʉ�۴�?����?���9Uq��uyb�'���ya@D!d)N"J�;��E5Yg��|��U�2_��������i���4
�O[R�*$�ۿS	D0T�n���d�B��x�'����d%���/���e��AwP�òh��J���H4�?�$�O��D�O˓Hg�ə�m�ni@Q[Fi�
n@��`2�ٜ���sy��'8���t�	����B4D�8�:A�M��SG/L��\'�X�I�$��oy�b��U6�S�rł�3P	C�&V��#ɕ4�.7�<������?��v�vs�'+�*�:A���˾M�t�O����O��D�<3�̿h����*���[\�C�'�*k�b�R ���M;����?1��Eΐ�b�{�K��>�j��e�TZ����ˊ�M����?+O&)�4C�_�d�'��O��P�A&~���Ŧ�&V�,A{�M,��O��dѷ+�:�t�'E|� �"S�]����"04LAm�^y��ô���'��'���X��X1[bF08�%D$$���c̄ p%B7m�O�����4A��b?�"ǣ� ����f�3N�u�CGp��C�@�A�����	�?=3�Ol˓���R%�B�SʤXǄ^�#�T�ƶi�8��`�$5�S���ӎ�n����Yz��xc��y���o�ğ���ݟ@s֊�����|���?��킀.�*(ha��b;���ĬJ�sϛ�',r\�${��X�'��i fm�g.���H���,�'e�F�h�O4�)Ub�<�)O��h�פ�:>"B� �Ο�~���0
��ē���<�����$�O�P8f���|�@	bM�Ff�(ia$��?1���'�2�O�|p� ��}���+�����i��8�y2�'���ߟ\;�or�#$�T����H���S��������D�?����dY�ěgQ
D|�s��!9N���o
���?1*OP��PA��'�?������[���t�B��T&\Hڛ6�$�O�ʓA�m%�(����K/>=y!�X#~��;$v���O&��rA�Z4�ħ�?����#�+5�����*}kTl�G+�h�Ky��'/����u7��$/�h���M_V�B�)	�����O�S�
�O���O�����Ӻ�ԚC].�jt�Ɋ-� %�U��̦���Ey��N�O�O��e���PZ	��m_�h��H��4�&9��?���?!�'��?����e��|(�86mX�����MS��Jp�|@�<E��g�/�Y[#ڊ'���Ԫ[�Ur��'+�'mj1Q5W��'��$*"$K�!��n����2���$9��Y�y�+ԩ
�P�d���O��d��a
^���o�Z}���	 y�(5lZ˟lۤ��&���|������O\�z�cWT�P��0b�5l�xMC��D|}�'1;�Y����ʟ��	dy2�S)(	qul؊XݒE@�s���;��2��OD���O�˓�?��E����`[<EF�
SI6J��Y�"���?9M>)��?1-O��u�W�|"2�G�X?�ȃ��=��B��a}r�'���'T�៼�I+X������
x�].4��bg�ߝD�tl�$�ۑ��$�O��$�O�ʓ9l������T)1?������D�D?���M�%z�7m�OԒO��P��}����S yW���1��9A�h���ДZ�V6-�O���<���ۼ_��O\���5&�E>90��3�&��=��J�%��ē��$ί���8���?�����\57D�%��+e���E���h��i�R�'�?��2	��(>7D��"�=l�����#<6ͦ<	W�X��?A�����ܴDg�B6��;`qީ�f��"L�2 lZ j������0�I����{yʟ �$�H��Px�O�"�lh*U�צ	(Gx	�����rL1�����h	-|xy#����M���?���ǁ�'���|����~�̿ta���x=<-�-Z�0�BP�H�6�]���9O����O���_�8��]�#f
M����0Z��m���lBE�	����|�����Ӻ�gϜ"�!��L��3�� ��X}R��hv�U��������	Vy2k��(p�G���(p���oďu��i��"�$�Od�-��<�� ��ҀC̣M{�,(q�ݟM(���d�2�?�-O4�D�O��$�<��H�
N󩟡K���剓9P^6<a��[m�I��K�	nybhU���+7n��DD�h�,b�� �ꓼ?����?�,O����P��'�iʥ����H���p��\B�Fy��d�<a��?Q��#��<Γ�?A�'y�9�G�Qyz�G9�l�۴�?�����ě">�L��O��'����^(S������f� ���N�!���?I���?Y� �<�M>��O�B` �%�!a����+z�۴��$Ļ��Qm��D��ោ��������(V5/v�C��
Ct<m1�i���'�L}x�'��'�q���:e�,�d���N��}+��i>� k��rӊ���O����"X�'���'[U�<I�O��>�ry��0J��u!�4[������Odb!I�y(=S�E*c�j,Ҩ=��6��O��$�Oxi�G@R}�U���ID?顭I$�ek�ȇ�A��d��æ9%�T�Rhn��?q��?aI��u��%�G��\��������'S|1�Ģ>Q)Od�D�<Y���.��y�P�c�(��%�ԄSLUT}����y��'���'i��'h�I�S�<�ˆ �ZnZPR@�	d` ��r�����<������ON���O��鄭�G��)��G8;��Z�c���$�O|���Ov���O�˓~yJ�X�3��@ 䢔�^� �(���5)PH�Y�i��	���'���'���ɴ�y��ŵОɚLF�i 
�g���{{�7-�O���O��D�<	�o�4d��ܟ�X�p-�1bSl�6���D�3UL�6��O�˓�?i���?�Ed
�<a+�f���@t�����9\��,���ͦY����'_�yK�N�~���?��'^��!k �Y䄩0��(fp�(i�R���	ş4��-3c\�'��Ĺ?��QF��3߸|�gD2k�tbc��ʓo]�]K�i>��'���O��Ӻ�&���z���jb��ECrͨ�/ئ���ӟH��m����yy��ɐ�G�Pc��rl��� z�f�D�j��7��O����O���y}r_��RwhփDu����)Il@� ��>�M�&��<�O>a��$�'BI�J͌ڌ|	�팜GF��t��j�D�O���'����'�����p��I�f �y0�my"��%�@!o����'w��r���I�O����O�k1�dct��g��VP����U��0�N��O�˓�?�.O����-������d���MxtQ�d\�Ry�ȗ'J��'�2_�L3R��Z*H�X$�Υ�z�a��G����O>��?�.O<�$�O
�DC Z	��҄
��֑��)Soj��0O�ʓ�?!��?�*O"Aڶ�M�|���ɠ���Jڃ[a��������'�B\��	�������I�AT����<:��Rd��-�V��Oj���ON��<a1LQ����'�4-�I'hd��q���M�����O����Ol��$:Oh�'[N$u�D�S�����&gOrR�i���'��	6=��ѹ��f���O0���u���i!�) ��}���[+O^�'���'�����y�^>�	k�k'B��c���s�`:�h�⦉�'߾5�Shs���D�O�����`֧uMXyμ��O9y*<i"ҏ�M#���?)�"��<�W?��yܧ1BT���;��Yc1��T��em.-��:޴�?���?��'"��	my���+dP�3EO�,H��#¦�\(B6퉜Fh�����2D`b�D�gr��$���Q��iYr�'���
�*�D����O��	&(��u�D(F?u:��Q�jV�IB 6��O�>@V��S�4�'YB�'��E�T�ߙ w�eS#+�-F�B��s�a���䖆{k���'����d�'�Zc���W��,�Z�;P�M9r����4�?��JI�<a/O����O����<���T�0 ���6��R�U6F�y��Z�d�'�2T�`��֟����?��@5�? Mpk0��W��R�y���I��x�I�X�I}y�B��+^�擾(	���b�> ��-ѤA��6M�<����d�O@���O�a @=O�i��E7ʝ�U�A$ r>��qGЦ���ן��Iʟ̖'��Q�tN�~����E.�9{v�(hǢ؝C&ԱB6I�̦���]y��'��'*()��'��I�s�R�>���w`^"7��H{ٴ�?a����d	���$�O���'���JYj��S��	8����J Lf>��?)���?����u~BP���'P���:��y���;�%�1�<Yش��$�:�8�mZ����ioZ�?��O����T�1�ݜ3�TY�D埡!��'9�
��y��'*��'dq�� '��u��Z�Ɏ_-J��$�iz�+rӼ���O2�D���M�'���6	� �w�ܤ[�*X[gZ�EGD͋�4^�JM��?�)O�?)���z|p�r�#�x��j��β,2���4�?!��?Y`I&��	Cy��'���`Ί-9T� 2c���	'�F#<�V�'��	8�2�)����?i�`��ѽA��rA��?��@#0h���M��4��uZ�W���'	�[���i�����8�>Q�8B� �1:(�d��YΓ�?����?����?A(O@�XR$E�@:�`���Z����AE�2D�Y�'���ҟ�'�r�'JB�A+
�V���zb ����%1^X(�'���'&r�'��s��fI6��D���҈s�ߴb5Hf/]��M{*Od�ģ<q���?��a�\Y�$"H��B�g=�m�!��(",< �\���	��D�IQy�F>-�Bꧦ?��"NAX�`��ns|�h3�ȣ_͛6�'���ɟ������:�j���	�
� �Aj�!�j�����^���ixB�'��I)�"�⨟����O����H����cMW�5�|m�����G����'���'�B-Y.�y��'���T�P(
�`��0#��9x�i��cĦA�'.����#s���d�O���蟌i֧u!\p�\�Fh;~�����޼�MC��?�0A�<���?�����O؈H e%T#�n ���*�-�ߴ_�0��W�iO��'�r�O�O���)�6�I����\L��O'j�oڭ`�*�	K�F�'�?�G�b��D�3$'�r���%Q�pқf�'r��'�j��!:���O����|�Ʈ�:W�(��c'�

=^I���w�ГO0k�aUo��ܟ�	⟴+d̉1�8��[�
��%��n�؟ܪ�â��'���|Zc��AC����(�pq�TKR?P��ڬOް���O�ʓ�?�����'<��
Uc�g�(�[GI�	V:�b�٨,6�'��'H�'��'�
�R�E4#�l̘���>@��@���yr^���蟐��yy����F擳az 
�#�+0���1��R��O�D8�$�O�D�Y���A�5В�zs�W�"Θ���زK4���'�r�'�V�\ �����'d��"�jS�hԸ\�@.H��<�y�ie�|��'d�����>aAʋ�,����� J��yk6˂ߦ���ܟ�'�&�)e+5��O��ɉ�.�b۴ė=w�z�)��2C�8}%���	�0�DL̟�&�t��j9���U��Z����L�-g�qm�wyBI�f�h7mW���'���6?9P
C1D��a��eY)��Ś�֦e����`*�e���&�(�}�R�܀	$Z�0@�-r[i�eM֦Aa�Ė�M����?I��%�$� ����`��0^ü���	T*1��o+S��	v�s�'�?�G
�N걑�����%��3қ��'��'H5��):�	؟8�)�8��S*��XH����B(oF�IBb�)R��?	���
�q�e�:z���ک(O4�ӻio�.:2GDc�<��U�i����$�&y �)�(��@�JJe	�>)��έ�?.O��d�O*���	�'L��}���B��\�� ���ǐQ�dd&����ן�$����ן�
Ц��{0�=;�#�`��!����Isy��'X2�'��	;@X !��O�6�3D�m�0����&m����O����O�O����Oz�/�y�ΈT� @ �獯d�tř�$�_	,��?Y���?A(OVt���Gn��4 C��F�L��6���,�d�F���4�?aJ>���?�o��?iK�t�1�J��>��A�9�T}������D�Oʓ<����e��d�'I�4���#����fB�A^�=w����O����O0�� �OܒOz��n�eQR�<����5 ҭH� 7�<A�jL,P��6�~
�������	�xєY4 ��#����%a�<��O���FG�O��O�>�f聽M��桓6h,TH[�!~� A{��^����I˟`�	�?uH<ͧX�����MO�)��וn�ms�X� �If�S�'�?9H��4��4��P�%���E�<;�6�'^��'��D��<�4��'T*�HnG���/��aѲJ��MS�2$8�)�O�D�On$��fр�@���+��N2df��Ԧ)�	4(pE	J<ͧ�(O�hQ&oա9.�Da�$]u��xE�x��'��I���I���'�E8 �Sy�`�sa ��֢�P�KS�8O����O���<����?S��L��a��̐h|����/r��U�<����?�.O|��O�}���$�V�4;C��t1�q7I�H�>�m�۟����`%� ��Ay.��M3J�r��Ju��:ޤ�&K_}r�'w��'X剼h��5�I|�Č��6�Hmt	P(H�i7#D�N���'��'����=. >��coä~�Ryi����F��7m�Oz���<��mUt�O���O>,�m�`R���g �<[|d)%<���O ��'[T�L�'~�Q�R"7�l�A�*�l|o�|y�#U�u�6-�w��'k�Ԉ*?�@�%C�:G윒,��P`�ަ��	����:��O@�DQ䓵_���S2�
�j����4	(x���?y*Od�)�<�OS��b!�;e���Õ䒖3LDܓ���>Q��Q���O��#ۇK 0n��#9�[�06K�O,���ONh�Ɵ@��ß��{?qeU�+�`s𩅡�d�(0	�y؞@�Iǟ����&��9
� Ƹ0#P���a��D2�4�?�5CJ&�'�"�'-ɧ5�̝�D�|��`�;L)&�ÂE���F�G�1OF���Oh�$�<qU�ęF�=���72���E��a���x��'�b�|��'�2��4�j��O��I��l�AG'wb�ۊy��'02�'��	�h�|��O��sK�I:11l%J�j�K�4���O˓�?���?���^T}�.
�Z4��dn.�4��C畇���O@���O>ʓS�	�U?]�I�Z�l
�-���ܙb�
2�F���4�?�)O����O��D��z�$�|2$-3Q�UcEiεX��ؠ͘�����'�[� B�#��	�O4���D�T���]!"���N�h�}�Y�(���|��qo���P��' �IU+��р�舕|�V� �%�4K��vU�,�����Ms��?������U���5^x��T5e�� p�mI�'�&7��O �dM�Q���d��'�q�� ��"���B�l�W�A�= ]�C�i"a�A"|�\���O��������'�	//�N�����-P	�$�sN+Q��K�4� �'��I�'F7>yo� q��!�c�||���"���p`pB�I�>(��W'eӜ4i�A��D*^��Dފjxx��oV��Q �,"vu�0�����`��@�c,z�`c�P�_tl�qm
J#���#�8
&չ��ʝ*�N  �
� ���0F&1f�[v��:�X���MuH
��w�Z�{2�b���D��%C:O*��'�C�-���PrFCK"����'IT�=x�% l��'nB�'��� �'b�0�f�w(}���$F�W�r��*�&� �y���J	�|b�~_��P����������J�F�V4��DQ�r�'��k�h�:h�����f����@�|��'�b��?��C�)�� "��(v*��+gk D��i��ٴt���kQ#2��p02h`����4�?�-O��˅e���'I哙'eB�ˡ�ӝsU�"�ʏm��[�)�����Iݟ��# �%"�%����D`m��S���E�h�UBK�0jL2�X1�G�(O��`CȲxj�rP��(j"��x`�&Q���˘$NT8�Q�I6���Ol�?i�dN�X �lYFB!@��uj��q�(���+m8�`��8NwHc0*����e�	"H.qA ��!S1(yԦ��8t:�Ie|V2�OX���|���� �?��?�HT�.����;	��ы⢗)ښ��,߲vJ��CP�I*�c>�dC0L똝�)I��,��r�6D���{�LLɰiN����)���(�x�|�Â�Z%Ĩ(5&/x�R �I���'��(?�<��4{�BH3%�H�l���ȓHn��6C���1�'�2�~\Fx2�*�S���9&��c��D����E�K��'���fа]W��'Y��'� ��֟�ɚ��j腱1���3���y����pHj�����]!@��Ơ۳����99�B�U�ָ��I�R&��:DA��<(�[�	٩j��	!R����OD�O����OH˓\It8@��>;Kʝ��$�	�� ��-bS��[�N/�8�4 K��+��)R�ʮ�<8id
����A	3�y�XD�ĉ*�iN3��<�$��y2j�w�"���ي�H����y2�I�f[4����fPf�j�c]�y��2$��tyRÐ/XZke,��yB��*p��iK�A(M�d%��y�Ǝ�F_�Yc�m�-�x9!�ґ�y��G
�8ZG���Z�ha*��y���q}`�s�]0^M^��U�G��yb��U=� �șOr�� �'�3�y��TTc\�J��ËE��t0TgO��y�#V�~��1��Í6���-�yR��y�TT�3�.0L�*�ŝ�yR�T�G���6�����i8�fA"�y�	��XgT-�%��O�����[��y2��:94���D�%wfrx+����y�-F
.ߨy(v�G�q��AG��y�k�4T��Q���e�֝�qo׵�y��0d�H��O�R) ���"�y�%�4B�5�s!���k���y�-��>&(�[w옳d�Ѱ��y"��U�q����,Y��P�����y��"�����N-K3�y�h��4�`���ńKf�R��+�y��xx�J琴�j�)A!�:�Py�,f}R��OܹU�h!�U&�[�<AF&�)� �{QfF2):��3%c�T�<A)UFv��7O�4���UR�<��S�%��y��֫P_&�ɦ`�F��(ڦiخ�N}�@fB^�5�Щ"@�4��gH<ɴ�< g�H�I<-��АM.�k��tΘ$1ј�>]�F�[����Ī�ݠ�x�O?D��	"�M.s�Xi+��+T�@�S�M�`���0���v0�H�F�i���G�,OT�Q�8v��	p�*� [d�P&"O��ćdbIЁޟ4�8� �(K����B"��D���Kw��)�p<� ����&:(���&�Y:AG�݀ �'�LY�$��cXnA���7v��T�n�+N䮅�,�6�y�A\e(<����	����Ap����J̓������i���r�I ,�
�>��o�zM����MG�p�X$�5�"D�� n"Gz�=j4�;kI|`i�,`�!p��̓�h����1?�|������.%f�69`,M-5�"��$��b�<��i����#p%	lѮ��c'�@��ZRX�\K��^�A�>��N3?��OB4CJ�o�u IH"TD��'��E�@P%UD9
�Y("�^MK"N�3�j��K�04 &�Ŕdb�2ס��=�Rj�%V�x`	�J�i�VHƪ�H�'�FQ+1�����z�m�+ %a��?��gH�l��(a3I�:E��"e#D���eE��G�:Ⱥ���Pƨq��}ӬI���N'�>���n�<�!�(�k,��,ܙp�pWZ@��U�F�!�؈ ��%1�ע2o��cu��s���
��N�,(��W��:�W?�p��d��"�Q �f1E���K�C��1�a}�D�2[��l��K5'�r�J��,An��nF%i��Qq�"G�D��0��A��L���+/j���3��?E��ҭ;ғ.]&�
P�7u�p�����b�������%!]�|�}r�Ñ1(����p"Ot9kgr��QVCS*�h<#�i��m��J<|JjiH+�'���p�S��5��Wm(E�� �`�j�奋)�yb Șx���mn�j!a��^�����0�R�26�P8��Q?�s����g�D���̡_,*��R��+Ea}��?
ѳ���GU�Xbb,EFh|��o>7�]sP��fFRec`��W���3	�9i��bK��6%cw*ғs��� ꌔERN	��␟�����)S,7/��d��DW��HRw"O֕c��0�nţ�d��2�ű���_�/aV=��@mS\$eM��S�I�2	���*W����Ԉ��תo��C�	  "$��c:��,�E![/;�^�(R(�&�qš�����%§���	�B�� ���.���j�,�BB䉵l*:I �� �؄"U�\9����@2�	pŀ]ΔA�鍕,�Q�8ʑ"K)i��;£ٍHR���E�-LO����Vi��ݠ��A�T��h���P$�Qҡ�{6���N�Fx��2��<�
���p���@V��<q��� �V��W��!_�09X������O�����[@�t9��<O�� 
�'��qR���KXJ����;l���8g��8���D�j<�����ة��'��ѐS�I$\�i������'R(� CU�t�l ˵�ߐ�|�[�L�TtI������×��R)D}�L2U���d�6��Ht�_��0=1S��"[Qn%����l���@�Ğ�Z�09�dT>��d�7�M)��8�A#�O��c�	�v'�1i`�i�Nēq��7)XNőu�M�xv��is��FfJ?�1w �6d �EՆ$e�屡�.D��{�*@�.�������A^�D#��-U�V�(xZ��m�O�"|�BF���2G��C0mJ�҂Db�ii@=D��a���uҲ��q�NR�FD�1x��)���:C�B���a@Lc�'�p-�B%H�s��1V���J�����'K�!�U�Q�P_�lb"@�� � d�%D��I%,�~$�"�G�V�tqs�M;6�`��D��x-�<�N>a��4*3�s��MqU:XA1��c�<	� ����}Hu�ߋ'����e�ɟW��9���鍟]=��c��2U=�dsb$�"q���3�|�N�&�&���r�Y�.	U:�8���!�	��ұ�M@��*D)��tk�Ze�R��dE7:��͓Q.��p�%O#uFFT���i�*��}#��bME�mW��!4H�U��%ԎN`VT��DȄT�:x@wA�)Wdp�*���: t��W���(����5�h)��BO'Oh.�sa����1�|J��1j� �P'�C�N��A�#\�� �O�"�i��B	CL�u�s�
4fԢL��d�/묵3��G}w�AaB%�]��I�4�#��>�jأm�dQ$�ѻN�yR�he�'�@-;4�Z�(�T:�����#�ʨ�4�U�^�~䢠K�+���8��(������_J:��P����Ԍ��)N,��0a��-{6��
�r��D"���S��.�=s�ܱa/��w�T�)A�_�g����H(xĮ���üRd�D���13*��s�<'vࢢd�1��\Q��+�Mc��X\�r MŬK��U!�� �^͂�E�g��ͻ	��c(@�Ԅ`O�s����ɻ]YmP5�	.�(!��J��0.����^*�aƁ)e4�I��P1{��K�
,�8!�TJ����Y��0��<\Đ
ْD���"�)�$Y����R[2�I0WX�3� �P&+��<%4�Jp`�(X��D�p�r��UNK�dǖ��#�X�O7��?�gNM�\s��J�9�$ �<����7SҸ�P�L
�!��?Q��#�bY�% �ÌX>�i1�G�Q�<�{ЇT>{�v�k�kA�V����Q���$�@Ǚ{4�EO<w�՘ ki��x��$D4$<&�<�ϰ$C�z��$��&��NG:� �0��`��	!�N̯3�a~��֛]2��y���<Z��"�E7r�v��� 3"���c�"�Pu!Ca� -q�1%��>����D��S衐�S=}�Z�`Df[)<!�D�Φ�2�j��c�*yZ����1��}Y5j�O��8 ���%�x��ɷ#���$ýߖ�3ɋ����sP"�Dџ|YRn�Ħ������V�.Ib�O�+�bx�g�;�8��	ގl�hCF"��?��" �-,0���.X�=�1kˇ����/}Xt��퉮�.у�� �+uHT�V���`\!�HL���:�z�k���y�Ǟ�"3p�B�Î)m��D 7Y����j��p������Kv[���L|2��εHd�!�'�����A�}0�����F)z֦�����(��X�W�2%Ćb�Ū�fL.̞zu��PMj�O�>��� D�Hb�'��\S�L�&����Ɇf�������$������YE65�`$w�	S�\�p�CE���~��<;&Ŏ�5}ܕ�@�'$H�J�$	nu�b�c̞%"�'�8!Kt�TS�$9R$~$������x����BV)s�<�`Q)�� Y!��vk,�@�*�2���h7bZ�oS�W�����fԔ&_�f�[�V��?���M�UԔȢs���Q
��CX؞Г6B>6V u
'i��L�V��&�4X������9z��}p�fޟL��!_�{2�X%�hP!�ȺYH@B����'�HA@��#U�4Sv�5R����<�$U_��8a�ݵ�x��cA�g�B��4>�&��شa�L`�� C�D@L�`���L"��2�H(O��Mk:���u%8S���TDĊ�O�yYuE�{��b�)	7r��E�����Y�d\�B��џ�@��>�O8�r�� CC�Q���` *5�'ÎP���7 �!(1�C;
}�$'��,C���6�F�xԚ����?�6��+.�l��AȚ��΀,g�(��x]1O�)��
,8� P���Nay��gy��*L����P�'l�q�LE-W�����[�^�{�>:��DI�A��L�q啝����S�qϔ�O1�Л�w����I׭8[��`5˥/�����g�>�اh�~�ٲ+�M^K�`�*LreX �>!�$Ѭ
�ȴ�/�v�����˟�$�Ȑ���Pa�P�E94���9w�:}r�݉v`���<�r�ͩ6ఠkw��Y�\|���ˤP��MrU�O+<i9�d��3	��M��E����4'�qGz⍚1��m�
"y����c��9�j���RU̓y4j���B�l!� ��	,l�湦OB7��c�8��H�� ���"�x@;���|��D��^
�@R��ב]�hhK�N��N��u� �z�ᄖ���	H?�'4��λ�t�	S��3N��T�ï�p�,��.ԎQ2U���@^�0�"�G"�>Q�#�H�d��+�$	�[ ��c�MįbĄ|�rO6}�JFE��!bZ��`QĖ��ɶ VE��}�%�Ѡ��j[>��)�ԍÛ ��<�OåxЦ���ڔ]8�V�ٳ(p4]�eJ���#=iqlK�*��IjG�
e�r!G_�[AD�!�,�ɍ`"��SN"���4��A��%�2�����ƶ	����:�XZ����0NN�E�����gs�m4 	�^:��s
_7&�~9y2�	�-%��''�ta�w�x4AU@G�b���u � z3�1"�'2*�P��&�)�'�p:��]�x�`yc棂=|X�O�����W%W�z7m�a�mi�&.��O�)�'~����ʰD
�>I���1D�O���pA%���:6Xf���D�\�	ۄA�k���ی"P\�ʐCa0ibs�.�2_��G0C�(9��_>U�IK%�\��㞤T&U�	��'��H%���祅�&�YG��1��`�t���5�k�����"§�	�����sV�0���6������ɩk�l��O�p��#�D-	W��p"��w��|"��O����Q�����I��th.���:o&@����0���� 	�͸G�޻I�D��>	`l��������'%�9��"�4u9

 ��J�h��K�4h� ],���hǧ�0�ا�ɛ�2'r���@�*���Iǉ�)�	k�"*����,,O�],y���+g'ā�U%D�8�T�{�L�13���I�}���/θ'���ff� ~�l��kY;F?Tػ�'E������U@��f�8�b�'�>�B�`��4KP��?�}���34$�s��2(� �%fq8�,H����~r���qp�(��m(��&��'�Ҥ#��'��W(��G;BeC5hA|7� ���d���F��/Y &��@*�-
nY��D\u��% �O� L�b7d@�E@\ՂQ�M�X?�x�S�i�,�4)��~2�G_���YS%?D���T`F�h�ȓ'F}��M�,�u(�(�Ext�ȓ9&Aҧ�Y&)d<Ї���tt ���*����y��q���?\|a��,�l��i�nS��Y�`=�P��P{�e�rn�5���dER�3�`�� �!�bF�.�q21n�O
���-��l��kK��l:���N�6��ȓ.��ݫ �wu~���ԏz،d��x:�)�$ܨ_����5E�GT�1�ȓ6nz4��d�3+�<yU��%@�X��43и�G$�	9�*uKBo TTn]�ȓ)$�J�P���b��$S�&���?��P�Ѩ��$��83C�EAm��B$�}a�/��/D|h'�[�ұ�ȓs�(��T�a'�XK�5ɖ5��.w|�ڂ�: .4@��HZ4�pm��d���CU/� `r���SB��z%�ȓ<� T���b���k�AƾC ����a��Z% (Qk-�j�(Q��F^�8s�ʾs B[���N!���ȓ�(��%^�;���B����7�Z���~e<�V���;�n�J�%�:X�ȓV���'�ȵr��)2���4,��ȓL�0��Y<	A6�B`ElE2�2D����.�LK�iS��<G�ѷ�;D���Q���C�ڀ�eE�W�ơ��+<D�����3;��5�&B�)�eؤ7D�xI��W��-Q��]�Zw6��G�4D�(ʳn�D^Vlk����-*���,8D��"��xj��a�ܣvm�Ѩ��0D�,��nL�?�:A��[�<J��)D�TR7G<n��`c��]�
)���;D���eʗ.6�>��@��hŪ`1�O9D�ȳ���	a:*�[ �C�'~H���j8D����
Ц��#w�,-XD��"D��&X,Z�����'.�0tP �2D����Vc�j����M�O�*xؔC2D���#��L��	w�ߒbT2[./D�2�ձ<Bxa��^�&4ԙ�f8D����!f��P��o��h��*D�H�!��,W�Y�w�B�k�A�*D���𧚾�p	s�`��><ƙ�4 'D�I1	T>�f��GȎ�d�����1D�L�Əۇ]���.i\�lz��߅~�!��Ү<d<�wf̛fD���D�4�Py�`M ,�!� �iV����j��yrb%xQ�&���b�B)r!/߽�y2��<x�F�!pJ�"��F��y�J�,>���l�pBʽ8�)��y�L�7)&����,ٽ���y� ��y_�)h�x��'�%�����$¨�yB��tUt��Gڪ
�R=Z�_��y�"Q#�������Ţ�C�yr�(�n�X&��)R�J�I�3�y2��)M����-��"j��BV��yb��:���8)#M������'�������+�OӸ;H�X�'ר���E�,%��-v�:t�N�<Y�"��=!Rpk�m��,�8JGiH�<)�o�Dݸ(��K�}���a���D�<�w	��
� ��dF�缵���E�<YVǜ�%y����m��i�
<A�Z~�<� &�(U�ۦ7 *���훅?W�T�S"O�<����8;�
�R��	NI8aK"Ò�P͞�KCBu���L@�UA�"O,����e�����ǀ@-<9���(|O^}�b��q��a��dP�oFT��"O�1����+|Z0��-��2g���Q"O@=����
���p+N�~lNU8G"OVI��*%�����  /�@8iv"OZ!s��	ƕ�s�D�]Dx��8Oz�=E����/M�L� ��|'L����	�yr��m���$�Z/t��l���W��y��Ʃ.m�y3F�oh�L*���y�I§Y�*��1Kb��x����Pyr&�G vp��G�$�y+2�<Q�].�! �1e�Ts6��`�<a�����B�#��0����E*S[�<	�FF=`��0�ЮЪ���1hT�<�cWf����q ��<�F�{�*�G�<����$h�TH���nU\�0���D�<���(F�h̛b��L�ν됪�G�<�rLN�=��и�CB]NmR�D�<�����f(3�bU����'k	D�<)qh�9���`�A�k�4�� �B�<A @�s/:�x� ]�>�����{�<�i�U�bM8cb���NT���w�<���X�mV u�
0Vh�=ɷƓp�<�毝�[�^P`���s���h#�Ul�<1��_}�4��� jźN�g�<��&v�
i;T�6P\����m�H�<ɲ�
R�􁙤l�4>���Ȓh�A�<�bmS8�(	�I�O������B�<Y*ٳ
�&�!SA޽'� � ��@�<yTB�, ��\�W��7QA�肱!w�<�V�ʨ�ȴ��.'����&��\�<�T쏓)�,�h$�B���HVdY�<1�aW�}r����b2~e����W�<��OC
~�`xiDڛkX�髣dGR�<1�I�	v&��oF�*����ëTv�<!�K��~Ȅ�#q���D �ђ5`K�<qGa>h��D#�f�H$��%\J�<��c�$fh.9�� ��"r��L�<��LT�r�>��t���^L�<&ߦ^�<@�F�Îj�T���K�<��#�1���A�y��Az��]�<�щڞ	]Č��-�By1��@�<yr&H�&z@9S�ǅK���p�UX�<	��U�#sʑZ�lHWo�(��Q@�<�]"3��2p$�7�NȠ��@�<�Ro�<lDÔ+��c�84Zp�[V�<y�aB���� �,�ҭr��T�<���_�z��h��
�i�v�$�L�<�v�[�qixy{p.�}�j9�A�c�<qc�T�`Gt��"&�#i~ A�z�<Ѧj<FX����`��`~��H%�Y[�<y7�\���T�MP�\����Eb�<�+�:$@�!f���iT:| !��t�<��tT�qdHa�L�S��U�<q�ě�5��D׌84]����jW!��qKh`���w�H����	�!�J�B�C�Gє�8D�-b�!�Đ������G�"B'R-Pb�17�!����p�7���	���� �0U|!�ĈT�\�P�͚A
ęx�� [F!�DY/JV��S�V1��6�P�e�2B�)� FE҅�А{�.���F|Ur`�r"Ori��� �\�
���8�^�;e"O�;g��<u��� ��U��Q�"O�� sG�&Da���piS���-Q�"OpLs�5D��m��gT?b�1Z�"O��D�+����DF�x4�4��"O>�p���4�r�Y��[%-�6n7D�<y�Ax�۵ �dd[h7D��@�!C6��(�׭}9>[I#D�\i�%>����N*� �#%?D�� �(	�-A�(�oљm.�c��On�=E��d��H�Rr'�xP�����?z!�d��@D�4���gQ:�!��L�$#���I�D��兜'�!�ڵc��8�K��`��{�N7uZ!򄛐O�r���ω�e�2�{�mOxg!�$^?<�֐��*P��a+T���*�!�D]$<��DI@���,�z�y�(�=�!���߰}��)R�.���aHŰQ!�$^�-����f[�@�D�����
Z@!��O��X�BJ	+-�Vu���Ȋ8!�$�"�D�bjG�N�R��B3�!�D�-\��@f�ƥ1�xL(���?f!��
Q�Dl��Ȁ�0P(5A*Me!�Md�)Ӂ��Q��b޶+G!�^12��%�&o��@���+]N+!��-��q�!��c�n0s����~'!�DQ�gT�A��p�)q�	
�2!��ի7L�eb��͘oY�(��ƒ�b!��V2��l�񥉏g&֭[��ƟSM!�N�H&\l���@u �8Q���d6!�$Z�Vc���a��G�e85$�p!�B^� �� ۷7�����!�D1J�P�� %a�����k�!��Z /���D�:1�P��d�:�!��:YMεe菋��ڇIQ��!�y�R�'nP�Nؼx@�E�LL!�U5Gw�U�ƅ��3�����'+!� "A��5	�ဴ_6���	$�!��]Ƣ���CY-mO^"" ��!�$�p��m��@n��Xp7i�!�D�/��q¡��$%Xv��o�?{�!�d�
?q�P�%�XE,�y���`�!��Zi��	w��;3�LPN��e�!�DFx�<mB6蟇<<��R�0,M!�$�<$��6#[5	�@�E�/!���W\���D1� �rs$]#!��\�X~�P�1��4��"��!�dJ2�Ze3�E�k��͋�"?~�!�DˉN�0��S�M�:Ҿ\p���q!�D�v���@b˙o������2o!�D��k�B�3mI"�8��ǄWj!�d&�\�9q��^pp�c�	 j]!�D�#�t�ǣ�7dc�+/�K!�䙧1T"�GITQTY�T�V;a"�O|�)� �f� fA�X��Yu"O��A	6m�����|����"O�,JN\_o�d��o��|�,�W"O��X��kS"�z��ӆ4{�%�D"O��R.�e���brU�g�Z�6"OƘ�e4"]��"-צc8�PG"O�)R�ʘ�{gY;�l�0w���g"OJ 薭��NY�\�P�M�!�(���"O� ����	��܋@�١�&Q:E"O� ��K&KУ=�8�H�N�tL3�"O���"�6 7ִ��G��p�p;�"O�(Kp�#<���(�_Z`Ÿ�"O��	X�e���R+��g#�iH`"O>�a�#���0���Jt('"O<�b!QL�D�&�k�`T@"Ov�sj!Uj��Y��"��7"On�iD�ُd�X};v�H�=~�5q�"O6�Bp�dB
,��!Y0Pĸ\�s"O���CxbЀA2^�� �q"O��@	Ǽǘ�pmO�F��Z�"O�8�'O�nZ��a�ˋ�w4����"O�Xj��U�|L����w��k�"O�5�	HNf���#T D)��"Op�@g	S�B)Y������	1"O,<Z�UB?칑p��< ���E"OB`H���1�p��
L���"O�a���9W�P0�Ɛq���Ir"Op��$�15t�QT����"O�p{��b��a7�σ)0�8Qu"O����JL��hH:�� ��"O��#�˶'m���Ƿf���V"O,�z��_�\���'�d���"O�%kX=��z�&�
�p=��"O.Q���_ $�D����ۂͨH�$"O�Mڒ�"H\r�x�C��D��5�1"O<�����8�!`#["jP��"O8$KCN�9g���L��y�"O��K�W�-D ����� ���2"O~�
��ʶy� �+�h��X5���@"OHD��A"=^�0@v���(�"O�%�6=��ٲtϊ#h*�B�"OT���.��c\�9�7���A��y�"*O6]��	?v]���H�|���3	�'�P�A�_�6MX�\�+N����'iE�j�U9�l�n���D�J�'6XtUE�fZt�2G�"/���
�'�$���A�7�ᘁ
�������'�Ȃ��B6\c��;DG� ����'v�f���t��t�I�r4��	�'/��"��N�L]��Ԩg]F��'v���$ek*5"��R;�D�'^���mߤ<
��@7����'J�� Q{RT�����0x��' �0��n�)Q�p���ɸH�����'P�`ғ�Еvռ�1)[��B�'���I��Ĉ-��5�qj�]:��	�'a�}AUBf�QF	�iW
H�	�'�.�Q@"\]T�����ȈP��d
�'�lc��_�`*�#V# ��	�'�
���C׆
f�2TR;j����'�E�rb��XUDKc�Z�i��e�'&�����
-?m*h��>]�0��'���*vXyy3�Y�0Ȏ�¥��<)�����Y��fk�H��'[A�<A%���7K�e �K�EÀ�c��<�e`u뚔9P䕐n`|�7�SD�<AbH�v^:�A7�&{."�h�}�<�'D� �8 (1E��{A���/C�<�G��d����ጟit�1��z�<�
Xd�ؤ� M��}a�ՈeXz�<y�K�T�WH޿)��D	��Kv�<A� F��d�
�:��� �.o�<�T����9�3	�(�ʵp�h�<� �݊���<7��YR�?���"O^�;u�5<�A��A�C-Z9�"O2�������^�`�"O��#u׏l�bݱdΔ��|�e"O�`�Ø$%��p��31�P
�"O&��'�ٮ:�����;q<��à"OV`��ȃ�����G��!"OX�f�Q���9�6��_��"Odi۶�Ƶц��t�֝f�Pq"O0�( ��!p*��iP6?~���B"O�����R�����	�eF���"O����l�:�y�FG�OO:`��"OBL�G��kG�`��Gޗ)9(RU"OJ�Xw�N'fB�9�L�4
v���"O���A�ɀ/a,@����9�2<6"O��uI_�9�0�2e%C��Hta3"O���C��_  T�Gk��`�2���"O& � *D/G&)rB�qJ��s�&D��a�ʧe����!B��aOB1�7E(D���ً��tSov6�ǯ$D�,�`��il���ϙ X]+�c/D�x-)ty��/�4Y}�����wI!�$ʒ`��!;�Ȁkv���h�4p�!�D��r���Έ��ͱ0�M�
�!��}�����"C�
�X�Z�C�-�!��8~�z���aܑ��|�F֙�!�dD#,h�p!�V�Q�V]�����!�9msx�k�Zc���T� !�DW0�����c�F���O�S�!򤛎7�����f�6Mn�q5�K�i[!���EϺ�#�e�1uW�B�U�(!�d�+Y����JNB*� f�(!�Di���TG@�h�&N�&�!�V:uT|�Za�W
%��"��!�EyM��o�{���R�Ď.W�!�$��)�
|�Ձ8�2T�DL�u�!�$�<�&�P��b��R�BB.�!�DS7+��c�*��%�E�Z�2�!�$�2�1JT�͹v�$����9!�d6y����9!��r��K!�M6�mq"T�s�,q��0.!���?.��ik̈́W�@�)��޶S@!��/m(�$�M�@I޸���:f!�d��/��B���A<�1����!��e�L�	�OTFJU�[�@�!�$H/i�6�s�L�X7|�	1NݍQ@!�>U�̺V�;>=(����*6!�ؒ��]�dk�]9�e�a�&!�$�+)�i
1�Z���V�V!�Y&i'0�hV#G%
n�5�4$׉=!��M%��H���{Zb��$ʀ}�!�$P�B �Ci��%Ex�Q��-	[!�dQ�y <yI�R#w1\if`O !���,-�� �s@�-#,&�"��	:�!�d��x9�ER).P[�/T1�!�]-7T(;�j��9^����/i�!��<����C�w*fL����&yp!��kv T����wv(�ԍݩsW!�J�<>�;%�T�,�媴�VGZ!��ef�2AG+�P��ỉE@!�d��<8b)� j�6Q���b6!��6��cO�^�r���,��v�!�dɡRD�9���%�v]�􈀸[�!���.1&D�� حR�pmb��܇=�!�� X���H�S��P'.;p�<x�"O�2'G�Qo�cs嚞D[�{p"O���Y��F@hS^�*�"O�����E�(��=8F���<�"OT�� U��)C�#�{唨pV"O����\�+���Bh�+=��}��"O��0.�N���JD����)�$"O�,�"H8+�	��	I2%���#"O��@��D�b z8�r)�7&*��S�"O��P�O7DY���qB\��0�C0"O�!Sk`����a�7��0��"Of�b#��.��8� S�'�=z�"OH8���H����n1h�1�"Ox�3�D� �:`g΢hV��"OY�އ+�歑��II�1�7"Ort���ޢk5��;��Ў3~0p�"O��֢U�=X�ȓ��� �y؆"O�L��N�=��#�����C"O�hy�)��%���G��$B(��"O�	gG�qf&�C`-��B�����"O�pS B�)h�U���X�3���G"Ov��$J�Eg�$��'}l�+�"OF�)�%ȞQ���2 ����g"OF�
�R�E��L�Џ�1l�D|��"O� 	E�y�Eʳ�$(�.��a"O��j֭Q�Ey�U���G9J��p[�"O�BD(M8s?�5�U�Ȼ.J��W"O>1�	�5��y)�(�
HS���"OL���6/Op�J@(ӍAr��"OƔs���p؎8�Sg�#�jUw"O��9e��]�$)r�4y�$��"O\=H�g�%BT&i�0oY�J��'"O ٷc�?Nsv�Pm߷3ȼ� "O�!��73�v�x5G�Y��"O��B�62�H��#�BGHIH�'�hܡ`��b`��-Q�Cv)
�'�|qP��Ĕ:+�D00�Їq�2�`�'�zE�C#˛J�E��+Gq�]c�'��1�C�*hH;q���|�[�'�v�J���N���Z�NĤ`;���'�X�u�M�N�P�A���f�b)�'�)M.B�00 c��<c�'ƠT����~sPk�Ѽ�~e��'O�d*U�u<�c-�$T(r�R�'�F,����;z+6��ɚu��]I�'(�$�a�Ũ1h�+�H�=i���k�'B��p�l� p$��(��iexջ�'�ư�v.���Ȭ��Øh�A	�'D�x���?jd���O�	�<��'w:48���+D����U��u��'A}Y(� �����H����0�'h� �m�9��4h�!�
�'Tf 8#�U�-���X���-����
�'JTd:V �9R$�Z� W�W�,K
�'�zP��#Ԯ���*�R��	�'Se ��E�,�!�c�:B2�!�'Yd�{���I��W*_55^p���'F������6"��@���#�=�	�'$-+T�N$4Z�颶�ձk`4��'��e�2K�b�� �\d�t�+�'�$���N�2���%�`2��'�6�P0�U:}7T�q'
;&��*�'dp���'�u��C� Y!�*��'�� �f�w������b��� �m��C]
�ic��n0L"OlЈ䮋�P�PH��A��8��p"O��¦��+����L�	��5 �"Oz�z���p��]z#�C�\���"ONT�&�<c4�]��C]�z"�!�D�=���1�եX�\(���!�Ċ�4��������!Ԧ�s�!�d�7=��%Qt&�d�1�D�2�!� %�>�K�\Q�.X�)˲j�!���Ua�JG(@X�5ɇc]S,!�B�\t�u���?B&a�C��Uq!���S���թ�� �mb�7iu!�䛄e��p+�>opɖ�ʊs!�$�@	�tHT�	�U�b�@��@]!���|��xY��=g `�j&�F>!!�䂵y�� �G�a��tqV�	&!�dڸr�LՆ]-~�ňD�x!�D�$0bF&C5L�:1{�iQ�!��4
f���GnՒ ���&�ʯb!�ė�zf�`7��q鲩J�J�V�!��I\�[���0W�R�*��Ƹ�!�$��L�� �7n `���:CS!�$��qDS ��,�fX���D	k5!�$X�:N4a�/I� �����Ɛ)3!�Ńh0lE�'�
E�*��f%M2@1!�$�;G�Q�:��LKd��<A!!���?L]���)�Ȝ�F�Q!�ċ>Km2��e��e�����N	~!򄂄i�^�p6J#.��dq�g߸ ��t��(�:\P�F���e	�*a���!"O�H�A�Wh��ДE�W@�т"O���A,ʝ���Y`��E
(�"Oj��oҋD��(�
TS)l��V"OQ����_��b�KI�	r"O�$��Tb���>Q��ڃ"O$�]�=�&�� �v�"`͂ b�)�'b$P�!@l�L���ǉ� I�$�'P�!戄:N�����).#@���'���/���b�I �����'��T3b�?YHn�)����,Z
�'`<��7c��t�`�P�/��Z�'Rz��g�����'B��4�I�'	��%�V�`�9+��$x�@B�'�:��C5+X�83�Ë{+�A�'�^���A6, ##�@�f3�]{�'�T p�AW�E�4�s2]����D4O>���٣f#t�	��I��"O�x�hI�O������E7
�"O<���cN�a�cе�`#�M!�dӓ @J��g��2P6���k�%�!�$sڠ1 �@�FN���+g�bO�X���Ld���S!߄a�:���"O��0������	k�J��^�dX��"O�(�%!f�$ԩ��l;�P�%"O��S��-�(`��`���"OL�� 0Nz�LSZ�8���<�y˘�iE��3T P��8�(�e^���d:�S�Ou(E2�:'�\d���A4V�)���xR��
;9�E�e玣x"�!KF6�yeZ���Ɋ�Hm�Te#���y��K@0	a�>e�6��w,���yB��A4ęw���l��j�ݻ�yR�ҖJ�YK!���vzͳ`Ǒ��yRڏ���� �c�(P�Ε����?Ɋ��� v�!�Q�r[�ԅ(,��%I4"O��@pE�N�,��&�R	i(�{F*O��2��2zr|���Q�߬���''������.[�1�SH�<��,z+O>���ǵo�X�Q�o��G�4� �Dٛ)�!��J�ɳ���uz�9����!�$�
r�=�TLX8cލ�F���3�R�'��O?ɡ��¾T�m����E
`���h�]�<!���s�(A:� �6h���m�2�yR�%/^d��q���.M"�'�"��O4"~�B��5̲���O�F1lm�uK�<�f���ubx�oH e`*�3q���y2�Y�ocV�3��o�4}A �y�c��;Lڬ"Ԫ0o5p�0Ņ��?���,ړ;������C�~Y�����\�j
�'�����D�u�B%�����
�'��0���
9$Z��[p͛�- ���'��Y�W&�"A�`*@'�z�\���'{���b<�98��M�H�a�'�$��sK։<��Y���$j~>��
�'ۂ����R9c�v}�u�+^���
�'��mF�Z�nJ�2I	�1��!�"O�L��`W&�ĠV
V:ieVx
�"ON�D�ҜI`��Ǘ�L<-��"O`tC���k�Ziൄ O-�M)"O���e�٧���z6�+g)�lB�"O�
��|�4�2�Z�8�Q"O����r ,����d�<�Q�"O~m�4KX���``��}�x	!�"O�[��5yF��7K-v��!�"O���Uǚx�)ٴ�D�(Ϻ�0a"O���`���9DH�UN�
W� �6"O�Y���'{h���D�<R��"O���dҫYd]z� �>@�Z"Oj�!�^�[l��-�f,؄36"O0x#�/�1cd���=j%ޡK�"O��Y��� ��2FdݍL����"O�@h#!R9"��-Hq�K�eQ�"O4�@A͠*P��S	H�����"Oz��Z�c8�m����-c����"O�y���b�v1� #v]�:$"O4,(2��	Y�����֬X�T��"O�1��)T�vpp��/�(D����"O��g挀#`U��Z�|8�D�"O �)G�_ Ev�]�K ����"O�*�M�x�b��j#`X:g"O�a��$&=�ȃT�Yg��̨�"O�P���Yg��,T�E�>q��"O�
�닒1?L�)�BC�̀P"O��%Gئ:�:Y�5c]�T0w"O�h����&^x�-��BU
AJ"OB�
GKT�;�d�%�� f/�G�<ѵ"V�X�� S�N�V�&I��+�~�<I�ɛ�b�^��a�A`��,b�
e�<��Y�:f��F�R/|>8�a��k�<i��$M\����O�p)����Q�<A�J/�@�`�<|'�i�/BO�<��'&D�|	tb�>>Q.%���U�<�$��K����%b04��a�Tl�<!`�������[�G���C3a_�<���B1
C����&�v(iR�^Y�<��c?B�q��F�0$�Y�<����@�4�b-Տ
�b��T��N�<!@�Q5[Zhɠ�N"	F`�v�U�<� �U�B�3B�z̩P��j)��{�"O��sJن|��EX5M��`$D�@�"O��a�/#~
D��]N�ʷ"ON�rvL�
Xpx6j� �"O�I�B�F�g�*(�'LN�"��"O���
!zyd��3�z\����V>m�sIߪ��H0��;iBr1A��2D�Ĺ��@�;���)6� ?5r���M1D��X��"��I�i��)�х-D���(4:��Z�#Y-��,�6J&D��Э�-���`�+D�l:�����#D�����@//!��oŨ:_4����"D�Ȉ�j.o|D�T�A,�d�%�.ړ�?��dV�B����&ک�<rF�	�(JB�I�!ؤ9a�J�w�.��̅�CV�C�ɌTPZ�{fFU�e0|��ߪ;�tC�(FЈ v@�!{��Y����t�
C�	��FEq�O�3Z̹���U��B�I�_����CCO���%�xSrB�I��|�ّ�)*�TMC5�;:Y^�?!����*(D%�e�Z�?�2�0,Se�!�$�'i��|HfZ{PT�B�ȸ=v!�$I��~hs�؎_^���G�!f!�Ā�X�	h���=U�١�]���e��(��ܠ"�Ʊr��E0eõ�t(�"O��B���o:I �$!��l��"O��Rnʯ�U';E��؀��'���4��Y��4�d͍*7�4��P�/D��H@b�&,�� A���T���#/D�p	��*"�xȐi�.w&}�,D� [��Ӫ@Xt���4�
%*G�>D�l�R�5��l��Y�v��؂�n7D�� �A�r�| �AY3R�8(f4D���Q���x"9�d�&MU� ���3D�(rb\�;)���S8K�D,�v�3D�`�P�J�06��O�0'>���/D����%̉8�`�;C���M#2pJe�.D��8#	
�#����4��L��� �,D�1�����[��^%z����)D�t���U�#�.��S��^�bY�B"'D�d���*#��0���9yT��'#D��HƊJ�#ʾ�HfPΒ�Ӷ@5D�,١�������-˯�.H
 d0D�@!0�*,.�� ��~d��Z�/D�ԣ�'��x�׬ܟ!���ע/T���'$=X�lB���R~�(�"O�U�@/F�pvj%� �=8N�(�"O0��E�,V$Pr�	�9U,�Uw"O�����M��f����C�_2�a"Ob=�n��9�"i@�	�;�TYg"Ob�M��?m�d
��;#� "O��4�-J��;W	T�g��� �"O�[�i��('�%�e�]7��"Oұ uGٌ+^�K#H[�3Ҫ�S�"O2��O�-1�x��c̣L��p"�|"�'�F��a���*LfPk��ÃP8ja���x�B�##� %(k��\�r�L�y��	��9+S��4��<0��ƾ�y��į@RE��O|O�+���y��4Y����%1p�ʉ��ޟ�y"R�`�����:d<:b0��'�y"�A�	b)AB�\14�@L��B=�y�Vze�X��8 2��-���!���'n�b$� ��	(Ā�i�1#��� $��R�]q�Hiu ''��"OA�'� 7�������(:�V\��"O�X�d͇"ӆ0�������|!�"O:��L-I��0��Et���"�"O&����M(Z���â�Tq�m��"O��b6ADZ����A�8Y��0��'f�ILi,)�B�V�Vg@պ���{fB�ɼ�\(e��:yT�@�Ġ-5PC�ɛ>�V|�J@%&f<��D�þS~DC�M+�-�W�:��#p��'@�B�0nAhmzfb_�,<�uR3�)�B�I�x2�a�1�W�|���PС�{˨��0?�a�O��N��ߪu���S��T�<�ć��.0� :GK�%K��R@�M�<�ÂB�~��0)W/^�XH��qU�I�<�2+�A	�O��Ct�i��H�<yEFF�x���sf�ŇJ<���b�G�<IwM���"�U?b��C�G�< )��>��`Z'ZD�nd�"�l�G�`����7�hIwA���p-y�'D��{�F�4i�`�$��I�l-2�%�D!�O���B̒&k��!��#�R30"O��ZvbPW�(�"���^�6��"ON�r3�F�e8���W"éE�����"O�y�Pf������9P䞑C�"Or�	DX�yb0�R�ȹM;
�*��|B�'_Lɠ6 �/�V��CX� �ݰ�'�r�Y�p�q�C���<���'g�l�Pe�=��a-�7���
�'fH��H�9`��(tj�.���X�'N
t��e�9t\|������
�'�B��Ʈ^Ț��)��6�+
�'ݬ�h��ɹ:��I�,�C�h�a(Of�=E���sZ��%�τ	�`���\��y�%K&C�(�y�L� 4�����<�y2�Ҏ#'��%��JX0O�5�B�.a������+(�ؤ�TĐ�N�@C䉌t��iq!�B"��C��l�LC䉠F=c���^��KʈF�C�)'`^`Q������G�EF�D�O �O��g�':p8��&�$|<�!l	)C2Ѩ�'r�R���qK����� �q��l��'s�Uk��$t�yt�zR4p{�'G�K��;G,Xt���T�'���'wR5�����1!���U&�i�'�f��PbȆQ=�\8�͊%�M�'s&!2����Y�^�۱L�-'x1����d�OF�S��{"Ђ)�dU�$,><(�� @�;�yB��f'F0?L�פˀ�y����jH��EM�)/}�y�v��=�y"�N9$َl�G�Y��	�n��y��w�R�(E*`���L͉�y�����҂��c����Ⱥ�y�i�:�J9��@Ǝ=�Zq�f���'�b�'���A��)��I�3cP�
�ɢ�'���u�X�.�4��gֲ7R�8��'�$՚��H�b!��E�'�v]�E�M������0�Z�'�zm)�M #S�[�%Q84� ��'Ŷ$� !R����B6���']�,yt�E�J����sl��7an���'i�\�TNľFzE�S��5�ft	/O���,Z���)wI�,T_����k��C�ɨ9�	���+h9�\���˓EҦB�)� �8P`�;;=���
�tHF+"Ob���Q�&�sdc�K*��J�"O,�8�=Xꅫ�"K`(>bq"OĕH1M�VDy㢠�,2#��^��D{��)��t|l���� �`ʢ�N�K�ў�������5,V:\�\�`�U��dC䉽�l$Iu�A���4� ��-�`C�	l��E�]��&�A,Q-�tB䉃[�:0٢IC�gD ���D;;�C䉪J�zeõ�
3k(�L�3;ҲC�I ��U ��T"�Wl
t0�C�I9S��I ��(E�0�ĜW:����q�P�'c.�8aGƲp�聁w�A!L���	*љ�" 4���a �uY�9�ȓW�Z��iՋmZ���@��(�ZQ��>e>�DhP=9��	b�(��9��n�2H2�C�A$���G�p�-�ȓJ��nI*3� `a��D-s&h��	@iJEۆ>P�Bē�|
���2�ɠ*�ƀ��MZ�2Q����zJ�B�I�9���!AQ/a��́��Xb��C�IC�N���$wp����O+�C�	�Zm � ��V�c>���$�߄\rB�I0� U
D/@!B}�i��Iû| NB�ɞkpNP3ɕk�J!�Q˅�*b�=I	�'d;޴CS+ַqDFp���#34�!�ȓ*�A�I��T�@�)��%Q&<��ȓs��]��S�K�֠�V�ݠGaH	��D#�Ar�
](�zd��V�q�TلȓD�TѸ�-��K%�%�&�	/\V���ȓk�x�C�K��˰�Y�� ��Q��l��I���պn�b���5o��5��NA��I��V�vڒm��E�<�jy�ȓaC.��G�s.Q�!F�#g(�ȓ}��i�bcJ�p� IG�Dm��U��xm�sa�-tٓ-�,9Ҝ��0��ܒ��:ܼy0���e��ȓM��j�C��lG~X�A�G!S<��}����'r��1�@��'S,X�ȓ��	�+Civ����#[3Fޒ���I͟��<����930�!*��`��b�<AV�S�T&����)�%g�D�c,�V�<�E]&��AA� �n������i�<��(�
*�Ԕpd��W�z�2�c�<م�����s�ʊV+d �roUF�<�'U=�4	�/�+�Z�����C�<	��_#:��K
_)	�v�z��B�<1H��0�{�O�E�Ԍ���c�<��T/iwx��3�]'GpȰB��\_�<Yw� PPN��׃W	^�Ґz��Q�<�pH�d$r�J�k���`��I�<Q�
?�&Qb1�S�W�Fm҇�k�<�A���LA��:=Z��B��m�<y��V8����2$7���3͛l�<����?����ɷ#�H,b��d�<Y�9�44��F�6����"l�b�<���1Z�Rb��*%��	�Ãd�<�A��E�`��I�(x���x�<�㡏�I^2���/j0�h���Z�<��-�r8��u�W$5� aF�Q�<i�F��Q�¨�6���S:T �6	�d�<Q4-�G��aia��/;��k�	H�<��S  TAa�#��XR
�3TK�}�<	�
F�{���=L~���D^�<� Ā�3��. h� w�Ѩc�Ұ[P"O�5�q��X���R�T����7"O|�7ES<NU \��ٱ۠�ss"O����

'\Ē�
G�) ��1"OH��-|�l�Z�(G�,-�1�"O���a�N�E�W�ג}��s�"Ov���D�uv i�@Π8.%"O��&ʢQF�!����t�d�P"O�tlֱb��u��YpK��y�,�.d�S��Z��������y���1j�$�`q�ͳ&��q ��
��yRa�0cL�I������P��ۈ�y�'�?o�@����վٰ�Z �y2�/`� �1akK�|4"�ؒf��y�m��r�v�!%'��m"�AJ�'�
�y�I'4&a�A]>SeZB�iT9�y�"�4��;S��BTv�y����y�ɜ?*�R�!���BeX�k����yf���� �ǝ:'��`��yү�B�QP���|�)��C�y�J��d��DÙs��9%���y2��I���0�҄i���2%�Q��y�+NB�d̢p9K�1
�S �y���+��l@�"�?ɂ0�QdǇ�y�aE�[�@X#��e����P���yҧI�M$e��ꂰXQ$�)��=�y¥�{Є��F�#Uk|B�'�*�y2��+
:�1���J)"�B���yÒ�<��}k�'K�G/��q��E��y��� ��ES C�\���\�y���%\�d0�@n��?v��be-�=�y��H\�ԯ�;��	V"�y��E1r�Ҍk'85^M��a���y�����f.�)�`�{3���yR��`�hi(ǧJ(x�l�.��y���q�x�#i~���"H��Y!��![wv����٧L�LEb5��#-!��;���+�FX/%��@2D��1:!�䉸�NPp�V�q�@��ܮr#!��ަ�N�"Ug�����jp�_�:!�d��.�ɠ0�b���tMO!�dQ<>8�IG��Gˊ�a��R!���f怄�sN��r���V�i�!�$�12�$pר�'9w��T�L�n�!��O7������;˴Y��ɪ(p!��1l�Z#Í<7U�����M�;m��џ��?E�aZ�'�b͘%bS�$�D�D%۬�yrEI#C�0肅�,Ed�"��œ�yߢ#p4� 4\8
�Y¤�5�yB��R�<��K�+�+b��O1�C�I98�ŒC��%r��#��]-g|�C�Ut�l� !�bq���޾��C�� �l�f$ �)RQ�\+b�C�I2�L-D�ܷ-��HI G�(	j�C��}����nC+A���t��O4*C�I�����Ώ�d��B��)8u\B�I�Z�ڸcv�
�Dmҷ#�^	6B�I�n�@�@7�#s8m�t#?��C䉞aFUX!	�i�L]���N�"��d�O��&�O�苦��VpB�眸m"a��"O�J���]�X�6�;}iƀ�"O�<;���L+ ��$+	HX�8��"O��rdl`W��	rM��Tɮ݅ȓl�d(b���-�ƨ!
v��T��S�? &ܩ�FS�G�T����?��ȡ"O��ct �F�S��L�f�g�'t�	C����L�H ��x�# �vM�H˰2D�|�怐j3��K�ΞD�h%2�O��NM�p:�o&8\a�-H�I���ȓc���#B/S� ���� Y�H=X��ȓ g2лt�ʥz�R�X�Ҏ_\��y��k@�X�
��t�g�G�%!6l��b�f���蕅M#d�1F���dz
��'���'��M�f�܅b4W�}>x���'}4)S��^W� ���(s�$�*	�'�ơ���;$,�Y�R1h1(�8�'�ztˬ84�G�C#f�t�'���ᓯT�'K���,Wl<��p�' ��%%ߟu ,l�&�Q�6�	�'�.A˵I�-3�h��Ȇ2�و�'�1��/O�8 ��T�ɑ%&��Q���?Olq2�8Ut%�R�-I��Z�"O6dѦm�� ���@�3i�S"O@����N���T��uT�`"O��iÔa��U�u�ߺG#R ��"Od�A��S�*pAE�rĂ�"O$hsE�1a{^�w��78��4
�"O�9�e�1J9y���e���x��'Jў"~�O�~�|���
�l��L?�y���-7��:�'2vq*+���y���A])�S.� @vܘ��M�&�y��o�Ε�D��n������yr-�*	�e����a�`!i�f�yR	�"��ђᄒ:n>�p�.I7�yRcN��p���iZ��r�N���)�S�O_МB\*r�j�㵬CLc܌c�'���(WML�#�� H6�ۇ=���'���Bc�^0b���f�~�Z���'�n]��y��<X��%�J�Q�'9�d��M��S |��4"�%�n0��'1�dcbZHq���ސx0��'����̘�)R\E�	�(	^|����?���i�60I$,�"LB&;��B̃�f�C��$9A�������-��\�i<j�C�	�s%4����pk�|�� JjC�	+X�bY��L�<U�����W�&9@C�I�{(�)� P��\ңL��4�C��w`�v`�'iv�PQqE�[4�=��'@��hADٝ��n�O�N��IU��Py��� %�@|م�'7T����0u��B�I.5C�+�7V����Y�s3z�O�����ZHr���!{���"O�=!!�Dп}�*	 p'� ��ȵ�B�H!�$X�� ��n�L����*Z!��HX������FPx�ƶK!�D�N���4l�'D��v�[�4��'&�f��~h�cCh�� �a��0b����Of#~��@�/A��I�G�ɋz�.�se�{�<�����'�"l�bھe%�Ы�y�<����\4`kA.�<���y���~�<�'�p�JPzf��'��\��-H|�<��`��i��B'8"�erF �b�<�e�s_*�M�9����`�<�mٰu�xpr�֑\�}��F�<�wi�3\Z��X�Ɗrr@��'J�I�<���>&٠���Kщ���b-Q�'ha����D�!��N�:��  �]��y"a�t$Z�ƌC�8�,԰�i��y
� ���2@U�	�hD����>c,Af"O�}h��
3 �L���eK<(U����"O�A+����O4��
�"WOJLi&��v�	O��A5*����M�/��Ih1�F�y�@)2�S�]~Tq���&�y��B:C��!�K�<�*F���y���'�� ��µ�R:��;�y��1���S L�|^�!�c���yR�[+0�$LcU#��c���5�y��,����lA*X����Q(�y�̝�l��U�шQ�9\r-Qq����y2k�'A���vfې5+&���g�y2�K��Yq��*�t����,�y�f\,
*k�'�
���%ؔ�y"�;k��!VK�o�b��G�ÿ�yR����	3�b��oq:At�]>��=A��?ɚ'�&�`W_i[���v���5Cܨ�'uP�C&.�I�H�犋&1;0�h�'��'cAK����F(.�.�
�'Pz�$�Űj�`�3��P�����'��D�f�/3�~�1�ۖD����'�lɛ����
��5%3D�r��
�'v��j�kT1ss*�ŮVH�ƕ`	����v�����
'�琴h�*�� �8D���T�O�k|�	�F���`��f`6D�ģ��M� Z���ױ`v�4L)D���f���] ϙ�|�n����%D�HP�b�ƕham���b�X`�-D���ď-9ʲ!3��9�R\k�6D������#)��P�%� a����WD:�In�'%�4O&H�ǟ/g�p�"3Y5��"O&�y���(ks��2F�
s:H���|B�)��"J�H�`C[1V��LХ�S<C�	j�F��RȈ�m�쬩�K:~1JB�	1
��\�����!�
�z���x�B䉫$�U(g� �[��U�r$��'� B��+�N 
3c�Y���)D�46��C�ɓL��]#�k�7p���4�
�=�ԓO��=�}�țk�<��f������Ɓ�s�<a�dY�%��сB�Y��ĚcZW�<� ,��t4 )��R�T��DRS�<��$�/v� �U̒wǶ�A獗M�<�Ł10��Pt��B��	�J�L�<���J:.8~��5@PW�h��`L�<����
�ڭr���'!^,QP��Ky�)ʧ3k�xSN�DY���}�h��00"EkR��,��Q�ċ�9R1�ȓ*�2<!0�Н1VP5)��B�-QE��6w�:�Ő�b���x �� �K4D�ۣ����+�#pV2��c�<D����߰x�J��7C�4u8��6D��5�d��c)Q.�EÃ�6D� ����:J�<�R�
�a������9D�L��=bM�@�'[�N\�4D����m_�-�$����,I��N.D�@���Rܤ��cC�V�(X��1D��P�o�%�5q��?*��u�0D��
4��1?.�&ٍG�p���&:D��i�i�cD�����N�J@"��;D��PQl�'xL�Gl[T�:����+D�H� D�?�,�k��ۑ5���T�*D��Q%�	.E��Q�W��;��ղ�A#D�Б�$H&v>� !��W��+EI,D��Ñ� ;Hxf�zR�� �t�"G�(D�� j@뵡߼~g$��!��$ 2��b"O\�Gɖ޼�sP��9�0�$"OC"�'b��K��T	���g"O�L�T	ĔBE�H`+��|"<�2"O�m����63,d(r)�n�,H� "O�ps ��G^J�hP��; t9��"O^��g%͸ ͤ���h�8cSV�)�"O����Z�R0ȣ���$��`ag"O`m���) �P�&�E${\x6"O��"f�� ��!3X>Ax��"O�I�4m��3�ӌD�ڔ�"O��� ��J2D�2)IE�<��"O�U�4�	����۱�Hـ7"OT��en�>=�N�;F_�Z�<�Y�"O���Ń&ZFn]���q�6���"O8�Ƀ��e��#a��[����"O.m1����g;�]C����|�{C"O�K��H�����S-O���Pr"O���)�:m��Ms�`�\�����"O&Q�/�8��@Y⮚�B�Z�YS"OZ�����g�q#�6z����"Ol0s��[S�8��,>'�|L`�"O��{gH66n��4�:\�(�A�"O~`rq�'!�̨Z��S�]�U�r"Oh�a싊HJpA�"�Dn�L��"O�+��K3MOPhQG�g��"O���A�q����f@XМ�v"O��SO�/|ސ�4��\�l%��"O�YUa�2g�Z� #K��&U��"OHL RB���R����g���q"O���T�)g���2�)�_��)�"O|%1 �3�L�h���~�����"O��yb۔B�>��lN��|aV"O4���Φ�|�x�j�j簔�G"O�h��J�g�<�����|��"O��P�o��[�8��H [�A"O��3�'J%?��8�5��1f]�Xqa"O���&ժ'�p@�C�/z~p�'"OzI�`�MZ�Y3P�@�#z�]�
�'�6pq7%� Bt�l����;���'�2��kT?��
WK۟;Q��'�����'�	~�6:��Z�A��� �'�43pd��d��<��-�N�Mi�'�੢�C�6>HXQ�ȷo�t@�
�'��,)�@1L'��PE��:g4*�P�'��uh�U#!iB0����z��'�!ץ����@c⁥a*����'� l��(H6{Ӽ��"m�7%�|���'l��@"#P4A��,B��jD�UZ�'i��T�ҝo�`���*��N,еi�':D�z4��H�C�W��5;�'>��P3b
o�L�AgO>^�%(
�'�)�p#�_�"��PfzE �V)(D����ٓTR�����f}c��&D�\�HH���p����6@� �p�%1D����GN�L$���p�Y�ڙQ0D���QiA4}�@�� _p�ٛ�l:D����K�&r~�hPr��.
���k-D����jݗ��Iq��{4�A���+D�H����dC2��ԋ(+�BІ?D��)(b�����R�
����"=D�`�	_73��yG9c������9D�d)�%�&0 B�"k�z�d���9D��إE�;�p��p�W#g�6�H��7D�� ������� �H��i��S�x5Y�"O�QG/ȸj��g(F���@W"OJ�r�ǔ �8L(J'c갺E"O��qCKD)��8!���Ia2��"O��R���[���$��#cT@hb"O�(���yD�ѡU(R��R"OR�7k��C���s��Ī\�)!"O"1�tE���"$�E�f&��!"O&<�¬�->���$H=[���"O����%!>b�(��v(���'w숈 ��	h~��7��E���'�nm"�	iy��:���(3<�)z�'������_�B*��h�lUY�M���yrb�+#D>ɢ��.
(��B�C��yǇ �z ��A�~bz���^4�yB ��U��	A��>Z D�dX �y��Jb�I��hŌm�ƙ9�O�<�yE�ߪ��@�ݠuz. �K� �y2�������	�Y�ͣbl��y�3�J�㔧��H��ay3Aˈ�y����4�����@L1� ��y�] R|8�F�65ƤH��M��y�oʻv�V� �d�<)D S� ɫ�y���RW������'��Ҵ�7�yR���M޾���*�������y�n)R,�ݱ��M$m���m��y�*��m�"��?	�2���ɛ�y��J,� z�$�)rb�j�"�y�/�^
��@�шh�n(r@@��ybn(�`��R�	�ru� ���yr+ҪJ�<�;i�&~�*�r�M���yR���3���qf�y2 uei#�y���,�0��g�	�z'���Q�y��8)��!�#!|�j�ߕ�y�E2����A��\qr֬���yrϜ�MOF]ɦ*Ƞ��6��y�_�%�<�E���*, ȕ�!�y��ڢqv S���}�
`t���y��=3a,q��O�D��Y3o�:�y�茝f�~� @�=JHx�d��yr� s�2��ԏI�	�(�wE��yңQ
	��st��
2�K��3�y"�8װи!��6i�/�y�ՄXP�ǅ�8wA04�D�2�y��/�F{��ֿt p!��-���y��r��\�Eဨ:e i`�4�y"l�%PBڙ"&!�';BSӊ��yRC�.� %�@%�0.� ��L��y��	% i�1�Q��F�y��I�ک�Ǣˋ&JHyR�y��Q�i_�A%F�u�4��l�y"�7~�l�Q���1�`�K-�y��2j���@�:r���w͏�y��?;�*�ʰɂ2r(lBkH�y���|����\=b��*��^�y2'�v�!�E�go�t�3#S�yb�����I�F�n�	����y��\���u�׫j� q�����yB�F�M�|�(N5jV�p���y��A�'�,�i���1T"je<C�I�/<x#E�]�=j��߸E��B�n�q�3O  6PSwS�B�	�@��A�Ď�6	��p��#[#B�I)lC���ŝO�M�振C\B�)� 4�;C�G�O �ySA�1l.�d�q"O��+��F�/=�Ț��.E<%"Ox�#�ܻWK�%CPĀ�c�	��"O����ʀ[�~dHd�����y
"O�i� �{止� �2s����"O�	둆ʖ�{%jμP��"O�谳j�<Y��)A)����"On�"!b�\����ƈ9��])�"O^R	.�HS �ŀ{5���f"OԜ��D��bP�Ϗ	w����"O�xp�]:@�͐�o!G:qj�"O�S����P�^��h�>x�\���"O�B3��H�xg��pYb��D"OT�@P���)nv$zT&� .J��7"O$0�1aQ�X�e�q=� ��"O �W��G�r12WgɹT��q"O�=�s�Q3���P&�*/� �"ODA�^�@������:�5�+B��y��\ V@��B����$柤�y2�D5f�zb��^����W�a�!��gG��6��xv�y�lR�E�!�D�+>�j���"GF�D�^7�!��Fz��wC�8b/����ʹ0!�$��(�I{U%e�q���T�?s!��t�0�PF�l\�{�hL�mq!�$��\E���Th���PeH�(!���yۨ�@tI����1�){!�Dˀtz����_�D�N01�m֮<h!򤝋0�Hy����9~c���U+Q/99!�D�3l ��2�R4D�i��M�u!��$&3z1��ǺT��R��3�!�$
�@.�x ��c\������!�d�n��Y1�K�xl�p��GO�!�C8d�(�[6�	&UW
հΔ��!�$\��� �CF8r"��i�K]z�!�["��qʃ��"(A�+����'F|;Iֈ:x� �^'a�6͙�'A��p���l�`P�DOͽ['�!��'�&��Q�o��d)���[H���'B�
�"��\'�lb�hٖS�j��'QNhqfW><�D8@�LSF�:=�M��m�W���0���z�;��
y��<�vc5�OP�n��1'ꅛ��x!#ςC��)r��d?�>��	ڂmx��cH�:e�J���d�b �O��N=?)c׍޵0p��%☄�`$x����4�=����O�20��6E��0�Qur� q�"�S��yr���6�7��rlh����y�aGw�"lsp�ԍ �r�k҄�	�y��ԛw=|(��$�mSh��iR��y�aI
�3$e�c4��#��D�y�
N�V4����Mړg,����՘޸'�ў��`k�	�,M����!k�S���:�"OD�� ���l���vI:V�&Ty�"OP�!�-$1�O�1-@���1�S��y��,_i�1�͵Ea���S��y�k�0�����.��)xg��y�@F���+�-9�yr��y��?](pu�7���'?`��E.Z-�HO<�=�O��y+vď�8h>�����7=Wv��	�'W�Y
'.
�BM"� :@�d]�	�'�����*�Y8��ӾdƬ�	�'<x�p���.;G�h�Al	ZP�Q�	��~��/3�I�vDJ?�P��$���y�`آ'kx	�ጟu9u���ך���hOq�� �)-ןԸ,AǊ� k��p"O��bG)�+( �hp���
@~� ��"O5sv�S/ad��qŐ|F`j��|B�'1�t:���<�4z�/�ʞ|I��$,OL0Ƌ�Id]��kO]4PY"Op%q�E�}�d}#���3�~��"OD�Re�	���s�iI0�B�x3R�tn�q���O�~��6ˊ$�������Y�j�'>4�V�s<��H�)UZ* �'�a�&w�:-��c�,W�ѩc)ݚ�y�,�+:]�dܿ"��&��y���l�B.X6����P-�y��"�����e�$���K�����yr��1~m ��m/����)J�M{M<鄧�>%?�O�Lcƿy�Ȕ��.�<��쀳
OT7���p��ubƥ�"1���Ɔ�i�qO�=%?	쏱!�p��DŘ-��02@/"�?�j"}���aV��4���Hu�R�Qz�<Qu���m��0H��DX4��3��y�I�A�Q���yҬ�1'����˺k�A+g����?yp���x�j��J&��г ғ:��!ʅ	>��M?�O>i+O��Bq��sd	�CI\09��#?с�0�u���o ��Dk�am*��&���M��'b�	a!�!��)E �hV<����O�b����$"�*��NqP�-Y��"ĤO����Q�a7Ѐ���,9��8r�����!�Řp�T��e��?v���bT�$�!��Vv��%�a$�{��HV���џ�F���͡�.i1��X�<d��1E����<aM>E���>P��1�B��A���C!C8�y��S5[om�"�reh� �B����-��Z~r-\�T�[җd/yM������8z�'-a|�n��Z[h)�7�S���1 �K��HO��=�Oޖ��w� .ol���i�oY4uh�'{Z�3���@ �� ��(I���7�S���)�x@H�Mv!���yb�&�|`i/�p^�P�1M�>ˡ��:j��&̇`&��13��2z�$)ғAU�&�D�=x�L��o�UL*���B-�'a|��J8�ra��?��ڐ甆��	Z���O�$yZ�+ǠA� !C!	!=�ĩ����'H�<b��pg�ɂ@�5<*���'�@�o؊�F��7��8�9�
�'8M���<�4L�P���
��y�� }�@���� �5��o6ў"~�%T6Dz# 
�^~�g˓&�t���H�-��kV`�ț�.�$�~e̓��?Q�ix��Q���HWz�7O�YB�I��Th�(U(e��X0���&k�BB�ɱv������]p+�	Wd��{��'�S�t�����O?�Z@�f&�	p�C�I�vl.�C�)Щ }���A�0ܠ#=�Ǔi�h}i�đ+_X� +Ҽt�ؘ �'�*Р��1�4�Bsi��j�Q�'�h�2Ǉ�,w��t�'NRq\Xb�'�NE���[V���'�!gG���	�'AШ`��D�Qj�7�}�a�(O�=E���1/�pؔ#F$e�p*T��y�ɺy�����ӇRmp%ɰ����'7ў�O��=��Tb⠨�n�v��8���yB�*�� rK�����DD��y���"��xBg�?b��C�Q���O��~j��՜����&��z^%p�Ok�<94.�(}�	��O=$����jy��)�g�? ���,�^�8�8�k]r6��s"Oؼ0�b��rr�J��uꤓ�"OV%�eOJ�Vd;��:@�(2�:,OE��X,{ʒe㇀&���5�q���'�<сm��<��R0��­ِ�'m�>@���m�: T�{����@���Ӏ��'N&���N9eʐ����@�����D'��>��݉ *C/8��0�a.��6��$�',b�)��	�l�2(@���l┬˝^X��� �	�W$fyk	����x�W��%�P����'x�A�.�&%����+C�D!)�'r�5�v�ͨ!����. c��D�ɦC��D����å���E��Y���~��OT� k��5��ɒ��osp�9�/�$t�5� �'�'m��*BF�=`�HY�&���-�8YT�b�@m�3z��OԒO)�� � :b��3��=��"OT�Y�E\�dPT�&ͯ�Y��74�P�3G^73����� ��R�M)��TӦ�ow?�*O?�I5}�a�/n��!�7#��	d�B�	fX�\caL�ꐋ���8I���~r�)�3����wœ>)
��U/�G�`��$�>���K
38���ҤG)YG�r�� �1�O���$��vb�2%��%�e�$�"w�!�7�(#`ϕ?ʹ;$�Ŵh�!��i�<۲�T�j�g�7!�D�
Zzu�BG�,ѼP!p(U8!��	�P9��Ƈ�(yc��6e�!�$�&G,�w��<y��x��� 7�!�E��D�r���`M�i����(|�!���$1y,�Z4EJ�T�O�]�!��(U�hz��� #�2Y)AoN1!��M�_L��`�CM1)���!�d��	��UZ��׺5Q��O��J�!�$��B0�1�$&1��B¨��$�!��0�HM�'C͐o����e�/�!�$�)I�d��,��u��M�E瀽!�dQ���2#h �b���	e�R�w�!���h'�L��;!�6!I�%čGI!���<H�݉��W�`�J�k�iȏ3C!�0>ND�8.:U;�i��<U!�B�'�$`+�n[�d��fնp.!�j��Q�g��]�s2�V!}1!�S�(y�e���46�xM��d��%$!�$
65�b {T#��	z����j�:7�!�J/C�B�y�$��3e e!ƮI� E!�$�!$݁C Î^L�X��Iq!��&"� ��C��$����	E�!���	а
��s�BT0b$O�!�$�4J���I2��!&�@ �Q=S�!�\fy�D1�ۊ,���"��!0!�D�Vx1Zp�31(|ܚw-�!�ޑ*�L�@DdC/)���!�ސU�<}��Y�����L%;�!����,���)���رfEk>!�DH�
QDaA֊Q�n,��gB�h7!�dN0k:��d��n<ɘR�^:C�!�D��f�8l���a`�������gja~2��2m*3���[5F1-m�V�h��4^pU���e�A�<���X2	Z����z,�%�r��) t��H_{�)��s�>����ҡ�"5�CϘj�E��dQ:Њ����R!ADo�,�8̆ȓ9�*���l�%1 =ᄊ�_��C��L���=[�Z��o�?��a��S�? @���dхp>^1��,�8V���T"O�+�KK�K4t�h@j��x�P�q"Oʨ�qN�$TwR���KϚr���9�"O�A��C�9N4�J�+��5�v"Opqʠ*ԛ5D�q ����.A�"Ot���,������9��@c�"O��1 �Θ�eȂ�w����G"O4�2&��) zL��h�w��bA"OX�HF\�E�Qza%Ž\y�pZ�"O�f��}׎I��$�	q�$)t"O��`�@N�#�0Jb$�4]���"O����. ��E1�d۶l<�p��"O8��g�!�N��pE�52�di�'�v��!ẻ&2cC�nv���'���ش@�&��0���%-�h�S
�'�r�R����##_�?pH��'V
]��ß�7Į�rI�8,��a1�'�H��L�ULzM6�Kq\��	�'�<QH%Q.�4@�@r��*�'{��Z�,@%B���	�Ӆx��b�'C�P�+\#'^���ݔp�u��'.N�{eS��᧩	 %����'��hw�F'h쬳eh���a�'�|�sFK��	�$A�+g�\��'/�a��`KT�����!�[c� k�'���s���?.mʀ�\�H�n���'�ْV,Ϩ&�� �4��(M%HU�'W4Es��]�|t4q�d�<X@M�'d|=�mM:{�(�J�H�$ժ���'�8��ʗel�������.�!��'�PS'�P���K��9Lt��'��P�ï��dR 0�0���j�ش��'��I���kaZ��Gʀ�\�L)�
�'ތd�K������I�6H�N���'��i�A��Ih)����C���C�'nR���A^S;��wR�G���:
�'����$'��������ܸ	�'?�ՓfB�3M~�b����:j��	�'���JGfU%_��ŻS�:G���
�'�pR�_,@_`��C���l��	�'*������6I|�Y�j�C��I�'��!!΃F��ay�җv�]�'��]��k��%��j oTb*$��'X�YUl*�v��_�ԞB�'�䩂N�u���{%-�'
����'�*���A�q2��T�%��``�'{e"�|��#�Q,
�h�!�'H��ů��lϼ���A�3�n��'�8I��c�MY�!�g$�'7v��H
�'��q���i�}#.�{���y2��F�0�@o����(5��y�.˙1�����P=��Y��A֚�y�L_i<��PǦ�	�D@�uk�yB��\�\D@�̟p�i��#��yB��gAyqB�6"7���7���y�@ͧ��u�`�#-��xD$ʔ�y҂ʂ\:X Fj͐��1r�أ�y���oTp�1�aR�?��a@��ξ�y��-	���lB�X�t��ԥ� �yB#O#���EI)Ur��4f��y�K��
���=H8��a����yG��0�65@d�6H�4 K��!�yD��RB� ޗH���$��y�<0��kA��0ހ���
=�y
� �0s )E�z��T ��G�l�BdK��'�P`�w(
EX�`��Ŗ.	�Ja��u�X)˧�/��[� :�-�<�{�l��?�%�Oa�*D���=��:�� 3��� �'��e&	Ε7e��2D)/����O��	�Fְj"Lu!u�O�A� ���1i`�N~��Nd�tx��M�P�l��C�W�<�$��L�(�.�|�@�]*O'$����Op��@�RA�	�б��ҕ����	3{�F	�d̝S�@�0f�>=����O8s��mJe�Ca0�:�ka���F/�)m�0�!&��-P�:�QP��n������	8	�t� 2�ێs#�y���E7���X��1q��X��I��JԳ@+� iv#[�c7���l�/�=�࢚�n�" h�#>��?� -�@��X���^&�h��Ɋ�� kL�8A�U��i,K�����N�B��L�$'���$e�탲OP:Rq�rH��n Ѱ��9D��6@E�7���[�N!sN�8in
H�s�'�0��'P�T���>4���sA`�#yV�t��V��84 ��Ɗ�Q�l��'����B%�0�Jq
�)����R (ā�p(���
	M��eɈ� �Z,`0*��[\���ϓ�:\���H+i�Ty��È�P�v��'D\Yۅ�i>�X����0H҂$��j�@U�ɂV�b�p/%f<@Њ�GM=~� SGFSM�q�C��	ya�	
.k���؄K}��'�S#d����FJˎL�*����H�{."
Vi�,o�����'��'���yw	��1�C2AΙq��IG@ٓ�p?I��'y�HBa ,������)I��¯���x��N�.n��2�$ڑ-�>IR1�*����V�@�M��b�s��pv��6��$h��H�jAY�0�e��Q���@;N����D��&8
�X6>6��!�$��ڸ��P,^
���� \M
չ0�J .$ ��B�?2��#>�E��%V0e�vFR�`֔e �@r?��i�6���������
	L�(�<a���2m�*�0 �'���k�O�EߎX*q"��&J(��W�p�,8a��(�O��r��D�~]����n��GZ�E�D|���ևN���ဠ�L��"t�ŗ
�je�D�?Y��wW�I�eb ���A�%��s����Y����T�VC�U$I���S`͑�8��ކG܎��!�<��ٱ�OB�]��
����M��󄊝\b���!�Vq�$Zj�,y�qO�(�6�iݍ�U��-zfA8�:*	� "aÙp�t*�`[F��2@� w(�Yg�Φ&�ԕA���{�'G�i&,1-ռ���@9΄q�fܓb̬�3g-�Y�&�ݎO $�I�FM�&�>�6,=9ߎ�Г�I~�)�l��lČ̣���J���`��&�ܴQ �A8a�1�P��U�c��� �
�#��"`D�ɑ2&�ؤypKA9`�!��hVHɰ@�,�󕈎(Q�jH��I!n��r�>��c��*��u�U2X�.��j� [9�L��_Z'T=��I��wP>��%��[�"���Z��3�)Y(N�r���#�~�;�!�	��h���4���� �8LV}R���!۠m��V���A�ŕ&G:�����'<�&h�c�P�%�Z1���2�!$/@�6L5��d;�*.X֎�����OZ AQ
��5V/١���੝�C��K���y����J��򣊣1�r����#����tn<�O��Yc�'A�Q3��!M`r�k�"O1bwk�7_��`�֟9���P"O�`��.�7t���t��iu�E#&"O�=��a�� ��8p�g�$|er���"O"�ZpDߙ+��|�4��\RM�"O~܈�Nۤ 48]���J#co0�3"Or0jD�Z���x`� (:!�W"O$��Dm9e�X�W�b����v"O�4�B���p��yD�;A�|A�0"O��qWbS�*n�9���c��2P"On9[��̡^^��aUG�;|���;d"O�:�V7I3"�aE��5�p1"OB�Ռ�[}l�[�ş�F�0"O���rBGt�����Y�?�0��e"O�x ��5^5�@%����,�H"O��� ��eӶ,��j�1_'��2�"O�5�#�2��\�"�[�$ =𓑟ԩ�R�H�z�е��A��[�Mb��
�eT3��>���)UC��ֈ9 T:E��HA����� ��y��B)@x���.E?W0F�B
��HO*��AT�#�D�[���@K�>�θ���]On�������y�	�%L�xё,�:F�6�0��K�M��i*0�b��>}���iofى4�E�<��y�c��^��4��'�F���,xT�9�͙������O�ԛ�LHjĂ�@ϓC`�e�Ս��t�Е��P�$
f$��I!dN �0�H�9�� T��G�LF���2���#Jμl�"
54�DI6�G3]�9�C��QY8%s4�4ғp��{#,H���?5���H*8ؙ�j�	sHH0R�'D�1gb�	b&:4HtmƬzDd�xe,e�H���Ņ��݈M��}:G"�O��R6��)B�uc��n��P��n;�|�sh��g`4���X;6��3 ��>	��ϖ[�ԩ���<9ԬL'<^f	[O>V�ѳG�l�HBc��"���W�qx��K�c9�1eV�xRv�[҇M�DVh�`�ChyB.	5�E�5K��)Jԛ*T�<���ha(�:J�">)�I�{�B�|*�j��␉��d|�&�՟��j�4��O���gܓ�P2!�
z�hb�݊)X@1����h'��"�JH#��"�z��慌p~�b�'m��z���X��Y[��yir�����1�QՀڂ|�����@�y�S�]!sC�
�!��xqg�+A#DB��&f� �"HN�@?�S��V,dB��R�/���1T��?c`�1�"�g?٤���0��8��/��A� գq.G�<�5 O�`;fmB3�N	&����	B=Z�,!փ�7��@�5�0̯{�'� �Sb��v�X�j�!ȋ?�H�X)8$)Q����M1���
�ڽ����7�C�@7i�@@�[؟�� ң:� �b���8Ӡ@1��-�I�*W���S�J��+�+J��OC��L�]{I���*8as�'�5+�<�x0�F�"8~��g.Z0%'D��S�W Rh� �۴0��>�zF�-q�ѫ/�8��L�7�\؇�_�L1��G]�(��=B� ڙI�|o�Dꘋ�E�0EJ�{�{�\�Th];#�(���J���=y'd\ _�p�e�OXd�J�����d��^3���"Ob�(e�I�wO�Y��"ɡ�dCt晰���h��I22��<Be��'���:H��"OƘ(�ȅ�Q�]0���B/&I�'�0�Vx%�|������%ZȪ�e�פJ0:�n,D�xK��J3e�>i����q�څ��y�0C���O�|�^�(��l6&��`��Ǟ(�yD�7����܅؀mr�Ȓ�yr��(�
���δ��i򤟉�y�^Ux�Y�ԢN�����@�E��y��M�������~8�J�'�3�y�����w��P8�7ț(�y2)Гl�q��7�����c2�y"�D9HD�Ҷj��0��t�S��y�!S�<�H E�Bv�*̂#�y�o�i䖱�����4�*��R��y��\:2�0P�@!�SC�͈�ybMO?��4+�A'X�{�i��y�
Z��>��K�4(90q��e�y�'\��y1�/��'���҃�:�y��ή�f�ӵ���V�@�Ŗ��yH�D�L����F��Ω�AgȌ�y ��"��Xc 
_P푃�N��y��hR�� ��4$ b���yr�X�Q2�
��J��l߇�y�hC$�+�m��K��0��yBHTsf ���Eب�d���y�3I���g	Y�Ƞ�Z�U��y����u�:� �kĦ	$��(�m��y2�� tڡpqʆ���T��yB��~��[�,J�)=�=X� ƻ�yr�
O+`}S�A��]�p4��G)�yBoK�a��r&n
�W:^�f%�yb��@��(��լO�ʠ"���yrL��Qk�EǪS�z�y���y��*+��z$MăkN��e���y�\ ���+��Q4�
�1���y���"p�:�����}%���F�Ȱ�y���E�tU�$N4iqĂ�b�1�y
� "Ax֦"K�85���W	z�T��"Ol�Q�C�P�hB��6$2�S"O�)�f�̕������țzN�T"O��ĮN:NЭʢnی��[�"O���	�7MH��1*�6��d�"O��)��ޗMIRH�	
$>�Z�R"O���F�t�ĨvG��"2���"O���/E��l�G g�L��"OV�x3���Q��u'�Lc8|��"OD�H2ə0d��H7�PA�Lx�'�8�k�g MJXx@@����	
�'�hqP�Nǅ@	��"l_��4��	�'D�!2�"���"X3$3
���'1�5k�o�V�ܸ��L֬Kv4)�'��]4@��2@Lp�'�(:����'a�H[d� ��Lȃ�;�
L��'����'Z/�!2K���PK�'RX��/�3_�U����#��9�	�'�����F҅&��i�C�+g�Ւ�'N�<
!��Ѐ�&�� ����'Y��!󨖥N/Pi�&��^����'��xU�Vy�h�F�ra����y®�>���҆�+e���b�gϗ�y��߹��0��%���`���2�ybI_�
,��)@�DU�fx���*�y¨��'�&��p�@O�|��ab��y� �(� �D̳1Qv]��IU�y��.?|�]s����6���9EO��y�%ާYe\Y��O�{��� �f���y� 5��@�㨃q2�@���)�y"�8p.X2%�i�z��5�#�y�A��2� �pHP���֫��y� �Wc��R�p����ŷ�yr`�_��T;�/�i٨l��FJ�Py��J
qצI��*u�'"OV�<�Ӯ�:82�
�,߄"��4va�S�<��Cר�J����)+�Z�pďDK�<AƮ��|�"�"�[�!�� �U/�D�<�gŉ>!X|��A��*jw�A�#o@�<!`���� jI�dJ0 Ðl[�<)d&kI6�f�Yz�gc�_�<qE���/�<M[���D;y��&�W�<�#�	;^�a��)�0e� ��1�P�<��ɏD��yWeZ�:�IT�H�<YU-Y�4��a랭@��4����G�<)'�+l1��)�FA�v��5a�LC�<)"��e!	[U�?x��-@�C�<�tJ<�l9�F�C�MdB��D+t�<�F ����$J�@��<�3Kt�<�@�:_��@��-k|�I�e�Mz�<��Ϟ8�FIB� [�I�]m�<G*E�)���0�ιG�8b��@�<� � '�` .�#Y�켘�T�<���_�P���UHL��h�i�<��L�^4������� MQb�h�<�@
�W�X�;�cT=C�|a��Jh�<��JǯO�����h�60+�yu��g�<ْJT��Re�vײz�>tГ��c�<�q@#d��iC!,{#ܸmPwj!�DX�:�{�R-�^X��ݥRv!�N�Vm*=kq� �v�b}!�4l!���vV�xS1eX9�$z�ǒ@[!��ȅ(��#c"M�@�,YӐ��:D!�$X~�B�0wJ��H��%c�60#!�� ���s�@�f�([Q8��"O�x1�dE<J���Æ�?W�8y��"O��RQ*&cԹKR-P#<��XK�"O��r�P�}pf�����4_��e�T"O,K*�x�� f�M� �є"Ov��#u{lQs&��8���(w��Q��U���h^���)2y�]��NE/L�!���8\?��#�&*j�+wJ�z�I7�Dy��y�)�'��i���>8yѵЎV��ȓ[���u#=�����	�rL�OZi�Ý���ÓJ�z�Ʌk�F\n$Y�`D�;w� ��I$�:����m�-����54��(��a�#� ��O�0('T�$�h�@��"r��d �CLQq �ΪdEZ��ю;�S�i
���&��,m�q��+mt�C��)w3�d{@ԇ �J��2A
3���ZgcH�VJUh)U�+&6M�_��������@��O����m�h�!�$���ɤ��= <�a`��7%ɒ�H��O��+��p#Ll{��'1��跈�	�<�g�����2�N��9� A5y�@��^�C]$�`�?a)��*W���Vz.�
�2�x(�i�\���5h�8*�P�v$A��l�Â�Nnb�����@:�Y!���uR��*:�1"ŏ�7N�͊G'N�3*���c8�O�p���K�L
� wkJC�Mh��M����Ks���9��&x�x��'����" �w>����e�;
����r����z(9�'S��z���
3�<�j�
}�>qsS�X�'��pа#	""�L��g75S��B"�9�(
�*D
|�:y[�'�e9g	�-D A�L�s�T��IԊC⥝7�C�E� �����2/f�(Z��T.�.<�@�^E* �2���tDŒa�á��#>�`m� ]f�	v�*=)��A~��J�P�߄iU
�BP��1p�^�)Q�m?�R`D�fܙ���	���k��c�Rd
v�\({�a~RG@/j|�ѣ�M8I#X|�Cۚ8q����8p̤Ô��-0�����-bp���;O)Vh�Zwj��]�a�2���@4<+:��
�	��B�I�v�!!��W��&G�
Ya<
�U�`� �P9ot��������)1��������	_k
�ɤ[Ȋ�������JA�,ۄ��/ќq�%,�.�Dcu�S*Nv0���M*�j�"��T3S�.��䆑OԴ���-�J#>�(';	*`PW��<"��!1 �L�'0�ZIO�̥8ROC	%j\<(�#�!"�|Mqt'�#�@9�%�h�*Q1%�Dp�(��'�����,�;b�h��/��iBD͹���>�s���$�f��f䔝����q��:c�b�0�o�Z��#��@�!�_�� ��FOƊ !�^�Er�8c��G4�¥��Nͩn��Ht�M�5�pa�]�ބڶP>����+snp�kZ���(�3�����E�^��IQUC(�O���q��G\l�	FA�6z��2$��6m��)�d�b�i�g�I�A�d��g�cu��-4y�L���D}2Y:WL����ǟ�� .Jf��N�8nkXaI��ӄg����C�&�!�dV?.1�te�"�"�Ǐ�2P�!�ě/V��m9 �ǳ�H�۴���!�[��DY���<�N��'�4!�D_K�f� ���i�Ak&���!!�D�t���	R�\j�l�G�ԁg-!�dР
��d���1QH�
���3!�$�8G�R,�t�Ɠ�V�9G�M�;!�d��kA��XE��ce��2t	!�d�>n$��MM�sH�s�
:"�!�$����C��o��X����Q�!�$�6��Ȉ7C��,�Z�iC�O�y	!��:)Ӕ�f�����)�!�,!�V�5� 'X�9<�h��J&!�䙼%�
�h5J؍9F��7��<�!��J�t���!���%�����-&!�ě�$���Z�` ��QfG�.a�!��4o�iߴk����e���!��i����gM�#vE�EW�m#���kE䚖�'�y�CNJ;D�B����ˇ,�\�X	�,�T�pQK�86pĻ�@O�l	j����+a�X�	�'-�9�1��N	�� Vk̍U�i ��d�	ʒȠ� �'��O��6*�&��`�ef�q�Q��� �HR�%/e���C�%D���iȸܠl��d| Q�O?7M�T�e�C/Իc��೦^4�!�䝫��9�㫛/nZEQ�O �����]ڈHjK �y�dX�lX��MC��Ƽy��J���>i��	�^�$��M��~( |xBfF�QBje�g�um�B�I1(&n�H�{#N<y��ϋvߢ"=�FE���$:t�/��ED\�ۑ	-��2���2��C�	�!N���Gb�+/��p���v~6�	7�\�(eE��)�'!L�I�R�d��2�O
p��5@�<"C�	�ˢ̹�,��W����ea�;#[|�d����$L�	i��9���r�
���"�;�УK����y龈��Ix��	��)�y�d�@�8� �"�Т�*y�'����tk�-@���OQ>-+�VR��!��X�)U�2�e�F�c
 ʧW\���'W���SC�(:�,�Q�>��g��T~�iL~�=��'�6��ŚSgB7+Qd����g��t��gՂ����Ѽc@��H%`V*_>���ɮ�a��� y�a��ˎ.���1�C�O|�Ё!��A�5�4'vڐ<�)B�gR�x����	��c�X�$k!�$
�ԊL��Ϣ��M�a��u�� �ȵyB�0��N�7A�[����e��B��X�gg[�'�J�hI2D����&��^ԠA��Fy���yc��R:�,��kڵw� ˓��2�*��{�'&��`dٹ����u��1��ۓ]�b�3�f¡}�>X���eN&�!�\
<���Ӵsx��`�$�I؟xP6
�9J��I�%�C�V+�����/�I�!;d͉#�2�,�*v��1��Oȶ���)U�c��j�8B�'�vm2BCّ0�q�b���L��r*֥$8�q ��.�L9cٴsW�>��"ݘ�%B!5�:���oK�F�5��C��ç�D�h�$;q�+W,Ilx��Hҍ�f%�{RhO+,��@����nረ�/�.��=���P���%��O�U��!_$ѭq���	lV�"O���0n�P�
�Ǖ�	y�m�U�D�x�d�;��B8�h�����i�)��#4�ԳJ`ʄ9"OP��r��>lH�ʙ�	a�<qwD�.��Ӗ|b�����2�vL�FF#%�Y�)D�l��"U6z�渹!HJ0C��Y��g�`�)���|B�Z�b��!��ש*�B\�0"\��y"@o��t��
!�
x�`���yrj�l�dr�O8�BQ���ߛ�y���2���)%Mܟ�bIA���1�y����;��9�ĤJ��PTEK��y2�D."e�A�x  �@"����y���ERD�"s,�x��d"R�9�y�K�E��X��Áx�,%��*�%�y��ԃ+`JH��F�(K��O7�y�I!y�|C��+n��4aΚ�y��"~��C� #$����ĕ#�yB�M=(#^�yũW�jm*Ջ��y�[%yQ�C4�L>'J�R�N)�y�fR�8=��3��;*� {�D���y��C&�lY`C(%4�5��L)�y�̞.8I*�H�&���c�K��y�#� �X|�Tf�L��pV�И�yU 1N�TS��7j���.t�D�
�'F¡�\���6��01u�X
�'��)��㑪6�5C1�)=H>���'�t��Ae-t��P�gnB�0t(���'{4��AEӞ*Fp�	���(.缝 �'P�U�Q�²v�n1B-S)�U;�'-�x�7U(02�vLA "�}��'[�0RE��*(�#v���^̊�'"���G�އ=�^0Xfg��V�I�'�p�Z�!�9U� Ui$k:�
�'
�����.�HE���T4��'H��X2�N�f�a�/ڲ\��2��� ��zc#Zy���SaJ^��H�q��'+�Q�irE�0��FJ5��H�z�(�7}�JN�w� ��A�O:f(R��^}נ���7;�XI;*O�Y��J�P��tj5���Q?�W�޳*e".��R�ʠ)�l�O�9�BF��r�� �LBɆ��)�
P��%�U�VLa�dZLI��#C
�����
)m�)�6���If�A>x�A��ж#/T�`�kd��'H�<YU�OZ8��d'�C����F��e�ذ�S:Jw�42΀�M���B�a�4n��5��{�H�X+�\`%��
�4mPCi�1��Հ.*B��)�kj0 � A�$���*_�U���V�@�$#�+|�T1��SaoN�Z��4V��<�!�UCj�i���qc�+:��4��*e8����Fb���m^�gN�	 qzUa4&��q��O���L�l	�@M�8����F�' �@�� ��T�}��S�O[�$�ތml*��V�=Șd+f
ĖC����&`�I-a��a�$H{ؠI5���<��Y��K���H&�T�`�׈oa���E��U`�O�%y�Q���B���ɲHJ�T�T-G��S��,cdd2V�V�}��|��"��oL�]�"f�c�l�w鎇L,�S�OK��ic]Ȗ�p�� 7.ERq���]f1��ٕL�H}��]�'E�u!*�j���c�;�  ���C��`p�,�~ I�-Ʀҧ'� �0|B�-��:O�ٓ���b]��;��П���$ڽ)�Z!���=S�� ��S�n}�@���w8� -�c�b@���я)��s�K�q��ulL>ɫே.]$�,��)�64��m�7��<
�x��U"�X��lK㋚�rH��	�F��rt@S�Sx$z5M��z�4`��[�G61�7�"W�ֽ����$՟�O��P+��cT��Xh�:�%�O5"nR%:a�P2�>��)1ʧ2��2�J�51������-.���!�'��]�'�n��r-M������O
��Շ"M�p2q�H�D�zU	B"OT��̏ If쨘�i�/9���p"O(YI��Y6yMtj�U�!�zQ!�"O�!wK��~�����O�o5���"Oܰ�(� ,����&0���"O��"��[��Y"CJ�RzE""O�`K���:��P!]�cd.8{0"O���� D20a��� -:Vڄ	D"O*x˳o܄)ݮ��aZ�"n9("Oځ�mp�1Xe��1��E	u�<���]s�-�#�fG���r�<i j_)'�&1J��W�`��@���]l�<iT��Ka���cP(T�<J6�]k�<I7n��~�
	�K<H����ng�<y0�9�*	���4tzݚ5��e�<�c/x�x�QpH�v���g�e�<��B�C��!�-�%G�\2��Mf�<�	P�h8�!����C�@����b�<�AɃVPt�p���,P�nG�<�υ��c� 5ݐ�I�Áj�<�K͋~f�� �ea�}yrJEf�<i�j̦K6�Y���lD�m�dJ�f�<�GoG=��(qdG;
�����\�<��`ǧr>晐F��qz\c�iL\�<���2{�*s�͛��tY7b�[�<i�aثs4��@M��y���4�T�<aWFc����jى(>���dWQ�<i�(�4a(�h�C��=����'K�<m�!^��s�@ʾxk��4���y���� C�!��5�� E�*� B��3f�X]��"Ub�LKr�:u�B䉩l��p)��U��ᅍ�ѺB䉝�*�h�b��4M�]���@�P�B䉏A��'M�&�N�+�-B�6s2C�	4g� ,�⣉5(e҅q�%A�%f$C��)3�|t(h�LՀ�[��2W�,B�	�H�x�{��*]�(�(g$ѩ3X�B�	�mRV��b��,X���gS�B�(6��LN�>�"pZ�&�+>�~B�I��r���nȁ^�բc��4bB�)� �MB�%w���L���d��"O(���`�/�|(ړ+�t�4��"O���C	V�p�0��A�Ə qN,�"O�3	�a5�8q��5Y��b"OV\Y!#[;9���Uś�vGvl0"O����;]�IR�M��r"��Ȅ"O�A���^{��sLI(�Ru8�"O���śU�~9Ise���N��p"O��#��.G�$-�oW� z��@"O�����_:h��*b�BX�B{"Oy�(D�R4H���#G�=�"O�hRV�ð~E��X�AD���"O�<6@�:l�� "�@BY��"OH`k�i��B
��1ԻC/��Kg"Of����� ="��yC3Y* ���"O@�0�>'&}���7E���U"O]R��C2+6`���.�|EY"O��%O+z�N�p��(Æ��S"O��2�JU������TF�[#"O�P��$�*~�8����z�g"O�|���Q�6��#���r��+�"On��v������AT�b�4YQ`"O�d�R@�9��`��b>t�`"O&��F��#|���h�.�UMJ���"O�H��� +G�<0��	;1I���"O��)S��.Znl�ĺI���:�?D���Ȗ�3&�Dh�BFj�9��#D�x0C%>�꼚�"�l�I�D�"D�(�����ZԘ�P�TG�0إ.>D��B����j1�B-N%;^��S->D��jB��/��h��Q�p
�ȇ�:D��F�[q���P�8ơ�v*OI�R)o޽Y�e��P "O6�),��\@���P��-k�"O8����<1����7@H˲�R�"O���AA�f�� 5ŀ�z (��"O
���+t1��C��Ve�pA&"Oh���Q��8�,3+����"O*<@��S }Ak�G)V�+�"O�$P���iZd��� KW���"O��A��� 
��` ����r'"O�ݫ��� PJb6���!����`"O�tv�&�Y�6- �m�"O�\d��A+q������ 05"O>u3���F��<;�A���2Ѫe"OfU����$r]F��j+l��-z�"O��aBL�'��Px�	�d�~tSb"O D�$"ն3I�q E��;>h&|�"OŉFAE�>�������w�bI��"O�q��eܳUJ֙QaHG"VHt��"Ob'd��-`�7�����J"O�HA�^<`hH� ŋsAڬ�"O��1ǩݽv/hP+�AI5t<^�XQ"Oܴ(�W3qV��q7gQZ�1�"OT�k�*Ң,�TQi���)E�	�G"O�]Ң,���^A�YH�Z�D�h�!�X� -�%M"�R�\�x!��U%x2ҔI�j�62@#��Ɓ1!�$];�%�A��d+�!@�X�v�!�$���%�� W�	��`���D�!�d�'4���Hv P�sܥJ��,m7!�Dښn���6C>�ȑja�6E�!��̈r�n�qc�>^�E�زP�!򄆊L;���+C�/W�q�%N�4�!�� � 
'
�_�i� eP�<�Je�"O2� JSO(�Ly�-�r�!�6"O�HcA�J�"����':�A�"O�)���!(,�����X����"Ol���$L	vd��hW�M��uI"O�y �ěrF����
6[���d"O2�BR(M0��Z�)�S�Z�C7"OD �r��[�����ȧ"�z�sb"O�l�Ǩ��c���I�l X��"O���DS
 �0q���QXVi:�"OD-1��"p�Jy�i�5V�IҒ"O�V�?T��0@(׮ut���D"O��Z����48tX#�fOZr`82"O���p��0�y���	U:\�d"O�=+��Q�b���JO�ڶ"O���E�Ek���"w���\�<HU"O 	ig��#U@���T���jU2�ʖ"O�Y�	I�Y&�h��G[�#^�Q)"O����(\P���b�$,ڱa�"Oll{��b���C:7j�"O���e�ͼ{����'=�p y"O�t`�EA:Nh��@Ʈ �J)��"O, ���
�'><ȓ�T$E���f"O� u��I��e�;Q/h��"O&�� ��ܜ����$�}2�"O¥X���z?�̢j͞
�B�"O(4#q�8d���	��P` �1"O��Oυ?Eм"g�s�:���"O~qs&��n"���&�{��ds�"O�ubU{ìys���:!����"Or��#M�J�(ʦ�إt��f"O�0�mN�nQt5p�l�K�֡�"Ou�u�Ι3�*��RIQm����Q"O�mI!�L�Q�䉃w��1��S"O��CFA�"P�QW��<Ӣ%#�"O��j�j��1*́D����P�C�"O�8;�h��z���f�І
{��7"O(X��g
:�,���.��y[8�;�"O<��B��~�h���,��3�N0��"Oh��[&rR.�Q�ʏ�N�x���"O�Ё�L�0<���G�M��	e"O�����9#@�ˤ��E����P"O�����%�����D�@��T��"O~T)r��f	X��C�=yn�8��"OBU`�C�Hz�� !>Z�I��"O48�7���|}�" �O�Oj,���"Oq�3A6
�rM�eO�3A�Ę"OB�qŭݯ#�H��]����sd"O��"���#B�� ���� ~�*0 "O��s�Αq �Uqc�_�Q�;0"O�� 0g�1]�@uiBl�+��9�"OM92g�:���`�d[�E���"O  8��"1����P)V4l2w"O������� ����3.��A"O��0jߺ=�ġ���+N0p��v"ONiq��J���P'�.b0Zٙ�"O�Q�pEQe芰�v�Y)aw ���"O�
b�]E�Lӄ�ϳF]"���"Oʌ�p"��3(��{E�:f["O|$@gk�SH��P���#U	ʴ�yҌ�k�ء�1�T4`��s����ybO��Zh����W$,�|y�I��y��@�VB����6�!�d��ye�2ލK�Ô��4#0&�8�y
� ��*�-�WS�4���>�P��e"O�$�"�1����D�f���"�"O�Y�R.D8n��ɣa�7e��u�"OR�*�	�
��e��3�t�"O���c�G�V��X��/l���"O��s�o��zĸ��;<o�Q�"O�Q�V��'�T�0�	i�iD"OJ�$��]?��� �4M[ڔ��"O�-hP�@�%L���-Ld�C�"O`�
�E�N���c�]�M/~� �"O��s��1F��f^�'���w"O��8���IƜm���4H�z�"O�p;��|.8|����
��e"O6���M�<��{�X�;�dE(�"O~�kE�?�Jt��`҄:�Q�"O���WcD���3�A.+V�2"O�	lʵ� BG�/: ��"O�4�7oC�n~��gG�[2�Rc"O�eӄ�H�@UX$h�G��5R�-�"O��K�cU 52�!��:u�"O��#�
�8<���Q�_�P�ٵ"O��9�g�R@��"�[��F��P"Op`��*������
kD ��"Oh���]	-PH�%@�:X 2��"Ob���`�2�����D�@%��"OP�C E�HY�j"��s�	��"O.D��N��L,�볇�%����"Of�bv�R�O���qD���b~�`�"OT����6�j�2ƇQ�"%��"Oꤳ ��g��嬓�^�^E�"O<��f   ��     G  �  �  �)   5  f@  �K  dV  b  =m  {x  ��  P�  �  �  Z�  �  .�  ��  ��  :�  ~�  ��  V�  ��  /�  ��  ��  B�  ��   b � D + �% �, '7 > �D 2N gU =\ �b �h �j  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>���f* 2���y�#W�@ݳ�i[)�d)�OЉn�g��|��?�u�)[�^�(p�
��`O��?��sY���ٴ���u>������\�a*���Dl"�i�T� b�h�Ioy�퓚[)r��,�6d�B�10�mIܴr��<Y���g��O�>"��	$oZ�a��Hb�ϣDp��O��M}��� V�P�&=O0=b�DݔI ��g! =���p3O����?� ��|��+�KW�՚�;����VxP	����0�'B�'�.6-ʫ1O�y��K�zM�ii#/17�t�ӄ�;�� ����O��}�ʧ)t����Ȏ��;��A�eG,��'=��-�\X����K�XX!�'�0L��]2h�ΤȃDO���e�%_�,�'���9OP�T�P�i��2�&@�5�5�d9Olmn�j�����v�4�f�a�`MkU��`+ J�7OV�d�O�dK9,C6M3?�O�P��eE�m!�m�:�����(tL��YN>�*O�)�O����OF���O�Y�����~�0��(P����<q��iP�C�'��'���y��  j&!{�it�Te('�C!<8j��?i���S�'H�
d�bnK�q�Z��&*S�ܕ��M�6���'5�*%F�͟l�'�|V�T�4��9R܈��٨m���(G�����	ߟ���ߟ�~y¨|�N)����O@%��������l@Kj,�L�O�Il�f��ПX���@C��К7tR�b%�7!D����BՖ$͂em�o~"/�U��5��_ܧ� �� Kx,��u��P����F-�<����?����?���?y����MS���pq���C�:�:��$|��'��nt����?}sش��?���bR�@�_
4@v��^h⤸K>A���?�'qɴ	bܴ���O�-��(Qb�@	EE�Vj��,_����ɒ�~�|�T��S��������*g�œ��L�W�t �����	fy��}����"�O<�$�O�'-MT�p�e2rR�ْ��V'
��'�$ꓶ?����S�4@R�'Y`��s���r�@@a�	$�x��.��q��T��ӚbGbeNA�5מD+gQ5� 1�
��Ԑ������I����)��|y2�j�x\��I ,�,��O>Y���H���-Q����O��o�[��;��	̟�����Rkf%b�kS�Rd��{�
՟(�I��nP~��T�Y���}���>r�<Lzc�R�G�z�:REE�</O���O��d�O����O��'Z�f9���C�0>t��-�2K�v%)d�i#e�3�'���'���y�z��.D ��	�j�@��i�%QB�$�O��O1�:��}ӎ�	�M2���%�<?�mBR�M�.�J�;�xã�'��0&�`�����'�m�5C��;��Ѷc�<aK�DC�'&��'.BP�\��4{'lS���?��0�Dh3G�<� P#�98���>i����'��Z4��4)6(��IM�"��DA�OPl���Z�Z�ɡ��0�)�#�?����Ol1�%�KbT�$�7�(W��ON�d�O����O�}���vil��!����`�@��X�T��O �oZ�{2`��џT[۴���yDM�/���/8���ÈM��y��'��'C� ���i��I�w��j�ߟ`�S�(S	J�t��DU eQ�X$-&�d�<�'�?Q��?1���?I��4�Rl_������S�������hd�Gǟ���˟X��"Ĵ_���q�o����E��"��۟x��o�)�S�|s
њ�mAG�|���d�N\��áE�u�+OFp���N�~��|W��Z%�Z?5�j5铄��U@.ui�a���D�	��x�	ş�Svy�r�8#k�Oʨa����L-P؊A4}��1&:OX nZK�
�������'��ɚ5��n�hQ�FR�jxZ�P�Kͅfٛ����i�@իx��d�[m����� h�R���bɪMq'�&�*��:OH���O����O^���O��?u��(V�9�P�k��>�~����Q֟��	ϟl�4��<�'�?y��i��'��T놯שO�JA)��3S��Ē�y��'y�d� }n�D~��ϸn��U{@��-�⣉G[l�}Y������@�|�_�������I� ��J'��X�vNN�,�xc"��ş0��@y�Nn�θx���O�$�O��'`N$d�Vg^���Qf��~��'�d��?���S�MחgӲ����Ǵ
A�|��ߞ[�t=x�W�~d�O��F��?�6(�DU�ʹ�"F�Dz�`[��]8E,���O�D�O���	�<���i6a���z��D��͂
3S��҈!���d�O�Ql�V��h����p(�n�r`j%���,cw����ߟ���d<nZv~R��Z�p�S_��Y!qf00�2'�V�qP���m��D�<����?i���?	���?/��#�n�M
h�X�m1��1S"���-�l�My��'}�O��a��ͅEb ���O�f�bg]4ZX�$�O�O1��̺&�z��I	����ӥ���҈*X���j:uB��'��&�`�����'�PT��t�x�P�T�Gy���6�'��'/"U����4.��\`���?�� ���갡M�,��q��FD(y�:�A��,�>����?�M>1Gf��A��@���l�eJC}~�(��5s8԰d�ib1��t��'�b"?a���24A%���g>%8B�'��'g��ȟ��o7�#�+�+h�:4����4�4-G�!X��?A�iI�O�9S��U��f/	�ш�@��$�Ofʓ6��p��4����30����Q��e�f�[�4p�������m`F1��<Y���?9��?��?�����<a�EZ
�LA�bD]����٦iQG,
ן���ɟ�&?����:��"U�B	�<�I�J�IcV���O��D�OD�O1�xa�5EO�8z�٫�ODN��P��B�v���δ<I$cK-��$������X�V3��Ss�TȠ�#��wy����O����O"�4��˓#��+*<�R
�B �t�/�@ԋ`F��yBci���0H�O2���OB���aTL�#�4�B2D2HJq�7m����� �����>���.�V�!2#��6@�c�A�"ǲ�	ݟh�I�|��ǟh�Ij��L�=r�"�?Z�um�<t���+���?���{�E������'��7M>���1I�h̩��B|�*/Q H�1O<�$�<A񊋻�M��OH#eMl�RX�7�фn�;<�x���'�N�Op��?���?���q��	�c�کcG�&kN�X+��R��L��yrn{�
��$�O����O�˧abAЀD
!`��4�����%�i�'�6듕?i���S��Z(�jp�0,X+@A�G��;0"���i�)$��M �O�	�4�?� �#�d��" B\�Q�@ *K< ���F8`^J��O��$�ON��ɩ<Ƹi}�k��A�(h(��.�u�`R� ��	��M��B.�>)��ZR��W+C!tlU�$�Y-!�(x���?tB���M�O��J�J��2N?a�B��mA�`� S�f+����Ho�@�'���'���'dR�'!�S;ˍ��N�Ezh8Q�/=�����iy�8@��'"B�'��O#r�g��n�'}\��GB%p�n��pe�
 v��1�)擼a�tm��<���N'&��X�TƵ,��0�lF�<i���J7j���������O����F����D߁���#b	�?�����OV�$�O6�nQ�6��\t��'�����&�HCWlėUl�d�Hŧu�Or��'ZR�'n�'ҥqČ�"(C��s4D��D(\�r�O��Q��c��6�U�s��'2S�UҮ`�wF\�],��t%Ee��'\��'l������͟'�U襨� ��(PD�؟�۴X������?�B�iK�O�.ԉ��z��W���&HE�
u��O����O02�&}���Ӻ$��(�J�D���q�b���My��4weڒO���?���?��?Y�j��@�!��#,��6O`SK2X��Q�4sBJ����?������?���$��j��)�P�P�J�5fb�I����`�)�)��*J95��a $�7]�Z��r'Z��'�t�k��
]?!O>A+O��#�)�� 9���(�2A0Ђ�O����O����O�)�<Y"�il�a��'K��Q��6X���bMH�EL��؝'�7;�	�����O����O�X{G�</x}�&�U�w�$0r�~Jj7-7?���'���I.�S���#��(v��)��A'��	avba���I��D�Iޟ��	�x��NG�H�D!{��K�'船�a�W>�?���?�c�ik�çS��A�4���Ҥ��`sF���D >Y��<����DZn7->?��K�7����p ̺#6�i�iN>.��83�*�OʬcK>)+O��D�O��D�O0�;�8\�W��`���H�.�OD�D�<)��'�H<9���?����i��L�lx'EH5$%��u�Xt��������O��!��?�b��rBAIV��*��1�EW)���,Ǧ-�)O�	U�~b�|"�͗u�����AHf|�'
^^�"�'r�'����P���ڴvPT�^�m�4��V�$��E	��?y�R�����D}��'7B��Ξ?z�.���-i�n��t�'�˶h��F���)z�*���/i��)� n�ië/*Mvm�����]���d3O(ʓ�?y���?!���?�����I9q����	-+t<���N���V�mZ�/BV,�	Ɵ��D�s��B���#C�)?Ӣ:'Ε [�>y�j��?�����Ş[�Mb�4�y2���7�.CF�=l�nY��L�y2�B'dn��	�h��'���I�8C!�,Zd����Sg�fi���	ß,�	�<�'=t7m�j�L�D�O��䎠x~���l�h4���Z�T��⟸ۭO��O`�OV�1F�]g�m3�����*s����f/9:x41��&2擼:}R&�Ꟁ�l֡ ��l����8�aqB���0�	���ҟ�F�T�'����'@�>0�	�tn��G�����'D~6��L�����O��oS�Ӽ��S�/�PXSq�c���I l��<���?y�r/��޴���)<u��'J�6�)��X�O}r���	!oXu��E3�$�<ͧ�?a���?�Ѧ���:n�,pTh��
TJU�p�a���'�V�$F�P2��'Q���������B��h�N�j����'wB�' ɧ�O/���S]�&؈�D��tq@�C�P$��k�V���e�4F��I�	uyrn 0�ŀ*�>t����@��08���'���'#�O|�ɪ�M;�mW��?�N�DV�d�'�:^���+�*�?�E�ig�OY�'\R^��* Dޒ$} iY�i\�wZ4]�͟_��el�E~bi6��@�O�w"d��䀕Ó:{��r�'Ȇ�y��'"�'A�'�����8)�|���%h"-�NH@����O �dU����u-YyB�r�@�O2���&�1#w�B��0x2�#���O��4�z�`#�uӂ�D^�Y0�Uj�����;VM�B*����D��䓏�4���d�OP���Q�����<� Qѫ	�(+����Of�>2�V���9�'H�T>��-%1����0Ax2�-xV���	��?�OQ�"ׅ�\��$?θ
�Q r82���� �i>�ذ�'F L%�"�A�?��ɓ��ߣ@�qC,��8����m����i�<���i���6�e
e����y��kV)Tk'�	�M��ƭ>���43X��[H�)�����}Θ(�D&�O��dC��6+?�;H�!���x�ʓS_�b��� 	��d�6D� ��͓���O��d�O����O����|�W�ݰ[�6���-I+��2�Γfk�6aX�r�'��T�'��7=�y�@�z.�˔)��$����`F�O ��"����"7~���������h^f�FX0�j�������hS�IKy��'��@�0w4���ɏ8'�v��'��$=�'�B�'��	�M+ $ԓ�?���?�#��=d�q�'L���q3�iՄ��'�4��?�����8:��ʒ�e�@�I��R?u���'���SM�;`��v'���(�~�'G�A����6N�(�E	S��q��'�'kb�'r�>	��01�^y�0�M� ����qMQ�>� ��:�MK/��?���}`���4��%Q��4J)�s�ܧ(��x��9OH���O��d�N�P7;?i��O�8_��� �6�jA���ӜE�6J��Kpy%�\����'�b�'���'� D:�ѣu������I�P��^���ٴW�H����?Y�����<�Q_�]?ո�,�D�0R�c������ �?�|�����,�q�F�~"(h`��f"9àH��򄁙c��� �p�O�l9��
A$A*?��+���s)����?9���?���|r(OtPl+	u��(%���'�G��{u�Ԏ)�4Y�	��M����>����?���{��Rg �<(;��SiЬ6�^H"�c�3�M+�O�<z#iܲ�����D�w���1
OH0�V�� �DT(�'��'��'���'���1�Y#"�p+!G�
`%��ia�O��D�OZTl��$"��8�޴��Do
4�c�0Ou��Z@�9��SL>Y��?ͧ16D�*�4��$ћ"M6U*�Q}A�y릈K.5�%�Q+��~|�X����ٟ@�Iퟘ8�N�sn�T�u˙L�髣��ޟx��Ry�li���4L�O��$�O�˧		"e��Ƕ^/����6q�z��'�Z��?��ʟ�)�`��w#>�F#��@�
}S�)�it9� bX�c����|����O��H>!T�~Ι�BoC�+��|��$�?1��?����?�|
(O"pmڎ������Ȉ�
A�	^�&ZMB�,�KyBdӾ�p�Of��N5�v��&�	u��	��ָ0Ԩ���O�`�s�p���h ɡ���V�O��հS�O UY��P@K�f^���'��Iퟔ�	�����ß8�IB�T�]=f�ܙge�FY6��5�N��7�ƥ��D�O��$&�i�O��mz�� ��ǂ�\,IXv��U��d9�)�S�<��o��<9@kR�sF�*#�0~�ڭ:���ybΈ�Um ��	�U�'o��ß���>[�bl΂����vCߤv���	�|��ԟ�'�$6�ܮvL����OF�Dg�r5����J2�Db��T��tӭO����OȒO@\�1�\)$c���@b�?��<�D��p�g�?s�}xI$�S�s�IDȟ�Y#틥UԤ�a����;	��k�NB՟,��֟����E��wo���"	E�������!VOR��@�'�,6��/��ʓ+Л6�4���'�#M���P������0O��D�<	S+M��M#�O�0�����'� h���gS�zM��Y��8ԡ?���<����?���?���?�!��1�� i��\�`�Y������`�L�ßD��ɟ�$?M�	�.�hQ�A�/�.1��-$�@A�O���)�)�@@�k%/�"�c�����I��*����<��l�a�|�D�/����$ހL�ʔZ��B�Y'V8:�n_;tz�D�O����OP�4�X�+��)ڪ	��KO�h ���II�:���XGc��yB�m�6㟰h�O����O~�8z%��їp�����l���.��$�{���Q>��#��?'?��� �5��I*���A3��	ßt�I����	Ɵ���y�'(�Aj�j"�'l�J���ԟ�����<1�4@���'�?a�iJ�'�,	���H;'����NX�a���r�|��'��O4�y!c�i)��3KltDb��O%"dA�Ī�1H��5LܧV��$2�ĳ<ͧ�?a���?�`��L�<��@@�� 0� �2L��?A���Mǟ��s��O����O��'kfz	�b�)2�,b���+n ��'\���?�����S�����[��Y$bT9	Y��AA�L0��L=YFF�#Q���7�R�V�	��4#�J
�k �R%��6T��I������`�)��by�a�x|�%S.y�<Q��H@�^>���R	>Z:˓g�&��AY}�'%bY��8n�	l���L��V�'#�).q�����֝8j����剸r��9��*ӲS��#��f��	Ry2�'"�'��'��W>U���>q�6Pϐ?0�l��*��M ��?���?�L~���u��w¨A�ʙ��,��sbɕ����p�'(�O1�����q��I�v9�F)*�x��E^�S�
��X�`���'[�1%���'M"�'>�1��
]��a�c��{ibmc�'�b�'�W�X3�4+H������?i��\��%�R	dR !�O�>��MÍR�>���?aM>1B[����W��\w>��G%�H~�  zF\�S�ʞژOqDL�I�ZG�*ڑ
z����+(Z%q����b�r�'�B�'�B�s�i���8l|<��*�xK�@wO�埐xڴC#�!�)ODmn�H�Ӽ�L��NyJ4ol����<y���?A��/d��ٴ��D�s�@q��'7	θ:�	Q{�EMG�lDa���,��<ͧ�?����?A��?aI9j$��˘t�j�����D�Ǧe ��M� ��ƟL&?)�	*��Ś���>4J��b`�$d��@��O��d�O6�O1���0��S��J6�Ղ�>�A�׬wJ��`Ր�x2�-,Y�b��Q�Ilyr�X1:�y�A(�P��l�vJ�#e��'�b�'��On��=�M��N���?9�1l2���q �z�hBG&�?i�i2�O���'�"�'DbKM�Pd � �'��f̊���΍2E�B]��i��I:7��Bc�O?��$?��ݚZbL�@Ў^�dQ{�B'%H��Iɟ����h�	ɟ���I��gt0�� A}`mrA��U6c���?q����V������'��6�#�D�F~;b$5h�$l��f��f�t�O��d�O��A�
�搟�؃�í:8TXy�%C�(Ĕ:`�I���?�6�4��<ͧ�?���?�fK�>-0h��'Q�`vj����ߟ�?�����=h�G�ğ��I�H�OK�,�3 	55ߔ�[�mL���O�!�':��'ɧ���-����rN�d۸Z�H�;>9P@hZ)l8�֔��S04W��IW�I�[e|ِㄞ&(o��x��o2��������͟ �)�@y.q� Q��kV�0�}�"��=AVJ5q�
ǭ�n�$�O��oZk�:��	��jݑB�� 3S��dU��۔CFwy���S��Ɲ�)J�02@�EImyBcKm8�"��=f:88�`IM��yrP���������џ���ޟt�Ot����#W1
8�����_�t)UDlӤm�u��OZ���O��?�������!x-�p!1E�d��31DB��?������"XH�63O ��V$M�N#��]�q��鳑9O��1�jU��?1go2���<����?�BM���\�"�.]D����i�	�?y���?i�����립�gW����ܟ�1ĩ�"Q ޹R�@��Mv�HU*�Z����ʟ8�?���H���ʶd��MԲL�W��f~�mI%75��(D�VZ�O;���	@a�x�zQ��6*T��p
A+%�'���'���S��Ȑb���0����IJ"%]�E�sK�ϟ���!٦,�'
�6�.�i�] ��P�*�2��BKG�$><��Sls����֟���DHm�D~�*�O�� �S�B&�<9��؈@�����)�B$ֱ�s�|�Y��ҟ�������Iٟ��%�M�}-��wG�.AŽ� �{y"�{��`�p&�<I����O�E���tS�_}ᐽ�bh�>q���?)O>�|b��#*0E[4��8O�j���/�i��e*!@�Q~҇_|�b9�	�#��'���*�jQ��f�<��5�b�O@���O��d�O�)�<q��ic�i��'���6,C��A��|����'�F6m9�ɳ����O����OPɀ&�I�V���
� غ��ub$�U+U/z6-"?9׉�<^3���4��߉.ԬÑU$D��R�P�<��������� �I�l��`��w�L�wF
�3��p)M� ���j��?Y��)[��ɗ�M�H>�"��0-tVm裣R�2Ĕ���?���|22��	�M��O��95� p�A���@�F�&0+�xz�チ�?q�)�d�<ͧ�?	��?S,��!���Y"f-x$" �p�!�?Q����dEڟx��O����O0�'o%Ne´ �:=yBpw��="-��'B���?����S���H�c>Li�3tCvl᧏�%(������������O����?y�G(����B��s5���/Q�Dp�PoG��$�O����Oh��I�<�·i)1 ;��aW����H"bD�����M���į>1�i�Y:��W�j��So� :
ɐ+O�9;�`���#Y� u��|�A*O�i�"PV�dT��f�%,�TC1O��?y���?���?Y����)̟H��4��o��\h��,�)a	�m�	;p��I�t�	X�㟤)���� �3��}��&SkS��e��?9����ŞS��13�4�y	�YC M1$��$�Ht	�F���y"�T`����䓫��O��DQ�>�eyڠg�@0�5�� C<������	񟐔'��6��A!�˓�?)eC����*DK��Tp��
ˠ��'GR��?)���)߰dSAE�i�2��p��=6�J��'��eiC��5I�n#�i���~"�'K�@��P��`�b��9�-
f�'���'z��'�>5���n5�D�ͷd�r\��,R�|�dy��:�M{Uo�?1�5ߛ�4�0P�C�ì\eQ�/�l$�;O��d�O��ѻ��6M(?YT�C#Ht��;����aɖ6R�F p��N�s�R�%�4�'j��'�2�'�B�'=f8�FkR�F�0a���-E�B �5W����4� -j���?�����O�n��K���n胗M(&ELXI���>I���?iJ>�|b��V�A��*��/0���� �m��4��D�;B@��'�'"�� L� �!AY	V�`�Jjn�5��ԟ��	����i>�'��7�ȜX� �D֫M3���O8��T{A�z`�����?if\�������I>�^�Q���B�>9:�h�b��r������'bX٣��?	�}��;Lh��h�24_��ȑEĄ$4,��?���?����?�����O���I�&+�\�@�� 4��R@�'�r�'�P�������'�X7�0�䏈E$P�°+�"A�����H�$��O|��O�I�%
��7�$?�#b	a��y���^����d�Y?Hk���
���'�X�'�"�'��'��X�J
�g��[p��o���yF�'��\�XZ�4>���Z��?����i]/P��VD&D��Px ��;�������O�.��?!��;4h���-�>����O���ԸhF�+�~��|�a��O��rK>y���uF+Ѭ��X��Hq���?)��?���?�|z-O|�mڕe�z� �O>3����������͟��I6�M�ξ>9��[�D��a�ytd�GEA$�u����?ylI��M��Oh`8�_�I?Q��j��Wc6�PvbT��y�V���ڟ8��ȟ���ӟ��O�@DN�IN�B�,>��p�"�i����'D�'k��yB$x��.�9h����*zd�a�r�1o����O\�O1�@�z���Ʌ\Ҵ���
��s��+�b�%m_��/�p�(g�'&�x'�Ȕ'���'&@	�S�(�������q<&5�A�'���'�Q��3�#vU��ǟ �	h���9�%�;����W͞�J��?�R����䟸%�Tr�N�pr��0�
X=Qf�hS0?�a.��j�#��E�'�`����?�qA��/�`�( D� KQ����(L��?���?���?���)�O>����KI:���/]�U��!j�O
�lZ������ӟ�X�4���y��Q�q;�ab�'��oPJ�I�d-�y��'�"�'*쪤�iu�ɔ(tQ ۟����2-��33O�b�<肥6��<����?y���?����?�%��0�\tÈ]�}߾X�&O��$���yC ���	ğ�%?��	*�0:��	&*�a*"jZ?x8pa�OH��O�O1�������lZ-��ې4�٥��"h�Ҙ�&��(p�H��E��Mk�NyrH�D�vY��g�
'�F�N�X��?Q���?���|�-O��o�a�T�	�G*4�j�ɢ2���8�L�'�D扠�MS����>����?���j03P&/Hm��/ع�Jlȓ&�-�Ms�O~���AG:�����w�d��"K�Xj�4`���p��y˘'/��'cR�'���'Q�"Y30EP2%iP@�ѕ�huX��O���Ov�mS��S����4��0'�qЁ&	 h������B
ʲA�'O��'���'�F�b6�i&��O���Ɓ�"Q�~4XX������NU�	14!:�W��O<��?����?���7dh\�eG�i�B`C�6I � ���?�/OF�l�_s,��I��<��g�d��l��P� �#F�d��6���J}�'V��|ʟP�f	C�^��hV�
�0��� A�v00
^�c��i>�*0�'�Y%��H���a���ς�f2��Fʟ�	ӟ��I�b>i�'.6���, n	��m�1t�*�� Ϝ6���`�O���Ц��?�T���I�z��f�٧2o��r���5)������D��=�&����g�Π�2��I�X��[��]=>��!���Z"�zyr�'r�'�r�'�Q>����@'g+��b@�K�n8h�B@�M�΢�?���?a��d�}��.�D�̺$gK1`�a��K�2���O��O1�n���e��� �9Z(x7⑻w�H��ܨ�7Op`!v�_��?�q�-�Ŀ<�O��}(��[(q���s��r��4��M��$�����O �Jbm���E�k���� �#�	���d�O&�-���-�6mC̃I�*�۵G��	|����Ηk��x$?ѐ��'��\�	�|y�� Q��44M,��Si�#t4C䉹e&$�� �75���$�*|FB���#�M��R"�?I�oɛ��4Ｍ�T#�4qVb,����\��a8O��$�O:�d:K��6m4?᠄�2�z�S�-���8WeĎF�UD$��&M��$�X�'!џ��wF	hw@%��N�=�.����7?�7�iU�̳ �'f��'��� ��:�v���A
YB���k�O}��'�2�|����E�ȥ����?���� �#��$aT�i�Lʓ �������%�P�'�Ĝ��� G�z82g��1�t���k��ə��?��L��R���d���,�h�;�*��<� �i��O\H�'�r�'V2��*�xP�QHȰz�xI�&a�.��R�i��	�}�8�8��Ob4'?��]I�u{& �)I���4�}7�	w����&� }�^����1����V�۟�	ܟ,��4M����ODB7�1���M&�`�!Q�YĖA��E�\���O�D�O�I5D86M*?�&B�	djdQk3O�La̩��.ߓi���ƶ�@'�p�'��OX�؃$K��<��ڧ3�T�����Mc G�?����?a)�̹�G&O�;��x1���a��������O@���O��O��#�U#��w�i���2W�hh0b� lB$l���4�(d3�'b�'vP��	�8hR8��bCآYt>�A��'���'+"���O	���M"��
*�0��p�I�'ˌ삓ⅶ!�H�����?ٓ�ir�O�,�'#�,�$>�r���&H�M����4�\Y���'�0�;Ųi
�ɶ���ԟ˓\ʶ�4�ށ}V�b )E�2��Γ���O����OX���O`�d�|ʀ�I:
���Q�V�EI�qz��E"֛��V�:<��'������'�>7=����&���˄���;a�iwg�O��� ��IY�[�6-|���+K�I�buKt�њ$�Y�!l����+�2DS��;�$�<���?I�`s!��,B����M�[�Iq���?Y��?�,O,mڮ<�V��	䟈���$�*�O�D(���<�f�PE�5�ɢ����O���*��۰r@F|�4�MG��2r%�+��	��ٙE��ߦ9�L~
#��p�I7T�δPaK�%�NQE��P�8����L��ڟ���}�O�B�@",�!Đ>��=��d��8"�e�lu ���O��������?ͻ��} "ni���9enP�H�E��?����?��G���MK�OH�֦����c�G�С��|����nG�>x�'��Iޟ��I̟�����I�1��Ⴣ�xP��R&@]�-��,�'[�7͐� �����O��d-���O�x�DC+O�aB� [A�jH�uo�K}��'�r�|��t.΢��	ÅQ9������R7
��S�i�(�<�X�Aȿ�t%���'��|�Rٽ0(��#�-L�N(Hr�'OB�'4����4V��۴l� !��f=�P�-�(f�N��g�
o`��K��jٛ����v}R�'^��'�\�I��0 ����.@��&���"Yڛf����Z�Wj�i9������R��?h���X.�r�B�ya6O����O"�d�O����O��?%yq)P=��r��"8� ���,	ӟ�����rڴo!�'�?�źi��'�8���H�9~�ڱY1�W�7E��!�|2�'%�O��i��i���0N~�	����6NZ���UwB�	s�&�������O����O�$�9R(8��sტvn��r�P@���OV���i۹��'��Q>�Qb���@p���1�J�x6�:?!g]�p��ßt$��'�)��Y�����$<���Q�ё6���ݴt>�i>�1U�O�OH0S�"�F��z�́q)�0P O*�o��B%]8��ʕL
�j8@���$	K0e�I�p��4��'$���?�a�O�c��m���5ILPN£�?)��,�-:ش���2^�Z���OK�I)f�R5�ab�%&�l����v� �	Cy��'� j�J�6a�2X)��ߪ��;cM�O(��]�x��z��G��w)�Dӱ� d���I�0����'d��|��d:��:O�MaIE�0�6dK3Ɲ�r̐-!�1OPd�q��6�?y�,0��<,O
 BbL]�I�ܛ�D�� (�A{��'��7M
3(M����O�����0�a�舘 (@58,�=��D��O����OD�Ot!����*�Z�33��4�&E�����8gb��jJzlZ&��
Ԝ���4�K��$uI&�¡H������0D��
�j��$��I�1	�1Q%S��49{�X���?I4�io�O�Wg��82�O	t�JҌ�l���Ox��O��2édӄ�\�4�W��?������;�N�Yɾ���^�Ly��'��'~��'5bf� ����"D�IA�YF-OA\�	��M����2�?���?AI~Γ�^%I��߂cW
����M�y�@X����|&�b>Qr��(� &|qC�)4f�9�T�l�Б�SH�2b���d���+��'nĴ&��'
8��ގQ�,��h�-���@��'�r�'�����[��+��w=�I�RmR��>O�l*5f�f*��ɛ�MӋre�>���?1��$�R4a���Z���e"C�JI��i�(��Mk�O(%a�����ğ���w��QS&�N�I�������-�����'3��'P2�'�B�'��D���!X7��ĐBJA�w������O���Ob�mڛ&=��'.3���|B�L?��9�fgE�y���rt��2H��'r���鏔L�V��*�ˇ9T44+�Ë�Xv�ɡ௑�{E��O>�O���?���?���w�Q���Hvx�Ie�Bm�y���?�.OjM�I1d\˓�?A,��U�L88���0$p�ٛ򒟐r�On���OĒO�2B��L�f��D��SkK�8��%#�J0M�N�n����4��m:�'��'l����-(��Ѱxd0ӗ�'!��'�R�O��I��MKB�Jj �2�F��D�Bů��8L���?�%�i��O
��'q�/K�{T�<��b
A�eƟk�b�'�&���i���,Ϻ��"֟ ʓ$0>�XVM��-���:���|f�̓����O����O���O�D�|r��TPM��a	" kL�E�­Oś&��;)�2�'���'��6=��<�6'"�0ŶhaA6,�; �'�ɧ�O��PJԵi��8�hEX2hu�\h3��
zX��V��Ty��3S|�O��|j���]��kC��p�[�^���+��?��?/OƖ�@X��;�'���'m�u+ж n@��1,>�C���BG}r�'�R�|"�L+\HP� ��@�J��D����dA"3�J	{�jW/!�1�nS�$�F���C�b��+bP\�W�A������O�$�OJ��$ڧ�?��ňkVZ%#c&��Q��h��E(�?��i0s�',rk�����1nA*(i%��\X�4[C���_�H�򟌖'�~�)w�i��	�5BJ0�5�OD*0A�N��x<۴.�Zp��qdSA�RyB�'�R�'or�'!�@:c����N�� �PDCV�	4�M�b���?����?1O~���YZfe�1��"'Zx��m�?^�~�Y�U� ��l�S�'�dУR`�1k�<\�6���j�(j�k��z�E�,O�1��(D.�?Y�:��<�p@R!�4��"BOԞ�da��?����?����?ͧ��D���%�7��ğ���٧/�>(J��� ��(�7,w����4��'����?Q/O����IYL�.qPU�[�:FP�q�$K��6M+?A-��{f8�������s��5LN����:u��0f��<����?����?���?i�����MQP��\?|�Ka�M�\b�'��dv�d%
��<!'�iM�'� 	s�(ϊ3hraN[�͸Hb�yb�'m�	�8@nn~R=sz����
�u	t#�$w������韔�P�|�W���ğ8�Iן\i��L�'<��a��a[t9�Bh��	Xy�m�Ľ�b��<���	M�Jq��	Q��`&�9���F~�	(����O���߀�)Rm�)3��isF	�L$��Q��.3R�����4��<��,4L4r��qe���jAa	[z уu�]�|_P��F�S98<`Pd�0B��5�6�bP�cbOR��B��V�P� ���^#T����#�'�@䑠�20x� ��T�YM��ʐ� ғ�Dp'�Y�p�"�j�.�N)hf�S:�D��W� �>	�UϮ
j�\��kq*R�
�Y��̩ ~���'E�,��uIS�*j Lk#��ug�}q�l��<ł�gڛU.�"�E�m��l��JV'2h��)�d�/O��)�2ހ]��!V��E���E��w>����G�.!?8B K��xsg�>�)O��:���O�dDNu�r�3`)"��_�ڵ��B4���O��d�O,�J���*�2��M�R��#Daԅ�4F�:"�Ԛ��iQ��ğX%�$��ğ����Qt?�ԡ��67z���DV0���m�D}��'�B�'*�I�|��h�\����?����@��@E	`S�,l��$���I��\Y�LB�T�hUS�cU�?�\����RP��`m�����kyB�?|\���?����Tm<��y���x�liC�x"�'�dN)3�O��Y.܉��������Gh6�<��N�f�'\��'��Tż>��OQ�\���i����� y�Mm�۟�IJ�"��?��D, 7I�a20��0Lzq���&�M�e�:1�6�'X��'l��ʠ>�*O�I"�a��qj���w.؁Ȧ�1��a���O��Gǘ
l�7�I(w*T��Ť@
f�7�O��d�O8E����~}"_�t�Ic?�5���w�2!YA+ޞQ�b<�q����$���&QF�I����͟��>.����aL�P�"I֦q��7�O��[Y}2Z����~�i�1��ɻ@���z�*>S�29�Rλ>I�����?I,O<���O���<��N�~G*���.ٴ��)�&�.12D �AT��'�b�|B�'����j�����A�%������`�2 Z��|��'�R�'��	�v��ИO^&	Ka�;d���ĈS5Q����ߴ��$�O�O��O8�x���O8�[���=_�	�p��5 �r�K�d}��'�R�'S�I.El�髟����=w�Y3u�¶G����@L?`yl��$�,��l��H<�	���P�M����a�I6��O��D�<١�8U�O���5��	��!S@B9�	�&`�9�����O���<�9O�� d���e�	R���f��i"�� ��i>剸&�6�	�4n����H�� ��ğ�P�4�h<�!�7m��P����Ο�[O|2I~nZ�~�S3D����Q��a�7�Qk��l�ퟄ�	��8�����|r�#�=x���dY�8�J���,��`�6�'���'�ɧ�9O����h=2��� �d����ĸ2�do��	�P Vf�/���|����~� PI�vY��8W�P��'�M�����Y��3?���~��Ӥf��Q��0��-���ǭ�M��EQ�)OZ�O��O$5��E�?P����a�.�e
�	�[�	�!��b���	iy�'r\�i $�ﴑ�!��-8|�U�V	A�	ҟT�	q��?)�'�����.�?Q�Y�f۴X���4A*�<A����O��
�d�?�!�K��l5�٘3�L�<���p�H���OD⟐��Hy����M+$�ەΰ�#@Ț�G<���WH}��'��'��	
lP
�hJ|�v�ң-�𘸣�G�F�t��"�N"����'t�'�i>��I_��O�e�j��`� �R�qF�{����'LRS�Z��ۈ�ħ�?���S!%�,j�N|�qk��[��T��.�[�vy��'������u�
�7;6M�#�a�����Q+��D�O~M�6��O>���O4���l�ӺK���"sQ9N��Z$
��ʦe��by�����O�O�r1a��ͰS� tR��cШ��۴+�IC�i�R�'/��O�NO�	I��P
��>L���&cߌDm����	͟&���<9�\`�$� �	� 2ʵ0RdF�X�0�гi"�'G⏁f�|O�)�O��Iz�L�� ֹ&W|�k�꒧GX�6M�O�O�\��yR�'���'�L�)a�E1(�������#����R�s�H�D�v���$����%��r�8[�� C+W�J*09q�cE<�ē�?K>������O�����/t\9�')=|��Ѥ�G�%�ʓ�?����'W��Ob���&�(R���j��C�N5�i�.���O���O���<��n�%��	�!&dHbǒ���͛��Ò9q�	ҟl�	l�IRy�O_����4�$�����H'���3�O\�ħ<a�=���,��Ā5��I���Pq�eI����
��,od���?�,O8��d�xr��,q�x9 F.t��MN��M3����Ozp��m�|���?)��c2M؏l�N�4*���@U�A|�	�� �'=��������6Jƿl����b�>^����X�`�	�X
��	��h������`yZwiN�ZT&A;<����bK==Ml�@۴�?a/O���)�)N� �@��C	g)P�:�gY	m|�6c�BI�6�O���O�)T^�i>�ņ7.�|)6�X� ^��ȃ�M����?�����S��'��z��A5`�!tT
���*�6��O���O`���@W�i>��Ip?��#� �d����z٩F`KЦ��I]�ɝ��9Od���OB�<_�,�@H�U�~5i
�����lZӟ(������|R���'K���"�1	����&�n�A���x��'���՟��	���'&B��(���fc��f]��#���!�O��D�OD�O��Ӻ3T�D�B��/�*��8����!��jy��'���'��	%>x�!�O/���ՙ�Kf�H$�۴���O���?1���?�b�_�<�3ȃ&b*H<  �|����SnfR�I؟`��ɟ4�'��=��~*��b*)A��6:H�g��YtxT�b�iI�W����ן �I�V@�nyRa�.(g>h
 ��$o'�X&�8�6��O*�Ĥ<��O\�G��˟��	�?�� JL-D���3#H�)��dc#�;����O���O$h�a��t�'��i8K�e��tN��1��>��vY����$�3�Ms��?������T��ݰ:���*�1J�y��@�F�67��OX�� �wq���f��'�q�l��w�F",��ui%�F�F�<d��i0J�At�~����O>�����'��I�K�����V>�����%>��a۴a|������OxB��%
>ݪ�A���T�2��4_��6M�O,���O�}Y�K�W}�Q�8�I\?�eT�\�ݢ!I�->U�Ta��S����Iby2%���yʟP�d�Ot�DT}�� ��L�-ۢ�b��V2��n�ԟ���F[�����<Y����Ok�Q�Q��c�,��{pBL3��	�;�`�Cy��'�җ�d���:�^ŉOg�Y����3/â����>a+OD�D�<i���?��f(P@�ucېC� 1r:(����K�<q���?���?�����ď�k�P��'+,*�A�J2V��"Y�%�^�n�Ay��'�����8�����s�x� X���%&(�sc�Zڴ�ckD����OJ�D�O���e!`[?�I�%6��q��-nc6( ���7�Pb�4�?)-O^�d�O����	��|nZ+6� �����^��MbTl��6�O2���<Y��^�v]�����?U�bjT.��h���A��b�z%����d�O��D�O�Lc>O�˧�?��O�*:��D�{�|E��%��L�j52�4��C��in��0�	џ ��������e�E\S!ϓ��Jǽi���'�v�1�'��')q���)B"��`��T�XP�lp%�i�,eH��p�L�$�O^���B�'��I�*�+uJN�cD/�0r�H�޴\��������O�ҭ4� �<YF+I�]�:0�G昆p��bԲi�2�'�U
Xt\����O���%�^��L���аP�O^~�7-1��'s��?�������i�<��Gg1X��� ��G	Jo��,H叐��ē�?Q�������gH�
T�kb�W<]2��fk}"OҌ�yRX��	�&?�culM)g4̴�cnJv}�]���0V��tiN<����?aJ>���?��$��E߂T�1g�=��d+�)O4�N�P�����OJ���O`ʓ&�n@�78�Lm#�nļ -����&�t�0�x�']�'@�'Z%��'��Ȁ��]�`��G�uT
��q��>���?����F�8l'>�aD떷O5j����Ѳp�x�Vh��M������?��<V�S�{�J�ޘ��t!'g���&�U+�M��?�,O ��FZH��� ��
w�)�O߿R��5��F�i|.�N<a��?	 .F��?�O>��Ok$�+�l�/-ë�F��Qȸ�@ش���I�#Ѐn�����O�	�h~���iU�H��Y�w�\E��.J�M���?!���<�I>����������kD�'�԰	a円�M+��^;p��6�'m��'��!?�	�5D�8�mC�r���R$��{ҐY��4*z�Y�����OS��=r`t	���ϰ�x��Q!H�t7m�OZ�$�Ol�[�Gn�	ß\�	K?I���.r�r	)�NDSL"���$�(b/?�ħ�?���?)��C!V]�!��Vk��F��J����'�~ �T-�I�%��X�!���&�� 6|ВW��.=u,��=������O �� �	C�\e�.�/6/V]���	}���Vʊv��?9J>���?��@�?�2}aՠ��x�|��#ri�l�����Oj�d�O^˓uZ<b�6��<�"�Ϯ�:���ܥ=6���R�������%������(�"L��d@��q�	�S�����	��S����'I2�'��W�|�5�P�ħ_�yi񍏸&�&D����$�`ks�iL�U���	۟4������K���4���(
]���|LTH��4�?9����"8" �&>e�	�?�Qņ٪��X:"I V)�1�� �ē�?i�=��Γ�䓞���$(R�*�k׈��u��_��M�,O�)��l����:��^���V��'�|�!� �K!��+���!�&x�ٴ�?���|!��b�"�I2��0�ơ'*j��Ջ��L�d6m�O��d�O�	\L�͟�AU�`Hth���\�nz�k�CŊ�MX.\d�?�����'^����a�X�h*eM�hks�r��$�O��$�m>U&��Z���	)�T(᧞<�H�!qs�����}��Ο���L���/ap��Mf���g�5�M���k�^�b7�x�O�Q������@MMda�os6HO��d�<q���?����4���s�@�dI:�X�EȺk�Y��ҟ��I��'J��'��d�p�x;�z2oE�k�j�(�m͑��'���'��S�09Ї����N
%�@9AŃ�|V�Lɀ�M)O6��<���?���<Ix�'^�z�J�.3��.�;`�P�O0�$�O���<��nM��̟�z���/�0��m�C�@�
"f,�Ms����$�Ob���Oj��s>Ob˧3^�\���A����	C�D.�8�ir�'��I#&e��ۨ�0��O:�	�{"j]Y�d��u/��pW�L ��A�'*��'f��\��y"R�<�I|:�H�cAָ�[,6܌=a$a����'�膃iӎ���O����=էu���?th�h����'��ݺ`� �M����?駣��<\?��	C�'9��\u��6[��������IlZ�����޴�?���?	�'H���uy�R-u�Ґ�m��Jy�&H*E
6�ʻ
���O�ʓ��O!�*��C<ah�o��3�̌���O�f�6��O��d�Oҁx@}�_� ��S?��ᐭA��w-P@%�,Q���צ=�	��	!|J�)���?Q�C� ��e6H$��GD�B���K�iZ���pT��'a�P� �i�� ��/Zy���ܺxrpH8�O�>�aNZ�<�+O���O����<AR$
Y�q�m�8DJɒ򌙵6�R�P�Q�x�'�U�|��ԟ4��+I^��%�16����X�bR����/g��'�2�'�2�'8�.��p:��X#b��zF�X 6��PdK�WF��'���'��'��P�DɅCn�6��e�1��k	�<Mvl0�S�p����8��qy��Q�}���FlycOU�2�c�h�9e����h�˦)���h�?y�+�g�'	����D.bЪɨ�_`�n�ҟx�	��P�Ip��O�r�'-����8aH�隬n�`��c�r��O�$�<Q1�U��u��4	��%⠏M3b{th��Z��M���?�iP��?1��������׃Ei&�M{%S�A����w������	sy�� �O�OX�⡯w��&d>�@�ݴC����Ծi��'���Oo�O��;yT �6�KL�~�2�e��L�~�nڙ?\�p�?I�g��?	��p1L��#Y�l���!'����'z�'��p!��'��W>��	S?�q"ߎw: ;�G�'$�����f���M|���?��|;��7Ò�����߈R���肸i����8c��b�h��d�i�1�@�yF��r��Ⱦ#����Ac�>���z̓�?����?�/O�y� �� Q�����BW�~�&u��lOn&�O���9���O����i���0��$-�����^*F�E�@���O���O<ʓ3V=#9�NġRb�7^���O��X����x2�'(�'�"�'g��O��������4`Q�V��P�U�����������I�^�DP�O�"c�&}G
�*�gR�h���#�L�0֪7��OڒO���<Q�g�IY\�K�ѿk�t���5m�7-�O��ļ<�"��,Zl�O�"�OL�T;���"in4�u�_&��t��w���lK��$§�n�� �!�נQJ�-���H�z�Z7-�O�dG�Y���$�O�D�O��i�O�����m �D�!YT���Y%YF�ȳ�iA2[�4�U�!�S��<J\���J,O�QSRDԴ$R�7��/8��\mZş�Iԟ��sy'�L�I�\2� F�\�
�6S�H� �ٴG#��Gx��	�O6(I�}Ӕ�S��Ŭdrd���Z�M����I�A��0�}�'<��?��M;��� �d
�d߱Oz����D�O6�D�O��rǺ#��U�S��> ��1��������'\���}��'Vɧ5�mU�G_欛�D;rubL�` � ����Os1Oj���O`�D�<iP
mn��+���/'�2���1w�������Ob�O|���O���t� �=��2�)ԜH>
� M%~?qO��j�]�#r�88v/ڝv�:��J�\�e�bF��$=����f�����H�J��t�
O�T@$�X��&��q䇢_�c$���.s�%��C D��@XĩT�*,<AHr&~5HIP�=A�f��$�˷/5t��$��=f7�`�D�T-B�[�ո{~"h�5d+u��%���ƭM�=���#R_~�����3H���Z�J�m�06� �#+Lo���̚CX��DJ$x�.�1UGGn|6<+s�R<\� ��!"����^vܛ3�Jo�Z\�	����A�'=�|���=��⡂�?�	�|��σe<Hv!��$�� �!�W]��3G $Q 3�Z'�tx�g���<���X�1�Ô��rр�Ja���a*�'����?���I�O�@I4�|�``h #l3���aB0D�48aX cv���Po�S�ؽJr�/O��Dz��-.��82��!_F��6j�+	�<ꓨ?�|�&�� %�?����?A�Ӽ�qJ�j��`8a�@"�$ɂVHɧ+�$8���@�$q����\�H��L>��	��<)Xa��̎��иY��	�����X����Q�D��}&����Ɲ�pw��G��
�
8�p��� �'p��|�����^����I O`���%@��W�!��F*:x� ����U3��QD��@��ɏ�HO�Sky�"6�hADR.�D��s:>�f� ��ߴTB�'}B�'#6�]џ��I�|wF�hz���� ̰|� �M�v����E��'x)X����'���J��!U�l	s�G��$d��(p_�*F�ң���<SbV�����!�B1#��8�HT�'�R��D�� iX�P���6�`�m_|�ȓ<~V�[r슟��y0� �7<A�<��U���'jVᒲ�{�����On�R�+s	����a��*�����O�特U���O:�ӜDeݴ��V�4*W��>����CϬ ϊ-�㉈;�2� �p׃� �H�E�?aH���V%<O,@ �'��'m�D#�
W���]R�L��K���'��8�l�36J`��&3w0T@�'E|7-T"rn=�2��7�h��Ōt;�1OJٙ��TϦ����t�O;��[�Y�� �+�|���ҭ�2	�4����?AW̐��?��y*��I�F� �ЂCP�c@6�rvB�%%d�'�^�s���I��z��CF��kw`�0l@�7%�Y��,��C�S�'f�&��V2<�\��l��I����΂8k�M�	 ݠa�Qd�z)�`��$�HO��a熻�`�C�k�*g+9�,�����	� ��>x�Rm+w�Nϟ���П���� O�׸�h�jȤ"��!�c�`��XI��I&<�|pE>?6�1��Z�/����+-<Ojl��ր��P�AE<�ĭ���'�>�����|��9SA�4���Y�4e4 �����y�I��o��"�dY�1�^�1���$M����0�tɓ�h8��"��NA���)�8�ᇦ�O�d�O�������?Y�O�x�2���uix����TH0��A���x�G#\�B6�W�ND�)���tO�x�'T��c�U�@
�(S4l��7�T�JD)��?Y�:b8l�(���, +����tS��H��R;,��՚����
�D(�	+��'��:�tӐ���O�A:F�M�8U�Q�@�Z$���8��O���t�����O�� 9R��;���;�b�y�bP���$��;F�xА��'�����D�j���6���v�Ǔ=>��Iy�)� �:��k���iT튕 ��4 W"Ot|�d��P���GG�o�*Mz�O��lZ�-d�:c��_��I�˅�3xdc��S�#  �M���?	ɟ�=���'�6���C\�X=�52e�:��'Knh���T>�+�< �E�)Apb��.I�6i�O�����)�^}̠#7M�;f� !�<G�.�'��9�����O-�@k ��7�{�T�U��݉�'"1��k[- M���E	R=|���ɲ�HO�m3��8"�8�^��ȹ��im�ҟ�I���9.q"(��ן,�	�<�]�������'
��a��+�� �<Y�%yx��a��J��M6�+4���
��(�ɋb������I&(�:U�΂B�q@C�� %c�l`Cd�Oq��'Ġ���z�6�yAH[6&2�r�'�e�UjJ�d=1��'(l�$��O�4Ez��ӫg��TkC�I��Y(w�1S�@��f��4-0����OB�v�P�;�?1����$*��u��9(���#�D]
�k� l�t�{�'��A҄�k$p-��2򄺑D>�x��2cnh�NQ�3	.����8+����?�5��F|]�q��'==�X;ub�w�<Q�����ݛE�I�r<z8Kt�Ar�ñO��	��Ц	�	ן�06`�j@�U��B*^=ʱ�Sޟ�̓k/��I�d�'I/F���^�ɋ�t�Q���X*��1�9��L�O�$«Qs�d)���ʠ3v$��'6�����Fv� ��8G^���D5T��ȓ"ؙ5�Ɣ1��X[f9��]蛶�/l��9�/�`�HB����'�
��3bp���D�O��B�ք�	���H��Jj�^(q�NF"(E�H��ٟ�Dh�˟ �<���d� nZP<���X�(�=�&� %e��\��Fx�����mζdh�$�T{����%���3���d*�)��p��h�/��P��p�vB�"�C�I��6����s�քq@Ks����w�'T��8�U '2��ȓ��//*�Yf��>1���?Q���(Za����?���?�;p�@�q`ړR
t�E��%Us�MrԨ�%%k~��2c_D����լ���n��l�u��4_�v�`�Bϐؖݚe�H'gKɛw��&x*�`r��e�g�	8+I��0�\2dob�*���_���	o~"����SK�'� E� N��ad�,�(�;���H�'�J I��(`P��bFhG1����O^�Dzʟ��~i��G�J�,�[��\�a8�}C��mx� ���?y���y��>���O��ӝ>D"�BC�Yb�-%�ɗ�F��,�X[!�1��h�1�� 5�F�G
ă�VC��3�r|�B��p 6��2j��Ȭ���O���]a�Nu	 b�yR]��MP!�!��R��K�i��lc&�)!��Q�1O��>��Ƈ7�F�'�R�G���i���4X�%�o�98�:O��E�'��5�4|��'�'fT�;ӏ��-� |�mɏz�P;
ǓenH�?�E���x���a�� B���Y Q8�H��O�O���G��Q�XM����ae��b"O(]���	�Z�h+f�Ȝ+2!уO֠mZ�Jǈm�U�eĠ�Qԏ��>c�8Ycm>�M���?Y˟��4�' =�
�PdņO�H0@�'��g2�T>���tbBF�,Y�g����O<pjv�)��(Zא}Z3F�yI��'ɩF��'�����ט��Oa�i��o�q m��RD��C
�'��C�� � ����:_XX
Ó1Q��L�$�,j��h��@�8x/p���I��M���?q�eA,�T���?����?ў��%V6�8�kā�Tt ����'���*ϓ��	xU�?]��z�h[<)����=yF��Mx�����M�'g<���ҒpZD
c
�[�tZT�)�3�$�5B�`����,���Ȳi�B�e����FW8vH�2r��c~����"|ҥ&��+�Vy�(������"��d�d���?q��?ɞ'��OH�Ds>��F R��۷�M�[�B�	��� ,,C�ɑeX�	����Z�FW.\ht�"-�xI�#vj���C�	j���R�9#��'�O� >0�g
'q��p%�5(	V"Oxt�v2���c�I&)�J�rV�$�Y�s���u�i���'0�'�����
�k��Z؂t��'��ɗ �"�' �iӟ.��|B$X�LJ犈7��R�狱�p<A¯�r��D0�	 ����sA'����I1b�~��.��7NuY�c-����膶�!�$�� �|�g��6!�H��!��]Ȧ�0 i�.�������oR(( �M;�ɧZ�� (�4�?1���im!��i���c��*���*�Aԇ0���'F\��'1O�3?)� /L����ߧN���NY�ͤyi��?-i e�	,+J�P7e'b��c�.*}����?Q�y��t�@���	5w5��rr[&�y".J�. �$+ 	B�M`ْ�K�0<�W�	3s��A�V�؀�:�+��K�}J�9;۴�?���?�W*�$faJ�����?���y�;g\��!؛f&���A�g�*�y�(L���<y����Q��%�R?E�吲b�Zܓt�؄�	��Ѣ��j�� ��ȋ�x�<9���ʟ�>�O�I�6�:T�L��2�,�m�A"O"���蓽fOZ�ꗄ��4zUˣ��Hy���ӘP��H ���V��DJ#`�h3 �|��I֟t���<)\w)2�'��)��.\�	Fau��8����7�R�"dO�ah5	ʚg>< ܃*��5A��K�!��ʛ��,+A�	�\%�*�� ��'����^�"�F��ІI�h�.T�F���y���T��t��Y�y�梊��'�`b��,��M+��?c�N�ZG���Sf�P��Ǥ	�?)�'L�$8��?��O �����i�����4�DeC� �H~����:B���n\�~�-h�"Tk���{G
0O�	{��'<�'mjp��A�,	hxma�dT�oF����'-�i�t�ХC�`����%e̠}3�'�b6��&�pe	4Ɔ�o���:�꒸Ov1O���U��ئQ���d�Oe�ة��uv�QAp�G�0�а��%C�0K��	��?�#�  �?�y*���� d�P�Y9<?҉c֦� ���'?�2�����{VH���L�z�hDB/U�
{�6����	k�S��x
8# ����s˅#D�u�ȓ4j$4����.�uɄ �$���I�HOx���_�bi+%�T�.�Jy���G������P��1�8��GeI���	�����iBB�$h�ڹ���N�J��Si \̓mђ ��	=�R�j4BMp���!�V GO���i��,<ORd��(��G�n����/y,]1��%�I.{, ���|B��9��σ,NZ\��eH��y2�\/��:�INJ�trՄ����dLc���.��F/YU��b�I�;@���T����m�W��O|�d�O��	�c��?�O���
�3��8����F8z!
3���xb�" �
d
d�R&����h��1t� 	�'�d�7��*f� ��_���:����	q����G'��@f��w��r�X�a�/?D��H2`I!_�Ā�n-%2�r@'�ɽ��'BXpiU�d�D���O<��%� \6:xç&�s,�Q&��O��I�j����O\�ӱkZ��d;�䆔��ᑷ U*<Y�Ԁ��x��-��'��l@�M�B�ʕ뱁.3�L�rǓ^0
��	D�&䂉	T�=�l��,X&�fC�3*S$!��`�$(��m`q7�B�I��M;&��.
7��H��]S̓W"]X��i���'���M���_�g��5���H�Zւ!��A��'<��D�O�HѦ��Ofb��g~R��H p("
A`n`5ò����"<���EZV?�d���7HL¶��`��^0o����,A�D�R�ݍ2>N�C�`/U!���E̔����j��"�9haxR�)ғqH��I���c����ĝ��	��i�2�'�"BБ1�/l���O��Df��.�WG�504O������K�xD c����$'<O�Ep`S�+Eb�S5�P$!^\���ړ&K�y���1r,+�E[��h�A-�!D�1O�x����������:A(�8"����L��S�? r��#�-d�����!��d�8՞�ؠ���"Ra����(Ӫ�f��"ۛz��1�Å��\2��	럀�	�<�Yw�b�'@���Ӫs�i<L�Z�{a��d'&4BvO$�1���J�6lՁb�q��$^�Z�!�D���-�������F�*3�~����'!���8��ʥ��m/YI���y��"d�i�<њ%�(����<a����%x؜0lZȟP���K���2��&�������>��$��꟰`T��ʟt�I�|�j�r$%��ㄠ�(3�t��$H̜{��3��,O@H���ߺ�'����R�у<� RCY�+�<�j
�Gz������蟬Y'돇S�������Y>�p��'9���SJN�[&��,;^���&C7^>B����MC�O�6DxK&�ZZ��ER"��<�(O��Q�����	ݟ��OT�q �'�Nh�.�� �L={2,T�j�J���'��/����T>�a}��DKw�1yƤ�6'�O����)��Y=�A�v���E��t"�O1P��'��������O\�1��%"2�y�qEJ�5zXh�'� (����b
��`��X�L�Ó{�����j�G4��Y�aVZ��6D�l�ֈƳ=�h����'61qC5D���!� 6������_���q��>D��t�_��r �a�˻w���#3( D��0#͒UÔ�@{8��g-�)�!���5wF4����*�t(��,ǇQ!�DA� �`�z�L݋B�f�VJU=�!��JnN�Ag��/��ӓ��<�!�dJ��TlJ�B�9�8�"O"�:S�<�,@s�Ω/�\��"O��hg�]/�\����;"�|��q"Opy3Ň�����c(?P@��3"ON4*�D�K@���p,��gL���"O�tpc��>2���ؕ�+�z͊g"O΄��l^Sx�C7�F?g�-)�"O��J1�\��)zE�ݼVH>��G"O$hh,�b08�q7��_th�"O�q	�D�CD�\#7��l�Zm��"Oj��t� 6ŘqH� ��l
��w"O�Qy��?:I6pbD��[���e"Od�*&k
Q�Q�׀��B�"O�m�5eƳ<Jj(\�}Y�=�q"O��@
�H
.�����$ES\$�%"O�x��7@,Xre��O9fH�"O@@c��mf�9�D*I���`"OR51�JۻjI��R��Ѯg �ŢG"OdIw�?��e2� �jh`�q"O�KE✽�Š�Oh����"OH���,,����&:=h�m D�,��ނw�̍�6�؈n�~�c@�$D��Z&m��3}:��0H�V�l01sN8D��C�-I&==7/['^�*����Gs�<A�ϝ� ������(:�t5�wLy�<��j@��Dtr�L^-H�4}�!&�@�<�
�~ABx�a��$\�U����|�<qS.�y�(Kǡ/��Ͳ%��x�<�g�?0��tm�m���Gs�<���ش�x�i��bVipLl�<�J�<sZh��䝹9Lq�rlHg�<�E�U�����F������Ec�<�p�>x�rG肳& B��v�<YǬ�gw���шC� ����h�<��"�#/
d�HQdѫK���&�g�<�b���-��l�R�L6Ak�<	��S�r�n��'� =צ�y�l�a�<ٗBݮ'e��T���zu���]�<� �d"w����F�(�,�?Z�u�c"O���5�?lc��h��\��(S�"O��CBN=�PO	
	����g"Ox��u��:}r�����t�m�a"O�B���(4�q,G�J���D"O�i��i؏=�-ca�G�B��M�"OX+� ^����b$c�Z�l`qe"O֐bN 1lM���4GeH�U"O�Ґ��
 �2!T8(a4	��"Ob�j�%�$r
v�rq��:%D2�r"Ox%�6�:�d�;�b+C;�<��"O����N�t�|lSa�_�3T΁k�"O��y2�
��MQ�"�Z:���"O
ӃB�<gĸ����J�m7V���"O�q넃L�.�tY���Χ3S��0"O��9�֍o�ňd��K>��"O1�g0 ���(S�H
=p��"Od���݆cq����x��qw"OT�6E�Z�d�#��.���Y�"ODY*����v���+��4�f5{��'�v;BH��F�����kՔ�B9F)����!ӥg-4��j��
�H�4d�.R�D��&+ړ(�����,�/	Qbb?{3��>K� �0�A�O�%��-*D�(  ��
a4�2f��R�m�`b�O�@�F.g��P�H�"~��o���|i+&bͨe��!�U�ԏ�y��\�R�e�P[�^����������FU|�:Aӹ��<�1$��&"���BL�*(�� (��K�9(�}���E	��غl�܁"T$��y�6�0�!�8���ē�����-��5b�/:����I�o�� �R�x2���?�'nC~Y�DnYV�85R��^�H&Pm��I!T���R���C� p����P�V��ъp�y�(A���[�S�O�P��`�ղ`�(4�Hf�����B\���#~B%�$4p��5D
�@Um���K�Z��H@���ä�J����N���	�+@�·`*n��U�n���tP�D@-��'�dp�'<�����Nz`�8�EE5o�� E�8�z4;��ݛzz r�'rѴB�	sn$��b���q^����#�<���pgFC�+�xX��9>�R�E�/3�$����Oq��+����8�P�"V+��p��at�'���
!"]+�򤔖]唠P��<:�Ċw��2Jh�QF
@�|ɧ�'�Ȱ(�iY���	zFi����>N��&A�n{�DӠ��9�0�}�D�Ј<q�[E��@�&r�����l���ѝ�
�`R g�xI*��6O*Ȃ�+��K �v��4|�m���.l��c�LY=�����/� IKǯϴ5�*ɀ��>�f 0`GR�*H;U�J%m7P���'r͒�H�
M�Р�	��/X�	 g�=T��-z����0A��D�(�?%?����'��t���F#؝��P���=!��܋%��ɀ\�f����R�$/�h@A�,-����cj?y5�'fh�ߟ���&y݉jD�>A��ثlϪA�E�-N^} w��x���~|[��ًOdn]����7J`1����~2V���"ˊ9Hl��I_ )�#k~�������&�0<��aYsgN�jWEn౫�#^�	��qO>��+N�M���3s���P.���'p��[�� �D�B�́u$�$��\�%��	No���#hg��H��=�CU.'&�9�򎛨 v>X2��A4%2qaU���b�T�'E�	�C���@�.��d��S�D1g�zXhg@/�O��W�Cy}rI�N�~D�q�S,|��d�g��8VWtq�.Op�ʑ���#���B�[�r����\Y�IK��%�G��,yE��B�
m"���IH����"((+Nv$;��
F����Ƽr�$��v�N�3J:�cB�ѳJ�~�)�B�	-�9�O�u�tk.�B��M���=AG��ghݿR��⟬�S��2unИp��B	��Ȋe���������Q����D-_U�f��D�Im}���'n�az2�O���kq�Z+n��J M���sT���VG.���`אd�߻I��Ɂ+-�ʧ[�$1�ES0A�]:T���a(�x��M�Py.�� ����U��$����@ ݳ'H9+�^DX����G�_tIn�Ѓ�m>-�3�i���;,�J0) ����#�*q"��*TO0�(G�p���{�hC�G�d�p@i�/L��1�T�3E�%y�DF(G���ش](����)�f0�c�:3�*�9�B�j��<��/x�F�Z���vNQ���-s��$�g��N��1�B�}��ya�X�?��,*<���$�J�P���ޝ}W��犛%a����[;>E���+��P�
Wڢ�ͧ�LQ�w>� NpZ@+H���5q"Ō?��"O ��2#٨(�bH[���/p6�H�H�H����&���N��k
�$9�Ȳ�?�	� 1󮌔gm�t�S N�XM��`�!𤔤����7�כ%O\���Ϙ*�ju�ӈC�t������'+~,��j�c�'�\y5��3��Փ�)�Ě��Óy0��c��,19#� ?�?	����Y�A�\�P�|HCCYc?������dv���.g�H@լG/+\��OD��6�A�>����5����S���0u7�$! '�!�0��V�~N]�"O��;��T�6��y
�)�f`
��ѣЉS��ThW�� ï^�wo�b>7�^�����\��@��=_lZ�B$'x�<!HL 7A���p���2(��S1b@Dq��i���d��$��9Ҭ�E�c���>
az����fMt����?�����U��x��] ��A�F�<�r�Ty(��I�
�pɤ�A̓o�Hqʢ�1�������c��ݛglɕQ?�e��"O�q�҄p���0�ՃK��*�7m�(�O��)��3?�����
m�tZ�@�/s_�e��
�C�<i��E	n��a���	Rh	�&iܕ���&�O� XV��
�@QP��YIdԸ��'���<�6��;g/�B� (�B�j���O�<aɚ�p.xhc�����"P�M�<���U��,h��cL<tʣ+�G�<��v�-�2�
�P����#�\�<e+8F�������<�#�ZX�<��OU�m�G:
�\�#c�x�<	��T-@��"�˭#~��7�Bx�<�����oz���>?������NK�<A�\�*4@�+G$� T��Ļ��k�<�`�K�z���ѩ�2RF�LS�i�<�R.�,��t��T��8{0p�<Q��Q&f���"��h�h�d��m�<񢥃�G���h���UޡӂgN�<QY��jeSk&F�@�G��o�<�`�B�[vh*�/M�oc�4Kd��v�<�G)E�J�"h�@�,�0����n�<�Λ� ������V�O	p�"��Yh�<��w��Q�K.����c�<��,��D��h�i~B=��R{�<y��̑
wҩ�g��R�։p�&��<�ueM�z�([K���i� �y�<As�ا|�r��c�j� �	��Z�<�W�����"珂p(��T�M�<�'�#L�{7Qw"�Č�I�<��`M�G�$�n�*�)`w��B�'��U`,�'@��%бB]�1i5"�l�6Y$bH��FD�#���T��sM6I"T@c�d�8v�p��=E��Jhb��W�Ko6�Q��J.ia��?��-M�V&,�D�$́�k4T{w�ޥ?����4�~"�۹/�>݅�	
e&y�GLW3;��Ƞ��ȌL$���B�~�d�O��>q��dG$�����ċ��N�MBr��F �M�!�U.ܩ���z1$Q�u��?c�R���Ly���S�8kG*��ا�I����R�(�[92��".��x��{#(�"���=O�큇� Ya��"��[� ģu"O���C�F�t �꒩ �,�PP�D�'����'�'��Q3�)����C��Ԅ�C��ۃ� �e[���d�-���Q���9� &��E��'����fD/1��ᤑ7N��4��'զ}���x
�a醅'Xi؛'F<����Q�0>ɅM?5)�8���O�x־���c�<Y���V �iэU�9���e�<���~jB���[�A!p� W�<��%EQ�h���	y�b��Nx�<9�˱$��+�?��rfD�<��	�p}<5��� [�\��&B~�<� dU���K�3��{gg^�IА"O��0�G�Z%&1���J�L.�h�s"O���i9b3��'H-=r��K�"O��p j�g��!�FH8|�:C"O�`��� �!��1 �E�<sk�Ia�"Ov$#d/۸p:��O�V,��"O���@�h��T;��'�H1�c"O�ysր)m����5V+ �̩��"O����^4���Z����f�>7�:D���{�L�(��ya ����9D��J)�y�\=xGꙮ1�⌀�	6D��;�G>������D ����h5D��	�A;@���Qn�;����d�2D�(���Ȣ6t@�c�U����0W!-T�L�kL
��C��U6"O ����-a�2 Hw�[�1"O�1sd�ײkۖŢw�Z�.X�I�"O���U ΍�N H g{kd�t�U"Or|)���H ���U��,�"OT�ؓ�̾=;h����?;~EY�"Ou��[��i�l%a��;�"O,�Y�jF.4�����j��i˔��"Od59��ڹ6�h�#H�&��"OP�y���E|��;H� ��"O���QgÜ0ybmy�	��h��"O��	'̒T��z2��y����E"O�xƕ�f��(GFHl�03�"O���@U�v���[�kܒ?]���"OP���Jv�$D	�Ɉ�uY ��"O^��ôb�[�n��$�RI��"O�`��:�6���29�B`"OPf��6����A抰 l݈�"O�����9,������%�%�q"O�X24�@�vLl�ʧ"ݴB�����"Op���Hк���S�	E�0�"O|;�!T0A�ϗD)�ə3"O� �Q��HDnX;/���K�"O�Բr�X�e�|(0�΀Qf!!"O��腨޳0[蠩 �+=�Ѹ�"O��*\c�RYa/Y�B80�B�"O��*�Kڞq�� Ch-!G����"O\�ʶ�V(6
]j���C`��3"OU��J�'d�2��ĉ�::~i`�"O(���ER6>� �e�э(8�i�"O���EK�=��i˅(_y#���Q"O��S��^ J�x��G��{����"O`&LH�H�B� ��e�5 �"OD�rV�F�C�H'��0N� Qv"O�������f��2BH N�u�w"O�e�$ň).&^I���86�01"OR,�v.B-$�<;�)hc %8�"OHY�Њ;8��,H!�<\X��E"O�LS��Q��<����c��|k�"Ozl�oI<�J]��)܇S�<�c�"O�=��lڐH�4���G�	M� Dz'"O4H��l�9,F|P�7	��F��� E"O��H�iJǮH�����lsu"O���a�/IE$����('�p�"O�d�D��'^l�"�.P�t��G"O�8�܅9&`sQH�6wR�#a"O��Y@��"=�|S�'�'Ze���"OH]�JK:HrX 5c�A�"O"��w�/`��bFD�@P ��E"O���2'�6WW�`sW+�*tc��$"O� b,��h��[�l%�@��
"yŐ�"O���s��ZX*�u�X�8B��"Oz�9"M\�3$���K�A
���4"Ov`X��5��تp'�(u��z�"O����O�[�9�`�߂[^�Z��Ik���IA�&�ΰ��A�JVAP"d ��!�$�w��U8@&A6666!K)��C��x���]��I��J�(�FC��S�V$:�)�	e���Έ�RF&C䉡9����N�P�,�fD�,d�C�	n�����%8�p���}��C�I�x�H��F�>v^U
��85��B䉀[��v�XeL^EzA�\�C�ɽ$��T��� �86G4j3N(D���'�VN�����%l�f��pj:D���J	,����S�@�tA:D��b�PIV�!6/A���C7D�,��b��=w��!�)ԴҔ�[�e(D�D��Ӆ�Hth�E�;�p\�F!1D��F�\�L�y��U�<Ik0D�|�K�F�qƄ��ZN`8� o*D���BJ�
h� (+���~$���"D���W%1�^�xQƗ�o�V����?D��`���6t�����S� �K8D�pS��
8�$܁�`�6e1��4D�@����4�B� R���j�6�<D��ؐ�H=w2�2����(�M<D�����4.�\�rG��w9��"%�8D� *Cw5,�pA��}f��ha�)D�$�RAǳl����)�5X~�H��,D��IvjK!T&¬�Q�d��F�)D�˗��?�ȴc���u�,i1%"D�Р�+��x���@��v����a�HbD�5�Obٲ���j��Y�Vn%LR$���'�(��O<]� �E��v,��k�$Z3�BU"O\�sB��m?�00�Ƕ(#lZ�	q������? �>�SG�?9���q��6�!��u��u����#QI�p�Յ[�qV�Ҍ��*�g}r�V�p���N�:���&��yҭ�8y�Ҵ�����4T[����?�d�'C��P�I��|���0�U>��	�	�9���`��#��Ą :0��%��'�ИF�N�L(!��n�m�0BŜ�X;�g�#qO~���IH�S�=F�v0��,A�L�J1�O<t.0B�	��L��S5-�+��w�-J��LS�'c�"}�'�6����
�<s�Tـ�FJ� �'m0� S�6�^�����|��H�'0ģ媑�<�Τ�4��=�ޅ�
�'�Ƅ��Ώ:]�:M��DF,6�@�
�'��b�I����)p�E�4S��
�'Cf=P��ְ6v�;�%D�(~΁I
�' hk��Y�,�h�-� &��p��'*�`b���_�V����.���*�'8��㬅�|-`�Ē���!�'i�@7�=��*C��Ů��'�z�J#��!�AP�	�(H��h��'�`�����;��A���Q �h�'���x6���(a�e�HG�'C�c�'%�lKwA<��U�"d��+]$���'�v�Q�MQ;"=C�H;��M�	�'�nT�ei�����)��8��I	�'��D���7܂`�-��Xx2�b�'���@2�ڂMd�=�Ţ�)I@.�H�'׺�PM��}B����E ������ �@a#�/f����`@_�6D��"O�a��^�R�R����an~�S�'��䁾s����%-��6 ���w�!�$+"z��(����n�C�Ŵ:�!�j��0{��J-B��fN�[!�䘆f�H��#�%c���@�7�!�Ĝ<]@�isȔ�F�(@ׇn�!��K�І� ��W�8���Ӈ�@�!��_fgp�k�a�T0�L�!��Q�tm�q{��$�P�B�@��^^!�O�&���㤊8��V@�iN!�$ջi&d����	l 8M��.։.�!���X:����U."��ݳ!#��!�$��!
r���cY�>������j�<	��]�ņQ��`D�B,h�i�]�<yP+�J�B-+bl]U��Ej�b�P�<�&�ީR`	����'��Tha��u�<i�ȝ�>w`p��ȝ�k�4�b�^f�<�a��CK"�s�%�>b���c�KZ�<�"�Ь;�p�2�mW�y�����j�<��Èe�05�/rD���m�<�d���B����ũ���x`$^�<Y��(w�D���kؚ#:���D VQ�<����8��p�v��s���*"%�s�<i���-iORlY��Y�X�Z�hr�<�q�C
uz�p雿>�Hh��m�<w�׃/'^=�_829�Q8G�p�<����;t4��R1�ڱaN��!%Ph�<1vMCzUȉ�㆑�p�ɳcBy�<1���@ѪaR6oR�ʐR��-S�!򄚟W���;�/K"΁��ŽR�!�$	̸�$��[W��B��@�q�!򤄹�đh���c�}�SL�9�!��$�l1(K'��œ3���97!�U�~,�"g
'��A��Ś�!�$B�b�V-3E	
�Ap&%6!����&��"͗�ܨʢχ0�!�$ֺt����E��(
��X�1�!�YL������R5ذ(V=|!�d< >�C��U�V#l���酟/!�$'5� ����!6@��B�,=s!��Bw�D]B�fΒC~��s�\*S!��'j�ι��!P����0u���1�!���5hb�B`�"If,Wޅ^�!�D�;fA�X4�L:jt�B�1�!�ԭl��H
�kېo��ƄW� �!�/C���poŀ5��,h���(K�!�DZ�(E�b�|ƨ�CШĐ'�!��%���7��1m�l%���1�!�D/.X�{��ޙ#��	:d�L�8�!�C����0� -�j͂�� 
"�!�dGB7Lp	�Z`T|�"�f�!�Y!l��c��\3s�@�����yB�[� - 2O�+|��Y�8C5�3D�,I�HI®� ��)m`�2#2D��ՉW#��te�I�O����*D�����
}����ԭ'$\u�P�+D�����%��H��k�N�*�rf�(D�\s#Ο<7�h`Ğ)	���d�3D�@c:V:�k aR,`9�(���&D��I#b�ZG�9�7j
�^�4�4F%D�$�@ԾD X�' I�/�ES�#D��2�慐OXf�;�Ǟ;k�\s�n?D��� �Lʜ���E&B
�L���<D�� <hzGD�>d�Ɖ{��$^jň "O�U�rF!�b��V���Q��D"OX
A��r&�|;��\�c���1"O��/A%�*���۸J5r�p"O����`U-W���x J�F�ȕ"Oe���H��`˱c�6i Ā�v"Ot������H��U�����yGJ��f�)M��aբOhC�	�)����GƃV��4A"$��8C�I�Fn��hPJ*�� �����4C�	B`�C�
=��"� ��B䉐nb���� i�y����B�ɟd��CqC�8s���/]5c]�C�I��8��G��e����&5k�C�`&�%�"N����゜� :XB�yӑ�Q��x(�sb+Y4rB䉌n�xKrl�~X 1�W膐N�NB�I�{�f�k`��9Y9܌ʅj��?^BB�I����.���"R��Y\�B�IK�"�0H�]Vb�s��X�_q�C�	U/�8�լ*��*riV1g�bC�JYFr1�B6FegI \J(C�	�I���[D�c�N�5�U)|C�1�)Xw.2q�v�Qr�F�B�I�D��ͳ�!	~x�4$BSB�B�0D$d�D��lϢ=���A�X��C�	�N*bP��M֭zw�9�5	Z"	�C�	�	��pƆ�q����Df�%w��C�/
�NH�6e��DrΠ�P`�-AafC��t�&�� ��U�,�J)�C�I3�`�:u��#�TY�Ȉ�2+�B��!Pb�S	��,K�DF�j6(C�K� ����W�:#ĩg��B�I�f+��-ֆ��=p#DجB�5#��Ph�EU�˪P� +8cn�B�I�"6��`IȨ?h�\#e".B�I7)0����0�N���+(B䉒[)hB�ۉ"u�X�@�,��C�I>wsְ����7�0�J��_�22�B�ɯJ[�p��!��e��h�M�pC�I$R���V��0#C�u0���:%�xB�ɯ�D�2 �Gd� ��=~)�C�I�j��E�%Z'v�N
ԌB��C�I	���a�� LDU�5@Ԋ(�HC�?mm��)��66���&MR?�B��u��ĐT��@����R��1\�B�I.Z�hpC�oU�(�	caE+Q�B�	MF>�#�BAB R�(�ȅ�z��B�ɚ!�<�Í�c4|�Q
3q��B�Ɇn[�)WH�~xN� ��^�7�vB�	�,4��k�Q�S�D��X�h�lB�"
za��� >mn���4B�6B��.�	h��t;X�S���?C B�.C�^qb��>1�	�A`�C�I9��Z6/��Y�B�+��x�C�ɩRRJ���C�u�Xp��ܵI �򄎥]z�d�!�tL�F�<�!���7�I"`j�&,��@�C;�!�����*�A��0!;��Y�y�!�U�g�MѢ��`����3i\�!�)o��c�H������蟣$�!�d�8Dp���(�"�� 3e�(P�!�D��+��UQ0�F~� 5���[:MM!���V�Y��	:v %)��zl!�� "hb�:E'��(��)-r�2�"O�9��O�9t��1��>u��yv"OB����Ы@�"�!ŀ�wE`�!S"OPD#��
�����`9����"O2�z��N�$:�r�(*� ��"Oܻ��=U <��W���i�"O~��i�0+�
��2l�+HP5P�"O��2���L&�A�J<9N ��"O�4{�O[`�:��P��76�>�{U"O"@�E4}^z���C�t`��6"O>�8�o\\)�5mњhQ&pz�"O��y¬�0vo���@�(�H��"O0�`��V�L`�;��=��(1�"O���"��sd0	P�V�4�؇"O\���OG�m��a�a	�i�ł�"OP���)�-f��0�ڂ
ND���"O��Ģ��lPܛD O
}�p���"O�I"v��56�x5*e:4�$ �A"O$\9%�ڊj�50F2CS���a"O �1D��=� ��s���҅"Oм��!,SvQ+`�+����5"O�Q�l3c��Iz7�X;��+�"O:<s��,��)��n׏n.�Ж"OT��1m�	p��x҇m �X�)JR"O��x���)'�,��,۴ql�A"O��2�2[��Xk�l؏&lvq�"O���v�L�GpŘ�j��]N�G"O��j�%�9.H	V�,�
�"O:Jp�̐����I�4����B"O�#a�VQ��JH�_��H�"Oj|+�"�9I���x�iֈغ��"O���S��k a� 4����"O��Y�AC�F�<�{��K�U�Z](�"O�0���֣0�]�$ψiu���"O�0�T�O<:8vp�s&V���"O��ݩ4U��Ѡ�� i�µ��"O�0�M0Vu�"Ȱ`Ǧ	k"O��i��1_�|�6��0��Y�g"O����k�	/.t"D Ǯm�.��"OԸS��ӽec,��/^)&I>ܘ"OL�� �?4͊�� ΄,I�P�A�"O����	�%t�k�G &^Ժu"O�Q�cR��Ȃv��u8��"OrTa�+����W0�x*�"O�A��&��_D~P�$�
�X�XK�"Ol��B��HK p���U����"O@�4�Dք��C� :��j�"O�]�G��t�l4���E0,-�"O!��鑴c�T+�'% ���t"Oh�:����f�h������""O���t�Q�ώp	�����Y"O��P��6��b�� V�ؕ �"O���RD#M3�l�p��
R��7"O�ɛE"D�c:Nq�"�ܶ=_<��w"O9ه�N���r
��d��H�"O��� �F.S6E�3�[�F ��"O��zF+���v)�E��LN���"O@�a�ɔ>=��h��ù0�kW"O���0od>��S�Ȋ3�v�S"Oܰ�1�)n9�RB-՛0z��30"OH��1$�����̕c�is�"O�IKf+X�M�����,L�N�l4��"O��`��Z�^������^X[�"O�@q�*�?X�]���
�n��"O� ���@N�A-�&�H-�ms"O
���`� �������&"O�j��,if�c��;��"O�Dď�8' �Qpa�`uyg"O8��� $j4Ԡ�/sެ��"Ot�!��Ko�" �,\�¶$�T"O���䍔)��t�Q�^/O���5"O��t��~��H��/�.���"O<���V�F��iW)l��"OD��q(΅v��[aH
�t��aT"O�a�5����0!���%tQjq�"O�Y۷ֱ:����'�w���7"O&ub�Q3o�`���گ=����b"O���VM����BAԓ>���A"O��������Q�"���l�v"O��D��gR����>����"O��HG�`�D��b�X8/�HeH�"O�Z���k8ԍ2࠙���e`�"O�I��mɌ���oQ%T�(�j�"O�ݱ��?t*���S�U��t#"O�Y�� �_���NF���<3%"On���T�p��� 6�H"O���/֏(.���]�1�K���x�O|9��ᔅm}�XԈN�~U�q�
�'��0d�O�C�%h�&t����'�L{0G��V�I�l"p\�ِ�'�	��M'(H��ڿR���b	�'�8)�̅.��lx��^�D˖xB�'+`�[�	٤?���]��2�*J��y��c����+��M�%c�����y��a��b�d�"�I� :��C䉄`�Ε���X�Ά��B�I�_�2'	�+i����;Y�&C�� 5��T�r͌IV���EҮ`SC�ɰ]v��5�ϋ/�Y  �'����<�J>�ϸ'P�!c�	��Oeܔ{�S,��0	�'D1󣄊h��:�nX�dd��'����C��P�-	�>	�Q�<1A@!�]�ԣ�9/ֹ�SK�<�`���g0TۧJ7+�is@�]o�<��F5_�v}�`m[4f�����_�<��O�"+U"�[��\�{n�2�J�U�'uџP�F��~���3��?*��)Fa�W�	u�Ă2�*s`�	�e�z��|�q�?D�<��IQ�4�ӖT�g�<D�XB�M�6^�����Mծr��u[�?D�4�e���?��={�AYFX��p��=D���4�N��jP�k�M0t�A�
:|Ob��y!��|3�xwDOb��s�6�	h�����:��a�gٗ� �H�+M^P8��E{J?Q�ԉ�{ô� �+���rXR��0��3�O�<��ɘ�UI��ŞS�f���"O�h��\ʮ��ժ�M�,��"O���̈I�L�$H��l���ǋ�y2�A�F>�( u((jt8�d���xRI�\��!��G��R%�7�۲s!�d۝g� �BjJ >������%�!�䁛1�Ɯ0�K	�"D�}�f�Ϟ2��OJ���D�B������y.���%�^�,A!���Nt�Z0m��$� g�ݿ�!�[x@ũ&� bV��84 @"_�!���2x��g�9J-P��(4�!��-l;D�(Ԇ
�C˘�C�ț��D$��|ڎy�
G��bG�X�n���3��S��y
� ���F�]����g�2kA�S��G{��)�~��5�"��?��=�#��3'!򤓻U��y9&���L�d���F�K !��j��R;k����F�c�!���x�T؀��
_a�#��V�!��.g����A
u4��ؤ"�4I�!�W�F%4��t*��?d�e���x�!�d.aㆉ#2'u�xJd�W�ux!�Dhf�����%��JYQ!�^MLq�1�9h�n�ʂ�Q�kG!�$�4�\�bT L�L��
`j�#%�!�D�:��a��U��+��n!��Į'�XеbŽpN�⢉ 'm!��
m��tk]
�:p)F�5�!�V3�H�Xt�18���(�2K!�>G<0��蟛n��]��f��_-!�86��S���q���a�Z�	!���7+.|�L�8���K ��[!򄌛v���xU�.vLİ���9a!�D�$T]�@Z7��B]ڔ� ٬x+!�\]�� �ݮ?�x�a��R�V!�I�C4�m!��W3�✨B�_�BvbO:�Qfo��'���ᱥ��r��T"O�1���3@	��9H�c"O��;f#ǖef���s��4�]y�"O4�@J޹��1K�̼f��|0A�'��I����pG�a�B�3TŇ�[^C�	�8 (�Q6h�'p^g�Є��� �@y�ʝ�`r�s ��:�9��<A���SRv.�DɂF�HT@Q$_3Q�B�I
;/dԋJɔ�Dt)�]�[��B�ɏ|�lxȑ@B��
�S�c�֒B�	�F�&m� ,K��i�V��(k�4B�I=���H���:`n��U<��B��	:��Ly �ؑ�:��E��4\��B�I(��HS���J��*�7�B䉑}5�Y#Dd��a��ҲKٳp�C�I�R�09�JX�'�p�ː��4J�C��rʲMK,n*")�tM�Z;�C�Is����T�G���#`��E�n�=çm+�di�IP 9M��;Ӫ�.m	�A'�4G{��TФ@�}���Ӷdy|��"@�8�ybLF1a:�Ÿ#�`���SAX�y��J+��XA6A~4s>�yr�Ԍ5�ȩaޒ0x"�U�y"��Q�B��T��p�8��_��y�(".,<�t��(aTH�x�����x���1:EK��ƨe�|D���FO!����F<2J����=��,�HK!�ޓ���×C�~0��Ū�l�!�d��a7�m�0l�Beny{0�1("!�Ĕ�~��E_�)-"MY7(O8[!�K)�r�/9����^!LJ��'��EC�di�0-8g�����X�	�'�<4B��Y�eqꬳՀG%�"���'�� �J�`	�J�)O�P��T�'K�i�)� ���+�/��e �E�A����'���A��{Xi[JuI`Q�'�.�P�e�Z��Hɦj(gϴ��'���� )A�FC�<b7���`�zm��'wґT�ڤq�"��v���@����'W���@��Z��{�hR68HD��'�5J���0�PF�� �`� �'=Ҙ���j��K��Dv�]�K>ُ��� ���M_�R����L	�3u�[�"O�@��$�6��x�+�{�V�	�"O�]	a�C3u���d��!.k�\`�"O !X��\+�59�k�WlV�0A"O�D+�O�4]�&��#ܛ_bt� A�'���!�`N5��Es��4g�83E$�O�J�>k'����l�ց�(i����+�h �
kI\AP�o� x�����p�	�q��z%��C3-&q���ȓ,%J��.}żA�To�#&���ȓ,.�y�F� 
<t�R��7 $m��t�$��D�X?a�Zy�6��Q����Is�I�
 f�@���=j�7��!�����	�<��$ЯI���I&ESch�)����}�<	�M��L�*�e�ypRt� ^�<a���X�Z�cs�ɒ/t����<����O2T�I��Yy���Tk�c�<��%�s<���`�82j*aq�*ZJ�<�d̱!�:�A"LQ28&�C��FE�'�?�J��!mt��1��-�x@Q�,"�OH�	1���G޴ �@5����B�	�D�P�1uf$?NeI�L��`�<C�	�=N���U��1�\16�EI �B�Ʌ�l�ec9_�q��X�I�|B�I�]r��	4HI�&�
/L�JVB�%{�zI����X���p�G+C�FB�	�m�|8���V	��У�-�(|d�C�	@jN�c@����T:��5IRB�$$=��(�(ĺ��U��HOB� JJ���@:�ā�s˅��C�	#;S�h��(�l�R�d�& �C�I�Uh����HѪ'�Z�Zp����C�I:�4h`�,|����'�M"�\�ȓm�``iq���;�Sj�2q��	D�'���YD�qkRB���?��p��'M��R��6�n�r�l
�:-��'�z\k��K9��X���6��ܢ�'�ͨ���j��aՋ�#(X�'&��a�7,����揫!���
�'�T�`���_�dU��k�$��	�'v8�0��Ґ.�@�S&=p[V�h�R� ��	�A\�@Ȇ��^�𰊥lK�Y�B䉫Mm� ��L44¬iS�	�_�C�#$=��
��k�l��DG�3~�C�	�`wR�X'#]F���A�F�-�~B�ɒls0ui��
�}&����|C�	�DI��%��nf8�����u�J���/�I1Sc�-	`e�L2ՇM�_x��)扪,�T%Z��@�4TBT������(��I
��XD/2k����J;E�C�I�Bx�, %0�.9��@G�8��B�IE����ҏ��6�Jd���E@��B�ɠTڸ���_/0L�&,�4�xB��;]@j�r�1��ó#U�4��+$D����ӧ7"V�§� 	w߬�8��/D�t�1"X�^����fߝ*�9��1D����	#~�`q(��X�<ud5QF�$D����AQ�8\���"�.8g\��E>D������,/[�y�W��b�(뢊/D��Z%����#t�A'��	�.D��@�@�$�u��P��%��,D�d�rDJ o+2]� ܄F��š�'-D��t(	)6L��t�� 4)���'��n���P#��:�U�Q�$
����'+D�� b�w��X b|b���4���W"Ob4h���EI����
��|��)�5S���bQ(�^+�ݻ"�D/+":C�I7
�,(�W*I�vS����Hçg�XC�� HE:"���r)��W�_�,XC�IC����'�2Mİ�]�4�C�	8+U���A�>h���G)ٰ'5hC�ɶ_o>XB�J�9<,A�D��8C$�C�	=
�x0���d�(mAI[!o���1�o2�iD�?^�z�k�6L�]�ȓ1�Q��U�8!و��@��D��i�Vɸf�1z��H􏕘8ɰ��+�:;�LO�*,��.��@�ȓW���I_�Wr|q��DW�<H�ȓ�,�QNB!$7.=����go���ȓ;n�\��a\0>�h�+���V`f�G��7J��if�ڵ�EZX��C�I�d�ԡ*��wn�A�,�0^�C�I3����1��'F��� ��W�8^�C�	�%Ϩw��.����AJx�LC䉳��9E�\k.���f;Ek�B�I�8�O�*}��,ƺj`�B�ɰr�̒�ϓ���I�D�>$߶B�ɂ&��$bg6G�" U�-����$�S�Oc���S����Q�`@�$�q��"O��1���?����@��?�쉣�"O�P�ce�/���1w��D"OnTI�fN�nB���CQ��`�%"O�Q2�ӎMp�ɒ��"l��(e"OP�s��v� \��~�D��U"O"��`'ٮ[�
5��#�N��D"O��2:M�'���Q��"O
�Rْa�z�rǍ�`�H���'�����h�"*�s��z�O���!�D���d힔ʄ�XЅ�3o�!�9,x~�9�EQ�H��L���ΦW�!���_$�u��>v1�u��p�!�$� Ul� P눗~U��@�
y!��ӆ<f� �4,�k�r�ȷ�ҥ!��(8�=�VGU-�>�pgI�ўP���([]>p�R+<o����A�
B�	{` ���:pi�2&�P�w[C�	 f��ٱ�*L%m6Q҅f��%�,B�	%,Ƽz��ߥr\�Sd⍻e�"ʓ�hOQ>��Q���Z6M��I�~��ag.ړ�0|2¡ 2�� ! 
e��Hóc�~�<�j�`�}��a�~�6H��Á�<qI��QB���!�<&�B�C�/�c���0=!H�x��)�bf�>���DD�\�<��C��:}�ɕ�F� n΁)@�[�<IB��&2���iSM�7l�� �e��G{��iӞ@��#�kV8S���s Ю=EBC�!PJ8F�v���ȆI�tC�	�k>F(�VM��� f*��Se&�=�	�'#����X�i�z\{�.}8ՇȓW�����AX�E�p�*Q+�r�B��ȓ�ּB@	��8�6(J!��7 ��O�ٗ舤4U<����N��؄�Y搲G
F�O������эWn�݅�I[~r� �5�\�c7!U�%�@]�p�Z9�y�^��>J�⊍}&�$,Z��?�'��$H�(�d�.�(�Eڋn-fi��'JZU����?Ҽ\����B~��'���)s�_�y\ ��C���Q��� 04u��=I������	\̬9�"O&<�+J.9�pC�b.xܑ!"O��˧%BaI�%���KA��
4"O�1�� X�P0�Q2P��3)��IP"O$�kS�?h��ȱM^�;(����"O�TɆ��Y�}R�	nX�8�"O,�1�Ō15�����;\D�Xu"O�u��k[� S��+A��\X|�"Oz�Y	��I��(B �K�B>���|��)�S�
WN�+𤆍i�
�ӥ�M
C�	-��X���4�w�1c �B�ɯi�
����P"|y6x�$�dM�B�I�"��頏�6Q��$H,�8N~B��3a[r0# �2;������M���C䉟��Ӵ�� ^T�� E�C�Ɏ;||�"B;7�H͒�c����O��$I�#��Db��OWr��S'k��.�!��ȗ.	��%'c4D��,VV�y"�I�6�^�J!4<�J��ƥ%B�2 y��������a-S�2oB�I�=��҆���xJ�h��H{�B�c���8t�,6�$�bV+qL�B��+X��T��#�Ȅ2���5T�fB�'[�D�#�A��|Q��5�DB䉢�|���!�z��i�7w�B�ɡ�n�Ӵ�@�BJX��� �.C�	�1Y��#��u�N�k҇V%%<�B�	6-�l:�f[*3�>�h���=g�C�I,���d���d�2S�L�)�0C�	�mE������".�D�4��?D� C�I7axe;�
\�0�E�$!�6c>C䉓|	�Y�>)�t� �*C�	�%�R�����6~C�@�%�J_��C�I
Pe�����6#��9a�7��C��#u����
V�zZJ��Di�x�xC�ɆL5�S��5:4p,ʲĆ.1lC�%jb4�
���������;^�B�	���Jߠ5`�Ń7-E�x�B�I�1�����엑ڮ�(r(ִw�C��3|��9�-V�*���ֆ��FC䉪D��p7�U�v�9��O.M�B��8�@
d#�-:fqjq�M�x�C�	�;U��jQ��55���c̣/���D{J?5��m��0�fep7nY�E���<D����aȸSYt}�B]o.�l�  D�l��G�e��9��h�O^BM��+)D���G�.x����>�4)�G
�O^C�Iu���8c���Z���c��� B䉼��<{�a�$ ܐ�G �f�C�ɀ����"��[Mh<Y���C�	i��#*	$�D(���mIC� �A�K�phδ5��1OBC�	6"ޢ��CT�r�:�I&i��B�	�7�:��W�[�n��p��y�B�Ƀ+��)��%ҙ )�X3r�O�,̪B��;"��hk�+��E�͊1I�B�B�T��2��:��5� �˘-ŸC��&3���F*_p��aqV�:~����5x��4��B48�h�S�`�3����ȓ�TÖ�� 
N�CE�R
6c��G{b�O�Xࣗ	��8��FMχ"\ �'yđ$�I�yZ��X�ʙ,F�N;�'����O�`b�8�h�hxx���'�4�R�c�5�<��e�M[v�E#���)�� �Y��N�r�t4��$ɜj�z�*O� #d�x'��"��B�_:����'�vp�F�?L���ǦPH ��OT�2��)QT�:�#t��ss"O.=��K0�����Β��-��"O�u���P�J��Б�0Ԋ�"O<ݰS"ȏm���C�sN(��"O��a�B�ܴCE`�kCf���y��U'y�᫶��$& :\�oX�yR�� ����5*L=�H=�+Q��yˑ	� �ůJ<jv�ۣ+���y�h۾,��Z�S��t����.�B�I�R�V@{sKU�=B�@DN8�JC�ɞb{�Q�I���QI�� �bC�ɖIkf]�a[�@3�E��Ě���C��O��q�"W��*��rTVC�I�7��h�GP,6�։	�h�+�fC�	;b��$�gN޿
��p��XC�I�D̕1f�[�]�y�r�YH�B��=6��U�&L��t����˥CC�ɿ^�.1H����ѵL6_��B��-S"<�iKn�ƕ� ���B�	:s�v����O�r �(� �LB�	���%2�(T����%B�I5n��-Ha_#����6&TJB�Ɏ�z�jb���k����:�(B�	�$(k�!Σt���#7̏&�B�I��
�����7W]� ���	��C�*����D;yz��H� �B�	6a�4�h!˼),L�����C��~�"�Q��4t=���d(V 4O���$8?�U�6-��!8�GQ:,)�X:a�t�<ib�ü���X�X���(��[[�<��ì� �)ŧ�
)|1�Y�<17I�2ҡ��.�(��`EY�<1�'@�[
x��D�0B�2� mL�<�1�>y��hr)�,(U𸓷oKK�<a����(���Y�]D�%�f�J�'[a�B'/��Sa� �J|�w�Z�y��S�p sՆF?�F�QF���yr(�,���o+0���h�	���yb`ӀDG�R�3y^�hr)��yrK\?䬥�ׅխ~d>��i��y�G��P�a���\5�( p�g���y��L�"`�M[d��q�����y�Ǔ�l�X0��a��ڜ�y���KH(\��I
)�yQ�̭�y�"��*�b��G~e#r�_��y��G(g�:���N��I�����V��yr�A: ���6:lz9 ����yҎ!Qȹ2.3L�9u��yҀR4�tx{a���Nj���i��yҍW*	$T���$&B`D�1�݋�y�#V����Y��N�SY|9�g��:�yB흯`���[צMM�=�F"�y2J֏#�¡�4��A�%�dH�#�y�"ߧ*��q�gǍ�3�V�S4&�/�ylB�U4iذ���V�FPj3DǄ�y�.��f�:T�B��U���Hd�5�yb�B�b� "�%�-7�A�	�'�^(ɥ ��r��-�-�����'�黧j��m�5+Ĕ^�a��'ټ���S��0���Bd��'�.��&�=61@�0;c�x���x
� T��b#�X�&�;R\:�k�"Ol4cr��	ru��3@���\W�e��"O
 څ�K4��m@�@:&`""O�4i� 	�Q6�Ko
-�*�zp"O���'i���2��C�Sn��S"O,rSX�Vr�*ݝUl���W��E{��)I$��c6Ȓ����Sʐ5�!��s�JP�#>F�tG*Q�ad!�d��F�����Ǔ�0�(�(�ɕ"�!� &Y��xt��3�2�:�ԙ�!�DC~���CGBњ	����ֲ&!�D��Tz�٪+��Dk7'@�g�!�E�bw���$I�,hŠh���0{�!򤆁�^��jƽ4��lC�@�;0}!�dɞ3l*��uB�;�t��t�B,!!���6:�N��@g['{��<�� ϸB�!��ۃ��A6�Q%�}X�  m�!�d�w�U�eێO�� �����!��W�x�`�5�Z7(���ct�P�!��ѮoC>��E9r���h2��t!�DIV��5��aĶ<���+־�!�D�����0��n�LJ��M��!�Lv��RĀ3oȺ�$�(�!��+wm�ԃu���
@ �,W�!򄐯}�N)�"�ּ�<�`&	�}!�d��laL��Ј
A�:� �%	�_u!��{%��q��+a�{���8jc!��w��c�ˏ�`S"�h�hۈ��OV���NXŖ �".�+,#�D�[�P��'�Fy0��_tDD
TEl�%8�'�n����\�@|�g�;��	�'9B)	2c�o���&e\?n!�e��'H��9%��?<����a�bL �'�L��K��{���r0aI�ke�`��'�
�Bp	��&�Z��Z1���kO>�)OR��	H<�eB �0hL��Gǀ���IM�����P�&t�� ��-c�����<D�����Ɓ7�0�X5�T_���x$:D�\�0.H+T��̪�H�)��`+9D�X	���-=^��Fk�&u��2��5D��W��6�Iq�J�X�����-��<!�' ���a��9}B@9�懞�Z���$� ��	60�H���@8#�x�s��'�T��0?��#��$���d7�l���A_�'?axR+ۖ ���1��z�޼���2�yr�p�4����t �c+�y��f�~M�@��f��	����yh4a�v�#��
��Dh��yr,	}���
�I�Y���8�䓏0>��b�o��-H��`�3F*���"O�<�5�ơ��:���}���"O`�e�@#)���+��B��kF"ON@K!C��.<���E�kJ�"�"O�"D��,
��#�H�]E���"Olx��ήv?�1���+W:�H�"O���D�vaS`�0[�jxq�Y "�!��Y$]^��Rh��$)�!���,�!��$V��(x��\�#�����de!���p>��⋌�'� ���,�@M!�D�s}614��=U�HU�֊��I(!��շ*G0H	RÁ:]k<	ʴk�2+�!�d9`�z��c�BhB�,̨_�!��Q")/.գ�R��`�v�M��!�d�?��,��1}��y�F��'0a|
� a҉�0
܌���ó���2��'�ў"~���V1sX�4*�銎c�ހ"�+!�y-x��x5͕4Tm�șR�
��y�d�Y��:�lC&A[��E��y��.�d]��!ݪ$��Hk���y�eW)�L�Cg��Tr< f/�&�yrT�$F��:B1�1�%����?I�b�S�5�FI��T͒�	�cۦ���	A�'9�1� �ݔ⒮X�@.np��'�(`B''�#H"����́;�T���'����&g�(�.�2"��5`�'��I
��A`Z�!�f����TJ-O��=E�t&ҭO�H�t��y(�:6�Ǿ��'�az"'��`zD)��of`��ZH$@�'zYHe�B#�bl 6�[(%d�4 	�'k"�p  �4��d{��Ў�����'�	�A�T� 銄(ډ^T��C	�'�pS(�:��R���R"(@	�'Qd|AC�ƱB�l�C$��+DS ���'�����C�Ol����C_��1�'P����2n��iǐ6���
���y∅�H�*���
"M��e�W�ٻ�y�� ?`|l�b���f�Y�W��ybI�q[��Z�^��ar@���yҠ��n�Ȍx��Y�$� 4��A,�y�@�v9<�F��&�z�M�*�yNV'w�1�Ff����E�P [��yB�H<�Rlb�Z<p��X &�&�y2�%t���߼7�`Y�,�y��V2^�,��e�ѷ3+�
&���y��r^-EL�b�H���D9�yR�<	2$� ��R9�XH⯔��yB肦1�H{@��CI���	�/�yҤ�,w�Du�gcJ$A��!����!�yR���<M�'�D7B}�����y"�W�?~�Rw�ٔKQfɱ�-�'����'�>	�)a)t峲��y�@M��h�O�C��C �;�<1l�\�!.Q�>|C�	�-�)C�*�X��!!Q�r@.C�I�W�ً�瞞Ӫ������C��3~>���	��K|б�&N@�B䉲i�VS��ӝJ�n�ڂ�V�O����0?�,x-����Q�!*p���DNx���'/�pǁ����P��L� UP
�'�hU���(D�|��e�J\x��	�'j���@�&�ɥ�W���+	�'��p�Ĥ�0��3��
 u;�lP�'��$0"��4�� y@Ѣe3Xh��'��q��oU$u�VY�ᅎ5:�
ϓ�Ol���]�J��M���G�a���)@"O8��O^ul,hI�R!�ީ��"Oڹ����"C �J�-E����v"O�ҧ�S ��y�F�]�(�Դp`"O�$J昡U_�i@���cq"O�TH�Ղ�`���-OpH���"O�j7,�	 ,�M��B�&v�IZ�"O.���+�mC�d;C�RUX:�jF"O6�2 H��u�D����ON���"ORm;�h~������L=D�����D�,�^�Kd�C�6�z"�8D�|0&�@�U��h! ��^�.Hxe�6D���@�F�
�Hc����P4�bb5D���������D0sj�$W�w��{Ҕ|ª́kU\�9�BȾ[T�䘡��Z�ў���3� ����˙l�����֏-4B@��"O��Q�%0p���D� �8@Z�"O����$T1�
��P9=~�[�"O����Z;M=�!�/Y�@�\�P�"O��A�#00���Bo�c�@i
�"O�]�R�Z����O� G�83��'ў"~B���6BLDS�$2Pࠋ�P��yb�гQ�l����62�>I!�N�y�ɔ�%���Fo�.�f�P�W��y2	�T�p�:�޽��M��y�H�13�nQ��ŒM��9��'���yBd��$����(�+>�� #"ƈ���=A�y�틳9x�б�J�L֍����yRŒ p�� �I�[��wIA�2�O��~�p�i\�#�v�!'
'[>��ȓo�:�XP�Էd���Ҩ���ȓ>�بq�R��*��N�o�v�ȓI���`���xl��A/I�d�Ć�J(d[h˦�F��Ă��_�YF{2�O#����1Y��`;����':Q��"�X3@���ϖ.���Y�'� ����<c���[�!43���R�'q��
�G� ��-���T?E�%[�'@�)�Lso~��C��Xt}[�'��Eψ5��D`�Y?2���'������Z1�!P��.��њM>������*��, ���k�$m��ˬ��IS��Xk7��3]�P���ݧ+�n4�=D�,#k���lQ�
�*6��T�>D�`sE=4����C�<�(�D"D����)�C��qD �3�e�t*:D�xZ��Nb���K_p�l	5D�,��]
��ly���6 v�˃�3D�� ����_jm���D�_G:���i1��#�O4\k�15��81p�ɂ�=C�"O<���u��@Wk8��R"Oȼ	ǃW�XMpI2�U�\j�[ "O��0�H=7��Q�
�p"O�����j����ԍ
 DYH5"O@�oR�<�(д*�l�FiA�S���	��H�?�}��N�a��0SCqNl����f�Q����yR��0��2t��1���f&ɇ�yR�]=~h�E
vmJAlԋ����y�"�{�e�aӢj��Yڵ �*�y�`P8%jR�f�Å]�ny�E��y�!=vD�t��J^�l�ldb�
�t�<QT�O�-��X�������o�N�<��g�:���U&� &bP�C�Us�<��%[���l��E����ЧFm�<Q�._�p��IwG�{I�X�U�DT�<�RݡD���C�C��I,�X!�J�U�<х�I�f}c� z��=)&��T�<���@���L�l@��CJ�u;!�D� ���7�̌��U;&��1!!򄏴e��m!�U�v��,��O���!���e P�c��6c�ᱶ�;�!�]� �x��G$�1���xY�gx!�ۀ@sR墐�_o�>XӠ�N%k!� �������"Vc8$�C+�Z]!��Q�(�	*R�Q�!4� cu�ӞY;!�D֗.��\�͙�@]��Ɣ)!�$\�P�����kY�_����0ƌ>p�!�d3".HJR7_��t�sk��,�!�-K�ZT�5+_�8	Z�$_!�� ܉ZC��*���	��P�ļ�4"OFM�&���"9{r�̄,��]��"OX��f)�oK~� �E�P��u"O���4hщ �
��S�N�F�^ȲW"OVY�T�]%�pTZb��3Z���"O������#���&)�D!*-�"O��c�.�7��p�2��P��@"O�=K򋃪fp��QƦمW-�h�"Ol�0(���ً�E7E�.!�%"O��cPL�{��"d��D�����"O��dOA"/���p���\~Ɛڰ"OL0��#�~��s��gs֥	�"O��Do5$ni�X�>ț"O ij���s�1�4�_�c��q"O�R��]�{�u!� ��T����G"Oh����ܢl���#0��?<����2"O�$���x]��y�f����ȗ"O&��w�Þ(���Z�$׎K�"X�"O����Ah��B�Rm㚴# "ON�҄�b���G�ZE�"�:p"O��а˴GL�Qs���6;r��3"O*A�f���j���G�H�t�"O6�R[	ߤH���>b(�K��M�<����hT����"���%f]u�<I"�"yE2q+d�	�j�����Jq�<���<H��T��EC�<떥�j�<��.�):�	j�$�2J����{�<�a
G�e���)#F�.&r�UKAĞx�<��oبh�$QD��U�h��6�[�<ɶO:' ̃'d	��ڽb  �`�<Y��ز!)(lk�]F6�qu�H[�<!�!T*J�T� cH�2nf�)�TY�<�wf�"W~�}sp�*�J<��i�X�<�T��k���I5DT36��P@�R�<�P� m�ш��O�8]�v��i�<q��K):7�B��-X�p|��Gz�<�6�=	2�� ���J�K���t�<qЎU����V�Tf��7� I�<)g�4@��B�u�vDC���G�<)G"�bͬ�FϬPb�*P�C�<i�$ݔe�B�8���BC䫑C�<��Ψ=���gl�1?�XT
0�H�<9G�q]0�A��)R&T����F�<	Q��!9nܨPe^w����� Rl�<isY?gO2�j��	����`G�r�<�⁁�=@��)�-w=J�%`�v�<! G�.Ⱦ�Pp��&m� ̹��n�<Y�H�6��P�_�<]����f�<qA�B��eYԮ�&�\����\�<����550���g6�p��]�<� ��?�$�p�<z��EY�<�2���F��Y��m9/f�˕eU�<�j�At�E���݋^�e3fkQ�<9���[i����� 4�� �ČSL�<�1�ʚo�2|�@��$}Ot��$��s�<��O�p�쌳c,�!6�R�2��Ir�<A�jأx���M �l�so�o�<����{��1rRLў}�Ľ(��G�<�A(i�N-
��nM¹��C@�<鲁U �օBD�N��X�Q��1D�xrUď�r&*
�K�e:�
�//D���e� ���m��ɵ}��JV�1D�8QFF�j����$i��r�3D�H��CG�Tb���C��H��а�6D�� ���@9E�h�B����ss"O� �KΙP�9��Ƃ]��`Y�"O�}r�	�[<)�@�FX��!:�"O
i��k��IPU���
�h�"O�<z�h�x�z���b�LY�#"O^,���8���EDT�&@�#�"Ot�f� p~�$�KK���D"Ol�*T��/���"ӈP�6DͰ�"O���7ʺ'(����f@t*"O�!����>-��F��Dy"O�=fJ7lR��FET�Lat��d"O����yq��Z"�Q�]��R�"OЬ�v�#��R�BŵdV2�R�"OF�'჆Q�l1sĂ�xL� ��"O<ّ�[:W�>��@��bD� 7"O�LR(�m���i`L7:9d� 6"O��2!�9ܸ���ˋ�8	h|z�"O8�٦jP�A���kE�F5(�H!�"O:�F�<9�� �1I��(��B�"O�P�@L ˖�"��>!����"O*�@�_#f*��ݷ�̫�"O���㓳pj\�����6@LL�#G"O�u#s�١v�4B�^�C�F�xT"O���w�V�$%�eW��4q��"OԱ�吢z���CD�pf5��"O4����n�j�y�Q�G$�5�@"O����,�9rD�V ]����F��n�<����>2n�i����V�Y�E�c�<�`�L\Cb-��/M�n�7i�]�<��M�,!b� ����97H�V�<!���%�\I$o�3E�R�+T T�<����~-z1x��*3-��!�EHu�<ђ� ��ݢP�	(Kst��!I�<)D#�"%W��qHڞ|��D�E�<��MG�u�pE���!f��D�^j�<�"��F����F��9J"%��ƍO�<	�Ӎ6Nl�(�o"Ep"��H�<) �ʭef΍��O�N6lV�n�<!��70p�jH�%��|s5d�j�<�l�I�x�i��?nT�u�qύd�<���Û*k���bƘ*��ч.�F�<Iƛ.otv\p���s6�e�te�<	��{=��!���
������P�<����@��XB4��!$Ɇ� ��t�<i�˒;\�8�Q��6�H�ԨTl�<��
D���Sn�!O��a��k�<��w���y��\�,ze2�A]d�<	7&�T:���^+\�Z�-Pb�<�e'�,}�ԁ�
�)x��ih�^�<�Q�?�}qѥR ,�}�`�PV�<�&�H�i�	rON;Ur�(���Vx�<9!�ť9T�)�3��M�ŏ�i�<����dV'��dcȡ"t��y�<q@�C�D�d'�v��Q�@Ox�<�� �.>�6�8�!�q�D���)2�$�W�V=F������b�&q��ne�}S���$
�F�`Y�ȓa��k$ޙ\�Z ����6v9�Q�ȓU���c�/�M�|�,S2^�Fن�/�pM3UO��	�y�С]0B!@�ȓa� ,+�تl1�-!A%԰B��!��^Ax;w��Q��A��%��N�6X�ȓ p0xC�Y.1���QMׇY���ȓKkt\zT�U=g�Ns0��^����S�? ����nCԆ��$%E��0DS"O�����*x`Q�U"[\b��@U"O,��Ԅ
�R����L?;E(s"ONA�ej�� �I��O�=8LJ�"O���⨌�,Dx�s�M�!$�%�"O=�0�\�Fy�Hr0G���T�R�"O�DUAZ�`�x)���ƹ.ɎPX"Op2�I?S0�:c�k��:�"OfIk��L�ƌ�*Z�T#��P�"O�M2��J%Ľ�ų=(�bs"O��c�U�� ��Cf�hhԍ!X��G{��)�-z��J孁�1���1�r!�$��^���V�vͬ��V��7e!򤞹J0n���O��)���͝/gT!�$2v����CK���@&����v�2}J|�'���"A<����c�Va1�ѻ�'Kҽ����n69ʡh�%L	�ٴ���}����P��K]�2��
U�q!5�>D���F��5(������'��@�.D�p�@6�}�F����G.'D��S�U��.�q��R����e*D�H�P�V��J�mM�'�f����<�	��`5t��8�~1!�˝�f���D��(�X��(�7L��X`� Sk�(B��0>��2����\����1hD������ӧ.W��{�M��l8��t&\+IO�C�	�8m X��Ş�}]�!�&ك�C� 
O:ћ��]�=[�����l��C�c�D	�!K�}h�|�wj�M,x���dq���>%?y��dP*��L�'�-n�:�O��'BZ����@��Jd�E�e��K�'������)7�@�F�IKv�8��$8�2�v\�s.2M����"̈́]zr��ȓS��加i�><�Ycq+رn�� ��=a��I��1U��L�pC����ȓ��aC�mN�%����-�,w������A���@�J��q�ƅ:����U��B�/ґ��%[�+C0ʎ�� ,O�QA�oҘU�*�k��wg����"O,�J�)�3&zh��+��VX4@��"O`����<	�b�B/I0i�W�K>%�$�G�G�x03oP�l�0c7D��07)@x�����Z�UubT9梟��Ӹ'�L�"h�b}d�9�Ν�X�ݘ2*O ���Ʉ3�<m��@^�Z�
�c���
�J4� P�[�
�hS��B+�����g�d�<���̧1:&H������1����<a��*mܬ1��)N�Z`���w�'��?���i��V-�q��"U�0��đ�&4D���VH�<]~��D�����У0D�@���.?[L��)Q%z���A#D���qέ4eZ� ���$K�*�&D��q�NN.[M����сB6ECf&D����۽"դy!�ї
�l X�/D���7��#�Da�	N4e�dZG�-D���I�4H���.�?0�+�A0D�,cs!���:����ib�R#��>э���4���#QFv�����^�C�ɕ@�P��(	�F�	�!�O�㞘�� V�Rz��I�I����[>4_�C�I��MQh˭|4����7^dL��f�$D�<��8yq$3p�(��SB%8D��0�`]:����BŘp��@A�5,Ov�<A�D�(��t@``��R`R|Y0��i}b�'l�|
� @Y�v� (������lG�(X�?OD�Ic�S�O�$I �˚�1�.��2�Ǽ2\\2
�'0���oP��`B��%�,)Of�5�Q�b>��vD�3|_F��$ �;t4���?�O�p �'�&����0@�����9)4���g|yr�'*���$+Q���=�^Q%C���'���&6?����Ξ6�H��A��]�āZD/���y2�|��d���VdPlRA/;�������OD����	.�,��a�H9D��0"OjQ`��|i�0cE�
6ec"�'U�$�.}mL�6�[5�d��b]�!\!�D\�U_�d�)C�t��AI	XO�O������~��/>
�w�W�O<���'�H)l���{
�'7�b�E1$G0qqD�Z>��s/O�ʓ��S�L��IA�:}xL�ؐI�7^[Tl��/��"�a0l�4̱�^k��C6�çF	�'��|�$כ?D� �Y��@H�X��p<�N>a�O�p �>hw�*rΛY=��P"O"���Ǥ�F�9J����I�W#�?�z�)��5 h��UD-N��3D��I4�S4����T�1���6D��m�ȹ��`���b4D�\�� �=R$%��<Kb-�A�>!	�Ic�X�T,nq~(��)\��Q��	ty"��Sa�a4��D���e O�y�ȩ4ȸ�h��W�=�8 {d����HOD�=�O�|sSc�Z �lC0Ì�Bϖ��}��)��$x&��sI	8	h=ʕ��2��d�[�'dўh���T�N
����Ѧ�5��	��HO����0>U8��6��| ���ٟD�!��ܭe��ѩB��e�(l2��Y����F���e����G�>b�t�p㞮�y��4�&	1���3����1�F��yb��;Pu�5`Ӽ3���;q燦�y�fP2BԀ�!/?f�r���&���8�O�`@�����u$ˬ��cp"O����͢.�X\����+��t��"O��	uK���ݢ�kO7*��I��"O���D�!XXiH�� ?L�-���'��O��Q$K��S��|J"��{���h�"O�����\�|%bQ�f�
��0��6"O���b���.u
s�ZJv���2"O�i�P�]�>��LJ��ڧ}�̉!"O6X�Њɋ5�f��5����ܚ�"O�(�%�I>$�r�{֮G�r�f�q�	^���i96�"ɛ�A��^�R�����!�d܊�Zq�e�׭��� �
/b�!�ڼW��7K��a�<1�D��9kca}R�>)5��2<R�
�鞖�����\��?�(O����TMIx��ݮ�̬"ע	L!�d� -b�ٕB�����Ƚ~?!�DY��)q��D�~�����`D'Q�H���'ux�S@Z�%�,��c��'gxB�d6�c�[${�&���D7��C䉧wa�+P�
��-�1DZ�HpB㉢%1zı%�U� [d�se�T*c���ȓ$�ze9�@�%2����`�"I���[�'h����X�	�A��ܱA�ux�'6�`�ú$Ǯ)@�/\':۪0�
�'=@e���iO �RWgց&���:�'m��O��<�8pi�m�=���(�i\�	��?��}�e=�S�8 $"R��4*@�q`$�S�HzL���1��-7��AK��Y3A��m��OY�
���]��朢 '��A�GN�(5��=����� >Lې���l\��&ɼE��mkR"O>���و6�4I��l@���h�'���9H��{�a]�(-�T01O�74[2B�?T�6-ۇ�����@V#
7&�B�	'8m6:탪1�x��-&�C�'t�p�s��R@/(4��	מC�	KFe���eF@��۷�d#<��A9�S��<.x�Ĉ���8&��3�y� �W^�	�`B�tw����Dܩ�yR�)�'h�L��g�=>��Ɗ�b ��G��TID�ՑF� %�D��{��͓Q�
��䇫C��p�"�.!gJ�ZE"��Ha~�X����Ȅ�21��
 ��\)�K(D�|ʑ'��vi8��G"�P�`'��b���'*fbu��@S�z��$HZh�݄ȓ;�J�sD
*OSH\����	�j���`8�8$�5y�0ܐ!kK%=V\���H�P�RHldp�h����R�ȓ(��:b�GR'��8�ʎH�͇�>;���P�(0�(�S�R<|��ȓ,����+ԁ��z�
7���ȓ.��xR4��4�U���j�>m�ȓ�I'�ߙB!j�y�o]�V�F��ȓZ�(���J8�D��.h��+�"O&(�ckӨc0����fA%2�L4J%"OjeZk�-c޴�R���"O�	#3�'�r�0� Jv�)%"O��1"�H?sF`;f ��L����"O��١�՛Y�HQ`C?p��"O����ڨ3�
�:R�E�&��"O�L⁧W�6���0���R�"O�djqI�]
ai ��&RPЍ� "OB�81i�g1jI!�c�97?b�Y�"O�x��&�%;��w�@
?ʔP "O�Fhȱgf��S�n.Z���"OH�)B$���Qd��H�: D"O�q)��++�����	&h̥A�"O`��HG&bk��W�(�0c"O��ڠɛ�Xz8Ԙg��J��	"OJa�ƾ<2���p�K�#+���"O�0b��wC�tYc�S1�Pb�"O�j!l�+=�pɳ`�q�j("O	��@b� ����D "����"O`���ǖh�N��EƐ!�r��"Op�B�\�p���D�>+�,Z�"O�c5u�z9رcT�|�䍳�"O #gD�0y7�yZ�Aη9�̄	4��uI
4뇣Z$b�@�S�'���5��/=����0�ߙIi2��
�'�x��e��2�6I:��R�@�Uz
�'���)s��D��YǪ�A���'$H����q�Щ�v[�>+��!�'7z���Ȓ�1��x���-E���
�'d�M�W�۠}��mc�_��|5i�'�2`w-��k�ƈi7$�9��Y�'3v��2 �������Ԯ���'p����`��d}n�X�d�21$����'�����_�i��fnګZϚ!Q�'�xl�v���,كe�@�J��C�'�rՉE/§|{l$�B%U-G)D��'X�"���"�T�{r�aU����'FTX[���+�֤!!k�v�
I��'������7]��:�g�m���'�.]BBg�/���bgUm���2�'�N��W�_�P[j�����MÀ-�
��� ��+���8�0��	�!!p���R"O��z&i˞{�K��Cb�I�"OP�(��]7S�1#��xdv ˱"O �jV
_�3J�H�!D
�1vޤ�f"OZ�Z�� �\��uc��xh����"O:��5G��,i�ĸ�ca��NӐ�yRmB�ז�X%�ى�>�����1�y�l�w��$�GޢP��I�y2���e�x�A�O+�-E���y§�+��U��/*�\	�i���yr�Q�E����hF�p�`͙�A��yb��E0K�	�M���ڴ!Mu�ȓ*'|Q��A >�t�Q#�_6Q����ȓ?�����	N��I����1�@�ȓS���+��T]uty1F%:`�m��f�{���)`]�Y���. A�$�ȓrߨ����,����%\���������c��	4`,k�/ۈoW�T�ȓ~v`I"7��9:zvb�M\����B�b�a��>�������!�ȓi��1�!~��J���*�^9��-�f���޵Ik��Y�|�*�ȓ~Zh<�C�;����B��:J�ȓb�JA��G4T;pF�53���V�������|��R��5�ĉ��N�&���Λ|���#�+�0|lF���Oa�Ċ��ڦS|�I��	�zt��R���%��1'�\i�Z8!8�x�ȓR8��XvoGCurI�F��A�\�ȓ��)��[������Ɖ�zЇ�&�mY��S8qhKBށr�����)�T
�O�=$��`�&��ȓ"k�� 2��=rz<�% �H�ц�Gm��2u���K4�*R ̥8���F�����<d`\�pD�Q�	����uO�ف���9\JN��7�ڋ$~݄ȓh��lңKB�[oQ��CZCq�<�ȓw�.e��&��o�.�ң�;^=�ȓTŒ�2(��,^B��s�Ը�����Q�HQ#��+C��P�ď��P3v���O�.��ѷ'$�Z@��aklȄȓB�.A�3��8i~
� u�@%Q�E�ȓ_Ӝ(
��V֐PHE��:%�&݆ȓp/>Sl��!�z�)D��7�h��9z� ����#�n�����J�̘�ȓ��ѹ�(W7/��ٲ���]V����6h�`f�`U
p�eQ�xU�ȓT�L�H$��lP�UY�!V ���2�7HR�T)�kyE�J"Onm ���~�ܭR�咋.L�
�"O�s3�Ҵ.Y��#ɋkl�jq"O8��H�����(5�	�4��p��	:�:³�S�_k0�၊�.,J
eJQ���C�	�8ð��*\1.��أ�5s�H7M�6r]J��?��s�����d�H(NI�PG��X���"OH���ڮ (�1ç�`Ƞ�OtigM�=ʀ��=T�C��ɂZ[�#�
�1]Z����+�dA�D��"! ��K���}���Єj�4`��"Ol�*� �S�jd������[�����i+��Vy��U3^�RX�Mn��S�T���PяB��F)Z�lTP�<	`Dx�	y�m��](d������ D���7�ڒp݆���b�>1���wڎ��fl&�>w�򜻣�/�F0j#
�
����"� �2�HM�GQ&p`�o�+<3@����	;��z��G��Ys�'�2T��m� 8m��09�<:U�K�OT����GÆN(�"��̫�#�	�xR��C��x�'��;�� ،�$�V< n<�c�DHN����3"O8h���-&P�|���(4��$�$�҂ ����e�O�ޝr���K`4P�H�,'Q��O�P*�w
���HCr����+m��J��E-�s)��'b���kAv���K��/���R���
� �ܿ��D4��u@&�0*�u��FҚsS������~�?�FOg�e
-1.r<��l�=`H�[U��/s��qxЭ��<���(O�={���O[�zBh��4�!ި4��0F%�-b�1u�(���ٔ|��M`�p�OU��
�!�/Hh�9k��ބ�ڙ���pDXj�"O�88��D1,:�z��K�N0(��a�M`�@(�bS�v��X��#� lZ�g\p����dFȼ;D������M�m�y3bI�R��$$癎4HF�����J�����ǘ�t	<#$�� &�Uڴ)ڈ;�˓U�����)Ҥk'�O�soY#V,x����4]�� 4���d�T��U��>�(|)��PG��nC�df|�#c��@�B��V.�I�<��`"�A� ��y�GǞT�-����dbȊ���DY�Q���p��AU`��K|B����$����V|��#��!)̠(	L)AmĺBO>�h�� ��	 �/4�sE�W����	��~!�"��O0�5�\����� 푚wf`Mo�*r��RhӲ���	��{sʉ�U��fl6m���זQ���xD�=��em�&Mۮբ�J�y�G��/��t�m�.,��<qq�F:n����
\1(8#�[s�'/�� ���7��qa��Fe�Dx�'���4N�6����m�.Z��
�M� 	83h��_�(���@Z�P#d T�U���\�h�0�CH�!���T����HBY��']��吲.X7sK(���V*�����وJ�hy;U�z��I�Ɠ~AY1�l�X��
K�}����� ^q��$?��� �'�0yM E*Q՗�yR*�v�9�;e�=񔍓�t�$��P��`�:���I2a�0�F`dBL�5���#�����^�<(��4*�,|�4��$ކ&�д�rKCbB�	��y��9qx(=s��:�\�S"J˒�hO���2�O�� 0R����i>)#�ž)e`#�-\`8ٚ&��0�T̻1Q0X����'��M�C�(sB�
���8�:I��a:,��g��f���c���A�O v;' ^q�06-�E��*M�~�J�-���"F9D�ؒs�:5u\a1M�]��4���W/<޸sc�vޔ���M�m�|��ӱih��'�� �FOv�)�Ɔ"H�� ��ƌ�;���:�3�O���O��5ez@J �&�P��K-8vx��%.MA���4�|�'kj�HяHT8�>�qL�[&���͞�v����¯�Q�'G~� VM�2M뇃�(t3��;s4��}�V�pF�#� {@��T�'�d�)p���9'���,�;G/G	_�T,�&�K�D��I0r�x��umD�oX�$�'���-�'e׬h!����:7$ϦlmZ$���R�j"<T �e�R�<ٳ�B�v]���ư8��P��$>� �r�ܹY:j�3��q��dʓ��|�O���;}��I�� ��db��-����,��ɢ8���BF		'��@�*7�:���G�
��H��L%\����I2�hL��G'��(���b�6�>)��$�t��![�P�H#���0yT�H�4��!���V�JS"O��Ԥ]�y��1j���F���]���V;%
e��h��?��,W$Zuzm����1b�F�H�/D�|�G/
T�D��Lߐs�(X���Q�~����a��+��	)��B�ic>c�<+��B�0j�!���`�*9� �8;�*�yF �����L��}��f�|�'��OD\M��&#e~��	�p�z&��8^Z��DNr=̣?ɱK��vPe�;��w"ƿx1ըFF�:Y�i��M��	k�7$��:׌��X.�$�ǁ��__�$����<a��W�j]�3,�-��s�d�	$M�c?U�����Qʉp��S�+���rgJ)D�|�`��D/
-� i�ZƴåL�
,.,sT"�1�y���M8Z����m�M<ye	E�_��$ 	�
E �� ��T��@QID6bAC�d
�Vu��)�CT��8�c�sF��A%gKE1��h�'���p���n��h�r�ΐ�4ݰ����up�!�M�"<IxH��C�)h*T��)�-	��c�
8Ug2вGE��x��f�Z��ب�z���˄+��$�a�6��V-���$���o� 8���܏m��$��q	x���c�"�y��2Gi�t�E�[D��K��1k9"8[�f�Z3�m�AO?)��N~�a$/񤇾y��:�[D���7@� (�!���{����!!Y�Hq��;V��)`��ၨ�I;ҤCE�)<OL�DEP �.!#��T��$��',����R�z$p��8*U�0�Y��t�[���9�m���q�<1G��
Y��yc��wŌ�iqo�r�<	r �1bKH�	Ү��
�����l�<� B�����/fp\y�$=r2��X%"O��*�)k]*����C:���c�'�<� �)��I0E�Cn���*���.�~%�B�əV�u`�ǃ~	@=!G�+=��c�81V�֪?�ҍy��S�6
փY�rP@8��K,1C��$(��I�+C
�!ö��6�P�(�`�Ѐ��L�T�&!�&��FМ$��MUh<ٵ�0[��1w
�(�l�Q�	�/��P�vo��
�N�<yq5���e��e���[LG����	g��U�g!ZI@���:S�e��αy~�hY�A��>V�%�ȓJs>��`� �elʄ��+CK`~�&����kB�Ll`��DG{�O����L�/�`uu#ý O��J�'5H0�1(Y.��(hՍϯ.�>��0��Q�*O����#.�3}�.�"�2��Hɕ|*�t�Q�Ў��xbDρ+zX 3t,��!F��S$f?��Ǆ2F͒;B�'wR��3�F�{�����LV��څ��{��������Ѝ��'�b��4	 �i�| �F${�F9��'�Z*q�X,C�Lx��
L�Y9�y�O�N�M���a�O��p��&U!�q�!I�R���'�H�ԢYI�;`P�A������K/��O���Y�L���ܼ=�2ҵ-]�X����L=D��ᑥ��^UDIˑ
M�YޕpPg<D�;�$�m|]��MPs�m���;D����,!e�X�u.U2gDf��d�7D�``� X�����D�o�T���J!D��K�΂�p/�a��́[�� ?D��[5�_�|Q��ٖ�\�w��m=D�@زn�Y�4 Y��k��B��8D�`�$��'LBm[EH�;9^���ׯ;D��hS�W9\Qd�K��F�NVnP�7D�,�v	�r�m��K��}�|��"�7D� �"@�(>��R�AP�"<a��7D�4�sO��&~h���o��0�fI��3D��ڐ�G1(z�a1�KզK�B�1V$.D�Sn��>���ƍ��+����Vb.D����f�8��!k4��7`�a�� ,D�s@��)v>0���a�
=8z���g+D�d
�AW tvtp'�bNI���2D����dD*�`骆IF,y�L�`ì/D���r���5
cI��v>�T�+D�P�Q�	B��e�&�Ėy\VP��b=D��#R�����ǉ֑|\|X��/D�����.a�*��uN�dRdjN9D�|�wm��j�,l��H#C  Чn6D��H��J�=jB8��!�LS�aE�2D���э�>Y�ݰ��	� C�-�E�&D�@�F��K��1+օ7�]҅D+D�0�	�2a
$�6�^�Z-�ld�2D��3�eѺ(2������Z� ��N-D�ti�i	��%8@��XCZ�s".D���@L� *��@oڷGȐ���)D���+M.-(�9��J��Y����E%D��P�σ7}(a����W` �p�#D�qv��C���"�A�.zF�CeL;D�4��A)�"#!�]�h��D�4D��r�� |庴x�b[>
 ��)1D�d�f��I���I�4��``o.D�� R
�<XL��g��&� �&>D� �Y,O�-�� O]ֵ���>D����p��Egʧ{��4�pb<D��b��3`�}#��T� y&�!D�@{���!}��S�;'���8�:D�D�6��!
��ŢJ�x��3�'D��ZcD p�:�A���0�"`7K"D�� @��F�1eM�ZeO
�pg$DZ"O���*F�b�� � m� V�� $"Ot%9P�
=:@��_�@�h[�"O:���	�PXЦOi\8��"O��;g�_�;���VMH�*T�=[S"O����^g��@���35� �v"OL�a�E̚7�('W9.�� s"O8 p0���b�so��viPP�&"OX��T]���9���)�>���"Od�����y;F�0FP�3KZ���"Ovy�#�����@F��`#�0s"O�Q;����?{ l���]�n,`hYG"O���0H��&k�A"O(���J��2�KU���	1"O���x�6��C���,3�"Otv��%F��I�<��|�'"O��R@a��X�D	2'�b��C�"O�I# -8qU�d{�G�$����"O�����@�Jq�,���ƤVy�ͳ�"O���ԭ�Z�~��R��+�"O|��%�ڣ$*j8i��X$��9��"O�Q)C��=B�\��Qě�&yt 3�"O����	�4T���CcV�DP�4�"O�H֧�� k��%B�5�RU��"O�Y����/��3A��%�xp��"O���!H�����3���(���"OjQ�Ѥ�W`֐@�ǚ +��t��"Oa��L�T���ʰ>����"OZ����=D���{1&^1�Pt�d"OL�S6�38�D�Ae���Jkt=Ф"Oh�㤍�ffڱ;��	�^�*�"OR�P#͌�R�IT*K� ;��k�"O\�Ð���S ��)q�Ös<�tb�"O:� $� *#�Z��#r�Śc"O.%�eG,v*��a�z�.���"O�ѕ%��DҜ1� ��t��"O�q��*�&rFvT���7MJ�)'"O����
��RS����DH#���1"O�����E�H���Qʪ�m##"Op����H.93�D�@���s"Oj�O	�W��Qa�Eh��h�S"O`uP4bX	+���)��\4��"OF�I.����M�2�Ё�L�"O(Q"�g��Q���τa��"O�̐ҩ��5/,h�!K�^�.� "O,�j�	�;?��a�!��$ݴ4qu"O�pR􊆶:?ݻ����l�z"O��+�=@�F	�C�� ��-"O�m�U�P�3L�y� �4P��C��8����R�@���j����B�	�^��u`�̏lM�L�#!_6+�rC䉮z����1��5�ڈF+�B䉜9>���ԇ�7v��t+�_�\��B䉵3F�$���F�~�P<��Y���C�I�HFȉ�Z�f�헿J��C�	�$3���s�mn��Y��ɺ�P�=IajIq��"}��#�B�vU���'������<!�����^	���I�m��������Bp�����9%�"~n�)l��C�ԅkD�4*Ƅ�f5�C�	�o�T����+c�Dr�.+O�~�I<fR� ���2w�az�߫*�xR��	�0ҒY�eNߵ�p>Y&-�;x��ڷ�
:�D[*�����L�x��F"O%�rO�EZ�Y���S��I��%Ѳ.���Yp�Yy%��@Ŧ�3��Q�S׼c��ނ9><���C�/��3whL�<� @x[�L\3t6b`q��ƭ(e"��r�g����'�fԂ�O�)KfY�5�,Y�y"�tEf�΂J���#���p<��K�9	 !�b��iP�"]>4n�-�a�õb6��RB0KV�ɍ	�%ӱo�`azb��+�hTC稖�j�9
3�W.����-wЮRtf��Yr<���囌h��)�<ţʻA�@���ĭF�h��G�� ��B�� qS`����� ZNR1�a��<�$p��w�<=�f-Q���$4@��S��[����'�~B߼۳hK�f�4�#L��;�#bP�"�O�)҈� S0�l���0ԫ	�%cХ�х�zǚh� ���ŏ,��d#%���s�#?[���A� BB<�?��/N���D�s�BS�9����!k�lU`��Y��݈�R��bL�/Od�Vc�,KP�z��b�-��Z;gTʈ�a�-��D�"h�mI���
���RUĂn�D�'$6��ǋT�,n8�@��9J�$a���30��'(Fqۑh@,��y�X�v��J��6���bH�v9�
w( /6-J7�QZ�]{}��m�!��K�}8��1�آ��l��*�O�0�5t�j���T�JeN�:�H�w�x�pV��d�ԯ��ɿ�~�	�Q��'���	�H�u���3f]�4�lM����O�qtO�t+ֈ��J��u�f�0��Ձ'�`��t�2�/���N�Z��0ӅG����<�@��I�wI�{�`��R�J����R�
Q%���?�2!��C�5��HM9ȉ?��٢V(��z��'���.�uA��e�ˡT�x�a�{�P�d;���e��v�ָ�'�V5��m>��D�&>�&mx��t��PF/)D���񏕀0n�;�m̧d � �D��V��׿F��tΓr�@�|�'��h��?G�^�
�I¹U�Ԕ��'���H�kIЉ����U#F�p/��O� p�6D�Z3��x�'�4ظ �0bP�%o�]���q�d�;���>4w�� c2-I�l�mLF�;�JW�nr�)�Ɠ��HC�Cvh��$�)���=�KxY��O�ZC�ߺ/��و�L*'���q�n�<�JQ;�>hh�-V/i��EJ��D.����BT�f���'#|�|�'������}��*��MTɰ�'H2��Ҧ�&x>�h���9.�i �d�.e�BgRu��E��I�dό��D�7̲�Ҥ�� ����3n�:A
��ªAp�7m͠C��Mz��@%�����,l�!��+T�h��CP;��s��]7u�O^)[�L�M�D7�,�'Y����f�T� H<�����,ꞈ�ȓ��pH�ț6���zR��,]��H�+��e���IL��~B�.#�Hy K�5!�,p��S��y���?*��遤��'Kx�����?��OOPR��7lO�x`�HI�V�~��&��.� �p��'܄eYT���l�d�[+*�B#��ZGLA��FC�y�)��ɒqӄ��xnu�c�W��(Ox�۳i.����L��i�St�!bN�"X q��"O��!�V�GM�T(��9::��!"O�l�Go��	^x���ӥ3����"O����5�����L�j�����"O�mP1e�td���Q�:(�"O���̝|5��!�˃�!�Q�G"Od}C'k�u�m�c��D�NL�bV7u���
p�Y�9�he[�D�,Dq��'�B�cN�E��d�`CY�#8�!S	�'�F���(0������{!
u2Q��]�*�+��_j@�GP&��yR���,Ɇ�RdY�w_�= eI +��O�,3R�f�aI����B�����$��Å˭%-�#�ş�qH��c	�'A��#-�'
$,S##�!L�p�+O�8�0�f��B�N�.M�`[����O8T����6dH��
Y�����'��ReBZ$a[6�BJS�0�[ԩ��V#�mrv�«&�>�������'%�:O��Si�=���� �D�]ъ��%�'Ж��ɍ��������R�[3L��%�ȹ!݂md]��Δ�0Ď���w�iiU�VwJāh�`�$�&�?��Eկ\Q�q�"�Va�����CiVԼ���N�uf���eQ$u~8�5-$�dyv�W��\�۸Fh�ѡa�<�2�Dj�����W�^]�=�u�ļ)�Fb?��㬚 y��A �F�'3�Z(4D����&G�{��0�Ԋc;�����S�}nx���i	�`fD���(I0��N�N<�C�r}���7�Ǧ��B c<��+�	�|@+J�9M?��9�o��DM��NG5`�����ÎQ�~4�	�S�? ʈ��`-xV��@��D��6\ �'��Q��B�?���`AР3 �4f�� ic�#��]B��
��Pv�<��%� �0���k+.��c/�p�<���I��z��H,��jd�r�<)��<� L!�_$����r�Pm�<Q@�=N�f�1����q:��x�`���s�#�$"���'��9*W�һy�V�ҁ�ȹ��'R�T�&%�'z����1��8��a�y"���	��Ib�e�O�$��e�]�(�T�s6�\�Xn �
�'����&�E���5)E<T�M�'���|gH�Q,ORyT�?�3}R�Q�6hyK�圹f�TUJ��˛��x���-\�uУd7�����I�9`����bE�8@F�Q3�'�*4����t�rÐ58��Kϓ	�z��C�6>��[�'蚨�h_�$'��� �#$��li�'�f�9 D &8��ȗ�^�q�!�L>��cޱ~��t��������葢�J��`�!M\;�\�2"Oޘ�h��2hպ�L�+B�[�b��n��e�V�� �.\I�g�UFP(����x����"��y�񄈛K�����7�N�[�%K�1̨��/Ѩ}��I�4�OФCӪٸ�4�U��2A�|�r�'� �%C�41F�h�b<O�A��CG�
V��5PPm1�"O��#!؂`�����͋��ppc�$M���dX3�M.���:u	"��~V@�I�m ����&"O��3���>e�V�!>��2�Y=B��d$� ��<y�hY�? U@d��.uµ���w�<!�B�F9��L�/0��اcF�<�GQ�4���FJҭ/��1�ĦKh�<Q�O	N6��A�$ !:���ef�<��䝄N��ÀP�Q��^]�<)beE"ȴm��ҿUH�t�g
�s�<s�L*? ����߮?��q�u��j�<Y�"�u�\�[�ʨ����KI�<�@[�]�Q�E�/�  �m�@�<�ǔ8PXp�/��-@�gl_U�<!t�V<�x8�ᄸ69��k�F�S�<٠J�<!t^�[�/,H`b3+�M�<��!ŏi��ò��	b��Y�g�J�<��!�4)�]{e�Yw�M�E��M�<ٴ�%}����lB��ʆ��M�<�&mۮ@�Ǧ�%;����mVf�<��i/"̩�eu��Y6
\�<Y��V-\E��FM�&Q9��G�<%'�2м9YWG�		�Ա4�Fi�<A�a�S���&�;ʺ�yF
�e�<I��O #ˀ���Æ�Y��i4�i�<�Gʊ"g@| � cN�	Dy�BAe�<�v-Ѧ#��Cgg@��=�fF�e�<��T�{�,�qr욯/���V��b�<�H� ���j@/G��I�U/Oa�<1�I�R�<Uѣ��'N��)�M�]�<� �=;��C�E!Ri�!%�X�<�eꇵK���HD�I�VO�aj7��_�<�g�C(3��iL=]����E,D��qD�D�M-�
�)�U4Ph0� D��1�V"D�@#��T�a�����I�$6~:Gͷe�Pia&(<LO��k�
th0�'�o��"O�)��� P�S�U�h�r�"OhU�w �3��x���P���A"O����s�� )�(8� ,y�"O�! ���6{�\j�Hڌ<��ib�"Obؘ � w�12$�����j�"O�qqe��+9.�dD���
��Ղ"O��!� ��'��H�&�];�p��?Or�'�t���ܞ"�Ή 5���u�ЍR�A���9�$ _�.;�l�*��'A~�� ̐r��S�g�? ,X��ƨOߔ�B%��;�YB��E?�V�Qo��w�R�0|jDK�b�)r�"�#I�����Ʀm�BL�E/X y4	 }��)�'����:|{�)Ӆ��	I{ta6\�W[^�˧gܲ]I(���gW榅#��O|�Q�NM&-���C�ވXx�#�ǘ�5��`��B�ئ�@y��Ocq�f��"�>���s��ʉt|��7H�9 �u�'&x��
�`>����L2d���ࠋ�u����e��j~���c�&-+�$��I��"��L�d�uU�A`����D�	���r�,�)ʧj��[D ϐ8��x�j�]BlL�	=E��}���^�4$	�&ȎI��I���@&9&��`l#�@B�b�'p�����<�J�o=D�D�Q";n��
��W��$���g8D�hȧi�#dŬy�U���E�<�S!9D�4���7k�J@�ň�^&$�{2c4D��S��M&�r(`�A�`�Y��=D��@�Ӧj��TC�G1kd����:D�`�h[892��E�mV
��1A7D�L�sN
���sJ����%�ǡ'D�����W[���H �U��I3��$D���g�ӗЭy�&��"�����7D��Cqǘ5d(\�E��(&�)�t�9D��"�i�)3��Ɋ��W�'�N�(U%4D�\*�DB$PQ1�
j$J�	a�2D�|�w�J4n�ГDR9��`��1D�la6k&�x=�3cR%6�+�C1D�8�gO�z+8���J9"ވ�c�3D�l��n�L���#��;g�`2i$D�x9e�ض�.3��G,wôԘ�,$D�����Ơ6���WM�$ex��#�!D�ܫ�.��N��|�B!�"(�a%D���i�2h7,� �W�xV�@e�#D����	��g�e
��#};�pq �!D���lA!_m�|����"D��� #D�Ty��9� ���"�&%4����"D�l����zڑ�5�C2a�4�E� D��'IЧ1O�p����)�h��f,$D��[�Պ*�0���Ț?A��R��"D������i��hֆ�)i@4��� D��;��K6n9��@�BHyl���:D����F_���M�o[�~�<���9D�<+�F�",��� bX0����Ħ9D�t���H:&]�,J��&o@�)�Ј"D����+'S)�Ed��;��� Q�$D�hqǋ����D$�/~Nt���k6D������Y@���i�3R�4A���4D����c�ZfV0�$g��H
p�4D��k��Bp]��)����&���k1D�h�:�4h_6Ch;��2D�H D��s���z�Ǜ�H�Q��$D���CcN7J�Y#��,�z�H4�$D��pr�9k�p(і�5΢�B5D�$�dFP�\�$��� )@b�p�E'D�����+N�DN�"N�xP6�"D���@-�k���hD�I���Sa%T�xR�&Zsv�Q�ˉV5���4"O�����0OT-��C��֔cT"OB�s�mLhY�����O4Hy��"O,}��I^Bf�X"�ڬ1S�!�v"O���7�Z����T鄑=<J�@w"Oh������ 8�k$�'	/��z"O`%�WELz���
��ƴHK�"O�-��K�1�<4�0)Yx�jp�B"O�� 
�54�p���E7Ux 	7"O>i����r��}���N+����"O�i�#��,~�y�"جC�"O� 0uH�n�-Y��8e.�#�(ݹ�"O<�b�W�S�.�[��އzjz���"O�-����<$��\[�9��"Opx3���H0,ps�oP�M�B�V"O�}{Rĝ� �j�9ro �5��x�"OH�S � %�&�9�CS�g͚���"O�]TᖥL;}��Q�Q��)��"O
�h�G�5 ��+�׶�(� �"Odm	�Xw�����Y#�v�kG"O��+ޞF�`���언y�X�y!"O�ŊtFʝK�	a�k@N��y��"O@��(d!�@��
t~:Ar"O���pdX�{H���ϗt�}��"O�j����Ih�Ң��8��Ã"O��@�Id���S>]ީ�Q"Ox\{EǯL@�W^�fRx�r"O�t�ӥVm����T�5zA|��"O�Lx��.X��%�5@�I5"Or�u�176`�XÀ�YH�÷"O$����O�P��N�&X�R�"O��㍘-,��Z�ٴ&��$"OLp0�
MR����q���"O�y���B8dq���6
�Vi�"O�z7���K4v(  ���n�z�"O�����RR�ƀ#Q�G22� q�3"OVMFHD��s�T)Y�����"O�=�`�,}ܨp�������"O��+w�2
X������$h�"OlI
1G�P�*�� .Q��/D!��ۿ�"<���8Cf6XЌ�8k�!��1pR�L�D*�(J�Hv��G!��<W��2l28�����q,!�č�NW��C`C9�\1�M�3!�Q�D��6���]��[�"X&(�!�ć;u-�E���iI�mq���t�!�O�xx��E��c<Ό����/iq!����\����>_*v�[&gɇbW!�dW- �|x1s�G�@b�"�N!��ڑ~�`F�Z�X{ejC�3!�ڹR��,z҃�gL��(c!��5M��@���h���#N!�,vL\���n 蠡c�[(!�%e�I3�o��8�1�*��!򤍸jt����W��EA�o�K�!�$Z�tP�g��3�p��wlM�6w!�$��m�\��� Ŗ����!�$�"Bd�\q��G0b�4����&$R!�D+dI>�3wK˰|�L��JH!�$ή)����� ��������ȩd*!�D�̈́���
)5�>��j�. !���o֮]�W�H}q����ִD�!���=?�&�#m]��ڨ1�(R�|!�ݴ2Dp��eU/O��9��'�%{!�c�����dޛT��ʧeJ�h�!�8*t�)��)چ$D24��Y�B�!��$~"��Y��U$)�:�He��]�!��^.-h����/^�=�����N�E�!�S2�܂��)yP��X��d�!�d֨c����`JC9O�0�`,!@!�D�.��! P�F�)�(�#&��!�D�?J6��A��d��X1�V�r�!��.LJ>���Aj�q�����!�D�r��(��Z�uȸ$�"lY�7$!�$O�(G%��`�&�0�<!�� `��*q>B,��a�&"X�q"O9��@{��#y|�S"ON��p��)R��A�J;]�)#�"O�<����S�����֑p,�G"OPX��fDK>TTխ(Н�A"O���ȫf@��I�X�Z��M�7"O�mSP�h�d$��`���8�"Ol�1cl!?
�C�J:8u佲�"O���c�x� Y�hK�� y"O�zB�%ȦMS�HS#ch�xz�"OV0�cJQ	���bUHƂee"O��z7HI�)�zЫ�Â	3K�E�"OV4�� hq�'�Ł?D�A "O��l��:����%M\	~�:�y�"Oj���N
IA(�ZuF��Q�tԨ�"O�,�4@!(l���A/�ΐ��"O�x�朑4��@�Dؿ;��S"O���P��/c��a�#��K�L��"O� v�ٝ߼w��o2l#�"O|`	b�ߩV'%;�F�~���"O̴�v	KT�6�g�=n4@�S"O�EH����Ps��ב�d��e"O&�B�cF �r��͘w���K�"O�x
f ��oX��юV�}	�ݠ#"O� q$�t�x��-A&x�$�
"O���"�ӯ^<�� ,ˆo��\y"O}qtd܍?0���sKؚz�v��U"O,	cOS+&��غa��2V�03�"Op�A1E}i8Qr��oQ`�ҵ"O�d�u�$q$���gX6 ���k"O���bn�XVx�0�N|�P��"Ox���%=����ŗ�L~lu�A"Od��a,�����䞮p��Pp�"O��9@��]h]�Ff5�j���"O6��q �C���2��
��T�"O>e�T�L)�<�1��I���$"O����"��=��!�pዊ��=*�"O�E �Y��PCOK�xv�c3"O­�B��. n�yq��b`��"O*Q9wB��!C��p��OGO��zE"OP���HR�s̲��"ь+�R��U"O� ��
lؔ1��k�r9��"O�ts누2&��SB̨l%Hu��"O�L�Pq�d�B��fÖ�37"O�]�$�ŚU���I-�@��h@"O ԪgĞ,H��3�FM�Z�"�z�"Oʼ������bF����#"Ol��2o�y4������?n�0��""O����z@�٦��e�����"O���Q�
S
,���\��}�A"Of�k�H
6�a8�!A�$�@"O�X����e|T�a� [����"OV�����+Z��)"�hS�NM(S�"O.�'[.R2n-Bǈ2jE�d"ONXj��I X���� ��4\�dq�"O�{@�̙~>���ĉ%q]�C�"O�LC���>ys��x�-\t��t"O� �:*F:e��Ֆ<r���"O�ț�$���ԉ�D�H=a7"O~D�C���v}�mC�HD�b�
�
d"O�� V%cBt����*�V"O��f�&u�����b���0�"O�!��8���
9����"O�K�̆fp�#��T9c����"O� 
�H�gɢ)�ȣG�v�̘S"O��ઋY�<�x�	���a�T"O���b Ϣ��q@Cfr�(��G"O|�����j2ѐ���!s���w"O,��F �T�����:l��r"O��{��J�QtD�Vc��D8Z-X�"O
9�S�3C`��3��U��ԣC"O��`�� �yY��WLiU"Ox+m��Dzڍ��/'4��"Oʼ5�*�*,!7��*d
��@"O`���d�x�(��D�&Èx�"O4��r�3��҅F��~�l�`7"O�4ɆE�n@h�'%��R}X&"O�9���:�^,��X��	 "O�3��2}�xQ�����"Oh�ѦHم;d� 	�eg$���"O>���}E�8 1FTRB"ODq:�__�X��1�0hi<�17"O�y���p���Q'r\b5��"O.�Ӆ�*5����&�:���)�"O�I��   ��   �  �  �    �*  �5  A  ML  dW  �b  Fn  �y  ,�  G�  ��  Z�  ϧ  �  w�  ��  ��  >�  ��  S�  ��   �  P�  ��  1�  ��  �  ( i $  k! + �4 �; �C M �T �[ �a h �i  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C�d �S�)U=w*����R�|cC��<H!�D�0@3�qJbʌ�h��K��I+ 7!�$O}_�%��h��F�h��d�S�0!�d��K�X�a�R9����Z��	A��H�d�ɀ�XfΪ܉�T�θ��"O8 ��)}�!pk\�'6.q�f�|R�,|O�Xѷ�������fE/��0��x2���&?-yN~J�ݩzGd�bp� E ��Q�
U\�<�������Q�ae�&
�� ��_ߦ��Ol �C������禡��b�3\����퐀h�މa�".D�$#!EL��8�0�R(n����>!�S�ԛ���3K�tI:�-�n;�q��>L��H��S{�@q�̴zn@`��JQ3m�v��ȓ	f
H�@��?%��q��V-L�V�ȓ��ґ�=�ޝv(^)���ȓ=\���wnX5o������&:��D��h�JQ���C:n�cn [���ȓ-�<s$��x����b$�F��O�7�*|Of����46`u#��
�����' �ɴXBDx���<WW�={V���KنB䉻���%13q��B���h�>i��	ڪ'�n��)\դ�B�d�/!���R��:1*  �#T�8��K��h����)Z n��1��ăQRD��"O�p@�� �K]�-)������<k�"O� �m� }�X܋�-�)c�T7"O^�!vB΋�����>#���Q"O� ��=tiztk��-g���"O�0��eLx��p(�G�~S&ȫ�"O���Am�N�d�R� i�`�"O$@�Jǀ\0Y�`�� =Y�� �"Op��#	8��Xc�e�䰸"O��x$��3��|�уSP�L��"OJe�����I|�0�4�3>��-;$"O�`�F)t�b5+'b�?��DjF"O8���������c�#C��`��"O�qB)�3"�f�9R����8a�"O�X�)7��0�g ��q�< :"O�YZ�׋i��zɎ5Yq��§"O�-�� �y"nta��be��5"O
]�ŉ�#x�R!Fa:�{�"O� �饊\2^�����J�cH��4"O��p@HH�s,�E�1B�!i�"O�ݫ2�� l�pi�!��~*DM�"O��;�U%�l�+n�1�6��"O��%�S�6����LN�o��{�"O���'�09k�8Xp�nF���"O�4�Ty�T�� 6x5Х�C"O��S��D���]� 3d��"On�H%�F�L�j�z�.߈w"��J`"O�Y�gJ"���E�U��Q��"Od���G�1�f�3��]%� ��$"O ,� )��zGLy�ѩW x���w"O�E�É�I���p���x�yv"O\���a\�Zn��!�.�-9�"Ohc�@�VLR��5h.2�9�*O
���<�8��t�[&��\�	�'�2� �S�0ȓ��˄r�L�
�' x�J�|�xԦ3~	��'Wl�9��I��h�����i�V�z�'�D/�3<���GT9*��hQ�'��p�ƍ'�^x�����(�t�q�'��� ��*7F��AI֮'(���'x����`Y�K�p��
P����'*t,x�.G�V�RljsC����Y	�'�f(A�0��8p��S<tdz��	�'%Tl;a��>$s��Gj�8s�����'�x3d$�*%~�	Rŏ�5�j}�
�'r�1���ty2-����)����	�'9|ɥ��GnZ5�`JA=	|�	�'馴xwl��)t&��W �7$��2�'��@��I��Y3~h��h�	�R��
�'�̘�4�E@�����/��1�	�'�P��ӬZ*%���E��#wLY{�'��bkZ�}�|D�#�@!@A!�'��84	�̸���%������'�T ��*�d�0/X/��2
�':������Z���y�/ҍG <�	�'7B�f�;A���h�m��D��	�'�N���N݋Ei����h,C �U�'Ɇd�VӼ5yX�B�D�H|��'�Y���?�<@�I�;�ZA�	�'��l���Δ�z�Mۤ�R��	�'Mޅ��F� N�(�R���[pE��'ڽa7CG3���ϓeF:�	�'��(�`	 d�T �C%5҂�K�'���G�7N��3C��&x�X���'9x�b��9[����S/?u��� �'�j��� X:V�Hè-t�0 ��'�,��"	�Q�X�����!����'���H'B��a� ���0��'���0��� GJ����I4e���'�@X��_-U�h�"��5AX����'܈���@��.���\!@j*}��',��#&�? ���"d�41��R�'"���u �)N:�˔(���B
�'?�H�$;�Xad�����	�'���1�!�5Sδݐ�Ɯ��Bh)�'�e§��5��8BtmI�����'�hp�O��C�vȁ������
�'xT�DR:p�����x�!�
�')5����J�k���p�^��
�'nP�#5f��%�� �"ɘ`��	�'z�|7�ϛ@/�(�A�9W�8�H
�'A���H�0h�p�`�#R>�,;��� N�)uj�+�ļ�㍙��*�0F"O�YY�GKh��Hq�_�1�r�9�"OdE��Swb�Tհwf�8�"O���j@�fj"��:g#�"O���KG�N表��49P@��%�'?"�']R�'���'I�'Z��'1h5x3��Z^��B�	bW��r�'�r�'�"�'���'L"�']��'s�)M���Q����6Ċ����'���'���'Y�'���'fB�'�xxK�� {��pO��
D���'�R�'�B�'��'���'^2�'��$�!������am��"�'�R�'���'���'nr�'g��'r��+Êd�([��Z�&��xS�'�B�'>�'���'"�'���'{@-�%�J\���l^E����'�r�'��'���'|��'O��'S����K�!����"�W�q��3V�'J��'�B�'R�'�B�'�b�'F�e��AK�g�zD�0NG�`�`��0�'�"�'���'("�'�2�'+��'<h����Ky�-�c�&<�Q�'��'�B�'$��'[��'���'��$c�V�L�3��"u��Z��'��' r�'���'���'"�'4�8�m���e��Y�L8��KP�'�2�'*��'R�'�r�'2��'����# �#c1dypd�)O�d���'}��'�Z.���'x��'i:6��O�����%�ΑW�Bha���@��S�%�<�����P۴&0P��F� '>
d7H˂�fm��&���M����y��'�aJ ���sN9ys�	x�.���'�����E4?I�O����+���?��@H�1,6E�&�K�'-2^��F�i��gǒ�"��V�/n�)�t.�5 �^7�L�~�1O"�?�@������͎0y�!3`�`fh�����?	���yBV�b>�$��̦U�h| �"a���hH^ql�y��y���O����4���d?Z+��r� ���F�tT�$�<�O>�Ծi�ę�y¯��s���K�kX�|)	�+�#��O��'���'<�D�>pm�>bx���t��8�%��"@~r�'������O���I)⎏�/�f�:��=n�X�G�*��by�����	�a�TA(��Q
�|��KO�qN��Ϧ�(:?!��i��O�	Q�Yz���E)�*�����
ߧx���O�$�Od�	x�P���	��d���(J����آ联Ee,Ez�C�����4�V�d�OR���O|���{>���#�^��9U%�>&��j<��,;*zR�'O��t�'6�T�w�6&���s��9}*�{���>yg�i��6�.��G�s�-����i� ɑP�!7A<d���XI}���e�r ��f���]��� ��"oz�q�b⛛Wt5/P8a�. ���Iȟ������S^yb*p�^A( �O�!CE	�3�U��ka6�K����̦}�?�6R�`�I��`�I+3�l���Ņ�4�J<�B`C�˓�c��7�/?	c�RQg��I*�D�pݥ�ݹj�x\Cb۰s��irq`�OJ������	��,�I���Ic�'U|�T!a�1A�H ˓,)J"5K��?q��囦��7f���M�I>G�!k"r�;�'M._$��	�N���%�d��ɘ��6m=?G���2�U�lѡA��)���>l��I0��O,O��o�Ay�O��'/ҩ��On\dᶎT;"�Wd]%�r�'��I��M�4��'�?1��?y*�����
�7t�XC���渂E����Of�nڬ�M�N>�Ow8��Rf�$Y������&�$�a�Å+��qQA=��dNǺC���O��.O�n�#���@�a`�N�L�&�D�O���Ox��ɥ<�3�iȈg��i���1���g���� K]p5��8�M#��>��O�,���k����O/*4�}���?�u�^�M{�OyZ&����K?U���ǋ
\m����N���EW4�M[)O��d�O:�$�O.���O��'/�Xi�)�HO��P后6I�����iMn�r1�'��'X��y
k��nW�D���`"�[<&S�I�+.�ao��M�L>�|��N/�M�'݌ a�
�BI
�pa���{���9�'��0+$�Pɟл�[�ܪ�4��4����O41?PA�@�*7r�8$ F�O�`�D�O���O��g<��� �9&��'<�"��E5��v��e�Z4�&ʚ "�O��'�r�'��'Rr%�d�'JR�ܪ�ʓl�@��O�8T��; �r��U��XyZw���	�BS�/$����=)�9;�iҴ7(��'Fr�'�����P�PB������O�2jje#u�֟0
�4Q�j@.O0)lZc�Ӽ����4#2��ra*�9F��W[����O����O���תa��B��MSA���M��+]0?�NՉ��N�mv���FS���Ҧ}���d�'�r�'7��'̴��O�=#)�ͪkX VhHH�1U����4,m��Z���?�����<i�Ұ)	B��12�.���X� A������	M�)��i��qy��˫W��]�Q"�$�"m���D�'2�!I�E�$��Op<p-O� mey2�CT� �1Pk��~����Sa��h��'���'�O��	��M����?I��Y;9~�a�Ϝ-�2�6��?��iH�OX��'� 7-Cݦ��O�l�@������$X~�p�`�����<�R ���='�����L�Ov�}�=� �xAQ�ɜ~�F�(�n�q�4!#�8O��$�O���O����O`�?��F߬]C���E� �f]A��ɟ�����,aشS�V�'�?1�iO�'�$�K�̆^a��4H*Pen��ę|2�'��O/�b'�i���%	�ҍ
Ag�,!�9�v�մc�
�����,p��<!Ǳi������	��4��F�Fq���Y��R� ���+�t�����0�'l�6͔������Of�d�|*��L3s���s�S$7[���#�@R~�˪>����?iO>�OY���'��H���r8���ޞ;�(���i��*��N@�~X���&x���AQ*o�}
�!�$QR��	ğL�	쟴�)�iyr�{ӪL@�N�\R�y�m�J9����e�~�d�OflmZ_��J�Iݟ�1�b w�*A!��؁`MN�kb����\�ɋ�XImZ]~b�]�JDJ�������]��)�A��f��Q��	C�Z-mzy"�'s��'���'��U>qH���uDh*N@
`*������M��M҈�?���?����h���͔/k�����/	ﶼ(p�Y�M+\���Oz�O1�N�hs���I�yQ�!����1��a\�o���	�b�}IP�OPʓ0ě�U�������s�E6�hȊ���*�p0c�N��\�	���Cy�h�HS���O�$�O���֣٫�M��e�OҲ@��]�n���dl�L�	$�&�z2lK?��A7���"��0�#ȋ8�M�T� �Xwdi���?!�Fڻd�Z�9҇Q�3����!���?���?����?���)�O.9�%΋�dU��ati��"2^���o�O6�l�#,9�I�l��4���yn��g�9��ԔJ��Jqo� �yr�'�2�'�(���iq���F�R��gП�`�pƛ�8K��x�H�$@s�HhBh�<�"�i�Ο��	џ���ܟ�	��J��r�L<��@� GM�J���'�P6�	xk��?�O~����:8�����!��Q0g?8�w\� �IΦ�<%?I�ɂۢUa�BL�6��<H�ٱ��lڠ��d �hϬYh�'T剃�M�.O� rElE�A~�l�2
ЪN�l<����O���Or��O�I�<�w�iH|�J�'��T"�M�/'#Tk�O�\h���'f7!��4��D�O^6��O��3����:��� h�3�8m����r�n7�4?�%�.����hyIk�)���P��SBD+t�@�į�"Hq��I�����x�	��P��z�'D9<h4����ܹd��CWJ�R��?��o�v�:_���6�M�N>D ��W�l�!^gB�!��,@�'<�6��Ŧ�ӵJ���m��<�B�,C��R��S>�=�	��S�R��僘�&�f�#�����	�<N�Iڟ�����h�	���G��(J����OV$���䟐�')��D+'��I����O�؀o�3<V�Ѱw��X�x���O4Y�'kR�'�pO���7z�����SX�BX��R7��P{���d�h>?�����E��Ӽ[���F�̼�fI�g����@��?Q��?���?�|�.ONLl�(���Ύ]���h�h�+��#s��iy��g�Z㟐h)O�6͟/�d ��L�4!v)ZU%â:C��n��MS�	�M;�Od,C��T�
M?%��k�3&�\��c/N$.��tC5��'�Mk.O �$�O��$�Oj���O4˧'����R�-7(9�7�+�0���i��e��'���'���y�Iz��N�@�(���z}R��"�/ĔoZ(�M#s�x���)Ȩ/�V5O q���mB�)��7#�?OtZ���?A1��<���i��i>Q�I�p;���ч^���[�@t��q��۟h�I��t�'#�6M1Rl����O �D�	r����� eRp\�ΝR��㟈x�O��l��M�A�x�.�3#��\�uB=�3dH�����R:z���+�",d�I��u�j^��H!��'8������9�8=24A6@R����'Z�'V�'}�>���	L�����HP�E��&��j��I�M�����D�����?�;d�@{�e��xhR�	��õ4[͓�?���AX����8��&�����Z-��� �̼YB�Ve�&E�uŒW�H�'�7M�<ͧ�?1��?q���?�%�ĤdPa�b)�K*ްǨ�>����=�"�U����I�P%?�	�l�Tp�C)�T���ϕ�0C�O��D�O��$�b>y�+B�l�i��I0 v�Ԫ%g�'��0�f�;?	EK�0DN�������V�-�'�
i�e�51���J�/M'�,HW�'�B�'�2���$]��*ڴ}����W�i��'�]���ҨBD�}�.n����_}ҁqӐ�oZ��M�SM̐+�Jk2�S�Ҥ���"�5[ȥ�ٴ���S�Lr�P;����S"�u��w�2,zG�,Y����: 	y�'p��'_��'�r�'�]2��yV(��݅w�@��n�Oz���OJ�l�8�E�'g$64��M�?��%Z�H�R	�0���ʞd��($�$k�4jz��OfT���i[���/ށ�E�E���!��^5]hεJ��_�_Q�oZby�e���S��O�]ȗ�T�J�HLz6@�2<)V�*v�ɹ�Mk	����OD�'
-ᤏ�!`��`�А��X�'x듫?Q���S���5D6m�c)�#L:�rI9?��0B�h]�X�R6T�擧t��H�B�ɐfN����b�y��p!"���c�C�Ƀ�M�GA�9�\����ܫu��X4FˬA��+Ȏm�`�u����8��ۢ[|�H�p���B�{娙ß$�	<L�m�\~Zw&�� �O�B���� x|jO8�`�"�z\�C9O�ʓ�?��?���?������T�%葠�MBd?���!	���UlQ��Y�'�B��T�',�6=�%2wGQ9=U(��Eh�+#���T��O���"��I�23�.6�p�p���p�2L�3�L�~0��x�@
�+��:�b��ay��'ҏ¨Jy���%��-[�e��Ё-��'L"�',�	�M�7#���?A��?q@I�9E�[Q�E�(�v�c-	9��'��듉?Y����E�hu�K�E� z��X�Q ^|�'�\@�D�Ně�l8�I�8�~��'��� ��-c�Ȅ����N8X��'1B�'�2�'�>�]�^ꄺ!Ȃ4.�ڱ�e�9.`5�I��M�Ն��?���f>���4�"�@("���V����e18O����O^�Ė���67?q�&�'~X���_�Ѕ�HT!��.O�\�$�4�'��'Jr�'��'�n�"�@|��e�6"�� c]�T��4?�����?!�����?q`�L�0�pE� 	�v��h"���a'��ԟ���Q�)�%E��d�0��"obR���l�r�*W�̦].O�`3�k��~��|�[�@q��_��>q&��4�,��%\ҟ���֟,�	��\yraӀ�� N�OdDr���'8�����[!r@�HX�?O�<n\�L��Iǟd��͟�cǡO�D}p)��J�/�䉴�7P�|l�z~�'�&l��e��]�'���t�LMS��e"�]��@bƌ�<���?��?9������q���7�N�/,I�V�O<��O����ۦ�[%� Gy�vӴ�ON�B�"��0,��Ta@� q�n4�d�O��4���Y��gӎ�R���aAϴEΰЙ�	�у2��4��D
�䓕�4�l���On�����̣������BN��nD�D�O,�_қ&BЦ{Gr�'�2_>�aI Bf��l�x���fd(?Y'[�<�	؟&��'��#B���8�4A���./A����1? ���4*�i>�Q@�OƒOfx�b&I��!�F/� ��U���O����O>���O1�˓?��voQ�N��u!�K�m�@��S-�5Wt����'��!vӺ�\�On��S�<��hJP��(!g�U�g��~��d�On�U�w�T�=��T�7ʨ?͔'�V��1�<U�B�\F���@�'F�I͟��I��p�	П��Im�d��z�f���O�qXC������6W Qv����O(��?���O�Tlzޡ1����HhJ��[�#�<�s�e��Ia�)�Ӱ1�*TnZ�<�*P�[��\y���;z��M���F�<���ƕLI���G��fy��'�b�ɻ.�R���%~�b��جU��'O�'9�I��M;���?����?��J��K��<��@Un�j4�iK��'v �[��&aӨ�&��+F���Vl9eK�[�|ᓯ*?�rJ�4a�����A̧9e��$߁�?9��T�^N8��\b�ut�� �?I��?A��?���)�O�`auA �(��0�.F�?p\�w�O�@l�	3��ɔ'��6�)�i�قvK��B_��#�kܽ[��d*�e��:ܴ.F���v��D���x� �}� ���FI�D�\�&Cc��5tN0y�䀐����4����Or���O�䌨RՀ̀tǢ6���)֏
N�:�������O`�?�ҥ�:-���..�\�q�*��z����'v��'�ɧ�O�R�	���A�,Q�׊D�L�����2$�����O��!�=�?9m5�ĵ<��lX$�3gfR7�D4�%����?Q���?����?�'��$�妝C�Ɵ����F����s�=	��h���f���4��'H��?���?Q�k�r�zlxƃG�a4�`��� y � �ܴ��D g�<������O�W�H=d0�� ���92jȡ�y�'[b�'�B�'B�����	�	I9Lhd	��V�h�0��)Oh���؟�R�?��ڴ��Bn�͡�ָC�"!��F[9}�`	L>���?�'b0��4���Rs�u��j�*Z=�Mqc�G�.��R�D�?��C?��<ͧ�?9��?�Ҭ6��rFgP�;L� �̉�?)���������/	ȟl��ޟ4�O;���7�ݜn���"��	q�l��'�"̴>����?�O>�OG$<!$fܼL9�a��'�-F��#���k���,�<ͧD���	N�	&30����a���a�op��A��� ��̟ �)��IyB�a�@ę��n��s�ܧ$-a�	����$�O�8n�f����OP�D c���,O��d����S�&ܤ���O��耎|��.?=kC��?]��e�7*m�� 5��w���<�*O���� <@��\��G[(R�R�diJk��po	��|�	�|��B��O,��w��c���1v"}a�ܲFK.�I��'AB�|��TɖH���?O|ԣ0mU�+���i� !�8y�8OT������~b�|�Q��'ZruiQNԣuanq
N�"<�ÓT���!F'���՟ �KV����=  ��HR�b��I��\��U��'z k�D�pb�v���-���Y=T�x�B@&3[R��N~����OF����gG�e�&W� ��D@���� ����?����?Q��h����W�6������5�Z�AĂ�E�d�dHԦQ�D��Ky"�qӎ��]7[$R�ËP!'!"f�z����T�	����Ϧ��'��PYD�^�?�H	� Je�DOL�G �Q�ҸZ�$�{�4��<ͧ�?����?���?��A�1F��[��ͼ,����
E=���Hզ%���������۟ $?��I4����"�I�̎H�YIt��O����OڒO1�F�sc�P��])"�
48���W��O@AQe��tA�܉��Zr��Hyb'��`p� K�	���i�'L��'�O��ɩ�M3ǐ��?�ac< "�qBŅ�<zdc�@>�?6�iJ�O��'E��'6R�� �A��Qgj�÷��3~�e+r�H�M��O��Y�Mŵ�z��4�wp�a#����\	Q���S's)�(Ә'���'���'%��'\�,�pl�9 Δ%a�-�4*y�:@�O.���O��o���$�'�6�9����dM�ic�Fz
��'޻��,$��I̟�7��PlJ~rG��&*ZD���T�C�l���JC�������(9D�|�S��S�����ß<��e��V��xBC�$Y�d۟��Ay��i�h)�&Ǹ<A����I�P���,����֭*�I�����O��D)��?�	w�әx�X�Kq��q�p'<-�b���I
*O�I��~��|RNY��x�;��XD��3�S�~��'�b�'c��t_��2�408T�Ʌ,�=/��G$�
-x�Õ E�?���U����Q}��'I����|����s'���h��'��9
�֕���<>n�i�<���E�xZ�t9B���b/(�a�M
�<�/O��$�O����O.�$�O8˧n�����cal{� ��Nh��#�i����"�'�'5�O%o���@g�<qcHS�j���JӅ?
���d�O0�O1��,[�CsӺ��=V�U�s��(aH,���ɵ!�.��A�'��'���'��'��<id�Jq��d�s�̬(]x��2�'�"�'��P�0��4�����?q��l�zN�"T-�X	&
,fyq����>y��?M>1a)�]�عh`�֪�r]�$�c~���U@�Y:NX;on�OU�E��9o'�g�Qi��*��!GJ�
A�$aX��'���'���ޟ��V��U�Π"T���0<Q2�۟�;�4hy���?i�i��O�Ԙ)wtQRT�d��-�c*O-��D�O<���O���d�J�Ӻ#a�ͭ��r�S�Thp#���+�6�5��(Ю�O<��?���?����?���8����J	��P4�%H,��H(O��l�81b,U�	x�Ig������DI�G��1`��Cn�,E饦1����O�d*����`&d5iB��3�x#�fL3L|�41��m���'b�a�ӆ�h?�O>y+O&��� tX(���	7_�M����Od�D�O���O�<9��i���x�'�(�CDNY�D� �h��9*J�I�'$�7m8�	:����Ŧ�i�4G��V'ID�U�����4�b��A
� E�� �4�i��I(\7�ir�O�q����.7�Xı�J�yq���VB��E���O����O8�$�O��S�'~
�(��Q�I�D\y�"ȭlR<:���?���" �b�G$�ɗ�MJ>���[@s$��F̊�3k�a��ћ?��'hұ����|7�Ɵ��a�&�"�t�x�g�;K�{Z|�C@e�?q[~�'f�i>e��������L��ə/ȸY^Tr�G�+1�ܭ��۟ؖ'�6m�*8��ʓ�?)-������^�<��G�P�DK��0��H#�O8���O��O��7,b��u��z���E�~�4y�&Vl�Ĭn���4�(d��'��'R(eY���D�1��p<����'3��'`"�O1��Mc��s�H�J��L�qm̫�@ h�����?��iS�O޵�'��&�Fq�$�pC��u|�zr�8K.2�'ʊ�ꗿi���?I(��%ԟ^˓|i�EB�&�o~9��^�$�͓����OJ�D�O`���O���|J�S�dZlB@M�31��uBꄚ曖CM�'LR���'�j7=�$I�v(��n̹�a[�tip���E�O���<��)�TF|7a�Ԩ'�T�p�$��HX�Q�Qg���L:��	QC�Ey�P��S��T�sZ܅��%���*OR-oZ�Y�b�'��D���j��`#��H%�u0��ӈ%B�O�<�'{b�''�'޺eҐ*ԅJ��c7�֦p��y�O�5Y�N��f�~���2�I�?����OVr�����)����5m� A3��O��D�Oj��O�}r�IG���f�$h^�Yc�b�0-s�����hD�/�k���'^�6�;�i�mp�dI�9��8�Fװ0e��@�q�$�I�,���W	�MnZF~�,L+?R8�S�%[�Т���,<n�I�5OĬ ���餕|r_���������4��ߟ�K�L�)o�4;ǠԡHܶ�)Smyhy�n���E�Oh��O���l��	EKn��=n?�Z��Ǫ-����'���'7ɧ�O�l��!�J�-Z�I�ae��fY�G&K!F[��H�OP��O��?I�`+�d�<�0�qN*0k�jϝF�@Ā��?y���?���?�'��D�ڦYX���ǟ�2Bb *g���i��d�Bt� n����4��'�X��?����?��gZWJ�t)�ږ@����b�l���!۴��DG� �N��' ]Z��j��M�FKdYS�M�>/�-�&��=S�d�O����O����O��D,�S�l	�ԅP�~���W����	Пl�I��Mk1�ӻ��d증$�𱖧�T�E���8@݄rի����&6-���S�v��im�[~��ڈ�� ���v�<�I��������LB�?'�3��<ͧ�?1��?a�o�0(Dd��3���Y��02a���?����D�Φ�in�ş����O-z� RM�$#q�RN>S|ys�OzA�'��'�ɧ����i�(�a�ǲ9��#'&ԥ_��8��l�"G�d7��ey�O2)����F�4Z�-��).��Gls��	���Iğ��	؟b>ݖ'��6̀�$$	�׹rP���Z��ZV��Or�]��u�?!�_���	`a@����	P���DA�������������'���p7#�or)O���t%ժ �x ��p�Z !3?OX��?a��?i��?����.N^d��/R�7J�L����)�RYn�>hb�Q�I۟���x��۟����{�)��;�r��3�߃M�U��M˜�?����S�'p��q�ڴ�y��E�@R���1�|}�����y24Lh��䓦���O��ąb¢��Pl�42bN���F@`�$�Oh���O,ʓZ\��J�1�'2Ŋ3&�Y�3J£)nt
U��^�Ort�'�2�'�'���a��6ո����ɢZxD3�O�q���Ǉ~)���F�<�)E�?�F��OĈQcO�s,()��ޛ0|�ë�O��d�O��D�O��}"��Db��<=�V��7�M�DQ#�Z���	���B�'E�66�i�*Q���v�8��F�	�p�P�l����L��+(8Tl�S~Zw� � �O�:���Ԁ�åkĈ2Ȱ �5%c��Iy��'n��'5�'���`ā 
�p�P�"��y4�;�MÔM���?���?1M~�-�6� �/�'a�[���h�Ա�Y�<��ʟ`'�b>i��e��)*t�p�,?���"�� Nn�=?9���A��D������d����0��&�ɲ��!|���$�Oz�d�O�4��ʓS��FƖA���Z;24�(�2�	j�����m�?8B�k�h��p�O����O2�d˔D�:C��[��6�C(%�`ٔ�s�L��x"��?%?y�����<��a³7�TP�#B�5m��ß<��͟4�	��8�I{�'d�T#���6>Z�u�D�B7
�xk��?��l��	���4�'��6�;�Ēw�ԑ�D]�}Q�YCA낢D�(�OH���O�iջXY�6m ?�$�պg��QD ��E�*H���,?nLmo�S?N>)(O����O����O������4�p�IwO��0��O��$�<�p�if����'}b�'W�Әc��H� ��}J e�%�5��R��	՟��	d�)��
�>�Ҽ[��
'`�`$a5!����1��Z��Ms�X��,?��$8��[�g�Y���ZR��{Gd��l��D�O��D�O���I�<���i?n��5&]v@p��a��h%�p���C�X`剝�M{����>yűi��5�RȞ;e��q1�\�7�Hcs�y��o��`�XoZO~���e���SG���{�~��a�62)*ḤŘ�2�d�<����?��?����?Y,���A�E�M�vݙ�`NV����Ԧi�E�������%?�Ɂ�M�;;Ѯ�憓ME���Ӎ]�;��ų���?�L>�|BE�ɨ�M�'�HP:���=a�x7'P\I�ă�'�.�٣&A͟���|�V��S�����i�t^�5@G� �<�a�h�����	П���LyR�x� �c��O`�D�O"4+u�̗-�����/L�1��8�&G"�������O��$-�$Q�	� �ZȐ�"��]�I N��-A��+b>I��'��I72���A�=�n���HC ������	�����r�O�b,D/e,B(��\K���4~��d��|y���OR�D̦��?�;fF��&�۶���,V�|>͓�?���?���	�M��O�n]�v< �)1������/I���ʁ�U��FI�J>�)O��?Y�`�Tj�(U$�+EF�P�
�q~�.mӘ�	���O����OR�?%���8�`��萱( P+�K����O���:�󉌖3Z�  ��p � �ׇE�Ъ1$oӠ$�'�>,cw�VL?L>�*O2E���ş/|X<��&ܿi���u@�OT�D�O����O�i�<14�i��3��'��Q��1r���*����X؉�'�27�4�	���զar�4F��6�L51�2d�f��S�R�YA�@�{S�}j��i��I!���Oq���N�,��4�#�
�L�bh�3!�}��D�O����O����O��D"�S�b�^����߄����$_q���'үw�2Q!�?}C�4�� �e�&��l��Q���7@��A�x��'��O��2�i+��p�2�Is�3�4t�ť�)("\��5`2LG�	_y�O�r�':b�×TL@a�`�(]���PIٜV���'N�I6�M�T��?Y���?�,�4�2'�1d�.u:��̠!$x�%��la,O���w�B'��''~�㖊�,I�H���BCT��pZ�G���QkVz~�O>���	�t]�'o4ɪ�-Q�n�!�Θ?VɅ�'���'�r���O����M�&�4S�i��]�l��1� ϔ�eK�8Y���?�`�i�O���'��6-W;rx���.R�Z�4���=q�o��MS����MK�O�*�Q��J?u�$IG:z�>��G���j˷���y�^�H�I�$��蟐�	Ɵ<�O"h&��,����r7����dӴ���@�O��D�ON����D���]z�x�2D*ٜ��!ǟO���Iܟ�%�b>�ZUA�馡�S�? j��`�#q�b$[�g�W	B�=OB<���2�?!�`9���<Q.OP�6�$l�<��ӫW�X���'Qx7�\�;�r��?�� I*v�T��QA��djQQm���'���?�����wn�gD�`��t�Á��+�XE�'�����H�^�r����������'�H�u���N���Y�"�I�Z<�
�'�P�C��@�R�J��B�m
g�'� 6m�H����O��l�Ӽ�s�W�e.�+w�YCFБ����<Y���?Q�TP��	ݴ��d��1t�h�O;�x�TF�� �4��[��ݻ&�|bY��ER�̩K�p�򎚾=�(T�u$ܤ��d���*qɗП�ͦ!��x��E*��z'���L��Q%�[4mŮ9�S������`'�b>�C�� q�(��n��,K�(�#]��o��@�>�Щ��'K�'��I�����E3J I�-�,9��h���T�Iߟ��i>)�'1�6mO`���L �hf�ƧGh�HH��3YB���ʦ��?a�S���	����	(:��i��f�
y8r�QPK�pA�+����'d@-0B��OBI~
�;�Ay����D=�e`�7/Z����?����?���?�����E��_4��9�h�F��p���0�?���?A&�i
���O��bsӂ�O(����T&~��2'
�B��"��O�4�:���s���Ӻ��CԮK�t�NY�A��b��0:�j��^��Ol��?����?Y�r����X��VI��G�ؐK��?�)O�anZK�q��Οl�	c�T$���k")}��I�����X}�'�b�|ʟ�P�Aڵ�d�ˎ;�`�p0�^
!N|r�'I;K��i>���'��u%����'�h�8��'�Zv "1"2�����I؟(���b>y�'�x6�Yk�M.&�jC"�7S;��1����Uͦ��?	CR��	�IǄ,��Y�t�c2Mׇ<�����:�LҦ��'��A8e��?e�����`�Y�:��80����1�(#:O���?y���?����?�����I߰T#�p�d���I�ɒ�l�o��R������h��|�s�h�����#�'~>�Ǐ,)>ĝuި�?y���Ş'X��8ش�y2J� ^r�$ �%�̔�˯�y�%׌QP ��ɫX��'U�)2HU*�vD�EJ$��BTTr�P!�4i���h���?Q��c;�0�A�d?�-�BD��:�
q[���>1��?�J>9���)��Y�`�1O�=�5�e~������iƞ��6�	�'�"�^[՚a4CZ".ռ�(�,V�R�'*R�'X"�S쟄b��F�E2�o���j࢐�R۟�1ٴ�b�C)OZIm�X�Ӽ���ˈ2x�d���Th��G��<)��?!��]��l�ߴ���D(=��9�'*#2`�W��@f�ҩ �VYA#�Į<ͧ�?���?Q���?`e�S�`I�%؟n�N\(�����ܦ� ������I��$?牬[B��T)��p���E*��1�O
���O�O1���0@�K�InDY��ν
d�t�������ē���T��?'2�GB�	Ny�`��y�cV3 �\�jV�XV��'}��'��O��I��M�	��?)���	н邬��X�0���
�<釱iV�Ob$�'�"�'A���\�D�""�-o|U��o�M[�O��V���b���w'>p�`7A6��&ݽe���'gB�':r�'sR�'R���B�#Ƭn���
��Ĺ>3�����Oj���O�,o�+|���͟4��4��XZR|�	H=5}`�`⧋#P_��M>a��?ͧjn"P�4�����|���˧Cm(-3u$��P(�IE��'����Ӳ�䓓���O�D�O��׏���0��ȩ%�!�֦�&Hc����O&ʓl��� �XXB�'�"Y>�)Q?G�R��]4��۲'*?9�U��	�'��'q�f�R�N )*�rrm�,W�ag,��4b�d�7��<��4���a��J�OJ��� �:��VH�4Y����O����O����O1�4ʓ4F��GR?N��`��L�2qp� @O%3T*��4X��J�4��'|p��?a�/��J��d0��;��c����?���\d��ܴ����:d�����#*O��
f��fJ^	��đ�J����5O˓�?a��?���?������b%����+@%<-��"�Y�[�m��H8x�	���IG�S������!��ex��h�dC�X(�����?Y����S�'Mp��ܴ�y���
���U�2V.�4C4j��y��ةY�29�����d�O.��V&*ո�A�mͧ3��m)�%��1�(�D�O����O��_@���U9c�B�'��g�<�laOW��'/�Up�O| �'�b�'�'�؜bԀB�Y��uQ !

a�D���Ol-��K&�46��x��L$�D�Od<�&d��4�h���=:"�$�C��O����O����O&�}����Y(���7��Ҏ�9	���$���� �z^2�'��7-)�iޕ3��ҋ@�bq��c['=�r%��$t�<�	��|�I�PA�Um�q~�I�\��%��b�I8�ݹJh��
�ԥJu�%bL>!,O�D�On�$�On��O���&C��3�`y�h�1	�=i�m�<ჶi��AR$�'Nb�'9�OLbM�
7�2�*���,��p ��K
g��?q����S�'ij��� �㠇��kp�p ��	ˤ�ѥ��Pp�'0MYVl�o?�N>1.O:�Qb��b��Xڱ`R?K�t`I+�O���O�d�O�ɭ<Y�i�B����'�qt	���x�ϖW���Q�'WB6-#��&���O��d�O�Q���q���H�(J� ��	B�w�6-??�,ا~U�)=���QcuBV6Q�v�;�kڮ
�X���`����h��ȟ����D�
�-[1k��U�`�:�pH�Fٵ�?����?���i9,�\�<�ش��^�%K�!ߑW2 �⧁D�@��M>���?�'$[ґp�4���W�k�laQ!�8$~�[�#�63x��2+T6�?1A�7�D�<ͧ�?��?�$��&1`�_7���@�3�?����$�ɦY�A�E�����؟X�OA8d� $ߘ,��MR!�2Y.��OB��'��'Dɧ��Y����֎H-�|l�ڏjJ�U8���.f��ղ����]���O�	02f�3�V�Tp��Sg�Ex�U�I؟�������)�Shy�i���� ��*�|��܂��; �`��`�O���]ئ�?W��	�#�2pI2.G*>�C�'�&�H��	՟���˦-�'U�\�a���?ͥ�4Maΰ�M��IA,I��-k�cx�ؕ'�2�'���'���'��Ӕ%�2)y�Ax� ����h}8�4^:�����?�����?I���y�/��T�Y3�ܾv��x[��_�zy�'�ɧ�OL�G�i��ʭ[��G׺ 7n�i�둵V���)^�+�'��'����|��^u��p��;Wct-�o��I��0�	ݟ��IП�'8\6
1�����O��Y�t:�W삣=A@�
���j��OV�d�L}��'���|��\Ŋ#�hհL0"��ҿ���ѪL!�A�s�F�z7�I���7|�d�i�N��V�ʕ�Д1�ER�����O����Ob��7�'�?���^�~�`i@d�Z�b��-��	��?���iȰh�c\��J۴���y�m쨋U��'��<ȑ�Լ�y2�'��'W��i��	�>;r�3u�OE�]�E�Qq�d ���,7�Ft����U�Imy�OQ2�'�r�'p�:-Pt8U�C,']�;���F��I�M�e����?���?!I~Γ��QSB�U�zcf�F�q�����g}R�'!r�5��	D��Ri�O�N� ��I�:�d�BAR��I�Z/�8��'-R%���'�P�`�
�3y,�Q'#F�w����'�"�'R���X�d�شFe�����|� *k_�12ƣ p/����B���$Il}b�gӀ�lڼ�Mcp�Q0d�PQF�pB�Y�o�j��a��4��I�T0�A����O
��A�
�����/%8~�R���y��'"�'R�'�B�I@�hK}Zf�@4�c$�X(T}���O�����uˀ��@y�fӐ�Ob`3��O�@��vA�_q E&Gv�ҟ��i>�#��M+�Od`�ͅ��1R��֛�ܫ2�5:Rx����R�n�Ot��|j���?)�s�2�P ��wRF)x���\|����?�-O��l��)�BX���	E������I��d��1�a�d����d�N}�'��	>�?�*�ȈV�Y��� e�����խ"Ќȉ!�]�5uZ��|3��O��H>�E&1�u���Z:�h���?����?����?�|j+O�!mZ�N4X�Q��ݵRDv�෡2X�*t*A�UZy¯}Ӝ���Oz��H�B�֡#*N�{`ʀ�,��$E�-3Ʀ��'*Bi����?��������zʸ{�N�w��<�R?O�˓�?A��?���?Y����	Ĩ3H�8©�;��1K$+��<nL:���ßP��H�SßP���oΉ0r����ն�2�� d��'�O1���AC`�4�	�;���P�fQ�(�nH2�/Ю�h�		4-��'��&�$���d�'�0Ⱥ�a� A�d5AP�^�>U�\�$�' R�'_"P��y޴4$����?��qx�Q�Ѫ��Q+%B �p�9��>Q־i�:7�H�I>%��I�9���fOr�H�q"��E�Q����|b��O��A�"���e �2k����B�K���q��?����?����h��NI!�,��bͪPR�����J�Ҍ���ɦ�4bJԟt��=�MsJ>��Ӽ�*�#j�|��_1��T`����<���?��[�.��ܴ��$̶pl��OAސ�4�	b�n�cgJȤy�f� ��|rZ�$��������i�Q
tñ^�h�B� ��C��QE�S`y��p�\0�O �D�O`�����.!Dr��Us��e	�`��'�2�'Jɧ�O�N��s`�06���T�ޒB�Ȱu��y�f$�QZ�p��Ɩ�P2�{��dy��J�榥y�.�:�0m&f\e��'���'|�O��I!�M#%��2�?9v\��`���+X#&�ʤI�?9��i��OV��'���'�r@��_C8�	�FIb�;�	���@$c�i3�I'NbLX�ԟ.���NT
ha8�qGɋ>z H:r��?��O����O���OJ��*��43��Uƌ¼�U$i��\��ݟ��I��M� ��|��U-�6�|P�BA�8�P"�A)R��8 �|"�'��O��9bs�i�I?Be`�Z�,�K��e�w�E���%L-5��:��<����?����?Y��]�)l|Y#a�J�E ƙ�?Q�����ʦ�iƆ�۟��	���OT��a�C�|A�5H�80.��Or��'�B�'#ɧ�� ty��X���������8 �3�A�g������w�R����ΝM?iN>�RF��}l<
�h��/�J���&�#�?���?���?�|*O,$mZLX��{�J(�rGdχ�R4Q�m��|�	��MÈ�ʽ>i�c��t�"�xtbc�!q��0��?"n���M��O�C�����P�d���LD��PP�H��H�,c�4�'!��'@�'.��'��8��t��쑻(���
���H4f��ش@�8Z���?����'�?���y�ˎ��1@&��<\x�Õk�Q���'�ɧ�O)�H���i���v�vX
Vh��T�HYD����D��@�,��'��'���t�	�^n����*��%�q���	۟��	���' �7-��3@��$�O��$ExH}��'�&>m��$�1%�X⟴��O�$�O6�O�E�B �W*x��%��!5<�������NP+6td�K&�ӯ6�K����ܷ*�p|�$�+YT����Dϟp�Iҟ,�	���E���'M���P�3#�طǈ=4��'j�6m"�0���O9mZZ�Ӽ[q�؃=�P��%�?�M3�Dw?���M��i:�*5�i]���&�	0�O��j� M^yD�aRf�!+�&��#NB�-|8Hq�@Z��ꐮ6�t{��q$����cW4?�v9ʢLG�1DH+�dze,)i�ē	�����K�,0�A�� &�ɰp
Z���(zS`�Y �%x��[����a�d7+��˳��1&�@�]� Ch1;-�6�l�¯���i��9�J�2��;2�B��a�Z�ɞm�Ҏ�R�+0��8�~T�Sk�� q`�����d0hiD�5�NP�
<��ik���,�.�8�hѕ]n1X�k�h�
Zb��6*A$�`�")Đ�hŮ��'baoȟ�I���S����X�ڴh��6�n�ae)�G��o۟��I�(���?�����)�ʁD�6�0�bE��?�ԧ��M���?����S�4�'/���Y����"J*<�t��G�x�$�bU��O�'�?	� C��e�P�b@��:�����v�'�B�'�6J��>�-Ol�Ľ�9���$g�r8q��Ǻf!N��'�	��^Q$���	쟰�ISv`K�")�� ʐK�&,Z��ܴ�?af� �	Zy��'cɧ5KD�"��I$���B�ʅ#��D�5,�O��OH��5?�Х� �r�B IN'=}�P��H�	�))�O0��?IK>����?��%N
{�Բ��H�Abl)�fԬ6��<���?y������=Y���.i�4��*�>m��r�b�2u%�6ͽ<������?���3&Np#�'B�b!G���!�;!Sv0�wf�M}��'�R�'��		.��O���_	zP
"�%���,c�}��i��|�'��&�.�qOF��.2h��:�N�&C��R�i��'��I�{����O�r�'����]-&оxa%�Z�\��2�,^P)�O���O��R3�:��JBV��1���"p	/#�"t�U�����'($���io��'q�O����p�<L�x��O�*E� A3�+�榙����XԮ�a���Ocr#c��^�����O��W�X���x�T��4�?Q��?������cyb�L�l������&��3�S�e��6-�^�����<�D�0�ç� 	AC�i��'�B+�!�N듂��O�I�L���He��7-(@�d�Ck0c� �$F�[�	Ɵp��ȟx���
,~ـ��I/�����A��M���
i���P� �'�r�|ZcfqF��<0�V���-��	�O�\"D%���O��$�O��-¸����!i�����J$ 1Af�˞����<i����?a���1s���+��I�b&98T���O��䓹?���?�*O�"A���|�p�/�iC!O��LT�t�q}��'*R�|�^��蟰b�n^���Źr��p,>�#��A���d�O��$�O�˓`�BP@!��4�F5J���&��E ��a�j�<7m�OؒOf��|r����8��і-ц5��e��敞PVd7-�O����<9��،�Oor��5V� "�p �1��c�ƕ�To������Ox�d,�9O��,��M[Pd��"%��R��΁6���U���d唭�MC2Z?)�	�?y��O�a���$l��MKB��O-��B�i2����� ��'��禩�$�ɚz�xೇB�t�6t� �iӀ�kB�Ϧ9�	�@�	�?��I<�'8MH����c�&i��ȯ3 �=z��i���',b�|ʟ��OJE3�N�	�$�K����|��P�g����a��䟼��'v�N�H<�'�?��'_����f�0S)�4*�f�to�Ecߴ�?N>��^?��i�����(�~HK᠂�}ux���4�?٤�����v���D�$Y����2鐣�v�#w�N<0�$'��)���Е'VR͇..|> ��`M�m�d*%ȉ�
����W���	�0�?����~�%K�!Dh��	3"����U;�M��kW}̓�?*O���A.����&���B��4p�Q�'Q�O�R7M�O��+�	؟d�'�$��4,�PтM7�Y[E�K�3��$�\�I[y��'��U�X>E��*B\u���?T��K���)��f�i��O����<1`��P�	�M��+��@�%-2�a�"I���6M�O�ʓ�?!�����Ot����k숭|�<��T-�Q�ޕ�!�ȃ(M�'��S��.(�Ӻ�td�IвL��kQ�+�$��N}��'#����'|��'Q��O��i�� Py�����h��Տ&�H3�i��P��"ׯ9�S�S2Z�r5r�iC�2�0�a��aZ�7-�{Ϯ�D�O���OB�ɺ<�O�r��ÆFn8���E_YP| p��>�4�r���Oeb�C��RX��c�f��aۆb9K�>7��Ot���O��v�g�i>a�IY?��/��'R͉�.��7\Ȑ�G�ᦱ�	j�	���9O@���O��5`��03�%+R����Ӡ4ڸ�l�ҟ�0�FE����|����Ӻ�1�D2@�@����q���� k��꟠�''�'��R�X��و@��J�MG�
,���L,ט-L<Y��?A.O`��<�;	"��ҭ�?�(t+�e�*}LmZϟ��'���'u�Z�L�%�����z��Y3S��/�H���,о����O���,���<ͧ�?)R�5
����@Z',�Ԁ7���S��'
"Z�T��,w�8�O�2�Ԥ2Z^����.�Q��ϪA,7m#�I˟h�'��%�L<���݃�Ā�6%�,Œ�!&H�ܦ=�I̟��'3��@w�!�	�O�����0QΊ)�h黴�06f,(0��xbY���i�M�K~�Ӻ�P�4~$�HB���<�Tm���XԦ��'��|IGk�$E�O�R�O���_�$�y�F�*@�|mZ3 �EY��l�Dy��'r�&�7��i�jr���G�%�t�W�-]ĥ��4����Ÿi��'�"�O^O�I��<�^-�D!~��z�$�*�L�l��^�B��	П �'���y��'�� ��\��I`u��:c� �qmc�����Ol�d�4^`�'��Ɵ���[c�a*���P�F`y��V�%�~l����	�L�5�s��'�?9��?ᇹ^4t�T�ûW_��p֮�$p��o�Ɵ�3f�K���d�<q���D�Okl fȈ�5�T�4���Iݿě��'>�4�'���ǟ��	ǟ̖'���9���mQʽ��ϋbR(�{�3f����D�O�ʓ�?����?�tC�_��lF�>�䈈�({���ϓ�?����?���?�+O��Ń�|��\2M2���P �"�|\��L�����'A�R���	�� ��
@|�	�'S�E��ǐs��@犇�(�l6-�O��D�O6��<�g
�9x�����@)�e�"�H(��3X��lQ"��7�MS����D�O��d�O�]#�=O��禩(�%J�q<h� O�?�Tlh$Nb���$�O�˓%;搻%U?��	���sIp��ǃf'\�9�/�" �!XƠ�K}��'"�'����'��	֟���W�t�E���O&��tϕ5�°lZXy��	3{�7��O����O���u}Zw	l�y��
����'g��Ua��4�?���^6�̓���Oz�>�c�"��U]��p���<fЎ����v� a���Q��)�	��|�	�?��O�˓�"-�e��X��X$�����`qкi.|x�'��'��n����*�H
�"�7jR<�U%�*T���l�̟d�IdO#��$�<����~2��8��y�E/n4�4r�T��M������P^��?��쟬��b謙�K�6`p�!���!�"0B�4�?Y�.��@��	ay��'��I���?��yyb- <XI����xbX7Mg��
0O��d�O�D�O�d�<1��ɔ"�TMP"���� �j���(H�]��'A�Z���	ӟ ��

V�)te�#��$`T�Ղq���i���	��I���_ybA٣B��(i��`��q�"|)#ɗ�c֊6-�<1�����O���O�y�S8O� ����6q9���F�/p���oRѦ���������H�'Z�(Ђ;~���/���&�����C^�}m���'"�'��L��y��'���Iw��z��
�k/L��"�@���'Ub]�\JC������O�����=���Q�1q��Ǯ	���bĤTE}��'=�'!��'��S����,��,!�/��[���9��yn�Zyb�`7��O���O\�ic}Zw=`Z��m���s%�(:yaܴ�?I�7"4q�����O �R��/ ʐ�I��9=��ش���ĵi�"�'���Oj����đ2ɮ�Z��W>8��f��>o*)l:b�����*�러A���2i��c��P��+��M����?y�x}��v_���'���O�X�C&ٞ~��b0��O
F��t�iw�_�xI��a��?	���?�CF�!	� �i�!�+#y|���oɛ6�'}d�s�K�>�.O8���<�����L	$u[pBB+�&�L����q}2̏��yBZ��������Iiy�-׵v:�c��@ �*a��ǒ�4� 9b7ϳ>�-O��<����?A�,0�,#�!�A����5(��)����de�<)��?Q���?Y���d*A-�T�'D�z���1N��ad��g�nZMy"�'o�	͟���̟�"!g���>Ĝx�U2˸����	�O�r��?����?�/O���c�W�4�'��ɍ	O��I2��Q��(��a�����<����?��V�6̓�?��'R�P�#Ƀ\a\Q�F$= b�4�?�����o���O]��'��D(�P����B�ԘQ��F���?����?�!��<�N>�OXZ�� ��9@�(�"5pM��4��;��l�؟���ß��������BTJ�[T,�7�!A�YѾi�b�'�x�k�'+��'&r���`����j�X�hi1�؛6��r[Z7m�OF�d�O��i�k�`�Ɋ�.Q�%�����\�����i�uК'�'��4�dQ:i%\�r���Y�*����a&� oߟ���ݟ� 섢���?!���~
� �)7퉯G�6AC�'Ai����$ϻ1��OZ���O���ܴ:P�a3��u��Qq)|X&1m�� s������?	�����S2�S8�j!B�!L(8�#�C}BD��y�P�d�I�����ByBbO
R֩BA�	�#8��ҧ�e��(�=��O���=�$�O��D�.�H�#�0�������6��{P=O���?���?�.Oʠc���|�#�� �n�h�I�AB��Y%��u}"�'k�|2�'j��+F��K�	-���@�ۂ1��I�^��V��?����?�,Ol�R #[U�� �t|��l�Y�I1�NYe��dJ�4�?�J>����?y�ʑ���'O�8����
���(K0RH!ٴ�?�����'o��&>e���?y��K������<$7by��-dA�OD�D�O>�D�s)�$$�d�?�e��)r��	�Q|0��C�tӮ��䌢��i�H�'�?��'����/`]�`��O��E���ς�\7��O����2�D2�S_U��y H��I�Y���(('\7&<�$l�џ���ɟ��.��'Q���jN�b�%JRc">@�!��xӐ@�w��O`�OZ�?Y���9�^`jqK}{�؄8$"��4�?!��?�V��'���'�)fZ�rd�R�.DEh�,����|��P�_[f�D�d�O�����p	K�J��K��2�eL�b�.Hm����ރ�ē�?������	߆&rF�����A�^��B�O}R��F��Z������h��jy�_G5�����:�z��@�H4J'*dx�,;��џp'����џ�J�!�@Vx��h�]��82�X�r�����wy��'�ґ��a�
cY�瓱v�,x�c�4yW��sh g��듟?�����?��0�����8o�Y���Q��U���02�͸PY���Iʟ���Ey2�Q$j�d���i5�5Fw�\b��+.<
�����%��Q�Iǟ �ɸW&H��a�d�jtҸI�a��t���!�bo���'��^�Ha -C���'�?��bt�R4ɂ_"�ԁǨ��ݨ@r�x�'˔���O���?DE�`�P���;��a�l؆��6��<a�%F3���˪~:���6��P�̙�-(��� �yؤ��Bi�>a����;����S�'}���萾@SЀ��
�f��mZ4�ߴ�?���?���U�������/R	�2�G���@�u&��?���d�'���E�4E�.�i��"A�q|Ӓ���O��$�6��)�	�O��	�.>�-�R�	�n�~�� �A`�\�yBHхJ�h�����O���m p�!��G�ptb�j] ol
@l�@L0�ē�?������ò�/�đ��I�"�����(W}}�HJ���'�B�'="U�ؘ �E2xX��(v	T�s#��l�Xd:K<���?QL>��?i䠑4a�Tl(ĭ Ժ(�Vf�#,�*�(��ӟ��'=�蒌���P(y;¸ђ
�&���k�
<B�'X"�']�'Y�	x�4퉰�k�`���		]����E�[�s��@]������h��ğH���s���	Ɵ\�	Li\��`A�i�܅�Cz�~pp޴�?�L>�����S�'l2�%�L�>f�f��w�m�ܴ�?q���ˀX�&>a�	�?Q��C��u�S'�4V��y�vGҕ�MÊ�9�����i�\I0*�(X��s%O�Z��y�ش�?���M�ȱ��?�*O����O:��ƴ0RFU	Z->-��C��F�E)�iCR�'��K!�ט��O���BgȞE�e#VB��7f>h��4-7t���i���'�"�O/Rb���R�ܙH�����U8a6�	ҁĦ�M�p�C�'d��DD�*�RB�ǡpF������h/$�m����	ȟ��Ʌ����?)��~��>�Z��ׂ5R:��lM���'�n�ӋyR�'�2�'�xȩӡ�~f}�J�܀����u�0��Źrf����ӟ�&�ph0��)T}�(Z��@i����%����ć"l�����d�I˟���ly�!G�|T��K��Z��3��
��0`q�'��O����O>�8S�,,;�+��l!c�Ʀ2[,b�$�	������	>,7`d�'2Hy�T��/\j�T�S>l��l�`yB�'��']R�'��YCwۦ�M�[	̤�b�H�#�i8��)Y$�	��x�q%�'EЂei0�)�'my�2�M�YиI��iȑ��T�ȓ7O���%ݍ�fԛ�J�3-�rY��j��dc�R��E!E�/p�b�/�C*ޡ�u	ZD��1Y3���.��X9��V�Y.���BB3�ܙIbi��e���8���U���`N���~���Y�mFFQ[DO
�l���l��KH,غӡ�0Xl
�c�`͠��� .��d�՗������w�j����8(DXw/�O����Odȹ&�@={�i�z-
E��H�\��hB�e�0����Dd��J��t��O�1�GJ��:�`��̟C2l%��-�?Q�4��鋴�0�qv�Z9/����֬�:��dے��wc&��񮋓}@L��Æ	䈸"1����"�'�)��'�dCO��Ux�ܥ`�|bD`��> !��N*%��+�Z�,o04�O�6u��� ���?�8@�7(���KDء^����ϐƟ��	}���N�̟��	� �I��u'�'>���=FHV9�B��'"&	r
��D�d_�C�d{Ӥ�8�b ���hOT`	�D��oԎ\���ʖ���1E��ϟ���MZt�;y�$(k��hO� ���!��04P�B�%�.��@	E�O�e���'R�Uy���8tB���K=�8d(#���y(A�7|�PbJQ���mHu%E"~�#=�O��ɇ.�VB�4@PȣB��#:�Iȴ��0vP,
��?q���y���"�?����H�+D�b�"-R�q��Ύ�KiN�s�gD1t��)��(/�0̆�	&��J���D��xXE�ãm��0{���-᜕� 	��cd����'���S���?�q��.f���m�6�z�{rJ�_�<�wD%L}^@��n�P�*�Ӓe	u�<"˞�4�H�b�?,3���D�<����d9(��'"^>]J�ݗt���G6�0t8gLՃ@�9��ʟ��I�[�����G�L)ɄQ�ʧ6����!�`&Ts�A�r�$`Fy��;�:�Ѳ'IPH��>-�7 ]}?��TDn%h��&1ʓ-m���ɟ��� (%ZS"(�t�ܭIa&���Ņ�<���5AP=[u �xQ�i��nW7h�bą񉙉�B]��ѮP%������\<0ÐAϓ�ܐ�Q����p��Ɋ!RF��'��/\�1Y�`�5!��	T��b)���ad��S�(t�^�T>-�|�	-:tJ�P�;e�z�q�K�9xZ�"�!��Hb��΁'��$��S��?�ӡS�8��|�P�pk(���ß0��r~J~�O>��b�+x�%�kֆ<���00�W�<�K��C��E�v�ѭ#�n��m�'�L#=�O�T<��ج	����0D�2#4�Bb�'�T�Gx�!�'��'|�dwݥ�	�H��D-9����S���I�#����0Հ+�O��q�d�/je�(��ȑ�]vDdY��O��J��'k�k�M�(q��I#�院3����'L������=�Ud�(���)ԁ�3��@�<�t�Z��"��QJ�`�D�Բ3��"|��6Nv���~�����"�� 'ܼS���<4��'ir�'�|-@��'��0�x8j�'��F>>0t��#����Ă��_��p>A�{y���T�@|��Ч��`��/��p>����ߟ0���|H�)*¡W��إP7��<: �'���Iğ��?�O놴+Q�6�r��h! ��'`���;]���s�,�tP��'�D��򄓮��lZ��H�Iu���#\\�AI��}�b�'fR�O�4ၑ�'�2�'r�ɚW�'1O��"`Di� ��|�բc۰*�>�<��nz�O�Ո#/'uz$]���R������d�;B�S�M��X�� �Yr�͗!;B䉃f�z<����-v䲜���S?m����j�IU������$�\�'���W���	��iH�4�?)�����;+��'��5�4�7ł?��!ʡl�3'���"��'R1O�3� ����rl�bMz�#iʥ�F��O?�D���(ٗ�A�E�\3�n�(?�t`�w��Ob�"~�I,f�� ��7�ܓ�ʍ)H��C��h��H"$o[}���MW�g�#<��)��KT/P3���d���Oٸ�Hɚ�?I��-��=��mՁ�?���?Y�'X���O����u�M�`��d�.��sA�.M���-�}B�^�7p)tM
�x�b� ��׹�~�E���>�Wn]d�����0O�v�h���L?q���՟$��I	c�6m�al�[BN��կ@B�<B�	�'�b���a�pg<�S�.T�����ᓾ`��Pp޴-�
��.?��tR嫘�4J�����?���y�H���?i�����O���?��l��䋇@<(R��ʏ8�N���ɳS*�d�~�	��ؠl���	��דn�a��3\O��D�O^�"�@rf�3&�4L�!@g"O�T�Ķ�|p�*[ X!���y�<K����[8hģ@���yB�.�ɕ{,��ߴ�?����IDu��à�V9	V�I��4{�Dx렡�Oz�d�On]�d��O�b��'����rgt���)��hGyZP�r��		�"1��`
T�
=��_�b�Q�f��O2�}�&�+WBN�WF۶j�|r +�h�<� P�*ؐ|0s��6{Ĭ�ŁKg�$�I<1��ѴV��dF�``���<��YK���'4�?�����O���Oެy��*
�����" `s`��4�@��>�|FxRDܙ�������b��2NPEJ!(R�)���ƃ� ,�!��ĩwؐ�E���bk<��	g�S��?� (0�(�+^���Be�%"X���"O�ع�$�9��%�_:CK�Bቢ�HO���8 �kf�X�d\�(��E�	��s���~�i��؟@�I��P�^w�w��h�ɒ=c�&m#�ӫDN�x�'���g/� U�ڙ��G,Oj,��f��n����FO�/��}��O̡�� ��i�p���v8��s%SJʼ,�D�?Q�h�8�ʟ@���K۟�ݴ3�����D�O��|jx}���3�DD�F�C,8�r4��[˒�BOM�`	� ��&�p4KB鉨ej���<yf@=Z��n�aJ���g��I��s�F�����O����O��أ��O���`>ũ@��O��D p7��ʃ�L�Xc*�sȢ4���:D[!��&�QB�x��"�nA<YSs ��:%��C��A�;D�z��N	�?)��/E|`�f�Qb�� ӣk�J�8x����?a.O ��6�)����;e�D�r�G܄b�B1�U�{��G{�LZ'��@i�� �h�8S♅�y� �>qI>� �����2$ޜbb^@��I�dy�B��T
��r�☶NdD�&�JxԼB�ɧzn���F�؆;zF�!�c�5N
�B�	�&%Р�C�si.}S�L���c��l)���mQ���MΑa8��g2 ��ZmF��/A�̅��+�ZT�&�˺_ Lp�휼Ts����J=����I�NT��)�U!$B�	�3o��i"F	�ZE��ͣ
B��4�^!cK��_9V��Fɉ�B74B��&J��+'b�d����d��-"��C䉛b'����'J�`Y2r
� d@0C�I)NRɨS���B���=M�C䉉d�D�1Ɓ͔<g�Y(aF�:b�C�5.O�l�3C�p���	G��bC�-�B�@�&�V�zФ�/C�I%@�RA@@L��� ȉ�Á74C�ɒ+��8J1N�ܡ���ʮ0�.C��/J^l�3��Tм)+���*o��C�	�ZJL��((��53���C�2H����½,�9Je�>K�C�I�T|�(��G%cؠl��J�7
|C䉟Wr��ĬG$u�n��o9;>C䉝'@r�A�bZ�9%D�@l�-�B�	>���t�M�+~`(`��4$�B䉙!�u�V!ێ.	��(`& �/�`C�IY����O�}�ȉr���	c�$C��5`S�=��	�^��a�I�GRC�əOк-	�`
e�FhP'�"O�(C�#qVT��g�2�)�pbL�(X����'��p ���_��h0oQQ8=a	�'�L� �h�Yo�ݡ'&��D��|"
�'ʬ��$HX����a
ψ:c1	�'t<@��0&�����ޯaG����'d�P�I��plƔ#V�\�p�pPLG	a���K��& ��f��P�: �� �*L�|܆牵T�* � �h~"��,?��,b�'��:��yI��y�-�{ӞԒ�G�b��
qAȧ��f��%J�Aɥ�0|��C�x���"���v�ޅ1B��<�5�F
I�Jh[oD�9#J0��Z�x�$�Q�@�g��ѪK�N� m�'���sʙ�@����qe�YJ��%�����eQ!�R�Y�Ɲ� Yj��$���f��B�AWX����0Q��yB�E_H��0����ϛ�$�8�έo�*L>D��Pi��]ib��残�:����Ц=����>����P�<�N�ІdZ�U���P�A�EO!��"OBy�́OZ��Ya�M(F]v};s*�J��'Uf]{���>�fi_�{�l4�� πa���2��Ch<	H�'��	q"�[<|c�}h��D1��X0-��0?��,�*�=Ga��r6�px�0A�*�?Ci��槀 ��	T��u�ؽ�U��
x�C"O�P�� l2ى�˙�p�pa�Ę�`�0��O���xB��/�֠�आ^hzա�'-�8BƊ�t� ��(�.\b.��	�'}��Ə�0o��2���;	��a	�'�Z�q�#)m���1��͌0�-��'�DK�ht���W�JV���'��xSņ�Z*�q���U�1rĭ��'r�1`q��."�Ek�̗ +Q����'n�s�N�!K<. y�n�)q�y9�'��\����VH���DԒ�j���'�VtXE%�3�L�Ģ��^��SL>�D���V�y҉��� S��@�B�������?�V���r�y�p(�I��uq3�k�0�ä'>$��J�
�%o�<��!*����>�,膜�r,!�)�"]8�m��;�4<Y�H�\B�I�8�D\�r� a\�R �W�� �Z�1!J �)�S�/"h 1�f�^��mP��_%kN@R1"OFt���hr7d	�Fl�0�d�N|��'�@5�"�<��5���b@��	�����uEC�(E>��ybQ� GRL	���s~��^���ؖ��{�S�O�t�+-P谼��ڻy����'#f�R�E�J���Q���w��@��y���:s	�a�
Óy���KU�0�r��(E�zφ����9� ��s�BA�0������{c��r���>a$��%�OR��ak|<�@�(.QX����'cR���g
��'����n� �J��  #��nR�D��,��jy�8!�+�}붠�`�1���ΫS2*�p����.�Z}B�#*��SW*+-O꼘5��$H*�١C�9X�>�q��|�<��a�&j�������S5�#V�V�X��ll�;:�ߴO�u�W"��<��<1Q��"�n�ϻ��2�kU�:�� ������I 	�`�ڤLL��L�w�L!i�!�dM	�x�L��!ö^�N��j¦)ϓiפE�P�ȹR�lA���R̓U���Aՠ=��Ac���>>F|Gx��ר/+�0P�#���6��� U�?��x3�x�@j��OdD��G�L�<A�1ϓhd&��BJܱx�DY�鉚&�E���<�g�Վe>��kV�I�`���U��#8�\�Z�k*?yկZ�g0,�ٷ��U������d\�k�j�<���B�,��yB�]-2� e���ƌt9�%�	XD�� �O�ʣ)�o�J�!���?YGkV�\Z��� ����Z�\st�١E�1�P�)��]R��"��]�nn�Q�@%�p:PiqqJI�<y.iK��Q�D�] ��7�����Y��KR-�50�PhsuBY����y����4��A��H��2��-^��O��IUi)3�T؇ѱ$��d��[��HE	�<0>T�vSd�xmA�B�.
T@0��[����C���6�0=I��V�*�XP��J&��*�cћtm��h���Eu.1�`ꍍ2���'U�-�q�Is/���O���U�� +��h���#F޹1�"O`q�ć��<@0EK�I [����
���`n6H��\}C�$p�M
�n@��u�2�HsHȳ	�B%@V��;9a|"�:ܐ�Uh�ML���Z�G�(��cJ�������`�t~�τ��,9��٢	پY�� %��'��`�t�C�'9 �h^�7��q!�� nd����@��{�����=?����U�:I wC�>4�Di7`P>*��a[���$2�D!�G�'�\��$���}t��Ǜ�*Ӯ���Ո���sHG!X��h�6�<��Ok��
R��4���E<	�5a܏�!��2�4���rgbP񇪚%:��+g��8U5��9��U,�;�w	 ��I�fpE�f�ŞC�8�s��]�/ԹD��A��=�����d�Rq�%�J�$�kH���[U�(�вO�]��O�q#,O�|�0��eO7yr.�����%7�8<B�NH�y�`�'h۾.r��xb.�As	�B�r�i@�Ţ/��X�#�:t���* "����=Q�h�+c�`�k��T��pb�$uF�6��0��H��*g�@D|�w��j�%ЮMc|t)��ڗ��ܪ�'��p�FG�D��0�&=\��5�����O��
��@<f��堃C�f`��L����6'ͫC}�pjdڣw�a|��C+P�1Q�I=3�-J�ʑV�I����>�p�OtѲVG�@t�����Y~�[��ɚX�D�4K��t;��H���">��"<Q���u1��a��iv����Eɟ�S>�čj'�� <^��!�ϣO����SÄ6�n�
�'a�A �ߵM�F`8uBB�"NLy��0D�\� b��$�+�����3?�缻��C!��!T ��p}�@m�O�<�  i{��y��2`cV�`�Zq����^r��C�f�ɬ���ŗ\}-�\�i��x��ǐo��Ѕ %�4��L��m9Ԭo��z�C��y*�+ �Sn�*Rg�G�����
ߙBR���$1f6+ `�i�t�޲$6�$p���ֹD.�ab�� �N�67�,I޴��1#�#� i��)	��/yPP�s�Q�X��C�ɽb���@i�1'���A�UM��)��JFq���.X�XTҰ�~�5aԁ�*���C5�ڥ?��H�������ٔ��U���ف����dL0}��T��(J;+�dy��g��ѓ�iy
d+���@���m>髒�A�6־�$� GΊ R�i�,y��A��-�I�5�`��xCN�|��j� O>y���6�)������?��d0�g��)���u�>+%���'��۔�<l���R1��<�t �I�xO
�{�"4��O�]��P&���)�:I�v(�C�,<�a���

bbC㉉k�$陵j�
h��r�ɁR�����B��#&��OP�*���i�đ��4M|H$J�g'v��%0�K�/C�l�
�������J��/1i�dA�����I7=��h�T-�,ߦ��Or�r�[v�	�X�8��)�}���c�
����+\�|( ��j��4B�+�"�S���Toj��s?$����Tk(��k��G 9!a!YGN�hV�|� "��*��Ȱi�0���P!�o�<!���=9�8�r딲C��̒T�.	��ї�n7Nҧ�����Wvb���7>#l���k��:�!�ʸq�x���'p�q��_���0Q�((;�/7�p=I���&��z�>j��!��My�P��@0�ڤ�t�i�Xdrd�z`]�и' ��ȓ#BN�X�J��K���iW.+k�"ExbeA�eϔ�����d�O��<�w�/�R�����O���h	�'�8��$�
�T)t�;J��A�ЇC�U�ҍ��]u��s���n�YĦћG�8$ԩ	�g D��s��q͚��G�.^�%9��h�8Ӥ��:��@��'�������t����d�];,8	�g�����hѩ
pdӂR�){f#2���~�VxBk�j�<��قƘ#Ȑ�C�BŃS��i��8���91�ߓE�<�3��i�U8���L��fOa13�=o8!�O?�:�h�"P56�˧+ Q�zA�����
�, Qk���0��Y��A��;K3��H�S�����>�\�<%D�F�G���5W�6�
�c�/waāy@	�)M1�QqcӉ`���������:�L�Xb�[�*��	�7er#<�S�N1�,x��/h���,�
���F��cA�DL21O��ƽF֖��L�	>�����MQ�'.������`�i`eـ-O���������L˗�� �$$��.�*��������0���|*D�ô�����x��)�:�ãJ���S��yb��#7X$��V�rD��BC�>��O�� ��0����#��X �F-y�B�	�&� �a�:K��DAK/-R˓[F�Ex��I�6g��))�H	�LS��w"�L�!�d��*�A:���N�����A�=�1O���V�'�$p,Y�l3x �ʙoM��@�'֎ةB��(�����μ^}���'�h�sT�z���g&ڼcj"I�' Xy
�̀�0��aW@O�V��Ar	�'¢�!� Q�P��HÆ��V�L�r�'���u3�MF�>-�|k�'�<9�����<'�H��oε2���Z�'�^���FB�P��3�&(�,�y	�'��q!G��7/&��Y�k8&���;	�'�>ٺ�V�w� ٺ�m�M(�a�'���s4�P=C@���IX��dZ�'Nȝ3p���;K�܀$�y_�1�'ct�;�nJ�ʬ�'*�!
dTc�'�ٹ׃]�`*�҇ɔ=����'�qbq&ӥ{���E#�w���#�'x�)ȐJ��t�x-�5�+q�� 9�'l��
�)�;�dIslʌr_��
�'����i˼,|RȻR/�*]�F�:
��� �1C#�� u�>)�����K�*�	�"O��t��.W�T�xq����I�U"O�9`�g�,:p�&�V�wʔ�"O��R	�>պE[Q�H�5�H�"O��)1jиI�Fp:Q�3hԜ�"O���R̈\�V�ӣe\	8B����"O��(ĭT�O6 �b��O�S=B!6"O���!&H�͐e�[ �1H�"O��bkG�[�����ҌA�<H�"Oj�8�����r��L`(ذ�W"OF��N�L�JÌ��Y%��3�"O�|Q�G=0��H�I�/m�Q"OztK![�TL,JTJF.<Ƭd�r"OP��V�'U�B]s�Iͩ
���A�"O���th��J�1q�Һo��<��"OX��۟~>\ض�;yp�eX�"Oh���<2�q���Y�%��T{d"O�u�E�ƽ19���0�W�z;����"O� 晋�P)P#�@3LI�q@�"O�5�@ᖴjo^�����v8P4�""O��6�ZDR��Z�%?�AI�"O��B�Ք-�����T  �qD"O8�X�C#��� �/I@��"O��b�������r`�լ
�R�"O" ��D;��8�CB�u� + "O,-C��vl�"�%L I0rI;d"O����f"@�Qp���#�PB"O,@1�k��&�k�䐍(�8�"O�c@ᆎ\oC��i��"O���L�����	=6晚�"O��ږ��:�ũF"Wb�!7"O|�ps��|Ff���
\�a�A"O�!%�{]�$��wg��"O��s�-B.�"���~��C�"O�����1,>%�B��s���s"O&A	���� �9SW�Ũ:��@I�"O�):@��9�|"��6�&��'"O�(��H�#*X�J2C���a��"Ot�;v��?Y��a�5d��B�f a�"O�з��ټ̳S"ĕ?��hr�"O��"�J�%?��;bƇz�4	�"O�`I"JH!P���q�4����"O��Z��\/l�� 8u�-J�����"O����D�Oa��ѭM:*Q�0"O�Qi@L�d��/Ձ��@ "O��B�ȣ~��Հ"/ҭt�|=P"O���c�ޠTZP3�͝V���9�"O�m�&�W�'� �Fm�5-�XܚR"O%�f�])c��p�l�9���"O4y���{}��T���u���"O� �N)K�X�&�(^����"O������?B� �R&[�u̕q�"Olp�s��h<:�8��ђQ�8	��"O��wEB<�Fm�$@ ��\��"OJ�I��ц="�msw��}�`\`r"O���%��%*=^ѢDI�;A<��"O��ǌ *wkh��T,���c"O��	r��!

���2ߊa���"O(d��!$(@�%e��7cL�)�"O�<B0AP"+�|��<4E��C0"OL���x�D�ч&�+#ڪU@f"O(�X�
�g���@4�^�RAx�"O:@�ũUWw�M;.� �v�2"O����d	
,!sM�s�|%��"O� �q�gK�S�:�He�V%�@�w"O
d��3�6hPĢރk�Z��g"OF�@7�3!f�ْ�A�6��A)"O��Wf��
��m�V���3wP���"O��P����1r2hB�s�b"O�ā�t}`��F�6b�h"O,���/��XY�2	�w�x�"O� 0cK�5}�h��Z��%I"O�QPD$�o3��FBS�KzlhW"Oޅ�P!	�M�|ƪ ���2"O���S G��Q�+W��)�d"OR�B�?,��I�J._ ��s"OA�ƫRG/V�zŌ�2�t���IK�$ �O9&� ��z�����#D�"��7?����ٓ
��@���!D�0��'�0�am�U�>��WM>D����M"Wq<���U�WQ(P`�k)D��{�ˇ�h�0�;�'YDj����%D�P�%B��?y|�b�ܨQtj�rƉ%D������y�ޜ3C)�;a��{��?D�������< ^$5�&rp�Aa�0D��c�EM��|�Q�I�)yj�-D��0��� � �W�F�%zbʔ�+O�<�ѫ0�ɍ&�[�ԧ����!¬B��� �`tg̳/���e�����'+�#=�P��3~�v�ҕ*� ������p�<�$�̂<�h���S3\Qq��_X�%�F��d�+xp K�kљ 	�*4�.I!򤖗+��Њ���jcHM��UU3!�$�9!�jiB7Ϙ;'y�%�G?q!��:\��$G�0s.�ش ��!�dO�=\HR��X�l��1bF悷*�!�
C}��k���-|�|(��8T!��/!���wG�D:!����h!�dxpIL�#(J-�ǂ99�!��<;ltyQ�D��,���E�e}!�d;^���. �9���x���Ky!��	�Fq�M�OS�N��ث!���!��� �1Q��8j�)z�JU1O����ʍ]�K"�@�Dj�8���%!��Cj���dO;T_(0Tk_ "�!��� M�����)�'q�@������!��;�����E>~�!%O�!�ρP"��#c��<6Bda���y!�$N	�LHw�_16uR6�\"m!�dM5�
�(ʠ\���pI�m!�$�H	�L�N��Y��X�"�Bp!��^fp�0様{�V�ɠ�q�!���
-7����]r�Xpȍ.u!�d�!ATA�!ɞ�f\��f)��+!�d�FDz@�'C�~h�h���4&�!�$?w?:�Qn�!j�tDi6U>f!�df�H�(�e� U�
�yT�gў�ᓄP��[p�?t���ª�5��C�	�@�2�v� �N��q���ˮB��'v�b8!e���X�#(�'J�C�	 A�4��cB����Ζ?v��IZ؟�� ��-g}�y���ݶL�R壡�;D��[��\�~��Tn��"���*O���ř$i�̰��)`�*�(�
O�7MM�#�$���I�MXEY�h݃th!�8�l�R)I�+��yC�!�D�r���W��`�h3�^m�!�3l�J�	����� �f�.�!�� |��c/OZ�Rh�c��	{,�z"OAx�c�4i��e�_y�Ԉ%"O^��ԥ��YT�M֡0jJ$�p"O���!b���1���,WX3�"O��@�*�S���Еi�+(��4C�"O,��G�&#����C�!|��C"O8�aE�S�7q�4�3��&VN!�"O
�)�2g7��+SL�u�x���"O���R@�e�l-+�לMȔ)�"O����R�d� X ��#�� ��"OJ�׉��YSzj����=��"O��Ql�#)�Шӏ��J���"O��d(�;���@
� �`�Z&"O���ǈ\�V���"oWO/z ���R8�(��Vy�X=y���H�8�JFE5D���2)4a��8�޶y*�)E�3D����N4��H�ǖ?�^=R�1D�|��$�z1k�@���)Z�##D�� P�W��ڱAT�H)n�5`�E?D���4耐'���JT��%+�N�3b=D��(�BZ��\aRɸ2
�P�!�D��'"�(1�#�����C�d�!�Ă�&Qd���T�)����ue�2
�!�$_0�J��ы9���J�v�!�DBx+*P��,~�yh%o��/�!�d�,a����]D��)�O�l�!��4xN�!S�2+�έ@��6�!��Ūo>�,���A�ui�u��Ǟy�!�F�OJ]C"'�m/�H��.J6�!�$�0$HbD81��A"8a�5N�"�!��_	{����!U	`1���U��h�!�E����Z�p���K�{!�� $J���K��� 4���4�!�$ӨxB�J��Cw�M�!��|�!� �d�(�a/ׅ!�>�[��	��!�߲ p����&�&+դL)���R�!�(��0��N)=��y�bO��!�d	Wx"ڶ.�wdF�z���!�U,����h�#G�@���h�!��$Os�e9��V�5)��Q"fӊ!�+���ӌɹ!�NT�GF�J!�$F(�@EQSN�8��3�ř5e�!��Y��s �/A�D`÷�юh�!�ғL�$@����4��e`R˄a!�d)Wؒ��"W�����!�d±]t��u�K�*�ҸĂ�!�!�Nmb$���%�4��A�_8'!��?"�$���B&z1��6L�!��M0�l����op��Q�,�!��+5�Ԝ:P��	E~.���"LD!�$E�.A�q�5EMR���@#!�J)P���%� �b�r�H!�@1(йz�GTW�b�1�%!�D� ~W��@/"B�T��!��!�DԊ�"W
534��'�2�!�$B3��a��O�Lِ�:�D�)p !�dIc͆�#���
��<ԃמP�!�d�C�0�Wr������[��'�&�j�C��8���*8�<	�'�z�$� ��,��fX�*�(�{�'�z|�*�6E߈� ���"-��8��'���+�m^����9G����6�'��%1B�T�#E�TʖA����R�'Jt��r'Y3��@���������� �`�����g�8gkILH�C"O��@	��z�09�	�K� ��"O��YEKO��y��gŅ�.���"O��%�&4���ၼ[w�k
�'Ț�i���"���'�J
.9����'Ofq�U��
8�X+'��pT��;�'*���s��@��炰4����B
m�<�����(缥(e��<.h��C�_�<��@6;Y� Eƀ^pT�tƖq�<����0ւ4���˿Af��E�ZH�<)R(6��M�"�C<B
�V�D�<�a'C?B�ɠ�̶4r�{&M@�<�m��Q��'Яw��Ip
Ny�<A�a�
l,���I.4�� �I�N�<�f)�rP���!	�9v̽�s��M�<1�J��D���'�ȣD���T�<y���W"��ʔ�\"gD��)�P�<���<�\`���*�J�[�/�H�<�I�2���:n��<����%
}�<1TP��J���(H=m��5�͆|�<)��WƱ!��;�6�1u�x�<ɡB�8R�,+�����֍Lj�<�d�I�4�W���k�V��G�Je�<�֯D�,�zP�LW	��I��@d�<��·6�5�����6��y↜�w=���s�ʈ:�t�J�.�&�yR挗A�p\�q��.ۺ��GbW��y��¼^��MBf�'�Py�&ӗ�y2������z���)�\*�#A��yr(��M�0R���	Ř4Z�����y�i�	�O4���Ehи�y""ԆV��cA"�8��(:5g:�y"#�.E<�q�B֚+XPi�� "�y�i��A��S��;n<�s��Q"�y�-B�8�P�6�Lf�,��!��y�g�q��qc�EH��;%���y2DP�#�l��c" 6<`�(�4�yrжv�z5�"�V+���H.�y��_k��ItB�� !@�qU�G��yb�W�w�^�i�E�Qz������yre���n�x<eֈ�5�y�K/@���BIC��(��.�y�LĬT[�
F�[�u�Z���g��y�!ۧC�xQDL+���J@�q��k���&�ȶ3��l�7�۱�RЄȓ{*�!���K�* 3@.���X	��7�\���ʘ9>��I(ƨ¨�����.�i����21+�h)b��$=z��ȓ'PPu�C�!�0��Z67�6P��OP̰�vK�=o���ʔ�;�4`�ȓ|.�!�Q��	
N�m�nA�E�ȓ�3u�S?D����iŜh�j��j��e��mʹ�QB$ːpA`0��iI�R��Rc@ sn��u���&A�V
31�C%�WW���8"Od�F��5䤜R�71p��"O�� SF �^��ĨO�A�0��"O����
�<��8��璑@�̉�"Opq�Fݩ_V�E���܊@�p�``"O�h���:yZ���Dd��]#�"On$sWi��(%�����"O��$�=8�� ��*ÛJ�4j�"O�W �9¤��8��E(���J!� �j�$Q�N�2~��LgM��,�!�� �y���گ	�R�3(�:䐤�"O8����^$9�Ԭ�P琪P*Z��"O����-�*(��� �9��%"O��pǊح.3��GOD1f$G"O��Q��R"����\�="����"O���撈=��99s%�&~Vѐt"O�Q5�E?�"<B��* ���"O���Aj���pgÍ/LH�(�"O�a2�2z�2`�hN}(ơ:"Op���йW#��c�ֿV�׃f�<	��1J��a�a��D�8�+%�
I�<�%�~�$Ty#ɓ�4�vds�!�A�<�3�P�,���q"�t.��!v@_u�<�"�3�T� `-��8��ܘF%M�<�!T9hX(v˝=HO�H�mWH�<�U�<g��@1
��	�Dip`�O�<�w�E�g����C�N�H�@�#�N�<	��m5�����H��mac�U�<���a�I�L̒Qg�N�<	S�۬e��s`o���)�H�<�u#@�<\:�B�iB�QFH�<�W)ֳ�z�C�(E-
��RA�<����o-�u��.��W�t)١��~�<��A�B�a2�j�lx�3��8D�����։MXޔ
�-�C3J8iR8D�x�ϕ8k�X!�f�[�'�ju�:D������{Y(L��e��4 U�f+#D�Ĉ�o=�����O� uh!#D�\�t�Q��X$��Z?Ǵ�y�4D��@���+6��E@�i�%�/D��z6H_7EE*=�ekVkr�ڕ�/D���%Ŏ_�FH�B�Pr6��w�-D��J��K�H<0��f�/g�&�4
!D�����W-*��]ɤ����:��>D�@sՌ��z�n$�Ћv�$�� (D���5@B'C�r( �@5;t�a�'D���Bn��1xn9�P����I�A%D�� Ú.!�ڠH����o��e��&D��JT��
�T5��aĢ6&�-��j$D���V�,'m������T�� �� D��@v�)2fr����5L�Y�`K+D�PY�)�N�l�9	^'��-Aa@%D�X{�&X�bYV�c�	^��E��#D��0�(Ϛ,����JR��S��"D�Щt�T�T*�0Rc�I=.�5�1�?D��y�+M'#���g[/#.�"��=D�@�4JR5u���
D�����` �=D���V&��u��a�#)%���")D� ٓ�2;v\Y����2�ĥ���2D���J0�}�rl�;�i{w�0D���@&��	�LШ67|�<J��0D���0�ŋ�\(r�#�%Vː��j;D��+��"�]��I�vTh�@��3D��3��HY ��&���N�Շ%D��9uL��IT��KR��PB|���&D��r�Ŝ|�~�F�_+$r7*O��i�kرq�ڐ�#�ۈl��y�"OB�`�ǦE\�2t�L�����s"O��&�U8.Q�XӔ픿4�*�P"O�L���M(k�����^�5s`5x5"ON�"bx��c��{f�!��"O�P�'��(N��Z�g�.cG�I�'"O���B��*_b�yiw�#b-FX��"OB	{�E�>��ȁ�є""��S�"O� ��Ɇd���Ш"lݢf��E�"O��*���!y��7�\!�ȣ�"Or�;D��#�C��)2��"O����H(�X���&	�2�
���"OZ���H3��LP�.BS�,��"O�Rրˮ$}0���[2^���Q4"OU1ulT�-o�!G� �h�h�"O�1/��g8�QA�O2��Y��"O�SGFQ�C$�m��ϒ�^�J��"O&���,��Q�Nʛ%�V��2"O�A��߾]4�$iG�{ h�B"Oh�B�dP�_-�)r�kA�U	�"O�-ڤ�]�X�|ɄK�k�*QP�"O���Tn����Ц��d�dт�"O8� ��U�7���@�
I�(�0ʑ��O���$�"�@!ړ)��e��L8���>%!�$��:����*| �u����;B��'ў�>I�qa��3x�ā�a�X��9���<D��+�!�u��� (�g)���*O8�0�ŋ<�P�B�J�/��i�F"O��!�Ő�N$���/.��HqU"O���Ř8E@��
 ���It�\�x�f�(�҉�cQs ~���,D��R�CמM��(�o�koVh���Oh�=E��+��S�Ҩ�'OL�Q2iF� �!�D*g&��p��EN�4"Ԡ�Y�!��'f8j�c��4��uHd �nq!�$�|����%@s0���^!��ۿb����a���CW�<����!�D��(�r �C� r��Ǥ<!���*`��A$i�Yo�eB��ʘ?5ў��aBxY@��8��h"Qd�
Hm�B�ɭ9k%����B2�PR%R�FB䉈NP��l*4e�T���%D�C�;�>��ꛡ5���Y��#9�B�-jlLٗ���DO��ۣ�(����hOQ>)��hSnI+D��o{����?D�T�BQ�s$,᪓	�Y� �w��O8㟴G��'��ɻ�%��p�ӴЃ��M1M>A��?�	�$Ezza�q�ڀ�7�-h�-�ȓBX�}���1��E�b�  �Ʃ��|+z�:ڰI["��F�j�V����rďd��[ j�@fX�	{��?)���ΏeVL(Q��&H����� �[!���-qHF �<%eV<�@�W��2��?�g}�d�k�P�R�E�1
@�`�@�TyB�'��D���F�h�4M��I�1f��'���53H��m�ãދeh���'�V�Spf� ��3�b��%��'�:�`ӌL�|���3��O	��'��ɓ#y漡����J<����'�������;�.݂��A������?���L��+���Y��������a i�#�%�D�O0��6O\���K��.��a�G�Ǭ �)@e"O���W)
%�x���$+��T��"O�rp�6�5R"���[�"Ot(���� ��]�A��'D�@��'~r�'Dɧ��8���-��#�d驑H��O����$4D��㵆�6B�T�ZF-�=�a R�0ړ�0|B6�B'� HQ��	}���w��\�<I1��)<��i��C6����	X�<Dh�:�z����.�n�H���m�<�B���"&Z8�vb�-}��rAM�h�<�.�\6�����Z���պ� cy��)�g�? >l������@%kҨ�@�͢�"O"x�'T�<��H���@<z�F�2�"O�1��lɭI��uq�m	(Pk1��"OĴ���X�!��b�*Ưbat�a"O8 q!����`JH�elQ�"OB��s�	rx��
�3oc��T"OQ@�O:,Gx�J�D/�����|��)�-a�Ĉ�΀FN�|ae	�-bj�=Y�' �<P���WJ��!wٮ����m���Нk�h� _o�1��+���K��B"J\�;6.�Q%�E�ȓ<�!c��S�
2�9#�,��[��4�ȓ� ؛���[n����N�=�B�ȓr�m�u�ѤS�P����
�<ړ�0<	C�4���� uI��e�q�<�m{�R c¬��k�
��7�Im�<�SFƿI�r�Z��M�
�Z���j�<aG�ڸi|ap�l��O���ϐ@�<I�(oz���
A/h�T 3 #T��ᝢEA� �C��9H�(��b8D����9g�8��T��;�զ6��K��<�b+XI��c����a[�o4D���qO��U��*�K�V:�3`2D���F�]=P0bQ Q�:�!��<D�l���
8x�i1��		7f�xt�?D�Db�h�s��aӌ֥g�:!�Ҥ=D��!wA��\��D�pkF@�ai:D�8ct@<?� es��/	�<|²O=��0|b�JݬD�
e�� n���pk�t�<ɒ�k��9(4��30#�����x���<���r �QW
N�"��gs�<a'�̝,H�܈��YZ� Q�2��U�<��N�
6�h ���Ƃ��E�q��P�<�p�J_G~m��IA�X@��)�u�<!V.Z�V�d�C�S�@e�X�7��t�<���@�ho)�g�Wd��Z�˄r�<�&�-W���B,��`��
���T�IK���$??)S��PPp	��޿)h6�w�@Q�<��D߬�v�@��pӸ)��DKF�<u�ː]��R�̍78*(��"�D�<�eoج�F�re#
�!��9S���|�<� �^�6�SFe2���Щ�@�<)��T�fT�7ˮ2�%I��c�<��NY�x�hT5Sp$˖�_���$��I2�|�œ3%����ʎ�B䉧	�ĩ'��1.��Sed��r1B�I�Hb.�hV@�1RCX�dd�r̚C�#�|��jC��J��Ο�9j>B�	�U���Nچg$�J�]8x,HC䉒kF��c/P�5y�8moG �C�	�F2��sI�?c���@��)�B��d���K��<E�XMӶG�C�����z"'�"g'XE	��N�Gq�B��!a" ����i�ꔳLf߂B�ɓ1�p�Ehґ9�hBȊ������<�'��!�i[��)�-T�p��\���n��҅Ȗ@�*�XP$ͷԥ�ȓք��g^�r���FY�<-��i�|�"�<[��Z4
�.O�Շȓpk��I_*
y�J��֍q�ȓG"p ��.T�x�eY}T-�ȓ�� v��oR�G���}P��I؟�͓P��ثT���S	 d��b�<b�H,��_cԨ�ŦS�?Nd��F��[ǈ�'���IT�S�g�? \ ���``%Z��K$,HE���'B�t
�g��D��Y�j��.���&)%D�x:tƃ<5D��Q� ^�b���#D�|csN�h��)`(ۚzŪA�.D�h�3͈"C�$�z�@XyJ��(/&D�d	WF\�0&�D00)��R"�`�):D� �AᄭG8�
�<w@��q�3��'�Sܧ"��� !*�4)�1�r�Ɂf*�EF��
�fĉ��C7�M�* � C�Ʌ,�}Q�#��z��Ц�*B>�B�	K;
��댍5�N���iΎ��B�	�d#��&뇔�6�1�+�(hB�	$R�rds�"�#K�4$jc]�q�츄�%0!a�Nr�9U(��3]lUD�'[>����iG�� �p]�=X��!ړ�0|r��"%���@уԂYְL�%L
T�<I�ǻ7�вE�ݼd�੺v
Z�<eo^�"��th���#?8z�1SJ�j�<�W�H�.�xܨG�Z�j&xD�5�p�<��%MĐ�0�6Sw���ŭWk�<w���g�Liӊ�&��!�S�<)��	*3�	A��_�X�"��N�<Y%T�|�F��!	��=z,�p�H�<��ڦG�r�Pc�ܴ{�xr� z�<����Kk����ʶj(� aUs�<a���
|]�A�28;jѱtʊn�<�I�:�\�s"���'/���,Vc�<y�훊I�ֵ��W**�,	A�G�u�<�Bv�¤�c�-��	PI�n�<�2L��|b��T�Q. =�xr�l�<i@ݰjYJ)� �+p-`-bi�j�<�bꀟmر��¤P��"�e�<��A]l )�@I�"�c�j�]�<Q�f=e�@!:�ےs�&�a�fq�<�H��[^�(r��ߑ/R���Oo�<	%�O2/�Ҍ��F�7/��T)*MT�<aGo<T��P��Z=f	��P�<Q�GH�?�N�����w��X7�w�<��"
�"��C��>6D����W�<�O
,x����H5��d�\�<%)Ǟ�p�['K�m�,�{'�WW�<�c�LKD~���g�[SN@N�IE���u��S�ҕ#Ѡ'av%��%D���g�pg��L�8{1BI��5D�X��װ���AfN��	��(D��pUO��`Q4�T*���XA`&D���tΒ4�l4$o=r� #��#D�[%�ǶJx����*J<� �a<D�DɄ���J-I�%��\l�f��<I�JZz��O@�B�M��B^�49��tD�3�X�wgT���K�4dŅȓ:6��"��v+ɂr�F�Qv��ȓY����F�d����1�Y�p�-�ȓ1����� �/�4P�R'�2��ȓ75����ݜz;��a�@Y�|�@��ȓi�PY@�,��^�9��+j�nh�ȓ�5K��,$��QA��3Lg�A�ȓy*��!Ǫ�oM��
%��/TYD���e�dZ��Ǚ#ˆ���¬-��ȓ.��<b��E)Q�pb�P�C9j���q�>�#����j�A�� N����ȓwNxE�0�_�������� �☆ȓ(Az�a�B�e�>���D�"V�1�ȓT�&�p%f
�N�hr���@.Y��S�? ��k��`�́pc��.l��g"O��!U)�a!������b"O&]2�'�.��E�!���a�+g"On�C1,�:b#��B�$K|��b"O�Y����-�B�����N����"O�,��ȳD�|x��O��s}��Z�"O��2$ϓ[	�AC�M# z��[�"O�Y�T���&���ȋVx�A35"O�D���cՐ�1֣�S�b�"O:�A�
�(��1,�= ��"Oteq���\��hw�	(#����"O��2B���q����끐2���se"O��c������L��P�T"OJ�J��Ÿ�|��o�%�΁1�"O�Qs��:�p�P#�RsꮡX"O��r蒒5O�T𗠛�����"O�YQˀ'|o�A�/@]�p��s"O���0��-zo:�yG��%�(�C"O05�v/�24��Ё׌G/#n�5"OݙӉD%M�4���@01�j�z "Od�� E
�1�.l����[��V"O�y@艈-��m���4�$���"O֔����A�(�k��=3�z��"O����_�����d]�Zg��7"OBH��ۥ5D��Hb#*N�\{�"OjX�Xh@�`������*L��F!��6Z�,��3`��r
RdK[9&��)�'|����v�M�.k��C�WFd1�'X��@G+�*
�2����N��Uj�'y�xq��@ 8��RFL�@�a�'x���@mYA���QM�:�H�'5dP��K^+����͇�@0R���'��I�O'`�`�ǌ�^���'�yB �E�z= \�ϸ ��hs�' ���&��)pB�	��[#r�ȹ)�'��A��BO#
��y����u�T@
�'"LA`�D�j�p+�^j�<��'�#NX�V�. ���9A@�'��H�C�y�
xq�h�	(ܜ8
�'��d�#H˕M͢��OV r�H
�'����2D��;,Tj!f,��OE��y���7���ԍ�9��l�Q����yB�\1+ �+T��dq���A�yb�ہT���9r����ҵ�N:�y�dX#� '#�\��k��y��;sN(��r�
��U�B��yr�A�[l^	��(܎`�&��%�Q5���hOq��l�C 5h��6��8�d�R�"O�E�uǈ��8�S�/��)�#"O����;��2�AƌJ��)�"O$�a��Jrɞ��s�[��i�"O��h�	�Wp�k7��q���B�"Oډ8��Ĕh�J���E�{�ZH:�"O>��Q��E��� ��ܭ8�
l��"O��¢�Ⱦm���X���Z�2��A"OV�l��S��'k�1��n!�$ֻ{*���&�;RF�(� I��!�$	�5)t��R��!F�<�g��9G�!�dF�ncn��t$�f�𰴏ǯ{�!�$�I�r��hE;{2	9��2s��5O!/t��CT�Yr����J�&	!�d�6z�,��e�]�[��A.H=Pb!�'�>d��k�=��t��#[�$!��*.ې��Bƭ�L(B�L�J!�� �p2���T'���$��lP��8P"O�#�=Vd`�kGD��5H�d80"O�a�1ND��b&-�l4�'�	�3�6ȓ"Z�1�Y���ç��B�ɜzP���U��k��6UXVB�I�VG�Y���N�v-��0+��
*.B�I��.Q��JG�V����%-�=GnB�	�/��Ղ ���� �1�ZB�	�~����C/�p�c��Ku�|B䉠~�|y�"EU>nx�E蓊�5�pB䉺�������3D�bE!��Ϝ!+8B�	�aL2�C�̈́JH�Ypȃ4P*B��|�򡸒�U*<8fd�f�B�ɂUIl�Pp�S=>k @�Scˬ��C��60��j�'ݿUK��a4 K��C䉨Vٰ�O�F���p�ܩ{��C�I<;(j r��9f.�sQ�3|C�I�S�T�J�����D��C�a�vC�I?4�vh����/�lLѕ�(E'8C�I
&�HA;`���A�}�����aJ2D�$��G˃3��C#�#,b����,D����@�0|�R-�5Ĝ�8��	��)D�,h��,)AV��v.Y9j��]���%D���m��:��;DH��>��q�vo0D��r�a %o�~ȉv�_4����.D�X�����Q��o�r��A��+D��(�ၫ�"�j� ٠]1 ���&D��%_�	�0m�@'V2���A&D���b��|0h6�	�2�6m�q�(D�Dф�2�X9�KF���P�.&D�Ha�fI.6����D$k��D wO9D�@Ҵ�@}4>4��)�cļ��4D����gL,I���`����vT��3D�X	F� �~�p�E
�I��4D�$��UND��`�fP��<D� K�/J�o���P�]�T�<�a:D������4!*����$�-	zT`F7D�8P��8���ՉKQ`zAS`�2D��� \�#���qSkJ�{�v1�51D���w��rd}x��
�E �+��$D���E�">��p9�DJ /-�B�.B�ɡxԦ@�A�Q�g���z�T�>nB��$	���@���8t nl-�#fuC�V�~l����G�<<��$�S�C�I�T���3	i�\�˒�ς) �B�I�NY(b�]9�HTA�M�?�bC䉾L�jaS�HPS..<�q�U�74�D�O���d�&��s����3�)�'|e!�Ě�F���hc͍�2�0=sg�8&V!����`��Н+�x��eRM9��U���ɧ�Ϥk+
�Xg��,�����%D�0Q��F7 ����/S>�n�8� .D�$3U�Q%0y�pRP瑃e׊���-D��A��N�*)L�y�C�aE��z'@�<�
�S��c��V6p5�����q��ȓ4x6rB��=�����֫(8��ȓNm�W*�Yr��)pR���ȓ�^4 S�p�|� ��#D��a����Dـ�P}�:����X�~��ȓ���u��0/	�ۢ��_X<�ȓ��)B��U�o�ʀ#���k>D��ȓ'�<H��)�@�n'A;<ńȓ��)�D	��X�P�RUɝ!{l
Ն�2EH�U�L��2QG@ZH���S�? �e����La�!"#K�+4�!!V"Oܡ�eM�*T���*H !�m��"OR�ň�/F���ҨB ���"O^<0��4$�dCF�H�c��e�b"Od̘W�ѣ/D@Hc��qg�pȅ"O�4c�,T�]�$�*����cc\��P"O�1��NY~ $�"��J��@�"Oȑ�0H�dv�\��Oͥ9U��"O��;���u��K.N�(	��"OT	?/ļ��RFޭS^Q�""Op=���.Ԅ�Ce� CoZ� �"O:���HU�)�D�iJ����"O؝���ٶI������?V�u"OT�BHȴ$�L<#C��=hZ��{�"O��#(ϧW,@2��Ͱ>�B8C�"OZ�Q��^2<d�@ �K���"O��j�ix呷OE��Tp"�"O\ �r&F��f��,C-Z�fAv"O�M���( `�\�ԩ��1z(�*b"O.��p���p�!FƐ/>޴��"O {"�K�D�V"�/R�&���"O�c��i�r���Kȕe{nQHt"O䠩6��=yS5X� ��r	Ȅ"O>d�ׯ��+jj�j�N��uN #��D.LO,�9&��1 ?<�!�Ne�� ��y���-��x%�¶_z�({"�Ա�yD�>\���j�SA���9�+���=y�y�Yu(1�G���N����v���'�azB�H�{�vX�U�6?o�L�1�S"�y�!�-�|�#%�6����D ��y�֫��%�5���R���hO��D)�*���8 �¡F�S:p!���*k��5J@A�.���j[*ug!����޵�iNᬑ �	�e�{��'^���<ZF��f+�3lt����!�!_��D.�D�a"K����Q؂-KP�j��>D��p3:^8B-ZٔT�@q�cM:D��BPԈ6�kRFՉn\��X�@7��a���Isk�JM���v���~�� �3!1D�X"$υ��b�Lќ�f��-D���Q�R
j���V,Ta�<qKĮ*D�4�u�֕Y�B�S��4r5.�j�l-D��)R �jD̻���h�J��(D��x��ӜothY2J�4o� Q�e�+D��I�#Y0%>x�E�=wn2=���O�B���A��xH�,B!����4/'�C�I�R
�CS�V�/STI�҅+_�C�I�~�1��MP�����&͆C����+% ت/��8�)ɻ#ZC�ɿ/r��AGoŏHe�	Q&͓})�C�		7X�,�v"��V��9Ko��f��C�4]�z�ˢ�
��x�i�B�2q�'Oa~B$R�h���qh�=`d%WG.�y2�N�?,<�Y�lS����,�y^�P-��n�v>�������?9���0?��[�CB_i��xZ�ƃ;H[!��A�	'M�я�I���3�ܬI�!�ۋB�Qav��9��B�Uj��'^�a��@!Ԧ��E׉$o�����'�ў�E|RgD0��0a߹0=	�)R �yb*Tx�#�.�� ��9��	���y��5\���'A�}�HH ӡZ��y��N�W��(��_�s�ܕ���i�!�$E� V8�0��M��|؅F���!�� D���n�-Z�����
it�B�',�O�Y�0ǈ�X�`,�5fB�)R�'o�'��3�i>U��F���ܘ���:x��Tj�<)Eg�pnh&bK�y��(aDdh<ɲ���}JD�a؜9�����%�+�?��'#��d�ǩD�h��ϓ�t�*���'@�-!Ч
fs,M3a}b���
�'��Z���8K\=Xë��vШ�{��?��'�0��i$6���j��*q���1�'�����qM��ӗ�F�t��@�'o�E!p���1���&��>t��z�'�����_�~eXȃF�4n��d��'�:�Yf'		����UA׷e#n��'o�����J�N��eM�/k7�hX�'n 0�'!�_V(dCGa��QNj�c�'�M��Z�
�iSf��E\$��'�<C�,]�l��J3��{��'��x����8<��'D�y�ZD��'�(�xB�\���*��lm�]��'V��HӃ�&����@�/�>��'��IB�M�������� S-��'���� o^�."�y�D�ͺ�0��'��1µE[4^�^���;l����'r�z�P�v4`Q�AO�2bYX�'3z�p5nA<��)�a�+#.�]��'O��D�x%t#�lQ�  �	�'�!"�'�^�t�n�"���Z�'$V��@F̣+?���w���8��	�'1�T��_�"uN�s� ��%$X�'�8��ˑSn�ͣ�X�1Fn���'�`��H�����ɑ�0��eS�'�����z�,4yā^'�zH��'���Y�J�!h>^�2��B>)�0z�'��{uON/Zd4��N&qĥx�'G��p��-/�a��#�J���'�8p���Q�D���cE,�Ll&m��'�<�0jـW�í_p�X�
�'��؀fkM�%@P�p4�G�|:�̘	�'��QHӣB>~ ���Ưn�q�	�'L�5�"ˮ[�.Ш'O;[S�)	�'N���O1N~���6o��P���'�:�R��!��D��K�{E�T8�'4� byN4	����e���q�'R�	��h΂)�����E¼���'���؄�Q�G��s@�Z�_�f�
M>9(OV����y( �ᰏ��>���(�jшs�!�DE8(Oz���1�x	*3鄳.�!�d�1G����
��Bz����6!�D�  Qb�5&��[_�M �FŒ^!�dC"Fy�EG[�HH��i��	M�!�d� N ����3ILA��I]/?J!�$�41��lڦI�-P��Y����+:r�'���'"�'���@�!%ֱ�� �
7�Y��'6�RrJ�+WD�i�d�xv8��'�zH� J���N���X�r�Y0�'�v�[U�ѯp����h� }P�'�"��a�F+�6K�K�Yun��'�j1��n�%�i3����L�����'�q`��(z�P��ԘM�XM>i���0=Qaݹ0��	ڴ�X�b3��
�m�d�<9�O.?�`��S̅ ������W�<	S/\*H�z��̇/z-����S�<��'I/<F� Aċ�����O�<����"�Us�j�
n�=rŋO�<� \८U/v*pPcg�F�4�!"O�D��hCa��s��:p�`��Y�P��ɀ0A��5^�Ti�oN�`$�B�I�|�1�B�O5�$i��Ϳ�B�ɨ}de�E��+n蜨���'L�B�<!��ə�!b��X'
�K�nB�	J3��y!�S����R���C]:B�	�к (4��,Rی8�͵FOB�əd�X1+�Ʌ��$��+���Ir<�@a�-V�z�p�MDx�X�# d�<QAƌ�v�.��KK>�}S!��h�<s.Z6&��ƍk�
(�3˔[�<	��[�L
�$��(K��z� �T�<I3�0}_>� Dbْ1�,j$cA[�<�Vj2?�tk��ގcx��� �m��^���O��d��ضR��UX �Whn�y��'�!��C�K���A�B�`�����%ƛ#^!��	/a� �!���pK<���AR!�d8R����W3:$%f�W'C!�$�8�TLJC��`Q���AO� !��F�ޝ����\*}��ڦM
!��#��x1P��q�V$Ӕ��:f��'�ў�>]AdNL5S��\�����`APQ�?D��F#�O�,4a&�Ã}�~y��#D�� u�T�@�`a��B�����h!D�̺��.Ξ"eΞ�%TB��;D�\�MD�Z
d����;�B��"I7D�谁�#���3�8q�`�!j(D����cEsW�0�pKT�s�p�V�3��^�'h��'o~�㗆@-�h§Fk�l�s�"Oxh!�o��5�i�`g�I��y��"O�m��)�8#3��hUf�
�$ �!"OJ�с��&3�^ ����HY:9�"O��;��t}aY��<�dG"O~�IP+HtO�QG΋�u�h�8�"Oz����8[���3�DpNi%�r�	���O��1�lCs*L �釴y��a��'��`�4dWe����rN�j�L���d7O�eZ'K�'�.�b��,���B"Or�Ї(�.�X��v�0zJ�m�S"O&�ɰ���r:Ѹ��͋D88xH""O�)��ˊuc���v �4�Z��WOI6EЯ@�j��ׄ]<qI����*��0|J�"���x��ҏ!��ĉT�Nf�<�A�޸H%�l�4��9�!p�K`�<qGF�,2v�w�"	f �$X�<aUȚs��Bu�Q!H�R�3�m�R�<���-�N���,�R�<�2m� <X��L	+���'�K�<�0A��k�[�l�$]Z�WHG�<� BS)�n��p������Dͦ�y��̍B�Ș
tn d)�����2�y�GQ�wD��$$s�T�+�
���yR	!�Ƶӵ ݙc0�y��-I/�y�a<
��Ux��ڻ_���iΆ�yr�
CQ�A�g�Ԕ\�(�`R���yba�
-���ֵ
1\�s����>��O4�h!��X�����g��T!�"OD�ggX�l�R����9�<R�"O�l��/�!Y���d퀞N��}	c"O��x�B��,��8H�Ru�
M��"O�i�D�ժ~�B|8v��?�R-[G"O�\���+ �܊���)\��!aq"O�P�a�ȲE=���Fn��c��pa"O� �I�d�S U��M��U�����"O�Ѥ���p9Z��ƍƙ@�J��""O�1�åީu���Vj�����c"O^���/T�R�d�T�E(0rd�Aq"O��8�+Y�QEx�RB��!e����"O���`Q:U�h�1!/�1iH6�J"O0U��������#�[1B3�*�"O��	�B߀?fE�o��"Ơ�"OL�����:��ճգL�Y�m�V"OV �R�����%��%}�4�{�"O�(z����nY"�2*���Q"O�dJGHф��:ĆQ*�Y�"O�=ʆ@MGrNui5%�<� "ON�HԠ�	s�����H�/Je� "O���Ua�7@��9i��ș��`;"O�@�UMR�r �<��.Ҥ\9�"O ���S0���r�N�"[�G"O�1ۗhS�C� �����Z؂��'����cĂ�\v��e!�'Y�L�'���U ݍ.�����S! |@U��'��P���!j�����ʠ}��`�'�X��Q���Sb� �iw�\(��'T.`���"T,��FDѲt����'��}B���C�r��J�x{(mJ�'FE��X/+�m��J[�s��	�
�'+��"b�	}jDJ2c)ZψL�@"O���ǭ��|�e�2@�J��"O�̙"-�s���P6�ӊ@�����"O�8�w!W=Z� |��,۪�H5�"O�X�#7����2&�=����w"OE���]�`x5�@
�Z���@�"Ozh[ь�:-�J�m�:� �f"O(�B�.vxi�snZ��jp��"Oj��PE' �����-b��d"O:聖M��|���$l�$+�T���"OX	ʄ�G+R��Ԩe<@��JU"O�t�Q恀��?�p�k��]X!�ޑF���O*,@�Q�b��W!��v"3a)��A�Eb߂V�!򄘭[I�X�+��,��-ˣ�� �!�Q���Ѐ��V��	�*ӗ(�!�D�=>z�B�	��Z�L�[��>�!�d
�Hdԥ�2BǽY��eb��Y�O�!�D�'W�`(σ(r$�Ȥe�"�!�D*)#�*��V�P�9�eNz!�V* ���w��=��H�Dn-q!�$Q�o��-��Fq�)�^�wm!��N�9��(y`|6��*s`!�˾Ur�(��b*�"Ė�O�!�d�2iL8(�E��J�rQ˅�N(Z�!��0����`�,m���5��d-!�Lq�X��1�P	h�k*ԃ�!�$�<K�zp'�"�����.�!�ʹMx���K�rt��(�$��!�$�m���SjA2otl<9�A�P�!�$M�P� �bϩ@g|�i���
s�!�)I��\����`(\!Ɖο+�!򤌳U]rf�?J������P"w�!�䅘2�����|�Bg
r!��U�9f�j	B����Ʀm!�$ɪDWؙ�BRsȤ
�`C\�!�ۙ̰
���R��Po�	|�!��S�,��v�TL��eba� p�!�T+c��t��jp?�ЃW� �!�� T1��ַ��+0��1@��yh@"O����\�nR��Hv�ܳd�b��"OA��-^� �.�;C@���"O�����_'A��E��C�NyL�A"O�m�F �>I� E�ua�qi��"Or=�I̊IL⩀��C�/Y@ՠ&"Ob��WA=s�>4 "�L&*�ʤ"OL����y/���g䙕U�%٥"OlX�J��|ܦ��"DK�H�Nź�"O���;�T�𶂒wH&�b�"O��Ћ�OF����B���"O�E�֤�!%�R!q`�Ǽ\���i�"OQ�$�-9?��u�3�z�s"O������[prͨ�D�T���y�F�-
���J-(��Q�V��yB[7T�TS�]�%_���jM�y�	TV�t�c�^�4P�x�����y�,�)϶yx�m�7/a�s�E ��y���,W��"P	�&Ƹ30$�,�y	ֆjˆ�� ��*5Εzr)�&�y���_��P�ԯ��9ٰ��'�y�ɗ=7""���JΔ��!@0G�y�$V ���'��C�=��̓�y�̀Cq!���P?�Ӷi\��y�k�r^�PF�T�: �8BV፡�y��/#b�h��X"*y�u�Ł�yR"�6%�|�a .\'KO�q4l��yb@[�M:}�pN��,�R����yb��nFn
 �Z�/��c�"U�ybE�2;���w"�;|�m2bU/�y�+GG=du�Q��5KU*q)q�T��y���n�Q�_-��l��yRf_��PQqA���p��d/@=�y������h7����0x�bnِ�y�U)	v�i���� ;�0AR�۱�y/Df倘HwoH.m�&��qcG��y�Cļ2�(����
Q'�h9��ӳ�yh�'W��b�؎yb���ቆ��yR�
L��Aa��t��9I @C!�y�k��F�y��Ǖ�>Ƅ��N��y�.�V%�i*��Y�g����W��y��D�e�n�f�_A��1�g̙�y��\�vrjX{!��a���C�)�y2 �+W=x����t��K�ʍ2�y�؂;�x9Ҥ.� ��g���y��$^V��� �J(b��u���yb�K#!͎�`�E*q���ek?�yRخ~���F�f�~�	&�M��y�dK�EP�b��4H�����cO�y��޻/ ����@��>��\�o�)�y��Ԓs�y5O��2�\������yRmX�:�ڈ����%-�����y��ɾi>�-Iƣʢ(� Y/��y���j�jR��%^�<c�K׭�yR(��n�"6 E���{a���y@�չ���C��:A&B�y2�Q?0�6�77vi2!"��y�����za�_ }�D3SB���y�HJ*(��WnW�l�,:b��y�@΄��8���f1����$�y"��A��i:SB@)ޒXx��S��yn�0q*���C�� Q(����y��}�6���c��������y�HK%�"���X�|�Z��F`ΰ�y
� |(Z�(MM|���N�v��\sF"O4�R��w4�T��
�U�0�c"O�+��=]:J�"�ƞ?fn-��"Ox�Yp!�!0�xRƆ��V��"O��Յ��"��sC�d�N�("O��#��!�9�HO�R��=y6"O���5��r��Hᒩ3�H@Y%"O^�i���d\� ��Ŗ(N}�-KG"O�,�E�\�*���;V͛ʔyk"O�-ҁ��(�&܁�gED�༚	�'���j���t����cJ�UCn��	�'���Q����0�R憩^ �y�'k�&�(K2Ĺ�M)@Up}z�'���F����2��$��>$V��	�'��\�q�
� łѸ)ϼ��@k	�'��DE�Ʉ�9G�͒��N�<��%͞�(t�="U��AdCE�<�Ϭ^�L�� � W��(�u�<�p��l�lp@�J25����G�u�<$NK�}���yBB�*q?(UbǮ�e�<�pVS��0�f&|!&�f'�{�<�%_+�r�1�%K�!��cV{�<!,R%+[f��Ġ�}�b��s&Pr�<	R*�13��t���>XI��DF�<A�fӮ������}��"��_�<1Q�P[(�!6�
��� �V�<!���6�x�ZL����DG�<Q5(�;�n,� 'U�=E���qeKB�<ӭ�v�ĽRwa\�<e� Q�ˀ}�<y�#@�j�閆
�`�*��BD�n�<��膑M2V���׭%-6r���+j��E-q4��Z�A�2o�*Ɇȓ\�0b���V-ȱ&.{Д��7�Q:$φb��}����=���� P@b"A�l8
�(�K#f�fP�ȓt��mib┰
�^I� S�r(��&(�Ѡcd<E�<��� �܆ȓ+����#I.Z�*c�	�u�a�ȓh8�`t�ŤH~4����f���\�\`R�#J��AV�X]�L�����H¶��J�Dx��P- f�ȓrL�B+;'���IP�h
���ȓ�<aCg�u���s&ʝ;8l@���J���p�gަ-�e���;@���ȓ HBiJO�-�XD���!��ȓ �Q �?YD��dQ�z�Jx��FH�X"c����a� �v�ȓxȨ��vI\44��Y֍�>;*<�ȓ]�$� �1:���@R�x�8p�ȓv�N�i�-Yt��Qiش^����ȓ{ hxBC
9Sj���w	��T�e�ȓlr�1����Z�؄�WI pL�I�ȓZۊ��G�P�ڈ�7d�!@q���j1h�J��,)ذ�ł�hm�ȓ ��Vj{WP(bD��M�@�����T�e��36�y�$WK����ȓ@�
S�x<�С����@�ȓf�d��u	�-}ԜQDg��@6>q�ȓv�@m��&X7	�,{�	�.�N-�ȓd�uHV)S�@�cVHs�e��e[08S��T�x��%�1	�u�ԡ�ȓ>,rk�![Tjl� �$7�L%�ȓYdm��p
(T*a䇟M"���J�v����j��QH~t���S�? ��B���6Z�4���=&r(�AW"O�B���k���ɘG$��q"OF�{�&��}kR��qd�4;��y�S"OН![	{�� Q�_�8���+R"OȈ��*Y&��%cS�c\�Z�"O��r�1�9�V��?�N�8"O0��E�8c��AwF�{ϸ$[G"O2�C���p'���p�X4�� �'����[3U���\4n��T��t��'h2A�(a�N��S'����'�ƭcf�91��$�sj��F���'�f9�Vd۸:vj]i�IR�JYV�9�	i���'����_�7 �1a�۝ 6l-��%��i0W�*��2����ow25��;��`��E��/4��� �A~�>��ē���4�<����q�ժJ�p�$�eH<@E�k�|�LF�b�4���K�<�+ \(�����?V���cd�D�<�R��)b�h�i<�pԋW�x�<��A��g����b�L@�x�t��q��D�?�����pq����4I����$G����k�0�p��s	k炇:e0��<���?�S���1�KP�G�Va��ـ"�C�I/˨t �h`� $A
1r�B�IKH���%�2�,2��'e�����)�I�o�� a@�=X����z索=1ÓMlP�z���yP���/��E�<a���0�WM��&V̠r��ؽu"O�D��4��� -��	l��F"O����d�+_���* lO�N^t�b"OrI�dc)p� ��&!ǶeơI��	]�Od��j�h��Mᆜ���\�9���'�d�+A��z90M:�	Ğ-E��s�'n�P�����x�9�Ј�K>���	]�]4��"	
#0Q4F_![��'a|Rō/	�ΠQb- �Zu�yz���O8�=�O�����ȚMz�i��	�8/�13�'����
�VT���gB�%�����=D��	��K+VX��T$^�1�h[E;D�4�"$\>&_D%c��� s�B�,�|���I��J!}�2a���(X��zǄ(D�x��I���Z� ѣ68���a��Ɛx2%^=b�Dl�"�[84K�xR'���y�n�.%N(l��k\�b�u�#^:�y �3*����V��Y�`:6j���yҨ5����g�N��q;u`Y��y�D(i�乢eۺGg@�D���y2�!b<�!���0Fd�17NG���x�j�=O�b��V�Ƃ[���s#���$�!�$U9+�s��N��8Q#bJ�"�!�	�_�<T�!h��x��IKG���!�$K�:�~ap��W+&����B␰s���x��d�gD�6�J�ǅ�R9H���
>D��P���$p|HC'C;aB֥3֭1D�����V^؀�� )���v�/D� ���>�6�C�mY(r�r�a�gL�<����S�`��# �!{�P@SѤ��o	��$�>ьy��	��I�Щ�K�2_q�l*S37�T�'�p��D	��с��G>l���c!���?��O��GV1&�x�fZ�2~`�#�^'�$�IP����C��	��̀%�C$a��]��,ړ��۸Oc4�K@�ϥ,1�) n^���tR
�'��kq�ϗba�!2��̇"�,8q��M��X���'-���S09n�kC���z��5�өXj���hO�OH0�S�? Խ��J�7�2�(3��
�"�#�"O��c/ݚK[���Т#�>AS����t���O�X����14�~š�h�?p����'*�����Q�3�p��(�4�VX�.O��'r��O�����/@�2m��%�x`�U `�9D���U���	��V>#n`u�Uyӆ��?Ɉ����'M�0�A���T� 5�#È��0<���$!���H�遈 �ƀ[�DO�K21O|���I�T�P$%߸yT*�]�v���hO�O8��3nJ���n�*\,�L(����D0B�	53�R��'A+p�4���Lܹ�ؓO����2�8	f��<W:��j�,�:}���:O�H����uY�0�3mŬB����<�S��y�/!"�{�%I(U� ��O "~��Cϊ��%2���P��}�<�GOr�<�6 �Y\�ہ'L}y��)�璇�٨)H��dm��n��Y�w�<D�̣��(65����qú�R�K����O$ҧ�i0�I�^B�[�ȫK���F����C�	����f�����"s�2'�DԨ'ͷ>�!F~<a�kU)�VM��ρ�@��ȓp��EQ2_�^�P�CP�+Pj)�'��~��Fc����MB gL,�+�	���%?����hO�i��͠��S� $����*�!���O�T�Gl� �E�i�U���p"O`�
�g�wN@��m�[V )0�'2ў؁v�ʌ5�h@z�Y�N���'D�t�!kY�:ψ�0�n�n서D	$�� h�$l�ɕ˒=\��)Q ��i�|B�I�0Dpu`��H�Mʨk'��,��ʓ�0?�Vܪ,��m��CUA,��c��Z�<q���K��K�>����k�U~b.��O>��b�vjt %�`�Ed�*D��HB$	���p,��<.�<�&<D� b��-��`��Ł�j�Ӧ9��hO�Χ�L���CI��5'�R�LA��`5D��2�g!WJ^�"g&�o�Aja'�<a�J(����&�d�R@��� 7ĜH�ȓb𘧭Uz�T�X�&��:��!�ȓp�6m1 ���H�,�qoƲn/*q��K�,��wM@*� �Hc��5Af-��N��j�˖�j�~\�椖;.��a����s����&>N�b(Dc\�|����E-D�����H�B�(!�1o�s��`a�m�Ї�I>	��A�ЁN�,�P�kǥJ%�dC�	�y��с֭��<�@d0��g2|C��?L��h�3�T�Y�����[�"<����?�Sbj����`��0
�<%�7h'D��С!{��,Z���m�$u)��#D��V�R?@܌�PG�HY�p%�#D����a�w�&�he�M�s�ФSF�=��hO��.*{�"������`UؑN=D�,���A�.Έ�Y�,�) :y�ǆ�HO��?yI�T����$�N�N\5��c���':��xy�L��<� ��k[��$�+����y�D57�FMBgR�	L�᫶i�4�y��)�3��@�n��/@��0���
�e�ȓY��n��o��ec� ��(�' ў�|�aY�/]
аnT�[�85 ��_e�<9G�g����ʕu��<���{�IH�̪3��6��}�GB ?u�Y6��<���0g� �gR�`\"�`�.Y�D��C�<O��I�R�$,�v8Q#��6?�ʓO.b��Gy2��2x�Yp��������X��?鞧�  uȷ#2мA�!�5ek���"O�4fKϹE��E��O�A�><C�'�Q�,��b?+Ŕŀr�^�wZ=ɅK8D�$���%3�2���I��K#�#D�le�*`n�IS��'WZP8�# D���t��3g!�y[��L�S�D � �<D�Avd� J��+��P�[b9D�x�!b�3��h�JN�j"��Ap�3D�8a¬V�B�((;F�J.Z�"ݠ2�-D����U_�А vM	u���!*)D���V!�+.�șV L)����!D�P�cM�N�u�I�)�>D��S��^<C{�-`Fk�<]@�!b D� :�)[� �|з#�-Q'tI�)+D���%^WᱤM1(R -'D��C��8��T,��*�\]�$%D�����v6 T��ܑ"1�Y3�(D�0	a�"p틣?W�fA��,"D�$�&��	SI�t,@�qR!D����ȏ-��u�D�ņY�J����=D�T�����(���Dȅ�UO���1D�Xr�S�t������v�� �s�0D�$C��7F�)
�H|����(D��"b���� �U).��ȉB*2D����̕YyL"�(T�r�B(4D��zA���u/��4��[��l"20D� H�N�v����"I��b,�y�L-D�����$��z&��{a�mɖ,D���,�'x��"��8"b��k(D��b2���lv5P���1�J�à�)D�\cA��v�.EA��5;Fjx"`�%D��9b#�"z@h Q���.��#�0D�d�b'��7�q��Ρ�4U�t�,D��	��^�	�H%��H24��r�$D��b`��P���#��UKF�I@.D��C����D�"$D2#��A��6D��鑻�hC�*�U Pa#u�޹W!�D�,7d�Bg��s�,q	CG�w!�D^59Y"LA!90�P��"��6�!�L7�H�x
-9� ��N"�!�$H%{Ϣ���J��F�y$�RT!�˭4u���˷Z��TQ��n?�\��B%	��I���]-E��#f���A���t���7ǝ�<n�݀�&)D���'�ݫ9a�7	ض�<8@�L;D�(�IX�iK<��EY�&����4�*D���E-&����K�LQ�w�*D�i$���\S�-bn�M<�e(D���4h��[H� �qf^(�&1@��-D��sFo��&805�B?�4%*g/(D�p�Bƀ�K
��E!�
��X���2D�l#�l�>�%՝3H���.T�Da(�
6�X)�c6}.���"O���H:U�@;�ĭ}�����"O� Z3�۬w�R$�V�"��"OnXQ���Lt���
_% .�b�"O T��@�^������n�)�"OVT� ���@|Qê	{K���"O����B���t
�;U�A��"O�T@�D�cB|PR��" �䈊�"Oʙ�1(O-$�@I�k��o��IY�"O�)7+��N�d(���N���s"O>e� 
�')�t�x /\�:��&"O��g#Q�q(�Mb1oЍ����g"OYJ7ψ�&�b�Q2��>
F��"O� T�WiA)����G� *�0�"O�@��7;nIr��D�(.ZI�4"O���nМB������T�Ab���"OLdCҮ�ϐ��1Ý
~ió"O���D�޶���Qc�f��{��'�r�@��x���-Q�h��m�t`k�KX�y �z���A�B�Y�@�BK-��'�J�zb��my��#b�&?�	q��8�V�!��f�L���")D�Hr�9JTIb�"'�&,P�I�"��	
�-IwA�K�>!h�Ox)'�G�& ����lH�J���"O����NJ�.Z��c0�M,]�� �I=^�(��'o.t��ǉ;I��F}��&}���z4;\�<y�!H��<i苹Y� 0�v�<�;�L�[�|��Q�lw��B��U��`@���.�OHT�7m�;;´�y�b�I���x�`�Y�|�0�O2����ڙ$�ŊL?�FŊ�u*I)���*]�s�%D�`�1��NXX"V�)4�����֖���P0�P��$L��s���$!ks�����M��Q�q�"	�`P*l�B�;$�P��I_�K�������\R��K�c�����Z�tX% (��]�'�	fV`k&dA��Z�jg� 'K�l��$�r�P-O� ��`>{H|��f<�u�� P�Q5����@��p?鰉�8�pQ*�큸~f��S6�CW�I�s���\����K�(n��#C�~ʦ��`׍J����CĂN�<�4�ɼH������8�X�ಣ�]��$]t���Ň5��O1���'4�i���:'�DɤL��
Q����'x^�K&l�0�v)��b�)8ؽ���D
����~&�$�&h���(��Z��(��lk�C�:e,�s�� G.bb m��9t�C�Im%�k�oL�-�n�����((]�C��&�4����ڑWؒ��力�|��C�	�5�@�i`m�B ��WŘB~nC��7 ��E)���7�&���5I�|C�ɠ1�l�j[4��u�1O
>B�	](�E�	Y܄c�bN3I":�Oތs�"γɰ<��R�q�Hp��W*��	�%~؟��g��$&U�-�A
(��	p� F��Q3E�r(<�!��56�'	�#��i���L�'��m`���bt�t�|
"� �p��N=*x�0k�L�<Q��[�e�dD��h�~p�q��c?���'&p(eK��+}��i̭@(ֈj�cQ1ws  ��jǪ-����D��(��	>nq���*�.4���8Wh�w�
�'j���.�q��D�Ď ���L�@@Є�Z�=�D�`���@���?�P�h�@]�`���9��Ȍ9�6��b��) V�I3ٌ��ѣ��c@ny �;O)�ab�G�YzQ���Ѣq:�	�!rX��P$71�*�#X0(]��L��g��A@����Ǚ�[������AsG<G����)`|���� .�\���D�~"�
�X9�v��0�H0\�v�ra��Z�2��]9�MD22�����gi�a[�1�1O����\�gG4	�c�M�B	�t�>a2FG�4���:��:ړk��l+#�Ҡd*��c�O�[`|<����^ -
&�ؘ2P�Ģ%�'O���P�1�f5�	A"h*��dj�'9z���M6��*5x�'Z�Xi���S9��7��}���[��6Cږh(V�?���
�kvnc?E��C�64���
2T=~aې �>���Э~S���a+�� ��ЀAÛ��)Տ^�2, �O�4���H3e��	{�(�5K�l��'�0�n	�E��;��ٗ����d��d�\dH�;Q~�}���M�a!F�	�D���+��GY�Mr7�X>{@|��_10��?	i]�a��������M�al�"/�h4Bd�^([� ��@�H49��#�!C��ҕIQ�	q�H��n�0�|"��)Qq^����غ>� �H����8-��b���R�c�k��vJ���r�,G=N]�A&��m�N�Q�$ɧ_�B\���G'9�ڤ��ҽ^M�l�Չ�$~��}���a��1��H�#�Ќ�G Ѣ$��Y2�o_(���`"�L�x5*��%c��-���N�!�мɧ�P �y���I��F70D��Ş,C�Z��I�7\jy���π6H�;u+M�.�bV�ɓ)��p��ذU��p�"�@�g՘��N�3B�U��,�,*��Ȑ/�&�N� �2�Xg(ƗA�t����I"��O �$✢U���F·'������ �X���T�U�K����aKM�/�jp�%�P-IN���O����L��,$\�����D�%/��ѳ%�GM�����J�$��I��!7��,��<{@��$qD�t�P�p�*�����3 ��t�c�G#U�Ҹ�ŏG
D�����8ql*EhL�Y��x� ;T�� ���ua|0;�_CҮuX���>�ԁ���l�"~3e�fa�:G���+��\�Z��C��j±ϻB}D�E��'0��ܙ&�횴Gz�� =%���"�Ǆ�p�謊Em�.'��jSk�2l�XsW��)_�>�B)�"2����6p�����m/%�뎍�Ϻջ��@��� uo���ϡ�"�B��vӸ$K�����Z�&��x�� BЌB��M+��K3^�>�a mB�EȐi�����@�R��%�C��*py�l�7,�;��,\�2�YP�	�:7p�B<g���5��!p�O�%[�)k�������y��2t}ℒ6�J?\��BGF�g��1�Ā
�]��[7[eT�Z����f@�Ǔo�x���O�����#�e����SN\��,�+��:.Ha Q�K�n�&XS���mZ)'�qa�w�Y���=^8�m�� #�0	J��3qϢ����ԪU��!рT*%(\eȕ�o�@�z���X�.�y�
�6�����ah��)��3L�* �%�.X�`�۝ �Z�"~�挋61�V8XӢ�	�(c�aB̲p+Ê6'���P.�3�0=���Ł#��&�^�#�J��px��F�߃&�Z�Ag�3Y�P�UC	/p�� �K >[3�=SS[�<iсK*�����nS�E�:�(�[��7B�ZhR��d�B�j�O��}C�+ԍM����$��Us
�'-p�`��_LO���g��
o���$��e��m�t$-�?��
����	
V1���n�����m�/ro8C�I�I��kd��i�]�5˘'\r�d�޸@�T���_��}��I�!^iK2l
M�`)�q�GK�T��$N�t��-G�I�^�	���+�Ce�
��Dh�eB�#�(B�I�&G���R�"JJ��p jk�OH���ޡimyR$�=�H�0����6(�$5��l��� �"O�)$%�;�ԁ�R��,�hٺ���@P��I(*|������g�\P6�b�E�����{��_�F����/D�����IT�e䴙��Ù�t`�yE�ԕ)�%Hf)i:������@<.tb$T"83r��@)Χ�ў֜�C; hZT�#921�������e�4�W2qT�\a�"O�C�1 T
�˖7O���'m�0Q�@çe�|AQ�T�"~zc�Ӊ ���B�dُb�X�I����y!Z����Cc�ϰe&��T����D�<Ɏ����ѯ����Ă���m��׆�D#�eH�@��'�T;���#���`L63|8B���%E���*��^��EbCacX���f�D6d|h'�ϝF���05C��V�͂C鉜5*��4gO ]{V��|�SB�$Epl#")'g{�0��\�'q(R ��Q�'QوX*򈕸'J�֥�32���	� �H�+����h[2�����,� ub�_6�}{�������G�>����3_l�"}�G�?��yK �_��,���i�ny�mA�|�l��"��P�ax�ɂ�d猸��LLh��s �N,��'�� ˗ <�pvj��4a3y�`la��,�0*'��1�`��.&�Od�Ά6:�ͻT�S�	�V�)�	�/,�D�q��d�x��y��>���Z��P�5�<!���
�K�4!��?qsI4���l�rl��$�>�h2�� ��"O�,�Ŋw�B�#Bf���,�
�"O��P�Z���!�%/͞H6( �"O|��I���$W'.8|p�"O��pr�R�U.��E��h�l-��O�@��}�$���*���G
OV݌Cቺ@t���2���w��e ]B�@��ċ)q%��2�O�	n�?5���P�N�!YV�哥��]�D��
t���r�'�����1	��yz�l	z갢O�4�TnX��剞��S�D �u���^�?���,Z��t�1'��� �����C?D�ؠ��<�Su�nȔ�+��)l��	�f�Nظ2��Q�1��s��s�ĝi�mz>�˅��LzD��AY�Xͨa��;����ğ
#��HɦaBQ�LY�P�=��HB

�h.�u-Tg?�UD���ϻZ)�t���'��l�c	H�m���iwkŘo��a��D�<���|�)§�4���`�#N�X�p���O�=x��?��%��.l�h�C�%�	���/[�BL�ɍ7=�Lx�Q0S�n�h|��S�~���o�,k,��&�H;��V�^*>�SO�Kb!�$ʖI��l &
PE �j��e�I1P��4:`Hf�JH��J�K@26��Z?qV_>�$c.���[r-\�UPBAh>�O���PD�>E�h�ɒ�ˇq�j��E�U>F"jq���Ԕ/_�THǫ*^���r���O*x:@D��`)�X9��B9�*�cS�X(-@b �1X��A�G�sx��j�K�'j֊ �6�'�~�����e��y��)� P0�O
,Z��S�� to�ѣ�i$�U�@�ʹy^Q�O�O��SC-,v�B�Q�V4�Ǡߟ�Zq����yr�VE��"�#H�<�eCŉ���U�KzE���[+O�\�qkHJ�S��!�(a�~�%n��X�`x�o���>�f�_g�$�#u��u6���i[�y>l�H��B�I�T���B��(V�]�E�Z�!��#=Y���(Qєx�/��9�z�9Đ�W^��3'��X�C�	8/�Fd����z$���ʭ��7�ԉ_�ԯ�%��)�禥���u� ��f��:1�db�4D�:�\4���rHT�
��I��>�q�@�\M�`�/<O�#�C,4���7��D���G�'����\0cO�!@rN_�twFm)����]�0"O`���,��t��@u+އL�F���I^ݞ����qأvf07��I��w�<B�I(B�x��S�P�"B�}��f�Q�@B�x\^,&i��&��A�Q�x��B�	(B$�l�)��mS��T8���m�>��rh�|[Tx;5��;:�`�ȓ����C�e�.4�
:t���ȓ(����S9:�����)G����v��a����f^-�D��).2h��
�H-�RA�4�@��&@?�L���=�
���1P�.YA�n�M�����V�J!SK�Z�صc�q�J@�ȓ7/���L�U���u�����{��Y3d��+�r�`cO	5	i�ȓwc$��b���6����aK�~p�ȓy���� �Kzp��)M�Vd��<�xSK�"0
��V�B�/d��ȓQG.����;D�]�&h�܄�ȓh"J3�N4(�� �e�)�!#�'�PcDܕ6�i��� �4���p�'�B��3OXX䎉 eE7"~6E+�'k�l�B�0m|��mU,�Z�#
�'���07`E5X�Х�čtu>I
�'<&M�4텨�x��e��vr<�`	�'Y8%�c�O	\Ѫ��N�':pf�x	�'������5]��:�&]�34 ��'g4���䄌i�{F+` 
�'v4t�WE�L�҂�A�ƾ��	�'=��"�)��J|��(�����yj	�'c��jAb�a�]z��TT����'����e�>Nف�H�=lhţ�' ��j�JAR)f��*�����'N�T�"kML9�+h]����	�'��I� .�(���3�-Ā���z	�'��Y�ȓ�nQ���X�|�t�B�'��`�؞^A6���. }x5R�'�VM�PeǏ\Glm�#Z��YB�'���:�-�'� 2�J�Ķ���'Xf�a!�1涑SA*��Q~�)K�'tj�K�f˳m�^QJ�
L0�X�
�'A�A���s�"��w嗯R��2
�'RD$�	�&s��sT΁��H���'��!�e���I�A��(�����'�>9�a�X�H����bkˁ!�`!��'	��	��|:��s��m�̈p�'.usb��/�v����m:)��'���釮�+�fE�Q��h!�'�,@�� `R�|�e@��A�T�x�' J +�H� ,VJ(��BgBT��'�:�� ߧU���끋H	4��'�Ԕi@"�	B7(�S�gú1��Q�'�~��Mڇm~xu怹sc�E*��� �\�fdM�Ya�L;d��3J�L�'"O@Q����[�L)����Q"Z)0"O����[�~	>E����F<sE"OZ0�%���Kh\iZt|�"!�S"O`���0:g�Ч�A�"��R"O.�r�m�:g��zt�K1��,�!"Oڙ�W��;���)���	a�S"O��3c��Wl���$T�	�,�P�"O,�+�B��_�vY����*l�:�"O���#
�)M~|�`�
=\�%2"O���%nct)H��ߚ@�V){��'���B��_�	4
��a��֝J�ށq�B��|�C�	%9�JL�,��V �x�g���L�'�D,��oLw ɧ�O��A�-�FIP�Z.6hL���'q*�p#���R#�(���@�J�d�V&�R��D�5g��.
!GzuHc��b!��4d�65�e�V�.%Є�'"�y�P���/ҁZd��
�"�d���Jsm�m�F_�  � ���Q��.B�2��a(eS	�Z����Q>����q�xq��Ӱym@)��������'�МҩV�
%\%�O>���$?�$���w[��tJ3D���Q�+As~<tkW�E­���K;'�_��;���U�gܓZt����-�(M�@���$_#�B���Xr������=� �^9Z���!ZH�bA��j����BL�fzH �@� �y����..O\8�#��!�œL�����9pSJA��rqk,D����xh�� �^7Y���d�/}�=l��Q��|��d�Y�K��!: ��	 @4i�E��y�d8h,��G�h���iA�/MqO�<��@_W�g��� s�ٷ4�1`����dB�I�.�a��E�,�-�'��YwzB�ɒO�(�������Q�T�c<!�	B��ĉ��$$����/%�!�đ�`�"�*4h�X ��ڭM�!���$1�����Vm���ŋ !��-�<�rڌ%�J��!!@�R�!��؎V�R	UIMzu>���",��'t:���bMlX�xA���E���B�D�Tݙ��9�O�<�Ҏ �0�X9�˞��-���ŤN�rU+S�%��a��@������7fR����$���H�T�i��c>%��g��74��O� ݰPA"D�\��
#�FPQ�ɚCg1 �����T��/E�S�>E�4n�"]���ׄG�. i��[ �y��ع{J@�H��C�4�ʁHq�����Jn@�cQ���{�ax2aғ6�貤� .	��A"���p?Qw�\�O@�h0��6R�Vi��`�٘�!�$�P/C�I�� �vi��	H<ܠB�w�l�>iq!��k�>�Є#��JM�RjQ�1��#%��P*B�B�xiaL�5�R��o�
?����a����7�I�}q�S�O�Tx0�K�y����/a�����'���G߼v�I��'�C� 
I�� I��`0�'�\j�.Ҍ^��ãdE?�$��D,5l�b
�{��x�A0ǬȽ
�&8�
O:��� ζv� <2/CItyb�ɂ9��Y��	��<��Pwګl����ä��%qO��qr�]�0<�BE�(@�R�g�;�b� �+�D<�bł�hǌ���6s�!@����=蜠&L���?�BFѵ`��T�'V<}Jp�
��H�'ֆ-j"M�[��!�Q�?Uɢ�}>����[/Yql�Ң��վ)l����o�`͡ejgU� ���d$>7��󴉎?�y@�,��^�I&8�DD2�r,���s���f�0�U�P�<2���a(9U��q���Z�4��X��x�s%�9�O҅ d��<����F�־z�
�VÝ	A�n���K����h��@�5ϟP�hi�dk_�H�i��wκ �\3/��ӎALƶT�	��˴%xP�ƌ_
����(�]´�L��`ĘE��=p��Y�b��'H��z�G�Z ��3GϹ?i� �V]:�� J͸��(V�a�c���������2E_�h�F��X�Z��R��É�/ �
U�S��*�>`�s�>4��r�H$; D��"o�$?=��#c	�,�HO���Ǝ�>uLƅ����I�Nx*�^�89wF�6\2�B!�]�}���93�*�ђ	�N��ы%\�
�@M�c��u�8E/?h�x\���J;��K�wo����	� D2w�z�l�7���#x�DR�R#���g�׺6SL ��A�H8�s5��z<r��6)Q �����Xr~�p�gE&�jB��6(U
�'m\�7��$�V%Ŝu�t3!w�ލ:cJ�k_F�i���4Bx�1�-ݩ2��4��O��P�C��(��uO֤HF�@�����p<��I���փ���~��R	0u�M�@���P�M"� s�[5�t)q��V꼤���3r�QGzb ���(�Qc��zFr@b7���'GvPJg$��%��A�ݑ`"`�D�e�������`O$	Z����:�
؅�	�"��=QR���J̬��bY�w��h9�.<}�iD�E�:�"�ݹ$O�9�F���F(K��SѼ�`�]�O�z�{��Lz���H�<��)K�v< �$�����r@ 2<���+gCAN��ϓ(5G��O�Q�d���PLBsʊ|uX1�#O�h�1W3ctHA�ӌ&����� ��~I	S���$�PB�/LO��bS��7{z����B*)����'yr��$��(-�=�c��4�N��B�0#��Uj�
�B�	*"O�L�!�c&aK#i�7�B��#�|� 2�Z�SE�Iv<Fᓯ3��1�^�S�V�A�?9�B�I!S5`�[���*C^:���*]��)R��F� ������OF��E�:�3}��Y��(���RPJ�J@�G���x�A�*�LE�%M�7�|�A�`����OU�Z�xMC�
�5azRk�:�P��!BO�6�������<���BJ�"���I��c�B�î٬rMDDba��S������"�y�dB(j�6��I��eʩsń����e��K�dIK"��fJ#ҧ	�4��A�8d���Џ�`�&E��j���H!��vԈx��T�k���,��yR�Hͩ֫�@���?d�R���ݪS�ӓp�a~ҩI9B��5K݁%��A�� �͘��� B��H�/���0?�J޳e>��!�?M�0LXT�^�'y�����Yl|\Q���Pznb���@,4���ؕ`!�dW�@��tZ%�(ԘP���� ��ͦQ����⍈��)�'qt����2SX�0��*?n��1�'��(�&�ٖOC��0�l]"O��H*O:�C��s�$u�c)O�R0bD9����$J(+�,�7�'�&����/�����;a�,8Z3B՜md~LX�F��y!��ġ+�СZ��"������ў�
�K!r�\2��l�'0��eʥb9��zq�^3��(��6�<b�d���2�ˏ%E���I#dFnP-&�p)���<E��hVaN�K#�~i����l�!�C������ARe0U�]��IiUA�!� t8`���ɗU�h<�gօP:�t��F�1=r����
<�����	_	ȴ�̚�2Xn`B���4t���'��L�e�$j�1k�J+)�����I]dT�Q�&;��9?$��"6K��
�X,��J�C�I�_��$�W��	$f���+I�׀C�I�y�h)�D@��� 4��c�I�bC�	8 >BD�f��]������0JNRC�I�I&R,�g�ĭQ�	+�i��nC�ɕ<�z�Rp�E�8p�'��I�HC�I�N@��J�#�L rU�<v&�B�L�z�k[!vC^��j 
hbC��#�(1�r#N�?�<4�sa�/x�*�I�s����'�~p��=1�M3�>y�x-(�^b��{�����?��LK�,�����b�{B�c�<qG�\�O{^|i���a��P`f�D���4��n8B��"}�$�,��0���*u�`ph�O�<��
�胭J�t1BA�
��M���� �<���h���؜tP(d�@�5�l� �
B����
d�Q>%Z��]
H��(J�DQ�ߊ\0��Oڱ�t���rE!�ۓ0��xpԢQ.�1���uQ���J92��B_�)�3��1-��B�~�VA�G@��i��Y��=FQ�)W"O�T�� ��\��G�\^N�ӕY��$ҹ}8&��2��J� ���,}�Ť|� l��5�ڥV���dCt+��1�'�^xy�n/����ъM���7-ǰR�>���Q�����d�=�􉢾H���Y n��F�̂q�&�"���e��� �l�Z��s�) '
�4܊i��8�~5�Ί�7�r��k��Ļ#�s؞h���̔"Ҩ���!>!�8��t�6����۶s2�O���(1̀����DA&�� ��φ,p�=����5K�!�dP'
]05�����`J�>q��I3�M�HɁQ@����������,H*�y&l�!b)U�h�a}bd��A�8�(�Q5k� š�F��]��T�!".]�Ɠ} �£�=� e#�ʓ3cܖTDz���Lс�a^�'U^@�TF�����F�8�f���[2�-��ܿ)q��b��(+���nڹg[����%ϾUN�S��Md��"Y����'��u�b@:'��B�<1�&�7y��p�Z-h��!B�e}��P�d];�G�Hx�
F䒮=� )T��T<�9JF�*�O�1j
�bF,1�C��*4ph �dէp�����*D� zT�8��P�o�&-����n+�D��H	�4�'�:���"ZWn(��D�bў�ȓ`�AJ��C�VF��gL7u9t͇ȓA�"�bҘ�+u	2j5��ȓO�4m��Fū$6����4e��5��*?�
��D�<�[�I�ST=�����DC�DZ��T�\+:�����^���ǯ6��[1�Š_?�x��WbR`�`Kٶ%�ܩ����jP�ȓG�H�#T���>�������2��Єȓ���#�L���*u�d��ȓ1/$���l�}Cb(��W��H���M
��h��x���w#&S����-*@a���0iH�a�����c1��G�yJ�)�_�}{�f>t�`U�ȓ2~�HQ�ĩD���NUT�z��ȓ�j�SɁg�r$襎�'4�$H�ȓ�j�H��V .��u �4Q�ȓ#�ک�R�ۈ06@�����'�Y�ȓhx���G�ڶC ��LI�@�JH�ȓg���&� 
vp���%F��ȓR�Τ�"�e�D�	
*v�*������<XO\@H�J\5��Z/���.u��HԎ��t�v������&`P�1��5���»\_ `�ȓt��!cD�
f�B�y���2M�|�ȓ6�"��s�&>u��X�)��h"-��_V	�p�ޔ�珎�`v�ȓ{��xsJW%BH�HuBr��M��\�� �4�ɏ���#�C\!J�$��%q��YMx
i�d�ZX�Jهȓ+	���&��mf��ϝ�Ln@͆�� �5Ҡ���K�s�N�ȓm��DYua�$�T����#���G|B-�/�0�crd���-�DT�y���hOk��&,��%@�lC�I0y��i�KU$�,Y�hȤ!q�C�I<p���P#n"�b��ڒ*6�C�	�0��[@�����R�X�^�C�	���6oZ��x�r��<!W�C�	�{�h���$��6�Hݱ3C�C�I9u�[f_9��������0��6jf���\�c$�A��A��DYz=�'��+)O��z��i�=H�Q�e_��*U;&M Mk"�xƣԛ[�1�Q�i�&��IĦ���B;��@t �/Z��U��m].���I@�D ��Ek���С�+�"%�C���6AV�j�	�*b�����8
-`D�즥ZU��x���i�u�8 �!K<\e��7ʊ*9d�Q��æa����#�D]Y� �?=D��¸("D�CJW0.����4��6`�2bԼ1�v�,[)J��h�'����%`��B�T�2D�?( �h�k���"4h�CUh��m�p#}b�π \	HǤڛ%V��Ĕ�O�8Є�� tM��Q�A�JN��D�˃M9a�4ϐ5\�q�-��P�l}��߹�Y�Х�����'���31���?�Z��!����)(�6���°�� �̀�JE9�a,?E�d�ԝ_�����B�A�(-�1oN�HJ��5��()*���"~"]wĜY �oL�2�.x9��]I��Q�م��b����ē����0�0�I�U1Ad���n133b���U쌌�0|Rd�\&dJ�S1�P���-6-F	�O���M�
۸��O >�y@nZ�LX�I�OD }G����'�Q�ѤEd�1O�>E: 	�) ��BM�O��Ղg�&%�s %�)��5��7/�����$ �ܠIP1D���7N�z*f1�B��j.��8�&:D�xKw���MQQz��DBلT� �:D�X�r��?u�t�L�AI��7D��RpE�05���K��P�h�i1b(D����
ڜz�nغDB-Z22n&D�(�4��/��؉aOɛQ�PI�/D��b�gH�$�yaG�)D�:ŀ�0D��Q�̔/�X��d�9�l0Bҧ-D�(�蔁]�N�Ypǌ$0@�l	E� D� ��Jъz;~5�&G��=��*�=D�4 �G�/�<�1&ŔW(�y�b�;D�d贄&+���B���7*<�p��9D�l�Ī3D��5��I�]9.P��A9D�Z�-�1h��9A��n��j�,D�|H���-y��)tǐ
Y�x�*eJ(D�\��iK�t7|PyV��:Q��k1D�T�q�J7X�����Z9cCHu��+.D���o¸U��0@Ģՠji��2D���lP�o��h2R��L_
M �"$D�0����y���k���P��tRgN"D�d(d��!Z�Y�q@X&/��1W�>D�D�Bʋ&:�=����\z���U�=D�0S�'@�N� CFh�?5���*8D�<{�h�jZR��)7��]���3D�t��I�R�f�G*6�ݹ�M.D��sc���~�`�Y� �ziC�E,D���2)@'��	+�	�8$~6d+�6D��	0�͸?.����/�:]Z@�#��4D�@j4�Ǩiq�1��!�-�&X�I?D�P�u�3pv�Ӱ����e�0D�8�R�L�&���1J�i��2D�T���M�y����L4T��8gO<D��r �Ê=2(��k�v�֬K�j:D� ����4d92̻WD��/q�\�V�8D�����G�~�h���+��U�h7D���½2S�|Xf"�LA�ecel7D��[bnI�+'��h���,Z�؋6�3D���o	n"�ĺ7-�-cn�K��$D�@X�*�a�c��U�^��$D�p���O�h����u��}7B"D�d�K� Zrc�K��A�|��%!D� Ӥ��?��C��"Tܰⵁ?D��hc�Z+S,����)3����J>D�d��'[�4��A�&�(�^hy�J;D�4c��%���G �6[\ E�5�4D��Sҏ�
G�bĒB��7>��I+3D�(�C��ZD�����܅1֌�I��&D�  �̐l�L���Y�)<tӨ0D��
0iH�lPSGI�4*�h�m-D����HN;-jDd* �*.�i�Q@-D�416���R�b9c�T�o\4���,D�@i��(@@̺�m�(o�.�ѣ,D�Xt.A�S�P��T�5n[:]I�-D�4c�S�ۤ�;t'�Alx��4(-D�� ��U�s�R�P��S=<�±"O~D0���Y�@=SӨ�F	�,Q"O��&��?~�ApÇe�0m�"O�!7��?����N?M�H�"O��)�^4)���Պ��zD�dz"O<���-߹i���*�G�`12E��"Ox�S(b�D��FI+�l�f"O0ٹ7,��6�tI���'Ă19�"O����۠q��i�j��P�~|�"O&!C��E�<��x��4{Mz��u"O��A&'�>G�tX{�m
&�ԳS"OF܃�&S�}Q-T�@,X�"O�y�E\�B�)e�օd`^���"O���w�\�;]:�h�P6�X�"O�I	6S�
9Ria���":�[g"O�<;�'~И�(͕��:�"O�0�,�>y~|�0E�'�h�"O
 ���S3�8e_-��8�"O� #�ٿqYv�Zs�2+���{�"O��#�f�s�����W�`ʙ�"O���Wh^�K�8�8��0@Z�]V"Of��જ5A�.d��
ݻ2A4���"Ot����DP���I�?C�B���"Or�J��Ё��mr�i�KO|5��"O�AS�@�4$~��!i�<���Q�"O���2�F��$(*�(� �Zԩ�"O����M�J)\e��.[h�X�S�"Ot��eJK���Ed�>E�@@��"OJ�2�Ӻz������imZ ��"O0���̤B�i0�h�7Yh:�"O���u �$so�ar�C+'OV] �"OJ@�ā�3� ��Q�UM���"ObL@t��"/���i#o�/d6!@v"OB0���@�iT1Ĉ�l�0�3�"O�$R��q,:5*�IH�d���"O  �1IZ�a�9�E�ʌA�F���"O$��Ҥ/�N���,�#3����"O����"A��8C�,@):DHȉR"O��ґH���l5���G	=:�A҇"O�� "��m<i$C�'J1zD"O��1��ƾ��}�C��=KlT���"O��3gDQ4a�P�Pc��N[��1"O��x�/	�BB�I1MQ�RLdQ+F"Or�2�M	B�h��K���@�:u"O>Lx@�H]��`�K."8�!h "O��80�N+_��y�ȞL�H�xf"O��8���)
�`W'_)mʶ�"O���"�͗�,���'�HɲU��"O��K'j��\FPyA'��Ag"��R"OB���*/��y`���rQZذ!"O���mR�*8<���.7J�HA"O����Z�e�R!����>e��a2"O��+1��;W�PP1�i��]/��4"O �j��rJ�
�nŇG#6�g"O��R��ڔyLT92-ً��HR"O��C� @:U7���ʊВ�2�y�H�+���Ip��'N
B��y�L�C0 ��%��7���XW��,�yb�^�l�����Fq�/>ڭ��>���8��Y�b���y� �Y�̐�ȓ�`�pE�+��)0G�4d�>1��Z$��{��Mj6p���7X(l��ȓdg���.ԗz����
vQ�ȓH�T�#�T)I����B�jV���S�? ���T�OMa 901�D`����4"O<�IC��:�"�*K�8�r��"O�\BP
��2
P�ЌlY����"O�8�7�):�:��?w� ��"O�qK7�P5�La�`�ƻh����"O "A�)B�r���L؜VBY��"O�`�!e��p}��Z�/Ut�P4"Ol�:ծ��H�������U;�@SC"O���`d�7���he惉+W.\`T"O��¶�P< �h�TeE�-D����"O��(3 ӵ%=@�c���E�ظ��"O^ � ��-�I�kXc�
���"O&`�$� =����[(�����"Oؒca͉�܈�FD�YN`(�"O��1ڑ3�zĘv�ϘmS�`��"O���R�F2\P�z+�5J���D"O�QC���|�F����G,��)�"Of,������n��_&�(�s"O�9��8'��d�ÂF�7w���"Oz��U�1�tف� �nv�pr"O6p8 �F.�6(�u�����3�"Ot@`P��&� �����6��g"O�$��S.
}0��؈`���b"O�=+�m�]z2�!���.��4Jw"O�Y�*�.P��Y "kJ�g����r"O$�Q3M�--�hQ�$*_���t�%"O05��'^�.}��h���� !"OjA��)ݑ^b�ɂ&�\�[g���U"Ol�x ��<�L ���V3*U�6"O��"q��7�~Q���ςL�r"Oby2S��*<���qf:+	FE�2"O�����b�2�A�θ�I�e"O\U#��� ��<��$/i��ˢ"O� ��E�W��ɺ�b^6��9�s"O0��eT&up:�1�bλ����3"O�m��Aӛ!Wmj����zԆ,��"O4\���ͼ:�Hhb�/�4�b�"OR�"H%R"��u!S��0'"Oy����CQ�|b��"[��Z4"O�=��L��w4D���$�B�"O��6�@��e`7�a�T�"Oĩ�,�5f�������"�d�(3"OF����*E�<�R �Q�i���1"O��ˆ�۳_�R�y[Ȕ�B,Σ*�!���
hء9f��%�՚1���s,!�d^4R�2S!��X)��*�u+!��2r�H�Qt���w^����=�!��V�Vv��J����2g���*Ō<�!�N7����h�@8���ΐ�!�D_�%<�̡u&���C�ޕ!�!�ȸN��|�WK�<FiX(��-�s!�ě �p���� Y�Xb�"��u!�D�4C�(��E�l04e;����tE!�^1A@��#�N�v*F=�!�ǹ9N!�$ҲU�Z�ss+ɋ) x�K�F"K!�W 3R��$�� l�*^��!�dxkz�+���.C@)i�aWN�!�dQ	Z8��R�F5�p���Ϥ!�;h�d���g(��K0���!�d� 2�����ļ,hukb�P3_~!�9*Y��ڑ�M�f�|2l��oj!��<��@;&���p�%�!8!��C��mT15�d��$U�u�HB�YQ ����P3izl����DB�)� Z�!O��¥#�<�0\X0"O��V�"㣁'��8ɦ"Oj|�#�ߍT{ � t��L�t"O�t ���*S?r��sJ�(bӎ��"O���d�[¬�[@�>����7"O���̼|gdؤD�X�>�"O�1��b�4*!"-F�!&�l؊"O��3�g?��x'ϒ�I6�lB�"OTU2jٕU�h�W�@e�����"O��`H�5M��a�#�*U���2"O&�q�EI<rY��)eˑb�6"O�Ya��Q8�$1��^�ԅ"O�U3�$��(������.�ą8�"O�ڕ���&�CP�<@�t͒�"OƱIp!��B�p�)3��"g���c"O�d�� 
  �6��1�R��B�	/)l�yG�:K�����@9�H����e��O�V��Y#�
��X�8��3/͇M!��.l�2р�@����a�0!�䑏m�$X�pi�*K��j�ڠi!�DL�A�����L�Q�Dd�F�   !�$�Yx.��g	�r5�
�mY�qD!�Ď�"��pL|���Ҳ�B+9ўK�D;�'L|\�5Z�""�1r��\�\�ȓƚ�3A�0XC6a���
6�~��!@b�Ĩw��a�`�oB"1��*ڴ��B�9�R���ɪh���ȓz�8�3�@�Lhֱ�fF�%o<���ȓ,�\]W@DI_B ۢWE���	*��#<E�t働�l)h��@=���銺f!�D��	U0��F���X�燞>T!��'|�l� @KP<%��`�a�E�*^!�$�?HT��̐!�����d۽6N!��$͚8��@J� �p�^�>!�D�7��"��7� �� �則 ���d��#{�`���Z�9�`�Cu!�66 !�� �a(�D�t�(��d��8[��0�"OFQQ2��%��3t��;��"Oy���
�� �A�A�Z���"O�@�@��,��=����B�h-���'q��h�'Cl�A��Q����&'Γ>�,<��'0h�@��L�Dz�ܫU��64�`3�'���Ў��u�h���і;1LS�'$��Dl��� $gC>�d�
�'�B)��*FRp����7L�l[
�'a���K��s�"��@��NƊe���ę'�Q?-�v!� s*�����Ȩ���!D���T(���ّ"�Z�
l���<D����I�����0����t�:D����#�	U|����K�l(�&�4D��6��$ȸ�:4���`DN ��	-D�ȢKM�X<8"���2>|���O*�r2�)�'5���7NIm�t8�D��V��s�'�6�R�M
?�*$X�$����'B0��O�f��q�΢4x��'wZ0��F<K����)H*�|�(�'���B�g���sC�߶�
�'�(�:A�7t��!�cC�Be��(O.�Pp�'n�ʥn�8H�v�b��3P�-��'�$�S$����BA��F����'�
�KCFT�
����1+RU��'t��X���<]4���aS.(�@Q)�'#�c�,V:�t1��N�$69�	�[������0��2-�lO��N��T���ȓtɼU�w��<&��<�BB�?�Nt��g��d�т������f�bNJ�ȓh�Dw�	@;�|ÑIU>~6v��ȓy��8�dK@օ��HP1fH���ȓe����Ʒ8��P6܌E{�F;¨�8)@���Iu��V�^.C`�Q�D"O�hE&ۯ`p�h�	�)c�i�"Ox�!E]�z���T�М+N���"O�����.J(֐�Έ6t=��i�"OI��Y.-JN��f�&<�y�"O� ��J̻77��#/\ -�.0�F�'U:A����*2��|�cEƲs��=��G>a��a��BغAҍיI�x2:d�8���?ስ�ոn~깹f�X�x!�ȓ6i�$ÙH�16�O/L@>���=�jM��."R��V��,T�$�ȓHbL9�!k\�Bn�����(7�Z%�'F��B
�	 ��a(�0L���w�L
;}VЅȓ���H�}ض,&B�8����oǏ WN4qf)D�Y�؄ȓ91�����[�h+��x��)˰���,M��Z�Li�5���P�bd����i��I�{G~��b�;It Ȣ�LV>ĘC�	�<{��i)s$�@ o��B^rC�ɀ]���K U!T�%�Ce(�6C䉱k���%�<k �=����)��B�	>+
vX6�+���j6��W�B��f����ކ+E�q׌#|\�=�F)]f�O����旬[Bv��CPϦ�q�'\��ݾP^���в9����'����h�,H���"&V�;�( ��'-��Z*c�|9 H�&b�LmH�'��1�AY�T��ؚr�G�.c�d�'��(qɗ�.[ �1iW�-����mh��Dx���Ą>���Xd�
�M�L�0
D< C�+?��5k �@�d�*rfǊm�C�)� �=��)F�0����Ѕˀ"O�!��	���!IA�&�d��"O,- �M�>�b@Q�!�Kڦ@;6"O�i"�E<J ��҃�V�cb��dX�|���0�Oj@i$���)� ��W[��("O`Y1���}h�i�dJ�6)2!"Ody��O:U	<e��$(0����"O�=�&��za1P�F2���"Oν�G��M�W"��U6��1�'��\�'�fm�'(�-:�ThS@�ك_���'��m�pJ�2%0��(x��iC�'��I�Q+M/Kt��WA�^n���'N�qB�l�
4BdY��kR5O�h1�'y�!�Q��!�x(W4?"�=h�'4�9ae=��Ȣ4�	-b�������29�Q?�IPf� r!j��$�y>�U[0c"D�(�2�W3���A��l�H�Q��5D�Lb�&1��y�����%�B9j�!�R
U�~q9C/Y��>	��cu!�жC*pҫ�V�,x��&�!�d΂(�0A�u��;g ~u �ʇ7��̋�O?��&�B�N�Rq��,V+cpD-�"�K�<��FX�_K�2���$�Z���D�l�< �L�D<b�0�'Юu��j�<�gB��F��Q����j���QF�P�<)b�{sL5�2
��8<��	P�W�<9��
# �p�5g�
n����Wy2�#�p>!��Wjj0���t� ��DDT�<�u���R�]�G��[Е�h�P�<��ʻvj	��J$.lhE-~C��0����K��8�˖H�M�B�ɩgX��"S~��s�G2FB�����9��3NP�(�L��]r���%",D!�D]�:X�(ր\�ii�ejaҟ>!�S�|S��"��7x�|!��NQ�_!򄐈S�Lт�D�5}.%H��"9M!���!��!V��ic�ő!m�32!��x2���ԩO/\b�kjէsў�; �!�'`��:ޡ�"ϣp#���Z�m�b�T�`���J�o����'��@&�QHX��cfݞTꠇȓY=������{���ѡ� Gi���ȓ=��w�ե%%F�v���@PΙ��z��&�Y0+-�A���<�B����}f"<E��j^�#X3��?R|�����]$RA!�"k��!�q�ʴKu��)S�b(!�9e��QNQJ��t�%��!�ѭSp�\��%�<z�Ԁ#��N�!��W�p,�6B�mj6���G�!��ʼ@�:�x��_	g��`��ޮR�I� چ�����M/��P!G�6�|�+����02!�ݟn1���7$Ϯ�ˠg��!�$� r��ђš{���p@G)K�!�$�(]��l�/7|�	���E�!�dGZA����Bip�n	�5��}��4�~�mZ}�܉�̓4���b�B_8�y��O�IµI#F^�w�>�����y¦�G�ܕ���8r$�H�,�y�D�7�B�c�I�p6�8�h���y2)M�d{\����@9�N�h�n��y��=L��� q̲.C�9CgΗ�hO<�I���$ʒu�s �9Y�q��L;>�NB�It
1����`�
��#�ShB��9�^�C�
�,Ij�hޔ�@C�)� �,�����J�k���=4�p��D"O�
V'��0�D<s�+�{��i�"On);FI���dY@@��� ٣��'k��0���%���C�MZ�5��]2�`�2����ȓm0�]a!�*v6���k���$���1G�W1Z���Y��<z38=��i㘨�����H�hV�J�x��ȓ
�fxsfP� .��@�e�N����*A�T�F��N�,����j�.9�'�ĄI�tV�A���M�xJnx��oL ��!��a�j�p� )�܃%��*�ц�b���0tCӝ?����4,��`��#ոI��O���kt�ߦ-�J�ȓF��	�4��>0��;�` IM�a��ɸ6�@��8 Ū�R�m�.R��b�	��NI�B�I'�2��"���*6B�	�8���H�������Yq��/,kB�I4wi�e%"��
BA�;#	�C�ɘK�=�mӖM�1�Tǐ+E�C䉡<Ƃ���D�
�P1��N�3�B�=��PN�ODY;b/
<d��l�@�/9B�'Z���n�LZ`u���I�r�	�'�j�������w�>�bp��'ӈ��r@�L��� Oĥ6�
�'$I8��QRT�97��2C�qJ�'�$�k$�֝y���M�0B�R ��9-� Fx���ѕ8v�A�lB>�9��(�s��B�	=eS>ʡ�?��#%��'��B�əV$	��[<'��i�u���]��B�	�q#t�&F�fN�`:$�DB�<D�����\�1��"p��>~��C��;5x��I�f[{�� ӥ�;�l��[��+}r�ϥBK��+}�&Q�U�������|ı�i X��ǟT�	��0˦l�U@x�	�+�A@VI���|b؄A^�]���";@�I�b�1؈O�8r�.F����D3���'f�H9P�DGf���2&�(�8TF|���?��ϘO��	R��*:�.=���XZ^��/O�������h� �5��#�L�O��}�%�<�g���;�l�B�+�=�����Xy��Ǣ4�r�'{�k�t�'z��C&s�r���7'�[�@X�	B)M�b3��rèƸkF��r�O?����Rq?vP[cM�0_� �Db��h�Dʮ�z��-M�g �\F�4�w�T��㡈�tD����y2)��?i�������\�$���cנ}��G���< d�.D�̩�	�4[�{D�GJ��Q��.�E��?��U�T"��uh�a�ѹ��O��'2,80T�z��$�O��d�<��l�]Ҡh�/|{]` ��rߒ���W��?Y��0x%�/�A���dB�5l:t�7��,7�lrֆN�� @�O�EQ���=w$q���?#<�D�F�%���疈�Ġ���]t~b�ϭ�?���?��2>�����3D � 7���F�tIK�"O*5�Rk�>E�*���N�q� �.���$��|�����$�Rf�X���N���z��;>��M���؇y�X�d�O����O����O���u>����2˦��ׂL?��8�aZbs��ف�X�ne ���ئ�B����|�*�&����0�∮w�B칇m�?�|����7F@6m�=�z����	q��zJ<!��	џ<���¦��=�Uڌh�ބj�֟�F{��I+���u���D	Fb�Z�B�	�kY�K�g\����Uo� ?�����'#�	/9h���*�$s>鰱�Ӿ4$q�ƈ��Jp����ON}�D��O(���Ǫ������G,��'{V�lZ����ύ ~�Y�$�F�Q�`��T�'��$�����Ԥӎ�:]~��S�	R��Έ2|�16n�<�܍��n[�%)�AM�	7#Kr�d�O�c>�I� Jт́�	�3����'�<
�G�.p��
��n���\�LXXh������D6prly"�#�P�����5�ɽ@d���	 (����Y���$:o���'By��[�T5bT�SOt>HF�'q9٦�ۊQ���Q���tD��!�~"��d'\��^�a��A�H��Б���'�y��Y�TƤ�ת
���B�aR;��@7�乪��B��i�u  �C�J��R�fl���*T=��;�2�'��)���Ot�)� `��6�Ɲ:�N%���?cz�MC�"O8<�XnFm	eW3g���7�	��ȟ�M���� w�R�r�Ã�DM&)[�+g�����O������I����O��D�O*��;�?qB�� 5�=�d��e�0HPM�
9��@3�#}�.!E3�$������T�d3ZQà���e�>A�6�T=`H�PgY+�f@��MS�H�Ju��S���i�����X����1���Z�,[6j�Ĉ F�g���7m�.���O���?�I�|rf-���^Y�sf�:C
��K�T�<YB�d�!�(wO�DT*]I��D�r�����'81O
LaW��p��q[�oE0���J�'z&���1���0r�� :xɂl.tI����`J\�@�F6P�F��T�[��*O� B�I�gB��c\-W80��'��i��N�P	��dF
��M�ȓ(��G��'���G�O�H8�Fb��r��*@+r:��\#�#�En�x���<WtX� �'HRt�'.B�'�Pв�&�?Uy��� �:9"2�h����FH�e�u�ΎX���V4��O�Q�0��<ТUyc�I+��z݁3��ϝOZ~���.�)Fp��QAS�7&PЧ%�W��'hL���?y�����)b�OR#;e�������$�O���$��~@�T�K� g��Q�G#ln�}��<i$�
.{j�����T�z���Ry�'=b�'Q���w掘3��D�1��E�6ɒ����y�'*��à��'z�6��dg�&N�����ɗ����O�0����#1ܬ�Ӫ��?r�@��ba�N�D�5�X牑h9����On���O�����t���(F���eN^�E�܅X���ꦥ���������<��Wnz�!�ʟk,ݦ*
��:g M'/?�<S�@K��m��?�򃏧�y��8�d�O��)�O��I6��%#�ϖ�g�&�x���'Y$�IK�O��ąA��db�,�/�?7��h��O�hZr,Q.D��d� &�#EC����'�=�	��4RD����	�OZ�������w���%
�W��L(� wT<��		_����Ozp0���O�I,S� �s���º+e��5W".����^*ft�U��d�U̓8V����dA��%���?!�'�N9��D!Q��բ�ˆ�0���@��y�n��?A����N�OF�I/j��s�`1C�n�&=�n�t�J�M�`����A	2�b`n��<e����M���i38�i̟��	�`�O��#�B��Wc^�yT,�r�����B��	�<Yׯ
ş��I�?����<���|R�Mڐ,=TuK�A�D���)��A��M��EF��?*O��d�O1���$_9@�E�
4=�;����BC�I��IJ��0���WgN�M듎?�/O�$&>��	]��Y� ��q��L%Q*��i#N�#=���T?�U-҃+#�5���Es��퀣k.D� �G�W	X�2�*7BN�5�i,D� ��
�~{����g�V�t���*D�l{��-�n �F�\:hx�'D�ȡ�ƀ�@{��Ce�F	:� ����2D����{�p,��ŔV��褩/D����G�Z�T9�(C�ah�u`8D�� A@�)R}���(N��i*A7D�\��ꍆP�YP� SY�؁�l4D�$ɅcO�G�̊�QVT�*�'3D���ū��w:z�c ��C<,�Zvd.D�@���Y�.:e��R�GD.Y�B�I9����0��K$���3@s�b�i�l�:�:���?X�@l��Պ�.�A�/ $*l�, ��҂~���1���i��H�d�:� ]��i:�������4n�A �ߘJ�6!�e��U� ���b��%��4#�^�IT�Y,����X�C$�9�bj֙N!b� !U�ELd��'哭��m ���oB����wӼ Q��Ξq�J�{��I�HʤHj��Kӟl�I>.�@�+�. 9Qtҧ�i�~b���iQfa�K�7�N�RD�T�ɂR ,Ms�m�;��?��� 5q8@�4 ����'�Ni ��'���'��4��¦��W��T�@���D@C���O���ǥu� 	���.�LMcd��~�x��/�a���ć�x�[1DG�ZwZ��'}��'�~1ӢJ��2��<�F�r��K�'�^�I ă.�ع+#��r�њ�'и1�pʜ�m��̺r �):=��'��5
`*�5�<���, C�!��'��&��*N�P�񭇁%BL���'����RA �F���]�$���1�'�f)���T�(��{pcӯ"td1��� �в��1RF�<Xo݁<��b"O�D;͕� $�5�d��m�`,Rg"O��'ޑLf�U"��K�`�p���"O���i�9�8[���BQ�l��"Or��F�(~�Q�Z�%7z=0"O�b䃘Bg��S�)
�H��M�"Ov]�!�U�9���s���Zt"O�i�/M!�F4�e��y�	�1"Ox	�Eo�F`Ւ�̒7hj��C"O.
0"�GDM�`%Fmp�z�"O�1�7�X�h��<��Y1b����"OF�v��+:0���#C�2�v�b�"OHaD��+�D�GIY@��!�5"Ox R�H!�Z�����5� 5[E"O��Z0CP;1ڢ�+�e
�k+�"O�<�`��o�4H���ޏp�
)bc"O��;4��X�6��d	3G}�䘡"OX(
��/�8A�(	�����"O�8����$) Ai�(E*�"9P�"O$M��*U�X\�B� �j��3"O�9� �O�!Ybܽ2�] �"O�50$	ʈwψp �@F�+ @� T"Ol����5G���o�P\�B"Oy!�/��Y�l��gϏe���ɒ"O��1���&51� 0��x��"O�l����-0�t<K"%A<F��eJ"O�a�u�F�/�!�$،)}�,R@"O��K��	�5-�H��"O���a�ߵ{�P���D��"O���Ҡ��e9t速J�e��"O�0�+މ��	q��6x ��Hq"O�`���'Sܚa����A����s"O.��W�����
���4����5"O��!&�&!'x��W���M}��s�"OtUБh��y��PX�aHs{`�x#"O����o����醔k��5��"Ob�B�dA	M��aH�Ѩ���"�"O��A�B�>nq���r��Y&"O0�s��+UA����7P���0g"ObqഉED�"�H���|�Z\u"O�`kA���Q�)��(�R�De��"Ov�)
q��5S�'܉(Ξ��"O$�����!�fTɒHZ�T��"O��	��ױ!������4x�j#"OREhԮB�tT�"#�X�f��Jg"O\�˷ ��.iV��CH*t��+r"OU*gƜ4�R��bg�t(h)�"O,,yB!܈b?����
����+\w�<9������GF�ub6����G�<Y����:���PĊݪo�I����F�<���E�OT��㡕(P<�SQ�\[�<1'�֑�)�B����r�XW�<�� Ed%j��ݡ,�:�d�K�<���-3�@"�JtR!�aH�K�<��K�m�8e���yŴt!C�KG�<ѳ�.-h�#��?W��!i���A�<�"ޗtu�|9�Ĝ g�hy�v�r�<a� #��M�"�P�0�� y0��y�<9p!�
 �a�w�у/v��Ppa�o�<�A�U�{��b�kO@��)2�Fu�<��I�W ��`���"	.�#���p�<Y�队iV)�BM��
��k�<!`��n���v�`>|Z�K�h�<Y"iD!OW2DB3^@���Y&iQo�<� ��Tďr8r� ��5��9��"O�9rb�R-�>�y�D�Xtʔ��"OҍU��)������Ϛ K���"OX!�KZ�|���C�";�Q�V"OnX��%�!x�z`"i�!�t"O�0���� |^u1�
�,��2�"Oz��R"����W%0XRuh��|�<�c��-c$0	����|�0s�Ua�<�1 �1	�P��q��7�(h�Gh�<iW�Q~���j�@�E��[B��`�<	���+0�JMD���1�|UpU-�_�<)�%P1F-R��Rx�A ��^�<	V�G�޲p�Mũq8d''QA�<!����R:�\�2���N�:tҠz�<av[�W"��wb"r՚�:�r�<���XF�ʩ{%'��j.��qv�p�<Ѥ)T0d��E+#�B<�����@�k�<a A%B��`�V ��F� 쀥��o�<q�I��ESB5Q�-ܪ��0��B�<Y��[-Ұ  %�]�G,j�
F�g�<�b�')�};j� =L*�Y�Ta�<��c�4y�Ƥ�����u�<��;9��\�g�?���	Q|�<a��z�V��tNC=D�]���z�</��#m ����z!��z�<��h� ?$�����6 9�p��j�A�<	���(�Z�"fS�2�T!ba��c�<q3釐E��I�/��DU��i�A�W�<i�Z��u6�3����!�$$��=��#Ȗ.ڈ���!��<?�b,���4��ݢ�+G&4�!�$��A��U�B;C�	3�h�!��W$	v<`�D��QV�W��#�!�$[5XߴXd��'$�6Iȉ܎C�	�A��x���W�^04�bKȌGoB�	��J���K-R*0��+D#B�ɸ[���A���XقƉY�C䉆q�.-Y�咗���s���2��C��c�40�u�X�Uu���̞���C��/Y!����k�.�hK�
;�B��  Кa�P?#�X��1ă,,dhB�`��i��j����ŐRn,B�7�|(�e��.�><��+�0Q*B�I�c>��8A���>価����	FwB�ɇ	�����ʔ(J�g⁊m}B䉴M2�My���uy,|zUE��DB�Y�\h��E���d"5iH�n��B��g� �Ae_�޾�Pw�Ġqn�B�	�	�2�ba,�	����G�/T�B�U<\pF��ln8Q�	&�lB�ɒ~�Ir��ҝ16�2�kR8#`PB�I=NS� 0�ʼG@�����n��B䉾a��됬K�,�����(m;�B䉾J�T�z���/?��;�g��fB�	�fJ����������Jh��"�4B�Ib�����G�'Y�t���W.H��B�ɇ>l�+��)����fԦ%	C��/d�]P��h"�=�LR�$��B�I�,5�� �-X���7�T�C��8AS.����	i�V���ũ4J�B�I���%*�BE�^6.� V�D�nW~B�I����1+T�f��V�C�(�LB��:Co�c�ǧa�qС��\��C�	�!�4)T�ߪ8>�M��Ǟ)shxC�)� �+�hF�u%���a��'pF�`�R"O,��am�}�z��TÁ�o'�41"O��G��7QP�R�M&'�tڣ"O>�����* e>�B%��x.��7"O���@�^QE�Q@��fp�! �"O�p�F���1��׃4Ɏ)�"O�x�Cřt���BG:v%���7"O�5�SM�����;2a�J��s`"Op(����Y��A:�����(�"Ofu�0*ܿN�Di��Y8	@E:�"O�0(F�$��Dۛ},h�"O*�!�X�8,քJQ�;L��Q4"ON���:$Up�c���~�P�"O�`��w�vD�MDv����"O�X�׬�7��l�c��)shx�2"ON�Th��:��	��LҬ��E"O����\�K?P�AT��
�t��`"O��`e
d1"򂈝40�F�*E"O�Q1��)��̲�!{�L0&"Of�z!��;gx���E�Du؍�"O����]o�& vHǽA��Գ"O���@%�)r���z��� �
Db�"O~qg�_9��@�ɓ1"y�H��"O���c�T��Rt)Ӝuո)Xw"O���/|��!f��)��`�W"O`��?12{�%��%�S"O��i�.E$��H{�����f�_^�<����R:L���±$V��K�h�Y�<i���t�<�F�
�]�4;� �[�<y�݋"���y��!Y�yA��DZ�<!��47�F���u/v�#�O�<Y��17��0W�\�5[vѠ�M�<Q�- \`$X����S� 8���c�<��A
,U����d�P�����N^�<�G��/x�
��t�0U&��d�X�<�S%-qt�!������aw�G_�<9TA���A��O(�����^�<��#�HZ�+c���-�X]��FCa�<�4�1=�̉�)��N~Н8��F�<1U�]�&��`��hQ 	��D�<�kATw"8B�c��^����z�<9D"�&'F�t�ug�:����ы�{�<A0B�-"����
��#�)��#�x�<)@iӹ&>.5hv摡1�6D�4��t�<����()$���)j���6cֈ�!�$t����'�W:����*a!��D,,>�)rDG	)�H�H���!�����
1D�' |h�i�睭#�!���܋� �`W��#u�!�d��6~X�
�t�� ���^�t�!��h�&� �
�"Ӭ��ƮA:+�!�$��;H�R��>d�bH�uB��!�RV�6ћQ��(ْ�X!D��!�J&��!���K� �������#�!�dq�	k"�K����{֯��v<!���"��9���&�����P�N!�	J's7�ȿ3�.��4�,`!���^1��s$���HV�0R�-^��!�I3JD�׌DU�I)�m�a�!�/JRPu��D?��KqkK�!�$ %o"�y� ��-�P)zs�#@�!�"�șL�&�*@cڤ&!���e��`B��"~Vt� h VF�lQT& Ĉ(��cM�/����$G����U�D�`�=B�L�>0�!�� �Ѱ��D�E,�����6�`�f"O& t~
�R�F��F�4 �R"O���������RRFD��%j1"Ov,�
�2R�xä�|ńC�"O&��1��q�V�(c-U=Z1J�S"O�%��N��Y�&L�X"F@g"O(U��*ȬSĒ#.B�lLaa"O��ۣ�NMcf�AЍ
�iWrk%"O�AA��0,�(1���WH�Ł@"O��fgZ����sq���:
��"OƽT���BSΑb7��#�A�S"O��9#o�22x�Ã��~��'"Oεc���6<�lf��.$m�X.x!�Gv-"٧�4�*�E�Y,!��)�`22�˼X�d�#
Oy!�DK�6�0˲b��:���c�T01l!�D�"h����(��ƈD�T_!��*�<��wƀ/p��q��OJw!�$��\��"㈀�;�,�!'m!�c�x�0�M�L��C"�� Z�!�Ѱ$2�y0�,���ؗ���!�΍OS�u#C	��UÚ��AC�n�!�d�3� 9�/�9)+n8@��|!���fz�d��Aˮ~�4sd��
|!��K�~y	�%I�T�֫z]!�$F X��9!�F��?;���Kۀ"�!�q6�8w��{'��cǊ�"�!��J�fH���SN4F�V��� �!���,�h4�K�;a�<�#g��!��4�~�i�U4=�p`@`��!!�Y����:��'Z-BІ�p!�D�fB�[CE���*���)
?!��{������wĜiC�
̕L!�$�2�T(r�L�`�
��"����!�dC)x�R51h�b�l%�T��W�!�$�Q���{׀)�^� �OS�!����a�n�
5�f���&�:@!�Dٍ E,�� GS�>%���3&{!��PI�	�����fy �y���MI!�D��w��I1�/!!	��Be��x�!�䋧OqΝ�6I�"sq��q�睐�!��4�`K�l�=Z�>���%B����8.Ѳ����
Qe�zG�T*�yF.-`�ĻN�?��u2wÞ��y�F��Ȩ��cAH9�%	wI��y⁃�y��i�K*p��ɫ�JJ��y���*[Pt���.�����(�y��ڵl���2'��G;�h٠-���y�GE�t`�e�J�l��m!/Ǒ�y�۲s�(q ��aw����nS�y�ux��S�������3���yR@W�\*b�����p�ś�L��y��	j )�s*�<xݜ�%���yF�2W��X���8pGn;�+���y"#� � 9S��:C�e�ԍÍ�y�.ڳw�0hp�b�Sa���y��ھp�B,�D��7�N5!� Թ�y2�ׇg%��(A�����%���yN� g���8guY���-�y2��<kV�j�,�!e�A��y�'5clZ|�V�L	w�б�o���y"�P</�,�HTi�"4�7iF�y3X���l�&=DN`�"(�y� �T�Ak"`��铅�y
� H��q·	ylH�!�� ��0��"O���1L%zgP���1�$���"O� ��D����3�hZ�'�PJ�"Oj5(�bW2(Y ��g	к1�*$��"O��B%�iBV��b��IH���6"OB�W��&�r�KΒ ��Y�F"O�i�� �r����s�щR�
��"O���vCJ�&�x�Ҕ0�x9C""O@P{��ٓ8�&��"/�x�����"O�����2���am�,�d9�R"O@l{���h�� ��
��v��Lq"O�ݱ����w$��3I�'yD:i��"O�=��M	�2&�`E���V�C"O:��0	sb0��i~S D�e"O4�ۄD�5�>5�'�Ob�ke"O�-�M͟r��÷�ˁs���a�"OxH+0ǅ81:!�@=D���T"OB�E��MXj���]�W_<4�"O�,Kbj�c�(��-N� ��G"O�\���H48~&�S3OT�� �"O�(a׀�0��x�`Άu��AA�"OjH9�ƀ�O*�@A�0 �zUb�"O�m`ȏb�*�R1ރ\>�50s"O����A4N��Ջ�h��"O�Ube�޶I^Q+Ł��$l�!�!"O(����"\�%�S炔3M2� �"O�X�6�]�"\�ZV�\�
dv-�@"OIx� �c�$+E		8���'"O��W�l��Rn��{�@�Q"Ox�1�Z=�X9��g�!�"O��&$X�X�lh�"� ~*N��"O�8f��;A�3��$r4�"O�(�sfS�Uz
���D\�c
�aZ0"O>�-Y8�óK��!N:� �kI�yB��U��۠��0dTh)�cy��hD���Y�5�vX��KԈm�,<�ʓ,�>���@�ےp�  ;>�C�2t�e��aT��j��Ϻ&u�C䉊Q�z����_ϲ�:sǚ!5��B�I�q���u��Rq�t(��+K��B�	�~��A�7�� ��Hؿ}J�C�	=-i4���i$�p�ss��QI�C�	�������7�<c�(�O,�C��2V�	��+_Kb��R��:I�BC�%��-Z�fI1"M.�s�G��C�I
=�`J �^�3b��#�OY/�4B�	k��	���?��yz��>�B�I�7t�c�S�x��@Њ�$�B�I"h�0�iVc���q����J� B�ɤ8�^�s�/�;�l�@cE4B�m��lJ6$ⲱ��@�c^��a�ĠC C�*i��+H6U�����c]����/�1v��br	��-����ȓJƄ9)�;W�x�z����IS��ȓ`H��AŅ�?����i�9��r�VM�1"\�PI���H� r�^���i2za+��S�h�0Sc�~��ՅȓI�e��	<T�3�@�3}�|�ȓh'^�Z���s�xɠAi"7T,܅ȓ6�d� 5�AM=�H��p7�t����-^B�,��`��cá
8t��`V������}'�9���[=J�Ѕ�ȓBe��l��y̰U�V��2ͅȓB�ZU3��H=V�T�X�c�N��S�? ���!�ϲf-�-���S�ڠ��#"O���'�)Z��= 6+�:l�v�F"O2u�U++P��j	�hŮ��"Op\1l�N��}�B�
~R�"O 1��뚀E�ĸ8�N������ "O�d��ip�@�%m�6�U�"O�� ��%B���Q��0i?څ"�"OX����ڐc.��X4-�G2� �"O��t�L��Z�lٗ{�q��',-"� ݃b9���ΎX^p��'Dl8� �ݍ2C�lJ�������'�:����ֲf�B��E��<��գ�'����Q�3�F!U��;����'�j�)���6�<�"_"��@��'q!Bg��?|��d��U��H#�'���@�O��v�cD���R,�'�Z�"��|_.��7�PLjb�
�'��`-��Y���KgM�Aiji�'}��:@̊6+.(�f�L�
댼B�')pH�s&�$/-�DI@1
�Ԭ��'a ��`�I�}����A�J���
�'t���eE�:1�$\+TR0CK�k
�'�:p;�G�j��D� #��{���	�'w�qb��2D�^���΂\���
�'�b��UGcƭB�FӕN_4���'Y
4Ċ;S9l��BI�B�8P
�'�z�c���� yb��ҕf$Rl
�'�x�
0L9U[X M��Hx80�'%r=�u��!_S�@�3((T���#�'�^�y�
#}*�Ȁ�Ix%D%�'�*PJ &��-�c@fݠ0�'m@�#p7�b�R�ѐb"�@@�'�\K�#��2�.�	��V�`���	�'I���ܪe�4I)Ҥ��h�	�'"r��b�?Vr*�rE��bY�a�'���#v���j��qe���	�'T��(eٵc����`�+ҘP#�'T.ٷ�&�4i���\�2 :�'�ژ(��Y"^H T�0Y���
�'���: ��
6���XAS�;���
�'�j(�T/L!и�pH�	D� ���'q8�'��N�RP��� {���)�'�$� �Oӷ�U�&�}��i�o9D�dq� �N	�p�� �����,D�	��E�o����a�/?���U�)D�����
I�bm����9�����G$D��i�l������:~���
0D���gJ��􃗣�.Y<� uh>D�d�7�J
M��!ѯ�8T5��'D���P-U
���"�R��.���8D�P�d΂ 0i�lY��Q�1��m��"3D�@i�Ȅ����2����+!M��'?D��8E���Du�(�Q�K�0](G�/D��x5��@x~P�F͟&�@��K-D��A@�&�0l�ANV3g?�C!D�  FOY�M�F�ӥ��r@��S�/D��QUE��U���C��_�=f(rN(D���aK�G�n�9�=4Hє`6D�0��G,(n����g�����T�!�$ٿ	�H{&���16B�kA�!S�!�D��l��Q�cĭlxT0W�H;�!����%��BV�<x-X�� s:!�$Ŝ>����60�}p��V�XY!�N�O8@Kc#>)���c�I)�!�� N= �ϟ+�i���� Rr���p"O�Z��D�{�n��U�	�?�VH�"O�	�r(q�>�[�&�?Pv��1Ǔ��2�u�K�.���a?<O��8�(M�4�`�4�R([�p`9d"OvpӉ���csk\>�~(S!"O������,D�tЄ�W�;����u"OFQ)wL�&Iz�TpJF/G�f��q"O� !&D�Fl�uK��o��-��"OXؘc�EH,hᑢ�46~H�8A"O�d#f�P�F��tzGJ:N,	�c"O8���O�#cp�!��鎧��T�S"O�d3'A��8&\�� z�AT"O
T�/��B<p��&Ƒ+H�T�c"O�!*�-�px�13U >�0]�F"O }�5!����Z�xLܛD"O��b��*I��DK��>R�JAc�"O�I�V��e�l��"P5|`���"O$��7ûg���Iw@��t���"Oh쓀EV�I� &	�d����"O�)s/��h�*��$'���"Oi�0B��gh (VD������T"O �A��A�����M!};4�1�"O��@��sx�����Ի=?���%"O�Z����llZ ���%j�jW"O�!���X�$�(C�L�D{J(:�"O�Q�h�$��+�� _r�up"O�QK��RGj�|�N��uZL��"O���6�چB9�A�f�y@�I#�"O6Y� ײh���uhXYB%��"O]�"fY�C�����EB�AA���"O�!���(�X�2"�,�9��"OԤz�f�>M�`���P�ML]R"O���J�IuЈ��!�>�+k�<��Q�4P 3��� c��i�P|�<�V �Uu-<�Д��C�<���L�pq��s�gC�� Y��C�i�<�v��e�����E�q�D�J��c�<!@�Oh���P�#�4G����G�e�<!5�٬0�4�v�Y50~���!�l�<�!���|� �&̊m����F��]�<�c��S6��+c��.,�4�����<�(��0$R����*:�Ν�PGe�<�@\!CVIѣZJ��8�+IV�<�F���y	$-�F�]�A���(�Y�<�v.�+\gFhs�I~lJ-���T�<i�-�Y��K���]����Td�v�<I���>
�����~fP���L|�<	c���2I��^R3lѰ���n�<	�a�Q,��c��|� �0Əh�<�4��&�$�h�H�(J�:\�u-V~�<������`q"f��?�����Ky�<�ƃZ�=���/ľta�ѡ ��v�<�Ǭ 5?ؼr'�B?��IЇH�<��$�~�l�i��0>p0J5g�k�<��b\��	���,	�bt�!�Dd�<���CvJ���
��-���p�J�<�&�T�;N�q� Z3�
ɨ媙a�<Q�
�h��yxv%r��h�+�^�<�Q��M/P���j�.S�<��	^H�i�v��//,�:��L�<�j�6h���;Dh�JRfhR���p�<�ա]�}] �2��
��|d
�d�<Ya��4~�N�*p	P�`E:���N\�<��Y� �d��ܐ�Y�r�Z�<� �!KCIŉx��Ťߺ;Q�9"O�1j����xdIӄ[�� "O��g�<aPm[V�0r���W"Oj8�EN�3PЍ÷����`���"O5��
�_Z�d*1&��}뒑��"O&�ڄ)�\Q�7��4t|Q"O� :�M&ޘsi	�Nh�!�3"O�(�"W~�=v&ؗL��+�"O�T�U˝*{�[�%��?"2��"O.%�W@�0=��-9�$��!�Ƞ�"Or��0�U����ɞ�t����"O�@�W�)L-����	��i�����"O�X�G#x3�%˥FY#rh��"O�!S`��T¦��deb1�C"Oz�[��0)\Ds	Et|q5"O������s����V$�@"O8�
#ۨl��֗3���:e"O�ay�c�3FJ��0�a��ZĈ��@"O�9���2�=	�/����d;f"Ojm�C+���(Y ӭ�5�:�#�"O��z��бT��	W�V�L�l�b"O��ҷ���'���6n��"O���f�\��A�DF5A��s"O*���AQ�?'nԓG�J?8���S"O&EAv�͡MbQZ��`���"O6����:
�a`@�	U�u"Ǒ��M�+�~�S#���:� �X�"O&QK�Ȇ�&߼�Y�fI�%o�!� "O>��c�R���t��*0b�Pb"Ot�鷏��M����BH���@�"O(��V鈧	p���21A�4� "O��{��#W"�<����^̤R "O8͛�*dj���c�÷�t��"O��c�,��$�.�I�Q"O�H!�.�� 7�b�y$g�<�!��;wP��I�o���³C��N�!���<�R��&�np5�6HJ�0!��4j}੘g隹^]�A�;8!�Au!6�"Fm�ظ�ɇ!�� ]9�ܺ�É�Up=���r!�<D�Ga^�1�P��Q�U�!�d]	+�N�	`�\�����!,�-CS!�,(t�a���Fq�d,��:#!�è&\��' D(��MQ䍙�|�!�D<7����I)pfةDB	�!�Ğ��(}�t�5f�������R�!�D]%]��2�RoѲlp��W;$�!�d��l��È���r�@��/�!��o��IĨF-�R`r�A17�!��F&u��m�5�ͥY��{���$�!���s���͘)
�~I ČW�E~!��V9Vc`�;��G�Fj^�S$%L�u�!�d�	�D�8��Y^b2���F��b�!�dZ;&S|��1#�GC*M2�V!򄁎d#�٣��,7(\��V���<!�>=�jLX$���d�\7!��W�zQbx`�"�8xl1C�`[�:��'�ўb?���G�X����W'� �(�s�"2D�(�c��/*���!� � :8��O.D� �3�'Gw8M2��߆eJ���@*D����jϮD��=�f��BD��J5D����oH
��ab�	D�\��i?D����j����Ǆ�B��A��J<D�Xqr↕P(Tщ�{�āCQ�;D�� @�h�A̮��i�'��3�N��w"O�p� A�1�XB�'��:��0�"O�I�(, 2؟rd����"O�I9K\ g��1 MR�&v<���"O��q��K��I��F8i_�D��"O�h9���d��H�~�Z�b�"OdY�̢n���6d�`��p8r"O��Sg�ɨ�E�r���A�"O��c��߉^�D�f��e��}�B"O�� ��ЬeʺՁ�@��I `Q#"O�%XJ¿ ׼�� o�2n��p"O��儃�*�� ���Y���)�"O2�93�&W�����F����P"O�P�K��U@%�q�8�6��S"O�E���۲X�25z-L�/�.��"O�
S)�=8�lh� �ڜY��"OB"�cH�"h��e/�|IE"O\�PT�Fz��Ijɒ0�. �"OڠC&㊚BlFGF�5��8��"O��B`�Q�O$���c��|!�"O@P�4�F�D3"�D��;u"O��6JQ�C��!� �%U�HUѓ"O�M����7i�u��@3Fm��q"O<M*��Y=Tz��=�&��"O^��Ξ�rn(	���8G�d@sR"Ob�8�Ǉ't�*�j��9��4!�"O� /UL �"́�@Є���n���y�h��e��: 05��dh����y�+�HB��cU��1��D�f����yշ/�,�`F�uT��%� ,�y�RV�t܋B���h�t�Ц��)�yr I;:7ڤs`�oyp����K*�yB��x��g�0�AE� *�y�LF�A��X���^�N0��[��yR��v�I��CYB�xȇ���y�ޓ6��y�eϩG��)��_��y�ۡ�ƌ{�#�Oײ���D��yRm��HPq󢢀�OS����.Y?�y��-f�|�R
�W�!zB�� �ybhK!C�� ��_c���H"ˍ��yr��%w����-C�D��a��+�y2'ҭ
:����7�x�*����y�Ȼ6B���J�5,�p��-�y�o=l�@����
fo!q`F;�y��"dM�p#R Ѷd;�=p�)J�y"ib��X!���E�DM�tcҢ�y҇�"un�+fV,��I�(M�yB�R*I|r�X��B#\`����*��y"�^�s(�1���P�bxY�%X�y��ͳb�ItBاK�����ED��yg�X�P�Z�A3@��y��;�y�D�*AS~�����5�آ6�y�k��$�"q!��ؼ{j�s3�_��yR��2�#q� � e���kU��y�"��M���V��5.�,�`"��-�yRaR
[��M0��#���Q��y2��*s����P'4
��ae��yb��$|�P`)��:AYx���ا�yr��H�4X�C�M2��bgCS��y�ҟ'�j��R"(�`J��ҋ�y�͂������m�Jy�7̝7�y�� 8(e���(h�z'��yB�X�S�6`�`"X�Y����6�E��yR���|�p7(����p�n�
�y
� +p���_}�	ku&]��s�"Ox�XD�7-(����N!C���"O��㥥�
>�r���ƫ6v��aV"O�y��A/�`��&#�ĉ�"O d)�J@�g�X�R��Y>���"Ol)��	څ�,�� �Nn ڰ"O�����ƕf��:L՞(�����"O���԰i�
�\�������#�y�jIg���h���$�x3�'/�y��r�hQv�N�q�
P&�V��yB/W+S�vئ\�}F�4*��T�y§��z�q�o�:F�~�{�\�yBl�3 ��ˆ&�@��������y��O��I�5m1,:ԁ��y��1l7����)��e}�	��(��yrj��QV�%a	7]�"�h�J���ybĐT*���ڈW�[��3�yBC�cFr��RdWWe�ESa���yRC�.U
�"���le3��H"�y�6��,���#	>XT���y��J>�cգE�,��i�<�y�<3ш���ٍw�j�A0	�	�y2���[��y`IB�m��X��`Ҷ�y"+�*Y�9��Ll�ZU��L�"�y�� j��4�pb3`�.�"�� ��yf��^6��:�"��I(p,j�P�yRm �5��U1U�]�H�P��`&_��y�m�i�Z��̇�u
��@ރ�y��ق%5�����دmT4�#�LC�ybm��ܐ��*U�f�.<��)�yrI� Eo]�7a)X���Է�yr��~Y��p�DQ(�P�B��y�/V �P�G�	VH����$�yb�z��xsC�¡0������y�	ň9��Ҧa8R��u��)���y��P"��X��J\(-ymƪ�yr�B(qLJ8�4ŕG� �+E,��y2ڵ��Y�
��<���W
�y"�O9J � ��X-��A�.�yB���v� �!��y�P�����y"WB
����7t,,dPFJH��yB��8f�)���݀f������yb�H�8^@ D�̖ear�ti�,�y�'D� �bt�r��k�(�@�g�%�yB��'7bIp�vp�p2-ϓ�y��S�<�JA�t�T���\��y2�P 37� �s0d̓Rʈ��yb�W,3d��Ӂ�$A�4q&@��y�"�^f��y��K��������:�y���34"Jѐ�dV��v�#Uj���y*��GR�����A
{l��4#�3�yY<w  %�ǧj�1��!=�y"�_�T�v���mT2�zi�fh���y!��Ms���/N^lX���yb-�)Fr���ӊ?Z)kt́�y�M�?D�ui���2�H�S���y��%F8�P��
 .�Ik���(�yR��L��ѹw�ѧxÆ�]����^A���JK�wo41C��Ѱs�ʌ��1�j��tĆ�@��ԫ�ZZvp��4j��toR�^m}���\#�t�ȓiyp��$L��[�"- CԔW�\M�ȓ@�����<��������D��A�Zt�2O�0z�N��?TT��S�? �Y�G�P=�(i舁&բ��"O���b���S�~x��'�%s��Mҗ"OJ�`���1��`)�Z�:�|̹6"O8Y`/^"=�`���ƈ#�v��T"O��Jr`�87���d�H^ꝳ�"On��v���G����b�̐LLd�"O����U���KX�l3\A�"OhH��V/���kJ�Ɩ99�"O����J^®� �ME�g�Ʉ�K���ҁ���:����l�v�f%�ȓG��i4K�tQW�Q��ȓX<<���_�|�Z�`@*���p��~d��iF�m�`�M�$`.� ��9n�5!FFB�i�ݡ�+�u䴄ȓ X�h[eO;zx���[�Y�.��xF��sAD�(�2L�TeZ1���ȓb����-��jaP�IW� �O�U��.��X6M�'YK�\��+��eI�<��J�ұ�EfS�Y�a�yjx؇ȓn����� \�A��aDP�|@\��ȓE�h`eF�% �\�qq�U�b�����o��I5呶ox�T�2�o-�T��$ �AP�E����^Y�@��ȓDzZ����fK&�G��A���ȓ@����q/�{e~��T+ކO�J���yU��i��(����B���'ў"|�0N��v�By&a��c:���z�<ag�}P.�D�W���=C�H�Q�<�0D�?-�ChD�!%\p��
M�<鶇ԋ%h)��B�R��:�Dp�<	1�X<����bN�7zQ(�I�h�<a)�.0H4�r
�(�#���d�<)wL%&���+����W�t��!B�a�<�u�^��]їI�do�47��r�<a0fp���7���W��d�KSy�<�W!ݞX�H8a�,1"}$��r�<�@OJ�	����nV���]��/�o�<����R�ȓ���s��x4�Jh�<���O"p!��ɖt�qA�b�J�<�2�� A�$�"5�	}��X��C�<Y���%@bM�WN�+H"b�ׂ�u�<��Bӟe�����"��8CΝn�<��%Q=ӆ��teT%Z��&ea�<"��+?k���t�ˈ)5��C�*c�L���,�3�t�j���{&�B�	�6��`e)��?�<|{��\*|��C�I]J*d��(Y8"���x��C�	K�t�Ӌ�b_�	('��I/tC��:Y�&�J�섋�c_ge�C�I�vU2փ
�L��[?x��C�5&�L	�w݊gh��@���6-C�"%Z
ųB�V!`K� c̃�h�B�6���pq�X$R..ؐ��݈H?�B�I�.��p8��	:Rde�gg�fҔB�	��Du���+[ U�X9weC�	�uP�m	��f�T���B�I��z���f��&c:��b��B�	�)�L���̰.�bh�� ^��NC�	�m\�X���*�( :�`�6�.C�I;��x��L"���%kf�C�	-�L��wK�4.|��Ia#E�b��C�	�^��<���^ c��
Ī)ĨC�	<-�d(��ǌ�b��,0Ʈ�#�C�	�T	:l��kץtx�uɒ��@f�C�)� (�[�O�5/�`3�ÉG�J���"O6�*@��Nu�1	������T"O�cU��u\Њ���+�XX�1"O�4�7'��9haW�+�A�p"O��9v%�5𤰱#�,	�6Uæ"O�,�u+��xX�ա(��h"O�)A��Ԭ!`��\[b��P"O|�jVl[�qF��jPe�?2?�)�"O�]d��%H��1�$Wk(�I�4"O �ѕ��'0���bз:�r�"O9A��� N&�	w!�C����"O.1��"Nt�z�� F�)���:�"O�	1e�ݤ���s�%���0[�"OZ�+��������ӛ<�Yi�"O^��m^�A9F����G�:_@��d"OPI)�,ˇh�
�K¤ʵ_N�PP"O��b�/Q %\m��F9-4��QD"O8,�BdB>��i .���5"O�J��O?��cf�8{����D"Oޕ é�<9�Š7"([���"OT�ҁ��K�쀺c��Y�y15"O D���UA%&�1��"܊DK�"O:8`Q�W8�v,��kɀ+�q��"O`�'��Ld�,��I;
�(�"O��0�R�8��%I£ٚ`G6A�"O�ͰG�[ ���GB 0K<2��G"O��e6����1V�dJ�"O��E	N�\p%GC�+<|\Kt"O�H�Piʩi�<)@�ʨ�ۢ"OZM��lB�7Z
�{pH�-p����"O�%�`nޱ*���3��4g�����"OP�&�)fsD� '�L�@h�%"O ���2�j(����M�����"O��[��
.M���k����ԛ�"O*u�Wh��pM��GU*G��}`�"O�Hu���OG���gg��ZT����"O�Q�e��C�0XI'&�.T~9"O���BLN6+
Q��=|��5�a"O�u�Dς��4�rE)�b���"O�0�P/P�u��Ě�c	�h)�!"OPE�%j(�Q3"i�=Q$�s0"O��1Iܰ,�6Zf�y�� �U"O��;! P�ِm�C��.�D 03"OdAŗH6۴�խR� �"O��iRΓN����� �kmNh�t"O:-⅍L������.��"O���'�(�+��ީg�b%;P"O�Li0"_�r�%5�)C�`�"O,Eh�O�X>驰*M�+��)�"O���Ǫ��Cv��r>�izs"OrQ��Eɒ�*�ѠKU�@َ��&"O���;=��E��F���G"O�x�%&%Z�̑�I�����~�<	��W(Z3�h6��Rx���Æ}�<���>�$\�����F�n��+�|�<�eBĪ,>�����vlf�#H`�<���F�{G��H9��Ń�S_�<���Ғ� ��A�O�0������d�<ٰ���PH�H�+2l���ڧ`�H�<��N�E���*��ҵ[�BM��<QW-؂;���0s�-t��+7a�S�<y�E���m^,c-�嫳	�D�<�鞥'sVp{Vf��I�n��6�X�<�gkK� ~�|0.�:��}�"b�_�<� �1C�h���$�*�M 1W�p���"OV�S�Cz�D�w�g�N}J�"O��&�޷��{�fώ4t�2"O�ݳs���8�T���!*8ɺ0"O���ъƠV��[1k�9L�8�v"O8`yB���6-�`��<-�q"O��%� =n��ț4)�B_@�t"O����í���Jq��?@�I!d"Ov͹�K�7x��y�®�&W!�Y�"O$�!�ճyVX)�-٣rzb�3"O�H�h�(7=�x�dAN.�s��O��k�ʇ��M��O?�	(}��4���O�R��ږ���~����G?I�&�P��8_S�u`���I�b�>����M�N������*&��AK�i!)���T_���Cb�(h���Ѡ�o\F����՟4?���c���?M�TѴ(-΀8p�M��ꧩ�O��d9?�{��M��6i��y駈K%5��h%�]|?���°>��"ϟ�>�"Pl���b�+�B8?���y"�v�6�$;����m�2+H�eh�g�Dp�l#1b�&����mZIX����(QɆDv�_E�! �Ö�\�BYSV�ɜXR�a�6B��rU�����Q�D"<a�,�)$&F%��a�:"u`�'C�0<�2��䓁.ޭ*��,u6�a�O��tIcHي	d��hu���5⟜6�Z�ȇh�2-��pN��?)��?��]���gy��'��	�w``c��Bli�@iу=0���D,ғA�#gI����Ҥ�ɓdv9TN~����5�d�.�D�<�F�ϫǂ%��ė�O8�Y��?_wh�B��V���<Q��_5�c�V:l+<!��%�ĮQ�"B)<��D��{4�xb�ʖ�1C�"?�
ܼ`��@���	���@B�(��Q����:�� #1�i,J���cCRh�VW�O��P�'����Q�U�_��y"��v�*�����J7��O4��?��*�>�P��^�q �52��M\�$��S�LH<���=<z��eэ;n�(�d�Y?��jf	zܴ��ě�5fډ���?����X-a��D/O ���7��So�5��Q��Iԟ�� ��/����[2zU`��$FX2d�)��K�za�c���]�Fl�2պ00����⯂�~�ny0�`�iW6ܐ�M�/�.�b�IG7Q�1���Us��#G�	퐸��П�ē������۴�?a��*�1A%P��#�*1�p�Ag�ߟ�?E���H���̹}u�	be��&)n�0��)�S��M;Vӟ�-x�
��S����d�4B��O<��S���m�	yʟ�Ox�e��(�*eiխ��q5���y��DS����e��\HD�!;�-x��I��G._�@�X�2g&4͚IXQK��M[�߷6*ۧ��*3X���s���uL�����*V�\c{@yE,�1e|le���<��Pڴn��%����Z��i�(�
��ļ_F���ubN-M� l:�'-�'�d��a'x�9�M�EDM���d즁�IB���Mũڮ��5��+T������텍Q���'s4t��	� =���'�2�'����M��y�-R�H_�p��b�GѼ��=0k��q�&5��
 _����Oٸ�Gx�@N2����`� An�H3D�e*��R��4AchG�I w |�	��x�在 <�-����<��bR�TI� i�&yJ�9�))��O�&�b�'�6����D�O��n�%�(P�9������{��І�`�'�@HEM^9���Ң�pCLQ�_˦��4��|Q����䓙5�FL<# |  �   -   Ĵ���	��Z�Zv��9/���3��H�ݴ���qe"�$�6@; <r�il��aDx!Ei��K��+uň);��6��ΦA��4H�{�*S�.��LZA���A��5�̴��D��O(I��48���Uɂ�;��`�F,^e�R͕'�ڥ�۱:-��
,O�pI�o�s�꘠[������"�v<�F��"�@�	�K:�h)Sl�C?��'}8ّA��W��'Xj�@!�� ���EϝK^�Ը���hdpDx��}�'\lΓf=\D�E��.���q�I��p}��%�0r�+F��'�&]��@�N��h�fQ�-6�5h�' �Dx�j��'�Z�+QeI�|���f"��.�n���,�&"<Aڪ>�7� 9����c*�gx~L��M�O�$K�Oeq�{2�`�����]
�>�(W� �M�,/O|"<a���2/(iӠBA�4r ��#L��>A�c?"H��o�j�H�GN�P��m���X.R��͖'�BAEx�ȘW�k6+ӡ�]������	��ʶ�,�)�(#<�!��O���Ԡ^�.F����M�M��4���dR�O,L�L<A�TU�8s��6DV�r���G?q�%&*�LO��98[$"�8�f�c�C�9ϼ��q�_�$�"a��i��?-��I�E㟎�R��8�N� �@�]��}ʖſ<�G���;�D�'�,H��K�8�tO����L1;轰��K	��� ^�tڱ�ɾN���R�+�x��h�oǇbhje#�B<D�����   ��ƊI�X�8��%�<��i4���R�'��'y�O�A�1�`����d�#F�����?�����Şa$���C֨X�K��,�ه�>�ȁ�\~y�g�$|o|��,r��'n��A��|3v�
����r�\&B����럔�IߟP�i>��'L�6���ys"�dҏF=��ᶁ¸;P����f,Y$��Xަu�?�2W�����X��\�^��3��AF�� ��P��u��ȦI�'�B��6!��?��}��ּ�Z���1��3kZ�����?��?���?Y����O��3���
mq� Y������W���I9�M3�jE�|��sA��|b'[Q�!l�*= 9��.k~�'�������ݹt��֓���6ÜRX��ϖ�M���'��!��O��O���|"��?Y��N��u��j�u�jY~Ah����?9*O��m-b���џ    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  ]  �  �  *  z5  �@  L  �W  gb  �j  �q  9|  ΄  �  ^�  ��  ��  >�  ��  �  R�  ��  ��  M�  ��  	�  K�  ��  ��  ��  Q�  ��  �  K Y �% �- �3 : �?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'_|#=�̋�/hNȉV!Õ0u�(�kRD�<Y/ۥG��P��7��`yW�C�<Y����:�kBJ��e��`�F�<�#�;  A�ц0��J�ܦцz���MK����gTl�xe��bx�ad�$@�ih`$W*Т�� ����A��H@H�a�1E|"F���'9�'k6&I�%ۙb��4����+e"���ȓ'�t�I�!�%jJ)�mW!v�H��	��HO?�)��A�bX(�h&H�\A2��O�<A��Ũ��a`�G(k��Rw RVy��5�O�TS`��C�����ȅ���<"F"O xS0/����x��F+k�H���"O�i�&m\*nچi��� k�P���"Ot�*BS�smK��8�!H�ż�y2�3^'L��1�A*q��'T�y"�u��ԉB��J������-L��ȓ:0p���U-
�ބ��DDOlZ	��#w~�HD��~�aUi<cl���Q��`
&+M�5i H�w��u�ȓMq�p�)�.� y4�P��ȓi�,�QDT�_1��㱬��n��م�F���@�l���ǃ�5
�rL�ȓ�R`!�,�f�"������5��}�ȓQS�}��j.n�j�@�n�
5 �Y�']�������J)�#��x�N�(A��x/���d]}���?� � �ۀT1.�HD^��y£�^�����ѽ=T�⃢Q%�(O�܈ç6��Y4J��n����ÚL�e��Ah����;����fA, 8х�v�������p=VD�!�
�&�j��ȓ&��ܣ��F�P\x���ɰW~���O�-�f� t��b�'N+ ������C~"@�Zt*q�S-�2KPXI��i���y
� ������D�aƈз#Df���"O���U���~�%��H��%��]�"O�]���/h���ƪ+���i�i�ў"~n��"ݲ<q�a«r�<aq��F��C䉹g|ށۗ)<U&伃��W	M.�Ɂ}��~bD�������ۗ>n-B�@�˰>aش���B���$�s$�l%���}k!�$ޟz�Y У�D�rE��F�-�џ�D��`�#��a��W�c�0m���>�y2LBmW�{4"ңUX���B�3��D=�S�O2��CX�{AS$,�<���y�/�6�+�W�����tdQ�Ƙ')�{���GOd���`�t!�p��J�y��	�<
 ��sz$E&�H��y�9Hƥ�ĩ spP%�E��+�yBcF�;C�}c�?��ɵ*���yr	�0_zA��	Փz�T�U�ĭ�y��çe0
��W�Ǩa��K �7�y��֫wnX��GQf��B���'xazek����F�� �b 0���yb��)($X�ʡE,f��Cg���y2��$�@�S��䁣	����j����>Ec�G�")R	tds��%a�K9D�x���ʞm��*� aX6���,�i���O Xa�w	��k���gj��?Z���
�'�
 0�Ne�!8�G75�8x��O����	�k�`)�b��<	\4��"OЃ�i�&	�Z( #��(8N QQ�"On��/;P2��#�W����Y%"O�h�O'N��<`�S@��c"OUA挼{4J�Ks�R�8P��"OL� 7i�ǜ���Ǌ<�d:C"O��2��թ[��lh�	Y,-``p�"O�Ube��u��٘V�I�����'31O�}�P�S�A5z��!�ofx��"Or���ptH���e��B��b"O����٣MA���1e�E��<)�"O��P ��b��7�F�MdLb�"O4	C�ӼRq��Zd+ ��s�"O�ǼL|�Qc�b̂��e"O��X� Ֆ�!J���9��a;�"OX�S`�D5b��q��w|�
w"O
IX���C�AqE��(�b�"O
��O�#%��0��?�<4xd"O\*G��|��	B�C@�:�J(�&"O�x�!��!�v��$�Q�$% g"O��J�,�t:₃���nȪ�"O�h�U#
�TS򇁸D}x��"OB���;@�J� 5&�Np
�ap"OD%��&Ӛ>E��UE
�\ff�)W"OZ����>���wҖH�
�b"O,�Y�C��C�"��딐[��=�#"O��)l�U�=#(��Z���"OF�ڔ���D��MJ�f�l��(�T"OJE�"A�[��a�C�W�q�$#"OxŁ �߭=TF$p�cI��F]"e"O�c���)CUv��6��q�"O�M���ıUm���/ rep���"O$��G"�W������2rH� "O��֎�?Y*�;��R7f�yW"O���W�\1k�E�`+�%Pb�2�"O���po�g�:t��,;��c�"O��� E�H��W�Y��R� "O�q� ���7'.Ց��F�����"O� Ќ(7�p��q���8�dj5"O�	����DM3���,L�'=��+�hѷ�f��55��1�'��؂�,A�_ej�c�W�9�(�`�'vd+�s���� µ3E�ܸ���?��?��?���?����?��2H������؋�jJ/UL@���?���?����?����?���?��+��b	-}d��r�g��C7b����?9���?)���?	���?	���?)�-��,sp�Ĩ���3
Ѭ(2�T���?���?y��?����?9��?��&�Dux4Gĳ}>�$(�*��4��H���?���?a��?����?!���?I��$��!'a�ÕhY�P��$��^ҟ���ߟ���֟\��˟��	��8��������:y][�'ˤ<�5h�/J��I�T��џ���矔�	����͟D[p���3X4�*֪s�ڱ8ӊ�˟\����(�	ܟ��	͟������	ߟ��r��?o~Q�E �-^`L��ޟ�I�������	������d�	ܟ<@JR���YAD�.Z�2%��ş,��ǟ���ӟL�	ПH�	ޟ�	�CP���@\~X  ���h�Н�	ޟ���쟜�	؟���ɟ��	ڟ���u�F$��ߺ8��$���������D�IٟL�I�����ǟ��	&.�~��d��ecv�<Y�@��IƟD�����I�p�����i�4�?���m�6�Іʿr�-�'㞁9�B�h�]�0��Ly���O��l�u.�yS�����#U� m(Q�Gg9?Y��i��O�9O��Zu��p`� �>� gT�
}���O�(�b{�D���(��OzR������|OЊ�`
+�%R�y��'�	^�OR���5Ƙ:{MAX�"13j�`�!�yӦP�u�d*���MϻeX�2�a1oY���hL�m�<Y��?Y�'��)�Ӥ'ټLn��<��m�)|��+Wo%�x)��<�'�p���hO�i�Ox`��\a޼�� F�L�m�0O����vL���ߢ��'��X2�	!�� �&g#� Ѵ�dT}�'�R1O��t�t�`G3Ğ��!��0a~�d�'j�KٓZ��tI���k�ӟpI��'�>a���@B��o�P�G]f��IIy������!9L�YziP�gʔة7I�;�����Ui9?9��i��O�G�-���K���>�jE�c膎:��D�O���O6l���n��������ZD!܃?0<$��$��{����O2�䓄�4�����O>�D�O:���h@�`R��M������Ւ(O�l�#����	ş��L�Sş@[�?$�l@�	)}L�lإ� ����<7��O2�O1�Z)��m�="�(�#JU'@+ܰ��%s�̞z��	�
�z����'D�U&�ؖ'�XH�2S�x���▪i}"H�B�'��'����4]��������J韨��Iդx3X�"��@��$�b�}�Z�x��O����O�Nܷ\�
��ʉ2j[��[W�bC(�x,y���^@<�����(�2H~"�;c��\;�MV�8�᠍8
j����?Q��?���?	����O�L��W�F�ֽ`R�¬d��ta�'b��'Ir6$Q"�i�Op�oZQ�	 Fv�d��ٶk�~�rT��M�N$����Ɵ擟,���m�[~���2V\E�g�ޣLdv��L�&Q6��u�UU?iI>*OX��O��d�O����0O�	K��hA8�@�	�O��d�<a��iT�TY$�'���'��_* k��X��ě2�/�������?�O��M��I�X]�Qa�A~�;�Y)q@Z�A$ˑ$2]�i>9ye�'��P$��Ѣ�H<q�䚔(J:X��d�Ac�ПL��矰��ޟb>9�'U�6�)���!Jȣa8�m���O�q�|�p��O���X��%��I�����OҩiB�S ���à�.|cdTS�,�O<��MZ��6m&?�;8�����'yc�ʓC�b�2퉹'3��2(^(HTI����O����O����O��$�|�$%��!P�t �9<����"�W~��N�D��'U����'~6=）�����A�'��'T`20��O,�b>��FC����q
�LW1�J�ue]/���P�EQ��O�չH>A+O,���OP��!j�!z��hDǛHj l
�L�O����O��d�<q��i��|y��'�DE7S�1!t��+�;)x���ĉH}2�'A�|� �!F��TB��0֪Y��$=���� oa�}�e�C4,1��y��z, ��֓N	��k��_[�� �a��-m$���O���Oz��>�缋�AS$5�1�%��1�B�@�I��?钸i��1V��*�4���y�F�r
\a�M!i�}a� �3�y��'��'|�(1�i��ɛd�h@��O��}	��@�2��)l��Dy�`�W�iy�O]��'��'|BfWq�V�w�{t���q�^�z4��=�M����?����?yN~Γs��}�qL��>��C�ΌLO�y{�Y������t&�b>uYAo��1^�i�v�K�=u�@�.�'�C�0?�"�W"3D��������#I�ډ�Nǥ:"�l��� �x���$�O\�$�O&�4��˓4w�6g��_�b�.
0�|xb"<|j���_BB'kӎ��8�O8�D�O���B��,��ˌ�/���E��B
֙��gb���b�) b�?�$?Y�=� r�� ������c�� �yr�?O���O��$�O����O��?I�ߧfV�-�3���DʽB�� ��l�����*ݴ[��.O��m�i�&h<n����%a�>D�ֈ�Q�y&����ԟ�S�.$�l�S~�	���%��D.�̌ ǌC-c���Q
ӟ�Bq�|RZ����� ���<�R7nP#���Y$m��*���	}y�Ff��#I�O��d�O��')!�p��BἉ؆E�
���'����?����S��l�s/�;a���v�	�]輨C�O.�~��`�/��4�N����,���Of�Y�n �F�n�F���xf����O��D�O���O1��˓AZ�v��2\��n�T9az3�
R45"sQ���4��'2듩?ɡ�ʾ	��ݨ���$��P� CQ��?��[ł���4��DC-s7�9����M�5��2$�!`��3E�0�y�Q�X�	ܟ(�IϟX�I͟�O��SpV+�`a�oN5����kt�~�A�*�O����O���Ҧ�ݦ>�ʉ���T�.�
��ME�v�Hl���%�b>q6�@Ѧ��I�Nipѣ�'t7��)�^<H�=�}�g��O��H>�/O�)�O��(�Ө[ڵ[��
�$��G��Ov���O����<Y��i��җ�'��'l�9�oПf�� T������u�O���'�R�'�'|��tj�B�<� P�(��C�O�y蒡J�B]��+��&���&�?y���O���U��E���:O�X�L�O���r��',b�ԟ�_�x���H�^�P�9�D[:!�n�dQӦ��e�˟`�	��Mc��w��z��WS�pq�	���IÝ'�V��Xwc�}�'�0�	*��?�z���\S΄��,b�����GZ>W�'��Iğ0��ٟ��IΟ8�I<D��6C�&"MH� �?m�ԕ'��6MM�7\����Oh�2�i�O ����oȥ9�jȤu<�@b �n}B�'#Ҟ|�����
��ۃa�Z�Nh�Ԥ2���{�i+��&��84$��d$��'`P�ۀ�^�j���vH�#�N��W�'���'�B����Z�Hr�4@��#�<���k�[�;�聻F�ލ}�Z���gt�6�ĐZ}r�'�	�[��� [�8�iw
��$A����M��O<"MO-�Bg�?�)��>�kf�&��]� D׎����<O����O����O���Ol�?�r�g �3U�`���[�v;:�u�W�P�	՟@
޴d����-O lZf�ɧ'��+� Lo�L� 
�`�xm&�(����ӷ!��po�]~��ɕ/�t��F��	LN�A`���?@HU��kG����Д|�[��Sҟ��I�H���Ҳu�$p�+��U��"�.��P�	Hy�	qӘ-�P��ON���O@˧i�� �-W��fū�C�5p��0�'C4��?����S�䉏�G�~Ҡ� O&��f_���{N��xi��O�	ސ�?� �)�D�W�h�V V�fmа�cmӝ���d�O��d�OD�4���D�OJ�F�➨yK ���/Ϝ=\�@��4a4�%���'�"�g��O��$�K}B�'��0ʤ�J<:����O�]|
 '�'Q�H����>OX�d͕ct~����x�h�v�"�
�d��I��@�1i�=7�d�����O����O��d�O>�D�|j"C�����$I8|��l1 DȊ>��o����'
����'N�6=�-�bM�T�
0���=F/����O��$ ��DG%z7��|	�兏�(�b�)6��4'��`?O�x
`j��?s<���<�'�?IaDF"p�t`C��1�r�+� 1�?����?�����צm��g�ޟ���؟�B"��V����RH#z���Un��Ul�	埬��K�ɧ^N29�p#Y�^��s�H�)e��x�RY�$T4�Mp��d�Ii?��l�>U���s�B#Tɓ�h��!;���?����?q���h����<b��|�tG��F��L����(����̦鉃,_y�}Ӱ���4q�f�K�kS<7mb�F�Zd������I���{��A즍�'�i����Yr�e�3;Q�H��-���sr���䓒�����E"�@�ĭ<����6��eo�I%�Ms"G�,��D�ON�?���$�lb�Y6˔�{�N�0��M����Od�d&�󉃮+�aJ�! �N��[�&#�����l�M�ʓ}��Xj���O4H>I/Oh4XGo�w�ʕh%ȟ)�ı���'q�6M
O�`��$���%�3JG�Â��x���̦1�?��R����ϟ��	<�f]�fnGJ��r3a͖Wr4ѣQ��m�'Y^��D��?�[��$�w&,s���t�y��$ 
7�\��'�r�'ar�'	��')���B�`���>��N�U�F�?����?y5�i>�Ma�Or�m�X�O\1�FD�Z���ک
+����4���O��4��a
y���W����@�ڨ*)��*���2o
���d���䓋�4�v�d�O��4A��ّ�I�V��$b���qT���Oʓ+�&��1z���'V�R>e���O�| �i�r��H���'?�6T�H�I֟�&��'�hF��*�l@�$"_צ�(���?Q�4��4��@Q�'��'p�#§U�U��#� +5]��:@�'/B�'����J����T� )۴3����
@�h�@�r�g�I��XA�/�?���Px�f�|�O����?�6��=8Y��[�qo���OM �?y��N1�<#ܴ�y"�'{>������?)+@U�� de�V`��J-�����M&'���Q�5O�˓�?���?9��?A���򉌬}(
ӊ"�=�׏��xn$X]�I��|�I[���p������hӄ^�\q� �0�/L��?�����S�'$�.��ش�yB�Q).������Ӏ5��{E��*�y�*I q<������4�*�$ض<"����J�Z�8� 橉�"���$�O����O�ʓ8ۛ#�E?r�'�"�J�QpN���i�f������RE�O ��'���'��'��l����Cj��y拀�\h���OРI���2s��)ҘO�Bx�	+R�r(F8R��`C�[Z$y���L���'�b�'�2��� �a-X%i��!�3Ql�4��K�⟘ٴ&A`�R���?A6�i��O��9g��A��$�ix�c�2|���O~ʓ�d��ݴ��D��L9�!���
g���j��
4�0�@��)[��A�d2�D�<���?���?���?���'�����	(d°Q���$��i���۟L��П��� ��h��2�$P�3���V(�+�����Iu�)�S8(��` �i�8
���!�c�:��As�� ����'����G�`�"�|�W��H�·��օ �I�e��y@��	��4��ϟ�xy��|�.����Ox��DL�0�C�-�d�(���On	le�ϟ8�O��D�O�N	�sl0(�(`����S<)4�"vӢ�O�Ȥ�e�?�'?1�ݜ~�"�˳AQ� �����A6�H�I��P�	֟0�Iҟ���^�'�(���� �̡&��� �J�Ο�Iȟ�
�4x�*��'�?)��i��'��I��(�2����қJ�J��|��'
�Oٶ���ie�ɫk����{�YR#CO6tB�O.1=��3���<��,�-{���֮��[��Ǣ�ODlښz��ݗ'��S>���Ꮨ+pP`��X'���É4?�"_�8��ӟ�%��'6�` IFABr4<�&�V�MS.�q�L��V�� §��4�P�b����O.�x���,SB�����0�F�"FM�O�d�O��D�O1�XʓS ��(�?���6MN�q�|�R�/\eW }��'�Rt���t�O����!Ee�L)�oP :�\�:A�K�^���po����4���Ȕy���'�.��bh8�L�*��ݫ"��(\*������O>�d�O
�D�O���|��I�N�`�y*D�@x�"�o��'b��g�&>�R�'/���t�'l�7=�|��f�E�U�`��&�(�F��O��b>��sM��Q�>�D�����e%F�����e�,�lA� v��O�iL>	.O���OTP��ԈAВ�	%�$V5��֌�O8���O̼��l�<a��i��(���O���'��	�gna��7d�
N��0�|"�'��I���'�`�ɭ[�iZe�s���'"�Dр���D1A�Qw8�HD�y�O'B��I4��#'b��!�ʛs����N;�y�J��fJ0��'생rgܡ�ŭ�.���v��l�Bn�<!ǲiz�O�NͷZ�F�H�Î��|ݢR��^��d�O,���O�r�+y�x�ӺsPY���Ů �,}����̝f����I̜yD��O˓�?���?1���?)�8��	� V��AA�Hh���H+O4o$dk�P�	۟(�IN�S۟D*UD��Zf$(#F	E��ҷBE���$�O��b>�P"i�;pF����	�:$X���� M�q7$my�j��gU ���@��'T�	3u�Z�9T��4-[\A���� h܁��ן,�	ϟl�i>�'>7m��d�1M�}��\��Z�Ӊď��dS����?��Q���	��I,;�Y��NX���8!kU��,��Ǖئ��'cx�S��?��}���u� \1a C�P�xH��#H~�̓�?����?q���?�����' +��*a�G�D���(��H�y2���kɀI��?)ֲi]ڌ�6�'�b�'��'������äK���c&劓<�x�ӈy"�'��'*�a��i��D�OLy��#�� ��DB�*��'�z|`��Jn�#��V��Of˓�?����?���	��h@�Ğ�v.^e�P�ւz�؋��?y.O��lZ$M6����|����b�h�aOA((95h[��y��'�ꓑ?i����S��Î�=O�ش,�,L���3N@?��C"�:ua2�B�_�操}�2�l�	+q ���rkƠEz6.U{��I����X�)�Sny��y�Z�PQ��$+�A�S%���h}�%��
d��$�O�!ln���Գ�O
��)���2D]�0��s�	=u0 ��O�M@��fӮ�Do$���ŷ?�'�0r ��,nV�A�Cؓ8����'5�	Ο�Iǟd�IߟP��n���S�����K	�T��-��66�Ӝ����O��D3�)�O$mz��x���*n����L�4�t���_���?�|zq ��M{�'�ą��\I����&C�&n�i*�'���p��ir�|2T���I�ث�N�u�j�e��c�pP)�)���P��ȟ��	]yB�x����O�O��d�O$Y���8�@ճ�^�"��ht(3�d�O���'�'��'8���P`W�0$(d���&�4Q��OLP��տ�h�.��W?�?��&�O�MQ��&\�t���N>��G,�O*�D�O@��<�OuR�'��
'G`�51�/C�g;�q�$�P���y���P���O���O��O��4����G�a w�218��¦��O����OZ�$�%2��7�e���I�eTp)�Ms�U�� �qz����V���3iA�w�B|��'0�D�<���?���?Y��?)bbM�Z,���m��-K��4� ��dM����p�����I�d%?�	��=��lS?��@!�?q$*a�Or��O�O1��䊄I#*C��+%��[�4h�e 6|1�2��`��ʘ@iBe{��Yy�ٻjZ��k
�(��1y��3�0>��i��;��'���w��R[^=���ĵJ��$��'�7-+������OT���OB	)&m�pQ6� �ٹ�<�cn��)�7- ?��o��Z@��I]���'ҿc�!I�.��x'��^3����(��<���?I��?����?�M~:Ζ((f�u�vF_s}�M	nK Q�N��*O���N���Ĉ�֟L��>�M�K>���ȑn2$ �@eL���\@��<Y��?��%��2۴�y2�'<�9��3f�0��X.�Da�+S/0�D(�	
CW�'��՟��	��	
<1k)�ȀO�>���I�� �'�.6��������Or�D�|R�4���3�o_
&$�;�b�Z~�F�>9�������8*�~4I�B) $&ybcn�7h���(XPd�*@g�<�'9j� ��(ڴ�4M[�>E`�� �ű9(�����?���?�S�'��ͦ�[�ō�+��=�P$5�̽ S�.� �'�6�%�	���O�xg��2y��š\�|���7e�O&���8*Ϣ6�2?��L��}p��i>�$c�z�>X���Q ��T
�y�X�@�	ퟜ�I���I؟@�O�nِ&��)�%��I��/+�=Scosӊ��%��O2��O����d���s��+âت���oȇQ�@�IQ�ŞX����4�yR �UP Q�(�%-�q�����yB�5��I�I6p�'��Iܟ<�	�����B�
��5s�X�a.�(�	�����'�^6�I�˓�?����H��!��L(�v��'����?ɉ�ϗQ���2�Z+t�Dh�g�ԛ��D�M蠴�v��)5�`�������7�����#@3|E�Ƀ�,�b�Ȧ�d�O���O��$:��SՀ�C��=�6V����P�5�?�ջirⰣ�Q���ش���ywN��:X�P+E�W��:�S��ӽ�y��'���'-�-jW�i%�ɢN��=�$�O��hr�V+=DX�^�pH@���V�	by�O�2�'�"�'r�%���i���s��,�� �
�I��M#��J��?a��?�K~�n��4
O�L����4�X*o��ѲW������h'�b>��M�F�Z��@W5<�vmc��ңA��iĬ/?���Q%L�n��X�����DЮG��U$�T�o��Lk牅a�,���O��$�O��4��˓,��� �!M�����L,2P-޸Dt�Dj*�2gӢ��2�O(���OD���9n��c.�\^@0����(�Q�{�l�6��PXf�;ʧ�q |�T�q�%u@L�� C�<���?����?���?y���lG� �,s��P N���؆E��T�2�'�-y�@��:�$�$�M'���J�	v4��.b3b @�4�֟��'2�1��i��ɽ>�t��N��	|��S� X*<�s���/��'�m��Hyb�')��'
R�5����`�.;�}�!�<��'�削�M�j��?I��?�(�<ũ�g
� �j���{vn�`����O����O��O���j7��G��K��� �˾D�(�vf3C:�D#?�'m��d����\�Z�Q�B�(1��Q���g���c��?���?a�Ş����mC�D�Mrĵ
��l��CgCݐ�H��'T�7m9�	��d�O�m3D��Zx́pf$�v�rᠠN�On�d�<p9l7�9?���t!���<�$��� ��@����$� ��yBQ�\��ҟ��Iϟ�������O�%���רdJ$���BH �2�#y�h����O���O�������V�������30r��n�=�����('�b>������]͓���:�Ӈ|�D�V��MuLuΓ"О}@�A�OY�L>i/O��O�t  (�ȡ ���=Q�!�j�O
���O��D�<��ib,��'&�'��:g��,	v��Ѹ#��	5��r}b�'��Oh,����aT8���c2sM0�PŜ�tbc���(DH�_�����S͟\��ݶ�1�w�SEڙ+PA1D�d�Ɓ �&�D�3�`�5k�l�A4�Rş�
�4o�n�����?�R�i��O�n˪6"-�i4?j�ij ꝼ0�$�Ov���O���g�x���b����7��?msV�\Cmڑh��s��k5E�d�Fy2��,D��yk�)MDx�H���
v��.�֩QB/����\��%�	#v����-Te���G������(��F�)�S�A��5
a%��b�T���� G�L�3�f[�\��'i2�@ڟXI�|_�X*6�
7��4F� ^��aE���t�Iԟ��Iܟ�S@y2	rӲ��`��O�d@$ G\DD0B�G�=R��Mh�2O�l�I����� �IП�a�M�!`J�Y e�1a_�u㵣�[�̑mZ}~�ךB`�t��Z�'�����{}sR�2r����B��<9��UM|t؂�'z�������Z�0E{-O��D��U�:��i �'����R�L0n��4�MŖ�u꒙|��'��OlT���i��i��
� ����ߔ�.���W��S�d;�?� �;��<���?����?����� ��V/o�$��1��?q�����禙�C�ʟ0������O�u!r�����5+ɵG��M��O�p�'B�'�ɧ��̽[��<E�~�t������=� ���ՠp��I�M�}y�O�����5u��'x(8��W<OL�h�C�Ћ-�,Yh��'L��'tB���O0�	��M��ĥ l�-(JĿ줱jP�R�X*O��o�C���I������0��S��BQI1������G��lZ|~��8�V��}�P+ٙT�@��F�.��B�.�<�)O��$�Oz�d�O���O�'j��)7�l���97�E#��
9�M��Mэ�?���?�N~���L���w�4,���V [�`i��T�aՖ)���'\��|����̑PE��8O���ǂ��`����00��}x�>O�ȁ����\��p�R}�@ z�E�.��=A!IF���q���Qp��T��1D�Ȋe�@�o'�XR��K�O�L�ņ�n���[5e�:�VT[׆ǯ9�gi�3Ik(pA�9m]d�!E�=�8�hGgA�YLP�8�Z���`��h	A��) �^-�� ��"���0
� �(b�kЏ^�B�pw��;� ��� GL�X��}S�B��N�)�@��iJ6��
����`ǘl̑ �(��rw� ���N�8�0=��&T
!nHܢ���B��TQ��^�_�m)�!J0Q8��w��
I����ñi1b�'�.��#�8�$a�蜒6��o}�t�1���Ov���	���s��}L̹�#Md�� �2��v���Oxʓ5�J�yg[?��	��ӉZPl�&�F�Wz��"J�4c0�O<)��?�'��'��i��g	���
M���dM^��\��r�J��M+��?���"�T�֘�\^��e��3�T����(l��7��O��$	7i��⟸�}��+�/"�\���OѪ!�p7��~mZ����I���ӝ��D�<��ᕪC�,	�HW�?�5�����7:���%���|B���O|�k�N_�Pd�PE�ɦa����զ���ݟ<��4-��@��O�ʓ�?��'�H��FV�& x	�	m���4��V��5����':��'u�=c��T 0�l	:�'�.��zӒ��V5R&���'��I͟l'���
,�p��Gb��a�D��.Hv�V��B����D�O:���O��A��ic���z���D
���*Ԙ"3�IVyR�'f�'�B9O�h�#/N#S�j<sJ�*\ �������'l��'��]�P��C���(�$"��A��hc����Kӻ�M�,O���)���O��$[�+���I�\d�٪�-�l"阔�ǒ���?����?�(O�B���d�4�'e�e�PM *���j4��
�tF�z6��O�Ol���O���J2�ɫ ����D�$a�"L��8[47M�O���<�/���ٟ���?��Gĉ$�H�����7���8"�@2�ē�?���G��Ex�ܟ�9�b�<C�;b&Ï^����i�ɿ?|qܴ�?��?��'G��i���1��v ��K�6 ��%�a�d���O�1���O�O:�>e�Հ��Ok����'cڐ�GMd��I�⩕�����T�	�?IN<�'4��ԯ�"uV q'Á)G6�}��i�b�'��|ʟ���Od�4���n��]ȼЖ�ő'B\l�����I�p
1`����|����~�.w���CsY��
}#0M �M����W��s���	����Iw�	���9\���XcN�G2Rly�4�?�⭚hh���t�'��'�$<����'�Ф#��0l5ak�g2��O0ʓ�?�.�2ʓ�qA�L�R����=Zj$	�7�P ��'�r�'�'��i�M�%�v���qǬ����*�na���D?��O�ʓ�?�a�����S�ZKm%�Ϭ-�t�Dk���M���?��b�'��	q��6�\�p#Ã� %S�u8��[�^5�'prQ���	?�,�O�k޳A����aتn�TQjce��D�d6M)����,�'-���L<�!�%5�j8:qFߦ{�!Y��[ަ��	ß�'/>P��2��O>��Ƽ�Ҥ��&s|�1��.D�rѵi���ٟD�	˟��IO�s���-��.f&L��b��q\��4�i�ɺ%�V��ڴRs��ҟl�S2���9O+��S��
�+�%ФʰY��Y�P��˟�J|�J~n�$ ��=�&W"��-���Ȍ1a�7� �a�^�n����؟��ӑ���|�獒�	d���bCF�h���FQ	�?���?�����S��OD�y�.K�>&����9��%���ݦ��Ih�I�]�4X���	,}�����@G)�,9xAP�
��\�"<�a���O��	k���X����j�Vq���j�P6��O��G�<i�R?Q�?�W�̄/���R�*	�Zp� �]�(�'�H�O��d�OH�Ģ<ym�l������.?�%��@w"�L�a�x2�'�2�|"W��C�d����'?�Q� �b�R6�O�˓�?q��?	.O�قF,��|z�ǖ�p�Y�j�=����j}��'�R�|�U��ȟH�«L7p0f��,8�� ����?y.O ��S��'�?���g���ơ�uVl�(R�`���$�O�ʓ
�� '���IA�e�$ب��F?}�amy�l��O���nؠ�����'��\c����r��4�z�Z�D��n:�,yH<�-O��$�O���$Pw���{����bO�L��a��i��I�'7��޴  ���T��6��� Z����'��)����Q�j@�!�i\��'z��'���d�|nZ�T��S�`�,l=Vz�	Ah6͊�G��an�ڟ���П�������|2EL�Wl0�á/�x���Vh@�'(���'��'�ɧ���pbSb�87CP�Jg�=5'�0Z����M����?��*�D5�(O�SE��UR�u��_�&] ѳ'�ětH�XFxb�6��O����OJ�sR�`�=���^�bdD�2(�����!>�v9P�O���?�(O���ƴD
���:h���.\6䃖�i�b�ʹ�y��'���' "�'/�I>5�d|�t��r\R�17���*���h�9��$�<����O��d�O������Rg�I�&"�\�P��M�����O`�d�O���O��!g�a��1���I�,�N2*0RVB�7�-�d�iA����'@��'��b��yB�٘XdY�p�I#>߈��b�Y+G'�7��O<�$�O��Ĥ<��cZ����˟0�Em��o�� ����_8؅y��S��M������O����O~�g1O��'x��J.8�0}iD*I����4�?���ݸ����OU�'���#ܤ7�t���ƛ|_ �����)(
2��?����?�(��<����$�?]�A튝V��:��Ny�
݂��rӪ˓n.��b�i���'�R�O�
�Ӻ��Ȉjc�`��,��Ip���L
ߦ��֟,�f�i�@%��}����^4\����^X��BɁҦU�1�K7�M���?y���*qY���'̄H�,ҿ2��]�bO�^\�h` z��a��4O��O��?��I�Hiqa�hے	��r�� ƴ�޴�?��?�ŋ�*���Ry�'F�d��C�$Y�p�H"k͐�H�<ěf�'剻w�,�)z���?�O���"�A�2D���2#�n=��4�?���T���qy��'����G�p  ��=�:i�$Q77-�O�|QW3O���O����O���<����\�*D������e�#'� �v�	�Z�Д'm"U����ߟ��	%b.��vj�h�
p��`��c�����)e�x��ǟ,��֟<��gy��V�~�8�G>��0ScT,r����U�rq6ͦ<������Oh�$�OFi��?Ok,�'�X�c���� $�����꟰���X�'�����n�~��' ��u�<~��س�f���R�i��^�0�	ןt��&����s���=^8"(�����H��S*Lߛv�'�bS��b������O�$��X�(t���/
�г�9a+f4��"�h}2�'�"�'��q��O�����Mn��Q�����mH\�i�
�5�M#+Op9��
�㦉��۟T�	�?!i�O뮇6,]��%AE!qHU(��N�i���'���y�!�~Γ��O^�;����:�8�D��|@��4b(t`�iy��'���O�j����oV���lĞT�0���B	��]lڴ0�IF�	q���?I7(Z�s��HP����-��� �'@����'���'�|�T̢>Q/O2�ĺ�����D
Bt���7~�*��#k�8�O���p0O����H��ɟl"�
UЀ@�MˊG� ���҅�M����m��X�p�'q\�t�i�]ڠǒ�?�����½9��k�>�n��<���?��?1����DL�V�PE�9�+A���-�b<�rA}�_�@��Ly��'��']L)�E+b��ę�"F���U�տ�y��'A2�'�b�'� �v�y�O��%3f�˳u۞,Z��%Z��ݴ��D�O��?q���?��(�<)fl�y@��%ؔY�ju!����Iǟ��Iߟd�'�f ���2�IE�b���f�\I�顆/G�i2(	mZڟ�'�T�	ڟ@ti�����Oflx#�=NHjP���'�8��P�i^��'�	�-24�K|r���#�J�!�z��Z��T	���'�'��e:�'j�'*��	�&����΂-+�j�%JґV��T���^W}B7mD�d�'3�TH4?�V��kj�Y������uB���O���O`��C�>�IS�'*WM�%�Ic����� <M	v!nZ��qr�4�?1���?I�'2m�'��h
�{Ė�ۃ��AMČs�	�,A?7Q�W`�)��8��Ο�[a�A�8H���0S��e{$�^��Ms���?9�� ���k��x"�'`��O*P��ݝy�
Dɓ�Y�-�d��i�'���Xr�1��O.�d�O2�;���v���+�������b��m�	 K��L<����?�O>��2�B����y��(���l?��'���8��'��	�<�	؟̗'!�����S�@2���
�-'�L��C�K�:O�$�O��O��Od����2m� �o�}�t��!.�s̎��<����?�����D ����'2��H�� If)����!����'"�'�'2�'��V�'y$��ѡ02TH�`f��Na>8)`+�>���?������$>q(Ө�y���S#��aS(��C��MK����?A��9*� ��� Z��C�o� :b=r���
@87��O��d�<u�Z-? �O-�O�8�t�G6G3���dM��29��q6���Op��e�*�D&�İ?QS�BQ �ݙb���*��d�n�T�p�Լ8c�i]�꧃?��O�ɗaԪ]a6i�$z�q�C\%/
6��O$��Y�\�t�$%�D8�S�/N���N�z�(��OZ6F7]��~�o�˟���͟���1��'I[�.H�G���@�eM�w�6�`Ft�\�(R�	{���?�D�
Ϟ�AQ5X�|�#Y�69���'?��'	�DbSI'�$�O������ ^�9�@�	-�R� $%˦px�XŲi�'�����%���O �d�O4��lW�����P	T�n����Á�����	�7B(a1�}��'Iɧ5��[�5�D��e�>w20- Â�9���E;L6�$�<q���?y���Z�s�eC�K�fJ���L�Isp|S� �v�	��d�I̟��'���'m��S���`^�@-D�0�\Ļ�����'���'x�i�oZ�ެ���5���� �QO���Ԏ��b�dlZ��t�	ş�'�p�IEy"���M�tl��\���G\5]R�z��Z}B�'���'���N��(�N|�`�̏45�A��DZ��l*ܶL����'%�'�����@�Ʃ!�i6pz�1�Ҡ�x7��Ot�$�<��� ��O"��O��9�����钁LBv�Qec4�$�ON���E�@=��^.B���
�%@Jj��X�Dk�C���M[�V?��I�?Y��O*8�SD�&;G��B��]�*O̝`��izr�'�����d5Ex(�/	&�.��5��j%�72�b�n�����Iȟ`�S����?�ÃԴ!*�qv�R3�� ����ۛ��X��O��?a��:���
�l�ʇ"V���i�4�?���?IԪ����|B���~�BF1%&���R�4H��݋D���%Ӛ#<�E����'��'Ĕ,�孑#�Ȁ�eP�TP4a�iӴ���:RP&��՟��IT���	v\sAd͑Ku$u���47���_`�b����ڟh�I����	w�����nL�rE���2��$*��Xy�'U��'p�'T��Ox!h�f7\�YC��cI�1�i&Q�O�$�O��$�<y%&܄k�޽p����ʋ�P�l����ԯ�Iן ��S�	ן��5-�b�C[H�sD��.��%�E;J͈e�'�R�'`R\�����@%�ħS��T�Fo����9*VMM5!�N��C�i�ґ|��'�����'Ɛ��"��[�d|2�Ƙ�Z���:޴�?�����/SI�Y%>m���?��raK��8�o+Xc$H
�':�ē�?���(��eFx�ޟT9�Q��a�D���I��/�)#��i>��s�6mcٴ*������ӈ���Nm'�\�Un�	�r�!O�u���ܦ��	�&#<ى��$J.9�����B�2Gn-H�	�M��'3q��v�'
2�'����3�$�O�	�����S��D�D&ro�M��_�	{T;�S�O��II�6fJImv�V\��	ƪL��7��O��$�O*!Y��Hv������	U?����Eڬ�⌆�1T``����q�5, ��<����?!��
���!��V��XD��GG�4	pV�i�r�(��O
���O��Ok�ƆH�D�KϽGo�����<���+�,c�D���p��wy���>oxj��m�Z���SE��@m��6���O��2���O����{���S�Bָn̝��� ##h�`����O,���Of�7XL��F2����qaK���h�&�,FL�ԟx��'K�'2��'�L��OfP5曠
2h�Y��ѳ4��0q@]�T��˟���Cy�G	56��F��wb�s�\�A�̖a|T�+�h��i��O�ޟl�ɯB-,c��قm��C���z����9����`�s�����O:�0h�����'��o
0��y�Pf� ;���u|�7Ͳ<�(O����?��|n��fy��EF��l�!�z�� 2�[;�~�\5�4"����{�D̤w�$� d�/A�� E S�y�T�G���ϝ�"�
$1�JB*%jRqt��(����,Cm�����V�@P+�M��6�Z�qgHE$9R"�ȥ ��A� ˕7@,m�WmA�=vj�*���gf��CE�s�>�{#&�4צ!�'%Ο#h|͑nF�"I � �1<{h�`ឲY�FHy�9G��@>6ʹat瘪'0b�'`��'�F�]ȟ��	�Jz�Ʈ#v"����:O�d��w !�"���,�j,�GK�?E��_%��EQ��߄	Ւ�FcZ!�ɣQ���UK.��S�T3pyd�xҟGy"��0�[$���zޔ��"�,�~�aݢ�?a��hO��{+b� �;h�`\c�M��8����/[���sU� O�|*���&gju	E�)�(O��#�����5JWA�����Qk���.L��J矘�������L͠0��͟�Χ:���7
��G5����AΙ�F����,��+@��ju6$@��Ǖ�X@#��~�}���: ^�U*��XO�~��o�=*��y��X�?Y��R�HeQ妍�6+�uґ)�X�v ����2�'VT��sE�Y:�P�1i^�[�ny�ȓ[��Q���K�M���Y��ϓ:���Ryb�ɭ3tD��?�+����@�d�2��aNJ�bnܬ�-	�p4r�$�Od��Ͼ.�@�zDኳt��T�O��I�0��]6	�
a�$L��Q��RʷHi�q1E�ѭ��O�۲��5�b�XÄ�4+�ȍ�	�\$��'�񟀬1��	}��[�%��w_ Qp2;O���
�nn�@�`K�6�����ىj�a|b"�C�X)�9�1�4t�x�cE��64��K�W�
Mm��$��U�T�7�?����?��*u���,�.=:�G'H����ܘ����*n?p�񶩕�o,�0@�-Bl����@����
� �� �[
<���W�DԢE�a�Q���d"�)��P���.��tO�3e��i(D��B�환tV���J��׈ը��1�e����'k�T�z`$�w�� 7$�,m���A���?a'�qE�����?y��y"���4�|��`��pGH)��DH-	"��OR8Z�'a�]
b��#mn|-����a��'���R�e�J��FH��S/$Mq��P>����A>̍��@���`���d�}��h	�n,���6"!D�ڔ�	-� ��,V��m�K��HO>qɄ(� �M˕�Q$ *(R�H`1�!�?����?A�'�b����?	�O'���?�Ȇ� �Y#�B� +0�rF�D8�0��¦<��G�X`�-�,�9r�԰ �}8��sÂ�O���_:	�,����̬$�Π6�Yl�!�$�v ��K��Y�\��	��`]�T�!�*�dM"s�*a�p�[�)Л'M�b��H�dޓ�M���?a)���Z��#�@���%"3�h��Ƙ~�|�D�O��K|D��'�|j@L�`4T��:�4T`$�^�'u�PH���H�B�����7U�&��� ��npQ�T�'�O��}�p�ٝW'��Zc�V
}5�t�3�N|�<!��ϋ�R)���e�4�w��o�|�L<a�+t�`ı�I� b0�R6N�<��QZ���'��?a�7��O����OZ,��٦P�ƌ(�.?"����w�#wgV�D,�|Fxrl,.��šݦ{a����J>?���)�����)I�$����{�����..2.z��IQ�S��?��KQx�:�Q�k�(��Fl|�<�7��%��Y+�� @�hUx�t�'P�#=�Ok��S߲Cւ`C�΀l�B�'���ƨ*&����'a�'H�$h��i��q���*����,2��Q7���~"�%��>	�I�*\�i�6�F-<�p3�E\Q?�`�Nox���Q���h&�C6�ƃ�BK����X0��O�����K��J&�ַ 1�T"r�#D��g�-U����NوB*���p#���HO>�bmÏ�M;U��-R����u�0q�l��h��?����?��'�Hi���?��O��ܸ��?)A�C�9�b	�Ċ�*�Xܪ���P8���-�<yU���	�!kW�0*�}�i�H8������ON�DA�t�����/'Hi���n!�9R��``.�p��V AN�!򤓆"�����f��w
Hk`�2���v�_<�Ak��ih��'��Ӏ
���Â6ȴ��ʟy=��4/���I㟘�%��ٟ��<�O��=!P�݌T+>�bi�5zcx�P��d��?Yaw�	.���@��	�B�le��+�B;�H�	l�O���"#NM.v^}*n^j�
�'�D�a��;ײ@h%��M����W&�'�x�Q��?x���`ʹ>W�T��'Z2Y�D�o��d�O��'}3��Iן���'W2����1�|��2#���PlH���$?e,I+@h�R��|����&*h�h�l�-hWp�j���,Hhh�fK�d�*]��:vd��S��?�@P'g�t���K)X�>�#��O+uR�������h���̵�G�L�y?�@�vmҍ�y"��x�zc�BԚl��%eν�OZ1FzʟƬ��JO�G�VAˀhV9w������OX�DF���`i�O��D�OD�$��{�Ӽ{ Cs"f����'E>T���!Vi?���U���K
�F�����]H��D�U�j��^�%cC(���=Q�'�j�M՚$:��iW����?9�ۤ�?i���?�gyR�'��ICf�`����f�c����B�ɆxSƵB3�U�T���L5��s���?��?!�X�`qD�yr�K(_p�s��D�<q�/�id$���'��<�Cz�<�+S� Q�!ci�2N�5��t�<I�&��l�����Dʌ���&�h�<�&� ���$��41~�i�/�`�<Q��0���R��цP��P��!�_�<	b��v�$m�@�B/�n�zPe�[�<!�b�M @J!G��g
�U*R�M\�< gZ=�V`�'ȃ-YA2T�Jt�<� ��P��,��iF��:�x4y2"O�Q�S��G"�DJ�J;�̈�"O65�ch[� i�F�!x����F"Ov 	��?xŶ��$ٻ#��"O���g[,�ր#���#ڮ�;�"O4H�*�}���P�b׸0��(p"O�H��߁' ��3�hɘ��Ё"O�(kb�6G	ڕ�&�J��"O�d���ŏL�A�&�q�2$�6"O��;��T�i��NPe�aK�"OLz��*r����1(H�.T�ٰ3"O�4!&̜u�A�R�N��u"O�T s��PnY�'( .P��"O��i���PĮɰ�B�o�Ġ�"O��c���}6ֹ!�ʻX3���"Ot�c�Y Z(�8�&yz,P��"OR]� )܈ST(�ԮٻU���r"O��S�I�*l�Ɛr#Ӑ�*+�"O�<����#A���XfK-6)3�"O��s2�XM��!�	� ��F"O�H�'�io�b�&���%"O�IW�"k��)�bL~�@8�#"Of��$d DriF��(@_��B"O�A33�بS�DxI3��%fJ�M�`"O�Aӄ�*uTy�#�'Q_<� ��'W,�`�'�b=�vJ�$~��K���*�<h�'�%f�x��#�V�s�ƍK��$�h��#~5��Yl\܁BCָ"J�_c�<Y�I��6:Txa���`�+�Hw��K�BG�S�O�y ���IfP:` D��P��"O
ݒ2m�/U4�1��E8@��ȡ^�(���h�L���2�j��𣅑W�TE��I9�ODe�I��8#T��6�:��3�P��"O��cÒ�P^� "`M3m�쁶��8>���D�^�	ɖ�(�F�>ҭSRǝ��y�B<
�ؘ8aϫ.Ƞ�Ff<����k��H�X�'O�JXT��AL !�:���"O���7Ɛ.Z6d��E�O��p�"OJ&�B� G^�;��]�ٴYc�"O��2Dm��F�XP%� 2u(�Yd"OB�:s%����j§ l�D��"OFS��qu^[GM/UZ�(��"O��:��~u�p���P�NF|!�"O��W ����U��4{0zt�V"O��aq�@!~��ʴ�W�E|�"O�|����"O�C��7-u��'�,=��	D�$�'����Y� .N\Idhz�^��
�'<�!"Jd ��pcł�ِ$��{;�x�` K&AP����sL��
=}7x-�IZ1�!�d�OŬـ�g�G&�Tbh��W�f�Ԝ>�D�*_��>�O>y��GX��P�B��ݞ�Ve�v
O,|�@T�(�z\zE�F�,а�h��6T5ʒ�Ƨ�0?�BH�J���F�N�B���2�`CW8���G�?�����c�H�F��cVmS�rs�5�&#%D����Ȼ"6]ȓ�N8S��y���!}'؟t��'A>�⩞���<�W�1=x��c��?D���j�i˚��4I՛� ���Qz���'-|Av��a�g�ɾ"�~Q�����^��Xy��+^�<C�I�W�P�ȥ���s�� �?$����F	��X\xx7�'�.X���U|j��(�-<(��Z�A	|��'��I�7.��r�B
L�BI.m��'����G���X�F��	�֬��'NX�(3%GD��q&,�5-|��
�'��a�d�
>4aH�
�*�3O21��� j��g�w�j;�1.P��9�"O��!��'tαJ� �&�Y$]���T@8��k��Я[�RՑ���\TQ@H;�O��&����� �&���$ �*�ޡy��4D��+�Oˀ9���U.�x'��a��4�V\�h$G۠yI��Q&�88���l���j�AO�o~ ��Z�b�=�ȓ7BE�4	@)1���)p������y'LH&)[���F�B'-e����#}λ `Tk�gQ�ao,��Ui�g,Їȓn�|�VF]�
�r��/¢f(HH����)A%Du�&�=o:�-i����|PJ$�A��\r ��*[ε�p2����X؁�w��$��)�gO�Q>(�Dh4xdj�1s"ߠr��%a蓂�|B�J�T�~Qd�Ĥ0��)HRcS��O�mi��ҥiP�)���	�vPQ��ֆ��eP�Kqj���%��$����1J��y2����JB햅W`���"� k��P�D�X+w	F1X�*�*6�`��~7* H3�E)2�K,=�8T�ǆ�s�<���K$U��9�#��Ie(�P�˄�*�ER犔�2(�V�Zu�L��S5.H8�%��1)���S�S��C���)��E��W�<Ա�Ǥ9lO8�H���
V55H�n�D��l�0 `BH���T�Ɂ@V�	�	B!f`k��X�F�>	(6���a��?㤰�6��K�i�$�s�.T��X�8�N��}���m��Q^���f˰}B��[*����+�f�j��4P�����}AGf�4s��4!��-y�8	J*�'��H0qB\3RN�А��c�+�74�6H1s�x�2������Z(Yb�� ��~}��X"OzS$:Q���BҤ�Y��s�W�<�K�>��'�Ҡ�C�D�ꑚ��q'kL	�nߨLx��)ezn�ʶ ����d��ɭYE�uK�L]�P���*8�<�kf�w����ʉ���=^�D�;�
g��ၶ�cQ�+���2>��Z�ƅ�}��T�"�I�p9 �$�T3sK�]�7`;W��O�zĝ�u`�ڥ��
Q���A�w��8YSƋ�p>��%������
�'�|�(d��N��}�D�?}-�x����Q��ϻE`C�`Ǚ4��C���F����iw8QU�})%�v�b�t�r�	c*�A�'��dWna�P���5�4p}U ω�i�5��+πY�Z��퉂&p�4�O+2`�����>N�p	7Ț���DD��?��G�`��pᅤ�;x�D�+�ɂ^�'f��ZdBܘl��Bu�n�m���e�M��5����qY�$Ӂ���	"u�x����W]����.��!PS����?1��	9K��@@�#Q��3����f*�32r���W�b���a���?E��w#tM�3�Ɲk���b��w�� �'�TX�w���Z�I�S�t))@D���?��f�$!^:T2E����t��v�'aF(����=L�JHr��ɗ��b�̾�j�� �p�y�	}��LCqI+^����mܘ��c �T$����>FL� �_��u�
�k �Xcp#�|���	@9l>�Q���O���\&��{ bQ#�"J4�T�#!�Iy���5
O�^��3DCȜC՘ՓS��#�e�Ag����;P��(��n��#��]k���t<`��G��w�!���z�ؙ�bj�C�P����V�n0�Ӆ�9h&�	3��.p|0hQџ�"=I��:�f<0�Mf�8
uX�����\�T|�9�Ŧ
_)�j3B@ �"Y�"��쪠��'1��YPˍ)<e���c\���$֔}�j�3����B�zM�N?�
�)P�z�l�g�y�P�B&F�p$��=��i�&Ќ ���sJM�0�L0̓��
^,��;�.O8 ��gyJ?A9ڨ1$�Qw�RM�K��#D�$�% 	1T4���<6��h�2�L2��DM�5��'�؉��9O�K�N��I���`v��Sa@	�(�"iᥬ�0�a~R`' ��'�I�_��R��K7[A�zu��5��D�o]l��-JV|�pV�G  �g~���%�� ���.N|!0ԇS��(O8���e�"����| 2Џ�?-c�&2��V-��M��W�YF�ڡc)S-]�ə�A ��<�aFG��j *�2����Ǟ�{�v�cp�ݍF B�)�ɹ������'�������L:&��Y͜<07$X1Qpb���44��ItFU%v�~0��(�h"��"S*��T����� �Dt"��<2��"�r%B�]����������(K4�<�2DB���7���m����@�F!<���yA(��_n��	`/Xz?-��`���7��$*v��K@��+��L<a�	I�+Ҵx�V���}�F�B��$��M�e~b�P�h�> tM�6S�y�����?���M�5*�jk�9[�R���*���#b裲.��50�Xtf���<ģ�;g�)��Y�A����.�/��q�@� ?���0;hb"��i�1Fy��Z
!�`H7�^�6�i�'cۮ��D�<�(��v�
��� �,P���R��ȃ����kG�� A1r"���O��_)d���qӆ�b�i��t�����#5)f�����-ғXe��JA�N[Jt���4s�|����_�(`�{1f�I��#�I�4RZ����|"�Y��~+̫qS�M���|�9Od��%�� 
I8���G:T�Iӝ>!��L# �t�P���s=$�@)4�@�>ɔ�B3<#�`.V���IQB�7��eHR�	�Q�0T�E�ͽT��|���'��2	�1�f�aR�&�13�^�a !d`�>b�Zas��q8�`����8=��g��PbpB��ka}H�5(��Bq":^������o~>a��ύP�2��D�0���N���0��,Z�At
��` 3^���EM,�/Ĳ%Yħ�N�1���T�1��$
�t��Hܬ�  �),`��\!�\���d́��.�D  }2�׮����̆�v쥃W&Z��~r�<c>T�k�/�rQ����cG-2�n�qbKT�Bv��'�<E�i�.�8����G�4��T�C �xr�ʛ?[={ B�_8���EB^<i��b��Q#r� ;��đR� b���Df�x��Ij$�臠
�;1���*�;.L���I+~L�@��֢�@ ���^�{� ��u�:�x�ϓ;} ��q
�zrx�pg�_�&tK!�;�-���X����7�Z]ht��gѿ/�@|�6�ɏ:��+�DO<p�@ł@��`S�x�O>�DQ�x�'�L3}q�T�~�
J������jؒ����ʯ\l�(�O�i�'��[9؝SBI[�x�UK�R��X��SbVM��0��%��mB�9�D��o?Y�&�.�
�k4�6LO�\�`�	��0*�@#"���B�
ܥ_����$�B� `�!L%J|*�$S�X�J�ݧs��KA�ۇ!�$`w�/n��C�ɂ=�~m ����%h��[�� غ4����$��N��5�>���[�L�nM@$����(O�}�
	�2�c7m^�YW�`A��'FEhGnۜx3��Æ�ՕV�
&ʀ*j |{��Y�F}�xK�-^� 2���җ7	�|��|%p�IR��&76�C�K��Ov��\�|A���{��qР��&4��O���J�2/�� �Rtܴ�a�'g��Q�7x6����O?g�jh�wΌ�z�o�/=��q"��&�?E��w�"L!&��>q(=3ĄO�� �'��Âձb!��R�/�&�;�(Y�z�X)��k�N)�`B�����I�mX��@ˆw8@Q����*�C䉗/�J�#cֶ��S�IM�+��C�I&@���;2(��SJ�t�V.W2r��C�IR�d�"@P�z��Q)W,JB0B�I4���
&�ѕ*�rE�q��yG�B�ə� �9�a!��R��։:��C��t�\�k�����Վy��C�I��$a�!i���sP�ߑHӀC䉀e?��A5
��{�p�����}�~C�I�*na�GnЖ̈Y�A�4`�|C�I�}֤1�s�ȧR�z���;
n�C�I#	N���	��}����Qo�0pw�C�ɏϞ�qp��ip�����&Q�C䉶� 0ä >.Vu9��O+jC�0���RN_�wRR���n:C�	#&�`RO�.�i$MT�/�C䉶�� 2��R-"!2�o�(V*�B�I�2o��c��\%�I��I"�B�ɺ$�8�0٨[�h�M�&)��B�� X��A�ER[��"�B�(Z�JC�	-0�9AVc�0P��{5酝Wl�C�	4p�U��җr��@X��ŽeO�C䉻l����7!H$��	�%0�B�	���giդs�z�� ՚.��B��: X�UI<�� �gH�c�>C��"|p��#���Is�[�!4�C䉃l��Ať�
�xHQOx!P�9D�� ��x��@���	_��Q��=D�`�U���d�)��V%e�8���n0D��{�e�\e|H���*�2y�)D��� P4=�}�U'�+ЫT�:D���AO
$P 3��l�BQSE;D���b�������,d�tQ'�9D� �Q��Zfm�a��D-T��(S���V�v�0��N|�숈&"O� $5��52��%�7�@e�~Q�""O�%x-�-A�M���Ĥn���A4"O�	�@R@&��{���q��Ś�"O!*��,=�HM!R� Lp�,�4"OY��e��%��!s�)�%=Sn��"OơhbJƯF9�LjT�E�I@�APC"O�,Z�%J�q��@+����:����"OvTX���(�0X06_�9 �p9S"O��r�mF�d�!�a�V� ��"O.ݲG�
:N!s�e�0r�*G"O\���M�+�(L�s��:]0��Q"O�x�aѦ_p��H�cNR�@"O�C5���S�ؼ7KD�Y��� �y�lÔz��b��?*wn��3�I8�y"��0)$�ҮB<�2)��A��y�fS�r�@!�(tH��a%��y���LQ�]��L�%c���R!K
�y��;�H��O/c���s�H'�y2�
�?��}��)�8	����+ٜ�y҅��#��2����
 )��b
�y���+F1�M�R']i(�'��+�y��Q1+�d��,�(p�6�zD���y����
�@ۡe�f 4�R��yCI"
(�Bg� LL��SS�W�y�H���z	�s'0�#�j���y��	!�\�	�z�����y"G��$�6�S�YH �A ϱ�yR	�2)���pc�:O X&��y�E�Q/�5�G���F���bD杋�y��<qD�a�
<I�%R���y�Jˆ{�Uh�gO�.��ʤ�V�y"/��
X Ļ��7YE�\���Ǿ�y�I{-�-���E&����#��y"י)�\<x1�P8KR����?�y�Q�kT"=BE@�D�d��-Y��y�G��7i*p���;&8�z�iڨ�y�;9JP�0��9uPM
å��y"��KP�脨���ҸA�",�y"�8����Rc�" �n�x�k��y �/$t$��A�s��	:�ڒ�y"/�61�H���kc$P���(�Py"�K� �Ǫ�/J�N�1�'H]�<)�)�&!v��c���T��Y�<y' �jO6�a�V�$
�/�V�<YS�M�P	И2X6�Xգ����B�	4t�EI��	qV8�ĭ(r�C�	� bx�� �d���h�Ǟi�C䉿d�f����
�u�@1ʱi��B�I7؆9�rㆶu�$RC���(��C䉻v����委�g�|"�����C�ɁPa̼��E+NU|� %��/SB�C�I�wی)C��G
���CSq�B��B���J�w6<�tO�3��C�I�z��Y1Ո�<�F�i�	�?&��C�0�L,�F$�|!���Q8q��C� j\< s�R�s�8�r����\��C�I+����fX-T�"d��^{�B�	���q��+'��xg��Z��B�� x<�ݢ�
HɞՃG�\�, 4C䉖����C֥z�<���X���C䉒N�>ݢ���L�x}�6$�Ka�C�	`���K=oT����i��C�IY�l��Õ6N�xe[c�I1�B�	6"�M�P�_��
h��Q�30�B�)� &�Qq燒3ǰ�`�L�=��"O�hT�E1N0ȋ��Ӈ+�F=!"Of�XS�\-�p�Gm�{���3"O�`Y���T�R��T�U�55�Y�"O��q��O4��:D�D�<*!X"O~X��#ܖ7�l��� U��c"O�Iz5���\��Mؖ՚1	�"Ob<� )��	V��5d�T�+"O�r��1+;�ɐA6 �4�"Op��A��I]F5)���w�Z��"O�Y�D�������D� x���f"OFe���V>��q�Cd�$P��X�"O�\i#Z�{ކ!{ い��� t"OBtH�D�	=EB1��R�-V%�@"OHӆ�X9;ȁ�SBҙ�N��"O�)�jT� t>���o�0�H��""O�M`�ePZ��`+�GI {�Π@1"Ot ڧ��2$�(�B�	G{���"O>%s�թ�bI)6E��|p(`��"OJ]�ƥN�7��b��ZvV�P`"O(�����'�>Ѹ7h9��"Op��r)$h���4�B@Tܙ�0"O��D(�2�~!��]�.�@�j�"O��BP�)$�b9ТY)z��h�"O:�p�d¾*�d�O-p_T`��"O%��dΰ\%v͉R��+&��k"O����� >�y0�h��P�"O��h2�"rV�`h�7\m��"O`��-t�AGi�(D�C`"O����B�[� 5��g���i�"Oک ���(�k0H^�Ob�}h�"O��æi��oQ2ё����iT���&"O�(��	�^Ö���'.7(��"O޼9� 2*wm#$��\R�lZ&"O ���Y*F�8*�p��#W>/!�$�pjp���W�'��4"V�K!�dU�YXL��Fh�^x!&�G�k!�d���,頴�I�m=.� 2a�-!��	�1n�����.#�`����\y�!�D���,��O��M\d�r�gC2+�!�Ā~΅���ؠ\��\�P	T x!�+IBjh�OG"2�L= 7V�g!���8�,��ػ]�L��f���!��	rڹ�$Hy@�Z�Ɣ)g�!�DGA��S�K.iX� ��+�!�H�p��w,�+[H\s�E�L�!�d��j ���`Æ�>�Q��	�5I�!򤘿IZ�Q �>$4}sF��!�\�u��Ti���Pdjaб���!��f����)�;f�p���Ţ?s!�D��	5F�	@�B�q̤�[��B�eQ�\F��oLM�y�תɤ0���(c�Q%�y��8r@i�� ��!Y���S��
�y"O��.����Y &L<��`T��y��s�0J!�]!f��bG��y� B�Q�,�����Z:�\ؓ�)�yr��
�$	R�ەi�`p�o��y�E�>!�b\�@�%\�~<T�S�y�@ ~�1a�-��`�Ҡڀ���y�,:~dH$���`'`��pkX��yS�B(�T�1C�+Q�4���/��y���"�-e`I����+�'��'w�{��/R�Ja�EL*�p�`S#�(O�5����0��Ԁ����L�pGl�1#�C�)� �]�GLD�J:<A�,����b�(A�Q�"~�	8f�&=H�bQ�y�����D�� C�	\7�T�����B~�}j�N�<r��I�,a~B��Ccd�P�ʏz�+��3�yBEͅ?��p��J�!X�c�"���y2"�!HH"�L٢)/��+"4�yT�&E&yvJ�o�f|���܄�y�82'B9���>:� ��0K�'�p?��OJ�A!F�sl�����`�n@�%"O$X3t �2�r,�`��>�Y0"O��cE�H61^TR�K��o���"O�q9��F�J���D�	� w"O�H����i�����P����%!�d\'p�D���@�5Ɣ|�7�	�0C�	 �$h��D�m���2x��B�I3Y�.��
�	\���D�\�B��! (���E?h)v��W�A�-�FB�	�bJ�mb��Ń}�����:*0FB�Cg�q�V.�4��b �F^<ʓ�0?q���6o��A��(ܶqk�� W��}�<���%c����D��5
srI ���B�<�䂚�ĩp�ЩI*� 6G~�<�HJ>yp}��g��o��d�Fg\}�<�L�:��y�IH�	��Y�fFr��@���O�8�F��xv��<V6xY�'S,��E$Kv,�	�#͆QY�!�'�8%@%�Q/�����X�=e����'s���&kʾ"K�0���@�6�*��'���6�ԍ4ْUI6�($���
�'�ڭԃ]*:�2�;�̅3.z�
�'�X%C4��'�$x��C,y�Ȋ
�'�t�����0K��u`�>?h��	�'���4N1L��;��5k>��	�'J�D��ŵ(�� ��}V�9�
�'��[R�ҝ�f���J��G��K�'������!q�BQ-����h�'ܸl � ړ�F�$L�#�Jm�
�'�&"qe�P��!����
ˊ�p
�'	e‮)1@$���6�n�	�'d<�i�Q+.8!�S`-
�'!�
3��	V� "�XK�c�'	d����5Y�d��g M�%zn���'(Vp�F���_(m#� F%x�%Y	�'�����$aE���F��'�ڰ˚�OY����ͅw�8|p�'ȎX#�J�ZN������s�*�'$��Rb\"fA!�%@n�mQ
�'��a�5k�.p��B�3f#�i`	�'4j��e�q^ ��s���M��T��' h40�M�y���3�ʆ��=�'-�܈'/.'���@N�=
��ɹ�'l xw������Ǉ�4BS�'k@�ЃOj��8��oƮ~22l+�'�}�tcbk:@��1	�'Y�(
&��P�m#�[7�T��'ON@y��Y�J������&UĤ��' t�
��(*E+�#ٮ	�$��'L�=��o[��y�1�W�zH�	�'�6��1�9k.�1FK����'+,|�拊-��@s�ė�y����'�qi���b�`��$��
I��k�'xT1�T78�h�SM�u�R���'�X��i�&G5�Q;\0?���[�'�, �h�	`&0xAC�-a�5���� L ��'�y�yCա݃Gbi�"O��{�D�]����� ��x��\�s"O����H ��1pc �>|�ʘ�v"O��Q"�� ��Ab��:	����@"Oޭ1�� �>0�$EW�a}4k"OH䩓�ԇCb�`��$РLn�M�"O���a#C�"V�铡��t��c�"O���OXZ9��������"O0h*w��%s��k�X��(�"O�I&�ˠdi"����fy���G"OMb-c0~�A% \�x�Ap�"O���C��h��&o�12P"O�ɹ��V�Z�� a�>+��"O�y,�8۴@�OJ(  <�D"Of#�*�7��=w��n��1"O�x)�F�|��d��,M����#"O�,(�5p��%��f�$9A"O��ʧg�0�}�b�0�i�"O�Ak"Q5̝�R"/$"�]�"O,%��#�5&2X���U�����"O�,"6h��
�D�4�ݓ��0�s"O�Dbd�]�k�����䋧�x��"O�lZ�o�!�lX��É�B�D��"O�,�w��5�`��=f��#"Ol�
�D�v���6��k�<�C"O�9��G�o�Xh�LD��L��"O&�ӕ�7E,` �M�c���2*O�yo_*EV���,�-s.mS�'�XAJd"g|�PBBf�Z�Xm��'3�)�u��W���a%R�i'����'�&��=y���RFm� o\���'C}ұ��E���f�R��i��'�:*udO<2��hiՍ�	;W$�	
�'}"��ҪХ)��P����e�h��'��@ku+ڦ▴�p�]�S�$t��'��5C#*��%����䌉tQ�L�'�fPaB	��hȎD��Bk���	�'iT�:b,ڲw&\��e�g�lM��':���`[�#�L�s ��W��i��'�z}b�!Ni��@��!O��s�'����
�`qV��i�\t���4S�ϊMx����%' d��ȓ+̂��F��?��[�LE\��ȓf�R�{�� н+�`J|.0]��@���ش�I�0/�K�>X� ��ȓyg�-�DH�^�8���Q�z�R��P�X
Fn��P@��)�4Zcn��ȓT(��E�'r�F1Z���/I��$��I@e�ԧɴ;��=���!P����ȓm����(MM:y93�ٖ7���j�j��GIR�50N\1�={�܆�U��};Yq�έ7*b�
�r"O���5��`�DӤ@%^��"OP��ǃ�g�V�۲��v/���"O���I���S�K�M+ظ(r"O�T��o�N�A�!�@z���C"O -B0nX�9�Z�B(�G�<1+!"O�U�� �}�Iq4iJ�9�ڬXQ"O��3��
u�x ���@ɉ2"O����L��i����H� ��3�"Oe�a��ry:���{��3"O�HP��^�8��)��X���B"O����Ն\��3�F�����)D"O	X$�K%bn�`w杰W���p"O� v�z�V�e���r��//��˔"O2\�b�B�l|np!��Ǽ �9��"O�QQ�NQ���x�m&�b�8�"O����I��B3p�p5��S�� �"OD�J�,�6)8d�P1I�1����"O��r�90����G�D��a�"O(����S�t�GX@=��s�"O�؉}���D�2J��P1"O��1����rjĤ�I��"��"O�����fά�*�IӗX�u�s"O��q�F�Άt�!#%)y洺�"Ox��&#)ڌ�+� Z>B^��"O���f��B�Y���Z�BȚQ"O������9}T�4JߑB���H�"O^L�������W�XQ"O@	�Tn�+q�P��W�<SmQ"Oz��rk�C���Bgf]�;E���"O<�(��
�o��0SÅ�3��m"�"OxC6�ˡ�F����j
}�Q"O�p����h�4��Ȅ5id�y�"OЙ�G�ծO�Q�GKHX�-�G"O�xu�H�8 "���	LT�,p2"O��P���-Y6��� k��B52��s"O��U�B'h�5��ԓu����"OX#�G�"b����
N��f"O��H4�8n�>��na��� "O�ѫ��Ȁ{���᳈A,	U�d+�"O�xQ$�GU���Q� �*z8��a�"OF�ZGڥ& �����!)���p"Ox���*l�#���,Li�=�ŏ��y��_rT3!�S6�5! a�/�y�� ���5˞:1iF]�W#
"�y�I@���]aU�Ξ740�+�T-�yR�B���t ׭@,5V�X0���y�(s�ȑ����0]DJ�m��-]!��o�zUٵ��,8�(��U�_�O!�d��&�piB��M7w��Uc�E`F!�䆠lĲlQ'�d�r��um?l�!�M�T���r&�$\���lފ0�!�n�X9�'ǢK��A���L�!���~�0<�FG>a���x!�M�^�!�$/7�
�� �bY�ԊW8?�!�DY�V�,�wc]�<�J�0A�c!���4�
|94�A=:y�<�@�̸u!�$��
8d8�-ס��m�uĞ�5�!�ƌc��4�O�,G��$�TF�$e~!��ڻ�h�	d�����i�p�rR!�dA:��j�a�1o�hc�tJ!�dB�<Tfc&���VN�i4b�^�!�D�$3�p��kC�h�d�p�ߵaa!��C{c���"Q9B�H��Sa�FX!�$�V�0	A�����X���hR!�d_�+�v��ɭKnq�)Z+R!򄘀xk���Ə/aJ�8��	;K!�(0�T��TBf�H��4P!�!Z�vh�`�/3E`�!�M!�d�6?�mh�C�'VR>�#%`��Jcў����p1�"B���j��X�ou�B��1!t�<��݆�P��R�=D C�	�8��h��A:Z�&h1��P�q�C�	� 4�%ŉ]���r�P(z,C�ɮ�jeyU��,Uy��!��O� �C�	�A����ړ%�,Mh�ڍMC�	m�b`�3/�d��`��QTC�)� @�6h��4q<��w�1�D��"O�Ѡj����H��'x��\U"Oΰ��	C�O�Zp�ɘ�h�^I0�"Oعh6Û�i��%H@Y��Hu"OT٨s� l�JX�Ag�\�U�U"O�h�F��8jt�S낶]WDX� "O8C��+�Bv�ϗ!�����	U�O��j��B�A)`�y�@�. ����'�9I�A-+a
M��ψ�T虃	�'�5� ��[����,g���K�'�؉3bfO*/���:�.6x$+�'�&My��E��!��(�^�C	�'%�A!&�,$�͢!�3����'W���I+.�aT�MUL�-Ox�=E��k�9]L ��G�4}��@�-C�!�I	����� %������ށ }!��!B����Nʝ:{�4K��>#s!��+N��4�@�=�J��g"�/!�d1X����n3fð�OO�O�!�$��ji������t/1R��}���Y�T���֍Y�`���҃�!�I^x���6�U�>�y��U
L���S��|�<���
/u�f�X� \�����*�]�<Q�"���4P9� �|"��AT,\�<����)H ��{$f	l�Xg�[�<����`��e1գM>t�08MS�<�)׈N)R,h� �{����PJ�<�1j�1hT"�3"��e^$���DMh<1%�՟K)����HS�Y��L���W-�y���V\�x�@IB^�8+w$�,�y�97V.�ʁ�Eq�:���*�y��]�3ǐ>j{|����#�y"�׫�Jq�@��_2`=���	��y�n[�'����F	*E��5�$��=�y�F����}����&px4`5��"�y�m�	u/p�SÎ�qל��D��yB�05�$ɓ�*�!�bA!e�O��y"�:	�U��D�pMf=�5���y2F�O�š�l��b�z�����y�����
��#�=j�x�������y"��-'�:�@c G4`ЅBd�3�yB�ЧE���2� }0;��KC~T�`�'�ў,R7$U*X�KE=i�p��%LP�<���_�%�@����D�l^�+�(�v�<yQiC�&Ô(���3@�jX��,�k�<9�m�'?�4�9E&�- Jf��`ˑc�<�#i�?#<�[UI �:X���[�<IS�z�<9�@�n���6H}�<��c�jq��#��!q�SF��O�<f����d)B��0a���t�Xu�<9���q������Ͼ~�ʗ\�B�I�N�š�dSe���-��D�JB�	�9 Z����"����R�y"��c�Z-�C#������y����ts�ȓ:*Ȩ�AG��hO��?�� źc���r&��	 �)۰g���<���؇(S|4 �I&u����2�݀'w!���~ �r�����!�KH�@�!��9{�H�r#�T [�.��AKm`!�D��n �k�������,޳Z�!�F"7����@$+����JK';�!�đ(j@�+%!�a��x���%Rq!�$EM��tL%��}���Ɵ?R!��R9&
X�d	�;n!�C��$C!�� 2��Oޏ�%ا␈d�� �"O��+�e7E�"�F���ف"O�C0�@q䁸�"�:���"O��a����6��P8���!c�L�S�"O���VgD�p�pt�䯙��܊�Of�;�S I> 	��K��N����4D����-0p�# ��"�5�.D�����%�z�B�M�2�t�Cql+D�d��ݎ��u@UXg�[�j(D�\�4%�.��j0h*d済���9D��a98RP�D*U���В9D��0u)�aG���򃄉Ђ�;�5�O��t���s�"7-~՛W@�Vp��'�ў�|��.��$.U���s��!��y�<�$n�ds����IՅ9�A1E,s�<�k��< ��E��%~� ƄMD�<���@*!Z<y��ѾT�(����RC�<�"4�b�m !2����'D�<�D��88�p8#!-���u�<��*B&aF�JF��U�Ҕ0p��m�<a�эi�f�@�%?��a�5��m�<��	\�) ���Rn�9e
>�pU+D�<I��m�|13ɷaBެ	u��{�<����J
��㭏3@���� J�x�<	BN�0E����
��%���Z1�Mr�<9��[�g_^q�P%� Q�B�Xo�<�r"ն���I�^�L8�����Rk�<��
;��
���0eޭfaTL�<�c���\kq/��t�)s��G�<���;W
���!��"K���e_L�<� B�:0r��D�y�$IB��K�<�����i��<��*;@����C��[�<)�̗�I�4%��iA�KJ�p�5n�B�<�uc܉iZ^�xs��
��y��A��P��|����$J"x��*�{a�t����gb!��B�ma>�QN�"�`:����!�$Υ�@!DM1j����7A�*e�!�Đ�L����A�d�@��ʰY�!�$zZV H0N�]�F	��
�g�!��I F.Ĺ2�;G��Y �l�!�T����B�B~���d������q��(��I����/0]�f��(3�#W"O|}h�"�.n���ˣN�G"O��3ת\5���Q	B��!��"O2CA��B)�!�W��չD"On�b��E
$����`º�ҭ�f"O,H�ak&ܘ0+�֎�Ds�"O�Tː)M�:�
��Fk_%@�pEh��'�2�|���j���b��A��f�ɺ��1D����Ά�xs���JP2O^5�b:D���L9c/��У�M~�F:A=D��9FLQ�lU� ˓��ehq->D��TΛ�.� ��Ɣ�v��Q�V�)D�� �,���x��S�^�"=��:D�pY&�V8D�B��a��Q�I,D�:pD�9��F�N�/��I�v#,D���A����S	ͼsn��a�+D�X�"���r���JI�ePr�K.D���L^ E\ly��j�H���?D� ��dǿ�*EK��R9?�:�`��3D��hmL3/(TsG�33��ӡ14���Ge	�Z�1�o�i��ey�$E\�<	bl�=:�9K�BU�s#�ei�X�<y�F�t}�h�Ż

���WI�<� ��c�XO��;&��3φ��%"O�4��HV+�p��.H6��uxb"O��7
��l��C����.�8A"O~��&�� ��X-W�}J�@�"Ol�	��K�l�A�B�M1��"O������f<�d#5
�%�t�A"O�AP�bC��ĵb����Xz*�p�"ODZ���/N:� BnJ+6�T<i"O`��AHΚN ��f��Pe��"O��@蒜X萉Մ�7J�<�Z"Ou�!CH����cׂ^�,(�"Oj��c�X��zع�,G>�@��"O�e���3:ΐ�����<�$	�"O����>~x�� ڞX��V"Oȍ�0��)���{Ah�QT�1"O��зό
�>a����NضHyG"O:�X嬈� ��%`di�ةu"O��3!�\�s(.�B��K�:�&�15"O:��T��%�A�6�J~P�XQ"O�xrl����+�
`�{e"OD��fꗘ\�lX@"��#PZ�I�"O��:d�.L\����Z�L�b"On@1�� � 1X�Ц�)`���1"O�U�H�Ӽ��c+)BF�ӥ"OjyabY%��r��J/ ��B"O� ����~=V��`f�s"O���7�
�+�d�f&kZ��I�"O�SWnE6�F����C�8c��ag"O�ᒳ�Җ\Z�����]�hn����"Omڔg��Vt�2��/0X�zd"O���CᏙ4�ڹ9'��x�|��"O�$���1B��!���o�`�"OtpP�o,/��q����$bt�2��'�!�&zװi:��#s*��I���Dw!�D\g ���aW�=�|P厇,Zi!�$�!����HJ4C6�)�Z�a!�dܜR)	݇��@իT�mP!�$W=M��Wn�e�]�
�.C!�$�$z%Q h��N����=�y2቞��z��_X�n�ʥ`I� 3��d-��zq	���x(���,�l�	@�,D���L�D�>]�g�P�,��a/D���q�]d��(5C$4�6�#�d'D���fmG�-bSE�0}%�US�B9D��Ã$Q���A�	Sy�mb-7D���p�"X~m�µO��-b�d5D�0���;3T���`iJ�m[��d9D�a���.X�����:EP�]���;D���*�Dm�=�#��$��8	�,/D����/޻m�&|j�iE�h ��"ag7D����^6��P/��Jz|�`A�5D��s&��g<�|�T钷"�hl�b�4D���TD���������o*�F.6D����%T�9N�4��u�D(D��t��<�5j�@�5���%D���Bo��)�2�P�L¥;K��!�#D�4��W�����T�}0�!D��ӑ��*y&H���S# �|a���"D��pw�7{����G��h��d+D����L �~Ѩ�B&v\L���*D��4�|�6H"��߬h�z5�d)D�$�U)�+p"Y�w��h��Z�1D��i����l�����!8���ick#D�HcL�{���5���vC�q�."D�� ��Q��A2p�X�c	�g!���"O�@su��*fB�Ph�lV�zj�X�"O0xS��P=�v`B�쌓W�M��'�I�2<�]Cŧޜ^���1�Ƥp��C䉑>��)�΁�Dh=��J�#9�B�ɟy�v��& ��l��wL�7�C�I�&��X5���Z�ӓ U�&�C��%���ڰ�Ռ"��5���Fe�C䉼/y����)ϒ{�a+���	~�C�I�)E�(K��ʫ]蚘	��ŪR�B��AM��P� �w4����?��ȓX��a�Ucȓ3�DL�'!'Ȁ�ȓN]%�C�wA�lif�} x��ȓ&�P(����2kR��R"h��Fȅȓ+}��*� �,#WRtJf놊�q��o�A�CX�u&�	ʤ�F�c^���ȓ(��\S�B�LE��9��l�����REhX ��P��4�3lʂ	�����_i4ɘ"��Iލ�6��f�ȓ{9 X�IS�X�� �P�����Qv�0�&.;�qЂG[1�R�ȓK�|�
ϨV�� �HX�%�.��ȓG�[�*�\�R]pʜ1�>|��K̵Sv�� *���$�P�^l���	eR���cH�/��sC��U����;a��Yw�[�#T���n�R��ȓTLdQx�EK+�f��6��w�����E֢0kӄ�	Hʘ��a͹CEZ����tu@�K�h�|���Bb�t�<qr`��%���w��1&.)��LIY�<a6�����3%1_�|@����X���hO�'�х�"�t0
�)=���ȓ"V��`v��n�����#`��(��L�f�
w�Ƅ.�]s%d�B�t$�ȓvޭq ��,��Փ���
�����+$�|���ۨp��r�S'��ȓ}�d�"�N�>^��-��,��@��t�ȓS�2L�a���)���R��T����ȓ?�a�	go\|jp�%N0Ćȓ���D�+&�-�A_�aDꭆȓb�R���G���zqў8�
Շ�h؀yZ�@�	^<D�K ��/'��ke8#�A�?xnzB�.&��-�ȓ)�H��E@�D����'-f�ȓ9�Z-HC(�%z2g.�tw��?��q�zTψ�9��X����"�V����*���)*"���O�	��h��"O(�B5E]L�ҵ��<@{b"O>y�i�.����2Z�P�A"Oz�B��T7lL�<PP��N�`qb�"OthpQL5W�r�r0��%C�~���"O�Y�&�Įc��L��]�z0�"O ��4-��A2�!��jԆ*��Q"O��A ���5�B8�j��P��d:"O����<��9���)����"ODP ��5\����`)9���s"O��í��Z\�\a@훊�L9�4"O�ЗgTt@��!b�7r�`a#�"O�Y0"��/!V�c�1
P�H`�D%LO&�c�kE�e�Ι�E��k|
ݩP"O�Y��Ŕ�k�0�M�Q^��Q"O��#�RS��	��+^�g>*�*f"O<4j�%Q&f���xg�)S1����"OH�����#ؼ��c	�*.r��"O� ͪ�,�"��(�-�|B5qE"O^�A�L+�M�G�J쵃5"OD���"LD*1�"Jԫ%4��q"O��X�-�'m���Y ������"OB=� �$+D�c���6�0���"O�m� ^5;�`��	�B4��&"O��8��A-��ّm�|'�d�g"O�L�'g� :%D�3$lb.IР"O0��0�՞i5P\��X=x(p�"O�#�̙D���J�%K5��iD"O D�u���l�|L(%�A�t��1��"O�Ց4�/�B�ђ��B���"O���1���"�(Lɵ�B�ь԰t"O��C�@իbG2<�'f��d��9sw"O@4�O�ê�jG�3 ���jW"OJ�Չ�+K|�x�`�$T����"O�Y���n�tt��O��4���*OЅ�&�#�B=����@F
�P�'7����J���<�9�W
7Bt���)��	K��i���X'k��ͪ7���yr�R-mA�PC��
^���t���y����= 䏙؆��h���y��Y6^�l�
U�.n:��Zw%]���'�az"��3.�8Ԥ�lj��@���yr�Ll��{c��rb�s���y��ϐU�Aڃ ��Z�|�k�[��y��߶�Z�p��2X���9$L�?�yB@�5 ��R��&��)������y��V���R�#�
H7)%�y�)��
)�*Y��d� ͸�yrH�<ڞi��86�qHPNR��y�� d��q�����RW�V�y�f #s➱�c��J#�Έ�|С�d��hW�:s��	j\�L�ƨZ��!�b��kSD�k��=CĨ�$0�!�D
��V�@e
܈=��)HPI�6&!��y���QF�9.��p���T�!�D��T���+F�ׁP*�9StHҒ�!��j�{c���^���P��!���?8�nBp"W �p��3�]8mp!�DT�(ȸ�':�� 
���<b!�d�v���k�n�r��UQ��'F!�W�^2=(3��G�������%M_!��A�h�+t C�~�� �F�4�!�dː6�fu�e��
�v�bߧe!��X'`�Y[���k>��Bْz�!�d0Y���c��&TQ�!�`7[Z!�$�U�xIb!]�?�p�Wo�hJ!��CI:F��%�#6D��9�Ϟ�2A!�DQ\C�I�1��HAh��.Q�[�!�d�{�09(��ˡ(����/L�!���-*Ԍ��NH�w=hIA�.	�!�d	�K��xƃ[B�}�!��}!��0w+T��@OE+B��e�_m!�d�H�<Hf@�>{$��1V/�P!�����c�ѱ#@tX�Ue�w!�DA�a`%(��İq�P����
�!�$��=�$]���;7�"��j�}�!��ĊD��4$+K,�L�3�I#|!�d�v���ԅS��U�5B�Yh!򄌞!�8Aq�a�6z�-�↪?e!�>'��ɂRh���IJ!�;Z�5��
0$5��.�Q��'R��K�.H��	$��1������ z��@�� 6���*H,x(�"O>��e-��E��ŔIUK�"O0욆�M;7(8���%��bp#��'��x}����fQ5�l@��D�!�Y�:�n�և95�~��F'ȂK�!���5</֥`4���l�@���!�䓦8��}`����M�dɶ.-B�ɳ2�j�c5#Ȇ (^)1�ǈU8�O"���вh%^�C�'E4����'-�ў�ባ$F�J!�ҽ
�.�1��
�" �C�I�X���b"@(d\��b
�U�C�	��b��0��+g&�)"���C䉼
�����B�)f|�p�G���C�	3^�V}`+J2C�a�G&ˬC�	3Ƞ��& �%?Ԩє�ƌRo2�OV���J��$�0H�O�����U�!��`�)�pI�/"g��3ŏY�!��R���1&,�)����G/�1�!��Gl�<�B���24��&.�!�D��b��8�t2<v�5 C��g�!�
2(�긒7*�cFpp��Rm�!����Q"�@��`�DPe$K~�!������JB;I:zGd^�[�!�ĞJ),-�qA�iX���TP�!���1�|��F.�R�	E�u�!��'��X�t��`Zh����@�s�!�cRQZ���.JVf�J����fS!���V�=Z�� 1C�u�6!þ!��Q�R��1���*'`�@�&`!��LO�V	���R"D�����nT�5f!�D�oUB�i���*W������MJ!�Z�L�VNl�fT�cj�S9!�0�T��eLMˢ�ٰ�	�pJ!�$�s��8 "��.1=!���m���F�8�1k� m�&"O`��!,|��$�]Y���Z�ODk�$ؠC�@�;CkڴW �a"�ID��K�	ʪ%ۘ�2B���t�3O?D�ܙ�&Fs�� 䒒X3��꤃<D�����Zq�`��JѬ�<L
S�?D�Th���!�sgA� ^u�IC� D���C��c�8 ⃞4&Q�q8��?D� #@�._2t!���[�.�HZ��>�O(�MuB��֢�	�"��Q�*���@����@Ԉ4)�	 ���(	~��]�$A:D��93�Ѧ+�b��f�^QI��C	9D�옃	��/z�E�D�R02h*+D���C�,o���C/	x��J$@)D�,�bw<!��LM;R�2Y�d%D�*fo�;<����ʋa�@�)6o$�숟�4��o�	[���Po[?jL���'�ў"~���1{�$]Q���"j���DFT��y��&$|5�t�(_�E������y�G��)0���`(N{��F��y���3_M,�$�O6A��a&��yb��o݆ac�*��,;��	��y�L��4*pƃ(����4��y�H�3ll��0ņ����D��m�<a�h����k���RcL�U�<�����\t���́�)��a��!WU�<1���#����O�>b��� �T�<��.�[�&�i�����P��P�<Ƅ�)|њ9%��=�rM�B!O�<q�D��f�~�`��_�D����@�K�<� �pCЯ�
|��Ԋ� %%�
"O9'N T��5�&!N)��"OP���T)2��1�C�/U�ИR�"O�����4DDD`��L�����1"O`�JF��Բ0���ǎޮy�W"OZXS��պ+̝�	��(7 �	�'�e�T*٪SS�Ԉ$���bR�=�'8tla��P�%�f��W��
�'��C`H �R_�����f?XlP	�'�iX3ǆ�Os�h�b�H	�'�:99�O�/+ ����F ��m�	�'��(!�U�[��ب�K�����j	�'l0Ĩ��^*;�Y�����.R�s�'�$��Ơ�M�\��+R�/�x	�'ddU��$P��%Q5j#D0����'$�(Xf#��聤*�;B����'<�����	�F� \9���#7�I��'ⴥk��@�YE���`^0�^\��'���Wh,��1�k.N�1�'�v�0�넑@�ʹ��HֻD�$��'=�IȐ�= �\5Q���
�lR�'d P��v��� ��NrT�
�'���Ǐ��E� i��BI%t����'����b�"q��-�6�N�U����'�,D
\� �F�8��H�L�&��'��� ��_�a$EK���>6�k�'�8|���	S���eH��"�(�'/�Q�SDH閕��N��%��M	�'����Ddh�͈2�G�Gp�<0L>����'Q1O�L0����c���8�v"O
ЋgMN
�+�,����#"O��R��Zf�<���U"s��m5"O �����B�̕Q$_=�x��G"O�$"W�	65xV��#L9Mx*"O�%�f��;`��"�UgE��P"O�h�#)V�/ezpc7���P"O\]R�/Y+[�Eޥe^�"���)�S��ě&E��p�ڔOY�Jœr�!��%i^ j%J�o:�0!��%j!�֋Tf<\q���
�Z)	Ţ��TP!�K�Jd�t�qρM��઒�9m!�䈥��	3�*ׯ�`�!V��F�!�$ �F��=�f�\�F�<l�W�7U�'�ў�>�h�(/M��zFc?/K QzU�(D��[�Lяn<���/`c�苐�%D��bg�ǡ.���zŬ�p� &`'D�l�g��%i<�pg�#���#�9D����.X�9i#�̃P�ͪ�e8D�|�� ˗B���
F��c��V�-�!�ğ�C�|�;"��;��aw��~�'�ў�>q:�eZ�=�n1����)��	gb=D�(�3C]9'D�ԃō8
jZ|�1�:D��2��ڤ"���FH�8x�L�a�8D��+���?�f� �X��2T���6D�4�%�I�̀A�!F��l��?D���m\�f�*��VfՌ ?�Z�?D�����ԙR�i��G�"Y��`R�)�O���0�O��9�Ņ&`<���M
��"O�Qȗ��xP���@$ߞ���(1"OTT`!�Z�,�� 4*�>4�P�0&"OZ�h��>R�������iU��`"O5)C ��^lz ���i�Z!�R"O�ˡn͍O��u�P��V��q"�"OH9��0�P��!,l.z�P�"O� �5�ń��8�:4h�H�KfLq�"Oh1�UC�����Y��p"O$���hC�(@�f�u^(��R"O2������dF����P1m�$��"O�V�<.�aC2X�,#T"OPU�%d�@��K@��	@L�$�e"O�����;oQ���ȵX*�� "O��Kߊv<�`{'�ǋ=$I�"O6�c�-N�^�nq��H �Č�F�|��'��P2j��:���7��r�p��'��pJ6��97L��D�g��}�'N��i�C�f�j')O�b̌X
�'�t�"��^>vX�f�ߟ*.���	�')�����t�L����.q榱�"O<�QWI�d̰��K����v�'�1O$YQ�M�.� �4ǋ)}� AS"O�t�w�P#I�Ա���\��,��"O�l�B��=�D�Bd��q���"O�0�c!G1*��@��#Ъ�.�y"j�.�ZL!%��3_k�����y���/Lh��d��_�4#�����D7ړ�O��8pC_&z��3��3o�hݡ�O �6`�8h��̑;/�M���,D���E����<�H���>P��!:�f5D�x[h/f�r�r�k�{�f��v)2D�<�OPl��e�}AD����=D���@^+p!���s�"{I�\�w!D�h�!
W���v��6g�� �J?D� �˝2��A�"����1�r�<D���E��u
 �9p�z �K;D��
�)�/BFy�&���rX3g;D��0W
Җ9��%��J"-5Lp��=D�H�f�ڛ7c��GN�#k�h�j�.D���a�X�($�m
a��0sE��&D������!c�lP�`d�%�%ZѢ�OܓO��S�g�L�sy,u��j������HQ��ȓx�8A�+°+�����@����ȓ+��#cÞk���E�މ'�P��ȓB������O�D�X��Yoل�>.�I�e"�a��IyS%��6��Q��\:�sС����Á� %|�I��Ot��s��֌7<�j�"G� 7�u�ȓ'0(�V�R==�I��̓��l�ȓ=6���T�%(���p�mj �ȓq���͜�b����1��y�ȓF�\��c��ic� � �O�U�����Z
B�[�N���ܡvb4P�~<�ȓl"L=��P<c�E	�\�pAl��wHXȹ��&���W�G5_9A�?9���0<�$e�$F�!W�]�N�<��[�*����v��R�@J�ɎM�<y���Q=%XM� [H�kD��E�<Y��S:/�8§�`���LTD�<)�
�°�8DՍ.�hy�u�<A��K�3��s�rNh��Є�o�<��̅�2Eƌ���+/�����A�<�"J�F@p+�lG0]9Z�b�#�@�<�R.Ei�����O& @�碒h�<Y"]B04��%�'�p����b�<i��_���ÓF	�3��8B�$�\�<�%Ы)d��S`�D���|�`�[�<�"F�0H��U��T{�4  c[R�<�ЁE�~1ܵ�.�!S�E��O�<)7'�8[KUk�K�UO�=��h�U�<� jE�'�@�(�J�O���+T"O.$���"xLY��o�1x�̛"Ot��)8$h�07�bWT��C"O*DJί���\;%B"�p"O�Iacʰ#B�d���
>92��S"O����H�*Nnz�����LlP"O*��!��&�E"�N�u�pcp"O=��ǒo�����Z�ah��۱"O��� ���/-���\9n����"O�m8�%R+1C*���b�=U�t��"Otൂ��J�z��#���x����S"O � ��+@c��YEC�)1B�$"O���L���X���"#~��5�v"OI�#"�f)�����e"OfEj�!�VnQ�3H�M�<���"O�=c���%�rE�V��'���)�"O^ȣ�ɏ�9R:�+bn��� S"O�m���2��`�D��B��D9�"O�R��T�U!V�:���19����"O`cWN_(6@���eŝ�S �5u"O�}��	��),�7f�X���R�"O�˶��A�qbUd	=�͐"O�pB�a=YN���"	�9�����"O�p��"M\&�U��,"�Xx��"O�1!Q΄�%ny��b�z���"O�X��d��	VR	R��
�v���Y�"OLP#�X$/� �15�U8=i�P"O�蚷e s�u��&V	'|uiD"O���g�IƌHؒƁ- �4�c"O��m�qu65RP�:���"Od�%��D-P&e¹x�!"O,�C�ѻ{���r�dO�Gb�`"O�Q[ׂ�!��4Q'Ç�T!"O4�)�.�w����4E:X�S�"O�����r=ĤK��#���"Otx2��:�n�r��['g��@K�"Ox�%�O�o�Z�G)܈3��{�"O��Bs@A�:�.�۰�B9a��D�v"O�����!d�x� p�1'���`D"Ot��� 49<@S2P�`����"O0,"����T�Bk��	`z��R"OB�れӝn.�=ՆJPI�l�a"O�CC�=9���̘ "��w"O���h�U�H�i��ĉyh<�("Or�#
� w������:w��ʁ"O�	8b��!H�(c�����bW"O�U�ߙ>����U�R� �@�"O(�`�n��VN%�#�(�@	�1"O@9�"�94��/ߪT�D"O��u���rp�$H�7�(���"O� �Ed�����邩W8��U�4"Oҡ���E@4J8
����A�މP�"O
��ԫZ�b�������s���y�3[��@�/��9S��Z�4C�I�~�5H%n���Uq&���:B��2Kb���׭�,^�=^bЁQ�"Op����9���hs�� jϔU��"O4p�ve\��4��d�A>��!)�"O�z'O�
Q� �0�哋e�ƴ)�"Of��A�cNN�1���S����'"O�e�'�� ���s�ۨ�~��2"OV��/��,��D�M�lt�9�"O��{�䖌Jelāc,9fh�@Q�"O��"4�+������4Q�1�"O� T`� �T�QF�}e�L�`����"Or4��H�v�
�*�"?x��y�P"Oظ�ī��e�xs��Ѝl��P�U"O��g�҂�.��go��Q��C�"O��P���
�z�r�8R�y�b"OfmZ5�ŁJN�j�Ob<E�4"O�q�@��J�N@G��E@!"O�i� EXN~%��c��g֘��"O�=A�m��<��❖9���Q�"O�(�,�.\
�7A�/���a"O(�p������8��X T����"Ot ;a�	Z/F�HōZ7!��U��"O�Ȣ�-�9$��""�](.����U"O�Ѐ�hI._Ϭ�Al0�rQ"O��DD˖gi�왕�رa��b"OKE�����EIQ5BIԬ���y�"��#{Z��1�̊
�FT�����y҇���8g'�nl�4k�k]�y����|�T�ʚ��ś���yR�F?[g�غ��A�e����EL��ybDSl�\5�a��-X8�EI����y��9oX @b'��9��e����y��+^%��95�/��$�#o���y�$�E�ܼ)d�\�'�l0ٳgG��yb_�+� y�^�7�q��T��y⦎z�0��bޟ8ʘ��"�#�y�I�.9/ |����'}J�j�CF$�y�A�>=�ı�@K�)��Б����y�	�t��E:EdJ�
�HjE��4�y����<�;���<}�L��T�^�y�93q܅�Q�sv0�'���yC��Yp��C��q����Q,��yr _#[)FJV�O r�@y��.Z3�y�!�D^XT�V�9qK�3U*Q��y��לP�T�Z5�B3m.�ش	���y�jW�0(A�ĆD��b͠䈚��y�	a2l@Ӈ�*~)VDq�U��yҪ^��V¦��o,P��#�ۓ�ybD��){�T�gя<�p0��S��yb!B�|�r�X)64H0q���Py��/~<�A4�,��{%��O�<Ѷ�P9���-Ď�y&'TI�<��@�I����!�68,��eSo�<�g���*䉕g�6v�A�Yd�<�7$���8 )��74^�����[�<٠��3�L�@o4X�����QM�<�Qh	)pX��ӫ�z	>�{$e�r�<A]%K��KpC�ِ֘vGGm�<�0�U�=1��"�/f0�eΊl�<�B�މK���Ӕ�Q)T��DWl�e�<iC ]3��c�e�=}���C���`�<���$����j�H2��%HAv�<��'�:b}4� d+Ǎ��q�	p�<q�@Be(��R������A�<��n*5D��燋c�E��&@�<�gغQ2����R�>�n@�� �C�<�#šVm�yh&e
=�HI��OA�<���W�� A��e\viE�s�<���B>88�d{aP�e����m�<� ���ɥ͊g`�0%j�<�b���`��p���?a��3��Az�<A5��t+'O�`<��D�a�<�P�RD%*�:�C9n�|K�CZ�<�FC��!�FCA:5Vl�a�Y�<� y�hǠz\��CM��u ��"O�l2�֑N�޹R�B
5~)Ӥ"O6-��/H�f��M��S��q"O���K�)qzTI!����YB"O�l����`͌�q�M# �M�r"OhAf��	/�iX�e˨ �x��"O��H�lU�=Tz(Ȇ���|@��"O�т��£p<�u������D"ON�)�F�	(�aI�C??��ȣ�"O>���/Q�0�PF"���P���"O���(As���ǚjJ!w"Oj]���<n"^��#��+���"Ol���L��U��M��Q� ;"O8�3��ņtX����ڈ �$�i�"O-� ɥ(�`:���t�Z�B@"O&%p��J�QMb�0�@�3r�iQ"O�L��
�;�x3�JGw���"Ol��f�(H쥀�À.E N-��"OJ�`Э�"Z��ڡ��S�$t��"O��b��Pu�8��0�Q���@!"O��9���:IK:���՞um��C"O�Q
S�ڂ0,�9�m� ��""O����A�JQ�$���j4���"OV���λ�i�#C�9�f�b�"O4m�┯���F�R"%��]2�"O�Y��h�8����*셂u"O�A�p%ӡl0޽AD���I}6��"ODa�!�*C:� ��#"ql���"O:2uN�c�lArDς�h\����"OP�1"Y�un֥X�D�(b�L��"O���4�׵'���S���5]�L�A*O�`��͗f X�A�$L#� {�'>9%�K��i�5AD�����'�D����˞��qc�͜�}��В�'�H;D�N%'yJ�ʕCT�'h5�'*R����:_�Q�	�S<H�'�
�3&!FL:��O)Oo���'i�X� �B�d����Jy`���'�f{��'"3�	3�L�޹b�'�x5$E+d�1B��=~		��'�@E���1�8L�T�s�(P�'��P�SJ��X���E_�b�\�
�'4�T��ΎH���jN�S#�|	�'նE���������>I�=C�'���b")ƴ&�Z�Ђ,͌7"�`�
�'3��1�lΠ�
ݸ��-y�!�	�'�h�P�Ý={��D0�FӶ|=�@:�'���)�n"}�pE��`Fzm����'��I�,ߘ4���Ba�k�r�+�'v�� ��:�pA�WJG�^�r;�'��A�� V�4����U'@�J����?�'g6N���E�2��|��M��&��}�ȓx��( 5׬oM��#�K�Y��y��t�7e�D�|���@�w�� �ȓGE~ȃ#�[�l�����'|C*�ȓ*a@a W��pˇ̿u�ի/.�O��'�r� e:�(�9�/F&o����'��E	�ሢl耒�S�`�l8��'2��("�B�(�q��L2�dZ�'�>t�
�;.��C�M�A��!	�'o������T	�2��87Vт
���'`�mZU@G<$<�%�5* ��	�'=���t�Ŧ,D +2K����y��ɬ�ē@;�p�k�a$�D�����S�? ҍ�C�3��y�rd��9�fp�t�	"�HO��Rz��b�(J�xcO�@�lB��2_.��B]�B�fp�sL�Q���8�S�O�rh��n��9�HL��+D;U(�z��'��	 �R�!�ǫjTU��*S,:5��D+�,Ȣ�	l�� �(��b}B!�+<O�"<1S�W�z�0�(�cZ��%�G��G�<y��R�� � ��98�KF WF�IU���O��m�e�����ࡇ�s"쐪�'��(PQ��A'��)A$�H���}2
:LOֈ�L�)]B��F�M�v�]�&"ODHӲ[�Y�����'%�< `"Oz�;RJ�a)EY뜐���'#�dY��[ "T�}H ��+mp�!�פ9D�Gbήt�0���o�-2��� �6D�pR�	�34�sC�	7,���,4D����jE)Pg�t���TX�����2D���RJ��A�8УR �?8H9Gf<D�`[�f��8���z��N�"�J�a�4D�4�S @t�`�a�/λn�=���&D�t0R`�&�����B4�Ru7�!D��9JSr��Ը���e����4D���E`�2H��q$	ͯ8�����,D���DDK&V��H)��J3/��(�/D�4y�뉝�֑�#��r�rx:�%-D�ĻW��Q-4��ƁUs�p�` -D�HQe����k��
�s\��+,D��j��ӌv �L+CO�G(|�-D�,;0Ċ+�z�
&��is>�*D���¶(�F�04I�N�6����#D��ь޲3u�9۳��KZ�@�5�%D�P�,@�b<R��֋ĜI��S�'%D�XA��;+	����Æ$�Z�дh�5��'��z�Ǯ	���� ���9�^�;ና�y�L��o�dY��+��Ё��:���9�O�ccGC+8�&`ϐy:��S��Ic��O�O�\x�!�ICXP<S����L� p�'�.x���
Y�@mK���nI2�s�y��'��O1�"C�䛬��xP$��L�JuP�"O�Xr�����q���re6l&�S��yr%.Y�p�խ޲*�:�&�.��<	�O��'��Qj��ܚ � ���`W�x}��	�'MDj��\�N�9�/�kd���J>1������b,c�Ğ$]X��cR!�=�.@$"OR5ca;<J���W�h'�Ȩ��	w~��d���np�`#Jf�NL��K��!���:6�^U��%��DfJ�
^�̆ē	�f����;D��#6��82����I4��>�tgBҊ(ŋL�0�ʝ[��+�!�*L/�-˓DV5�������5ўl��	�SȚXqeb٦ R%��!��p>�B�I},�l����-��<�5��S/�IT��MʟHO���z���<	��<H�C#d!�T7Wv�)��&]�<����4fP�I{���SC�;v%�AL�@Qa)lOT7MH���䔣x"ᑲL�bQ���5i�#S.!�$��<L`�r"�W$ ��(�s��+�'^�'��Ļ_�u���G�$���u%�Ii�a����<���]�t8�I��[��
m��K�<�'
8�j��5`D<K/`i���p�<1��\�(�\91�G4�r�c��A�<9����(HrU�;oXH���y�!��h}�A�4��V9�;��Î.�!��A>o�ta:t#Tf��Y!E��?-qOrb��G�� ,<��Z�M���A�O�{CJ<`�"O�����J̸��=v:���C"ON���K�0Z\�1bO�i>�,"�"Oh��0�Q�D` [����c0P��"Ox�A�m	/L�0�s@�� H���"O�-��,J��*�9�f@�[%"O~U�SO�L0{"&�7��&"O�RecˤRgISׄF�I"�Yc"O���0G!�tl�`��/Y粹ط"OlA8�,�7��,Cb�a�*-;�"O���񥝤0�^�)G�_T��X�"O�<�m--j�3��l<>m��"O�arf�ĄR<\A��A�,�xAu"O��!���2�e���H��"Oz�Aa�?i#Ҡ��	%��"O�Dp���,/,j8
�G�5��j�x��'F�z��ɳb�^
'*�-'�ճ�����>��OV��"RU&���c@*4��[���Ħ%��I}srɨ�ƍ�*��a��˸]�HC�	.$�E�� �M#�X� ]�y�t��4�<�d�+G�2���lF$B7�UA� D���fL�%n�2�JD"i���"�J D����nU�n����Ai�ؠRp�(���+��y�$P��scʆz��z�4�y2��p��#�����!�@��y���*��1�ɔ5b��l�����<ib*4�ɲ6ӸT:� k�|$k�'�(�����'>�y"`�2
���DDZT	��I�Tw���a�"��ӆ`8�)D�[��ӋR�����
��mP���H(�ə�yB�0#��6zZ8p���
wiRX
��1B����q.�e�g��fn���M�($1!��I� �VD�F�)��J�|ay®F��T"��s5n�fX㧐�=��P�']ў�|"�h[�8-�H� *��O㦄"fcy}F�J�'���i�	, C�tR�bN�<2�x+�SO���O����8�*Ѱ�AՍ�M��9fщ'K���\�~*��u�b�1�Q�NI&|o<�"O�?��x��>�rD6j�B݌���M�,�Q�F�dM����a�-�i����gZ��y��Ӟ\��P䄛��ZD��6�y⫌"QI~Tc�Ɯ��V�{����ē�hO�I/}2B_8R���!$����xQ��y"���,ږ���r 0�N�#��'�r�I|�Ş$�laU�� ���2�TL�ȓ_?h��Ĺj��;�c ����'����O.��D���x8uj�1%8��wD0_�!��CX�A�W)+*�I9aM��rC�	
0Hr��v�q�TH[��I-rC�	�1��}wK�f^0��`�ط��B��#{i�u-��jpA�$fڂB䉞.0���ò3 ������P�ZB�Ɉ-[���n��I'��S�G�#a��C�I%2��lX��Q W`�%�5鈕w�B���)�gA�U�T����& &B�I�Dv�I���81!�����vLC��&:�n<H��ęb���+��.�lB��.� �mY$΀��r�R9Q��B�ɪ* �a@�V���#`�ΔԖC�ɋ� S%�f�8DK���;.�B�.lK�5���ڙ!&r��"��B�ɹ{=P4�9�Ι�7��KJ�C�	�"�&]35.�&�=����<<�jB�	Yt����K�C|ID�T�A�^B�)� \�@���@���#�	"����!"Oh9����/�����&΄#g�у�"O��QB��(Rr��4�8q��Y�s"O�%!���w$�� �X�/E��G"O� �Ĥ՜dh��vL��z/*��e"O�@����<F�A�ceޗ^��Qc"O�� �Q$^�,)�m%Yʶa�A"O��S&͌O���	�L�o�&�'"O��b�KE%=���:�j҂G���q�"O~�`�_�)C43)� xT�1�"OD�IF�W�UB�qh�7ns�0�"O9҉��J8�dȥd{,$إ"O(%�!l�/ LD$�í��Nu�E"O}c�c�U������ʋ�a�T"O6 smա1� "ՠ��fd(�A"O0��f��
҅���"�r���"O�\��e@�[�&��U�\�O�D�@"OԄ��#�)tT{�Jg�d�G"O$��,����S���78��U���'�y�ԉ֋b\���>`/V$��.yJ�2�'Z�4�'([��a�� U��dZ
�')lM����P���Q!�W�%7�l+
�'��0O3"�MSP͋�.�M�	�'��"a_6\���Xp%΍ia����'v��p��Y�0ޮ���*�&j��$��'��EoH�;���1n� U}�D��'��h��=I���&VY�u�
�'I\HA��F�3�8x�a'J�W��[�'��0��°+J4��R"� J�P���'9�i��h�$oa�x���pUP���'����Ad.b��q9&�N�r�\��'6ܝ��D�y�J�
��d��,�
�'� �"���\1X�' �t	<#
�'[���#��N]x��VZHxщ�'g�}�왒��M���ʊC�����'�@�a�Ymf81���0z�D�'Vݱ���u4΄��2�9Z�'*�0�A�])3E�V&*��2
�'7��+Vn ~�)z�ʅI^�D�	�'������.'HN}b��8�u�	�'��Uyg�\9�3i��)�`���'�r��*"Î�p2l�7�����'Ej�rw�H�p񄉋H
Va�pY�'�V��R��Τ�S�^�V�H`
�'hx��Ύ>T�� ���[l �(
�'	"d��f6�Xm����B
�'~��`�`A�]��`1n�[D�		�'����G�̈J�
ЂL!�*���'~b�����t5NP���	�*-��'����������Yd�&I]y�'�y��ʮXiV���f��6���'v�,� a� 9-bĉӤ[%�����'��l��P+v�mqso�-hϴt�'�65�fh����ч��e9�1�'X��2��.&�����#D/�D
���+I*N-���!�U�##D�0��N�o!p9B��'qʘQ�"'D��ل�W�6@��)˵L��t��3D��IP�<a�ry�g��YYH�R�-D�8R��@�TS��؆�ըW�L!��=D�X�O+ЈC�l��"쀤2��?D�TGBYRu�,3D���ܠC��=D���N9I����Ԍ�/;gĄ�=D�|!�L�[�±
Mr?�bu�$D�� ���e�K�nU��;0�Pu|���"O�ݪrn��G�~]������G"O���tؽ&���x� �ll��"ObL`WBŨo.�mvl�
/r�'"O)k�e����$M	nzⓟ��OȚ'1qO>��ĶCs��(fC+2.�Ɂ�'T� �an@+�-�b����� |rƞ=��0��'X�����S:ib��;H������x�pC3������E@,�Q1��A"4�N���o-�O��a�O�[pܬ�E ɐK�䢁��+|���Cf�. J�O��wHWn��!G��D��'�I��ƒ�L���[�SZ$�#�O p��9����J�"}z5LΉt��L80�߷rV`8P��m�<yCBĥs�ZT�%&��j+���dEL���� ]�B���K��g����[.#S2���`��K����ɂV �����Kr��+��וH����Β�n?$�Qv��3_V ��$�X\I��5fvu
�V�V����B�J-¸i�든l���J��i�!R6��XX^ay���#]XM�p�4D��;w�D���<9���,S�� �E�>��DI0Mxh��UgP- �ȍ�S�RJH>��R��,Yz���f
�}ب�9(2D�,����b���a��5����ޣ+� 4�j��W�V\x3A�=b�쓟RX$�xb1cU�<xe��4i�h��I<�|r#��J&D�J�Z�>����)ޡ�$",����E.C<�:��	)$�d�;����:�y�_����(.<O
��N�{�&ԹȎ�&�b��$��*�0i��M'Ģ	��#����xC�(2|V�Sc��((-r��9��+ 9B���;O: �b���87U�c?��JD�:�޴+'�_q�h�z��=D��!���WJ�p0��I2pA6�[�K��^L d�P�($�<G�Jc?�ODܻV�T ��"��#�`��O����-  �X�m��;�a[N���� ��hs0�6B�}:��4Oz�JT�1Q6@a7cO�M�Pqb��'b�|��nG1�L���܍Y��ȅm�%�dq⨀v������]ڢ!Y
��G��e��� ��ؕ��A��&�|[�ߪ,�G(@��IXGဌ"�����5�4d٨)�2$;��h�GĪ�yr+�Z�����v&�x&�����ȕI�r����R�e������19c��	�c����*���
U�v��C�	76�*]����2L�~y���H���R5l�� �tj�r�ػt Q�~� Eӎ���2,4��Ї��28<4I$EayR�ϭajP0���N��c�eFĂ3C��z��G!�6����c6F� cD9�O*)[ ǒ�@pzx8$ǚ0#����$�|���!���A�� x"�!t�D~�r�?�����p�Th �P��8���!D�����c�<�(���"`�zd+�?l�pX�,�@d��JҠG�E�,�?�x�H�<��$X
T"X�V�Z5JW4-)�J�b�<ْɯ5.�*���X�n�HS�!)l���7�ï7k����o�09Ң��n�'P��UkV�1d>pX`@�Q�<H
ӓ2> ��)\��B��VA*�b�t��ѓ�	�$�&PYeDB)5�tH���5&J���S�P��E�⯆*?ڔ�D�w#UoO�%qR�_r��<�篊���ӹD�l�:��Û>���K�ŖF;�C�ɯC>�M�ů�(Qf��P�C��"�*�c�X�~�e��t: �!"�g?I��?i�)�N֘@�ҟLPhB�ɪW�����T�cg�p����+Mh�I(>��3��'��H�Ӄ�*FL@"�D� Nh�� Ll�p�kӂ�3���y��H�\�@�62�!�'Њ��҉؊/@�J��ܑ�@��jA�yE�T���J8�� z`��L��y�c�v�|���;�Pp�f�܂:� H�,G�iK6�;H�"~��������jļt!��XUU\.B�ɮ6��قDd�j�<��vj�y�F��$ ��|�E�ԷQ�azr��<�0R��3~�N0c� �p>)�l� l�u�T�Ǧk��{'�1l�[U�B�m�d��'��0Zr��3ZZT������2��)���Kq��:�fԲX^P��}�Cg��S��l�����l����DH�<i���xFqɓ�zLA�r*��&f,ڷ��9�����Tt?E��u�:-(&�^�Vի���1 ?n���S�? D��r�e���A.��M$����O����w Dr�D��0<�N�i�Rq N�P%�xH4	�X8������Cd���3�=ue�2�`Q�q���j2jL�Tdx�{wO�u����"�l��a�I�5ᐨ($�	! ���BS��V�n� ��dG�%QϦ�s��{�ࡳ�Э�y2�7<	�-� &�hܦ�uf7�?ɳ@�3	jz��f�����sӔQ�@j2 ����
͑-�)c
�'�F�s��\HՌ�CF��+���H����3R81Y�'��|qg�Y�*�P �냍��p;��$�x˃%2�ک���b4JeK!΄3$��	c�=��(SJ���b�L�Q��7�&�R@����ϖ��O�4kt�D�Q�@������!��'�%��h�S���g)�/sվM�,ONQ����ΓOQ>���L4=|���V�Y���qBA-D�|3�Ð�=�r�@�H�J�WJ�w�II�@� 
6�3扏���p O�c�LiA	�}�@��$
�VR�qޱؤG@�eW���"|��1�=�O��2��8�\�xP��/�<{7Q�(c1��)�8�'Q¥��Ċ�4�&>�
p�� d��#�V�M͘<@5D����[5y�m�F�҃q�t�[��_}R͋�'���c��OE(-0g�9��d��(qx��V�r��{��
�2y�~R��j����a
�e����Ѷ`6ީ�˟�L=@A�O��QΜ�^�����P _���4
�c�f�d�dTQ���j�I��Up���Q?�R��S��I��?h�¥/[�ǐ�n�g�*��$�/7/R�ҴF��� ��E�L/7�d�'6�T=��iήa~�I�V�$�A�j�%J}�O�ƴp4��Y<x��N��0i
�'� tX�`Ѩ8΀����j�ll��J���i fzu
q��#ZL��L�;����I�>!��>b�t���oJ(]�y�Gi�L��X�B��XR鏓3��V	�eCx	�n��� Y��T�(��؆v�pD҃	|d��ގ ָ�&ŋ��O�P���Э*��8"ͻ<i"A��L���Â�I'lLS@l�8(`Ѐ�4�x�@݀ou�����Svu����x��/^)�����[Uy���ή`�Nj�J\l:5: (\�!�d4eQP !��1q�����bS�(�d�'�d���ͅ'xUl��O����.&v������ϱU����'�����ΛH#��f��KzX@T�N�!����$OJ��c�+:��iG� 2Hpy3�"O�� �T�<�T�P��X13@�@��"O:�G��F��B�tޘ�6"O䐊V΂��L�Q�#�7�����"O*�4�P�>���iҢį`r��PP��K�����OJTڧ)ƣ*�
uS�ֿ\�¹�A"O���e^;"-�I"��3�TE�F8O��"߅#p.���F�<�a;��m��r_�y��6^l�k ��<4h7-�����c��Ui�t�Š"~!�)[�]����?��<��`�]�O��W�(9���	��7S�jG�?E؝ڵ�ʧ|_!��<�^	�q��I�Lܡ��P;��m�si��@B��O��}�Pa����)�,#እ��cƯm�x�ȓE����@�uS.BMJE   �I��JP)��� "�a{��ɬX՚�W#ʤo�2�c$ق��=����7J����i�Z�*$�ڎe��4⁤mw�A�"O<�V�3\��BP�Ia���d��#�"(6m�"�H��h9`,ݢ1�Hj"/J�E
ր1�"O��; @��]�%R�O��F���Iq��� z��u�b��"�g?іŌ>2\pC� T2�;tK�F�<�FK�i"��9��P(�&'��<��!i���ߓҴ  !`�+��AV�L�]��	y81f1O�,X�"�80�|��8 ���"O�P�S��v��H��3o^(! "O��ˊ�+��+s%A4!F�"Ot ��$d�$4����~%P�X�"O��cTs�ё�d�v�
U�&"O4+�h�}�r��$�o �IQ"O� <�
V��R�:�
�@��"Ox����ЬD����� (q��R0"O�����)f����a�ǜG^\�w"O,��aB�E�j@#�l��7"O@y�Gț_H��X�cp&�"'"O�e�VEB�z;B=���M�8q"O�a���S�rz�aU��h����V"O(����H�<V�T c�<U��2�"O�ᆉ"Q�]��?~�k�"O �kD���]m�|�ק�w��v"O�0{P��UT��
0�[ (q���@"Oj��f) $��}�����?J,!��"O舻���[�&�@@�\�H	{G"O���B��I�ŀQ,e�^5c�"OR,���8~Ԍi�Lôk�@PA0"O��S���sh �1e�u�L���"O��U��V�
t��k�
d�:��"O��J���
������U.���""O�t���+E���g
I���"Ot��F�{8~����Y�����"O��Ȇ��R�m{%�W�d��ݺ@"O��BW�P	2��$@oJP��m@�"O:��hڨ|����@�%?�L�s"OR#�iI"t
zI9pσ���c"Ox]�0�V�q3>Ay��@�40"�"O@t�f* �O9}����B�t,x�*O8�SS���u�4�;�nL'Ds���'�Xxy�D3â��0�[�< ��'�j���V
>2X����FQRX�'���T�guԙr�Iʊ
P,lR�'�d �ƛ��t)�,�';�L��'�py�/[,�蕫e�[0{5pa
�'an���^��*e+e �-��p�	�'����BŇh�>�J��˖K7���	�'n��5�L*�j��j'D��U�	�'hTp 䆔�N�k�ȕ*��	�	�'^8�z�*��G�J4S�MWt�Pc	�'��@�A�9j�(�cC^�{�Fl �'�ZyX۹z�"I�'�z���2�'�,�G��D6�H���],,�6���'�|)C��?&��(�`ѣ
��H
�'5v��ǝ6K9D|�3ץv0 c�'�8 �Wl,VrY)3Nձ%�ڭs�'����E��~��Qp������'�(�R�A �|�`q�G�E�2`��'��h2�H�L�:i� �Ǫ�҄Q�'䤋R��Sl�H���K�J58!�''tebPcM
VN���Vj��
�'$$�ql&N)�a	�P����'$�h���9xܨ���N|p@{�'NE�.�4���0��=LD|C�'�@�r�Ȝ�I&2D��O٣=��L�'�x��d�ĝ?��1�T�^�4�iZ
�'-���Ed��S�n��'Ŋ#p��	�',���B��-7��%k��]0�'���@HŮ.�1���7\���'�\��­4�M[S�U�D(�5A�'z��#B���T�2�� �4Q
�'���#7��n���.�"{�����'�|�x�e�@�R�g�k ,��'���t���@�� �.`�`�j�'\�Y��]�x]�@��d>*���'���!��l�Dc2Ŗ�h0�y�'}L�!�#�%\�8�P�@�c n����� >�q 
�dF���H
k�j��w"O��h`��,�n,SS�2e�\� p"On�@V/hj��l�sR��0"O4�J�*+y��8�ˌ�/~V��a"Of=3s^�G0��u��-R���6"OR������(!Qɛ)XjT%�"Oڤڠ�ܺ�j�"дueZq��"Oظ�g�4Ih���R!:o��� "O4��S�Q�N�5�e���~�~9����({���3.�qO>u��I�7)��y���:_�4Q�Ռ7D���4�ԫ����e�2<9ux&� ���2><aX� O<9��I�T�fkT7b	Y���'QZmBv�޼{���r�gG�~� ��f��M�Rы�n����+� Y���n�;�0�)f>�_�%��^
v�ؓ� ���L>kNN���ɀ�>ᒭ��"O ��h�B��M��畱"�\1!uV�bU/�&;��		ǚ>E�dD޷Ju8��Z�h0�6a��y�L%m�E�F��P����%b�R��A�,1q�E�"����'��'N�%���C��^ K����إkX�[羡���,ʰ�A���C�M�%�;�ON�*D/ǅR�e�B� `枳����w	!޺4C5�����B�Fa�t�����۲���y����d���!d�K
v�������D��A[�L��ߗ��)ҧ6{�����L.�ʣh��h�F��ȓb��`֪�&\�:L2t��4�)%�H"4U6�
-��	�A�DU���[�"��ǆ�5��B�I�@�@q���%"��!1� ��}A,��h^����1W��5y��M'J�l!I��<!�$�1{L����av��L���~�!��)Br��m4��䠑 Ё#!�D��~��l� af�!&�]% !� �Vt	V)��<i��BFT�\�!�d f�Щ ���$@�Xr��I�!�D�fV��3��F�d��py��Hd�!���3($�X��牕U%v���d��N��|�oޒ$<>%�I�y@�9�HN�<�6eh�cīYy��'��Z�a�ᆒu܌��邨4�t@���O�5���'�bM��Sl�L?0)���S��J�*ЉrT�:D�䣦���i3��+@��)Z��ھh܀�����S]f�:D�#G���}��'A������\�q�/XY�Ұb�'IJ��ę��|�31���rɠdT>D��p�V='�iPm�����}��I!�V� �@`�M��{���
�X�d����� K�<q�H 3�aN�-�����J$���;��'�B�x`�!$*8l�FF�3b�����b�Wq?D�؁`\�@O@@�D�M+e���*c�)ˠAlX8r��4>�FB��/Y��3'��G���ȕ;;�4�A8uX��*!��)+�D���L#�'�y" V�UV@��A��.Q����!�yR只{�~\��%�`dY�#(�]�G-�']Q�hpA��;�v�	����Ov �
;bZ�4�����`�,//�{��[��¢"G" �6D�%��J�l���o��\�`����X�fT���'̔�Y�-Z�Y8E '�Kqf����̾g�=C��[40�,d��H����<��u�%�[�1BB5��\rB�I�6\TPas��Y$	v�M�T!a��7�H�d`%�<C�S��?���Wu��U8d��8�����jJd�<i �)G�R���:��p�i�Z�<qI�]ͺ�#��j;��ðm~x��Ӑ-�>6���Ǥ~�n�ȅO��{8�����ybn\�.��뤀_r��Q�5�ɛ�HO�\g�C�|27dK9N@�1D�ׯW��LT+Dn�<�����>j�h�4D�eºH��/��z�
���fJMF�٤O?���e��:@��,9���	P셷<!��_�v6����S V�a2v ^&<������R̓��0=���?�z���ύ5� �aEC8�����ݚ�/�>�ti�4�J"u0lT��/�&����S�? x����S<t�n�c�"�3J��QsU創U2l�����v�f�k�����Ό�W&��}�<���̚��y��/*�{�o�m����4@xj
��R'ӹ1�u�f�	�~���'� h[�i�1Z�(��%�Z�EdK�'��(Y�
Y���!�⇚1o�i�'�b��V��5��9s��{�8V#��]l�ց�[�J}��'�On���*��hd(Ƹj���
��8�&Mҕ"���l���'{ȝ��*_#nH8PX�$ܚ$X"���$�?���2UO4!"$�|�D�(�����d�Hy�o��<a�� .�وRk�v^�uA�#W��0��^�-��;���Wy��	 �f��@K
��E�%��@��"�C��>�2�͝�n�NL"�*�'$ʀ�'�6���ԸKN�	���4Go@�
��~�V�p��k����_�.��9խ��Am����L h�'9%ۀ��'����RhC3]� ����i��Y���ߗ@��: %8�V�� �b� u2b�[�o.RB�	6`P"̪� S�Utr�(�.%ʓL�R����H��S�Ow�� �n�p��԰����t�'ۂ�:n�+6Փċآ)��Qs��|���#+��Ac���y��R��y#�hF�E�� �W��;��?)##�	Q��P `�:RH�(�i-a�4�P�̌� ���D�1���j3K��y $
�^i�,4vd���A�hyrɝ�2�����Gⓞ;�2� O u2!��_���B�ɴ/��#MMT�̌��.�
8xlI�'h��R�fE5p�T��C���̉l�Ƚ��O�I��ծUFi8���U�~���'w�27�A����K���+&���M�����H��e�d͡'g (dd��OZ�������.%K!�ޯ?��b�I�j�!�0�Ӱ�����pm;p�]��Q�	�Q�ZQ��b�č�a>�OڴJaM3=�5h��/Ae�=Ғ�O��A-@ :�`!î��Lxs��j
����$��w�<�i��a������(�y�A�(_�X�sL��MYXH���طkj�I�b�jl�rbC/
ȪA��P��4D\��-<zt��K�;:~}���G��<��I+?Ƞ������Ŭ)+ZeS�FىF)rt��*�
]���'�J$b�S=W џ���蘂<|tY�a�ߣkqBY��1�{��	�c��-�.O�-*�ᐛf�.�3��%����&�/7
�a�'����2�"���a�^46�`p�',m��κ]����[��}��Si����8�e�[�<�F�����FE��8���e�����u��	�k
C�3�I� �ؤy���6��3G������Ȗ!����Z��<X��L�����T �zC��:[9���!>�Z���\�&�C�I\��L{��.O�\ ��*W<4�C�	pKZ�"���vtd�w��rB�I�o�6����@P\X�CI
V�B䉊Qc6��wb�=B���)���&�%��"~�	�'��0���p�@��ּ4��C�+�nQׅ�5@��pA�`��x�Z�	tYI+TiOW��,z�*�0 �p�BR)�2	~�Z��6|O�!��W)F�`%r�4G���a!�5Sбs�a@}�d�ȓD�9P��3!�����V�.|�?��-�ʥ	3�.ҧ-�)�Hۃ|�Xh��R�(T@��ȓ@�^L�i�	&�$p���`fd�"Ĭ���@�>Y���O��I�/+_�\!J��C6,���p�"O����'˦t�]�Tg�a���'��q!r�K�.���퉴z���'E�"@��Ɋ!@|���Đ��(bd�ε�M$�����U(�&�t@�� SZ�<q�V�)3��ǡU�QY�i�V�_:m�BB	�Wb"}Jp�H;}�^pA�g�2mp���5O�X�<A���F��3C +�;�'%<�"��92铘h���Ӳ �j8����Ԁ�2 K�H�!�Y
��X�q�����}qT'}���RlZ K=|O��A�0`�aٲHKb`���'�&%��)��<i� V }�a��E�$.$	�	�U�<�f���~j$� �3��]�tn�}�<� ��i���;s���Ơ�`"O� �F�Y4�����-ެ3�"O@��5����1|>��b"O��r(Y�j���A� `C�8��%>D���v��NUذi2�)8
Y�El>D��y!�E�$����ƛI|ڕscB3D�`"D �d4|4+�f�"�FEiq�3D��qS�T48�T�c*#2\�y�H4D����(P_��� ֪Kj	0�5D�L���<5T���3Ʌ�Ah��gN,D�pS��P�'5�$f/"O����g!D�t��q[��� T���a�.>D���a7`Yq�+�|�i��f(D�h�� f�XH�e�+��2f!���g�iCB��[���W� qi!�dۅW��eӧ�!.vmBR%�PT!�Oy���F�-�X��
Z�
"!�*)<0�pEnY:e�>�jV�S�!�$��#�<!#S؂B��ti�Y?6�!�	"�0@�� u���e(�*D�!�$�)\�<����6lg�l蔈G?m�!��H�����w�C�:���(Wg��@!�ŃD9�c1����X�b)ȫ3N!�dP���'���|A0���%O!�P�E����T���H�.ə`�Y,^!��� B�mJ.*RJ��dl�Q!�D���I��9(���)PeW_a~BKH��:P�7�N�)s2���k� =�ջ�#T��ybC�Tat�!�P?��dpHQ%�yb@
]��5�d՗J!,����˭�yb.�(c�fY*Ut<���f���y�&�	���ƈ�t��������y�@ZVH����p�R��M���y����x�N\<m��ܘ�dY<�yb��QF☺$JK�`Buu@��hOR�E�d E�]�q�%��Z�*��4<R�#����bEX�iya�&�&}�@Xse�P0ҧ��-`��
5�d�oG�wZ�@E��b�%��=�6d�1Q��iǨ\?/*d�S�
��lB$� �v����
�'`��t�a�J�P�*e�!���I��h	��7� 5���=����V>�ᧇ���]ȱ,�$,��C�K�~{*�9���0M��.�0`����CŎ���*e�I��ƕ3�>@(A�H��"5�B�$lbX1�Ow�l��B�N&Ty��(="�M�gG��>o"�t@al��3♄�u/O�8Z7K�	MǦ�@��(��(T�ONl2&èoRAѶȥ<�~���:Y�yU�$� !+H�f�4��W$"Lj�LЁ�?a��	�)�m:��H[aFY�<YC�(��`%Yr$�4'b��E�ӵt���*�<E�d�*T��� ��d9�'I�<@��R%��n	���!9O�}��'o���2&�Н:b,D@�.�?V� ���M�c�
١�'����$0�L$�8��`��mǐ0������A���In:��qEd��0|��J�I�z�	󤆳e�Y��_��~«'4�)�p�Ҹ<������(6��2�n�;���E+Yֈ�j3ρ��<���Y1\�p�)��S�T�OA;$#	/#��|д�ю�@Ŋ�0C3�ʓF:
&�����k؉<\���&Y� �`���Ziy��ڠd�|r��J>��hʸa�橃���A'fyC��"D�8���ڒJ
$ĩ#-��h 0�V�?D��#J1Wx���S
{�)�=D�D@4F�� ���e׎w4}�`,&D� 
w!�i-�,���B�򈙵�%D���Я� ��`22��<�sf$D�l�Q�]�4��yxCK3W����!.5D��ˠO9<my�c%Ϻ�*�g0D���t�@c̜Q"ʂ6�lx ��*D���DOτy]~U3v��>j�N<���(D���gb�*�|H�f-�=��ą9D�$�1�[�V�����l��La�:D�� ��[ƥ�C���s��tL�e�5"O���pÃ�w�&-����7��i�"O��x���%-��4q��S43f��#"O t����H�Q�A+�.�2�"O
M�4$��U5�9;�+B�p�x��"Oz}��+M'��L!��[�$h�`$"OL�M51?저�J�	OL2X�$"O��"f��@�\%ȉfJ���E"O�����6%�`�*cȞ0l>6ٱ�"O������ ��`����-\�pt��"O��"�B��r<�iC �/"��ȱ`"O�u ?�0К#/ſ�`�2#"O���E���5�@(����ad %��"O����H�% ���l[�i�z"O�U5�ʰ_��a�id�x�"Ou��dښ������R� G�zs"O.IRO�4<��s3f�@v9h'"O,��rc֟x;,�@w$�/W°q�5"O��bF�ä$2<R�G55�,���"On,E�\����
Bl���"O 4��Ľyv�QQ� �xh8�#�"O�H�F�ʩ�و�`E;5��|��"O��j A�DS��i���]��U��"O !�t�²-aL�I�DH�Q�|��"Ox�P�bN�^H�c[�mX�  "O��P5ixe����cd�h�"O�0�Q�O8d1T��fcS#_8Ц"O`���<d�th�#A@�DS8T1"O�tbG'��nNR(0��>	���2�"OL��Ņ�/��P���J�ڜh�"O�⃊�Ux�!r���#�hy��"OT�k��St`��	�Y�2�H�"Od8��ť#�V����ǢD���"O���逌|W�a�V��Ѳ�"Ot		�һ�$����l�S"O�E��g�7n�@�bUDM��(D��"O�*0J �Y&$�6⃈tO�HxW"O.��N�`Y�ScT����"O���@�.��	�+J�cԄ��"O��%Gבj��s��ޮiUX���"O.U��EΏ1�1B�A�-M�$kG"O���,fn�Q#A'3"=V��"O��UL\�cj@x���I9*�g"O4uѣH
:��YVΝQB��"Oص;�Eۼf��!jB�N�1Z�b"O�I蠏 �m���:�����q"Ob����M"jhQ(`�;l	zuȲ"O�}���F����(V�h�r�Х"O��ja.֫Fz��QF��3��d"OX�R�#O�y�Xa.M�Q:�91"O
$z��߯�<� ��:I�|��"O�� 1�\��rD�g��!T?�Q��"O ��GW9+��+U�F�S8�M*q"O�Q�p���3
 U�4�J=V��[�"OJ|��_/j��YF�N;v\y;2"O���āI�~�6-�B��)p���"O�P���ֻ:,XP4��#d�Й�"O�x�1�'8�����,1 �C"O����F�~�>��A��`���"OΨC�
O,�����{�p�"Ot��v#��)��i���6
���"O�,q��[?ʡC����X��, �"O((��mG>�
!I����tX"O�����2l�c�Zy`,@T"O� F9 b�G��3��� w2i��"O� f睴
� A��'Y�G{����"O��@�%��Z�� ��]�-s�ta�"OLM�.A�n�8( �PXm+�"Ov�0��"v? `����)$����"O~�)4DK�c�����ݐjmf-�r"Oґs��9R�Ր���v�0a"O�����<M^F�B����x1cU"O�x�A�0,>�`P��W'�j��G"O�(���Cp�p5�D��
{N�m"O��p	�$H89�kH P"mc�"OL4Аkח~{&���뚬S����"O�!R�)^���u���ݎa��"O���u�G�+ ��)��\Bg"OL��%AT�Xq�d	�)��3�"O��)�]J,{��̷A@Z|��"O��*�Ε
^$D���G�=^�4"O�T�%ϞL)(l���i�"O�R�� x*�4�k���0�f"O��Q%��Jv\���	D���X�"On���.��I�F�)p�M6B_6��p"O����Ѳ2�@[� �[��5e"ORy󆃉"7wXMAF�_�l�`��"O�������M[�.O "���&"O��x��9��b�L�G��Ek�"O�y���4:!BI3�J_�C�٨�"O��A�I Lx&|��]F�$ѕ"O�h��$�f'D%G!o8���"OZ�A��#Y��$���ЗlO�Q�"OF��`R)\��<�aeB�	ؔ�B�"Op�퓻[\���0�Ȫ�~j�"O����1ll�b�4�r��V"O0s�n�a� 9���&\�(%�T"O��[��S�c����p���;5"O���^�m{�)���Ď>�vD��"O�TSQ���?=�b����;v,hP"O�Ĉ���a���R+�.��!F"O�AZB�' ���Ɖ#an��"O<}:#P*{l���
R[N���"O��	D�I��1AbU�&��Ě"O��E�ĢJ�ԩe#�}�jIE"OR�� �3W8�$��#!R�"O:h4�-�~���&�A��"O�Y�e
��Q1�ׄDr���"O\q	�Q:�ś�AQ�Y��	"O�EC��s`*��
Q�8b"Ot58�Ɗ*����e VR4 �q4"OT���L˳zČu3�I���{�"O�ÃY$3yT�z"iLF�ȹ��"O\Tz�gU#�<,�CQ�Lx��j�"O�1���0%�F���k�r�F<Ҳ"O4*wA��bA(l(�A�5�A#�"Ol�H������d�	'�(4��"Ox���)�j�%����RI#�"O��B�K2:����EՌ ��+0"Od����-,�J���E8x�؈�"O�� ��N �3g�6���t"O0�	a�q�b�3�&�:��d�"Of5��ӳ�n�� �\\��|�%"OX�����2�VY��C�]۞xC�"O������6:49&M�����;S"O��K���6LW,��n���2v"Olh�ti�*�Fj&��`v��X�"O�!�ugǹaC�Aڱ�Â:I�)�"O�  �g�����F,�'B���g"O$X�����l �kWV�X��"Oh	jp@�wN�\U�.l�ʳ"O��� 5$N�Lؐ!_
CQ�0��"O�3��B�tIP^iv�0D@SY�<Q ���JA�Ο�
t
5GS�<����/(%�5k�b]�I�l\f�<�MD�'֪�� 6;��9F��b�<�Q��3���ҖΒ��j1�w�`�<��+ܞKע��2���Mh3��g�<���N`VTzR�8ᢕ��Fx�<�i�&T�>X��#�Q財�%��w�<��c��Qh(}��L_8!��pဢ�h�<��k4pF���e��6tE|A�o�b�<ٰ��	^���C���<91cLH�<I(E�?.Q3A�R�ETT��RN�|�<��G;Pr�苇�Y�W����u�<i��-0{���jB-m�6EZ6�n�<��K�4���6�M+N�,���R�<��g�UC0eG
�H'�)��P�<�EnU�\� ���T)l��aC�[P�<ɰhP�C�ܜ5���f�@�p@	X�<!��\E���U3J��@���P�<��*Վ9ZMQ��Z&�m`�Rq�<�'d<A\�
� _3Y�tYp�Ix�<y�`×\7�q�-J`�.9�Gt�<qq�8k��{�ד@+��*Ls�<�1È�j�Z�땋G � �d�Iu�<�j�/"�u��P��4Ѡ��g�<1ҩ5��`���>eL��H�_�<A�BZ�W�Z!�c�	�<�[r([�<Yq	B�2p��	���%�8�Ӈ��V�<���,*���vHY�|�<��e�z�<q���3.�L��DE�DcD�� |�<Y��\�t��L̝~�8�0��Wx�<� H҇m�XY�꜖bU\!ڤ`�p�<�0�93r�MCr�N>e�q���Un�<�Ì�U���2@ ��
b8�pU�g�<�ҡ���݋5gΟOP�!�2�y�Y�z���0�k�"Vș�Gǟ!�yR�S
͡��	G�`�h҃���y�L�[���W�Ǯ@Ϝ �!�6�y�펇,BX��ɒ>�|�y��5�y�,I~"=�!��]�p!��y�b�7qn@�3�� J
�8�C���y�$S���S�X�o�����S�y�'�#L�L��D��cx�J�C��yo�� �I2W�W��M��`�yMr��)�ģѴS�&y��&���y�e�T5<��P��b��Y�CDG-�y"�O9S)*�� F[�bV�M�+ރ�y��^�:��!߻`�*]���5�y��=z> ��E�Nn�M����yr��>J��F�ÆyQ؍:���y��G<T��8���#n+VE�sDؓ�y�)�:ZP������3#�Ȥ�y"��c p  �P   �	  �  f  �  3'  �/  �5  <<  ~B  �H  O  EU  �[  �a  h  Pn  �t  �z  ��   `� u�	����Zv)C�'ll\�0�Kz+�'M�Dl��$?O0=;��'��+�j�c@9�[�F�h��wiX�.3�p�bę�wwђ�Q'<���3  b݁����?��g���?�8AV	g0�%O\z��63�x!w�V
Lx��M��g�‸�ʒ{� �;g�b���'�?�j> ��Ũ���:Z�p"HD��ޑ_����I*���m��%���ݴ�h�����?���?���nD��JG�Q&��h�ě�b��y����?�i�2X���� Kh��I០��;F� ӢZ�|M�I ����x�h���՟�ӯO����w|��D�Y���?U�C&	\l��e�E佘֡^~�<�v�߭r9ԭ�K��8XG'@|}�>O⟨sKU�=�'�
�)����i�̝�W�?bȎj���?���?����?���?�.�杗��)�p�_�K ��c���Ĉ����4c�ve�>)&�i{�7��٦�R�4�?q�� �l݃e� 3ѢIR�mՒO���x����' ?RPzF�f|�����$(`��B�#U�#a�9 ֧M��z@n�#�M��i��3�P�
c�ï	���Bh��Z��8���1o)��'� ��%kX�@DxXs���?��a�B�+Z�� �bf�>hnZ��M�f��j߲aے�\�`�c��Y-2�N�5"Y654�a)b�it27����,�$0�4�� ;g�j�`'Bx��!�<�\CsB� '��q���5.� ��`�+�M[´i�6mU�`�I��'����V�3Y^:v�ˬ^Q��� J�>&�a:Fb�⦥#!���R#�D3 �J̚�����X�?��L-z7�!�,X���'-U�,��Т3� rU���k�HTo��?Q�� : Z@f�:?s֥�	]���3�@�r���A����Ҍ�ȓ�! �ѯ35�9��2�:���&`�E�Ԃ�-0��L��[�_*���ȓ��n����f�* F�9�P��a�<�ï՚{�4�p�%�J�H6
Ri�<�'�A1}jHl
�L(i�0�� �|�'��)��qA
�Y�D�C�����'�9!��� ���M��2�H
QE1c!!�$X3qd1��5��L�Qŀs!��Gj��9X��P�e�ND�Ƥ��R�!��Խ,��ݳ&+�٠U2��A�!�DP�*��a;UF�1Zk�Y���!Nx��	�O?}��h��p8f��%�5��p' U�<��!Z<6	2�B��Aa���R�<R�H�J<����l �cT؊��C�<y��S�����!P��`�z��y�<�@.[fB�Hzv�Y"���Ӕ`�<��ޓ,��eP�-EF�P��k�]yb�N	�p>�A��s����\�_{Y��l�Y�<����h0��CM.t�ԍ�e�V�<1���QBeř�X~�@���j�<�U 	�rH�)"�C!&�,J .b�<���޿. �R��d��I��IRGx�4:��� �M����?���#6��a���?WBT������?��
l����?���6]6���W`�#������+�H��x�L�(�2���{@��'3�#?�Dŝ�}�ԭ�T�B��T��'�"��"# c|�H#�ކ>��%A��(F`�<�r�ϟ0��1�Mk�GN��č�:�r�#򭜄
@l{*O���<q���i����QJ�.yB��� ��)��nZ�y�`iKF��(�հ�n��������شL��x��?�.On�9O�[�lij�A���z4�3!�B�$�p�8���a4*�)§Iֈ��үFĶ)�N�$j6	�'�b�
C��@�S�O�T�s���N�.͙W�ޚ1:P���OvU��'Q���iL)d�:�����	�X�6�F<9��'���'�2ٰ�d�(.�he$�r��܆�I��h���y�
�&ae�DiUL	:'��`��KhӮ\"��<�fE��B�g�'n�����q�"�q6oM8$>�|Y����,�'�< "��ǎ�Ϙ'h���eJ�`u�	:W��1���T�L(�	�5e�"W%,�3�ɧ�(B���+tʸ�	vd9Y���+?�3���|��@y�˽!W������<�,���!�$��������=E&��������HO�	�O��t�b)�B�5nW���ā:1��ٲ��<���p���e�j��5Ҳ ��T�A�B��?�ЖML;+�D�A�ڑv��$ۑ�&����+���ɥ�&qȄ�r��ɶ6�4���Z���P�J;t����8N�g�!D�8�d�i����K�L�0�JP!"���e$�<{3g�)��!a�g�=��2&fԆ�B��IVy��'��'I>e���,�@	�W��@M���� ��yסA,N�H	�Q*V�m�|�W�'�/���C�
��k��	GZ�)6�Q!�tf�XC��?X�x1+�OD��ORܙe�'7B��Ԫ�O�*|��1���"#�����!��O����*{�|(A�J\� {:h���H�2�O�ɀb@��N1|�c���x�0��E�'�Ƀ	PF��ش��'��	�O,���ַ[�.�P�#G���њ�I�O��䐘rN���B�۹3�P-�2/�[���2s/�� �r��nC�n	��{��s~ZMi��:��d�z�ل&��dM�X�����E��p�d��qZ���k~��ޏ�?Yu�i�:6-�O�#|�QI�?((z��A���c�R�I˟|��I�t��p@���4+Wz��׋�G,�?�4�I^	�KW��P��%�J��E�ݴ�?!��?ѵ�ݷE���A���?9��?��w[
�YPaD�P���pjC<h����/O@���;�d�����.�Zъ0 0h(܈s�\�6MH�*X�2z���u�1����D�3�s�[���5�̗,�Ҥp�R���3����:�<���po ���(�,+x�<�=.*Z +O��=E��dߜ+��%�3Ď�v�&�"C�
��$�֦�a޴���|b�'����$��%&�L��%*)C,�}�'l�!2����O���O�O���'�2Irn��Z�X����Їn����X?N&`[wN,O8�C秛����`�I��5�ʙ(T��� �g�L�`)�-Җfо�ۗ�
�t�צl�������U�Q�DS%���*/�!��ƩO�H�A 8�d�OЉn�ȕ'<�_���O,!x�I�y�80cVkk���K>q�Y�Eٳ���tuAԁ �>עU�I0�M���!����'�1�rO
��dC#��I����43�RY�uJ�_�!��1�+�U�7���s�ɶVF!�䝡~,����X
�*`��8+!���;>�AA� [��I��Ȁ46!��3:8 I�0��0�~�j�T.e{!�S&�P!!����(D1r��0Arў4:ch6�MF��CWA$�:���v:��ȓPx@⦯C2m����e1a4��G֨z��:rȝ�n�"��-��|71bT�߰MU������'��ф�i�%@�J�Lz����TO�Xl�ȓt��!Q�� k�ʸbg�� I�J��ɭJ$#<E���|�v�'ꃄ?|�v��3+�!�č+|���RW9|噀2 �!�D#;��\��H֑Ռ��u��W4!��
(
�B���CW�L� ��AOL�h!�$
�C�J�1'�!S�H��Ã��U�!�$�zf^� E�O��8�t#���ɞ9�����??�ArK�_~��d#��K�!�D�J���R3i�> |�!x��"7�!�ě�&�6��jŽh��G�6�!���-�I�R�O�U@�(c�G1J!���'.V����� ������K�*T�}bB�0�~�d��P��}�3�<S��y��'>�y��ҧA���� ��
YB9��܄�y��0gY�{��ĶR�����yaS�C,�Z�.U�� �AH�y�bP�	[TAI��Zw��-���G�y�� sN�A���?q�R���M��hO�����5=�ja��\g��[�)�f$C�I.A���H�7n�,|�@�A�C�I|@"gd�?Jq�2��7C�I�!�؋Ԍ�>�D}�4�F�	�B��>ql��i���>i`Xq��剈S�B��;<�@�@�WT���L��/ϔ�䋱��"~5��a�*0I�D�F��K'� �yr-_Z)
&炙p�h��'Ϙ�y2�;TqJ!�b�L�n�x���W��yrGV�~eV�6N��=;6�h�֋�y2�J<b��rn� `��iC���2�yR�D =��l���W
��)`tgL���� ��|B� �P���ӀH��H7���y
� �$j�&�4DK��h�'�$��@�"O~�A���v@���R7K���"O��2]Y	�QE$K!>}� rC�X�<��+O87��aJ�E�{8�H�6��zx���E�� ¥ΝG�����s���h8D��"��ˬ��Īm�L����f,D���d_<"<m�6��5Ug��s1�)D�tR�DY�{G`e "Ύ�2��	��C'D�X�KN(Y�Ct�K��& 'D��!n�2���R�*K.����C1ړ:ٺuD�������F��_� ��"B�y�cT p�!�1̓)Ԅ|I h��yr-VuS��q�"�2paj���I��y�
�~��gd���X<@'���yr+O�V��)�#�U@4�,�C����y�oM�&�HQ�S?"�e�����?��f_k�����(��*�0a�d �MY�x�H��A>D� +%�D�m��/O_�e��g;D���&�.ƹ 
�cUJ��5D�TëѶ3���b��Z4tW�]B�/D�����ԡJƨ��(�
T�)9�',D�Ҋ�+h�,4hr����K#�<I'Oz8�iaF�g���k�����A';D�Pp`��/]#V!���C�J�*�f8D�p����z$D��8��Bb8D����,�8[K4�{�bCr~V�(@7D��* ș
+	���U(�#�J�[D�6�O�1���O�=*w��`�fX�S��P�`�`�"O�;g��@�Xm(� �i�&i��"O��1D��Z�|�5� �HV����"O>�s�@ܧw����A̿/���P�"O�����r�d]�.B�=�.�HQ"O��O�<�0 "�޺PP���P퉾:��~�g�я:hj���
+�۔�~�<�΄<�T��6�ײd��5�իR�<	�	�'.\��a%�6:`�JV��R�<Aᢕo��� 
[U��� �V�<�`F~k2d�m���ցQ�<�Ѥ�/r��I�+�4 ��ͫB�y���>�S�O�FH D�Χ%<�岵,Ҵ9�����"O�)�_�I�P���%ˤ|�̭�"ORt!Ǆ�8�`�Q�I7����c"O�Y�+��=$-����9�d���"O��!ڭG�b��O�Kjm�"O��
ՁD>GD8�!��{msX����8�O�x���R�$`3̀k[ ��"O�u (��<%��J�A�t:��4"OJ��c�A*�r�9��ʋd_(b'"Oּx1@���U���	/e����"ObѤJ���ї�N�Q"e�U�'�ܘ�'�R�;�Eg�ƹY�̈́U�ʅ��'�"Љ���? ��e!�-@�b%f٨
�'��ISbMf��=�ĄgL0��
�'��q��, ��ы�FF��b
�'�F�S7�p�ޘ����"�,
�'Y0��Ro�X�F���,��X my����sQ?-HsmE#^I�h�VF��t��3h+D��K�P�U�Bm3FNʛ2��sV`5D��qp�(1�6@s��1��aRb�1D�0&gV�drĴ�玍�e�(�B,D�$��!>ک��#�����zsn)D��`a�#J�A���$d��Cf��O��y��)���8BF��$'�rf���M�Z�I�'D��R�ĎL�`LZ�)��TdX��� �ђs�6g�vL��̔�s��	�C"O�S�J5�2��Tk���>À"O�5yV�Y�!�|��i־-ݶ`""O`�f#�<*
�Lr2������S����&6�O�9(B�	)P�RA�5
<:ϲ��"O�M0R-�2��	@T	�q�r��$"O|�%�`�̀�g����B"OF��4F�|�����ř���K0"O�%�T
U�2�`�У��8��'z��y�'��+�FZ��4ň��̾	����'L	��4]G�����5��P�'/Ґ��G ơx�jͬ*�d��'6�Qؕ����pKч۷�6���'����1�ѧ^�����Ź?�}	�'�.,�)�(!w�	���b+tpp��$�t�Q?�����7@��{�*�-&%�śC`,D�|w��
Lxh�y!fY�,�j%��K)D����P�B����eU�B�RQ�'D�k�)�捻͑"�J1�6�&D�`Q`F/D�y�� ��5�G'(D�L�%��n U��oN�5�ȉ�f�O6!��)�'2qh	Y�+�A��h:0��'����K�:�x�b�hR���'DިJU$[����yR%B�KI���	�'�d���e�.Q{Zĳ���J$�R	�'/�z�χI��1�dԖF�̒�'~l��E~ۊ��b�#/����*O��1�'u؉�vjߝ[��P���+ق��	�'�J�L:"]`P���((\�%�	�'c�2�ܮ2����Q4��S	�')~+�C��+[���U�@*�����'�6��cDВy��XR�(9+fn���T��=�-!��5���G_,q���;s Y�ȓ|Bf�;�/M�i�HHB�G��h�ȓ`���+�l�j�j���G����ȓ�@1�U@["�t�4��,]ұ��p�xp��	x~X���P����d�FE�DlUc|��A`�C%㰜G{��F������P ��
3&�/"Xd��#"O�4*�K^�=ؼHC��'���"OB�����0��%z�:��<��"O�E�DO�(�j�s"�����"O���PAZ3z��5�![����"O��C�LЧv6MQ�ϒmq��T�'0������ӳ\��k@@٢ l��������$v�����)LC��)5G�V�zɄȓ[m�$a��[#O���ce(T⾠�ȓP �{׉O�uZ����
\��(�ȓnv2˳9C�����ZM�ԇȓI׮�YD�t�"�)P�HI��'��-��FW�A@��F�[N��� �����pӸA�"���ۺ<����( gy���<u��+2��=9 F�D6@��!�Qa�Z�HP �@PU�ф�yL����U�:�&�cA�D�݅�	-;h�I0��8e�Q�ƽ��e��B�	�2�b��R!���n@�X��B䉙b�����G�� �;⬞�tB�	�U���o�:wM���K�2C�	
�-��^�PS�t�U-݆+.C䉐%��$�B�D�9a�x�GO�2a��=�Ӌ�Z�O'Ѕ(t.��u��2��9��-8�'���&�4����g���$=
�'N�K��!�8E+�.y��<c��� ��@��&���ϝ�2�e7"O��)� Í�%I爔V�Q2"O>y����1�D�cw(=Z�V��`�'�A���S�;��D�pϋiU��9�A��:l��ȓA~>@��*�s�.mQFʛ����ȓÞ|� �)JX���O�X_���Q:| �!�JPp܀1��6v���ȓ@1�� ��:S������Ąȓ^)��3��>V�ʹ� ���"|*P�'�h��w �(x��T��qRΜq�깅ȓ �x	� S��B�,k8-� �]�<�S)�ɒ���L=�P#熛[�<I�͐�@N�BR#S��zp��K�<��CҰXE����EI�	���@Ix��Y�輟TxF7j��4jsJ��s���B�#D���F�*�������hÉ'D����m�_�4�C�
�YTB�R��/D�l膪�xf*u�фG9m��c�f*D�(�(MJ16uz$K�)Z(�5M)D����a��؄%�/l�rĀ��;ړ�H�G�4Ę&d�XH�)^-+?����/W�y"ԬM�lq�l�;�1kW Y7�y���b�Y�@�K�H%�F��y�jֱVkRM(��ۛ@�ū��>�yrjL&S��T��gM f������yR	��-�.�K�B*g,�h�rHG��?!5D�����8��ȓ�l �mX8�`*��?D�|�Q�mR��c҄��P�n��5�<D�ثd�6~5�U*Z��X�08D����$�hH��YS��d��p� /7D�k$M��L�jaAb$ӛ�$@ȣ44���ӃAu����$�ӣ'=���w�e���	/$X�����	�Q�°`D���.u��o�:>���'���'��g޻
E�i#�jG"�@�TnÇW��)�s�����$�^t����3�"D{@���4(�]���S�?�{Te �Z�b�o͂SO�,��A=�}������d�|◡Ӹ&g�:W�K;��!i�Yay"�'� �`�/& �vMq*�I���6u�I9f7�x:�E @��A9�
�j?ʓ9T����UT s����i�Q����Or��w��%3-�&�g� ��i�O�K@F�J�Yz犄�_��\�7�R>����S�<3d�q� �8l��橂v��D ]�؉2��J��Lm�T�t	��i�?v4SQ*�G�I"��c-�1���'��)��4?IgL�4f��0�dOѴ@F�eZ�n�<��@nH��D˙6��	�t
j�'WL#rCn��� !3�͈Ya�E0T�3,��(O�9Iu�զ��Sǟ�	{yr�'����ܗ��T�_}H�SgU:C���e766qk@"!P�1�O �O���#�	�i��j��P
t��&�D�{V�ip�f_�B�nYT��#Lw��e�&z�:b�8'�k��G3n��0�'I84;���?Y����'~�H�]���s@;Q��"���<a!�$ї4���Ro��M��xy��7R�1��|�����$�.h���B���#����څWl��C���Od�5��Ol�ĩ<��S��չGf�� ԧF;m|eC2�M;,B�9H��^���4���[�m�c14�Sޒ$�1JV�Mk�D+�$L(Qb�QU���hm��-""<;�H��O`,���'���IW�ږZ���1v�W�1$�](a�'�ў�F|b菨`�n��B! �|����Ñ�y�� �m�4o��y�J��nP���Dæ���`yo�= k6��-@Z�d~>�p��%S<�X(!�m!�-J4�O������O���O �h3�'@�)�̐���4�@tA'K��5�B� ٞ.��y��	���c���1m���H|Z�!�0^�0T��fv���Zj�'�0�)��?Q��� �0�L��04(lbB����<�O:����ȷM,q��ś���y�Q�''ʓ׌����D7*2<�Ѫ6 ���?1�&��'���'�R�j�Қ#�ڨAb��jx-y�'â��g��,	:�z (�Xh�P�' j]�oP�E	�Y�׉����t��� 6�Ӧ�U�t���+ ���"OV�!�/�=�6�ñ	�Vi(�@f"O�$���?��P(�1y\����-�O��}���p��kB�X͚���ú]�4�ȓ&j�!roխd�~�1�cКX' �ȓ.|(p�&��S����(�
!��Y{�!���
�}mԜ��'Ep�p�ȓ>w^���Y:S�d� 'ψ3Gp��ȓE�~�E%�%>b� �%O<[-���!%�,����r� ����0)Z�1Q��.?�!�d	؊Ejb�ߖX  @�ů϶ul!�D�]G SƋ����(��f�!�d�J+T��J/7 ��3��x�!��ZR�.%8C/�lA��c׻�џd�g a��|2� Hێ�i ��?Z�ސP��g�'D��p �WM�O�0$S"ъ�8�(�g]<���I��DRU!<�ˊ��Y�-�x�C��{�&�JU@Y�8��<[���O�8��\4�� C�ۃ�\�k���2/5��D�O��"~Rci��0�YSLP0V^a!W�����>٠W� �ES""ܻ��
:���xu��<���?����?�L~�/O4��+��@w�F"P/(jq��h9O��=��N�-��a2�R1@��Z�HDr��M�N<�r�8�5Nc䰈P䁡+�p����O�],�C���8]��S��'��q�$'G�@���<$�V�JwE��~��I/���$M��'(n��)h,� q�Q���*D�a�Dj���ɚ�~��s�<��a$\��i�cM�r����Kץ��'��'�|E�I�l��R	{��"m�\��ǈ�({Vѩp�'��%*I���C�.�'|���W�N�n��S����A8�M�ȥOL��O�)XP�>q`�i���Ӧ���U��5��!"�@��*OB��'�>����7B�uS���*ǘ��!�:T2A �'�6Q�I���<yR��l~�,��Sr��.�02a�Z���Sn(}B��6����>�H��	��J�/_,:A��8�h���'�XT� ����9O�� 1�O^ 7�^�Ƞ	��Z)O��|�s�'�\��	�e)x��H�%���@��PXB�	;M�2�����JC�i�Lh��b���d-���E��O��禙s����	s %��M[�SdL�5�>�K>	�������'8�Niѯ�5fc(�(�BH�s_�'�ўb?�E��/.R�3��>�p�6D��)!K���H��P
>T�Q�8D��i�*�'t�� �L:
��}��#<D�8� �Q�\���ʾu�it�>D����JK>Np��� g	�R�=D��P�nS�B�,ԫ��8/��q�O9D�`��)�&@�M�"Y=�U���9D�t:$`	�x_���0J������v�6D�0{�l��32�(����̥֦6D�p#�N�0ǔ0Y��.W���B�L5��hO�"�I���	߄M�����#s$C�	(��� eA "ar���㛒6c���ͅ@�Z��#����Ag�e\�,�+�.1p�qui�d�j�!��Ҽ�9�%[� �&���Lz���KV�)(j�P�o�P����'&��3�LxB#o(Rl3��0I��q��NU���B��3=�ys��C}-�Gi¢v��:����{�j84�C�c���f�l��ҷ��G��u�����?��	Fj@���Ib2́�G�S�� ��[�ʧ��I&/���"��
�]v��Y��	�(��'�2d�@�V�7r��C8�'XfB5����8s�,��;�l2���/R�'T�>�m�6?������hx��D�x18C�	�*��x��J̫U�@ �VLF�
��U�'�d�x��\�.D�Q`��E����O����O��d�4�T����O����Ov��w�@y�-��%�(����;�R8;��+�� R��Cx��䰣H�$�Bc>Y��Od�����r�V5�'m�8��|�eEM���Y��i�����Ę {�pb?�@�OP}+�_�M�� �'�S2i�,�	U��l�'-Ԉa��|z���-��`0$M�VA�+�����!�d^*y��k�#�Ea1���#�V����S֟��'��R�m��c�X	d�#4���'Z�q�Â�_�(4 ���!�x����� ti�f
�9��z��T�fp ��"O����H!<i<���O�F�(M��"O�PS@S o�[rI��^�v��c"Oj�+r&��5{"�rFV���g"O���EM�x���;(�
0��"O���  R�9`塕%�42�"O���FM�*u� )I�ƊR�6p�"O�!{��À\�����e6c��P�P"O�|p0ċ	��R����"��U�"O�Pq����b�(��%m�H�l�"O:�lO��D���4��L��"O�!@Өi�͐�jE�,�d�""O�����K�~��pSR��*R�p�x�"O`;��<x ��uϗ!{�=9�"O��S��+6O�5�獔�zW2��"OX�t�r�j�?l Ie"O�A��Méd��LRe�C�n�n�c$"OPђ����c�$�J\��"O6THQ�Զ\��Q��0{��u"O.�hT�Z̑Q��� &��"O]x4�1��`�ҀA�2� y�b"O���`�3 �th��'~���:�"O��dBA54�Z��.CU����c"O%����_�*�l�7DP���#"OJؓ���5H����+�#mR^Ear"O�����2l|Y�*jE���"O�%��c$W�
�RdT=H՞@"Oԁ�QgƇ=%�A � 6Y�fI��"OJ]x�Ȉ8%'�ɨ`��]����"OZ}�J��T��\��F�@p�P�"OD�h5�� 71@�9ՠGtkX�X�"O���O�!a��Aw�L�Q,�J"O@�+pa��k�,�����5��H3"O�ЀtG��,����!�-�����"O"����w�D%��a�->Q&�t"Ot��H��q�F-�!�����n:D��pTO�?��D�aE�z�Z���7D�8���/y9�	U J$ �(��6D��xD�R��uKS������8D��kG�+&��j�O>1A:)z*7D����!XP d[  /|6��G@5D��怞�7G�A[�F�;
�,Q+6 !D����Q��0��ڸ'�V���D1D���}�F���`�6D�:�!=D�,�C���=2�+ �4���U ;D���늂��(BϞ�^"i��%D������8	o�X2t� .�qXsk#D�hw��(7��a��α^���0  D���R��9$ '/�&� ��ы?D��P�`�R!��°�ަ�6/#D���l�0�h��&N�&UR���?D�8駄��g�H��L�FT0ف�>D�d�ц�,S���:6 ߾.d� X7�'D���2ι? J�X"�?{��j��2D�y#
��O*бsȝ�{��P��4D��crD�k������]�N���5D�$��	1ɂI9�N]�ް��s%4D�h9 �o4��F'Φ 9>h8U�3D�<���;`L��!���99��t@%D�Xd�S),
���H>����f#D���B�>�.QG,ƆDTJ�F�4D��/C��F�IuA  �Ҽ3"�2D�l� @Шh�
Q���)3u{Nub�'��ݐ��>�y�����+��5�
��� x d#Д\Y�83&��aCjp9V"O� ���{���J4�Ƣ{.���"OPDyc,Y<!�v ����d,�R"O|L�6dQ�4Q�%��(�.mvth�"O�����Q !�*����"G��hp"Of`�q��0%A|��'�
 [�"O|�(fL�$��0��ׯL���"OL$���:vv���D��8	¸)�"Ob�SNB2&�#RM֥Hg���"O"iw �x?d�@��Udf��"O҄3�.� 
6s��ܐ1a�aY�"O�]�񆎫�l��W"_�:?�+�"O�����B$��2�Z�:�"O�xH���h���� �2��(K�"O��Q��Ӓ��q-B��X��"O�E��O�Q{F)���U�M�z��"Ot�q��[�w�A�E�x����"O�!���y����J2,���d"Odѓr�:E��IA�I��.�A�"O���eMX!Z	 �ʒ ��lcV"O�8Z�(�6��q᷇R�Z{��"O�e��ѧ+S��c���!c���"O 3cN+y�p�v��8+UQ�"Oz�� $ײRF0�5#�yK¼��"OZ��LU�1�]���(H�9��"O��
�(wx��h���=V�hH�"O�9p"�щ<�~�q"�M�KCj�p2"O�Y�0`� �
�
�y\��j4"O�ɓ4C��8*Fm21iC�SRaHg"O��C�ęm�hA��bN�fX����"Ot(�A��Z�a� ϵ=��Qg"O��27K� ��� � #��i�"O.�d
ۚR�-��/Dwn��V"OD%�a���谉s�ƞv�&"O�8h`��-\��K!��1���1�"O�����\�½�sB��\uHs"O�C�,x��Q��6i�B�"O<#��Ĳ"��\�5̂�},��Q"O�±C��?V]�� Lo^<Ӵ"O��s�* ��3G���x�ۑ"O
 i�Oŷ].<@�^�9����p"O.�ڔ)!#�XѠ���*�Nܳ�"O^%0�*�-6��A�� � ��`ۣ"O4԰6�Q�S]�Ibb0(���D"O�83Ԧ�w|nI����s��M�Q"O�`�Ш$B��0��I�C��kR"Od�Q�b�Q�@"�"' x�Q"O(�c�Ӿ6e���"�,D�f�1�"OJ娷۵l��armٝ��(��"O����)�f�n��Ζ�Y�x�R�"O��6��op~Q�2G �a}��+f"O�I���%[̥0�f͐�*q��"O
eJ�%�:��)�5L�Lz�3�"O|�ȁg��Od6@x�/�"ya���D"O(���j� l��*'o�>x����R"O�ȇO�-/0I��L��&��C7"O�XRsҺ.���ڦ
".�A�"O|�rb�1 �p���Y�t9PYc"O��2����
I,8!"OzEh���~-��ڔ�*��e"OB����D�x^HZ��"f(��Z'"O���G�Ԍ�Xq#cD���e1"O�aXV�8F�P�a�b��W��3"OF 8�@��,x:�Г+�@c"O� ��;��ƻy;r9�a�D�j3�s�"O,-�@ ��b]��Ŗ��	�1"O`فᩍ^�蝩�A��dF)"O�pR6��0}���c-Iզ�H"OĘ '��e�@ϣ^"���"O	!W���RD�y���:dx""OPͲ`JO>޵Y��d��T"O6b��%e�q;�o��;P"O�X�t�W oY�����R��`�"O�eY�'�%�<�5���lA u"OX�B#�l	���bD�(]���s�"O��Z��=
�����)A�@T�u"O��`0dS�ӅVV��Y�j�A�'� ����e�x���Uk�)��'���aHQHh�@�ua�0_��H�'Zڜ1JL� _���	<Q�Tl��'��a�P�O2��4��|Z��S�'Aj 0pF�qI����d!?&����'"��
��R�؁(&��:��Q��'��E��!0uL��6j���'�z���m]2����B�5?RЈ�'E�P�O���=XT°#�����'�N�#���*s��i�sJ���J�'�(M!4��O��u�tj�'0��
�'��Q�c
�V]hu���Hv��	�'.\%b���O��"��7���B	�'���'CUN���e�*���)�'��ԫ��<bΥ�e��?*�q
�'��0*D�b)TYH�H٠#����'���碊�d�4�y��D����R�'�@�[3�W��� ��ʑ|���Y�'�l��QJ��dc�h�|���!�'^���������%�B��5��'p^�� 	�Đ	2�B�7H@�y�'pԠhuNO�foZ�z��(�<)��'�����ַ3�~�¥��i�����'����!f�8[���tM�Y�T���'peұ�5xv�0�B:K��T��'�x�C�+���~�"�#I�n��'L%2�BU�M=�@�!I��ʙ�
�'Ͷ@�wHI��Lsa��(P����'!�IY�L�XM�]C�Əx��8S�'����0�`)�)�([�j����' �r�C�8n�Q+K��3�hYK�' ���O�? �8�C��6wb����'��,0��3ͤ��������V�?D�H{0�1�̊�AA�
�ʁ�1D���"H�B;F,À�C�� ��;D�ta�R�d�����6<�q/D�x��ߤsh�B�I�z��	��2D�x+��U�y��F� B�|	1�*D����U�0D�&�Ŕ��Wd&D���C�"�����A�b%4)�I:D��т$ڥ28����
�=:� �;D�lH���a#$�f�`�;�/ v�<�D��5y�e+ិ(���!�)t�<Q6MY�K^f�w��0*F}�!�t�<�!��l">��a����F�%�Y|�<��F3o�m���ٺ�,|j�@z�<�&JY�[��ƝNw 1g,@v�<	6�U{�f�{��Mw��X����V�<Y����"��J2DS�M�<��n��/Z��i�����N�<a��P<	��x�H(<s@k��HM�<� F��s�S�l�R jH����"O���FEV�PUtt*�@�d��P"O��� ���u�,�Ё�ʫ!
��c"O`��t'� �H�[��ߥ?�,�0"O�sť�.F�	��B�8�����94������8�v�qKE"�,��C�	=�r�1w*_�7%�nm�#n�C䉤�@R@�זmN2���F2q��B�	d��A��V�0�h��2JB�ɕz~m!񊝐yaJd�W�՛jLC�I�n6��j��
7/��L���0t�PC䉭?�F�(u�D	m-��
��%D�B�ɘ
Z��0&턁7����fÍ�,
C�	V݀�P��I?j҂��G��?e�HB䉍 ��@RHD�tQD�(bkU748&B�ɢy�����ܞ���*Ԃ$	�C�I�>N�(s���)�|��c�6�C�1��4��k�
s���e�_�LV:B�I-Q�r�P6cH�P�z��b�[)d�B�I�Q!FC�=}�NDȢ�܅D��B�	&L���I���Ufb�ɖG(D|C��j�`9��s�X����Z_<C�I�nl4�ˣl0e[h=Y��Z� C�	�L3�P7G	3c`DU�3d<�C�ɶ-q�	%jr���qeV5"��C��8=��@u��ݐ@m�1f�B�	�q����0hR�>tU`��Y1�B�	XiA�c�F�m� �!�Yn�B�I�+�R�8�-D0!�0�9wDC�ɴk�Ҙ�+.9Q"ԑS��8�jB�ɿu��T9u�f� �� �ŦponB�I�j�!��bR��8Ip�,��'~C�	3HN�$Z��Ӏ?,&����A�)�HC䉳:��)F[�9�F8�l��u�B�2[N4���
ϑ`�d ���2�B�ID뺱#" ��"�B�JWh��vj�B�	�z�a��P�aE������
4D��[$*Ŭ{\�� ^$C��c�/D�H��"6i�Y��F�j\<qB,D��� ͋E޼2s�.]�"�Q�2O�pK�'�!+銉@�MS6kOH��
�'Q��S撀sE�U�Fǵ:�a�'��4���R�8�q��ߎ��ĉ
�'9�hP�%WY�Q!*P	.<E��'��]��cZAo��x�,��L>=��'܌�e�եTB���8<���x�'&���@'V(�m��/�n`��'gH�b��ע\w�h�����L���'�򜠡��O�2@�EW��¹��'���FȸlZ� ����r1��'�R�S��ƟQ�v|˄�V�2��
�'�*�y'˖%[��}���S�N�p	�'ǤU�χY➠c���L���R	�'`\�Y�'ϱd����0�GD=����'D�(�0+^:s׀��-Lغ�
�'ql��L��;�qC�ЀXl�݉	�'��Yx��I0-�퐲#�!O���'��kH�P��U�K�!rR����'8��I��,��` p�ݿo�	{	��M��hٔK#Tp���R�}�
�х"O:D�cdC�Th��K�Dپ��"O��Uʍ�`�R�B�� m2�u"Oj|����E⑨��"A��2�"O�1�c�F��TK'�Y�g���"O� @+��@�YfH����ilX���"OZ�9U〖}6�(�jT8L>��F"O�X�b�(r�P�`
Ԕh-Q�"O$j(�^DP���2;)h��t"Oju�A	BŮL��P".���"O�� FH�	2<m��l ����"O� C�,(s�4�G�%q�Y�"Oz��!Qm}�$`G���^h��T"O����ձX�`��7V]pu�"O��4,
�	/� �5@љ7DxUZ�"O���k��. `A��" ��� "O��9�@ҕ-�|P��(�\�8E"O��
���	%�(=pȂ|���S�"Of}�l��x5aC�]�,��"O�h��Ùf��)�C��V*|�
�"Ob��n��&��r�$R��"O�1��D��v8^i� �?�"���"OV���UH� 8� ο<B�p"O�i�G/��pz���ٿS�=��"O��S�T!s?�U���&-j }�r"O� �F���!����A���"O1��MފO$Z��­˟)�b��"OR�*%�֠&����8t��`f"Of�;����y��X�c[,L��r"O�,�f�-6��X�	�5)��;�"O!�gc̑MD���Z�	(بf"O4aYD���Ē�����<���"O�0�ԅ�"X��)G�+8j�I�"O�䙕�ߘ���CE�.1�Q��"O~����_	�MB�A�,���"Oڥ����n����C�X1$�1�"Ol��`�T�~�����a�>7Z���"O�Pa��%D��H��BұY'�8��"O�$����ehl��㇂*�RC"Ot��d�f�$����-,)��"Oh���,ѯx]�F�� nݸ"O����R$]�A'"�z$�"O̠�âG�Iȩ9���H�2�Y!"O�X��gٯѢ<
��Ϗ^&��i�"O�k�D��3��{ �M����p"O��a��z�����ݦOvM;"OHa� F!3]����f ?3 �x�C"Oh���*�0��T(K�Rт"O��yN$�x�[A/K�>l;�"O�!��M#"� ċ׎�(TP��"O2��gȝ������,\�p�'/�Y��_>�����e�'52"�x�'QB}���ʞOT�y�.dF��[�'�.�*S�G�aDD�����ԣ	�'l�h��6?<�$�Պo��#�'�hiY&(гJ��B��	�$9��'BB�kp�M�Q�2�� �v����'�����"�!d�H�3�j� '�[�'`��JW΀�O���(&ϬB��Y��'}�d�&m\W=(åȏ�RG\�	�'̤���`Q��"PI���#P�����'�"h����*{�U�t�C,@c�p�'5`u!E-��ݛ�k@F�@P!�'��U C�I\p�G��7C���	�'':D��J�����v=�A��'���ThI")~݁F���f��52�'�h}Ƀ�1=l�` �$�b@Q	�' �a[��gN �q���2 q�J	�'Q@��J�+�v}����;��hK��� ���0�\�YȄT��Z�p �"Ov 8���(;�jir�샂:n��R�"O��X��k����$X>�J "O$@3�B�t��KS��.�p�s"O^��`�q��)3����ҳ"Oƌ@ƤM�\S�`24!7 ��A"O^��7��z	$=٧��%w ����"Oft��E�fR��C ��<���"O\Q �h�h�|�"��W{X͈�"O��Y�l��u�p��/U�Yв�2�"O�����IF�����n6'x���"O�ْ���6U��%.F�e� ��"O4�GH���mCCP�!m���V"O�4-%��8\�r�f|��"O&�Iԉ�m�B��VD�x��"O��hJ<F��LJ��Bg��Q�%"O�9��*ΣqŖ�*��C	��!"OR���(������o�)e��傰"OQ�ƫʯy*�Yǩ�!y��11W"O����K8,���A(�&�D��"Ot@՜7�Ll�]	�J�2��Qp�<ɢg�L��;��ŞsB�Prfh�M�<Y�	�]"�c�eO��� D�R�<����./��r�H�a��|k�� u�<!�.���s����Q
�E��Lv�<��MY�q"�)P��&7�|�AώL�<����j��$ab��w�)�祋O�<��I�G �XRl�x�<�2��M�<!Q�׌lC�����A+��Db�<�Q�ڍ9��4�s����lYs��F�<A �J�����K��F�p�B�<yV�Q�d9��"�>IL��#�PS�<!%�x��ZT������l�m�<��A��Y����	�P�k`ODm�<�����$�Ѳ��f�ڠ�C��C�<��`"���@�`B+	����IA�<�"&
I��$�$��	� ����u�<��ɛl����'�AsDؐg�Kr�<9��(, P&���;��x�4�Rd�<y0ҿ��$%�^0VH&�]�<1&��%+�ҭy�J�8��=I�N�x�<)7Fܷi�D���^�Gr�ؖ��s�<a���?v��۵L���DX�fFd�<�@}���1�ϯ4��	P'�~�<����RZh������ua�`Pz�<�w�Po< h`&/_��#�_s�<!b��m��R�-2'؀C��e�<�a؄K�Iv�\u$t�cĊZ�<`�JMx�ڄb!/ȱQ���j�<�Dł� ����#OLDٻ���i�<�dƜa�Bp@�I�`͜eC��@�<�E���;w8irR!�G���q�͝_�<�+`����D�N��M�P�PY�<!��"p���CJ��RT���Y�<�"�΁`"I:Pb���S"�X�<q�BZ�njy����!A����W�<��X����C��<N����g �h�<yq��s3F`;�Ѱ�L�H'�Ue�<�7��H�acܑg@��A�H�<1��$?��!K�@Nf�`�p��|�<�Ă%-y>�j�s���`�Q�<���������~��-ZQ�<)���(XV�;6�IZ�μ��jZP�<�I�'�( $�-xF�Z͂F�<� >1a����x,�]x�L���N� �"O���뉘]�P�A��]��X]�a"Ol����^�x�X�#�NS!w��T�&"O��:��J*'������u$�r�"O�(�@�5[m(�	���n��J�"Ov�����=�(���']0�s"O^-�f"�10�H�PL� e8��"O5{T�ӹWh4�NA�'"hS�"O��CD�;Ƅx���_�g�8Qs�-44� �%�R�FRp#��f鮉��H/D�ԫ�^�8p
��'�L�\�q�,D���ᤂ?��(���'�(0&�,D��󡆉�'�P�'e�	n�h�D�(D����v�S���'l>��v�%D����6s�T����ʄjD�(D���g`��b��$H�:d�x���##D�,r��7�U�Th�)=pc�C=D� �(6_�\;�	*vZ�m�26D���!�՜dM�ڣ%��X�240d�1D�s��3e_U1 � x�*�:&i1D���.���"��A�b� �G�0D�4j%�� )dE��\�*���/D��CAK�%��`��G�]&șw-D��1*'��=hQ��.����7D���˚$�v ��/�D2	�&2D��+�è{�4����x�(��#D�<���
* �����I���ZP�>D���&\����xM�H�t����yB�ĕ�4�*�m�7�z�x1�ܔ�yb��0v��pf+K�7XQa�ν�y�H 3]���+B#_7tB��U`�8�yB!Q���h��B,2��}�E$��y�.x	�VLX�&&�������y�CIx~T	�/��HQ �
ӹ�y�ɗ#F���*�e��e&���y���.E�6ݢ扃wZ�PQ��F��y���	�n�Xt��DzPX���SF�<I�
�!��p3�L���l"d�f�<����(�i+��N�Y.�h7�c�<!���)VdM�¹j�d]���\�<���-e�������-
�]�p��<aU���@Z82%/�Or}J�}�<��Qo�d�з��'L�La�V��@�<	��Ȟc!P  �߈<��4��M[w�<�4_�wS p�Մs����j�<�񡈁q�.%�@ʇ)V�PA�!�p�<����3��l�f*N�f��e��So�<)�
5.Q��C���/K�0rւk�<)�HC:j#H�Dɞ�x�Ԥ���Qf�<�å�?t{����fd�QI�,�i�<�+�,V��:�-�J��I$�{�<9�
y�Xs�ևI|��V�z�<Q�ݔ;.�l�!S��ZW�LP�<�l�!%Z�hB�ĺI{8H`#�_v�< a�;¢�����q��y��"Or�<Y�'�PT�Z���)i*l�XF(^l�<Q�!��@>���(}�`�ৡ��<i3*�6F1����ω3AF`�b��<A1�W�a���&#�*���{��}�<��,��\��Q�wT�	� ��y�<	���)$�H�kE�[j���h�u�<d������C@�v�PAbd�s�<�c�_�w�Ͱ�mL�|9B�p��l�<�p$�	����$^.�v���n�<� ��kE�nad��7�͒@6r�""O����������Z�AK"O�CU�^��N�6�(�qa"O"$�q��q)��J�Dܢ`�b��a"On�I����p�āϽz��<xD"O�4���q&���Z�p���"O�p��T�K�)���&i�麧"Ot�nF�)C��'�R;^��"O�(�g#\�:�铉(���"O��٧X��c��k�"O8���oR�`J��;W�]�5"Odur���
5騑IDd��t�f"O�Mq��#�.!K��Rm	�"O �cb�WwIN!!�_b��"O^�yG�·X�B���MWW�Dj�"On��CÖ7'(p�b/I�UB��"O�m��K�_ϴ��1n�&'EAs�"O  ��a,j��/$��	3"O� ���G;9?4r�
X!S�a�"O�	�u�$pO&1��F�1ad���"ON8 4��t�(J�Y�.T�A+�"O0�Q!C�����"��5e8�8""O�QI��;����΀8t&��"O%�,�=1�N@�!��s�z�Z�"OZ�:�I]�!Z��t;�4��"O�}ڶ� >"8�M� ֢a�"O��y�꓾:���׮�_��#"O�@�F��w��LO�B���(�"O~����N�Q�<����f;"OT���g{�s&�fD�bbj���:�fx�'!U'R����D�!t��T�ȓ.����,�Jn.}����A�5�ȓ]vA���P
Ҍ�F�M-���ȓ	�q�2 ]4=��1@B�V�k(��^��t*R�ڀ�8Y;��
"`�ȓQؠ��U]�p���E"!Jԙ��;Ӓ�m��b�	 !�:1��`�+ �������Y�Up���YI�0�I4_d-����1��<�ȓ	.��!/����)_sEC�I�A%8�Ӈ��mC��J��H�ȓ]l|]��oW�~TtW�pD�ȓ}i���P
_�V@��茷o���klX� �؀q.�i�J*E�R8��8L�ܚci�NUܭ��N�)V���ȓ$wl��b��N�&������1%U������"aۈ�i����(}�ȓ$���E���{��	#Ag�Z	�ȓ'd� I7���j\��A�ӻj̢̆�*�,8��`�'0t�wF�8I��ІȓW��3�@�w��=˔F˝W^�Y�ȓ%D2��c斻.���D�i����ȓ_U�d`DÔ-
h�����/D}�-��@4�X��K�^���JV$L�f3֔�ȓOf@��dR4d�H�Q�I�(�u����ݑr��j?�a�2��&q̬���/(�! 5B¬��ذ����e㰽�Ɠ�l�b��\��<��
�'��x*'"���Ԓ�+�� �~L)�'(FD�̕��xM��������'Sf �и53�� �	?�fDI�'��,�2BV�C��U�VBX�$�K�'�pC �+BH����ٴw��8�	�'6^!�@�� d�>�[�m��x���� �Ţw��e�xq�C%�|��T�"OA�+F�C6Uæ���"Of����	�DJ���gbV��"O�5�LÌ
���p�+��^�(rR"OF�'��yGxp $E��*K����"O`�ҁ M+r��&MH���"O@T�@í*��XF��@�ّ�"OzaK�̥h,񀰧D�� �À"ON��VJ��B0q��d��4+j�9"O"�hR�;:�H\pr�
�un��"O�M��������#+��L�a"O��X3&G��@{Ce�?�J�Hs"O$�c���o��}x�DD�v s"O|��˦�>p�I���T@	q"O�[' �)Fӊ1yeF�7U��( �"O ӭ��P���>5�օؑ"O\�Q�_�
T$�&�C�I�� 9�"Oz0�oԊL&�|���q�(DC�"OhY�Ѩ�<~
�Uy�`I6���'"Oni��@?"'�E)V��p�(I�"O��d��7e�@yeI�w����`"O~���a��x`֭�2�R�d"O����CA-��t�S��wrT�2�"Oj(+��+E�X�*Ņ��P�ʔ[�"OB�!V�Wm�u��+`v�C�"O�Q��6.���@��	)}S�D0�"O�h�J�%��i!��܅VN��H�"O��sv/Ÿ4��6�	�rP�4��"O�4"���2�0�[PlMtU|�@u"Oܼ�\	wp �S�ǧ㢍R�g�L�<���ݨ5@�ت��#-ƶ:ѭ�P�<�D�Ȟr$��C.��>���@��M�<e�=UUBo�� ;��U�YP�<QT �� �Ƥ�w�Z�v�Y�g�JL�<�R�}�Qئe�"VϤ�q�E�H�<�_ d ��
[t�h7'�A�<yK_�P�{��ȃf!�<pmB�<�w��GY|�Q�W�wTP�R��U�<I#i\�&|b��e�Υe��xh��KS�<QI�5E��I;��&weP�3��S�<)c�
N]p�r�A��5�DQs�+R�<�R��'%��m���U	��Q�<��� �4��e�
!NT8���\D�<�v��&zk0�2�[�(Pe[��@�<��?S�la�d�\;>
L���ē|�<��m@,ڂ<��%�.^Ш!@MZM�<u��&>0}���O��r����YI�<!T�jMZ����߶i=�m�p��L�<�Pս�:TJ��66�\�#"�H�<A	�;���� �ܱ.,~���G��<YSb*e��a�-X�D���LJ|�<	U�<f���'M��T�� �M�<A�*[ w�f�����QԨ2�nKn�<���a>�`kV#R�FA�yz���m�<�T+�$,Ɯ
FS�4Lb�8T��0�[��[���*O4�����y⃍^]b�{�➖'U.qVG��y�-G(NN�����1Lü��UL�(�y���#��r�����	��y,��'l0yS�
4H�!ĠM��y���1h	��װ6^��e��y�����6ʊ�8��]����yrMB�Z���%�G�6�P���`��y�0֒�R痁=cN}������y
� �����E7��A�d(4j�Z"O���D*)���v�(Y]���"O@<+!Q-B�>9��b�1=K,"OVpa�R�K�.���"ٔ1�T2"O��QN_�.�V4 Q�S�LH!"O�"t��^X��W��o>�Z"O~It��7 ���r'��k!v"OԀx�hߦ;�T�q�g���(HYB"OA+��DU�Q�0�U?*�	ʡ"O���O[�XKsǐ��@q�"O@����2f���C���.�[4"OD��.�{frt�(�'9c�1�"O��A�%"(\�ǖVh�R�"Oxqi(r������\y;�"Oh9��(׾wQ�(�M�,I�)��"O���JT��\��U�'��Y+6"O��ۢ�LaXڡ�GA�u�p�1"O� ���qh,<�������"O����K�m�lӡp\����"O�i�$�]�k�|��r�-dL�1"OP�Sv���р�*uJ� 6Z���"O��@c�'g���hF�$Rn�u"O��h�c
�1��p��L�%-A��b�"O�C0��CQh����ND�˲"O>�N 9%�!��,ֳ	/|Q�"O<�jtJ�3C�Q���S*l�0c"OR�h6�K�ʰ��*�Y�9K�"OH0#E��))�Bqb��"w]|��2"O�@�JA4#¤� (��F �R<D��SGa���1�"�S�+�|!!�8D����픟)����P��|�'�7D�(���37����D�-V�T1iu�9D��B�\�&z�HY��T) �4ɓ2�6D�pJ"�H"Iq �&=+���dL4D���d\�N�Y �O*j�\��3D��;��߶T��T��R��P�I�%2D��qc-�	^Q�{V��8lB,�G1D�T�PLӘS�~$�VP)+��A�k1D�0`��0"P8�ÎZ�Z$�	�&-D����G�<��"�ϙ�V©�0D��"�d�E8�N6\Oj�aA�-D��1�,6B�0�͕=	Bt�D�/D���Rf�C[��(��H��`-D��*��t�����G�"���a��+D�ۇe/B:�c��$ 3���pA'D���_8C`�9g�,F�d�a�#D�8˳a<E�0qs��^$&���(Ui#D�4C���*5�,�A蚙rЦ`��?D��P�F�7���	��Z<Cռ93C<D� �'��
z�p3d�7q�^m�ѡ$D���L˚%G�c��<j���K�-D���4U��Ss���hX��r�.D��`dɽT�BF��H�@u�!D��JC���*�꠪̋s�D��,-D��0֋�&�y�m�B�:4(E�?D��H�)S�qVZQ��B^���mB->D��S��vy`��6�#(�����`=D�䳰/�N��M97�E#M������9D�j�3q ��I�(p�8D��BS&���� � ��u��"D�4rB��0]|@l�M  4�x g�!D�x�Q S�%�!����4�T\(%�>D�d)�F�tal�૏�fH�%�<D�fB��
zUj��75ӊ�z�&D�� �9���Dڤ��TW�z����"O���g��[5@a����.�xd�"Oh�& �:��D8t.{�d�%"O��+L9&�����S�MY$Q��"O�Qb��-�J��/G��DA�"OXL�o��o"킲�H;q��Ij�"O���U�ЫW��B,øh�ҁ��"On(��O�I?����z��$�w"O� ����@�!����N}�2C"O,�Pլ�@�L��k�df^�3�"O*���,H�d�l��pVb��"O�0���3��JC*Ӱ]�j)�"O�c�#Ns�M#I �c��1"!"OB(���,+Â�1��C�82:%q�"OJha�i C4Ib�G�D"O�x�k�"\� �ݤz4\ {�"O��4m_�e!��� .R� b"O<DC��M%d�"ކy&�i9�"O�٠��J �hl�" ,kt�6"O���D���� c��.��qs"O,t�%Nނa��t�g#�>w~X �e"OZ��!V�x�M߭Ky&�1""O�e)1�V�yRn-���F�YY^�{"O(��L#rx���*��u�6�J`"O�s$ً^����>K.:�q`"O��se��T({TA��B$.c�!�$؆|-z)��� �.tq�_5$�!�D�6{�$a�� @�3І՞J�!�$ Sq2b��'eHl��`���!�N�|a*g�ەH@��6NA!�䕖l�2q�F(�L⢉crL�eS!�Ė� ���w��4��\����jP!�D�b� x�\u\�T3bI׺@�!�$���h0�6�\�@!c�BX!�$��;���s����@�:���`x�!��/^H%��\�_4�Pj�
6�!�D%:s���3��.c$��֍"�!�$�0����IؗO��ن�]6O�!�Ġi=��B��>C[d�I�*�-\!�Da򁱃�D>TA2呰�D!�$�:dN2��c�e4�lq�g�H�!�d�,H/���I�{�	t�M<!�ǌ��ݸ���(U�䜻�� �x�!��F�ac��� n����.W!���֭
�J�!8JBP�$E!�DO�#��٨�-�)Cd�c���K'!��G�-� Y
Rvs�B	I!�d�%+6�؁6��kG
�(��C�!�P_���P��f.H�T#Q7$'!���
�|�Q�$M��\S�[�Y5!�$\lZ¼���F�1��Qh��b!���r�x2�
���x`�a$�B!�d�
HU������D���1�!�$��^�p� C%:�ʬ2�J-�!���hrؠ�!��PU�J��z�!��K��\���Ÿ;?�,y��&"�!� lBLh���%2Jh򥤑3 �!�ċ1H����J�
4CF){r!�dF�E`ʐ ��C����BŚ=!�B75h��@�Gպ�($H�#h�!�Ę=)�d���z N̓s��!	�!�$1PĨ�0ek�\��qgA��!�dM�n�M���G�z�ڴf�RR!���f��D�vB<фM`�Õ��!�� T��/�N��4뛇HLP��"Ot1�4��C����g�p"�%�g"O��c�Ʃ�2(
6)B�S/h���"Oj���\4����H޳#�59"O�a�� �5RTҧӳ4>l��"O�(s�#Ĳ$6! u��$z�"O&,d�X8���Al��[KF�R�"Ob�%�pj"!��e"C# �@�"O.=��ϙ(Y.9�2�Ϊ9j� "O�B�-�a�Pr�n.<��"O��˄�����b��w3@��S"O���K�@m8=���.1h�9W"OѪ�.G��i�҈c�L�"O 0�%�C�D�Ԅ��-ɏ �f͐�"O�]@��-/��,����VG���G"O�A�O�/��E2���K4��`g"O\�'�m��|Q�%lxR��"O�\
6�(:��w�KZsTp "O\i���J�iĝ{�)q8�"p"Or8��B�+h*AC�
�q���"Of��
�Uڼ�C�	 �j�X�"O��
Q��8E�JmbG(�2+�(9�"O����]�S��}��E��)Е"ON� �ɭ) "M25��@\��x��'�mX�7kC�ey 	�:+�t���~�b�}e�!�S�Жx���Q���y�jé1��E�"��a��q
��yb��#l:<@6�V\b�2p���y� ^hD�91'�	x�.���y�铬?�m0`���#�&a0�"B�	"~lI���9���j�̷_Z�C��%Qx&�壎�иJP�UzB�	?F�J�eN�	�`1 �aN�V�LB�I8S* P���Q����3�Y�^�xB�
O�6�9%(�=)i81�F��
/LB�ɼh����!G�N�HY���p�B�I�*��t��`��-�ZM�S��$M�B�	�!���Ss�X�Nn\�RM�blB�5b�
��! *_Vd���6/�2B��$^!�����DFH�f��9�^C�ɐ��@�EK�h�<l�Q�:clPC�	�pr�A2=h�x9pV�B<{bC�I�?l*��ʝ�ِ���1Q"C䉤\"�����  ~�@9�0c�B� C�I;#�L@�A�@�h�����:�B�	�V"-x�&@&\�[t�Y�YJ(B䉮>������Aָx��'��C�	>t��PUg[� ���I��˰x�C�	�5p���b�l��k�B�xdC䉩r��L�Ԣ�Df���"��$�0C�	�W@�̑��8"芠"@
2hC䉉z���P��&+����Xo�u��ve�$��F!	+&�'�b0`���YS� �V*Y�]�BT�dDW:f�P�ȓe)���E�	&r�N�#�jO��0Ѕȓ,�L�� F���%���ް;!��ȓG�4h���T:���SM�2Ԇȓc
��*����L�6�8c@��������X�Bٓ$2��%Nב,u\��
6��RD�Ś���(��!�v��*i��r%���d���U�:y��Ĉ���ȿT��L���N�ޘԇ�T�$�s�3A���
�Y�^-�ȓV��`�7]�vГ�.�}����S�? t���:��:�h7|&jl"Of�
˂0�P�j5�Y�.�Ȣ�"O�} j�|�T���η�5""O1h4B��>��`��*�$�"OF���oL#:W�0�m^8S�İ�"O���s#H%c����Y4@�c�"O0$���ʙ��)V�~��"O6�e-8D�IbAx=0zG+�y�<Ѧ�OgiP�X�Jjδ�e-u�<Y��x�(��Ł(Y�,m�<с�r�v"�aN�pG���Ff�<��O�0�*q�5�.)�J�H`��I�<����_Z0���!��`���@�C�<��#1)�x�%�S�)G.�����}�<'i�H�
Ta���\k�%y���u�<����J<�cˋ�����n�<!�CŴEFl��,ɏ�l����<i�(��,���g����dȧ8��{�G�#B����
�AT���A�"!~&�!�i�8$f��?�k�	:`i�x#�IJ�X�l�
w��6?6�AU�hA�Q͚d��0{G`JY���'�3]T��6�U�y��-Pp��G�,�1��'X!���'�B6P��Y����g}��E���N����H�o���(O���D�+�:� �ƅ 0ܴ%��V��Ц���4��$W��SXy2N;=U�,K¢�R��4ۅ���^,��!JC�$/�y��'_�e�RL�?X�(qw��BpA�cҝ!�
�)S2"h���N9bYD~2��d����Ͳ��H���Š!p�@�g �+*F��B
�9>��S�a4Io^-Gy���2�?1ݴ��`��J+3�س`��d 
�m�����<���?AN>�'�MsC���5��Q�AH� Y�;X�<��G�t�DL�DK��Zd���۸|r�F3Ivv7�O�eo��:؊!�YwzB[��.�?'��S��ә����D-�W�qO���D�S�2�X+�@QG`>j�� �O�f�@�K;s�P�Y 6��ю��Ǭv�B��ҠN� ���̜!� ��'M��) ҡ�2
p��@�.gWB�FzBb�&�?��i��>-c��B�= P���8e���#*�����K�I�u�(YC�bQ���`F&���dFަA�4�M����2��0.0N�8t�
Sh���7u2�C�iR�'�哵!��	���n�/3����~8X �Rm4�V��C$�h/0$�煁&����O��y��S���Ovkl� ��E�+ڥ����A_�5 �6�Y-[A�ݺ��ϫ �J��	���� �Ki�����%E�ܴ+bi�Oǔ?�=�R�Wy���o�,~���_���X-O�O��s�Z�K����[�@�F�D4K��O����O��ĸ<E�$�W�!`���b�b�>�����(O�}l�'�MÏ����@@�ˏ�[v|��?�j{��ay2��y7�6M8,O��Ce ԟwȼ�H�s��1J�,F�g�]0��ו �|�kU:$������T���s�F��8hd�'��Otr���M	��M���<��Tz��
�mr`��O9�"<���N�lCT$f���x&�йn]�dA�"gi��<:���՟8�'�n��'�
/.�ʍ�@H�:V\���HO�A�Rg\�C�e(�B!CU��y�ګ�M%�i�'N���O�剥J�4a�R�Q�FGPܻ�Hh�*1�a\'e_����D�	ǟpu���	̟48sGR	s���CWC[�(���A7��3F�`�#AQ)(���ٱMC�`�'���;�
a�w���TI����AY� �a��2����W L#K��-E〫/����4��0 w��/��Ԕo�B�ܽKB %��jD�q����s��w�����r�X�Ķ<������Ծi`0���3ɶ�'��nr�K� ��I		�J���M�f�x��*�P�攈�>O�V�}��ۥ��dV�&��Z�    �   &   Ĵ���	��Z��t�D�8,���3��H��R�
O�ظ2�x�I[#����4Gf��BU>[,L+�l�(m��bZO�Hؙݴ���k�0���Iz��	����Y<4t��Q�&�҄X0l#�ox"<��~�^)Q�K�H]4� 1���>V��U�̳����cYX�F)?���>Y8H7M�X}�"/Y>��1q�ڧT���A�J���9g"[\y�f�O�dXb_��uW�??a (�6�����"�*td�3��dЬ��vd�*/3��
e��bٔTQN�4qA3ON"�i0�"a����Ehh�3��|r��|�'nN�$��趣��I���eNNоXw�s��tቊBl�S�g
E��y� Ƽ-�8mS�ŏ�OH�������$ �a�>�r�!_���Ls B��v�+)�"<1`�:�I�|NL�DBE��X�C��j��7��	�O�Î�Ğ������fQ��a5�-�"�t�K^#<Q&�6?铇�$A ���'+*�5X%�Mmy�M^S�'*�5�?ɓ�&�N���*��#7�x�2J�.CYN#<)b�4:E���לJ50q�&ڱ+̽�e�^�7�1O2����Z��Kр�K4؛Z�^d�W��z�dx�&� #<���'�Q�Vh���"9��,HPOΐ�q�IV��ޖ{���㤻iX��t�	tj��Ɵ./����t�ܱ�㞬9��Ʉ5��m�n�i'��*��<����]
q�'+f�Fx�js�'����GM:\�����h@��',~��@ ��0��Ia�<�#J�8'S��%���Sdi��+a�<��+�<���X��	�8$ir��^Y�<� �e����5)f ��.�{�6�Js"O��at��m�x8���]�(h��"O���� K�_#�=0��C? �b�"O�|�"U�p��(���{jp�@"O>��m9&$bE�2 �1Lf>�p�"Ou�*�/w@F�ʖ�Z>%x�"O��:�E!+lx[%��7�<��F"O�82��/i�����Z|�i�"O��jlӂz��У�MU Q(�"O~<iQg��n(<��֣����ps"O�Y+0� �#1&�P$��=����"Ox�קZ(_�܅cE�@g���"O������r��9 s�[<��A"O�Xg��}�D�#�\���"O��'-��T�Ţ�
S�R'|��b"O�	��iG�rH:��f�Q"Oܰ�ЊK�2�d����ƂG�8}Ä"O�s    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��     �  �  �  H*  �5  �@  SL  �W  �b  nk  �s  �|  R�  �  k�  ��  �  _�  ��  �  0�  {�  ��  #�  ��  (�  ��  ��  �  a�  >�  ��  � I = 
 �' �/ .7 o= �C �H  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H����<q�I�$3Oj���O�~��PeZ_�<�6�E�>�acfY�l�����S�'b�)ڧA~9��A86��%��(�0�b�ȓC��s䇜�`�f����|:��'%ў"|
�`8tڬ`��]cN&��e*�z�<��
�#b$�!��N�k��uO�ty��'t��X��K$3��" �M�pr�';�	��}
%�p��[v�<1�X� )�� ++�&��`�Nh�<1&L7p�5�1��J��E�jNg�<�φ�_TB9Q�� �Xl�q��͟�E{��I@�}��d����}��	#*	��B�I�}b�r��Q*-����4��7JH���p?1$�ҷ9�*�`��3����wDX�<�j��K9tH�Z<�n�6�W�<y��i��鲇*(DR��S�e�8�y�ᅾ��ـ�f�=��x8��Q&�y���1:Fp���KD��� %	��y"8�M:��@lbV�)d	Ӕ�y��[��Ը��M�g���CN��yb��1�
�"��[�<x�BI°�p?��O*p�M�>Jt:����VT��q"Oz(En9k��ˑe!�߰џG��G�v�c{V��``<H!�B�	;�}!t/��f�3��L�{q��hO>�  ui��r\`��!#�b6��C"OV�pA /�ڌ�@!�PTDru"O��fo��>�L@xRm�!;���"O2"�=_�h�l��_�,�C"O�Z�
�Su�	�U�, �lT1&�	T�����׾�C��
�Z� � 6ꍖi�!�$�,>�� �k��x�\\i�bA�
1O��=�|��ΙQFh�5�N�NcBгKZ�<q7�U���T���=�v%cs
�Z���0=ɳ�ܙh^���W��--�8�l\U�<e��nG̬�0kQ�-�R�����P�<�b�����sS��876�Fk]P�<�2#V?x9^�;�&�8r�ޝ�7G�N�<Y!�Ά;�2d�E$nR��A2N�<i#�Ŝp��+Ԇ��T���J�<�V�/��(�+i��,i�']|�<Q�@B�F����:��p�TKd�<��GE+�~ݹpI��q(���D�Ʀ�X�'(��(vbL�����߫KFh�9���'�y�@BQ�?#�����U�4��3�'k^8��AR����L�d��py��$=�S�T�����,$u+��C��y�@��5��p�IN�P����PyR��4S�a�.H�<�:JĢ�t�<em%d�ؘs��ϻ�<�S	m�<)]x�@VKh
FQp��=8�܅��Vy2..'.�ZC��/o �ADK�Y�<qç�8ւ�#��
�*�!�  �X�<��� ?(\x頡�^rUF4��)�n�<1�"�/N2�F��
\*�QÃ�E�'d�?A�l�>=/rY#0
�;�v�'A&D�PA�gL
0��9!�dP���h�<mZP�')ў �7�oض�� ?�-i�o<�O�0���wG�J�� 	���"yф@�'�}�
@	Y�ա4X<����4D���䒭
Qnms��\7}.����>D���sG�`�P@�i� f��a�;��-�Sܧ�v���βY\v`{w��&fH�������d�&㲈K�$��>��Q�D����A�h�a�ĸ1&D���n ��Is�ۛ~B�X"�
�6d�<����,bA�'B~�w
�5Pa�	��I]~���# ^��s%��4NA6%�y�%�\�>%�RS�>�,�������yB��yL�� �I��G����+Ƅ�y�J<JTmB#nSt�ui����y2��fq����- ] ��gd���y�̌0t�\��/X-�N�▧I��y҉��N�ִ��99�vH	7N��y��{�L ҪC�0`��vI��y�B�1!��i��Ҩ��yK�%��y2!Sd�����B�����y"�W*X�r ̀#J9��(ޤ�ybFZ��&I�u�ױ�Xi�C��"�y,H:}D iȖ�^+L��bꞦ�y�n�l� V�OF��M��(W��y��<CƑ��ڊO�&4+�m�y�N�Re�FO�*�uZ��E�y�R�k�J	7�ӟ"I��!ƫ�y��?~���y����i�� L,�y�a�*j�X��O�9��(��yB�)lb�#�MM0��B E��yBG˒|�BݢE��7��0�C��y�V�*D����b��@6O^��y
� ��J��E%��e�Z����e"OF)	#���=| �����ޭ�"O���2��8>����h�" 6"O�ȸ�.@ �@��R'4��D�"O����1Yu$u�T�	* �A�"O� (C����}X@%A�h��"O������%�����?M[�i��"Op$p���<#@����(T��3"O����&8x<�JY�,:V"O< ����Q^�*�(ߥEfD��A"OjP��.M�<�	�t']�Lja��"O�Y��ٴZ�D[�&ZZ1�i�"O���#��ai���%&�W}n�a�"O�Q��C��JErUJ¥ݦCw虻�'��3TjCT.�i)�!�82����'����dJû}�t��G"[]eH�'٢�� �4dv��d��]��'�r�p�\�FhQ���M82i��'��!���'t/4=@2��
3�A:
�'nt��5#��Z�p��q�2�F�
�'a�툦�ޔ6���`rg��%-2�	�'����Em
�O!tQ�1��*$�|��'�D���O�p���4����'��Q���!�X@��gQ�0,By��'�z�3��]�S��a�Dh�2���
�'JҀ��i�.� �ĥ�=S��tk�'R��� d�2����4L	MZv��'�r����$d`Њ�o�C:�ٙ�'�̡�H��r�D7�90�촡�'@>`*  �*�E���])t��'� ]����*Π�`,A�ilvQ!�'�l��`�
��*@�'�x��'��d�SjȑM1| �����4����'@][�L�$�\���1VDPM��'�ٱ�b̶u��6h��F��%A�"OT�"��@ʰu���å�n�Pd"O�LZ�+�~UJ�#0�U�1��i*0"O���gF�q��@��Aɀ+�����"OB�9TG[6[�@�Wc�ks����"Om�7�rQ��X�"C.p�̼��"O�`QlV�eST�R<��I�3"Oh���E֒l7,9�����5���"O���vJ��T�"�n{o(��"O
U{�DRVn�%``��R)��"O\@I�e�^Cr��U� =l��"O �9�HT�kVRA�f��R����$"On�V�B����	J&_����c"O��x�KE�AxPHD��xX�"OEjC��"h��ٓG(H-5��1�"OdIy����\f&,s�	6�,��r"OH3���@I����ʙfL#�"O�<��Q('�T�	���"4���S"Otݛ!MS�R{>6ブ1?.d���#D��a5�V�]��XbԀĒu��:V->D��aS�R��: �@�p�5��	=D�(�C��V�(M�t���t>v��?D�l���l8n����-L�\��=D�AL�!=�Pi���f,���N<D�lەaAx+�y�D;m0�x9E�8D�`��=�����$�}��h�$D��c>[�:���`F�L�*O*ѹE5ZF���TE6R���"O��K��(�@�D	E�<;W"O����l�l8<�ѣ"O� ����Ꙭ	�<���B����"O0u��M�&_�ta+ 퇣L���rv"Oz�a&'��daH�j�E�f~�qs"O:�ă�-�p�a'�xR��rp"Of����ݕ}�Ɣ:'�Y�V�:���'���'{��'w2�'�B�'���'�`�:�b�t�h�&��C�U��'FR�'s��'R�'���'���'>XE�P�O�F�
�9��w�=r��'nR�'�B�'z��'���';r�'>�H�!:����P.�2d�>���'���'���'l��'�2�'��'��=�@!�J�Yh���h?j� ��'p�''R�'��'���'(��'}I��rDc�n^�C1��C��'(R�'���'���'B�'*�'Pά��MB�g��:@˃�"}�0�'���'��'���'��'8b�'���Q/09҂��4��Ȳ��'z"�'���'���'9��'�b�'tN8�@�1����o�tx��2�'EB�'��'��'o��'r��'Kr����I�l,ȓU��RE�'�r�'�r�'�R�'���'��'�	qW	"F�#vL�o���X��'*��'��'��'3�'�b�'$,�h6Έ;'�R�� IJ�^�N��s�'���'�R�'p��'�B�'���'��Q�u*�;!<�J��&�D���'���'���'Y��'��as�V���O4@ 6�@+԰�[�BD}<��_-"��?�*O1���
�M��	t�œ'� 5W�0�߀I\�e�'��6�<�i>����\�� ;l������C�A�Qc���՟����#���n�]~R?�:���C�)�:;�p�(��=2D�VᏻP1O0�į<ɉ�I�j�����N3d�}0G�ҁ���l�\��c���5��yw��CN�wa
++����(D�W2�'�>�|R��A?�MK�'��-���K3�^�raIF
XN�M�'���蟠���i>��I/8+>�eN��Pܘt�ğ�~����<�H>��iJ�$j�yB*R�F����Ł��|����L��On��'���'��d�>���R~�X[s䒇QNlaxpCX~r�'��`�����O��d��v�@�+N6JI��DSp�(`b�4X ��Kyr򧈟�D��@]�|�F�62��u�I���������c4?!d�iw�O�ƬqRFɸ ��	y�R�B/�9e��d�OX���ODQ�keӼ���Dn���ט�*�E��CSu��"��B�|�D�O����O�)�O����OL��O,\!�&D	�P����J&\&T	����OR�$M�R��K���OH���O�tlZ 3G���ß 0R��*� ai4L�T�����ڣ\���	Ο@�	���S_���'��H:Bq��q�i��e�����c�^5i�O��$�!Pǂ�J��7"<�O��U�h	a�Z�#�Ʃ
�j�}������?����?�� �*��(O�n�h�b��S�(��3���+
� ����Ɍ)�PM�I.�MC���D�O��'�2_���R#ӕh��X U�̓n� �H��/dW�l��<�����J��JY�*O:�	��z=��E�@���x"`%9��p�9O��D�O��O ��O��?�Q��t )�4Gڊ6�h��m������џXڴmu|�ͧ�?᳸i�'3��Z��H�&<*��(�r0���|��'��O��w�iI��8��}'���b� ���[;Obb$���	�q�r�JB�	Dy�O���'�!��L��R&�^|��C���K��'3��M�  ���?���?+�>P ��sĊ�2Ĥ��k�B�ʅ1OJ�DLl}�'_r�|ʟf�)�M%�^�蒬�"q8\�@֚B)Z�ҍuӊ�����T?aL>�Ī��'�
�K���q�`m!�IN��?9���?���?�|�.ONn�&3ȭ���&�<XNU,خ��G��˟ �I��Mc�2`�>�,9���C���+���x���6pX���?�1����M#�O�abc.���V�� 3�	k�|�pIٜ�8���{���'r�{��^�N)�0�6���V���*H�h��7-�U�L���O�d7��-�Mϻ$v�l����$������L�B�և�?����S�'2��۴�y�G��N\0q���3Zt*s���yҥW�	�������O���Z6U"�A3iP�ro*��eǲgn&���O��$�O�ʓOK�V�W/7#��'�I�o����R�H�B�62�O,��'���'��'��|��E��d�#�/W@ъ�O���Ed�+Ft���󉖫�?���O�)�vM��Wμ��U�p5�H3��O���O���O\�}
��LY�1p�Kѩ�\5i�̐4�dm���i����3&��'��6�:�i����<`l~9��+Wkr���h`����ß����{�2LmJ~r�՗\tp-��.R�,傕�ԩK�T��Aa Tm�%���|Q���������I��8���W�p#��gCˈ|N%���py�`z�6� aj�<�����O*�5xŮ�i�
�!#��y �2��>���?�H>�|��D�	gy	B�;&� �_�^��q�t~@�D��m�� i@�'�����$A� !Mآ�Oя�����'2�'���'��P�l3ݴ��;��dR���-b�  ���B(�S��r����|��'����?1,O�!Y��Z��������!n�P��`�Q��7�d���##�]S��OV��'������ ,�s��R}��U+L���h�5O*���O@���O����<�O}ĸ��-&Ɛ�	�&L,K ��ڙ'�R�'c"�{�:�"�İ<�i�Q��+"�Z�|��dN��^'�bf"�ߟ��������Ŧ�͓�?qW��%G2�qd���4o�y;2/Ȳ��;Q��O"�I>1)OB�$�O���O MXS��ݴ,¬T�m�N�J�M�O���<� �i�|��0�'��'$�Sz�,YSg�Hk�f�	5M\�e��=��IßD��w�)�P"]�wQV�
������ h�0%�E�"�G7�Mc�O��ʠ�~�|R�Б@�f�s��QRTx���]�,^��'s��'k���T��Qݴ0����,�FV�p-��J�j4��(�?!�Û���u}��'���D3q.��-W�!��T�t8�
�����'@��󱧒�?�pZ� Xp�׷6>��)�9!�L���jp�h�'�"�'K��''R�'{�S �8!ӑA�(w;��zE��"eT��a�4 3�,��?9�����<���y��E5ؾ�k��Dqj�jd�\���'�ɧ�O&����i4�O�!���!/!T�B��W+XP�d\2�bj�a||�Oj��|B��R�|pt�JH��X���O�Fa�����?���?�.O@-m�&s������t�	 Im�C�JC�4��egO��[�0&�H�I�����O��2�U�%���4%��3㌜ф�S(��	*'�9p�IǦ�O~�������	�' y���B+Jʹ(`1YI����՟���ٟ\�I{�O�"�B�G������ c����(ne��	s��O��������?�;;>�{�)�؝2��Y�z=͓�?���?�'���M��O�e��W��2�� 3��3%a;N*���o� 1�O(��|���?Y��?�ܦA+  !2H����9E����3�Qgy��k��%$�O2���O
��6�dגX\��#l�2�p�Rc@	D}�';��'ɧ�Oi�ԉ��2-�n=�&���t���a�m��f���:��	5U��5���<q��	L����BH�6q�ܠ3E�?�?A���?!��?ͧ��ğ���g�_� ;�K��e��%�#�Y�,�@pK�+���޴��'����?���?ٴ L7=]t�8��@�3�x��`�3:,(�Zڴ���׃N�()��)���,ӥ�!�,܊��]�
�
��>O����O����O���Or��@�(RgڭO!D�0EA�p�`���͛ή˓�?Y��iO*0y�O#��'��T��c���/3n�z]�ffY�v0��?���?���=�ܙ�4�y�'�ظ�uI�K�����e��2��y@��D�@e��/�'��	ş���֟���"9�@Q�l�j��vf^�*���۟�'��6���6M����OV�$�|Z��@�a�����&K�. RHX|~��>���?YN>�O�z�R��߃IWZ�y NN�sZ$RǪW'u4*rE�i��i>�� �OƓO�<�p�э;Od��wgۓ;r����O����O��O1���4#��#X�j�4!b�;Ɯň�o$o�ա&Y����4��'ʜ듇?�2D�>Q��eCG��0�h �����?1�%߼��4�����H��U�'��S�X(%k�HK�UÐ�:3�pb�	sy"�'��'���'�V>�[Fi�5i��	�l/V�I+�Ȓ��M�7&Ɨ�?���?O~�r1��w��XcY���L�a[7�����'b�|��4iܒ(2�61O�q�d�B����õQG��q�9O����˃��?Iu�,���<ͧ�?q�(N!A�,�2�/x'�l�­ɥ�?����?�����DDۦ]�D����	�d�K��
�A-��W��l��d��v���蟘�?�d�� m����C�.���˰��f~�#)�����b"��O����I#�2I
H4���Ќ�-ܑ�����b�'���'K�s�1	�
%�	����gDX@;E�RП��4}�����?YS�iF�'��w���-� Z� �R�C�Ϟ�C�'qb�'=R͔N��F���]ۚ������
�!�:D��H�`�$�	kc�|�P���Iџ��	՟L��������)H���G��N9"�CLPy�/�N�`f��O���O��?�a'りC�y��E�,3i�H��jJ����O��D3���U�R88�R�ΫMq�`���Fq�ኄ�()����(��'[R�%�0�'oʅ����$n>�:-2���k��'E�'�2����P��jڴqN��Z��|�����B����`D�:0� ��Q8����K}2�'���'?~��Q�D���޴d��(9�gP�y�b��޴����l�V�j��6��v�.���`���¶���+�߯vl���Ob�$�O��d�O���+�S�V�2��ǒ!XUJg�`�'t��pӈ���?9Q�4��O=�@ʑdPerON�!����L>q���?ͧc��� ޴���S�1k���!{MvE�7[�e��g�S��~"�|�Y��������	���g֟	��P#�eJ�µ���J����I{yrik�bUZ!��O��d�ON�'��C@h�7c��1���K<�@��'�&��?����S�d�͉}.,z�Q6�
�����L��$���ɫM����S�'��$7��ə/�H��F��*q�莾�����O��D�OH��)�<���iH�-!�r�](�n��D9�Ly��>@��'�6M'�$�O�m�'P���Jh�M�I��`8�ᆬrN��'ޒ�	1�ik�i�%�BJ�?I8U�� ���W��8���U�8m�}��6O6ʓ�?���?!��?q���iT<zI�p4!�5�z�` U�]e2uo�-J�$�����i�s�|J���"���N�[�N�� (U�.��0,�O��d$��i[Z��7�i�3G&�>l���n�`��iyc�0�Ã >-��+�V�yʟ����]���!AW�'�tM��'>6�υ|��O��D�)yJ� ���]n�E ������ ��O����O��O��(a�^6�\ȓÈ;<O �`��0�0"�����A�j��
�2A�����2��3��Ń���&1A��"D(Xȟ8���|�	���D��'{r�۷�^���l�sk^�,L���u�'p�7G�azj˓&-��4�E#FA�<z�0����'Y=N�k@:O����O����=��73?��I\�����-�8�6 �/D��3��z����J>!/O�)�O^���O���Oye'+5�ԝXf���Of�i� �<���i���d�'���'��t#�L�2�' �Tk�,�#�^`����P�P8#�A�>��������'����<7�2��A�49�PA��TIv�$��*�Y�	�SC$�y��'-j@$��'D���#�ȏ4w�L3�.B/2^�1�2�'��'����$Y���ٴ �\t9��)0�=�b�
H�ҁ��_=�ДΓr4�F�dH}��'h��'�����>��	q���s����5�~ϛF�� �RAV6D�������qȀ�E*������6�ʬ�":O^��O��D�OF��O8�?`�*��YR�M�u�K~��$�O4������RAy�c�j�O A!B㇖Z�0P��7�~5��3���O~�4��t�4 a�F�HP�Ј��.D�|h1��o������N\ ���������9O�m�oŖ`cR��D�X�:�ة���5�M���T��?Y��?Y/��}
A�֐��H���'
�+c��,1�O����On�O�S�f�%�B΍�(vq��勎tf�h֋�U�f�) �uy�O P}�	���'�����N�1��0(�"A��`ԁ�'��'db���O0�I,�M�G&�?�$pp��(wdD������#t����?��i��Oʑ�'���MO<���%/V�GF��; �k�I�E]�o�j~ң�%X�fQ�S�H�IY���2n\.<��!��m�"��IOy��'�"�'b�'|�]>52���h��Ma�)�0���F�-�M������?���?aL~�cᛞw�8�R�N�1�Խ"�/ǺAj���e�'B�|���*�m/�3On���g��W�̍�M�&���E:O�9��ʞ��?a��8�D�<�'�?�Yw�Pdq��R;sT���� �?)��?i�������iB��h�	�@/,fM��/��l���S���
h�?�"P�L��ޟ�'���r����%�hv����5_f�	"h��,��b�ۦ�SK~�ᥟ��I�SDA����a��@�IFC�����ʟ���ڟ��`�O��gΦ>�aʱ��b��cD�1p�~Ӗ�A`�O��D�٦)�?ͻy���q�(x~ݻ��R$�P��?����?a�k�M��O|b�MU��
w�A%O����ܫ;��T��@��O��|b��?���?���Eu���p�.5JX�d�ݭK���3.O��mZ?�lQ�I�D��[�s��D�".CH%�O�Fj�#����d�Oz��>��>'!Q�FC?/���I6d�h!��0��I�l�D5��'j�m$�,�'�N�"5�\&R �X�RkC��E���'�B�'�����tY�l�ߴRB\����F�95i�-thd=�g�Mj�����F����|B�'�&��?���?	�a�>���z���+B>���R�,&��ݴ��$O f��y���o�N����!S@��ѱjI/��!`D�d����O���Oj���O���#��R���+�)on�Ha&yF@��	�� �	�M�2$L�|���1ʛ��|Zڤ9`@��[�.Q��j�#K���K>����?ͧ2�V���4��DO I��"lM�x�R�8E�<u�|	!�
�+�~�|�\���Iӟ�I��|�C�`!L,X�T�6����U��"�
���-�Mylr�hdʲ���h���O��)��6a80 �V;�b��Ȭ���x�5O@�dMc}b�'{�O�I�O:��i�
<(Hf �5rw�x;�E��-�%���c��ʓ�Z���O�)
H>�
��w��9��C�(h@2#ό��?1���?����?ͧ�?����$���;�!��h5�$Ӣ)bZi�-DGF@ ���l����Д'��Z����;��XH���N=����h�t�x(��ϟ� c�[Ϧ]��?���0E�p���f~��2Y�I�7(Ɲ=�u3G��,�y�Q�H��	`aB�4~}��zo�#����4@0���?A����OR�6=��A�)M�1��Z�x�b}c���O�d0��	����7M|�h20��^�t�[�Kf~I��Em���J:uj�d+�D�<���?�cOS�����7nS=�v���?I��?������d���!����?���ԟ�rt�D�ɢ�@�\��9zY��&���	(����Od�d�#��S��IVdY�w T� tx���ɒds��zp�Z@2�D�'J������`��' m�#lvt������]<���1�'�"�'[��'Q�>��%��,�ǁ��G-sf�I�AX��I�M�
�"�?���e_��|R��y��(/s���o։;)t�B#.�y2�'p��'' ����i���
�����۟� �K�N^�3%����F�
�~43�3���<���?���?����?y��;ƞ4{�,J6w\ ��ל����q�!Ɵ �Iϟ�&?-�I7S �x@	U�B4@��V�6Ҭ��Ox���OޓO1��q�?�`4�K�J�=��c�=i,��q�<��E�z���Ɖ�����Q�ֶ�bp�U`6`��@Ig^�d�O��D�O6�4��� ��v�D3��l�9H����i�szʍ"�b��#�b�b�>㟀�O4��<Y��-#��2'�� r�ie��#��޴����Y4B�A�'}�\��Z���6�@�&h�!6���c��]}�d�O��D�O ��O0��>��\�N��͕�2צA���D���X�'#�n�¨��?a��4��C�dYY���3,ƩB��C&Ka����(�i>�1�LΦ��u�΂ sd��Ó�<�f�6�L"7�'��%�X�'DB�'��'�t��d�^�*!����q�x䘡�'BV����4!3�l���?�������C���ku�+([��8��C7�I0����OL�d>��?�uIS�y�6|kRm���,���nE�_�4A�0 �&�^��|2t��O��ZH>��F5!�|��5�A�a�,���j���?Q��?����?ͧ�?Y�����Ϧ�QJ�	�"a�$̝�	�#6(Æ���֟hq�4���?��R�`��8&�PŢ��SFU0华vqz�I˟x�"�XЦ�ϓ�?�JCF3��i��dӢeE�ر"˓=�D�A�9�d�<)���?���?���?*��h"���L�|�� �"�����ɏ�1x�*��X����<%?�	9�MϻnF�+a�^
g�
���%O�m����?aN>�|���Q��M��'�h}s��eŚ�	0NU�,i��'n`�[6�؟�B�|]��I�����E�!!�숏mt�4h����>4p�&�_yr�mӀ�Ce$������O:��7@E� ��d��cƅJ%�4�2�D�O��'����>䥸JԪV/"�iG��n����O ����ޕ�T)���<���~U8����?y�A�?o�(@ՄE�.8~EF�۠�?y��?a���?�L~�u���?q���3aEV�I���a�BТ,���z�F�Tb�'�|��y7�k4F���%M5fӠ `T%l8B�'�"�'����F�iZ���O�A�7��(H�k,��Mdⴁ�N�>��-s��ÿGg��N>A+O���Oh��O��d�Ob(�R��EE~�dL׭F
��2Bm�<)d�i�F�Z�]���Im�ޟ����[1"����֫Z��}�6.C�����O���3��)Q<u�8ѱ#�K�$b�� �X�g����>�*ʓc1*1��O��J>+Oh� %K���90$��DJ8� �O���O���O�<��i��H �'jDP#�Q'�ܩ�S��,YI��'/67�;�I�����O2����� �I<(�s��$gh�I�J߆�M��O��������k;�	��N̈T�XVx �2�̑
���1�7O��D�O����O4���Oz�?�k�b�c���Q.P�h��tB���d��͟��ߴB�F��O\6�<�d�D��qf�,K���� �TҒO8�$�O���#S�7�8?Q-��18H�@j�JAT%��<I� ����t'��'���'��'hp�prn_?@��DiN��l-�yX��'�BY�\ ޴�<���?a����${#\p
��}�|�I3^*������O���4��?Y����Og6<�Ġ�+u~�����5iؐ)���J"��|2���ODzM>Ia�z]�xA��)^��kV�L0�?����?Q��?�|z-O&�l5+�lE�0o�#�=J@��|��Q�c�TyR�cӄ�J�Oh�$4Զ4�/^w$�X��̩u���d�O�p��yӎ�)Mų���B�O_蹢�L9��4
����'���q�'�I����	ğ����P��a��iˁ=F�*eK7.x������F��6L�K�f���O��$3���O��lz�����Z���h�F�>|��(��M�����K�)擆��im��<�&N�"
�n��lZ�v��E�ckB�<���^.I̮�IL�	eyS�� $�0�lI� �mB�j.'O�4m�
G:R8�����ɮhr<[ #�+����$�� �4��?��Q�<��˟�&���t�Z"E(>T�rBNWR41�7?�����HD�a���'
�F����?q#Ǌ�4(��A�@c��#��G��?����?���?9����O��RR�×4��$���ęe�6�+���OL��ɞXMF�D�O��n�I�Ӽ�l	�Z�u���U�PP*BO��<���?A��Q0�l��4��$�=4��Գ�O-���I�s�>1��)@�b��B�|�U����ΟP�	џ���ߟ�À R*R�b��6� p�O	Sy�	l�t���O����OB���G=	)�{T�K ��p��Z�:-��'���'�ɧ�O� T+�F���a�p��:߮�A��R����O�]Y�b�%�?�76���<�@��R�fR4H��su�A"`Ir�����Ř��ş,�b��c%
sd��*k�����Ut��4��'��듕?A�ӼK�l�5X�P�F	34��)�r�ªtͶT3�4���ʕ'�z4���T:��^�NK�@\�a��&d:d� '��$�OZ���O����O~��.��'+N����
?y�.be��n m��ߟ���.�M�T�K�|��e曖�|�O�(�yz��
?�"}s�k]�F��')����dGK5C��&���]�� �Fo�-L"�3f��
L�I�IB��?��;�d�<����?a���?���"��{c�ڻL[�M8Ԍ���?���W����(؟�����O�*��3������#�OP��'�r�'Cɧ�I��q�5� �O�000�3�ځ������|�>6�1?�';f��IF�>�t�"�!A� =�k�F������I����	��)��wy�.j��a�i��������N>6�X��cn�:��˓'��$O~}2�'�Td��!M��G�Kk )w�'J�W/d���� !�kH�~ �$�~"CB�� ��@UF�/$`�z�$D�<9(O��d�OB�d�O����O�˧a,d�����?W��%hAeߞ0)6%��i^���Z����s��˟\����� _�u_�<�r���nI2��.�?Y����S�'?���2ٴ�y2�<�����/U2��6��aHhjB����$�,�'$�	 	��T� d�=/,���I������Φ=Y������I�`��nP�}d���`��U.D��c�G��m�I�X�	H�;Ĕp�K͗}k % ��'SF��.�b Z6�ʸw����N~����'J�~< ���Μ8�ϊ$+`�&il���0�גs��1����L])$��'T}��fz5����&e;ҙ�k�k#�|30���.�d�Kv�L�CDa{؞��᎒(y�&L)� (;b��@.k	�iY���S�I�s�C�к QW#��?^�A��ǚ4��,!�	� ��5D��N�{����c�@���B ,��*��ۖ�΂>���j#��8a�ܿg��\��a�T�P�����(t^-ҵ�d��ۇB�m��	c�g�yU�m�����_���$�<Y����;!���eɌ�C�'jV�LQv&�V}���X��'���'�W��g[2[w&p`cD�#M��J'JB+���O��?I>����?�d�j@P��q�ǚO�3G�@)!n��<���?������P1/�TY�'x)��d*����A#�DV/Lw�}mqyr�'��'xb�'�FU)�O`�yWE��:�Ud��?:+�kQ}��'H�'B�I��������]:^��{0��#o����s��&'�BTo�՟�%����՟I��Uܓ*ZI��B�)��x2d!ӥЄ}m�ԟ���Vy"�Ƀ-��'�?���rA�.yhN��F^�n�Ld�M�6c6�'���'Rv�1��'��'����/z�45q&�9!+���K)k�V_�H�!���M���?y����\��X�N:L�:��&6Icr�[#Ua6m�O��d�5F�(�}B���*��dK�.݇�f�ben������@�!�M3���?��z�]�Ȕ'�\a����B�<�(U��0qt�#�y�n�!���O��Ox�?��	��ĩ;CG�b��%s��$�����4�?a��?����[��IJyR�'����brp�YR�_FM~����h��O�E!:���OH�$�O��)�d-Jz: �ǥ\	F�:v�צI�I�L���0�O���?qH>�1Q�"f猆|�B܂�ć�]���' ��y�'*r�'?�I�K"D�Y�$<����@N;C8ݓ�g�/��$�<�����?��U������	��|�����X�dN���䓁?���?a)O�P��O�|����{��؋��G�I)6h�@I���'���|��'����m�$#�$l
E-�?��5�VӞ+��I�L����X�'��-�`I�~����p��c�YFm0i�5(�|���iY�D��؟x�	�a?����dH[�+��\�*�T���ϟG����'BU�*!����'�?q��c��!<�Li�B�Kj��2���ͦy�'���'L2�'J��yZcŸ��ȋr}L����@p ٴ��D='�}l�����O��iG~2	I�8)�ⅻ8DJ��)�M+���?a���?Q$_?5�'��s���2/O�v(@�T�8<-K�i�R� ��'5��'c��O,�)�2���T��A���>H�����@�>d��	b"<E��I��X���o��|"�'��Y��7��O��E����,O��r�$�<N��=K���=�� ӑ��6(1Dx2�:�ݟ��j��Ub<Ҫ�S�)�k��umZ؟�R�euy���~�RGȨ4h2Q�u�C/PKD�x�޽JvOhu�$�O��?5,��DF<\a�B�W�,���H�:�@,Oj���O��t�	t?	�G�!o��I��n,W��`pA�ܦ5�B*���'�2K��:���O4b�Hd3b'^R��(� �����'ER���O�˓y�l�= ��a��Q�p*��#R v�O����<a��s���+���dP9;���v
s�ڀ�Ǻ@�Pao�r���?Q.O��!w�xbD��ZNYCCL'k{��a�0oZӟX�Igy�%ȑU�D�����k��(� ��,ǩn��#lz�'�������	G�s���
8��m���M�ᒶ%�)HT6��?i���4�?����?i���*+O�O"O�T|*�\.��Q`(�-����'$�I�<Ɛ"<%>!`�AЦ+o���Vv��i`�t�,<�d��ᦝ��ş����?� L<�'���cI�wc��i%�%k^Bq��is2�'�r�|ʟ�$�O�����"�n�c�ۧ`=���G/Pߦ}���t�I����K<ͧ�?Q�'��,y�MW	4�P%{����4�?�H>yU?��͟t����(y���Sd�� ���������o����I��7���|B����z�� ,*&L��Z�!"��oN|s��x��'������Ο̗'͞�v-Ÿ&RM�B,�NOH�$d];`?TO��D�Ox�O��Ӻ �?+����Ǆrh���������I[�����'=�̗�T���E
+�([�o\�}��}ðO���&�';��D�Ov˓r�Yo d���e��{�G�cV���?Q��?�*O�A��,�b�ӱ��h0�MƖ �V�x�]81)�4�?�J>i*O�i�O��Ox��#�×06A`Sᑝ�a��4�?�����$N���Or�'���;~L��ʚ(Zz�;��R)����?����?�"`��<aM>��O�L)ś�ZRB�Z���E�F��ߴ��D=n�T!nZ�$������������a��ς�Hܜ�4�1g�h2�i��'"89�'K2[�l�}��ðZ�X�0d,!6�,��d�ʦ�0$l��6���I�H���?�#�O,�Âi6�
 U&lht�N Jp[E�ii�[�'�T����L���Cӣ�^P�%��J�6����u�i]B�'��� sF�����O��	�< 1ȴ쉏D��z���X��6��O�˓L��S���'YbޟN�0HA�NwxMzdf&� �KӸi�O�2Iw�����O�ʓ�?�11����
�r��LI�����'�!�'I��'2B�'�T�l�'l��O���PE�\6b�Y���h�d(�O�ʓ�?�,O���O�dS.hV�1�ElD�7m� ��)�j�xQ�5OV��?���?Q)Ob�t�U�|
���8�4Hpƛ�F�:	3�!HҦU�'��X�P�����ɁX��	�+�~�{T�-'~��p�[�) �ۮO���OX���<1��/'�S���{��V���؞�%p2g�%�M[����O.�D�Oȭj�;O��Y�1�,mX�����$+$I�E�d���$�O�ʓ.z��X�]?���ʟ���4ly��Yw%��{�lM��`��?�p���O6�D�O���A�4��D�|�����4O�FDB����3~'����㗡�M�,O�傂�ܦ������I�?Y��O�΅F&(�$N!Il�`�o�I��^�F�'cX�Ø'� ��<���4�߿"^�X���G�yݜ�͐&�M��A�m�V�'w��'��$b�>�+O�1�HO
���E��_�X�@C�Ӧ%s��t�$��Py��i�O����b�x��p5�X5tH��a�Uͦy�	��I�;h�U��O��?1�'߂�����5�h1����8J� @�4�?���?QB,��<�O���'6,/���-�?��i�׬�RN$6��OZ�Q�GBy}bT�0�I@yr��5�"[���D���2~��������M���6	���?A���?����?�+O
��#M��4�נO�Z�ͫ#Y�g1"��'v�I��'w��'��ک%�ViX��W#��NH<`�P��'E"�'���'�BT���P*���ĨU9Q��ڲ޼9�p��@�2�Mk*O$��<a��?���x�O�H8�6J	}���g�׎��ayݴ�?��?A�����/Ky���ORZci�1��*�=t~đ* �<nm�ܴ�?)/O��D�O������	v?��n�!`��	�GF,U|�C���������̔'���z7��~����?���U������8��S�Ν�G��d�vX������8�	C`@�g~2ݟ��{�ʡ;P�(<DL�i��Ib&��ٴ�?)��?���<�i�q�g�)�(�H���O�$�p�fr�n���Ox5�;O�L��y���K�o9���Sp�m�j�4|ӛfό�`Ԛ7-�Ox�$�O���s}B[���A$׽��e��,A�b�.9���2�M��.Q�<����>�S�����Q�#;��"TA�)�0B���M����?���{`P��[�Ԗ'�r�O$8���ВWǴӧ�]�FGj�r�i��Z�\��+i���?9��?�����|�ĆФM����C�Q�
,�F�'�^u�4�:�	���%��(Xz�����V�)Tk��5`<�iD�̓����O��D$�I�$).�ՙu蘪���6�7#eȰ[�b�]쓂?H>���?��N�U��u�H��WX��B� ;d�\5����O���?�	ƫ,�@��'<���;�cK��L��y�0��O��O����O��b=O��S5�i�ql������H}R�'"�'��	 x�-�I|ZGd�P�<�P�%R�wt0zAi���'��'�'P���')�Y
�{�h��I��h���C��oǟ��ITy"�������D��*̣�'��5R�H7oրx..}��Ty��X�I�v*�k��iJ5�M>��m�MшR(��t!�𦱕',�0K��Ӕ�O���OR���<\��J�	ՄAȆF2閝n�ǟ���}�`�Is��pܧ�`0ŝ"o�l�C�(B�{�8n��&e��H�4�?���?Q�'o��OݘC��ns2��ü1�"��f��Q�Ս�`$������"dy� �_�q#1.��4�x�!%�i*��' �JP�4\�OJ��O��I��
�Zb���������f7-;��A�'��&>M�Iϟ���BSpI�QE�+R �=��-�k���ܴ�?�t��[Q�O���4�����7��2�Aq�4��Ѱ�W��c@�ʟh�'�r�'n�Q��s��0�h�R���f6�Z�][�K<��?�N>���?��AU�@�`�H�D�i�
�*��p�p̓����OR�$�O�˓J�H ;�(+���k{$��ҒN�:��Q�x��'��'���'Y��9��'��� �Ui�H�##͊<����!آ���T���ǟ���gyb�Og��ҷt,R�$�42倔-��r���ʦ��I\��˟����<�0�W�D��o�F\�Cc��GP��j@� ��&�'Q�X��11cߍ�ħ�?���C���\�A����!�3d�a����O.��?a��P�I Z�A�R��)�@��?ɀ�F�?A����$��$�?��T!S7�"|`Ή�U"z�� �d�(���<�&�y��ħYf4��򩘿q�:���#�A24lZ�m=<��ߴ�?���?���d��'I�m��Lj�Y�7���E�9���$�Oh�y`�T`ԩ�W��j[�`R��T�������4�	�|I�x�N<y���?q�'�����]2;gP��o�r�&���?)��?i� 7-,,���'���Z=����'=�{r�#�d�O���4����@�@�D�Gp��@�T˼�RT�$�6�?�˟P��ş��'�~J�dG�
�fP�A���z�)χ(4�pO.��O@�O,�$�O�l�'��.�x�B���9 H>e8@!XM/1O��d�O����O>��-1����.&��@�5Sg��ya�C�|L@LlZYyR�'�'4B[�|c7Kb�%!e��q:9��}]%�2l{}��'��'"�.K���I|e���x�4`rC+��q4,W��9��'}"�����*�ѓ��M&:LR�L��Y�����i>�'"�'�����'��P�@������I`��b!�\e�r����M<�������4���]�\����o<ɢ"�\M�>7��<�V�Rv��~�����`��xy��5vJ�$�VLM.pJ��։wӘ�d�Oh��q�'m�����%V�? Ry���-��n�$P�l��4�?����?���q�'��aG;m/��Z�@ߒ\(�5z1���$r87�Zp�"|���5�D�Ĩ�)=0$��*�":*�S�i���'��*��Y�lc�0��b?�A�U�8����]�e�ܽ�Əf�]�d��<y��?���WA�i���ˏ$N�!2�)ߧ�,�#�i����D>8c� �IK�i��9Bo\	Q��j��L�𬂄Ȣ>Q�]̓�?����$�Oh����G*m��C��P!S&��I4�҃)�Xʓ�?���?�I>����~BĜ�d����L?�m0s��<�M�eKD~b�'���'��ɒ�i؞O�&�@��mjT���݉(�:m�Ob�D�On�O`�d9�� aH�h��^�e"8|�wۏL�H��?���?�,O��ѤL�G��$���ȓ���]�w�;j�z��ݴ�?�J>9��?i�!�|�kf��雝t�D9J��T�Z�oZ�(��hy�!M�3<V��������BGl�2�����I��Ir-v�	�����'�"<Q�O��,��.,���1�*P�5��	 �y��\C�F�F�����'(.xA�OdiY�cA�t��3�e,jz�"O,�j� M�6����rI\���*0�⣩O=g����W%�0@�b�bI-$��$���faJ�c���$,9��:C���vU�͋S���(y�PQ��G�	0���ҹ2�R)hR�	?�V����ˇZZm���Ϻ��FJ��V �Q�B�*���h��4^�Uzt��,45��u4������G��?1��?��4����O���0�`ͬ�@i��P��-[�L�l�`���Q�"���hc��넝9@�9����&��2{�ȳΖ�xȣȍ�j;�hc���������XD��$�d��0	Z��@eR���>;�`�	�a�^���O��=I.O�hV*Ϛf����a�&m0�Qp�"OV���@��h��z��T&\�� �ZV���ɿ<AF�@�4'��d;
��`T�M2xX���'[8C��'F��'1�U���'�b�'YX ��<NB��9�f�)��� >X�D;w#�+�p>!�+��D�N����y2��R� ��X�!���Xń�I������O^ ��ɝ+p�� e�Y� 2�a�+�$�O>��)�$:��Ͷ!rpt�A!��6�yթ$_�!�N`��Ĉ!k
�)�H�VI� U��d���IXyb��KR�ꓽ?�)�Q8�:1od��/��X���*a�G_a��D�O����:%��x�d�#!'�)���G��';��$���H�l_��Q��@4Y�&HGyҊ���t����L^>&e ���-L(��x�I7�z=:�k��(Ou�'2��[v�9؀j��]\�#л�Q��'��
�5Q�m��ѭ�P���0>ɠ�x2E���v΀�4'2)�C���_�*��}��qCsZ���	_��er�'3B���Q̔a��JD�6�@r��n4�4�V��Xǈ�H��R}*�Pc>�ħc���0�3�����B��( @<C������RQ�������On)j�ᄝmf^=p��.x����V#w ���O��S�^��

D>�ەN�T�ν3��
6 B�I�R�v9X�c�[e���3�z&�"<���)�d�R��uk��ĳ�.�3լ��<�p<@z6�M��?i���?1��i��O�ʿb>-J�+��;d�TI�+>$����h��}"��)�Ѫ7��<O�����#�~Bl[���>� �4��m�-L��3$Ɲ�[�����O`q���'��{@T�4CI٥IH0/��}�����y���"R 9Y�� (�f�h\�4�#=E�TeC)2�
7-��J�@�ʗ�<��1$�
.'�$�O���O�*ub�O���}>�b��O�d�H��St!Y5L�j�r�+�|r�ǖ���20"bc�,/��]+�O^(��|-X?�?i�t۶��RB�9Ay2�E

53F2\��X�<���%$ܠ�A�@.� �ȓP]�4 �u���!�!R54㤼̓_ұO��{c��Ԧ��	���O:���	K -�!�' Fd}�a�'�J
�r�'b�fҽK���T>�3�Ƅg���S%h'\p����;ʓ{&`�D��gR�c���!D���а(�T�C��8d{b�>#��XQ�K��<�5���V~C��O_֜AG�A7��݈�C��df���k�	/o����$\&Ez��@��к73X���tmZش�?����)�AOd�$�O���3U�,l���3<f ��K�>-*&N�O>c��g�'1���w��V���q�E�*2��c�K��"~��m�rE"�C��\��1��g'j%�i��,W�T�<E���x��f-לz��c��' d��G Q @�0����/�N"5Fx"?�S����5{�X4ct�Ł57�lJ�f�A�"�'�X�:Ӭ��dh"�'���'5���؟��2Tp�a؂k� bT�·,{��	�,����d[�;8`1��I�QrU�q �2kn�d�*�}RG+w� X�c`���(�wEB�~r@�?iߓ[���D�ڥ �g��E�4��ȓ1׀�q�(B�R"�d��3�����)§���	c�i\��jW�>�H�x�,��O���'�2�'�rk�xVR�'���C�%�r�'��Y����6:�A�"� #
�	�w��'��q"`2m���&i>zxv��	�J����I�X�qD̏xzTҀ��=,��c%D�`��mاl69i&a�?NY�-�!(%D���uχX���3���Aт��m����}��©$�6��O*��|
7�Q�P��7��+��xVa�iraA��?���oR�����Ԙ��)�.UF�s��Q�H@I��	Q�L("�4��A�B�����*�c�7|vDy����?����'G�vxr�lҪC�X���Ӳn�!��5J܈����2fiJ	I�a|��/�D�;���%J@;Z���3�,20�$�*m� ��'s�R>7���?���?i�)
HL~�ڱ��Pr�L1����|��7"�*����a¬7Ҧ�)�tb>��L/R�b�+��<��m)5�J=N?̴[&i�:1�́ɒk׍d�6P����O��x̒F���`��;�l�c(��~�'��)�I"��-J��d��h��J���cp�!�G%l�*���f��*s-^"�8���?�#�b=0T
*�J]�r���1��J쟔��2���qG`ݟ��	���!�u��'�"o�"��R�N��#� Բ%N4�~�*����>aE�@s�j���o��D5�l��H?��Dx���W��h�0,�7NȊk1�8!sF��\ۄ��OZ���Q+&��%�&H$-�5�vo�l�!��C���pw��S,n��ŝ�z�©Fz��i�>�8PoZt�����E�D�嬌'oj�0�I럼�I����2i�������|�*����	�s餘�F��e���E��<~����d�"���[�����f�
�;��PV���b��'�~��MԦ7�TCw�,<�*)�
�'�fU�B,ܸX)��i�U�P	�'�~aBQ
@<a2l�#���N�n�x�'Z�c��16o�M����?-����%#;g�	RFo<E)r �3'�!2z���O�$E�
��'�|j�펆F��5� ��Y� -��L\�'PH@��I�2mY��2�Ë�Y���ʔ*SQ��Z1%�Or���O�ĵ|z��L�KԚG�%k DY�����K�S��y2�m����ߥS��1&���0>aq�x�Mv��R׬M�=o�����y⡈�j��7��O��ı|*q��?����?yB�Õ����U�f�|1��E�/����������ɇ[-�瘚P'����H��f}pC��{����2��{2d��5���.�X1̟<S�x�g�'n1O?�� �u���#Dk������jAq�"O&$9@뀈��0��f���@�"�HO�:g	`�Zq�Afg�qQG�V<v�������v���p�nQ����p�	ޟxY[w�wf��$N!g�����VG�PQ�'7ԉR�qL���j��l��b&c ���t��m����2�p-�K^�
�<xɧ�Q�i���Z��+|O�Y��`��Dy8M��J�_�n��7"O.=ʶ͊�J�6}�t�Ǳ6���{u\����T�椒æE��)�:���0�ғC��Z�ğ���ş|�	�g�m������'`�ʁ��Ɵ�ؕ��-(��(E*Tx�kf�!�On�)�X�	7��	kA�ĩcj*@ =j��2�On���'N�� sV�۔C���5+�Y��y�g$D�P��2��-yRT��`D/�y .Y�.�a�˄�lDfP��&��yR-��a �Hߴ�?)���)^���`R�?Ҁ���k�+��y�%�O2��Ov��!��O�c�ʧjA&x򤭏�O����$�S�|&��GyFT���|�Dh�
Gđ:�'
n�����I NH��=ڧ`hݺ@���=�`��1�̌�ȓ4 �6����9r��N�����I�ē��z����{�|<aׂ��fE0��8����i���'&��/#Ȟ��	���I�TF �cB�9n���iA蜭S�e�U��O� �<�O��Oj�؀㏘l�8�AQ啦;}��!1��=T8(��K>�)��X�GI*��y3!��─�`�%y�\���IȟxF������Ǆ�)��Ըp�\�	J~!ϓ�?9
�\��Sd!�:�ֈ��O�LV�Gxb&5ғ��G � ��(��^��d�D,�2N����O(��o@�5���d�O����O�`���?q�W;�șFd�(��M��B1u��'�
-�)���9MF{��+	�@12J߂U(L�j��R�u�D\.�,�Ɇ�R�5��hO`�� �fm�mcl\"�ֽ�$�O<8k��'�R�|��'�R^���%�M������9,�IF�?D��ـ*W�KJn��]N�||b,@'�HO��qy��#c46���*�� @��R:���aX���d�O��$�Ov� ��O��$v>�r#��O��d�+�F��e@�+�$Dz� KK��|b����?� \
��ڠ����R�:��|R���?��&���Jf-\C�^d�uGрkS&ԇ� ���0��]�*�����I��Ն��ȓ$��=vFA�r�̀����=fK4����O�	���G榹�	��d�O���g˿:�V�κJ�${�gN>,{��'A���q��T>��F
4݂"&~�BAPj1�#��yD���ǝI�j���k�	"������<�(OF�#��'��>�Z���XSFBTq(��I3D��0��)��P9���J�6,3�6�O6�%��K!�;a�:�2�薟c�<Tk%s���V%O��M����?�/�XȨsk�O����O��#3����9�
E�j�3��X.����*�|Fx�D²���3���<Y���W$��RN����)�矔�u.�?/V�0ץNQ�e;1mF9\�"���ϟ`�	���G���$�0�
��Y� �4��#k�Γ�?��19s�)'V�ȠFS��	Dx2�&�S�d�޵0����MO:(�	8R��9r���ʦ\ 1VN�N���M]��!�SV`
�\�a��)_�U!�D[6e�T���#�t�`��rN!�D��a	DЪ��ӌs@��ز�0E!�,��lɤN�?6h����k!��$���k Ҝ 0�$�'��w[!��,
=<����%�IF&J�u!�D�3@�I��H"���F!�D�j��Y׌Y{Ҙ*u�,4!�� 9h�K�K\�&	��@H G�!�d�':N��Βj0akt�٠+�!��;��DR!�=�(=ɢ
OBP!�D��~t!�f8�$�R�H���!�$X#+L�u��+sƘ��甦V�!�$�;[�F��Wm�3S��t���	vy!�� N�z�#3�]��j�=SzB�E"O,���'�b���U ��z��%��"O��V�A�z l�S�\S�yz"O̘PQ��?����ƿ�f��"O�8�1���;FD@7��;� ���"O��H�#8��j�'D*^��"O��h'�#'2u�R�ƩP�Ju�"O�}��b[�>�V�0R�p抭"P"O��#G��"���ǅ_�A�����"O�����X�09���L���$"O�}`���$�q
�G�F���"O���A�1:���MK+��su"Oд�c�ڴ)�:����ޕzQ#��>�������O꼄�r�-kڒ�����!����'β0���Ȳ%(�UcB����yB��Ns�̈́�	9|�6XEΰ���řk�nB�	<6��#�!�+�Ў#�T�S�� ��}b�@��>A'��1�pY�C�N'�����)�I�В���<R����5	����H�<�s���P5L�iv'�Zo!�$�hJb��@8X��ت+;�I�0������fe�E(�����(�&^���C��:8X���p<�x �h�8m����P)
�Cx�CC˙%T6��K�q;p��]�g̓s�qdc�>�ȥ�#��5�hɅ��3��p�҅ۦI0T�X6�1���:7�[jݸL؀Kԯ!��<��I3<Z�*�f(a�tͨTȖ�HT����@w#@)"cW�>4e��5Ot����B-=4:�r��F�f�l�v"O�P
Ee^)���d�%����᝟�1�����l�|YA�!W�O�Tp�i����%�14K2���'#a�0Ώ����蓎vӼ� �� Hk���'
>�j3�-�Ϙ'�V�JRĀ+x�J�H�ܘ/��y�'?V�H��'J�XÅ#Md��{��-��|�c�������
Ğg*����Åw�nm��	=��=Q�G��>���cr�,��o���b��b����G3D��zǋ�b�<·�X,
��a��#�<�� �&"1(E��S�P$��F����n��RqJŲU��
 K��yRD���Iz�c�_����S�Y�j��`������M3�#��*0�W���}C	%h2L�Um� ���	�*��?A!,�2
Pv��ď�=�H��I��(*��(�cG�|牄?���	�k��H��Q;6.��'B�=`�"?�rN¬ڀ�u�x��W�(gzI t�I�V�Qz�O6U4�zG"ObH�$D$g�n�)� NSDk[�8p�\�D���&�'�$m�*b�>J��܊RI�l���Mn�@Sf�>D�hA�LM
���9F�̓!됙1�B���Ģ�&���?��9S����{L>bA�'6��zCD�9��� MDn���f Q #�A��ES>jn�y�m����Q6
�|�4�Q�7\���U�'�P�7o��}ƐA[G�K�`k���
Ó9�d�1����Yw�5( �A�G�Lb|��+8侈�Yt��B�	�w?�5���O�')6I3R�$�ʓ���� %�-��QF��/;�~q�S�'{�F����	�L���ǧ;���V�D Ub\��p�Bw��  Up�b�FY$�Ɣ��S� ��'�	�4G��'ORq�O �R�4��	��q	�b�����W�S=N JF
Z��IӁ(�)�z9���4ᤠ����]r���'�2I�mIQ�z��1,}f��J��Dڐ.ˢ���#E�yh`�1'�G�)�d�.p�)�Ǚ�;�X���Y�����'t��* ���s���s��n[���O�������t٦ŀzj`�X���vȋfݜLB��At-�|��xB�"O0)B��8fw]�u�)?:r��4��b��ar��e}��ǆ�ħ�,�𧛟��d�J/i1��`"�Y<���;�O���`��)\̎����ÍD \��$�F,,a������
i�<�J ȕz|���Ą�M��.z��(���y��\x��R6fS\e �$LO.�PF!�i.2j�W]N�b�AƷ���R�M'=� �k�,@
��'�ԕ[ 	��'�	˵i0i33���B�K"��c�1OB�I*��#�]�	�s�x�]��>E�Tk��=���Q盜1첸�׌P�&�^�����CN��"<pK�JMV��Aj]�KF,��@7$P��l8[$քx�l4�?6#Ҝ[|�7Ms�� �u�`фC�-��	�1�l���X�T�7�_e�ؚ�!ڱ!l<�x�� �i$l���*�D�X���1��I{��D92���Z���3��/Su�1S�<����P &�� ��GϪkZ4 ��	3� `�o�m���R�iM��X1��KP�;�<H �eTD{��9�t�'Ó�aB:�S@�X�G X0���I
T\����U�@QPV)޷�h�(���!4BQ��b� -�� �����%7a�T{�Dӑ^��m��<6��jP�7�����_jn�aw(<,O��rQ���v�Xm�N)���h}k̎�z �qB�}&@`���/~�F��#���Q C�ٟ�*W���j�hB�Q<XG�MVMĚ?� �>��;��_;n֨�7��t_��h˘cY|4/M+��B��Ll�
��'~ٯ;Uy�3��#�y�B��F�
b"��@��[��0?I�N�����Ul6x��2�JM��رiZ|�fa`)O�4 Aoߖ	�p���]%^��͡�\#��I3Q���Q1|�M����)X��#>i�+Z�>!�4�&�_�i1v�9����"5#Ul?l�X�%�E1`@�2���Ū�5!��`�4�J4C�d��ቂfa��x��̎Rɮ��v��,e�I�w���*��
�-W���Vn��&�6mS�}e\ ��"}F	�2��HHF��J!��ᔱ(�'?zEV!�	I�pm�q��/1z�Y�G4 ���'�*����@5�b�r�>�	��ʿ*nx���
s�XI���',$��'@����%r��ˎ7Òq�G�=�𤌁�ԸI�B��]�$� ʟ�m��I�J7��{�e!zv`E:!k�X:�">)R�V�5/�m @���dL�CW�<��Ѽ,}���Ď�	E���@�:����o�l(�R�� �1�����پd�� E���)�]jG�PCy�����v���6�3��ɞ$C�4:(�n^0\*���$̴��r�M�c �����wF\��ã
�Cj
����'A��	zc�U8���PWh�7F8`�w��a�i١p<`4wn\�(\c�`�"P�¶4c��
_���X5���i��	��'�$j�	���(}k&G�#Ul�J<TC�I��KaD��f�1�mWd�'�� ��F���ʘ8��}a�O�9h���5X	��h�"Сe�<:�.��6�Z\��h_�v�X�#<O��K��U�Zh0�*5iM=�*(C�FH�4HZd��È������$�ax����.I�K��n���AG�̠�y��ɵX�Υ���u
Ra3M]6rϞ]���:
��(J�%�5Y��]�bB���'iO `?�H�ħ��e������2��pV��� �r��SEC�x��z7���)�fq�,O☩c��4>n�����Ä��U���	Q��xg�� ;��sd�M*y�#=�W��h�^���l�=&�8��.�j}�d)N���A�=1Ó��	>�֑�p%P�[Ԁ���	�0�fEc�爯ls�����-W��"<���9Z�J̈�`�1Y�EI%�]�����!��2D�S�]|10uF�(7(�B�ɉF�bbHQ
gn����2z�|��UhTf��u�(+h� �s��i��?y�D�6J���#�̥ ��Ť�r�<)�G�"�*F����)K���q�<Y7�K�x-���S��!��cE��w�<�6�u�K��(Vx� B���B�I5�e��M?+�8q�T��~7�B�_4��ᨍ�
]�̳! �� �.C�	�#�z�H��["վ|�H�z�lB��V!P�D�د<j�����%i�B�I�Y�r<3Q	�76�p�ULE�	�C䉙&t�j'�\�/rP�2Mΰb�C�ɎV�еb�cMpm�΍5\1�C䉚cF��a�WN�рG�&5�`C��<.v-rR�Y@G�� ����@d⣢L5~إ 7�#A R|��+� ⦪�t@��S�"oP��ȓ&wp���L�%iиxG䞵S����do�	��y�S�OҢ���@O�	ꈉ�ѬK_�Ձ�' �d?��m#aDɟn�$0�N�����;�^i��"�z�1�ٕt^����S@�����1:�x�u�A,c��db�x�R �FcY�.O
B�	�`�HԘ��2"���'��[@�>Iv�E���É�$�[s�v�p�Ԯl���Æh��y�( ZO��s@_<]�l�$��~�lޞ���Zu�|�����I��"3�@m5j_�a!�Ĝ�6��@�l� �t�!)�36�&	�DCS���<���=E���E�$EX�9R�]��@�$�p�l%�!��u$?�S�d��K�� %H?R��=@th�5U�.�����t� z�Ǌ��5��Xt�&{s|�����t�hsA�A��S��{�'Tn��b0�G&P3��yG+�T�F���P퀷�@X���;���C�&e鶑��%6B��"�O&	7��'���h��aZ��G5��U��E�I1^\xUZ�4����6�8��T�{�ƙG��@�B���+��-X������I�YS��W�'��%hwL[�D�&�)mE�y�d)so]�rϤ����F��NA���gy���,��"�H�� c6B�>�氋��'@��Bb�8N����BkV�X�A/�"LG���ēJI�0SE����&�Y�1���EBL�3\��~�D��(��	;1���q\�Y�bQ�<I� ��Gʜ���N�9d~9sG�
fy҂9=���=E�$	�!2��Z��jj�h C�O��yr �-�dP��ᑜh����̦ޘ'��Q2�-,O"���c��A�m��P�}���ku"O�}�$W�6et|��b�8W���B"OhXP�NK��(s� �6}�Lc"O���D��&�|�� ҟlw���E"OjD;c���n�$��$Gt<��"O���G�4tY�i��5N���%"O��!�	4G�PW�@�P��Ѷ"On�:��[^��Xxހ�Vœ�*O�͠�D�0/9d�fË�w����'84iz҄M&}��`k�Πq�'�=�f#�<�^t��b.��
�'Ϝ��E.��_9X��n�c�8$�	�'uM,9EN 2A�L�D8�rf��p�<�#/%E'���r�O(+�&T�p��l�<�@NB�ke� %)�R5�ta�t�<��J�Z�x�ǧK�}4-
Ҧ�n�<y7-�)!\�P�g��"H�ţ�O�<��R*)��,36��~~e���P�<�v
ӓ{p�������� �E�<!��@:�(��3$e"�Y�'�L�<	W���`�-(�t Yg�R�<QT�T�K�" ��ʨb��b�Qu�<15
����}	�EB�}�ll��+�l�<���_�eO���'IB,b����&�h�<	Ɔ�2Q
��r6 �)(_��:���<�[hq��̍�#����'��\�T ����$aˉ=6��{P!���ȓrҤb5H�\@$܁�̉�Z�¬��yR|�s��߶G��й��V,�����g��� RC�f�����_>C�*]�ȓw��J�i5wb2���O�:8<�ȓJ���S	ك!�2�� ���R����"�dM{��Ղ]�r 1��oZ ȅȓ*�V��T���b���g�O�Fs0(�ȓ	�*��F�3
��JF��->g�i�ȓB 8r�AD�sɦ�A�c\+k�`��M#�qC���D�B5��(dن�w9"]�����l*����1l,E�ȓJ=�=oאM�HMU�$���1D�X����
+��(��Z0:*^��n"D�<w���s?�Mk͕J�*����>D�$z6�:U�r����<X��S�<D� ��H�����+ ��M	�;D��bb��Zn8�a5����s�7D�T�Wf�/\F�a���M3Cڪ�s��?D�h��)�rR24{ƌT5����+<D� ��+!_���4"��ss����E:D�8(�I�*#x<�#薱�X� ��2D���6d�3t��l8����($;6%D��1��6%W|E�5đ���u�#D���B��9P4�xh!��Tv
 D�� b`V ��R�h�C����3T$���"O9����P"ԧ~�T|��"O�zp���`R�=�T
�"O��\�>�2T�@�H&Ar�Pv"O��[�e�Z,��ɼ8Tʼɓ"O��iQ�GOV`s6��ZR�I��"O@�Z�F*?\Yp��)^Q����"OLk3� �\�b"E*���"O����*�i^���\#�Du��"ORA�oŅ,�С�a˽��M)�"O:uJ�)M�p��P�0M{+��y��*tfA���.7��c�D��y����C����+p��	�a��3�y¢Z�X9�pr��R�g�v%��Mߎ�yR+ϒ!z�X�oY�c[0jA�F�y�D�S��b�/�;l�ȃ�H��y��"_��
����hd�x�g	�>�y҇IT�.Qy�EExTy�J��yRiB���� q�Z5�L�hP���y2i'o�tٙ0�ٵ�(�gͪ�y��S��c&N�r��%8�#ͤ�y�D ���GꉮbBTS�+��y�qۮl[�ȿL B�c�E���y�}-�h �GA>Fw��Ї
��yR,2I��qO�C���� �y�Mpꀻ����A��(0���hO�����J�y Ȑ�i��$s�
�� d!�d�>�t(�l�]�d��)@�j�!�h�!c���S뺼A㎸_�a|��|�"X,&GNd��嗐iƠ�� ��)�y�)2p��U#s�4O�Q�!⅀�y"�̜r�t����H%�����M��y"h64����B�N<�X����{�<I@C�!dH� Bb��>��ȩa�<qv�-f�Zh��% 	n�� o[[�<�VhIv�B�2�S�N	�4��S�<W�ڀ
$fI�T#�"���&j�u�<�`�է:8�V�\�.)��Q}�<i�ᘱ?c (��C�%I���!l�a�<�ϛ>{.6��E�O$"�x<A/�]�<9M&�4�k��:[�\��ӋX�<�b�U!ͮ����ƸQ�<�q�MW�<�g�>P��ϼ�V%����]�<�w�1;D�ԣC@�=O7�A�ǧW�<�'
	]���yp#��f���-�U�<Q�e����=)l"�V�KO�<���EZh�2K� N@��Y�)�K�<�f�E��}Y���pR�i�J�C�<ɷ&�4'�.d9���>q7�|����B�<� �Pp�$G�_�^ma)T��Q�T�d!�Y}���/8D���`'�3x������tD�B)�hO�S�2�t	 ���>| ����3dlB�	�LЬ&��Jl�@�@B�ɖ{
�=�N�n]�+�;A�zB�	� �T��t@�*�	���	3B��#$�ɐ���H��B�׃��B�%;��d$\n�$���E�Z\�C䉎;"�0S�mЯL$���-B�b	*�;S&*"�<D��C�C䉴�E�����Xyp��-��B�	>}��b���;)�-�:�B��"$@�[��L)�Xa���3��C�d�xr\b��<�3`���C�)� .̛�đ3\�LHs��%<�&U�"O.|1�$�#���)pC�m�q"S"O&%��E�w%x8SFb �8�Zu"Ox��L�,C8U7!E Yҩ��"O �iFk��&	4�rр�,<�Q��"O�m
0��?M�zi�� 
)<X�l!�"O�T
#X%P�(-��A�
sF���'��O�usf��% �DN������'�'�=P��&,( Jwn�-S}�����2�H�nh���7x�&!0�P�O#�4�ȓ{�^�G�AjX���'�fф�'[��BS���ZLz���E�"?"��k�p�0��Ãk咰��������Z��"'�
P��bҭTg��ȓf4�B�)i��	R��+�̭�ȓQVnHS$'˩oz��%%&?�a�ȓ)UZ��7-�P�r��Ǒ9z�昄ȓy�x�G7;��I��Y��J݄ȓi��ӷÝ�W	hM�l2 �~��ȓtR>�q��9���	�$9�2�ȓH� =J��ܚR�Jm�!H',��ԄƓq~t�8���&.���1e�?��1R
�'ZM(F.��j�(
�]OȄ3	�'Iu�j��8|���L�4Z� L��'p
 �#I�A��칆���e�x� �'2�hq# S�)b�IAk�`$�r�'�~e��Z k�$IH`�2B��ab�'_z!���,[�d$�`F6	�B�j�'e^Ș�L��a�ɛ���)qQ
���'�N�����冈iaG�:g&�xp�'�����)X� n�e��'�<4 '۟sg~x�e�R!h#�'�B�Sjӥ��%!��D<�)�y6��Q@�Q� 2��@�y��\�H'tpڅ�Ez��x3�
�y�B^�8�
т�s���Q���y��S>,�F���bn(�쀠��%�yB���eS2͊򉈢_�F��B'0�yB��@$�$$J�T�4 �c��yB��8��|(��>BzHRP'�y2m&E� a�a��
8�mD(�y�#ư=�,�ҕ�� Қ,
�@�yB��d�H��A(�u^��Ud�>�y����Ej��Ć��a������	��y��N�BIabY�S8u����y2(�z��a8"E%8�V�Ѵ�����>�K��8��D^7V9Y�Ę�z%�q�AJ2D�D1��# �1�	�ɖ���/T�HS�'�(^R=��
�7�$pYs"OLH�@l�4k	z��`�_�*�ZēB"O
�UNN����B��)�,���y2DW�Jv����i� 1�6A���B�yH?%�h�j�m�7�J@�Ҋ�5�y"��
��T��/���r%l]%�y�M�$�p��1C
;����#��U�<qb�O<r��E��x"��K�G~�<i�cF� ϼl��ڗeԔ��	�{�<�E����S,	s.�����m�<�$Z�t *�xƉTrȈ@8YA�<YT�-i��i�>Wn�P�Bg�<�U�� ����gΊl���X�<	eՔNT�;���yY|	�&�SR�<١�At@�@"R*�v$�U$Ms�<� ��RI�5#q({�6ء$�v�<� ���RjS��L4;��C'a�%��"O���&�|j�5���[���E"O x��kNnUf���c׭>>ޡ�P�mӐ%�<��t����|�!qR�ͫ3f�Eړp`!���Fm �Xd��C�f�3�)DF���/�����X<L��)㇪ :,�l3%�**C�z�	K�#�杈S\������HS0�)4�Ók�$X�!�&?A���.�p�ɷ��{vHa�^?U�xB��0T'Dd�4oQ3~�.��0���.˘B��M�z�#b�Ѥz��5�$K?\�<B�	�Tv��r⊖{���D57��C�	}6Ri9��d�LȓTL�/T�XB��mAR��d��
i�K�%@RB�!��a�J�r��]I��ʼxjC�IA B�[�'ڣ? ��@caǗDtB�I�6��Q�rHW�a�P]"��;N5jB�I}g���''X<�6!�V�B�e=*B�I=	��h��m�tF> �r߁[��B�!b�*	Rg��+6zIa_�\e�B�	�+t&�kW%�cl�r���5O�nB�I6�z�ࠅ��(T����%a="C��5� ��i��F�r�+)BB�I-QB�t�s而
s��z��9�B���n�!�R��U2�ߜ8��B�IrѬ�0v� ?��s�*�
(��B�J�L�q��á��Hp�Z��B��vi�E:k�$D+7h^�b/�B䉓"��h�4+��4'��B�J�B�I�3��	��ņE����*U!�B�9h���8�H|�T1@�Ŝ,�fB�I$C�v�cgC�K�ꡢ����<|B�ɾ?�8�����p�De���&B�	(O�Ԭ� �TGP,@��ݎg�C�ɝM�Y�F^�k�X ����"}��C䉱JX��F�8-��J�.��i�C�	7g3������2򽒣""{�B䉄d��i��IE�ڝJ�"A�*{�C��8{~��+�傍C��}8dO�<3LC�	B��QX���a���[20C��F�R���+_���T�G�I5�B䉩Z�Z)��H��vN���t�	�3jB�	�X��(��J��M#�t{�I22TB�	4l\�CHvӺDb�+�t�ȓ}�,ѡ��Be�95duxS�OU�<1P��4�n@jFM�,7���FPL�<Y�M�C'��w�^.`����˞�<�f��	HjS�R��xj �~�<� V3|1v<�D�T �$)�-Vt�<9-�I�v�1�O�g��ms1�s�<!v��?l|d��k�9j�H����S�<���9>Ƕ����5� �a�N�P�<V�:Q�U.;���uN+�~B�ɲp�`51�·���	r�؊ xB䉘]>z�v�^	�~a	��<ZB�	�:���t�-`���偏:	�B�	" �.��T�X ��H�o��D�B�ɗG�@�Yp P�OO����� iB��w�`��6J�!-(��S��(��B�	=C���#a�0��0�i�2E�B�	�h����$�7[nH�"J����C䉆LP��KІ�>*�rUQ�$1��ȓ�.9)T�	�#�`<�&��i���ȓ!<r5b�Z?#+�8HE�?v�t���bQ�zbCI�>@�&�� Z(�L��S�? ~�kp��,q�]�w��6zl�"O�a�l��!m���f �uZ�IQ"OVM��oՕr[�%���3S�=q�"ǑV�����t"�z��%"O�48��!LaQ�!$��d�F"Oh�B��\�:@��į�QE��!"O�F�$;"J�+a�"O>�1EG5d)5�]%ުQS�"O�9:UAǱ\M�$@��S���"O�\�����n�a�M#����"O��G���`p��] 10E�b"Ox}�7�+<�p(�l� bR�KF"O|��d�E"Ⰲ#�-V0Є��"OX,��26���V�'����"O`�:���Ge��1�F1y�3�!��^8��Z�铯:���j4��0n!���|���b�Z�"�VA;�/[�/h!�D�M��� e�J�o��)�T�	n!�A$е�Â�),�p!"��[� �!���B�|�-	��.m��LV�v�!��"޶�U\�5����d�B K�!�D'Z��fEZ�њ`	ꁀT,!��	%�  �"B>hʀ�5��!�!���
L���=;'J�e'� 8U!�,��i��	�g#�|b�F�,R%!�$Ìj�4��Azv@�q`�K>X!�$���,�R�ƓSdf`)t�V�l`!�$���Ĭ3�l�1CG�q���5/\!�ď�4�yZ��a;��KrB�N�!�D֧3��0��Lj2��(��
3^{!򤟲y�P+�Mr+t!	���MC!�$�H
 �PnL�Š���)�!��Dg���h���#k�h�V+ڊ	S!��#<����7|�.��&��!��L?q����R(��q�����)�!�$@V��)v�V�zu`p-��mk!�d<Lͨ�AҎ�m�>@��)�f!�d�@r��a��5yA�ɱJۡ!S!�� nЄ;#�Y�z%��Q./!�d_��v��1,	�����$f�s(!���8r��x�����D�"!�ҷ-a�Ib1j]�lZ�ɰ,>^!�d�F�4�H�cA�D�^��5K[�z�!���0t�3���=�m�J�
V�!��d��;рQSPd�z�
'3"!�dԨnyE��*
�NA�zd,�67!�dр2�� F��09����z?!� Fp
0&�ԼAȽ�C�ʁJ?!��,���K��U�A���C��4HE!�
}f�]b���
������4:!�DÈlj���J{a���VwZQ"OL�C��,|��0Kr,�b�.���"O��FhJ�]�
P�L�R"O�Y"$f�*_�I�,ĂDx (˦"O���W���D�Z���xo�0��"O�X��fL�:̹QcILD����"O��j��%�J��󈂚��]A7"O���t�ݨyvl(@6����� ��"O P�؜d�.���]��p؀"OdE{DDBŤHSe!�/�Ҕz�"Op��H�n��H���	�^��C"O�݃`lM�@�Б�C3En�A��"O�ҖAJ0-|WH�L_�EI""OJp�Q΃���	��Z!bV�M�B"O� (L�3hQ�!PJ������yM���"O��A  �u� �!a�ߦ	�n��V"O6���Ҟ�N@��Gk����"O��b�
�ga����C:=��S�"O��hP���pH���{��S�"O�����3V؅�`�Ww�P��"Or��F�kP$
�'��Lն7+!��'�b1�JJ�fq80��KH)`�!�D���u�D���<2���6�P/R�!�$��!$��g�� öI۲�Ĭk�!�Ğ6y��� �ȃ�>���CB�o!��[|��a��)tH"��r�ֵJ!�Y�BOH��+�B&�h��ҩ`�!��¿<?LYʱ��V�!���D�0�!��\4
�$d����1*����D�I��!��V8���Lu.A���\�p�!�d�#iv<9G��8Z �3�ڄn�!��C�.��јVnկ��4�˕�2�!��55ǐ%.5�Љ�7I�Z��1K
�'��0��g�,�('�$f�H�	�'�Q���\�J�_T����'�zi��Ĩ���ڗ_yD���'�t�	�5	(����!6h��
�'뤥�s�=.r�|b4�Q	��qH
�'纀p��-/*|�Qug��	�<�	�'��Q*S�]�XpMs���˘��'���[#��;o�T�s�G�F[����'�.�aWb5`�ha�2I�Ѳ���' z�a(ѯ{�R���[�z ��[�'7�`2���H[BA3aE���8M��' ���7:b^��UR��'��z�bI�
���OD�=P�<��'�(�;aPW�t�'�Ă���'� t�eǎ,��s"� �z���'d(�
W�Vch68�3�ѮB�T=��':8`� �2t<��TB_6礀1�':�Ļg^�� A9'i:�����':.`rr��!�� h�OW0�65��'Ц9�a��=0�Ѫ�� �����'3fppq#�#<iXU� Sf�|ܐ
�'S�¦�8��Ԩ�O/��j�'�X4"� ^�<�s�_(�2�x�'\�5�P"�b�������8�'9ƕ�1�P-':��I��1��'�@���X6[z��7d"on!��'�b8�(�%�hf��~�D�a�'��lX��� ��$:eH�#�}��' p���cX-;t��J���$O��']��(��֔?z��0JҦ! 0h�'�v��aY�.;�Uٷh�A����'Ȏ}�$	�.f�6A�6��`di�'� %�7�Q�#�%�%�ÅV� �'�Ri9��$R0��t$�=a�0��'��A��`X-^������
p��Ms�'���.2�!�ClP�`�'�})d�6h6���-��iŶ�"�'N��S����>Ju�'O�#_`,	��'��Q`�30``��3*�va��'�ڱa��2v�Ve�DÞ.T`��'3 =�4%ҸH���Bd��' �>1��'Eb�IE�L�B�A��ʚ�G�:�S�'>� �w�"p?(��@�L5=�&	��'���a�d��gvJeP��?g�L���'?�I����XM�����u���� ʡ��/�5F�zY��N����`D"O`�1BE2K{�m�AQ���"O�C�Ǖ�$�L@��=-&���"O�A�DU2N��B��L&� 8�"O�t{$��e�t�들�03�ؼSE"ONyP�@�x8�g��!lu��"O 1�#��q�ި"�e`n&��U"O��@T<����޼Lc8�I�"OYw�Kq� ���Ȁ�m�8�S"O�=h�Ĕ�[�X�2b�V�:D�"O�����'$��B#��|4]I�"OXaqC�69�2�:BΘ�q����"OR�s�NP�8X𩙔���E@D"Oh�kԥ͗Դ�P��Ms�p��"O�y:�0|k.h{��I�^ꎜ�"O�aUgA����� '�z�.P�q"O4�i0��e��"��!]� ��6"O��C�HW�������f�"O"�	�n�o�|�a�{Ebm`�"OT4�����`S��Ե�S"Oġ�A)�����N��B���@U"OXI��'/�Z�bE���s8n��D"O,h�'!�@BCG��	bR"O��Zei�
x�� ���L�pBc"O
-��)�/(>ʼʖ�R�n�4�е"OH�8�j�<]�p"�gI�5�8�P"O&X �ܘF����ť�75Y��P�"O�8�F�f`Xa9�A;	M��Ӕ"OȰ�4��[~pJD#I�PC�"O$lp�@u�P`��\!�18'"OD��"l��Eu��@#��i�zͻ�"O�� �._�Q@�'�(:�f8��"OT�[P�/�.����U;�)��"O�͓�Ň�#��!��E$[/�	T"O��;�G�'hS ��2Α%Z�#�"O�]�  ��6�\�8��3\]�a"O0X����dgĠ��ۜM����"O܉*�'W�g��\����C�*�R@"Ot�"�D�#0��E������2�'8�M�t�֗G2L���ۧX����'��9b�� �#M,�E
�<Q�9��'�t�f�T�q���qk��H�L�
�'^�)��;�^PApb˵?)��*
�'���T�Đ5��p#G.�7���X
�'�b�;��ބL��P�eM�cGf���'���6���H9���$�M�V�� �'Dj\0�ݶ�p����EV�0�'
��UB%����C��88zbų�'��k���X�K		�`L��'0�QA�φFǖ��+��:�'���2A/U&�4xBIָwH��'�p���ľư�	Ҍ_ N�謪
�'��8�،(� h�G8N��5��'tb!� j�NZ����xb�-r�'��9�B��F}����딐&t����'���ʤO*x*��t�� .P�'{��"(Y�j#"a1�d��L��`��'�f͸6�Q���QD��q��'�H�����
	pQj�9F&V��'�)��P.td�P�F�Cج, �'��c�ٟL�\��Ȏ5����'6(�R�,���]SFn 5d+�D�'��4�L�7^���EJ�������'��t�]!
��X��8G�1J��� \:�ͦL��ACAO+V�I�"Oj�p���8�� �-M� +�"O���V�� ��0�c�1b�����"OU8 ���\@ڕ�g��W��%�"Ofћ��?�n���iO
�M��"O����óY��c7�q���2"OBL8e�ހ���:�dٛczإW"Oh�ʢD�1}*����k�eF"O8	@F>v�P���≣7Z�2�"Oĉ3B�Z��̉DP<_G�	�"O�Xj6�γ�Ba�VNk*F��"O޵[��^"G\���d�ǮTY��'R��� N�'��+7d�*!�X�@��6D���*
%B�,�[⭛�o䵉�� D�T@̑,&O*x���/:��q ��4D��/}Lb<��!�;]7��*�����!�S�n�!R�[�`F4�RD��+�!��<��h�a� ̶�����67T!��X���)�&��!�+S,>�!���3PgT�p�_�_
�x�E^��!�~�¨Q��"d�j��'e�:�!�D��Y@f䃵��
|>p#�L�n0!�ZU4Z��2$g]0E9�eG�/$!���/4���Z�̊OM�u U�$�!�DX=4R9x��<��� �Y�C�!���X��1,�8'�LZ0'Ϯ<�!���4c��!���&c!��Q��KD�!�č��������M"n�3#�� �!�Ф~� � ��4J{Ir���%S!��	q�VF�<,z��x�σJ!�^VX���?p^�-c5�X�}/!�Dj�Rx�􋟗"�x��� l !���$ �X��GR�w�\�w'�0Mg!�B"�6��b�C+3c��vF	�W�!��!!n��T�Wč)$��!��(+Y�u��+$C��Qq디�!�� 	c��@V��(�YHT�=�!��F�{���#+ڱ�� ��!��H
16JlyCDłdk� ��)�>�!��B�-R"��f���D闅v�!�X";��	r*
hk�5a�3t�!�d�qbR�ʓ�ƿS��z&���A�!�$��SI�$APM�
xl$
G ;w�!���o���+��(\�<��m#b6!��4�y	q��>�H��T��>!�^+�^A�`�_ �p��p� -!�N�.�Tw�[chy����F!��S�H�1 e��X�ܰc(ź+�I]��(�&�+Y�e��AbSI�m\|�"Ot@@sF�fH�]Ca�K�:%�c"O���#d�4I@l�����#���+p"O
���ꁹJ��DҒ�Q�3g�m�f"O�) � ̋U�X������QP�"OfL���5)�بF!	y�!1�"O
����XE��X���ߠ-��"O �[�R0��ZF	��G+��"O����+�WR��b���+q>-B�"O� �@��fҸ���FL�O_���g"O�ԪC{@̔a�d�w5(m��"O�=(�ΚH�B�Z�$=##̴�D"Ofqq7�_M ���]K���:�"O9�pi��*f4Ⱨ5l��� �"O�d`ã�!&� ���!C��e��"O|l�dO_�ril�����5|���a"O� �1��M+l=k���+8�<[2"OHx��i�8�����(q@��"O��zG�N��N���ID�T̘�"O���ҋ{�ġ(��ܦH���7"O�Uۑ�L�c2���@	¨.��(�@"O��C�L�R�d�#�B;��<�"OH]�f��+[��P��Nؖt��"O�(���B5k��LY��������"O�qAGMқ-�]2��U&s���s*Ov�{F��h�zݨ���_Җ�Y
�'�:�͜8�(<!lRU3\I1
���d7W��d��ME7Z$�A'JÄQ"!�D �G 9v M�7P��� �؆	t!�ć I��)��P����i���!�d3��D�F舖 ��%㧉P�!�!�J�����u�C�B��+pOZ$�!��&30��RtOH��d����!�DK�U0 ���/�|8�Jњ��}B��/}G����_�r�H���!�$Q�k����g̷K3"�bbI&j�!�DђBU�H��c�:����!B�!�F�.�%z�KE�~.P�ǻR�!�F��iie#�Wc��s�ʕe,!�O�Y=h)���A�3aʭhP�Ģ1m!�dU�����#@�c��hP�
�w�!��҄	�"� �	�4/��O��=���٥�D<�iy�*W�L�� �P"OJ-8�������Z�J�������"O�(�e� ��@iߤ���"O�-h�BGC��E	 n�'��9A�"O��cd���5�lZ�B>\�F"O�I�u��Iڄ�R��Q$�rG"O��Zc�P
X��(� J+{օ+�"On�§���&aH�!ц�-�(�W"O�Q*�(ȊVxx�t+�?�d4��"Od�7B���'��)o$h�"O�9e%W�=xTQ����hh�i;C"O�U�f�/+ɖ5��U�P]�-��"Ob8��-Ñ1���CcX?PR.�KF"OP�A�a�.G�u�6�
iY�1
6"Ofy�4D�93ICpƖH(4��"O�iYn_�KԪ��C��);8���"Oz�IFڎ	2��1��]�{�T�P"O��pVHZ[����^����s"O�K��صE"N�i��_�^��@�"O|���~w�p��ޮ\�ձ�"O20���H��$�p�i�3$ժ��U"O$��E邖GD޼�q����x��"O&h���ۖy��iP[�<�d�y���m��1%G�|� ��NN�y�
���5��M"$��4�����y�㚊�ȉF�T}��#J��y�M�F;\C,��H��M3ӊF!�yR��=��pAa!�;E�ike,X��y�?7?�d�#+�9Ҽ��uō�y�NϒI,p����.@l��N���y2Y7e��-9soSm�>@ ��yR%���F���C�%c�����n��y�h���vL�ԥ\_h>�k��V0�y�Q.M���I�h'O�媄�Y;�yB@�2x&�Xb�e!�*�-;�N�a�'1J�ءK�H����
�3d�A��'����ԉ�1^`�$��/�P��'���Y�-\�:�-c�B5%	Υ���� �`$��-���&�+tհD��"O)�ҏ�(5J��eĉ5ѴU�"O�yk�Ʉ4�*3p���`(A"OP +�@�^�D�AF6N���X�d2LO�	�l��@�8(qB�U�V�\i�"O���ŭ��@���!����S"O*h��Jw ���w��$6�D�"O��dD6C�������u��Lc"OT$x�g�0G���AJ�>��dR"O�D`���2%��RFiS���9f"O.����<x��@��DV���"OЈ��_�'s���%,VI"w"O�9����5T������&8��С"OV��>i��)V㝚m���q""O��!\�VH(��*��(�!"O��V��D�"�2t�\:���c"O�q;��޲m���Ca�H�%FE�D"O�єH�:���KgA���1ۑ�II�O�ܕ�TD8:��RH�{��h �'�$p�V�X�4� ��ӊڅ	�6�a�'�$DYg�J1b��#Z~~�]��'�ְ�w�_6E��� ���w��l@�'��y��%m�j�F�inN�P	�'��dqp��={Fx�ڀZ�,�`i	�'�Թ�a ��H.��ceß+�JU;	�T� ��'��iH�
�<	�b)��U1=�ɢ�'J�8��)_/��Q ��@'�����'��hţE"kx��'F�2V��r�'S��q�L�9�т�h҂˜�@�'�p������eY�
�*5�2���'��9�TI0=����	 	4���'�F�S�_P�B�Y���9	�u���r�<C��Ы4��L��j=2r���ȓ/>�8yg�ؖr��0ׯ؍G��لȓs�M��ڔV�8,�g�U��`�ȓA�����	8=U�y�W螞+\f��ȓB�8M
(Dђa�"�$4Z؅ȓ7sD��&!���������K�����	�����O/y������R�F��ȓ�����L�&����PN�1����-�r��ӡ/t�D8�a�7��q��J��}��釁Q�����L��j۴\�ȓ��y�@��R�L22�/X��d�ȓ ָ��V蝔p'��"gݩ)��݅ȓf4���3
�3Oޙ�VkB�`~�Q�ȓiJL���. 9��R��2�j��� �����M5V�*&�F9�e�ȓ
d.��t"��1��	��
��ȓ!F��p��H�\d��cI�w�j���}l��SFL	���+��V�KrL܇�>���vf�56Ԣ|��I������U"�����),-�s2$z���ȓk�ܭ�T�)txD��d�	8q�l��Lg́U�J-�S���d1�ȓt�0!�@�(pՎD����VẌ́ȓE}V�ۅ�B�s��%һz�����P�#���=g��q�l�8,K�L��C(|0���;]��iEn�3��0��{uJ��H	!s�t�b�0"�M�ȓ���h%�5�)�э�~Bp��ȓ#4x�G�G����'���� ����`Ÿ#�v4��P�j@<�ȓ&H�Z%
q3���؁X|�$���i�� �n��e�ϗz�Շ�S�? �5+�Y�f3.a��&0Zsx���"O*%QW.��JL;�B�;eN��"O�e�&l��ă�rP��s"OЬ��l^T�F]'T�D��"O�����i"��R$�%(�h�"t"O��R�.ؼCڀBe)�VB�3�"O�� �Վw�ԭ(wF]���h4"Or��I~3�i�v怮X�4()�"O|�!�f�X�|�/U��U�%Ξ�y�MZg�(���PM@��I��y���	���b�+���ԡ5F���?�'	Z)p�JOj؉�EP���	�'4�݋F@H�I�fP�0���I�X ��'���9��fJVQi%�M3:�J(A�'HyA#�3�����CB/�,���'��(y��,�U�4S�Nn���'�n �qᏺT�A��e�*@��+�'�ܵ� ��;�S�l�$I��'������cq�@�`�9j�h��'S��ڴ�E1r�t�!�	��lPE���'�$	��ꩀe�7l���'!��� ��2�Є�N�N���
�'�h�a�A7s�r�#�hU-8r����'�t�E�3O��)B3�;X�u�"O����9w�	��D� ZG��	"OʝY�ՙЅ�V
^#u?�t�"OT!:E�C=T�!XQ��q���c"O��0�˼w�Z���.d�~��"Ox�귭�/���R�	�P��%�A"O��c���#,FPs�G5g�&�Å"O�M�v�@/S��A�E�"O͓2�xy��[�k?/T(+�"OZA��4���
�@�:JdD�K�"OPȹ�

Z����ga�,n3�J�Of�9���F @�A/<�� D�PZ���]�DY@��u��R�k3D�40�s[��Ǘ�7��)`�D3D�����4(��#עF��)p��.D��!��Vԑ��Ӷ`�=��+D���W#ηZ�*Ȉ�D�
c~�����=����$		��%;0(�7��D±K	��!�C�ar�dj���x�b��.'�!��T� �Wꗰf��Ȫ�����!��0C<�cЧ�'��	����`��}����ǐs���%jI1Z����7�0D�T0��ͤ?-丸0��>LƁ"!�.�O��<�d��Fb�-~%x�@V Z�K��ąȓ�䳲mE.= �����D�ȓs�0Q��CQ�`erq%ƺ1���]��4��b�
b��jr/3p�ܝ�ȓ7ш���l�h�Rā���,V�ȓT����E�չG^�p�M�1,i�4�'�a~rLJ%~\��G)��)4hD�ƉG��y��[����Cc	�c�uYei҉�ybC_=E� 	�d�(nX��,Q �y�.e�-��
����*���5�y�@KR�F��`9�`������yB
"OՀ���6):q��!��yB.Y4T�ᆥ�<'6������y�Jϓ�3Nb`ee�&I	2���"O6�ӗ-���θ$RLpp7&V]�!�d�i����rm�*#N$�EW�d�!���f鈔뗢@�t�I�E��
^�!�ί#|���/t@8⣋�K�!�� �5�ף��d� ��B&�LKc"O����1�*���$q�,u��"O؁5N�7n໗I��L��"O�m�Fe^�0$����q�R�1���5LO�PHN��{�*#'�M�E��"O�H00%�$��I�6e�6~��a"O���Kq�¹S�H�0s��c�"O:Q�-�s�.�bC[0S�4"O�,s媇�2<Ys"�y��qz""O�a��g�R���Z�B�*R�ԅ�"O�m�ӢN43�TTx�L�x@�u"O:L�w�'j�I�bX�a�9ـ"O�[�
����qdA.��%yB"OJ�)Dϒ�c9X��
��"O���dƺ|�y��P�3�bIQ�"OBy�ߋ��� @L�ղQ1"O�𒳮�w-�������hA�"O��1�ԩM��81�@�p�5"Ovlg�юP���Z�/ͮh��1�%"Ol���+?� �xGN�7xpX@�"O���@�J��c�mW�9u��s�"O0A�W�U09U�E�ď�^�Yz��'��?O0=ӆU#D���.�  "�E*a�'	�	�`4NYydX�y,�Փ`�,a��m�ȓL#��цn¸��)s����Ѕȓid>$�Ø�?�>�R�%2T��,E{��'���'eԢ+������^�"�)�'4u���Bm8@ʖ�c
���'��
҂�Q׈P��@W�*����hO?��l^�*Ԩ��Lݬ;��P2�(
B�<1���
vF��uJ��|)�@�Q~���ΓE焨���-���uF��D�����S��!�ۼC|][�>����(I���<T�4;�� �Y�ȓX蒌"A[���`�[eR\�ȓa����ĤiȌ��l׉$�����^�]�B�D�=�$�ꎋn����ȓR�Nٰ�eكMXՉ���8��'ў�|�aOhx�"ҬȖb�$���,�_�<1f���D�&Q�a�C/��p$f`�<q�HD�#׈�ڢ�w��ݰ�́s�<Q���	J��4��m�z�p��O�U�<�1iP�H�
��*.���V�<�aLSo~~Aa�Dn̚�I��NԟD��[����ɻ+��lPp��p�@�ȓ
�xl(E��"�8tz�/�~C�8�ȓA2�3ƠC]�v�#@"�kKXȄȓTjx�`r
&X��seJ>�&1�����q��	�$�→�@Q���:d~XXP�ˬr�W�(Ժ��1D�`���c���,�L��#D���dS�'4���-��c�����!��O���4O�0��gAy�� ��
��Q�"O�h{�&X+JÜ����4�^���"O���!��}����	G��d"O�4���k��ث�"���s�"O�y�D��\��!��k۲i6֥�f�'p�'/�)�'2���j�L�&o��6��*/ZU0	�'���9���lE��#�jѸ^nYو���O4"~��U�`b�;ХL�c&P�(%OQN�<���
(M
��5C '�}��fJ�<ip���|��Ȳ�F]��U��M�}�<a�'��^���*���UU���1�ZD�<�� F�&} ����rw�����v��hO�|�� �W����㓠� ZP���� �S����]vb-i�� ����]�D�!�DMr����g�6��1HWI�%|!�DW�\,����W��p�i��'i!�Z?�|H��U�"�{�"L�h�!�DV�S�M�p�¡^]�Ca��K�!�D
�"�p��$����T �ў��'��y~�l�4P�fؐ��W�~<j[�.F��y`��hሹ���J�cNP!e�"�hO���)��A6B<�HN2d�$s�IK�N��g������U�uut`HS��..imB�J'D�����@�.$0� (�!B�0@�&D�(�G/	?�L�Q�.���ء��#D�,z���-F�\P��)�IZ�mʓ!�O��>ڙdb�)l��l� ��6�h��YM�L�B˘Lc�ˍ
f���ȓ`$đ��D*6+�݊��/���'�a~r"X� n�)st��f���1P��y��6^��Q�sc�0/�d�h���y���2��c�I��'��-�&
���y�A�=��qzpk� �0E�v��6��>��O��!ECTc�p����]�EӐ"O��y��G�/`�d����.�M��"O> ���ٱi	�pF��G*N���"O��at��+�����s>(��"O�"��CU�,��l%y�b�U�<�iL���8�����u}�𓵣ON�<	��=�|!�BV*6�XtH�J�'a�4�J�f��:@iԸF��\�����yb�3l�Q��"89��9Y��Y��y"�H80^�m��E1��f��=��)�O>�أbCY*ѓ�Ř� �n�Xc"OJX:�F�2_��=PB��
8�����"O*�1 ��+W�����@����!"O d[C�M<%�,�1,�`s杲�"O$�`%��X�⠊+�d�(�ɗ"O*8h���rh�1H�V��ꕋל|��D%§-�lQBsg��U��5�F`
8J6a�'B�	S���IAM�N�8b�L&""& k��0D�8!��
pp|����͒��q��l0D��x@~0�0�Ɍ&Q�5!�!-D��Ã�-�L�fn���&����/D��hE��@eSb.��K�<|��,D��##��>V�t�u��/^��f"*D��	ЅU12�BF�W��t��b(D�\Y$�݉,�z,����$�\R��&D��@�	G.>F�=@���
q�	/.B䉸J�V �Ҋ�@F�A9��Z��B�	v���*F�["68i6MK#4{����&?!��N�!�Lt�m��t��H��
v����D%ړ�����*����W�@�Mm`�����ğ��P�!,� ���h�\�!�C�}`��t�� j�P��\�X�!�٥
�$�"�hQ
kwnd*�'�0�!�0h��X���ө)jT�� 7~�!�dHF�N�͌'<e��b�!�nl�	��?E��˕�{d�c��ֿ>�2][`��)�yB`�`�q5hR�FL��q��ޗ�y��[?@��T�60qZ4��M2�y��3h�����&"&:����Q��yQ*���+q$R�cҍ���y��e>!3���8� U��y��
o�ШfD_�}�8 t�Q���D�<AO>E�T�۾;  $�W�0l6�S鑯�y
� |�)d��v���RPK�]R�P"O��ei6G���I�)\/pB�eiv"OB(
�H4d��}����2�8�j "O�{�J�4��\�fZ7.�:U""O�J�FW#f�J�E_�ZL�"OF����W+�����O2�b^�����%��|�����:قQJ�ܲ`Ϡ��So�r�<�αd��yR�)_��#�KW�<��O[�PQǭ#AAF�:U�Tm�<Y"J�T�cOOH�R���A�k�<��V��q��MR-<њ`I��<Y�
����J&�Q(O��!F�{�<9��	�Pq45�Q�(�R�ɤ�y�<��"G����B`�L�c*����z��hO�>���V�T)l�b���JE�|�����:D���0͖&�-��C�;]$��j�Zv	��mӼdAA#Z�t�ȓ2�����3G��7OA*;���H<�}�4)� ���V��vxX��ȓ7����g���|��I��Q�؆ȓQ���l�j=�FꋆZ����?a���~�&�K�In�8 pb؏&��q�Fbk�<q�F��;&IZ|�V�1��h�<9�j�u�$ܡ�&�Qޖ�D�[[�<��Ȍ4_��U8g�_:}�����V�<��ʑ)`����T�ʊb�"���K�<94��<�&�%ʞ�Bin5Ё�N�<�j��_�Hu�ч�$E�哆��J�'a��CO3�6Eѕ/�,zD=æ�ƥ�yrKXH��IB𩟛6�<;KR��y�H{��D�e뗄/.�� V5�y�׺�n�`�,�//0ݳҦ���yb�M__p��q@I':(2�����y�g�<	f�1r�hs��2A@�(�yBmA+��!�C�Z�pxPh>�yR��3qV-V���a��.�y�M ��y��$�#JI�ēg$F/�y�kW�V�b�@T�[2;k�" L���y��Z�1!��k
�1ؤ��N��y� ٣;�0����(��L����y2Z�<��l��FL�o����L��y��](%�Ӣ���<�� �9�y�/~��\3�0\�~�tM� �y�%� ҄ô��( F�e@�(�y�� �!h0�2�O%%��t�CL���y�Գg�� Ѥ,		&� �h# O��y�J�,qiH��.24\���BS��yo�>|ґxq�ŧ-�8��$�3�y�LP��ɩ3a͙"/2$�Dg<�y�A�17ό1��j�UZDO���y2j
�)�ث2�ޡ
z��V�ݏ�y"�?h ^��CoÏUg��a�H���y2�&P�DX#	y"�2c��y�Q�G��� ��+_�h�[!�Z��y��˜Y �Q�ǎ�PԆ���y����l���u��F�&I;1E�7�y�H���i���9ʨd�`�"�y�H�I������P-�>]c����y�M��?��#@�6�30���y�%]1>��ٺ��G�3��R �:�y"���B]��dD�|��)�D�ybDM�UT� V:|�la��P=�y��ƧC�2,y�
�u�<hZ����yҢ� v�͘�B�n����d%�y
� ���uX�[�����?[��Y�"O�������(��잉`���"O������<�a��^3e����"O���&��j�mSaC�����"O>���M�-�j����!]��5��"O�t����CH�����7y�v���"O���@�����G�ft��!"O��h�OHp-�%���ӿ/k|�S�"O m�ХF�}�࠲�_;��"Oj���kўEѶ���� �$���"O�dK�J�b�3A-�%$��be"O��"��fL���m�E:m:�"OT��F�Y \3����L��/��(��"O��ĥ �Oְ�H���N����4"Ox\�2Nѡ#/j]�ɓ��
� "OXC�\�<stuc6ʆ6�,Q��"O:��6%N;��C�T�ܴ��"OƄ�t���E�(���	*U���b"O��0 R4B��Mb���7"6�A3�"O6d��JU�T_(��F�LC�"O*A�P匽W�����!8�Y�E"O�\	�fV� ���1��� p"O�|�#��wh5�)�<�� a�"O�٠C�HzƲ�8��I&Hsh�#"O���u-7K���E��^(�`�"O�P4��7C��DP��6]>*uA�"O�uxT��`�2j�i����S�"O�X ���'Z�=�PI�!�pe�"O�dZA�G� 	(כ-Ѵ8��"O l�ō6�B�t��6w�zt��"O��"S ��(@���H�BT�7"O�<�"% H(���Ϛ<����s"O) �Q<�x��h]�+���#�"OڵY�J��`$�)
���$�"O� ��iX�T����V:�z �"O�āt
:}� ��F�
�a��"O���@î��q�
)5��w"Or����d����)ȫV��̰7"OVE�C�b���	V�R�"Or,�v�M����(Ob6��xb"O�4R�� � ����r�@�S"O֩�V*�N�J��7���g,�P�"O���7��_��yC ΁�m2�P"O�ڵ-��伻�Q&�@�"O���Z�o[�O�fbL�"OLK��,1R�A=VI�Y&"O�H�욈A&����C� B���"O�	c���?�Xpy��Ƌo���"O���e��ʝ��`�L4]�"OR|�p��,Jf",S��yښ�
G"O�pH��'��@�#�G�Ò!��"OxQ��[%Le�V"̔?��}K�"OR蹶蓖2;&�h����ܳ"O�@"����6� |r�aO�<�&ah$"O���W��;���J���e�
�!��]%I��[dNҨA0�%�(X!��,x{���l4TțF�=c�!�d�B�{�c��N8ۆ�A�c�!�dG^V)���X"U�\BWcS&f�!��S�;���0&���M��� I�!���8V�CҤ�.���R��14m!�d#U�&��� ��~�� �I�VM!�DS�G}2YI�a�]v��FLU�S/!��ԍ-_0���kH =��*�ۥp�!�� @���dE�Nj��q�◶J�pC�"O�u�Ȓ�D��cAʞ����"O���w.��Dj�L�T��s��Æ"O�����T�B�DS� Az�"O��	��$D �m�"jH5�!��"Ȏ�!�E�,-�P$�R�㺄2a"Of��wb$���׋�t��"O0���͒Co�p� ��*�^��"O�	��C��Bx�Qɴ�r�J"O^ݡ�F�@`v���՞e��)R"O�m��d�5G����� .�x��0"Oډ��*4�Z�%N�%��Y!�"O�H��#��dh�4��$�	��H�"O^p�M�|��j�A�]4h�"O�} �L;G:fݲ���+n$I�"O�U�A�>�	�B�F�c�Q�"O���^��)��`�M�Na�"Oʐ
�
�b��5�����(R"O�%Rw���y�\ih��O��]�"Or1�I��,{vEڔV�& ��"O,���^����<%h݋�"OnQ���)�>|����P;|�a$"O��b��E=p!���c��>pQ��"O��h4�ɲB)|�Y⍃�4T|�Ã"O`E�u��)X��eLQm'��{"OhX�,�r�����ߍ�nZt"OBM
�Lȴ�)�'ɒ3���#�"O���r���k�)P���E�N��D"O���
�7���d��-e���"O������s��Y�j�SF���"O�кq�M��V�ŏ6=�}����yP���TC�4��B��y$֓n��P�L]�$����&.���y��߲/����s�< Fq�栌��y���4`�8����
Xaq)���y���i]-�F�X?��Y����yR�A+;��"7�����i@��y�.кXv�C �N#��DJe��yb��%q��
%"��	�����yb�ސv
�U"��c�IP1�@ �y2ᙀ�v��M�]q�E!���yB
k�4��� (�홗��y2	ݖ
�(lX��6f1x�+�!�y�d�Y�(��o�-#��z7k ��y�G3�l�
�*,<�&%lO_2�yR@T^��{���'j�q�+Օ�y�b�%v�;���B�M+�yҠ_�8k��{�����@���y�d�YX����
�,��R���y2h�Fp�( s(�/���
��yb�A>��@�K K)��1$��?�y2ʔ�R6d3c	�IV�%�Z1�yB�?`xX���9J8�)�я_��y�]Ud���Q�F���ځL��y2��'��T	��ʐ'z��i@�՗�Py"A�R����@Όn{�8��@t�<y���>����#�J�<�I��ʟK�<1b��9?���z@$�008�qy��Mb�<��^!^��iK�J&<qtcT�<9��3BΎ�8�j�%n�؀+�`�u�<�c�
'Ғ� C-^�_���I2�Fo�<�mK�r�� ��9�~yQ��C�<)��7.\$���PT@@�%KAB�<1$Lj>�h�΍�\�\]p�.�u�<� d�ڦ�	W��,!N�GkR��"O���d�!H]��O �0M���"OLl(v���b�ĉ���3�"O2i�������gC�gV��"O�t�g��)Y�X�k#�l�.<JW"O��q0#M�A�$���GG�,��H��"O�9��-?��|�&��)7` Q�"O��u�J�"ě��# 3,-�"OԽ��YT��q�����7+Ό� "O����Ȏ�c X�AR�N:q<��ٷ"O0H��d��I|́��>"Nn9�r"O2�Q��[:!i��U=i.�	!�"ON����+�L���\���Ѕ"O*���X%���*���F���0"O=��l^�X�A �A��H�� �"O��r���#2���'�d䒀�A"OZip�Ə\T|��E��>@��s4"Ot���A�z��	��°ư�)u"OH ibݧer���V�ŋL���"O qp���/gt$�Dō(<��"O��c&G����1�X�T	jlئ"ON�z ��D< t� �
��R�"O0с�!{˨��� �	�~���"O�l�p�Ӽ}JXS�@�1�Y�"OZ]S1���6��4"/��b1"O�` �*�F�LkV��:�`�@�"O�a(�/�7��̒ܳ��H�"O��CHG�lt�#���"���H�"OФ��웑IO$�c�*�����"OR�	�
�g���9�
�)t��!�C"O�2� Jexڀ�c�Hc��y��"OBqz��ƄAC���Q��/���"O ���@
�uB���_��h(S�"O� ��P�K���`��h��4"O�$gB1��i���` �<��"O� ӌ���Ɇ�M>|�Z`se"O*���K�e$\���NE
E�p�y0"OZ;��H%UxMڵу:АXc�"O�-jՌ�%G�P ��@8<�8���"O\��1ϑaYM�@.X�R�H"Ot��g���Hyx�x���1>*��R"O�e�D�b�LM*m\�-��[��'q�'KdYh��W����R�(�*"�(�j�'8�0�1�Ζ'�4�z��fDBM��� �S�$��r��a���f�F�x�l�yR���Y����	^�Ơ��Ƣ=E���x�{��E)w���8�ZV)��g-ؽ����D|Y83� :w����?	�!�O?:�(��ʿs@�գ��s؞�l�_�ɒI�D���d�<qg���[���C�D��� ��<���兘�P�HC�8Y�N���>_�`�w�B�1gH�1����R��U�6T��B�I�l�4���
�B!"��2��	�fB�I�iP�03�&̈?A�C�"�8P$B�	/#�dQ96��|!�u��&+� B� <^<�̑�EP���.��C�I
+6�����\�D��a�;6��C䉤ue�d�,
A�l� �d�� ��B�	bM�
�����#e��dtB�	nb�[��C�4��,����~B�ɜ��h1&�2�8��G9(�:C�	���݂�D��<�Z��U7�B�I�h6�� �3&�1z�|��B�)� tEy�* �pK*hxMQdۘAkS"O<�Y���L͂�"DAg:I�"O\mS�'ɱ0U��ip��K|1�"O �A�Q�;^�ɠ�O WfT%a"O��1DHW�l�h�7���w��l93CH<�pɆ$<�(
S�J#}J���Mi�<I�%Y�����!z5�	���n�<Q0�ǔe��P-�P�Pao��FyB9O�L���iи)��\�Rj�7 �	�D!��!򄊪2x�q	�`�"�[Q��+��I�HO�>	�CM��@��׋4�P�k)D��:��	p:b��$�X�[����'D�b��
i��S��W�Q��`+e�1D����+)g V�C�c[�G���ySA/D���Ā8l��peL97nZ`��-D�\��g�_�e"w����я*D�$�"��%.�Hz���
~����,D��I���I���"T��	$ra��+D���!��%�l�D&E$����)D�p@���=븨)Q��4���
2D�8�C�H�/�L��$$�* �����,D��0���N��@�d 9`��� )�OO�aK3Đ�@�ft�p��pp����"O�`V^�P��N�?hT;"OZP�t�S�uE$�RR�>I0�\r"O�|@˚�=�d�k�PXâ"Ov�Y��)VT�k��Ԋ#��O��5��_ԄZ�ÑP(:$�b�&�|���㴔�s���]	N�K~���t~B�OV��6ǂI�*|{rܝj����w�⦙�'����<��'�.��G�	�S)�JcmH�{��ɚ�'��t�a�K52T�ۧ�4���7E%4��֋�-���j�[CS�-Ӵ�+D��X�A�`����ė�y���;1O�����'6ފA�Ȕ:`,b �Eo�-qX*�OF�I覥Fx��|Ή#)S�x��d�9K� @���ʿ��<)I�ȕ'fZ��s�D42�p�̞3t)�]*OVʓ�hO�Dnj�
����̝#��#4>Y�>�E���E����B����D5 �mp� �	�HO�܇��s�<uRi��"��1�)��d��	ӟ\��L<����#��e�Ҩ�A;� D�8	�ua�X��(X�0�Z��W�N���t�<Iߓ3$bC.ٖ)����
\L��R≽Z�^�{����rk�y��� EXB"<)ϓ=�Q���J64����T�_�isDyb�|b5I��X���+QN�*;Oa�r��y}"�'���E(��^a^P�C�g�Z�����c���q��(/j�Yb�/ٺ?F@B�	�Y_LxFM�;����eZ�w(�O���DJM������� ���͖T��`D��.ٝ),�]����8Rl���O���;�S�Oܘ��b�t%����I�ǌ5���D1,O*�)jZ/$�L8(�g!'n���|R�'��R�޺X���C�t�>�"�O�=E���	=�@(3$?�@@M7�yr̔r�\]B'�E.3i�'���D.��O�I3SI�]o�0�A<P��`V�If>��U���`Qb���c3��z��:�$%�S�'^�y�A9}AP�D��jF����/*ܪ���& x�D��*Y���J��"��*����8~a�ȓ y��]�d�b�ڲ��R�<��Ș:qh
d�V�������ȓ~^�q���Zi�BQ�c)v�h���S�? ��y���!���X�HNG�hY��"Oz1h����
�i�%P�a���qǒx��)��DB,�k��U�0yĄ�@��I��C�I�	�yrD���<J�y	��*;��C�I?ز�@�d���e�7��(��C�	�6i��  �Av�\��B�+�C�	�u48&��,�ܤ��,�f����d�<��4��Q��ߘuu��lGu�<�A⁲M�dx��k8T����u�'O�?q�N׎,�v���0�°�<D������F�.]�&���8��9D��:2��?MP&�k�@�z� L�w	+�Ov�'IR���,��A�a542H\�O%����S�)� X���&)p�Q�Tʆ �(#=	��T?��C�4�����%id���>�*O���$��egl`�I5u���ɚi�a~"bM�j��ǜ�)�R� &eąi������Р�y��8P��u�è�	lNn-� �O,�'%Q>���a!"dz��W!h�Pi���=�O���Kylq�6=��X���)MNv5D{��9OZii����C��p�`ٸC�.ӗ|�>����a{��1e�/I��"��x�	�<a	�nj<*���p`HI�p+G�7A�=�k�D QQ�N�V�2髆ꞗ8�p��
@�0�7��4Gu@P0N_�A?�iD"O,MP��ɂy�N��c�
�AZ5�@�'<������S�#.\�y�l	�"�*�+D� (� P*mZ�l���U�}���)D�P󢥄��! ��M���%D����(@�
m�ٛb�A4���$�N}"�i>�"֣��p�@ �7l�)`����#D��HU�E9`���#�*�e��H D�0`p��_��-	Y3|�@�2"O 9v+		�|#%d\�qBQ��5Oz��$;(*�$��
�' ���GUx�!򤘞��-1�#p���R��Z?bD!�䑃Z���cp��,�Z����!���M�L��%�tQ��Q�j".�!�DUdUx�7�_���t�Щ]*�!� 0J~� 󦉥F�Nh�a��M�!��OK���7�DX�I۠I	0�!�d�|��88r��@,hYT(� �!�ĝ�XwZ��e�I$+�����@�!���.3���,r���ȃ�O�!�@�2,�p7��{��T�q�
�!�3~G�䑐c��!A�F��.C�I�+M����R��A:iW��C�ID"��3,��jdMt�)�B��a�`� .6� C αk��C�ɇ.��iZa�Ù!���uP�.�C�	<	8q�N��kHܴKs�̢*R�C�ɥ:�@�J�P���Rf�I(w��B�	E���t�O"t�`A eDE�L/�B䉕1�e��C�\Z6�h�f��&��B䉮^�A5A����D��("RB�ɸ2д���(�&p�����^�]�<B�I�J�t�#�� ���i�G ��:B�ɍ Ԏ�a�E�!4��%�s bfC�I-k�*#J�7f��!y*Ʊr�PC�I�k�����-�_��Y���A-=�C�I�%s�̰�l��4F$`r��@<�LC�ɓ/���aW'V�F���
�� �!<C�	�F[<���H�,p
ԮӤg�C��;b����ԀÎ/�"p�R!ҞwM.B�)� �1됬[�I�����4�jPȂ"Oz�����? ��f�6t�f��u"O����/��T��8�&6J�cs"O8�)��ؑ
��H�"l��4���"OF�I�bW��Z���KI�$d��B"O�;�CC<etT���&�h���"OvX:��I�g�U�8�f"O�u*P�ǊAŲ�F0j�ɚw"O���j�)����G��k�"O$2R.���5f�7��	H�"OTt��L�Kݾ=�E"������p"Opy���G�45�a΀a{����"OY�L�*��0<P���$P�yǺ�8@�'�,y �a@)���K�%,f���	�'i�q��-@�c8 I��)%�z0Q
�'��5B]�R�0�����8��	�'I�lc�
��u���I@�B�'�0yałR�K'2D�!-8)�~I��'�� ��oY4�R8y�W� �j��'����⊤M��a�2#.��
�'�Č��hȥY�f|P�@������	�'�tjU	�U���2��p���'2����	&F|$˂�κXA�Ԙ�'����.�*�@U�V#�d���'������2ڶQ2e,4H\��'���4h��l$�PXp�6g�(��	�'�0{a̅
7a3�쟣UE ���'�Jp� ��Z�Hu���P�_�\�*�'[,�yA�Զ<�ڗ��Je��h�'���1�N�!�2@ 7�B����0�'Ř��~��x�bB�;8-n�1���O�<�4��#O�Z�q !ʳB�TS��AA�<�"�T	/��8�R�J�b���E�d�<�.ÿUD\hφ�E&f���O�\�<�4�<lxz)[��PI�x����a�<avd�x��U�@�8�ٰR�X�<yt�X�+�ʁ�v"�:qkH�Ȗ#�X�<!'�]�AŨE���ȣB!���l�<��k̀`������R�Vs m�g�<1��(P14,�F'��U.�i��#�v�<��Ž+,,���c��[�x�p��8�	5)Xu1�Sv"�hTֈ+��<�h�=o߾B�'5��� ���h�4���-�,��mz�!�������|�'iBp ��w��Z��F�C$p=��'��u@r�� ;hp�&gőf���'�����Fw8� y�" ���a�.�n�i{��>LO�x��2ָ���'(l@��c�#n�����	g�$T��'�$ɺ�g;�>��aD�S��IȎy����V��y�6�l�O@콉���=�HP�#�^�=���Z�'�Q0PB�. } �!Ղ*r6���"���O�x$�3?���L+;nD,�SJњ!�ʬ�b�~�<i�!/Nx��ʈv�$�"\�Wd�9�"�y����$T+(r�y��lN�|oq���,Raz���3�����ʖi?�a�:^�"�ʐʕ�<<u�S�D�<���٘mm����Y�g�zع7i^�g�p��G��K{��~�������̕�p�u2/LT�<��ˢ��b3'I~z��0ab�}l�<:��|r"I���$G�!\��p�
,'�Q��;%!�ܾ%��P{��?��t�M69����k����I%^�n�kS�Q3ye^���M�<C�	�k�
�a"'�2N>5���	��B�I��,�� #�	3R��xDF�6\�B�	�'5Xu��́���؃���#�B�I=��HP�����?�\�j��y
� :afL�=N2��ғ"W�?zn�p�"O�1�W�_�i�TA	"*[�]l��J1"O�a���!e��ų�$��F���"OXY�#NOhn��`hY�R�����"O:�Q���lM�§�l���r"O ip�3wג��� vf��"O�����Y�ڙ�Ƣ�-�.���"O�XRlN}�zqITa�0z����U"O|��d�J�F<
��Ӡ�4?�u�d�|ʹ>�q�=�}"�%�?P���{uA�'\����D�	R�<)�/^� ��Ơ�b�HS� �fU�Oj��OP&����E D���)+�PADF�{ m����E&H��U�Ϡp�Ci��W�*l�B�&J8X���l��=�a}�8�N��%=�	#	���O��FBЎ�t<�!��	Ir~�S��֘ �莬K\V A� ��B�ɽu�@uZ�錎�ƅbK6��Ld| W�T�\f���d�Ǩ���4�I�ڬq̃:F:
��"OY�w��>{�Fk�F"�I�#cQ�~����g��m�ΕZT�::�g��lx9�B͇	��Y�L�
aԅ�� qB0�aŗ 0>��2��e�z����B*Xfn!RCc���B�A&�'!�����!a��c��2y�(�����VT�z�LV~�}V/Z�2@�I�&55
QǪFs2Nba��_T!�̺x��;Sg�6)�pba��(rP�$K�1p
I�1�	$Jx�j�E��{��}
�T h����ě!�)���~�<9�.�R	p��4�tp��8B�������;L d�q��N�${��(�.�S
��Op,�-f��r�K3d� R�'rYt��+&�O���CX,]4t��cU�X��8�g��.�pts�BW4Fy�u�́~\���Ƿ�?i`��&_����AU�,�r��>1'���T	T����J�O�������r��x�c���g��0���F�A�'�:d��4١NG����)�;n�$b�ϺEÒ�O�L��˶ሣu��SÓ1�$*��L&:j[�;0K�9�ɠ ��!�W3�v�[���2�("�O8b���94M� YӠ� \tPQ㥮��
�2�g�;	ހ=�%��u<���C�t��ňwe�wx���$�
�,`Si�~[�-+g瘫F\,��j6s��ŸǅX�rt����D���}��
U��5����^����iX=D��{rK�U���ī�S	���4B�kaz�8�HB�l����FI�M%2�Fֈ�0�vNO=l��訔b1hgp� �؟�I�J��,4�����;����d�����ȴ`߈ih@j��t�]�,o> �%'�D��&I?x'03�� 3�byZ���v��=~+D�;O�蛇��]�B��(	�.�}�X�@�Z�Y*��wO�b��䓯�*�2��	=}�[�^>I��ja͉�o��H1��
-b��t�E�Ϊ�x�c˶>
D�Z�<��5@ݦV9�|�������� H��P�ez��K6=	D��.�>��"U��'Կ���ٺo*0�qEc�%xL���DW0��=���H�h-��j�;mI� �S�4�,jJ�O"
I��L"8ŢqAs�3r�����M�0�lZ5��g}r�C	H��8�#�]�T���ʾ��'��A�c̈́�\aQb��o���V�?����\�^��Ԃ�zq4��W��O�}��߈I-��7����<1�)_�4+��B䆐?Z��v"@?Q���-Fl����@�m&�G��'\ �S6$t�1ḼcU�� �CϺ�yR�/��:7`�M��tJF$���?���	)pب�ī-lO~Pi��٨��cU�W�Q>�K��'��� �]%>rb�@�P�	���)e�P��G���y�aےd���C�4Zd��茅�(O�P��![�e��#}����L8�R�.H�i#�
�i�<�S�X�`���x�Z(K |����T�K�\'�"~n� _���D��R">��B���B�I�]:��qc���C�
]�5���i�����%(��PazM�w��8:qkEq��8Xua��p>���Շ0�`c"�ݓ6��ܘbLs}��b����]�FB�->�~D�1	�Hy����X_;��<��/8�fl�aI9§2�6���"5�(R�Ϟ&c� q��X�8 Vl�sM��9� �? `E���Ke��9a�OX���OfI��L�W����7�r�X��E"O�!£��Y��&ꉍ��e�"�O�)���4WEb�ӓ�T��Ӯ�S��T
�l�;Ӵ���_�`d�B�:���U�I�@^A6�//p|@�s"O�y��)�L���BA��,3��2��e�ga_(�>� �C�.�t�QL�}�l!Z�F>D�� @E��a�!J�.e#��.j�4�׸iX>|�ڤm�ɧ����m�r߰���瀛/��+��K=�y�)�+ޜ%'!��PDd3R
����D�i�vH	ۓ~�T!P�5�!IЇ�E*)��J�d�Cפә*���уM�KF�`��I~�r��ǅXz�'	�j�0�ȓ8���dC�1z:�*�@�$�,Շ��ޠ���8z�,q���<r1E{��6�`�i0�DuXh��3�>ls��&ÊC䉡�$)�B��+�����Q�BZa�3*����!A�}}�!@.L�J��23E_�H�͉E�>D�aE�M[m�%Z�aZ4+d�0�z�걉0M�G�2P�ō:ay�&ܞ(�z�����lj����N��p=qc�f$���3��us����dM �x��Z�f����S-��xbl��PqKv���S�8EF�� �'��c� �;f��HHDʚ31��V����>OΑ�0���b[BEc�"OR 񢥖����qD��M���]��b����!4g�������<��
J;c:A��O�d�^-Jc��T�<�l3I�1��*JH�X��.//�\-���09=���DdM��ay�F�5	�M�!nɭWE�����5�p=I"Փkbx���(�,x��G��rm��:ABҿq�^�ru(���0?1�S%?p��gG׸Z�<�A�)Y,q�	��.��,s�Y0�ϐzqz����\�db�:��;+%�QUW��DAF}Rf(Q�T��B��6yY`[4��*\�f�閥��}rJP�W�7G�r��5Hv�@�W�<�Ec� �8�9�D��&�fm�"�I�<0*S J�BbO6}��)0kv�4�4-={�̲.â���K O�����K,Z�azr�����S"b�5X5|xᆊS��ķh�~РB���ēn�~����OjX�	�v�C�\�qty��O�%[�2����,J���SO���Vd�U�F�v��IAT*�F�
-(I<��hT�5jb8�D(��C�(�����h�h`�!E|���0~�`�cőUܧ5��:D��-h�=b��X6B�h�h��_�@�ݦO٪��Y���!(Q�%�ܭ c꛾fCRNb��p҈�	6���#��>E���Uc��hq�&� ]�5�����M�@ޖ/+Ь�o?h�)W�N�+�>`���|����'U�e�T��8�f��<�t�8�d�{�����H�R�+�1����V��%�#���$�����P)�d��@�ޙT�xZ�
O*�{V�A�A�܍�!�|�Vx��	�fA00D��x�'E�@e���x��D2�O'�@��ȓ��S�ׅ~}���6F�R"���'�*�����w�S�O�{ �8Ĭл�"t�t��'��l3!ė=�	Q%C�&�����'LD���^pH4D�)�D��'RY	�@J�W�>�Y�&M�%yb1��'d�W�=b��*�>�p�)��4D�,���L�Kh��(s	�%J:�� 2D��#'*˲P�
���ψ�D`ԙk$M0D�pҵ�H�F�d�7��gsNu�C�+D��EkT�2�(:�-�(�$�-D�<�G%��1�{Ў�0dP��閎+D�0)C$�]ݴ1H��@�?��df�"D��	�),ra,=
�j�qܨ�n#D�Hا�O�t�hQ��%_(��i��� D� �斚"duzM�8��0{��-D�0����q�4�pe�)|�f��I!�Z?*$\����N�0�%��?#!���y�F��eL�x 0xJ3Ƒ��Py�c�{V4��3�ӻ�Ą��Z��y�@K����@�-X�e�(�6�ybD�as8�0� Ӧ)�l�X5�P��y2�G*:���b�])�PȚ�o
�y�E�)�T)Q�V",�H�����y�mA�`tr�JA6#3f�3����y�G��]xQ�Wò��K��y�i�'.p�)�`زR\��Ӣh�=�y
� �)Ag� 56��V��4#\Q"O��D$J/	|������W$�""O�%��8)<�DB��X�{�"O��a*�e�DD���Y�!�d"Ot3�$U!k\A�`�#�6U�"O�-����?&I��O��s�-C�"O2$��"�����c��DN\��W"O���b��|_����_� t�ȓgb�؂B��-OX�۶����<���0� >6z�A���&of8�ȓ(�j����ٞ�iJ�L􆰅ȓF.�81�A7&NL�y���#�^0�ȓFW\�3
� )�'įt�"8�ȓ(�[�f«s�Is�Ì?|6����FYh��_,�r{WKБ?�ȓF��`�Fe Sd2��ҫӥ��1�ȓ7LL�%�j@:V�]fu�!�ȓ)�4j��ɕP��!f�S�oE��Fo�(;�JD8�]IëG:RBe�ȓm�"�����5�ƕ��MQ�r����ȓ98��"L�+qV���.���^=��q�\i���N����V"�؅ȓp�-3���E�Ryu`�\�D�ȓ{��r��5-�a� �l��݇ȓV	�-#�V�WJ:��Ca�x/���"ޖ�����R�z�+4e
�x'px�ȓkZ����&Q/��'CQ�x�`!��iBuaS��U�&y;��"o%TԆ�=΄�(Z�3$+���5I�`��Gd��ؒ%��e���1r�j���fW�3�k�);��� y�������.H��IA��ʇ :�ȓN$r��# )P�^��w�Q}Nĝ�ȓs��Œ�B�*����L'vu�ȓe�t#����$	��gB�s�Z��ȓ�=j�CX F�}�w��e(`܄ȓ!�$��&�D�X?̩@�X5��E��27&��Mq��I�BP2uB8�ȓE�rL�W�S�r�B�J�6�"u�ȓv�$��D�
�Nz�N�<����h�%�\�h1u ��Z�L��ȓb����փXG��P-F�����>�X2�ʔ�����䔍� ��y��UZv-,l�ܴ u�� n�C�	?v`X��"
J�"@��G�sg�O� sT�̥��F;�d�Q�P���OP'lE�"O�4{6�'��Js�G�%����2egt%%����<!��8m�>��GI�?����T�<�@�L?�AJ@������ِ�p��c�%V���dݟLK�ᗅ}h�� Ώ�$�az�KB?>�h@���R?��K� m����M�<��a��n�<�K�Ex8�,|��d�7j����<�W�5l�����D+�'j�|� ��!o�����J(X�0T�ȓ*9���1��%ej��5�S����b�,&��'�:�я𙟘AUf�S0��BaY' d�1�)D��J�
͍B�, �+��c�b	�V�+���8��	�r��|�*��+G�0g��3����i��0=� %��x�t ��J3hS%��0
a��'ՒXAD>D�,�$�@_`<D�Qb(g�����?�I(f����I�#I�Q?}@���6\��1�G��Dt$xqf:D��b ���FS
��U�N�D�;�aث��bL>1��8�gy�/�1W�@�ғ�R�J���)����y"!	�����R�ިL~�I�$�-�M�`=XXH��ןx������E�4 �ʞ+r�!�� BpZ�a�7i�� 7f@��ֈY�"O,T:%���rmtLpP�[�$?�AJ�"O���0`O�D���Ä�,,�(4Y�"O�� ���tX��3��tĶ�k�"O�ty�
ǬW��pSa�r���T"Ov0�w�O/�bAQ$���x����"Od<p�X<���� ?fRH�t"O���[N�f��Q�U� N����"O���Zcu���Q�Z:?RP�Q"O"Ē&��MX�yf��jLx#P"O@�{7H��{�.T�0�GP&�-�"O�4*R-�z���g��
Dp	3"O&<��G.I���5Fo<���"O��Ql݌o�V\�AŖ�@��"O��,X��^��*� $̄�"O��"�9w; |QwjB�= �Qq"O����$ص6�v�q��F�mpt"O<����%bb��iG��	qF"O> Q�	JBѴ����C1\
�!rt"O�-(RLG�_ЦEa�CMQ�j�C�"O�!�f��	A���h&z�X 7"O�\�A���k���Hvr���k�<���%M�	�kI�Y��I�Wy�<	�M�3~�0c�=����v�<)�*�5q+Z!��B���@\H�<a�� :��s%�	n�P�[��RE�<9�W�m�B�z#�� %�t$Ii�<	V@��*�G�vo��K���d�<��e�1k��+�ǂ[�`�9�x?A��ؙ>�'�����Ӳ�5���'|���O�P%�i1����n�1�����w�l�AED,c���`s茝
��gdB�8J>4j��*6��̉P�ϱzC, ����O\�BS�,��>Q�Z�y�ؘ�ڸCp���G�
k��W��MY� �4B��	WH�4�O؎%8e`�/h�D�(���\�NM����Q ��V�T
`����IT�0<y�CE�<D S�T3Q� �ŅڝE.����4ZS��ԥ�.�Z��[ e��@�shA�5��x��aK�R$}�`��f4�aR���x�"�H>�f����@�f���?�����i���h0+Oi��DX@�J1�����p��O����ޠn48�j�i���E�ɭ��=�f�_��G�h^���5f"Yb �a1�
P �
���Yi�5���Y&��@@*sT�����,O8���σ�&w
1`"���Y3�$��=a�A2QGA�<
2n ��#lڴp'#�s�1�u�\�d�!�F�	q>�U�ag��^{��56O��
��b���q��4E�ջV�S��8����m��OJ�O1F)���I�~���j�x�4Hr�z9|�i�'ȵD2��7��A<i�C��c��@� ��4,���V�
�N$���K�3P¸�[� b��l۰���(3UlK�|zVe܋%�
L��D0��������a����SŜ
q]p�Gfi���ED��6,�����:rfd9�����YFF���/s_r�?�=K�l���14��u ԁ1H���?1����Yv� �M�bj<c?A�C��'�T��%3[R9��OZua���_�R8�u`��<At���8L"�P:*:�GʘFъ�ۃ��!p"��h��dV��[DW�!��e�� !��Q�Э�E.��tw����0]��A�;^���y''�A؞����C-0�����K�FI�f"�OU�gꂑ7���X�.ĈCg�����Ȩ�`׼/�!���z��Ğ?T&`9�K52�������?K��j��$ҧ�0�`RC=P@���R蔙itvфȓ	��q����#BA��@lڞ1'a����u�)���q��G#Tq����/MvKq  D�4 $%M5:�r� �#�y�4س㣟����$���'m���slI�4�&x��O.j ���@��!�_�2���`
U A)� �� �@˗1D�D��o��. B�pP�]3X
$��o/�A��l��+-%F#|�Rʗ�2��AS󈇷����A/S�<qB��عٴ�\�9~�qÓJ 'v�%��i��H���O?�$VV�őf�K�����l!��G�-�ΐQ�NJ�)�0w�:	���̫tX�| e���0=� p(#oT!نyx��>d�Εz��'��]z��<����臰e�f�ks�J�3�~�	�.Hc�<�ÂO7T����((zP% ���Z�'mڹ��b�6W���E�dj�
P��C#F�"��#G��-�yb��_"X��.^�&k��¦h��M����i2���K>E�ܴl�zh&Տq��p ]�<���ȓv��jB�$~vBE0�S�ZL�@�'���5� S؞@P � �z��򤝗K�A�e4D��ٰ��9�6 �o["f蚕��5D��1[e��C�G3?�@m��0D�X�-J'�>,+Vl�6�*%Z�*2D�$�� @��W��Fa1iԇ6ړZKj8� @Ю���CC��<rw��3g�ۜb�: �"O���"	ئ2� �sv ]=B�|A��	,��yc��:e�듟h���K�B���v G�����^*�!��3�uٱ��4�,5Bѥo�v�A?,>����F[$EN�9��J�f$�s��	:��\"�D�4�х�	�/�(iE���F~<1��l˭{���G��'u(���B�iz�Ԇ�T1@%� @[o:�Y�f�Hl��=Is�Q�<ވ����TlÉ�T���)�L�ٱ�.e�&�� N��yB��!u��q!Cͽ�DPP"Ɣ%2-2ǌܔ=��Ca�OfXa��Y�|q�F�7�zq!eF,uM����3D�@Y$�8M�h�7gſMA����l�D72i�#D$|N̻�d��<���	!�F �'��V�L�2�X_������2H��bv�c!�e!���s6p5I0H�i�D���F�V���h.��f���@�G�H`f��R�B<pׄ1�r�B=sߐ��f	�Sv<�$F6��;]��a�j�z�s���i�b�>��n�+�������P�e���1� ��H���UOR����X&je$��o�<�ċ&�gy�G�Q'��D�Byz�z ���yb� L�`����j��S�z���2��4����a�0Ÿ�HN�,�`y�KQ

4���(m�v���B˿pz��[i�X �	�}�䬱S�3��'���	���C`n	�t��� �L
7$^x�Y��)Hnx��	�&0(�S4�{�6�)�@��fPF�x�.��M��xҠ����Jݖz�2#~R�)I�(M�\��dM 1<v��Dx�'(>9��Eȝ.��}.u��AK�Ά(P
�|��F3|�εIcΞ5&�n�'�.�G�,O�)��\T#B�W	Ѣ.���Q�3O��y���w�9�J�"~�Bf�ekֽ�PȀ)/�B�g
ʦ�!�̍;��I2�49Ó�)a�M�6b�,}l>�R�><�V-�<Z��b�8�vmE<[��	�~��qy��5���[ �«9G����U�"0L_�y�PIj�Ň	"�):�h�1E�YI`J�d(<A�kP=Q�uaS�E:@.<�#1b�|�'�U�C�]7��^��@	�80�F�iRÊ*rF��f"Oz�� � ��hؗ��*B]�1�uZ� �C�EqO�>��$ƛ ����X{v��d3D�,��
'bT:���Xl�R�Y�3D���ë�S�61Y�g�+@�8�0D�� R�w\f���ۗ�D\{V�,D�4a O�31r����-b�^9�g9D�h�ӅK,o�R��^�Zx�B`8D�Dr4,�%60�_�3-7�*D�l:W�;;4��i��\�u������5D���$�Uv���.I>
��)1D�T"���*7��h�I�vؑ��.D������$#B
�p���;��¥� D��Y݃Kzn�@IјF��}#v-*D�P�f��4��A�w�O�l��1���6D�RX�SN`��`��2�#2D�dq�a���AR�I�2��H��0D�PЅ�E�:8pC�$=�i�( D��֧Z�1MdPɐ�5\�|P��d?D������ʽQ�ĕ_�FH;
;D���I^!w���b��QV�9 �;D�H�'�Ð6��q+Y�z� �"7D�$�犼l~iq�V�nr(��"'D�� �j��çLZ:�DjUm�\�d"OH���M�@DIEV��$��"O��"b�l�X#�h
�gk`�Ґ"Olh+F���;����C�Ms�@1�"O��(�
�[�ex�/K�ph���"OdI����	Yg���qH�c��዁"O�M�e�O;`�Vm���19�8S�"O�\ڃ�G� ��Q�f*�w/��i"O��TM�:=��"�	L�2j�cW"O^�҅���J3��đQ��P�1"Oj0c7�[l�X�0�Ȝ?{"�Ъp"Odq�ԧs�8x�&K�\	�H�u"O\S�/P�7m4LACE�*��]b"O�8���5k�(�
ㄝ!@���"O�y��N�W��$��T�uB���"O�����S�����nJ37
,M�'"O��`t+��uܴ#vmn�vh��"O���g# �x�4tѷG�%N�V�S�"O�Bǀ|G����GQ/XrVݸ�"O���	�F�����C�'tB=��"O �s	R/0p1�Vi��ykK�1:�>�z��A��n����w�)���+���e��]��R&^� ��8,��\�΂H�)ڧ��Md&ӫK6����38�po�Ag0�ҡ�|��i٥U��5s�D�$_�@���,$��YR��s≫YI<�����<�íW3�����fy�Z�%�4��ˍ��xםK�>��Qx�F�rW���NWjy�L�4�Y�+\�ݨ��7m�?+�1f.	m��y�G����c砕�FAN�rק���DW�͸N��J�*�6�>Y�r�q$ވC��)t� l[览��^w�t��tdĦ@�pٓ䃞Z�<�Cdj��IFDhT(׽I?���O��"}��O��x�)ݐ	��8��U�P?��T�G��	��/[/\����H���O*H��e\%�P�1�١I[H�2���l_�!X�Auy��0�ɇ<g�$�S	$��P��?�,�X��	��1�`�d>��a��ʦ��"!��0|�eE'H��Ր�M�S�ʩ*◢\W�u���ͦ��a��U�@�Zç��5++�#!��7�D�j%�b ��O�9�`�y�J�F��a���iGv����;Ъ�A�ޔ/RX;tD�+K�8�k���D�I�r�O�>�ӵ[p�e��7U�Ȩ�ψ�&rJY�G�X<|[��y�a2�4��<��-�ƁړEW~���@�N)��8�M\(=Xvq���'�����K*
2��j�[�HB���'�Ԥ����.��\�RnW�A����	�'ĔY� !�@�΀HR"�:2��S�'S�J2�ܴG� �,��"�|��'Yl$������m���Z�4V���'�r0�WDӬAxD�KB[�L��'���g��&��)��$�!�.�C�'�6a懙�(t( ьB�'@ܻ�'�"8`3�6��3�n�b���h�'��ؠ�k^*v�K'�,[L\���'�d��gW	Ԓ�8��Z�Op�� �'C������P�zЙť\�EP4A��'u�m��$�#NRjp"�N�A+�D�'�����\�i����ģ=�
 "�'z�K�X	��}��#�m(��h�'[XP��l�'m^���s���aX����'*��Go�Q�3�܇Z�|���'
��	c�!u�ԭh��E���'Q�P��Ё&(ֈ�a�Mcb���'��:6o�"$F5�#�Tw��DX	�'ix`A���Ё�3@�vܢ|��'<���o�2J��Tr#�،\<$��'�t�hQ-F�$#H$�b�[:���'�x찃G��X�8�'a��
��':f��E��1�$1&e�>�rt��'��|���Ιu��ɫ5I��#����'�p���Hn\8��٥,;\x��� ��o�B�؄ 7�l>�-V"O�QQ����h��e����I=�|�"O�틀L��q�P��1��1#D}��"Ov|�EG�>�di��
p' ��"O�,q��PV��,��hE�$��"O���I%{E* &! p	���f"O>-��jV�u�́Pf�˯�Di�"OJ�p#�m*��¦%p򞉚�"O�y�S��P�x�K��1�ʉ��"O.�B�� {�AC�F:�ءRc"O!aa�2�6U��lYe�R%bu"O�p%�9�p�Kí�5��|H�"O4�h��κU]d�;�l���b�#"O�MY��K�&��u�^���ܺ1"O2	gg�,Ю]J�K�c� Ur�"O��$��< ��A���t��	�'W^�ӰJ��q��5�&��q#���'�,�3�Ё_6^��拎�8e&ٹ	�'ް��M��vb,ͰE�E;)`ب!�'�ЕZ7��M�th��(
.m �'��I�2�ͭ�y�C52x�`�	�'�~��0?3�8��&��\�Aj�'=vt+��*O�L���ߌf*֤i�'*�t a,ظa�
Pp�oZM�Y!�'��!��K�h�~P�4���>�89�'�E�g
�VY�	c���#|eD���'�v��foE#"�D�����
9:D#�'�R� E̗�y�9IѠ��f٨
�'�,��s���c��У��|�[�'�F�k1�I1f�B���"յ��${	�'���(Bۃt���j�A��e�,���'�E�dm֖���Ç�enB�`�'�`���$�	_�iu���y���4:u�)	p���o����ʂ�y�D�D�� c���{����d���y�F/Q~ e;����k���/H�yB�E i���	��I\�^E[Dɖ�y�/�}T�t*���k���Z��y`�*&$�]�d�˧�R� r�͝�yr*	�)��hC-&a<�9�����y�ŋ�nvH���/����j�"Ƃ�y��E�I ��f�*~0�3�Y2�ybKT`S�᷍S�C$�m9��7�y�	G�pp� ��2sSt��dW*�y�,���x2��e�Π�WiĀ�y2��{H�#��0�6�����'h��sk��%��!���KΨe��'�\� ᎑=2}LARc�I�Eę��'��ӱ��+yx8T"͜E�^��	�'?�E)0�05�̸��\�:����'K��8k�Y�P�_�����'�� 3F �4E��"�[W@���'_
!i!�>f���>�����'��� �Y�&��`�nP�8���S�'��'H�q���~��,8	�'�>I���a�a �ۘ}(�l��'�����L�46!�!�	��@M����'�,�!`�'^��m�&זk{�`��'�d�0c�*����6��c��s�''� �@J�**&Y�$�M<a��Mi�'��0P*��W�(�	#��#����'��}bD䥬�-vY��NV�<����K�@�"�D 
�Z�x�(�|�<10��"m�h8R��X
?���#Z|�<� H}!��"_@�� ����� "O`|���
Dm!!\��<��
�'���`���;#b=P�mʴ	<��'�������1Trf\�"(3	˖�Q
�'7"�#�j���xYd�.rXP�y�'���[��*O���^�{$���'��|3��C$_��a�ėfdT��'Ɔ,0��EP���`G4Ű���'��I�6oMg>���+�>�e!�'k��P�V�I�zt��K�
���
�'`����)Bp�)Z��xH6"O�(���f�80`�(Y�~
�"OB�hF��A����X>H�Рw"O���N$����$n�:j�X�f"Oj��$d5NiN���-M4aox�(�"O�V��~Ta��, �d��&"O����)�p��4�*v}�9"O��D��U���	$MK�_c~�+�"Od<��l��ܲ�I϶t#,�"O*��B�BU������R	�8�"O蔂��Q��h�SE��9��r@"OnM��ۖx/*XK�d��~W�0�"Oġ;7g��'�pD�tM��X I5"Ot裄'*��K��ϯ;L�S"O��1����̋���K�(`��"On��pD�H�������!?�����"O�a�"�S�D��O�A�D"O�h���(Z�}���h��s"O&%�#� yP&���Ƿ,����v"OB	q��h��`:'����0�"O@�ʀ�_
_�� �AKȩ,t�a%"O@�B%eӽdԐ<�DI��Et
��B"O�9��<�Ȥ��&�:wτi/!��N�A�<�i�CT!RN�Y��-_�!��B&[,A�t��N["���[�s�!�D�;	 �rc��Dƙ!�A�!��ԋ[����i�=f�.uX4�V�7!��<zrc��J,"A�>�!򄒭s�����k�DhE&��	t!�I�ODj�*�9fތ`{�c7W[!�Ĝ:z5���q	��+��D��lޖtE!�DZ�E��,k��خ��$�A,E �Py�L�+����'�
�Gfv���@��yr�ޚ����/W�9Q��ӕ�y���L�N��D�f��F���y�/ݱ5�j ��b��,,m3e�^�y�+�k�����*
Ai��O'�yr�$��9)� �������)���yB���v:~�r@u�I��.��y2猢5Lz��(�;U��B��\�y�л,h����G�}Ir4��K��yb�El7ȅ�����kvb�s�n��yR��g���W�H?A�%�U� �y�F\�<���nҕ	��)�,���yB��.x;�4��nT�8����sS4�y���7WN�J�F@/2	�4h�)s�!�>d�t,�Q��k�� ���.?!�d�.Z��=��h;43P�IU�
=!��A�$L	���8CD���6'��	8!���pu�}��(��gB��S���N�!�$O�.�p�x���U��!�/_��!�$(J^\,C��0ۼ|���0qO!��5Ƥ�A#K%]�t�:ը�-!�d�.}ڵG��+%����%�9A!�� �4�3�B@��]�򃁝X�-J'"O�-S��=_Ж�A�̈́�k���o0D�p�G���P�wY�m�<��Wi;D�XIQGO�U���jg`�L
va�V-D��r�ᜌL0� A!��:3�d骑m,D�pb�b�T`�رQJK3u29�,D�H��	S�(�4���!��U�hɐq�*D�PcqI��(d���|�T��Q4D��z�ɐ/;	$�Yt��#qDx�X6F0D���&���1HsC
94*p2��/D��C���M@��zr���: � �+D�����iڔ��v)Њz4�q�&O,D�4H��P�2��rGDJ�x��)D����MK>6��	�g�;r�ڑ���2D��0mS�|�3����nܔ���/D�@��H�NU���.9�q��g;D���C��zP�V�Ԟ@�*l�;D�L��̂\UdىbaN. �5(Q#<D�4x�j�)���b�:z�ِ�l;D�$��؈H �d+�`�lՂ��cC:D�|#Ƃ[f���̛�B�U-;D�<(��G=bz�Q��'r�B�*�:D�����6 ���0�/�s��Ѱc,D�t#W���](\��dV�,��[�$>D�����S0:�,}�� �;��ԛ�0D���e,�9 Z&�XwEB�)�t�V�.D�#Gt>��P�]�l�a�/D��Xb���gu� �寜;"�(��."D�0�'��8g>��u@5P���I��>D���)N��#�)#����3�'D�p)@MQ%�RĨ��"j�$qTF#D�P�qEҴGj*��k��o��ś�J D����gI�v�:��5��+����A4D�x���--�:Qkf3a��@��1D�ȸS��*VÌu���»<s~����;D�\q���S��P��tv")0��8D�4��J7>u���	�be
ţ�8D�x���w�u@�mJ�9���7D�D�g�W!xUh����|��9�Ĝi�<��*(����L+	a&Ă���\�<Y�'�:έ`�ͤZ��tZ�#�X�<��L:��ň���$�Y���S�<����0(h�H�E�1��bU�<�K��.����OS�Fh��R�<���,E�XQ��ǈ�p���pI�f�<9�H	C��e��0�BJ�Id�<y�H÷v��	iƋ��I k�]�<��և&�Q`q�Q�*�:�hD��t�<Q��až���k��x`aڱ�Dl�<i�gZ�s�逡���m�4�!���h�<17�Q   �P   �	  �    �  �&  q.  �4  �:  NA  �G  �M  ,T  nZ  �`  �f  <m  �s  �y  ��   `� u�	����Zv)C�'ll\�0Kz+⟈mڄc� 特m`�DB�6%p� �f�q�䐻"�m�|Mi+��.�c`e�	��IuJ܅b�"I�;0�4���'Y8��J��}��1c��)U����	��l%ʡ�bC� b�Ԛ�@�����B&� 9� ���X`�-��H���9���=vr�,��$�3b��4�WEXB�b5���1���G��z�*�4yir���?A��?A�⌽�g�X���`�r)X�������?��й0��F[�(�I)es2���O���؊\����6&���� T(�����O�ʓ����O���'	���O����tI���R�~��AY�8�O�牐�>�+�&�)������۴0�(��y��,���I<Y�D���ⓤ9>i�1ӑe��D������I���������q��?�P�wB���Q� �$/��5R��'~�6O��m��4כ��'=�6�	�y�޴`����'��3�
��K���{#��<���*�� �G�?}� �Ϊ'�0�W���LF�IX0�����@��m-m}[��i��6��1����u�?���lY�Ik^��5�<"�J�A��;:Ȕ7mP�K�V�i@DN�Y6��PA�,�D�tk>E�mn��MG�i���Y���` �="�5�j����B �ŷ!��7���ec�4v� ˃G�)�j��!ǔ(���@�֏�V�K� AO��Y�*M
g@x��pB��\��	�´i#^7͎Цu��\�Q�qR�,� zR����G(3~M"��ڵ��p���_|�,�I=^5��u	�"s��31��
d<|���U��sA6y��N�i����9=�6][U����2��'���'	���O����K s�I��'xD@�P �-nY�T��N��]�R�:Q"O�mA"�\�VƁ!�Ə�7��eB�"O����96��3R��-��%��"O���#ȁ1�И�F)��D��S"O��Jq΁�.?�	�R�7/��,	A"Of���Aif��Aj���j!;F��fU��~Z���<�n-�4i��	��y�5��c�<!v�@�U��y���G�]t�Ѣ�v�<�f�3Y4��*ʢK�H�!ʞt�<I�͝�3Ft(��͠q|�02�I|�<g"A�������ic�c�t�<	�mS�f�(�n�>�h�AR�����3�S�O��lٱG�;C"�,�B�:.�ʧ"O���a�ލ+�D*4��:�F��q"O(�#�>�:��R�� ���6"O0|�D�K�%���*�M&��"O�峕�O?CMh4�LZO_��z"O�ep'��8j�XaP4+�.2T��X�<�r�.�O(�LN �0�"A�C�(��"O&	���Rvސ�AaJ�M��%�V"Op8��K�3s��
0��[�Lpu"O����MD�ufp��Å0����4"OB�a�m�d�x��з��G��<y��X�!��������J�x�2O
$��3#A�O�ʓ�?����t��$0�npʂM+s��!C ���2㟿e�X��B�6�t�)��I�F�J:c�M=���� :B�rL�%�z�:e"��C,!s�,�z/�� T�ɏ@�F���O�4oZϟ@K2�žM`�V;dI�Y�3GSy"�'��	S�OO�Ɣ;� �S0	�K.Y; #��1!�$e�����.\����G*s� `P�f�Ox�D
ߦMr���ß���sy���y�2O�T 􎐁CJ���Ba�>�XQ��R�ϳ>qO>�ف� �3ܑ�&�^�K��i)��;?1*Ƨn���"|R�O�F����N�9�H@�ľ����q�j�D�O�c>��N'bhR�Z�o�J<�r$4���O^�����j�
tV�na
3���a�џ�Q���L�WMJ,{Şb��c���$2K(S�O���	k�,@@Y�~ni�%�Ҩ";<B�)M�Х+0��\�>��"��:-�B�I,}c��zu"��c��|`V�P��C�I�=��d�h^�+J�]��I!�C�	��lE�$�"V���#���
��C�	����0�˟.I�Z�ASKT(��KeJ}�Ć�d����P��*O&6�8׍v�p7�?����	<kD��"�[;����W�c��C��=
kN=xw�=T$*�j2�Y;s%\��Ӣ�O�̇�I	|%P�8�@
02��M�r'];��Ǳ*5��h��'eI��a�h�vr�'�`6-1�D�=o�`�$?�a#A�B���z���o¤�Q���OV��?���?���>׆$�'�%^��s!��� ����ۖ4���艟rb��*s�4�G8�l9��O�^b50��1eڽ�Tgۢ �8��0��	f��1.����Ox���'�򚟘�� �Ca(�!��7	rte��A%�d�Oz����T���A֫M1�89��+]2�O�O��(�Ȏ}��S�B�_������'��	$O��2ڴ�?�����iI4��Dд2O4�
���(_�0RR?���D�O\��c��Sb�z����(�T>E�Ow�(�`�f��s�k��+�\�X�OaRT�Lw�-r�Î֨��tô�F�v�t����2 L����O��lک�H���)�7<��ѳah�"X�r#���XB�ɖ$1��X"h��("Mh��[=?�N�?1��ӆ!�B%'��q�Hd��E~��8lZ���'��D�a�X�$�O��$�<	�����	���RV*Y�������8.:���\5T�N�(���)BS�	8�䜁�*4:AF�2i%~��0j���	 |�� i]�!�1��ORP1-�4_N�a���U���C�'k�6��O 0�*�O c>��?9�%Q�+� �	� X&xC�j����d0�S�O)X�V��>o �b�d]?���I.O��m��M�I>�O��	=vp	��K�d:Jx ���}�z�*L��M����?9���|2�O�B�pE��f�% ��Hb�ٽM��]����Vm�ق��N�џ�\c	J3�$Ul����J��!�X��0�F�jm��s���iږ����%5s��Gy"'�u�+��
F�d�I���0����?�b�i��R�@�	Qy��?��TI���V9`��Y��*��6�OJ��"��7<�	1��	�(/���'�6��OUm�ҟ��|�	�LF�H�v����d�B<��Xj�J׏� I�ȓ�T]��n���GC�^���䊵� ��9��=;�F�"p�ȓt��gC+7��� �[�Qoj��ȓ~�^%��(�,(��S5PB���o��P*S)��Hf�
!�XR�F{�'D�̨��9��^ }Ŝ��A*��wR���"O�ܛ���O²`��7m4��c"Oȡ�r2-lI#�oÎ+���R "O>$���B��0q��Z�`�� :"O�T�0`�Q?�=�Fni�X��"O�Ճ�i3L����-�>��d���'a��8���7$� �#CҬJ�R�8&`F�n&���Exybe+I4%���u����o>~,�B�͇~onA����P�4��8�BL+e)�1 �UY`��� ��ȓ$^p@{�;w;΅`������ȓK�^�A�S(M)0p�ە9�n9�'^�X;�)%I�de��8�$�7g_�-��A6�Y�3H�	8T�zj�
 �Ą�`�	(���:+L�" �!�D��ȓb�ڶ@�p�-Ąe4:���c�R@#rG�.��сD�ԥd�Ņ�	5��	4��Ȁ�@�Rs�� �U?�B�	8"<R��3\_�1�6�Wt��B�I	P|��VI�C�8����U�TB�B�I&�<��%o���G���a�nB��0JJ�$8�"	(�[�O�2x �B�3%"�s�����ѵ&]ZȞ�=��}�O�:ܸ��j�&�Xs��=>&�B�'r���B��J_4E3���0�&;�'�
�����p���pKԺ ����'� ���ΰs{�e��l�;i~��'14�X�+��g��C@�-��c
�'��)y�$�m�(�C�R㖝��X�||Fx���I/\��,�Aj��5�u�U�8�C�I�\�Xb��ω(�^5Ps�S�J[�C�	Pl�I�튦a�Hkmѯ}�&B�	4>�`�1v`چ/��D�P�mPdC�IjwvM۴�ʈ�&Q����&C�j�*��5N57g�{"LY n6˓R+"a�����(c�*K�*�"��C�)� ��ZĮ	�&4S�n�*4���@"O�9Z���24ҵ@$��*+�P�0"O"0kA�&?74�Kc��.t��"OP�� a5^�[��H�]Ӗ����',hP�'j�d�s��%^L��u+��4��'�hr4EY<E� Eo�bO��3�'�H��I�l#�'�^A~���'�FpE��7�|��D!#?���'8�U�ax��U�cF?��T��'����C��am��2��Q�v>����d��Q?�h�����(���L��aZ�!.D���d!��U{��sd�L�fy��K�9D��y�����t�4��"6��1cS%6D���e@�#"�U*�HM�6�~���6D��B��!�heHV"�a�
YR��'D�a�L�_�& �flG;-1�D�P��Oz-��)�'!L(��_<F��)6`�',ҖDZ�'���DրE$�"�D��:�a�'��|�P���_��,He([�<�2�[=|%�DR�e*��k��TW�<���d�]��f��ea�T�<�T�Y"8�
U�e׶O�\5x���Ry��+�p>1 -C���ʆ�ʵ��)f]N�<��+���D�χj��i�2�DH�<��اs��12EoT!,q�3��G�<)�e�,t�j�m��aB���&X�<�5�A	/���:��8AU6��⪉Wx�H`E��8��_�6�Z#\?��;A�4D��	q��$��)'��FƆ��e3D��c%�8K�Ƚ�g��,�z�"1D���v��U����C
';Uh4�� 0D���D���1�l���Ʈt�*p�Ec D����.	-gNb��P�)��SEG*ړVK�@D�$/�F��4w
�}���G���y���;>��a#�W	n�s����yr� �Fd)�R�/Pت�j6 I0�y��P�v� 
���O��e����yB�Д6��p n4L��1["�P�y�� b��q4-E�/�xҪ���?��F�h�����Ո�π20 �o�@���"�g%D�`�ƥ�� ��r�mK�F��o$D���*Q�PR���$��MJ@�J3�"D�(
��##t0�kG*�B��>D�����Do6��7�@�?jr(�A<D� ��+ʸ	��7��d���<���C8��A��ݍC(� Z'�� aB�\"�(8D�$X �M\C��Q�̡U��SrG"D� ��K4�R\�sb��{ي0A%�!D��z���n����
l�p�>D��C�!��erz}���_�B���R��:�O$-� �O� RF%���>��0.�9;v
(�#"O������A���P��a�s�"OP��d�_8J��d"�E k��K�"O����!O�/Lxsu��t���`�"O|D��%R
)pDE�$�
lO��	`"O�A�� H�m���F֌6�ځ21�	�o��~��F�I�(M@�2_�LҒ��B�<Q������0���^��� ���v�<�p��>e@ܨ�B�� :�*]�ȓ|0�y+D��~���4H��n���>	�Z$�+{�t�X���
|$�ȓ.`>�gb� � �R*Ɖ3�9�Ʌ٘#<E��N�1��lPj��r�$q�S�	�!�$\,E�ʱ�d&�����!T�
�!�� ��)��!<Bp⇭��-�>�y�"O.���cǚ2>e��͉�cw@��"O�hQ�G?+!���E�*`�S6"OVm+���6Ծ�3��"�yQ��  '�O�)��Mê2~<��E���M�"O�͑WG�d���u�I�a��9��"O����V�M8M�D�4/�@��"O�]13(�)$���AE	H,2���"O6�@a�"y�biI�N��Щ��'�.T�'~�<��U���{�e�-u�\�y�'f�mz5咽O�~D�fH�0��T��'3�m�S䖰W+��*�.!�&�s�'�t!�@%�z�ąkENCJ�
�';~� bɇ(+���ڙ����
�'Ǣ���gslr�˴'N�ڪ�+��DW�Q?�#�,ȋEg&�2�:yq k(D�|T��q���b����{	*D�$�F�(I�y*G ��:~�(b�+D�LZ���#�"t��E �)Lp)��H*D���dI�l�lE��\(W��8*�"+D� �ٝ{���4�A6�Y���Of F�)�'f^��q¢]>n�j��s�RU�����'c�mK��[���#�M�TD�x�'����'U�Y|E�@zkt8��'��3��Qp��07�P(h4u��'�.4�R��J��C+X%xdB���'�L,yk x�8-�d
e�l+O�C�'�h�����13�}��Aèl�#
�'⁓D�G�H.�� $nzǮ<�	�'�su�1Y����y���	�'@���T�O!P��52�]�v�\Hx�'�j�%���%��!�R�&eff})�������Aք�=���s��{���ȓc��A����3��`{Q��!���ȓ&c�Yk0 ��~B0��Wc��,@�ȓ[?��b	*Mو��c��SU@���cm���IB%��{`c�\T&q�ȓp��ㄭԃ^�@u{�"K?=��mD{B������8tI[�P�jy���^��"�rE"O�Xs7�[6&�i���'ͺxK"O�L��`��NÚ���P�j�"Oa�tm¾$��Ac��A{G���"O<��-�F�D̊�&ۜ��ɛf"O4P@#�$�UI��V���e���'�Dݻ���@CX���m_�� sA"/�B�ȓN0��+��J��8� M���Մ�$��r� F6T(t��,9
q��fۘ���ԈCm��HO�x�@�ȓsLLр�kW�$�Ƹ� W$?�n��ȓ�h��OY�U(�=Y�/�[��ї'�\S�I��	V�?f1ir�� ʡ��	#(�S�V)H=�1�d�^��܅ȓx�x(BC�CY Vjb��a�A��m���#��>E��4qvO٦El�Ɇ�I�:,��H@�Bu�-�s@]�k�����h:��*Yx�!CS!28}R�M �C�I Y;��H��͹K5��!E 9
�C��0l���g�.�n�PsF,	�vC䉞rD<1�j�2T�Ҵ!�&6B�ɡ	e�m�VIR=�:ܲp�K�C䉪y���於��P�ǐ�_)�H���0�z$���;
����rb�D�ȓ~�"h�"¿?�8( 'řg���ȓd���� !#y�4m�� L+�@���S�? ��R���M����FBWY����"O*\���A�p)��^��L�q"O,<�W-P�w_
m����t�2�$�'*������S5k����FR8����%(s�8�ȓxo@���_�3�H���i��B��Q�ȓY��:P�T	Et�[Wk�� ��ȓ<	�IS���<�����r�P��ȓ?�� �e��]��,�g M�!2N���9`iy�͜	�6�i�C�76h,�'�ڹ �g��E`c�!&��y�g����5�ȓ>��=����/5�TŘ���m�2��ȓr09� ����X�Ɗ�3�\ȅ�%�\5��D�-'�:!�l��ȓ]=�@P���xJF�[�N�?2���I�M��ɹ_ܦ9PV�j~�5�vHɖBwB��* ,SN�k~��e��/C#B䉦a�by�Ff�C�Iس��')��C�ɤ;�u���N=���s�� �C�	�z=ҙA�˗<Z|j��F,�6chC�ɩM����D%�16V)���9A���=a���S�O�`Ʉ)34���6�( ��'�H㗩ֳf@<�h4�
|�L�
�'n�5���T�'��l�@�^$yT�p�'TT�a̙6A�[Ã�;k+�� �'^rQ��h�lHZ ��a����	�'����HT����R��L�K�x���#v�Dx��	$5'4̹!��
*�`p�C�U8B�	r��A�
X&��]�+,,\
B��M���ޑj��=�Ph@>P��B�	
}�2	��{g����C
63ĪB�Ɂs�vL�g��,2��v�y�B�I�8��|B���2E�T�̒xc>��=1H���b�J?9H�x�w��06�CqN%%Z6<a��	Uy��'���'DN�ӣj�����o�9Ai�Qb󟮝K2H ?p���d(D!Z�t����!D=Ե��^-r��I׭\7cd��r�C�� �&mE�H�]&�����-T�2����I�f���O�b>I�����.^0D��΍�>5�xKSξ<��wu�aҏ�
aE�LCc�}�j���	����ѩe�H=���jP�5���W	9���!|�^E��ҟ���d����Z��'�j�R��C4���G!Q6����'E<j���P��R7�DO���T>��|b�N�md:]8�L� svJ��2���<Q� �D��d��߸�Z��I�>q\��A��h!1�X2 M�d;!R�'��)�	:?A!ˈ�!�z�D��:	Z�����H�<��FL�JI$�*Q�	 �e�P�B�'��"7K^�!��+PB_9���䥎��?)���?�3hÔ#?�r��?)���?�����d�%�����B��rp�_K��������Ò41�)�4�<Fx����Y/����< B����d����':z��8N��i͟��DK�%(d�����I�`��)5?Q!X������?ٜOp�Ԩ���,w��u�5	[:@=�U��'�f����2A�i�NO):^Ȝ��0A���Sٟh�'a��@�鈶2�2����A%*-@1&�9
�L�(��'�b�'s��h�������'q��Pa��;\��rM�^]���B��%)P4�ǅ��X�F�'�h� ����=y#��q\z�@�y��V쟁�� cs�*,O��+�'oy��/� � E����]��@�P�'����3ڧO=
���	�;��ZD&͚K��	�'��X����x²uZ� �!HD�I,O��)�Ir�:�~䥟�p7H�	j���s'��L_>��@"O��`�$&��Ex��T�bkz�Iu"O�SPo��8�<0��F�=}6nYX�"OTX�dI�:g����8º���"Ov�҂L����+�dĪ�۳$"O�hr��/~T���.f��t���D�+q���O6z�:�ٯ[&]���V�E�\9b�''$H)����a`ˍ�6�b\�	�'�P$p c5\�J����6qd=`	��� ��5Ђb��Qx��PY�EV"OЬ�ѭ�$}��5�2�.{�6�!4"O����)j�0u�!@A�28\P�@�΢�O��}�A�f��D�I�Jȶ�C���ZF��>��kB `�|5+@W�Z؂8��	��5�&���A<Х�gf΢44t��(��5�wL��MC���#�(u��ńȓR-��b�'@ a�;��>)�h��ȓXX�����V7q��EM�W��<�I2Q@���d
�E�R��/'T2P�lZ!��9v�䃵L� N������%�!���~���K�w�ʤ+_�!�$97vbPKa�� �8�	�m�!�K��q�����%2A��џ,hf���M��?�O�� *�[�@�$��ӏY�]��K��^�H�Q���?���\�B�˦	Ir�d���ITY�6=�2���L�O�Ș#W�ޗ3������7a]v�I�+� c�"L�1aU����!��127���4�b�LK%x��##��O�#|���Վq���CS�ӔAI��c�\�<�� ��M�EM�JZZx���.OZ��=XB8�9'CE
��D�#V���Οؖ'�O���.�P�0���rT�Y"�Q�Pׄ��:�|%��C�-Y�,yx#��[Rn��?�4�ēA�8b>A���Ԏ.�hdq�6z�y��(?��O��q#�>��y2DJ�@��{4E�41��Z��ֻ�65[㓟p�I���.}Rk/���ck�8hUƆ�n��t�!-^�C�ti�I��a�'��>�	KG0�C"�$dߔ$�ƀ̋aHx�dD>}�"}�`	��I�����pE�-3сv\��s��A'Ę���I2�N�*R���F���cb���6�N��놫�?Q�(@��v�$ɷr��V���.��B}ތ����)�$����)��$��c��sQ�?����?A^HQp�2Ad�x0��{��I�/�ҧ�9OhT���*�&�5H^�ʶ��`�T�⮃�to"T�'*�mJ�O��x��)�r��cR*D�;1��AIɸy��@C?��MN~ʟ�dSq��$@+V�9!ꈁ}�i��8N�2�_؟x�uD�<u2�)���A�R>��2D�.D��)ai��q]��h�
(��lm��4$��٪���O��4E���x��E V��k��^�Jh�&T��$�tG{��	{���g�H(�C�0P�d���"O�%�P#�\�d��SD����
E"O�#��JV�-�d�3{f-a�"O��k�#�/���"ʆ~eP���"On9�W�M����!/�5\v�4"O4A*I-+n��b���"O���៫(�h�3-:c���(�"O�L�d�9Ȁ�5+K�6"O\Б���<k�0���+ި���0s"O4�	�Y.Yt��kC��#R�0�"O^�JtM��`@ ��d͎�	�"OXh�i�>P98��ad�/\T��"O���Z�I������,{��D�dZe)«^���=�FN��<X�v!V�,��}�gꍋ	"y�QL�sͺ%"�֬k���8�C���<��*V	&��쀑=J�ٙ�K�O�J����۶_�&\
�� E���1�0I�|1���îF<�Y��J�P˷l�(�$���t�6h ��j�>i�dqQ�%�=[O�m�tc�7x��B�	X�lL{�	�<��@�K�G�hB䉍:G�H #�Fֈ���l�2�C�ɼV�
�%����9�L�Xp�C�	/M�0�AB�F�݈U:�+$-�B�;R�L���-����"��+vB�	� 	���h�1B�����x��C��qc�� �B�m'P�J��^,;ΚC�ɫTl�IQ#b�.f_��#���bC�����yPe�~ �0+g(X$�ZC�Iu���h�P7(����ɿt�B�	.7Ťd�!�ǖ������E�I?�B�I�x�Ɲ��"#A���ڱe�8{!B�)� xys�w@�����
��#"O\�z��?i��	vLQ�|�~���"O���'ď$���K�7A�:��`"O���`J%z��S��;]|�x"Ob��Q�K�y��H���7�<��""O���`bB/Q2�)BW��7�H�2"O�P�*�T|���ӮH��Ss"Oh��q�W��p�u��bD 2�"O�y�ai�4��"	�7C�}Z"O ���˒+-�ry*RF�#8��%"O8M��y��\ �ZEs"O����;O̘a�K�$5�U�"O�vH �����	��q�� S	!�F�"�Tepօ�!�&�yQ!�q�!�D�6@^)a2�ܻh�"�)��NL�!�d�F��ѱ�I�)�N�P W h�!��/�la� [�XЬE���0q�!��
t���&�lDR�b�2�!�$V�(G�pC疿u-�}�5O�}�!�d�h�ˤh� L�x8�߄�!�d�!UfV��C�^�&���)����!���*l¤��2|���h[�8�!�V�S��(7!ގES�@��gOi!�ݽr��)$�XC��ArM̞Z�!�d7D%P&�E� ���P��ս-�!�d�Jl���K�C�,��3Gو�!�<q�,أ�~�<P�fV9Uk!�D\#Z��hfA� +����μ^g!�߾J	X�AчH|�� @*[��!�$[�z���E��dj��xц�t�!�ΪU�\��&!��ze�4�ckB?�!��	T"��p�䕑:�v�jBj���!�d��d5��hM�'�q8�+^*�!�	�}�d�0���N����7��}�!�d�@2@���ڷ���D��&�!��\��H��
�J�f��	�%�!��=~F<<q�ʕjmde�I�6�!��&2���h��7&V/'q���"O�!-%�Дӵđ�c>Q�
�'��ժU�է_�� �fU7����'T�8Pe��`2�tI �)b�p��'����G�3J��Y���R��<��'�4���#�	GT!@�(��X��'���H� \9Q��ǡ��mR���'���`�Q �B�ҡ,�h2(tc�'��<�$�X3Fm�l �È0�R5��'���(F��r�NN�QV�@�	�'G�At̏/o�0���-xC��H�'(���`啪*U��PR��*#��A	�'$dɱN�"T�4PP��H-j- ���'����/7��<j�ɂ�`H*x�'v�����Ύd$����)c���'��]H�BP�@>���й`8樒
�'Y�HX���C����)X�h��'�L�����T�A��}:�I��'�)Z�	_���Q[�ɍ�|��|+�'^d��'�1_FE��Oc,d��
�'��1��Ї�x�S挐'!�
�'�$�CBDR G�PE�0h�
�d$z�'�ƥ���]���E�;m�~ػ	�'X�ܓ�k�:i'���`���;N�1��';�J5'D;k���p��.��h��'�^��Rh�3#��ʑ��,��
�'o��'ˣd��P�Q^4<�s	��� ���K�Gft|2�K���"O���a�����bg¢ ؈�"Or`9W"�5�z����>��r'"OB ��Ԑh3̨*2���T�)"O�I9f$��
��qri�+��`"O�!�(S3
�r�����T�8�Ys"O<���g��X�0�`�*�*OXH��`�\��:�g6@��P
�'Vr�fk�/=e��ҕ�?�z
�'��Xq2$V�zش2rD�=�<̺�'.p����9}���4L��.��9!�'�=@fI��yAoܘ&�ތs�'����B%��0�=4�|<��'��D��� 2�u�� (�fE��'�XU��b	����Y��B�ꈡ��'B@d�G��;JF���ĉ�j���'��Y�Fl@-��QP � ~��<��'��<�u���4@�)ҥg�h�h�'�,�sB�U0��$��g;�A�'�ju��B��BPY3ˀJ�.���'�����H;?	H5��BH�>7(h��'��u+�J�K�=F[(:��y�'0�$�LZ�`ܚ,X�X;
�'r6��L�L ��)!�S0[.�q�ʓy�xą��,���B�!������3��I�<�X���f��&i�ȓ] d@��������j�*C�ćȓ	*^�b��F�;
 ����ц�� ��I�T�%�d��MÚ����LU��հ0@�|�0��5j����N��H� �4܀l���'^�6y�ȓh����,į;^V�����\��fe�����I���G�	�3Q]�ȓ0(f��q�9,���:�냭D�"	���}c	A�E*����lH�l� ���pXe����~U�Iz`#��>�ȓH�F�`ҿ���I��׭q��ԅ����j��ѝn� S�.N#�Z�ȓM* �ЫVÜ�&Ό������gm�4���`ü%F�݄f���ȓC��ʀi�"ڠ��	Z=	�e��tڤ1��c�N��)sΚ>&��	�ȓ^m��h�0t�����>~����|�h������Y���̷GNP���:8�h�\�p�6���5r��ȓwĠx��kN�S�9�B�'x�"Q��D�Q�#�*ihuu�[�JH�ȓn���yB�VF���DL�v0��ȓ@��L��:/*���� ��E�� H%�b��4r�H�Q�1#q��ȓN�X�s�>�0a)&�FLj]��Z-�xi�\�Q�v�*Ba_�L����ȓy����>X^�j�疳>� ��*��r)�.�Yt��M�x��v��(��dݏ9:=@�=h/�a����`�uꉘo�0ĠF���q�ȓ.6Vv�7]6p��t&�A'�܄�K�B}�"L*%��SEHN�E^�Ʉ�M�\m@��2�h�&��S8΄��}m�!���"��L��G�7̴��#
���!+}��m;g�^2��ȓ?Y =÷ ��#�
\�ၙT�Z!��y�dيG��/]����_�R5x �ȓdF�ծ��r͘#kQ[�j���S�? �P�,��JEN����(\Ș0f"O2�:c�IYB(�e�q��٫Q"O�A�f�?	�B�Y�bNd�"�;P"O.X+�d�(�vDrrˈ?+��U��"O�z���<~͂ܨ� �>����"O��B��B��\�4NZ�~�V�qd"Oݚcn�X��5	b�>޾�2f"O��L�"/Ў�r�j�2����"O��``F48��BQ�W�^,�6"O ��&�ր+ D%�"���x��mP"O�y��F?q�\Հ	]�()"O��&�^ 8��m#'ϑ�Z��"O��k3+؅n�*u�EG.2��1�"O�(�k���O��1�zR�"O ����΋h�<K��m�Aq�"Oz)���)T��I+��=p<l��"O�9 ˀ+���b`i�%��"O�=IG��H�������W.Yr�"O
iQ��ÈyD�suA�RQZ�e"Of��Q-��a�(�Z�/�?k��$��"O���
�;��a�`Q�=�����"Ob�d,� b�tq�J�G|xU��"Obq���юd�$Dqīyu���"O�	�'Bۡ*�4ܻ/
 r�̊�"O��R�߷$�����o��qzن"OT��"^'HlH���Ƭm��ca"OV$� �"H`���"�_�f:�"u"O�9�6�.B�Z �eKGd-�"Oh�2����T����<;E�Xq"O�+��զ\�Υ��H�o�L��"O<�AVGq0�5���W�|b5��"OH<���#�X+dgYx8P��"O6 ��J��n�&`��[?��#�"O���o_��Q���{/�)��"O�4z ��Z���ҧ�����AC�"O�� S�=� 䂲�D2�j��"O�1�"��O6�(�bϟr�N$�7"Om���0����_� p`�S"O� p�O
Fr���U(�1Z`�x�'"O�����"R��xg� ]"���"O�p�@N�X�*-�pe�~o�Ty�"O��Q`��^rr�i!D�0fz��7"O�U�1���l%��آ��eZH<��"ONdB��ҜnojU@�W7F�L��"O��ؤ�G咐� �zͩȎ�y�Ɔ�S\ �##N@;��`h�A �y�� B"Ver�ڶfۄAJ@"��yB �%F�h��PŖe��X�K��y���E�Pԙ���,� j��
��y�H�q �ؗ.X� 0q3#���yBNθ7��H�%��`��x�U��y��� N����͙4by|���%F(�yr�(K`�}�6ȃZj��H���yBh�0�M���5T�V�P�L�6�y�M
�dnБsC�M��U۱���y�>_�D��t�@��P�ƫݙ�y�g��>}8�!ɞ5<5|�21+V���'~��Ȁ������!h�,�K>)�!
�}:d-��B>��rmd�<� ��>M�I*A��K=_�,��'�~		F�Ր7tQ�c�
;\x� ��'���l�+N�<PZ���%g��'l���$�T�IP#�gѶ��
�'\YT&�$c�T���Pv��`
�'9�Q�/��r��4 �ȣ=�<�
��� &Dq�hףdz�2�!��+ژH@�"On	&�M�-h�u!�4��,�"Ovɣ2M�1��;�g��m���B"Or��B�ڣP~��ކv�P��"O��"
�>�`�O	�vfҨ�"O � q_�3'�4��-�r��9Qw"Od�D�PF�d���앻
wLi�""O��m�m'�$�0# ^��x�"O�U��4E84�c cɐ- ��8�"O�1�1��C���Z!�ݜ@�\�q"O��ǬśX�V����9u���v"O���P�T�] \����6�:��"OP�q"+�-lf���g6��4��"O��Xd�3[�Ȝqvb�p�q�"Oм�oR�X��I���*|hx�"O~A�*�@��D�.�."��""O�u�mί����UǍ	"��c"O���2�D�K��yӰ��].D�g"OԨa6ȁ�K8����c�B�4"O*в+\�C%xqs�dǸ�""O>T�Ҍ	)ܼ���]�N_j���"O
�#���n$�9���1��X0"O����V�Wh6D�@�T�#"O�����E�`l��C�� �/!�	V�Q���7��1#�!��XC!��0+�̰��`!��b����!��_&q�Fف���uk:I�g�Z;4G!�$͕=�$��ĄnV"\QԦ�$e�!򄝺3�FDy�m�"HK*,i �V�!�$� -��V�^�eWJI[$��#�!�DZ�fƎ��-� T� 4�W�޼/!��4l�MK�E�$�b!���I�@�!�d��eh�q�5~>(��E���!�^�)����D�2V>�P��M�%�!��a�����D�x���7�!���a��,L�!ihI�n�c!��ÏE�Pt`�HвL�h��j�#v)!��d��@5L�^[���`Wc�!�$ˉW8��p����nEt5���Y`�!�D�~�ԱQ,ڰp�m@7����!���	_� v�+wOH�q��Ѧ&�!�O>�Z8k���B�)zaKF�$�!��(ꅬ�(<P-)��Ȑ�' �%��>�𼛓`V�p��h��'�\1�@U�<^U���ѳY�l@��'i��R�?8�UA M�q��'ɠ�UǘYq��HVAͭ[t���'�p�xe.S�d��x����Rj�x	�'.V�H�(�(0�i�¯C�]��'K"�A��0Y��!�bD2u��%��'�� �V��!Jޒ��4�CAV��#�'l�C�O�"��T�a��-��4�
�'���1Td^T
��c�Q� ���	�'j� �w*Н c�N���%n�}�<���jdL���J��i�͋R�<�A ̀=��!#��[�`R1���m�<9p%Ԁ���������H�e�Zu�<9B�!����6��wi��&čO�<9�/�{#Pa �Q$�wJ�<�g�E1M�`���$U�ЉF�IG�<v-3��А �P��%:Q�VC�<�(��fuR9�wF�9zD�Q���M]�<����F@0�a�@�2Y �I�C��X�<�� ��v��"#�)-%̨�LF�<� @�Pq��7D� p7��Fv�1�"O���'h
^<{0� i�t��"O8�"�"	(k?�Y ���6$�!�"O���ϐ9~�� �ַ2�^��"O����Q4 �8��Ņϸ���0"O�x0G�̹}���%��Q� ��U"O���lQ&8�F��@���t��"O$$��IK�7�,���@�NY�"O�Y�V�[6~�Se�^����k�"O �Uh(������@,F�<-�u"OU3$j��W���Ĥ�=s1P"O2}ZƆѥfGָ��O#bh��A"O@Hz�+P�p��-[�͆5W�aju"O~��f�����	G"�f�@�b"O��[�#�!L،8��2r�`a`�"O�����Jt����HŁ��4"OΈ���Wv��[�
 &��Җ"OD�sJ��%���T���dX\K"Oj��%Z�9�V�Ď^B=("O��؇���(�;�MT�kG�h"O�� ޘ+V�����C�D� x	�"O �x��9U��`Ze	3�8X�"O$s3O"Р5�4k2'�H�"Ot�:୊�O�����i����(�"OL(�2۝]������W��()�"O�͓E`��?�fL�7cܑi���j�"O�����>���85�m�"O�H�
1{�N0y#�P�*��5"Ob�S��>hO���C�p<Q�"O���PÙ0f�m
�J
9�4r�"O��k�C�%&�����/�t�ñ"O�,cv-݆�H��'EMV��AIw"O�#�)�6�&��s)�==�;�"Ol�#n�&"�z�k�h0O�Z�*�"O���6��5�L0I2�I�.�XHV"O�	��B��Q�(��3-��|�u#�"Od�z)�t�5y5#�9�`���"O�p��*�,4#1�
1z�� Z�"Ort��V�&�*��/��t�"O20��׎57�x;t�¯ij�e��"O��Ĥ��mƲ��4�	g����"Ore���+%y@8#@��;\���"O�H�-@�F���oҠj���G"O����$[R���ΜR}����"O:D%��{XD �3�S�Vξ\J"O�P��O<1M��#��2G(�(i�"O�M��� H�V�z�eG7	^�X�"O0�S�'�y+���W�
nL�b"O.̋W(�7o �#�*�,EQ~���"O� �)�n�}��#� i�X�#�"O�arGM'�����,�h���)�"O����*�8�����8f�P"OP��T ��j����a(��2���2�"O�(���]��谛��E�8�t�c"OB5�P�Z"!�^i��'�]�x���"O���5��k��,�v	�g�.4��"O8 �KBM�(��"�S%I���5"O.����M�n1"	ۑ ��$Y0"O��@sM;��<���L:$��"O�Ԙ���]�@��Cd,��"O��ˢ��
%;D���G ���:�"O����Y-'����g�-j�DM�"O��y��[:�.u��޴j�"O|9�[�f�*�srJT�"�[�"O� �`c��A& }��������C"O\��3g�3e�\([��X7Vh��j&"O�K��Rx%45��acT hv"O6e��̛(
� ÈU��"O��j�Ë�\z�`'H�m��Y�e"O51�I�4N�%�l9M��1�""ODT2�#����Ӡ=j�(4�S*O9��ʇ+�T[�FpM2�'HI;���J�t�1eŔ4���'�0\�6B:6��T�!fa�B��?DjZ]+�'�*��=	fJ�$y�`B䉾3���B�,�2anE��S�|��B�ɰ2p��W�
�M���QCаT��B��5>pj�⡯���d0G�"��B�ɺo�|2�G �@'6X�B�	�Ni���'V�.������A2ԚB��62�>� �R��P��#F.pPB�I�)I�\2�-�0�4����=J�\C�	/E<m�-�]]J�P��?k�B�I���}23��P��y���ʒ&pC�ɑD�VaM�Ll�������P� B�	�_�p1��F8�x�apmQ�z�BC�I�C��@��
�0h,nAGL�&C�I	CNMX�@�\|�p戕j�C�	�[��	IEBޯ6� ,@
W _:�B�	0k�
�gl�#!O�MT
�~��B�ɧmd��cH�?f��i��װ}֜C�	�<(8��앎c��쩓���RB�:h:+�='QV$��ՋQ{��P�'k,�c�H"`	F���O�4�̼y�'��	4$�:��H������ޒ�y�`͡[���Q�	{hp�X�B��y��A=v����ٹteĨ�uI��yB��M|�05�]Ѧ������y�M�Rw��� ��%��[�GP��ȓ-@���B(�l�8�0��g�rh��V��Թ �p�)��ȉ]ӌ��ȓd�D���\:�B�3fo�)�ȓl�v�HcIW�WvQ	U [�qr��P}dU�'��4X�zy2�I*����'�,�k��
lt%��_v�����!�h���PU���ŇU�VM��,P,Ms�W&�&������i��.���gg�duI�Ro�t� ��ȓt�KǢ�4"J:(�0��e���ȓ]]v���h��t��@�t�n���D�4L���0��Y�2��D��W�r(1��?��9�j�\Q�Ą� �@�[T(��)̰�B͝�b�fY��nB�����-U�@��OC5$H���Bې$�c(Ӗd�����
3K`m��'�"TP��^l���Z�-	l3�m��v'�#�n �VM��N�1K�,�ȓw�i3��ME�.�2�K
u?J�ȓl�.���@R�C�d�8�K�K�
Q�ȓ??H�)2��t�*��bD���,��ȓq�@B&D9��p(�L��6<Շȓ-? �{V� ^�Ni��'//�F%�����`��S�ipv�!�ì��%��ih`<Z�N�6`�r�G�V4|l����X���������FC;&��5�=�#�w���%��5X�$���f�	�-�,	����FȰ&��5qC�I�}d$T���H�.Z\|��76�$C�I'X�֔�l5#(�E�!Y�C�)� �ZQ�<��a�v��%*p!�"O8T"B��q�� :�.A�~!Vp�"O^���ɖ[>�+��R�;9(LrQ"O��S�̓�T1��t,
_+xd��"Ot���	� ܢ�%;.6��"O�0x`��"��A!a��M��52E"Oƽ"�ߴ#���a��)�����"O.Ԫ��ݵK�p9Vb�z�]�W"OfqX&ʣP�bL����WbA��"O�D�w*�%P:���O�Z,Q�"O@��� )O�mH��pF�S�"O�M�AdX��I3�P�H_���6"O0D1Ɠ�}J���g�>hOV���"O����14�XY�2�T�*6|���"O`��ꁻ{D��X Y�:#��H�"O&�I�uԬD12h�<�)A1"O��B\?,����W�I2"OEر"�12�j!��>#��V"Oq�L˹@Z�뵯��:L<A�"O:Ta�G��39j|�c B���ʈd*!�D�q|�+�$���J�.�+�!�?N~a��V��%�����!�d��5y��1AI�(M2ɓ�|~!�d�4��䧓�$��AzW�*�!�d����aXtc�x�hp��CP1!�$L�&�����^29^9ӧ�լ>1!���	-��H㮔y.���wh�%!���
d�(D0�/S)� Y��8R�!�Ѷ>�}z1��
Y�( V�)r�!�,�.�je'J�f�¼��DVV�!�DO&^h��s�O�jP�h31m^6xZ!��1L@��N�I<�x���C�x!�Ď'za�#�N�#CXP��!J!m!��/�J=�Gb��N���#��Ο]l!���|,����;�D�82jɐ@l!�d,�ݩ[!"� d�U7H�|���'wB��*�ޕ��A�8ʥ�'C(0�!��c���#��4��(��'�~X��zL���L#.rpy�'-xxr�2e��A(�o'\�F|�
�'�P@�#�̂q�JDi�)	d"O 1�ˑ�v�J��\��
��"O���nO���a2���s	�q�"O�����_֒eA�� g$*�Xb"Oܠ�
X�c������E~���`"O a1�ڋ0F8q�e]�>d©b"O�-��
�,9���%EU;G^�)G"O �cS�*P��e��M�%�T�"O��S��f;I[c��hm���"O�<�"�Z��U��FA�pÆ�r�"O�l˷+26:Yw+O�\\f5p�"O|u��^�gN\�9�꓉wʵ�%"O:�CD��#������$Ev���e"Ot�Caڀ2>�usq�1);����"O�)E@��JC����p��8�"O08J È��pPU���R�5T"O�M:IG�b?2�:a�]�f����"O�1s���W,��U�
-�H��3"O.LP��%XC�\y�IY� �M�"O6@�g%�Y�jܨ�����D��"OdyZDe� |����/�xI:,P�"O�$�����
���Α#���X�"Oz��@��î���2V�2 �&"O�	�#� Z6"ǋ��I~|�ѓ"O� N��>'�=`Ԭ�Yz��z�"O��b�mF I����TA>~u�@95"O�`�WCW���xtIĊ���"Ol+w�ˤA4}�Gԟ]�~���"O�ꖩ~i��#Bgkq8�0�"O�Y9���H�V���P�@`
P�U"O����J�_ � X�Ꞙ2T���c"O�8�(�NZج��,̽��pu"O���,)z�.�@��X9:� A��"O�ܨQ`њ+0x)�r�[�D��exA"Ot��`N�T69���2*�"Obp"�oH @�AiCmC�h���[�"Op�h��'YW.�k�k���Q"Oz\1cM��f�V��1@�?���7"O�����|�`4��!�8�"O���D僧#��mi�/B+ֺHҒ"O��9�(�q��M�/�6I+~M!�"Op�(B$٣����Aώ��z��"Ol q6��9<tMb%o�!r&��"O��1i��$X�I�YYh��"O�p	T�\�t���&ʴ\eV���"O�OGZ=�h	��4THP��"O�7 G�b��IKw�X#<hM� "O$A����#,@�xa璯^8<p(�"O0�4��9|d|E
�"M��35"O^��Q��x)Ԧ�	����"Oܱ�!�G����rfͨm�T��!"O�I9�'�2��R%�#.���p"O���6kL�R���p*he��"O�<KaD�S3��ꄠ��m���:�"O��C#�A�ne��ؖ�$�{�"O�T�!�7r�>��/۷j���"O���S�Z�&KBE�B`P�!"OJ���G�^lX��ڹ��a��"Oz�Ca�׷�DA��q�@�g"O��UDS=�ju�F�o�"�d"OԴ�W퇤6�N|Hҍ./����"Oz����Z;[F� �q�����"OΡ"f��$� �96���&|5"O�$�eA+Q�J��B��ٲ�"OҜ��EE�m@��mJ���)HB"OP��"!�5:��M�Uk��%���"On�&�%���s��3/`lEh�"Oh�
�Ry!��JY�zD�Y S"O��I!g��B�0�	G$���� "OT��o��$���iP��[#0���"O�ɋ��?+nNTʄ�
�	1f"O��0�0/X��z�E�{�Dkf"O3E�ۅ �4ӧ�Y�%�x���"O��0����R ����.�v"O�1�fӐ|���U��L8XJ�"Oz�	�U0i�e[�İ_ї"O�!؅���lM�pA�� 2}�B"Ol�Y�M4M��Pf�1]L!#Q"O.|��K*n��`[�6"�\��"OB]PO��R�n5#��,w���"O�(	��X��p���F��5�$���"O �:��V�l�9:wkJ.h�.�8c"Otu�q�Q60{Z��#�7vrH�""OL[eO�x�2������]h8m�u"Olh1�&]$��t��L�q\b���"On-� ���� �A�K�5f�I�"O̐*�-��dp:Q��?\�@��'?�DG7Dv]bUM�R���C���%R!�� ��f�B�^��rm�?TE��"2"O��Ԁ�	U��ƍ�*o9�I��"O��!c�F��dx�+Z�����"O� ���8� �t��j�R\�t"O���i8T4�aÏ�l֚��"O%8�&h�H�
T@4��4p�"Ov(@�kG� ��Mkq�>V����V"O���V�T�XD�B��˟a����"O�pKrJ��k���(D����y���;��"��T�B�L�� ��y�6Z�Eqs��=֮�B#f\'�y�-W��]����DlQR�U��y��X�j1>�[V��4.�Qq`:�y�C��Đ,R�#��{������y�P�Ix�(�"�R���B�yN5��ʓ�M�|ָ(	Sj�y��Q:R���u���s��A�b�L��y"ғ`��x���V�W�4d�&	Ƙ�yr �� �6�:i�"O�$��ˌ�ybn�Nv�� � �K���ZuC�?�yB��*`��=�vi� G��ɨq��yRi�6F%��
�ǅ�B��L����yR�ۀ)XL*�L�A��1Y�iѩ�y2 ��(���	T1Ì�q�N��yb�+��- �Iw��8��һ�y�C�[��ɳE�Hk/\,�v��y�l?nNĺw(*^�9�RD�-�y��)Ť\�'MGD�`���^4�y�bV�Vv\h�����D���k_1�yR.��[��,�B	D�\r�T��yrf�7`G�q��`;
x&HH��I��yB��$���i3���*��������yr+���ˆ*+^�s7�P��y� �[䡓t̗���m���B��y�膮�0���J�C<v�Ӑ�_��y��?>~��GA.5;>�@��y��T*�N�(�fЧ43,iY`���y��r�Uh�!�DL)e<�y�AI!s!\ jrE�|�L[Q��/�y���\Q̘`O��AH�� ̖�y��6O�h��⭅�Mp@-�"JR��yJ�(x%�ys�J6V/H��(ҕ�yҠ�=]��)�@*�;}ݨ���E֯�y��[�$+����x��h�϶�y��>�������6#p�q�W�T��yR�ƫ+c����^�{��#��G��y����z'4�� bK�U���qL�y"`�N��RA�J\h@�Q=�y�����(���^����_�y���_�L�w��"��"��y≔�3���Q��M8��	��y2�ќ>������5j�m��#�y�#��;D����W�=X��)�9�y�MS�1���,�/�a�n���y�J[�l�f�砏?)'�MY�`���y��G�� �$ا(rV�ӥ�׊�yb���&m�$ZA�\� �Iه���y��X�ع� U6!�c���y�L�� �˂�,�u�N��y���#�\����eGlX����:�y2A��Nꓨ�d:Z�Z��@��y2�[�}��%��*�0]����eڹ�y���<-��2fnZ�Ud>Ei�����y����p�ک+&�N�xTXQ �-'�y
� ���%��	B��
#.�q{1�7"O��#a 
F��bb�'6z�x[G"O��2�Ϣ%�`��a�h~H��"O�0s��M�b@+� %"}�<�"O�X@!.U>Du���f��b�b�"O.8q�E�h&@�$ωzY6�%"O�L#���\v\��� L�T��"O�I���Ѹ=�x�*��[e@Q�a"O X秇 hd�$�&���0`�}Â"O�H��D�5"~�IB������"O�ڢ,�ms聱2�L�u���3"O��s`n�N(V�j���-j\�w"O}X��moj��D�O�Kp�"O�@r���
'mĔ+P��v=H�� "O�Uxr����٥�D}D��*r"O�d���ŻB�NM(j�h�"OƘ� d�>c�bx[�T$���'"O��(U�
<WYHDx�M�  �8W"O�3J���8`�i�y.Pp"O��Icd�k��	Pf��(T�|飥"O~��핃K�p=�Q
�&,�B�t"OV �V�Þ}J��IP�N���U"O*���\ Y���#e��y��J�"O2�9���#Va�}�I1s��"O~�(1M�*U:0�5�$�
�E"O�2���"s�R�:�j��܉(�"O��A$](Fx�T��c�k�����"O���t�@
j��
dɇ1b�Yh�"O\!`��R/J���)�.�"m����"O��T��p��1m
 ����2"O��I��B�ᶽ�lC��Ecf"O�xC-Os�fêD�4�Qˆ"OR)Q�gM��HQ:��\z~Ř�"O<���+`<^�	2�G�A� �"O�yeH����٩D��v��j "O)hdB[2�J=P$����6�JV"O�A��[-*f�@��9.� Ʌ"OZ�D�;t��\[���$�B���"O�(YuaЦ;�p�ȏ�g�zMڤ"O@���շ]]:m�R烂Q����"O��sF�g��0KF]-�ͺw"O�,����T1'�	��"O�qJRaPoc`4��΄��D��"OL�8u��]���C�	�}��\P�"O4�#b�5Y�lp�Ē�Z�t��3"O*9� c[)>0�ãM	|���"O�Mq �:e��WMK,z_� ��"O�8���	�=2&�I\�
T"�"O�9���J�7�P��AkD-P3���"OƐ�e��'O�4Q�H�?G1 �g"Ol�g��!`T�1�C\�@�'"Ox��C�*.��s'R�1�8(�"O�{Ќ٦LpB�[� ʬ��T�u"O�A�QM��hP"�-X����"O�=3`/X�m�^X����"�A�"O ������aEG�1��E�"O�0�v��d?.̉sg
�=x�X�"O�[��
�"e�&�s�(�"O�iyG'0\J�]���A"Ox��C�&nS�K6�#up���"O�����j���s���b|�x�"O���D��-[�Hh�˚�pH���"O4乢H��O{0�T��F:��"Oz`�b�	6aYP��Ӯ8�Ep�"O� �����n�x��+^�x�`"O�}���ws�m�F��+g`XM�P"O��(w�������S!*R}J�"O֌z6��'3>��k�/�7F�$a7"O�M)EI�\�j`�vDF�Iނ���"OBL���t���x�<�f$� "O*�i689[�(�!q����p"O�Y�%o\쌲5���;��1{ "O
#��K����K�i�ܕ��"O�ڄ��3�q��f�?D#�90#"O�y��'i�$@a�c[�o�5��"O.M�Я 	Jj���p"�
�*D�w"Ov���ӛ'��$�� VQ���2"O�Z��[�R�l�Q�7s�i�R"O*�Y/��̝S�8��qD"O�]20O&9�DM�uc�-R��k�"O���B�E$�H����/?�1�b"O�Q��RIBH;"�B�5�ճ�"O���+��2a� ���Գ9��ܑ�"O<�;�����s�\��F��"O��)AHǕ1r`�8�M�'Px mB�"O��J#E�][թ�-�'m���%"O��ҁع >�����kN")��"O~���j�>\�㫄�<Ne�7"OLHZ�Cy��@��GkC.��Q"O����G)4t�a��B-`�"O4�@�Qau&�@g�^���ʢ"O�d�FnȲ!G`S��B���a�"O��"�g�hHF���B�.(p�"O2X���)S��pq��Ԇ|��D��"Ol�3q�k�d�.N#U��h��"Od@���3{z<�sa�I,<�Vl�%"O:���M�x����W+Ιi�p�yS"Op�;V�P=*�<T6K�#BK���"O��a#��:e�,b���+����q"O�E�� �Gz��ҵP+���U"OP5�+ֲw��3!ݣX��m�"O�aIA���f���(�E^�:tP"O�Ts��Q�"Dv�u�&+~��a"Od�i�bɺ��ҷ���Π:"O�8*aJ�:}ڈ��n74<���0"O�a�bɌ9o/M���kW�=2U"O`1 ��!A���S��$� ��"O�a5�̒9�*p��'P�m3�!�C"O���̛�vM)��_�x+���"OH���,2C.�{G;����b"OHd� Ȳ&������Z�у�"O��k@G"��i��� ����"O���$���� ��GI�\�rmZ�"O�!
��A�d���q��[�"O�Mst�;s�TP��D��,���"O��S%C^/24���^�z1��"O�dbU�P-���j0G��af"O���!�[?T��2�(C�T�x��"Oz����6_��"AF�N���C�"O�Hi�O�A�c��
PM�d�a"O�Yp�
����(��[L?��a�"O�d��ᔙ��5"�m��_�-��"O���c%5��Y6��*e(�	"OJ(@&��(����1�Ŵk����"OH(+�k��ʐ�	���}��qH�"O��s�a��J�)2K��@2��p'"O� f/	�9����J�	:.rm	2"O�� 7�C
oKHЈ�A����"O� ��2���"*�ȉtM�!g�@��w"O�dȂl��f��ӟ^���Ae"O�mX���.��Uk�e\�Ht�P�"Ozթ�i��"�$� 
�Ҥ`�"O���(��k�r�b�早[؜=Y�*O4��4�I-+j*�S�RD��*�'�E����E�EjӃ�+�<��'�*Ƭ����B�KrސT��'��ҕ�^,.����OҲdU��'~�]�s瞉9D���ٶTB=��'�n��팬l�����f�&�>���'f=��s�,�p�戄=!j���'�����W-0�e�"g�^ɎQ�'�rs��!�V���׌W(�1
�'jrm{��S'�*��Y�N�Y�'�52�L��X�p���*Y��}��'6�}3�mJ�V/�Y�U�O@���'��-@)��5�V����J�&���'��U�q��!�|=�CfMpT�+�'��Q�E�D4���MY�X�D��
�'N)��G��j�����S�~�Y
�'y�]:4(��N��)�6���Qφ�
�'�dʲ�Z9*�]J��9��	�'���E	�X�~��!��-+NH�'��wf�U���rCD�V�`]��'1`A�B"��n�<�{&�UeJ���'kTղ0i+�މ�����[�p�x�'7��3���u <X"g��!I��
�'����+��Ed�,��l�:��YJ�'�Zt��N*DP�[7�A�	nn��	�'�&ă�%�g��m�`��0ș�'�����@�a�f���~Ѥ��'����d�4�z�q��N�s��b�'����u�0	�|�@� h��`�'{ DZF	�N{x�7iF	����	�'���W�L�r&ӆ�5cDe��'z��1�l��qʰ��DH..����'��-�&o2C*�U����*��Hi�'Fh�m�
x�\hd�Ϫ���0�"O�X��&b�\ �ȑ=:�v�s"O���F+"���1jT�$V�:"O�ic�JQ�k�Z��q��;��L�"O6,�����<�f ��g͌K��`��'3yi�
�_L� 33 �,`��'�*�3��3w��y V'S�k���'V�;4�ۃIF{�*ưcD<�B�'�n���ٔ#0R�"PJ�'M�$�:�'`�8#!�Ո.�d��̯-z@��'��<2ЮA.���bD��*���h�'2�H��,+*@�{e���ԉ�' ���>nD���ɵAF�
�'c��+��K5��
%<���
�'/����K�ޑC�����1�'�pܻ�_�!Č�)AD�`v��
�'-��� ��7I�rDK�J���'����҂F%�0̚!=yʡK�'7���&n��Y0����Ϲ%tjD��'�ȤZ�`	�iY����p70 �'㞐@��,B���ޔv�D�#�'�D��f�=15��X��3S���'�(�1� =4���G%D:|@��'�*� S�D:B��)i\�.�`�'�h� �+dED��s��4S~���'�RI��CI�.�V��Ɖ����x��� ��0�M&�� �
�'��"O�<��EW�qq�qqc�G� ��Y9C"O�k�*H�I��+A�6�Ae"O	�r�ě*�,���3	� H�s"O��s H#��2���{�½H����,AS�LN��iũzl>��%�M"�dJ�GA#g�qO0����SL�A����8�F�s2�=~ȅB�O<�+�������bpO�.7�������̴9�]ڢ�x.��$h��g��p���P1&˼�)�(�+q\i���.-�H�r@J��b�`<�"a�<)����t����MS���)Ǻg,p��%}HcǤ!Ȱ�ʱ�'L�O£}���$ΆP�eE�pHƝHP�T����Ğ٦�(�4�Me���)8�q�LT;%����$#�w?�*W:g��f�'C�)�L<��/�"m7�]S�
C�iV��2��G.,�4�Sݴ]���	�i��f��e�Ţ��O�����b��w"����Ȟ�i�n lZ�z��,��'X�[¾ �2��;6xȜ`�d�,�>��%L�kl��j*�h`坘F8��:�ቯ �MC��?i����O,>7��?+x�2�ᖈ
Ұ�$�W#
����㟴$��G~R�U��ʨr���_: ��L��(O¨l����j�4�P�$�48�
q��]B��]�pr4�:�M#�|���x�g_	N��f�J_�d��NE�����4`�RĨb�Դ4��I.�OxQ�A��=x�X%R͌�\E4���"ۍ/t�}����|�%�],�ݐ��Y���*b�n6ܕ��4��j�<`�LE��(�!-:�`�DQ��g*�O��Oe�r�$W�p"�*ؐX�nA�2�")sjS����hO?�ĉ�wܒ��Eӓ"g�U�Á�(S�����4K��Ɣ|�O���W�x��	�sܬ@3'f�w�Q &H�L
���Fʊtx�T���lr.6��^�����/�3��5��'C�<�R�p�	�l�:$H�(]�o�"?i���
{ހ�ׁ]/ ��xE��𐪥 -��{AB�1Q#RO�h�伱/Q'#EXt9(O�����'_����5���ɵ���{0LH�H?�7-�Onʓ�?�(Oxb?u+ ��r���އxN$�ӥ:D�TK�4t��@�!N���zRa����ٴ9�6T���׻�M����ħA�5Z�j�MDD cGS;����=��X�����(ܲb�P�A1�O�ڱ�vKz>Ţ3a�4�0�;Q@ߦR���k4ғy¤E���R�b�M)�ɟ1Qr($��,V�;3>$6�5,��a
"��Uè��R����5�+4U�H�.��t�	ܟljٴ�?����yBj��:����N�e���f(_ҟ�?�|�K<�F����ఁހZ�pm�4��g8�	ݴ=C�6�i
xu
wĔ�I2��R���P�@j�'�R�ۢ�v���<�'�zL<���uz�u
V�M�Sg~�ڴ��;��)�!_�pZ�y'�3yd�x 2�Z�'���8����F�9= ���s�^�$6͑�f����I�A��b4fE� 3S��"��åU*����hi�E�3�d˂,@1u9���7�i'x����Z���<%?q��M�&�;E"yXW�L�i�
�-s�<�GU->$�MR��^�)��ӓ.�y?1I>�p�i�T#}*[w���� �ց`�a+D��>�~5���(��9lO��9`�  �   ;   Ĵ���	��ZP�viė:&���3��H��R�
O�ظ2�x�I[#�x3۴|f�v�J=|L��gJ�'��l� j'�6-�轢ٴ.q�$0��\�I�F�p�� I@��4��X����f$?�!�r#<) �d��&�R�~��� p�<
'��`�^�xQ��A�Μ��'?����6}6-L}�D��$�A����36�̣ln*�c�CN^y�C�ODcs�ʎ��9O4�y 
�/��cEI�6\��L���X����b�8��D�`�葰1����'H$�n��$iq��%F��P���q�'�dS�	�lu�'�����K �R�	�7
�j�h�'B,FxBDH�'I���vjƓ4�T����ܥ/I���O5Ku"<)pI�>C䆚�J�PMV�M���/�H��OT�R������'s<!��m:����)�*rY�8i۴;WH"<	s5�Fa�*�Ɏ(75Z� +|�;qh�Z�>��#<1� ?� �B����P�¦.x2�Kc��Yy2��~�'���?I��ؗ	h���'��MY|[Sj�?t"<�e8�2����н)����B�R�]v���s�C1O<� ��$����~B���p�� 7|��ukƐ���lT"#<�m5�k(:�R�^6V��-AfՈs��x��o��X�K���i��mGDq�����|y�@�3z���*��$�B�<a��"T��P�<�2k�3Uo�O�2��>R��#%
�f�>I�s\�l���I�-C��Qe�:2z���P�:Y�I�"7D���'K
   �a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  '  �  
'  �.  B5  �;  �A  H  aN  �T  �Z  >a  �g  �m  t  Iz  �   `� u�	����Zv)C�'ll\�0Dz+⟈mDԤ�57���DB�������$)�9�R��<5G D�Eg�  !Xm�@�߶>���VƐ=-�I��~)�U2�'Wꊠ���(I��A��{�>��`��H�t)�#GJ��x�R�<2�¶^5���Q���������,���0c�Ш�aA�H���EbN�R]e�pJ�8Q���5 ���"J�9pX�q�4gn�<����?!���?a�K����_#>�xؐw)M;9
�����?�1�i�*7��<���hܘ�'�?��v���aD��[2�%��_c��X����?S��Ɉ*48!�	�fl�l�p��A7�̠$�.r�F� A(�,q(@����<� d��1q������℅�F�g}4O�㟬���R*-��'��8�Q�B�s%���Pl@hܼ����?9��?���?i��?�)�,�ݾ �j�[4?S0���%C�=m� �d��a �4(���i�����nZ��M���i��fg֌
f	�E��+ZŌ#=!v��s�O������9Ahd "%.��#0�,���[Q���EG�u��� �i��7��ԦY�Ӯ�RdK:*��X@f�z�Px�E�I�lQ\{r�t����P�[�.�s����h���I�Dk�7���޴�z욁�X�E΄��r�ZRːH�𢅮)���5C�����GyӸ�lڶ ��9s��%{Ӳ���D�<(tM�gힲE>�Lˣ.�:yע	=��i+pcϰ{�I�ߴ��/o�L�X�g���Y���� cvO���`�ϒ�d��CĪO3d�܈�iZ�dz��N�`xv�a���AR���'�O��aNIa�+r��R�
���g[��� �f
����شj����O�4�;Ć ���@+"��l$����ވF��i� D��'!�D�h��p1�`�V�#�25�!�O�W� U@�G�0�H�֯��!�$I%Yn\�PJ%M$v�&�O ,m!��JנxXҁZ�,��cl�:=!�$�0@V
�bağ^���yeL24ў r��/�NothP��'u�(y���%���"�X ��-���#�Z $~�ȓY\��CHĨ}�x1� �M�r����=�u�8l�]cco�b,��ȓo�$�D�;��\��?l��d��@���:�遌|w�!g��72��	b�#<E���שrm$<��%�"l�Lp��ږQ�!�$ۢh�n�iUÍG��\��NLA�!���#�QN+���5�F#�!�V�=��M"`�A�\ 8�,��!�d�3H"�B(�_�P�	�`R'�!�dBn&�C�Kg�PR�	C�)`�ɑ2˺��ĉ�s�(ib����0R�y�B	��js!��(&��x�Ņ4���x�悚 !�D� V�����=B�&�CE�	!�$ݘW����I�j��8C��܇/!��.q7��i0痍i���A�����yB��>d��6��O��N��B�y����j�c5��$�O�H���OL���OF�p0��O�˓�y��Z�uÑG͙t����A��0<�BnU��h�	6mz�		��M+���N���В�W���D)}�2�'x6��O���IB�L��xd6R$1X�%�<�4;��O�d�ɉ-��̣#�OhQj��ܓOcZ�QSD�2yx8�qd��*��|J��'�L�	<:�dRQ�I 1x�������!�����O�˓�Γ�y��7���6��(e�M������$�`g�
�{��	S/m�>�2��ڝA��q�q$�K�	%� =ʗ��S.P����%BU6 ���
 6`��K�� ��ٟ�%?a�|����O�����Ul�-� ��k�����	�q����ʣj1��ň^EF�?)���A(|��@пD�hEz@��>X�H�� ���3ʓW�����/�(*f�$�<0���/� �)y�bܲӈ� <��z�\j�̢~m�Y#sL�3�����yZ؋q��cr�$Ӓ�ŌBv����&0���Gݝ.�	��^:E�H�Ɠh,`�#q�&Xk�Qņ�.;-n��G���<��q���]Z�L�p�T>]EZ��D��z<��#p��)��wL$i�ā�}�ֽ���'p�@�"˲Lۀ�	b�"����B����� �ز�R����e˹v⁇ȓ���+0�ʉGR䢑\ ;�,�%�Y�4���� ����N�;Bt�
&�O�l�L��w�@��?�,O���O�����,�\���e�.�.�P��!D��� Y��&����(1���ټA'f<�}5�l�ab ����J��Fd\1pq��!XO(�"��N�/�3�BN ��On1�`�'��u�"}?8����m��2!*�D�O��(h�)���'u��1�D(z�����O�yH�f�aI�!��xq�T�'p��O.���4�?I����9H�b������Ԉ�7n�d`JF	��.g��'���r���t��ɣ�@Ը2���T>U�O�|,�@*�5�m��K@H�O�JWO�(�\�h�֖\w��}J4�U��!��F�R��h�F�e~�鍢�?���h� ���0��88�kR�N�>C�<-�iʷ ��g���,*Pq�����h��d�Ԧ�St��&���4�g#j����<�wS*P��'"�'��I�H&\ӣ��	MӼ Z�a�z�>�d���b=���P~���d
�K�d�O���O��s���0�@1I4@�
$c(,��_$7Vx+�L��1��܊rL�~�UFI���F��,$��p2��$�?�´i��Dp��Y���	�N��8����;*a�����.ٔ'�ў�Gx�)�>R'���U^��`J���$cӞ���Ozqn��(��ꟸ�O��%#�)�-9�6�kF�ܰ6#4�b�ሄ*�6�O*�d�Oʓ��Id>���_���1yÊ��&���'�;���"�Ͱu�Co�@�FrJe�5��+�.8iꁣ�"`#lR-�=r��ˇ����_�+W� ����(O�E�D�E�$�1U�~ĉ�B!j�b�'�6M�O�ʓ�?i,O��'[N�]#iL��Pe9�,G$R�%�l����}R@& 9����ނC��������M�����?YC���y�5F�F��׍ _���� B��y�kҙ���$��5mzy9׈ ��y	�T�P�Aci�!�4��Ù)�yb��~���2�
�;�L�����yR�\�k��ѴǏ��(Qk�I"�yr��(Et��� �={�(0����hO������&!�,PmV�\���Kp ]�8�C�I�
���cAL�v�j��v�گ&�C�I)ee��K��0@`~-Z�� o��B�ɣ>��рh#���7-E�B䉆CVZy�'덡m�,�`�ҵ:�B��;,v20��\9~U�aQ/us���ܬ�"~� �G��t�ڳ���:ǔ��d��yj��
��c�� 2 �c�� �y�b��c/���A� �}�i�A@ۥ�y2G	�&�����jM�
Q�U3��B�yr�ТiF����YkP��#D��0�yR�I�^���XP�_�c&*4������
�|R̀*��B	1Ea��flW��y�%Q���Q���&��0��bF�yb�_��b2���Q�.��e��ybKq�,x�5>�`ti��V��y��Η,D`Cf�$n�n-�%f����>1҉Nm?Q�%�\u��e�)]�ڡ: O�_�<��(�,"�6*�I��X�6ِ&(�C�<��R�#E*a� !�䀐�<y$)�CO�� �K�� �2�+�ov�<)A��;,4�U�Ӝ+B8<c ��r�<�1ǉ� 4E ��A�"�0�Vr�'6�1����>jT���Pe����J�P!����a��F{��rn���!����!*��X:4Xzx�,Λ"�!��t����K��>���t*^�!�$�o#��6��=܊,c��D~�!�ą/.�X�ѥ⏬-�Na0CF��&2dZ��O?�J�"x_$�jĤ�)Wԥ  ��T�<)�m�E��ҖL�Kl���k�M�<	4�VH�8�2��jT�1H�H�G�<���&6Y^Lk�� ly���� �]�<	7�S�|���pEWc�h� �\�<�F͗�%dH��B	}�̸�Uy2l���p>	��p�9����&�^����6!�� ��B�HƲh�:=�-��N$�9""O`1@cH��'K��D�E	�B��1"O�y{gǁ�3�܀��+����(�"O<�c��ҡ<Tu!@M�='��"�'� ��';ƘpP���f�{V�T�}�
�'vt�ڐ��:c�v(���S��)�'a$���G6� �vK�-I?+�%D�z@�Z>�ȍ#%n��O����g1D�T�EC#��I��E؇eq��"6f$D��;�ۻDx8c�	\�����.�D�AG��gZ��T����s�M��ݝ�y���?L&�m��[�'��)I��y�	��V��-���K��B�"�ybMŶQ�YĄ���}؆$��yRV)��ǈJ"y�Y�����y���GG���`��0�~��TeǑ�?��W�����Kr/�0d�"���a�h��o���y�"Z�I%���dC�
 R�)q% ��yb�
�t̠�)��u/��p!���y���
3J2h	�)��v��o�4�y�-Ղg�e2���^���헣�yR����l�O��[K��"�����D؃*��|B��%�:��d�CH,�[ƥ�y�HE1��J�2D���v�ʷ�yb�Xb���qdű7��M��&3�y2�/t�0-�q��4�tm�����yҧ�n�0��B�[� ��H�������>	sdWu?���0`�i��;vtҀOB}�<Iw�F�F�81ƍ�?P��h��z�<�TO�G�ޡ�2�Ć6��E��s�<�cD  ���h��
�T����j�<�r��5����LǔVT�Al�<��h�>P���@�i�n�1��L�'��š���L2R�D�Q㘜A�0�[�o'!�)Nנ��u�W�`Z,"�cҥr!�Ow�d�F�*&xǌ�9$!�$T=Sz�+�8-�����(_:!�D#�������8���zTA��R/!�J"2����� ޲�ˑ�Ͻ�R��'�O?i �PSK��3�h��q���@�H�g�<�nW:DL�	��:3�R�x I�b�<	�ǩe'��G!�8>f~+0�Z�<�VI̸n�������5K����ΌR�<�5 Ҕ!��3AW�8�bl�vʟP�<!T�Sd;p��%FhqRĪ�Qy2N�(�p>�!� �c�:��e%R�>v>�a2ɎQ�<Q'���P��'��s~�ę���L�<���� �§	kn$����L�<��*�Hݰ�� w��R�%$D�X��ł>+D��*��%-|�uB,�O�E��O�9��-Z�Vİ�ȖM��Y=�y�"O�]&�Է|��Hp@4�!c"OV�����A��ʕ�k��؀�"OB�ʢ�<M�A�O01�hPs"O
,�P�X�.�NUCb�z4���D"O�mqe#Y]�d� ��@�iE�DB��	����~27@X0e�ؠ��A�O�\���g�C�<�ǃD�2$IWS/�<Q�"l�g�<A��ןo|92򍐑K��8���}�<���ϦQ=��Q�
$����+�a�<���9̢�iˆ+V!2e$�`�<��oR!Q���'�Ļ>��Y�fEß���j&�S�OI4��Rep�,ЧO�Bc�M�4"OX`�,B�B��<+& (�)u"O� �XG��$��x3n@:a�.q:�"O��`2���ex�J=G|��"Op�rW�L>S�����;4�Р�4"O�hr�n�Q�΍(q*�� x��V�d��M;�Obu 2�ͳ
h~Y��IB��c�"O.pr�Io�z�#���%����Q"O����&	)Wb���&H�H�q�"O� �X�0�썒��[��Y�"O�UM���+͊(��T���Nx��e��"�n
���ZR/ĿW����3H!D�)�%-b%bC���dp��`�#D����⑓��C0�IU��wA>D�q�O�yz��CE�WmB� �?D��{r�6bL��$� �3�F�M=D����Ϛ ]�.,� .�
o��E=ړ
�D����`>�T! 9?Z(Бp���yG+V�I;'#��9�M�l��yBÚ5�|4�E��(]�`��DT��yR �*JB����[3"��Nޒ�y�"g��裌��H g����y�R�d2� jE%�^`r�ܑ�?��l�]������&��"bi��Bu�ޭ?۠�:��'D�l!m;/K<-�bG'[�L���'(D���HO��
ࣧ������*D�p�#��'h���D�BF�1@6�3D���-�d��ɳ.T8*��]��`0D��X�G�$E�(8c�7/r>d���<Y�Sb8���ч9I���ф9 ~���)D�(���-��Qr�9�Z���(D�(�.E.8�2��mQ�xeN��4D�$�2.W�I�,9����H)3o4D�4��j���`H���5Ԅq�g3�Oz�p��O��rԤ56�����JQ�N`x�A"Od�0�����M���_{��ɀ"Od	yV/�NH�a�M���W"O����>1���"`���""O����(!f�Y,1�Q�w
̎�y��Ξq18e(B�����d�&�hO�CD���:�h$�E�{�V���W /��B�	�\>xܪvdN�l&K̅b�V��1"O�����b�*0�0`ȶ&�8Di"O��Q��_���$�P��t"O(P�7EΤ"$9(���L�9�"O��	��0g�$8��5h@�d�'�0������Vk��P���
�2��� h<��x�]�ޅ&�1��C@���ȓ^f�P8e�bD��R�Go	.���QH�)k��L�'<�è$f|��ȓSX��� �X4X�B�x��ZC"��gt��4��4�l�q$dԜ	)J��'�.I�e��@@��68��X��W&���ȓt�Jp`G�:zG�YCc�@�oʝ�ȓP%������+'9����-�P�
E�ȓ=��,�!*F5��4�U�G8m�=��X.�8q�^�%�Z�2�"N	c�<	����}��	8
X��OR>�bJ�5��C� ,0��5l۬ļu�� ?w�*C�	�+XZ����:(�H�'�1Xt�B�	#Plj�j��G�Q0H�B`�ж|�B䉩�D�:�G_�&}ZQ��a�a�hB�cU�E1F��2P:��BV�=�)�j�OD�[Ƃ�4� ��tB��;�@I��'ۂqj2�ӬL�h�B�1�v�(�'�Hl"1�%I�@{���}�J�x��� �Ð�V�f�賓�*Yܪໂ"O� ���6j�F�� F�@L�t"ODL2w���z��p!N�C��%i��'x�R���ӡ��\C�ȇ6~�$L�I�+C�|��<E�	:�I�Aߢ�L�4�^̆ȓYҘy��!�#��؃�R�dԅȓVi��ע�$m�|K���;�&I�ȓ��zC�G�
A&�q��O�q�*��ȓK���΃6���KL,��'�$��W��*r�b���Qe��\��ȓ������S������ۥ�꜄�dC�y	���+��l
3��%򪑄�O\Ea�i`OV�26���i�ȓ�Ф���R�<��Z�+��p���	�m~��ɶR���H;7�Y��@�7M:C�	 v^�� %P"���b���<C�	*+��m�F�פ�����B�\�|B�		�;�T	.p�Ѐw
xdB剷=ex��w���%W��2��V�@�!�$[��=���XT�2`��_�ўаt/)�5�~�xR�e�px[5$W?v�L�ȓ]�PP��{lB�!�M\�uT1��9?Sq�j�E�Fg�
>ε���Nl!�����	�$��&���ȓ�2��%B&��m(�չ\5N-��!�4R#)��C��ř���3=8|T���Jm�"<E��CL8�S3�ZMc&f�rh2"O� Iwb�bT�A���s�!Sb"O���⏿E�u�r��7���E"O�s��4 _��)֋��E�4�t"O�Y�B�%������D�OPp�F�ޠU�����/<�z@!�f���'{��n�,��'z��z���B������� 8#� ѻ,O`���OL�䐠G����;=�2��	'@������!B�D`���L��I�]W��">���F?�TI��+U$ �j2�j�U*ld�eb�rj�%T1r�S��à�(���jD�$�Oc>��pj� �s������V,�<!�hp[�e8;�[�8�H���0��D�j�@%�#�"4��#%兪T�剟8	&\��ԟ0�'c��П4�I�!�<�Մ�4���: �g����ɷu"0\9 �~q `ī`�"�	!��u�O��� DCO=9�(��D�Ν�`�'d*�@L�!|���P�(L,؈ )�eB���x�}�`=&�(����%*p����<Y�����	M~J~*�O�sTAM8 �dQ���jޠ�E"O&E��Ǆ�T5"0Q�*�i��]!����ȟ�`�d�}،�ʹ-�lK��OL���OF��C��(<��d�OL�d�O`�)�O&{`B�k`�C�Ş������Q�1Oem9fiZ|j@F\�*;���O�b���G�Kf��R�D��VQ�5`�[$G萰� ��H].c��&Yt�'x�x�)6,i~��G�.��]zGLZ)-"|e��D��dX�Rz2�'�ў�� sщ��T��)�+c�)�� %���fM�'A;�A��]�S>��I��HO���O�ʓV�8"�8OȲh�� �媀����7y�ڀs���?����?Q���?9�����F�����')��DU�	�N�-���8Aa��*�haGC�
6��&#�H�'D8i�酞A��]!�l�1g=tE ga�A�Qiۇ0����E�@x��q���O��Ñ�'S h�wd�����F�	fE�yzD�'vў�E|�����[�:FJ'oH�o<R�ȓKyL��dJԒV�����Q�T2Bx�'��6M�O2�\�9��N��i���4�\JЊ����_&��B�_-�?a@���?q��?1Q�2ۦ0��U�gH8��|�Cn^�w$T����G�x��1G�[H�')bH���Rf����Y�C��8�*tH�	YoS�M8 �	�7�4���ORc>��F��d��ط�̝US�(�b&�<�[��!a�ϔ}yx����l&q��I��d�-c�F�C��1xI��	�H9[��O�4ِ�9���?�	�K��v=R-��YvJ�$�C��&��c�p�uy#�;�PC�I?I�8��p��l`�E$	�S��B�)� (������huRb
�z0��B"OȌB���B��юV�0���
�"O���m��T�A-�)�LtR �Q�O^�}��W��p�b
n�13��+�䑆ȓHg�%�F�X�-6N���7�
@�ȓc�n�A!�N�1D�Yۡ��N�F��ȓ`y��P�LyI6i`ceٱeT��ȓ!��kPck�X���/)Ϫ��ȓo.R���:p��+%l�6.p���&>����$ۊe��	I��3ΰmƦ��C��G�=��*��L�x0��1|�fC�	<�q���ɻ4��ك�6YbC��'e�L�ȀGH&3Ȫ�(���u�VC�I�7�ȳ�A�A�0��g����	Z�P�'N28�N�
f�@�n@�r��U��i�'n�d��'w��'��h�u���~?�iK ���a��7-��uw�E:G��pW-_�8�����m��O����fekA��-�p��)I0��*���E����0���(6��  ���On�d-擔6��[Hsj�󷥍�PI��0?�p�-���R	��
.ȵ�V�U@x�H)O��J  ��m�-��N�?a����^���I�����|�'������� ������JMm��	U�'�ў����ʄn��z��X�?�l�!�
:�Ɍ>�Oxb?�1��6��	{c�@4xЊ7M;?��OԂǒ>��y�M�x�0T�T�ؔY��$�$��Lk��8�O���@�,}�� 񩄒N583-�I���g�ER�B(K���'��>牎^D@��6��?Rɒ�[$DT,����U�+}�h+}�������i�h�@
�m��\1^�a�F:Dh�aK$��ɍr�Т� c֤j��q���J҇�]�?Q!��S��@��r3�_��,���L�%���p	TⓂ��:$��`��?5�"���CV��r`����XSv����~�$	���|�fL�Z���?��n?'�)S��JV�͑�a�7M�d�'��H��O��B��i�8�z���պX�r�yrc�_�mV[?t�MS~ʟ��T������8팯[c�1�ԡ�>k2ie؟�أ���]�������,P��5D�4��>`����Ĉ)���e�4ғ��'�"�'�Paɳg�~�ap��X)/�	��Ʊ>�K>1��T?��\M/�4Ys��/ZHX�
�M�y"b"F(�(Q��|{��Yw����y��Q��Ь1b�������V�yR��0
����!���Zgm^��y����X�v�֕��`6�U��y��?dZxU�0JM��Ys0���y�O�!ҹ�w�>J��5�FN��y�Bߙ�J�[fF0,�,bvl��y2�� �FAqf��?W&^�yBM9�y��fL ��g�RI��P�fA��y�n�r`���XEN���!�U��yB!��$�����-g����f؝�y�-�:��0�&��2	�6iy�����'n�}¦l�-q:����m�!r���"b֎��7a����̀>њ��͎�X��@�
��%�4��Q,�?�48��b*�8��Qˍ$,�jH�0ʁ�!0N12L�!?���b�L>`���h"�7gp����
'*���fiɓ϶���6$^lq�1�'T�j�O��&Ď��*p�c£
�ؘa�IBx�X� Ϥn��Y`�ƥC�Ĉ�'.D����a��L����FR�ZLK��*D��8�ˌgY��2A��(�l���&D�0HrKM,>� �����Ufh�A:D���-�=NZ���Al8}"�6D��A6���zV��x��A5D�X�a�'7#��;Gb 6���HT�1D�T��,˕1�VP�H�U�r��u�-D��{���Q"��J��c.Bգwb*D�`XDA�)i@�r�CU�HWڰЫ&D�8�#-�,qF,���2 c��d�#D�P���ѮVxz��Q.(d�v��+#D�� �d���K�?�r��O�9���"O�1*�c��z�����i���e"O�0q�/��Haܵ�W"z,Y�"O���ōT|�����v,�1{#"OV�K��.ঔ�vA�;����"O`HЊP�\���h@o�!o�&��"O��i�˲8�EKȗ'���g"OT����>Q�M���M8p�d�y'"O �P1��� *���.,-:x1C"O����D�n�x @��Q"O�(��$�1}-N0DŒ�N�aQ"OL�`b�Q�q���S:Z-���U"O�(��\"��� GŮ/ (�"Ox(P��I�2�QO�&2�T� "OЌ�E,R+ e�M�;�*�"O��з=l�3�^�v�Y1�"O:� ���0��V�]-O�0�h�"O,�)�j]�s>a��	33�"O��Ħ�ck"M�'X�c͎h�s"O>�S0-N|>����׆�b�"Ov�h5��0s�����0�J��A"O��9�b"+UJa�����a"O~����&��!���A����"O���3!}Luk�	̀��]C�"OHa�@Í�%]�պ��\�m7T��"O�Y�if~�u�'�V��"O.AS
��O+(� f╖��ڑ"O�E�*讁(C�W$+O�"O���P�ӧh����HQ�(�c"O4͘�JW>�<�k��/�x�"O�Q���k�8hKed�lG���U"O��B���NV �A�BJ�J��ܑ�"Op��`c�$����ʠS���*a"O`s�V�p�T���W?{����S"O`���# ���h"�t���"O2��U�R���0c�� D����4"O�ѱ��8&^`�"��>m"�ݨ�"Oz��cOC�*�$ɣR�V�IT+w"O�=�@CY8@��O
�)���a"O�l ���[�(Ĺa㛃V�z�#"On}�A�C�R��$A�4�T"OX�VF��)6��86bׁ_p�yC"O����%�GY{��X�eD`M�5"OzH1�ㅅ��A�" P�q�-Q"Op(s��2;j4��W,��G��K�"O]rRo� ^j��&��CӾy�"O�Pq�b�&E��@
!'}
"Opa����{��8�&k��^4� 8�"O�y2Vㄺ���E�?��J�"O�ev�_�d[49:���dĳ0"OV���D	)C���eش&�x��"O"�3� T�/V�C�ot ��"Od@c�I'C�	LY`��"O�D�$@B��y�e�D�ȫ�"OO�դH� ն��gA��y�Hʐ%������C���Lkf$��y2F̛X5�)1g۲|��ı�$�y�!�*n�0�Q�b�+�|�a.�+�y$��H�~YA��n\��sH��y��/}Π�Hs��b=�t"$ۚ�yrl�.�dD�QIюU5lK�+A��yR�7
�h�b���L�,��'%��y�Ws�~��&L����7����ybH�W�N�2��_B������y
� ��P2 �Yk�%���ƈt�~���"Oލ���'Y�Bq�2�¡Q#���"ON��	ڵ7��Q��Fdaː"O|�3l˰A��PS�ζ:i�)"OVѪ5��%,iR%q�nT�tc���u"O���Z!(�� p�+�%��)�"ON�R�e��jg�X�
��V�`l{�"Oxq�J�g�@���5��Eڐ"O�$��>���ףĭ$�b�H7"O��* MF�G�u�5h�o����C"O���#�P~ ,�(4�ͮ�HT�"O�T����-��,�t��O��mE"OZ����ւU1D嫒cU�t�$�s"O^����1$��y��A~�U�"O���g�A���{��
�{F��"O�������H3a��"CV000"O�U2�^�>�B�Ceꑑ\2�x#"O����P?lq:5��O6��"O,�����(�J�RL�5Z/�X��"O�hR󀑴C\~,�jߪk���@"O�չ�f� Bh`��)��7�LԘf"OvK��&-v�:���9�B�8�"O��'��OU\��ՏFK�483�"OpL"��)+$T�z��:@��z%"O:���$B1eAZ��6*�p�<�[�"O�T�t��|t`4I1�Ƚqˮۂ"O�\Z�\9CA�YHUO,Wa
%3�"O����ރXb �@.�(#�(�"O����GZ�v�X�C�Q-Ӛ )a"O��O1�>Pr���W��)"O&ؚ�ƋZ������3|�p���"Ol�A�k՜W��G�)*��â"O�a���rWT@T�&�v%�v"Ov,���a��D�o4!A"O�Ɂ����Qj�
wރ>C�-��"O8�)g��*\%�
@]:���"O���"NF�gj88��Z�k�ȩ�"O��BC���a��8@��* ���f"O����n�n��'��Z����"O��!��h�T1�G��W�д �"O�l���B�Y�<-zD;��	C�"Ovy�B�X6&	�5��#�P���"Ot�#��U��� x�̯F�-�v"O�`���G�.!0@��8'~�k�"O��n'��tcl�)s��q!c"O�h������R��ǻBB*��3"O�D��Eՙ;L�X{egՉ)4x��"O���'��Z�2�[�^�=��Cb"O�$qC->A�5�C�(F��p�"O�����2*H��$�K6u�t�K�"O�M��EQ�q�5�2ۜl(�*O��'邉=C����b�W\+
�'Dv�r�E���gI�!xF��'�vu�q�ջ�.�" !�����'�F=j�M�-W�Q���ދh��j�'�����=u=�q�ʼft���'��% EQ�ڍ��mޛV��Y�'�����@�_�fe	��P3TZ�-��'˖C�
�O,���V��B��C
�'uR�ӂ��'&��aN'�r����01펩Z���h�Ϝ[
�'!^�ze*�.
\�BqnZ�\n�@
�'��t� t��|����&o�Y	�'HD��V��?fLm9S��F���� @�`�])^2�e�d�c�"O�ȑ%�3�L��PТy�F��"O�<�t�L�a�pdM�|-:H�"Oz$�bO���C���<��B"O��p&�=��RTEʓy�T�q"Of<�b↑4�"���M]���	S�"O(-1��3$Xm���q˂��"O�d�-���3�ǴJT>Hh�"O������3*��b�l�wD:�`�"O���4Hú0��I!�K7�[�"O܌#0�Ӓ�(P�@j݊=�p4:�"O� �b��`>T�J-8@���"O��9e��5�Af/N�W*0q��"Ol!�CM�d�1�/	�D��s"O�1���V�AmF,���()�x���"OnU��)���i�(��M�"��"OH�C)�-Q�N�'R�<I�"O�%�W�� 0H��r�&�\�"ODIٔK�m0��Ci�<Y�v��"O��V���	�vD�3�ˢ9���p"O�t ���+}�R�S�~�,��a"O8�Q�˥@�2a٦�FH�\���"O�8
��$*{2s!�^1d�h�H�"O��y$��
3��*���/{`]p"O�+�
SUt��m�T"O�!v)V�T��y�3�[0-_* �f"Od��7���P6>0��Ù�;��)A�"O��Q�X�(ȅ��	YΜ�:�"O8x�bW [����@-��,�C"O�m�u`�+t�@�MN�fL"ZR"Od�wM�-ilts���X7J�"O�p����n��ِ5mT��H�A"O\�j�BU5��yUꎗ8�h�"O��Xu`�7 �|R��4m�ѩ"O�@{V�U�"��"Ā���Ѷ"O�!6mַ��Q��%�<��"OP(��_g8�(��b:�d�C"OBm���R=w%���1BE*z2:TS�"Op�aC&P�>�"�hG���x�+�"O���0��2"(��2W���.pPI�Q"O��R�� W��q�S���h_d��"O�p"w
,{�6	��ϯ,Zp�:d"OT4*���Z�ֱ0�%�}Qp=��"Od�(�+�M_ �q$F�>���c"O8ݩ� �%q(W-I���q����yr̦V�U�Lď.���k�G�h�<��P��j=R�.�C4�x��.�i�<y�	Ȓ�\9ȥG��AP�Hq�<	u��*rK��p�`ƪӒxy�-�o�<��R����'�V�h(��ۂ��n�<y1`�g@-�B�<�L ���h�<ё���3U�@��J+���t�f�<	�H(p����X�<� �1&��y�<�'�2
L `�ڢTa)���a�<��JX�����ݜ*I�"�_�<�J�li��pbAN��QdI_�<�#.sZ�a�⠘���XQ�Q[ܓy�Ԭ�ЬE8�����'�,�%��i�삌i�P1%��6x0��:$'/D�@�b�:2j�ܑ�ئZ�Z}Q�!D��`�o�Tx�a�G����*O�l�F�O�{�YPB�� �x}��"O.�q `�0ā�,@���2"O����G��С% مq��`""O���t+�v������| �*���y
� 0�@fH� Le1�Ŝt�B��t"Op��%�d�"���%֭tߠ:"O��X�ǔ��h����#!�I��"O��pB�� E�ڔcD������E"OX=��M��/ڶ���*�	J�q2"O0-(u���R"��8
��2���Q�"O8���M�g�.��ЃZ��) s"O�p�'���?���b�CP7la�I�!"O�}C���+,I��HJ�xE<}��"O����c��|;�Ua�����"O*@��oX�L��\�.�&l�ԍ9"O�y� iƘpQ\�"� 2T��=+�"O�yzF!�	G�t$�W�� ����"O�iچ��|�\�Y�BJ�r��Ȱ"O ٗ �%m#�8�@C/5l�L�X�<1��R*u�豃޸^>N���c�\�<2LR�G4���
�9�4M�t��`�<צ�!?�\i�"� �<�qS�
G�<iǠ�_6�5,���2���c� B�	�%X�eҷ��;_� bu�E?B�d�p ���4.�b�X<'0PB�ɸT�
@:r�˦q�L���,.gA�C�	�o%HX��}�p(@�tŘr�'*l�0glI:Y�1Rc��OުT�'G��#UL°ilf ��JNL!X�'�<�K��aϖ)�5�ȸG��9[	�'G0���&zdd��M;L4�a�'VF��Deڴvqx���H,B�T4��'�"�)uG�� ���cW0>!8�'�-c�/�k.e룁�"����'\���Ǉ�5c7�@�F֞XR�*�'��8z��X[tU�h�1:���'�@�G�?9(�W�ܜ7�!	�'>���V���r�6qj���1���8�'�X�aR般Q�Z��рNP萫�'�\��E;ޖr'�9ox�0��'{<y�e&��T Y�HW�d�ʼ 	�'�N�cc�m����sǎ�nV�Y�'���a`��J�����Yz���'rT]��&X<����	�O$��	�'�z���L�}},��-_ L�Q��'���%��z��a����B)�|��'��K�E�l�`5�`%)�B���'G^xU`;�l3&^2w���q�'E�D�"�$CH���,m��'^.-h$cW�^�~)��d�4A�0��'Z��D�4�� }r���
�'A�8��h��J��f��o�Ȩb
�'��r�N^�)�`X�AB{�(��'B�Y��'�-u�8	��쇷p�^���'��t(�hI�65
�������
�'֪�r^� j��S�l�����'(��;��D���]x��1^��}y�'��t�d,��A��AcF�\�����'ͦ}��
Ì���!c�=Pzyc�'O8��ߛaU~��E犢is��'�|1SM+-K���䣊�DA���ȓv��z���1yǰ��`�B<h�lЇ�� dkTY3p�`L1N�Af����a;Q�БTH1�u�͊s�D��s�9�6I��Ĳr@�-C�6���W�����À-;�j)*�X&'�T ��E�re�p, 5'a��I�#j@���^+l�3`Q��-a�.��{��͆�S�? �D����SH��Г�T'A�|��"ODt�m����h����\���b"O�QQ�aוe�ư�˞&~��s�"O�h�1�No�p,X�#�
#�tX�"O.���h@^L5xc�.=���*`"O�IBFb�4DL�yv���tY�5"O�ly��/��Ԩ��4��"O���W.9b�2��L�=�D��b"O i��b�#' �1.@�e��-�"Oހ�@��J|z�K'l�gN����"OZ!q�.V4;�<�"cbTa�F���"O��ѱ@�8$��,�GE�X��m�g"O m�6jI<I��1۰aF!EW�bP"O���dc�v�� ��02��1"O����6 �������$*�2"O��ց�M�ʁ	�̓(#w�p�"O4a��GU!e[��c텦D�|0�"Oܽ�b]�yC61�`e�
a���W"O�!�M�y�(�if�D�J4��"O҄�3b	��D4@b��Q )c"O�C4욃f�4���I�J��"O��2��ɹ{�ZM���*jR�# "O��#s�^�tRRX;DK%bj4I"OB��1BU��Pacr��IM�@e"Oj9�*ީ'za���q��Xr"O�<)Æ �,��	��]6E_�p��"O^X�'�P4+�YABL|���"O
X�t�%3�-qUA�Eʴ�P0"O�Ը�m^76�L��'V���8�"O�$Ƒ�2�z��� �K>��3"OP�;(XXH4[�E�
pj��"O.�s5��	��)���T��1#�"O�I�H�U="9���/ߴ�s�"Od�#Bd/�:]��0<���b"O��0G!��LE�|�ŇϥP0h�kt"Ol�� �ȍ��(��d�!	7X��U"O�US��_V켹V�MR����"O8Q+l��:xX��"�$��v"O���7ꂚ��1�D�P�J}�8p�"O@�W�S�<����%6�4��"Ot�H�	 V�d�H ��9bf"O �B��⺵�眃�J��3"O�P0��t�U�U%�2!�֘��"O��)ňr,$+��7P�H�7"O>9c�dw�~-qAj?Q"ୢ�"Oh�r��؆h�tE+�(I�pau"Oez��7N�#T�Y��`�3"O,�i4��1.JQA�M+I�b�� "O"����Y��@K��	�e�na�3"O�xJ�2R�ah5�
!k
�E�g"O�t�AdKj�t��왕t(X��"O �2	B�~*�)I"E��]b��pU"O�C�F]&9�j욲ˋ�d=���"O�0�AC-pcr�� ��{|=�%"O�8��)M<0s�i�@�r��1�"O�)Jp��1f�*7g�.Y�D���"O���%K�{D��@�E#��j"O:ؠE�)R,�p�O��Y6�(�"OlQ�`��{?�l�Ä�y%�t�"O$=��^7��!󇢊�M@���"O� (Q�&wH2�1&��2L�@�"Ot�����~Ā�v�"B|}�"O��Z���Z���X�`X����"Oj0:M�	If1��cU$,_hI�f"O� xl�@�f$�E��Q�TB��""O�͋B�]ۘ�X@��f�YH6"O�-�����怙�S(�&}��"O��9p��3`�@X`��2;V�"Odm�4��(BY��^=+mH�!�"OJ���D�h_� h�N)T9T�u"O0X��'�%V���4-]�<34��"OTA��X�E��@�F,1TŐ�"Oܘj�)A2{�D�hV�T�2P�ȓblܱ��!V��P�%`ڿF��|������щ6���y�eć.���ȓ2H����.r�$Tw��n���!Ӑ���Ѐoa���vh=8�`�ȓD�H�!�)m��8a��A,	\���ȓ7��BR4�tY�SI�*Q↩�ȓ{l�;�հ�ĵ! M�R��(�ȓ�T�����;��Ȃ5C� �ȓvǖ���f	qx�q��|9��}����$�/q�*컷mҚ(6h}�ȓo(d(�KĢ#��[ ���@�ȓh�����*r�2�AC<�ȓZV|�[DE@>L*�jd�@�j��m�ȓCx~���d�*re��H�� {T	��04�Rp'�����S�/����+����U�N6]|��dO�0ʐi���"��U�V�s����TeL�T��-�ȓ(j��h�M�n�&�üi�*х�7v9p��S��1���K�$�ȓ]�2�tp؂H�i�c�`�ȓU�V�cCJ�1m.����Ԓ/K�e�ȓq�Q�!��~#�M��A�Bh��V�( #`bN'G����1�Ss���ȓڂHRĬA�T�HP��Ї��i��Z�$���(�+��Y����4l|���5<T�D��`�A��!ɚ���1�R�3#.��کP�A]-�Ɲ�ȓb=��$���ȳA��'��m�ȓPQ���gA+TR0xs�Y+E)��Lx,�FTq�(� _t�ԅ�K��֌��d��s��
L/8���P�8��(� ���"CTB��ȓ_�`���/*w|��񃀟1i�d��,�. Pv郅E�H���K��*g����;�Tt��'%%�`��B_�-�Z��ȓb���Y�A�0-���A6#����d��i�F:(Z,J�,� p*����Yr*`Q�&�y�V*�m�m�������giԧ_� ���x��5�ȓw#��s��m�`�R�� )�Ň�n<$�'��5H���C����ẍ́ȓ1X)�P`Q�y[\Kfƃ�v�*u��@2,iz%O	, �6���f�8�d�ȓK|���¥�~����A��`���{X���-��d~���!�T�0�ȓ*� �SkU,�0�"�A1Dh�ȓ�֕3f�Ɠq��Yp��96���l�N))�g��03��h\+`���XΤw�3vX�@@�̞=�p͇�q�έ!(5	�Jq���`[.�ȓW#�� 5�3��XPwB��,uL��jy�Xe�X �ə!�ׇ2���=���K� �Q��j�:�b @�I�\�	�g��A����?9J(x[�K`�C�I�F^ȸy�A2pQ�Z�I����C�ɐx�7�H���}��,9i��C�)� n�@1'ZG1<	�1Ĉ2v����"O�zG��gj�Sc�]AFL�G"O
��K�FIl�ۂaS�*<��G"O��@��	6��lx �-����"O�I���:|�� �E��J$���3"O4���ɕ 2D�PnHP66��"Ov�
 �1C����mp'V��"O��� 6N{��r�e�BL�!���+~�٢�d�nc�T���T�!�d����s�-�(-]+J˚$���ȓ<Fj��q��:#�P�j�犑{�*@�ȓcl�{��oT}
v�]�v=�����!��Np&e�$�@�2�d���!�p���~t�t������a���ڥ�wf3.Uj�	1j�:>w���gF�Z�	�(j�z�*�K��J[a"O�7�^��@L��`�o�̅ "O��B�*!�Ip�����s"O�U
4��^(��7Ξ�E*]!"O�Er(���a�'k�)d'�<K�"Oċ����V��j }d`�d"O��	��
g�P��D�ñ?=*�q�"OL�zS���G���(�=;���"O�q�F�]6�u�#R�B/�%�S"O`��֮�k�yCU��Ы"O�{�ʘ/Q��7��<_�٘"O�E����4�L�G�	�kSV���"O� � X����#��8:�t#�"O�����*{,�P�ac�?p̕�"OJp����$�d"`�1
�$�&"O2�#��$]����vR�}�h�`�"O8ȓ�d�#�UaQ������	7"O
I��B�I%Jy�`�C�A}x���"Oz�e�?ÞM���L�e��"OB�O�	�5cHXԖ(�"O��	\�t@{�j�
L�ʉ��@� �y�#ֱDŲ�;',�*@����y��7�X�� �f[ ��f�՗�y&�*�T9*S($/?d�a�́�yr����N{��-)��A �,�y�I�'u���S!�H�6�B��y|�@�\(�J�KF�nK|�a��5D��!�lL�f��(��mD�qz��ZHB�	�7�2H��%C||`�ch�5}2�C�Ɏx!�͙�gV�g&L`��&"��C��;qu��� ��F6dq�k˛��C�	_��b��~'�@3�Ŋ�RlC�Ip�b�*�C%s�p�!�J `C�i�� V�@?���W!��U�m��'rz�S툼n�()7ŏ4���'4x�1�g�<�8<�'�A!u�,A�'l��`�F�?� !�J�|�����'x#�!uA��K�o�Lb	{�'�B���1S�L��ECT'�m�'�\x��Q$״̳�
��Wu*-��'�z����%:h�B�ՖR��|��'9����C�c�Z� �d�;%�Ex�'����Diو@���4e�n �
�'l��b�-D�oݶ����оeB<��	�'�jw&�;h>���
Y l�X�'a�M3�Iscԅ�&�Ĺ�
�'l��悍?���`��t��);	�'�b���ŢU��K�
;t����'>̭���7v(�B�F�x8���� D�C�՞>؎\"�B��$���['"O��"D�6L��� ��*Mʠ��$"O���P�����b��_�ڡ�A"O������0Z�	K�E��I� "O��,���1�??Fz�#"O�@��nF�T��T�@l�㬽��"O���R�M�B-hƭO�����"O~- '�#A�~l�"M��?&���"O�� +��3��@��[��Ÿ�'�t�PCn�1'��;�I�2V���'ܔ)�͗�)�F-S���<YF�h�'��bA�4XKvA_:Xv����'�.�LO6Y�$�Vc�8J�8��'��X�mɉ�}�����LQC&C�I8�d�+�� �TEy��ǜo?�B�əY.E���D�3+B�$d��6��B�Ʉ_d3�Ĕ�D�R�U*l4�B�I=$��0�&HI��9
�	�>�dC�	A����B�8^?�ո �$o�DC�	�M����dl\\jP�0�f��y�h�,� �A��Q�"-G�4�y� �
؈$i�D�
O�����7�y���+�D�h���^/�M�s���y��߁xQ�鱇*P6[8����)H��y� � PyD��!\*<���D�yR�¤n���S`"�=�� ��
O�yBHR)H[°r�Ț�5i��A3��,�yr�4D�l�#B**2Xɓe
��yLF\tA�1���zjxГN��y2�S�*�x�*6(�8lDIᢄ���y�͑��
��ƫչLu�d�� ��yR�қ/o�M�ե�;@hIs� 
�yb�^�Lz���!�L:D������y��sQ��4IN�`��ҡ����yB�=
�D�8�gS(eb0�t��3�y��ʡ���C���$%ҹb����yBT�S��]��'�3�phB���yr�'�r��eUI��@#��-�y��ԣ]�N<���:.~ET�ھ�yRj�"[l��チۃ@�:H��HD��y&�=v�^���,2A��ra��y��U;(|u���M-�Ȍpc�Ґ�yBD޶*L�$@3f)�f������y2cB�2\0��!�S�P�J���y��,Q���Cʸ�$a:3�J��y�*F6�|M3Vʍ=[MJ�K���y�-�wc�a�j��r$�2�u��jb6��E�$��eG4�.mE{��'e�<�EA��b��"�.D������'��������<|��Ɠ�K� 3
�'͠T�g J$#���8���F��ِ�'v��K��uH���@�˭;�^|(�'r~0�!�Is�\�0ē1�䔚�'ƴu F��0SCE˗JŻ;����'�L���d�&e_� ����/߂a�'4��"�柼<U"u+���j����'b�!��ȏ ����#:�L��'v�DA_�C*�� ��^�7��
�'(nsVB_�3PNtc2H^� !��'��)*��۔+`F�c!hz1lX�	�'�@=R���lD	Q��E����'n��4�Z�y�R�c��R�Iu�Tr�'~����4�����˼,�\���'�ʴ��kF$x���2#b�9vIZ��� ����2(~�}3�E�%F}�Q"Op͒4fV|
��z%�O-Nu��"O@��T��[jDMѥoSO��(`C"O�b��0I��m�����b#"O�T��'I�����=�Rq�V"OΑ��F;O F�lǘ:���w"O��؃IĤ}J\@�X6ry���"OBqc��A�#C�끊L�,��9"�"Ob5y��w�j9����O�d	XT"OzBB�̜����3�Ƞn�ԵH�"Of����n�AƩ��k��E��"O�!�a��)�B!BFW�n�.T0�"O��h�,Z7v����V�*��yE"O.D��Ϝ1V�b����9y�j9XW"O��Z�@qS|��R2A� ���"O��J��t#�#��ԅ.�j�@'"O�F��L������3�f��d"O���b-�X2h�"j�$|�X�J�"O.����yY�݀�		U�r�R�"O\4��P�V���P3*I*F���@�"O( 2'����j�O΄Jä�Ȳ"O.�I��Ӷzܜct���K�0Y[E"O���ܲD#l��B����`�q"O6=��I8RxC�+ʹ�`	2"O�����͜̡ 'k(d�|t� "O8�;� XE
�a���\(���"O�h�!�O#Uy�pbŗ}�(�e"O$D�kQ/sT"�"
+� �R�"O�U�e���Fo�����!�"O���P�7�`��E�}��@y�"O���ukA� �>zP�ƦTR"O���?PJޝ1��NM�y��"O�tB�� 
a��d�U�I(�R�"O`�{S���12��3aX� �8"Oh��F*l�.��D#a��a"O�hk�&IY�D��/�/Y���"O��i�-
�c��@� _�t�r"O
�$%@�J�d���P�(�ޤ�$"O�Hr�S�Ah�X�c�:����"OL@�B��Gr1�r�D$�<1��"O���S��^����GO]$`����!"O�%�pe1��0�X�u����'��,1�рO$��+��E�:zT���'��=���˯q�4e�th@,
pdh�'�>q����`E�����$�9�'�L@�Аt\ĉ��͜	E�d��'�^�D���r�|#0�֒v*��'� �X�oX�9���<YL���'�e@�#�5� z��S�3�*x�'�t!�E�-?��x�`��%S�Ё�'�Z�
�jW���H��"ـX0�'��P�)8����F��d���'"D�GiT���Z�+HJ���'��U�h��'�fx9%�����'�\��H��0����̘�2k>���'�$\R���.�f�+���.?X(�	�'�Z,"`��?Ш���D�M�($��'h�e"!CU����r�[�K�Uk�'�T%�i�-1��K�K�P�Z0y
�'b:�@�-��"Ud�W�Id�y	�'�2 `�'�x; �ޟLA�'�,�g������7���z�/6D��b��P#�,X�D�:i*��2D��I3h]�upt2�BK$i#���+D�� <�2���!%P`�%�@;q[�m��"OV|�в2ǢYB�B%l��"O�$�#ШJ�v��BX�i��Y1b"O�h"�
��'��y5�I���!�c"Od\���0�L��D"�C� �J�"O V�#tR�`�b�C��x"�gLj�<a`Ş�\�b�	�1]�1
"ʝf�<ө�	&��d@�g��h�V�kł�L�<9��_9/ (Q��׼*$D���D~�<ّ�U�lϤ5����5u�jt�6Oo�<9gJO==��8y�-������R�<�7�
�#@���� Z�<�a �%. @�fnՉ(�ȝ	�N[M�<ဢ��@)Ze�e�Ӌ{Zl,��Qq�<�,S��IZ�`�/q�A�J�i�<	�� �&P�R��ۄ	�F� ���]�<ц�*Y� i�6<��T�G�[�<I�ݾ'�ݒ׈��%�r�`�T�<A'��yF`鴪��lŶ �g�[�<�g�'Q΍��A����"�Z�<a�	���ji:�lL�B"����BR�<��,�kZd�FNH�5�[GI�<q�h�
f}K'�7.����ƊB�<�]�C�� 0�kݱh9f]څ'YF�<)�x?<,k"�P�5��Q�!�}�<�2�H�'��)��Z1x�����_�<�cEċTBQ�lR-fu5�@�_\�<y���?f�N��ɚ�;
�!��T�<�gH	�4�^8;���"=+�X)V��R�<�P@G5;c�I�E
�%~���Qb��h�<���N� �� �Ŋ!h�,1�o�<a���?����%�G�a'�Hp Sm�<�ÅFG�,�#��D�CnTՊ�,�f�<y���B����eL@�JH����G�<�E sx<��5A�	4����D�O�<!�/,-$���
�#H<=��lGW�<	P�O%8�9Ο�#��R"M�Q�<���0ftq32,�?>�I#�JN�<��b�uׄ(pV��@��U��j�H�<1e/�_gp�E�hi�#�E�<��#�������^��ഈ�}�<a1��Q����{+d����M{�<I6�ȤW�\�x��O5���c�s�<�s
��v��1���2*Ѱ��I�<��b��K��:���+	a���"
[E�<��j�+:�Ma�.βW~줚�g�<��KܤE?<y0V�L�_��T
GIZ�<�&F���5-^=��8�L�A�<)o
�q���eOe)"P�N�k�C�	Hc(��"�#2q�p�ңr��C�I�Hz!SF���@�u�7�P�GۢC�	����5�� d�)��B�4E�iS���M�ָ3!�0��B�ɘq>��M$Q��;��[�u�lB�ɪ@�����aHQ�U1aO�k�.B��%FyP�F��`�v�Sv�L�>��C�I:lKpU� $]3+J���-׳-u�C�I	V!�1�*��l�(��3��n��C�	�Mdq���2{����b���B�I�]18��7`^9�d��Ə}��C�ɀ#�,��J�vo� ��L��7h�C�Ɏ4^�@�WJ̝X�fL�c_!nC�I=��0�q�E9iTi��۠@A�B�I�`[F%����o'��*p�B�)� ,Qs��$[�X[0E�(h�Yi"O��rˊ1�{^͸Q���¼�ȓYZ��/�� ǲ�0vNA?�J��ȓi��H��'g�& ��ٻ�D�ȓA����яĘt �U�Uc�:Z$����:T�а��޾?Ղ+���6W��TZ���C!PS4iR�^�����ȓVad Ⳮ�	%���5�˾Cc���ȓz�F��`��
\�oǠงȓ!���0k׷b������݁eB��ȓ�d@է�VĜ���λN�Pq�ȓ)5�s��*j�Tېƚ:jD�t��C�IA�0zf��rU�L�rZ�|�ȓXy��!�;B2j��S%�?Tie��&RTQ�fKn��Qg�7O_}��%�>�C(Z(�XuL�
v{ZX�ȓK�|� ��1n�0�iC�LV��ȓz�;���pϖ��D�a�ȓ?��y�s�"q>"�yv�KZ,9��@т=!�@�������q็ȓZ?�!�uǀJ��X��&^p3�ȓ5�}�� a�Ń�Ij0��MR6��%ČSlH�� j��i��|Y@,Eft-�aQ6�>}�ȓmɤ���c�'��=�q<�<�ȓ�9[�(�+� 2�	1
d����83慈E��7B�m�d�22�����5ΰ� ��A�P#
O7� ���$��<Z�Wk�b�@0�Y�6k�܄�F�P�
~:�I##�(Yq���ȓm����f��m�Ht��ƌ�@�2������g�ַ!p���ǥP�:�(-��BRj��$\�7��9�MY�LK,��v�d�SwmH�s0Ґ�v��aR$��N�"�a'm��7-Z`�A��?DzB�ɤTy��I���->��y�lA�/n�B�I�nK���G��:U�La���]<C�	�{N���K�?#(<)�萧w9�B�ɑ9 X���Ǝ0��a���Bj�B�	�d�F�@�o�l��%`b��B�I�a:r�c�k�+��-(P,�f8�B䉼=�����x#���fԶW��B�	7L`�M���W+T�xᨳ+�j��B�ɹ`��$�U�ۓH�)6!G+f�ZB䉽g2lY���"�"Q��㊈3�HB�I#L�hP�#��2�ElH:T�NB�$mERI��-	j2�����Ĺ<�LB�ɗ�~��`(Z���0N�6��`�'�L��G
��t���u��tX�'ހP��H�[����@��h�lm�'���wÉQ�i��?_���[�'-Ly����n�|0��@��5
	�'e�5�R0P�T��"�25�2��'�l
�_<#���n91��l��'���&�
<F��V+=�8,{�' �|*t���S��-s��� fƴ���'�N��6��l�a�&m�3t�jl�
�'}<)T��;a��{�Z�Z�pI��'�,��m���V���e�j�'`�x�  �$��a���
[�.��'�Vu���I�b�H�BQ�_	Z*a��'<���t�Z�A��2!
����'�(�cثp�"xPcS��Ԑ��'�v4#C+禙ز�AK�A��� Bm��@�=��ةV�P�Z�����"O&�"���a�|<�@ͷA����"ONA��NH>�y$c�p3F��f"O��'��!�B�����wD�z#"O� �@U,
>�33�O���0"O��j���H�ް�a`F(y���"O�����@�p�*	���>��т"O��ۇH58t��@3w����"O�+%�п4o���2O�0�\�Z�"ON�zwG��w����-�.H�쨋�"O6	���
k��5���Z$QB��"ON�#��	2K׌ ���L��|���"Ou���B'{ƪ �M<3��R"Oz�K��
l��a�G�K�"O�����]�^�)��#'��q"O��q�͛�Px#PG��Y]"�G"O,�Q�N�'je���.1��g"O��8�p:��ڲLt�チϸs!���@E��e�?-JB�f'o�!�$��k�!8ݩd��Z�\�!�D�-XO,5r���Y0�y�@�l�!򤞹k25���Х`ݐm9��"B�!��4+�8h�&^�*�0f���!�J(H����Ą�G��M!F9U�!�dW�i��,�7mB�Z➽��-�9�!�D��h���E�N�8Φ���ݙ#�!�$��"��9���'V�ʴ�޹v�!�d�%>�r�P5cB�J8���u!���~�8�6¬r���� �� e!�d�q#��� �B�W3rh�7�>M!�Ϗ��P�!�'6mf`U tK!��F�j���uC�����	5S,!�(,V2q��_
>���_!򤌸)��ݪ���]^�p���a�!�䎚:����\P\�vlb�!��/Dh$�mߗCx��Ta�4�!�K4��-xp�L�0(�|qQ��)e�!�ӆ��PD�߽�{W��	H�!�D�3'L�́��ɝ
K��De�!��ոMXdmi  � 0���@�L �j�!���zݔ��#�ʻB�xX5,��7_!�$_ |Ʈ]��J�;�N� ɍ�!�Dt������z��!'m�3�!�䂆G� �������#�%�9X�!�$w���Qnͤ�6���%�&�!��dp�1��!�&x��F8,�!�$�c�.��V݀v���&��V5!�W�e�.1H`h�	���Є̃I !�$ޗKR�`�J��w�N�K'!�l!򤜷5��ꤋ� �j%���C�D"!��@K�@p��VL�A���I�,!�$Ҫ�f��
�g?j�h�7�!��C˼����B�m����\�E�!��� pV��x3k��"U��^.$�!�Ĝ�V�)5o�\E:�C�Ѻ�!�$Q)��5{A#y2��
�S5!�$=] �	��-K!�	���!�Or����	�I��%B�`#|�!�ă�k*:L�"J�`�x��`�c�!�$V�r͢���)^"�Bm��Y��!�Dʔ���x4I�SR�\���ēy�!�d��9�q��Ą�t2�-���U�P�!�D�,6��Ұ흽6u�2Ύ�h�!�ET�T+@�� �*�LN u!�� �(��F� r�`�\��-��"O��!�@��$���Yؚa86"O>8�b�6D0� /���@p"O��9�(�m��8���M�!����"O�m���ӻs,�5�5�y��3�	���+%��<u�)�&�$���)pDj� @�7qO ��9Jb4�և�X�.���4u` �O�t���1Yf�K4�	wY�����ĦpR�Y4B�8��Hɡ��@*$��_:�9q��/uf���)�M��-���I2%����O�nZ�(�O�P��+J 5N|hPBj����E�a	�O����V�{}��hj@���d��ۤ��p>�w�i��6�f�8૱	� 9��ѫWb�4N�$�a�
�M�fV�p��	qy�O��4�x����D��d�#�9t�7L=�¬/{=,<���)z��ڂ#ܨ��O��;-�`�����9��� ۓw]P�lZ�FM�5h��=A��ncC\��I�<"k�t�|��sj��S�׮r>Yk�J�d>�o:}h����ٴ�?����il� AwJ�%����-�.���'tBT�t��	<rL�Wb��DSD�3=�#=9�4Hq�֟|�U?���I��I�eA��N:H�Q�������'{04�lZJX��@��ƂLy����-սs�����b�&����$P��A����/��H�'L1#<�Æԯ-�8�e���t�Rt�!�ܷL�Q���I(e��E*5N=)����O!�fO�d��'B>�q�3�a�&��kâq"��OJY�0��O4dlڰ'N��<�����d-+�T0�� ���HQTBѴQ�Q�P���6@��m���xiv��,uq�M�t�i�7 �����X�����$�����Q��G3��1���ox���	��P�ȱ�ٷ)ab���oMƨۗݙ+�`X�h�2n�
Š'�� J瑟@����+T�V�Ru�5+�"���a��2����LX��c�'�+��h�ūN�)'`�h��Iڦ���E�E%��5��j�jy��oӪO����O�O���h�(��k��h��آ={"	��OF��d�9^^�X��/�1T�\X���y9���	��M���?�C�i�BL�q%l�z�d�<��89_f8�a�]|��MҖ�oRT�l�ɷ Gy�1�ђI�tBG�ܯC�x��A4��a�צ`��B�AF?���i��	�C��A��]*~z܅�c��7O��;XjV���̇]��DR��?%��@��cJ�OrHi`�'-��nӐ���~B1�ֆj��h�eJ�O̬TZCN:���4�"=)1$-,%n�r��93f\�v+	z8�d�شM��i��2,ߨ[F�u/��(\���'aLĚ�jy�N�D�<�O �']�aJ&LQ>��,R H���L�.Р�ru���es|PJrCϹD`KY3�q����w����t�I!0�MV�;� ���4z�6���(9�hI:`aW=cOl��6�	:'���|��5�Bp��J�澔ˁ킒��`mZ	�����O }��r��i�ZU�eIܛv�0-���ĀME@�'�b�'��P�z��N�XLX�H����~�Q�ߴJ(���|2�OD�N"<�ik�OR;;�A��!��9�$�&����	K� ��   ?   Ĵ���	��Z�:ti�-���3��H��R�
O�ظ2�x�I[#��y�4g�Բ �I�n-s�E�_�]	p7m�䦕��4E�� ��q�	x8�Ļ��My�֠�B��H(�Qy��7U�#<Q�
~ӨP(&m�r��xp@DB4F��r5X�T�$�����1?�E���/��7�f}2*,�1��l�?)��0��0L־�iP��uy�`�OvԚ6F� ��9O��@qJ��0~
�rt�
[bZ���(��L�@���'�,��$�ȄyQ#��!Ӹ'=�TΓ�|�YՌQ�����fn��hJ�$�<�ቭ!�'���#1���{�L:�I�h$�'�Ex��|�'�!�f�N	^PH�$$��}��-��&#<���>��I˟R��X�H>C���w�Y�D���O(��{��]�Jr؉[�B��K1�=S�,�MSV�1���"<���	��pˀ�8���(��[�HI�>q�	)?n��B�9Bw��2b^�H�����<�fȕ'5��Fx"��N��|� �%�L��t��'	��F'|�1 �?�@�"<	(�O�e(����.��L8��Ev�����$Z��O�D�O<q�	�W�؜1�O�"
�j$�wL]?y�3(o&�O����*�1	�D���N`!GK5F���l~.��>(��4w��	�/^5� �O�h�q�סe�8��F.[e�0�X����M b�\c�0�'�ǁG�'�b�S�������$�C�2��ۨO�����d[3�OL���LR&����f��0��:F"OL�y��  �~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J }�<�u��i*�b��ϸg�.!�'|�<�� ѼG��2�B�.���G�<��HM&@���I�%(�xC��Is�<A�̀?��\ a�)R�
|��k�<Q�,
2CCv���V�/�H��iM�<�r���0N���*ʙP�{�HBd�<1�-�><p��Zv�ޕ{�|%
�a�<���g���f�1P�$�Ǉ�[�<6���EY��j�^�4�h�y��|�<���8�቉�Q�M��	�`�<��'ӿo:QS�	�|�35K<T��Ң�չr�D��#�i�z�`��?D�X�ʣ	��=���\�<}�b�=D��jD9W��B$�N-`�&��!A=D�\j'�B�"�AhvL	= �Y�ь9D�9�"�.]��3u�L������<D��*�X��DI���9eʌ��Q�%D���S�2�H�@��\���(���7D�컦�R�*�Z5�s(�>Y[f���"D�� �Yuo[�I3������Q0�"O�\"�k	�C����D[l����"O���ĥ3�� r�E�>!�J�"O��2��<7Qv�!�MS+t�t��"O^u�E��'i�� #G�1��T�1D�0zē�zx ͜#�����;D�� ��H�8��cͯB� D�T*4D�T&'�R+���L�
�����3D�p��M'T|覇	�PnDiai'D��I�M��3�deꅉ%u\\z��&D�X[��Z�PQkwc��/���/1D���6��x�R�7%���gM:D��(��䐭4a�
Y�pM�0�;D���uM�G���C�P$XnA�� ;D���D(#F�PA��L:�^11..D���F�#�R���	S���q���-D�l��͊U^PD�g�΅R�R���!+D�d���	k&�TB��xB ]S��(D������)=p`T�ۮ���{�9D��ґ[�W1*[�N�&��Lh�	;D�T���\/3�֘P�I�V"p�kӨ$D��bn�<Ry����p�d��2e"D�bs�ǀ>钄peg\?P���=D�lX𡛢�n�i$J]z"A{�):D� �K�m��%x�\�0�EJ&=D��dΠ�.��,(X�2!+:D� 8���E����(J�M�e8D���o[�XK�a�!��d��,IC4D��{PFM,�B��I����>D�h�LY�G��p�%`�Je@a2R�;D���7��w>���ȵs��tZ�9D���#A�u�����4OQ��Xr�*D����� ��̐�LC�#�l� U�)D�H[B
ϛK����F�B�8�����%D��+s���3��8�P����#D�8��
1
�d�S�&`*0�&D�@�1d͜6\ddZ�]:��K��$D���@��شa�C���"cm/D�(���ڌ~��uPF��w�`L�3m#D�Dp�+���eek�+�H�b�%D�����{�v@�c��
(�S�J(D�XD#+_�5���H s��U��)D�Ѓ�B�&��UHH���H�
+D�P��/U�h�]���!x�x��N)D�8�&@ל��#j	Y��t��G)D�$+2a��M��`Q�F�
HDM+V)-D��8�
]�ZM�$'F'�;�o�<i7�V���S�,�u8�KAT�<Y��rt�1��L�\Y���J�<	ai��<t�T"�ŌA�����AI�<�*�,�����+�&8q!a�<�։R#�N]`�FL.�(� B�A�<94BK�2��R�	�"��1��B�<A� `d,h
�D<Y4��5��U�<�E�/y��5��2Y�r�!2�FO�<���F��ʆJ�t��w�E�<�t�X�\������*P"���Az�<	�n�/mT0����UZ,����m�<Qu���e��4���,B�KVh�<ѵ�<a n��0���A�˞f�<)wÏ.$b�hD7I���a�e�K�<U�#��@!�Y52�0đRoJ@�<����:��[2H$0�"�<9$�ϻi:�Q�ðlr	$C`�<� �K$jS0S��t��NX�@
�"OP8�f)x{��;�
�:y�����"O��T�8M��5��DD ��"OzD8aM��hb���7hD0V;���"O|�P�GB�x `��R�74��I�"OLL�`����aE/K4X��"O�r��rh�E��"�n�p�v"O�l�T�M!^耽a��6+ap�"OR�zp�e�f�'�̭tT@5�"O��uk�,nu���E"U����"O`�2��D����u���@iX��"O��A�O��h���d��s�"O�á�Ϲlid��ōVd�Y��"O�%*�ƥ}XVl���m�h�4"OD-a�K�	p�H{��U�IW�Q��"O���t�v� =��G��@ac"O����ڟx�%,���F�P2"OF0�dNR�Y�$ՋWj� fF��"O� Qd�!]�x�@jM�~1č#q"O�t�@)��f��Y"�$�P�"O4�L�2��AUCܢa��yA"O
y@c� (TZ�����@T��W"O�P���݁w;����Ļ94b��"O���Q �Xd�CQ�F�
/�AJ�"O`�0�d?nB�D����\� ��F"O�IreEϛ'���I�X�"O��R�,U�fe�$� 0BY�"O0�������Z%a�$ɑ21��r�"On �Ef�`c�$�P×�M.*�1U"O<u#E�\�~(9"�m8�Z�"O�$��m	xb�h�![	=v��"O���G���nĠv���~ZM�S"O^}�4��%k28�F�VV��V"O2�+�F
�)�0|R��g�����"O�a�Jϒ:���+ۏ(��ԃE"O�����D�Ĥɏ�{`�@�"O�8#�O�b;48�m��lG� ��"O���5��/�
�R�=(A��ؗ"Oh�� �Z�x �$Y�a�2Rz��"O�x$�0�� i��A�P ��P"Ob�"쏬$��W��U0�:E"Ou�a�Ki�4�����)?&H5ʇ"O6|��B�8k�Qx@�8k�>}�'"O�Ik� ,��q���ǹ!{$��P*O�gCҥc8���$Z�G-b<��'���Q����A�h-�`J	4{�m�'�DLC��BB-�*�7�x=��'b�s��-M7
��V�ʛ)��p��'	fU$�0F�9
F@��m����'֔����&W����	F��@�p�'�$���C�"�<E1�kX�}����'ب�(W�&q�е0�/�z���b�'8�!��]����$�:��8;�'�LSF�(m�N���
%5�����'�P�C��,j�^e��.a(]Q�'B���#�N(�Y��*P�\(-��'/�\��>w� �!�JC�SՐ�!	�' �Cb%X<����*�I\K�N�<I��[�j���Hۇ/��HX��p�<1�h܎I��u¦�#7�[]f�<i2���V�uA@��9f|�3"��z�<a��o���"��0>v�dk�e�p�<	� 'H��%�r'BVE;�k�o�<A������!R�əs?�h��b�s�<�  yd���<�k��>�^���"OH ��H�p�l	[JBf�8��"O<e�P�+GB�`/��� �"O���gf�Y���vn�t��`a�"O )�m�t6��P�Ix��a"O����"ьi��=�&��[6c�"O�hb���	
��$��a�M�"O,��墆(��)򍀶�j�#"O<ܸ��[-(�.8��	O�h���"OL��v�A&c�F\s��+�r�hb"O�x��2��,X5̖�}�BѢ""O���T,x��h�j*J���q�"O<���䀧j�A��hn}x�"O����I%U\ait&�D+h��s"O�|���20t]"���(+�e��"O����E�:�򈠃'�1B�Q��"O,H�aឨE�hH��R1f�H�"OK��ƈ�a��~-��z�"O�����@-ޜ��p��9��"O�)� �#Z�ּ0���e�ó"O �#tC	6$�2�ˇ��9=d�Y�"O>5)f��Ia:.�M2n܀"O�L��U*����MH����(�"O�����=�t�b�� t�`<��"O��w��z�6i�1k	_�J��s"O��A�H�*q�|� �M�M��4��"O�hZ�X"D(@�Q�_Ev�x��"O��e��4,,0q+�/eYN|9��IFX��Z�J���(7��� !�6~!�D��M��y���&
�����������(��x��3p��c�D؛d5���"O܀9�㐮G�y˵Q=5����=O���d�=?�(-��&	�uy��Wk��y�N�<�U��$K$�|��PX�#@�9�j%��+iW����G0%���/x�X���$�G	�uoZr≅	�Q���t�4�O��+nÏ&�X����]l�<�%�2�D��L��f٣���\�'axbT�'P��i�aoXU��@	��hO>���	�a~@D�ԥH�L�86:{!�$W�`.V��pd���MR�d�V_��)�'G��[��C,�(p��A�^��
�'h���1BӸ#2���m�=r�����N?a���Op�qȃ!(���Ő2K�MbDG$D�LJ�%'v�Ti2��62�5ӷcߤ��Dv����+�4���T�*����`#72��C㉙d8��Q'ǁJu�IR��S�t��	�ȓ���i�bA?jt��Adhԕ\���ȓ��pp���	-$ر
�Y���	A̓jFD�y'#B%�}�P�sE���?����~Jd�V�RMx�0?6-@pnWo�-F�<�|�@hO{S�}�Ʀ�k�V<rcll�<ѥ��P�L���ς
x@�
��@ܓ��'p���])��R�r�$�sG"�G�<=;"O��(S��x�q �"1���Y���?�S��1�D4*C9o�T�B��5��B�I�,��I#�Q�[���w�e��B�I��t�A�e��Y� ��nB�!Xq*�'�U�n��y���Nx�B�ɟp벸��@_�8��;��O-"N@C�I���u��/R\I����P�C�ɰ/�v��$�F(�ɱ��#SX�C��)�Ѫ�m	N�g,Ψ�C�	<f��t�7�P�DM�! �?wZB�I�X�R��BI�)a4!ZPCB]iDB�)� �M�"Р47�$�ƭ̎.��3"Ob��1C��a��Uh�ZW���"ORP��mi���Fm��*=L�q"Ob��D)�419�����ބz%�[��',qO� �6l���҉���,�1��"O�����د����)�4Z���"O�����"f2���;Ƞ(xr"O�ٔ��0QmF䓔�¨w |�Yq"O��D�ЏW�](���9t�C"OH3tg]��h��#GĝZ"��G6O6��D�dnLy��I�[jP����iX!�䂳-�D�т8J9�yZ5���!�"R��%ѥ��(~�*݊�cM5u�1O�7�.�S�'\0�jV�D�r����F����	O���Y~�Thn@1�T� �Ż[�D=�O�p�7J��u��0�G
�k�����Ic쓣�'L�X�Cue���I�E��D��Q��?��;�Ζ��{��~�T��yTdL'M�8R��=�wm�Z��ȓ�,x8#�����@!5��	pj�ȓB_*5���6%~���Ю���ȓG� (;��6в�9f�)a��T��U�������1�Phi�H?+q$ ���K���#P��ز����+>���+_"O�,C�Î.��0��!�!����"OB� H�&Nl�@o�~�
)Ҁ"O�"׌·8��xH�.� W� ;@X�L�'�\�FyJ~Bt��P1��e~(z��Fn�u8�$�a���*���Bq��mϛl.����5���<1�@� ,�Pr ű8>���Yr�'��aG���0D���k�N� Iy6<�N0����'�����J��T���^�D�s�'�ў�}�s�
	�0��6.��ѱ�`t�<�d̩a� %�1G�08.2���y�Ud<�<��������0��oҙ%�бY�P�E�!��`A_���pG�F��@��	,��SЋ��G?���r�[�|��U��ɺ-���D;��V�8 S��qՄ�B�D�n�qO!aӓ>�|�COֲ
T#�s� �Fx��?�lZ�wk��A��Ҁ,����NO�RC��("&yA ���a8&]RTO�b�����5JY���7�Z)��l�:�!�$[�!�(��G�K�
�%ǘIQ!�dǅ.���� N)	� aK��!�d�#U}t�&fSy"�}��7k�Op(
�H5 ���i��+�^<@��ĽN�����N�x�	��̴N�&A볅H$U������`�K㒘����=3�����eW:jO���I{N�O\x�EkԴ�6���E]�Fx�"O�E�-�d;��6Fڝi�
 ��"O�t@����ie�lA�z;�Ź��'��'���	�i��Q�µ�Q��7"�@Ղ��d9,O�������2�L���l�<5z��Q"O�i0��a5J�F�-"Oh��V�ԉ3	�icꐕ���H��'j���6�,E�Ay�knQ�a�"�.D�y ��F�%cӕ-���9��?�S�'`>D�T�-_�Va�7�^�w0�X�ȓ?lpْ�"�)Ä�6��|'���I��0=��	�����#�1���B� �p�'5�y�E@;? d��LU��$暭�yB��F<��C�k��5���K�.O��p<y����'Քx�dN�?]u18��F�Z!��Mʾ�A�#�7dX���ӊm�!�� ��.1���㧃S�.\��'E��x@���?N��i�.��0�p�Ə+D��!f�eqpA�r-�F�TpzV�	V~�2O��)��<��J��,�]����0Mkj8���]N�<a�l	1K�8Pyf��)����4d�F�'A�x�aU�6gvoK�H��qWb��y⩚;����D5>;��������yRȊ8��qBk�;���Ea��yR��]�d����!g��icm�)�y¡U4�`ɉ�S��ј+�&���3�S���>!A!��G�^�	ӄ�'&|z]��R�<Q�H*& TH�BE�S3�1T#�N�"�M#�'�qO��p���٘� �y�54v�H���7����z���':�|X���X��hO���Dŋ�XpG߇V]��Є�B�Z�ay�I�1�)�R���Q�P�˵8	�C䉫J}��3cΔGx�ؔ��)M~#=��0BI"Т��h�N�P�	�z��G�D�FbĹI-�p��`Pn��lE�'^�?7��:� �L]�&���K0d�8/!��T�H�����V���!�)i.�d@��(O?��v* Q�fՉ�&P"!]n$YB)8���*�BPl�0u��ˣ��)1v���[����=�'`ȹ7�
�t��8sft��BO�<q$�0�PUK��>F�lX��ZO�<�'�԰$� Y֎E:��y��kVL�<��㆏J0��!.y��(��H�<a�f](�0[G,�-PT4���@�<A1���\�!� �=/d���梁c����'�
ȣ�* A�6�=��pP�'*i#n�$n�xA�̆'� �'�޴�5⛜�R0ɑ�5�T y�';�5�����t� �H�>Zz�� �'�	��HO�no���@!D�a4n��'Hؑ�������0%[�F'N@y�'��@2D�[y�(s`*�7[���	�'▉qTO�H�Hڀ�]e��	�'�(�;7�������(`���'�J]IA��tmȘ��G�8ʁ�
�';LR��
>_�\��)�$/$��	�'mnh�!T@���T"����I�'���c-��H��΀��R�H	�'����ʕ�r�ģ�+5� ��'5�]��!�@�fq4@�,4�0 ;�'���j)SK�Q�`8� c�<�P)նI�.!��B�8�����\�<���O<�>M��Z�P�>m�djU�<9�$Ϙ~$&�Hb���M+ē#�>C�%t(�H�AL�>�J�Ͼuc:C�	2<�xx:g�O�b��h��e�*C�!8��5
h�".V�IwE �[�C�I�O�����Ō^�l�2��ڄC�ɁV�v� '��,����B9i�4B�?��3��վ;"R�)��0v=rB�I?��Jiћ0W"Y�w���C�ɶ;W��iV��h�$Я��B�I�'���1�NX>JBF�RI�S��B�I�ܱ��C^u hi,�	BB�IW�L����5�,�96�3��C�Ɏ}B:|B��,�P�pk�j`�C�ɰi���s�D1&0��ia��)��C�IKFY��259��a��z�C�I 0���F�1��8����p�R���˻{��Q�h�-J <��W'T.LLb1�'Ԙz�!�� ��k!*��|���ԍ�H���"O� ��A5]sr`�E�'�&�r�"O�`X`�I%Q�0���,a�Ay�"OR	��NB	o/�����3b�F��"O��S�(�NP6   qk���#�"O���EI
�* �k��%N��	�f"O���E�l�0��<8�vT��"O~X��ͮ,�����As�q�5"O���u"ƈ&���F坂��q3"OF�ICn�@�`h�*!(逼yq"Olm2�/��P�r��.�Bya�"OZ9�����B���G�H`�"Ov��O�6T&ڀ�=���d"O�3`M�w6jhr�V3�� �"O ���#e/����ʕu�` ��"O����)y���"T�*� Z"O�E���@+r(�T��dߟy�tD�&"O���&ZV�E�R�[�F�
�'���'JQW��a�f,^x���'^X�mA�J�����F���݆ʓamH%	6fA8��3��Ӆ�N���giv��pcR�1E��+�a��^\�x���U��O�,hCUOɊFr�1c"O
x�נڊe�e!#�_�|+Txp�"O����3�m Tl�{x�!��"O
� �
�o+$�m �!f(�Z"O�|S�#d��4r�'�;H>IxB"O����J�~�:4�7�ʨS9н9u"O:��ɕ�g�2}ysFNH�"�"Ol���*�r���F��".h�0D"O�!�F�Cs��qᱥ��f���"OB�Z���	�qz ��[��u�A"O��A��U�Va�U�\�k ܑ�"O
����&l�hrG�R�N�8�"O.���!j�����3>����u"O~8��.ě9w\a�6���s`"Oʁ�SÚ=�FQ��Ѝcڈɚ"O��sqV�M��Y��ǰ(˘�h2"O>���52�>!RU��!�,u�6"Or雂k
6:�~Hq@ķ�nU��"O���eZ#v?�}�� [7�X��"O
Hv�J�`�u�fN�aif@��"O�A���*C��#Ql^�A6~�"O�A@υ�	�Ƞ0׫ߐ9�&�s�"O����b~�%+Pi�X~�1W�')�����,I�'J�10�nh ޼H�ǐ/ �|1��'�r`�#M̩A�Xz�EN*8�eK�O�%���Vx��N�"|
�$�Z��W�0��c�m�<��o@jјr
�7^���Qc�:dtU�'�l��fY�ϸ'w�dstaՠDwr|�J��e���{��6s�D#�cՐ�x�����T�I�;.2B%ٱN��0?��ދY��I�'[�*���K�'-lA8� $�xIH�?��G���:p���Ѩv���Q�-D�L���ˊG�0@�7ɏ<}f�����<�P�^&9� ��'�0|ʔn C�>%1�DjNj\�pB|B�	�K-�mI¨��L��D`��y!l�����<!���v���M~�=	ƖD�D0�!�U�Գ'�e��P*v�O���ȑ\�Bv�U|�DY�Ȁ���9os�d�$��/P����`�� ���?I��u�N�b��1��Iʇ����&��e5U#���~!��Y0(������;*�ɛ�j�1ly��?s^��g�Չb��S�ϥ�ϧ3���8&`Ԯ Y�H���^�<�c�:9�f9���إkFT��'i�:�'GP��)[�g�g�d}��T���+d�!N<�B�)� ���⃷T�)k�+� �6��s"O�i��%�|�Ǡ��8ɑ�"O&�S��ܖ%�0�"��. ��!"O"Yx^
��M��o>,���y�e�����GJ�d^Ա���:CZr�(�{�(a���Ğ�s&P���C��a�j��{!��J%#6@Ka��Y�`%��_-=`�\"�C�$(����"8�iBbI�	�~�0�S�cV�x䉉$�*���-Np��"~
��r���JP�E�B��5b?�C�	 EP�Ѳe�_3��c�#��;�nDKUƗ"L��"��ob�C!ɇ�"2~Q�A�O=(�zC�	�����U|-~��g�ͰB|��A�)�~��?i�	�S���{�IښrZj<��G�'f� �"�=��?��ژw�`��Ϝ� B�a�#E���ǀ�h��Q�P`$�Oq����Q�6�����$:̸��	
xuPɺ`��8h���V?-آ`=vU8����6�rͰ!+3D��r��%s�����١���v�`y�GĔ"�UKjZs�^�D��oV:f(����!1�t9�B��yr��5y�%��͋(HX؈�+Z`E���=޾��`�.���(��y�#=��F�2a��T��E,��;�n�~؞��(��}c�	˧A�>0���6,ݹR���s��^�k�l����<i�؍;��'[������~0f ����T7h�{R�E�	���-�4�T�A�Ѕ�X��OD��,�<�����7@��qz�'�ډrW�J�6JyQ�# ��l����*r͠�y#���9�J��=�(�h���@���J򔭑��R�5쮍��s^�b�$��oL���B$�9���EQ*SAܨ�$؛/F��3!H?s\�>�cӽ8��`�)�3h!�B��xbE�͆].8��W�N�naH��ۖJ�bS��"K㐁RQ�����}���rP]�B_�4��e��V6żd�=�'��dR�5�ӪB�`�n�)n�	~��G3��"�Ȅ�9�T�0"DQ�Ն��	Ó�о�&LKB�$Ht�b��28� ��`�B�"�"h��Wm�O|�	�Wj�0Id'�aZ�-AQ�ĩb��C�ɔv�*8�%�ٶ#���(D�$�PI7_��}"���9�V�)�A�v�R*Y7! ��&��C��C�J螜�ħ/eL�B�-lO������kY*�1�@WHm>��e�
�v��ibEψ�Ge�<�$f�9]��6��1O���҈,,O�<(e)"Y�X)p��-���
��'QR�2���U?qu&�(Fa�]�PC�Dђ���Y(^��E
¬�K̭WV*A!:)�Vh��C�P����*[_��%�E��yP��`��	-@(�H�H���0Au\��2(�/D,�t�C�	
3Q��X�k�0{N<
TI��zz�|�h$"������%e�H��2MĀTLF�)��D'F�PyV��,�J$(�E�QlFlZDN�T�'RiB�'��<K��ΰJd�����'<�4���Ð*��6α˸Oj�5��H�>2]��Z�@��TԀT�Սڿ��3õiI�Uj�/��Y���*U+H�� ъWd�c�](>y��B�bĨl
�� 6}�O��P�៌����)S'\Xڃ�E
(�^�; MU�z����Y$?���Y�1�T�5	�E��d���T7���B-2B`���C�y��0�rS��a�4��%y��H�i�y@«�m�����'T�}�d�$hN���2ǌ�g� �`B*`nV���D�<9!Ƌ6>�:�&%}��)�����[��\�U�x�5Y�Q�X�)����{��ӔB�������Q0�5{U�čm��2�l�;V�M������F�����P�R���˲"��0�0�;1d;O�;��>�BA��O�D Y�,�C�Y!���ls��H�0w�`C�	��1�UB�)r&�4e9Z��Z�X�cA� ���G�w	hŲ��*��O9��%����݂��٪Q*�u�
�Q(�}��#m�|<��e� �Y�'?z�Ͱ5�'Y�ఁ[�D~ O?a�$��>l�A�u�0L���b�G�<i�(،+�$��Ƣ�P�Ը1�cU~}2!���L�R��'U@��T`�<`�`I@4&o,Ip� Ӓ��T!ݔ�8h��� ����>�:pA:D�LC���;4���������a�<	rC�=,�ć4[��D�� ����X�a�.Yo��!���<�&yK�"O���-�.)�H�j�E=B��@i&�X;�V��Ʌ-%�V�;Ċ��g��XO�c�,q
1�Pa�	�07�ة��1�O�ܹסу�8� �{���h
e�:��@�>	����7nJ��N�h�3LO�9�s�!O���ٕ�y���	.!���#�&S����p�L?��b�,��� ��aPE+���Ó"�Px�Q"O�p��$p�񚦥\�r^�xz��i߲�Tnߡ]Ժ��NK�Nk��D�3J��c?�X�{~XH �KŬbF؉�bH��B�I�Ux�Ǐ7Qp���\�f]B�2� фTx�xSŇ�ZFڵS���?��c��+?1On8����<[��� a�*`��ag�'��mK獜/�M��&4I��y+ç�DA�m�cD̓~c,X�di�0y�]`4$8\O�姝��bͺ�G\7<��<aቒ&Ϩ���ιP�����I9l{%i�l�>�uǤ�"u�i�7`��N|�)�v��y�ݿh|0��A��@j�0I��ܵ^��������aJ�p��M��s����C�o���B�Ҩ �:�f.D�P��K؆+}�B�"P�G��53Ճ̈́\��m���^)p'�4*\�V7��F�'��I��ޗ�<��i�uB�N��+"��}ꜜ
�����J*0[�h t�%x�4)��$m����I)*����]�y���5`L	F��#<!��>Q
x���ʸ*�,)�e� ��	A�@,$����2g=�ՈX�G�!��ف@; P �!ܷA��Y��g��r��(����M{��7[r�׈Y�A9$T�~λ3*��	�3whQ�S�D����	M�u�28O �5�@�wR� pC�ȏy�J�QG@^� �I'%H�3m���g�Ńr��vW�<0�{�Ǌʪ0(宀� ��kբہ�OX|��Ȏ#��G�R���L!V�r�я�D���]�oR �&��.@�p�ěs+���� %LO<�(wŜu	���e*ъ&>pBe���q�^�i�`Ky�I�?�g\�$*j�j���
�D5�"\!6���B 猞9"y�I՘b4��ȓ����MI
�X��˛Y�j�o�2] �������uYcۏq+��ۑ
�]�P?Z�_xu��#M�c�����#L��{B�L]�����æ�� ��7	�-��k�����a�
���s �?q�d��̏+��'ݐ䡣��֧z���J3JCk�1*EfKd��O�xQ �\�I�,��M����`Y:Y��UZ�%\�6/�)��c�0�>�q+��W_��@����6�)QsJSZ���1�b0�|j��G4&��Á��/��A�#����ɷ]6��slFN����F��q2�U�㚾w�T�e&�Jn�X&�86���ȓYj:S%�ɵ*3Z�АB9����	0W��p�ԍ� ���=Zm4C��/9J���T���ZH�#�/�����M�;��=a�Ocݪ�v�z�ޠ�#�[(��!8�g,R�H��ʍ�9w���7(���)��<�Qz4@��K@`��r@��k�'�)QuhW6%��>͛�;O�ҵ"B�/j�>���|���c|U��W4��y�e����ғ˜�'�b�p��F9:M�(�=E��,�� �N�s��dQg���?8���ȓ�~uy��ݾ-�$m��Oƨ&�9�ȓ���{��o�&8	�)F�M�x��ȓc@ʵ�P��C|��1�+-�@��ȓ`�x���Su�dhT�R�q��Ԇ�sc�`����Cg�YC�x�ȓ3����/J�@%�T&z(4���o0��Y �Ę(M���B(����]�Ҁ��S�n��~��mh�#�e�<"(YĒ���ԧK�$���[]�<y�,A���B�h�:#	��.W^�<�$�j�,��l˨�p�)�+Br�<�uJY��8ت�*E��!��Im�<Id�*Q�� _&-�$UЅ�n�<y7	��JD��:�� Q�"A\�<�� �%�j�Q�� <��I���\�<Y��ڦK���e�iq���Tf�D�<��AV	P�dH!����A7)C�<��!�v���s�+��"��7���y��P�`��i�Bh��a^�{�
!�y���y*��05j4�tĐQd�9�y�*L�VY�Fɛ7*��Q�T8�yrm,�5H�Ȟ�)��%"�b�$�yc�%O��p��k�|� ī�JL�<���7f^LQS�YT�r�X�/DM�<ɠ�Ru8�9��b46R0XT�D�<	����T�hѲǃO�9�%qe��@�<�s�Kg�Vђ�g��X`�8a��<�&ƛ�,L���11���@2&�z�<� XQ�
Ʋ'�3��H$L9Q"O~�vo��D��*®Y^�8�"O����X�2& p�m��M
t)�"O � �훣m�H{���o���!�"O�Q���T&V_��b�HS/ɚh 4"O�Q��Zh����'Fֻn�l�:�"O�D���-�A蔥�J���"OX�J�V|,�$
R�6�6�b�"O┛��\&y��#B
��d��ܘw"O�q���%
��3&��w��+�"O�@
���]x(�P�hP�Gb��H�"O��������h�G��A7F��G"O&ՈEzT� (]%�䋥"Ox�c�BאZX�a��J�(�I��"O��A��Y�}a8��A&ܔ_ ��(�"O̵�v���q&�(ivG�����"O��$*��z��31C��1��-�"O�	�Gn�%QC@d�"/�nQd�V"O0 ����\�l -5?�f�c�"OB��u��Ka�Q3'�7E�~xk�"OP�v�[70��rH����uX�"O���bE���X1f�S�{�`�"O =Q��C�N){歉�PҢ�5"O@�Q���<��܊fL�E-R�A3"O���C>
��`@j9_���3"O�t{sʉ	lXl9�iU�G��Hac"O0(p�K΃-7�����	H�.�r�"O�p��3qF���ǫH�@�PiA "O��S�H3*p^s�]:q^A�"Ofڰ
��X��yPB�$ɫ�"O�[�L(v��p3�Ĵ���cC"O.hq�$T<��C�C	=�,{�"Ov�p�U�L�$}Э�0C��Ka"Of���G�&�R��C�>� ۆ"O���0G�g����'��~�<q�"On��pd��@��ЮE�R�iS"Op�S�GB�}q��z�h��%�n$��"O���`P������?ZٶI0"O,`�[(y��A��r��"O�)��'Zp��qWA���5r�"O�ҡ���<�Dh@%!I���g"O��q�.X*|�J"WF <a���4"O�p�HΒZa��Z��[H��m�"O�l;�A������+V�2���"O�<�p���MΘ��1�ʱv8����"O�|����O�$����H�(�	��"O촓p�×
���K��Y5*�T�R"O`L��	��;�r�ه(�2��b�"O���֫-s�U�D�*������'����w�R��'�~H��
��D1��`C�֋O��H�
�'Լ�
u�Jq�)�kفU����O>,s��3��)@O�"|�4�0<�L2wjݒ
R]z�'�X�<a�g*s�)ѣ�!ZL�=�7�%x⥖'�l%��h�ke�ϸ'�0y�ǖ��[(ɱ<����
��-�<Y����1c��dK�����4Ӄ��^EJ5c��L��0?i�-�"S�"�Ζ""9��9O��6��y�<)q�("��Q/d�&%��k�%V�Ls1�s�<q&"cH0槗+E����el�Pyb`X�[�
�R�KV07Aa����fpx4�
�	[���b`��y"��<J(3sJ5��-�����s(OP�l�5n��qO4aW���$!"�O[�Z��}���',!�!P��@����q�H�Q�����:`	UH�a~∑� ��p#%<`
]����?��O���"M#��9 T�.U�J%5���SB®8�F�Q%�h�<� �	x�EةG,�#��1�p10#�� H��F�=gd�rp�>E���N=Ux���d\�S5K ��y�A3]�VYc�@)]�ϊ5�O�4�
����NT�
�'�>����7G��^�p4�ȓ8�����&�p4�@�U�26 �ȓ&��p�۩d�l⥫��-�`��,�*\��`ϣ<~�8
�㚎+�&E�ȓ9�2u�K�<����g��A�܅�f1�!H��̿9KXP�A�[踹q6�^Bܓt�آ|�'�N����
r��#u�S�y�z��
�'�T Ae�
\�D�����t�" �uՁQL��U�'�Z@ �#��.�0�h� `��{�LL�l@ #P"F��eH�O�d���@%gT0[RFț'-|h2"O��Z�L�f�=�H٘_
���w��`k��ѳ2�  C/��ȟ���m�H�D)��e�4@��-�4"OV�+C ]>A���K1(���zD��7�=�0Z�Y1��V!��g�y�PĀF�%!�xD�t`ì������/{�@�8Հ����@�gS�aY��ju������`�'�*�BG�N+H��V�Æ'-P����D] 9�8�:P�Y�	��P��N��TDˌOp�ḗm�-a9��ђ"O0���5Ģ�1�Κ)@�҇U���F�=g�P�J��?}3"�RnhjX���	C�h##�&D����T� �� �ѣZ)c�Z��f�);gB�
��=��
�.��k\ ��ԑ�HOL�[u�H<U��'L�3��	�'��Y�3���"@�x7��V�� J[�d	��k��B���8�IPr����I�����jV�$�F�:p�̲@v����#�fI��-/T��9�g*T�:d��G&(��6l��ebD�1�f���C�I�4(ād(��8���s�E��CK���{� C�8v� �!=ʧ�����*�b�@Q�σT���⋏t�!�$��V̌��4�D��2�𡂪 ���H��I;O�X�ѧ��� ��Q�h�F}� �4�.9CcN��@���7+���p=����,���r�m�����Q�^K����	��:Y����OC{�-ɕ�'�y�!!��QT�F�:�k7	����'ީ���ڿ�6ɀ��Q*���.��'8ȳ�bE(90bp�R(t�����+�=Yv��O/&]����jl܁�Z�aq`Y꤂R�z��ؑ��y�On���	V���3�n�L���8t���mSJC�	�eITi�s��.?U��h#�7H�^�{��7>� ��S%�4�H�T�8eKO�=W��$���#�%o��w�L�K��1���>lO�I#	�?$;Zك�,L�ȼ*`�o����k56��1��	M)�h6m_�53r��1,OJ�hq�X�y�JR e�P�`@1f�'����a?�&C
1'`�1^�H�Hd ���Ő2�*"�*��;%�F����ɲNB&��I����d3��5!�@7$�B%!L��	�O4����(EF i"�
s��ʰD�!Z����U�(J{�8�q�@�Ee�T��'�Y#�'`P)�m�<p��T�ԽxD�����X҄�g�A3H9T����?=�p��|���4}��9^!�ql�c�rH��ѿ�(O�;��<V1���T���Yk��e��y
�`I�^<n�����^�^��)���۷-Cw8��Bo��-x�Afϕ�>���5E ��Xƙg�Xӧ����e�X]�	�[�D�q�/
�HrX� ��|<��'W|�"��
O�A�ƕ>�I�a�*���B�O���H��Z�0�'�¼��C����O�	
�GY���
�C�o�k��|"�E�hض�ӲE�ڔ��ci@�?���E�����?�������]��ӧ���h��U�4$���-��/ty���	�[��98 �Ԛ6&>I�Em
yu"� A�	 ��a�/?�c��.� �6O�H1Gk��s
�b�d�7�O�qg�L!�I/p�di��>����\<U��B�)S�|>BAU�ܠ_�,e�v ֐�0C�	�S�@�z�(��$��D��FƳk!��Ec�1	���$���?��9:��)��O<�
"L:v4H<ӂ�A�(
V1�Op�80����M���"zd�!��e>���HEџ$�g�N; .!�I<E��+28{��?M\� �)CH!��&\R�����&	��!�)�� R��\�$a��La��P O2~�Q'�
O~��R�(�O>U��L�@h !�xC�N'>,VEzT�B�(ÔH��ϔ(ɀ���,-�52�8[w�\GyR�M4ŀ ��T�O02�q @����Cʸt��l���� �ɪa�ƦxD�08g$�@�a�,Az\�D�qt�S��?9gI_�vq��D��l!Ca��k�<y7 � "��	
�#�����.{?A�ּN_�4��M=LOr	ĥ��,���=��j��'��\C�+��Dy9dHB�J��P��cJ.,J 5��A[�<1��1_j�([્+	���� �Y�'��qQ�3[l� G���v-"��tH#tn�Q���(�y��9-�v��Ϫ��d(0-�Z��2�א(��I�"~�	�l�f�p.�)Kn(�h�n�B䉙���T吣a�( �&�>p��*��g�� �p=�FAH.j��Q@�<���.�{x���6nE;k�VM��y��O�!HxH�Sn��y�$�'5���b�ʄ&"\���C�y�Bƍ$(ȉ9�b�&(��#B��y���2aY�K5m�W�ސ҃(��y2�=|�FU�E�����r�	&�yb�@%{�:�*�,W�@ac3��1�!�d�*m�Ä-K�m���#$���q!�DV�cL0�"�nF=��)����
7�!�DĀS&|��a�\�2�X��"��.�Q����D�R$x�E�4�֥D����-T���9)a�\��p>A��1s��	-t��x�芮�H����=Z	��R��Y
u���:!�>E��'C���s&�:�1c	-� lJ��$��Ol����,�'I]>h�0l
�fJxyw�CBE�Ɇƪ�S�dW�r"T܄鉃 �`���N�0YD0ۣl�!@�@1 ��>K��K��&?�@�GX�F�b�2p��,0��8�c@�G�D��$�=`@�,�ȓ)H��D Ů^y�b��r=�ɈBBĊ���.�X��P�а/D�xT��lyJ?P��|!��T�^|�pb��6|O�A���F#1b	@�4�D�ه�AOF�{�H1ej
�j`Uz�ԡ�Txy��D@BCڛG:�|XF"X-��A!�2�I�*�q�@�G55��>������g��M��J����9@l�O�@��ۧ|����1(9LO�%����3�.���3c˫��~N�͓6��&	����U��9��&�P�w�]� $��gQ1���C�y"��Z.�2'��GD���tÉ�?��%R+v��A��	L5�p�Pf�X(�j/O�$T�l�!�I�[(b-��[�::u���y��a�%U���I91�����B�\�^B���$ܙPM��Qc+}��9O$ ��a���S�O ,7N��	VD
<` ��Y�OlI�)J�WZ�U° �Y� ��'P.��r풆�a{�j����c��ڑR@�$PI�(��ı��_�Ƹ������-�|0c��
8�� �̇��y�ϛC�AAJ�0kX@��C [%�y2!P�# HB5��ai:I�!	��yF�T#��;�l��k�f��PF��y2M6��QF��[lv��� �;�y�N�3��H���CWQ�<Ң獚�y�N$>(MA�ԐO��x�a�á�yr埿c��Qg��&=	ԁ��iŻ�y��M5���c��D�[ъE�y��� #�jqX�&��i�zz��M�y��HW��;���1� ��Ɓ�y2@ΫQ!��h�G��I�C���y�BE:jX����*��lp��:�y�/ur�K䔿"T�ǦO �yrmN�ْQ�`F��A��C��y � 
��{��-n�X7)��!��S�I�h�P t�*��1욢'Y!��Y��� ��i��<xR�T�$�!�$*Fq��2a���UwD��#,�!򤒙Y��O�q{l)t�Ҽ	�!�d�I���Fd�R"���6�!��> �Pe���)[��bg�
9h!�еh��tH�)~D4� #E�	�!��9�@���L�D���TCK�c0!򤆲FGܴ󳋘@zlC�T�|!�� ���(9�.xJ����E���3�"O|E�:_�L+��rZ���"OШAå��L�P�gޅ��9b"Op�GO�W�f1{g(X���,�%"O�D ��x��<�5h�,O�$�Q"O�����.[�ݱug�A7RXs"Op���L��W� d2ed <-�� g�'�p��uKV6a�|��	V#����GF�j�k�'�L���Ѐ/�t�I!�Q03(\��'�H�!U�#p]DMѰm3)�h��'���g�,ԁѦ��+T�k�'���'J=�ƨZo� <[����'�����%$�A�+�!�Iz
�'��XQ����z�b��F�L�x
�'�����}��K�a��%-Rx�<9�Ƒ@"ι�v��C��ᯟ\�<9.�#z�نGĨzE, r�Z�<�Fn�6SV-E̅(i���S@ɖ]�<I�M��@Q��H檃�/D@q30�s�<ٱb�%��KX=s��)��Gg�<�"ER�9�2�C˶,r�a��,Xe�<����c��U���P��6U�OHi�j��!�'K����*G�{��y��37w`E�O��� �O���0�q����&�? �������2Ю�Qn���Z�:�(l]ر�_w����'�$})E�N�1��A�֪U+N%b�Ru� s�\4k���X�R��~�*�
Y���uMذ���q�\�.����k(]ֆ	��O���)R�7�p��t���$a��@.'� ap)�Mf��5p=y��IS�)���`����ɁD��Y�%���0, *�O�@t�ەq]����;�b�}�*M�`�� ��/2+X1��ũ�?��.�!��*���c_\������m#T�W��Ј2��h~��-��BdxQ��OA(������1�>��7��%HU���,���J �P&��q�T$�'�N@���	�|��NL�bAp� 9B�6�𮖙��'4����~��/��G*��;5$ܵA��KKU�<A��)ƀks�;QX�� ]�<I�޾#���z%,�::EB�d�t�<�@��oc��f	!JR��I\�<����%j؍b&^6@pXG�HY�<����nF��d��&~}�e"V�<�q�Z%�z���@Y�,B��h��}�<YC
��!8dY���q{�H��x�<	�BӺ0��(X��-�D9���p�<1FΌ=*�Hd�1�O6C���'Fj�<12 RM�h�E�8xGp�Cu�P�<!�'��R.�KD �1Ek�a�DN�<9��N�Q�l�DD��#e��fa�N�<�U	A�����*��)�c]o�<�t(PE?f(s���>�����li�<Q�,%h���&@��޲A˗�`�<A1�D(I8���%װ�YC%ZX�<	ģ\� �9scX<��1��Y�<���Z5�<}۲�	�<s��:�/EV�<�0 B��֩kӉĬ�4H�2�Al�<��ML^Q�C�īB�
ܩB`�`�<IV�ǈMg�<��L>7*����LZ�<y�)�7"�A���B�H	C�`�<!��ǅJp�AeI�z)��h�s�<	fІQ(��w�K.�nUH"n�k�<�$�H�����v�t@$��U�h!�ȓj��Ƀ"�·M�� �㉖7�~�ȓ79ЂGCŶ.���"A	_�h���'��y¤ 9 ��à�H�<Zd�ȓD|8�ԊO�hs�`�uE@p}��w�T�Y�gҜ_�dCpk�L�u�ȓ*�!�O� +*����R4R����S�? ~ec��<"�T�s�酒;�vy`1"O��ui� N�A��yږ`Cf"OV`�a�ӏ@3��[ȃ8����d"O��c���'!"�\(���>��\�#"OI��b��
Z��I/Ƌ�����"OFu�!�@}InhxF��=#V��"O��G�9c��!�tl	�88���"O���T��0Z��8�>�bU"Or���"
T�(�Z�J��oy>��"O�P�b���Ze���^���a"O��	�!K�IqبP�ˊaX��sC"O䌣��. |�M�WZ��
�"O r�Ҍ@N��a^�/��q1"O.�Y��1��F~��`�"OXIc�,�X�n�q�m�(&�@�T"O6�����X��|��&��0|b��"O���!�����!'G��h�8��"O�0�S�ƭR ��[�x8�"O u6R=#4@HuǓ,#��i��"O:܈��
�GfR�jRĉF�t��S"O��LG��(�"�R�e�Xl"O�|��N�^�R|�U$.���$"O�A��W�ͤ�8�H��9`"O � �I�F�~	IP!ߕ���*�"Od����F���1��]˒���"O>	je�3d�}I"h�k����"ORX��� @٤�B'�,�Xe�F"O�� Q�ؑ3��s��
�"��P��"O&�xsɥp6��(�dI!od�hI"O�l�P�l(���Wf=�w"O��J6��:6�,`³�&n�#"Ov���ĎKj�c��9jd s"Ox0VB��R2lC���7�`P�"O�@[B"�&�����ʁd���"�"O`rV�׃, ��'��pӢQ�"O��6��!ڞdH1/�X�jd"OҰ�Vo�+|��	�N�N�N]�S"O.8I�͘�@��*��zi�� �"O��؄�"L����6N�I�İ��"Ox��\`�e���CaqգE"O�\a��4`(ܪ7N��uZ�j`"O�|��RЭ��K�u#֤�"On]����	&��U�O����"O�} v�Oj�9����
�P��"O�@K�/�6d���Y�E_ .�<�"Op�p�뚕OA"�b��5�l��"O�h��%F�Om  ���M5�u"O��b����A[���F|�R"Oށz3-G�v ����
]$D����"O��9񎘺|���2�h�7�Xu"Of�����&J�X�˄�J�d���"O6\"��:T�����K�h�,�h�"O��ȇCB�|� �{�$�2f�<=0"O4%i`	�1�:|"7����<P�D"O�����D��A����<��K"O`@� d��ɱ0 �9�\��"O�4 ���4s��y�Q��:ɬ�Q�"ON�J���9���GD�q�4��U"O�𙤇��`��5mD|�@���"O =����wu�c ,̤t9)�"O�S#gB�	���LC<p���d"O"h.eD�1e';P�F�B�mǳ�y2
�-=�Ƅ���"P� ��6��y����'�p8��[${�Jw����y
� *��2,B�M� �d�W4�X	�"Op�A�"��p�)xS/�bf�
�"O�E�e(B3
�(�����RXH1"O�30(�sC�x�v�F�|Pz��$"Oι�RO�@�U[5�3%<R(	�"Oj5��Gf~e���פ%r$"O��a�M�8�V�$	�	�T"O��S���	����^y"O�=��F��:P��g�E�Dct"O��f�׭+��|���5A����!"Od�r�Y�tŨ��S(Pջ�"O��V�h:�ö"	>l 8IY$"O��u 	=:T�x��^7�x��"OڰX��<4�2��G�X;;�#"O訣��,�Q�$.�QsT�A�"O�$*j�8������*n��ڧ"O(غ��T����H>n�:��"O0l��(�*]]�yQ�╺d���b�"O4�S`&�=z�(y���*�<cV"OfHS6n�H0���`�<T|�[�"O:�h�=g>�����J
!��[a"Oxj�A�ub,�^�a��)"ON�sY�b<��-�c��ձV
4�y�i�$G��T
1�M`\Х��A�y2Œ	��Djv�$X����5�V�y�U�\�|pv�_7!��QV��y2��H�0i& E�B���5�-�y�f]�#Ų܀t�<�`x�j��y�@424�d�7
Z�3Z�}�$D���y�ٕ+�\�@k �%eF(:�m�0�y�A����\2�ʄ>H"�[b"���y�M��V�"�0��Q�Fk<8"Ql�Py�&��sr&�V��U7�0��X_�<)g�V8�@�3g�F.�R�Y�<�e.�<B�������1Z��p��Ya�<)1c�60��\��+n�� h^g�<!�����R ���0,U���_�<y ��{�쐉�HQN�Z�Y�� Z�<�	��Ո�R��a؊&�S�<�C�N�0ș�M��k��x�f`�O�<iB�z����
Px�d�0��Q�<�qBɞn?�} �k	x���j�SR�<��սg�F�x�A�p��K@�QO�<�#��Ccؘ��EE�l� ��e��H�<���1����W%[?,�Z"Õ@�<i�W>l���3�b�9�����Ac�<9ċP��^h�[B�5p�D\�f��B䉕0�ly���Йw!�Q��+�?m@�B�	�{ݲ�S��>)��!�r��s��B�	70�*L�uJJ(&��`)��w��B�I�@��t�����L���� iK-�JB䉐!���Eq�Pmh��ƹH�`B�<5+�1�2��?4�,��iF
hd$B�ɠ94��a�K��3+D�8çE�i�B�I(ow�ԋ4B��+�ظѤ�/�C�	B���-
bG�-yeb�B�ɄF����2��Z{�}8 )Ыa�bB�6P�T�G��:p*����C��C�	�-(ȳ%`O�T���g�M}8�C�I�a��@ �Ä�]Ŝ��Ԭ�'4*B�I<T�<�#���X^�͐�`A�5k�B�I�:��!zbeT}�T�Q �C��2e<B�BT���V	X�H��d�~C�I6Rd��
��Riؠ1&Z�H1�C�)� �����<�81���ܬzWh�c�"O2)A��K�\�BE�![��X�"O��
�Zz��&�(CMб��"O��Q`�,z��(cт�,n/\X�"O�)�p���J,�����"OX��NCh΄�dB�k� �"O4� �H�.�n�Ňʭ}��P�"Of�4�? ���&H�<R�T(p"O��C.\/&��FEˠ=<%S&"Oy��J՛;`E�bmN�($r�i"O���4�\d-`NBV���s�"O>ᕅD K�(�:�	�e��%{�"O��
ǩ	S��
���9V��ɠ"O�Tpe-�>N��ѻ�EVr $�"O��A��3̶X`���02P��&"ODq���>2u�r'-KrH�V"O� �aE%V��2K 6�P�;�"O���J6 $�|�PC��M�6�p�"O�e��V��*(G�L�Z[�"O��B_�����ǻ�6�"O�؀��l���r6�]<,l�R�"O��1W�< �b٨���a��"O���X�F�\u�E�0[KB��"OV�I%E 5kX�����ǭ=z P"OX��W��oO1�J׀@1�m8$"O�pA�F�b��)�=6���"Ort�%��Z'b��GnqZ�"O�P3��z�9���ȅ]�Yۢ"O�!Ԥ�����S�/f��"O�hkp���NN����$"O��"O��f�F�Z�!԰Mڀ!�"O�F熩߆���n��D"O�A�2Y��|
%m@ն {�"OR�3N>��Qb��K(a�xܫ�"OH�e%#&�xk�j�-C��lB`"O�q[3o
�~.��rήF�5iQ"O�X�   � O�  T�  �  Y�  ��  ��  D�  ��  ��  >�  ��  9�  � (	 � ( � $# g) �/ }6 |= �C �L V �\ �d %n u a{ �� � A�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6j�V����2�81�8	q�G��Q�O/�yRL	0���(%�B��a�B���yb�'nP(7'�7@��*T!�/�����'�$ģ�ȑ+�&4�3iйڐ$��'��HSB��&-"m��+�1~�=��'縜P��5f�0r��
�g���J�'��P���Y�X�kG�`�6%X�'l�e�&/oøBu��@(�x�'	|x
��P�2�9���-o�h��'g�$�e�|[z�Bd�)j�ҥ��'б���͆;R��І6`�6�1�'IBk�ݚDA¸�`-�C6`�ʓ!
���s(���@F ����J�RT�HĆR�B(��h^0*rB��ȓ`&6�h
�;5�Q��Q�1�ȓY;��2j_���d@.6$����a%,����7&���*��S�p�ȓ�dp�Ã���h�E����@ ����c��!z�y���=�\��lb�����'�:X��W;x�F؆ȓe"�� ��}�K�d�1T�����IAę���݀}��3\ib���"O����AB�X��S$�P�E��B3"O���C1eB��7���A���!"O �`�-���ӣA�w�h5�"O�R�ļbi �b��=����"O��S�H�]ں�a��ޞ�Hx�"O�eq�bֶE^�%�5N�$bv(�ȁ"Oʐ��HU/��؁B$�#��m�<a��ߔ$�q` L�	\$���d�<� ��"U��%�kR4+_�Q13"O���g��H�"���	qx����"O��#Ukܔ.T����=Uu ]�r"OT������yK� җ!�"\h��"Or]ѣЗq��Jwa��pZB��"O�c���#}5r� ���ES\9�"OT���,�*v��x�A�m��`x�"O�TSp-μ'*qB植�w��Pi�"O���&�H�p���f �U?��P"O��Ň
d��J���8B6ta"O"u����
C��ҷE.G�����"O��լ�"M�����$�}����"Ox���X�l�$�����/Ѵp"O`4KR��^�d8s�&�r���"O�<��O�E�08y�B���"O�J�`C�;���_.J�H��"ON�3��&��HT��0�z1�"OD8f��J\�eȜ
p��Qx"O����Iƾc����� %�:��"OFPAw�+kvȰ�ߍ.e�䊰"O4Q����M��S&a�*2ƍS�"O��HJT�c�x{���$挊�"O6)%F��
z E�cϔ-gxK�"O��Y�nˎqC��Co+Bʰ\H�"O��J��jENUz�IE�:�`""OT�PC �t���"S���P���"OȊ���9���b�ɛp�D�0"O�����oh1#�)�&�>���"O�܊aoO?���3E�V�����"O�pR�"�[���mD�-4(��"O ���ꞏ]�\r'M 7�@�T"O8����+L�ȱ�ʐ�$�$��1"O��ۗ$��,J�ç7+�X�"O��"A��Lk0P��f_�Y��ɸ�"O���*�*���'L��$��=�"O�ua�i�8X�*����^=-M���"O� �e�P�a_
҇�KX��u"OX �e��:����X�a�R��"O����ظ
��q�B� z���CF"O½{�m�V5���A�@�T��"O�t�cI'9v��*H�gK�PC�"O���@�sa5i
�#�¤8�G�'!!���}j�0AO:[o�t�Q�]f!���A�⨘���TV,�P�I�|!�#c�,����_ � �&Q�O�!��&~�TC��Z���D� �!�dPG������
��3�&��5�!��U�^(v��x��)p��~�!�L�X{�iJ���<D��!QE�1I�!���mƬ�{��ց%d)�z	!�	�U�4L����M���U�S��!�dЗM̅8��	��j��	�3 !�D4@@Z'E�䚵`O��!���<j?��������DK��kV!�pW�Lʀ�֝{�:P2QiI�n!�3DB����_Td����
�C�!���M͉�I��p��É2�!���Ȭ�e�`K�(��c�
6�!��(= @�`��?|�6���@*4c!�$�6�,0�'� B��C#��qV!�	rl����3>܆�P��fU!�dE�C%<\�k��
'R�q%k�F=!�ĝ�2���Z�kƢG%�iؔ�?M:!�dM�j�"�Z�H�,��(gl�I!�� �=�7`�[����N�T$d���"O }��(�4��p:�)��c	�tj�"O�af-ðTm�|`�(:.آ� "O�t�4��-x�b(r��[�ʁ#�"O�����$0�0Řu�A�@%�e�'.��'���'q��'���'���' �m��m8VddP:�l.-�N ���'b��'���'�r�'r��'�b�'l�M'-efb9���&Cd�%Y��'���'��'>��'P��'nZ�MG/
*\����JʤN\�<���ϕ�?����?1���?���?!���?����?��+�
��ӧ� &ZL1 dN	�?����?����?���?!��?Q��?��NM��Ų�ȣ � (� 
�?����?����?y��?���?���?�1������S.[�|����?���?���?����?��?I���?q��H.ZA�EI�N�H>��b���?Y��?Q��?Q��?����?����?)��N�m�"�'��?C%�a;1J���?!��?���?����?9��?i���?Q�d]�I���6�,�Up0�(�?a��?���?I���?y��?!��?��	V}�ųŇ�UZ4�3��H��?����?����?��?���?a���?��j�d:tH�N� - �'��?���?9���?���?���?Q��?��&���ҢC7c!��S��?)���?����?���?!��hb��'rH	69|�A��R#8�4m{p�R.' �ʓ�?�,O1��� �MӰ�S�x��a6J�&]OƸRì�?u�2��'��6m-�i>��|�JշF��s��ŵ�\:С��(�I�"��jӎ�����韞�O��Qcq��-]$�	�.�{�~��y��'��Q�O�$���U�]�p�i�eK�T �c�u��M����=�;�MϻYb���$�@�!(���-
%d!�Ț���?��'��)�S�0l�%m��<Q1ϔ���Bt"� ݤ�1M��<��'& �d�!�hO�i�O��ì\�����E��g�,LA�8O�˓��Vq��B����'�`���^W�*2#T�wK�(kc���X}��'b2O�SP^`$���+V�`ɲ� /���?Q��^�%�|R���O�%a�A$X&I�#*�]� *=+��D,O�ʓ�?E��'�X���Кr��0��mv���'�t7��V���&�MC��O��{��B?^��$kƃ']�čQ�'��'u�lT�撟�ͧpb�d�n�p��"�٤V���
B���u$�������'���')��'2�c�*U�~�` �'J���R�p�4�p� ��?!�����<������i�MˁS�
5��h�3`(�I�M;�i2O1��uY��H��ѥ�.�Z���"iy@&g��Q��KW|��ui�GT)dt�n�q�	���$ ��3-��h1Ȗ�O^�`�$�O���O��4�<�v0���Z$2��cݸ%��eU _2��y��R�F��{Ӷ�D�O��o�
�M���oK`*���5�,8�k�oa�١G�.�M{�'�`�-;˚�4�~��$>���;H
��롤���Љ�ւ@�'�����?���?!���?����O��,*%RH���Aß9bvU��'�B�'u�7M_�|\˓;ƛ֗|��� hd��5J�~X�a�)��'�������3sp�V��<� H�^���14`M�|$�ӵ�@7!�&q��Ox�O�ʓ�?����?��z2��4��+"`�Ԯ�#e���?�����d�𦩁VC쟔�	�<�O����M���S�i�ijFDP�O�)�'
��'
ɧ�I[=H���!�E��!�$�MEzL�Ճ�^
#�6LGy�O�@���Q�����
$:����1	\�H���?	���?��S�'��d����+�x��m�#Gw������]����,aܴ��'t��?��L�#�����R�.�F��(ߵ�?)�/�䬪޴���Ȧ�,��O+�ɪA^�����d�b\�i����`yb�'"��'���'�U>!A �� �`�QkX�.�E�f�D �MS�P��?y���?YJ~�7қ�wLzA��%
*6���/ƿ,��(����Oz7MDf�)��d1�6Mn�d*�&JP4�0mP��Y�d��a�o@CiB�J_�ICy�O�rd�,��Y�\%-@]-S#����?a��?y+O%o�~��-�'2g��h���yƩ��--ƥ��e��fu�OȄ�'@�6��ۦ�O<�r�2j݀�Q�)s��
P��{~R�ń y����1טO=
e�	3WPa���y���"H���c�V5��'���'B�sޡ�b�9[�0=�pFX,,�`�a�ȟ�Rܴ+
�p+O.xm�k�Ӽ[V��;!D|h���ۼqB\@��M�<d�iX�7mЦ)��bЦ��'�Ԃ����?�p'Ŕe]0���X�jK��B
�S�'O�i>�������I������Po���-P�<8�s@Ւ-n�'�6��:�����Oh��=�9O� E�V8D(EC0�
�V��eK'b�K}�z�h�lڷ��Ş�xqE���蓠�6>5z��2jKaP ��'yj���ןhz��|�T����[�g�ꤹ᧙�]��Hs@��T��ϟ��I��Sqy��pӂݘ3A�O�����	f�^`�5�ʯfZ>��6O֙lZJ�j$��=�M��i]b7-@�$��Y �S":�PCBDC.Bqf���l����ɇ\�`���Oq��� *�x@��@FL���-IQ=,��g5O�$�O��$�Od�D�O�?%��l��=0d����>"x�8�.��$�I؟X
�45gha�OR�7�2���y�hR��M �*A�a�80$����¦�'H�x�nZP~�����AS����8H׍�?:/cA��؟h!!�|b]��S��$����40�B�e��Xa��)A�舳�-�ʟ��I\y�JqӦ����O���O�˧$|�}Ӆ&B�TD��2�c_�iH4�'������o�d�%��'���b���$��@՟�U�1Ȟ�M$$0&Am~�O�`��1Z��'ڲ�q�m5c"��bMP�5��K��'�"�'�R�O��ɤ�M��;I�9*�MI58z͋B�J�W�z��,O��l�T�38�ɋ�M��lA4jp1�s��rLa�A)�#ΛFm�H���n�2�h0 3��d�Oƪ��1BX�jG��bq΁�zF4�S�''���l������ş���E��Ϛ���M�1u��f艘Ȁ6��;3��D�O�$1�	�Or5mz�%`�hL|n:Q� ���`��)��BD*�M˥�i\$O1�J���mk���	>1�䤲���z�`�a�T1J�\�	+{� ��'�'�J'�������'���2c�$J�@����T	JC.���'��'�V�p�޴.�����?���+��L��I2N���a�JCa�`��k�>���?qI>��F�>�Q�k�a
V����D~�F�#A� �iQ���4��'����o]\0�ʂ/1
��Ӣ����'���'�)�'�?�#K�nKZ���FP?Y,��zRō�?�t�iQ���w�'Ld�(���8mƅ�Ȇ<W��@���4hpZ�I����ϟ|�Nܦ��'>P$9r,]��I�*������ͺ�Y��W������O����O���O���Y�V̋�����H��Vm,ʓw��R!(��''2���'�M��:y����JJ�$S���C�>����?�J>�|��e&K� ULŶT`ВC�Q�XZ��4!���"�2��r�OB�OJ˓�|��N�(��P���S�jx����?����?q��|z,O<n��Oo>��	�3�$���E����̘.&�FH����M��R(�>��iz�6MC٦1◌R�j�fa����;�� ���$&#41n�|~bD7���t�'ǿS`FT�/�"q���ʁq��D�wl�<���?Q���?������O�s��,�d=٦n�')�lA���<��x���d�$���QӦ�'�,)VC	���S�bMY���˳Aڐ���?���|ҏ��MS�O����J@���A�L�&�k�O�%G^�DQ��̒O���|���?1��vl`Z4c�z��Hӳ�I[M��*���?�.O��mZ�l2��������o��nۓ2/
�cc��w/pe`�`����Ap}�*bӖdoډ��S�d���e�կG>z�,ȉ$S��#pe��kjz���O�I��?�W�:�dյ<��	dԌ�� �{�`���Ov�D�O���<��i'�Y�%��UJ�ٺ��>'=��)_!剗�MӉ�>�S�i��c��]�8*��c��tD��a�~�d�oڿ?N�mj~r띖!,���r�)C+�H]B�K+a��t�"$܄����O����OX�D�O����O@�D�|B���K�d���*I��1aS.Z� #��I		(�r�'`��O���P���i�Q8��!�$�5�Ǎ&Z��&��?9ٴ ��I�<�S�?���+uP��m��<a�٦��p)��z��p�(I�<��Ǐ:�F������䓻?����t�'�mRe�1^�A�a�K(}��2�'��B�'�Dy)�'ZBlw���LF�?Q��՟p�vBWI�A�f�&�
��s�t�ɻ�Ms���y��'��6�i� �v�O |qh�;*|��f"�z���c:OD��,4&܌ a �:2����?�9�� ׺;�'vmqҫ�N��H �~4�)���'�R�'���'W�O��M@�
˳6�HM��
1x��D`�P�q�Rs��E���O���O�O��4�u�O�#[��B��+�"i���Od5n�)�M#ײi#��rñi����O���'	|k,E�e}�,�4����բ��״i`PN>�,O�i�O��D�O���O�Lz��R=ou���I��2m�7��<��iʲ|���'k��'y�Oi�ˎ�/Y�=����""�Ф&����dl�&lr�Ĭ%�b>YR27ay�pI����Hf~��Pb��&$?I!JW!"��$O�������5I�a�+�� J(8�#��>p����?���?�'��ď̦9٧��� �S�0*����c�G�b�`��ɝ�ĳ�4��'Ψ�hǛ�-x��m�u�FK�
=Bk�g�n j����e�'�Q���C�?��}���r����Ŕo��� +�k�Z���?���?���?1���O�Rt	�)^p�C��;z�j��'"�'��7M[-sq�S�M;M>���� ���jEDC�r�H�7cڡ/\�'%�7�F̦��~��ll~Z�p4LE$��H �ڲa��a�A�J�O�@�Č����4�����OJ�Շ+X��XcfI&"�t50D,�Lu���O��$V���֞,@��'��P>Uƫ۱=gDXٖj�:g��k�H.?I�]���I��'��yr��+2�=K�q�Gǎ�=��H�'��<��T(ߴN��i>�9��O��O��$��?.��\6�Y�	h@���O���OZ���O1�˓"X�&.ZNr��0��#3�Hq jZ���tW� ڴ��'?���?���}, !��X'k��������?��2Fށ��4��(C ��O��)� �)�ŀ�&�r50u�~p:���?O<˓�?9���?!��?������ a��H�e�I4FR�rf&ވ+��nZ	I�1�'����YȦ�'=l� ��#Y�(�z�i�����4��F6����p��7s����.ܺQ�΀�v�K���֊t�����km��l�INy�OQR愨` �ZU �Y���@^:5I��')B�',�	��M��H���?i���?! %�>uق�j1��'b�:#Ŕ���'X��5ۛ�*|��%�`ӔɃ
2��\���p
D��' ?��O�!`b�DP̧���DF��?Q��6Pw�ĬR�R�:�	δ)�b�'MR�'��S����fmԍ��(�B��M��!�����)�4_|�9)Oio�_�Ӽ�E`1?�\��@fU�g�p@K��<�a�iQ�6���q�%LŦ�' 1�i��?�"&EI!>��rEX��@�[Fƍ�^S�'��i>%������͟`�ɇ7"��Y'FV0�a���76.<�'D6M �eԺ���O��*���O���}�*%�Y�8�R�a'#Q}r tӜ�lZ��S�'	�]�4隈N�&��/F�x}�HSцO����'����f��ޟ\Ù|2S��cƭԓa �XRjۿ]t9"%@�X��؟������Ay�/`�̴� �O6�:���<"A�1;���t�X�B?O,�o�u��T��	П��IƟ8H�J��Ux�80 �*0j��t���b�o�p~"/Ӆ[���'�䧅��N	%=���0�W�#��t�$��<Y���?���?	���?!�����1�چ���*;t��9Y4��'D2Gg�|C6;�r����%�`��.\(<�*�j4�ɥz��kv��f����d�i>M�c]Ʀ5�'��
���q�x���0D�媃�G��������d�O��$�O����*ܤ�j ��� �ӂ�3�2���O��w ��b�n��	ß��O��DءF�>K��@��ho�ш�O���'��7m�ئɓI<�OS�-��W�Gj�aـk	]���sd��I
&q����4�"\��,Zr�O|ЂG$�'Z+\ h���k>��p�G�Ob�D�O��D�O1��ʓ;��VeJ�lm+�&�?P&&�!����I��MS��b�<�ڴ�J�)��#Tޮ2u�I�u�^�81�i��7͘�Y�6+?AƎ��Xں�I+�i <�`����<1�}*���y�^������P�������ɟT�O�6�P�AL��<#�L7u|A;��d���
�)�O���OH���D	��݃[�ԌY��v�(�`�;�`=���?aI>%?�R"ZѦ�ϓ`k�� b��5e� �����$w��!�Y�N�O�M�K>.O����O����~�T-�A$ڵ_�`����O��D�O��Ĥ<��'����?���e�I�n,_���@bD�] �(�RH�>�i�L��(�m���k�|!ty��Ɖ�;��I(f�B4�3 	9Q}t�%?��'wt���6)�p):*)p��Å )�\��I�x�I�����r�O���?fZ���VJU0`�p�`�Π��!mӂu��<��i�O�.N�lM��bѫa
�bb�� #���O��I���C�ئ]�'jٱw���?Y�V�͜2'txjR�	
��������'�I����	�H�I�����:(��4R�gj�3��vժ h���<���ivzܢf�'��'��O�����-���7�%��i��<}ל����ӂ�'�b>���c���lp`�ʻ\jL<R�e�'HO։���.?Q��ݶB���$ӝ����DS)!7Ɯx�䁹"&��*# ���O���O��4��ʓL������h�rO�;6'Z9׫�$��۶�Ʉ]�B�u�b㟬h�OH�m��M뇹iKBѻrS��9���P�v��3J����X &��R����)���:������x6�U�	箩#=O2���Oh���O��d�O��?)���٩�U9E�c2�"w�X⟄�I֟���4P�Zϧ�?QS�if�'\
��BH�9F�xj���0�,�B� �D��A���|����Mc�O� v�O@&���J\.�F����W�"�i��e�ƓO���|���?Y����г#̑=�.H��	�L`�-����?y)O�qm��N��'�2Y>;2�ˮp�H-��@_#|Hf��;?��W� �	Ѧ�O>���?ղ1�ҀuO^���OO�]�n�ˣoW9'.��C�9�v��Ef�O�� N>Q�`�4U�d���Y���-�?���?Y��?�|�(O��l�)[(���RM�(d��T�<9A @�Ɍ�M� �>q��iZ�U��E\VGDBf�c���Ч�zӬ�o��s!�Ao�a~2\#V^L0��T�)��,`��!%=��d�K�'��d�<!��?���?���?�-����WI޺,�4�0운n�$Ԡ�'P�����BџL�IƟ4'?I�I��Mϻ"��0ː"Y({X�T���db�!(���y��x���`��9y��4O�����J�T��*��m#b�9O��8@H��?�6�8���<9��?�AC�99ĴBB%�9M�����?���?Y��������W�˟���۟D��D�1�$��WkN�HQhf��
+��ß��s�ɉyF��Y4��f}��`���R���l�zۃ�:�M����&�L?1�J5��ҕV>:�(X����#6=����?����?I���h� �d^�>U�7Hޤn�Ա  �[	&H��DZʦ�����x�	�M���wc^ac��B�3c�T�j�:�'�"�'$BH�_Л֚�� � <��� �L@�.j��.�7��m�eK ���<��?����?Q��?9f�_�:�6u��
K�G`Fh*B����$���I�`ȟp�Iޟ�'?y�	��P�Kצ� I��q�5R#, Z�O���O�O1�2M�Q$���+T��]`v��"�	
X`7�Oy�kQXR��������-_Gv�7��n^P�2�H
p(���O,���O �4���������۝�|B��"��D�pkN�[2��aӮ�{�OLPmڅ�Mӡ�iI�S�g!��� ����h��
ѐtΛ6�����N�i����i��y�4�	:j�rhs�gZ!zPk�<O��$�O ���O���O��?�J��B������(6�X�������Iʟ���42���O�7m=��F�;"H��CЃ"r�l�V	�j�z<&�`�	˦�D���l�L~��0�L�c�Y!���зcܭV�(��� KƟ�R�|�P��ڟl��ןL8�H/�3 �_"5�я�џ���iyB,a����<�����)U$aeL�I�:Ւ�2ԡ��A��2���ꦥ��4`����߁9i�Z�"�p�a9��?H��8�&�*�|�����Ӑ^Uv�ɈL�=�ĭ �8��d�c-�d��ҟ�������)�ny��t�l1S&�T�`����#)���c�D�YSF�D�O��n�^�a��ަ��C�\r	�>3�<����J��?yٴ=�.hڴ����� ���n�ʓ|�U�N�_�V�j#`�������O*���O��D�O���|
�%�1I��K�)C���L!4d���K+E2�'�"��$�'��7=�v9��$3,���B�bÔuӔA��M�5�'����O��DcE�i+�d�K��P����r��`�*W����%D�y��e���O�ʓ�?�s�:H Rf�q�� Jנ�p%hA��?1���?!-Ojdm��8U�'��a� \���+!އa*�Z#���O̕'��'[�'���	�a�t�e�K�7����O��9c��gl
p�A�4��@��?�A��O�����+��]� nFތib
�O���O��d�O�}λ�2����E�R:�Xه�ʎ3ݞ�r�N�֧E�+�R�':`7�3�i��aS�?[N��r��kĜu�hj���۴3\���z�
-2@'x��Ծ8#�������3�ڙ�ȚNK�	�D�R�����4�����Od���O*�d�I�>ۆ$\�L��a��
>5��T��M�'Pb�'����'J�����"hqm�kH�KQ'�>����yR�x�O���Oм8b �8�:D.��=X"��瘹7��b!����d�~��$+��F��O��&�~�B��D� 0�bU�t~����?����?���|.ODHlZ"c�r ��6'���T�Y0:��kT$!7�:�	��MK��g�>���yҶi�Z��O�&ɴt�qȵ\"�a�cj
 G�Ɛ���&f�'W(��I`�����kJ$}�`��1���?�v!�Iy�@���|����������J󃌆e���u#���"䂧+M��?A���?�2�i�D@�O�2�fӤ�O�Ȃ�O54�LM�� �����(a��l�	��M���J�b)�MK�O��R��-3 �J��q� 	�&jTA����!���O���?���?a��R<u�'�X�p�ԍ�*U�2@Vi����?�/OX�m�3ظ�������IX���I�m1B�qei
Y(A���7��$UH}�Os�6<mZ���S�D�S#VB� �K�%#X`����c�8�`��*r�dQ�O�)$�?i�@$��˼Cl�̺'�δO���&�X5F�(�d�Oz���O���)�<��i{�2���TgZ,�p�S�%St��΁�c�R�'�<7�*��&��dæ�Z��P�>���Z ��(b��z1,���Mk��i�`+0�i�	�?~�z��Ov�'?����^�AC�Gn�':������O��d�O����O��D�|�tO��T}�G!�D&�0Re�J�o��66O���'����'��6=�.���X�C_v%x���%�-ٔ��ʦ� ٴY���O�� ױix�d�>(Oz1#g��tĪ�Y���11�|r|�p��P��Ot��|����01�R����H�`	�;4��Ep��?���?�+Ovdmڔk&��Iߟ���3.W����
׿Y�}�b�۳MV  �?��Y�,�ش/-�vi*�䆼$Wz�B2��4w��M��L��`��ɂiu�5���:K˜c>]��'����I$!���gB�B�zL��G(2���������I��|��a��y�/.e��X`i@�l���I� _�BjӼ�J0�<6�i,�O��W�N�C��)oQ�M��o����ߦ�K���McĢܹ�M��OU��S��*�O�?/��l���*c�V|F.�9w��OP��?!��?���?���&��(���N�p��v��5B��*O�0mZ; 7����֟��IF�֟��
*5Xh�o�!D�Y!�f�'��^r�֤�OtO���D�ie>�
�d���P(�R�@7�8D�fb�e�˓-��� %�O�-�L>�(OB�e�	ҍ��c��L�Q����矬�����	ß�S\y§t�x�T�tޡ��^�5��i%�T΀%�%;O��nZ@���	̟ �Iꦭ���N3a����2,S�oNf9{��Gt{� lZA~�왈a2��-"4�Oi��ġ*��<Kæ��L�%���yR�'A��'��'����
�p����j
&#���P�@+��D�O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!6�D�O���&�i�O��nz����j
0mb �(�Vy�W��%�McS�'���t�O���iWBW�V:O�И�F>���Q�l�
/wh�y&>OnD0bh�?�r�?�$�<����?�pD�1|�%8�#�/�0��gC+�?����?�����Цm�1�̟ ����"�;pp]SW��*����w�m��$���	�M���i�Oz��3�U�&&��2ª
{�U*��D�%������.�S��RϟL���oˠt��d����e��GM�����T���� G�D�'��@�2��=&���cD�N�v[�ٱ1�'��6-�V���PE���4�n�+sG8Z�-Yp!�u�8�w�O6�i��m�l٨�m�M~��\�Z��S�;�*��Q�=Ю�@���/,�n1��|�Q��Sٟ���ӟ�������X��Ʀ�v���Myy��}�\�{���O���OH����ܸ:��vƈ]}<�w�C�����'�D6�ӦU�H<�|���o���bCY_(Й��ԋp�܌�Ѐ_~bߏ�&���>s�'��I�9�*a�q!F�fEz���$�:���ʟ\�I��i>!�'�f6M��w�L�Ю+�����+I(v �jV&V�8�����=�?��^���ݴ(���(w�X�!$�8m¥iqEضv0�:%��(}6�%?�Њ��`��'����1  ��<m��3��[�L(��r1o|�����L�	��x�Iޟ��bT�U %��5z�I˛q��(�h�1�?y��?A��i�x�:�ONAs�T�O©9��݈g���Co�E,��]��Ovo���?���Y�B�lZm~2NM�'�NŹR$�A�g� �>��4��ޟh��|Z���I˟8����Z5���r�� �㭛�Pa2,p��\�����fy"Dr�Rt��$�<����Iׂi�s�ɱ~� �U����ɜ����Ǧ)k����S�A�
�0�7/��hZ6ܲ����o�� H:A<���$Q��Ӣ0�b
�V�	�!R��)�$Z!�����1o�y�	������<�)�ay��`Ә0���Pz1��l��I$5���	-e�V���O~Qn�`�@��I��W�0i���VxrQF���?	�4g4\�!ߴ��DK�)rde��'<�8�H���-�m��YV�T�B��IΓ��D�O~�$�O��d�O����|r�扳Z'�| A�Ěiʮ4hch�#T�V��%�'a��'R7=�D=)e�3L��EÝd��i�F�O���4��	Z��66�e�������|����&x$�p�l���l�(	��.�d�<���?9$�SѢ�1'�ىb��%:7Q��?I��?Q����T����r˄���	̟��7�� 1PJ*l�%�3,�x�[��ş�Iv≐h���"`Id�U�n_�o��4���+Ĺ1�PH~r�k�O�)~�P��c�o	B8�5-Q���?q���?Y��h���d�$oDX=Ѓ��6Jz&M�%��.���̦���k�埀�		�M+��w��c	�A��)m�	9�r�J`<O,���Ot������6M$?�uB���S�y�vL�.	�  �'v�P$��'��'U�'�r�'�����J/�Nmi�F0K�v�Z����4��]/O��4�I�O
|�W8;mX�r��E�tTc�KGg}��'���|��to��i��I���#�b�a� �(Ԙ��ihfʓYp� P!���%��'SL��A �)�@Ekf ?���C�'m��'U�����T�p�ڴZL����wDm�oG4+�~���dxL�8k���$G|}��i�`9mZ9�M���\^�P��BP=vlƼ�禋9R��c۴����t�r���'��O"��֪��Ta���t��t�r�8�y��'�b�'���'����W0D*q�կ�4آ,s�!R�p�x���O��D����k�K�oy�z�0�OL��*R|���7�B�L�k���z≽�M3����T��C^�&���Hg T�t݄0���Nč��
� �fyjw�'8�$�p���t�'���'�n�r��[,)�B v���d�'��P���4O7P����?a����	D9sN`�kR�'��x5LD�Td�	���d�O�7�A�|��ʛd�`u1�-��$
pY���;0����ɋ�x�
���l՟D���|B/JB4������L��+؈i�B�'J��'����X��j�450J�"���th2�Ї:Ĵ,S�� �?���j+���D]J}��'���@+/%�֌q���=����e�'�-)K������OI)5g�ɽ<��)�=Q��lS���KB��<9-O���O���O����O��'��-��/O�7s�}��?���M+�
�?����?	H~�� ���wB�Y-�f|����˻(����$�'���|��$��%T��=O� d0�f�	d�����5LjL2v8O��@4M�8�~|rQ���	���V��]���y�,:t���5�����	ϟ��Oy��p��U+�Oz���O l��� �jF@�����")��P�O �	����O���?�$J�9�L貢�;%�~,\��A�O�S�.cض6-AF�\���O�����H�9�K����A���O����O��Oң}��.|2Tab�I |"53b��9H_`Ձ�� ����2fE"�'c�6� �i�ݪrj�y������o�p��q�8�ߴh#���{Ӏ��F�m������xe���f����7;�*���ͮK$��#ʛ��䓏�4�^�D�O����O2�Dک,ײ]	��'c�>����C�!+��>��v/:��'�����'p���n�dh���3�EWb�$���>Aa�i�\6MU�)�s1g>�&T
�oY�h�(��3�߬�r��J*?��^?T�������$�f� :�k[�c�P�)�Iu�����O��$�O��4���@�F.	�Y
RS��� �0�@��	�y�h`���
�O�hl�?�Mk'�iY��+s�E�]�xH��+�}(�Fٻj�曟�����k����i��(0�!IӼǒ�a�CĆL�dy��:O6���O����O����O �?����^-�7�PC��k�O������T�ݴj�J�'�?��i�'�Zz���'2�9k�H�,�،��5�	��Mp��|2U	���Mc�O����#P.�����o����&��#?� R�5.*�O���|���?A��(���AbĜ/�F�zJ۸/�L�0��?q(O,4n�O����	��	W�4i�d�\pB$��[KLİa����Q}MӦ�m�?��S��ȹUi8}ґ���:8xñ��e���Y�+�:tʀ`�O�)�2�?Q�d'��B�1\��q-�*->���F��>=����O|�D�O���)�<���i'h�ɖM�.t���H��^�"u��l���'��6�:�	 ����O������aI�c�*�G�,��Ģ�O���I��B7M6?!GjPL����wyB�T_ժ,��k�Nv�h�����y]������4�	���؟X�O�V��f,ܛyz!��Q�"D�i��rӔ���A�Ov�d�O�������]_��<`�)E��pcĭڢ
���ݴG���%��iK
M��6�h��y��6&�f���� sV=*��}�xcba�I��`�c�	My�Oib ��<,J	��L])t�
-��DwQ��'��'��ɜ�M�6�Z:�?y��?� }�T��f�:X��r挹��'e��S|�v�m��<$���gF�ri�xI�"(74Yp�3?�l��bަx��
Nv�'lݨ�DO6�?IWƌ��� �'呴C����'�R2�?A��?����?��9��Y�fߠ2�ƥH���4�u�v��Ol�n�{t�'��6M6�i�I��Β@������>�J�Cc�g����4s�F�oӺXh�$v�j�@2���&䟔�閤�Mx�9�`�^9>��� i|q'�������'��'���'w<���#T5���X��N*0x��V���4Gl�qJ��?������<� ����Вl�2~ �[�g��0��l���S�S>(A0$�jZ�2נ�qǠ0����Q�^�$�b.88;���OTI�O>-Op�9GgF)S�0ڔ)����P�&�O��D�O����O�)�<���i�X�p��'S�T�%]2g���b�

�6���'l�7�9�ɔ���զu�ش,c��
��Eb����^�PK�<�A'&z�� �i���q����O�q�P�.޹��e������h{垾B8�d�O��D�OJ�D�OR�d'����@�d�0>[�8� ��4�|�I�$�	!�M����ߦ&��*�M�!C�
$M�t�@a����h���Gy���Xn�D6�"?U�R���\��b�7$p��y�#?1իE*�?	�-)�ļ<�'�?Q���?��W
a��1g�)�уԅ��?����$[ئ�������I֟D�O������]<yp�aG��좹c�O��'��i�ؓO�S�1Xq�K�	_��H��^hx�۠ʁ	m�fSPe!?ͧ�$��˂��W��("��m(�P��)���y���?����?	�Ş�����Rw�ĲS|�BTC��zt(R��/y�L ����j�4��'���fJ�T�)���	~ n���V!�6�����`2a����'�E�q���?�&>���V27t�yB4G4���2Oh˓�?���?����?���;>ժ������4�/.�HoZ(�������	A�s�<����+�鑤a���p��1
�bek����B�2�iFܓO�O:G�i���!�����͕}\��H�æ��O]��P���A�2�O���|��j�<a�$@Hp|饏�
�0�����?Q��?�)O$��	< ^���O��`��|pw��.D����@ܛq)�tk�O|��}��$��3f�	t�<���#�&�9��??a#�@�yr��#3B�/��'}q�����?�R�N	t!\)6Ҿ! du��(���?Y���?���?ы�ik>=h���p^��s�� ��,jB�O@1oZ:l���	ܟ�kش���y�@V�l
m�dɻtܼkĂ��yp�,%��ۦ�
�%_����'}�Tkd��?m
ч	%cD�0	G!�;����s��e4�'��I͟d�	ϟx��˟����<�i�f��+B4
�k�J�V�`�'�p7홞,T��d�O���5�I�O&�S�\ ����Y]��Rp�EO}��v� �Io�)�xl�� ��E��&׾x2�@G:!v�MI6�U�]e�����1e�Ob�!I>/OJ	��
�X8 ����K���:3��OV���O�$�O�<i"�i	PUa�'�]�PA�>����]�B[ ���'!P7�7����$����
�4Ǜ���cV��b
AtZ���HU�
���i���"U�F@ZR�O�q���Xt�����lj�XI )܊ry��O����OB��O��D6���T�����T�t��fl�5{�D�	؟��Ɋ�M{�#A]��du�B�O&�0.��e'>dz�$ VE��i�M�����lz>Y{4'J��-�'ht
'�E<h*PbvK�
mF�+���3\���'f��Q�앧���'���'dJ,�Z?9:qh��=����',rP��i�4=�x���?Y�����10|��h�4\��U*raY2v��	���d���ڴ ]�����bAD yS&*G��R��
#_�2����;@)a�b����v�R(�;P�'���e�9O)� j�D��C	B�2�'2�'D����D�'�Bݑ5P�ȫ�4H�tH�	�I}P��dG�\��@F�
�?���?�M>�������%�2��,&��ڣ�E�YÜ|	`�0�M��ic�1 �i�$�O�l��g�P-�̺攟4�&D�IF �M�/x̃CMo���'��'Eb�'	2�'��ӽL%��H�"
�l������7��*ݴ,�@���?���䧶?aѶ�yGG���,a��Ҭ�'FA�t��$l�|�&�����(�nr���ɺ}Y�����E*LӀE+ӣ=A*�I�:@\��D�'7��'�����$�'�0�Z�)�.c��s�Z�]Q2D�'�B�'wbQ����4~�=���?��7��+5��I0٪��_�]i���>)�ib�6��H≥P������Ty���T$xK(�#p�J�W�1��T�|�5�O�T���`��=b���#z$�3�N+2]����?���?��h����M�8�r!AY��@	Q�G���$���Ѕ���I��M���w�l�K�>/X��X��t�'P�6��æ�#�4?b����4���193�-���5V�
A��hP���B�	˸�*�B%�d�<ͧ�?A��?���?1�%�1y@��ir�Ӯ4��y���H�������������I��(%?�I�-I�}�!�u�`	+���^�ɪO<�o��Mc��x����k�"��EŘ0m�B�5��V�9U$�)����3N�:��V���OD˓gfx5	r@��,Q���rʃ2~����ɇ�M�v�+�?��G�FfKJ6>�^���*�;-:��/�M��Ȭ>i���?����*��W$_�hp��@�Y*,��U$�3�M��Od���
ĩ��d���w���3��@��'\�]Bl��'��R�R &��Q�
p,�r͋9n0�I�q޴7��u�O�6�,�$�'ws��R�DÉP�r-K�bU�|�6�Or�d�O�)�32�7-0?���՜S~����j��$�6,�@��6	&����� $�̖'�O^�*�K�6�^�c�F �*w�Ɂ�M� �����O��'�����,
$)q��b���d����'m�ꓤ?1���S����*BHK������\%,
�\��!��%�<�'t�	~�I�d�2ȉ�bY{�T�@��G�BC�	��M{0�B�*5Tő�!�2�N ^X\��o��Ċ�1�?IZ�\���و�BA��V��,���Y�qC�)���`+�����9�'�P����bJ-O�*`-�'mʍ8Rd��$��9q?O����=���x�L�:��Ì�@
���UP�����[b�Iß����yG)��m1@p��c^0e�($��"5_��'?ɧ�O��}�R�i��d܄���U/Z�@�h�r��Xp��*�'a�'��	؟���6Z@�0�`E�f��/�Ow~���ǟ��	Ɵ��'W�6M�~�6���O��$�/:V ȃ��J18��Yp�KL#G���ty,O���xӆQ$�\�f-N���`�D�Ό4.�:��"?�t	
-�|�r�U�')��$�?)DgJx� � )L].|"��ŏ�?!���?q��?���9� ��m|~��
�9�y�ׂ�O��mZ�
�`��	����4���|λoY���"�27T6`�e[��ϓ�?q���?���*�M��O�س�����f��V�
�*�kZZ>h����l$�';�Iɟ��	⟰�	ڟ��I�R�T��ŋ?B!$	e��x���'�p7-E=���?�O~�]X��K�a�/����T[�Q�U��Iȟ�&�b>eP��Zke��O��o.ҍP�Y��|4o����D��2�1��'X�'��I�60�9q���h����%'�N��	џ�������i>��'K�7m�9l&��D�&�Շ#
' ^��a��.r�p��*:�V�|�Odp��?���?a'��Q�� ��+JV�A�c�WOZt��4��$�5n�i�Ol�O&'�*U�$q3��8N0{d:�y��'�"�'Yr�'���)P�B^qX%f��=0�����?�5�i�����O��r�p�O���'�}��q ͂K�4Ey�8��O4�4��Dswӌ�c�&�鐺��Ql�8&���� ZO1@��OT�Oʓ�?��?��!j����Z&���i�h�`Y����?q)O0�o�Z�1�'�B]>�1��ЎED�i�0�ڤ-�0`�G,b��������O&�D&��?� ��H��Ϧi�9��F5(�8��a�
�4F�!U�cӞᕧ�$h?�I>iUB,�F(��&�2 (B|��]&�?!��?	��?�|�*O�elZ�=��(2��T�X����U�W�u�ƫ���I�M#M>ͧ8��Iן�Hg�I'8��xC`�ݻk4\��.�ٟ|�I�J�@��F�=?���e	��cy"[!�YP���x�P��@\��yQ���IğX�I��I؟��O_�H�W�\4
�������+^1�3_�Mk�_����O���.�$����2�N؃���!j�<3aBېY	�-���('�b>]S3��Y	�	�HG^)���,G��aU/�/*W��ɢK�`�2�O�O���?i�D1D���F �A������]�p�������?����?�.O�LmT8d��	�����1�0c�Ȃ�G�����&��?)�Q��s�4=��f#8񤇟hvŁ���<.e��+��/�Ɍy��dy����x3�b>	YW�''����V� c��²L�-�\�I��,��ɟ���O�O��C11M��C�S�BHP��'���wӂuxgJ�O���TǦq�?ͻM�@��
SZ���4gQ�<����+��F�|�6�m�C? `z�8?��G:0��������4:g)�j���E�L|	�H>�-O���O����Of���O�x0gCN�zA\��ۦo�8�ŭ<9��i66b �'o��'��Om2�G�zj&II3���Np" �GI�5*�~���eb�8�&�b>�p���=7�ԭ#B /�&;7�'85*�{sm5?v��Ct~�d�*����D�G����@^�B�Y q�T�i4���O��D�O"�4�D˓A*��'Y"92�Wrt<آ��$� �����y"gӐ�V�<Q��M���i�
���!U�|��܈`țsh؈`�ؤEP%��O���[ ���d�w4�qBtb��I%jmB�G'�N�Y�'&��'NR�'��'�<�D�H�� �3�	�8[Q
�O���O�`lZ�gqH��P�4��{�VuK`��;˺�@��5!�����x�h`Ӝ�lz>�ta�e]��y�>t�f���re1�ډ(�-�P�a���U�����4�����O���]-���� �c�\̊��4����O"�2���PM"�'"�U>yv�J�#G�y�C� WM�( �8?	�Y� �I��(J>�O�>A3+�p�H� q����|鱖�c�N�$�Ĉ��4��x��a,�O�d����'�����ٍb2~(�d�O0���O����O1���e�F*��v� BpgJ�Z� �#H�$��aa�Q�Xz�4��'�Z�"���8$2��eM_��@D�n�6MGæ�r��rr��l�+�f����O����d&�;�J��SC�?q��Þ'd�	͟������	����Ib��(<&�P5�Ȩ<�L�6e�#Ɗ6��$6� ���O���1���Oؤoz��*�Ɏ%{�,:�߾RNrɨ����M�C�i��O1��|15lt��$@�0�s�>b� L��Ɍ�*��� �fw��s��S�ΒO���|Z������-^��`9:�I	���Z���?)��?q)O��oZ-e���	ʟ���f� �uH�@z��c���1W���?��Z������sK<��LʒJ�nY�dc�y��㴥�k~R��1��AqeIK��O��i�Iw�ܑ%`�Y�#K� ��D
�@Cr��'���'R�s���!��Y!���n�����O�0��4 �qi���?q�iO�O�Ή�r���j�dX�H���d���-�ٴD5����NE^��O���|��S�a��X�Ӄ�-�5�T��%��EQ��|rV��ȟ��	ޟ��I���`p�@�g'��d�"m���h�IFy�d�vh����<����'�?y!�N�Ҋ��Ԃ�f�R�)��  �˟�oZ3��S�81���B�C�|��h�/K8���A(+/<��]�U9���OPLiL>-On�B�e�[�BE� ���t�8�,�Op���O��$�O�i�<��i9�[&�'��<�$̔�9�'.+�Y�'�Al�⟸ �O��d�O���Z�l�tiR�Iؒ3��U���H�UM>��`��&��I�n���ݟ����R��u�b��$j��U駡��n3���O��d�O����O��$9�S�F��P��a�'��)˔�8�a�'��t���8�.�$Ʀ&�T�uNº?���A��]>59nd����e�I���i>�Pf-ٝt/X�J�NI�W@O><rU����m��D���هw���G�zy��'���'�ҏ�?n$`g,�?n� 5�L�.�"�'��I"�M�Lډ�?mf��$�|*�]�J`٤ D3Xr��#@b~B
�>����?�L>���M�sL�6��Z%cǍB���D)�:$�ؒ�*uz�i>���Of�O���$O��v0	T�̯>�i���O[m�Ɵ��	�b>�'6�6�Z)DǼ���^�p;�і{�< el�O��d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q6Q,��M��w�8���D|f�04ʖd�2�'�b�'�r�ča�:���O�Aِl&���@�T�����T�3������R��'����$�	Ɵ��IƟL�I�j���Xp* ��Q�K�(
�P��'��6�	I�N���O`�$4���O� s��~Hѳ(�
��aI�r}��'�r�|��T!�)�>)�%f(&v���ƞmK@�cɓ�x*�	<;�iq@�OƒO�ʓ��a�F�W35 ��d�~!�M��?!���?���|b.O��mډEȤ��Ɏ)���yCi��g!���rm.���	��MC���>���?�;�B��dG+R���+ʬ�Z!L�:Hv��'V�YЅ�RIbO~����F��@
\"������(>�ϓ��?Ї���Y�$1baL&�����O
umڎd56�'*I�֘|�ë8�����Z�M��2� � O�'�������77G����O�`x��37��	�M����mk�͗M�.9S�'��'��h��9E� ���I!j���td�7�Fx�eaӖ�c�<����i��h>��W
N1>VV��$��$cE�ɓ����O���3��~��B�?��H�KA6+�({��'^nD�۲fE~��D����O�[?�N>����jl�(��ގ}�H��ՄR��?���?����?�|�.O�oZ2
/� Ӧ/WsM~�!��_�g�V��5�J��	�M+����>���2v�] d-G�x�8�AŞ=S��@*��?)��1U���'���	V�Br/OƔ�� )�$l�5*�^�B��5O���?)��?����?����I��d�u ҃e���� :����Ld�p�B�#�Or�$�O���D�ئ�]<�n�0��,$�0��:H$�	ޟ�&�b>�1N<:���2rL��HĊu��PC@���F] 牬~�D�Pg�O��O~��?��d5�a�LF�/xP�舚��(���?����?�*O���	�y"���O�( �by9aU`�z13��:��$P�O�}m�:�?iN<!�G@�6!Z�C��E�:�d5�M�x~�f��&}�a��&Q,�Ot�I��$Qer��z���'mΤK|�h�Ê�I��'�b�'��ퟬ0�!��a���2���0YN~��0�ȟx�ߴlqƑ:��?�@�i��O�ʤB���R͆2�~U��!��l�DP���Y��M�e.��%�
��'�(��0�Z�?=��!VG�ҁ(�=m��J �ܜ/V�'n��՟@���L��֟���%�tY�!3o���4�A ^VL@�'ʹ6��}�l�*���O��󄜞RP��o+��eHsO i����'3d6mƟ�$�b>�Q&ˤ{a��[�����`�]�#x=����iy"��w���I�F��'�ɷAF|k�e�.T�.)(#����ڌ�����i�n����~y�'k�,���f�O@kP��<���*')-7�J���#�O0�m�W��Sh�I��M+��'��L�1e �u �F_Y��QC��@�����X������i���F����.�.��]�'�[ ��%�V�A��$�O����O����O��$2�S�^�5ѵjR,��)1��V�EhR$�	ҟ��	�M������Ǧ$�X��@N'�t��Р .�K��%�ēa ���O�4�P�Y���O(]�!Ǟ�%n��ڝob�5P��՛P&�E��2�O���?����?	������GD�=�H!vk��H:���?a+O�������D�O���|GOI����J�$��`uZc~�n�>a���yR�xʟn��@��w��5�p�ϐG޵ 4�F4���#��fn��|�&C�O6��K>	�e��B�j���+k[�h����?Q��?9���?�|r/OЌm��H^<I��_�C5xxa5��#�6)Ia��ҟh���M��R��>Q��i���QI�D�3Q�&P4���D��O&6M?S�\���H��*�G��$	_y�J\�E�	ct�}��!�i-�yRQ���	��	П8�Iʟ@�O�~��񃀉kq*���A�;.�i�np��p�bM�<i�����?�Q��y�X:{�r�!�/��~��n��%.�o��M�7�x��D��(*��,y�'�J	�%EL�5l���N�R5|	A�'W�X����)E�|RW�����JR'gOr��VAN$iࠆ���� ��Cy�H~��	;3g�O�$�O�J�S�%\�2d��N�@<�a�0�ɇ����צ9�ݴq��'�L1�ɝqK�ఀ���F'X��O��ea�1�
�x!��Q��?)!��O�B��CJ�U{%��-#���5��O����O:�d�O��}"��v������;�v��vAE�&N8��j0��Q~���'4�6m:�iލ�#��.�%�[*X�(X��������OT7�¦�pC �?��,�`� ��0P�l�7tjHY�ŋ�T�z���a����4�|���O����O��d�'E��D�3'��Z�H��w*�j��\�F�F S���'q2���'�xd��:l�9j����S��PB0j�>Aa�i��6-X_�)�S* �,��!��q��$�,N'��4 b�1HJ�L8
�p$�O��hJ>�(O�h�1K��*u�!$�95Nq�(�O>�$�O�d�O�i�<	2�i3��
��'#�d�U"E��p�� �D���)�'V6�6�����������۴g�� ؀�IWr�s�����=rA)�>Q!��� {T�R�1���	��ʔ"���0AxT\`���%�2$��5O^���O ���OP�D�O��?�d�7?�Z�8�ՐZ�)�T���d��ϟ �4�Nͧ�?YP�i
�'n؊g�ĩQ �"en�)�djb!��L�i���|�φ�;�F��'k���M�64@yh�)=�H=��؁�q�	�v��'��i>I��؟d�	�lt��Dk%t6TP��^�#�P����d�'�6-�3��˓�?�*���{�GM
i"R��s�U�v��5��X
�O6�lZ�M��xʟ
�*�J�'!H�T��!x�mB&@/?�f�	4��DD�i>��c�'��T'���e.��Vh�1$�O�V�kcO�֟��Iҟ����b>��'(7-��A���9,�-����%�Q3.��̬<a&�i��O���'I6�D�N�DU�B��WI��y�O;�Mn���Msw��m}ޥ�'�.4#AL�?���&m�󦓅PiSB: j��57O2˓�?q��?��?���3G�ʡ2���:i6)�,S'�u��i�bQ�5�'���'���y��d���\�[��1�a��P۬q���lU��n��M[D�x��$���m�`��'W8U �F��Xl�G�н*�ϓb1Z�pi�O݃H>1(O���OX��$#E�,�hjE:M;�i��O*��O�Ī<ᒴil2}+��'W2�'��8��Y9tn�zE�Zt[�d�K}y�(�l#��NV�%Zd'�kxhMڕ�[�'�L�'�𼘤j�e�5���tSٟ���'�|�C�@�0(<�JT$��Ģ)	f�'X�'��'��>��I
4\�l����bOS!J��I5�M�S����?9�j�&�4�t4��'�<^褠���b9
��=O��o�<�M�D�i"���ٷ��$�/98�3��jxB<���Д+�L	�`f��m`f����J�VK�0�.�9
�yF�<W�����%[��a8⃖�yH6�t�M�Js�9`0J�<>�DQ���m�vp�ϔ8�,B��LϊQD��$��e��2]�H���@�[�恚���4OD��A+�+B~�T�ݣP'���H��Z��C��U�5㚛/�����N��Dn֨d�=X�e�7Q$���eJ6��
όp���8Y	D����=W���M
���s���Q�l�0�&����Q�2M14�pd�s���F�,~,}�)�)dZ�8�T��v�4s�̙7-���'���'��$	3?ٳi��H*� ɛ|�[6��I�'kP�������={���"�BT@Y�b"דp���	&?F6m�O��D�O���H�	@����,�<���t0Ȁ��:�M�fku�����$�
y\�hKDH%FW��3'�)&, �nҟ��џ`�@��ē�?���~�#�)T>�]r!��uĄ�@�F���'���y��'+��'�P���!�,X�t���~Y��k�2��݆y�>&�p��۟�$��؁E-T���B��蛡{v�Z ���<)��?	���H�@�0	�M�WH e�1�N�wv(���
P�ܟP�	\��\yrC_X�2ĉ�$ĕA -�j�|��1�y��'���'J�	?��Aa�OE�����#�dI3���Z��M<���������;��	�"�6�s�슘�f��V�H�|�H��?����?y.O��a!l⓸�XY�֍�Mm�NB�-D�eP�4�?������<	�O�L��O2���/�\t��m��DU$ɘֶi���'��	h��)�I|R����G�I3��RT�W$1ٔ��%f�)S�'c剒��#<�O�H�B�k��d`2���l �<p��ٴ��#J��m���i�O���T^~�	�Gx��Wg�e�%������M�/O>�;��)���*>x�G�	 ��e���{G�7튵s�H%o������џ|���'x�귫F�X�"<{��S�\�h02�zӀa�6�)§�?qT#ޭ^8V�X"���<��,�-��V�'J�'N��5I7�D�O�d��@���(_F����ł}�83#�2���R�&b���Iʟl�	�"���y��܍	@Jl*`��8Dw]��4�?���)�'r��'sɧ5��Wk�����m �6"`� �ʠ���əsY1Od��O��$�O�*6�r|�m�DFP����A�m�,���䟰�I˟$��N�	˟ ��A��*Ï4h��cW��F��Qo�.���?����?�����<�?9����El]ҥ��5��a��*�,5��'�R�'%�'�BU�T�!�}��A荓'Z��ˤ��9��P�`���\�Iݟ��'�ց�Op�&P*�F�1H
E���c�	��H��7M�O"�O��d�<bb�d��]�}z���zʠ9!��D�Z��7��O(�d�O����"{��d�O����O���#),<I���¯)�ٲ�+��%�<�$�O0ʓ0���GxZw�$�ȡMV�04е�����1"tP޴���1lZן��	Ɵt�������`JP)K�;A�Ar��6a��=���ib�'��b��'��'�q�FђWgӼ��P�I�_^�dB��i��T���a���d�O��D蟆8�'��ɰ:c\TX��@	5�NX�DF��4B��ٴޘ �b���OR,����$�� ҉̎|3>����¦��ܟ��ɛ3W��@�O���?Y�'`r9S#g�q��8�$�j�����}�cG���'b�'5�L��|��sv��]�F0�cؿ%��7��OQ�+
H}]���\�i�͘�+�
����B��.@`q+0�>��L!�?�)O���O��<i�Ѓ閡q�'(t�F�`V	�#fm�9�^���'M�|��'L§9� 
�ǯ]�V6԰��͛�T��P�3�� ���?��?a-O�1
Q	�|�!'ԍE�)p�˗3��y.�ܦ��'�2�|�'����O�����$�|ИU� B�P8PtL�)��������쟴�'�H,�æ�~J�$�����[�Kմ�����&$6P�&�ibB�|r�'c��ݾNPqO�)��@�]�D��a"8�Sǵi��'<剪.��Q��p�d�O��IV�(��^��`
y&��$�P�����z��8���4�.o�����C64�L9S�@��M�-O2��vJL��]�I�I�?�R�OkLəG�T�#��S^~D���.=���'b���sx�OJ�>�1r�צsY�QQ�ԬG���@�"d���f.����꟨���?%y�O\�{�f�Ab-�9P2ii�	A�������iN<�d)��ӟ��@��i<��枂@6�%�7���M����?Y��|�ZYb_��'x��O�}�𫊾DPz)!���:`�lzQ�M>����?������Ծa�tՈ���
���ռic2�=9����D�O4�Ok�����j$Dh�Hj��U(f_�		�b�d��֟��	ky��Բj�3�EG�9�!iFjՁ��!j�>�)O��$0���O��d�7Ry���H�\=R���K #b����5���O����O���^���3�Fa���{���DlT�?��4�CU���I���%�ؗ'0~TaR�'X���Z��(���L�)��:�@�>��Ӗ�6�'�>l*9K|�gM];I�ָ�ڝoRp��"K�@��&�'��'��I�����_��{�<�A��9b���i�ad<6��OPʓ�?�V����i�O���k,��D�5��x�	AS�ǵt�'���'�����lW*�����E�4B��IP#b�$�x@��'��	ϟ�w/�̟���ܟ��	�?͔�uWaP#̴BU`%=��t*�5�M��?y �1����<�~bЎ�(	&�5�� ��8�$�b�ئ�Cv���t�	џH�	�?�����ȨFQn�����d5�S��\%�6xm��9~FͣgC9�)�D������C��(�QM��B� P��i���'"��� ��)�I�l�dm�8O��,=T��)������'�
��.8��O��d�O��uk
�Jy�e3tI.D����E��I͓u�,��M<ͧ�?�I>�;��	�m��'a��*u��ts��'(R�*C�'7�	����	��ؔ'������=W��qb� ,��O����O6��?�*O�͏!Y�1����"��cԁM�Š�D�<q��?�����䉶r9Χ��m���D&2]�0�d�] ��L�'&��'��''削F�Q���m�v��iG"H8	SO9+�굱�O6���O@���<�b'DSb�O�=
��5�`g�2q̉�E�m����&���<!"B�:�?�J?M��֘|�F9{!��f�����y��d�<��i��� *����OT���\�#��9�P�*�fF98�\��xB�'q��)"�i�y���%H�5�F�����q�f4p�i��.}�����4O�S�<�S����ݦt|���H���)c�*?7F��^����#��1J|I~n�o4X�N���X�)#ig��"bӜ���%F��e��䟼��?e�N<�'@�2��	"r�ǈ^?u^��i��(���'��^�'?��pz�H2t�R�z�Ċ�6�m�a��M3��?��'�H�מx�O��O��tkC�%p0����3��AZ��i��T�d��T1��9O��$�O�ЭP�*ݸǯ��7r�������q��l�<�e`N����|*���Ӻ{#��.ta�]Rp�hq� O�z����P�����O�d�O����h�NA�u���3�-O�ص���Ƕ�'��'>�'��	�$�h{g�Ԉt���q��9\�)�QG��� �'�"�'��P��RT�����I��+�N���e� 2��\���9��D�O���2�d�<q�jʸ�?�t�Q9z�Ѝj��2D(�5�ŘG�'#R_���	&eVV��O�"��y��=���N܆�0
��4��78�	����>Eb��e-?��C<cU:$Z��S�7��J���ʛv�'��V��Bw�����O��꟬UY3D@�e��ySg�F+dP��P�-�k}b�'4��'N�,�'�b�'	"ӟ�iS�w�r�ę��n�$�M[+O޹�t	�ᦡ��؟<���?�+�O뎔&Z�b��
s5���L]fڛ��'CjV��y�L�~Γ�Oqpрd �#a)z��".M ��޴q8"�A�i�"�'���OĎ���D�pUحJ7�վm{���'�!G�!o��b���	W��{���?��-A�� s�2LtM8�1M��v�'hR�'�z�)&&�>+O��$���j�C�c���0R.�A@ĩ2��>1/O���g��������֟�P�(�#d�x��ܕ&��쁐��Mk�f͎�{�T�h�'��[�l�i���BMy6��0Ç+*��>��NA��?y��?Y)Oj!9���\p�A�fN 8�b�2%�9o�8�'{�Iӟ<�'z�'LlHO�Xu��qΑ���,^�ؼ�O��$�O����O��h\��Z�6���S��ä<P�`��Dd6����i��Iӟh�'���'L���?���������D��Z$KV�S53����';��'�rV�hj�ɋ:����Ok�gt�pa�Q�<�j�!S�ſrp���'0�Iٟ����0�pe����y?� :�I6�[�$]{�j�? A4�#1�i���'��I�H�脀����$�O��)۴_lb�1��j�T���ڌu�v�'���'�B�Ν�y��')�	nz���x\��)�]�� R��̦e�'����2ed��D�Oz�d�V�ԧu���!� ё3�I���;�L��M����?�&n��<1����� �ө1��� F*�F�ط GW6m
�Ho�֟���՟��Ӽ��d�<Ѵ]X-�!��(-tu�7��).���d"�y��'�B�'����JT�1�a���� �-*G(�m��	؟�Rt����d�<����~ҁ�#nS�� O -Y����M3,O����f��?��	��x��#n�n��D��&0�@�A��0�Iaڴ�?Q�&�t7��Vy��'���֟�ز|��܉��	H�.q�uJPA���Eϓ����O�$�OH�3`�M@�� ~�Z5�*����!���4}w��jyR�'�����	��h�c�'�b����I۲���Y���pyR�'K��'��	-}�"a��Od��3���@[H A�iƦ�@�4��d�O`ʓ�?i��?��+U�<�gh�
/������
-�52�+J�?������	̟��':��XaΥ~���/���02�X)�t���a�ʄ获�M;����d�O����Of���?OR�'���c�X4L��I	�d�9K�F��۴�?!����@�\w���O[b�'��$���i�
�X'.����ڇ(i�꓀?���?Yǯ��<!���D�?)�灨�"� 0�F�'嚭��g���Mh9��i�|�'�?��'Q��	�r�m[�O�V�`�S��˕5R6m�O���I#Y��$&�$0�ӱ;9��c�-Բ,JR���l�= 7�G�L��nZǟ8��şp�����'=�@�M��}#&4�q�	)���djӂA��<O��O��?)��;a�L ��ի|`^y�rڅߴ�?q���?af�L�'@��'��Ċ;�I#0�֗ ���� ć&I�&�|B�?r����D�O����EQbFB�9=�8�"jɊCpo������G���'�|Zc���+�D[഼{��	}���Oт�5O@��?9��?	ɟx
`əa��Y���P�jQ�� �͌; n�O����O��O����OJ�/	�r�b-�R�&8u�$��e��+���D�<a���?I����	ƾ-{��A&z�@��] `!��F�J�O��d7�$�O��$-W��dG$�E1&s.� ��_y�'���'��X��{��E��ħaQ0��0J
���v�Y)��ʀ�ix��|��'y�	�y"�>�E���O��ݳ$�ݼu�@i������I󟸗'��5�b*�)�O����&RlM��GU�I ���\?AH'�4�	�����ퟬ&����L�����F�~���!'�ݦ*4�n�^ymϥq307mWo�t�'���l3?Q�7A��[&�U�j�l��#Ҧ��	���"�&�͟�&���}z��� 3�T�z��N�K���ɱY��	xP!���M����?a����x��'L�f��̪@(Wh]K�d=�+���w��O�O��?���7wԔ@���]� b����+X�;GZ�i�4�?��?����E�'B�'�����N���4LR>&��D+�2+���|�X��yʟ���O�ā�1�Р	�jE���
�⑩?��`mZڟ�������'"2�|Zc&��##  ��X����S`a(�O�h2��O���?���?q*Ofi�$�1:�@Z��S�(H��D
K"d$����̟ $����̟X�p@�꽱 ��c"�4�7�6a#n�IZy��'���'h�IdX���O[ �G�Kz �x����q�ɉM<������?���.Ȉ��u�]���<X�P�W����R]��������zy�j�J��� �V�J�R���ǉ1T@������	n�������4*��=y��,H�8�qw�
'o����]��a�I�P�':���!6�i�O�	�,d PqsU�� a*ʙ����{TX�'���I��yb�a��$���'A����EԞOk��%��u�4oyyB�ǲx6�p��'����'?��F�r���B!/�vd��/	B}b]���I]�S�S�-����1��CP�%�`���q�6M��w6l���O����O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J 3��b�h6��Op�d�O�����D�O���rG^i��	�C� 9��;��LN�'sb�'	���b��ʘ���ͣS��Ԛ�lT��!0$ &#�f�'��g�/=��'�r�'���'yZcn�93p��+7����Š
I�dߴ�?��4����Vj�S�g�? �HD�P2զ�)�,X�3��a�i.Jls�zӴ�D�ON�����T'��/z��e"��
8�>��b�3d��(�4'$)[���Ϙ'pb��Q�
�#�ݏFmʉ#F�N-Za�6M�O����Oh%`Bk�<�.���d�����`R�hM27�۠a~8���2��'�حb�	.�i�Ov��OLR)F��`�J�4{����ئ����S�R)�N<����?�N>��~�Z��M�z������Q�c��\�'"���y��'��'��I�����OI-r��(�Tnν]XX+��ē�?	����?��*<>�IT.Y^�h�T�P��Ȑ����I̓�?a���?�-O�yRB��|�e��9��x�g�J�{]\��du�I͟�$�`�	͟�hp �>Q0��6�����P�=x(@��b�r}��'�B�'z��|�b��L|�s%�1c*�ɉgvNAPէW՛v�'u�'b�'".�s�}B�>�!Qr�N( X�$@V�A��M����?-O2훐aYM����(��3aMǋUTn�����D�)J<���?	��S�'e�i��a��)��K�C�*pCfEZ�d˛&\�| !���MC�\?E���?��OQ� Ą�?���ۥ
}��ib�'F ���I�E�������ø��q�<Q��&��0"�6��O~�d�OT�I�[�e�
�AO!-��Dk�*��(þi�Q��d$�Sɟ����(&EpKG`اI��Y3��N��M���?��7���&���O�����p�I)5����t��W��c���BK?��������r��ҳM��Ha��M�)@�ՃqDE��Ms�]o�� U���'�bP���i���G�-l�����h��/H��Ia�����t�Ġ<��?�����$^*1�L���"[�Pɰ�m��9�0 B�_}2Z���ISy"�'�R�'�� �H"a�@�B��^=�uȅJ?���?9���?����V���l�'z�6���N�4�^�У��$V�&5ldy��'��I����ӟ�B�v�d���`*�b���l�Y;�*¥����O����O,�Gw^=xER?y�I���	�
�.�*� \譢�M��M����D�O��D�O�$Q�?O^�D��x�dM��2��
�&,'�5�lt���$�O��=��a�P?����H��1W6 ;MJT)v��>+�p"�Ox���O*��ʃFD��'��?�"��T0t����3��yh��S)g�2�1��+�i��'���O]�Ӻ3�#h$L:�I��δ�!�ɦ���ğ��u�q� ��Zy�I�381 �th�J�~t M�.`�m� ]7��O�$�OR���a}2P� �!���h��*��C%U��u�ڑ�M��<�����$-�Sߟ(���H�!dȟ�P�x�hʙ�M{���?��f�=�wP�ؕ'�R�O�I��*�55��2�*�%�@�i4P�P0&n��'�?����?��
#)
ܕ�����JܝH�6�'�hBo�>�,O���<����Q���Tx�gE�r�AI�x}�E��y_���	ߟ�%?�B��>UKpS��K�:�JH@�ꐃ^��	H�O�˓�?�(O��d�O���K�>m9	¿��p!�R3p��z�<O&�D�O2�D�O��D"��a���x�®B�3�$�(&�7rQ�J�e��M���?���䓕?�-O-���iL��P����o8�!
�4��L
�O���O4�D�<�aiF�C����Ps��T1��2���7�V0X'���M#��?q���';qO��(!�&��]��U)�ZLX��i�2�'|r�'ª��q\>�'��T-�7
���D��#㤕 5�P�.O��D�<!��Ko��u�+��A�5#b�ܰ*Vnύ�M����?Ap����?��?������?��/F����^UZ�q��(.#�o����I�"U�#<q��4k3pUqF!L_��H��S��?����,��s���0=	�2�Fm3��V�"���[�<��`�5?���ԭ
�.3Y��[�0k�	S� L
Aɂ�J���.I�թre�?+9�t�U��2t�2Q^�$C�����U01�`)��DV=��՘&�>LpU�����ZLuq��X�2P@�P:%�0��a'Q!ܠ5X�� *d �#���[4:��g���Px6�Ĕnv��k�
�?���?i��Z��.�O��D|>��A(V�S[��	ďRI��\���N�8C�	I���P��͘�-A�k>����D���N�� �D�e0�� ��ph�/T�.NH@���Φ�#��9-$!4�E���@J<y6hFW�¨넅R0��[2�G7J�(H�	��TE{2���M��A�14Ԕ���bM/'!�֟pt�-;���<<���Ȅ�p1O4!�'��	D=�aB�O �]�2mb�0��+l�$1�V5^`�$�O( qi�OH�z>�I���9'�ڝ03�خ�~��'�2�Ѣ�"o^ � "O�p<I&��}��� ��K��Ӆ!/�k׃�}�����a5H �x��]��?�����d�am l��/�;M��&T�	�1O���DR�
n��0��F/�r���9�!���!۲�
Q Р�0k��~a"��̔'�~����>�����	��U����Q�KG�-�샞q�ƼP d��X<���O�`��)d�AI��ͅ0�?�O*�S�4mj��#��#�!��o��G��'�
7	Ҋ8�i��  7A�>)����'`�n���՟5H��d�)}b���?���h���� ���R �\x��נJ�<(�G"O�9rǃ(l%�1�դ�,��P�'�#=i��Ɉ!�Ȁb��x�0/��W�����@�I<M��T*aŎ����	韄�i��F�c�N=b-���@E�_t$�A�^�L���@�b>�O6�@��*2�$�E�a��e��tc�+�O6��Ɇ�и��a�H)���D�A�,Igɣr�������$ʒG��O�ў8���?np�⠅�l�ZCe=D�7e��(�jm#D$�.��kpM??!��)
/O&! #�ǰT��<�1�D�9.8��K\>����	�Oh��O��D�к���?��Oz�Iᇏہ;Zd���̆�]�D� ����x�k�&ɠ�x�E�)8������*F��@	�'Ψ��vC�3H��Dާ���@��!�?��o1t}B�N^M8��r��	o��)�ȓc��TKQ��p��(���X�dS�`�<I@�DP��l��t�I2Y=L)z�J֓x`>�kƪ	#"z`���<�`����	�|Bq�����'����^��YK�O��1��$O��� �Ĉ3m���0e*T~�1���Y:�x�C���?�N>��X�C��t�!��?D�����J�<���O'	���
�o�\�z\@b*�_<y�i�x<YӣI�_X8!B�P�"�,[�yB��&�듓?A+�������O�����0-q��;1�[I�=1�	�O,�d�*$W"����S
#�:\:�f��$UJ�O���*���Ɉ}�.��v��;F,�'����+[@x����٘*�>�PBI?�/2�X  ���U ,�LG�<kD�'�F0p���?1����OJy8$�D)7��$�p���F}����"O$�ڷfܫy��E�D䄽d2	S��'�"=��ɝ"i�)S����>\�V�M�.���'��'�H��)N�'K���y��N���8�cd�+ag �*�C7.1O�%K��'�(d`d&�/&�v!�eGZ�xM�{�� ���<����;&�p��)�="6�P� �.��'1�P��S�g�nM6T+&ܠD�!�kֵhC�I�9r@���F7w�Q:�+L���ߑ�"|"u�T�Rr*�c�I��u��c���72�+@��5�I��p�	ݟ��_w�r�'��	:*��:V&�#����1Ό@!����Onu[�/�B�6�{t�~���e�NM���'~$�G�֨E����#��Q�� �r�@�?1�Z΍�wE�C
z�3��D��ȓ`ߤ���v�9��ZB
"�I���'t�ŋ�m���O�<��	�5�L�5�F�3E(�%��O���� �|���O������'�W�+JXy:���2'�4�A�/��x�E���'[jE�w�ϭ���� #L����<�Z�	D�ɷM�x�It�˵{��HK!\�M�~B�I�( 8Z5�V�3YPc�x%�B���M3��A��0�⦭4 xٓ3��P̓UZ�h�#�iM��'��,s��0�ɯ,�|��6dI7N?V`Sb�w�^��	ן4���<���D�!+�@���*u,��P�o�a:2�Ex��A��uIJ!�ߎ{|�Id���ɾ��<�)��&.#x�[��� _,Ż��Z�;a�C�I	
��ȡ�����2U0!M������r�'�Ѱ�+U�4}�<�u듾w��J��i�B�'��n�[Hؠ��'d�'��w��!!3��:��Ų���E�<Q��i� OP-�P���_M�S=*�1��'Yl��RP�?���U)�I&�����B��	��ȇ�j�T��DU�����X�,)	ׁ�?�`y����'��"�i���'^��C��d�'_��'"��'t�T ��|@$"��F䰔btO� �4ƍ�EFe����r(�8T��p1��d^}rX���	@�t�CΙ^��q;5!̐\I�D0��şD����L�I��u��'\r�'B֙(�0f�pxD�63e��cT�z!�DD+W�,H�t`�]e,+㎗�(�4��F�y'�ؖ��h؞��5� "l���5�ٯnx�X�Q$L�R���d�O&�&���Iɟ,�?��_�K�
M��&�Hwh�`�$�]�'?H����0I"r��#�pd�%Q�c�6wfx�O|\m�Ɵ�'��*�ê>��[Q�5B��D��l�@���Z�,�i��?��b��?������n� ;B��#��h���#V�6g2��S+<�,��K�<����9%������)?� ��D��:�p�	�D�6z���b�1�@x��'�0����Uś�>)�N��$��Y��҇w6�=�� r̓�?1�S�? ���CƘ*
�D��jͩ4�Y3FOulڮXq&��$߮6D��RE,E3A���IG̓�MG�,O������v"N<A �D%�$�P"O�e�ņ(yL�����15���"OZ�r�$��a8�b���x���1"O^��s��PH���	��dF��2t"O،���^e\4\@R�ѩT1�t�"Oԙ˵B)s"&c6-��':H@�"OV`��S�eX h�Ǭ\Cx$z!"O�<b�E��3��\4��$�@"O�s'/�b|	��j՘||ȕB"OT�"�ч�$z	Ɯz�)c�"O�T�G.�k'd`Sw�;<�v�t"O�Rrc+C=P��Wf�)��u"O�a�'j ������I�6��"O�أ��, ���)]ְ�a�"O0X�H�)�(0"�b��X�.�+1"O* �H�.0�%�Uo�"P֬��"O�,�S		 d��W�ϮX�"O���0$�7/`�}r���"� �a"O�]��C�$<�1��D f�2��T"O4�$f ;S���9��o͊�"O�Qu@�)W�$�̟\M��T"O6(��mE5Q�d@���_�7O��!c"Op�m�%K�(P��W(B�y�w"Op�ǁO:䒼�"�B�����"O����ȏ,v(1��O+/�nXk"O���d�V4V����wLJ�#�Lec�"O�`���%P�� IE���X�"O�5ۂH�.m&A�e��4+�8Yɦ"O]�&���u:�ad�V�z��Qv"OhIg΍�M�:a��]'f�D�D"Od��+�K���%��
K��2"O�� v�
+/Jؘ���٢g���0b"O�p�/A��MJ􉍢~��̱�"O��Rg��
�p�@E��#'�n�$"O���� ��Xh������+y�]��"O��#�D�'��S�PE�x�a��8XD;B���t�/�g~��ԗ�tqr���6G��v@W�yB[�&4�&c��ID2�9�. �wL�e��aCn:f���)�����^�*�@Ra�L{bͅ�	b�J 鰈\�9���ɣO��]R�E�d�zi���)K��C��/�(ؤ��G���",o�zc��ӄ".k�j� �#�'TޖHB��)��M��Q�S2���a¢�ys�Plpeh��A�`g��R�,ۚ3�q�'��@3��0�^�Z�<�7�*$�j2D���[�3��+0��YN:!��͹zr�x� ��;�����$Z9򜃗�/vȉCr�4:=az�Ȅ?���s��y��C7L� �K�^P i����y�&N`�p}	�jL�fr�-!��'�v%2%-#Ed��A��IK�N@�1%,�.����C��x!��˨[D��EI2޺ЊD��<�����D\��'zq�#|�'��9Qe��c�J�����y �i�'j���ŝrb�����Ml8s#�"�N�i�F�0>I�!I�}�4�E�8x��D�T��И"l�	됩�Ek��p�i˝hٮP��`H�M8]:�(D�����&�R�Ӂ��	�LXj�*��
�\x*e�˃.#~�Ă	>R���j��c���X�o_P�<A�b�74�� !0�U�/
����J�<iF ��V=� R��$!}�t#Ch[�<��NѨN�كa���5��h�L�<!�,�0?�`(��D!cT\y!��GR�<)#� <�j��D��Y�a��L�<�tE�>,�5�A��!�di�'ɌK�<� \=K�?l��ّ�X�����"O�aХ�N�Sp�%�I"p���Ƀ"O8aևI�[~��#��>���q�"O�]�g
^�����w��A�Q"O��{dj�:��P��>�j�C�"O�pf�-|!�,�3�_�����"O=�p�^8M�R��f	�	�|�R"O(ě���m^���V��4 �����"O�M�2�	q��Y�b'�"ai��� "Ozܚ���8�0��֏�!gNr"OdT�Ջ6ɞ�Z��!6(:|zW"O|8����"��;p4�U"O`5!��S%`�@Han�Ct��0"Ob�Z�GX���1G(z����{�!��%A�����#cK���n��%q!�Y$��X9Ff��:8�����\W!��ƞ:��1��ȝS(n��P'� ':!�ğ�#>2����ǜ#
���f��O)!�D�-0�fH�Dʅ�;Vnd��,!�_(���q���>eCr@	ep!�d�M��ˡkI��D����� ��<����'pB$��!O�P�2�b���8CF�
�FL��I�=ƪ��aًD'����Ҝn�z����&0��' ̪����z�)����w�ъ���^���J��I���p0!�I5x��q��2Vt�O��2�4�)�.�ꎾ R @T�])��'�=@!�)�'v��CQBʀ8��TQ�Q�7\T�!�C�T��'�D�G�,O\��go�7���BEQ�Ig�D�C�O��A�O�צ����M&�p<���ԤJ���a�M+�ʄq�(�y+^l�p��=Q��#?��&�B���qbB%<~,}�ʂ<�l�UN�.,$t�c�3�D�l�$u�g��`,,��C��m�ԟtȠ���?�@9�Y�!��y�D剥Ld��3��;�`y4�� fe ء Kc �-����#ȎbR�]��e3
�|O\��S��cH��S	il�)b	S,X y�̉6[D<����G��M��	$g��)��@�`�ɽ{骰ZS*-Č8��I^����u%�� EĘ�[�`֝5fw�EyR�]yh���A�&�2�5�B"����ƈ��pq(�(��\>�`J<�T�A96}�Ŭ
�\z�)�#Ư^Kv�:�����	����|�pݨ1l�s�#<��.!F)bAS@��d�!&�\�Ed�Ȱ)�c^�+��f��O$��Sd�+pL��i����V�6d@�D�I?��O�>��-υN�����W�:��,)p+G�T�X�u��?jq>T���iP�>E;bA��U�+6!J�eF�Q�'��0�%H�M�Bs��q��ϻS�MЗ@њE۬ԱF���Q{�!�y�4�Ko���10�w���S�v���ω1A��lq�G
U+ 4���'z��d�6Wop�R1��"٫&d�?c�@��'�3>�t8qNў,.�#`)�|tr���A��͉b�_9�RO���t�7Jz9l̘��jM�L@�O
����֬)�:���L�$Ty�#<�*�6.+�����][����-�|P>���!
Ypu�� 
��O����QTܨ��ڇ�:�"@Y�擛>��P(�	̒E�7Óc��p$��Df��RTjA�4��D���I1��DnV�s�-��_2y�L���Ѡ.dft;s�"A���)�S�yW%<����A�T���e����5�*B�}���	���a�X��;��99���d>yf�т��Оs���_w��D{���1�Ä@[;Q�e�M��t����'�z��/ڲjB������	F�9	���.y�x@*��#�z�\�)�p���r1�Ys�X�����*}=S)�f瘸r5-���1�R��1A�b�	��%����ZF�R�3�\��J?����6 ��`�bS5q����u�#�ts�MCҀ�2"&uS'h:���45��KSi%k⎐�R�5N�PM W��TUP� �oe�PD��O�Ă`&N�"(�a�2N��VІ}���OZ4�ʔuJ<�¶��%�0|!L����1V�k$&q !Ц�Y�#ɅX���f��� ���I,R��x���SQ�!r��^1��b�(�������K�¨�ם~r��3Wx�R��C2E�I �h�\z��Gn\!� 4��ǋd��p�cEBæ(y�M�3
��5pw�ÜZ��Db��C����^����*Ҹp���� 7d�d���2qhNt���S	c��E4������Rg��*���(�NŊ&�^+2	UV]� �D���R+ԭkt��Q?�V�>����m�fś�������#��w�<Q��/+��X�㜘�>�xd�ͦ���m�{���5��U��y���T��&M��3U� ��=1��	!8&j��D�g($@;@��KT�R2C���Ԙ�F24�� ��Z������W��8Hz�Ѓ��_�X��@c� �Q>=I��Ҹ$����*"��J�+0D��� , �U��ev1��a ��>���'�Ȑ�q�D�i@Ο��|���.o���x �'P
8l����@��,���,{�0�P���B��"ѡD1*3t��w
RQ7��=E���s����W�9���1f��E���G}�`���nً�dD�zdQ¡Gcr�kea���~��9b�8��4V�x8��IMƖ1PK�u@��	�j@:Hr6�)�)r�K	�qH�牪s�q����.Che� �ə\�.B�I	U��@sgπ`� ��F�/>��'� a�aA�Wl�k!j�X�S��mC�\s����ګZs"l�$�3�p?�aLK�	�b�X�R0i�:C�Մ-G��Zc���a8<%��0�)���ґL�>?S��:tj�,S��5!���ͳ�%�n��VV͑�I2'J�zA̀5K��'����əSN8�kF�Id}8D���I5X;�mbC�"�)ڧ~:�8�߷,n��˘%u̸Y�ȓ
�\zu�G��P�C�"W'�ႇ	@>���	�E�Z���G�hND�+a��
�'^�������"�R���+�,q�� ;�'fv�b�$]�h����e�y���dF"X) 
R���'�lQ!ІCZ,r�*�1!���}KS� � �4 (`Cb$9�'��%�0ɧ=ɧh�<��%�*����W�U�l��"OƩ�l3�И:���Vu��>q�]9 3���
�Ƕ)�G�Zj�F��0���y�@���2T�L<�&ܑ=b���L��^�Jĩ��L��=��)k0Hɵ�߈xЮ�	��L�M-�mG}2��X��ȇ�	T�Sឱ���ɫi,��mH5V�!�$��2��W�XF��cs	)Y�^���r�x�rrG���S�O���� P)p�z�C�k	K�f��'�&�@s�O;F�F)���.G����L<���r)),O��Sv��(*(��	 �$4���U"O@�ʃ��S2���(�ho�t�f"Oș���ۋ"dVPr��� ~�P�"O�Q)4�[�p�A���Z�$5�"O,0�)"<q|�*r�� 9�D"OV�� _��P��BEy"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��   �  C  �  �  �*  v6  (B  �M  mY  3e  q  T|  :�  �  �  �  L�  ��  ̳  G�  ��  ��  �  ��  +�  w�  ��  ��  ��  x�  �   [ � � ! V' q1 ?8 �> �F �L vS �Y �_ �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�'��7mL�2�p�)2N�&g]��*ϓ�Zφu����P�ݴ�����'�¯�'��SF�=�����df���'QVL{q�i��I�|�A�Ox�\L���5�C76���v�M�+���<	����7�'�l�� ԐOE�I�`AͶGn��aQ�i�0��y���ڦ�]!¶Ex�C,v�tX�کk��d�Iԟ@͓����ʏA��7�a��`��q�L�I�1�0��ǫy�͓o��z�����'Z>��$�R�1�&�8�o0Q'&���'��I��#�MӲ��Q�
wp�� �.2�l�3�\���ܫ��o�>���?��'��	 ���r!�G�{!��h�Č3���?i�ND�f0$�|j�n�O2$�,��H�
H�48c�+D�`�*O"˓�?E��'0��sΘq��a�L^�ke�Tk�'�7�M��	0�Mێ�O���$ƪa-čp��N�5,z���'���'��øST�F����'_%�T��VT��se��<3� ���K0��-%������'���'�2�'���s��y<�qw�C�]��M�!X��޴W� ����?�����'�?!��?)#�l�e��_�P8!�Z��	��M��i�O1���i!SiT%S�X�I��H�D錍n^ZDb�0O��д���V���@�d�%XM����W�0���/L���qk�6�.������	�� �����}yk�ޕke��O����ݪ1��S���s�B�qR�O,�n~�s��I��M��i�h7�Q��n1YP!-�"��ӇQHi��_�7�*?IT`A�J�X�) ���`�=�]#9ebԛ̊5��R��I]uT�	���	����	���D��q��`�#*�Fcj�9�
4��� ��?1��LśF�$��I�M�L>���<R��x�`[�aB����jY�'��6-N�� Uú�mZ{~�MK�y�8�CP(�n7�aq3�E����c����`�fS��+ߴ��4�����Ox���;D	��
�2�h$�����d�O:�l3��%Њ���'^>Y��M߹e��Ͱd,�;}=�@�??6Y�H�	�CN>�O�� hT�K�`���\7����rNϤF���*������޺k���O�k)O�չA�����!X��]ۥ� LFn�D�OD�d�O���)�<�4�i��y1�D�d�D]�3�_��~��r� ��'�7;�	���s�8��&��9o!�})2��"��|B�C���"ߴ_a����4��$�"!�q�'��S�z��`�U(�1>�j���� `��$�ߴ����O>�D�O���O���|2	ˏ��L���ًs݌�@��
?כv�CI�����,%?��	�M�;e�r��J��dtx����$4ȁP6�'��F@2����FS9�4O�uC&�ՀL�=��E�%�:u(�0O\	`���?	2��<Q5�i��i>��I�17$Y��据c�Ȋ욐6u��Iß��I�8�'1�6�K,ZT�$�O����T� !+�\�u�����ۭ@7�㟰��O�5o(�M#��x�M��\4��B�g��H��.N����'|�t��HM�H�S�O�譻KiT���2�?�Aǂ~�(�(��!p�����CR��?���?i��?y��)�Op�:��D9I����$�#0����o�O:�nZ5������ �ݴ���y*E'6 \��C���6,�Sa��y�eӈn���M�����Mc�OvT������7{R��0tj�Z!�m)R@ª]�˓w�F_������	��|�	��D�15�P�`uC�~JĤ@��iy}Ӧ��0F�OD���OH����^*"��I��
<�P R��S#y���'��7�]rL<�|c� .o��Y�!JT�}��҂Ȃ�WҎ���}~�%Q#K����7{?���M�-O��CE�?[b��6�,�,ȪAd�O���O����O�<QF�i�H(��';�P�dMU1:�Ra�N��J��'6^7�!��1��Ėަ!X�4K�V!�+zuDQa-��(Cդʉ�rAxW�iJ�d�`��TY��Ɖ^��t@�:��ba�� ,uJ�dT >���s�H����?OD���O����OT�D�O��?1�w�� `��ش���qI
0�m��?q�i�N�	��' ��'#�'б��%V7G%=j�EX=m��)��A}Ӿ�N���a��i�7l��6�=?��N��]N��87#Ƨb3�d�G,U�Q�
a����OP|".O\ynfy�O�2�'�� �<'{❑�n��&��uKaτBqB�'��2�M����?���?��'�� �Ƞ)�R�ؔfH�s��<�a��<�������O�7�K�A�´�%
x��ӏ��E�@��DB�N��TZP���*��'�T�]
+�\��;y���yW�� 7�\l����8:��@l=c�"�';��'�C�����aF�I��ugjêkZKT�WN^����ZQ�R���':��
~��_�擅�M3������V�F��em����W�<�6-]��B�˦m�'�B��EB�?����(���  0P��[����i2�/���'���'L��'���'���?k`���e�t��k�>���4&��(@���?A�����'�?9��?�;��5�5 d�[$�F���Yc��iq�7��Ȧ)���O��`�p�i��䙯`� (�P�ʿeF0�q��O�P�������k��k_�ʓʛVW���������p�R&��,yʔb�e[ןd�I�����oyR�h�R��C�<i�w�Z��o��F��W��?m2�3������O��'a�7���޴����.;���х�֗}�Q�mI���I�/��{5,��r&.�\^���b�>��%�?q�h��*=�h[C��R,h\���H �?A���?����0X%6��̴e������O���HR(3S��¾{亱��L�O^�o�5F�版)(f�S�X�'ݤ��O�;��� w�\+��|��1o�╸0�'w�7M�ߦ�Sڴ"��(�4��Ğ�h�����h="�1x0dB��� ��{ ��O���W�e�����'�"�'@��'V�	{D�Y�X^B���`܆!H,ը�V��)�4G���R�F��?����rƁ/�?y��y0��'Œ_A�i��f &H��QS�� ڴmj��	b�|�D����7����ώ!��q���(Mcw�����01t]���C��Ӓ޴���F<@�f����dRH�p��@��$�O����O��4��V�&&�)q4���:J�Ua&�M*�z��θ�y��~�X�h�/Op�dnӈ<mz�d��"�R��T"K8VV�ɠ0�3 ~�LoZr~r�B�ZԀ��u��Gź���*��5 ���#K�"T����1��ϓ�?i��?���?�����O~ ��� ܔ
ͱ%@5 *�\���'
R�'h�6��:�����֖|2cʌdp2p�Ҡ�-_X� ���PW1�O�m��M�'zh�	��4�yr��W5��@f����\�ヂ"[D�mk�-�N����Q�?>a�H���?1��?i��@�BƎŀu�&q�2Nн[7��a��?q.O�m7�B�	�l�Im����}>bԚ��,t�&��$�~y��'��V&�T>�b�Mh�xY;D�������+� .B�|Y��C����|��(�Ou�K>ɢaC~_|�ٲ-Ш �$���3�?���?���?�|�)O�xm�(���46
2 ���`t�PA�0?�3�i��O�'�V6��\"�L�7�+
m	(G@9n��M����M��O�HQ%"Q+�rK|J�&^k+2�Q@J�>[�L[�ay���'p�'^r�'2�'��S�c������Mp����*	9�^U�4�@=Γ�?i����<�v��y�h��mc����T�L@t��G��ϲ6m���0M<�|:�@K��M��'��P�U�)�b��f߲���'VZ�����q�|R[���Ο�CD��.brt�cdI6D���UNN�D�	ϟ���fy�
p������O>���O��##I��/�ΡT�%�lmQ2,����D�O���(��*`3�pQ� �����K�+��N����衒ԭ!q�r�&?ɢ��'�r��I�;�Rm� ��)7�ą�E��%�@I�I�0�������f�O�R/��lƼ��c��j�j�K֣�B�R�d� 5�G��Ox�� ɦA�?�;E��0��^@�ʄA����f��sț�OT7-CN[�6�*?q����J�)N���ǪT�F��Ņ65�>��M>�-Ol���O*�D�O����O��:�M�0I�M�C˅���h3è<�v�iZ�F�'E��'���y���Ra�Q�+JfT��Z�Z�
���f��O�O1���rU,ž5�$��G��1�h@jT)������H�<��O�Iu8�dͣ������7�<�0ag���Q1WG�=�\���O��D�Ov�4�n�c�v#�B�bE޻ N@)W@�9�y$lB58W�Md�⟬8)O����O�7��;L��h����60:�#)A�,��p��
aӺ�AR˖����:L~��d�E�v�K�K �<B�"�!j�ziϓ�?����?���?����OǢT�g�T���a�)�v��7�'{��')7�-��)�McI>�aN�7��k�?M���C!�'��6-RΟ�I�3¶6�9?�aN�7l
�U@��$*G�D�BԎrM��� �OhL�H>1.O8�D�O����O�!0'��~v����^+X@�Eg�O
�D�<�@�i���'���'/�������F�<���ě:g�R	���Mc��'U�����O��͚i�ZA��B��4	�2�kǋݐ9���A7b�.��?���'�Pp%���cHt���B�/'�������ʟ�����@��ڟb>U�'Zn6m8OS�xj�e�77C8�(!�5_�D�%e�<��i��O��'��6��x�2�KF��5|���JQ�&Ql�D�e�Mצ9��?���[�
�N���k~
� j<� #4��`BE&���;Oʓ�?	��?)��?1����iN�:������-�x�#�7kўTo�y�:u�'���)����݌� �
/H�JCk�f���4 ��6�'�)�"��m��<q��S#ED�hP��{`X��D�<yD����$������4�D��pĴ���G
�Y���-;~����O��$�O��	��f�ߌ	���'A�
+�Mq@�.qÀ$�cV�8��O���'�7��ͦ1�	ry"��Re�j�ŝ`v2H�iA����;��%"G��<n1��)��0nF��H����1�-!�ʭ�Γz��$�O��D�O��d/ڧ�?م��+f�D��P�I!}V֐���?��i���!�_�,��4���yW�ڃQJ4��e�=B��
�{v�<�5��Nc��dʗ"��7m8?�IH�ju����(7:1��
%;��=���)&&�axK>�.O�I�O����O����OR�钮�T+��(\�&����7��<�u�i������'R�'���y�ړ?Μsd�Fj�ZTId��9Q��c7��e����t�Ob̜����)#�:pYâ�`��-��$�6|8\�2�O<��`�4�?9e�3�D�<��kJ�&����Յm56�
�0�?A���?q���?�'��D^ܦ=��`x�\�Peĩ^�`�N�!������w�x�ݴ��'�z�U@�6MgӸHl���\4Lƌ]u� @�
��l2��*P����I�'����6���?1�}��;՘����޶Q'�� �U�#���?���?���?A����OQd1"��!Pk��b���bc,u�'�"�'v47m;h���&�M�K>�U��=Fc�Ỡ�[�!F���Ǐ.[ĉ'È6�Zަ�.	B�mZc~���{���b�N�"^�u�� �{zz�Y�Ȟ��)�|�X��Ɵ���矠`�:I�&u+�/L�g��y�$^˟��	fy"f�O��+�O�$�|�73: ]0�Δ�P�u3��@~bɽ>1��i��6��N�)P�F�\s�5��LA;j�d���O�9U������K�
4��ĥğ(hT�|2���4<��r`�7<ɴ%�q%l���'2��'���_���ߴ�(�����2��p���W�Q�؍�q�N������?��[��ߴ-���q0��U%���뛁�L؆�'Q��*L7ћf��(���, ��@Vy�f��\��cA��.4�ByYW"�,�y�Z����ğd���\����X�O�H���˛��I��u�	0�l��cSc�O`��O����d���]3����P1y�2��a��YR�شot�x���]�E��4O��1NR.p����������̎$-��R.4��Ɂ�y�\�O�˓�?i��e 4�X`Z:X.�zv�"�����?1��?�+Ol�?�N���ݟ��I�(�����L��"��Kڣ2r��?�V�(�۴+�x"�˚a��qȃQ�Fƺ�)V��2����,���EbT������e��$߈JE:�XӃ�tVddIBJU�E�����O��$�O<�D9�'�?a���U�LL�߈"�Y*�-^<?�rIxӄQ�A��O������Y�?�; �&���	�� �@l]�8�q�Qy���O�7m���\6�<?�`lL14�����'������sy� ���2�<�3H>(O�D�O��$�O����O����2,L�lp�`�"��0)f��<9�isX����'0b�'p�O2¤�60l��CI�!(�-nL��Q��[ڴb��x����P9/� 1L�bT�)g�ڲa4`���G�"k�kC����'��$���'����݅v�`��
өoj:�8g�'%��'����dV�����څŜ���ѵˊ bY�L˰&H<X�IC`gy��޴��'	��h�&O�Op7U�s�P�:�'؝Q�A��զb����k�:�U�����	���IL~Z��Z~��bԫN�i���bY=[�v͓�?��?1���?�����OSz��D��F�l F���j���b�'B��'��6하u-����MCL>�6@ô����_�܈��4�[	o�'g�7-_Ȧ�SQ�flZ~~2m@�i�`�����W�茠�Ð>Ѣl�0H�ן ze�|rX��SПp���ɴ�Ĉ(՚��a.])X�:�I�ß<�	Ky�kd��\�gb�O^���O�'z²�c6 �&\�ȑ+�cZt ��'Hf�$w�F+�O O�	���]{�'�Jd8MB�kݻ#�\��ݵzdy"@��$~�F��B�I�O�qSO>	3(Ŝh!��pQ��l��#��X&�?����?���?�|�)O�o�g �b'� �oh���A]�V�,�A0" �t��6�Mӊ�b�<iشs�%cg��4�"�"�K��{��&�i��6���1�n7�k�����:�0ݱu�O�|��'u(��G��	a_��� ��.5~U��'�I��d��Ο��Iğ���^��@C�<����	P��h��$x6�6�K�!�8��O&�!�I�O�mmzޱzR�Ý<�8:�g:,� ������M���'$�����O��ě�C�F9O̐K�΃��%�t�>������y�AN�BI�I�'
�	ğ4��_�U�Ae�4NʴQc����k�����ߟ������'B�6m�$G����Op�$��e�2�q'�*Jƴ�u�r\��౫O�lZ�?�I<q��>X�lZ@DK�jD(=��jU�<9��DT��bJ��T�~51.Oz�I(�?Y���ODu8�`�
(U�����Ⱦ�P��O��O|���O�}
��`T�B�]�ݲ�L�'��U��;i��g�#[���'�7�/�iލ� �_4m��t"�d�&>eD @,��xo�5�Ms��it)
S�i���O8������"�� �,A���[(M��G޵kzђ�!$�ľ<���?����?����?Q��L����Ѝ؝$���JF���E�%(`��䟀���|$?������y⭎�X��h�.Z }���O��n�&�?�O<ͧ���'Rಀ�qGƉJ��a	ܕl&�V�C>'wL�.O�W���?�q�2�d�<aqű(�B��.e�TڴO:�?Y���?����?�'���AȦm��'ʟ��󭞨]�B	���ΘI?5K��{�d��4��'�v�q���D�O�6B(�z�� �d�!c�����p�Ǫx���� ��/��S:�*xyb�O�h�Z���⠏�{'�hï
�y�'��'�b�'�R�ɘ/W�<�9�lQ�B9�%H'e�����O �Ć��5��t>}���M�I>i�E��s���i�L���P���'��7m�˦y�S�x�>�l��<�������'��G;x����X?&,[�E]�RwN�Ś����D�O��Oj�D��!�*���{0̜ёJL�p�"���Op�/���d�z���'mV>�*d*�m���R���+K�@��!*:?�P� �ٴ)��&;�?�	�/34�Fԑ��_w-` e"�`��$���|2���O\�+H>s��*"s���g��U� ��N���?���?���?�|")O�l
�����ΠD����̱oqj�pt��Yyr�xӚ���O�0nڹIu-#!犱7��QGb
��2��ܴa&�v7C�6��3���76��~�Ф)p֐��b5]� �7�T�<�(Ov�d�OJ�$�O���O��'.�ָ�0힎o�H��1(��(��S�i������';��'U�O9*`��n��e҈0�cH�(,��r�	̱q�&-n��M�x��T6G��<O��{��o%�1kB
]����<O��"Rb�3�?�Q�(��<ͧ�?��	�	�`:c�_�}_��g�+�?9��?q���dG��ix
Q{y�'��)�;Z2)�� �8��-�d�t}��~Ӵmn���@�I0���U<�[ծ�%#�u�'&�ha�17FL��� ؟d��'	m��J�j�nL�6Bɓ<�$]�c�'�b�'u"�'_�>1�I�^���J�O*wdA�D�']�(�I��M�Cb�,�?�������4�t�y���u�Td�%!F(��8O�l���?��4!!�"ڴ����YFb����Cu�	4|���T-�)82Hq�&7���<���?���?q���?�sV]`	��K��0��7O����ަe��-�����I�%?�1aN�R3-D��j=��ƌ0N'6�8�O�=lڻ�?�L<ͧ���'<n�e�#�]&F�3EM&#��m������#.O�dj�E�?a��1�Ľ<���̾a[����'Oq��Cc ��?����?����?ͧ��D\ͦ�[@/�ޟX[��4����-Q<A��.����ߴ��'��˓�?���M�4[z-H��4e����
�Y0ܴ�y��'������?qZZ�����ߥ���ɺG��Df����R��}��������	���	������JQh��H�7u��}��D߷�?���?�־i����O��LqӬ�O00)@F/;��[�k�� 5&��S�ɘ�M���i.���C� ƛ�=O����zd��rR$qa�hb�źa|̚g�X+�?�6�D�<����?A��?����j;|E�⯋�@�dP�ҰB�����4�'d�6]d]����O��|�`��. :�����/8���g��v~�J�>� �i�d �?E��!��>��x�*ހG2�+����jSO�"-����i�����$�|���;.�E�9G�R�'$VB�'���'e���Y�� ݴ ��#�@(NɎ1"���wG}��KĠ�?���O/�V��J}Riw��1�(X	C�e��h]	U�����Ɛ�%;�4?�$�B�4���ى�i��'��S�E��{�$��V� �����9Ќ��qy��'���'�r�'��\>��E΋W9JX��/�5Oٴ���ψ��M���	�?���?yI~��r������L�9ToN�Y.���eaC�B�i�"����jL�Q�g���	�'*)Ed͕���G�׊2�D��#PR����'-z�$�Е��4�'VfPr:z�<±	�T���`W�'��'��]�� ߴ/��̓�?��\�b�� `�0T�`Y�+݌{fZŋ�r`�>�&�ih�7�n�ɯ|����7h�m���q���⟄q�cڛ[B�'+7?1�� � ��W.�?����=� `�MX�r	�ț�G��?����?9���?��i�O��y����r��8�VB�G�"�~Ӽ�0"�ON�D�ڦ��?ͻzz`!�c�6mQ@Ff�4&�$8���?q�4`f��,՛gs����3lZ�t��Ɏ���:w�ʅr��x*�	#���$�t�����'4��'���'L���R��6+y���Kn�@�V�\h�4>�6\����?�����<��Z�1@ 웡pHP��a)U5/��|�'7�릅�N<�|Z�
��/��a҂ex2N��U��0�����~~��={
m��;|[�'x�ɜ(t��7�Dd�H�AMN(ޔP�	ܟ����i>U�'��6-N�AK��d�.Ep�Y��V���L�%[I��dXަ��?��W��;�4����iӨ]+-�=�\h۠�%���z�أ1��6-r���	�]t5�&�O2�����;[�8����k��A�B!0,�a̓�?����?Y���?����O:�YE鎷8�6�H�̩:*ʄ{�OP�$�ȟp`吟D�ش�����w����|c���Tw����x�Nc�P�mz>qIF����'@a�� ��&��5��ubem�+v.��4�K�?	`J9�d�<ͧ�?Y���?!D�Z0c"�9`eU�m~^�r��L.�?a����DҦq�	����	��$�O=���u�� �2L25EŚX��Op�'E�6��֟�&��'V`Шr� �(�DK5���t�R�*Q�eÅ�C���4�pQ����P�O�9���.t(d�	T�N��I���O���O*��O1��pJ�6�ɓ8�*��,X�p�az�I�$m[�,�3�'���q�4�8R�Ov m��dyd�yd��Q��<*�!A��	P��MC���	�MK�O�02R���z���<�1��43H]��FLj����U�<a+Or���OD���ON�d�Oʧ\5bzF#C������X�&�*�i�t4�!�'���'��O�r���X5�Ƹkrs�ոs�˳!��ilڐ�?AJ<�|�G!U(�M��'Z���7�����жO�$��'��PySJ�<�4�|Z�H��ΟT��G�iX��P�ظaKݩ�ӟd�	ȟ(��ZyR�r�`� D��O����O��z�L˕�$��ێ_L:D*>��=��D�Ԧ�
��ēV�����LN�:%j�b��=at �'sJYe!	1�¸ U�����ן� ��'�
lgd�.U����4oVU��a0�'[B�'��'��>��,Y�Q��ҹ,�h�c�
x���ɚ�M�AE�!�?	��!����4�ċ�+�8_ڂ<��T6�½!�6OҀoZ �?q۴���޴��D�N������"��}K�m���*���'�*��Q%3���<���?Q���?!���?��E$T�``�IgObtsd�'���9
R��by2�'��O��@�wIp�
�(� �Б#ݦR�N�l����O�O1���x�I����TA��a#��aL037�u����<1s,҆<���d:�䓾��F2W$f@�D��Z��
�k�]0����O�D�O�4����֯��2r���e�Ƃ$2��y��=��Aq��⟤{�OV�oڳ�?1޴��t�g,E�`X\�î� �� A�����M�OT$����,1�i���I�/}C<����>���O����O��$�O���5�N�Ta�/�R�rC��+�P���՟��	"�M%�R�|��&��|�`R���)s�X)Ju;��À �O@�d�O��$ų���$�ԉ���Ĺ��P'edr�����\@PQ�'Q'�P�'���'�"�'�!��h:���կ\�@�Vi�W�'V�P�(zߴ�����?�����I6B0�`#�W-
<u����:Q��������	�����S��kB
G�❹��  ��a�আ�5�&ds�g�ϐY �_�擘n" �m�I**DV�zA.m�w�	T�Z�Y%�����՟���՟b>]�'� 6�S2���Q��JK(�f)��_V��7C�<���i��O (�'��6�Y
~��!=9���X8ک�I�y��H��a�'9�1�pK�?���X��h�)�,��Y��U�2�8	�a�Ė'�R�'��'~��'f�&Z��r���Z�L��A
�q���4�ڱ	���?����䧷?!b��y�a�~X��@��_�RK��"U�I�6=�6�Ӧ�O<�|������Mk�'D���ݐNQN���J[/G@DQ�'
�a봄�ٟ�rđ|�T�����wmR�G!d�k N��Fr60�'H�˟������iy�ay��P��*�OH���O؅3b&	�C�^,��(M�`9�����<�����d�O6-�c≎L[�lx����f'����#�5D��A�xYf��"!�H�|�VB�O�H���B3��Y��7``� $!J�v'8�A���?���?���h���;3�"�"��ρ�
�"��7��d���]�$���������Mk��w��X@*�� ��)��7x�@!�'d�6m@ĦQ��4xʔ��ڴ��$Ҷ\o�\��'Nj z!نF�L	[� �`�s'�&�d�<�'�?	���?����?���� V�|�#�Zi�UqT-�4���	C��J�����%?�	���`d�!gK�T���	i�:� �O�0oZ=�Ms�x�O/���O|\�b��8��:Scf��1�H�8Ȁ�O�� �G��?��#�D�<i�ɇ�t��y8`�_�2z�M��I� �?1���?���?�'���Ϧ��oP�lZ�*X7^_:���*O+ ��I�'o�柘��4��'�x�vC�&-�O�6m��{؞y�SEB�"�"�Q�J�p�3�j�j�E�ʰ+�"���T�J~���0!T�+%�0e���h���2pҋu���	��`��������|�: ۴M��ds���G�,��cC��?����?���izf|�͟��m���'��	:�̓,��1/�8p�o��Ot`l��M���=�1yٴ�y�'���9!�ҭo�
�ÓuO"Y��h�78&��ɤ0��'<��T������	=I�$��_�VF�3�b�>���韴�'W 7�'Z�F��?+�����Ɏ������A��1Uċ6��$b}R�k���IE�i>�S/&������΂9 P����9b��O y�VD�CcGy��O���	�1U�':�]�6�R;<F�5��ò t�R4�'7��'B���OG剁�M����9�U�\�K��9�r�&#�-���?a�iQ�O8i�'D@6m��d��/7'��&!؉>�l!�MCM�M��'[BБ�p��S2	���5"L��Ѓ�
�1*@{�j�IRL�My�'B�'/��'�2U>Q�g�a)��ퟱ2 �%��Mcլ�?��?�J~Γ���wA�i���A+���$f�)Pch	��"��Iy�i>���?�y�o����S�? ���1�?7��JU�A�Dj�>O���wϭ�?�4i=�$�<Q��?��K��$�*�6�Y�������?���?������������ǟ��I��!ӬU�|۰lB�MEJ����o�$��ɔ�M���in�T������%���k��E4�еp�|�ɖ�d�p`(]2���j�;m�d8�?��OI���`?N&�#sJ�?���?Y���?Q��I�OHaG͢�ļ���X�9� �O�<o��
r��<�f�4�bpiÂA-7�,�10�Ԉ�2؃R1O��nڻ�M�$�i5,x�iL���OR�s��=�â�,/�Y���X��2P���v$��O���|*���?����?	�9=�0S"j�8��A"-F8�B+O��o�T,���ڟ�I\�s��R#�o���Z+Q,[�Ր���Oj7�o���)�� �j���0���:���|`�ه˘)��hr㘟��*W�S���zy��-�xZ�ɟH��4��I+V�r�'	B�'��O$�	��M���Y��?�F�F��E"�Iz�<D�+@&�?�3�i'�O��'��7M��XmZ����T6xB4�S�H+����צ��'�`��I��?i��w)t��V��+b�8���%���{�'�r�'��'��'񟰨ð�5VfDu�5`T.K'��O �$�O8�lr����H�޴��Nx���T��y�R��܇���गx2Hh��8��&m86gj�
�Lx��`�f���Tؒk�)ӛ�nZ0\�ն�M;RA"���<���?Q���?��l�M�ҵq�T?hv��{�k��?9���d���IZ��hy��'+��^E����n"k���'��tA�	��M���'u���	�e���	˖t�, S6��4����H��(9ͫ<�'t�h����w��آ.	4�4C/SCDD���?���?9�S�'��DZ馁�6G��eoJ=Ц*�5a<b�2@�
�$.6$�',�77�	7���Ҧ͢�aS�Z�Z<�F�G�k`����Δ�M�v�iD�\H`�i��	�[ZX�6�O�L}<y�U.A$�10���&;itd͓����O��$�Oz�D�Ov�Ī|2c-
��D���ӄ:&tH2l�-��6Ͽ2�'B���'��7=��H�ʈ��Ą0%�*�$sW��Ħ��45#���OD�%�¿i%�d\�}0^�HA,@X=sQiU�Z�D	Y$��:��T�O���|��)9�e��F�}�pyچ���h���?!��?�(O>qm��>��ğ�I0D��Y G��+fVmS�I6�
(�?��V��H�43U�69�D�  $I('��
g���R\�y:��O8��҉L�jЊT˧��d�m�2O����ZrH���~�J���6S:!�7�H�4�����ܟPF�D�'���j� ��#�&��Bρ1K�xA�'>�6M��n^��:B�6�4���h�� ,"B���%�<�8M�p4ON�nZ �Ms�_X�(�޴��d�7�|A��'z��C�ֻoE����$5E����#)���<�'�?!��?Q��?�s)�l�9��m�h�Zg�!��@���b����8�����$?=�	� ڈ�$m�/cn����[8!��OhlmZ:�?�M<�|ʓ��'0�,����l������O}0J#�:��/G���6뾓O ˓�X�B�,ݨo/�]�P��+� Z(O����OP�4�zʓ�F���@R�@�p�91���c��4�y��yӨ��C�O��o��?9�4=��`h�d�@ވIJ����a�sb����M��O�iS0l̰��t9�	���@�˜9)�!���ۂ<���&<O����O���O���<�|�!�maS�[ .�F�Q�/I"?<�����?���:��fdÁ_8�	+�M�K>�r+����u��̥�%)��'vJ7�����E=�6�&?�r+7'�tH���n�,�!.^>d�<p!�O&�L>	)O(�$�O��$�OX�F��g���IJ�� *�k�OX���<B�i����'���'}�7_�`��$d���@��c �8)�n����M���'������>�����d����U�D�`�@�<C8�t��Ny�O���	�s�'��Mq���p,�b�5� و��'���' ����O6�ɢ�M�cA��dVL1������b�#0P<j��?1Ǻi��O,��'�d6M�",�)�dA�7R�)��.�7 �	Ҧ��P��Ȧ9�'��@�0N��?�sU�h�B��|����@�.戤Z����'?��'�2�'"��'���,�f�*�LS ]A@9"��=8=��4q�$m���?�����?���y7 �	j�X̊F�LK,�;TMZ�1c�7m�˦�!K<�|���V��M�'ݴ9�!�^D�(�S�Y�<�Xhz�'��)B,A�ɳ�|2\��S���!�N�O�i����i��|�ՃL۟�����	ayb�l�~�"��O���O~UӤ^�N�fH1��v\ �f7�	�����ߦM��4Lt�'1�%����9����M	����O(�5m�#��g�)W��?�g�OL����AH� &�߮Dp�e��O$���O����Ov�}��&�0��5�^�(�pN״f���1��Bg�֪D2m�I/�M3��w��9�O��c� <p�f�Z�<�2�':7�@Ħ���42\��4��DL��(u`�'B��4��0��A�7q� ��JKDO���|���?���?��7���2�2\"���ʁ?�b��+O�m�:���ܟx�	o�s��)�	B�t��BJ�b��}�W�%��D�צ"޴K����O}v��� �y�k	�i7�7��
�t�
���|��ɘ����e�'�)%���'��wd�*�j����5�,�Ȅ�'{��'�����V��4D�`��qx��q�7�X,�C��<*@���e��V�D�i}ҭv��m��Mo�Ա�����F.;�}���vt�)ܴ���@�xN��ĺ3����w
��z�d��yHasd�˿v "�B�'M2�'���'b�'_���*\=��D=���QF�5V 2�'gbv��E��:�������9&��Ȱ� w�h�h��X7B��<x����ē>���j�O�	(=��v���Ȱ� �@�EZ#�E�H����$[�a<��:��'&X�&��'��'=b�'�������:l�-i���i&��j��'�RW�hXݴ{pN� ��?������٦~.Ri�S��1(�8��Ѧ��	����榹�����S�.��>�rQ���<��rgB�B����B�En ��pU��S�3"�G���y04���|���B��D��������I���)�by�Bh�$�:�A��Zt����ȸ�DP��ʓi����d�l}"&w���"�$O{
��6I�M��"����ܴ4��ߴ�yB�'�"�ٳ	F�?�h�R���J�e�޽��U��@�r�|�T�'���'���'wr�'��ӣ|r��6*�.LF�0�'����ݴF�΁���?!���䧂?����y'�K#<2*ţ�]�^4�@��7L��6MJ䟼'���?Y�s}\�P�i��$	��x�$F�W@��Z�D�%����IV����8ҒO^��?)�*]�`�vH�R�ur�G@	iK�j���?���?A.O�o�s�8��I���k�|����4�Ƞ��I�$� �?�T�P��4j�xRl^^�ʜi��&=�J��i���y��'_ �уe�*�X��X�d�ӑN���?�R�-���)a�<�pyJ!�ɘ!n2�'���'Z��'bT9�׷C�"�'PAͺҘݑ��R28�6�RP����qӶ��7OZ���O��D�<�&�	�8�(x#��&!wPd���,Rc�x����?a�i�x6m�O�pT#~���Wc�|�4
���lS��!����cA,Rؙ�Hˀ����4��d�O����OB��I.ddLe��@]+�ttC�bK�5/O��o��}*Z|��ޟ��Ix�ޟ4�2f��%�����[��O�0����?����S�ϪPhu�Au7�����>��܃҉ʨVh��'�`L�î�䟜iÐ|�^�D��dʧkp�bJA̴1`*�ğ��Iݟ���֟�Svy��n�� ��O�]A�D�I�֜0��P�di�B�O�!n�X����#�MӢ�'U���Q_�lT{���E$
Y$Н"����iO��1@���Cd�O�^�&?����Lo��$�\���GиE$F��۟��̟��IΟ��	]�'(�%��C�{�D�7�^{aPX����?��n��鈒��$�'X7�;��"ɂqBD&W�P`ï�/��)&� ;ش��'s�*q�ܴ��d"B�⌙�n�'K!�pb��Ѯt�J��H��?�'��<����?����?Q���P"i�7+�3lPh�9��9�?���d릹�g����(������O�|�&J9 L��,��)[�T��O���'��6G�� '��'�x��FeW�E�5��
�'/���Q�
a���T$[���4����k���O�L�u�Ŗ54�P9R��(d�@D��O4���O��O1�`˓9כG<V��0������֎A� �>L�qQ���4��'��
���b������4�X���G(�Dn�p�C�h���zrXhB�g���L8,OP�p��οM���ôE����K�;O�ʓ�?Y���?y���?i���	��z�M�b,�M�W�*N�R�"ֵicN]�'�R�'���yt��J%ee����kؤXO���ɓ��XnZ�MC&�x���@�@��?O�B�,]�3�N���A�|��b63O�U�1�	�?��8�D�<ͧ�?qBm�K��;􋟄�ށ!����?A��?	���զy2kb����ܟ�J�h^�$8��S�g�$<?�prC�h��yK�I<�M���i��O�us�!H�(�ry"�G�<�"�>O��đ�c \@�kD�E��I�?�� �'���	�#���n<	�Œ)����G��O~�$�O��D�O�}��?����v�O_���A�o�%z�`ݩ��qÛ�O��7�b�'�
7�<�i��b��)��}qP���w �B�(k�Rٴ�V�}ӆ=�`�
��ߟ�j��P���Ģ��_��(xWO1���`=*��%������'f2�'���'	I$&���x����|b#Q��Rڴ"�������?I���䧋?�G�>��5�ДLp�(a
]�	��M�B�'������O��O���1s֏M��1��"V�>�tX@6W��	�X��г�'�\�'���'��U��ƮEAb��_�wD�A�'���'����DZ���ݴ�$a��}Cj�iC���N�4q�g��R�����Kћ���u}Mr�
]�	Ц9Zf@�&%���(�@J3�F!h�h�5A�hmZd~⠕�y��A�ӫxq�O�������Q�aȊ��y�OV��y��':��'���'��)"[�8b`,�Y�BࣴlZ�Z�*���O������}>=�I��M�H>!��/k�/ѺL�h���@,2҉'Y�7-���)�	6��6m1?�*B�A!�\�N��SR�QxNHr���Oj �O>Q*O����O|���O�Y�íϒ>�8"�F�X��TZ���O���<1�i������'���'~�w�Xx@�e�0���L�`�g��	4�M���'̉��� B�y�"�h�N�ңNӳv�n鸓�ěO(���Q�(7����|JC��O�(�L>�����K"U(�=҃����?Y���?����?�|R,OTn�6}�20�Q�?N��Ď�Zmlɡ�����Mc�r�>� �i�8	xPm�ML�\Z�ʕ h�[�
�O�6�#Z6-$?���&)V�iH���9<8��S$�9�Ï��<Y���?	��?���?�)�"œ�S>SdI ���8=X�y�U��GJ쟀��ɟ@&?��	��M�;G xs��
?�,͛�H��{���r!�i�&6�Na�)�S)}���l��<����W'��hmp\P%�3�a����.�����b�Sy�O��(�� /��e�W YdJ�AK�����'n�'��	�Ms1�ج����O�с���t��0Pę?e )spB?�	�����ڦ�j����:������ԸM��d����6*ޡ�'�����|�T�C����Gڟ�CP�'D�hR�oG1ވ�
�j�s��3p�'���'���'W�>���P�3]	s8��B ʙ["}#C�'��7m+#T�j0�f�4��Ap�*`�(��c��u��:O��n���M��lì�Rڴ��Dh��y���'����ތA�`�f�Ƚ�6!V=��<�'�?����?y���?qQǔ3��(yH�}'80���T���d񦭰��������ȟ8&?�	=6��O����U�q������¦��4�?)��3�h*­�6�Pሄ���z��Y�F�"���!���A���O���M>I*O�D�M�^\
��@&q^�{k�O���OF���O�I�<�нi���U�'��p���@�4��k�4���'��6�"�	��D�O�.B(����t1d�&Ѕ:��X�$�T�8��iC�	�c+�����O�q��n͋�ȹDnVYI��"F�T*\��OX���Ov���O���>���(ᢱ�O5�dpQC�(b"x�����I�MS����ۦ�%����N�l�ꅛ�
V�Jm���ʟ�'�\7m��ӓ']|�lI~"b��:2��5+M $P����� C�b��`B2�|Q����I͟�B��	�W��	�V���U�c������`y�i�������O�D�O�˧"p���3��&vt:�q�m\ O�\�'��PM�VNn����C\�'BdS�D�$dx�P�~ؠ	D��#��D�TW~�O9@��	�.��'�ҥ!a�&b�p�R/_�t*⬙��Q���H�	۟b>Y�'�Z7MS�w��Q9���D<�t �U2M�DC�I�<Ʌ�i��O�t�'��7��>$fÌ�v@4S� 	���lğ�r�aI����'�T�A$��?M����7/6p^v�Z�-Lv�T$G6O ��?Y��?	��?	�����K*@��k��L�x!����%`�l�Ddt%�I��A�s�8����+ւ��;�u%m�5-��!�*L�2,�v~�^�d�<�|����M�'�R�R&P�B|���5��iƢب�'`�#���d�v�|�U�����DX��fp���!�5b��ş��	ҟ�Ivyb�k�@�Z���<1��c���6o]� �@�i��߶k��r��<����M���d |�� j�
+0=�@H�ñ*��IVvx`k����cLc>�s��'U���$B������1R�rDBփ�� �6��I����	����q�O��H�8U(��: �I�#��uzp����Ac����a$�<�s�i�O��ӻ5��0Y �\�n6�X�M�D���O�6�O��jA$j���"�(�Q"���`�WL_4�.\�V-�l����CÖ����4��b����O�d�O��b�A
$P<�0Q �5@�t�Ѡ$�<%�i1Μj�S�p�	e�'�`���"ݱ,r-H�- �zà@�[�\������Ip~J~�q�&8�$U��"�C�RMO
ϐ���iQM~� �9���u�'!�I�.�6�҄�:~j��.������I�\�I柘�i>a�'��7͎/VN���
�U���xA��MމU)V,2�D�ͦ��?Q'S�<ٴ(����'� u�g�P�X�[%�Rk��������Ju��A��t�9��q�� r����ڣW� � 7OJ�$�O�D�O���O��?�Ɂ�SHO�%��̟����hU�
ܟ|�I��)�4m��\y��w���OT!�wD�:D��Q��l�;!�a�Ф�O˓5웶Fs��I��6�5?y�䜑B�P�R桑�ut��CL$+�d�8e��O(�PO>1-O���O�$�O
Hx�AϑP0:���N-�v�p���O����<9Էi�D��p�'F��'��"ƞ\	��5p���b@]%�|�?�I�MS'�iXr�'�Zm\� �i.�i����(T�<���畗d�N�vc7?ͧ>�m��ʰ >Ɂ�M��!� Cg㙄@��hXV���o�0QgI9j
湨%���sy�[��8+$��Ŕs�8�Au��*��E�h�H#>��L���'-���F������죲I���#�J��SW��A�k+�&�[�
Z7C��)'j�N�C��s��%���S�le�vnɄ���tW-w��Uh� 
V���oA6e^2����ab���~��'��!o߲ѱ@(4θ�cJʠF��+���  xֈX�D(��}��Ӕt�T�!��#�\�񄑷N���Iy2�'��'F"�'T�$@@�Ιj���b�ޢZ&b��QN+>�'r�'K�Z�����F�����M{�� `�$o~�����M�+O"�3���O ��4p���8p�:ѣBf,I��-�#FQ�wP<��?���?�*O�PR7��u�T�'�:�Q��44ƴ 0��d(NT�V�|�t��<���Ov�d8�^�� � af�
�G���@,QW�%y��i�B�'�ɩ_3��(��0���O~����d�\�ڂK��V�K�;k���$� �I�C,J����4�� ���Y��� X�F�6/ڝ�M+,OVܺ$B���A�I������?��Ok̛ &Ũ,��-d
P�i�����'�Oа�O��>��D�ebH����M�I��c��4���̦�������	�?��Oʓ8��HH���
�Щ��K$@��i� ���'��R�O��?A�	���er#��,Ҽ,Q�'�/}�d�4�?���?9��� �Ifyb�'2�dH%X��TM��ׄ(ሊn��V�Ԭ���_�\��'>=�I�����,�lXKg��:m�ڣ\8���޴�?A ���	��	Jy��'0�Iʟ��
� ��e�U�r�-#��Bf��!�K>)��?A����%Lh�#��Ǡ{>t�P�eH����&Up}�[�,��b�П(���x��mj���>:�����JD�����g�	՟�����'|����o>��2cZ5���x5��%t"QeCj�l��?	H>Q���?释S+�~JGM=����U?>�����݃����O����OʓR󊹪�W?)�	Mh�`�������	���54r�iݴ�?�N>9��?yb�Ë�?y@i�Q}�A�$V�0�$��`	H��"J��M#���?I*OƬ��k�k�S�L�s�qb̀�[��uY��)��(�Ќ#�$�<�Ε��?�N~r�O�b�#ѥ�	`L�	�	�u`�l�ߴ��[�<I��o�����OZ�I�z~2�AN�RB E�y�.�Ɇ�6�M#(O2,z0��O�a'>��O��d�ZS����Ob��)j�W�5%�F`ݲ8��7��O��D�O��I��i>њ�c���@&N�s]�ɨ5F���M���?a����S��'��3��u.ݭ~Ų�$�ŤI1N7��O����O�U�%)i�i>���v?��k��HT.�1'l%����O\��+��|�'��sӰY	1ǜ�.����$� ;Eގ0'�i1Ҁ�s���>���)�	�9�Z�	�@�-�L
�@�s�Z�J<a��^g��?*O �$%+Zu��V�$|(���'	�2���<!��?q���'����;E�f���]*b*4I&,+v��V� 3�'�rT��I�E-Z��� Kb���ޅ�̜�2.��k�ʡn�����I���?1)O4\�E�iC2} ��H����fIռW��8L<A������O�ak��|���)�P��	�\�b�']t���qļiW�O�Ī<�%Ȃe�	�)�T�S����$Qʌ��%S��7��O���?������i�O��d��k�ӗJ�ҥ"����<W�}I g� |Љ'x�P��a�*�Ӻ{�ț2;�z���U�_�dk����}�'�erD�x�r`�O<��O���iz\<� o\�IД�@ͮ�h�n�Ky��'D�A7�i-��i0,��S-��@�e���)ݴ\��qB��i���'u��O`�O�)AZ���Ƭ�֔	��G��n�o��,����L$���<��c沜H��A�~H
lhe�Z'$����P�i���'��KGW�O�	�O��	9�^4��a$/��!�%MڞDײ6m�O2�O�e��y��'�r�'�^���'J�jR�\OpAH�)n�T�D<oLZ��'�������'�Zc��Yփ�)M� yv�_�G'� �O����;O��$�O����O��d�<�'N�j���"ŏ5��ͪ��+����P���'A_���	� �ɳ���4�ރ\���ï��tD^�C��w�$��џX�	��l�	By�XW���W6.��f�_�rl���Z&T�T7ͧ<i�����O����OZX@8Ox\���O��-���Y�!��RЦ������	��X�'RD9zt$�~������H
h���KD	��k. ���ئ��I^y�'�b�'���'�I6k*]i�M'\ ��b2��fm����NП��IjyRo�5��'�?q���:�H�\�4@��1(�0��4�S��I�D�I�(��*n�0��TyRڟNX�"��,U������)Z����i]�QI����4�?����?q�',Z�i�Av�sk���G�0u���#Wjl���D�O��?OF���y���9y�}b���(�P� ��۟cI���,O��7-�O����OT�	�s}BT�,�S�F���A23'�CJЩ!�(�Mk�ȋ�<�H>�����'�V$It)���6�˕�J�@lJ�A��~ӂ��OP���!B� ��'��I�L��c�`��윔c�I�2�_s�h�m��'��T������O��$�O`���8{�V���47]������M����Z�V��'Z�S� �i���F�_��.()tFA�����2¬>�ᮑ�<�.O���OR��<!B�D�9��hf�H�S��b��K280Ȧ���O��OZ���OR���^�"�$�C���8I:��g��2@�<����?�����۱b� ϧq6HP�Fΐ=1�b�)2��cc|�&�@�Ip���D���+@
���J�Q�2Z)f��#Ę5#�O@�D�O*��<)G�ˡ'�O��x�N�>�$!i6D�%lԀ��6 }Ӑ�?�D�O����)B���R�P��cA�;t̞TPv�o�f���O*�-8�����'"��C��6��udY�m	�bV��f�O���O�P52O��O8��C�$�P`l�/xt`��@!M`6m�<�"eDw��~��� ��`R#�?PG���`E�b
��b�h���O��@�=O^�O��>� �UqU��50[^�����l>��i뚝�vkӸ��O��d���l%�����R�8e �n�DQ���C�.~Ӥ���4&������O��ĸK/t8cPgޣ~~d�启_�7��O��D�O��+��Cv��ߟt��C?�E/]�*��;�Ɩ ^��F�HƦ�'��S�%n���?��?A�"Q"k��ِ��� aѢ�ʆ�Ƹ]��&�'jP�C:���O��d%��Ʈ��R�Ѫ´�a��S'$�h}�1[�|��Gh�(�'X��'�T�th�#��eʞ�(BD�J�F�c��Z�}��B�}��'��'���'L�h*4�Ŗ.u8�can�A�dh���y2W���	�X��\y��On��S��
�'��g �B	�0�^��?	���䓾?��b������\����E<%F�%J�K79�Q��Z�0���� ��vy����kL|�CC�)7��	ޤj���Â�}��&�'��'�2�'nD�Z�'�V�\y�HM�|�#3�XS��mZ̟��I~yb��8��������\B �0e:��S���^e���/[}��'���'}�50�'��'��I��L��>lIŭG�o���Q����D˘�M�X?����?m��O��*aI�.%2� �hƙu��LB��i$��'�f�y��'��'%q�b�`�mB�i��)��+#�T��ıi�&u�6�p�����O"�D��>Y��9b,�Q�H�jߠ�3s�	�'�&B�>�OB�?!�	�z�37*����5%k�]���4�?���?���W�E�Od�D��4�"�R�_(�1����#)�9�|ӂ�OR��5O�S� ��ԟ�ԋe� �uN�.!���P�W�M��j~��$�O��OkL�d��E
3��^�`�6�F-�I$K�ޤ�Iuy��'�"�'��I"#���V;1K�����7K� k�
Y���'�|��'��:C�$�[&��(J"�"�)��'a��ݟ��	̟��'z"�(҇q>��fǗ/#�(�3`.Ȳ}a� �w�>)���hOL���G����/u)�H��)�Q�#��>h��0m�ڟ���Ɵ���ZyD�B���He�P�i�Nܳ��GG<*�1��W�G{r�'�h|�!�'���O�M$h�kpxb�Xej�i4�i�"�'��	�{�$�	L|Z�����4X�f�E�K�����Zv��>��;�����S�t�?&X�\��G.ļI�* �M���?Aׂѷ�?9��?���:*Ok��13��L��Qp�}�r+݈A��v�'�b.��OB�>�X��U��[�Ϝ�+J�Y�d&��sr8M���)� �cԹs	���>��H񳄬�Q@,:2��"'I�ȓ]���Kc��m����'���f>X�BuOɸ>
�i9FJ�u��(	� C$N��|���y��!9����z4�M�2U�L��t���B��n	�w?*M2�J�Ck`�!��F�%�΀� �)y������2�;Cm�kz�rH�F��S�O�i82�9�Cȿx�Z!b��@2l�����?���?S�����Oh�Ӿ5��hC�R�	B��ࠉ�(;�,�B-s��-����;gF��)��O�%BWĚ��Z�kqeS����z7 S�=D��8�j��22� sIW�Mj���"������{aJ�s���-Q�qx���V�h���O��=1�r��n�\XB��4;�cA@I1�y���#�ܴ��@��D����Ҙ'���Ğ5dh2$�'hb�F�6��Q	pB�~�p��wF�F+��'�, �g�'w�4�P�c-��n��<�e��F%�6�8VND��G\~��P"��o�x"�ɃE:$KSD�/s}ʼ�B�iȼ8�b$��5�&���ꙹt��<S�;������ė'�xA�� d Y(&bY�|� �yB�'���!#ٍ�zT�E��w���9�'k�6��$1p�k�Ĺp�*�#�R��$�<�ѯȷ1��Iʟ��O�,Mqf�'�b<�W�xRT 5�"Q����D�'�"D�j�F�o�n������O��g����h<|�`���_�\}��KG��I�T��a�
�<�2�@^�O��Qѡ�SL�i`���@} L������Od��'ڧ�?�GG��5K t�!i[%��]��`�`�<х�@�6<x���҄r<��7�x�H��dM�<z�����^�Mr4�g,W"X��mן��Iߟb6��?��t����d���<�݋
Z(�#�L02�S�b�}��s̚��I�#�|����%�3���s$�W��Y�ȵ+��/]�bt�X�F0�s��y���?�3�/Lk�0�!V�nE ��4��L��b���<��t�g�ɿ���q��!>l8�Z�Ɣ m��B�	�n��\�M1'}���ӣV0��e���"|�0�ŕYRڀ��%+��Pq��T� �%���?!���?��'��n�O��$m>Œ�c�	j����o@�uQ���zR�,��ŁtŐ���Nx�`�Ƥ�P�Y2�	�)a�� &H׃;OD	��<#�jsU��Ux���À���͉J�:��^�K:�d�O���0�	_��~��d9��1�D��!�C� a���ʙ�� �gX��C$F	�N?��<��Y��'z����ab�'4��˦�eJCB:s�>UY�Mzr0O.y0�'��1��+ �'�ɧ� j��f@j>�Ń��͚4T��RC�'RvI��2cͮ�`���$J�]�jI��Q��p<��ӟ�'�,�d�	
,�� I�}-�9 �h:D��yVj�� s�G��ƙt+>�$��4ix@�U)$1x��dLA�!��)�<����"�V�'E?yࠌ�Ol�hэ�9Vs�(����}璘�Ջ�OX��N+���)�|�'�:��V�@53ʄ�5(^�`��M��pf�<�S�'슥�V���i6�!a�+�L�O |��'1O�LP�q�ʗ�.�P� �T��ɩ�"O*2c�=5B�UIǁ�I�����'8"=�`ĝ8֍��q���΋>M����'�b�':��ũ�;{b�'��2Og�ǵ(�J��ѥ�?{�Q��n��Q�1O�����'q2�(F���uT�@��(��]�{R(I���<�aAD�p�fT8��i�P��H�#��'�P��S�g��-|��@U����T��d��b�C��GalU�V�߷z9���0�{!��
��"|B�h�:�L�q��P�K�-�a����iߴ�?���?��'��O6�Da>�c������� _Fƨ�U�Fv\�B�	&&�u�5��D"�yc�O�<_ �s��=�h�5�H�P	[wMO�q�xu��DڜP1���6�Opm �W�7ji�6iǭx�FI��"OJ���"�=�P@q��%�$����D�`�{;>#'�iR�'�,�3�[D:S#Ąxl�pd�'s󤐙3>b�'���щmv�|�pz �H����h�����p<�֥Ts��M�.�ZEFI*��b�3n�����sx@��(��O�a�H�e(W�o�2Q��MӽUL!��T5Q[���r�I�hc�FӾ��sO��lZ$R:�QI!� TaN�SA�O�b� h�eT��M����?1ΟN�ڳ�'��Q�G�Γ���Z�řp�B4QR�'�鑱c���T>�q,x�;OCB1"g/	�P�N��O�8�)��.n4��	�E�?��%��UI��>���[П<�<�B�+�K� ��	Kr�T� g�\�<	d���Kj��4��R%<<"�@n�����$ab}��F�7�~`@6��El��L�	ޟ�)cF�����	�|���<���?��DC��R���֭M%ڍ�����{A�y��~�lƿe��`ʄCu�E0�{�牡��<�w�	�^��a�7d�![ 㔱�'c�!{�S�g�	�L~ɰ��
w,���m�B�Ɂ4p`��G�_��x�)�32\��JA��"|J@�=�Te�3��A��c�Α�N�ctLJ��?a���?)�D�n�OB�$y>!3�)�wJ)��m�#c&p=�7�]��C�	�  ��%����<R���q�����/����H&!� �&�B������'s��D�O"�O��$�O.⟼	TI�	�,����K�H�h+D�X�s�I��݊�O��J������'Mr���d9R���n����I(���` ��Q���D`;H��	�<!A������|Z�!<*���G��$/$���L��_�6dSaW���zc悧@���M*x\�z�-��(��xv��9=R��j%�&=7j�ȧ�ܵ�(������Io�ɽb$�AOX�Z� �#A&��;�C�ɧ_�m���3?�����jφC�	�M3��Mb4#���
)`ʈ1��VC̓gx�y ��i�R�'!��!����|2\0Cw�N�f��FEy�����O�8S��Ovc��g~ �V�S��� @b�K���	�;J�3o���!�*r?��QH��G�$\i�j@i3P<¦�"}��Հ�?��y���CΚp*����4{,`  �F���y�Â)g�VbၦpȲ�k� M�lў���HO��U��6Z�@�V,�X�A��(Z�����|�	���]��럨�I������a�RlN0:`�Q+���DU�\x�\f�g:p̅�ɶ#�L3��S8��!׍�A
�㞌��)<O2qP3�X�a�tq� ��p��R�7�ɻ
x���|�,��g���+!*�H��Q'��y��P&�Rpz��ܖX�4��o#?�)§�5YǨ� ¼H��jߡ"����כv�t	���?��yҰ�8���O�ӊk���j\*nH�6ОuՖ�: �'����� �@�s��q���1 "�J�$�\�s��9p�k�M²��	ec�%Ȕ�$"�O���h�e��A�R��� S"OLp�d�=��\���5�ԭ3��di�3��(U�i�"�'
�i8s�+=�f��aH،l�6����'��V!�2�'L�i�0�h��0��H��B&brӦ�7bګj��AŢA�����'��C�[�"�F�$��^��fb@/p��X�d߀=H�i�(O��p<Ib`�ҟ�%�{�	T�.8|h6Iύu�N���4D�`�'ڲ|����o�,�<��v�3��޴���$.	J����Ŧp�<yd	���f�'�2�?	����Ol����@*u!�h�h�����O�����U���/�|�'��hk0��ra{&�_?I�$M�N�0�5�0�S��IZ氳W�̆B��M�G���|��Oā�"�'%1O��	���U"�
�j޲���w"O �iTX�Pzv|ڦg�G�Pq��'?<"=y��G�	���"9ʦ��Bf��FG.$��4�?����?�a�T�{?�e����?���?�;0].@�FU�l��	� -ʖ\�21!H>���`�������$��9q�9`a
#�� ����RI��'�1��2dVU#b�I�٪���'�z` �%t*�H���]�s�N(��g���n�ʟXs��蟬�I~�'��i�'̀؋SMӡ���n®�B�'����J�7( ����煢R��9�O�o��M������?)�Z˧4c�-҃I�*#d��s�'J��-�v/5�������?���?ᑱ��D�O��S-c����I!$�	�BF�`��P�2$�+6�Dk!JdD��C�'%rd���Y.@~�	鴤]0�5�K��LXD}���| �(��_8�|	�͊��L����� *�(Pr��x� �D�%Rܴ��'�c?�8��7:-��V]X�,H�.=D��:�d�3!z�|�'�ӐP���Ǆ<�	���D9�W�ө{��=�g��,vYT�)�$��U��C�I+n�ȝ� G�u>}�� O \	�C䉿2�l���!�\���R�}��C����di�o��h��c���C�ɹjA�@we�*���5'�k��C�	0?����]Nf�hP�Ο�r-^C�I�8!hx;�oļ%{����'\XF�B�	�}�d�v��*����/�vB�I����#%/O��p	۸&�@���.,-R���H�`�h�ν^�°�ȓs>���Jf\��d�R.yʸ��:����Q�|�px ��TC�����^!X�J)"�|@�� :t(�x�ȓ�xIk��`129��+9x`f9�ȓ%��@%W6d�J Hg�R3!P=��.���(��H�X@G֚q�I��J $ 9l�9�*�Ö���S�Q�ȓHS�(� [T&tC��݊lKxL��QSZ �R��<
+&��Tl�n�⬅ȓ�T	S3�P2/(z$�uc�獡�KQ>��i�kžf8h�@_�c�!�䞷s̚�:���"x�:�5�Y�`�!�ĕ�<�^�BeqB��T�N�l!�$O�h�$���F`��Tp�ʑx�!򄀁���p�^�uب�q3�Y.Q|!�X�Y�$��o�0w�0B�]�[f!�$�.o*�s��J��<(a�޾H!�dH��� 3i�55��Q Ԃ��Q8!��Ȉ,
E����
���� A	+6K!�$�lπ����	�U,�t�M�u!�䍂F΅��D�:A�* ��n������=��z��~��Z$�J<�%�L�؁i�L��y��[,1�N� OO�@�j,����?Q�=����Dѣo^L�h�5Ad�E�`��N	�{_��'���D)y��4y5��-{�D�Q�'�D!�&d5Bђ;�K�6v�x �B�H��F�tC[���Y�f��ZX���
�y
� �A؂!�1bq��
ҧJ�C�҄��)<�=)���O2)+$�,Z���I�`)<dj�"O0}K��A�����ʓ��|@��'Q� @)�HX�|J�O�1@/p3Ǉ�!��a��>�Or�|������'t�yа(�,'X�d��d(�sӝ<��Be�C�9� �ȓ��\��L�f�*�B�P��D��3���;�C�2�xx�l�lJՄȓ=�p�BwN�#2����� ��9���dX SJϐ���_m�����91��)"��L���rK�����aQ��JJP���AM�k�`q�ȓZ��əA�Q�N.N��,Z'�t�ȓ!b��&Ng��p��ސ�ȓ0�,��O3 *Հn���!�,�S��4qwصi��[0u��$�г� ��h�:X�c&ʣd���e휅�J6 E�QD��1�6؇ȓF�Ԓ��?�.)R�N�;�>I��}�Pq+a&�TP҇A��"s2���� kl�
�dU��I��p1�ȓwCZ���!Ƅs��`S��D=1�T��:�dqqf��Z<;�9h���i�Z���NJ�cq�	# ϛ� ��ȓx��in�A��,{���&�~�ȓB�(��KJ���RDB>4h�ȓl�ٓ�N��^�:ĠD�jthԄȓ57�(pq�@�^�^	�Dl8ԡ�ȓ)C�����?D�0��]�D P�����!B��dA�軃���ꘇ�X�����p=��a�h`��7��"�ϖ�/�=���	���ȓ�"�А�K�n�� ���(=��a#)[�h��!��-��F�j݅ȓ
�%��А?C\`@�R�G%U��,(@�3Lģb>6�N'(|A��'C0(ʃ�A\�8�3H�jC��c�'Z���Q�������"�&$"��
�'��슐)Ӧ[����K,kz�{�'!���B���	 �}�bj�G2Je �'�p�'HB�p�����_�T�У�'�X�h&���c����Ɣ3�'�ni���6|)��0 j��!�;	�'6���爴O�q8�GS
	vH+	�']y���[G����E�lP�s�'���&N���Dٕ��e$ԁ�'��`��/@��ͣ�ğ!Yz����'t�C��	l`��O	=T (\�'d�X$)H2 �2�� �V��4��-2H�A�$ (KH��ě�]�~ݘ�	_G��a�I)E�axr��.H�"@x�m�
EZ�AN�Y���n�ER$�� gͲ����&�hg% ��d��O��|���'H���� w�8�{`�1�l6�
w��j%��8㣏.-����3��$�t�X H4>i�d㗭m�r,s�LH?��%�|M�c8�3�'0�}ڐBݱ[.X�P�g:\C�� #8�i�1bL[*
����.�ƨ#��$+�$�%����>�@n�ȼ�Eo&����g��b�Ȱ��,~��ITDG<���T�-���S%��gQT���ZF�!�DA�M�����P2wor��f��M��ɣ`��ĸ��W%��	H��i�Q�@���5uÀ����4[�!��>>U��nI�U��(� �D�/��@�a�Rg}�E�D/�]���y��T5N��E��:���0�F%�x"�PO���A��b�tD��*Nv�Pw�),j�h6�!�O0�kЂu4j���g�	ݜ�R�'� ���k��:�xl�f��>� �� *H.4TN@9v$�"x���G"O>�c�JX���B��2hȒ��$`!�U+>2D�%ą�ȟ ��Ċ*Ni��J)�1�j)CA"O`	�kW�\��@ǂ5��݀C��T�f��'0�Yd��Ϙ'^z8q���� ԈtB0L��h<�VX<�RÈ�&�¢W�:ux'�.
p^�*���%$�q15�'��zbTg�6%KS�I6X�j=k�_��c4)X�nE����[���Q懂[�Рf��ES<A�48D�p ���)B,��Wj��?_�i@��4D����P��j�kIi��d@v�7D�pr�26�x�"�A P	¤X� 2D������C����E�ߣG�Ҩ8g�=D��"W
K�d���1�b�S�n1p�.!D��x%��sКA�F*c�9��@)D�����	;V0�b%"\��d0�+D�p�畽Ms��ɵ��8i�� �PH'{qN���'�h�ӆ�'(vY+�aԏk���Cn��nd��H>�n��jl�(&����|R��o�b9�4��!IEl�QBMZ�!�p�"OH��F־?&��T�#ڬT������nϴX��+)9����ׄ3��rD��n>�3\Լ����FEj5����;612C㉕i5#7&��C�����6c����iA6뢹zbC�)��j�Θ�mc�&#�i��y��ƣ�|�{�,ݭQ"�IK��N���<9,ܯU*�i�O��ٷ �"���J�D��X�<q`���y�H"�D�`���#�7F����3�ɿ�؀s	Ѕ=��dyPcG:�O�D9�cO�'f�e{To,r���؇M�?Th���F 'k�\5��Ɯ2z�N��E�Ό���d���87m�-���[�c��Hưh�yk��}�V�+7��f�ї����F��4��y �m8���V��9uȎ�1�OT!$��bf�u�@Hɐo�rK�j�"&: �*`�C�oD��!O�$)�-a��[�g?a@� )*zr���^��X�
fN�Jx���7_���'Sl�	 ��+H��PtE8f��7Ɇ� �z��҅�9%�d�`�%�*����䞙$�j|�w��!EI����`��a�'A���'`�sܓ$���P6���h7L%��28E�h�'O��x�a�	\�x��!�_���DT�O�Ɛ���d�J�o�0T��=�7ʐ3|b�|�0��L���$k�O8��w��i�G4+����@.�xr�P�'��Y��Vk�h}�� _�����P�a�D�`��'az�2�O����sӴT���]�t�  �D�;M�Q�"O�M2Al˗
@ҕX�ֲp+&���R� KSj��B��T�k�0hAY�����V
K�8�Aw�2��"��,G�*A�ϓ������N�L���s���c�<rN��"��!L� |�㉵:p��8�ùy�h�x��!2�8[��"D�@]�y�ıe&W������"D�Xku#�)G��Z��U)Y&��>D�D�#���L8��g�5�`�=D��`� ���������8-�2�"=���:)���>=�@�Gu��ӧC���H�);D�pp,��PqJ�( �*Ls�<��:�I�#��}��ɭU�r��'�1Yʴp[C$�:�C�I�&�L���-M:')���c8��)�ȅ}<�Rl38F |@�dFU�Hŭ�Vx�\ 1dGF̓Ǣ�KEg0���� !�/�e��;���v�D����&by���$����b@�SܧY�\sfF�3U�� �ȩCX��&E��R@�r�h�`����~�\��?QSO�	�0<�����0A0���	&�z���!�Sh<��g�>��c���DRE�_�H��1�'^����F� �4|'l�����ϓ�$\R�yr��_-T���n�?d!��4����y��Y�L=�!�˯W ��ãE�0��S(������FKCh��S�*;}fI�7f���y"�E�g%�1�UjKr+��)��'�D`p��'����B��/(�P{OH2h�T�K�'�©V��9�BQ��3^RY"W/��x«I ������Ť|�4�Цן�y
� 0�*������"tnN	���:�"O�к��YD���FoL Q�08Qb"O>�S��ˬ]�W��%j�L��"O<��B��	WH�凅�H�!��"OP�W�Vfy��y��
&��d��"O$����Ŧ|^Dhf�֎H0Z�q�"OP�a�֤�|9;��Ѻ'PL��"O�����A�9�j=�"�Oʥ"Ola8�b 3":�]{U 2o�̛�"O �խ,��{cc5ٲ�93"O��4���O���M�7�Р�"O*Lز@�q�X�J��ƅY� 1�"O��a����ii�e�FO��}	�"O���
�
j����ٸ9�<��0D�1���j&��W��1;�)��B0D�� �m��4ے *���+��h��1D���X	�Mq�$S�H��Ӄ�:D� R�d�
{^ыѤQ8i$H�C*O�� ��'2��qK�G���Ku"ODAX�D�a�t�A�EP�M�ƕ�"O�tB�H�D��U%D(H���	D"O�yS""��a��«9�fT� "O6�;�S:9
�e
U��V�
�pa"O���@uhw(��N 4�R%��q�<у �^����s��j�gBd�<ѓaU��6�����zg��Y�<�t/�b�B}C�B?X���ID�Z�<�QnۓF���EߒZ�d�i%�l�<ّ�V�~�Bd�BE��=.*tA��~�<!��î%��p�ïP�����'~�<a(5r�	��A�?@�|��KQO�<��2���4�	5a����J�<�Âʷ�椐�O�.�W�x�$B�Ɇ [4lb�M�Jn��U�A4xM�C�I�I��@�O�+�45��C�H��C�I�e&0`�AIt"�*���g��C�ɇc�p{�^�%b���֪o C�I�x�w��n��`pw�	�?;4C�	NCʸ+��E3>�� ��nƎea�C�IxD0��k�1`e��$,��($`C�" �����9A�`�bb�.&^C�I�!�`BmC��n�ig%��nC�	�V{��UD�X�>@�U-%�bC�Zx��r��G-/Bh�4"��	�JC���N)!�:����]�8~؇ȓt�~�2�/Ѡa��*���w�: �ȓ0�zD��CI�N� x��Șn���vm�,��˝b�"��DkM�y��$��.�f�{��V5 ;���U��Յȓ{�șd	ȺR|\4 �gA�,�i�ȓa��(b�5[e�K�kC�Y�ȓ$�d�T�B�,>h����H�]����VEl� G�Iz-8P���H�r��/3}���|)��'ʊ�[�D�ȓ)i*�Sa��L_����IĞh8�ȓO�&Ay��{&�����7���'����D�� sv<ag�\�}�f4�ȓd�(�@rL����Iqg�$f�@�ȓ*�5��,*�ȳ*&��ȓM�B���A�9Wۊ��!�Ժ@�|]�ȓSpH�eBU�Z�x�PQ�؊X���|��ɦ�L*aU��Pf�}xŇ�(W��YoU�H��ѳ�U(CT,X�ȓKV��p� _���ۃn���:$��S�? *8*�'׉�
9AR"�1�"h��"OUyb�
���*�@�wy>Q�w"O�A���V�(l�P)��@��qA"Oܨ*uW.T��5Iv�ؚ'�>��"O*�R��pl`e�����ҴXe"OX����`�
\�t��?���r�"O	Z�ˮ�qD&X�8�8���y�U����D�؊�4��g��y�����ɉvT�w�\�he�v���`v�ـ�L2@u�P��˧M@L��YdP�8L��r}�H��˺u���D��橌�"��a���"0_�!��_��Lca� C��f�2���ȓd�D�C!� �,�.$���8/���ȓ9��$&£Ң���J�>�n���~H����^� ̱%ME�#����,����(�&�*��
\�bJf���[�r}��͔9R�-��C�J�Э�ȓ |�y�$@�-�.5��ɍ�m52ŅȓBPl;#)"�p�j@�e�L��ȓ@d��p��Qsp�+�ŀ!��E�ȓu�UZ��:"�,���'Vz8��'�V��ek�8���c�,��5p�̄�mU ��u@	]Z.� �bą~d�l����肣r}��fYHu�ȓ�x��cR83]�8(S���E5
8��x�Es�i��F7v|��Ȑ7��U��.jH�����1I�ĸ禎�+i��ȓkٔ��5Q)dj�5���y���ȓ=�ya�@�cmDѳE�BX���ȓ�����G�1cB�c��+1�C�	 �����̩tK��� �HB� yt���_,]���H-gTC�I�O�(�C�/w��IT*ڠ.�B�	�;!dD@��Y6�Ԁ�§9�C䉎ip2�a@W'Z8����e��sZ�C�#`�k���<M��Ţ�
ʏK�B�	>Y�l�af��-�`���ŝ�!�B䉸,Ʀ��E`%M���K��N0݂B��!���!��ݵoL�i��&�7_��C�	9I|l]3��]f��h��VfzC�=;St)��'>���b�Ԅz�VC�%6D60"�E%K���XVL�#< B��4}6�`F#�O\@��� 0;۾B�ɂ��(���B 	j��Nњr��B�ɿhS)���˾:�4I궫
6;u�B�	O�u��c�� P��fK�u�C�I 2l9��d�4,06K�7tk�C�I�}s�AV����K���t�C�ɮB��$�(ug2�PBG5u RB䉤V��a�k�8nL*P�UH�1�B�I'!֡��:�@[�/����B䉾_��s�f��3���hy�C�ɀ�`��G�)*d\񥋂�[�C�%�ܹx��J;4:p�C�[63�hC�0yjUP�+�
Z~c��3D�����T(�P�iR�]<h��h��*O��+@�g�����a�r�h�"O�S��Ut�B���S��C"O^8�tg�Vp ��`B��z7�4�6"Op��â�V��q��26�e"ON(��W;�N����F�H �01�"O�Xpv�	�V��$�e�a7>ݡ�"O0TZ4h�'0�pq2�v9P�"O� n����V e`r�cA@«1����u"Or�aP��Cj��ҠW^.2@��"Ol�p��>k��<�f��n�H��"O�Agm�)Luz���&�>r�
ЩA"O�5"5F�b�]�E���Z�"O�8## 0p��� $
�d��<�"Oؔ�K�\C�h��$@�X��Jg"O =Y�l�F��u�@��L��h��"O 5�f�MNH%K�T�y�5p�'��CC��0�F���zYK�'�1�� Y���uJaX�e�E�)��<٠�O0)NtT˅˜�($�C�@�<�d-�r���:��C�e!��ꡌv�<�Q��=4�m�3b�C�x�jҡ�W�<��Ґ.W�L��D?���,]U�<�7#X>*0�1�3-�<����K�N�<�$� Z��=���8���km�J�<��^
�R�����,!���-�k�<�Qϴ/�0�F�C4��i�3�h�<1C��- �%�WM�I����BA�`�<�$g�9nsF����j4,���N�Z�Ǧ�oZe�Sܧo����g��>jW,q�Κ#0�Ņȓ)fXa�'�0,�$�ހX��������?�'3�����qy5Y#��TB��'�`���Gr� ȗe"~�T@s���$ �O�i���#���:��Y��8ٱ�'6��&���	<N�y��h��\^��?D���2�ԛsj�H�j�v�N���)�I�{'�#<%?=xd�H1Y�
B��u��p`��<D��a�n]��4��q=5�咢*8D��9A�γ]Zb��'�N�Ȧe3D�`Хb�0F�r�����DM� K�l2D���3n�
%���h�\%#
��I��1D������"d�ZF��z��YK��3D���qK�?"��q0a������/�Ic���'@n�ЅK7O��
��IS>��ȓc��z&hH,�R�B�k�+Q�)�ȓj��y L R���a�M�]��,��U��Xq@��,bC�Tڄ�ۍKN���ȓF��<BQ'>u��]�
2��ȓL^���)���j����.58�ȓ- ���ÉP1��<��j[\T��?�b$��X� ���B@�po��ȓ=���R�g�6����,/�4��Ojx�3�K��I$�ǻL���ZP"O����ۇ8{(p�\ "Ohc!@�C�Z�	��:  �A��"O�J1�� R�Z�C 6g���"O�l�dT�*Ѥi��!���x�"OJ�8�"�%Tǰ��$B�9v�hd�!"O���`���g�ty)�!ʨ�]�g��nx�|���זijxI��B:���A�.D��c��6��L��NL�ݬQs��/D�<���6����/��}㊱H�	.D�����߂Q&>9�[���+D���7워vC��JgL_�2��bW�(D�8v�%|��`��?WC\A�Ѕ(D��(t��X(�0��GV}��:D�LA����.��j�g�8&M�� `�7D����%�I{J��D��5 ��
0�"D�����ξu��A%
H� �2D��q��N8+@a�1�\%=,��-6D� ��%:s��Y�Х1�EA��'D�H@�n;b��� g�/x-�Q"�#'D�� Zt��c�+Sw!��B��fR.�R1"O� �c��)���JA^�l� �)@"O@��v�=mz��` [������"O�M�T5HV
V��ō_n�<q���)@,8���aB�J��\E�<A�����*��IлꙠuWH�<9��@.�Ab�H0l�h��!N�X�<�2�Z��\��W̜�rG��"4kAI�<)Wl�v������l>^��'O�E�<�#��'����&�A�ySf�}�<i���!w�v�ӄ�
�H�j�q�En�<�`��Nv�EK$/4�@D��(k�<��i�L��k"�3�pu�_d�<Y��M7���Ā��Ĉ�\�<�#��Z���)^�Q�f�� U�<ѡ�$* tl���DrZ�J��S�<����TZҩ�v�1B��q:�]{�<qw'�:u�1�S�/K��;�.�w�<a�E��'O�A�@��}���J`Gv�<��N�!
�B�+�"�1X0`a�E�[�<i`͈��f�� J*y����b+�V�<�E J�)�d=yt��.�rPCf��T�<�F�@W��TAToaP�� 'T�ܢ@f��j,\��$�=��h�� D���aC�F�ʤ��ş�i�J�� D��SE�l���xFJ�� ��l���$D�HsBj9�v
f��^�65�E$D�|�	S
0<�\hBb���.D�Pɂ��%K�Q��JXz�
	��L-D���զU$'�Dp�O�{/Ԭۧ�5D��S�LJ^��s$�Q��T�SN5D����K��0,~ث�J�e�����2D������_���j�h��:��,D�,��D�V`4�J��]&JP�U�6!0D� �A�W�< �X8^c��h.D�0�� ���DB��D��)D�p��t�܄(�$���:-�'D��:��*H�j��~_Z  ��:D���ׁҜ~����ń�TX��m9D����Ę�{�l��ˁ����7�8D����EJ��0���e��X֞�915D�dz�O�%��ivY� {��2D��ঀ��I��Ր5�ݝ0Hl�8*%D��9����dh��p�`��J����%�&D�|K%�ɤV���J�j��FjE��	:D��s�f���z�&�[c/؂�jC䉳J�����XI5B�PG����*C�I�xJ���k���>��Q�$[�C�	4Zb�0�r�Ӛ,��|�U�� +��B��&>Ո}���#,3���R��eQ�B�	>m����G+m���kP�T=�C�I$c�^` �j��m5�ћs����C�	�g���q��&f�4�c��CU�C䉆@qdT�E,�k/\���ڳ)�C䉨"m%ZW)߃N�ճ�D�`�PC�I<Z��4i Bޔ\���q!��!B��%�9P�S�<���HSĻ��C�I?V'�0��
��S>�<:��N#�C�	�DFxMH��a��bv�N5�pB��Kf,��%W�ʀ�V�N�g'FB�I�Z�.2@ϛ=Z��B2 �6�B�)[i�P�,R.oԤ�+��·��B�	�OX���鈐rڽ�B���x��C�I�-8�w�
�N�l�!���C�)� ����7��ZD#Q�m�X8��"O�1е�
�`T����k�]"O�I��a��-�t�x0A�4���3"O\�S��J>
�X�G��u[R"O��7���m��;DO$v�"OХ�� �/)u�t��?����t"O\�.J�;i�A�m�(&��L�"O�0 ��h�X�K�j�)yd��"O����1q����6L�y\����"OZ@�pbgz�!cLV��҉!�"O HV%��K���� (r�(k"O�����ZQ]9Q��UO.e�b"O(��#Ű9]x��[�=�!P"O����E`�Tb�FN�f�"O@A2wg:&
��u��p�����"Oح���O�$lY���Y��8(�"ODlA���6t���?!��K�"OvT��]2!/x��TA�5o���f"Od��&ڗH�	uɁ$a��܋�"On)c�a\l�!���:1��s�"Ojm��f�jǊH���f���2"O\��c�L�j�p	�����;�"O��T��@��b�ژn,D��2r���(�$�#��H"�VA8B-D��Ũ�:��͓� ��o]��&�+D���UL��b����ܚf�k�)/D�4�R���w��S'f4SI��s"�,D�p�F�HCdÕX�Jr�y�`,D�� c�k[`�#�/^������4D�S�j(l��x 4���*�Jd�/D�@ɥ�B�ЮɒW�e�	�$N:D��S��Љ^�y���N����)9D�db�i
,C���g�V�>��e�$A"D��@��u�J��Ԁ
�+N|e�B� D�0�����^�B+J�yz ���I=D������a��Ȁ��˂"��dm(D���'�A/|��a�$J
�?��u�+D�P�0��D���nJ=4:��2��6D��2��5��pۅ��9E��� �4D�tȐ��0/X�UK]��ԠhCo5D����	X+b͚��X�lzs�'D�!�En�US��ͻK���k%)D��2FN=a$L��$�,W���R��'D�tQG��P�,l�� ͙jDPT�&D��X��أP��Qq��V�Y�z�9B6D��r�!��w�@aYiӧBD\���7D��`qJFu\epŎP�K�\)��6D��A���Rt, m~0��>3�!�_�<�|�`���!��D��LC!�D���t�5���j����P*!�d�,����C�&�AkT��#t!��M3+=�9;'-�;�I�f����G4bL�����f�IS�3�yR�+Up�pm�x�N|s��ݔ�y��Q)6$� �6IY��䥇��yB+��1Xh�,�.$b��H�h���ybo��#!�KG�"y�u�#!D��y2D���V���ֺN�^u�Ư��yR�@4(�y q�ʃ0[$�b ��y�"�x�nD�D�^�vd�9��C��yb�Z]�6�r��E��$��B���y2�^�A��e��_�t|aj��y�I
E� ��*<�UX�^(�y�I'۪�J�&�7�lp�[��y
� �X�n�7�䉄��č��"OX��%d9P�BU�g�U�ͱS"On���O�n�B����z�<"O�����T�����ƛ����"O��i@�G�WЌ`���l}�5"O��ru�߽9���C��! �� 1�"Oja��N�e0��aD)��{�E��"O�}���K>�ig(-h����"O�M9�a��l�܅��ɔ:�d�"O�TKթ��DհU0�XL�"O�-��$�����+�/
�(�*$"O�E�6��"t���U�����"Ox\��m>9"�x2����1�!"O&�qլ];=�\�ʳN�(b�L5�'"Ol��������ZvO�����4"O6�jA�_'l�����N<El�墀"O��a��6R;^ ��섨1/�P�2"O|�C#�O�QQM�6'Lу0"O�aS�N1,_xh�����:$""Oq30�^3>���Eќ+��5"O�q�`��u�j(�Qc�(%�lY�"O�\CBo�k�pɄ�Sl�\��"O̹ф��QQ4B�X1�hB�"O�����'"v|PK�GN8�䐴"O6!+׏�\���
7��X�90 "O���a�ǁC���%�G�85�X��"O"s��
<x���ȥ/�~$��kw"O��{F'���ib4��3]��q��"Of�6(�X���e�g�0�d"On����6��$	��=ID"O ���(-v� DC�0nb�!V"O ������4�2��Q�[�"O���I�2��l��W�&��r"O�1aǖ6(���Ѣ6Һ�q"OҤ�c�΀n����uj^R6��C"OB��������C���Sk4ݫ�"O�X�ʚi���`�0dlbS"O�QY�
'e*|9���4����"O��Iv�ׂ~� ��rP���b�<��]�c��t�Dn���UH�<����&(Q��<-��P�%�D�<���"ᾴ��T�J��@ R}�<��A_8#tVmK��Ê>a�A��%|h<)�c�(`��P�T�$�Rؑ�D���y��̊]�R�p�#ŧ5���ܐ�y�nJ�==6`�-���4�Q4�y�C,B�=.Y��P��IgZi��'�D���N$G����*M�IhX�
	�'�p��HV<��B,F�.��q��'2U� �ٯC3����E�|��b�'mȽ#L��X]0d�e��=bYRH>)�yC\ɰ$��,HA�&&ڝӎ%�ȓC!�Y�G��M��zE��tL���ȓW�`����=ɸ���@�,�nA��(\~�"�c�J��}�!
(���* ��I���,Nm�@�Q�q*`(�ȓi���
�,��J[�li�����ȓW���d�#I�o�Z�ȓ� 
1&T?Zf*QR0� n���[
]#�B#O�����جE�"%���
����1,4�9��`Zޙ��N���!S#&�H1��m_�y𲀆ȓ{D�$FˆYs�n9t�&����zW�=�2Mͪp�%i�=sE�B�)� ʍ �1{s��P��ƄP&�L;�"O��ʱ�ӛ,�x���jX�Hr�tH�"Oؼ[�G_�VG���ָ&�@�"O����僝�x������RT"OXx��)�0ZT|{�E�����"O��
�%L�D]3T�׀,��tX��'0�'�"��>��&PZlza�֎���傀�z�Ih���O+�@���1}ڕP�I=\d �	�'f����O�7k��yf��D5�A	�'Zid�F���Q��%B8��)	�'��KbC;tt�3�@���D���' ��C���#u �x)��
�'X I �DB`����W��xCb�
�'�@cF��9(��`��lܪ�B�xJ>	������O��10UE�"s6��+T"�|�8��'��x��5X5kb�ɠC�U �'�rL��m��8��ҍďB�RY�'��|C6�#K.�a�MT4(��J
�'��`�!c�$(�I�TEP$1�.U�	�'��k���.*�4\c7�Y�/S���ʓ*xAw"�]�H� �,L�a��Gy2�'9�Oq�����Q k���LA��5*�"O�@�#�"wm���t�\*�jh	"O�+�� D�	JS$W�z��`6"O�q��}?�9Hр�S�9"O��(�i�\X����ܮ`J����"O����L"Lh%�ѡ� ��њ�"OT�S��5S�X�2��:[����A"Oxh���Fd,0���Ά>ftU)d"O�D�$�
$k}Z����[�)�jԒ"O���fV����R���4�����"OnHa���f���*D�T�[�V= R"O����`���d���S�X΄D��"O~m�B�X�
�喡Y�t�{�"Op��BB�M��3�$5F�r�S��'�����y7�m )}����L�\����5"O|�js�ڷ^ܔM��6I�X	X`"O�Ѕ������љ!��͢4"O�AC��ap���f�9�"u@�"O�a�ը�/=v��"�o��)�"O0�{0��1�T� R8J��� �'�1O��6�X�M9B|�#)��ة���'
���O\"����(��QS�*Id����^=�H�7o /VV	Ѵ�8��Ćȓ_���%��<�̘��&��\.2L��~/� �:F-�!��P5�ȓ��X1�Y6~bN�p���G(�8���
i��$i�4��2�Ԅ�ٟ��'�,�˗*���0�@%�ve���?���?�*OD�Ә'r����ߴ@I؅ZU	������'9�ճpb�pӮ��
R�fa����'R(���N,3_p@SͼV#pJ�'�ȁ�U�
����2�Cy���@�'��AK���&����Ȗ5&H�'
R�RF��m8{���9:���ߓ��{���+÷.0x��ٷF��tz�0�d6�Sܧa�6x���DN $륇qKh��ȓn����]*Ed~��R��U�U�ȓgrй{1nd�����q���y�:��sBNSZ^��S��Y���7�i�g�ޒ��ؐ�P2)�����D�9�u��_��0��Φ~v�F{B�O���dN*|`���VOǇ�0�
�'/F�K&Ռ
�j�&�۽���p
��� Q�B�œ>\���#JЫb0�8Zs"O���! �|:��f�U�)2���"O��ӭMe{��Ӣ�63�l��"O4x �	=G3H��G9�x8"O�K��\Dl�*�!שn|L�D�d,�S�	/eb
p�+9N��&/!h!�]��dh��65�D=��D&6-!�˟4]�qh�/F?����+'!򄈖ʼ�R!F�R%0��e�; �!��A�TD�U�9%lUMG�+!���2�*�!"� 1&�6���!�D@ y�z��B�C�8��ű���<kў(��Ӯ{.Ԛ!mO�j���D�E�a�����O��OĢ}��OP�h�2�܉WtX�I��Qu0��ȓd�v1�0E��%#�U�ޙ�R�*D���Al�?�蚇`1v[�	kA�*D�@� �S�Nl�to�3�T��A;D��aD�ė<Z�`6+�+b!  ;D��ad(� �B��N����Q��F>D�t�6 @�������F�C[�qpV!�O8ʓ��S�4��3M���k`a�8;`�QP��Ԧ	�!��?hq����23Fr��!�P��!���O�8܉��I�'- ��)��,z!�ĉ]9�90% -,T�hĘ?<!�.	 }��iB
�|8P�F�3!�_�~�R����T��h�E��B0Ofq�u��P�8@��:P�\�u�|�'U"��̇2*gHq�V�C���*O`�=E��\�$�a��άX)0M C�����'#az���Ɗ� �b d�D�С����y�I�
'x���L�J\�i1�Y��y��E�|ؐYY ǽS�z)��8�y��\,ft�R�ů;����Y���xR홼$��F�F=`�(�^�O���$@֦ ��LXX�P�T�Ͷ2x!�d���l����`Pt`0I�r�!���:�
`y�g�X�b����.�!���)[n��0`)���a��*P61�!�$̻T΢�6H��F�����B��!�$_�4<��BFL?ti�����#K���Ą
^����%��jʾ�He��b�C�I�]ġAanB4]ŲX(�nߦ+;�B�I0@Ö=q䯙Y$T�`t_�vB䉋\��Px%�Nt�Jl�d��f�.B�Tg��
�3]�B��غ"��B�s�\����@<6��R�|T��"O��X�H�n�{��Ԥ+S�5�P�'�ў"~JԠ�3]r�2vΏ���! UEΚ�yB�E+*9��s�K�	̬�*fښ�yB�U?)=R ��g@'T�`C℗�yZe����C��p�6G��B�	��� ˳.�-&��JF%��~�B�%KCX]´o��H`p��7��C�	�i����e�A�b������̃C��=!�'A"P�0B��$p�H���%�TD�Ӷ8L��sgݼ��i��F#AhB�	#>�$�Z�,ĲQ|a��ņIWB�I�X0 �&]�L�6���%��W��C䉧��TQ Ա6Q��R�	��C�<0*��)��@�_NX�E�[)�C��Dd �T�xhr� �pG~C�	�#�"P����j�(�Á��@�O����O���)ʢ(����hف/�Pr��ה\�!�D�l���S�˞�.f�k�h:|!�� 0�*ҪE�S_�xO�2�Ƞ�A"Op��Q���Y؄hS-O�Z�L	"O������ A�t��+W�}�	 1"Ob�R�� �@Pj��Tk�.a�Ԛv"O\zg���o���˲i�F]�u�@"O4���C�+���"�և���a"O`�zS)�PV��W+H##���`"OH�+�I	y�����JܺT"O޽��c8o�d�2I9?<l9�"O��ʠ�L3����I �(�kw"O�i�%G&Q���id��*�J�y"O��Q�b J�&!ҫG#�j���"Oh�!�K�a����J�E��4S"O��P1�@>(u����a[)���"O΀ӆ/L�n����!N�}�4���"OT�rtK�̐y1u@
=J	>:�"O��H��]%��B�O,N�8�`"O��[1&���8e/ˎ9���T"O�`��BN��X��ƖJ�iV"O�PSFY-A� �A�0C�6�;T"O@M`$�,F�X0�.л^rbEb"O���BOR���jvm&9���Q0"O.���,�<:�.Qb��p�l���"O�@"pgW;#p��
��L�{W"O�٢��޸V��	�FXg���R"O���$j�
H�p1�kT4�r��"OJQQ���>L��L��D�0��"Oh0YS@�,\ڦ��֡D�;�p9Q"O����E�	V���J��QZG"O.�XWe�!l�,�̅�(۔t��"OX���R5'�BN��$l�"Oz�����?[���rb��;�}"O\�hwB�9BNѹ��81�$��f"O�JD�Z%:�t��gE1�P�"O���ț+P�v���DK�(Z)"O(�	���]�<pY0��[F�q"O���v��:
��c��G�L��"O��!rBցseZ�Z0��V���"O��2���f*>%�Bf�?>�t��"O���� �:j@na�ń.J�j��"O^B�� b6��͟�h�,��7"O���+
���P��iB��3"O�����m�����>>iHE"O2	K&҂y��XB��.��sS"O��2����*�����ڟy�h]�%"O�[�D������,b�Zq�B"O6�#��LW�С�
�-�1+s"OȼA����"�uag�(,M��c�"Op��W`U������bM1.1�)��"O��p�Z�X�<!cB��N�J!	&"O�!�gJM�A�FDy3��$�Ej�"O���L'(�4�a�(:0�`V"O¡�!A�0]x�	Âw/ �F"Of��.^/�f�b�*&&!�(`�"O
U�&䉇<y�ywi�i(x	�"OؙT��L�@`����f�6�Ps"O�͢&�1N1��@ ��1o�1h�"OI�gJ@�UX�@jg˂3m��$"O��C��Ln�V�8�Ѣ:@�hA7"O�A2��B�B1�&)C�^a�4��U�O�*|;�D�K9��s�F3��,	
��yҥ
jȡR��2O��J��y���]U6�:�V,�ޔ����D!�O�ԏ��a��p�G��}��Z�"O� D�[V�H�4|P83��@?�j���"O��:�kW*H��Œ�aĎ�~8�"O�����΅W�<�X��&*���+�"O��!�`�={j�S���)u�~my!"Ox�a�o�)d�t����?9z�wS����	�L�I�֦_8j�:��	���Z���Od˓�0=A���JW I[V���^$*8�7�A�<��f�-l�� ��c$
^¹��ď}�<Y1f Bv��� Ýd��;2Wd�<���L�@;�g�-f�򬳱�b�<��t�n�AL��dU�I�b�^]h<�@-��h����s�)z=VLZ�F���?�/O���ėCR�D�q̓�}�D	 gH�)Q�'�a|��Y��BTY1ˎ�u�uD�:!�D؞=�Xb�.Ͻ0��E�'-!�Pa�6�)3�Pn�"Q!�Y1h��bsLȞx�4�*��!No!�DJ� 0u�b�C�:�G�.�!�DI�W4Yeo�p������ lY��w��A5���b`�Ԫ�^�a���J!�5D�xc!�*|�jŭ�Q�2YC��2D�����=$��h��J\�+�$=�d�"D���r�X+$�IG�v) Q��#+D� ���Ҡ$�¬ۑM��\`��`�<D��S��Jc�l!ʗM���[��9D�2Í�Pi:����Q.���@�a8���䓘��@�y��<А�'�()� �	D�!�d�&eD40ڷN�Zh�|���ŋ~�!�D����n��mY����X1P�!�D]&6�D�l3sP�L��MR��B�ɓ>�����l�P���i��$�B�.G="�C�q��Ac�~�vB�	D�B\&N���$}�&��>8�
��D{�Os��B��e�G1,&�`�@�?�!�Ej�H�v(uʈ�W�
d�!�
5u�y҃v���/��w!�ܟ^����U�5H�L�6���!��U�y����¨V�hy`�.R$;B�'�ў�>����I�u[Px�q�T66�d���&D��h���%�\�S6҂$���U,#���O4��!�'�?�sB�<"�탵 Q;D+��a3鐴�yB*W�,��}�6F�,;�h�H�J�	�y�_0E�B��O�.z��v��
�y�ET9yY��Su/S;/�k&�P��yb�0��
T!Q�+K�|S�Ɛ�y�jښ �p7Iȕ&�D��y�!
�9��)x�F3>�5�A����O�=�|Z��T�=�B�~��HZD�y�C?}
�*@L�+^�!
r��yBdO�T� U�a���O,C��A��y�A�3�tI�k��P �a���y�N�8j��[4O���kΥ�y�D�C5��F�W?�@M��@�9�䓜?����^69� �%�Ƿovyk3j��xb!��ϻ&��`3�d�c;~A6n�>cj!��J�%6��KΘt/��H�+А+k!��J�:�q2���/V
Pb�钊t-!�D�18O���%�|�'Zb�!�dXc�pت�OҶr�j�t��7�2O����eԤN���B#
&r�򜫷"O=:��L%������K�@�r��t"O"��K*Z����3Ii�Z�
�"O lj�S�U���n]>� k�"OllIwP.Kt�i�D� =��(6"O� ��r� d��bBmմv@&���O>4#1�Q��}hdd�	i�z���(D�L�G�A�x�^�c7�:X�>@Q�!D�lzcb�)m+n�y�l�2U��P�N ��ƈ����AȊ)S�bX��N�,7XڱP"O$KE"ږf���g-ϓs:��p"Oލ2CU%���h���TZ�E
�"O�T�F��g4hN��[B��u"O腹P*������'D�p���'!��_�Y��X��͂���(��/sm!�D_�ʖ!&`̅;���QҊ��kaxB׎�?Y�y")ܙ�@��H-_~�a[6�n��'�� �0�ћ
Q0�Q�.1�{
�'��I�T�F�(Sw#�.��A�
�'��)��N,�T}�FkU*+=��
�'׀��Тn��`��I�	NfJ9�)O�����!I4K�,δ6c�Di�	҈K�}���q1�S_��X��w�Lz5"�$�<)�.�eW0(K���?��������yw�K$]�&U���ZUH�����y��A�@N���J�4�b��y≖j2����N3����:�y��D x��P�դ���f��Ү���y��P�e6N_�|���!3�Y��y��W�'�5�$Oۓo��#"�.�y2Jؘ	����Հțc J�S􏁫�yb*�l��͚����
��ၓ�C3���hOtb�İ�M�jr�����"����v�$D�|
��S�L�N�:A@K�Z� �%D��sf�ұI$�(�T
K�FQ)vC䉟]A�E�rK3_�N���#�+P4�C�6z��M����;Q�V�Z��C9`��C��6:f�	� �4\��q���Y=�B�	�Rt\��c)��G~��
��u�0E{J?��p�w�� �E�;$V���"D�TB�o� 4�ʵ�`�F�w<�R� D��*��؄68P}C'��%jA�(X!�$�B��@c��ԲrC$,��V!�[5M9$,X�j��tG49�4�$>rO���e	�]~RT��cC1�|�h"O�Ը���!��!�P�m!e�˥&�On�=��:p�O�C�(��I�#\Ty@�'=�PnZ'b�h�w�J�,gN<#�'ꄌr���&rA��I�M9����'E�:CB��Z\R����ơ(�'�:�p4�Q�Ӑ%��(����@3�'o@(���jop�i4HT_��'��=XL'm�m	�B2u:Hȍ��'�a��`�����E`�'~���*�%ۑ�yBEf�@���Q�xY^qQu&���y�� �\!bSJ�"ot@ ਞ�y2	��(����a�/Q�aiw�Ɗ�y�HR	T%�Y2e��HyTmBg�W��y���Ai╠���uV� �f���yr�Ӡ+�l}I�dZ�;� ��v�Л�y�� 8|����,8�]!�fU��y�B�	� L�e��p���UK���y���:!yf�#�aT7Y0��� V'�y"�p��[U�V/',�I#���yk�S���fB�&4"D�܎�?	�'�|�z�+�:S�r!!a�,?g�h8�'��GI^�d<ɲ#/�=?yF�B�'�\��#�&L����)3x�h��'$�#��1D��t#Q�^�+�����'Ҡ���b�)E�1A76~�Qc��� ����Ɖ(���h-X��p�FV�d��}��GSe������]J,0�C)D��&@�$F)`�ӔjW:6�t�S#�,D���S/��~W��2PI�=v�E�v=D�4��B���f����e~�`j9D�H��]L)p��C+F)T@6D����/�L\[u��'T�#P�3D��G�QA`����-�b� ̲<����38�
�,ٗ-G�����(����H<2i8bN����a%�h�/RW�<�U��QeL	�S՘0H��amR�<I���P��I�C\��,C%!�V�<�r%_ X}�
U�Y�|!!f�ɍ�y�F�1����6
:.��;�#���y�+?�FXч��/�N��̐���>��O�A�5GD5$+�:roZ6�M�"OzYhOA$L��Q�N�*k�0�"O��ٕB�Da(��snM�{�^X�2"O��Yw��a�Jy�Po%u��=�"O��땯V"cF� ����+����"O��K'�^�$Ҽ�����.��u"O�H;��È\�l���:PT��"Oؙ9���x��k�%x���a"O��s�۾ej��Ґ J7`�B��#"O�� 6�<9��H	OB�Xy��"O���W��*zt�Y3w+W�P��j"OvIW�D�+%>���A����c"O�U�#�6F���bBC�*z�!�"O�d[�j��8*��L�'x��A�"O�9�c�M:odNE+�i,d�T�&"O4ؓ��>$<R����ʏ!P�10�"O�� �jPc�FnT D�'s�����YA���ƌ9DI��/4D��#��O�B���� _wS5�ǆ6D��Zu�^'�� �L�uG6D�p����{�l�JTA��X6(TH3D��{�aVi\����_Z�(āW�+D���"	��
B��6��WLPРqM/D�h�!΄ 1<�1m�3k@E�,D��8`
ܥP��4�'B[�)� �Q,D�\�S�R�>��e#�F,��:�%D������P��`7��8q贡u�1D�t ��C��ܹFg�6xiv�I#D�,3��t�&a�A,.hNE`�;D��H �ŞZ���D!^n`�2�L8D�0�g��5�@5K�b�w�j�Qu� D�hcs��~�H���ڊe�-E�4D�8���ÂN�ة��!	:��fm3D��j�N�s���bbÐa(�;'N1D�Y�НzTB��P:L��F�O
��Or�$�<�O�2���b�(ӌY�0`Z!9FQ��.D�t!& f���%�V-��a��'9D��I�&�6 gl�V&������#<D��95-�)���Vg��sA<8��;D�pc!!�)x "4bN� I6�iW�,D��Xc� *JG<AȆ	����RB 'D�؈㡟9kf��u�ų\�ބ8�c�O����O2�O�3�	�$n��ΊG�R���2=tPB�ɫ��#0���F����>v�VC�I�xl�) ԩV�	0q�RFJ�Z�@C�I�Y��Q�F��>p"�#fe̥\��C�	-i.�Lj4 N4;���`N=
jC�I"gʒ��G�ƚ�̠��j���C�ɩL�X���U[3�X��$H�˓�?�����S�π N�j!��!,2���$�>ZEF����.�S��B&�p ���ԸkD�D�����!�D�}� ��D�B(�&� l�!��).4Q'Ϗ}����\�C�!�ĉ4f���;Op��;��s�!�$�q���ʥd�]���Ss'Qw!�W(:��L��o���f\� l!�$�i쩑��ӫk�2|���r-�'����i��I >�&\�Po�a��%>)4!���0�fȂCb
�$5�X���ݩv!�$�vX,Ax�B�$-B�gK'U�!��H�XԈ�eo��A+�Y���B!�ZJ��9V�w5DX���:)�!�P�e���$H$��$Q";�!�����Ij���	���e$�%�!��8]��Mʅ"0f	 �(����>�!�D�?)�xba�[>-:f
�
(p�'�ў�>�TH�(6J*=x2�?(W0K�.D�����P%zn�P��]*��8��,D�d��;���ř�8|k�O7D�Q!.	�飧�m��Q1�0D��%eڬb(���En�u["K.��-�S�'d������F l�x��E�J�00�ȓp�m��お�n�"��4)?X��-�Ԡ�!MW�P��!�)�(A1�y��ڙA�×UO����5���ȓY��ЈC��2W� )�E�x2J�ȓHY����9S���H_�P<���)D��!k��^v�:��x%��f�<y���ӂ���� ԫR�%'U�y�HB�Ƀ|����Qv�:�q%����B�	�"N<�ϋ�aZ����H�B�	�mq����#n P �Q���*>C��		�Uc�%�L?�S0���1�C�ɜe&P:�MR9N�����h��Hq:C��+��t`��\m�j���(�;k�C�]�dHC��ߢa`*�9�ퟚN��C�	?P��x�⢊%DC 	[�
\4#��C�ɣ�N5R���=f�ř��<Vl^B�I�� |X�I&Tr�2��'m�DB�I�Wipxzd�ǎpQJ	��
���C�	�h;d������w��� ��	*0���=�Ş�����|P�1d�/�Lb�	�3]�!�d���u��-5[�D��	\�r�!��+s��9�0�E��<1�ć�;-!��2�TR�p<X��T�g(!�Z�$�
�Cc� �%�Y�U���"
�'���R��dxv��ԗ}*E
�'\�Q����Gn:�P��q�,X ��?���O�лU�L��Lܓ���6(ກht�"D��e�qjR(#Q�W�FvT�Pe^l�<��*�%�����]!@�j���\f�<Y6@�PV ec�'��{ ���x�<��þi6�s���<g��=xVo�<5��Zx�b�G�JXJi�.�k�<���,G ̘EØ5-�� 9��OyB�)"�O����c��kQ����!�
`SB-A�"O��IF _|	�A�p:P�*�"O�!r��r������+RG��W"O������v�fQ�aNQ�4��-z�"Ob��$��^m<q�wMܗ� d��"O���Q�Y�Mx�D1�K[�m�-x�"O��w#-M�t �D��������'aў�ST�'����O�(#�.8�U抶Pd���� �L��D�%^�>�ITH@;X��z��	ßdF������
92)ݏ8n��I��yb��'�0�'���c� � �	���y�GV�R���[�hQ���ܺ�y­]����"�J6P�B��G�ŵ�y�U���dA��W�@zX�����y�����!���J������y� �;7&̀a
�4?7V�� l_��O����O�b>��Q�	�<u(6 ̢[�RU�	2D��:�퍚0Hx����x�8!�s*/D���ڦ�"��H�P�X1�sJ"D��c�ɊZ�x5S��+9�VM;�!?D�4� ���H���0�|�Äi)<O"<A�&��mʃ�\K�d��+^u�<�%�(��Eg_) �嬘|�<)7�L`�`�E�=y�<LCf�Uy�<AE�^\� [�nX�
�&�J��y�<)�M�>�P��3d�*iz���o�<MJ&2r��pv�j��z"Qj�<!�N�o��j���EFD��M�N��k�'71O��Qr��Wt0��2�=�|%�W"Oָ�����y;C�dv���"O��Z��
�JE12ĭ=�� �"ObH(�%�"yV�A�@ �0ء"OV�hϚ O�2T�vK���Y[T"Of���Ĵ\q��+��� y�"O|Q�V5�������d��`�4"O�B�`�8��b��+�ȵa�"O���dk#���ʄ�Բ䆥��"O>��D���0���ꑳq4hs"O�T�#(Ww��L�QmJxZ�"O� U��R�uc�kرCe���"O"����*�P��
�_r��4"ODZ�DE
C�H8QT�[�N�L	��'}��%b�ʎ,C0��, ��b��2D�����*Ϛ�@�&l�$��)0D��SQB_�{���Aw
R�B�T���+D����W10�m�%MS��,��+D�$�6��]� eK�(��N�$�a�6D���e��N (�D�ɑf� ���A*D��0�F7��qG���6I�a&D�Ȩ�b� �:4���ghE���#D��I$l[%�:���đx�Ez��"D��@�Ss$��V)��Ϟ1b��!D�lGIN�V� �+�hA.R���a,D���ІQŊd�fG�"S�� �5D�����^!�\�W� �^-�8h�n5D�`Ö.�,J�2�J���G�n���>D��e%W�6��e�2V�@Dy��9D�,�RG�*f�<`���;t���`*D�� #&\�vE����|�>-*��#D��i�&��}��b�B��%D�4��*��,�6��eI
'z����$D��Y����d�(�(0k�)%�ּ&&D�`����i*���GcA61z��1�a$D�X��k��tQ��j�%��V^��Qi"D�x���ŚlW�=2�e��=���!J?D��)���&y"�9��"��]Q1�0D���6�R
>{*�P��0� rG�0D��i���Eڈ�7��)���A��.D�ْ�Tr.�rdB���dz4N-D��( ��:o�`���*�~)����*D�\�R ,5���aq���6����&D�ēBCʤ�9X��\5R삩��b#D�� �����!t�	QG�P�V�L���"Of  %J�cuX]C#��:���R"O�0uC]�!�DAh��#�
)��"O��aS`�c�!��.M#x��
f"Oh!4���u��u�t��7f�""O����A
g� ءf�:lQ�
W"Ol��5��
A�*l�`,�0@G�<�A"O` S�-ܩm�8\��a�E�"O`S��D~���E���	B��"O�|Rd �&=F�0�	кMS��A"O�M�Ε�b4&m��F��[<DlA�"O��cR�	�?#Z�`�fՄg�G"Ox%����#5��}D� E�6X�"O,�9���:�N ���?�tB�"O����n��'�Щ�3�U4�ذ�"OtE�P��(��\���
?�Zu��"O<�LJ�Gwbi�[�,�`XZ$"O`���ZL�R��R
�	J��	q�"O���%��	[.H�j��/ Ơ@"O
أ�@"6l
�货\���\b�"O�za�V��yHWǟ��$�""OL��u

7��Y�%�X8YyݐB"Oda�ƛ�T�(s�Y�,xj���"O�!��䏫f��M ��@r���"OA�d��
;lh�)�� �?U��q"O�6���~�V�Z�	
HB(H�"O h�
r�b}J��*M]ȩ��"Ov=��"<��hT��,fa4ȋ�"O$����
�^M*3g�>Q���w"O,t�G^�DP7��h���"O����	ˡ��dč=L����""Ob|��2u�� �@�(t�"Oވ"Q�N�#�`���N!n�X��"O\�P`[�
�d-Qg�T�W��X�"O���		Jb�8��ڏJNP�"O05 �/Â{9�@R ��+��P�6"O� *B��6a���{�hL�p"O���3mDO����"E��D����w"O�t�UBK�v�Z"p��G[	A!��6I��`�A,M���
�u�!�U+W��g,�`��`�e�<X�!���KTl��C-W�H�õj�,�!��94r!ӵ(ʽ�Tz��w�!�$[ ?��ġqNӬp���x���o!�@$(k�tz��h�j��@D͂}�!�֯+�k���(fbd E�

!�D�y�[�FO�#X�M�4d�&�!�d�.��!�%E I����b�0�!��?��%5�V�gH�Y�F⇸*!�$�����xi�5,)�Lɢ�I�N!�[�1{���� mP�ڤ	��!��?d~\-
V�:e����gI�u!�:��U�D�D-7��� 5-W!�Db�&�J׋��FU�'�#QE!�D� �<��Q�6������O2H�!�A�A��!��O^�ˬ��7�G�C~!�DCH���B&$����ѵg�_z!�dR� ���٦[�}1e�!"!�dJ-%P0ї胻 %��Rpd�q�!� �Fx���*R
ޜ(�M�<R�!�M��U���X3�����<�z���θ4J�A��
NV�;`E�]�XՅȓz�D�q�/�W�"H3jKq$� ��0@�E�ߢ!x~%8��C�ȶ���S�? haP��9M�����ω)F`��I"OPE�P�������N�:["�a"O$��b,���SS�_8C]�"O���FY
l�P�{�[&=�ʽ�p"O(�@*ԏ����J��l�ђ"O4$�`��D�����(oM��"O��A�[�K��ħ9���"O�f#��rՈ�矼=%^<�E"O8j���n"
!�˜;)���)D"O���dbT���W�=�b�`7"O�� �"&���)ж)��&�y�K��W���)V�ORkEQ�ڷ�y�R�zW�9y� G�D��fm���yrͿo�č��+��6ھ �Eo��y"L�`�Px�4�VE\x��$��y2l��%׾��T5
@&�T"�:�y� c��uSį�-��!�L��y2g@l2���Ͼ&A:4�^� �'T���t抖[�z-a��G�i���a�'���r��.y(��x�.]�v$Ԛ
�'B�Re�iG(9���7��	�'G���
�;Yb�#ݿb�l2
�'�ա KL@�dA�*�3GH(��
�'B��r����qpW�JU�~xp�'���Ca*�;zI�g��bO��'�l�Ą'v@9qw�ɋp<�=��'�F-0 )�	���֢ÀW��q�'B0�����M�� ��MS�Z����8{�t,s���WҰ���W�<��ǒPqZ���	O�j��mv�<q�م9����ι{C4��HDj�<�Ǉ�+mIZI��әmIڂHe�<�@�ʯ$F����chB�����b�<���ߖ� dp�BBEVёC^F�<�PٱA��1�5N�#YQ� J@�<���ÿ0��`�	]�R���)�x�<A�oֺr�fi�p�J
�b����G]�<�vk_LP�����:���2NKU�<�Dnĭk��t���?Q�FL �A�O�<��"N���a�I�V;\qx��a�<A�A�y�0�Q ޲G�`���eT[�<Y@ޯ���ԏ�0�P��T�<�!�X�NQgi���5�S.y�<S�Yp�RD���M<j��Q�7�AI�<�Sj2���a�	6<5����dp�<)�܂o�@�(3.'{,re��h�<�Uܰc��h�ǉG }2)J��<	� I���z&͐�}��-9��Wz�<YRBŜ^e����mN���� �'�r�<�a�~rqsu/X�k1bшp�ID�<�fWKj�����$g���H@\�<���H�R� ��!Pi� R�<YUb��8,u�S�t�fX��d�<	�FD):�1S��� U����]�<� �"z9��)D�C��{aeTe�<9'��0��Dl�-T��x*6j���ybM��L��Xe8��DB�߂�y�/Յu���fB��Y	v%���_�ybL��=�d0�B]�|�����y���--]��HK@&����U)�y����C;L�y%F4�H�@"�4�y"ޕo0U�� ΟzU�����!�y�']�L�Ќ�tl0gAN!�y"�X�J�����
�����J��y
� |� �Ef�"�P�b� 3��* "O6���˒�)�f5c�����"O8���� %P�Qy���czn$�"O��P���I<4Ls��
|��(t"Ol����׆>�@vi�^z�UPc"O�IxQ��O<�;Fh�p��M�"O�C�i2z!	�]"c�:�7"O8���A�&^X+eœ�)}b�"O&�0��*�H�	�V�FW"O@�<��]1��w�T8A7"O����O�:�q����.C}R���"O���Vި�E�I߸I`r8ۀ"O�� !	��1�RU��MB�\e��P"O�ԫg�%3�]Ag핐1��
"OF��A��:8*	&&9(^�J�"O�;��@K�[i�NR"O����Ѫ65H����I�o�LlC&"OL��ꗍLZE�7c��;�`}QW"O.T;$��x���2��U4�zy)��'�Oڶ�/v�^�z������0f0O$!��ɾi���(ҲAF@��PCS�����ZV�	2]Fea�cL
��mr�%�zB�	�6����N�u�X�2ѫߨ2X�C�	�pҦ��ƠI�;�L��j Yz�B�	����%	�D�8�@�dN�B��}x�сn1`�Fl�sĄhxLB�	�_N�ВM�U�"<��� ߀˓�0?�3c�?N,��@�Q,: (���W�<q�* U�"1�H�	r�@�@FW�<����,]�6E[��=((�vM�T?a�����s6�4IO�; 4�0a��!�$�2u�rp��MZ#��A�+L�"=��9O��*%�`�螒p���AW"Oތ�6��<>5�D7q�"OT`�U��(9�J�f%6^��2��IB����^$WL�t�r"��P��ꃅ�!��ͯd5t��"�74g�����
o�!�dɆZ�U�VeM uYir���> !򄀵#i�!�5��.9t�@fm��!��(�d-
�kп)'���&m�!�dI�3��e[ԃ��)
��q�E^�y���Uf�����VM�i����1 �jpX�a���y����i$��!�H쀐P���'�OH-KhL���{�@�31��M�"O�(��8l��D�H������"O2e E�����86�_>L�nL	�2O��ԅ�I�Xt4�#!
	���N9pp�B�I;l�t-J�(�>�N	�Ŵ�XB�ɣ	�~T3"JxabT$2,V�1"�#D�Lk6K���5����8.�h�l D�x�7�ݕ16�kg�U!L�,r�,:�u؞h[��@�MrU�%�U$j��m��&,D���R�e_�-�#'���Y�0�<D�,3�Bŷ6��TIpn׼R���R��.D�,�� T�%_(u�c$��䊡17�-��`���<�Z�{�%ӄ� 4C�H�^��d�ȓ8n�q���BUJ �AD�h��]EyR�'qμ[7�V��0 �k��yPzڴ�hO�	,�Q�T��a�?l�De�
�[���/4f��LҎ?X4գ���m(FX�'���G���'>ơ�gm��m���ꝈG��F��S�W���t���ik'��5�V�hF{J?�k���	�,��iƝ|�`U�!��<Y���S���J�*[�6���PqE��;��B�)� V9�B��(. $I��V�@�
�"Ob����Ȝ{$T�)�
���"O����Ŭ`u���W$~�bSB"O�!���ɺfK4��C�K�n����'�qO,�e]�0&��#�	��&�&��s�؟�E�ī�'��iC���[Ѭ��t��*�y�.L��4�p�ץ$R��j4�O�y2���;����-�+�:#�hY'���ˮ̰>�"��b��ݑwB��Ju8<�r`jx���'h�{�Ӱb2��Kd�^�x��	�'�H�#���XD���%��p�9��'����M/%K:5�B��<c�~1��hO6-C�c�/|l�W�摩"O<�hOp�R5����J��[�"O. #�.H$���%$D	&"O.�i�*/�H�o
��"�IlX���O����W�0����"ٗt�#�O���T䖽!��Z�#R�0d���} �x��	�^��-"�Ԫ7��p#�[�>!����?�@R(�����Ĳ�C���06Z$�Oz�=�J��?-�
�Q���6nZN��n�F�<A�Ό�m�\1�Պ\5nf�Z�d�}�<�q����3����7��z�<�CZK�d�ңA��%+��EN�<9b!5n�"�
�CَV�mh$b�b�<�আ�X��!ԭ�]���a5�WG�<�@'L��rU���:��\��_�<qK�oY������i��mk ��}�<)��k���)�b܊Uj1� ��B�<�1M��BQ�B��	1č��FZ��p=qD�=׺D�3
Ős��ȢQ�0eV!�F7���mB�G�u:���
�!��1c� 5:5�S,!;�E�G/�,ax��	�h2��ץҵY��Z2���P�:b��F{J|�ν?�ܤSWnهl�Pa�E�F�<1cJ�-��s6�D�}�����~�<��(���JH�gz��Ô��Yc��K8�8�R@Y��(	z�ŏ?GԐ ʢ�9D�$����
�ȆD��G�x��BI6D�LBWJſY,�%��9+ )S��>D�8�<}��U��"�+D̀d�>D�@�1K�X���Aa����8D�Ȉ!���k��:�ȸ�7�5�$0�O�T�􎂉5����#�Q�5���� "O�E�e��7?p� 5e�5��"O1(w�H�U�\�J5,M7}�<9�"O ��)V�m[@,�^�r�ʒ"Oh(k�%�S/B�)�K4U���f��x1��)�'B$0t`��ע!��"-٨t���g<�/�6� ���'�bu�V"�V̓�y��$\��ēo1PyЕ��9alB0 Q�rj|i����?!�)��s0Ԉ0"�Y%6�P%��Q�'�ў�'t�����Qx�	zE��pS�a����t�&Ɖ+�n�Y��HB5���ȓ���D�ѣ_�⸃��Y�<��	|�#�Ű'��bR�ĈT��OET���OZ|8���/)�h�#�3��>q�����1Z��9:��M6^u��x�
"�y�F; ,�0 ��x3���y��P)w�Fom��x�`')Y!�yb�@�xp�dƂm�4}�V�C,���T���O��H#��%ոx�v��94�J��a,5�S��?a�$��%-n 	 ��O)�Z�,�S�<��iM�s��qY� �D�^���K�<� �x�G�M�.��sbJ�.��A�"O*� w �{YNu��I�&>`�q"O�\���ţhh.��EH��M"r�"OV$[J�<�^ q��c0<�YD"OPs���"��`X��5+��+b"O�P*�-T3'@��Y�C��h(�a�4"O��&I�B��ur��
�}�=��"O�hB��_�X�*�A@AX/Wq��i��'��ė�b�l�C��9�#� *���L}R��ӱ[5�R̚ '�V�
t�Ͷn_�"?!����u�����G^3h�,��A�>0!�º`\��1�R�½�rL�:8��A��(�ԁ��S�np�%+�H\�w�"1X�"O�Bv��P����D�+O��0ѱ�d"|O��j��x!���1'��JA��O�9c"�Ï]�����CC`�XW�F�<Y��O�Q5t}���0�<KTË~�<Q��#~�����	]�~5}�bT�<!g��##��1���G>5cXU����t�<Ya␺Ohr�V��[�&4�'��r�<��X�F&e�KB����Jp��p�<�BA	�V^��_2g�D�ŊZk�<�D�Z�o�n
����vo����Vd�<I�M��~��;��X	]֩ca�^k�<1FAFnƢ �`�Y�@�Ա�aHd�<��&E�Ĥa�I�`��؊ �`�<i<=&0�ʓ!Sc��Xq�MR�<q�8��	��_J��ɸ���D�<����K[��P$��� ��K@�<��͙�{D��eP�l�n��c�v�<�#��7h���1S��ZQ�8���t�<9хљ�@��Ь9A������(T�t��� 9&�8�	iW���v�8D���� �q.\�#��А[eBm{f�:D���p@�=t�A�pL:/�\e*E�4D��Kӭ��&|H�*���W�:y��$D�HP�ҧf=�	��c�y0"ё��?D���ɝ#�P["Y�]Y���J>D�sc�+H���Wf\)N�ؘ���;D��
7I��1�h�����C�4D�Xc3BÌ5�����J�aϬ���3D�̫��D2;�kU���\y�)0D�t���@;�tA�W�%A<7��V�<A�%�+�+��
����h��S�<�lF�4��E�d��#`7\l��Dz�<)��θV�\BVH9
�ԠPA�q�<�p��.E@=iD�51�Rб&�o�<!4섉� 婀"��R��ek�<�&�W.��=���� *(�&�RP�<Q��� H�D���H%H|�k���K�<����$Xv��:��>Dd��A	L�<�Q�!d�,��&->�̡��$�|�<�eˀ�RG`���ŕ�f�<Xr&�r�<Yժ^�e��l"���6\����j�<��A��F��ȣ���-!�4 �w��M���
�Wj�C'�$	�ո�I�#pmC2gԀ��8ǀ>D��AЉ�#�((WMS0��ҳ�=D���a�.��`,Q/_�ФP�9D��Q$�P#�X
S�B;~��(ӧ9D�|�צJ�	 Xp1��@�BЮ��Q))D�h���Ʊ`m2 �c#��y�nX8D��ufDyنp�J�b�R`)f�4D�� �(�4\���EDX�MFQ��!'D�P�����[l}���L�0m��d&D�� ^��LM$"�ƭS�EԦ���"Op%�w.U
@�H�X4Jj�$R"O|��ͺ"T`$���
�X�>���"O2�qu�Y�%P�8y3�/Q��l)5"O���I=�2����5w���b"O�)�cM�=^8D1���0s �ۤ"OnM� �ș.��鉡#S>z{�z�"O��`V؉ע�3�l��Q�L|�"O�5���>o��iY!�^��Ւ�"OДl_�jƊ�0郑��Ȑ"O�,§,�s���[��ܯ@��T�E"O��B�� ��ٸ���%RV^�W"O�4*0늎wa���+P~0]��"O  XR�	��:12kʃ6�8�"O<��an5�<�Ҵ�K�`L јt"O�����θV��hi���,2��=�s"Ot�i�N�Ze�C��/�
���"Ot�b�`�<|.�p��J���e+�"Oz�B�$ �naq7I�=/��t��"O�$j�!����g��Dn�Y�"OI�ӆ׵A��B� T
~N�]��"ON��HN=	�����X?�D��"O���qh�H�ܽig+K<`�P8� "O5!uX�Uw�RWcRi�,�c�"Oj���LJ4	I�%p7B�2sǶU`�"OZ��v֗gf��J@"֯+���f"O��«S�e>�{w��.�"<Yr"O�ĐS��~H��*�R�<��"OT�2��0o D�K:ln��7"O�X��"CڕIC�W$W<�T"O��y`��%:�p`PJ� �:�"O�ĺ .O�^Jt@S6dK���Q"O�T�ү^�Х��r�����
��yE1N,J�{�� wWt}��(�yr.��1���历>?�>�yЇ�	�ybb�w͂ec�AC%1���2�)��yR��1~�̜�ᓽB��s���y��H�$��g�<9��	�I�y2�I:0k�(ZJx���y����N���0!w���bFʳ�y���=JB����v����%�	�yҊH�}�K�:1�vms' Hv ن�}=\lx'В8��y��ɖV�"%�ȓ-x]s�BR�@�-o�g/�Ʉ�S?�=�eBւo�BPO�q,-�ȓ1�p+��V7Z4|�ڃ�� v�:����V�GQ�D�شj��9WΌ�ȓGKj�PGՐ,�$��AV�o�����O�̓WLY�i�2'���@X��ȓ%X���ԇX���a�ggA�k�`��ȓ@'t�Ȫd@"��%I)6u��/�A��)K6I���Ӊ�m��B/��kU�͠?��( �"L5���/�D��2Kc�'�K�:-Ɇ�<��58�ۀJ��� ��M~o͆ȓK���J�Y�}	&�x�L�����R��(���`��q��S `��M��@>8���ղ�X!��#O��܆ȓU����
F4d`:�U$�%�XA�ȓx��ʑ�ǣ�����据:����P�p��CY����� j��|��>��`j���;1��� ��Ʉ.��ȓ
aT����șh�={`S�C�8��mJ�=iC��p-��C�(%U����	=]In� 
�1��� t%���ĥ-�� aRz��!
7"O�!#�aK��8���P������б�����Y3p$�}��Ş�=�����ײa}�e�DI�q�<I�,�?+S��P�.��a,���K�2w̮��B�Kd��dO�]���?�'�8����ȜU�;D┾X=Ɛz�'��H���F�_ h�fR �(�I�J%�z\��A�(f.��Kʍ���UCd�lR�_*���@n�\2���Y  }���\�fy�� �R1�a��DΎB�B��xq��	Ҫ%ItH�F*�f�Op\����~!�G� y�$�����Ԣr���HV'T�6X4�чfu�<�C'�6����cG�h�y���=x&]S��I�8q� 0��u�����Ox5��BcOr��5���>]�EORl��؜rg��h���O�bTB4+ħ_���y���s���F$Ű<�� �9aP<�@�	���4JW�Kx�8�n���(r'�	�9�%yQ&X6]��*B�e^�5@��!��݊Z�OY�������
o|M�<�����jtY��b񀩒 �IU�M��5�LR���)C���^!!�I/uZD��@J�c�`G��`���r�5:�T�A��ƟT��<yҨ҇p�%Vm�m��n�}�<q���0T鲆$�g
�;���Gy�K��|=�ehPn�NX��1E#?�f�X��X&���`;�O��ǀ�eZ$*�fݫ,�����Y������e�"�Px�n �0a����`� �ES�H����I^u�` �_�'?����D�3> �z��Q�r5���	e+r\�՞|�o٦3�*axǁ�y�؀
�K���~BIC�9���=E�*�!mHZ�S�)~��3��C:�ēR�<��*�<Q����O� ��0�V݈�:d��KG(l�O��%hX)=�����*N4���"�
M��Y�����`(d�pjd*����O��"�E�W�b%~dVcGB��IQ�A �x2ş�V�F���$�����yp�1u��<q`o0_zX��P�(A��� ���?A��"I&&(���%A��d�!,OT�fo��M�P�&�X2��]��@��j�$���p���|�)����:��dZ��?}��i�NS���a�. |���ҡP�r���O�����P,r���t;2����:��+e��蠂KU�b�谨�m�:�]�z�2��F�@z�d��IzҚP C�ɪ�LTx�"����	�2���B!kDV)���)�S�^��#�->lJ��2��W+9�$�Ł{� ��A_hH<���+QML���¾X	�̒t+ ��?�DD<&�� O�K��d���TDT��PP��*�0�p�;�,#"^���˕��Ś�'�X��!���-`�{�A�"'�������RiB�rT�5T "tn�uK@j�iy����c����܌s,咕뜽N��+�)��'�p�%ʕ;�L���W�y�0$>�!�`�"�k�K�4=�����p0��Y�JD���)<O�}Ye��x�8�%ǁWU���0���V��Ep�6Ub H�O�qq�
��B甆>���"��K�7=ʹɲ+9N�Z��*-�y��S!����ɔIɐ�SBʒe U�ى�X��T�X< �8q��F@W-���I�x����rL��k����e
�q�r,�҅DJ؞H�s.��!Z�� !E����9��	�0ɖEؖd�ȔaXQO�"z┈3�����ɼD��5)����]��f�H�س=����'�~�pb�q4/�(j�
�C�"ΰwa��O?C�Q���jr틬wP���.�>���iZl��
�6@��J�(�HH;��ҽ_l��AS��D���E�q �����]�'{�ܜ��&h��`���� $�"�᲍�V�6��"OfP�ϟ)n�N��G	�<x�E)��E����̅�|�h��GY�A��n1������(΍9��#@"��~1��	"qB�W��+�=�'� ��	a��?h��P��Զrr�!0/�_��9!B�N�°aq�o�L�Q�'�<�1�?!�Ƒ�wA^��p�R�5h\s��;��E�rm,��v�֯C���ʅ��	�a}���7���Iw�帡H��-/e�ӣ#��ͩ1���t�r�ч?9lX9r*9�g?9RÃ�;p�0 �������m�'�`5�A�]�O�@�D�V�rlP�f���pB�'Ar0���(�mX��ώ&џ��g�<J~4�Ӆ�3 Nazc�p�$�۷�N����ħfB2��f�y�&�#G�d=�r��ECRQD��:q"d�	�h�Q"ц���d��#�61vh�'/<x��C�<��Ӵ� �H���FM>T'?I ��4O~N�z�2l�����=�On��g�:�?Q��3i$6L3a�9I�U��[ݟ8�f�%(�ご>E���²C.�dZq�Ig��`�0SўD���K�π i�!^�7� p�ҫK�z5t��>�V�h��$�~$��F/Đ5
*UQ5��'!���"a�� ���2��YUKϐ}!�$6O�r��&��"�@\{�AR&y!���Q�J}�e"��4�t�Ñ��8�!���IT��Cn ����D7h��'�������Λ/@�Iy�ǅeU�5P�E�i�!�d�(�R�8Y9Acj�,� �+2 ���L<��_�3 j��AnE�H*�$�4@RH<�g���w��c��V|��O�dR΄)W�1�OHd�����laT`���j�z��'�)�rH�s�I,G��\����a��X@�BB䉸(�j�R�lh.
�H�Y�N/4OZ�!n�2帧�OP�ESf�	|wjA�(��$�b�����3f"}2��^�%�v�RNG"U�@��X(¸'z��%�4�3��Õ<O��tψ�3H���B����]�B��+�{���I�3��L��e�(�LdRe/��(8�k+�����-$`Ê�x��� ?At�����P�{P^��W*�-9Ԅ�p�ÝL�a~��$u�,̃�蔚��@{�/�m�@r���yR'E?
��E�Țn�Bh!휣��O츸���8�(�n���J]�nQ��̂�$`��"O��E��9
�̬;5�9d@���v4O~��/��Ҹ����@�
\l6����S��=��"O��a6<����A^��	c��>$cC��=����6�0 ��J�A���ʸ�!���(zf�T#�f��d�R0K��!��@�&�~}i��rZV=9���z!�@!z��"��TM�����
m�!�d�$?t ����b7�3s�̆SV!�ę�L���H��0����Q�!�$̄8�|1�d�	h޴�a.xs!��D5���A"G�p��� ���}!��-�n�[VE
5	��$�v�!uj!�
�$?�T;�(�/���`�*>&!���[�:qX�DZ��2x"�o�>P�!򤐊pbx9aU.Z��h��I�C!�$���<h��H�2��=�ѤB	%�!�ă�k�ju�rS6&7T���cɋ �!�� ��'��O��"S��!�$��1z�+2%O6�"�bI�!򄁠NGzuq�g����$�á��x!��-Tz�blY�X��@��Ék�!�)�����4-ch����<�!��	ʕ��]*D�� ��.P�!�D�W�Q��$^�\Ԋ�r⯛&�!�$W�9�F5p��`,���/]8*�!�J	N���
̷�]��ɑ�I�!��J�c��`��`W+��D�j�����P�:��5 �+�@��������ȓf�f9�G��aZ�8�fl����a�ȓf���!�F���5�lj(�ȓb����Sc�4l��B�ό}%L��>�(2ϐ�m�����!����>\n�j���Ğ%�C�K��؆ȓaB���`^�Z���7��"q�4�ȓM�,�R�_�"�D���L2f���?:B�:��[�5DV���e�8KH��ȓ`Phe��"!(��]��'�A�~���TB�%��Ǜ� P�R2gM�����5K*��+�+S2�t�&��RP��ȓ^�9��AB�U�~��%��2�H��ȓy=ʴzEiM-/Y`�b��]�&D�ȓro���6��*��;A�D�k�J��S�? �Yp��`����7��,�����"On����
��Ĭ�����"O`ۃK�2E����$��H}x�p"OL�#��	*��I��-Z6d�[�"O�Q��N�j%䌜�r�P5"On�al���,k��`��D"O���A@�08,2�0�C<~vt*1"O^�ʆ���z,Y���!.�5�"OD��',�+sr�U�&d� φY�V"OL��5`�4l¸�ׁWWQ&U
�"O�l0���N*��)S
�)Q|v�
0"O�8!R��,F��q�S�"jh�{T"O	a��fƞ�1��4I䍠B"O���t�Ў}y��ٖ�2M�-�!"O�X��O~����a"�O+��V"O$���ѐn��d����i.�8:G"O�iPLR02pA#��� A. D�"OXݡ�j��3N��\r�(N״�y��˅l��X��`�6RFFU��k���ybI/$E�1��gݱZ����f�&�y.��}��c�%P"�j�$5�y"� �> �ePWfr �&m@��y���)�Fy��
�Vla����y���M��|`T,݉\7n���ˊ�y� ��6)~��5�Pi��y����yOJ�7C�H�gV�Q��Z��>�yrE�V��-"ՙ<+� ��yB&�=o CDnH�8��k�	[��y���v�jD�� �2�Z�aE��yBoN-��y�HZ˴�Y����y2��� ���j`��=Wa
�P��U9�y�C��-�H=���E���`R
���y�l�2:�9��+�j0Ȁ�m�/�y"A�<;�̀���u'�L�q��%�yr���B����ug��҅G1�y��{���Rj���:Ŭ��y�n�G�l�BFNƣo� h�u�O�y�
�d8���C��޽XrI���y"�%_*��fG��q�bM��yr!�7n��'��uȡ��H��y���tn{��ȜkdmHQo"�y�n�6=(`�S��ͣgiVٹ@"���y�(��I5�i�mܮkU��q� ��yR��m8T���ł4��2�(M �yr�w/�4�s��(�N��Ǥ��y�k� D�iv#�,uzV�3�Ǒ��y2�7/�B�8t�5H��Ձ�yR�;	�l%���X-=��q�q���y�lPF�1rT`_��,�+�M��y���1U.���ߕ���Ӵ�yRNO� ��d曋H<�H��c���y�-�=\��� Ix��q	�yMȥt̤��'��8W.���&�yB+�>O�l�d�4�<II"聁�y��Wg�\�*s+ϵ%�x��f�%�y�%V��]@���b|J�� �yBa��nOHL�1']�c������/�y�c�:`q
%O��!���Y�K �y��ý��bC`�Vu>$���ؘ�y��Dz9pC�Z��Ub ��!�y�DЖ���+��U���0�����y���88 A�ŬM����gU�y�I65-��,�����pw���y2 �Gx� �C�������L�y
� Z`���H��
������"O��G�4:�i��E�8y�Б��"O��Ð�VDp��KP�{7�i�C"O$e�e�ѣ~}&-��C�H�hД�'
`�@�@��#0!�J��񠂄��S��#�/��n�ډ��$0�IʐlZ�w����W�4&`�<��A>1.thR$�h��q�D͑ P[�ea�rҦH��"O�4⃇2M��(��NV*j5�V-��"9v��[N?Yq�7������b�&O�Te��[�ω|�B��4
���5��4_�����K�D��a�0�	_�*e�U�^�(�a{jB�h�R�I���f��5k��*��<Y���`���/�&�"<�v�>K����3�ϯc�̩a�O��y�i_?3F:�,	e�D��Ñ���d�l�CC����3DС"��V+C@ӾpN5;��/Dg�)�"OvD�рӎ"P�}cK�3Y���F� �xr�&2�@=��`ُ.���aO�� �ِ}!�$�v\&O��̅�{�2(p�O	���0���]�(`��� ��@*��]za�5�",OP�K�`�����䗼+�p����'���W�(�~��P��a�E:0��8���#	�iI�4FO�dH<IŃ�	a��3�F݈��M�3�Nɠ�EZV;���Ɗ�hⱟ0�@W'�	��)�Ul!V'u�"O�X�jĉfҨ4�TkU���]q�5@�L�8�K�M�\m��6Q>˓��� `�'UuT݂��N+��ȓQl⴫*Q3h�$$�a��$@,x�'ϨY�0,�Uh���ɦ�l�ã��9B]�W�׈6U~���W4Spq@j�%M���b�%2$���/I�HU��'l��Y�%�(�a���J%�������16��0 0�/��;k9 �P�F6q��!�G��:B�I9=jh9�`d�S��tQ�O|F6�I"a7��ӸF��� eʃH
M{�
�f�,B�	%H���1hD�*'�ƣG�c4؜�΂�0=A�,�$����uL �8DN>�O�08$���G���Wg�k��h��kҾD ��X���xb&4�I��]�C9t�*A	�hO���B�Hc^h`��4lF�B;Pa�R��U@@B��y¤�7+����̙1��݋#�?a�BX�Dش!�=}���+Y/�X���ō*�Τ�����BC�	�I�\�E���ʴ��CYD�r7z ��F������A�&PB"㎧p"Ҩ��,տ>����dW3V������ 
q^�+��P�d�H%�"�Q J��4�@�%$����Ȓ�/t|�ZA�F�M,��˃&5ʓ=l^��g��*|p�J��l���<2�%������J���y�"%X��xR��ѐi�+�	�%)�-fuy��N�i��)�� $��Z*\����=:"���+D�x�O��g���DQ�9�ڵ
��4#��D�!�����0<O��W)"h�`�F%5�b� ��'��<�A�ݙx��]����a\إׂ_А��\N�<�V�R�=<��ÈA�~�"�FK�'b����Ӽ94�F���>^��4�VP �x��&�yr.��q�x{�f��2�v`�(�S�@3�NJ6$h��!K�"~��
6P�|Z�C�����!D
�d9C�Ig���y�ڵS�D݃Wf,�P��{��;$���I�b�����L�V����&�����&����4B��l�3!ݮΦ	�D�[: P���ȓ�2{���!�%)�ąSqj�C�i���S:�E %��,9P��;$�:D��#�OX�#(U��,1��T�0�=D�h@J��G0�Y@�C�AqF��� ;D��*`��;Հh`��hY|]H�,;D�H�eV)e�\S�۔"Yp��,D�@�c��^�(1���s> P�E�'D��A`�G���o���M���&D� T�B>����8mb��ؤ�'D��J5�A7kT�CĸK�����o%D�� .@@Ku��% K'����"O60�̜�zȎ��B1d�����"O\ 0�C� 1��s�#�%Ir����"OX
E@I�e˘U"�ūk҈��"O�8A��R.h�����䁙nI�3a"ODL���L�~j�ղ��� ����"O��A뒭U�̘b��3����"O^��c�2q�B�+uA:h>䴒�"O���e��7���@�GG�m"��Y�"Oq��̾�Dp�&�Sh�ʰ"O*(� ��
R�L(�Cf܊.Ph�g"Ov��W��8��ĸd&J0!�<h��"O��
 �=�8Q�'�*�uS�"O���!��5O�����X@�"OF좒�F�e��z#MC�"�TX�1"O^%Bϓ1�4�k4��iI�=��"O!�C(�y��8�#'2U��"OP|�4L΂g�V !7*̵i.���W"O�ͣ���2�v�c�Iņ'�hk�"O��Y(Ԋ+�*M�����w��Ճ�"O���@ٷF����Ў£l���O�<��H;O&�JF�65�6����J�<�BڈZ��=)dO ���eB�<��m�0����������(�g�<a�i�,� A��6��� !
U�<�Q-�0�L���9Y�ՂAEi�<���H<^ $�dL�=�j��Veh�<	���;A�h��m�9A)�P���h�<�S�$8�@PQ��LC�r%�c�<��kH�T4��<"J`R��Wq�<i���=(�*�� �,���W[�<9��āS~�dsE�	�_X ��e�|�<�W�H���Aō	�bAJ���~�<��ꃓS�#Ɵ�݂i�qh�\�<ɔ�x����ŞN�F	�2�Y�<aţ��,���FeC"-�\͹IR�<��ct�h�p�� �n�!f��S�<1f��y�P��6W�5kaO�u�<���ȸl����LZ9����Zs�<Irψ*�4���8]2,;��K�<� �ۏ�F�b��A�����G]@�<y���XA $#'d�t���`�!ZH�<2'�Mfv3 �����b
G�<9���~&Ƭx�@ĚKe�Y!�O�|�<i׫R;{h��r��E$|E�el�r�<!6!�b�p�q�%J���8r	@j�<�4+�>B:���c/juX�kGb�<�W&6,$64�jR$��1����Z�<�aß�LtS2)P4�\����DC䉺S�Z�	�/��r�S, ~C�)v��t���H
u��p�g�Թ1�JC�Ɉ)+�!�+ݚ*z�C�k�+{t:C�	�lk� 3�6�Z0A��ØE�B��)^J ���u�Ɯ��@_;E�(B�I�oڜ��4�Q�kY�t8$� �+�C䉩?ؐ Q��?�I#*ҫ19�B�ɟoI\��g�3d��҆Aл!6pB�I�[�D�D @Z�&�{�&57�VB�	PL~���:n�Q�]�,B�	�u�Y��J�&�,LqB���C�	�>.�Q'U�Y"ɰu)¾J�C�Ƀ&蘴P��*������"T
�C�I��ek��A�S����tk
�k�����B```���6vӔLPe̌ZN�+�K҂= �[R�Ϲ!�!�� ��Q	ʝ��=i�̄5+�:Q""OX�Y���E�������g��Y��"O�Hq��Φ]L�H9��њ*���b�"O��(��ɜ@����͵(d�M 6"O2���+*��hH�ATvh�E"O���qZ('����fH2{7n%�"O�b��G1D��LhƌE/L���"O ��!�K�/�2iX�*�%x��iU"O�@E��iV�ǉT>[hU��"O6I��v�~�Е(��pO���"O(���NO��(�Th��D��"O�����K�xfSGG�q˞�!B"ODX�`��� &Y�v��q`5�'��0pn��eL�R�*E��,;���F� r�Ì�x��i�Ɩ�b�4��g�O z^w���
B�iΙ)�*}CB�L�vf9�ǉ�b�䘑2���$���d����5/�p��F85�tԠ��Q�W��]���>�QaU#d�P��I��f�x�b0u?�y�7*B�X��'�|��2O~�"�}��b�bLQ�CA�u��РCCP�'H8�)�b�N�S�O�`�X�nD1�h�{�����+�O������![�1��K v&�Zbɖ�ѲC䉃D�z�a'�#���B�.'��C�I�AX��A�˕)T��ys�IG�Y!TC�ɎY�$�Rb�_8�$Bse_8�"C䉬5�0���	�7E�L�u�҅|�B�	'%:Թ�7MF�!��H�є��B�24�:��2��A��x���,��B䉘�3��ÖTz���<YU^C䉡6��`�cM�*	������
�HC�	�y�`4JTȈ5ch�s�G}�C�	29��I�ǂT������fM
�C�I������ �:�\����*B^�C䉿GS|���L��ߊ�M(nC�8d� ���K�V�8!��ڞB�I�d����%�%t,�q�6;�C�l�D��"��U��a�䊙@y�C�ɩ~f�����7��Q�h�8\��C�I:S$|�e�s8tyz��ǘC�ɕY2�S��
�
�p����!�fC�	[�޸�,k�,��h i`4C�0m2���w�X�82�`?C�	�{�^X��낁	E�0-�7i�B�ɂP��Ŋn���I,"��B�&QP�i�O�#�T����
I'B�	�t�Xǆ��;�4lZ�oZ')C�ɤ:(���wA�Lf(�R��=@.�B�	� P���aD$,\2¦�50�B�I}���iBgҷ�!JfB�	�"���F�4m%��o@b�C�	%<|�1ua��P��гF��+�
C�Ʉ~f� ���[�d��Qa��\i�B�ə"���Qō�F��T�K�;@�B�<g<\bU���d=3�����B�I%bѤ����I�i�be���-4��B�	�z��t����b�:�I�I�i�^B�	*`t�P�S��&q�Q	C�Q,�C�ɜ	�~�xP��7i*J�A�^C䉏	"�� ���cT��U"C��"M��L����-����d��;;C�	;u{��фF0'b�����Z�C�I#�t��p�ۜ2X�X��N�5
�B��;q��u:U'�>^�NA@���:%�NB�!>�@�����@8���"nT��ZB�Ir��1�"׬_0�` �Jթya�C�)� ���PSJb�c�4��A"OT�i��l������L/ d��"O$Xc�[(2(H��K�u����"O���d .TǪճ�E!vH���"O�)[W��o���A��'
=:E�2"O|�j�&^.;��u30�e$�e�"O �NI!��r n�:E#�1{�"Oҍ�PÂ,'�B��}ȨaG"O4]9��$���#�L-���"O�\��[�D��,�/s��<��"Ol�a�K����(X�r������yBg�]D88�
J4���$-۠�yҡ͚"W��;�OB�7~�q�y�aGj��.��5���y2x�LA�H�X��T���yB&��� 4��A)��o!��	$@hЬ�Z'��;�� MV!�d�%-ΐ���X��Q��}�!� pGr� `��9n�
H1�DT�7!�S�S��Q�M�ʭJ�nF/QD!��΂Jq*�P�i�q{�!�.ZhU!�$<DBTT�pl�,J�n�bE�^.!��A5AҖ�k��N�X��-*�!��h!��K�P��q棎�V�"]: �/!���H��i�c�:h��RL�}�!�X	C �@�*^�px9�iݷ@[!�D�gcH4��FN,�%��)N!��
X��U�_*d_�h�ta�.�!�D�!�~����ͅi}�uI6� C1!��ǘ�
��f�P b}��X� ɗ/"!�2jShq�'ӓ	h��+��2I!��\'U��4�S�z��Q�τKf!��@�}C~���Ú��.�BC.��0A!�R��n�p !�?�D��f�-Q?!򄖟W��0��o'�*Pc�)��S�!򄁞?��p2�a�<�� �O�!�D�:����5E���"�S��Ww!�	%� ��H�Y�Fi�#�x�!�DیB�F�����W�X�7LCaS!�Jh���B�� Z��!���>8!�D��nŖ�3A�mb\!H�y$!�d
�7��5��#YcT~����@!�
�S� �Ж ��X�<���E�d!�4T��$3B��#��
E\/c�!��[ U����CN!L����Q6�!�dŖO� �S�ݲO⎤ �Ϋ�!�$�$l�P�����
pnh �̆�!��h�
E�����h���UIQ;t�!���{���1���g.ҙ��A�`!��̌3Z�|��B7�D���a�&G!�ȔM-�eGτRvh�<!��P�Zx� AABϮM7���P��.;!�$6_CF="�%b��P�4&!�M�Ԅ
�nJ$K���3�KV�vb!�ټbL%���[�|���*i !�Dk�V�<b��0 j���!�d�#C�T�%W	���si�$}!�׋v�h(�Q�ϼ}�����!��Z.�� ���_�᪔%��e�!�䇳0
��h�k�7y�S�bU�NS!򄞎l�y2gb
2Ba:�AQ� ���dQ1��c�lط09`��PBۻ�y�I
m�$�9�G�/����l\��yR˃6"���d�0�ցK&DK!�y
� �؃D`ٗo��� �ć�2�<XRv"O���$jIg��	��F>\��f"O�`�J�a"lx���9;ԅ4"OP��+*B�j��(��AT���"O$�f޻P64<;�G�jBXia�"O��!���8v�9���м%Anx��"O"�r/!@ X�-53F���"O�)R-�W���b޸X�bi4"O�y��9�(����^MR�A�"O:��g�y?� ���K�!J
���"O�) P,έR�D����8l�
�"O�s��ۼVR`���E/>D��"O�+����"�V���O-�nyi�"O2�D��65_�9��ӹb�Ą�U"O�X��Ė0|����A��q��"O�����(W�L�K��M6 ��Y�"O��r�勲";�q�\64�|k�"Oؙ@�hZ"W���cP�"h��E�"O����Ԃfs~e�$&\�{g~�a�"O^��b��?{�ziS兗:H��˗"O���g�^�e���p ��*��w"O.���!�<���#4,��m �ab"O�Aװ�ȑ�0ʫ[^�xe"Ob��ΐ `��Zg�B/+��p�"O��`��Fo���(�,)h�sU"OV��ŀ	R�$�c�3<XX��"O�q8G�F�7��1��G	H��"O��#r�E�1�N�A����]�d"O�0�l͎^Zh��!�ѤR۾|a�"O*!�!,�6O=������L۸m��"O<H�% � D�H��Γ�
ìhsC"Ofŉ5�M�I���m�2|�:��""Or��5�2&�m�@-B��-�"O|D*F�C9^&Q���Z�~��e"O�5Y��ɉ>�XPS�+ר@W���V"O�\����3�l��e
�$g@�i 2"O���V�®:�D�3�ȇ�i����"O�y�%G�#|ea&mN��� c"O�Yc)W�j)	E� %a�&�)�"O�(Y��?��9 u�����,��"OX!�U�2w��H��V
^fB!��1ik��̀�wJ6Mcߢ�!�D�%{�JQs�%��B�@�T"C�A�!�$U+�8��4n�q��D�O�L�!��0_CȄQ�ȘF�������%�!�D��|8 �*E��JEҒ̆��!�dM {=<Ó�>Tmn�3*��8�!򄍇,���ÂE��,��*3gUJ!��E�"`ak�h�30�x��@�0d�!���>}����دa�N���	�z!�dߴwĔ��S�w��0!B�ja!�*	~$M�#�ۡ��;�*W!�$�P(cE��eѬ5��I�6J!�$�;C�.U�5���d� !4bR�#�!����+��ř8�!؃�߃a�!�4��t�EN���|b��۬,�!��F���I���p��UqO� c�!�^w����t�\	2H��R�R t!��Z;\�� G' N^�`@�V�<;!��&nڐ��ڷy\:a�"��-!��=Ғd��G��M������?'!�$@�Su� K3�Q56hV��r�K5�!�ÏA1�ܺp��%G��u�+-7!�L�X���1!AP<R�r��G�Rg�!�� ��I@"ٜcLxA�D�?�պ�"O��3c��^4�ū"A>:�PȀ"Or�I#���T������^�)�p"O���B��9&"���ӎ:j%��"O�tVG�S,�9��/��H� "OH��f Y�j|"�Q�)I41��a"O �.�wƴzv��^���"O�p�3��7!STE��31d���"O�ͣe.&�zp�S� :�!"OF��7$��i�Ⱥ�M��B�8x�"O>��v�Bt��p��.�,�%"O��G��#/R&�S#�W�ƸX�"O8x:3#��8$�H���<a��,��"O��X�!˽#s|4��׿xR,��"O��ѡFJԑ�"C�1����G"Oz0�D�)r3�@3���X��|��"O�A��+�b���)�>5q��""O�[An߀�
��Ǜi�b�"O�}�G�[�G��|�. 9�r���"O�8Xwϑ�_<P�s�G�ʂ�
�"Op�"4iI �4u"U��v��c�"Ot�#��N�=QL�k�	��H%C&"Op�p� �,����gS�;J��#%"Ox��Tl�a��}�Q,-VӦ��"O�\���W�-B�k�>�6Ix "OH���B��R+���lP�\�2�Б"O� 3�֥^���vK� ���"OP݃ad�z�q���۫o�$��"O��a�   ��     G  �  �  �)  )5  t@  �K  �V  #b  Tm  �x  ��  p�  �  �  x�  �  ^�  �  )�  l�  ��  �  ��  ��  \�  ��  �  l�  ��  M � � p V �% z- �6 �= WD �M U �[ :b xh xj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>�z���瘝 C��rs��i�99�E��^� �O��oW��|��?�Q�952�b��d̔��&*�?1��MO��y�4��Dm>�������sXT�0�
L�VeF�˂�̕(�c����Uy��S�:��MB��v]G�\f�[ش0�M�<����Kw���?�m3Q�D��	��F!�X�$�Of�	`}��ʀ,r�F<O��(�_�S��kejC3&�	Ie5O��I:�?	a�;��|R�-�`�P��O�]F!: �y�,͓��� �$�զmp-1扉��Zj�{3. ��.H62uj��?aV��	�t�S�Fٴ(��A
���N4���������O\q���%9�1�\u���9����̨aSJy��[k��(ɵ��=v�ʓ���O?牟uhq�:)�J�ƥ�m8�扉�MC��i~R(d�N���,غ�$?Z~e��'ש/d>���H�	���QiT٦�'��K�?��@�V8]�|��F��mK^�SE·@%�'O�i>M��������$��7"�0������={4,�>Y�\�'r46�=G�����O\�D)���OP,s4�5ز�r���1���vdZr}��'B�|���� >-��N	(p����ÞE9���V�S0������^H���e�ړOZ�Z1�|�d�$����@�B|B�S��?���?y��|z,Of�oڑjv���I�.��6�$;ް�������x����M�J�>Y��?9�=?��+Ӭ ���p���Za�穈)�Mk�O˄����z����wYNcC꛳�p�ͥ6I de���I���I�0����
��7!%�0V�D�7	��?����?���i�H��ȟ��n�e�ɘUl���h���Z	���S�4�%����ß�(P`Ymn~"f�[���Ca�h���z�ֶ�N�ȐJI~?	N>A-O�I�O��D�O��ɖ�C"�,e3r���a��م��O���<a7�i4�aC�'���'��ӟY ��`��jx�q��߼^���z���̟��IN�)*f��_1��!�	/A��5x�[�3a�	�dd��:B��R.O��?q�j0�d͹Z�����Ǌ3�HLږ�ޅG*��$�O�$�O����<���i�+��|u��&�)��j�����������ڴ��'P���?ѢGG�e�v�����
!;�%E�?��m��5Pڴ��D��J$`�c��d�A�v8��;>I��4����y�Z� �	���I�����0�O2|�`���,��
G�)��	��d�LE����OV���Ot��T�$�����%n���: d~pٱ�T�,�*]�I���'�b>5qu�צ�MČ��L��tJf�8g�Ȼ[��͓
�d�۷��O���M>�/O���O���f�d�U$Y<�TQ�Y��<��ʟ���FyR|�t\��"�O<�D�O�Pz冁=i��M	f�1F
�h��J(�	&����Of�XBt�џ|yɵJE�dj���	6?�����.�T�#gS)��',���S��?a�/�;rڭ��#� =�@�vo'�?���?���?Q��	�O���1oni��(Ͷ`y4�{�A�O(�o�3Q�������4���y�g8wY���(G;���u�̗�y��'��'���ـ�i���"l�~�1�՟��w!�$T4,1�wU�+����!�d�<�'�?1��?����?��@�wJ��Ĉr2Y2�A�*���٦��$�����������gKCr�ZA����!ud�9"�&�����柨��Q�)�S�7H��f�Z#O3$@��BГg	2�ߦ	+.O�<Knֹ�~|R[��H$��	���X�`�<3@H�#��ş,�	؟X�����@y�NiӖAS��ODu��j̀)�h1�ţ	�Q}$qa�*�O6lZo�0�I�H�'�`ÈݾT<�pP�A�%iL�ժd!J)	ߛƛ�4�6�R e��/]�S��� �ez"fB�.���A]!;��+G9O$���O��D�O��d�O��?YȔkĘ�hǯS����R��ğ���ȟ���44^R%Χ�?���i��'�����J� $I�(t<���y"�'��I�F]0@mZd~�+�������H[,yb�O�`����ʟ�$�|R[�L�I���I�(Jde��2a�@�tÆ�;�ִ�ů[���	Qyrmr�j�� ��O��D�O�˧9�D����j�� �L~\���'.��?����S��DȜQ�,c3AͤK� ��EɁnK��Տ�5F�d�O�i]��?�$�0�Dψqԥ�+�����o�=gq��$�O:���O ���<�iz�JP!½!Fl)�w�;e��u�!��:r�' J6M;�ɶ��D�O�)0r����aQ�-l X9����O��DP��F6�&?��F�kGP�I:�dlL�|e�TK�v�bP�`,�yrV�`�I埘�	͟���⟘�O��$k��H]D��!c׳1��tk���ɫ<�����'�?	A��y�e\=2e�;�:����!�Џ9R�'�ɧ�O����R�if�� >��rEd��G�H��w ��]��DZ(MD��[�� �O���|��#���� �ʃLV��+�%N>��!A��?����?y(O��o�0w�1�	��ɨMY��(ٛyІ� �m^8cn��?�@\�X��˟�$�D(a���w5h�ħ��j��u'5?�gIJ�%���4ޘOHD��?��B���y"�&=w�萇�,�?I��?���?�����O|�SiE������/}U�e ��O0$mZ2���'��6-"�i�!��C�2!��m�ì*������f����~yB�Q������I�(��C�T%Fd�����]>�0�
E ��U'�4�'���'���'�'S������}$��.�R��T��ٴA�r�����?���'�?��j
24A������;o"�:�#����؟\�IY�)�Ӎu>�9��A$x�A(q�8xFE�2��3G4��'��E,ݟ4�@�|R\����F
	Ab�iTI�AF-X��]ݟ���ğ���֟�Lyr�u�vɨҮ�O���¦�P��L��&y�ҙ�S��OTdm\��h[�IΟ��	�����D�~�+2�M�%U�T	���.SR�\�+���RE���>��*ix����Ҝ]}�<S�%�.F�F��t���P�I��p��K�'s:h=�7�7y���.[-<����?��Hƛ� ɔC��I�M�L>)�BD�C�eK��U?h?�xRa�T��?Q)O6@s�r���+(��C�:]�����Vz6*XZU!��<F���@��䓾���O����O���"cfm �N\v'�𑑥Iw�b��O�˓;Y��!ޢ�R�'W�T>)�W�3e�Ĺ;��<; xH��� ?�PZ������ '��'Q���0��^���3HĿ9���eJ�;�f��˝j~�O(��	9Ua�'c��f�L(s�`���K>��V�'w�'���O��I��M;�o�`S6�a1��<k�.$�����[��u���?	��i�O���'�OP�^�>�����( Y�P(�!W^��'�LS`�i����~m�S�O\�:����E�E,� �f!=JCv	����O��$�O����O2��|R��_&&n���+�(oS��Sq�I
H���eC2w\��'!2���'�j7=�f��t"D!Ml�=c�����%s�a�O�b>�2���=�mDT�uM�w�ڑ���[�zA�1Ox]#@�\.�?�n:���<���?����%�=p�
A�K! )+Pf��?����?i����$A¦�Q2��@��ҟ����8�J�QQ�I�JD��(�"AK�g������h�eW���IŹ%�
��1IS��sK�$	��0�M�&��DKw?���:�I��#�;z���` * ��r��?y���?����h����7(�<`�2
�� (zѲ&�IJ�d�Q�$E�D�ɔ�M#��w'��C�*��]K7�̢u�X�+�'�B�'��)��]F�v���]�u�\��3)( 2�ƹd�%q&�[�5��Q���|rU�,��ϟ��	ğ$�	ßD@�Λ� Y�� E�3VDz����Qy"q�Q���O��$�O^����ɫ�����@�gO�ѡ4׽. f��'G��'�ɧ�OM:e8v�^ M��tX��0��pß�k%����X����q�D?��<q&J�u�N�+�K�"z��=��G��?���?���?�'��DQ�Y3�����q is"��E lA�!D�| 4������C}B�'YB�'��, A	M�@���"Ք���(����f���g��,%�4�	��R�e��,��%���Un��LI�6O,���Ot�D�Oz���O��?�Q�F�	�J����#�v�e@�ڟ�������4�&��'�?��i��'b��y���}����װ	����y��'�	�^�t�n�c~2���z]b�e�d3�U+_�)���Xh�~I�I�dz�'���ޟ���ȟ|��N:0{@BȌ-��� +�=7�M���x�'a�6m� �$�Ol���|"V&N�[�n��d*�4o��5KV~���>��?�M>�OxJ�(�*�����O/W�:B���!\��i����|�a`��l$��Aa��s���
,�ld�%%�͟��IП����b>��'M6��7S������Q�0EWS��\9uͽ<1`�i��O�Q�'�� �I���8�͔28f�Yg��G�b�'�҄��i��iݱ9��T�?�Y�W�� r�����=n2�q�E��rޞP(t7Ojʓ�?����?)��?Y����iC�^�����,�{FrEr�ߒuBtm��U�	����G���H����`&�=CDV(m��g��?����Ş��Y��4�yB�A�>#���Wd�)�j����T�yb��|U�a�	�xD�'Q�Iџl�IU���Z�$ɌD��/� S�,�	�����ǟ�'��7M�BG8��O�d�Wtڀ ��%<ޝ��lY�h( ���O�$�O֓O�Hsg�̡��E12	�S�,�瑟�ba:0��LXo!擿0��oAП|P�B�/�t "�iP>�l���ß������	PE���'����f'�#k� ���c�HȠ%�'M
7͚
1^~���O�oS�Ӽ3��$��h0�K[҉�����<I���?���J5�u{�4���Ӗn"�d���S��%�ִdI�8��,��o�`��,��<ͧ�?q��?	��?م��� Ƃ����g��5L@5��D���Ґ���	ӟ�����%�@����qc|�0N
6|��ǟ�	y�)�*�<  +�/�(Њe����Pyq�K����ٗ'dN�Cń���"��|�T�x�F�J�&��a�2,б���C �U䟔��ϟ �I���S@y"�b��)�J�O�d9$e^�z@�yzV^({[e��7O�o�w�|��	ğ��'sd�BC� �.�yF&,d����і8��v�����R��TH y����mۄn̻-l�;��_?8
���bp������Iğ0�������2K��ݢ0A���/q�KZ#�i�	˟�	5�Mk@��|j��9ț��|RG\�(	}i�< �����l�Vq�'L���4�����V����&J:mB���P��0�L�C�eԊa&(��v�'�
'������'v��'�R�ӣ�=��5��Q�q d�'��\��:�4I���I/O����|2ワ$.J0���T��j� ^~��>i������F��|���|�2�I��V�h��@uҦ���ƾ<�'���������zhP6o�=y�R��#'�2ߤX���?1���?��S�'����H$�O�2��]!�R��1p̕���D�	՟�s�4��'X��?��@�UV�����#V���Ղ�?I�e�R��4����T��K���/O�m)q�͏�hJw �k8�T�#9O�ʓ�?���?����?�����O>�\�8C�� CU$��C��m��\f
h�	ş��	]�Sşd0�����,V�̼��V)������Ζ��?�����Ş)�"�ڴ�y����Y�I�r�c�ݣ��]
�y �.�$U�I?��'���퟼�I�pDXxPFg�(Į��I_3�Q��֟��Iџ|�'a�7-�ր��O0��ŰX�� "&G��P�،W�-&�\�쨭O �D�OܒO=ke�0fpQ�Ѩ��e�ЪR���ԧQ4f�Vl,��'`�l���<����.bv��I��$:N&����R��<��۟���̟�G���'f���ҍW�:���E0���C��'�p7MW�|;���O:�oZm�Ӽs@�Y$I��;c#ڿ2XrxɇD�<����?i�����4����^�%��O���AVE,��*����![<(�ӛ|�P��ٟ���ϟ�I��+�'�L�L��%x�=��b�jy�f��$m�OZ�d�O���\��ތt�v��6`H�-��D�%�4cW��'���)�>�zDsW`�ek�|8#��p�l�i5�I�uV˓d^�����O�AO>�)Ox�xQ��)x�z)Kg@b8�}9GC�O����OZ�$�O�I�<��i�~q���'
d��O�_�d�8V#ʠq0���'�6�<��9����O"�$�Oά3�C �L$؃F����3��@q�6� ?qc��9�D��V��߭���&RZ�C�%ߟB�|��4�u�h�I��I����I����#BǎV����@�˽R��1$ߪ�?A��?���ikD	S�O�r�j�>�O��w&S�>W�aa�Ɔ(^�rD) ���O^�4��a��o���el���B]&/�T�H�/�8�:�0ӥ\"3/��	X�	Xy�'K��'Z�'K�q�Q!t+�8+PJt��Q :#b�'��ɪ�M�ׂ�8��d�O&�'���)U_���	��X@��'�2��?��ʟu����n4����	#X��(��Q�+{�}Hq��* ��|�ׁ�O`�HJ>�t�K�{��ːg������?a���?���?�|2+OR-mZ��`!8��#Dt�Ŧ5UhdQ2*�4��
�M��ͪ>��NR⊙�'�<��3Ӟ�P`����?I�b�=�Ms�O���nK���L?�HB"B�'�^�2�V=aȌ�"�l��'���'{�'&��'�哜3~�9��!�8��aB�I�D�� Y�4S�����?������<Q���yW�^�
3�%� �N�k@���w2��)A)��7M��ɥ���!	���-Y	/Ű���#{����3
�[_�	sy��'E�FO�,+��6�ψ]��Q6�N�8>"�'�R�'Q�	��M�W��.�?���?af�W'�֬�4& �A|�i����'#���?�����za6E��H@&ڊ	ѦD0x($�'+��Ԅ�;�x���D�џP�R�',5�TI��@��U��Ȯ0������'���'B�'�>��$XL�RoРʀY�F,]+]�@�	��M��K0�?q�x4���4�x�P��C�R��6���W���>O|�$�<Q"��Mc�O(����Й�z�� tqh�
� }��#b웋�l�9um>�$�<���?Y���?���?)2�	/͈	��Ƙ1O��7`���d���]�1��}yR�'b�OfR�ƎMAdTS�"֩:�Z�"��0H~j��?����DC�xY�%�%�C�8�6���;�(�94B�P:��$�@8���'	B�%�4�'-�
ƨ��jƁ!돴y�P��'���'�����T\���4u��LB��`=��`�#�h T)��)=��̓}<����O}��'22�'��yB�ה"E�Tї!͡�����������R2�¶w��!�I������@��b����+��<.n<�R3O����Ol�D�O~���ON�?3'��8�0���7.�f:�N��I����۴b?\m̧�?)0�i��'2Jt2A��id�̸ �Z7ze.a��|�'%�O�n�ʇ�i�Ɍ�L �dL�{>�b C�I��9�u��L��0��<�'�?	��?1 g6\&�Mq�mJN�����_��?I����DĦŠ�![cy��'W�*xr�A�Ⴡ.R��[`�%IPX� �	ş���d�)rE'���('	(�9c-VtFX�"��L�� +O�	8�?A#%������A��	�dL���4H�d�Od��O���)�<�d�ixV�f�"jA�%�K�F��-	Í�l"��'��6�:������O���KՎ
X�P!JU�rj��:��OP���<|��7�/?��'X�X)��wj*˓)%`SF�]�� po�	�M����O��d�OJ�D�O����|�W��o^����1�"�ض��b���lŞ|�b�'�b��t�' �6=��\���G�z���6 �h<�(���O|�b>%�DEئy�_���9`f�l(�#����0�f�0��&�O��J>�(O����O�@A/ j��,I��/*��д�Ot���OX���<��i���z��'���'��q�@F4��x*��� 
�,!��$�S}�'��|b��\�XT�g 
h��LJ�`ĉ���@.�b���oш\1�t����\����%l� ���Y�N�XDГ��70�����O���O��:���b��	V\Y�H��P�(����?)P�'�^����?1��i�O�.�6���&g��p�DJ9���Or�D�O�]�mӨ�4� 1Bn����l�v&Q��E�B�����%H�����4�����OH���O��D�c�6�yC&51��E[��]!P.˓	���g?�"�'����'+H�jү��t���5'رz� �ʹ>����?�K>�|�T)�
{�Z1��+Z53������n4p���Tf~���j��I�L�'�剆@�6)¥��;��iF���:pJ!���L�	̟��i>y�'
�7-��8�<������������"�/�`0�$�a�?QbX���I����I'`°!rCI�,�SU/ʍC�Px[@#�¦��'5�B�HX�?�E����w����gF��\���ȃ�(�H�`�'x��'���'���'��1�.\%���k�����&9�?���?���i&�Y+�O��Kw�$�OfP#ʘ+]�fHX�lĎk�Z�hcm7�d�O��ԟ�@"u�i���� ^D]kg�؀t�@�sRl��=Tl2$F7vR��~�	vy�Ox��'���Աٖ�jb*�F�ԑ��2�'���"�M�M��?���?�-���3�N)��y ���u iS矟x�O`���O�O�SKz"��Ҡ�5���ԁ�0T�M��"%�:��*?ͧJ����E�\��h�\餽�@X����s��?����?y�Ş��$��?�(boJ��Bԑ$�Ӭ���h��� }�F�d�_}�'�,�A���e�]� M�[�����T��r�mզ��'�TQ��?��^�XȤIK���H4ꂬQ!�h1�w���'��']r�'p2�'k�S0qh��\ vl����Ss_��޴"yV�+���?����O��7=�b�s����|Ԭ�[& W�h�J4Ѧ+�OX�b>%�g��覽�?��02#HI�
�K�$ޡ0�θΓ3�����@�O�BI>�)OR�$�O@��pF-]&9ۇOۭq�0s�/�OJ�D�O����<���i�v�ɗ�'Y��'����lϯ3r������1���"���HV}��'��O��	���G<��C6e�H6�h���@��oJ;d������k��8e������
�E
c�at��yW�La��U�h�	ӟp��ݟ�G�T�'���'��6EhaCu��:�D���'H7�O�J���D�Oؕm�P�Ӽ��Dޏ|�B�ʠ\'*Z��O�<����?���HΙ��4��DJ�~,T�{�'|?�A���04p����bTe9��<�'�?Y���?)���?���/'�����-UW����������,A`r�'B2�)6$��T��L�$O��r�.F�BA�h�'���'5ɧ�O8H�sՃ#�U25���(�v����(ؙ�O��V���?�3E �d�<9%с>�"�j�)8L!; kG�?���?���?�'��d̦)[f�C��h�aE��j9b4c�1u��E�o�Ɵ�ش��'�6��?����?Ƀ�[�>����YSM�ҊZ>�JA(�4���K+B�$�����O}��۸V�l�R
ռ5Xt�E&���y��'���'U��'�b���$L� q牕^ ���ҁ.�,�d�O@�ĕꦝ�a}>I���MSM>�PG�&o�����L��Ji-k삵�䓪?i��|ƥ�0�M[�O6ԑ�� �U�憎i �'���b�;`���?�6 "�D�<ͧ�?����?91(
?.qM�w��<?ऺAa�&�?�����Φ��ǡ�Ey"�'4� ��A��%�\Y�f�)��[I����8�	`�)r�"*J�~�HX�VeA�f+��ڰO9h�����@�џ��|�e�+A�H�vg� �a�H1NyR�'Tb�'��^����4z��\K�eR#He�<�4�3I����/���?���6������l}��'��-sq�Ƥ?[�h3fCR;VC�!fU�������'�h��e��?�c�P�ہk�5|��t;wA���M/t�P�'�"�'�R�'�b�'���w��|����	N��h��TX޴QJyj��?�����?	D��yGEK!;*r�h���&JZ�B#)ŀx���'ɧ�O;Hӱi��I,eABuh�%�"�Z�z��JL��T�&[|< �'�'=�	ǟ�	�ı��k�,:$X�P`
u��	ٟT��ß��'^,6��-ʓ�?a0"L S�<"&e�	-%���E�H���'@���?!���_c���'cת����j�
�@��Pi'b�5P�&Un��'`�F����b+S�6�"�oJ>��7��x�	矈�	�hG�t�'¤�	B��W� ����(h����'?�7�\�<���Or@o�O�Ӽ�e�L5^�0�Ǥ� &�� I�N��<���?q�HL�� �4���I>@z�3�Of�䒁�I�PJ��s�P+���Q��|"T�������	۟x�	��4�&Β.r	j����%_�:�Aw	�Py��j��Bǁ�O��$�O@�?1UF�*m�D��kJ�v7�:#g.��D�O�7���6��1���<DC%(���n�v�d��O��<'���'L��� &,��"^�~�8�3$�'j��'o�����W�T�޴x5Jz�� �0�Q·'a��駡M�10P���N⛦��x}��'���'+8#�ȅN0���BG!o��K���������Q�,�����	����:��e������g'��ȕ6O���O6���O��d�O��?�j@d�I�H�Z�v�� �l����IٴBz��'�?I�i�'8����B���x{wa����@ɢ�|r�'��O�:�葶i��I=hR��=��qs`�ޜ�L��ȥ���2���<���?1��?��&�O���y@*<A�l�'(P��?�������f`���������O��$��=*n<�e
wzD��O���'x��'cɧ�	���Ł��%3�F�U�L'(�2XA ���Xb#���S�(bF�H���
�����J�jx�bS���)�I��(�	П��)�Gy�aӼ�8�#�'v�n-a&!�A��9����#>���OlTm�t��fW����4k@CőXau���˲"�mh��M�<�I�r�.tm�t~�$VF��4�J�)�	b�0��C�Z|&���T5LR�d�<����?Y���?���?�-��y��KR�zq��y���;Z�hT�tm�ܦ��BNԟ@�IΟp'?M�ɳ�Mϻ`V̀p��P�O�!�"�Ҏcf�
��?�L>�|��F�M۝'�0U* G�CF|+'�^�'�A�'r�1%��{"�|rU�L�I�Q$fUh��Ŋt�W�'f��CGZٟ���$�	wy��V���k�<I�[0��F�@���*V���a ���>����?�J>i2��8[e>���;��q��~f�5w��aǓ��O���	uL�f�8Ĭy�
 	i)�Xyf�ܩr/�'���'A���۟�@���n�D���\5�=0���͟`�ߴ@�U���?	��i�O��(j��u�܏J��H�A w��O��$�O��)��s�0�4��t�ǥ?�Aq��-=�5�� u��N�Ay��'Zr�'+b�'RFʄ(���2��.��xP���@*�ɐ�M�u/�:�?q���?�K~z�2W���ԅ1x�l!�֜>�z�TU���	���%�b>=�`K���2,[�2���9��,7���Ka�)?�s�Z\oB��������D@&%�P�X��eDD 2r�٥ �<�$�O����O�4�l������f �I�����Bvʟ"\xF��H�B�x�J㟼:�O����O8�č-"h�����-�4��O$rr����u���=}0��s���4�>���~b$����n�:P�T�C0pOt�I�����˟��	؟8�	i��)\S勑�wP�F�-0��j��?!�vH�f�H����'6�<��'\ ��q� 0P$���1O��D�OX���}r�6����< N�2���&
��ݛF晫�,�!�G^/BN҉�o�Iny��'���'���T�;�T@փ�?7�6UIa�$:���'�	�M;⍄�?���?�+� ���+ۮ#�� i� s�hy����R�O���O��O���	ȚᚂN�1'� s��^�6 ����uS���b+?�'���Ė��`��� ��,G.pI��̺*�b!����?a��?a�S�'��d_�)rAmE�~�i�D.J�-�p\kC��T�Tt�'�6�;�	�����O�1@��F�\j]�`dƷ7&��QU.�On�d��
4Z7m&?��qBU���2&�L9dp�)�8��5���>��ϓ���O��D�O��D�O8��|�P 1m��E�.WB����N�9)�& �5m��'�R������;A�Tĩd>R٢��
E�9�I���&�b>e#1m
�u�S�? �iso�>*�l����>�Q��;O���G��?��<�$�<�O����CND|k#��n�����o����162�'��O�/�.�Ir�T�d�`S����s��O�|�'Cr�'f�'�p�1�6@RL`��� =|�5R�O����Z?Ŏ\;�C9�Iؿ�?i�c�O��˕
7�l;Tk�4�$�5"OH|��n:r7H��
²&`}	U	�O�o�s�VU���|�ڴ���y�j��o h�5N:���cf)I�y��'SB�'�F��i�I�5��	B�ԟLA'��gbP)��P�,��QJ��=��<q���>+>��Y�m�4y֌�KC�ɽ�M��O��?����?!���VU��D&V�q2�A�D��l��?�����ŞC��e�Qf�rY$K$�V0#����M��Z���,X$-��<��<�hC?� Tc�`��+�l�Fd�~��IٴW�$�3��7#�q2f�K�
!^T���
{~D�c�D���d�Q}R�'6��'�@�b�j�q�v��Ӊ�=�,��n,�v���� F�2��T@�j�S��M2�K��T��k��
�X;���Ro�|��I�?;���Ճ��O�xh0�	2,����ߟ��I��M��W\���s�@�Of�8s� �D�1w֕s����)&��O �4��kPCh�D�"Na�G�)ZD�kD��F�%2g�My��	q�	fyR�dl20���٩P�����͡C��XYݴi��q���?����򉎏!<|�[f�M�@��	�P�	����O(��7��?���/�3��+����]��L;h��y5BԦa (O�)Y��~Ҕ|��N�`i�m�t��1y���:��Np��'<��'���\����4	
X����X.���e�<��Ч�¼�?���{\�����W}��'{������'=���(�$8���ѷ�'���F''�V��4��M�6��)�<ya���\��dE��sw��g��<�-O��d�O���O
�D�O�˧(?t�:!�(} �S`M�G|[3�i�$t
��'d2�'T�O`B'`��.ͣ0:����\إ�S��2��$�OT�O1�f���ad�x�ɴMd����&yC�Q���X!��	*M/�|�w�O��O���?Y�6�څpLM�^0�IC�`ߴ$X�Y��?���?a+O�o�8hӦU��۟��*[L~�-�����aVcë	[�?�Q�$��ʟ�%�X���W�Qk��[4�W)L��P�P�/?�h�j��y�ݴ5�O�0-���?��o۬ 1 �k"��+O�@��1nW��?Y��?����?���i�O�a�%��״�xf)�>?3�(�$"�OP\m�2g�.���ܟx��4���yg
ٵ��9�#A�?T�K4mO)�y�'���'��ً�i0�	U��ڟ^�YeJ
�Rs�@Ȱ�9T�>����,�d�<9���?���?���?y4�֌A�E���P�~�@0sM�����٦u+���꟔����%?��ɹ"*];3 �^�|�J��آ2� p8�O��D�O�O1��ax����v�!��_Ҩ�ha��	f��7��\yR%D[�L ������8q�sV�śp�����ڊRɠ��O�D�O��4�8�4��o�'d���3�f�$��*�h|J����]�b$fӎ����O�$�O��d_�H����jM�'�ܑ��j�8.������j�x�y�8�z���?�$?��ݹZ����w$W4���'X d�蟈�	�8������	@���]Q� \jD`��1e�H���?������������'C 6-'� �Mk���j3Y��=0��R�A��O"���O��ܴ$��6�:?	@d�<B�IB�Y8L��ݨ� hѣ���$���'82�'��'0h)��گY9�a��/�D!(��'��P�lٴUb�����?�����$�fmQ!)YB�����f�4a@�����d�O��$6��?i:PI�8e����#�!�fH���Ŧ�d(�����1r.O��|~�&�4"��Y��1�O�+�2x�ѩ#��Bٴ7��ܺE��o2���`�
5���;#��-�?���f�6��C}r�'SLeK�A��|�-I��	���"2�'���{@�v��|�d�fO���<�G-� .p�`�M� ���0F�<	*O�����`�QH4�N�p� FE��S~�o�/I������|�	c��t$��w� %��E�O��L�6n� elݹ��'��|�����ʛ&2Or$q#�
W���I���(S`�[�2Oꨠ���?�2%?���<�/O�Tg@�� \l����x��B��'�7�Ğv���$�O���5:ة�p�O�p���r@���qY��<��OX���O��O�0*��H�,�d��Z�T�&u�s����/�,x�l���R��Iџh�3l�=*�H��^+�|A07$$D�Soԋd�jѓf	�vBE�E�p(�4~2�()��?��i�O�n�1�(p�A�Y�$���OOl^��O���O�(9Dw�J�H��s��?��d΀�.������t��m
BGn�y��'���'�"�'��9�xsF�òE�޸�� )w�3�MCcaԭ�?����?�O~���W�4zr-љy*~��V��y���\���	ğ$$�b>e#�L0� �!��B�l{����Js�����
2K8�I��>9�S�'�p�$�4�'��e)C�߼:}�����I�B��5�'jb�'i����TU�LQ�4!A"њ��f��r��'�ZHI$eL�6��b��L˛��DLr}��'��'+��ڱ�WQ�D13L�1���J��6�����JT�ޏ0��)#�	��T�fH�h�KF��e�E�4Ov���OT���O,���O��?�b�#��n��@�X
2��0)��� ���H@�4"%@�O8.6m"���"lnX�x���]����%��_o:�O��$�O�ɗ�	�7�5?���B�2�G)��C�ҵB�B��I �T���8'�D�'��'W��'�29�BEӿX��! k̶
֦����'�^���۴*yj]�(O|���|����7o�p�˷i�Żc@�p~RE�>���?aK>�O����&ݳ/B���c+w�0Ex�K�_�^i�úi����|"�ʻ��$�������5p�R#�Pw¡�Vݟ��	����Iڟb>ŕ'
06-��*����$Ȱ`�dr#K��F��r���O������?Y�Y���FiP=�#BZ-x:}(��T�$�r��Iß�bY���'���*�O
)O��2�	�a�6Ts��w��hv9O���?���?���?����	K�rm�����q��L�^��s$&k����O�O����O�����D����q8�e ��ԥ��e��n���IޟL&�b>��II¦�͓!�45���!%Fh��D�H`1ϓAX�r$�O�$XH>�*O�I�O�9갌�Jr��TI�+��+A��O�$�O�ı<��i(t��'���'�&{�EQ�n�6���fu8f�_l}��'oR�|")� zW�X҅ɍ=^ ��ߤ��D�zd�SU/U�L�1�@�{��I�&�d� �Ę�O��c�ö�}	��D�Ot���O�D'�'�?�4nW�j�L�5��� AX7�S��?)g�il��R��	ߴ���ygj�:�:�ze��,n��[� �y��'��ɯx�
|lX~�I
���S�:��-Q�*�Rb����A�������|�Q��������ϟ �	� ��fR1g$l���tjNd��Kuy.k�@t�g��O����O����D�3�xdi���Q*j�2H�'����s���p�
�Dn�D��?k� �!N�e�0ʓ*��!p#��O���J>A+O�E�� �(��|�ǛoJ��L�O����O���O�	�<9&�i(��PV�'J�,s��_=؞᳣
U0y��X��'��7M:����D�O��MTbY�畧t�M(W�R�J��@y'ʇ��M[�O(����R�)4������,[?�\����0���3O��d�O�d�O*�d�OZ�?U3�Ϛwm��Y�LK�M;(���D�����ݟ�ݴU����'�?9��i�'��������҂�!z/:���y��'��I�"_D�l�P~R �YM�\ �9�,QR��r����ğ���|rT�(�Iԟ ��؟���	S��e��L=�ي���� �	ay¨g�p�#P��O���O|�'oo�A��OBK�f�%N��:K��'m���?�ʟՁ&�ΓNS����B�� ��QsBܤ:�z;���|"S�O����H���x����V�`�3H�"�D��5�%��H���!�l�@C��Wwf�)��B*��z�M���К���?;�j�Jg�7ze�jF�q�d�ٓ'HM�l���*�HO���ιm5�ș�$�%B�8�2>�l(�!��ȷ(�*y�(��ɋ�B85��S5)H���P��!}����'�!�ƅ2�#�99����(�'BP(�r�H��r�(�bWΓ�C�
��ET#a�\)���)x��Tʋ�n
���u��B��}K4(�w��%;�n�	#3<$���#����3��4*���'�����&�d����x��� L��,P�kR9���bb�Μ]��&�h�	ן\��By�bh��	w>�P�ř�I �O	�K�^l�-uӾʓ�?M>��?����~�K��&�̳��ŀsJ2�����d�Oj���O2ʓ9y��XG^?u�ɝ&�P�����b5�zGD+/5T����$�P����\��LaܓtlpZ�ᇔi� �LF�2�lП��I@y�ꇞ6�>맂?)��b�	[=��� 'C���`dH9�'7B�'^Z�Z��$�?u��
��@g�H怟
jż�zU�`�X�_�rU�ѵit��'f��O������Q�a��s��� �c��9��������X����OW�Y��FN4��	�4_��} �i&��[��s�r�D�O�韄p�'���);��W��":2.ܐ��Y,�\���4^��y�����O�k��F64:��8��τ`0� X즵�I՟<͓� ��O�ʓ�?Y�'p���f�1]L��q�GYA�$�ܴ��u�`L>���?���f�P��}COX�gu���̦I���)ЯO���?II>�1 �`q��cW� aXcCO��bh�'<�����' �	���	����'0�y��cLT�Ȕq@`C�<���r� U���꓀�$�O��O���O��P����T�~9����~~�թ��WTᲒO��$�O��ķ<����*2�L!h���hC�R���:��R�\͛V]���	a�	۟���;~�v����K0R�@&ղB�����b �<��O���O��Ĺ<Y�#I�����*˯r$�5�#�QG�%2���M���䓆?��pD�>�U`b@�1e�&R��	������1�Iʟȗ'�@"0a'�i�O����lࣵ�ԑx���f��O(�@Pu�x�]������$?�i�� ֡��g�8Fg��aD.�
DHmCu�i��.�V\:�4Z����8����DF�i�xպCj^'��L(��ԑ%n�&]�4���qK|jJ~nځ/����OёZ��1�	�	6�GQ�$nΟt��Ɵ��S,���|z�O?2�n|��R�)0'M�jۛv�'�2�'�ɧ�9O���˭7�,�[�m@���T�l�g���m���	џl:������|����~2��:?�F0 gD�2~P|Q��V�M3������3?����~rm>,��e���=tG�`�tR��M���0mdx�/O�e�O �O�aa�mʹM�(��!,�n�HP��+�D≑m"�b����]y�'ӄlHƅ�gvh���Ԉ'�
���d]���	C���?i�'Q����#�=�����  �H�2u�ݴiʊ��<9������O@0���?�j��i|�mz�DH1 5/m����'y���Oʓ;m�HnZ�7�4��'�σ2�~��3�@h1H��?���?�)O�KA�O��5E+a�5\��p�EE�E���h��p�^�D1��<�'�?)L?��p��G���X��
�t�!&hm�`���O���&ex����'��\cβh���f�E
� (a(��M<�,O����O���������������X�Ļ� �>���4������?!��?��'���T%	���b̚8Rpx"eS��i R\�|8��$�S�S=^u
qY���+B~x�Q���NI7�X=*�lZҟ��	ҟ��s�O�N�C�ne�&�J�@x�a��Jw���m������\%���<��Ytq��Y�6��q
�����s�i��'!�.68��O��f�OT��T)L`�, �)?}Pտi)��|b��~��?���?��%���AC���Q0_/����'�7+�d�i>	��v�B#��Ӄ��<�R�ӂ�G� ��-�O<�����?q/O���G����!lS#|�B��c� ?-$�S��<���?����'��䖨S4�+DF	1cE85�Bɚ+����U��$�O���O�t,གG8�ڐA���d�2���C�8X�Υ��V�$�����&� ���4�'#^�9u�Ī>��#&G�c�u��j*�D�O^��?Ѣ�[����O����Q.2���u$@�xĤ�bA�Ϧ%�?����ğ3�'�A�r�X6U�dDP! �N�H�9�4�?�,O&�d��$ɢʧ�?������ph�lxvA��&����}�>�'�H�	wy��O��R]�t�� ub`��GI;\����H��&����������?��u���*6�<�� )W�K;������MS���dR;Y��Af�G�9�Pt{u	Y�i�*��'�iz|l�ky���D�O��D� '��2CD=:�l¬]M �
��Ik��K�4�?���?�I>��y�'���F�*�L ��)�-,>��
�d����O>���I@�$�����K��0q��Q@����%�4��ulZџ8&�먟��O����O�0)����Kp�)X.B&{9yǬB��9�	YM���L<�'�?�O>i�E�s"��	��ѫX����bs��'�BW����П�I]ybE��M�$H2֦Y��T�Pw(�<K�>1�� "���OT��!��<�;f�2%�C�/4�����M�P��8nZ�$�'W�'��\����/�����%P�1j\�QA�)?����؜�M�(O��$�<���?1�~�$��
c���c�-K�Hv�؂{IZ}��V���I����I]y���!ꧾ?��#%Yg"����b�����CK�]}�6�'m�Iޟ�����\�хg�ĕ'���1ƕ-Pu�A�T�Q�hR�Y7aӄ��O��m!��X�Z?1�Iڟ���Wy�)�L	:Ĕ��$��$z�O����O"��άw`�IYy�؟T�ӡDțm��q�j]�F|�Ʒi;�	��h���4�?���?��'	�i�]؇H�*������Q�8�5Lp����Ov��B8O�	��y"�i��|' �t�Ӧ^����E@f��Ac1�6��O����O@�)�]}�U�;Q�B	�� ��'�����G��Mc����<�H>1����'oL\#�Kюwq���Ƌ2!R���b�<�$�O��DT)=��\�'q����|��e(�kS=mLl�� ��sO,XlZ��d�'�$�����O��d�O�e���K�B����F ��f�`�æq�ɡP�
@�O���?(O���Ɗ
wjF�<\����X�<p{�Y���f�Ė'�b�'Y�O�f�;Ajԙo���.E�Tƨ�����*\@����O�ʓ�?9���?�FJ߄�bX� ℗�| ��f~�]��?���?!���?�(OT���D�|"t,�8"O�x�r�'�*H�F����	�'IbP��IП �I�Nƈ�	�qFE�!���'J4�b �-��1�O����O0���<�f��2R�S��@�1��
�yनܷ3/F��2ŉ�M�����D�OF���Ox��W:OB���Y`,,e$E�G��1�J2��h�:���O�ʓYmH(A�V?��	����5�����'˾iΈ�HQfF�Z�ڮO����Oh�X0)��D�|Z�����l�74��=C�V�caH�s��J��M�.Oȸ�QbB�������8�	�?�s�O��7���@D��A��L�ui���'RI
<�yҞ|��� ^� ���i�r��_�V����7-�O����O��i�}U����J���ӄ��:� ℎ��MSсD�<�I>q��4�'Nn� R��s N2n=��Y8i��i�iNB�'T"��1U����d�O��	&lz����ǵ"�E�t6�-��F�W&�?�����p��}���ᑫ�
	I2���ao�ҟ�j`�[��ē�?�������/�T�pc(OL�qrƊ�}}"o��yrX�(�	�%?��V*Ɣ|8���8&窰�W@όl�`�BH<I��?�M>A���?i���$����	ĳ.>Ȣ%ԫ)�V�H����$�O����O(�=޹�u=��$h FO�e�D� ��K���xb�'
�'r�'��`��'	���R�U?6�z��¨+T.QP�#�>���?�����Xȸ&>�r%/�?�PiCM���֢���M������?��'x�j�{RB�.:�P��q^�F"��VF���M��?.OviY3F�]��ٟ���*:�:�����c���@�L�c�̛I<���?Q���?	M>��OER�0(�s+V�!�%,Ġ��4��d��/Hh%mz�Os2�OL����2!�][�*Xۀ̎1�Fdo�����	4$��	I�	Eܧo�����/^�{K��Rԋ�?�o�n���pٴ�?)���?A��j-�O��J�%�	�8q�)WnX�3R ����"@��$� ����3'�ё��'@,,T�D�0F�L�3�i��'�B��\� O<���O>�	$� Ab6 �2M$��)֭��6M7��G6aF��%>!��ڟL�I.H�z��0-�����S�{���Rڴ�?��d� D[�O��$3���°*�Né4ʽ�]�m�:���R��s$��h�'���'��O`�'C�@�޴�O�G���p��|�rc����v�џ��ɸ4,R����oA��V��)�,��1�����'^"�'��V�������4���N�C��1��DX���d�OJ� �D�OH��9|���ʍcų�%��tmb����])N�LH�'?��'�rR�D��M��ħG�h��0e�1KS,]� f�i[W���	�h��TF
�o��X50Q��I�f߉0|��%��u|���'kV���"��'�?a�'8Q�\25)��@1��:�Ė�l��!&���	ʟ�ASg~�&����
�8Eے�>Qv� �̀�`0mZgyr�� 0� 6�S���'/�de ?���R `������"��,��IΦY�	�����"Z����OIX\h�OJy�����m{�`��4P�JM��i��'�O/�O2�$B�|c�-,L�H9�̲m��dlZ+���?���$�'�P3��01hr��Ɨ'uV�`� S�'i2�'�l%h`g �4�8�'��=8��:px�hA��<���ߴ��'���f��O.���oml�.�tdH��c]"yt\o���J`����|���A����`hY��\#6�X/b4�'rY� ��ȟ���ey2@S�H����b�ԗuX����X�lk:`��#-���O���Oʓ�?Y�U�%����8S�`��e�V��t3 �[d��?����?9-O�p��]�|:� ˟dp����ř<<l�M�U��A�'�b]�D�	����	.Uc�����b��8���g�63� ��'���'�Q��R%���)�O��Z���)>�6Tb�M�t�Q;1h�Ц��	Byr�'z��'H��'�哱SrR�	�˜9��	3r���c;�| �4�?9����5�:��O���'E�T&�/S����#C�	"ՅA
zwl��?��?Q ��<�+Oj���?q�p�C{ݬ	�N3<�
$+z��ʓ#;
�f�i���'�r�O:��Ӻ��� ux1����>2�{�ئ�I{tw������"��Gv�� �,m\��a��H��6�4�f�lڟ����Ӳ����<q�$����f��:I�t���ȡP�O��y�'�F���?y�	� ]�����Ɏ�5ڲ�3�'E�'ӛ��'?��'v���r�>�)O.�����H0#��{���6��$�8r��x�v�$�O���˴P�?���ҟ����d�B ��-��O��	�&&�Y�|�ߴ�?d�5=���Ny2�'i�Ο�����8׆Ӽ1��	1�$d���: �����Ot���OJ��t���o�S p��������af�U��	gyr�'��I矐��՟\�E��
?���٨_-|`���Q*)Γ��d�O����O����OdȪ7i�OV��@�˄��
W�Ўn�f�xR��Φa�	�����H�I����'����۴t�� �̱~Īer���UF��'[��';"R����X�ħl�����=xԥp3�Ť%,"-A�iR2�'o�OIy���
)FpI�.J h��tBX�z��6�'e�'�B(U+R��'"�'�����`).T�Ǣ Vp�X2�"D|$O��D�<��NA��u׺q����Ea��Z�$g�� L��v�'�Bl��"�'���'��D�'�Zc;R��ǲ�d0�4�B?p��Sܴ�?Q.O|��)�)�

�a{Ŭ��|���o�*-�6�Ȩl �7��O����O��	s�i>���A��z{�=��͝Bc䰫r؛�Mۧ�'��'���y��'����$�:L�F���̥UH���1�o����<��	���d�<����~�a�i��W�^ Zb�m�9B"#<ɰ��T�'�B�'}��ⷡ�46-������P���o�4�DQ خ��>Y�����sB5_q���c@�,�N�1��W}"���'"B�'mbZ�hr
� �u���?�� �[�iǼ d���O��D#�D�O��Y�31 EC��5�je����s|f�`���O���O*�@0����2���bg��7\R�A�ɨC�f%��x��'��'n��'ۘy��O�m;Ԣ+�<�r%�K3&��Q��Y�\���T�I�����|�H��Iӟ@�ɠ�͉5G�%K	6dc3�C�Q�q��4�?1L>�������$6�'u(�c���q��qy¯Ly�j-�ߴ�?y�����,��&>��	�?�c�mߤ�%b,�6/}�aW$%�M��2b�5��.��i)�ȸ�i�3Ċ����܏pI�1ٴ�?���j������?���?)�����;�l�!|H\mEa=7ڞ$��i��_�D*�&�S��J��\A��b�� ���*l7�<8��pm���Iʟ����ē�?!�ԩi��ƍ"���lɃ���"	�O>�I�4ϸQqs�E�%{�	c�k��A��8�ݴ�?����?�����O�������6��l�����\�dT xA�7�ɲ�b���I������>�Ą�v��g�Yx��̍�zL��4�?yD�"wl�O���?���&�(�A΋	�Ε�K�k��hvS����<�I�����X�']�ՍW4�F��t�����x��	]%~c���M���� ��0W\�pa*�zpd���k8ҩY��=�I�"�"�	r��i�����d�UP����A�.��0���Ӎ)�(�S%� Q�x,���ۖk�C�3fM�%Ǥ愉�B��#$��$(�	����ؐ˯68��-ƐX��x����rP(��L��,E�҈[�HHҮ�H��+pJQ�%� 1�V̍����i7�A�8���9Q�g���	Q��|�\8�'*H�?�Y%�8�dL��v��t��oE\Y-
����&`Jh�S���
hq���Za�-KQ
����R�[\��CR��'-�i[##�="�I��T�*B�vj*�̉��C�p�4lA��?K��[�>Yp�M�5��´��!&�`���4 k��m���<d�ҝb��J
%NL���Q8��#�$�OD�}���M���cb��xTK�,2Ĭp��g��S���a��B�@�0*K����I��HO���@;8A�x��j�;,�Sg.}��'f���@�d���'A��'��w,����*�%�g�� S� �+��&Htp�Cd�O�����ߥ21��'Z���#+ �!�,8k
ޱ�N�;SG��� Q�+�O@�j�	Y�����RD���
�a߀��CC�Uz������dF/��O�ўpp�"!�h1a..,ތ��%D�T���W.��L�	�}�m	0�!?a��)*Or�Q��ٖ	�:�p��1��x藯�9!!��Z��O0��Oz��������?��O�ZT������ �Ĉ�he�؉��~��B�ɜp"N���Hۦ0r�M�(`2$C��¹(�,�&��8�Xj4j؞����-ê�&��(r�X+��)�`���Op�=�"݁ ;�a`�,ٞ6�̚�Z=�yb�^���Ek�aKZ=���"J�*Θ'�j��������lZꟌ��t��p4�-D�<�2 j�2Q���<y������	�|J�e����&�|���U<,8���=9E^tC��#O�Mѣ��.1����2hT����k��xB@F��?�I>Ae���uc!��V^Ę �Ν4�!��d�������z	�h0�=\�!����m�CG�<9���hD�3����B.扟{�ع��4�?1���i�59Qr�5"#&DFIܯy���C��F8^�2�'�JA��'(1O�3?���	�{��L�⥉�/+D�s��Qg�$�;��?eó望Hz ���KpM1�	-}R5�?�y��$�-Z���з'�ft|��Dg���y2CÊL��k�\?a2IX�] �0<Q��	kw�Hæj��<��Q��YO��ڴ�?q���?��(B/"Q }���?��y�;E�&)�g�bE��C�/.B��l1�	�g���U�|e��ò�AzDs�cѨ�qO,���'M����2���3q�ž' (P�$ſ'��L>�7�B?�N���Q�`Q��@�)�~�<��f��^6�e8AȪ/(�A���x~��=�S�O(.Ѱg˃�^�ŁTi�FJ���l�=V�0���'���'���s���I����'B������ۇR�jy�u�;�h��na<�Rm�X$"X�q���F�����A�A����[ "ljkE�6?c"+�
�$9_.>��!�O�8f�\��ֱn�6 d�	s�)D�\��mߗb��I�v���f��('��9��'L���T�l��D�O�l�P쒊xR��4GڏAF` ��O�	�2s��$�O��S(��;��q�����G��ʕ���?��x2gr�d��Q#`)��l�U��UHvA��p<���B�`&�� xE�я�]E���oRZ(p�s�"Op��6��s�hP[���$E�4��O�nZ��q��S0�Urd�&%^^c��*2���Ms��?�˟��z��'ʬm���f���)&hO<J�	�'��kW�T���T>��H���#/l�P+�j>(�)�OV���)�ӈ�<�;��A�P�(���F�.��'��Q��ۘ��O>��2ˇ4K��e�t�E=�X��'r�eq`��6{���\75�u�Ó$葞�F�E/��X ��P&̙��C�)�M���?���o�D Ed���?y��?y�����a�@�����`���I��'V�9�ϓX-��!ܾІ�E��<5Z��=�PNYGx�Q�-��L�%��M*Ya�FHQR̓]q�)�3�d��T��h�T1Q�r]�4��;�!��U%_d4��r��X����&ɍi~�ɢ�HO>��4	�/g	��0��W$Ѣ���h�
�B�o�̟8�I� ̓�u��'��<�.�K�K"M��xs mUYR�X'fɯ[�!��9{&@9�M��b�ܳ�@s^%ON)�MOy�blTҎm�
f�п���'�xa�&J��V)���Yz!C	�''��R-�,@��cA�2%d��{�y�H9�	�~�~$Zڴ�?��v��b�&{�RLh�J�;�b8���y���?������=�?9O>�voǁI�����N?;�6���	F8��A�,�I������^�bz��zBB���d�2x���|H�Ġ�@H�r�`Q��Y��y%w�q�!�(}8�5AB!F4�x2bj�@���\$C+�<�$;r�`q�dŤev�n�����Y�Tj�%�?9P��( ��c&�9%l0 G���?�>&�)r������p	&e�	\.8�*&}�h2�7}�X+�O�L�����A1���=!T�l��>�"DSΟd�<�j7c�=G��#�ʓ�dnY��aW^�<�.�"����8 �qWDR�������iO��``�)L@�ʲ씂N���'���'��qѢ��'���'�r��y�G:cHH�WM]�nލ���6-޲$�c�o�}����qC����|���>i$�|��B�=7a�S�[%�rm���=b��p��-�d�P��L>��`D	�D�J�F�@X~����E��?!�O����|����@�N�||ʡ�Bi}���юd!��B0^	$)���=qplL9��ST����HO��sy�R�L|���㇌Aўa1"W�m�|q��GO�;��'mr>O��ݟ�I�|�7�#j�F���Y�e9��9  ńY������I��['/��q�*=p͎�}�"���Wf<ag/�)}zp�5�Fs��`
�A~�\�	t����qj�by�d��4*�0� D�`��2=,�AQ�R!ODX�sѪ(扞��'~�j�|�����OR)�0�D"o����t�=�]� ��Oj�I4�x���O瓳X�`��7�d�z�a��L<� ��啟��x�-����'Xfe����cHy6�F7{�4��Ǔ4��%�	J�I�}�� ��/�����i���62S�C䉽.���A���"Ĭ��#Z�DL�C�I�M{����@N~ seĨ>��3^m�%[�p#�iD�'K�ә�����}�,G��:^�� �d��.E����O���f��Ob��g~�Mʕ'~֐:���;9��K�����@J#<����UK&���E/1���[�CO�DÊ^f2���� |F��Y���)��/��KX!�� 4�򕆖�m�����-W9DaxR)�S����QC���Gв|�0!5�i�B�'��Ĺ���A�'���'���w�c0!/͠4�sOM����󤅊/z�y� �;ovR$2��͐:�� rG̴��'/N���3�l�I�W:
����
O���J�y�I
�?�}&�\�w��iq��z�j�tI�X��4D���$�q��@va�[��-�� ?y��)§*� �`���p����23�ak������?���y¾�6���O��SB,ȍ��ZZ[Ѝ��XYP�<020��a#�R?q
�:EL�z�l��F��6��C��> q���6 �F�Q&�@%�ū���O���� p�����z�xq�6�^��J��"O��bω�	>j����(w�p� ��UW�U�4�iŽi�R�'�)*K7}�������J�
���'��$�$���'=��,K�R�|���AK��тY#\����fZ��p<qt�IR����!��m��c�`	`�DY��\��	�g��d!���)�ب0j�?23��qpF�r�!��\��͚Bl�xzdk#ţW!�$��Q#��C2�SQ�G�B`g�%扴rQ�h
۴�?!�����L8���K7^�h��7vl�	]��b�'K�� �'�1O�3?!�ώ����'�A�YŘr��t��?Yc�ߥi�A��ߒX�(����3}�N׿�?!�y���g�$IV�"6�C2u�|��3g�4�y��ϼs�n\QQ$&p��Pe���0<�鉡`�>0��"1��2'Æ,G"�ڴ�?Y��?�-� CF|0��?����y�;2�����6E<��"E�H*LԘ�y2)E��<Q��8��afl	�HӸ���$O`�J�Ԅ��qD$`�ѫ�� �[bA�� �4�<a"A�џ�>�O6=��۬Y�qa�J]b=��"O���֎��c܌|H&@�5�Ը2�������5`/���7o[;zy����iT~h�9��ԉ|����۟����<�[w�R�'L�	�4e�ZIɰ�R�]z�#v)ךZ��J�O����ؑ]P`Q�NܴU 6�[�G�4!�Dؐ]>@����D<%�,y�.�*�L�à�'/��%U&BB!��n�'�<=ؠG���y"�2��p���!�F� d���'|�b��P*���M[���?!�`�)�+��D�6`��
h�9�?a�'ϢU2���?��OUX�
����3_Ҵ`�2&�V0Jt��g�>l��	�g�P� 	a��iִ��t �\��3�;O�I�2�'��'��	[ҧO58�NX���L�z܆|!�'����3JL'5�8��ڃ(p����'7-ȓ	�QcLB+~��X`	Mx1O����K�)������O���Y�k86��� A�e �0B�#)"���?�vĂ�?y�y*��ɵS&���@KE��jq	�|y�'�������S�b
0�G�TO�;H׷)��'�����o�S��ᰄ�F���
Y��AUq7���d�<l�ċ� �-i7��?l�%��'�HO�W�m����nL;	D�����Ц���ҟL�Iw��)R��ϟX���������B`���/�=
P�ن=�n��E�l�ݶ9�牀?b(�v�9��ݐ��!]�x�ԒAM<<O��{4B��crm���d1��.�I�����|R�� ��hx'CU{T,�$��?�y�a�M����	��P�F%k4�ݵ����}���Xa���_<�����b�4e�׊H3�ѐ���OF���O���캣���?��O7�}a��	�0�R�3'"��k����x�����b�@���Lit�7J��	x
�'���zgI�yl�h �ڏ[�r$�aݢ�?��3�LL[�`�]��H�g$M��m��P��a� ��ZHB���Ϝ�Ѥ��<q���I2n�ȟ����2yF=
�i@|�@���μGRY���<���������|2Q�M���'�S6E� I��9�mC�AH��$@-O����$^.g܀�#�
���I��e.�xr�̎�?�N>�үN_,�tSq��9.��)�A��l�<!%�@�c���6A�(�s��c<�ֺiJ��1n@B�r�o����юy���7-�O��$%��HП�ڂ]H������5ipxf%���	�}����IG�S��Oި1Q�U�1�~(�1��Fȋ��Q��ɔ'��?ŻDl��=��;�ET#��{��*}����?�y��d��6A��� �4>�����y�l]'eHN1q��[�;�L ʧI��0<���I �n�[d�X�Xް���ݭI�:�4�?I���?��ߓ@�,�:���?a���y��oa���u�	����̜�<�����y�(����<鳦��|������ϘO�TbծEFܓ,!�!��	�����T�3S� �S�	��<��	ǟ�>�OT��GoR:#SlRc�94�*�(e"O� rxSb0W�$�A]�s� L�ѓ�T����Ӥ)=�m��+��sW�J�4�Tz�^�����I��h�I�<]w�2�'��	ٛMFT��֤_�>aD��gϟ�p�8�H!O���fP�cN.��M�7u� a
P�!��P�c���CE�ѲzV�m(6�ІwK�H�7�'����H�:/X�'G<�R=�5\��yb$,�n�0�����,�1�K��'n`c��+�e��M����?�@D�.Z.��h�SQ�\iسa���?!��J��p��?əOh.t�������0�B}�♒wvD�#�����W&yXRH=�D�8����];g�xR�ÒOv�x��$�?Q���?���n��}x�`�.Fk@�G%�6L�.O��<�)�',=�,�Y��i�PgZ$���S�E��.�#q��z�H�	�y�Y�`TDA��M����?A-���Ygf�O�)!A'"�@�6�� |�����Or�/V�P��8�|�'	Ȅ�V��ň�L�ʞ��M�J�"5�S��=�c#E�f>"0�!N?y�P�OrT
 �'�1O񟰵�a�<.k�|� N�LM��R"O8��eƟ����9����?�����'�#=��Ԥ\�x�Pf#	E����p�e�<Q�
Ͽ&�j��hS��A�JH[�<IE�Y7]'�<�#ꕄ{���'��@�<1��vA��8�>e�D���DJy�<����� ,�����(F�4Ɣu�<� [�q쎝�0ǚ'��y�q�<)��عkp���hYi�N��v
�D�<Q�LY�< ,9#��#D�-<�TB�ɷL�^=��%�%)-��FIZ�Xz6B䉁~x�j7%?G�$ W�ԙ_�FB�Q�^�R#�w۴Y��a��Q�
B�'Qz� ��"p�ppɲfVOgB�	���ɱP�6�A��^"��C�	D6�[q��^�f�G$���C䉿�[��I�*��x2c�&m�C�Ɋ>r���0_��c�̜o��C�I�Y3h���n�,Z/�	*�I�H�C�ɝf����R)θ|VZti���p2dC�ɱ_hk%b��r(�2��{�8C�	,$�Έ�@�)r|\����1�jB䉵v��dѕDE	0u,9hua�y:B�M1d<i���9E�����Do@�B䉍7�Pi&�;B�ۤ��l!�B�I�TS VXMI�q.Hd�vB�	C88�@#��v�	�#��1t(8B�	�-�� �Ӧ��\��S1c�:"B䉽:pR���U]�(��A�1��B��4���'�]�~`�pBiϋ-^C�4�D���6!��$���7y!�ȳ'�a���}I:�`�@4i\��^��x�ؕ�ܗS�%�q�R0�y�\� �H8SiD����`!��yB�܇dq@��U̙��E��Ȁ�y�D?I0 1n�&H���Y����y�Ѥ ��5� 圳/�ډP�����ybcS�줬�ӫ�7TA�²K��y��i.�'�<)Fx�F��y�l��H~b�Q��|�Dl��@B��y�7D��	A�S5|\�qA��0�y�g�3=�4c�O#z���1�H˶�y�m.O �jamW�"�J|l�y�
M� �|��¯�'��l@�P;�y�kE&(R��V
jqzҡ��y�ʖ��e��A=[S4���L��y���/L�d8��3VD������y2��5s9�P�E(FTp���9�y
� �9�C�*��Zg�,w��y#�"Ox*��0`*��ꢀڧZ��( �"O�8�'L�Qp�0x �ʊ_�b�Y1"OvEa�n��i������N�9g��1R"O��q�ħc����o��za�%"O։��}
h4SnR=`gR�a"O��*��rK��� ��J�kK��"O��a*R���Ap� �L`�z�"O��(���]�t���O, O<)��"O5�S��)�P�2&IȞ��q�"Ol@kU��(Am�F�ʍcr	�%"O�x@g�� �A6�Wh�*� T"O �Y�
F2��4'˔@*y���'D�GIʭ_r�� �q~�qb�!3D��j�Ŏ�`�dX�+F
b&xI�1M%D�l9��1\���c����l8v9�-7D��`�mR�\?<�,��^��5�4D��)�� �<E�xᤌ���N�C&1D�\2ri�3?b���ηzb�d�e0D�L��C�:���u�J)Mr
m�r�:�OM����?5ԭ�c��O�� #�8Dw�@�D�hh<1%�C��,���*�2ՔA��Lm�'�\i���/<`��~�boU����#2ᕒ:��t��	�c�<��MW1Z���b�ؔV��j�J�۟4�EhQ�)��m��>E�TLM�c����qo�3H���J��O�!�&pU& ��B[��\�QI6���	ieJ,3�F&@ay"ɪo]9"+�crT{��tڀ��V�<§,l���$���'��4�iHB��ɺ=
�'���he�@��Lt��ўm�L̓RnHQ�%�1�u��O���&ΐ}�Y�U�'��Jߓ\ͮYb�L�>I�D��/g�a(���*f*eR$%�<��f�������8�7�۬����cdK:���!��dQ�<L�E��HϴBx�J��H�^(������$�Ǌd������k���T�'K�ɡ'-�H���Qj�	&P�50�~�1O�Z�OR��p�Y\%�b�IB�a�>Ȣq��2f��T���K,�졄�����u��KW�r��B�A4�(!�\Y��pMA
';*5@��2uJZ����9/���>�� a�3s�Yp1-QR`��K�!\OLl��<�剫U��pooK�,[��� 8o&�YCg171F��hѢu�n��n"�Ӓ/�4�&U�5CS$J���i!B�{�dL�=��!ԿA:6�E��N̈́JjFi�kN�U;,a[[a C��|�Fh�gV�5��`X%�6PD�Ї�	�>L�hH(� ~�<�s1�� g�q�[?1O��{�O�R �7� /7���!� �z1"��JRв��ƚz���e�m��i�U4Bt���Q8|�8Z��-AY[�#U�3���ɝ�U J�B���5��U�2�H
�\��RT�c�;/h�5��{ ��ʰ�Cr���������P��V����ְ;U���΢ʈt�g��?���U)t�^�[PH�?�����кCb/}B��4�z����t8y e��9��'��q�7�	O �3��;l�򴙇��z|�0��`@]�E��-_�9�j�����X����IAJ]ax"�#�T�5![�P z���N�qb�|��Xr^�3�BU ������' Α�'�+c��|��gl�4^��$ �ak�}��o��t��$1\OU1C��2"�P�Vnʇtp8�`�@@5s��a6�/e�}J�cQX$��)^��S���:u�=��T1JY(�#���2�Ґ�9p��IV��!w��c�P5Q&}e����>271O��� ��xr DQ�q�S����7-�!u�e�W鋰/	0Qa���J����56)��3%Ձ,*�awK�CG6���FV�d= ���;67��r�l��dTH����䖁c�hc�x�ׅ��f����)�h'�ɢ## ���9�̩�!�]��l�'dй�f��kZ��J�*�9m]���A�;P��I�Q��I��I�0$�2�d�obT59�h�:!+FDG
	SϦ��"NE�C���j4�|Z�%xmRpbgoG�C�,5� ߁T>�H�'�����9b$�3S�˙w�8|�c��01Y"N��?y��5|��(�	���T����q�?�*����]��@�� �yl9�O*��%k�."]�\8!��A���h���-`6� �MߧW��p�ϭvY���޴̪ɻtJ"�?����c�YDu*9��(ԕ[ن�	?{Nj����-!��pD��?Zz�B�)=:x���N�Vt�)���
�? �������UxH(0J��״
�̌����3<��ɏ)���[�E''�ʰh%�P�̧U�P0�}>� L�C�V�R��A�E�`���jP"O~���̎$�zRo��-pk�m���JǛ�guf�؆���n��b�?�	����0��+c�Λ�f���H2L�!��3p�l�k�G2Ҝ�ƯI�$�zU�.�]06!;�+ݙ*|��K6�O&��1	��Obd�'�?Ţai ��?��P��'��(*[#I\ �k�`��� ���WMb����e~ ���o�%�~2M�*�Ї�IѼ��$"z�(��\���'���U�F9Jd�&*����V8���*j>)2�o�z�G��)x�8g�ͻ�y�ř�6�ƀ�va�+%Z��Qj� Jڜ�h'b�,����p�b�VY����w�!�M��Nm����I�,e�
�:�'�=�"�D�]n����Y(�l���3h�N�Y��n��{򄂄7T��bg��TB�C�Ź�0=�7M�-j!�RTg���o�~A���$�:���R/k_�C�*?�X��#�8=�@�`�4\fb�@�h��f��G��>ki���m��r���2�$0�0B�Ɇ;�d�s)�2H�*}���)J:�l�'DV�ēt�G��O�Ђ��Y`HBv�I���4"OhШ�M�Q��a�$]�E��H���:��5��'/�M��Hڶ	�L��y���דC���pI<���Jج��f��o�%dH!��$oT� "�F���43ƀ==4!�]�V������ j��pO�f!��ՈUFR�Z�I#�̉b��Q&~�!�˰kV�ȡj'I�&�x�#س5�!򄋥R���pc��!� %z��Q�a�!�d��VdA�ƤD�[���c�A !�!�5V��4{�ՎF�
�P�S+&p!�$O���Ի$�;�������!�@$8pp�;pl�cb�џf�!�F���=��G�ye�9��QX�!�dţL2����>X�t��ֳv�!��4�t��B4`���צ�7q!�D�?Q��R�Ѐo�L@�FSw�!򄃓:�d1FE��������9|�!�X���0�G�+����ˀ�@�!����Xh�G�BȞ�2��O!�D�7L\�x��*_+���h�+Y?D!�d���0	���Q���x�+]�~�!��#"�*�ছw���ۂ�[��!�8�I��̺,Ąx��� �{2!�$�PR<��e�G�z$q0*+*!򄃔�������z�ڥHN8�!�d�0h_�,e��̨!gm�%Jm!�D�	$��y2a"t���͈�PQ��{�E����*�5��s�8�+"�T3F����e"O�)���%�
Aٓ���E�*���8}�W���O,A���B���ˮ%�fuH��ݮ
A
xz��ފ)H��}Bu���ظ�8�I8q�4�[��'@X<ibGװ/R�s�o��Z�dĊ��đ"~d-H>ɉ���S�H:r�̓!`TZ��X*>�@��=Yi���Dmt$�����'���g~��I /�0���.O}}rc�22b��'�8�&�Щ�.i����[y�L��4OsNa�g��<ɰV�u3ʝ�F�0r���B%c�<tI�|�`"��!{x�+�I�}mp�r������N�pe�[� �.IH�#�[���"O��RE����U����C΀����/aX����|r�����xn0��5b��4���03	"D�H)�m�;{q�!���d�J�3 ~���' $b��dģ`�8���bX�b�
@�a�!�䀣0�� ��S>S&� ��V=3�!�\0@$t�Cu��{q$���]-!�ވB��Q��ʴb^z)Vo·�!�]2[�QɡH���l쨃��,`�!�U�
ib�����@���R��"!�� b]8��ͦ>�0��ML�HŃr"O�QbtKԫC����nS�n�@kS"O��Zϋ`�I�U��
0}Ba�"O�8֦�)<�ȱթ�2��<��"O��jb�*p��``�i4rh�+ "O�EB�,3�(8�&�P0V]0�)R"O Q�aDC�,�#��;V�VY��"O�d�`O�^Eܜ�����p��r"O,�@e+N-t�:-��Q,S���f"OYH��7TM(���m��U����"O��j%"$+ɞ �w�I#8��U�C*O|!ʠe]�4d�Q.��>�|��
�'뼶NF3H��l�%F�aq��a
�'�f8he,��OdV�%���&�	�
�'?rL�r�4o�<H�)���8 C�'k�U�tAI�`�ʭ��#_���'�>4�rb��;��|�ר�0a�'4�	�cO�X2t��'E?�, (�'��pw��q�J���BH`�'Ov��(K/i�i:e䘿�<T��'�\�H�T`L	  �
#��@�'�R�Pd���hS��v��{{~���'�$3�ǂ1	H�0��m��Q�'R	�cϗ���S��a��H�
�'���!�E�H Q��KJ ��'p����Fb�9`B��x�D���'�N��n� /� t)`��#��Q�'�����'u�UyT��0@i
�' ��ufQ���Q0�b�6'���'E�e`��A�ud\�T+��T����'"��cRMS�8��_p�u���y҆R�[�^`s�.�r`�%JKL��y��+@�nU���i.nq��/@��y�$R&}�^���\�Z�ؔ�.�y׉Q�^�p��4R��D�y���H��H� 蓫g�Y����y2�W�\B���.�p���.Q&�y"��8׶l����s#ԥ�y�G,T����\�@�@R� 2�yÛ@^j�+�9���AA)�y�E
.����V �� y^=h�� �y���`�(�Yf���,�nT�ʃ%�yrk
r�
���[\��x�4��g�<��o���7�V'z�� ��r�<�@��=7�䔠�i&A��� ��\r�<Q�(N!o��"@��#Yxy���G�<PCO�O�\�9F$��paȀN�<YpK(��Xc�D34�S��	R�<A��V'.�2`��K�?`�N��flI�<)��-e��T���A�B�8��bF�<�@��S��	�G,q���a�F�<��)J��xBiے\*� �D�<9V$^�k$ҽ����M���v`ZD�<�@H�o���ʏM�F0y�o�}�<�0�зP����jÉ,
�	���^�<r�D�(}��F&{l�h�+^�<1w��L9>�Z�&O�R_�� �C_W�<�T	�|��I�P�������G�S�<alT�g����v��12���4��N�<��˄(Tz��zF��.�ݠ�a�c�<�BNI#a�V�q �� &v���X�<��/۲E��F�/#��3�d�}�<�D��z�@Y
�n�>����VF}�<�u㜱6��(��\�(](�� �A�<� ���!͈;ntK��]60.��07"O�Z�Ȗ�E�vyz�蟹s��q"O�1�v�&�$9���q,���"OJ�%@��.���`צ^�%����Q"O���Ε�9Q� 	v��r��;4�Ip����Mm�H5h
5kLЙ�*�!�Ĝ<?BV�"�O.p�Y���¢C	!�j��(��=Y�E{�鉹0�!�d�G�a����{nV$���˪vA!�D�~��J�㗯S^2h�(K�g,!�$Ϙ��5��S�&{�8�(�z !�܆X�Z�釂��7d0]��	�Q&!���-
�)9�	�*E��3&�%!�$�7Th6a@��$:�*feE24`!�F�)C yS'��l���C�->F!��RI.أs�ZRG�M�B�8T!��0r�r 9G�?b)&�IeO"�!�$_�-ްy�&ԒP��I)��ߣ �!�DVv��(u���Z`�R`��q�!�$�mkh��@�^2OxJ�z֌mq!���!Vv|-9 �A�%p��"!.$�!��J�� � ��I�@�tLh7�X<	�!�D�A8��X� N�s��	vh�?�!��߻W:,�Ճ�|`�@��
#j!�$̡E��u�!O>��d��8`!�$�p��1s� H�`㨎^_!�dʺ@��Չ�C֗I�h�p��JI!���7X:$����׌�T烄N%!�ʁ1$��ŕ2|�d�y�l�4&!�V0���H¬6�tqp��5w!��ϒ6ª���4C� y� �]�lm!�䏥iPR��k��ZD;��>e!��\�{���+��q�V0�dςgY�䓠>ma~r�qt���sM�.Nx��q�Y��0> �"}blD�9�F���X�B���:�N��y2%�p�X[�l!6C(�H�`:�O�C��O��볫�LOj���Ž>���'/��	>E;0�I(c�V=��%PT���>�b�|�mȢɦQ��*P�ȓ#����UeYva6����8�X��	$��?��"�#M𢽒�B��%�Q�ii��t�c E�N?���'Z���E��DD8�(�o�� >z���'�����SES��B�u�iÌ{�'��zc����X���G|�q{4a�b�i�"O�y�"ʋWd`� ��,Rڌ�C�n�'�"}�'ʰ�y��G/c���IWÇ��a	�'�6�с���K�d0��KЬq�
�'N:9�TE�9Ħպ!n��,��'IdѪ9�p<���+V�a�'�Hl���N�O���� U:A׸8��'�"�[v�S+M&M{2$B4?.� �'���X��Ѹ;Ni�QA�C��)��'@�᫑CE3�n���ڌ@���	�'>H�;��ɪu�\˃i=��h�	�'���b��.������/0h�1@	�'�p������^�
�5(ښY��'�Hy0�A�v�0Y�UA/z��ؙ
�'�A
�+̵�F�r%��!1X�k
�'��:��Xq�����)e3
�'�ڨ��LΒ+����X�Y1fP��'*���E�M�mt♂��#z�t��'�� ��%N.2>�����u?,�h�'<���7����rH%|2���'��	��L".Yf5��B�l��M���� F��5����V��O'� �"OV*E�;*�n���*g�����'#�$E�����Н[Ө�$��g!�D9|�e�Fm��+�d�hPMӨ1n!�M�mZ�*���;�B���Лe�!��y�h�եֻW�4��/�@!�䝧OGЁ 1��5e�@��@F�!��Eb<�l	�,,�0ϙ��!򤐳6��U@�5�"��=}�!�Ă7�FE�v ��?����k�:}!���hz�q���:}[�	��m!��,m�X��܊'e�iO�=e!��7��Z��n&p�+���5e!�F?;�dUX�� D'nE�-�!��D�F �Y1o�	D�(��*D��!�Cv̘�b��nd>��6
��!��~F]��I�`d*qr��1b!��*.����&[�uD��XE�ɗZ*!�d�9`ޤ�AO�;I?�0@F�1y!��ǈ4��XP@�>��Ԉ���=�!�D�O��Q��G�}��Q�!�V�qJ�����b*T!!Ȯ �!�D�.Y��e���[.��ұ�\�L�!�To�5;G$Q�H�0��*�{�!�Ǎ1g긁�[f����2$!�7dH �B��8.��֍�
�Py�B�p��@�m�t�P '�։�yr"K>� tRe
�)t �0�*��y��"Tք�2`�t�9�5���yҩ�#k��	��Ǳh����u�[��yb�V:���8%hB�5hH��샜�y",U�@d����u�Y+�L�y����H��G�~����yRЭil�@��	z{BU�`�ߧ�y�@ߢZ\��H���>2�py�����yr�S�&�l9w�7G�@S���yr�D�w�%	��=�VV�.1|���.�jĤ	�r=*�Q5�U2L��ȓJ�:��J�_|��sp��/H�&ՄȓL+��w���.�@���.e�,��T谨�,T�A�8B�h�3!���ȓ
��#�3<�l�br��:<�ȓ'��}2��݈zL&��O�in�D�ȓpi��kEP�x���&�Զ0�0\�ȓ!k���e"_�q�8Ë�0z�P��ȓV?�B�.J5_� �"t�4}C�U��Q �̩te��A��=b�a�
- H�ȓ|��aPK�Vg��	7�mת���;���� \�\U�I�΅�-[p��I<����h"�e����>�\�ȓ8~Q�ì0�����
�3=�2���9������68,a�,w0�����S ���9��I 7gӦNĄ��	a�'��E��C��&I�W��n�^���'����1@�����6(O�X�v�
�'9�t����&a�*Mt�H��BК����)S��u���ʝU}��ȓ+���萞M�|��%�Ix��P��Ѩl��ɛNy�`�C��T��]��F��{�bȪn�b���ϨyVń���-Y�)��iR.\�H�4�ȓD`-��].^���h4�5�☇�_���1��VU�F��?[�|��-�p�f^ e>�h�V,u�x��S�? ��B���?@m7���.OH�4"O���vHW�3�z�E/�046R��`"Ou2S� Z���Boөk,����"O�Q�F�'S��)Qm�m&Xq�"On�J �%W�1C��9Xt��"O����Ƙ�<��5z�a��N@���"O�x�(|�n�J�%HIM�"O� �a��8s�r #CCBE�'��lZB,V�!�Z@�#�Z� �zŃ�'l �� ���R!�E,^�J���
�'���	��ϒ0�&[�dǷ
'R)q
�'�fd�đ�UƼD�2�A� h�$�	�'���1`�2eٚ��V={K	�'ӎ4�E�@ȝ�@���v� �'٘���C��[�^�{@/%�r�[�'z���U`ڥ�
�'�Z�wp��'!�L�c@�.�p����j$�X
�'1���P.˓x���U��P���X	�'��k�F��c�V8��Em̤��'+\�а�M�7
h�:b���9Id,�
�'zh�R��4a��ĭ�2���
�'���Ye�Z(fnd=�D+��y����'@�˗d5o8�L��6�:�'��ir��/
ظ��L	e�B�"�'˰�"���R)�Hՠ*����'�
�<F 4�� cY�MJ:x	�'qt��g�Uq ���.|���	�'��AQ0���'��'�I�#�!�	�'�N��,G!�@��k,-o����'�D�0&^>f�Ա���Dl�A�'�*	�$ :LO
4S@�+�����'���a!��n�1���������'�ʰ��E��u�O�� �'�j����B� ٠�&-5
��D��'�����$�lq��":
!�'���ԏ��K9�����<-h�<P�'6l�R��>��6V17�\)a�'3����m�
w0Xi���/%�z���'i�͑t�
 �f4�C�#m���'2r�2�F�j�i���<n�Zi�'&�iX7H��T�#dE�<"�8�'΂��5I5nr�`c'�3:P���'zF)���޻{���S��4k���'R~�Vi��w�T$��`�:��J�'3<������;�`���B�d��'�,��@$J3ex���=B5�'����U/H9���B�a����'�l(��۔BoJ�x��#c���'vN���g_m0������.0=��3�'��<������P#�ַ!k�"�'��i��nO:`���`eN,�9�'J�)��ĺBE��ևծM݂�r�'v��"b�	>ML��u��L�f�p�'�v��&/O�&P���� PK2~��
�'�6�2�Ad �SCS<���'�r�腮�.8Z)��@��g�V�x�'�l���_�|f032��!dM��I�'qd�Y+[�S�l��B��
V�"��'jX=[�:w��|	��Y<UFV��	�'���v�A�N�3J�M�n3	�'���'Te
.` �o��{�nU�'ʲ5s���h1^�����\�3
�'�l�B#Ӵ<�<]X�kX�~#f��	�'�vLPSl�	Mު	�ʔ�qI�}���� ��ʢ ׂ�^a�7$ܶw�D���"O^ԁe`�*��,�1���w��P&"O�)aEĤ*�D9L\�`Ǣ�x�"O���$CP�gnbTy 놎g⚌�V"O~�AAa���Y*����sl`��"O�T0��2d�m�b(~d�$��"OHE�#�ޘj���S�o��IR�"O��v�ŌO�Z(�Mǭ?RL "OD嘦�H_.��b׫�82J2��s"O�ۣυ_JZ ��N���]�q"O
x0$	�)!ʮ�۔������q�"O��r�]��!���\�(�ִ�r"O�dQ��3b. �4%�z)�B"O|�ˤ&T�Ȩ�v�&�j!"O~���>kwB5��E�=%�ur�"O��C��*d6� �
(�m �"O��3���m���n6�#"O�Q�Ƞm���#�H7w����"O*�ҧGK�F�P�hF^�#H����"O:�S�,��? L��$ʉ4"FJ��t"OJU"LӼ�r����-k6�B2"O,�����T�^11��[4>!V�"Onh`Av]x<�AF͘c�� �"O���''��)J��$EǳlYD[ "O����+��w�($x���(�@<�u*O�5S�M"��!�ܝ5�,��'�2��v� �<g^��b�9k��Y�'`��y�S	����,�@(�'��`�W"�	4RH�1�+X�:��2�'t!����x�QV�Z�@a*�	�'��`�p���wB(�إ���@$��i�'^ӅBo�����Ƙ9��4��'��,Am�<�8�Q��[�@.�
�'�:�S�g�`�j�kq�� 2���'���b�I�/`�`���E�;dp�@�'Mxۢ�ım��Sa�G~�x�(	�'3dy���¬>���n��jvv���'�D��L�U���A'��d�tȳ	�'�1`�fW�N�Б�w-B�q����'�V�]�R����&H�A���@	�']�d��&]�Hx���׃
�GfdX�'�����d���(��GyVԘ�'d�\���/B�4Ӵ>�ji8�'��H��oT$�����?_��ч�\8�,
�c�;����5�����ȓ ��{Ԏ	�&�`����*��@�ȓ_l���gت3���� hަ(xD��h.M�A#'�X'�(v ������]�a#E
Ht�y3�&7h$��5�R1so�9�0�#$�_$I�	��0D�Ր�ѝ#c�Ļ�I�@` ��ȓ]~�I�ꛐ�L" Ћe8��s��CT��5u<��W뇄9G��ȓ�L�C�3b���*�a�>Z�4�ȓId���"˩gI�Z���:6�U�ȓ
	@}Q�%� ���r��:4T�l��<���g*D�ĥ)`���0fv�ȓ53�������d~�� ^[�<�AH����Y�hߩhQ�DӁ B�<	h�&\��U��]�s�����{�<1�Կ|
��"�*k�X�h��r�<$bW9cɜL �ѝEzL�C#Jo�<��MH5�4[��B0=4�В��j�<�$ŀ���$ �W#��x���h�<� ��0��ۑl1���i�up@�r"O��;w����}2�>�8��S"O�t��i���0�B� ܱ"OR�cw�JA�4���8�P�I�"O���aM�$�Q�aB�/����""O� @틦���#n-_�H黡"Od��(��P����-ɤ;I��$"OD����
`Ҿ��JD���|	�"O@� ��S�~4y��M���ɔ"Oڕ��/V���a%��"OP�AO�PPdY#��)g`�(�"O�yZ�I� ��`[��6hT��C"O<9�Q`�#�nu���='�i�"O���f��NЬ 3��Y�z�z�"@"OF�"���DśЉ�;��a�d"O`�X��]�$d:�I��#�d�x�"O"��Oؕ0T�10�͈�S��m��"O�|:r'��]� 1�'��~q���u"O�ݰ�� Z�6��6N	�`Y�Xr"OJPT	�6@���[�VK^s�"O��EBT��UZ#B�|&�$�"O�T��� 9�N���D�4)'"O�$�! �?8�\�y��@;Y'f!�C��F�O$|H)��>N��lx �����	�'���X7��A������Ǝ��	�'�"P� &W�8X�hI3 g�J	�'Z�ui��: �L���"~YD�ʓq�H��-S69�q!C�&}`ȼ��v�y� dW�Iњ@����(7\e�ȓz�hQ�g�`�J)�
0un�ȓc���A0���p�պEϮ=��͆�	2��wF��!��4��.>���ȓA�.��v�YT��A��z�ŌG�<�#�A&:�xIǞ�b��e�D�<�%��P�~�%���0�J��Ɵ��'aɧ��dJ��u
��@Ws����  �!�dȯi�x !-)`*E�c`D?V�!�d-������L�d�¬q6j��Q!�D�K/���,ͧD��`'�
l!!��*%BEY�C3Z�&m�� :!�G�.�&�w�э#&��:��Ͷ2!�d�E��%��P*M��b[�~ў�D�I��4��pr���<�#��k�'�a|B�ςs\dU��D�;w�h��(��y�ɟ?j�t 'f�k�t|rp�@�yB��|��|� �ʓRg�d0����y��R&�0@��Έ�?�1h�,�yD�G��<Z3@���:��ÄQ���=1�yR^]^ �
�nE�Z�`M ƦѼ��'�ў�Oi�ԑ�)�,�`qzE�[�T��a�r�)��È�[!ZM�s�Kd�,������0>)SÒ�^<1��D�vP�͌J�<�h�Ysj�z�5'<b��0*n�<��͋�����'|�����<���m��C�IT�)Np%8�ɋwh<Y�ڸ`���b4L@68)�F���y"�X�Pe�a�2��.3 ųꙄ�y*
	$�.�	!��Q֜A��Ƚ��'�az�JT={�
�ׇ�7���+�Δ�ybа�8����.��4x��˴�PyR���t��ĔJA"��%AR�<�ӊ\�>�(�G
�> =a��M�<�u�V��Px�p�I����`TGy�i>��<�掝�h�@���M5�LRp'�{�<� ^��r�Ap���R�7f�Q�]�8E{��)���}���Ϟa��L�c���!�# P�(�&�@�z����O!�ęw��;%d�5$k`�{��Ǻ?C!�d(��{A������N
H!��$ �x�sC�:�´�Vh�9!�UVo�����N����1�!�d�*J�:�c��זwu*L�c��2�!��N#� ��%��O����ue�N�!�DҐA��;%	��[R(3�Ꞿk�!�$�H�<�����;1�]`�&)�!��X�^Te��%�O<�M���ѕ!!��J�tt�Gτ~��|�qG	@!�$�g;�I[э�}P�}�U�1�!�8`蜥k�j̦]0(@!��f�!�D۠?3`�d��J,)�g��'Pt!�d�O�n��]��r�#�.�=`!��K�"��+ŬU�vCGd#T�
�';"�$�%�|�DYf�H�'���#%>�� �&M���x�'��걪������+ֿ9�����'
��!K>O�@��C�.#� ����xB��Qج�#Ѩ��Hql�0���y��
�ܼ(�N'QAV�Iu��yR�ߛKM���#���>���+�쇆�y2J�%~Un�@��A�^s�l�r�:��>��O(�s0�S6dD�a ��RE���""O$y��9;,qI��9=p��c�'�!��7lV�]zB����|��1��_u�Ii��(�0�c�))�`3u�M h�E��"O4��mA��lT��߯%:�a�"O�1���즙�en� c@���@"O�((��P9 ��@����q%"O|�Dɕ�F>�k���%{(�B7"O�%���-q�
���j�	h�}Q�"O��s�)^-cEv���α]�t��"Od ����(8t�Z�ϒA_R|�t"OP0#'-e%ZчLܢ[W��e"Oz��t��#3q��)S-E2�"OFa�7-�<U��4)��?8t,�V�	h>�1h��0;��1sD���� �d6�S�''��v�Iq�Ա��}�朇ȓw�X��R�ǐ5J<\���{��!��)@�)���oݰ򡅿A�.(�ȓp@@����T ���#e��A�ȓ}�2����h�*iK��Y�~_�ȇȓ1��d����7k�[�}�,X��7v$`u"��6W� ��'��_�<r�'���Á�T3�����Mp����'���0w�Hp��K��If���'�0��_�AH����ǗJm�܋�'�L���fA1��x��P� �Y��'��1s��;!��j��>���i�'H�-��ā<EP�X�Ïb�J�'�4���'�-jݸ�9� (x��4"�'ϪI"b�����4a���w��٫�'l�~�)�' 	:�%Ǩ�[tE5n� ԛ�'r��XeM�̸,�6������'EָP��R?N$���ku�l�Z�"O�]@�l��sͼU���
���rD"Oؼ����[~"�Q )L�g�Ne��"O�4��M��A��I��>5�!�"O^ �Q�]:5w�tqṽ�;�v8�S"O���&b]Q�V�j�A�M� sS�|��)�3� ��	C�C�L��%pF%��I���!"OF��ЧEI��1�~�>���"O�%�*����]ѵ�Р��D��"Om�ԏ�b�8�c�#� up\8�"Ofq2r䎌vN(<��`�<�"��B�'��:��uBD�#�L T;n��$�7�O��h�tC�f:Z�0b/Ɯņ�_V�U!$�Q������E�mL�d��w���h�B�������
�EbQ��C͜1�H��j�9g(��J�P"O��Y#
A:J̄��@�fi�W"O�y@D@�U�p�rA�&N�X�T�'B�'6+��S�v�X�ZW��3s�Nȱ��'$���tŁ��R',��e$�9z�!�DVO+pɋ�,�G؊�ycNY�F!�$/uD���G�"t���LIk�!�)V� ��&��!�z��jG�X�!�dĽ%�h��&��)S�vY�"H5,�!�O,D�u�`��2l��Ő� Q/:�џ4E�T�;j1�)�G��t�~�ʧe����?q�'	2e�"�A@�aK�gA�z��Y
�'=l(���`���Q����ֵ�	�'�@I5b�&JP&��d�q���Q�'�*��4�ݹ�~���f^�y���'�8\�1l�?W�4��I[
\!���'xz�Q�@_� �RC�� W�؉��'~Ř��^�ǳ�$kA/�^�<Q��V��H��G�	��jS��^�<a�gͨL��!����fT�02��W�<����!`:�%��M�61GRm�C�CW�<I'��|�8A�e'�5q3F��h�Q�<�U$@�L �ݩ�)ʳ/�	ۃNX�<�b �+N��ш�i��2�W�<��):N(��� B.t�܉�&��Ux��GxD'�P��Gɘ<P���*œ��yB�4h�%���D�K��|�S!5�y�b�Bg�PJc��C?�`aC�Z�y���#$��U�޹h�̡	��×�y��H�jF
�j�́�l��  d���y�i[��ꜱ��._�t�"J ��xB�9HP���z�||9��I{��t���ᧂ���r'p�йZc,D���GN�$:9%O�(V	�Ã�+D���p��:`6,�Q�T�� `g)D�Њ�g
a��������k<D�H:���=t�P���^1&��9D����L�u�:t`$�Ȳ\P�Q��K8|OLb���/��/�"�R)P=��H&K4|Ob�ф���G��$��ďoU���O2��k����եB�fwB�R�ˍ6X�
�JfH1D�𪶌^?5u���!k�
��c�/D���rC}��P�f/<����S�.D��а��o=�FjKh΢qKn-D�8�N1.�!���Y�l�(,D��
���Z�4���"x[Bz��)D��i���&�4,��M܏�� ��"D���C�$@�-�W!ږ?��� �,D�)`���Ɖf��po�!�=D���b�Y�F���R�&"Zd�1��(D��z0a��r�[��S�C.�sŦ&D��A1�{��5��E�&E�����"D�XOQ��tCf���H6�	�'�"D������Q��ͦe9Do�A���0=�t��1)>�i��Ԫ�]k�@�z�<� 6y�p�	).~U{�@-)��Y�"Ot}!e�Vj80��N��D�q�|��)[*X�`�dc�$I!FO�yL0B�	�4����V}�<�Վ�	�jC䉻5�	PRM�5V��������C�$9Č���s���T�53)dC�}-��d���`���6C�-�*��͉42�4�4CE�m�`C�	k�����ho�r�ñEH>��D&|��87��[5�5�T��8����ȓ>������r"�8+��GM��=��V]����3�t��pB�,'����&�>MsӬW.A���֥1�����r4��@��R��A�Hx���q��8��>�2��#��l��+6A��x�^�a5�γC3�`Gb�sbd�KE �}�P���*�DC�<1�PY�U�;|JH]�f.��7C�I#<�`�rȚ?�KA�F�*���"O"�ٲ�ײh��xCq��A[�!�"O*����*ɨh���\:Wl��"O�� ���mI�[5׀WF��x�"O�8���WL���K(=rDJ"O ]��˓�#�d����
�g1��J��'�ў"~�e�$2E^}�Ҁ�<�@�1A�P(�y"�O�K��PZwÓ9�����j\/�yB΀� $]��%�=^-Ԕ��)�y���wB&P�B��(�8Y�uƒ%�y�8h�h���P�W�QbE��y�W%QB	��(]I��!#��"�y�2���)�b7@�PX��L��yrL��L���ⱋ>iv��h�E�&�y�U$ܜ�yv�-��&�<��?ɘ'n�i��ዪc>�K7� Or,��'Z��x#l��B�>��n�~2}��'j2 B�d�-uh|*�a�!���'����D�F�m�hG����B�' ����OǪ�v#�<�"�B�'�T�g�Y�/����O� b]�'���(0n�x�Q"E��ma~�k���2�^$��h�#4�8�L�J�j��r"O�#����䩐j��y���S$"O�,C	�J�����E�����'"O��rv�V��p@'�s�l*4V��E{��T�U$+L��I�5h��,Ɛ E{�O���͙.
t;6��{�2��
�'��y-�$0��x`蘰}��	�'��!F�b�&��P��>nvRih�b�'���	�ƙ�X���WJJ���'!D���g�L�ZLa�%�J��I�'j��s��&%��es6�� >�|���hO?��D�:S �0��_�Bٞf��ȓ,p� CB�ɠ��,^.��ȓ@R̭X@DխG�`+�&�ktbmD{�Ot��)v.N&��V�W�u����'ء8��g�8�f�b�#cΐW�<QM��ai�,RW,L%���{�<��`L�i�R`;"gʎV���0t�<�S���B�c	1h�\9�#Fpx�4�'v �7I�0o�,�P�v,I!��k�<12���w�(�ӏU�F�D�
��o���ϓ�dH��~����Lզw�h��ȓCO����Ó:D=y�ʣ|'f,�ȓNr,�q��_��X ���
J�!��S�? �EVOX�0���b ��uv��R"O�X���0��D P��"]�5"O%��͛$#z}�S��9~��%"O�D�Ee�'`Pњ3(	�5u,<'"O��IGm��$�"�� �y	��2�"O��<mTY	1�x��
�"Ob9�D�*^^���c�0�eʂ"O�}���uu̐���C��S�"O�q���ۦF׸e�D��T6\�e�|��)�ME}� חd\��X@�I5�|C�ɔ$��)���:b�!+���p7�C䉟~T��W�.^����n2?��C�� dd��F�K.^d�P֮V��P��F�"�"W�
���(�s�ñs����	/��Y ,�n�x����T�ȓo�H�����N>�͙r�\�(L�i'�|����A�k@"ؚ�9��:��C�!E@|[c��b^h�{�ˋ�Q�x��d'�*�ԋ�*�X]g/�w����0�8H�sd�^�Pb� `�艆ȓ���sj��a����fOH!�ȓq��5���ƧyV�����2a�.���+f��h���R���/!��ȓg�2=�w \*����*8��t�ȓ#��H4 ؗ@֨qQcX�"��-�ȓ#�Ԑ�&iV�{�^�i�M�1q�؆����"JCv�Ε��c�V;^\�ȓ�	y�k��[ޤٹ���,�ȓl4R��GI��8{�E�-ED:��ȓ]m\�Y�J�B����F��ȓf���ԧ�H%�=)Q��M�2��ȓ=�40H�)�/�D!١挌Z�d1�ȓubX�-�!��Ȑ�TT�$م�#�mi�o.lhx�����m}�H�ȓM�^aG���3���xf`���&��ȓ\��bI9�t�b�č86䁇ȓkMܱ1bF٬.w� CJ:JM�e���v�yI�<Od��1�]�	�8��f�P�Hg%� 11��&˖�C�,��ȓR2j̑�l+b<đsHZ|�̆�<�z��#�()���`����1�ȓ<2�H��'�q��e��8p���!`"���(C ��� 8_H�r�)�$ã\ �LZ���L�ـk��yB�ޑm�� �cn��+��	�Њ ��yRfɣ:�*$��B�'V����-�y�C\?g(Pu2b��wȲ\��ϖ��?�'xJ�a��Ht`�!Kȍݴ�@�'����E�8P�E2��ˏ� Y��'}���A�E��`Q�(�:����'��M��I�2n?����[U^U�
�'i�:%��*�de�6(�3�E��'a��Ϗ�?t���vj� �2-��'��M���?^>\;Ueݵ��b�'M8�^!^�FU�'�z�f��'�|�`wEG-8�^�W��w02�B�'h�{��;	窭�d�l�ⴃ�'�.U��̌O�(��˘�4.�	
ϓ�O����N�bÔ��E%�>P����"O�H�5O�x��*4���VGHԃb�	R>yp���-0��f�1�<K��#D�Љ�c̚PM���c�@�p0|<��"D��Q���H�6��k�z6B���-D���D偡icb�� /)I�}���+��w���3� \��Sd�,�0��OW�|~"@��"O�����7��EH㨏�Pq�#�"O�	� J�����%�].Sa���'���C	(c��������B�;D��)��!*�d�q���t?��w*OX$���"Np�6�Y�\�q�`"O�0�� +���!�O�Ty��c�"O���V �o3u�7��Dy�Dr�*O(]A��9dj҂�	6���
�'��0"%�[=Νx�1;Y0�2�'���Y����k-8M��Mŷ<a���'�8�x�m�<��D�l�5�@\�ʓWT��@�x���Gƒ���]�ȓh�����&=�ru/�<t��ȓs���s��fh���>�i��QA�AY7.����E�â]�m=.Ԅ�/�kD(E�?��a��e�/��-��s�e`�ƞ��j���j�-i��ȓB��S"!	�,�����G�>?o~���09°�1t�6,���ضu�V��ȓ�v�*"�L�E�ZEɷ�]����ȓE��� �%��O&4��E$@0�����M�Ly�m	�	�
)�`��s̀��"4��2 [��t��1͍�b��ȓKĵb���qA��ѤkUF���W+��x�*
$ު��ݞVw�A��@�LQ�$�
8Cԍ�Y}���"O���J�V��	��
(2^�q@"O�󡭝+}>h�VN�>�H���"Op�!��N �@���,Y",��11�"O,e{�&�X#���JڵS�T�a1�'��Ih�r���#W�����8��C�	�"�����"tk>����K/��C�
7,�Y�R�-�
�Xf^�E�rC�I5l�(��J;�5��'^C�	5s���`�
[~eȂC˖PBC��.]��i���%}�H�	u�DMZ\B�8-*&�P�*�^�0��^^��=�'sZN�@
J9xeBL`��C6N����Qw(4���یGB���2NO��찆ȓs��0s-Y�8�� ��dG4N�ч�J�4��D\ ~8�g����-�ȓ$�밀�^p2��Ѓ���ȓNZڼ�@iܢ~�����]^�5��!뾍j']�-��{cS�*5��G�0�EB�(���ҶM�/7ՀT��Mk����/��;Kɹ$�� {��І�}=�����0Z�K�>����/C�$9s�^���Qᡄ�<UOf`��ph`�`�Ğa�yQ#�Y�� �'kB�X�d�$&���[�`H�j^���'�){�	�RBBa�nޅg���x�'+��B)ˤO�LТ���a+z	�'S:|  %á=�Z�A�W�V`�P�'�Fy�ӝ>��M� ���"O��B��b�:h"N�-�B�z "O`4q��q*�u  gƯ)�Y��"O�ca�L�g��0�֣J�.k�"O^���E8~��Cf �N�4�G"OR�ٱ/B�H<5zQg�8UJ�)�"Of�!�9<�|�:#�٘D�)؂"O��z����ٲ�A>�X��"O�mcl�{x�R��ع`�p*3"O�T�gղF�pm;�O�<�p��',!�� ���s�הq�Za)7�vT� C2"O �H�(/��%�F �|,3�"O��" 
d�K��O�b�����"O@`�q�%CsZ!6c��it�x!�"O
�����-<�QD�?XevtR�"O�M� c�!H6N��V
�7S:��T��D{��iý@���$$�0BH�ԃK�<W!���-���A�'6>?.����B�!�V4������$19L�|�!�D�	�8�v���+۲H ֪�+c�!��ܲ�jfF� s�@�����}!�΅* ��+Ti�â��@.x!��V�[��Q�pWk�%[!�Dׄ	�N}-���SN=&ۼa
�'�y��O�/
S�֬��	�'���G����@ҋ�Bl�
	�'O�\
4n�=0�iP�@�Uc�'���BÌ$�|T��(��0|`P��'ƺ8���;BP8�bT�#f:qP�'29�F�$[��:ٙf�B��
�'�ʤ�&#Շo@�� ZJ���
�'�L ���
��m��-NZ���9
�'����D.Ո(����� )��ib	�'na*4�3���s��kD��r�'Nذ�I�f�܁��KYOi��']\%2ҵj�*�{�)� �=��'5li��
�Z6����ޏA���q�'����Q$�,D2��'n�.��ݓ���/�z�!��@)P����1`�0�1�"O�A�%��<߼ ��@�W��$��"OX�9�݉Ϙ
я�7 �n��4"O��������z��`�"O8����6_<\�b�@پ���"O�,1`���*t�xt�C�`�!�"O0Y���=$��A�V#W�*��Ֆ|�P����K�
|2'MW�E�0sfJר84bʓ�0?) �5u��brj�3��8j�B	I�<�t���5��0�b�/9E䔰%�	L�<�*L�w�А��i��IX�V"\E�<�$N]�l��q��+O�
����^@�<���Q�d�:l˜}l숓&@�s��UyB�ONx`E؉W�Ȥ@��2hI�qsN>q
�'o(�0!�`*}��\�V/�I�'�a~bM�'�����A
-A楒En��hO"����\0���wo�� M�����$�!�䁔k��8[P��6)E(@���U6�!��0v�"���|>Z�� �{}Ȇ������/�fgإ�#�A+?
`I�ȓ<o@��b�u��@a��]#<:�t%���I�xV���iI�ZD� ��S>~B�ɯF�t0@D��7v�����N�g�>B䉼E�-A׍b�q���
��<B��e\`�s�˶a��Ҁb�7d�B�I�<7��Y�aX���Q�Z�C�	�X8��ӡC�\���6B��"��C�I_���%�B�de�[s�ԗZ�C�	OCL�B%W�(��R2M�,C��;@�X� ��i���[�-R�p��C�	�& `��指]Fe;Ŭ�[]hC�	W[�԰բ��+��k�B�)"�B䉀D�x`fϗ!�� ��=��C�q��I��Q-Pΰ����v\�B�	-[yx-�3��/>�e���ڤPoJB�	�a�,�M[♃U�Y�#$�Ox��� ��遊�
?���[�H"Τ�1��'�ў"~BC6,����O)��M���ͦ�y2-Q�b޸����M)X�@�Z�M��y���1qs`<��M��S@B�b!�\�y�%��lɀ �Ս�"I���ѧ�ݥ�y2Cw>X��썊Bڼ����
�yR�]�W�*���䎭?��Hg�=�?��R�ӫvhT��v̺@���y���3Y��i��	u�'r&0X@HJ�g�t8q���g�*5��'}*U���)S�%K�D߷^����
�'"�-�2�\O��p��N�O�=1
�'��Qm���	Q�B�K��8�*O:�=E�@ǫn�\�� Ƈ_���+����'�az"N@1�,�p3C���p����yR�D�M�:�I�3p�v@��y"D�;L��J��Q�}�h���ۙ�y򂌅nRą�t4	4m��y�E��5��y�+�:[*
��3����y���a� ���F�L���G�y�*�9\����!���ad���y��&�T@�(��/��ۢ-����?Q�'E�����^��!A��S6�����'���@�N�_7����a%� ���'�@�j�1U=�����>g��
�'�4A�Dg�G�1G�H�
d�b
�'P��SfI	!�&u�Q"��O_�T�	�'pe#1gV��)�G��Hr�9)	�'J����H�y���<����'	>B&(0 *�<�AC�)HFa�'ạ9�¤8v�|Ia�J3/�%S�'�-g �2���P�*��O���'2jl��W�$���g5���8�'
b��N6	���ǁ��*�z���'��9��H�-f8ef,X�8�lh�' b1��L.�����ҵ,%t��
�'���ӱ��,�r()R��+8<�J>���E�d#E�_�h�F��EG��'�T�d.�t�eE%c~�26��.��(D����霴x %A9���f$'D�����OK���G�
)�p	�c�#D���ӡ�J�Wb˂u,%��"D���3�#X�rɑ5)�LQ�p��4�O��!�bS�=� ��E"�/y�9��IX~"&�`�\@p.[&H&I	�y�hR)l����"�	-$+^�����$�y(ߙ��X[�*T#{� ��iB��y�b�>U\!�A�ɟ��4IDǆ��yBB8��m�u�@&uh�A
$���y�L�
� �y2�܉lք�bۭ��<A��$A�a��蓨�8��ke$J!>!��7IZD��%�)P��1tID!�D4u۾Q�mX)�,�Ѩ�;!�_!��[����UB�m?H�!�$ҥ@M���M�{��%/{�!�d�4Ra^@��m��(�ȡ�S���}!��L1g2�Qf��bN��3�+ܭ(�!��L(CG��#@�D�o�< &+W9�!���D�S�θ2��h�J�2;�!�
�Qf\!��^b���C#ǉ�!�DӘ-��%��*.] �{�oN�]!���B@���'�N$;�r���7*!�D��F�pb�	�g�*���B80�!�$*抉`�����|B�K,�{R�|B���qY�]"9�F��3��{+ўd��3� ��3�/X,Fuv���h�.�t��"O���q�
v^����cꎬ�C"O��J�� E��Y��Z� px�"O�Ik'ŏ�b�����1&�ҭ2"O�pg"�'a:8�b���1}�´��"O�9h�N�8g�^�i$�Һ��CB�'�ў"~Zw����љ@�	&7Yz�хi5�y��Oo��4c�:*h�m�&�7�y2%®��`J�<5Kޑsԭ���yBd�h��%t���x8�3/��y��v���P���V�H�B����y�8$����甪P0$�`�	 ��=��y�+�+?z:��+��BԾ91ѧ��y2�F'h�� ����<�[��(��>��Ob��H�oRrњ`"J�����g"O"e��c�x��c�5w��a"O޹��j��.<07�N�"��-x�"O"�%��h xb�0l�n�A�"O�L�3�0s��Q{V�l���i�`�'�a��D��)���%Úma���t"ʜ�yr�S:��Q�wo�k��"��I��yR�BM���f
�]�&�`'��y�� ��� �^�L���������y$�5GRD@��E�Da�UE��y2�P2~�d���Ӓ7�vY�E�Q��y��"��J����(,#��)�䓣hOq�%�����A�2Q`�1;�5��U����	1\N��p��M!5t�y٧ǐ'qQBB�	�[ZVq���иr�ʈ ֎NPJB�	Wޑ0DҬ6ޒD�G��[��B�	�e(ģ�N�������?<B�B�ɣQ$����b͟l��$Sw�I>VՊB䉸F_$��bY%Iu������u2tB�ɪ>}��eh�/;Uz���j��j�`�O��D?�6���k�L�e�c!��_+gT�� ���8?<���I�!��/�${ �K�_�Hp�q�!���)ٕ#r*(X�j�((v��t"O`p
!"�J&J ����&��+�"O�xp2��cF^�bOb���Y�\��՟h�?�}2e`��3ݰeK�M.�}Qa!�k�IZ�����y�[� X�70�S3E�4�y�H;i�H����.8*�}�@ �yR%�:6�r�[3ň(+�"r@���y�/� b*��̌�.l�����yҬ'`tV�L�-#�hGNL9�y"�!>����.E�2Dn`3G�1r!�$�c�	j�Y�6G�d��ΣB�!�P��wa�xQE�*"k}!�\4=�h�C�ܱv?ZXӂ�8l!�D�r,�"&�;n"��	_!�d�{H�$�R�>TxQ� 'oW!�dX������.1[~d��n7h!�$�*k�2<�7�U��x���ӭ%Q!�Q!6C�QD��M������}2!��:l�d�'��5r@��2�V!���)q0��4dǎpj�9r���-n!�$��O銙���|O����oR w�!�DF�d�N���ק2����j�!�d�+1\�Q�T��n�Q���.w]!�d�9HA0�(@e@�R����哪pX!���ò����H�MH:dϻ"�!�$ѭ*���a%����a����?�!��
�{^XiS�@
���r#7Xp!�� �=��N�^	���Tm�8�,��"OPmp�&Gxh��b%�Y���J�"O�mK�@܅w)f\ s�I�t�j��"O읠��71m&��G�88{\9hs"O��`m��f;؀k��( \l
"O(HA�-F�Y$\ᖪU1`AvBt"O�`q��#�`3ǈ^ x���jS"O>�KROРd��/�b}Z6G@�.!�:A�,�Ɉ81�O�f�!��:��0q�"�7d�	ǀC�	�*����M��05�-hC�I�^F���e�
f��ꔅٻSS�C�I�^������)�����G�f\lC�	�9Q����u�Y�� [�@C�ɰy�!�+-^���S4nR�e�C�	�ZՊ���#��戱��*eƴC��C�"�g_=T��zR�_��NB��n�PE!�G[�n�z����JB�ɠU:8)Ȁ"��Z����2,D.��B�ɐU��	H����s��d�4덐�C��a`����H.N���HBC��,K�2�F�U8`h���R�C�b#�(�̗�s�䁑�mѽw�0C䉛�� �7������� �z��B�v�1wB��6�X��� S5ŪB�	>M*���p��M� ���i�%j��B�:!?̂�ęA�,u��Ǌ�C�ɰy,�5*6hËB0m ���PI�B�I��!���U���%P�O�:��B�27�Da��#�[�d�h0mP�z}�B��+K�����[�R�rP���8 �B����4EFF��LYӇ
4%�B�ɿZ(���B*����ƥq�rB�	�s�~��& ܟ2AFu���^�M�fB�1"�d1z��ޓ0ze��.��B��/@������"x���W�f�B�q*��bլ�<|�9k%�2so�C�I�/��;�)U,v�Ѫ���_<�C�I�bd�r��*uS��B'_�NC�I=UD�c�)Z37���7�ޅ�ZB�I�#���jTI�=��T�e`[=،B䉧a�����E�detܲ�i�$�bB�I;�m�Peӌh�  ���E�6B�I6���A��1G���C�ʸJ�TC�I#a(h��u�R�}�>D��ǅ[�fC�ɨ)�H$�":�����!�C�	�"iԭ�&�7c�N'_���C��&x�^A4�͔y���@Ϣ~/zC䉖5��tK7��	��M"PB�B�,R���5 Gu �<�'��(V;0B䉀:��#�ZFy���Y�kg B��6 耀�CƇ.� �@�ڷe�B�I ^�D����)^#��hV�� {�B�	#�t �$̈�+j�HR$�6U3B�	�Cn�y�LO
GR���N�>=2FB�	�U�)`e ��\�a�P�^�u��B�I�u 2��^��x�Z�̝� ��B䉁fR�lq郴��YE��Q��B�Ɋ
1�̊�i�����Q�`[�C�	� �z��mG�Y����i%2��B�ɟ����A����,�$	5|�B�	�e�����FϤĹf(_�{g�B� N���Q@������ uEBB�I �.��&O�%����2�� 9�
B�)� ���ϭ�Pಯ[�B$�5"O�ɲP�+wp�<ږA����yK�"O4���E�2r�	I ���dC��'"O��9�'^'��ˀn�:{^�]re"O��	��M"Y�m�
�4\嶵k�"O�a'!R�l�0 B���mZ$"O4��)֊^��9�(Vl���"O��zS��u�X�ѣ�M�A�T�:�"O<�s�hR*)���Æ��!'D,`"O��0�O�*�uq����uf�� "O>�lZ/*<� V���"�"Ol���jM�T �P1�V�$"Oڭۢ˚�z�0�H�nI0�V�8�"O�$ r��sҒ�ِn�_r��3"O|X�A�(G�����^�����y�gCCr&U�ҥ̑o"`�����y"�L&(S^��R���fPJ�����0�y" Ġq����Ae�\3f�8q����y"fT7`�¤@�L[_��7�^��yh�
�`׍.�����N��y����(ÂH�fr���2|��mh�'Ƥ	P%L	<݌���]"r[����'a����f� Z&����dP�pdx��'�jA��A�錙��$uB����'M6���Ə�@0Q�� �#�t��'� @�.�5�}J�GɐN�ؽ�
�'L>A��U;BBtbp���v	49
�'��
!�ӧn ~Dl
�'�@�ڣ-��>�������z�= 	�'��a��
"y�蕊Я˥B�pdS�'��`���O�q���&���&F��'.$����M� � �G�$D"���'����	9�J�y�m�	��"�'TDy���O�!�OU����'����cĝ:C��LHG����	�'�0���ߍX�ɩ�k�r?jP��'N"�'U�.<�Ыk�	;�4���'��2���E��dbR,� .��1)�'Z�i�`�RF>��­ �'\bA*�'����f �d���q�\�����'�tB&ńwf�ʢ����2�'^VDX��݌Z�l����2�*�`	�'Dę��ᖎ��1!�Up�ݪ�'�L���C�X8�&l�Hi�	�',*%�g��1���sI?8�<1Q�'�6�*���%/�y��ʯ<��Q�
�'<t�$�� J���<�.P�
�'Z� B�63��*��vV�S�'�t@���H6aF�}ؑ��=�����'ΖhÖ�ڠu��-r���@)�'��(�@�Âp"�J���f���'���ʝ�'��{�:6�0M2�'S��*���`�"�blT?,����'Q��zU�U�7���8��0s�I;�'ޮ}�Ǆ�>l����ʯ'>a�
�'y� b���2A�Vp�v.L#Cf��'��)��@iI`�-���Q�'����D����"�B�X���`	�'�4�2�H^��;AeW�O)����'�N�#❦\��1���Z<$I#�'|NI�IX�]z��b�(Gt6�1�'c�t����By�LjA�M�=�|T�'��iڢN@� (���Ȓ3���Y�'��X1Ǩ����	�A���D��
��� ����aY05C�f���x4"O����w^B�+Pa�&  ��"Ob���
W�@��A�� }��)r�"O�`�%LUgE(��G�ӆ>��� "O��3��G��"\kE�&E��4��"O����Ȳw�P�����\�@(�%"O>�Yjނdg\@q���4}��!٦"OZ��/�9@��X����t"O��i]R������=���"E"O�H
��3*�̙p%�#U� Hx"OT|h�,�� �X	���Cɀ��\��F{���-ph��U&�!��T��2-�!�DV^u2�1#H�>�L0p�@@#�!���s�&�;f��f�L�%/�{�!���x� (��H�o�����Nĭ!���q�$9}J|�':@4�g@�������p�(��'�J ɒ�8O��t��G��c�6���4���A��@��!�?�xh3�LJ�",jL:D�,�A�Yʈ��an%d����c6D��C"��o:����Z,)�ps��>D�X1�؍cW(�"�Y;O ����0D�����][NT��m@hh�Ь�<�
��v�p��Z?�$�;��S>\qJ�G���h�6az���(C �[�H^5;�~C��4c,��%4��l��!�?5]R��ē���S�,fչ�#8 v@��`��m"C���q�CH�9a>*�s�b�@�DB�	?u` jE6_1
���C&�.B�'Z�D�T���m��щ��BdT0����h�t�>%?�"ǍA�>�ҽؐiZ�{+D�U�<�O��'v
�W�� <p����J6-�d���'�Pt��/`n�8���E5�L\���d8�'~����'�
G�	@Rc)�|��ȓ_�1��7n�4��IF�A��܆�,�©����~L�%z�`_G䍆ȓ��ȑ"��p
���c♄ȓb�e�p*�%&��f�Gd&0�ȓol�ͱ��J
t� j�KϹ���c��?,Oڬ���X�!8aU(A8vԴ�b�"O�,`"*�,�2�b! �1h�!�K�_�<�Q�Q�=OL|S�+]h�ў|��ӄ�zt��e�	fГ�DʀC䉱8'��+��F��*@BF�r�T��?�{R�	�'7�ppRN=�0<�0��%	BC� {Q�x8��g�܍�DZ�L���n�a}��G5{x*�B�#��X���<�K�ؖ'Z8�˶��(��TO����c�@��y2ʉ�������@�  ��(ިO0"�d@�0��0��"Kr��p���e�<�Q.ؐ\{��b�"Xs��h��W�<�bJ�()X0(q0,�4��X�SR�<y��	�V�f��J�T�Q�C�v�<i�ȗ5$��!�e�!�0%��aSo�<yt�ٮ�v���X�q�J�:b.�l�<��� � ��I�i�����h�N�<i���,2r]�tC߷5Ah�����t�<�����L�2���_ͼ�%fKX}"�)�'4Z����*���
�f�!,	����[t0�z�鉌0[de2�ě�r�u�=Yۓ{=\Z�j�"j@�3�ĕ�)���M���R:I�#�	ǧn�q"/�~�<�����B��N`H,��@�$0�Շ�K�`�Ѱ�)kp���m�.*3Ь��	\�'�8$���J�^(���
X�j%8�O�-�O� A@��!@�*P�RDȥO
�43O���J�S�Ov،�Q8��#5�6v%����'����B�7$�$����v=*�(OJ��$HQ�b>�@�ݣ!*���`�8ud��<�O�`�'W@����/YV	)%�	2���;��yy��'}x ��Z+.}9�`�x��Y�¼i[���O���H��)��u�׫�w@��z�'$�$����5$�1Ȧ"�@�"@�,�(O?�$�/�Ɂ
H�
{fY����?!���g0ڨ1�@<i8��Cʻ)���=O�i��&?�"ƣL��U"O~�@����EM�5)"�M��9�$�O���o�g?I�.ǲgB�������T��8���9�y���2Ҋ�`0(G�NZ �	7`#��$�<�H>���ɬl�d�y�G�KBPDsc�r�C�	r�e�EǗ�l� ����
ѧ�ē�p>�'�
SK�d�Q�P�C�ƞu8��$��'njI��d�%�f�I�^e{`�m�<yT'�(Qgx�"'+2Ƹ<����h�'� �F�4���3�h���`�N x�E(���yrÀ8�L�z���8S���m,�y��Va�T|�Ѡ'Q
���u����y�kX�/��i�̑#NA%��6��D.�OX�VZ<f�. ������P��'��	� ?>�B�+	d8��`�⎧�rC�	#Zb�ѳ�B�9(�����F�0"=���T?=s�B<Q����(}���P��"��F���'*JV]�U�#m�ƅx����( �H���F{r䐋`�Ё�'��=6+��ɥ
��HO��$�MSmX3E\�_�q�U �#,�!��hT+�H��{p�pwOX$��hD�ԩ+}!��zU�	 �b�ZG�S2�yr�B�PV6��c[(�Vl��A�y�l� %D��#ӌ8"X���O��ybJR�$
�9,�&���V����%�O� �\�O�h$3D�L�
i*�Hc"O���Ξ�G5 �����,t_x���"O�D��͝<]f�R�o�>1�R��"O�%���A�m12o��`08a�'Y��OLԨTM̕kJ��!N__��@�"O���'bD$s�tS��D�(f�s"O �r%�53��1ɖ�H)f$��"O�)b�	� |�`�P�u`��X�"O��{�$�
H�b��a�à2?v%Ӈ"O���	��gi�ۅő�mB�8���s����j�E�4�D�CR��sC�m!��M�oj�b�rY� pW⇤�!�Z$��Ձ߭@���p@ԡ~�a}ҕ>�E(�I�
�(�o^�h�s����?�/O����(l�x��/16�d�r��:]�!�DWPC.��#-h(��֪N�D&!�$�v���ۃ��\�"]�	��IhX��&
Y&�P<� ��j\���e+!D��Q�O@jA�pF#>-R�{�h)D�sugM8�lR�˄;&�h�H$4��C#�,U�����S�p�lC�h
E�<�¥�B n���$�>A�5#Cc�~x�TExB-\&U�͎�&*�,Z!����y�V�c�MX�Q5j��mS��y�� 8�9b�\�,? =�����xr�ii�i���߻>��mc��I1&X�6Y������'�v�>�w�ۉP�	�B�гP�@����'LO��#zyr��L�19�`*`@U�:!�'t����	�?��xJ�ܳ$��,S ���D{J~� �����{���W�ΌN��H��"O��p��� ��A�-�TyV�R��	}�'��ɳD��5@5H!Q�dis �N;�B�	�g�V	B������,�%h�B��rI�]#��N1)/X4�+�.d�B�w8�Y	�A�e�L,��F�X"C�ɉT/��Z�M�E,��j��"<q?�S���Y�IP���gR!P����T"���yR�F;/v|`�Z�_�*��7�=�y��)�	z�����X�Q�U[b[0��ȓK69!p�"��!�s��M��%��R����R��$�^�� �*a~�W�P���7
�xth�l+d`�c$D�L���:B��h�G��2��5S�$0��{���';wҥ:U
S	\zp0�"�:��ȓ6��4`�d֜\[��-��'����J������p}��;� O�"��w���1eU$f%4�Cר�J<���ȓ1p�D�5���+��%;:�B&"OI�e*
(7���$υW&��#�"O�8"S�&��р�0A����u�6D�X8��%U��PR7��I���S	5D�,r�J>"*  e���礜o3D��u�B�t]�,ID
<#*f cqa,D���WN6����U��/T@F$y�+,D�<d��)V���*uC��u��ɦe(D�`Z�I�
&@��5�m޵+�h'D��
T�R�_��)#C��3������$D����H�0uziƃ^_��Q�3�$D�Da�*I �H�2f�F�{�~m�B%"D��xE��C��qD�@C���Q�:D�����	B�|3v�
���Y��8D�c����%j��҄:h�A�$6D���� ��(QhU�w 5E�� �5D�����X��NF�`iz���'D�ԛ�&�6d���9���j+ qj J8D����F�agJ�ԫ�]���Ja)8D�����Wak���I��7D��sv�L�y�| �_#Dt�"�M6D�|�ԍ�0*�v��ě�Ql���63D���%̞ R���vE�9a�@���1D���w�� k�`��f@W*3��,�'1D�Ȫ1/J!�q�2�Ӡ}w����3D�PqQ��$S���x�+�-Zo�0c�,7D�����<V�Pi0��d<�dF #D��(��]�!��3��x:Jx !D���w��8�LR��9����<~�`�p
��]�#
 LOt��6MB/t2���I�� 	Z�BT"O��* ��2 �ɴo`x�"OEp-P�R��@�l{^���"Of�J�-ѽ�Z�CT[�[�i��"O��b("��Jc�_&P+qkP"O�Ջ��V3_�c���z3"O�`�n�o��U��d�7��8`"O�p{��@'H��́hy�؉"O����(>$���ϐ�F�$ڑ"O�i��W):�3�O\�1�6���"Ol�C��"K�q�7nJ�
���"O�ɐ��U�2QP���D�$��6"ObP�gL�u���3NBxvv0�a"O��c65"��Ȋ�PTy��"O�0V,$A���Q��=^^nĲC"O*M�匯Q��Y'�VATq��"O����X�b�jhQ@$�,X�l��"O� ~�ۥ`ƘF��a��	4$`��E"O�؃�?zt�t�6�D0@�"O�4��R�a�2!8�T�}�@�R"O�D��H� ����S�C��$q"O┐���i���K��Ǔ/ߠ��#"O�J3"�3Bhl��Rn��n�"p�"O��p�O�Y��ã �>&�Źp"O4�r��Xy-�I��6;�P�"On �e�N7k^e{`ΡO'xXK"O��DB��:�Pggø0K��S�"OB��r��H H;�L�+�J�"ON�� -"אm�b����*U��"O�@2W��gT)3PԳH_�}	�"Or��D��5�J`�5
�+f9"`�"O|��p�ɒA�<�P�V�W<lX�"O,�	]���l�1�s&��p"O$%�(S�k�ҹ�MZ�ic�0�"Opm��Y\�;��S7o�h(�"O����A����"G)�)~y���"O.Uڶ�m.�����g��E"O.����Z�k��X�2F�N�h��"O��`��3�d����Η9�b4c�"O�U�0*K��\8Q�dI�A�,���"O>��F�*kDڱ � �:YxhM�V"O��iạ̇̄
�"���ܴfh��a�"O^U���%4�ᆛ�[Z�Rt"O���&�g$� s���R�$�{"O>5�&&} hu��L,2�j�`'"O�����X��U���G����$"O\X�6�zW�-�R�P[�"%�b"O��C�M��1O,�
�I y���S�"O��EFN�$��&FPT�x��T"Of����M/��c��0�H�Q�"Ox�4nƧc�¸�C��8�l��@"O��� �U�"�@$����B�:1"O���n&F�h�h�>v�朲�"Oܙa��9z�0$�g�X*�	@"O4E	��L#�6aY��T:Eʶ"O���KȨ[Ѩ��3��m\��v"O�xh$�'K�(�+f�R���"O,��a��F����(9<��0"O�m�S�
-Me� #2#(��U"O��
�ER�x @�Ԗ�7퉠�@q���S��!D�](x*Z5���/+��B�	5md�%	bn;���i��P�f�!�`̡��0}���'�`X2,B�\-��J��[��U�'�
�+�n�<d�@\Y�f֛d�*�+�"�B�[��ĔWm`�YV�",O-���m��H[�.������'*m�ECW~� r�CĚh��x�ǐ�y���O��TԠ��
O�ة��˽E�qy���8����T�dD�)�2yGη,�8��-�S�sx�I��:A��[��6=HB�	��r�U��]j�SFH�,u{�q�G]��ðֹd��Z�'���v�M~n���&�ѿ]>1���^�,��UKw�Sz�<!�ތs�Z��4�)ADp`����:R���0w�J��Z��7Il�oڽ℩�)S]ܓ"�P�pT��%|�@:c!�,nz����I�c*��F��8��=YB�"��s�`P�h)� *|�5��a�WL88Eo#�����tJ��j��H8O8W�1OJ4:B��S�
 g� �Z�J�����#�D,�9`���	WqFLI#�@�XD�0��<�!�F=Z�&����Qe���a��{�n��u��+m��IՆOcf�JG>\�2��!�?��3�t���$Y�CC�PeeK�~P���-2D����(4~Æ)*���)\���a��(��t�g�##��I�t�ő�5zɐZ`b/�I�bPf�"3n�\�n�HE�����L�<t��!#�'d�+��]��8���N�3n
�y�"��*�b�����`C&љA#��	ӓP�X��&�	U7Vu���[
��'�j��DA��v�A�
v΀s�J�+O:�T�P� PH�u�	����reV�!s�4"O�D���K�o�$��sN�
az&1[��H'Z#�Ę	��=��8����g�X���n��d�b}(-k�1�l�́{�А�!�x R��'��t�Q�R��E�oάn�>��掟��]`E��+����6�n���ѡ�i�A� �^�_�qO�������u�!V8s���J��n�'��-��/��]�؉��j��<�����	̞�\�(�IBL��ٻ)�7&���i��'� �n=�p=11��0w�(M���C�b5�d"�BlyM�
є��ɪ�\䫕�\�H�vh��O����@kĽ^��j�v�N���L�$�IS"ON�s�;i:�V�Ѵ8����#T=3p�K�fӍb�Y�S�ً_>D�o"u�p��[�����/�yG,,���A1+��Hn�h�Ǣ���?� �	)cj!�N���@}���ӑ
%��(�旰��#q�7J):�@�j� �P��3�Ji���|��2��!9B�S+E�n9;'ϐ��O�ز�ȼL��Ŭ\�=@�u�P�̝u���{!)�-59q	f%�2;���H4b���ʲ(����Ĕp�Q��N��bc�`@eO��2��(Z�����Q85$\}��IL#��"I�*$�x�㑰J.�tfH�N�t���wh<���0df��x�.ǌO>��

F�'�Zu�& Ԝc��D{?�`�+)�	�sCv(����+q9@T�B(�.$!���}���R(R�O]H�'K'_L�7��(�:-Ä�d�p��<AǤ�n_H����j��]�M�d�<���]8.@���N{�0y��:@
���%���R��M���<c�� 5����4,�UZ�4����v���1)��-A<�!M�30�l�JQkB�g�N���b=�"��64�|�R.Hl���!���%�x%��,�I�x�ɩ��wF�xC�-��M��Ii萺G����@�8O��B�	�r|�5�˘t	�|Ȇ"M����J�A=]��G�B�$���(��I5 ���	�aO�IJv�Ih��C䉺o��6f´-ٖ�
C�
�$�����J��ji>|�2��1��z���)��)�E�Ȁf$DX�p�H��p=) ��\> SrLܢ�M;Wl�>��PFF)x;�	�V��v�<9![�ݨ!r�(Ӡ|�:�Ӷq�N�����l�i0|G����6~��ڂ%�8��[�ٶ�y2I����q�I�(n�^�iG���x9�!�]$���'�>�I,�����N�_�t�q��{�C�_�L�'���~YhP׬Y����D.y��|A�K��=�d�k����ɐ��do���0>� �^�^$��*dJ`�¾kM(�r�GZɖ%��Z���$!V4K � � ��N�QDy�	�[� �F�t��#`�L+S!^�FN���ȹ�y"O˿|@1��9H��xiq���y�E�E(n�j\��m���y�嘗bW��*㋃�Mf
�k�)��y������c�E�,�H���f֭�yBm��K��|�`('5V��h� �y��̀~2VD1��?#�@r�]����'C�r��K1B�4 ��m��L>�S,թN�$�IV|=)g!g<�s���;tP(�U�yB\�*�◂E�"p�C�G �R��D�.p-v!PϓEn衔�e��(��\�E��U��ԣv5�CƁ�j�!��U�^|ظЂC�
�]�w�^H<����?���(�OL�f�\��3l�Dy�#�>5�E2Q&O�a��A��5q=��~zDM�5 ]& cI'k��P���G�<��*���Lx&H�#e�2��C�����0nχa��-Rvi�
:h�h&?1zV�x�Ѫl�X�wfP�%��j ����?ك�Q���=�ɸ�NɩN��<A��$R�Zh�@l��螀���A��@���~e@9yD`-q�V*��U�^ >�?���W���;�(M<T�t��4 ޛS�M9�
�p6i��k�6{����&�1$�̋b���:�[��BqЉ��<��]&o���.�,_��x�G`½��c?�$�D�$����%CL޵��.4D��yw�S�+6$�	��W�Pc��$-�tA4]��Bs~t�+U&��CԌ��~�#M<Y%�L�X�� *1�SQ�б:Q+�m<QhB{.�J'�������9oC&�
�g(vw�p1JM�#L���m���
�EÒ����@���IIz4���_qD�
ۮ=�4��!R�A}��� ��U�ޑ10"Oȍ��B" /�L	�eQ3f.)�"O.@0�Ϙ��bd[U#I�li�@�E"O� f����׆1��+�W�U�c5"O�Q[6l�"#�a�n��C\t�rw�'Y��ˁ����ɵz�$����}˲��d�	�6C�ɴ3��r����S�*=@�)O$L`�b�8P���Ne�\+��S)p��a`P�_7�ҁB�&�BB��=�6����
t7���b*:d�K`�S=���e��!��L����������ا,�\@���/4���U�U�)�B�zo�uN�^L��1"�)�6a��D���f�$~dڠ��̓&_���M�}n�L�%Z��	�>��1/W�؂$�vO(h�B�Ie�*pZī��8p�O:J邏O�,HG!�9L༽i�"�f���Q��R< ��t!Z�+�Xm��g+R�jQ���B�|`Ȉ���v�T��B��'< D��>�gϟ+e�Q9B�N_��� �`h<a5$���<�+���,8���@�-TG^)�Ў���T��
�{4��s�ٯD��H�AɅ�z�牯E��T�w�	��~�ΓGk
�B3�0\��д���S�"Oȵ�#AY�t� �A*(�R�	���**�X�!� ����
ܩ��Bjx��ɀQc��
�'�Tx�fW?i��!�	X�fv.t��oDr�O,|��Y�4#7�Ͷeݾ4�5��&9:��!D�\�'�H|@��)��'8���C:D����|m�Z��ț �����9D��(�@/`�z%k��P�yP�0�E D��#f+O�?��ip�ѳ2 (D�V�!D��ÕJ�*�8����"�H��+?D���B*�1dn���C�ub�y�6�=D���`F4[d��Pc�
���p�<D�$�F�R!Z,ڥ�4�F=1,RPZ7,)D����-�N�� ��!T��3�	'D��bSK�n��  ��<K���$D�<���:A�J<(�ȑ)_`����m1T�P�t�"�d��F� Z���"OΩp$B�(g����x���"O�XqeN9]5�Eq C������"O@�8U�(q[xm�_9(�� #"O�$[�B�7?��01v$W@��Piv"O���f��	9kzy���O�x��"Od��#��a`Ri�b�;N��uqW"OH��#dJ$u̰S�R
�
9h�"O��!�R�q�,x���La�� �`"O����ę%Ot �d^�E��U�W"OV��$�4�r���Y�BK׌6�!��,�4*V*�*U�Z�Re�+�!�dk����D٩�6liG�A�h!�d��L����q���h�pp*�"λg�!�$ķLt�P����{��5 �=	�!�D\�tnB�A�:L3��ZN��!�D�5q�Z���ݯ 5���EN�R�!�䋺	̠XJU�J�d2�y����b�!򄍼G&yZEN֥B2D�o�e!�D�s�y�*�/w���YA���h)!��ΌX����ŏ�LA�]�U��!D���g�Ɩ7���^�t�2��U/z!�dߝCK��i�)�<�hm�č��!��v�1�$g/U�̐U%V�|�!�d�2dCD@���	,e\rhr�KA+�!�DC�J�J��ɪ[Db�2S
E	�!�d��9����V�JHr��c��]�!����Hf�$.I������+�!�V�b��R���\"Hx��iJ�k!�$��rY�QI0/���(C/H!�,sπ�)�@E(M������,n!�B]}�E���xZ�Y)���b�!�� &qS��̸��� $�<Ŏq�s"O=phρc}bU��A3m,m��"O �f�&*�}��)Bl�1�"O 1��LT`�t�5l�J4�%"O�x�*P�X��]"�b��I�Ř�"O0��b�X�eX�9c�Z
�lt��"O"���Ŭ&��B��T��9��"Ot��7.�p��X�I
~pp\Y"O"Y���ʒv�(��!� q��q"Or�J e�3z7��V��Ujx�j"O:��4.��a��<�b�ŭ0���"O���L�A�$S��CV�!a"O�AbZ-PX82W�S�J�ؼF"O�2p��n̻�
�1�| �"O\�9aꎩd�`����
��)"OX��ɏ�{M�ZA��;���P�"O�`�f�LC�1�Y�}�^%
1"O���lD�؄��!W2"���`"O$�'�P�q�$Q���R�ĩw"O0��fK�NՖ��f��@��JT"O��BA*O4��#l���d�;�"O�8"HQ(_�: B��P6r���E"O�)�h�)Z�@L���(+�Z�"OZ�����sp���T�����X�"O�I�'K�@�F�[rc\7[�Ԡ�"O���p�I2�@)$�.`���U"O��QD�I!T}��^�$�:鳣"O���qjS�:0��6�Z�\����"OL032-�!
DiA���6�\��#"O<�k�b��K���0� 'SO����"O��� 9�z!2a 
�67j@3P"O�1��o0~RS	�c�|��"O`-��锫4(.Ջ`g�*M�$�"O��91!�=~�������N�f��"O��@�׏	���*S�+���T"O�%�c��U��QP!AؠV��\@�"Or���*��w�	�$"4�"O���Y����RNE {��"O�{FK�i����®��:��#F"O��Ro�]���� �
3�H"O���L���P(���56�f	�"O"]Ck�%�L1y��)$�2�ل"O<�v ��\\���9��S"O����h;��9(�L2���[�"Ozy@�h��j�D�`���9g"O�@��*��$8�A(�.�m�H��#"O�B7斩Io8��-��s،b�"O��:v�_�T�ġ����+�n�sG"O����*���A2P�^-��"O��)���2<�hsD`Đ9�L�[T"O����=`wp����B$w��Y�d"OX-�CL�7#���A�X#.ǒm�"Ov��d�����2��/#��q"OLdJ꒳d϶d��F�5���6"O�к&+h��;��D0&�.p%"O���UΏ�j>��_�ɱ�ՔN�ў<���9>k�>���!Po������;����*1D��6�۴*�����C�6��ɸ�Jkӄy�eXz��O?7�����EK<!%��Y�{(!�,k�V�)�%�8
x��3$ӧD����).g�i�O�0=y��]-^w�Xq�Y>u�}k���G8��Q���6� [w+������V��9�fhS�K(q�!�D��BH�a�a.E"V��q�$�ΑR��a8����V �'E@��f!d`�'?��;q`����H�b="��]7G#�Մ�S�? ��ɠkSt���h"ǔ�k���ɳc��*ag
�&uD��O�`���B;Ubf ��y�m�qwQ#���40w������p<id��"����cקlGvh��L f[�)H�	C̾��ǨW<S�J��:rI4(6��D�azb.ű
�J\+&�*�E+����dP1Q�S��>�܍h��҈i��i�<y1��_)�(��P zЌtd �d��C�ɓd��H�����D�B8�b��i]d)��&`Baq�J#/��d��Fg��P����@�	�-5�21GV�@5���t��V��/��"�35M2�xgf'&��\"��V�
o�v�S��gi2)	�K����\�H��,k�i)�={�vm2����,��͑�Q�qp��?��)и$ڪ$���G�AO��I�/ީ\�V�H����o/@��^;���-O��h E��z��z��Gd�|y��V�Z�|���)��XvTqR�=E�<!�`�8[��'M���TH�G���[q�5 x:��Q�B6@)����'+bL*�I2'òA@�/�,.a܅J��%q�J=KR��������F�*.n6��fL�םJ}��e��c���\��p��o��:���˧�>�O��S4�7~z����cO8e�gɱ�X���0�a�� |�}ax��Sn���'���)�CH1�|��$��d�`p
���T�#�> �e��gH���id�^w����U��&�3tn294x��O2%�𯙢u��u�	�dm�:�`U l)dL��	��0�n��'�Vذp��L`ɧ� G� OfL��G�̣^*�0ZC��6tP�b�Y�Fw|��O��`��D��pA��h�8�@�d�4}y�HGl�8��O�1��hC�|JeȐ:�
HįI�O�:`C�r�<	�� �q�f\���U�ܰrMτS� l!���l;�A�'��XD�,O�( �Vm>���l_�-���5"O
}�rO���\�%�we���P�+�4����N')VZ�H�!<O\�	�f
�B�x��π'�P����'���c 	�.-�Y#��P�A�\���EF�:^�����w�:q�',�qS�jӞ Ȉ�UI�/&����{Fגz�u��Z�T��I���G�	%�p�'��_{�t!G[��y2��!������:%�=�7,+D�T�q�
X8[�¡[�'[R=F�,O��1�@,2��N]�yE:���"OhոF�
d�kt�+p>t��֍9gD�6gкC�ڱ
דS��(�T��w�t��S���&\O@�J1G^+��E�!
w��1��:0Fp {V���]~Dp�"O�D��@����Q�=��d�Bvu��	S�Ox�>e���]_�}2g���S���2D�6D�������TSA'� J�QRD��(w�1�J4��	o��~�éI�rY�%��0G01�g\��y2�T�r� i�I��c`r�@Ff�
�?qG�e�
�&'lO��9����B�:��w抱x���AD�'V���N#C�Bb�A����+�!d�������yR YjrJl!���$������(OȘqp`٘ꈟ��që8,�B��$遃�N���"O��bg_ċR������A`"O�E��̙��Uk����GLԩS�"O 	ʒ� ��������f�xR�"O��kN[� �F�[ōҟ;�}�`"O*A�wgQr3*�A���?t��m�"O�4P��  u�(u��'I�} 7o�to�pG
"Q�:|�
Qq�q��'W|P�G�&"&��2�N�4��'Vx@�$,�>F�Q�#�G�/�.x�$N��X���K� $=Sz$�H�&O��yB��c�(49q�K��2)2�k����O�e�� ,{l��hP/+|M�Qf�yP�L4O��xh�v��/02��'N����]C:4��Fа;k���.OT�P�D�����J��#��-+W�ő��O������!LB��F�ī3���;D��+����E�p�@�N[�<�y�hX�4�<b�2⾵����(�������K<A"͔7qS��)$��n��4��&�g��tjR��4\�!��@ʲR�45Z�Ě) �� ��X�0R rB��*��'�\1t�Еw�ҥ��(��U��J�����@]�*7jO�FXE
��H�7]����-}�z�����!h��pc�ɼ�xB�O��@#�-o���p큄��D�-�$��RC�����91������D-t0�գ�F+5_�0
2�y�(�0k����a�..��)����>G�<��m͝�b��"�x���KL~��<��,t>�;�郳`=&,�2.|5���[n��1�Jn͌X`��Q-\�$�A�Y�A��ȆL�6X�����<� r�!2��*sf��`���l1&�'9�ĉ��Jl�����]b�H���ޠ������ѢmT*,%%ZK�<Y�d`�]����	.Ļ�#�@�<!�2��a�iB���	`��W}�<e3ghB!Z�GK�]� Ly�<�o̍~����N/%0P�I�������	nD�'q�)Y�%=v������1pt	��'X�Ā�L�5	�(�V�J)t��`��yB�J�v��t�ƥL�O��y�/�f�Q3J�S����'�L��O�<��My� ��s�$��4�\��%�+O�ջ�2�3}�B�cd,Ōqr4�'�����x��vtP��ՎL.4w �sunV:Q\$!*�G��[���bS�'���q� �V�8�Q#��a`0\XϓS�𑣇�gj>HH�'�,�rf�]:&�*�;�mQ�^�a�'r>�!�)U>!�J�������zJ>��������ӈ��%��!'~��p��ڕu>*��F"Oؙ8��5|#~� O�� H�@���U4DA�R�(1TBD�g�d��|���C��XMf�R� �s%��D�!�蕁��H�uKd�ҰD*A<l�P��]���i�&�O���w�O�P2��B�?��@"��'Q6��c��<��T2�3O�Y�`�1Z$�a�D� s�+�"O�����\b�0��OǱ6f
���<��ݾY�HG����Pt���T�׾s7ƕ��]�y�D�Z�4"�@��^'\}B/[�$bN��e�!�ۭ�(��ɪN�㢋_(��Bq
�i#�C�	�T��a2�*΢F���BmS�[�TB�ɗo��QVb׺Bz�CҬR�'�8B䉒_{�]PT�L�!�ܴ��ǍG��C�|&��y��Y�vD� S���C� AA�T�� �= .�z�H�e*tC�I#%���k�1W�Ӌ�60NC��3�"��ř���!��2{C��%+�eʱ�C7X`&$�^Y�B�	����W�@�i� t����(C�B�	��	
�ǘ:m��������B�	�˾�90j�	i��i �"R;"�B��	&}X\��?<��@B����B�	N�t�n�/b�Q���i��ȓr�hl�e�B"G�R8��l���ɇȓ{N����*O�ab���Ԅ�ȓ3A`���:����L-����9B|9�&�D9���g�I;�*���Z�ĐסZt��O[���ª���%��oȀ���/��x��^ՠ���K��
Q�U	@]���ȓ��C$�_�!�L�A�#4�D��!��(wi	�Y�΀Y���xɸ(�ȓ-�
]�T �	���Vڹ|fZ��ȓ)*DB��G
.M�5�̶;�b��ȓh����O;4��D�$0z\��ޢ��`���c�Zq�a͙�GX���p��ud.�UE�99��XY��}�� ����c!$(��9Q���ȓhL��c�4�R}�!�_8�Ze�ȓ?)JE��θ:Um�:놀�cB�����S�M(Tڸ���Ɍ���K�E=[�O=o�C�6���h�Io�6���')+/�C�I�aVv̘0cǁ@~uZQ��0M7zC�+/
Hl�TN�����صJabC�	�.�����ͤW�R����{�B�	#r`��Kd�_�e��D�&I��:��C�U�%�[�.4Ա��L%xuC�]��7�
l�A�VY�t�Ny��'�L}y�����{�B[�'T� P��Q��0�v�OE���JE�H�%�>P�zb����� ��Y�F�Vst<�w����7��]?���>��4E�=�0|Z�E�XG������=-,��Ɯ�-�ˈ_�T����%2���)§��dŇ�Q��e�!�[�"(`���3RW~��6c��p0�b9���Yi>%���,F`Ԍ�$�;(���sF�M���jf��Y@�f'ő]}�,&>�}é�00�|��b�
�nh �8%�ڗ0���Y������,k^a�4��;DNXb,Ѣ�J̀��3w��	"E ����M�g��S�'��PQUh=)d&\�0��Y��m�Bz�M)#��)��O�3}�*P���q�[��f5#w�Z.�?	������"~e&٣#�܌�U��l���ɀPg�92
�'g
\��"�
���}j�*7H��y"�U��()0)��"�0�$E��y�ǈ�%���� �@�f� "B��y���t�hibB��:�n�b�l��y�o\�S�� �d`��Z�Ζ��y��I&O�QC�T�PD!�W$�yriP�Rkp�#PO�GoȤP�^��y�ŎW6�ÆE8c꩘s���y���|E"�'f�����yRȃ9(jf���K�ؕ����ybl�,����2I�-�jY��c�Py�'�-j�$=ۗMQ�o�$qz�@�<��ҸJ��]kfJ�>C��Љ�T�<���owv�X'f��#�pٖ�P�<AR�+/��v�[�'H��Z�Q�<)���0Lʹ%��eW�U�P*6D�N�<Qu�Cc%n�I7%��-=r9�nFa�<��X�2�-�S�%��)j��Q`�<�ы�R���(Q�CL�	ԃ�Y�<�2J��i��t$��
Oi�511��U�<�$ �%J�l�v�	���*�]�<�a@�@����+:�L�0'*�d�<Q���7F�P]৹B9�e�Ŋ1f�B�	�ag<}�%�]����#�D�I|�B�	/j��#c6Yu6� ��0�B�8�Lܛ�$G���������O̒B䉣;�b|�s�@�q�tt�E�A>h��B�I7D�\��#�J�^� ��C<.��B�I1d,��@�V�MvL8�uc��.{�B��.8$�� ���En(���$Ҁ��C�I*"Z��@i�}{"�X�AN#�C䉜JyȀ��h��RS8x����\�B�ɖ	����2p�e� 	3?�C�I Ӧm����iNܭk�%�	-��C䉓� �`�Iȹ��v �C��"T���`O�<�����[^M�C䉔D}�i��\<"�XH�vB[1��C�I9I`����J�g[�x�)!:�C��2��L#�`]�MB͡��
r��C�I�Y2+F��^�8SAF�)V:��'m�A�NE	�x��h�H��H��'f�����L�8�	cCP�E�.5C�'��q�����eF� 0R�:*_z���')�h�!�J
93����n� c���'���0m�m��y�@�V���y�'���KehO�3朹��F:; 9A�'���T�K8*FXD�҆,v���'���eW�H���bC邷T��3
�'+rx�"�)�����T ���r�'4�2���l�(I+6�ߍ_����'U��Y�a[:!@�+YT����'���3�@^��k����`A	�'�6�����O|�t��;�1��'-�ɠ/�%8�yP�nW�;�<���'�cSD�w��\%ޔ0e������ �͊A@�T�ƨ8CBT$67�`�"O�s���)R�j�� оa")
0"OL-��5 �J��N�
=��JC"O��b��%p�����"#�Qp"OA��GK�0�ݐ���zl�"O�hr$�<0i�U�H<["�X�"Oڌ��J1�0B��$ZP��"O<i�	@�>T�e�(at���y盇jLt���� ��h
0���y�N�d��pY� SG�v:gA )�y��q�J陲�
�2�^�����y"g��^���˘�W�)P���yb�¦���A���N]>��A�م�y�(B3��,*���>*��A��y"�_ a`��{�DI=V�����Q��y�J��3L�0�BY�`��a˜�y�ճ!\�(����2G��yB�Ϳ�y������,)dh�1֨�sRÝ�y��	 �%a�@H�, h\Af�0�y���M��P��	�8$�����y�aD�E�f�80BB�6j��K
�y�&�7hܤ ��e����pxW� 	�yR`�,��4���+
0��e�_��y2�ˊ~"V<����U���9E�(�y"/�$H��R�U� �����y�P�46�PAifI�L�0@E�ȓV����G��d�f��m��p\�!�Ũ�en�*b��?[E&9��uV���g�(@��rS��N�<�ȓ	P��"�]&F��-���֤z�D	�ȓDHp,	�  �s!�i��FHyz�8�ȓs)�t*�%��$K��Xc���G<��VkF�H"�`%����ȓl~,i��n�
�b�4�ˆ>;)�ȓ�&Yq�#�lA�@H+�$�&��ȓ	U\s1(�IQ �+�·{��}��goJ!��`@�F�I��Ǳ'"�B剐g�"i{dO�iִt1a�& æB�I\@H�4 ��,�XhrS.7�B�	�6#b��NA�f�P1萴.>�B��R���*��Ƞ$�7D�]f�B�	<���V�DY;���ӛw�xB�@�(�&ַkՂ��A P/Y�lB�əQX$K�cT?$���-��B�I�e�jl�W�W�#����V�T�t}�B�	�g���ꔧB;�Ї�*��B�I=etba{2c�Y�"�q hR���B�I.Z$��zv��$/��6�.<�C�ɯL�D�4�C�j�5*���DA`	�'�$l)�nȶK�E#�! tdY�	�'��\8��ɟG�f��Kt��	�'}�5z�'�*k N���N�2�
 �	�'�,=�OD�#��VP�SdP��	�'~����aI���f��R궜"
�'`ZEN[��^uL�2-��'�0��b[�n)L̐%���>�h�z�'+������8�H50��<XD��'����A��-u���/## *@Z�'����e��:ԭ�+��$�t�>D��{6�D-��|�cmũs���Bb:D��yP�Uv��@�"�ƎiP��+D���͇c�V]R�K�$VXF|�2�*D�T��A�gT!q��_�~�:�	s$D���	S86�f�afd�&pM�2c/D�� �|h��<8����KS�u�:�1 "OjMs���\cd,���!?��Q "O���Ѧ[�r���T)��|pg"O���BZ�(�PZ��84�@"Oܠʷ"$j��5ڒ��ܐ��"O�8q�Ɂ3d��x�����Iq"Ol�Æ�� @�$,A�w�$�"O\�I���9�p4��J( �6�;`"Or�y�Gˍ{�$x����H�N-9�"O���3A�,
��)A&:	��p5"OV�3JR�H`����G�Ľ,�y�JZ�6P���̵L�>��%��yB
]cqj�"s��Z���eH�B�<sZ$4�̍��ʝ�K���P"O��Q�_�Q�p�EW���� �"O֝����?C�j������@H�!"O:\�'��.�����->@k�"O���Y	]@�H0q�!z��8`�"Ol� D��!)hu l[f
@Q"ObIRp��f���hw	��Q����"O�E!&Y%��9R��>�d�@4"Oplsѧ	�. t���g��?Ƣ�ò"O��q��v�21��֊9MD���"O&)0�5 f!⤣�0L�Mj�"O���4�� ��0h���J6����"O4����ΦJa����[=)>��"O���A�ݜh��$�#�ۛ/	H-�S"O�yS�
Bn~<5����sd��d"Ox���
M����t�IM6���"O��Iec[��\���IK>����"O��`R�G�<��L�G��;���a"Of�×�P2-p]��H@{{�m�'"O��0�-ޝtЄ�ѡ��_hƐ
�"O���J�+�r�bN���)J�"O(�ÏS�^|���&�e���q"ONYЁ��h���֎��
J��"Op�K��F=cpL�Tl�h]R� �"OȘb��{5,1�M͍/3���'IN��s�N2lP����M�:��#	�'��h5��9H��y��<W�Pa�'_��9�/�0�t��<��
�'����"Ӗa�,hK��[�C>:�3
�'�(�#D+Y�]���0>� x!
�'��8�"�<i4&��I�i#�@	�']d�P@E�m(����R�L��'�j��QC��w����A�*M��S�'+"��p�-E%��+Q�U�5�:��'g��a7F��g8Erqك:T�%�'`��jw�
#P�&๠��.k�'�0�H��	�*�n��#�VeY�'�JYZ�F�tX�H
����t �'y~l{�'�39;�a��P�V\r��	�'�� ��*~���*THĄl^��'\n$r0kĩ\����X,"H`�'���3����N1M�*x��7D��;Ƌƙ�zIj��Ǩ#M�ݳ#�6D�\04(�8��-�A���<���t�9D�Сg�meX9�Jc��,�ӭ��y ��cb
�#K�<��� P$�y�K����"��EJԙ�r�Ҷ�y�b@�[�v� �I@�B8 �����y�GΫ\���"F�H Ȭs�I��y"iX�b��d�����>���.ʛ�yR"ԝe��	���E�����C��y
� ������d�p�'��1R��x�"Of���+�A3PY A퓭_��7"O,���	E�j�$H�E%�5/.5��"O��d��q���Pd��#E aP"Oj���Ӏ. �4�w�7'��a�"OJ}��BM��p����P�_�q��"O��T-�EY ��<z�<�U"O 3�c� ^|�Agk&KΪL�"O����@+2\IF�@�k��u:�"O�%�w'
:����2
v��l{�"O�-��Y0�S�Jh�`"O����GT"^�P�2Í�3A����b"O��{�g��:�&�y��ʦ����*O�y��JG���b/G'H�Q�'�ܠ6g�F�b��%X1Z���'g^�
K.'�*�`ܘ=���K�'�f�bI|�<���Թk� !�'������s��İ�E�^gB�*
�'����f�d�"0amY����	�'�bպ�KU��B�X2���V�Fl�
�'�jx�  ��